PROV|1|1|Приповісті Соломона, сина Давидового, царя Ізраїлевого,
PROV|1|2|щоб пізнати премудрість і карність, щоб зрозуміти розсудні слова,
PROV|1|3|щоб прийняти напоумлення мудрости, праведности, і права й простоти,
PROV|1|4|щоб мудрости дати простодушним, юнакові пізнання й розважність.
PROV|1|5|Хай послухає мудрий і примножить науку, а розумний здобуде хай мудрих думок,
PROV|1|6|щоб пізнати ту приповість та загадкове говорення, слова мудреців та їхні загадки.
PROV|1|7|Страх Господній початок премудрости, нерозумні погорджують мудрістю та напучуванням.
PROV|1|8|Послухай, мій сину, напучення батька свого, і не відкидай науки матері своєї,
PROV|1|9|вони бо хороший вінок для твоєї голови, і прикраса на шию твою.
PROV|1|10|Мій сину, як грішники будуть тебе намовляти, то з ними не згоджуйся ти!
PROV|1|11|Якщо скажуть вони: Ходи з нами, чатуймо на кров, безпричинно засядьмо на неповинного,
PROV|1|12|живих поковтаймо ми їх, як шеол, та здорових, як тих, які сходять до гробу!
PROV|1|13|Ми знайдемо всіляке багатство цінне, переповнимо здобиччю наші хати.
PROV|1|14|Жеребок свій ти кинеш із нами, буде саква одна для всіх нас,
PROV|1|15|сину мій, не ходи ти дорогою з ними, спини ногу свою від їхньої стежки,
PROV|1|16|бо біжать їхні ноги на зло, і поспішають, щоб кров проливати!
PROV|1|17|Бож надармо поставлена сітка на очах усього крилатого:
PROV|1|18|то вони на кров власну чатують, засідають на душу свою!
PROV|1|19|Такі то дороги усіх, хто заздрий чужого добра: воно бере душу свого власника!
PROV|1|20|Кличе мудрість на вулиці, на площах свій голос дає,
PROV|1|21|на шумливих місцях проповідує, у місті при входах до брам вона каже слова свої:
PROV|1|22|Доки ви, нерозумні, глупоту любитимете? Аж доки насмішники будуть кохатись собі в глузуванні, а безглузді ненавидіти будуть знання?
PROV|1|23|Зверніться но ви до картання мого, ось я виллю вам духа свого, сповіщу вам слова свої!
PROV|1|24|Бо кликала я, та відмовились ви, простягла була руку свою, та ніхто не прислухувався!
PROV|1|25|І всю раду мою ви відкинули, картання ж мого не схотіли!
PROV|1|26|Тож у вашім нещасті сміятися буду і я, насміхатися буду, як прийде ваш страх.
PROV|1|27|Коли прийде ваш страх, немов вихор, і привалиться ваше нещастя, мов буря, як прийде недоля та утиск на вас,
PROV|1|28|тоді кликати будуть мене, але не відповім, будуть шукати мене, та не знайдуть мене,
PROV|1|29|за те, що науку зненавиділи, і не вибрали страху Господнього,
PROV|1|30|не хотіли поради моєї, погорджували всіма моїми докорами!
PROV|1|31|І тому хай їдять вони з плоду дороги своєї, а з порад своїх хай насищаються,
PROV|1|32|бо відступство безумних заб'є їх, і безпечність безтямних їх вигубить!
PROV|1|33|А хто мене слухає, той буде жити безпечно, і буде спокійний від страху перед злом!
PROV|2|1|Сину мій, якщо приймеш слова мої ти, а накази мої при собі заховаєш,
PROV|2|2|щоб слухало мудрости вухо твоє, своє серце прихилиш до розуму,
PROV|2|3|якщо до розсудку ти кликати будеш, до розуму кликатимеш своїм голосом,
PROV|2|4|якщо будеш шукати його, немов срібла, і будеш його ти пошукувати, як тих схованих скарбів,
PROV|2|5|тоді зрозумієш страх Господній, і знайдеш ти Богопізнання,
PROV|2|6|бо Господь дає мудрість, з Його уст знання й розум!
PROV|2|7|Він спасіння ховає для щирих, мов щит той для тих, хто в невинності ходить,
PROV|2|8|щоб справедливих стежок стерегти, і береже Він дорогу Своїх богобійних!
PROV|2|9|Тоді ти збагнеш справедливість та право, і простоту, всіляку дорогу добра,
PROV|2|10|бо мудрість увійде до серця твого, і буде приємне знання для твоєї душі!
PROV|2|11|розважність тоді тебе пильнуватиме, розум тебе стерегтиме,
PROV|2|12|щоб тебе врятувати від злої дороги, від людини, що каже лукаве,
PROV|2|13|від тих, хто стежки простоти покидає, щоб ходити дорогами темряви,
PROV|2|14|що тішаться, роблячи зло, що радіють крутійствами злого,
PROV|2|15|що стежки їхні круті, і відходять своїми путями,
PROV|2|16|щоб тебе врятувати від блудниці, від чужинки, що мовить м'якенькі слова,
PROV|2|17|що покинула друга юнацтва свого, а про заповіт свого Бога забула,
PROV|2|18|вона бо із домом своїм западеться у смерть, а стежки її до померлих,
PROV|2|19|ніхто, хто входить до неї, не вернеться, і стежки життя не досягне,
PROV|2|20|щоб ходив ти дорогою добрих, і стежки справедливих беріг!
PROV|2|21|Бо замешкають праведні землю, і невинні зостануться в ній,
PROV|2|22|а безбожні з землі будуть вигублені, і повириваються з неї невірні!
PROV|3|1|Сину мій, не забудь ти моєї науки, і нехай мої заповіді стережуть твоє серце,
PROV|3|2|бо примножать для тебе вони довготу твоїх днів, і років життя та спокою!
PROV|3|3|Милість та правда нехай не залишать тебе, прив'яжи їх до шиї своєї, напиши їх на таблиці серця свого,
PROV|3|4|і знайдеш ти ласку та добру премудрість в очах Бога й людини!
PROV|3|5|Надійся на Господа всім своїм серцем, а на розум свій не покладайся!
PROV|3|6|Пізнавай ти Його на всіх дорогах своїх, і Він випростує твої стежки.
PROV|3|7|Не будь мудрий у власних очах, бійся Господа та ухиляйся від злого!
PROV|3|8|Це буде ліком для тіла твого, напоєм для костей твоїх.
PROV|3|9|Шануй Господа із маєтку свого, і з початку всіх плодів своїх,
PROV|3|10|і будуть комори твої переповнені ситістю, а чавила твої будуть переливатись вином молодим!
PROV|3|11|Мій сину, карання Господнього не відкидай, і картання Його не вважай тягарем,
PROV|3|12|бо кого Господь любить, картає того, і кохає, немов батько сина!
PROV|3|13|Блаженна людина, що мудрість знайшла, і людина, що розум одержала,
PROV|3|14|бо ліпше надбання її від надбання срібла, і від щирого золота ліпший прибуток її,
PROV|3|15|дорожча за перли вона, і всіляке жадання твоє не зрівняється з нею.
PROV|3|16|Довгість днів у правиці її, багатство та слава в лівиці її.
PROV|3|17|Дороги її то дороги приємности, всі стежки її мир.
PROV|3|18|Вона дерево життя для тих, хто тримається міцно її, і блаженний, хто держить її!
PROV|3|19|Господь мудрістю землю заклав, небо розумом міцно поставив.
PROV|3|20|Знанням Його порозкривались безодні, і кроплять росою ті хмари.
PROV|3|21|Мій сину, нехай від очей твоїх це не відходить, стережи добрий розум і розважність,
PROV|3|22|і вони будуть життям для твоєї душі, і прикрасою шиї твоєї,
PROV|3|23|Тоді підеш безпечно своєю дорогою, а нога твоя не спотикнеться!
PROV|3|24|Якщо покладешся не будеш боятись, а ляжеш, то буде приємний твій сон.
PROV|3|25|Не будеш боятися наглого страху, ні бурі безбожних, як прийде,
PROV|3|26|бо твоєю надією буде Господь, і Він пильнуватиме ногу твою, щоб вона не зловилась у пастку!
PROV|3|27|Не стримуй добра потребуючому, коли в силі твоєї руки це вчинити,
PROV|3|28|не кажи своїм ближнім: Іди, і знову прийди, а взавтра я дам, коли маєш з собою.
PROV|3|29|Не виорюй лихого на свого ближнього, коли він безпечно з тобою сидить.
PROV|3|30|Не сварися з людиною дармо, якщо злого вона не вчинила тобі.
PROV|3|31|Не заздри насильникові, і ні однієї з доріг його не вибирай,
PROV|3|32|бо бридить Господь крутіями, а з праведними в Нього дружба.
PROV|3|33|Прокляття Господнє на домі безбожного, а мешкання праведних Він благословить,
PROV|3|34|з насмішників Він насміхається, а покірливим милість дає.
PROV|3|35|Мудрі славу вспадковують, а нерозумні носитимуть сором.
PROV|4|1|Послухайте, діти, напучення батькового, і прислухайтеся, щоб навчитися розуму,
PROV|4|2|бо даю я вам добру науку: закона мого не кидайте,
PROV|4|3|бо сином у батька свого я був, пещений й єдиний у неньки своєї.
PROV|4|4|І навчав він мене, і мені говорив: Нехай держиться серце твоє моїх слів, стережи мої заповіді та й живи!
PROV|4|5|Здобудь мудрість, здобудь собі розум, не забудь, і не цурайся слів моїх уст,
PROV|4|6|не кидай її й вона буде тебе стерегти! Кохай ти її й вона буде тебе пильнувати!
PROV|4|7|Початок премудрости мудрість здобудь, а за ввесь свій маєток здобудь собі розуму!
PROV|4|8|Тримай її високо і підійме тебе, ушанує тебе, як її ти пригорнеш:
PROV|4|9|вона дасть голові твоїй гарний вінок, пишну корону тобі подарує!
PROV|4|10|Послухай, мій сину, й бери ти слова мої, і помножаться роки твойого життя,
PROV|4|11|дороги премудрости вчу я тебе, стежками прямими проваджу тебе:
PROV|4|12|коли підеш, то крок твій не буде тісний, а коли побіжиш не спіткнешся!
PROV|4|13|Міцно тримайся напучування, не лишай, його стережи, воно бо життя твоє!
PROV|4|14|На стежку безбожних не йди, і не ходи на дорогу лихих,
PROV|4|15|покинь ти її, не йди нею, усунься від неї й мини,
PROV|4|16|бо вони не заснуть, якщо злого не вчинять, відійметься сон їм, як не зроблять кому, щоб спіткнувся!...
PROV|4|17|Бо вони хліб безбожжя їдять, і вино грабежу попивають.
PROV|4|18|А путь праведних ніби те світло ясне, що світить все більше та більш аж до повного дня!
PROV|4|19|Дорога ж безбожних як темність: не знають, об що спотикнуться...
PROV|4|20|Мій сину, прислухуйся до моїх слів, до речей моїх ухо своє нахили!
PROV|4|21|Нехай не відійдуть вони від очей твоїх, бережи їх в середині серця свого!
PROV|4|22|Бо життя вони тим, хто їх знайде, а для тіла усього його лікування.
PROV|4|23|Над усе, що лише стережеться, серце своє стережи, бо з нього походить життя.
PROV|4|24|Відкинь ти від себе лукавство уст, віддали ти від себе крутійство губ.
PROV|4|25|Нехай дивляться очі твої уперед, а повіки твої нехай перед тобою простують.
PROV|4|26|Стежку ніг своїх вирівняй, і стануть міцні всі дороги твої:
PROV|4|27|не вступайся ні вправо, ні вліво, усунь свою ногу від зла!
PROV|5|1|Мій сину, на мудрість мою уважай, нахили своє ухо до мого розуму,
PROV|5|2|щоб розважність ти міг стерегти, а пізнання хай уста твої стережуть!
PROV|5|3|Бо крапають солодощ губи блудниці, а уста її від оливи масніші,
PROV|5|4|та гіркий їй кінець, мов полин, гострий, як меч обосічний,
PROV|5|5|її ноги до смерти спускаються, шеолу тримаються кроки її!
PROV|5|6|Вона путь життя не урівнює, її стежки непевні, і цього не знає вона.
PROV|5|7|Тож тепер, мої діти, мене ви послухайте, не відходьте від слів моїх уст:
PROV|5|8|віддали ти від неї дорогу свою, і не зближайсь до дверей її дому,
PROV|5|9|щоб слави своєї ти іншим не дав, а роки свої для жорстокого,
PROV|5|10|щоб чужі не наситились сили твоєї й маєтку твого в чужім домі!...
PROV|5|11|І будеш стогнати при своєму кінці, як знеможеться тіло твоє й твої сили,
PROV|5|12|і скажеш: Як ненавидів я те напучування, а картання те серце моє відкидало!
PROV|5|13|І не слухав я голосу своїх учителів, і уха свого не схиляв до наставників...
PROV|5|14|Трохи не був я при кожному злому, в середині збору й громади!...
PROV|5|15|Пий воду з криниці своєї, і текуче з свого колодязя:
PROV|5|16|чи ж мають на вулицю вилиті бути джерела твої, а на площі потоки твоєї води?
PROV|5|17|Нехай вони будуть для тебе, для тебе самого, а не для чужих із тобою!
PROV|5|18|Хай твоє джерело буде благословенне, і радій через жінку твоїх юних літ,
PROV|5|19|вона ланя любовна та серна прекрасна, її перса напоять тебе кожночасно, впивайся ж назавжди коханням її!
PROV|5|20|І нащо, мій сину, ти маєш впиватись блудницею, і нащо ти будеш пригортати груди чужинки?
PROV|5|21|Бож перед очима Господніми всі дороги людини, і стежки її всі Він рівняє:
PROV|5|22|власні провини безбожного схоплять його, і повороззям свого гріха буде зв'язаний він,
PROV|5|23|помиратиме він без напучування, і буде блукати в великій глупоті своїй!...
PROV|6|1|Мій сину, якщо поручився ти за свого ближнього, дав руку свою за чужого,
PROV|6|2|ти попався до пастки з-за слів своїх уст, схоплений ти із-за слів своїх уст!
PROV|6|3|Учини тоді це, сину мій, та рятуйсь, бо впав ти до рук свого ближнього: іди, впади в порох, і на ближніх своїх напирай,
PROV|6|4|не дай сну своїм очам, і дрімання повікам своїм,
PROV|6|5|рятуйся, як серна, з руки, і як птах із руки птахолова!
PROV|6|6|Іди до мурашки, лінюху, поглянь на дороги її й помудрій:
PROV|6|7|нема в неї володаря, ані урядника, ані правителя;
PROV|6|8|вона заготовлює літом свій хліб, збирає в жнива свою їжу.
PROV|6|9|Аж доки, лінюху, ти будеш вилежуватись, коли ти зо сну свого встанеш?
PROV|6|10|Ще трохи поспати, подрімати ще трохи, руки трохи зложити, щоб полежати,
PROV|6|11|і прийде, немов волоцюга, твоя незаможність, і злидні твої, як озброєний муж!...
PROV|6|12|Людина нікчемна, чоловік злочинний, він ходить з лукавими устами,
PROV|6|13|він моргає очима своїми, шургає своїми ногами, знаки подає пальцями своїми,
PROV|6|14|в його серці лукавство виорює зло кожночасно, сварки розсіває,
PROV|6|15|тому нагло приходить погибіль його, буде раптом побитий і ліку нема!
PROV|6|16|Оцих шість ненавидить Господь, а ці сім то гидота душі Його:
PROV|6|17|очі пишні, брехливий язик, і руки, що кров неповинну ллють,
PROV|6|18|серце, що плекає злочинні думки, ноги, що сквапно біжать на лихе,
PROV|6|19|свідок брехливий, що брехні роздмухує, і хто розсіває сварки між братів!
PROV|6|20|Стережи, сину мій, заповідь батька свого, і не відкидай науки матері своєї!
PROV|6|21|Прив'яжи їх на серці своєму назавжди, повісь їх на шиї своїй!
PROV|6|22|Вона буде провадити тебе у ході, стерегтиме тебе, коли будеш лежати, а пробудишся мовити буде до тебе!
PROV|6|23|Бо заповідь Божа світильник, а наука то світло, дорога ж життя то навчальні картання,
PROV|6|24|щоб тебе стерегти від злосливої жінки, від облесливого язика чужинки.
PROV|6|25|Не жадай її вроди у серці своїм, і тебе хай не візьме своїми повіками,
PROV|6|26|бо вартість розпусної жінки то боханець хліба, а жінка заміжня вловлює душу цінну...
PROV|6|27|Чи візьме людина огонь на лоно своє, і одіж її не згорить?
PROV|6|28|Чи буде людина ходити по вугіллю розпаленому, і не попаляться ноги її?
PROV|6|29|Так і той, хто вчащає до жінки свого ближнього: не буде некараним кожен, хто доторкнеться до неї!
PROV|6|30|Не погорджують злодієм, якщо він украде, щоб рятувати життя своє, коли він голодує,
PROV|6|31|та як буде він знайдений, всемеро він відшкодує, віддасть все майно свого дому!
PROV|6|32|Хто чинить перелюб, не має той розуму, він знищує душу свою,
PROV|6|33|побої та сором він знайде, а ганьба його не зітреться,
PROV|6|34|бо заздрощі лютість мужчини, і не змилосердиться він у день помсти:
PROV|6|35|він не зверне уваги на жоден твій викуп, і не схоче, коли ти гостинця прибільшиш!
PROV|7|1|Сину мій, бережи ти слова мої, мої ж заповіді заховай при собі,
PROV|7|2|бережи мої заповіді та й живи, а наука моя немов в очах твоїх та зіниця,
PROV|7|3|прив'яжи їх на пальцях своїх, напиши на таблиці тій серця свого!
PROV|7|4|На мудрість скажи: Ти сестра моя! а розум назви: Мій довірений!
PROV|7|5|щоб тебе стерегти від блудниці, від чужинки, що мовить м'якенькі слова.
PROV|7|6|Бо я визирав був в вікно свого дому, через ґрати мого вікна,
PROV|7|7|і приглядавсь до невіж, розглядався між молоддю. І юнак ось, позбавлений розуму,
PROV|7|8|проходив по ринку при розі його, і ступив по дорозі до дому її,
PROV|7|9|коли вітерець повівав був увечорі дня, у темряві ночі та мороку.
PROV|7|10|Аж ось жінка в убранні блудниці назустріч йому, із серцем підступним,
PROV|7|11|галаслива та непогамована, її ноги у домі своїм не бувають:
PROV|7|12|раз на вулиці, раз на майданах, і при кожному розі чатує вона...
PROV|7|13|І вхопила вона його міцно та й поцілувала його, безсоромним зробила обличчя своє та й сказала йому:
PROV|7|14|У мене тепер мирні жертви, виповнила я сьогодні обіти свої!
PROV|7|15|Тому то я вийшла назустріч тобі, пошукати обличчя твого, і знайшла я тебе!
PROV|7|16|Килимами я вистелила своє ложе, тканинами різних кольорів з єгипетського полотна,
PROV|7|17|постелю свою я посипала миррою, алоєм та цинамоном...
PROV|7|18|Ходи ж, аж до ранку впиватися будем коханням, любов'ю натішимось ми!
PROV|7|19|Бо вдома нема чоловіка, пішов у далеку дорогу:
PROV|7|20|вузлик срібла він узяв в свою руку, хіба на день повні поверне до дому свого...
PROV|7|21|Прихилила його велемовством своїм, облесливістю своїх губ його звабила,
PROV|7|22|він раптом за нею пішов, немов віл, до зарізу проваджений, і немов пес, що ведуть його на ланцюгу до ув'язнення,
PROV|7|23|як той птах, поспішає до сітки, і не знає, що це на життя його пастка...
PROV|7|24|А тепер, мої діти, мене ви послухайте, і на слова моїх уст уважайте:
PROV|7|25|Хай не збочує серце твоє на дороги її, не блукай ти стежками її,
PROV|7|26|бо вона багатьох уже трупами кинула, і численні всі, нею забиті!
PROV|7|27|Її дім до шеолу дороги, що провадять до смертних кімнат...
PROV|8|1|Чи ж мудрість не кличе, і не подає свого голосу розум?
PROV|8|2|На верхів'ях холмів, при дорозі та на перехрестях стоїть он вона!
PROV|8|3|При брамах, при вході до міста, де входиться в двері, там голосно кличе вона:
PROV|8|4|До вас, мужі, я кличу, а мій голос до людських синів:
PROV|8|5|Зрозумійте но, неуки, мудрість, зрозумійте ви розум, безглузді!
PROV|8|6|Послухайте, я бо шляхетне кажу, і відкриття моїх губ то простота.
PROV|8|7|Бо правду говорять уста мої, а лукавство гидота для губ моїх.
PROV|8|8|Всі слова моїх уст справедливі, нема в них крутійства й лукавства.
PROV|8|9|Усі вони прості, хто їх розуміє, і щирі для тих, хто знаходить знання.
PROV|8|10|Візьміть ви картання моє, а не срібло, і знання, добірніше від щирого золота:
PROV|8|11|ліпша бо мудрість за перли, і не рівняються їй всі клейноди!
PROV|8|12|Я, мудрість, живу разом з розумом, і знаходжу пізнання розважне.
PROV|8|13|Страх Господній лихе все ненавидіти: я ненавиджу пиху та гордість, і дорогу лиху та лукаві уста!
PROV|8|14|В мене рада й оглядність, я розум, і сила у мене.
PROV|8|15|Мною царюють царі, а законодавці права справедливі встановлюють.
PROV|8|16|Мною правлять владики й вельможні, всі праведні судді.
PROV|8|17|Я кохаю всіх тих, хто кохає мене, хто ж шукає мене мене знайде!
PROV|8|18|Зо мною багатство та слава, тривалий маєток та правда:
PROV|8|19|ліпший плід мій від щирого золота й золота чистого, а прибуток мій ліпший за срібло добірне!
PROV|8|20|Путтю праведною я ходжу, поміж правних стежок,
PROV|8|21|щоб дати багатство в спадщину для тих, хто кохає мене, і я понаповнюю їхні скарбниці!
PROV|8|22|Господь мене мав на початку Своєї дороги, перше чинів Своїх, спервовіку,
PROV|8|23|відвіку була я встановлена, від початку, від правіку землі.
PROV|8|24|Народжена я, як безодень іще не було, коли не було ще джерел, водою обтяжених.
PROV|8|25|Народжена я, поки гори поставлені ще не були, давніше за пагірки,
PROV|8|26|коли ще землі не вчинив Він, ні піль, ні початкового пороху всесвіту.
PROV|8|27|Коли приправляв небеса я була там, коли круга вставляв на поверхні безодні,
PROV|8|28|коли хмари уміцнював Він нагорі, як джерела безодні зміцняв,
PROV|8|29|коли клав Він для моря устава його, щоб його берегів вода не переходила, коли ставив основи землі,
PROV|8|30|то я майстром у Нього була, і була я веселощами день-у-день, радіючи перед обличчям Його кожночасно,
PROV|8|31|радіючи на земнім крузі Його, а забава моя із синами людськими!
PROV|8|32|Тепер же, послухайте, діти, мене, і блаженні, хто буде дороги мої стерегти!
PROV|8|33|Навчання послухайте й мудрими станьте, і не відступайте від нього!
PROV|8|34|Блаженна людина, яка мене слухає, щоб пильнувати при дверях моїх день-у-день, щоб одвірки мої берегти!
PROV|8|35|Хто бо знаходить мене, той знаходить життя, і одержує милість від Господа.
PROV|8|36|А хто проти мене грішить, ограбовує душу свою; всі, хто мене ненавидить, ті смерть покохали!
PROV|9|1|Мудрість свій дім збудувала, сім стовпів своїх витесала.
PROV|9|2|Зарізала те, що було на заріз, змішала вино своє, і трапезу свою приготовила.
PROV|9|3|Дівчат своїх вислала, і кличе вона на висотах міських:
PROV|9|4|Хто бідний на розум, хай прийде сюди, а хто нерозумний, говорить йому:
PROV|9|5|Ходіть, споживайте із хліба мого, та пийте з вина, що його я змішала!
PROV|9|6|Покиньте глупоту і будете жити, і ходіте дорогою розуму!
PROV|9|7|Хто картає насмішника, той собі ганьбу бере, хто ж безбожникові виговорює, сором собі набуває.
PROV|9|8|Не дорікай пересмішникові, щоб тебе не зненавидів він, викартай мудрого й він покохає тебе.
PROV|9|9|Дай мудрому й він помудріє іще, навчи праведного і прибільшить він мудрости!
PROV|9|10|Страх Господній початок премудрости, а пізнання Святого це розум,
PROV|9|11|бо мною помножаться дні твої, і додадуть тобі років життя.
PROV|9|12|Якщо ти змудрів то для себе змудрів, а як станеш насмішником, сам понесеш!
PROV|9|13|Жінка безглузда криклива, нерозумна, і нічого не знає!
PROV|9|14|Сідає вона на сидінні при вході до дому свого, на високостях міста,
PROV|9|15|щоб кликати тих, хто дорогою йде, хто путтю своєю простує:
PROV|9|16|Хто бідний на розум, хай прийде сюди, а хто нерозумний, то каже йому:
PROV|9|17|Вода крадена солодка, і приємний прихований хліб...
PROV|9|18|І не відає він, що самі там мерці, у глибинах шеолу запрошені нею!...
PROV|10|1|Син мудрий потіха для батька, а син нерозумний то смуток для неньки його.
PROV|10|2|Не поможуть неправедні скарби, а справедливість від смерти визволює.
PROV|10|3|Не допустить Господь голодувати душу праведного, а набуток безбожників згине.
PROV|10|4|Ледача рука до убозтва веде, рука ж роботяща збагачує.
PROV|10|5|Хто літом збирає син мудрий, хто ж дрімає в жнива син безпутній.
PROV|10|6|Благословенства на голову праведного, а уста безбожним прикриє насильство.
PROV|10|7|Пам'ять про праведного на благословення, а ймення безбожних загине.
PROV|10|8|Заповіді мудросердий приймає, але дурногубий впаде.
PROV|10|9|Хто в невинності ходить, той ходить безпечно, а хто кривить дороги свої, буде виявлений.
PROV|10|10|Хто оком моргає, той смуток дає, але дурногубий впаде.
PROV|10|11|Уста праведного то джерело життя, а уста безбожним прикриє насильство.
PROV|10|12|Ненависть побуджує сварки, а любов покриває всі вини.
PROV|10|13|В устах розумного мудрість знаходиться, а різка на спину безтямного.
PROV|10|14|Приховують мудрі знання, а уста нерозумного близькі до загибелі.
PROV|10|15|Маєток багатого місто твердинне його, погибіль убогих їхні злидні.
PROV|10|16|Дорібок праведного на життя, прибуток безбожного в гріх.
PROV|10|17|Хто напучування стереже той на стежці життя, а хто нехтує картання, той блудить.
PROV|10|18|Хто ненависть ховає, в того губи брехливі, а хто наклепи ширить, той дурноверхий.
PROV|10|19|Не бракує гріха в многомовності, а хто стримує губи свої, той розумний.
PROV|10|20|Язик праведного то добірне срібло, а розум безбожних мізерний.
PROV|10|21|Пасуть багатьох губи праведного, безглузді ж умирають з нерозуму.
PROV|10|22|Благословення Господнє воно збагачає, і смутку воно не приносить з собою.
PROV|10|23|Нешляхетне робити забава невігласа, а мудрість людині розумній.
PROV|10|24|Чого нечестивий боїться, те прийде на нього, а прагнення праведних сповняться.
PROV|10|25|Як буря, яка пронесеться, то й гине безбожний, а праведний має довічну основу.
PROV|10|26|Як оцет зубам, і як дим для очей, так лінивий для тих, хто його посилає.
PROV|10|27|Страх Господній примножує днів, а роки безбожних вкоротяться.
PROV|10|28|Сподівання для праведних радість, а надія безбожних загине.
PROV|10|29|Дорога Господня твердиня невинним, а загибіль злочинцям.
PROV|10|30|Повік праведний не захитається, а безбожники не поживуть на землі.
PROV|10|31|Уста праведного дають мудрість, а лукавий язик буде втятий.
PROV|10|32|Уста праведного уподобання знають, а уста безбожних лукавство.
PROV|11|1|Обманливі шальки огида для Господа, а повна вага це Його уподоба.
PROV|11|2|Прийде пишність, та прийде і ганьба, а з сумирними мудрість.
PROV|11|3|Невинність простосердих веде їх, а лукавство зрадливих їх вигубить.
PROV|11|4|Не поможе багатство в день гніву, а справедливість від смерти визволює.
PROV|11|5|Справедливість невинного дорогу йому випростовує, безбожний же падає через безбожність свою.
PROV|11|6|Справедливість прямих їх рятує, а зрадливі захоплені будуть своєю захланністю.
PROV|11|7|При смерті людини безбожної гине надія, зникає чекання людини нікчемної.
PROV|11|8|Виривається праведний з утиску, і замість нього безбожний іде.
PROV|11|9|Свого ближнього нищить лукавий устами, а знанням визволяються праведні.
PROV|11|10|Добром праведних місто радіє, а як гинуть безбожні співає.
PROV|11|11|Благословенням чесних підноситься місто, а устами безбожних руйнується.
PROV|11|12|Хто погорджує ближнім своїм, той позбавлений розуму, а розумна людина мовчить.
PROV|11|13|Виявляє обмовник таємне, вірнодухий же справу ховає.
PROV|11|14|Народ падає з браку розумного проводу, при численності ж радників спасіння буває.
PROV|11|15|Зле робить, як хто за чужого поручується, хто ж поруку ненавидить, той безпечний.
PROV|11|16|Жінка чеснотна осягує слави, і пильні багатства здобудуть.
PROV|11|17|Людина ласкава душі своїй чинить добро, а жорстока замучує тіло своє.
PROV|11|18|Чинить діло безвартне безбожний, хто ж праведність сіє заплату правдиву одержує.
PROV|11|19|Отак праведність є на життя, хто ж женеться за злом, той до смерти зближається.
PROV|11|20|Серцем лукаві огида для Господа, а хто в неповинності ходить Його уподоба.
PROV|11|21|Ручаюсь: не буде невинним лихий, а нащадок правдивих захований буде.
PROV|11|22|Золотая сережка в свині на ніздрі це жінка гарна, позбавлена розуму.
PROV|11|23|Жадання у праведних тільки добро, надія безбожних то гнів.
PROV|11|24|Дехто щедро дає, та ще додається йому, а дехто ховає над міру, та тільки бідніє.
PROV|11|25|Душа, яка благословляє, насичена буде, а хто поїть інших, напоєний буде і він.
PROV|11|26|Хто задержує збіжжя, того проклинає народ, хто ж поживу випродує, тому благословення на голову.
PROV|11|27|Хто прагне добра, той шукає вподобання, хто ж лихого жадає, то й прийде на нього воно.
PROV|11|28|Хто надію кладе на багатство своє, той впаде, а праведники зеленіють, як листя.
PROV|11|29|Хто неряд уносить до дому свого, той вітер посяде, а дурноголовий розумному стане рабом.
PROV|11|30|Плід праведного дерево життя, і мудрий життя набуває.
PROV|11|31|Коли праведний ось надолужується на землі, то тим більше безбожний та грішний!
PROV|12|1|Хто любить навчання, той любить пізнання, а хто докір ненавидить, той нерозумний.
PROV|12|2|Добрий від Господа має вподобання, а людину злих замірів осудить Господь.
PROV|12|3|Не зміцниться людина безбожністю, корінь же праведних не захитається.
PROV|12|4|Жінка чеснотна корона для чоловіка свого, а засоромлююча мов та гниль в його костях.
PROV|12|5|Думки праведних право, підступні заміри безбожних омана.
PROV|12|6|Безбожних слова чатування на кров, а уста невинних урятовують їх.
PROV|12|7|Перевернути безбожних і вже їх нема, а дім праведних буде стояти.
PROV|12|8|Хвалять людину за розум її, а кривосердий стає на погорду.
PROV|12|9|Ліпше простий, але роботящий на себе, від того, хто поважним себе видає, та хліба позбавлений.
PROV|12|10|Піклується праведний життям худоби своєї, а серце безбожних жорстоке.
PROV|12|11|Хто оброблює землю свою, той хлібом насичується, хто ж за марницею гониться, той позбавлений розуму.
PROV|12|12|Безбожний жадає ловити у сітку лихих, а в праведних корень приносить плоди.
PROV|12|13|Пастка злого в гріху його уст, а праведний з утиску вийде.
PROV|12|14|Людина насичується добром з плоду уст, і зроблене рук чоловіка до нього впаде.
PROV|12|15|Дорога безумця пряма в його очах, а мудрий послухає ради.
PROV|12|16|Нерозумного гнів пізнається відразу, розумний же мовчки ховає зневагу.
PROV|12|17|Хто правду говорить, той виявлює праведність, а свідок брехливий оману.
PROV|12|18|Дехто говорить, мов коле мечем, язик же премудрих то ліки.
PROV|12|19|Уста правдиві стоятимуть вічно, а брехливий язик лиш на хвилю.
PROV|12|20|В серці тих, хто зло оре, омана, а радість у тих, хто дораджує мир.
PROV|12|21|Жодна кривда не трапиться праведному, а безбожні наповняться лихом.
PROV|12|22|Уста брехливі огида у Господа, а чинячі правду Його уподоба.
PROV|12|23|Приховує мудра людина знання, а серце безумних глупоту викликує.
PROV|12|24|Роботяща рука пануватиме, а лінива даниною стане.
PROV|12|25|Туга на серці людини чавить її, добре ж слово її веселить.
PROV|12|26|Праведний вивідає свою путь, а дорога безбожних зведе їх самих.
PROV|12|27|Не буде ледачий пекти свого полову, а людина трудяща набуде маєток цінний.
PROV|12|28|В путі праведности є життя, і на стежці її нема смерти.
PROV|13|1|Син мудрий приймає картання від батька, а насмішник докору не слухає.
PROV|13|2|З плоду уст чоловік споживає добро, а жадоба зрадливих насильство.
PROV|13|3|Хто уста свої стереже, той душу свою береже, а хто губи свої розпускає, на того погибіль.
PROV|13|4|Пожадає душа лінюха, та даремно, душа ж роботящих насититься.
PROV|13|5|Ненавидить праведний слово брехливе, безбожний же чинить лихе, і себе засоромлює.
PROV|13|6|Праведність оберігає невинного на дорозі його, а безбожність погублює грішника.
PROV|13|7|Дехто вдає багача, хоч нічого не має, а дехто вдає бідака, хоч маєток великий у нього.
PROV|13|8|Викуп за душу людини багатство її, а вбогий й докору не чує.
PROV|13|9|Світло праведних весело світить, а світильник безбожних погасне.
PROV|13|10|Тільки сварка пихою зчиняється, а мудрість із тими, хто радиться.
PROV|13|11|Багатство, заскоро здобуте, поменшується, хто ж збирає помалу примножує.
PROV|13|12|Задовга надія недуга для серця, а бажання, що сповнюється, це дерево життя.
PROV|13|13|Хто погорджує словом Господнім, той шкодить собі, хто ж страх має до заповіді, тому надолужиться.
PROV|13|14|Наука премудрого криниця життя, щоб віддалитися від пасток смерти.
PROV|13|15|Добрий розум приносить приємність, а дорога зрадливих погуба для них.
PROV|13|16|Кожен розумний за мудрістю робить, а безумний глупоту показує.
PROV|13|17|Безбожний посол у нещастя впаде, а вірний посол немов лік.
PROV|13|18|Хто ламає поуку убозтво та ганьба тому, а хто береже осторогу шанований він.
PROV|13|19|Виконане побажання приємне душі, а вступитись від зла то огида безумним.
PROV|13|20|Хто з мудрими ходить, той мудрим стає, а хто товаришує з безумним, той лиха набуде.
PROV|13|21|Грішників зло доганяє, а праведним Бог надолужить добром.
PROV|13|22|Добрий лишає спадок і онукам, маєток же грішника схований буде для праведного.
PROV|13|23|Убогому буде багато поживи і з поля невправного, та деякі гинуть з безправ'я.
PROV|13|24|Хто стримує різку свою, той ненавидить сина свого, хто ж кохає його, той шукає для нього картання.
PROV|13|25|Праведний їсть, скільки схоче душа, живіт же безбожників завсіди брак відчуває.
PROV|14|1|Мудра жінка будує свій дім, а безумна своєю рукою руйнує його.
PROV|14|2|Хто ходить в простоті своїй, боїться той Господа, а в кого дороги криві, той погорджує Ним.
PROV|14|3|На устах безумця галузка пихи, а губи премудрих їх стережуть.
PROV|14|4|Де немає биків, там ясла порожні, а щедрість врожаю у силі вола.
PROV|14|5|Свідок правдивий не лже, а свідок брехливий говорить неправду.
PROV|14|6|Насмішник шукає премудрости, та надаремно, пізнання легке для розумного.
PROV|14|7|Ходи здалека від людини безумної, і від того, в кого мудрих уст ти не бачив.
PROV|14|8|Мудрість розумного то розуміння дороги своєї, а глупота дурних то омана.
PROV|14|9|Нерозумні сміються з гріха, а між праведними уподобання.
PROV|14|10|Серце знає гіркоту своєї душі, і в радість його не втручається інший.
PROV|14|11|Буде вигублений дім безбожних, а намет безневинних розквітне.
PROV|14|12|Буває, дорога людині здається простою, та кінець її стежка до смерти.
PROV|14|13|Також іноді і від сміху болить серце, і закінчення радости смуток.
PROV|14|14|Хто підступного серця, насититься той із доріг своїх, а добра людина із чинів своїх.
PROV|14|15|Вірить безглуздий в кожнісіньке слово, а мудрий зважає на кроки свої.
PROV|14|16|Мудрий боїться й від злого вступає, нерозумний же гнівається та сміливий.
PROV|14|17|Скорий на гнів учиняє глупоту, а людина лукава зненавиджена.
PROV|14|18|Нерозумні глупоту вспадковують, а мудрі знанням коронуються.
PROV|14|19|Поклоняться злі перед добрими, а безбожники при брамах праведного.
PROV|14|20|Убогий зненавиджений навіть ближнім своїм, а в багатого друзі численні.
PROV|14|21|Хто погорджує ближнім своїм, той грішить, а ласкавий до вбогих блаженний.
PROV|14|22|Чи ж не блудять, хто оре лихе? А милість та правда для тих, хто оре добро.
PROV|14|23|Кожна праця приносить достаток, але праця уст в недостаток веде.
PROV|14|24|Корона премудрих їхня мудрість, а вінець нерозумних глупота.
PROV|14|25|Свідок правдивий визволює душі, а свідок обманливий брехні торочить.
PROV|14|26|У Господньому страхові сильна надія, і Він пристановище дітям Своїм.
PROV|14|27|Страх Господній криниця життя, щоб віддалятися від пасток смерти.
PROV|14|28|У численності люду величність царя, а в браку народу погибіль володаря.
PROV|14|29|Терпеливий у гніві багаторозумний, а гнівливий вчиняє глупоту.
PROV|14|30|Лагідне серце життя то для тіла, а заздрість гнилизна костей.
PROV|14|31|Хто тисне нужденного, той ображає свого Творця, а хто милостивий до вбогого, той поважає Його.
PROV|14|32|Безбожний у зло своє падає, а праведний повний надії й при смерті своїй.
PROV|14|33|Мудрість має спочинок у серці розумного, а що в нутрі безумних, те виявиться.
PROV|14|34|Праведність люд підіймає, а беззаконня то сором народів.
PROV|14|35|Ласка царева рабові розумному, гнів же його проти того, хто соромить його.
PROV|15|1|Лагідна відповідь гнів відвертає, а слово вразливе гнів підіймає.
PROV|15|2|Язик мудрих то добре знання, а уста нерозумних глупоту висловлюють.
PROV|15|3|Очі Господні на кожному місці, позирають на злих та на добрих.
PROV|15|4|Язик лагідний то дерево життя, а лукавство його заламання на дусі.
PROV|15|5|Зневажає безумний напучення батькове, а хто береже осторогу, стає розумніший.
PROV|15|6|Дім праведного скарб великий, а в плоді безбожного безлад.
PROV|15|7|Уста мудрих знання розсівають, а серце безглуздих не так.
PROV|15|8|Жертва безбожних огида для Господа, а молитва невинних Його уподоба.
PROV|15|9|Господеві огида дорога безбожного, а того, хто женеться за праведністю, Він кохає.
PROV|15|10|Люта кара на того, хто путь оставляє, а хто осторогу ненавидить, той умирає.
PROV|15|11|Шеол й Аваддон перед Господом, тим більше серця синів людських!
PROV|15|12|Насмішник не любить картання собі, він до мудрих не піде.
PROV|15|13|Радісне серце лице веселить, а при смутку сердечному дух приголомшений.
PROV|15|14|Серце розумне шукає знання, а уста безумних глупоту пасуть.
PROV|15|15|Нужденному всі дні лихі, кому ж добре на серці, у того гостина постійно.
PROV|15|16|Ліпше мале у Господньому страху, ані ж скарб великий, та тривога при тому.
PROV|15|17|Ліпша пожива яринна, і при тому любов, аніж тучний віл, та ненависть при тому.
PROV|15|18|Гнівлива людина роздражнює сварку, терпелива ж у гніві вспокоює заколот.
PROV|15|19|Дорога лінивого то терновиння, а путь щирих дорога гладка.
PROV|15|20|Мудрий син тішить батька свого, а людина безумна погорджує матір'ю своєю.
PROV|15|21|Глупота то радість для нерозумного, а людина розумна дорогою простою ходить.
PROV|15|22|Ламаються задуми з браку поради, при численності ж радників сповняться.
PROV|15|23|Радість людині у відповіді його уст, а слово на часі своєму яке воно добре!
PROV|15|24|Путь життя для премудрого угору, щоб віддалюватись від шеолу внизу.
PROV|15|25|Дім пишних руйнує Господь, але ставить межу для вдови.
PROV|15|26|Думки злого огида для Господа, але чисті для Нього приємні слова.
PROV|15|27|Зажерливий робить нещасним свій дім, хто ж дарунки ненавидить, той буде жити.
PROV|15|28|Серце праведного розмірковує про відповідь, а уста безбожних вибризкують зло.
PROV|15|29|Далекий Господь від безбожних, але справедливих молитву Він чує.
PROV|15|30|Світло очей тішить серце, добра звістка підкріплює кості.
PROV|15|31|Ухо, що навчання життя вислуховує, буде перебувати між мудрими.
PROV|15|32|Хто напучування не приймає, той не дбає про душу свою, а хто слухається остороги, здобуде той розум.
PROV|15|33|Страх Господній навчання премудрости, а перед славою скромність іде.
PROV|16|1|Заміри серця належать людині, та від Господа відповідь язика.
PROV|16|2|Всі дороги людини чисті в очах її, та зважує душі Господь.
PROV|16|3|Поклади свої чини на Господа, і будуть поставлені міцно думки твої.
PROV|16|4|Все Господь учинив ради цілей Своїх, і безбожного на днину зла.
PROV|16|5|Огида для Господа всякий бундючний, ручуся: не буде такий без вини!
PROV|16|6|Провина викуплюється через милість та правду, і страх Господній відводить від злого.
PROV|16|7|Як дороги людини Господь уподобає, то й її ворогів Він замирює з нею.
PROV|16|8|Ліпше мале справедливе, аніж великі прибутки з безправ'я.
PROV|16|9|Розум людини обдумує путь її, але кроки її наставляє Господь.
PROV|16|10|Вирішальне слово в царя на губах, тому в суді уста його не спроневіряться.
PROV|16|11|Вага й шальки правдиві від Господа, все каміння вагове в торбинці то діло Його.
PROV|16|12|Чинити безбожне огида царям, бо трон зміцнюється справедливістю.
PROV|16|13|Уподоба царям губи праведности, і він любить того, хто правдиве говорить.
PROV|16|14|Гнів царя вісник смерти, та мудра людина злагіднить його.
PROV|16|15|У світлі царського обличчя життя, а його уподоба мов хмара дощева весною.
PROV|16|16|Набування премудрости як же це ліпше від золота, набування ж розуму добірніше від срібла!
PROV|16|17|Путь справедливих ухилятись від зла; хто дорогу свою береже, той душу свою охоронює.
PROV|16|18|Перед загибіллю гордість буває, а перед упадком бундючність.
PROV|16|19|Ліпше бути покірливим із лагідними, ніж здобич ділити з бундючними.
PROV|16|20|Хто вважає на слово, той знайде добро, хто ж надію складає на Господа буде блаженний.
PROV|16|21|Мудросердого кличуть розумний, а солодощ уст прибавляє науки.
PROV|16|22|Розум джерело життя власникові його, а картання безумних глупота.
PROV|16|23|Серце мудрого чинить розумними уста його, і на уста його прибавляє навчання.
PROV|16|24|Приємні слова щільниковий то мед, солодкий душі й лік на кості.
PROV|16|25|Буває, дорога людині здається простою, та кінець її стежка до смерти.
PROV|16|26|Людина трудяща працює для себе, бо до того примушує рот її.
PROV|16|27|Нікчемна людина копає лихе, а на устах її як палючий огонь.
PROV|16|28|Лукава людина сварки розсіває, а обмовник розділює друзів.
PROV|16|29|Насильник підмовлює друга свого, і провадить його по недобрій дорозі.
PROV|16|30|Хто прижмурює очі свої, той крутійства видумує, хто губами знаки подає, той виконує зло.
PROV|16|31|Сивизна то пишна корона, знаходять її на дорозі праведности.
PROV|16|32|Ліпший від силача, хто не скорий до гніву, хто ж панує над собою самим, ліпший від завойовника міста.
PROV|16|33|За пазуху жереб вкладається, та ввесь його вирок від Господа.
PROV|17|1|Ліпший черствий кусок зо спокоєм, ніж дім, повний учти м'ясної зо сваркою.
PROV|17|2|Раб розумний панує над сином безпутнім, і серед братів він поділить спадок.
PROV|17|3|Для срібла топильна посудина, а горно для золота, Господь же серця випробовує.
PROV|17|4|Лиходій слухається уст безбожних, слухає неправдомов язика лиходійного.
PROV|17|5|Хто сміється з убогого, той ображає свого Творця, хто радіє з нещастя, не буде такий без вини.
PROV|17|6|Корона для старших онуки, а пишнота дітей їхні батьки.
PROV|17|7|Не пристойна безумному мова поважна, а тим більше шляхетному мова брехлива.
PROV|17|8|Хабар в очах його власника самоцвіт: до всього, до чого повернеться, буде щастити йому.
PROV|17|9|Хто шукає любови провину ховає, хто ж про неї повторює, розгонює друзів.
PROV|17|10|На розумного більше впливає одне остереження, як на глупака сто ударів.
PROV|17|11|Злий шукає лише неслухняности, та вісник жорстокий на нього пошлеться.
PROV|17|12|Ліпше спіткати обездітнену ведмедицю, що кидається на людину, аніж нерозумного в глупоті його.
PROV|17|13|Хто відплачує злом за добро, не відступить лихе з його дому.
PROV|17|14|Почин сварки то прорив води, тому перед вибухом сварки покинь ти її!
PROV|17|15|Хто оправдує несправедливого, і хто засуджує праведного, обидва вони Господеві огидні.
PROV|17|16|Нащо ті гроші в руці нерозумного, щоб мудрість купити, як мозку нема?
PROV|17|17|Правдивий друг любить за всякого часу, в недолі ж він робиться братом.
PROV|17|18|Людина, позбавлена розуму, ручиться, поруку дає за друга свого.
PROV|17|19|Хто сварку кохає, той любить гріх; хто ж підвищує уста свої, той шукає нещастя.
PROV|17|20|Людина лукавого серця не знайде добра, хто ж лукавить своїм язиком, упаде в зло.
PROV|17|21|Хто родить безумного, родить на смуток собі, і не потішиться батько безглуздого.
PROV|17|22|Серце радісне добре лікує, а пригноблений дух сушить кості.
PROV|17|23|Безбожний таємно бере хабара, щоб зігнути путі правосуддя.
PROV|17|24|З обличчям розумного мудрість, а очі глупця аж на кінці землі.
PROV|17|25|Нерозумний син смуток для батька, для своєї ж родительки гіркість.
PROV|17|26|Не добре карати справедливого, бити шляхетних за щирість!
PROV|17|27|Хто слова свої стримує, той знає пізнання, і холоднокровний розумна людина.
PROV|17|28|І глупак, як мовчить, уважається мудрим, а як уста свої закриває розумним.
PROV|18|1|Примхливий шукає сваволі, стає проти всього розумного.
PROV|18|2|Нерозумний не хоче навчатися, а тільки свій ум показати.
PROV|18|3|З приходом безбожного й ганьба приходить, а з легковаженням сором.
PROV|18|4|Слова уст людини глибока вода, джерело премудрости бризкотливий потік.
PROV|18|5|Не добре вважати на обличчя безбожного, щоб праведного повалити на суді.
PROV|18|6|Уста нерозумного тягнуть до сварки, а слова його кличуть бійки.
PROV|18|7|Язик нерозумного загибіль для нього, а уста його то тенета на душу його.
PROV|18|8|Слова обмовника мов ті присмаки, і вони сходять у нутро утроби.
PROV|18|9|Теж недбалий у праці своїй то брат марнотратнику.
PROV|18|10|Господнє Ім'я сильна башта: до неї втече справедливий і буде безпечний.
PROV|18|11|Маєток багатому місто твердинне його, і немов міцний мур ув уяві його.
PROV|18|12|Перед загибіллю серце людини високо несеться, перед славою ж скромність.
PROV|18|13|Хто відповідає на слово, ще поки почув, то глупота та сором йому!
PROV|18|14|Дух дійсного мужа виносить терпіння своє, а духа прибитого хто піднесе?
PROV|18|15|Серце розумне знання набуває, і вухо премудрих шукає знання.
PROV|18|16|Дарунок людини виводить із утиску, і провадить її до великих людей.
PROV|18|17|Перший у сварці своїй уважає себе справедливим, але прийде противник його та й дослідить його.
PROV|18|18|Жереб перериває сварки, та відділює сильних один від одного.
PROV|18|19|Розлючений брат протиставиться більше за місто твердинне, а сварки, немов засуви замку.
PROV|18|20|Із плоду уст людини насичується її шлунок, вона насичується плодом уст своїх.
PROV|18|21|Смерть та життя у владі язика, хто ж кохає його, його плід поїдає.
PROV|18|22|Хто жінку чеснотну знайшов, знайшов той добро, і милість отримав від Господа.
PROV|18|23|Убогий говорить благально, багатий же відповідає зухвало.
PROV|18|24|Є товариші на розбиття, та є й приятель, більше від брата прив'язаний.
PROV|19|1|Ліпший убогий, що ходить в своїй неповинності, ніж лукавий устами та нерозумний.
PROV|19|2|Теж не добра душа без знання, а хто наглить ногами, спіткнеться.
PROV|19|3|Глупота людини дорогу її викривляє, і на Господа гнівається її серце.
PROV|19|4|Маєток примножує друзів численних, а від бідака відпадає й товариш його...
PROV|19|5|Свідок брехливий не буде без кари, а хто брехні говорить, не буде врятований.
PROV|19|6|Багато-хто годять тому, хто гостинці дає, і кожен товариш людині, яка не скупиться на дари.
PROV|19|7|Бідаря ненавидять всі браття його, а тимбільш його приятелі відпадають від нього; а коли за словами поради женеться, нема їх!
PROV|19|8|Хто ума набуває, кохає той душу свою, а хто розум стереже, той знаходить добро.
PROV|19|9|Свідок брехливий не буде без кари, хто ж неправду говорить, загине.
PROV|19|10|Не лицює пишнота безумному, тим більше рабові панувати над зверхником.
PROV|19|11|Розум людини припинює гнів її, а величність її перейти над провиною.
PROV|19|12|Гнів царя немов рик левчука, а ласкавість його як роса на траву.
PROV|19|13|Син безумний погибіль для батька свого, а жінка сварлива як ринва, що з неї вода тече завжди.
PROV|19|14|Хата й маєток спадщина батьків, а жінка розумна від Господа.
PROV|19|15|Лінощі сон накидають, і лінива душа голодує.
PROV|19|16|Хто заповідь охороняє, той душу свою стереже; хто дороги свої легковажить, помре.
PROV|19|17|Хто милостивий до вбогого, той позичає для Господа, і чин його Він надолужить йому.
PROV|19|18|Картай свого сина, коли є надія навчити, та забити його не піднось свою душу.
PROV|19|19|Людина великого гніву хай кару несе, бо якщо ти врятуєш її, то вчиниш ще гірше.
PROV|19|20|Слухай ради й картання приймай, щоб мудрим ти став при своєму кінці.
PROV|19|21|У серці людини багато думок, але виповниться тільки задум Господній.
PROV|19|22|Здобуток людині то милість її, але ліпший бідар за людину брехливу.
PROV|19|23|Страх Господній веде до життя, і хто його має, той ситим ночує, і зло не досягне його.
PROV|19|24|У миску стромляє лінюх свою руку, до уст же своїх не підійме її.
PROV|19|25|Як битимеш нерозважного, то помудріє й немудрий, а будеш розумного остерігати, то він зрозуміє поуку.
PROV|19|26|Хто батька грабує, хто матір жене? Це син, що застиджує та осоромлює,
PROV|19|27|перестань же, мій сину, навчатися від нерозумних, щоб відступитися від слів знання!
PROV|19|28|Свідок нікчемний висміює суд, а уста безбожних вибризкують кривду.
PROV|19|29|На насмішників кари готові постійно, і вдари на спину безумним.
PROV|20|1|Вино то насмішник, напій п'янкий галасун, і кожен, хто блудить у ньому, немудрий.
PROV|20|2|Страх царя як рик лева; хто до гніву доводить його, проти свого життя прогрішає.
PROV|20|3|Слава людині, що гнів покидає, а кожен глупак вибухає.
PROV|20|4|Лінивий не оре із осени, а захоче в жнива і нічого нема.
PROV|20|5|Рада в серці людини глибока вода, і розумна людина її повичерпує.
PROV|20|6|Багато людей себе звуть милосердними, та вірну людину хто знайде?
PROV|20|7|У своїй неповинності праведний ходить, блаженні по ньому сини його!
PROV|20|8|Цар сидить на суддевім престолі, всяке зло розганяє своїми очима.
PROV|20|9|Хто скаже: Очистив я серце своє, очистився я від свого гріха?
PROV|20|10|Вага неоднакова, неоднакова міра, обоє вони то огида для Господа.
PROV|20|11|Навіть юнак буде пізнаний з чинів своїх, чи чин його чистий й чи простий.
PROV|20|12|Ухо, що слухає, й око, що бачить, Господь учинив їх обоє.
PROV|20|13|Не кохайся в спанні, щоб не збідніти; розплющ свої очі та хлібом наситься!
PROV|20|14|Зле, зле! каже той, хто купує, а як піде собі, тоді хвалиться купном.
PROV|20|15|Є золото й перел багато, та розумні уста найцінніший то посуд.
PROV|20|16|Візьми його одіж, бо він поручивсь за чужого, і за чужинку візьми його застав.
PROV|20|17|Хліб з неправди солодкий людині, та піском потім будуть наповнені уста її.
PROV|20|18|Тримаються заміри радою, і війну провадь мудрими радами.
PROV|20|19|Виявляє обмовник таємне, а ти не втручайся до того, легко хто розтулює уста свої.
PROV|20|20|Хто кляне свого батька та матір свою, погасне світильник йому серед темряви!
PROV|20|21|Спадок спочатку заскоро набутий, не буде кінець його поблагословлений!
PROV|20|22|Не кажи: Надолужу я зло! май надію на Господа, і Він допоможе тобі.
PROV|20|23|Вага неоднакова то огида для Господа, а оманливі шальки не добрі.
PROV|20|24|Від Господа кроки людини, а людина як вона зрозуміє дорогу свою?
PROV|20|25|Тенета людині казати святе нерозважно, а згодом свої обітниці досліджувати.
PROV|20|26|Мудрий цар розпорошить безбожних, і зверне на них своє коло для мук.
PROV|20|27|Дух людини світильник Господній, що все нутро обшукує.
PROV|20|28|Милість та правда царя стережуть, і трона свого він підтримує милістю.
PROV|20|29|Окраса юнацтва їхня сила, а пишність старих сивина.
PROV|20|30|Синяки від побоїв то масть лікувальна на злого, та вдари нутру живота.
PROV|21|1|Водні потоки цареве це серце в Господній руці: куди тільки захоче, його Він скеровує.
PROV|21|2|Всяка дорога людини пряма в її очах, та керує серцями Господь.
PROV|21|3|Справедливість та правду чинити для Господа це добірніше за жертву.
PROV|21|4|Муж гордого ока та серця надутого несправедливий, а світильник безбожних це гріх.
PROV|21|5|Думки пильного лиш на достаток ведуть, а всякий квапливий на збиток.
PROV|21|6|Набування майна язиком неправдивим це скороминуща марнота шукаючих смерти.
PROV|21|7|Насильство безбожних прямує на них, бо права чинити не хочуть.
PROV|21|8|Дорога злочинця крута, а чистий прямий його чин.
PROV|21|9|Ліпше жити в куті на даху, ніж з сварливою жінкою в спільному домі.
PROV|21|10|Лихого жадає душа нечестивого, і в очах його ближній його не отримає милости.
PROV|21|11|Як карають глумливця мудріє безумний, а як мудрого вчать, знання набуває.
PROV|21|12|До дому свого приглядається праведний, а безбожний доводить до зла.
PROV|21|13|Хто вухо своє затикає від зойку убогого, то й він буде кликати, та не отримає відповіді.
PROV|21|14|Таємний дарунок погашує гнів, а неявний гостинець лють сильну.
PROV|21|15|Радість праведному правосуддя чинити, а злочинцеві страх.
PROV|21|16|Людина, що зблуджує від путі розуму, у зборі померлих спочине.
PROV|21|17|Хто любить веселощі, той немаючий, хто любить вино та оливу, той не збагатіє.
PROV|21|18|Безбожний то викуп за праведного, а лукавий за щирого.
PROV|21|19|Ліпше сидіти в пустинній країні, ніж з сварливою та сердитою жінкою.
PROV|21|20|Скарб цінний та олива в мешканні премудрого, та нищить безумна людина його.
PROV|21|21|Хто женеться за праведністю та за милістю, той знаходить життя, справедливість та славу.
PROV|21|22|До міста хоробрих увійде премудрий, і твердиню надії його поруйнує.
PROV|21|23|Хто стереже свої уста й свого язика, той душу свою зберігає від лиха.
PROV|21|24|Надутий пихою насмішник ім'я йому, він робить усе із бундючним зухвальством.
PROV|21|25|Пожадання лінивого вб'є його, бо руки його відмовляють робити,
PROV|21|26|він кожного дня пожадливо жадає, а справедливий дає та не жалує.
PROV|21|27|Жертва безбожних огида, а надто тоді, як за діло безчесне приноситься.
PROV|21|28|Свідок брехливий загине, а людина, що слухає Боже, говоритиме завжди.
PROV|21|29|Безбожна людина жорстока обличчям своїм, а невинний зміцняє дорогу свою.
PROV|21|30|Нема мудрости, ані розуму, ані ради насупроти Господа.
PROV|21|31|Приготовлений кінь на день бою, але перемога від Господа!
PROV|22|1|Ліпше добре ім'я за багатство велике, і ліпша милість за срібло та золото.
PROV|22|2|Багатий та вбогий стрічаються, Господь їх обох створив.
PROV|22|3|Мудрий бачить лихе і ховається, а безумні йдуть і караються.
PROV|22|4|Заплата покори і страху Господнього, це багатство, і слава, й життя.
PROV|22|5|Тернина й пастки на дорозі лукавого, а хто стереже свою душу, відійде далеко від них.
PROV|22|6|Привчай юнака до дороги його, і він, як постаріється, не уступиться з неї.
PROV|22|7|Багатий панує над бідними, а боржник раб позичальника.
PROV|22|8|Хто сіє кривду, той жатиме лихо, а бич гніву його покінчиться.
PROV|22|9|Хто доброго ока, той поблагословлений буде, бо дає він убогому з хліба свого.
PROV|22|10|Глумливого вижени, й вийде з ним сварка, і суперечка та ганьба припиняться.
PROV|22|11|Хто чистість серця кохає, той має хороше на устах, і другом йому буде цар.
PROV|22|12|Очі Господа оберігають знання, а лукаві слова Він відкине.
PROV|22|13|Лінивий говорить: На вулиці лев, серед майдану я буду забитий!
PROV|22|14|Уста коханки яма глибока: на кого Господь має гнів, той впадає туди.
PROV|22|15|До юнакового серця глупота прив'язана, та різка картання віддалить від нього її.
PROV|22|16|Хто тисне убогого, щоб собі збагатитись, і хто багачеві дає, той певно збідніє.
PROV|22|17|Нахили своє вухо, і послухай слів мудрих, і серце зверни до мого знання,
PROV|22|18|бо гарне воно, коли будеш ти їх у своєму нутрі стерегти, хай стануть на устах твоїх вони разом!
PROV|22|19|Щоб надія твоя була в Господі, я й сьогодні навчаю тебе.
PROV|22|20|Хіба ж не писав тобі тричі з порадами та із знанням,
PROV|22|21|щоб тобі завідомити правду, правдиві слова, щоб ти істину міг відповісти тому, хто тебе запитає.
PROV|22|22|Не грабуй незаможнього, бо він незаможній, і не тисни убогого в брамі,
PROV|22|23|бо Господь за їхню справу судитиметься, і грабіжникам їхнім ограбує Він душу.
PROV|22|24|Не дружись із чоловіком гнівливим, і не ходи із людиною лютою,
PROV|22|25|щоб доріг її ти не навчився, і тенета не взяв для своєї душі.
PROV|22|26|Не будь серед тих, хто поруку дає, серед тих, хто поручується за борги:
PROV|22|27|коли ти не матимеш чим заплатити, нащо візьмуть з-під тебе постелю твою?
PROV|22|28|Не пересувай вікової границі, яку встановили батьки твої.
PROV|22|29|Ти бачив людину, моторну в занятті своїм? Вона перед царями спокійно стоятиме, та не встоїть вона перед простими.
PROV|23|1|Коли сядеш хліб їсти з володарем, то пильно вважай, що перед тобою,
PROV|23|2|і поклади собі в горло ножа, якщо ти ненажера:
PROV|23|3|не жадай його ласощів, бо вони хліб обманливий!
PROV|23|4|Не мордуйся, щоб мати багатство, відступися від думки своєї про це,
PROV|23|5|свої очі ти звернеш на нього, й нема вже його: бо конче змайструє воно собі крила, і полетить, мов орел той, до неба...
PROV|23|6|Не їж хліба в злоокого, і не пожадай лакоминок його,
PROV|23|7|бо як у душі своїй він обраховує, такий є. Він скаже тобі: Їж та пий! але серце його не з тобою,
PROV|23|8|той кавалок, якого ти з'їв, із себе викинеш, і свої гарні слова надаремно потратиш!
PROV|23|9|Не кажи до ушей нерозумному, бо погордить він мудрістю слів твоїх.
PROV|23|10|Не пересувай вікової границі, і не входь на сирітські поля,
PROV|23|11|бо їхній Визволитель міцний, Він за справу їхню буде судитись з тобою!
PROV|23|12|Своє серце зверни до навчання, а уші свої до розумних речей.
PROV|23|13|Не стримуй напучування юнака, коли різкою виб'єш його, не помре:
PROV|23|14|ти різкою виб'єш його, і душу його від шеолу врятуєш.
PROV|23|15|Мій сину, якщо твоє серце змудріло, то буде радіти також моє серце,
PROV|23|16|і нутро моє буде тішитись, коли уста твої говоритимуть слушне.
PROV|23|17|Нехай серце твоє не завидує грішним, і повсякчас пильнуй тільки страху Господнього,
PROV|23|18|бо існує майбутнє, і надія твоя не загине.
PROV|23|19|Послухай, мій сину, та й помудрій, і нехай твоє серце ступає дорогою рівною.
PROV|23|20|Не будь поміж тими, що жлуктять вино, поміж тими, що м'ясо собі пожирають,
PROV|23|21|бо п'яниця й жерун збідніють, а сонливий одягне лахміття.
PROV|23|22|Слухай батька свого, він тебе породив, і не гордуй, як постаріла мати твоя.
PROV|23|23|Купи собі й не продавай правду, мудрість, і картання та розум.
PROV|23|24|Буде вельми радіти батько праведного, і родитель премудрого втішиться ним.
PROV|23|25|Хай радіє твій батько та мати твоя, хай потішиться та, що тебе породила.
PROV|23|26|Дай мені, сину мій, своє серце, і очі твої хай кохають дороги мої.
PROV|23|27|Бо блудниця то яма глибока, а криниця тісна чужа жінка.
PROV|23|28|І вона, мов грабіжник, чатує, і примножує зрадників поміж людьми.
PROV|23|29|В кого ой, в кого ай, в кого сварки, в кого клопіт, в кого рани даремні, в кого очі червоні?
PROV|23|30|У тих, хто запізнюється над вином, у тих, хто приходить попробувати вина змішаного.
PROV|23|31|Не дивись на вино, як воно рум'яніє, як виблискує в келіху й рівненько ллється,
PROV|23|32|кінець його буде кусати, як гад, і вжалить, немов та гадюка,
PROV|23|33|пантруватимуть очі твої на чужі жінки, і серце твоє говоритиме дурощі...
PROV|23|34|І ти будеш, як той, хто лежить у середині моря, й як той, хто лежить на щогловім верху.
PROV|23|35|І скажеш: Побили мене, та мені не боліло, мене штурхали, я ж не почув, коли я прокинусь, шукатиму далі того ж...
PROV|24|1|Не завидуй злим людям, не бажай бути з ними,
PROV|24|2|бо їхне серце говорить про здирство, а уста їхні мовлять про зло.
PROV|24|3|Дім будується мудрістю, і розумом ставиться міцно.
PROV|24|4|А через пізнання кімнати наповнюються усіляким маєтком цінним та приємним.
PROV|24|5|Мудрий сильніший від сильного, а людина розумна від повносилого.
PROV|24|6|Тому то провадь війну мудрими радами, бо спасіння в численності радників.
PROV|24|7|Для безумного мудрість занадто висока, своїх уст не розкриє при брамі.
PROV|24|8|Хто чинити лихе заміряє, того звуть лукавим.
PROV|24|9|Замір глупоти то гріх, а насмішник огида людині.
PROV|24|10|Якщо ти в день недолі знесилився, то мала твоя сила.
PROV|24|11|Рятуй узятих на смерть, також тих, хто на страчення хилиться, хіба не підтримаєш їх?
PROV|24|12|Якщо скажеш: Цього ми не знали! чи ж Той, хто серця випробовує, знати не буде? Він Сторож твоєї душі, і він знає про це, і поверне людині за чином її.
PROV|24|13|Їж, сину мій, мед, бо він добрий, а мед щільниковий солодкий він на піднебінні твоїм,
PROV|24|14|отак мудрість пізнай для своєї душі: якщо знайдеш її, то ти маєш майбутність, і надія твоя не понищиться!
PROV|24|15|Не чатуй на помешкання праведного, ти безбожнику, не ограблюй мешкання його,
PROV|24|16|бо праведний сім раз впаде та зведеться, а безбожний в погибіль впаде!
PROV|24|17|Не тішся, як ворог твій падає, а коли він спіткнеться, хай серце твоє не радіє,
PROV|24|18|щоб Господь не побачив, і це не було в Його очах лихим, і щоб Він не звернув Свого гніву від нього на тебе!
PROV|24|19|Не пались на злочинців, не заздри безбожним,
PROV|24|20|бо злому не буде майбутности, світильник безбожних погасне.
PROV|24|21|Бійся, сину мій, Господа та царя, не водися з непевними,
PROV|24|22|бо погибіль їхня нагло постане, а біду від обох тих хто знає?
PROV|24|23|І оце ось походить від мудрих: Звертати увагу в суді на обличчя не добре.
PROV|24|24|Хто буде казати безбожному: Праведний ти! того проклинатимуть люди, і гніватись будуть на того народи.
PROV|24|25|А тим, хто картає його, буде миле оце, і прийде на них благословення добра!
PROV|24|26|Мов у губи цілує, хто відповідає правдиве.
PROV|24|27|Приготуй свою працю надворі, й оброби собі поле, а потім збудуєш свій дім.
PROV|24|28|Не будь ложним свідком на свого ближнього, і не підговорюй устами своїми.
PROV|24|29|Не кажи: Як зробив він мені, так зроблю я йому, верну людині за чином її!
PROV|24|30|Я проходив край поля людини лінивої, та край виноградника недоумкуватого,
PROV|24|31|і ось все воно позаростало терням, будяками покрита поверхня його, камінний же мур його був поруйнований...
PROV|24|32|І бачив я те, і увагу звернув, і взяв я поуку собі:
PROV|24|33|Ще трохи поспати, подрімати ще трохи, руки трохи зложити, щоб полежати,
PROV|24|34|і приходить, немов мандрівник, незаможність твоя, і нужда твоя, як озброєний муж!...
PROV|25|1|І оце Соломонові приповісті, що зібрали люди Єзекії, Юдиного царя.
PROV|25|2|Слава Божа щоб справу сховати, а слава царів щоб розвідати справу.
PROV|25|3|Небо високістю, і земля глибиною, і серце царів недослідимі.
PROV|25|4|Як відкинути жужель від срібла, то золотареві виходить посудина,
PROV|25|5|коли віддалити безбожного з-перед обличчя царевого, то справедливістю міцно поставиться трон його.
PROV|25|6|Перед царем не пишайся, а на місці великих не стій,
PROV|25|7|бо ліпше, як скажуть тобі: Ходи вище сюди! аніж тебе знизити перед шляхетним, що бачили очі твої.
PROV|25|8|Не спішися ставати до позову, бо що будеш робити в кінці його, як тебе засоромить твій ближній?
PROV|25|9|Судися за сварку свою з своїм ближнім, але не виявляй таємниці іншого,
PROV|25|10|щоб тебе не образив, хто слухати буде, і щоб не вернулась на тебе обмова твоя.
PROV|25|11|Золоті яблука на срібнім тарелі це слово, проказане часу свого.
PROV|25|12|Золотая сережка й оздоба зо щирого золота це мудрий картач для уважного уха.
PROV|25|13|Немов снігова прохолода в день жнив посол вірний для тих, хто його посилає, і він душу пана свого оживляє.
PROV|25|14|Хмари та вітер, а немає дощу це людина, що чваниться даром, та його не дає.
PROV|25|15|Володар зм'якшується терпеливістю, а м'якенький язик ломить кістку.
PROV|25|16|Якщо мед ти знайшов, то спожий, скільки досить тобі, щоб ним не пересититися та не звернути.
PROV|25|17|Здержуй ногу свою від дому твого товариша, щоб тобою він не переситивсь, і не зненавидів тебе.
PROV|25|18|Молот, і меч, і гостра стріла, людина, що говорить на ближнього свого, як свідок брехливий.
PROV|25|19|Гнилий зуб та кульгава нога це надія на зрадливого радника в день твого утиску.
PROV|25|20|Що здіймати одежу холодного дня, що лити оцет на соду, це співати пісні серцю засмученому.
PROV|25|21|Якщо голодує твій ворог нагодуй його хлібом, а як спрагнений він водою напій ти його,
PROV|25|22|бо цим пригортаєш ти жар на його голову, і Господь надолужить тобі!
PROV|25|23|Вітер північний народжує дощ, а таємний язик сердите обличчя.
PROV|25|24|Ліпше жити в куті на даху, ніж з сварливою жінкою в спільному домі.
PROV|25|25|Добра звістка з далекого краю це холодна водиця на спрагнену душу.
PROV|25|26|Джерело скаламучене чи зіпсутий потік це праведний, що схиляється перед безбожним.
PROV|25|27|Їсти меду багато не добре, так досліджувати власну славу неслава.
PROV|25|28|Людина, що стриму немає для духу свого, це зруйноване місто без муру.
PROV|26|1|Як літом той сніг, і як дощ у жнива, так не лицює глупцеві пошана.
PROV|26|2|Як пташка літає, як ластівка лине, так невинне прокляття не сповниться.
PROV|26|3|Батіг на коня, оброть на осла, а різка на спину глупців.
PROV|26|4|Нерозумному відповіді не давай за нерозум його, щоб і ти не став рівний йому.
PROV|26|5|Нерозумному відповідь дай за безумством його, щоб він в очах своїх не став мудрим.
PROV|26|6|Хто через глупця посилає слова, той ноги собі обтинає, отруту він п'є.
PROV|26|7|Як волочаться ноги в кульгавого, так у безумних устах приповістка.
PROV|26|8|Як прив'язувати камінь коштовний до пращі, так глупцеві пошану давати.
PROV|26|9|Як терен, що влізе у руку, отак приповістка в устах нерозумного.
PROV|26|10|Як стрілець, що все ранить, так і той, хто наймає глупця, і наймає усяких прохожих.
PROV|26|11|Як вертається пес до своєї блювотини, так глупоту свою повторяє глупак.
PROV|26|12|Чи ти бачив людину, що мудра в очах своїх? Більша надія глупцеві, ніж їй.
PROV|26|13|Лінивий говорить: Лев на дорозі! Лев на майдані!
PROV|26|14|Двері обертаються на своєму чопі, а лінивий на ліжку своїм.
PROV|26|15|Свою руку лінивий стромляє до миски, та піднести до рота її йому тяжко.
PROV|26|16|Лінивий мудріший ув очах своїх за сімох, що відповідають розумно.
PROV|26|17|Пса за вуха хапає, хто, йдучи, устряває до сварки чужої.
PROV|26|18|Як той, хто вдає божевільного, кидає іскри, стріли та смерть,
PROV|26|19|так і людина, що обманює друга свого та каже: Таж це я жартую!...
PROV|26|20|З браку дров огонь гасне, а без пліткаря мовкне сварка.
PROV|26|21|Вугілля для жару, а дрова огневі, а людина сварлива щоб сварку розпалювати.
PROV|26|22|Слова обмовника мов ті присмаки, й у нутро живота вони сходять.
PROV|26|23|Як срібло з жужелицею, на горшкові накладене, так полум'яні уста, а серце лихе,
PROV|26|24|устами своїми маскується ворог, і ховає оману в своєму нутрі:
PROV|26|25|коли він говорить лагідно не вір ти йому, бо в серці його сім огид!
PROV|26|26|Як ненависть прикрита оманою, її зло відкривається в зборі.
PROV|26|27|Хто яму копає, той в неї впаде, а хто котить каміння на нього воно повертається.
PROV|26|28|Брехливий язик ненавидить своїх утискуваних, і уста гладенькі до згуби провадять.
PROV|27|1|Не вихвалюйся завтрішнім днем, бо не знаєш, що день той породить.
PROV|27|2|Нехай інший тебе вихваляє, а не уста твої, чужий, а не губи твої.
PROV|27|3|Каміння тягар, і пісок важка річ, та гнів нерозумного тяжчий від них від обох.
PROV|27|4|Лютість жорстокість, а гнів то затоплення, та хто перед заздрістю встоїть?
PROV|27|5|Ліпше відкрите картання, ніж таємна любов.
PROV|27|6|Побої коханого вірність показують, а в ненависника поцілунки численні.
PROV|27|7|Сита душа топче й мед щільниковий, а голодній душі все гірке то солодке.
PROV|27|8|Як птах, що гніздо своє кинув, так і людина, що з місця свого мандрує.
PROV|27|9|Олива й кадило потішують серце, і солодкий нам друг за душевну пораду.
PROV|27|10|Друга свого й друга батька свого не кидай, а в дім брата свого не приходь в день нещастя свого, ліпший сусіда близький за далекого брата!
PROV|27|11|Будь мудрий, мій сину, й потіш моє серце, і я матиму що відповісти, як мені докорятиме хто.
PROV|27|12|Мудрий бачить лихе і ховається, а безумні йдуть і караються.
PROV|27|13|Візьми його одіж, бо він поручивсь за чужого, і за чужинку заставу візьми.
PROV|27|14|Хто сильним голосом благословляє із раннього ранку свого товариша, за прокляття залічується це йому.
PROV|27|15|Ринва, постійно текуча слотливого дня та жінка сварлива однакове:
PROV|27|16|хто хоче сховати її той вітра ховає, чи оливу пахучу правиці своєї, що видасть себе.
PROV|27|17|Як гострить залізо залізо, так гострить людина лице свого друга.
PROV|27|18|Сторож фіґовниці плоди її споживає, а хто пана свого стереже, той шанований.
PROV|27|19|Як лице до лиця у воді, так серце людини до серця людини.
PROV|27|20|Шеол й Аваддон не наситяться, не наситяться й очі людини.
PROV|27|21|Що для срібла топильна посудина, і горно для золота, те для людини уста, які хвалять її.
PROV|27|22|Хоч нерозумного будеш товкти товкачем поміж зернами в ступі, не відійде від нього глупота його!
PROV|27|23|Добре знай вигляд своєї отари, поклади своє серце на череди,
PROV|27|24|бо багатство твоє не навіки, і чи корона твоя з роду в рід?
PROV|27|25|Появилася зелень, і трава показалась, і збирається сіно із гір,
PROV|27|26|будуть вівці тобі на вбрання, і козли ціна поля,
PROV|27|27|і молока твоїх кіз буде досить на їжу тобі, на їду твого дому, і на життя для служниць твоїх.
PROV|28|1|Безбожні втікають, коли й не женуться за ними, а справедливий безпечний, немов той левчук.
PROV|28|2|Коли край провиниться, то має багато володарів, коли ж є людина розумна й знаюча, то держиться довго.
PROV|28|3|Людина убога, що гнобить нужденних, це злива рвучка, що хліба по ній не буває.
PROV|28|4|Ті, хто Закон залишає, хвалять безбожних, а ті, хто Закон береже, на них буряться.
PROV|28|5|Люди лихі правосуддя не розуміють, а шукаючі Господа все розуміють.
PROV|28|6|Ліпше убогий, що ходить в своїй неповинності, ніж криводорогий, хоч він і багач.
PROV|28|7|Хто Закон береже, розумний той син, а хто водиться із гультяями, засоромлює батька свого.
PROV|28|8|Хто множить лихварським відсотком багатство своє, той для того громадить його, хто ласкавий для бідних.
PROV|28|9|Хто відхилює вухо своє, щоб не слухати Закона, то буде огидна й молитва того.
PROV|28|10|Хто простих доводить блудити дорогою зла, сам до ями своєї впаде, а невинні посядуть добро.
PROV|28|11|Багата людина в очах своїх мудра, та розумний убогий розслідить її.
PROV|28|12|Велика пишнота, як тішаться праведні, коли ж несправедливі зростають, то треба шукати людину.
PROV|28|13|Хто ховає провини свої, тому не ведеться, а хто признається та кидає їх, той буде помилуваний.
PROV|28|14|Блаженна людина, що завжди обачна, а хто ожорсточує серце своє, той впадає в лихе.
PROV|28|15|Лев ричучий й ведмідь ненажерливий це безбожний володар над людом убогим.
PROV|28|16|Володар, позбавлений розуму, тисне дошкульно, а ненависник зажерливости буде мати дні довгі.
PROV|28|17|Людина, обтяжена за душогубство, втікає до гробу, нехай її не підпирають!
PROV|28|18|Хто ходить невинний, той буде спасений, а криводорогий впаде на одній із доріг.
PROV|28|19|Хто землю свою обробляє, той насититься хлібом, а хто за марнотним женеться, насититься вбогістю.
PROV|28|20|Вірна людина багата на благословення, а хто спішно збагачується, непокараним той не залишиться.
PROV|28|21|Увагу звертати на особу не добре, бо й за кус хліба людина згрішить.
PROV|28|22|Завидюща людина спішить до багатства, і не знає, що прийде на неї нужда.
PROV|28|23|Хто напоумляє людину, той знаходить вкінці більшу ласку, ніж той, хто лестить язиком.
PROV|28|24|Хто батька свого й свою матір грабує і каже: Це не гріх, той розбійнику друг.
PROV|28|25|Захланний викликує сварку, хто ж має надію на Господа, буде насичений.
PROV|28|26|Хто надію кладе на свій розум, то він нерозумний, а хто мудрістю ходить, той буде врятований.
PROV|28|27|Хто дає немаючому, той недостатку не знатиме, хто ж свої очі ховає від нього, той зазнає багато проклять.
PROV|28|28|Коли підіймаються люди безбожні, людина ховається, а як гинуть вони, то множаться праведні.
PROV|29|1|Чоловік остережуваний, та твердошиїй, буде зламаний нагло, і ліку не буде йому.
PROV|29|2|Коли множаться праведні, радіє народ, як панує ж безбожний то стогне народ.
PROV|29|3|Людина, що мудрість кохає, потішує батька свого, а хто попасає блудниць, той губить маєток.
PROV|29|4|Цар утримує край правосуддям, а людина хабарна руйнує його.
PROV|29|5|Людина, що другові своєму підлещує, на стопах його пастку ставить.
PROV|29|6|У провині людини лихої знаходиться пастка, а справедливий радіє та тішиться.
PROV|29|7|Праведний знає про право вбогих, безбожний же не розуміє пізнання про це.
PROV|29|8|Люди глузливі підбурюють місто, а мудрі утишують гнів.
PROV|29|9|Мудра людина, що правується із нерозумним, то чи гнівається, чи сміється, спокою не знає.
PROV|29|10|Кровожерці ненавидять праведного, справедливі ж шукають спасти його душу.
PROV|29|11|Глупак увесь свій гнів увиявляє, а мудрий назад його стримує.
PROV|29|12|Володар, що слухає слова брехливого, безбожні всі слуги його!
PROV|29|13|Убогий й гнобитель стрічаються, їм обом Господь очі освітлює.
PROV|29|14|Як цар правдою судить убогих, стоятиме трон його завжди.
PROV|29|15|Різка й поука премудрість дають, а дитина, залишена тільки собі, засоромлює матір свою.
PROV|29|16|Як множаться несправедливі провина розмножується, але праведні бачитимуть їхній упадок.
PROV|29|17|Карай сина свого й він тебе заспокоїть, і приємнощі дасть для твоєї душі.
PROV|29|18|Без пророчих видінь люд розбещений, коли ж стереже він Закона блаженний.
PROV|29|19|Раб словами не буде покараний, хоч він розуміє, але не послухає.
PROV|29|20|Чи бачив людину, квапливу в словах своїх? Більша надія глупцеві, ніж їй!
PROV|29|21|Хто розпещує змалку свого раба, то кінець його буде невдячний.
PROV|29|22|Гнівлива людина викликує сварку, а лютий вчиняє багато провин.
PROV|29|23|Гординя людини її понижає, а чести набуває покірливий духом.
PROV|29|24|Хто ділиться з злодієм, той ненавидить душу свою, він чує прокляття, та не виявляє.
PROV|29|25|Страх перед людиною пастку дає, хто ж надію складає на Господа, буде безпечний.
PROV|29|26|Багато шукають для себе обличчя володаря, та від Господа суд для людини.
PROV|29|27|Насильник огида для праведних, а простодорогий огида безбожному.
PROV|30|1|Слова Агура, Якеєвого сина, массеянина: Слово мужчини: Трудився я, Боже, трудився я, Боже, і змучився я!
PROV|30|2|Бо думаю, що немудріший за кожного я, і не маю я людського розуму,
PROV|30|3|і не навчився я мудрости, і не знаю пізнання святих...
PROV|30|4|Хто на небо ввійшов і зійшов? Хто у жмені свої зібрав вітер? Хто воду в одежу зв'язав? Хто поставив усі кінці землі? Яке ймення його, і яке ймення сина його, коли знаєш?
PROV|30|5|Кожне Боже слово очищене, щит Він для тих, хто в Нім пристановище має.
PROV|30|6|До слів Його не додавай, щоб тебе не скартав Він, і щоб неправдомовцем не став ти.
PROV|30|7|Двох речей я від Тебе просив, не відмов мені, поки помру:
PROV|30|8|віддали Ти від мене марноту та слово брехливе, убозтва й багатства мені не давай! Годуй мене хлібом, для мене призначеним,
PROV|30|9|щоб я не переситився та й не відрікся, і не сказав: Хто Господь? і щоб я не збіднів і не крав, і не зневажив Ім'я мого Бога.
PROV|30|10|Раба не обмовляй перед паном його, щоб тебе не прокляв він, і ти винуватим не став.
PROV|30|11|Оце покоління, що батька свого проклинає, і неньки своєї не благословляє,
PROV|30|12|покоління, що чисте в очах своїх, та від бруду свого не обмите,
PROV|30|13|покоління, які гордісні очі його, а повіки його як піднеслися!
PROV|30|14|Покоління, що в нього мечі його зуби, а гострі ножі його щелепи, щоб пожерти убогих із краю й нужденних з землі!
PROV|30|15|Дві дочки в кровожерця: Дай, дай! Оці три не наситяться, чотири не скажуть досить:
PROV|30|16|шеол та утроба неплідна, водою земля не насититься, і не скаже досить огонь!
PROV|30|17|Око, що з батька сміється й погорджує послухом матері, нехай видзьобають його круки поточні, і нехай орленята його пожеруть!
PROV|30|18|Три речі оці дивовижні для мене, і чотири, яких я не знаю:
PROV|30|19|дорога орлина в повітрі, дорога зміїна на скелі, корабельна дорога в середині моря, і дорога мужчини при дівчині!...
PROV|30|20|Така ось дорога блудливої жінки: наїлась та витерла уста свої й повіла: Не вчинила я злого!...
PROV|30|21|Трясеться земля під трьома, і під чотирма, яких знести не може вона:
PROV|30|22|під рабом, коли він зацарює, і під нерозумним, як хліба наїсться,
PROV|30|23|під розпустницею, коли взята за жінку, і невільницею, коли вижене пані свою!...
PROV|30|24|Оці ось чотири малі на землі, та вони вельми мудрі:
PROV|30|25|мурашки, не сильний народ, та поживу свою заготовлюють літом;
PROV|30|26|борсуки, люд не сильний, та в скелі свій дім вони ставлять;
PROV|30|27|немає царя в сарани, але вся вона в строї бойовім виходить;
PROV|30|28|павук тільки лапками пнеться, та він і в палатах царських!
PROV|30|29|Добре ступають ці троє, і добре ходять чотири:
PROV|30|30|лев, найсильніший поміж звіриною, який не вступається ні перед ким,
PROV|30|31|осідланий кінь, і козел, та той цар, що з ним військо!
PROV|30|32|Якщо ти допустився глупоти пихою, й якщо заміряєш лихе, то руку на уста!
PROV|30|33|Бо збивання молока дає масло, і дає кров вдар по носі, тиск же на гнів дає сварку.
PROV|31|1|Слова Лемуїла, царя Масси, що ними навчала його його мати:
PROV|31|2|Що, сину мій, і що, сину утроби моєї, і що, сину обітниць моїх?
PROV|31|3|Не давай жінкам сили своєї, ні доріг своїх для руйнувальниць царів!
PROV|31|4|Не царям, Лемуїле, вино, не царям, і напій той п'янкий не князям,
PROV|31|5|щоб не впився він та не забув про Закона, і щоб не змінив для всіх гноблених права!
PROV|31|6|Дайте напою п'янкого тому, хто гине, а вина гіркодухим:
PROV|31|7|він вип'є й забуде за бідність свою, і муки своєї вже не пам'ятатиме!
PROV|31|8|Відкривай свої уста немові, для суда всім нещасним.
PROV|31|9|Відкривай свої уста, й суди справедливо, і правосуддя зроби для убогого та для нужденного.
PROV|31|10|Хто жінку чеснотну знайде? а ціна її більша від перел:
PROV|31|11|довіряє їй серце її чоловіка, і йому не забракне прибутку!
PROV|31|12|Вона чинить для нього добро, а не зло, по всі дні свого життя.
PROV|31|13|Шукає вона вовни й льону, і робить охоче своїми руками.
PROV|31|14|Вона, немов кораблі ті купецькі, здалека спроваджує хліб свій.
PROV|31|15|І встане вона ще вночі, і видасть для дому свого поживу, а порядок служницям своїм.
PROV|31|16|Про поле вона намишляла, і його набула, із плоду долоней своїх засадила вона виноградника.
PROV|31|17|Вона підперізує силою стегна свої та зміцняє рамена свої.
PROV|31|18|Вона розуміє, що добра робота її, і світильник її не погасне вночі.
PROV|31|19|Вона руки свої простягає до прядки, а долоні її веретено тримають.
PROV|31|20|Долоню свою відкриває для вбогого, а руки свої простягає до бідного.
PROV|31|21|Холоду в домі своїм не боїться вона, бо подвійно одягнений ввесь її дім.
PROV|31|22|Килими поробила собі, віссон та кармазин убрання її.
PROV|31|23|Чоловік її знаний при брамах, як сидить він із старшими краю.
PROV|31|24|Тонку туніку робить вона й продає, і купцеві дає пояси.
PROV|31|25|Сила та пишність одежа її, і сміється вона до прийдещнього дня.
PROV|31|26|Свої уста вона відкриває на мудрість, і милостива наука їй на язиці.
PROV|31|27|Доглядає вона ходи дому свого, і хліба з лінивства не їсть.
PROV|31|28|Устають її діти, і хвалять її, чоловік її й він похваляє її:
PROV|31|29|Багато було тих чеснотних дочок, та ти їх усіх перевищила!
PROV|31|30|Краса то омана, а врода марнота, жінка ж богобоязна вона буде хвалена!
PROV|31|31|Дайте їй з плоду рук її, і нехай її вчинки її вихваляють при брамах!
