PHIL|1|1|Павло й Тимофій, раби Христа Ісуса, до всіх святих у Христі Ісусі, що знаходяться в Филипах, з єпископами та дияконами:
PHIL|1|2|благодать вам і мир від Бога, Отця нашого, і Господа Ісуса Христа!
PHIL|1|3|Дякую Богові своєму при кожній згадці про вас,
PHIL|1|4|і завжди в усякій молитві своїй за всіх вас чиню я молитву з радощами,
PHIL|1|5|за участь вашу в Євангелії від першого дня аж дотепер.
PHIL|1|6|Я певний того, що той, хто в вас розпочав добре діло, виконає його аж до дня Христа Ісуса.
PHIL|1|7|Бо то справедливо мені думати це про всіх вас, бо я маю вас у серці, а ви всі в кайданах моїх, і в обороні, і в утвердженні Євангелії спільники мої в благодаті.
PHIL|1|8|Бо Бог мені свідок, що тужу я за вами всіма в сердечній любові Христа Ісуса.
PHIL|1|9|І молюсь я про те, щоб ваша любов примножалась ще більше та більше в пізнанні й усякім дослідженні,
PHIL|1|10|щоб ви досліджували те, що краще, щоб чисті та цілі були Христового дня,
PHIL|1|11|наповнені плодів праведности через Ісуса Христа, на славу та на хвалу Божу.
PHIL|1|12|Бажаю ж я, браття, щоб відали ви, що те, що сталось мені, вийшло більше на успіх Євангелії,
PHIL|1|13|бо в усій преторії та всім іншим стали відомі кайдани мої за Христа.
PHIL|1|14|А багато братів у Господі через кайдани мої посміліли та ще більше відважилися Слово Боже звіщати безстрашно.
PHIL|1|15|Одні, правда, і через заздрощі та колотнечу, другі ж із доброї волі Христа проповідують;
PHIL|1|16|а інші з любови, знаючи, що я поставлений на оборону Євангелії;
PHIL|1|17|а інші через підступ звіщають Христа нещиро, думаючи, що додадуть тягару до кайданів моїх.
PHIL|1|18|Але що ж? У всякому разі, чи облудно, чи щиро, Христос проповідується, а тим я радію та й буду радіти.
PHIL|1|19|Бо знаю, що це буде мені на спасіння через вашу молитву й допомогу Духа Ісуса Христа,
PHIL|1|20|через чекання й надію мою, що я ні в чому не буду посоромлений, але цілою сміливістю, як завжди, так і тепер Христос буде звеличений у тілі моїм, чи то життям, чи то смертю.
PHIL|1|21|Бо для мене життя то Христос, а смерть то надбання.
PHIL|1|22|А коли життя в тілі то для мене плід діла, то не знаю, що вибрати.
PHIL|1|23|Тягнуть мене одне й друге, хоч я маю бажання померти та бути з Христом, бо це значно ліпше.
PHIL|1|24|А щоб полишатися в тілі, то це потрібніш ради вас.
PHIL|1|25|І оце знаю певно, що залишусь я, і пробуватиму з вами всіма вам на користь та на радощі в вірі,
PHIL|1|26|щоб ваша хвала через мене примножилася в Христі Ісусі, коли знову прийду я до вас.
PHIL|1|27|Тільки живіть згідно з Христовою Євангелією, щоб, чи прийду я й побачу вас, чи й не бувши почув я про вас, що ви стоїте в однім дусі, борючись однодушно за віру євангельську,
PHIL|1|28|і ні в чому не боячися противників; це їм доказ загибелі, вам же спасіння. А це від Бога!
PHIL|1|29|Бо вчинено вам за Христа добродійство, не тільки вірувати в Нього, але і страждати за Нього,
PHIL|1|30|маючи таку саму боротьбу, яку ви бачили в мені, а тепер чуєте про мене.
PHIL|2|1|Отож, коли є в Христі яка заохота, коли є яка потіха любови, коли є яка спільнота духа, коли є яке серце та милосердя,
PHIL|2|2|то доповніть радість мою: щоб думали ви одне й те, щоб мали ту саму любов, одну згоду й один розум!
PHIL|2|3|Не робіть нічого підступом або з чванливости, але в покорі майте один одного за більшого від себе.
PHIL|2|4|Нехай кожен дбає не про своє, але кожен і про інших.
PHIL|2|5|Нехай у вас будуть ті самі думки, що й у Христі Ісусі!
PHIL|2|6|Він, бувши в Божій подобі, не вважав за захват бути Богові рівним,
PHIL|2|7|але Він умалив Самого Себе, прийнявши вигляд раба, ставши подібним до людини; і подобою ставши, як людина,
PHIL|2|8|Він упокорив Себе, бувши слухняний аж до смерти, і то смерти хресної...
PHIL|2|9|Тому й Бог повищив Його, та дав Йому Ім'я, що вище над кожне ім'я,
PHIL|2|10|щоб перед Ісусовим Ім'ям вклонялося кожне коліно небесних, і земних, і підземних,
PHIL|2|11|і щоб кожен язик визнавав: Ісус Христос то Господь, на славу Бога Отця!
PHIL|2|12|Отож, мої любі, як ви завжди слухняні були не тільки в моїй присутності, але значно більше тепер, у моїй відсутності, зо страхом і тремтінням виконуйте своє спасіння.
PHIL|2|13|Бо то Бог викликає в вас і хотіння, і чин за доброю волею Своєю.
PHIL|2|14|Робіть усе без нарікання та сумніву,
PHIL|2|15|щоб були ви бездоганні та щирі, невинні діти Божі серед лукавого та розпусного роду, що в ньому ви сяєте, як світла в світі,
PHIL|2|16|додержуючи слово життя на похвалу мені в день Христа, що я біг не надармо, що я працював не надармо.
PHIL|2|17|Та хоч і стаю я жертвою при жертві і при службі вашої віри, я радію та тішуся разом із вами всіма.
PHIL|2|18|Тіштесь тим самим і ви, і тіштеся разом зо мною!
PHIL|2|19|Надіюся в Господі Ісусі незабаром послати до вас Тимофія, щоб і я зміцнів духом, розізнавши про вас.
PHIL|2|20|Бо я однодумця не маю ні одного, щоб щиріше подбав він про вас.
PHIL|2|21|Усі бо шукають свого, а не Христового Ісусового.
PHIL|2|22|Та ви знаєте досвід його, бо він, немов батькові син, зо мною служив для Євангелії.
PHIL|2|23|Отже, маю надію негайно послати цього, як тільки довідаюся, що буде зо мною.
PHIL|2|24|Але в Господі маю надію, що й сам незабаром прибуду до вас.
PHIL|2|25|Але я вважав за потрібне послати до вас брата Епафродита, свого співробітника та співбойовника, вашого апостола й служителя в потребі моїй,
PHIL|2|26|бо він побивався за вами всіма, і сумував через те, що ви чули, що він хворував.
PHIL|2|27|Бо смертельно він був хворував. Але змилувався Бог над ним, і не тільки над ним, але й надо мною, щоб я смутку на смуток не мав.
PHIL|2|28|Отож, тим швидше послав я його, щоб тішились ви, його знову побачивши, і щоб без смутку я був.
PHIL|2|29|Тож прийміть його в Господі з повною радістю, і майте в пошані таких,
PHIL|2|30|бо за діло Христове наблизився був аж до смерти, наражаючи на небезпеку життя, щоб доповнити ваш нестаток служіння для мене.
PHIL|3|1|Зрештою, браття мої, радійте у Господі! Писати вам те саме не прикро мені, а для вас це навчальне.
PHIL|3|2|Стережіться собак, стережіться працівників лихих, стережіться обрізання!
PHIL|3|3|Бо обрізання то ми, що служимо Богові духом, а хвалимося Христом Ісусом, і не кладемо надії на тіло,
PHIL|3|4|хоч і я міг би мати надію на тіло. Як хто інший на тіло надіятись думає, то тим більше я,
PHIL|3|5|обрізаний восьмого дня, з роду Ізраїля, з племени Веніяминового, єврей із євреїв, фарисей за Законом.
PHIL|3|6|Через горливість я був переслідував Церкву, бувши невинний, щодо правди в Законі.
PHIL|3|7|Але те, що для мене було за надбання, те ради Христа я за втрату вважав.
PHIL|3|8|Тож усе я вважаю за втрату ради переважного познання Христа Ісуса, мого Господа, що я ради Нього відмовився всього, і вважаю все за сміття, щоб придбати Христа,
PHIL|3|9|щоб знайтися в Нім не з власною праведністю, яка від Закону, але з тією, що з віри в Христа, праведністю від Бога за вірою,
PHIL|3|10|щоб пізнати Його й силу Його воскресення, та участь у муках Його, уподоблюючись Його смерті,
PHIL|3|11|аби досягнути якось воскресення з мертвих.
PHIL|3|12|Не тому, що я вже досягнув, або вже вдосконалився, але прагну, чи не досягну я того, чим і Христос Ісус досягнув був мене.
PHIL|3|13|Браття, я себе не вважаю, що я досягнув. Та тільки, забуваючи те, що позаду, і спішачи до того, що попереду,
PHIL|3|14|я женусь до мети за нагородою високого поклику Божого в Христі Ісусі.
PHIL|3|15|Тож усі, хто досконалий, думаймо це; коли ж думаєте ви щось інше, то Бог вам відкриє й це.
PHIL|3|16|Та до чого дійшли ми, поступаймо в тім самім далі.
PHIL|3|17|Будьте до мене подібні, браття, і дивіться на тих, хто поводиться так, як маєте ви за взір нас.
PHIL|3|18|Багато бо хто, що про них я вам часто казав, а тепер говорю навіть плачучи, поводяться, як вороги хреста Христового.
PHIL|3|19|Їхній кінець то загибіль, шлунок їхній бог, а слава в їхньому соромі... Вони думають тільки про земне!
PHIL|3|20|Життя ж наше на небесах, звідки ждемо й Спасителя, Господа Ісуса Христа,
PHIL|3|21|Який перемінить тіло нашого пониження, щоб стало подібне до славного тіла Його, силою, якою Він може і все підкорити Собі.
PHIL|4|1|Отож, мої браття улюблені, за якими так сильно тужу, моя радосте й вінче, так у Господі стійте, улюблені!
PHIL|4|2|Благаю Еводію, благаю й Синтихію думати однаково в Господі.
PHIL|4|3|Так, благаю й тебе, товаришу вірний, допомагай тим, хто в боротьбі за Євангелію помагали мені та Климентові й іншим моїм співробітникам, яких імення записані в Книзі Життя.
PHIL|4|4|Радійте в Господі завсіди, і знову кажу: радійте!
PHIL|4|5|Ваша лагідність хай буде відома всім людям. Господь близько!
PHIL|4|6|Ні про що не турбуйтесь, а в усьому нехай виявляються Богові ваші бажання молитвою й проханням з подякою.
PHIL|4|7|І мир Божий, що вищий від усякого розуму, хай береже серця ваші та ваші думки у Христі Ісусі.
PHIL|4|8|Наостанку, браття, що тільки правдиве, що тільки чесне, що тільки праведне, що тільки чисте, що тільки любе, що тільки гідне хвали, коли яка чеснота, коли яка похвала, думайте про це!
PHIL|4|9|Чого ви від мене й навчилися, і прийняли, і чули та бачили, робіть те! І Бог миру буде з вами!
PHIL|4|10|Я вельми потішився в Господі, що справді ви вже нових сил набули піклуватись про мене; ви й давніш піклувались, та часу сприятливого ви не мали.
PHIL|4|11|Не за нестатком кажу, бо навчився я бути задоволеним із того, що маю.
PHIL|4|12|Умію я й бути в упокоренні, умію бути й у достатку. Я привчився до всього й у всім: насищатися й голод терпіти, мати достаток і бути в недостачі.
PHIL|4|13|Я все можу в Тім, Хто мене підкріпляє, в Ісусі Христі.
PHIL|4|14|Тож ви добре зробили, що участь узяли в моїм горі.
PHIL|4|15|І знаєте й ви, филип'яни, що на початку благовістя, коли я з Македонії вийшов, не прилучилась була жадна Церква до справи давання й приймання для мене, самі тільки ви,
PHIL|4|16|що і раз, і вдруге мені на потреби мої посилали й до Солуня.
PHIL|4|17|Кажу це не тому, щоб шукав я давання, я шукаю плоду, що примножується на річ вашу.
PHIL|4|18|Та все я одержав, і маю достаток. Маю повно, прийнявши від Епафродита, що ви послали, як пахощі запашні, жертву приємну, Богові вгодну.
PHIL|4|19|А мій Бог нехай виповнить вашу всяку потребу за Своїм багатством у Славі, у Христі Ісусі.
PHIL|4|20|А Богові й нашому Отцеві слава на віки віків. Амінь.
PHIL|4|21|Вітайте кожного святого у Христі Ісусі. Вітають вас браття, присутні зо мною.
PHIL|4|22|Вітають вас усі святі, а найбільше ті, хто з кесаревого дому.
PHIL|4|23|Благодать Господа Ісуса Христа зо всіма вами! Амінь.
