COL|1|1|奉上帝旨意，作基督耶稣使徒的 保罗 ，和我们的弟兄 提摩太 ，
COL|1|2|写信给 歌罗西 的圣徒，在基督里忠心的弟兄。愿恩惠、平安 从我们的父上帝归给你们！
COL|1|3|我们为你们祷告的时候，常常感谢我们主耶稣基督的父上帝 ，
COL|1|4|因为听见你们对基督耶稣的信心，并对众圣徒有的爱心。
COL|1|5|这都是因着那给你们存在天上的盼望，它就是你们从前所听见真理的道，就是福音；
COL|1|6|这福音传到你们那里，也传到普天下，并且继续增长，不断结果，正如自从你们听见福音，真正知道上帝恩惠的日子起，在你们中间也是这样。
COL|1|7|这福音是你们从我们所亲爱、一同作仆人的 以巴弗 学到的。他为我们 作了基督的忠心仆役，
COL|1|8|也把圣灵赐给你们的爱告诉我们。
COL|1|9|因此，我们自从听见的日子就不住地为你们祷告和祈求，愿你们满有一切属灵的智慧和悟性，真正知道上帝的旨意，
COL|1|10|好使你们行事为人对得起主，凡事蒙他喜悦，在一切善事上结果子，对上帝的认识更有长进。
COL|1|11|愿你们从他荣耀的权能中，得以在一切事上力上加力，好使你们凡事欢欢喜喜地忍耐宽容，
COL|1|12|又感谢父，使你们配与众圣徒在光明中分享基业。
COL|1|13|他救了我们脱离黑暗的权势，迁移到他爱子的国度里。
COL|1|14|藉着他的爱子，我们得蒙救赎，罪得赦免。
COL|1|15|爱子是那看不见的上帝之像， 是首生的 ，在一切被造的以先。
COL|1|16|因为万有都是在他里面 造的， 无论是天上的、地上的， 能看见的、不能看见的， 或是有权位的、统治的， 或是执政的、掌权的， 一概都是藉着他为着他造的。
COL|1|17|他在万有之先； 万有也靠他而存在。
COL|1|18|他是身体（教会）的头； 他是元始， 是从死人中复活的首生者， 好让他在万有中居首位。
COL|1|19|因为上帝喜欢使一切的丰盛在他里面居住，
COL|1|20|藉着他 ，上帝使万有与自己和好， 无论是地上的、天上的， 都藉着他在十字架上所流的血促成了和平。
COL|1|21|从前你们与上帝隔绝，心思上与他为敌，行为邪恶；
COL|1|22|但如今，他藉着他儿子肉身的死，已经使你们与他自己和好了 ，把你们献在他的面前，成为圣洁，没有瑕疵，无可指责。
COL|1|23|只要你们持守信仰，根基稳固，坚定不移，不致动摇，离开了你们从前所听见的福音的盼望；这福音也是传给天下一切被造之物的，我— 保罗 作了这福音的仆役。
COL|1|24|现在我为你们受苦，倒很快乐；并且为基督的身体，就是为教会，我要在自己的肉身上补满基督未尽的苦难。
COL|1|25|我照上帝为你们所赐我的职分作了教会的仆役，要把上帝的道传得完满；
COL|1|26|这道就是历世历代所隐藏的奥秘，但如今向他的圣徒显明了。
COL|1|27|上帝要让他们知道，这奥秘在外邦人中有何等丰盛的荣耀；就是基督在你们心里 成了得荣耀的盼望。
COL|1|28|我们传扬他，是用诸般的智慧，劝戒各人，教导各人，要把各人在基督里完完全全地献上 。
COL|1|29|我也为此劳苦，照着他在我里面运用的大能尽心竭力。
COL|2|1|我要你们知道，我为你们和 老底嘉 人，和所有没有与我见过面的人，是何等地勤奋；
COL|2|2|为要使他们的心得安慰，因爱心互相联络，以致有从确实了解所产生的丰盛，好深知上帝的奥秘，就是基督；
COL|2|3|在他里面蕴藏着一切智慧和知识。
COL|2|4|我说这话，免得有人用花言巧语迷惑你们。
COL|2|5|虽然我身体不在你们那里，心却与你们同在，很高兴见你们循规蹈矩，对基督的信心也坚固。
COL|2|6|既然你们接受了主基督耶稣，就要靠着他而生活，
COL|2|7|照着你们所领受的教导，在他里面生根建造，信心坚固，充满着感谢的心。
COL|2|8|你们要谨慎，免得有人用他的哲学和虚空的废话，不照着基督，而是照人间的传统和世上粗浅的学说 ，把你们掳去。
COL|2|9|因为上帝本性一切的丰盛都有形有体地居住在基督里面；
COL|2|10|你们在他里面也已经成为丰盛。他是所有执政掌权者的元首。
COL|2|11|你们也在他里面受了不是人手所行的割礼，而是使你们脱去肉体情欲的基督的割礼。
COL|2|12|你们既受洗与他一同埋葬，也就在此礼上，因信那使他从死人中复活的上帝的作为跟他一同复活。
COL|2|13|你们从前在过犯和未受割礼的肉体中死了，上帝却赦免了你们一切的过犯，使你们与基督一同活过来，
COL|2|14|涂去了在律例上所写、敌对我们、束缚我们的字据，把它撤去，钉在十字架上。
COL|2|15|基督既将一切执政者、掌权者的权势解除了，就在凯旋的行列中，将他们公开示众，仗着十字架夸胜。
COL|2|16|所以，不要让任何人在饮食上，或节期、初一、安息日等事上评断你们。
COL|2|17|这些原是未来的事的影子，真体却是属基督的。
COL|2|18|不要让人藉着故作谦虚和敬拜天使夺去你们的奖赏。这等人拘泥在所见过的幻象 ，随着自己的欲望无故地自高自大，
COL|2|19|不紧随元首；其实，由于他全身藉着关节筋络才得到滋养，互相联络，靠上帝所赐的成长而成长。
COL|2|20|既然你们与基督同死而脱离了世上粗淺的学说，为什么仍像生活在世俗中一样，去服从那“不可拿、不可尝、不可摸”等类的规条呢？
COL|2|21|
COL|2|22|这些都是根据人的命令和教导，论到这一切都是一经使用就都败坏了。
COL|2|23|这些规条使人徒有智慧之名，用私意崇拜，自表谦卑，苦待己身，其实在克制肉体的情欲上毫无功效。
COL|3|1|所以，既然你们已经与基督一同复活，就当求上面的事；那里有基督，坐在上帝的右边。
COL|3|2|你们要思考上面的事，不要思考地上的事。
COL|3|3|因为你们已经死了，你们的生命与基督一同藏在上帝里面。
COL|3|4|基督是你们的生命，他显现的时候，你们也要与他一同在荣耀里显现。
COL|3|5|所以，要治死你们在地上的肢体；就如淫乱、污秽、邪情、恶欲和贪婪—贪婪就是拜偶像。
COL|3|6|因这些事，上帝的愤怒必临到那些悖逆的人 。
COL|3|7|当你们在这些事中活着的时候，你们的行为也曾是这样的。
COL|3|8|但现在你们要弃绝这一切的事，就是恼恨、愤怒、恶毒、毁谤和口中污秽的言语。
COL|3|9|不要彼此说谎，因为你们已经脱去旧人和旧人的行为，
COL|3|10|穿上了新人，这新人照着造他的主的形像在知识上不断地更新。
COL|3|11|在这事上并不分 希腊 人和 犹太 人，受割礼的和未受割礼的，未开化的人、 西古提 人、为奴的、自主的；惟独基督是一切，又在一切之内。
COL|3|12|所以，你们既是上帝的选民，圣洁、蒙爱的人，要穿上怜悯、恩慈、谦虚、温柔和忍耐。
COL|3|13|倘若这人与那人有嫌隙，总要彼此容忍，彼此饶恕；主 怎样饶恕了你们，你们也要怎样饶恕人。
COL|3|14|除此以外，还要穿上爱心，因为爱是贯通全德的。
COL|3|15|你们要让基督所赐的和平在你们心里作主，也为此蒙召，归为一体。你们还要存感谢的心。
COL|3|16|当用各样的智慧，把基督的道丰丰富富的存在心里，用诗篇、赞美诗、灵歌，彼此教导，互相劝戒，以感恩的心歌颂上帝。
COL|3|17|你们无论做什么，或说话或行事，都要奉主耶稣的名，藉着他感谢父上帝。
COL|3|18|你们作妻子的，要顺服自己的丈夫，这在主里面是合宜的。
COL|3|19|你们作丈夫的，要爱你们的妻子，不可虐待她们。
COL|3|20|你们作儿女的，要凡事听从父母，因为这是主所喜悦的。
COL|3|21|你们作父亲的，不要惹儿女生气，恐怕他们会灰心。
COL|3|22|你们作仆人的，要凡事听从你们肉身的主人，不要只在眼前服事，像是讨人喜欢的，总要心存诚实，因为你们敬畏主。
COL|3|23|你们无论做什么，都要从心里做，像是为主做的，不是为人做的；
COL|3|24|因为你们知道，从主那里必得着基业作为赏赐。你们要服侍的是主基督。
COL|3|25|行不义的人必受不义的报应；主并不偏待人。
COL|4|1|你们作主人的，待仆人要公正，因为知道，你们也有一位主在天上。
COL|4|2|你们要恒切祷告，在祷告中警醒感恩。
COL|4|3|同时，也要为我们祷告，求上帝给我们开传道的门，能宣讲基督的奥秘，
COL|4|4|使我能按着所该说的话将这奥秘显明出来，我为此而被捆锁。
COL|4|5|你们要把握时机，用智慧与外人来往。
COL|4|6|你们的言谈要时常带着温和，好像用盐调味，让你们知道该怎样应对每一个人。
COL|4|7|推基古 是我亲爱的弟兄，忠心的仆役，和我一同作主的仆人；他要把我一切的事都告诉你们。
COL|4|8|我特意打发他到你们那里去，好让你们知道我们的情况，又让他安慰你们的心。
COL|4|9|我又打发一位亲爱忠心的弟兄 阿尼西谋 同去；他也是你们那里的人。他们会把这里一切的事都告诉你们。
COL|4|10|与我一同坐牢的 亚里达古 问候你们。 巴拿巴 的表弟 马可 也问候你们。关于他，你们已经得到指示；他若到你们那里，你们要接待他。
COL|4|11|称为 犹士都 的 耶数 也问候你们。奉割礼的人中，只有这三个人是为上帝的国与我作同工的，也是使我心里得安慰的。
COL|4|12|有一位你们那里的人，作基督耶稣 仆人的 以巴弗 问候你们。他祷告的时候常为你们竭力祈求，愿你们能站稳而成熟，充分确信上帝一切的旨意。
COL|4|13|他为你们、 老底嘉 和 希拉坡里 的弟兄多多劳苦，这是我可以为他作见证的。
COL|4|14|亲爱的医生 路加 和 底马 问候你们。
COL|4|15|请问候 老底嘉 的弟兄以及 宁法 ，和她家里 的教会。
COL|4|16|你们宣读了这书信，也要交给 老底嘉 的教会宣读；你们也要宣读从 老底嘉 转来的书信。
COL|4|17|你们要对 亚基布 说：“务要完成你从主所领受的职分。”
COL|4|18|我— 保罗 亲笔问候你们。要记念我在捆锁中。愿恩惠与你们同在！
