JUDG|1|1|约书亚 死后， 以色列 人求问耶和华说：“我们中间谁当首先上去攻打 迦南 人，与他们争战呢？”
JUDG|1|2|耶和华说：“ 犹大 要先上去。看哪，我已将那地交在他手中。”
JUDG|1|3|犹大 对他哥哥 西缅 说：“请你同我上到我抽签所得之地，与 迦南 人争战；我也同你去你抽签所得之地。”于是 西缅 与他同去。
JUDG|1|4|犹大 就上去，耶和华把 迦南 人和 比利洗 人交在他们手中。他们在 比色 击杀了一万人。
JUDG|1|5|他们在 比色 遇见 亚多尼．比色 ，与他争战，击败了 迦南 人和 比利洗 人。
JUDG|1|6|亚多尼．比色 逃跑，他们追赶他，捉住他，砍断他大拇指和大脚趾。
JUDG|1|7|亚多尼．比色 说：“从前有七十个王，大拇指和大脚趾都被我砍断，在我桌子底下拾取零碎食物。现在上帝照着我所做的报应我了。”他们把 亚多尼．比色 带到 耶路撒冷 ，他就死在那里。
JUDG|1|8|犹大 人攻打 耶路撒冷 ，夺取了它，用刀杀城内的人，并且放火烧城。
JUDG|1|9|后来 犹大 人下去，与住山区、 尼革夫 和低地的 迦南 人争战。
JUDG|1|10|犹大 去攻打住 希伯仑 的 迦南 人，杀了 示筛 、 亚希幔 、 挞买 。 希伯仑 从前名叫 基列．亚巴 。
JUDG|1|11|犹大 从那里去攻击 底壁 的居民。 底壁 从前名叫 基列．西弗 。
JUDG|1|12|迦勒 说：“谁能攻打 基列．西弗 ，夺取那城，我就把我女儿 押撒 嫁给他。”
JUDG|1|13|迦勒 的弟弟 基纳斯 的儿子 俄陀聂 夺取了那城， 迦勒 就把女儿 押撒 嫁给他。
JUDG|1|14|押撒 来的时候，催促丈夫 向她父亲要一块田。 押撒 一下驴， 迦勒 就对她说：“你要什么？”
JUDG|1|15|她对 迦勒 说：“求你赐我福分；你既然把 尼革夫 给了我，求你也给我水泉。” 迦勒 就把上泉和下泉都赐给她。
JUDG|1|16|摩西 的岳父是 基尼 人，他的子孙与 犹大 人一起上到棕树城，往 亚拉得 以南的 犹大 旷野 去，住在百姓当中 。
JUDG|1|17|犹大 和他哥哥 西缅 同去，击杀了住 洗法 的 迦南 人，将城彻底毁灭。因此，那城名叫 何珥玛 。
JUDG|1|18|犹大 攻取了 迦萨 和所属的领土， 亚实基伦 和所属的领土， 以革伦 和所属的领土。
JUDG|1|19|耶和华与 犹大 同在， 犹大 取得了山区，却不能赶出平原的居民，因为他们有铁的战车。
JUDG|1|20|以色列 人照 摩西 所说的，把 希伯仑 给了 迦勒 。 迦勒 从那里赶出 亚衲 的三支后裔。
JUDG|1|21|至于住 耶路撒冷 的 耶布斯 人， 便雅悯 人没有把他们赶出。于是， 耶布斯 人与 便雅悯 人同住在 耶路撒冷 ，直到今日。
JUDG|1|22|约瑟 家也上到 伯特利 去，耶和华与他们同在。
JUDG|1|23|约瑟 家去窥探 伯特利 ，那城起先名叫 路斯 。
JUDG|1|24|探子看见一个人从城里出来，就对他说：“请你把进城的路指示我们，我们会厚待你。”
JUDG|1|25|那人把进城的路指示他们。他们就用刀击杀了城中的居民，却放走那人和他的全家。
JUDG|1|26|那人往 赫 人之地去，建造了一座城，起名叫 路斯 。那城到如今还叫这名。
JUDG|1|27|玛拿西 没有赶出 伯˙善 和所属乡镇 的居民， 他纳 和所属乡镇的居民， 多珥 和所属乡镇的居民， 以伯莲 和所属乡镇的居民， 米吉多 和所属乡镇的居民； 迦南 人仍坚持住在这地。
JUDG|1|28|以色列 强盛的时候，就叫 迦南 人做苦工，没有把他们全然赶走。
JUDG|1|29|以法莲 没有赶出住 基色 的 迦南 人。于是 迦南 人仍住在 基色 ，在 以法莲 中间。
JUDG|1|30|西布伦 没有赶出 基伦 的居民和 拿哈拉 的居民。于是 迦南 人仍住在 西布伦 中间，成了服劳役的人。
JUDG|1|31|亚设 没有赶出 亚柯 的居民和 西顿 的居民，以及 亚黑拉 、 亚革悉 、 黑巴 、 亚弗革 和 利合 的居民。
JUDG|1|32|亚设 人因为没有赶出那地的居民 迦南 人，就住在他们中间。
JUDG|1|33|拿弗他利 没有赶出 伯˙示麦 和 伯˙亚纳 的居民。于是 拿弗他利 就住在那地的居民 迦南 人中，而 伯˙示麦 和 伯˙亚纳 的居民却成了为他们服劳役的人。
JUDG|1|34|亚摩利 人强逼 但 人住在山区，不准他们下到平原。
JUDG|1|35|亚摩利 人仍坚持住在 希烈山 、 亚雅仑 和 沙宾 ；然而 约瑟 家权势强盛的时候，他们成为服劳役的人。
JUDG|1|36|亚摩利 人 的地界是从 亚克拉滨 斜坡，从 西拉 延伸而上。
JUDG|2|1|耶和华的使者从 吉甲 上到 波金 ，说：“我领你们从 埃及 上来，带你们到我向你们列祖起誓应许之地。我曾说：‘我永不废弃我与你们的约。
JUDG|2|2|你们不可与这地的居民立约，要拆毁他们的祭坛。’你们竟没有听从我的话。你们为何这样做呢！
JUDG|2|3|因此我说：‘我必不将他们从你们面前赶出。他们必作你们肋下的荆棘 ，他们的神明必成为你们的圈套。’”
JUDG|2|4|耶和华的使者向 以色列 众人说这些话的时候，百姓放声大哭。
JUDG|2|5|于是他们给那地方起名叫 波金 ，并在那里向耶和华献祭。
JUDG|2|6|约书亚 解散百姓， 以色列 人回到自己的地业，占各自的地。
JUDG|2|7|约书亚 在世的日子和他死了以后，那些见过耶和华为 以色列 所做一切大事的长老还在世的时候，百姓都事奉耶和华。
JUDG|2|8|耶和华的仆人， 嫩 的儿子 约书亚 死了，那时他一百一十岁。
JUDG|2|9|以色列 人把他葬在他自己地业的境内， 以法莲 山区的 亭拿．希烈 ，在 迦实山 的北边。
JUDG|2|10|那世代的人也都归到自己的列祖。后来兴起的另一世代不认识耶和华，也不知道他为 以色列 所做的事。
JUDG|2|11|以色列 人行耶和华眼中看为恶的事，去事奉诸 巴力 。
JUDG|2|12|他们离弃领他们出 埃及 地的耶和华－他们列祖的上帝，去随从别神，就是四围列国的神明，向它们叩拜，惹耶和华发怒。
JUDG|2|13|他们离弃了耶和华，去事奉 巴力 和 亚斯她录 。
JUDG|2|14|耶和华的怒气向 以色列 发作，把他们交在抢夺他们的人手中，又把他们交给四围仇敌的手中 ，以致他们在仇敌面前再也不能站立得住。
JUDG|2|15|他们无论往何处去，耶和华的手都以灾祸攻击他们，正如耶和华所说的，又如耶和华向他们所起的誓；他们就极其困苦。
JUDG|2|16|耶和华兴起士师，士师就拯救他们脱离抢夺他们之人的手。
JUDG|2|17|然而，他们却不听从士师，竟随从别神而行淫，向它们叩拜。他们列祖所行的道，所听从耶和华的命令，他们都速速偏离了，并不照样遵行。
JUDG|2|18|耶和华为他们兴起士师，耶和华与士师同在。士师在世的一切日子，耶和华拯救他们脱离仇敌的手。耶和华因他们受欺压迫害所发出的哀声，就怜悯他们。
JUDG|2|19|但士师一死，他们又转去行恶，比他们祖宗更坏，去随从别神，事奉叩拜它们，总不放弃他们的恶习和顽梗的行为。
JUDG|2|20|于是耶和华的怒气向 以色列 发作，说：“因为这国违背我吩咐他们列祖当守的约，不听从我的话，
JUDG|2|21|约书亚 死的时候所剩下的各国，我必不再从他们面前赶出任何一个，
JUDG|2|22|为要藉此考验 以色列 是否肯谨守遵行耶和华的道，像他们列祖一样地谨守。”
JUDG|2|23|耶和华留下那些国家，不将他们速速赶出，也不把他们交在 约书亚 的手中。
JUDG|3|1|耶和华留下这些国家，为要考验所有未曾经历 迦南 任何战役的 以色列 人，
JUDG|3|2|只是为了要 以色列 人的后代认识战争，教导他们，尤其那些未曾认识这些事的人。
JUDG|3|3|留下的有 非利士 的五个领袖，所有的 迦南 人， 西顿 人，以及从 巴力．黑门山 到 哈马口 ，住 黎巴嫩山 的 希未 人。
JUDG|3|4|他们是为了要考验 以色列 ，好知道他们是否肯听从耶和华藉 摩西 吩咐他们列祖的命令。
JUDG|3|5|以色列 人住在 迦南 人、 赫 人、 亚摩利 人、 比利洗 人、 希未 人、 耶布斯 人中间，
JUDG|3|6|娶他们的女儿，将自己的女儿嫁给他们的儿子，并事奉他们的神明。
JUDG|3|7|以色列 人行耶和华眼中看为恶的事，忘记耶和华－他们的上帝，去事奉诸 巴力 和 亚舍拉 ，
JUDG|3|8|所以耶和华的怒气向 以色列 发作，把他们交给 美索不达米亚 王 古珊．利萨田 的手中。 以色列 人服事 古珊．利萨田 八年。
JUDG|3|9|以色列 人呼求耶和华，耶和华就为 以色列 人兴起一位拯救者来救他们，就是 迦勒 的弟弟 基纳斯 的儿子 俄陀聂 。
JUDG|3|10|耶和华的灵降在他身上，他就作了 以色列 的士师。他出去争战，耶和华将 亚兰 王 古珊．利萨田 交在他手中，他的手战胜了 古珊．利萨田 。
JUDG|3|11|于是这地太平四十年。 基纳斯 的儿子 俄陀聂 死了。
JUDG|3|12|以色列 人又行耶和华眼中看为恶的事。耶和华使 摩押 王 伊矶伦 强大，攻击 以色列 ，因为他们行耶和华眼中看为恶的事。
JUDG|3|13|伊矶伦 召集 亚扪 人和 亚玛力 人到他那里，他就去攻打 以色列 ，占据了棕树城。
JUDG|3|14|于是 以色列 人服事 摩押 王 伊矶伦 十八年。
JUDG|3|15|以色列 人呼求耶和华，耶和华就为他们兴起一位拯救者， 便雅悯 人 基拉 的儿子 以笏 ，他是个惯用左手的人 。 以色列 人托他送礼物给 摩押 王 伊矶伦 。
JUDG|3|16|以笏 打造了一把两刃的剑，长一短肘 ，绑在右腿上衣服里面。
JUDG|3|17|他把礼物献给 摩押 王 伊矶伦 。 伊矶伦 是个很肥胖的人。
JUDG|3|18|以笏 献完礼物的时候，就把抬礼物的人送走。
JUDG|3|19|但他自己却从靠近 吉甲 的雕像那里转回来，说：“王啊，我有一件机密的事要奏告你。”王说：“回避吧！”于是所有侍立在他左右的人都退去了。
JUDG|3|20|以笏 来到王那里，那时他独自一人坐在阴凉的顶楼。 以笏 说：“我有上帝的话向你报告。”王就从座位上站起来。
JUDG|3|21|以笏 伸出左手，从右腿上拔出剑来，刺入王的肚腹。
JUDG|3|22|剑柄连同剑刃都刺进去了，肥肉夹住了剑刃。他没有把剑从王的肚腹拔出来，粪便就流出来了 。
JUDG|3|23|以笏 出到门廊，把王关在楼门里面，就上了锁。
JUDG|3|24|以笏 出来之后，王的仆人就来了。他们观看，看哪，楼门锁住，就说：“他必是在阴凉的房间里大解。”
JUDG|3|25|他们等得不耐烦，看哪，楼门仍然不开，就拿钥匙打开楼门，看哪，他们的主人已经倒在地上死了。
JUDG|3|26|他们耽延的时候， 以笏 就逃跑了。他经过雕像那里，逃到 西伊拉 。
JUDG|3|27|他到了那里，就在 以法莲 山区吹角。 以色列 人跟随他从山区下来，他在他们前面引路，
JUDG|3|28|对他们说：“紧跟着我！因为耶和华已经把你们的仇敌 摩押 交在你们手中。”于是他们跟着他下去，占据了 摩押 对面 约旦河 的渡口，不准一人过去。
JUDG|3|29|那时，他们击杀了约一万 摩押 人，都是强壮的勇士，连一个也没有逃脱。
JUDG|3|30|那日， 摩押 在 以色列 手下制伏了。于是这地太平八十年。
JUDG|3|31|以笏 之后，有 亚拿 的儿子 珊迦 ，他用赶牛的棍子打死六百 非利士 人。他也拯救了 以色列 。
JUDG|4|1|以笏 死后， 以色列 人又行耶和华眼中看为恶的事。
JUDG|4|2|耶和华把他们交给在 夏琐 作王的 迦南 王 耶宾 手中；他的将军是 西西拉 ，住在 夏罗设．哈歌印 。
JUDG|4|3|以色列 人呼求耶和华，因为 耶宾 王有铁的战车九百辆，并且残酷欺压 以色列 人二十年。
JUDG|4|4|有一位女先知 底波拉 ，是 拉比多 的妻子，当时作 以色列 的士师。
JUDG|4|5|她住在 以法莲 山区 拉玛 和 伯特利 的中间，在 底波拉 的棕树下。 以色列 人都上到她那里去听审判。
JUDG|4|6|她派人从 拿弗他利 的 基低斯 把 亚比挪庵 的儿子 巴拉 召来，对他说：“耶和华－ 以色列 的上帝吩咐你：‘你要率领一万 拿弗他利 人和 西布伦 人上 他泊山 去。
JUDG|4|7|我必使 耶宾 的将军 西西拉 率领他的战车和全军往 基顺河 ，到你那里去，我必把他交在你手中。’”
JUDG|4|8|巴拉 对她说：“你若同我去，我就去；你若不同我去，我就不去。”
JUDG|4|9|底波拉 说：“我一定会与你同去，然而你在所行的路上必得不着荣耀，因为耶和华要把 西西拉 交给一个妇人的手里。”于是 底波拉 起来，与 巴拉 一同往 基低斯 去了。
JUDG|4|10|巴拉 召集 西布伦 人和 拿弗他利 人到 基低斯 ，跟他上去的有一万人。 底波拉 也同他上去。
JUDG|4|11|摩西 岳父 何巴 的后裔， 基尼 人 希百 离开了 基尼 族，到靠近 基低斯 的 撒拿音 橡树旁支搭帐棚。
JUDG|4|12|有人告诉 西西拉 ：“ 亚比挪庵 的儿子 巴拉 已经上了 他泊山 。”
JUDG|4|13|西西拉 就召集所有的铁战车九百辆和随从的全军，从 夏罗设．哈歌印 出来，到了 基顺河 。
JUDG|4|14|底波拉 对 巴拉 说：“起来，今日就是耶和华把 西西拉 交在你手中的日子。耶和华岂不在你前面行吗总”于是 巴拉 下了 他泊山 ，跟随他的有一万人。
JUDG|4|15|耶和华使 西西拉 和他一切的战车，以及全军溃乱，在 巴拉 面前倒在刀下。 西西拉 下了车，徒步逃跑。
JUDG|4|16|巴拉 追赶战车、军队，直到 夏罗设．哈歌印 。 西西拉 的全军都倒在刀下，一个也没有留下。
JUDG|4|17|只有 西西拉 徒步逃跑到 基尼 人 希百 之妻 雅亿 的帐棚，因为 夏琐 王 耶宾 与 基尼 人的 希百 家和平共处。
JUDG|4|18|雅亿 出来迎接 西西拉 ，对他说：“请我主进来，进到我这里来，不要怕。” 西西拉 就进了她的帐棚， 雅亿 用被子将他盖住。
JUDG|4|19|西西拉 对 雅亿 说：“我渴了，求你给我一点水喝。” 雅亿 就打开装奶的皮袋，给他喝，再把他盖住。
JUDG|4|20|西西拉 对 雅亿 说：“请你站在帐棚门口，若有人来问你说：‘有人在这里吗？’你就说：‘没有。’”
JUDG|4|21|西西拉 疲乏沉睡了。 希百 的妻 雅亿 取了帐棚的橛子，手拿着锤子，静悄悄地到他那里，将橛子从他的太阳穴钉进去，直钉到地里。 西西拉 就死了。
JUDG|4|22|看哪， 巴拉 追赶 西西拉 ， 雅亿 出来迎接他，对他说：“来，我给你看你要找的人。”他就进入帐棚，看哪， 西西拉 已经倒在地上死了，橛子还在他的太阳穴中。
JUDG|4|23|那日，上帝在 以色列 人面前制伏了 迦南 王 耶宾 。
JUDG|4|24|从此， 以色列 人的手对 迦南 王 耶宾 越来越强硬，直到将 迦南 王 耶宾 剪除。
JUDG|5|1|那日， 底波拉 和 亚比挪庵 的儿子 巴拉 唱歌，说：
JUDG|5|2|“ 以色列 有领袖率领 ， 百姓甘心牺牲自己， 你们当称颂耶和华！
JUDG|5|3|“君王啊，要听！王子啊，要侧耳！ 我要，我要向耶和华歌唱； 我要歌颂耶和华－ 以色列 的上帝。
JUDG|5|4|“耶和华啊，你从 西珥 出来， 从 以东 田野向前行， 地震动 天滴下， 云也滴下雨水。
JUDG|5|5|众山在耶和华面前摇动， 西奈山 在耶和华－ 以色列 上帝面前也摇动。
JUDG|5|6|“在 亚拿 之子 珊迦 的时候， 在 雅亿 的日子， 大道无人行走， 过路人绕道而行。
JUDG|5|7|以色列 农村荒芜， 空无一人， 直到我 底波拉 兴起， 兴起作 以色列 之母！
JUDG|5|8|以色列 人选择新的诸神， 战争就临到城门。 以色列 四万人中， 看得见盾牌枪矛吗？
JUDG|5|9|我心向往 以色列 的领袖， 他们在民中甘心牺牲自己。 你们应当称颂耶和华！
JUDG|5|10|“骑浅色母驴的、 坐绣花毯子的、 行走在路上的， 你们都当思想！
JUDG|5|11|打水的声音胜过弓箭的响声， 那里，人要述说耶和华公义的作为， 他对 以色列 乡民公义的作为。 “那时，耶和华的子民下到城门。
JUDG|5|12|“ 底波拉 啊，兴起！兴起！ 当兴起，兴起，唱歌！ 巴拉 啊，你当兴起！ 亚比挪庵 的儿子啊，当俘掳你的俘虏！
JUDG|5|13|那时，贵族中的幸存者前进， 耶和华的百姓为我前进攻击勇士。
JUDG|5|14|源自 亚玛力 的人从 以法莲 下来 ， 跟着你，你的族人 便雅悯 ； 有领袖从 玛吉 下来， 手握官员权杖的从 西布伦 下来。
JUDG|5|15|以萨迦 的领袖与 底波拉 一起； 巴拉 怎样， 以萨迦 也怎样； 他跟随 巴拉 冲下平原。 吕便 支派 有胸怀大志的人。
JUDG|5|16|你为何坐在羊圈内， 听羊群中吹笛的声音呢？ 吕便 支派具心有大谋的人。
JUDG|5|17|基列 安居在 约旦河 东。 但 为何住在船上呢？ 亚设 在海边居住， 它在港口安居。
JUDG|5|18|西布伦 是拚命敢死的百姓， 拿弗他利 在田野的高处也是如此。 　
JUDG|5|19|“君王都来争战； 那时 迦南 诸王在 米吉多 水旁的 他纳 争战， 却得不到掳掠的银钱。
JUDG|5|20|星宿从天上争战， 从它们的轨道攻击 西西拉 。
JUDG|5|21|基顺 的急流冲走他们， 古老的急流， 基顺 的急流。 我的灵啊，努力前进！
JUDG|5|22|“那时马蹄踢踏， 壮马奔驰飞腾。
JUDG|5|23|“耶和华的使者说：‘要诅咒 米罗斯 ， 重重诅咒其中的居民， 因为他们不来帮助耶和华， 不来帮助耶和华攻击壮士。’
JUDG|5|24|“愿 基尼 人 希百 的妻子 雅亿 比众妇人多得福气， 比帐棚中的妇人更蒙福祉。
JUDG|5|25|西西拉 求水， 雅亿 给他奶， 用贵重的碗装乳酪给他。
JUDG|5|26|雅亿 左手拿着帐棚的橛子， 右手拿着工匠的锤子， 击打 西西拉 ，打碎他的头， 打破穿透他的太阳穴。
JUDG|5|27|西西拉 在她脚下曲身，仆倒，躺卧， 在她脚下曲身，仆倒； 他在哪里曲身，就在哪里仆倒，死亡。
JUDG|5|28|“ 西西拉 的母亲从窗户里往外观看， 她在窗格子中哀号： ‘他的战车为何迟迟未归？ 他的车轮为何走得那么慢呢？’
JUDG|5|29|她聪明的宫女回答她， 她也自言自语说：
JUDG|5|30|‘或许他们得了战利品而分， 每个壮士得了一两个女子？ 西西拉 得了彩衣为掳物， 得了绣花的彩衣为掠物， 这两面绣花的彩衣， 披在颈项上作为战利品。’
JUDG|5|31|“耶和华啊，愿你的仇敌都这样灭亡！ 愿爱你的人如太阳上升，大发光辉！” 于是这地太平四十年。
JUDG|6|1|以色列 人又行耶和华眼中看为恶的事，耶和华就把他们交在 米甸 手里七年。
JUDG|6|2|米甸 的手战胜 以色列 ； 以色列 人躲避 米甸 人，就在山中挖洞穴，挖洞建营寨。
JUDG|6|3|每当 以色列 人撒种之后， 米甸 、 亚玛力 和东边的人都上来攻打他们，
JUDG|6|4|对着他们安营，毁坏那地的农作物，直到 迦萨 ，没有给 以色列 留下食物，牛、羊、驴也没有留下。
JUDG|6|5|因为那些人带着他们的牲畜和帐棚上来，像蝗虫那样多；人和骆驼无数，都进入境内，毁坏全地。
JUDG|6|6|以色列 因 米甸 的缘故极其穷乏， 以色列 人就呼求耶和华。
JUDG|6|7|以色列 人因 米甸 的缘故呼求耶和华的时候，
JUDG|6|8|耶和华就差遣先知到 以色列 人那里，对他们说：“耶和华－ 以色列 的上帝如此说：‘我曾领你们从 埃及 上来，从为奴之家出来，
JUDG|6|9|救你们脱离 埃及 人的手，脱离一切欺压你们之人的手。我从你们面前赶出他们，把他们的地赐给你们。
JUDG|6|10|我对你们说，我是耶和华－你们的上帝。你们住在 亚摩利 人的地，不可敬畏他们的神明，但你们却不听从我的话。’”
JUDG|6|11|耶和华的使者到了 俄弗拉 ，坐在 亚比以谢 族 约阿施 的橡树下。 约阿施 的儿子 基甸 正在醡酒池那里打麦子，为了躲避 米甸 人。
JUDG|6|12|耶和华的使者向 基甸 显现，对他说：“大能的勇士啊，耶和华与你同在！”
JUDG|6|13|基甸 对他说：“主啊，请容许我说，耶和华若与我们同在，我们怎么会遭遇这一切事呢？我们的列祖告诉我们：‘耶和华领我们从 埃及 上来’，他那奇妙的作为在哪里呢？现在耶和华却丢弃了我们，把我们交在 米甸 人的手掌中。”
JUDG|6|14|耶和华转向 基甸 ，说：“去，靠着你这能力拯救 以色列 脱离 米甸 人的手掌。我岂不是已经差遣了你吗？”
JUDG|6|15|基甸 对他说：“主啊，请容许我说，我怎能拯救 以色列 呢？看哪，我这一支在 玛拿西 支派中是最贫寒的，我在我父家又是最微小的。”
JUDG|6|16|耶和华对他说：“我与你同在，你就必击败 米甸 ，如击打一个人。”
JUDG|6|17|基甸 对他说：“我若在你眼前蒙恩，求你给我一个证据，证明是你在跟我说话。
JUDG|6|18|求你不要离开这里，等我回来，将供物带来，供在你面前。”他说：“我必等你回来。”
JUDG|6|19|基甸 去预备一只小山羊，用一伊法细面做了无酵饼，将肉放在篮子里，将汤盛在壶中，带到他那里，在橡树下献上。
JUDG|6|20|上帝的使者对 基甸 说：“将肉和无酵饼放在这磐石上，把汤倒出来。”他就照样做了。
JUDG|6|21|耶和华的使者伸出手里的杖，杖头一碰到肉和无酵饼，就有火从磐石中出来，吞灭了肉和无酵饼。耶和华的使者就从他眼前消失了。
JUDG|6|22|基甸 见他是耶和华的使者，就说：“哎呀！主耶和华啊！因为我真的面对面看见了耶和华的使者。”
JUDG|6|23|耶和华对他说：“安心吧，不要怕，你不会死。”
JUDG|6|24|于是 基甸 在那里为耶和华筑了一座坛，起名叫“耶和华沙龙” 。这坛至今还在 亚比以谢 族的 俄弗拉 。
JUDG|6|25|那夜，耶和华对 基甸 说：“你要把你父亲的公牛，就是 那七岁的第二头公牛取来，并拆毁你父亲为 巴力 筑的坛，砍下坛旁的 亚舍拉 ，
JUDG|6|26|在这堡垒顶上整整齐齐地为耶和华－你的上帝筑一座坛，将第二头公牛献为燔祭，用你所砍下的 亚舍拉 当柴。”
JUDG|6|27|基甸 就从他仆人中选了十个人，照耶和华吩咐他的做了。他因怕父家和本城的人，不敢在白天做这事，就在夜间做。
JUDG|6|28|城里的人清早起来，看哪， 巴力 的坛被拆毁，坛旁的 亚舍拉 被砍下，第二头公牛献在筑好的坛上，
JUDG|6|29|就彼此问：“这是谁做的事呢？”他们寻找查访之后，就说：“这是 约阿施 的儿子 基甸 做的事。”
JUDG|6|30|城里的人对 约阿施 说：“把你的儿子交出来，我们要处死他，因为他拆毁了 巴力 的坛，砍下了坛旁的 亚舍拉 。”
JUDG|6|31|约阿施 对站着敌对他的众人说：“你们是为 巴力 辩护吗？你们要救它吗？谁为它辩护，就在早晨把谁处死吧！ 巴力 如果是上帝，有人拆毁了它的坛，就让它为自己辩护吧！”
JUDG|6|32|所以那日人称 基甸 为 耶路巴力 ，意思是：“他拆毁了 巴力 的坛，让 巴力 与他争辩吧。”
JUDG|6|33|那时，所有的 米甸 人、 亚玛力 人和东边的人都聚集在一起，过了河，在 耶斯列 平原安营。
JUDG|6|34|耶和华的灵降在 基甸 身上；他吹角， 亚比以谢 族都聚集跟随他。
JUDG|6|35|他派使者走遍 玛拿西 ， 玛拿西 人也聚集跟随他。他又派使者到 亚设 、 西布伦 、 拿弗他利 ，他们也都上来会合。
JUDG|6|36|基甸 对上帝说：“你如果真的照你所说的，藉我的手拯救 以色列 ，
JUDG|6|37|看哪，我把一团羊毛放在禾场上，若单是羊毛上有露水，遍地都是干的，我就知道你必照你所说的，藉我的手拯救 以色列 。”
JUDG|6|38|一切果然发生了。次日早晨 基甸 起来，把羊毛拧一拧，从羊毛中挤出露水来，装满一碗的水。
JUDG|6|39|基甸 又对上帝说：“求你不要向我发怒，我再说一次，让我用羊毛再试一次，但愿羊毛是干的，遍地都有露水。”
JUDG|6|40|这夜，上帝也照样做，遍地都有露水，只有羊毛是干的。
JUDG|7|1|耶路巴力 ，就是 基甸 ，和所有跟随他的人早晨起来，在 哈律泉 旁安营。 米甸 营在他北边，靠近 摩利冈 的平原。
JUDG|7|2|耶和华对 基甸 说：“跟随你的人太多，我不能把 米甸 交在他们手中，免得 以色列 向我自夸，说：‘是我自己的手救了我。’
JUDG|7|3|现在你要向这百姓宣告说：‘凡惧怕战兢的，可以离开 基列山 回去。’”于是有二万二千人回去，只剩下一万人。
JUDG|7|4|耶和华对 基甸 说：“人还是太多。你要带他们下到水旁，我好在那里为你试试他们。我指着谁对你说：‘这人可以跟你去’，他就可以跟你去；我指着谁对你说：‘这人不可跟你去’，他就不可跟你去。”
JUDG|7|5|基甸 就带百姓下到水旁。耶和华对 基甸 说：“凡用舌头舔水像狗一样舔的，要使他单独站在一处；那些用双膝跪下喝水的，也要使他单独站在一处。”
JUDG|7|6|用手捧到嘴边舔水的数目有三百人，其余的百姓都用双膝跪下喝水。
JUDG|7|7|耶和华对 基甸 说：“我要用这舔水的三百人拯救你们，把 米甸 交在你手中；其余的百姓都可以各回自己的地方去。”
JUDG|7|8|百姓手里拿着食物和角；其余的 以色列 人， 基甸 都打发他们各自回到自己的帐棚，只留下这三百人。 米甸 营在他下边的平原上。
JUDG|7|9|那夜，耶和华对 基甸 说：“起来，下去攻营，因我已把它交在你手中。
JUDG|7|10|倘若你害怕下去，可以带你的仆人 普拉 下到那营里去，
JUDG|7|11|你必听见他们所说的，这样你的手就有力量下去攻营。”于是 基甸 带着仆人 普拉 下到军营里带着兵器的人边上。
JUDG|7|12|米甸 人、 亚玛力 人和所有东边的人都散布在平原，如同蝗虫那样多。他们的骆驼无数，多如海边的沙。
JUDG|7|13|基甸 到了那里，看哪，有一人把梦告诉同伴说：“看哪，我做了一个梦。看哪，一个大麦饼滚入 米甸 营中，来到帐幕，把帐幕撞倒，帐幕就翻转倒塌了。”
JUDG|7|14|同伴回答说：“这不是别的，而是 以色列 人 约阿施 的儿子 基甸 的刀。上帝已把 米甸 和全军都交在他手中了。”
JUDG|7|15|基甸 听见这梦的叙述和梦的解释，就敬拜上帝。他回到 以色列 营中，说：“起来吧！耶和华已把 米甸 军队交在你们手中了。”
JUDG|7|16|于是 基甸 将三百人分成三队，把角和空瓶交在每个人手中，瓶内有火把。
JUDG|7|17|他对他们说：“看着我，你们要照样做。看哪，我来到营边，我怎样做，你们也要照样做。
JUDG|7|18|我和所有跟随我的人吹角的时候，你们也要在营的四围吹角，喊叫：‘为耶和华！为 基甸 ！’”
JUDG|7|19|基甸 和跟随他的一百人，在半夜之初换岗哨的时候来到营旁。他们就吹角，打破手中的瓶；
JUDG|7|20|三队的人都吹角，打破瓶子。他们左手拿着火把，右手拿着吹的角，喊叫：“耶和华和 基甸 的刀！”
JUDG|7|21|他们围着军营，各人站在自己的地方；全营的人都逃窜，一面喊，一面逃跑。
JUDG|7|22|三百人就吹角，耶和华使全营的人用刀自相击杀。全营的人逃往 西利拉 的 伯．哈示他 ，一直逃到靠近 他巴 的 亚伯．米何拉 。
JUDG|7|23|从 拿弗他利 、 亚设 和 玛拿西 全地来的 以色列 人被召来，追赶 米甸 人。
JUDG|7|24|基甸 也派人走遍 以法莲 山区，说：“你们下来迎击 米甸 人，在他们的前面沿着 约旦河 把守渡口，直到 伯．巴拉 。”于是 以法莲 众人聚集，沿着 约旦河 把守渡口，直到 伯．巴拉 。
JUDG|7|25|他们捉住了 米甸 的两个领袖， 俄立 和 西伊伯 。他们在 俄立 磐石上杀了 俄立 ，在 西伊伯 酒池那里杀了 西伊伯 。他们追赶 米甸 人，把 俄立 和 西伊伯 的首级带到 约旦河 对岸，到 基甸 那里。
JUDG|8|1|以法莲 人对 基甸 说：“你去与 米甸 争战，没有召我们同去，你为什么这样待我们呢？”他们就和 基甸 激烈地争吵。
JUDG|8|2|基甸 对他们说：“我现在所做的怎么与你们所做的相比呢？ 以法莲 拾取剩下的葡萄不强过 亚比以谢 族所摘的葡萄吗？
JUDG|8|3|上帝已把 米甸 的两个领袖 俄立 和 西伊伯 交在你们手中；我所做的怎能与你们所做的相比呢？” 基甸 说了这话，他们对他的怒气就消了。
JUDG|8|4|基甸 和跟随他的三百人来到 约旦河 ，渡了过去；他们虽然疲乏，还是追赶。
JUDG|8|5|基甸 对 疏割 人说：“请你们拿几块饼来给跟随我的百姓，因为他们疲乏了。我正在追击 米甸 王 西巴 和 撒慕拿 。”
JUDG|8|6|疏割 人的领袖回答说：“ 西巴 和 撒慕拿 的手掌现在已经在你手里，因此我们该将饼送给你的军队吗？”
JUDG|8|7|基甸 说：“好吧！耶和华将 西巴 和 撒慕拿 交在我手之后，我必用旷野的荆棘和枳条鞭打你们。”
JUDG|8|8|基甸 从那里上到 毗努伊勒 ，对那里的人也提出同样的请求； 毗努伊勒 人给他的答覆跟 疏割 人的答覆一样。
JUDG|8|9|他也对 毗努伊勒 人说：“我平平安安回来的时候，必拆毁这城楼。”
JUDG|8|10|那时 西巴 和 撒慕拿 ，以及跟随他们的军队都在 加各 ，约有一万五千人，是东边的人全军所剩下的，因为拿刀战死的约有十二万人。
JUDG|8|11|基甸 从 挪巴 和 约比哈 的东边，从住帐棚人 的路上去，趁 米甸 的军兵以为安全的时候攻击他们。
JUDG|8|12|西巴 和 撒慕拿 逃跑； 基甸 追赶他们，捉住 米甸 的两个王 西巴 和 撒慕拿 ，使他们全军溃散。
JUDG|8|13|约阿施 的儿子 基甸 从战场，沿着 希列斯 斜坡回来，
JUDG|8|14|捉住 疏割 人的一个少年，查问他。他就为 基甸 写下 疏割 的领袖和长老的名字，共七十七人。
JUDG|8|15|基甸 到了 疏割 人那里，说：“你们从前讥笑我说：‘ 西巴 和 撒慕拿 的手掌现在已经在你手里，因此我们该将饼送给跟随你的疲乏的人吗？’看哪， 西巴 和 撒慕拿 在这里。”
JUDG|8|16|于是他拿住城内的长老，用旷野的荆棘和枳条责打 疏割 人。
JUDG|8|17|他又拆了 毗努伊勒 的城楼，杀了城里的人。
JUDG|8|18|基甸 对 西巴 和 撒慕拿 说：“你们在 他泊山 所杀的人是什么样子的？”他们说：“他们很像你，个个都有王子的样子。”
JUDG|8|19|基甸 说：“他们都是我的兄弟，我母亲的儿子。我指着永生的耶和华起誓，你们若存留他们的性命，我就不杀你们了。”
JUDG|8|20|他对他的长子 益帖 说：“你起来杀他们！”但是这少年害怕，不敢拔刀，因为他还是个少年。
JUDG|8|21|西巴 和 撒慕拿 说：“你自己起来杀我们吧！因为人如何，力量也如何。” 基甸 就起来，杀了 西巴 和 撒慕拿 ，取了他们骆驼颈项上的月牙圈。
JUDG|8|22|以色列 人对 基甸 说：“你既然救我们脱离 米甸 的手，愿你治理我们，你的儿子孙子也治理我们。”
JUDG|8|23|基甸 对他们说：“我不治理你们，我的儿子也不治理你们，耶和华会治理你们。”
JUDG|8|24|基甸 又对他们说：“我有一件事求你们，请你们各人把所夺的耳环给我。”因敌人都戴金耳环，他们是 以实玛利 人。
JUDG|8|25|以色列 人说：“我们情愿送给你！”他们就铺开一件外衣，各人将所夺的耳环丢在上面。
JUDG|8|26|基甸 所要求的金耳环，重一千七百舍客勒金子。此外还有 米甸 王所戴的月牙圈、耳环，和所穿的紫色衣服，以及骆驼颈项上的链子。
JUDG|8|27|基甸 以此造了一个以弗得，设立在他的本城 俄弗拉 。全 以色列 就在那里拜这以弗得行淫，这就成了 基甸 和他全家的圈套。
JUDG|8|28|这样， 米甸 就被 以色列 人制伏了，再也不能抬头。 基甸 还在的日子，这地太平四十年。
JUDG|8|29|约阿施 的儿子 耶路巴力 回去，住在自己家里。
JUDG|8|30|基甸 有七十个亲生的儿子，因为他有许多妻子。
JUDG|8|31|他在 示剑 的妾也为他生了一个儿子， 基甸 给他起名叫 亚比米勒 。
JUDG|8|32|约阿施 的儿子 基甸 年纪老迈而死，葬在 亚比以谢 族的 俄弗拉 ，他父亲 约阿施 的坟墓里。
JUDG|8|33|基甸 死后， 以色列 人又去随从诸 巴力 而行淫，以 巴力．比利土 为他们的神明。
JUDG|8|34|以色列 人不记得耶和华－他们的上帝，就是那位拯救他们脱离四围仇敌之手的，
JUDG|8|35|也不照着 耶路巴力 ，就是 基甸 向 以色列 所施的恩惠善待他的家。
JUDG|9|1|耶路巴力 的儿子 亚比米勒 到 示剑 他的母舅那里，对他们和他外祖父全家的人说：
JUDG|9|2|“请你们问 示剑 所有的居民：‘是 耶路巴力 的众儿子七十人都治理你们好，还是一人治理你们好呢？’你们要记得，我是你们的骨肉。”
JUDG|9|3|他的母舅们为他把这一切话说给 示剑 所有的居民听，他们的心就倾向 亚比米勒 ，因为他们说：“他是我们的弟兄。”
JUDG|9|4|他们从 巴力．比利土 的庙中取了七十银子给 亚比米勒 ， 亚比米勒 用这些钱雇了一些无赖匪徒跟随他。
JUDG|9|5|他来到 俄弗拉 他父亲的家，在一块磐石上把他的兄弟，就是 耶路巴力 的七十个儿子都杀了，只剩下 耶路巴力 的小儿子 约坦 ，因为他躲了起来。
JUDG|9|6|示剑 所有的居民和全 伯．米罗 都聚集在一起，到 示剑 橡树旁的柱子那里，立 亚比米勒 为王。
JUDG|9|7|有人将这事告诉 约坦 ，他就去站在 基利心山 顶上，高声喊叫，对他们说：“ 示剑 的居民哪，你们要听我，上帝也就会听你们。
JUDG|9|8|有一次，树木要膏一王治理他们，就去对橄榄树说：‘请你来作王治理我们！’
JUDG|9|9|橄榄树对它们说：‘我岂可停止生产使神明和人得尊荣的油，而行走飘摇在众树之上呢？’
JUDG|9|10|树木对无花果树说：‘请你来作王治理我们！’
JUDG|9|11|无花果树对它们说：‘我岂可停止结甜美的果子，而行走飘摇在众树之上呢？’
JUDG|9|12|树木对葡萄树说：‘请你来作王治理我们！’
JUDG|9|13|葡萄树对它们说：‘我岂可停止出产使神明和人欢乐的新酒，而行走飘摇在众树之上呢。’
JUDG|9|14|众树对荆棘说：‘请你来作王治理我们！’
JUDG|9|15|荆棘对众树说：‘你们若真的要膏我作王治理你们，就要来到我的荫下寻求庇护；不然，愿火从荆棘里出来，吞灭 黎巴嫩 的香柏树。’
JUDG|9|16|“现在你们若以诚实正直立 亚比米勒 为王，若善待 耶路巴力 和他的家，若照他手所做的回报他─
JUDG|9|17|从前我父为你们争战，冒生命的危险救你们脱离 米甸 的手，
JUDG|9|18|但是你们如今起来攻击我的父家，在一块磐石上把他的七十个儿子全杀了，又立他使女所生的儿子 亚比米勒 为 示剑 居民的王，因为他是你们的弟兄─
JUDG|9|19|你们如今若以诚实正直对待 耶路巴力 和他的家，就可以因 亚比米勒 欢乐，他也可以因你们欢乐；
JUDG|9|20|不然，愿火从 亚比米勒 发出，吞灭 示剑 居民和 伯．米罗 ，又愿火从 示剑 居民和 伯．米罗 发出，吞灭 亚比米勒 。”
JUDG|9|21|约坦 因躲避他的兄弟 亚比米勒 就逃跑，去到 比珥 ，住在那里。
JUDG|9|22|亚比米勒 治理 以色列 三年。
JUDG|9|23|上帝派邪灵到 亚比米勒 和 示剑 居民中间， 示剑 居民就以诡诈待 亚比米勒 。
JUDG|9|24|这是要使 耶路巴力 七十个儿子受害所流的血，归于他们的兄弟 亚比米勒 ，因他杀害他们，也归于那些出手帮助他杀害兄弟的 示剑 居民。
JUDG|9|25|示剑 居民在山顶上设下埋伏，等候 亚比米勒 。凡沿着那条路，从他们那里经过的人，他们就抢劫。有人把这事告诉 亚比米勒 。
JUDG|9|26|以别 的儿子 迦勒 和他的弟兄经过，来到 示剑 ， 示剑 居民都信任他。
JUDG|9|27|他们出到田间，摘下葡萄，踹酒，作乐。他们进入他们神明的庙中吃喝，诅咒 亚比米勒 。
JUDG|9|28|以别 的儿子 迦勒 说：“ 亚比米勒 是谁，我们 示剑 人是谁，叫我们服事他呢？他不是 耶路巴力 的儿子吗？他的助手不是 西布勒 吗？你们应当服事 示剑 的父亲 哈抹 的后裔！我们为何要服事 亚比米勒 呢？
JUDG|9|29|惟愿这民归到我的手下，我就除掉 亚比米勒 。”他就对 亚比米勒 说：“增加你的军兵，出来吧！”
JUDG|9|30|西布勒 市长听见 以别 的儿子 迦勒 的话，就怒气大发。
JUDG|9|31|他悄悄地派一些使者到 亚比米勒 那里，说：“看哪， 以别 的儿子 迦勒 和他的弟兄到了 示剑 。看哪，他们煽动那城攻击你。
JUDG|9|32|现在，你和跟随你的百姓要夜间起来，在田间埋伏。
JUDG|9|33|早晨太阳一出，你就趁早攻城。看哪， 迦勒 和跟随他的百姓出来攻击你的时候，你就全力对付他们。”
JUDG|9|34|于是， 亚比米勒 和跟随他的众百姓夜间起来，兵分四队，埋伏攻击 示剑 。
JUDG|9|35|以别 的儿子 迦勒 出去，站在城门口。 亚比米勒 和跟随他的百姓从埋伏之处起来。
JUDG|9|36|迦勒 看见百姓，就对 西布勒 说：“看哪，有百姓从山顶上下来。” 西布勒 对他说：“你把山的影子看作是人了。”
JUDG|9|37|迦勒 又继续讲，他说：“看哪，有百姓从地的高处下来，又有一队从 米恶尼尼 橡树 的路前来。”
JUDG|9|38|西布勒 对他说：“你所夸口的在哪里呢？你曾说：‘ 亚比米勒 是谁，叫我们服事他呢？’这不是你所藐视的百姓吗？你现在出去，与他们交战吧！”
JUDG|9|39|于是 迦勒 率领 示剑 居民出去，与 亚比米勒 交战。
JUDG|9|40|亚比米勒 追赶 迦勒 ， 迦勒 在他面前逃跑。有许多人被刺伤仆倒，直到城门口。
JUDG|9|41|亚比米勒 住在 亚鲁玛 。 西布勒 赶出 迦勒 和他的弟兄，不准他们住在 示剑 。
JUDG|9|42|次日，百姓出到田间，有人告诉 亚比米勒 ，
JUDG|9|43|他就带领百姓，把他们分成三队，埋伏在田间窥探。看哪， 示剑 居民从城里出来，他就起来击杀他们。
JUDG|9|44|亚比米勒 和跟随他的一队向前冲，站在城门口；另外两队直冲向田间，击杀了众人。
JUDG|9|45|亚比米勒 攻城一整天，将城夺取，杀了其中的百姓，把城拆毁，撒上了盐。
JUDG|9|46|示剑 城楼里所有的居民听见了，就进入 伊勒．比利土 庙的地窖里。
JUDG|9|47|有人告诉 亚比米勒 ， 示剑 城楼里所有的居民都聚在一起。
JUDG|9|48|亚比米勒 和所有跟随他的百姓都上 撒们山 去。 亚比米勒 手拿斧子，砍下一根树枝，举起来，扛在肩上，对跟随他的百姓说：“你们看我做什么，就赶快照样做。”
JUDG|9|49|众百姓也都各砍一根树枝，跟 亚比米勒 走，把树枝堆在地窖上，放火烧地窖。这样， 示剑 城楼里所有的人都死了，男女约有一千。
JUDG|9|50|亚比米勒 到 提备斯 ，对着 提备斯 安营，攻取了那城。
JUDG|9|51|城中有一座坚固的楼；城里所有的居民，无论男女，都逃到那里，关上门，上了楼顶。
JUDG|9|52|亚比米勒 到了楼前，攻打它。他挨近楼门，要放火焚烧。
JUDG|9|53|有一个妇人把一块上磨石抛在 亚比米勒 的头上，打破了他的头盖骨。
JUDG|9|54|他就急忙叫拿他兵器的青年来，对他说：“拔出你的刀来，杀了我吧！免得有人提到我说：‘他被一个妇人杀了。’”于是那青年把他刺透，他就死了。
JUDG|9|55|以色列 人见 亚比米勒 死了，就各回自己的地方去了。
JUDG|9|56|这样，上帝报应了 亚比米勒 向他父亲所做的恶事，就是杀了自己七十个兄弟。
JUDG|9|57|示剑 人的一切恶事，上帝也都报应在他们头上； 耶路巴力 的儿子 约坦 的诅咒都临到他们身上了。
JUDG|10|1|亚比米勒 以后， 陀拉 兴起，拯救 以色列 ，他是 朵多 的孙子， 普瓦 的儿子， 以萨迦 人，住在 以法莲 山区的 沙密 。
JUDG|10|2|陀拉 作 以色列 的士师二十三年。他死了，葬在 沙密 。
JUDG|10|3|陀拉 以后有 基列 人 睚珥 兴起，作 以色列 的士师二十二年。
JUDG|10|4|他有三十个儿子，骑着三十匹驴驹。他们有三十座城，叫作 哈倭特．睚珥 ，直到如今，都在 基列 地。
JUDG|10|5|睚珥 死了，葬在 加们 。
JUDG|10|6|以色列 人又行耶和华眼中看为恶的事，去事奉诸 巴力 和 亚斯她录 ，以及 亚兰 的神明、 西顿 的神明、 摩押 的神明、 亚扪 人的神明、 非利士 人的神明。他们离弃耶和华，不事奉他。
JUDG|10|7|耶和华的怒气向 以色列 发作，把他们交给 非利士 人和 亚扪 人的手中。
JUDG|10|8|从那年起，他们欺压迫害 以色列 人，在 约旦河 东， 亚摩利 人境内， 基列 一带所有的 以色列 人，长达十八年。
JUDG|10|9|亚扪 人渡过 约旦河 去攻打 犹大 和 便雅悯 ，以及 以法莲 家族。 以色列 的处境非常困苦。
JUDG|10|10|以色列 人哀求耶和华说：“我们得罪了你，因为我们离弃了我们的上帝，去事奉诸 巴力 。”
JUDG|10|11|耶和华对 以色列 人说：“我岂没有救你们脱离 埃及 人、 亚摩利 人、 亚扪 人和 非利士 人吗？
JUDG|10|12|西顿 人、 亚玛力 人和 马云 人 欺压你们，你们哀求我，我也拯救你们脱离他们的手。
JUDG|10|13|你们竟离弃我去事奉别神！所以我不再救你们了。
JUDG|10|14|你们去哀求你们所选择的神明；你们遭遇急难的时候，让它们救你们吧！”
JUDG|10|15|以色列 人对耶和华说：“我们犯罪了，照你看为好的待我们，只求你今日拯救我们吧！”
JUDG|10|16|以色列 人就除掉他们中间的外邦神明，事奉耶和华。耶和华因 以色列 所受的苦难而心里焦急。
JUDG|10|17|亚扪 人被召来，在 基列 安营； 以色列 人也聚集，在 米斯巴 安营。
JUDG|10|18|基列 百姓中的领袖彼此说：“谁领先出去攻打 亚扪 人，谁就作 基列 所有居民的领袖。”
JUDG|11|1|基列 人 耶弗他 是个大能的勇士，是妓女的儿子。 基列 生了 耶弗他 。
JUDG|11|2|基列 的妻子也给他生了几个儿子。他妻子生的儿子长大后，就把 耶弗他 赶出去，说：“你不可在我们父家继承产业，因为你是别的女人生的儿子。”
JUDG|11|3|耶弗他 就逃离他的兄弟，住在 陀伯 地。有些无赖的人聚集在他那里，与他一同出入。
JUDG|11|4|过了些日子， 亚扪 人攻打 以色列 。
JUDG|11|5|亚扪 人攻打 以色列 的时候， 基列 的长老去请 耶弗他 从 陀伯 地回来。
JUDG|11|6|他们对 耶弗他 说：“请你来作我们的指挥官，好让我们跟 亚扪 人打仗。”
JUDG|11|7|耶弗他 对 基列 的长老说：“你们不是恨我，把我赶出父家吗？现在你们遭遇急难，为何到我这里来呢？”
JUDG|11|8|基列 的长老对 耶弗他 说：“现在我们回到你这里，是要请你同我们去跟 亚扪 人打仗，作 基列 所有居民的领袖。”
JUDG|11|9|耶弗他 对 基列 的长老说：“若你们请我回去跟 亚扪 人打仗，耶和华把他们交给我，我就作你们的领袖。”
JUDG|11|10|基列 的长老对 耶弗他 说：“有耶和华在你我之间作证，我们必定照你的话做。”
JUDG|11|11|于是 耶弗他 与 基列 的长老同去，百姓就立 耶弗他 作他们的领袖和指挥官。 耶弗他 在 米斯巴 将他一切的事陈述在耶和华面前。
JUDG|11|12|耶弗他 派使者到 亚扪 人的王那里，说：“你与我有什么相干，竟来到我这里攻打我的地呢？”
JUDG|11|13|亚扪 人的王对 耶弗他 的使者说：“因为 以色列 从 埃及 上来的时候占据我的地，从 亚嫩河 到 雅博河 ，直到 约旦河 。现在你要和平归还这些地方！”
JUDG|11|14|耶弗他 又派使者到 亚扪 人的王那里，
JUDG|11|15|对他说：“ 耶弗他 如此说： 以色列 并没有占据 摩押 地和 亚扪 人的地。
JUDG|11|16|以色列 人从 埃及 上来，是经过旷野到 红海 ，来到 加低斯 。
JUDG|11|17|那时， 以色列 派使者去 以东 王那里，说：‘求你让我穿越你的地。’ 以东 王却不听。 以色列 又照样派使者去 摩押 王那里，他也不肯。于是 以色列 人就住在 加低斯 。
JUDG|11|18|他们又经过旷野，绕过 以东 地和 摩押 地，到 摩押 地的东边 ，在 亚嫩河 边安营，并没有进入 摩押 的境内，因为 亚嫩河 是 摩押 的边界。
JUDG|11|19|以色列 派使者去 亚摩利 王，就是 希实本 王 西宏 那里； 以色列 对他说：‘求你让我们穿越你的地，到我自己的地方去。’
JUDG|11|20|西宏 却不信任 以色列 ，不让他们穿越他的疆界。他召集了他的众百姓在 雅杂 安营，与 以色列 争战。
JUDG|11|21|耶和华－ 以色列 的上帝将 西宏 和他的众百姓都交在 以色列 手中， 以色列 人就击杀他们，占领了那地居民 亚摩利 人的全地。
JUDG|11|22|他们占领了 亚摩利 人所有的疆土，从 亚嫩河 到 雅博河 ，从旷野直到 约旦河 。
JUDG|11|23|耶和华－ 以色列 的上帝如今从他百姓 以色列 面前赶出 亚摩利 人，你竟要占领它吗？
JUDG|11|24|你不是已经得了你的神明 基抹 赐给你的地为业吗？耶和华－我们的上帝在我们面前所赶出的，我们也要得它为业。
JUDG|11|25|现在你比 西拨 的儿子 摩押 王 巴勒 还强吗？他真的曾与 以色列 争执，或是真的与他们争战了吗？
JUDG|11|26|以色列 人住 希实本 和所属的乡镇， 亚罗珥 和所属的乡镇，以及沿着 亚嫩河 的一切城镇，已经有三百年了。在这期间，你们为什么不取回呢？
JUDG|11|27|我并没有得罪你，你却要攻打我，加害于我。愿审判人的耶和华今日在 以色列 人和 亚扪 人之间判断是非。”
JUDG|11|28|但 亚扪 人的王不听 耶弗他 传达给他的话。
JUDG|11|29|耶和华的灵降在 耶弗他 身上，他就经过 基列 和 玛拿西 ，经过 基列 的 米斯巴 ，又从 基列 的 米斯巴 过到 亚扪 人那里。
JUDG|11|30|耶弗他 向耶和华许愿，说：“你若真的将 亚扪 人交在我手中，
JUDG|11|31|我从 亚扪 人那里平平安安回来的时候，无论谁先从我家门出来迎接我，就要归给耶和华，我必将他献上作为燔祭。”
JUDG|11|32|于是 耶弗他 往 亚扪 人那里去，与他们争战。耶和华将他们交在他手中，
JUDG|11|33|他就彻底击败他们，从 亚罗珥 到 米匿 ，直到 亚备勒．基拉明 ，攻取了二十座城。这样， 亚扪 人就在 以色列 人面前被制伏了。
JUDG|11|34|耶弗他 回 米斯巴 去，到了自己的家，看哪，他女儿拿着手鼓跳舞出来迎接他。她是 耶弗他 的独生女，除她以外，没有别的儿女。
JUDG|11|35|耶弗他一看见她，就撕裂衣服，说：“哀哉！我的女儿啊，你使我非常悲痛，叫我十分为难了。因为我已经向耶和华开了口，不能收回。”
JUDG|11|36|他女儿对他说：“我的父亲啊，你既向耶和华开了口，就当照你口中所说的向我行，因为耶和华已经在你的仇敌 亚扪 人身上为你报了仇。”
JUDG|11|37|她又对父亲说：“我只求你这一件事，给我两个月，让我和同伴下到山里，好为我的童贞哀哭。”
JUDG|11|38|耶弗他 说：“你去吧！”他就让她离开两个月。她和同伴去了，在山里为她的童贞哀哭。
JUDG|11|39|过了两个月，她回到父亲那里，父亲就照所许的愿向她行了。她从来没有亲近男人。于是 以色列 中有个风俗，
JUDG|11|40|每年按着日期 以色列 的女子要去为 基列 人 耶弗他 的女儿哀哭四天。
JUDG|12|1|以法莲 人被召来，渡河来到 撒分 。他们对 耶弗他 说：“你去与 亚扪 人争战，为什么没有召我们同去呢？我们必用火将你和你的家烧了。”
JUDG|12|2|耶弗他 对他们说：“我和我的百姓与 亚扪 人有极大的冲突；我曾召你们来，你们却没有来救我脱离他们的手。
JUDG|12|3|我见你们不来救我，就拚了命前去攻打 亚扪 人，耶和华就将他们交在我手中。你们今日为什么上我这里来攻打我呢？”
JUDG|12|4|于是 耶弗他 召集 基列 所有的人，要与 以法莲 人争战。 基列 人击杀 以法莲 人，因 以法莲 人曾说：“你们 基列 人在 以法莲 和 玛拿西 中，不过是 以法莲 逃亡的人而已。”
JUDG|12|5|基列 人把守 约旦河 的渡口，不许 以法莲 人过去。逃跑的 以法莲 人若说：“让我过河。” 基列 人就问他说：“你是不是 以法莲 人？”他若说：“不是”，
JUDG|12|6|基列 人就对他说：“你说‘示播列’。” 以法莲 人因为发音不准，就会说成“西播列”。 基列 人就捉住他，在 约旦河 的渡口把他杀了。那时， 以法莲 人被杀的有四万二千人。
JUDG|12|7|耶弗他 作 以色列 的士师六年。 基列 人 耶弗他 死了，葬在 基列 的城里 。
JUDG|12|8|耶弗他 以后，有 伯利恒 人 以比赞 作 以色列 的士师。
JUDG|12|9|他有三十个儿子。他把三十个女儿都嫁出去了，也为他的儿子从外面娶了三十个媳妇。他作 以色列 的士师七年。
JUDG|12|10|以比赞 死了，葬在 伯利恒 。
JUDG|12|11|以比赞 以后，有 西布伦 人 以伦 作 以色列 的士师，他作 以色列 的士师十年。
JUDG|12|12|西布伦 人 以伦 死了，葬在 西布伦 地的 亚雅仑 。
JUDG|12|13|以伦 以后，有 比拉顿 人 希列 的儿子 押顿 作 以色列 的士师。
JUDG|12|14|他有四十个儿子，三十个孙子，骑着七十匹驴驹。 押顿 作 以色列 的士师八年。
JUDG|12|15|比拉顿 人 希列 的儿子 押顿 死了，葬在 以法莲 地的 比拉顿 ，就在 亚玛力 人的山区。
JUDG|13|1|以色列 人又行耶和华眼中看为恶的事，耶和华将他们交在 非利士 人手中四十年。
JUDG|13|2|那时，有一个 但 支派的 琐拉 人，名叫 玛挪亚 。他的妻子不怀孕，不生育。
JUDG|13|3|耶和华的使者向那妇人显现，对她说：“看哪，以前你不怀孕，不生育，如今你必怀孕生一个儿子。
JUDG|13|4|现在你要谨慎，清酒烈酒都不可喝，任何不洁之物都不可吃，
JUDG|13|5|看哪，你必怀孕，生一个儿子。不可用剃刀剃他的头，因为这孩子一出母胎就归给上帝作拿细耳人。他必开始拯救 以色列 脱离 非利士 人的手。”
JUDG|13|6|那妇人来对丈夫说：“有一个神人到我这里来，他的容貌如上帝使者的容貌，非常可畏。我没有问他从哪里来，他也没有把他的名字告诉我。
JUDG|13|7|他对我说：‘看哪，你要怀孕，生一个儿子 。现在，清酒烈酒都不可喝，任何不洁之物都不可吃，因为这孩子从出母胎一直到死的那一天，要归给上帝作拿细耳人。’”
JUDG|13|8|玛挪亚 祈求耶和华说：“主啊，求你再差遣那神人到我们这里来，指示我们对这将要生的孩子该怎样作。”
JUDG|13|9|上帝垂听了 玛挪亚 的声音。那妇人坐在田间的时候，上帝的使者又到她那里，但是她的丈夫 玛挪亚 没有同她在一起。
JUDG|13|10|妇人急忙跑去告诉丈夫，对他说：“看哪，那日到我这里来的人又向我显现了。”
JUDG|13|11|玛挪亚 起来，跟随他的妻子来到那人那里，对他说：“你就是跟这妇人说话的那个人吗？”他说：“是我。”
JUDG|13|12|玛挪亚 说：“现在，愿你的话应验！这孩子该如何管教呢？他当做什么呢？”
JUDG|13|13|耶和华的使者对 玛挪亚 说：“我告诉这妇人的一切事，她都要遵守。
JUDG|13|14|葡萄树所结的不可吃，清酒烈酒都不可喝，任何不洁之物也不可吃。凡我所吩咐的，她都当遵守。”
JUDG|13|15|玛挪亚 对耶和华的使者说：“请容许我们留你下来，好为你预备一只小山羊。”
JUDG|13|16|耶和华的使者对 玛挪亚 说：“你虽然留我，我却不吃你的食物。你若预备燔祭，就当献给耶和华。”因 玛挪亚 不知道他是耶和华的使者。
JUDG|13|17|玛挪亚 对耶和华的使者说：“请问大名？好让我们在你的话应验的时候尊敬你。”
JUDG|13|18|耶和华的使者对他说：“你何必问我的名字呢？我的名字是奇妙的。”
JUDG|13|19|玛挪亚 取一只小山羊和素祭，在磐石上献给耶和华。他行奇妙的事， 玛挪亚 和他的妻子观看，
JUDG|13|20|火焰从坛上往上升，耶和华的使者也在坛上的火焰中升上去了。 玛挪亚 和他的妻子看见，就脸伏于地。
JUDG|13|21|耶和华的使者不再向 玛挪亚 和他的妻子显现了。那时， 玛挪亚 才知道他是耶和华的使者。
JUDG|13|22|玛挪亚 对他的妻子说：“我们一定会死，因为我们看见了上帝。”
JUDG|13|23|他的妻子却对他说：“耶和华若有意要我们死，就不会从我们手中接受燔祭和素祭，不会将这一切事指示我们，这时也不会让我们听到这话。”
JUDG|13|24|后来妇人生了一个儿子，给他起名叫 参孙 。孩子渐渐长大，耶和华赐福给他。
JUDG|13|25|在 琐拉 和 以实陶 之间的 玛哈尼．但 ，耶和华的灵开始感动 参孙 。
JUDG|14|1|参孙 下到 亭拿 ，在 亭拿 看见一个女子，是 非利士 人的女儿。
JUDG|14|2|他上来告诉他父母说：“我在 亭拿 看见一个女子，是 非利士 人的女儿，现在请你们给我娶她为妻。”
JUDG|14|3|他父母对他说：“在你弟兄的女儿中，或在本族所有的人中，难道没有女子吗？你何必在未受割礼的 非利士 人中去娶妻呢？” 参孙 对他父亲说：“请你给我娶那女子，因为我喜欢她。”
JUDG|14|4|他的父母并不知道这事是出于耶和华，因为他在找机会攻击 非利士 人。那时， 非利士 人辖制 以色列 人。
JUDG|14|5|参孙 跟他父母下 亭拿 去，他们到了 亭拿 的葡萄园。看哪，有一只少壮狮子对着他吼叫。
JUDG|14|6|耶和华的灵大大感动 参孙 ，他就手无寸铁撕裂狮子，如撕裂小山羊一样。他做这事，并没有告诉他的父母亲。
JUDG|14|7|参孙 下去跟那女子说话，看着就喜欢她。
JUDG|14|8|过了些日子，他回来要娶那女子，绕道去看狮子的残骸，看哪，有一群蜜蜂在狮子的尸体内，也有蜜在里面。
JUDG|14|9|他就取了蜜，放在手掌上，边走边吃。他到了父母那里，给他们蜜，他们也吃了。但他没有告诉他们，这蜜是从狮子的尸体内取来的。
JUDG|14|10|他父亲下到女子那里去。 参孙 在那里摆设宴席， 因为这是当时年轻人的习俗。
JUDG|14|11|他们看见 参孙 ，就请了三十个人陪伴他。
JUDG|14|12|参孙 对他们说：“我给你们出个谜语，你们若能在七日宴席之内，猜出谜底告诉我，我就给你们三十件细麻内衣和三十套更换的衣服。
JUDG|14|13|但你们若不能告诉我，你们就给我三十件细麻内衣和三十套更换的衣服。”他们对他说：“请把谜语说给我们听。”
JUDG|14|14|参孙 对他们说： “吃的从吃者出来； 甜的从强者出来”。 三日之久，他们都猜不出谜语来。
JUDG|14|15|第七日 ，他们对 参孙 的妻子说：“你哄骗你的丈夫，为我们探出谜底来，否则我们就用火烧你和你的父家。你们请我们来，是不是要夺走我们所有的呢？”
JUDG|14|16|参孙 的妻子在丈夫面前哭哭啼啼说：“你只是恨我，并不爱我。你给我本族的人出谜语，却不把谜底告诉我。” 参孙 对她说：“看哪，连我的父母我都没有说，我怎么可以告诉你呢？”
JUDG|14|17|在七日宴席中，她一直在丈夫面前哭哭啼啼。第七日， 参孙 因妻子的催逼就把谜底告诉了她。她把谜底告诉了她本族的人。
JUDG|14|18|第七日日落以前，那城里的人对 参孙 说： “有什么比蜜还甜呢？ 有什么比狮子更强呢？” 参孙 对他们说： “你们若不用我的母牛犊耕地， 就无法猜出我的谜底来。”
JUDG|14|19|耶和华的灵大大感动 参孙 ，他就下到 亚实基伦 ，击杀了三十个人，夺了他们身上的衣服，把衣服给了猜出谜语的人。 参孙 怒气大发，就上他父亲的家去了。
JUDG|14|20|参孙 的妻子就归了 参孙 的一个同伴，就是作过他伴郎的。
JUDG|15|1|过了些日子，在割麦子的时候， 参孙 带着一只小山羊去探望他的妻子，说：“我要进内室到我妻子那里。”他岳父不许他进去。
JUDG|15|2|他岳父说：“我以为你极其恨她，因此我把她给了你的同伴。她妹妹不是比她更美丽吗？你可以娶来代替她！”
JUDG|15|3|参孙 对他们说：“这一次我若加害 非利士 人，就不算是我的错了。”
JUDG|15|4|于是 参孙 去捉了三百只狐狸，把它们的尾巴一对一对地绑住，再将火把绑在两条尾巴中间。
JUDG|15|5|他点着火把，把狐狸放进 非利士 人直立的庄稼，把堆积的禾捆和直立的庄稼，葡萄园、橄榄园全都烧了。
JUDG|15|6|非利士 人说：“这事是谁做的呢？”有人说：“是 亭拿 人的女婿 参孙 做的，因为他岳父把他的妻子给了他的同伴。”于是 非利士 人上去，用火烧了女子和她的父亲。
JUDG|15|7|参孙 对他们说：“你们既然这么做，我必向你们报仇才肯罢休。”
JUDG|15|8|参孙 狠狠击杀他们，把他们连腿带腰都砍了。过后，他就下去，住在 以坦岩 的石洞里。
JUDG|15|9|非利士 人上去，安营在 犹大 ，侵犯 利希 。
JUDG|15|10|犹大 人说：“你们为何上来攻击我们呢？”他们说：“我们上来是要捆绑 参孙 ，照他向我们所做的对待他。”
JUDG|15|11|于是，三千 犹大 人下到 以坦岩 的石洞里，对 参孙 说：“ 非利士 人辖制我们，你不知道吗？你向我们做的是什么事呢？”他说：“他们向我怎样做，我也要向他们怎样做。”
JUDG|15|12|犹大 人对他说：“我们下来是要捆绑你，把你交在 非利士 人手中。” 参孙 说：“你们要向我起誓，你们自己不杀害我。”
JUDG|15|13|他们说：“我们绝不杀你，只把你捆绑，交在 非利士 人手中。”于是他们用两条新绳绑住 参孙 ，把他从 以坦岩 带上去。
JUDG|15|14|参孙 到了 利希 ， 非利士 人对着他喊叫。耶和华的灵大大感动 参孙 ，他手臂上的绳子就像着火的麻一样，绑他的绳子从他手上脱落下来。
JUDG|15|15|他找到一块未干的驴腮骨，就伸手拾起来，用它杀了一千人。
JUDG|15|16|参孙 说： “用驴腮骨， 一堆又一堆 ； 用驴腮骨， 我杀了一千人。”
JUDG|15|17|说完这话，就把那腮骨从手里抛出去。因此，那地叫作 拉末．利希 。
JUDG|15|18|参孙 非常口渴，就求告耶和华说：“你既藉仆人的手施行这么大的拯救，现在我要渴死，落在未受割礼的人手中吗？”
JUDG|15|19|上帝就使 利希 的洼地裂开，从中涌出水来。 参孙 喝了，精神恢复。因此那泉名叫 隐．哈歌利 ，直到今日它仍在 利希 。
JUDG|15|20|在 非利士 人辖制的时候， 参孙 作 以色列 的士师二十年。
JUDG|16|1|参孙 到了 迦萨 ，在那里看见一个妓女，就与她亲近。
JUDG|16|2|有人告诉 迦萨 人说：“ 参孙 到这里来了！”他们就包围起来，整夜在城门埋伏等着他。他们整夜静悄悄地，说：“等到天一亮我们就杀他。”
JUDG|16|3|参孙 睡到半夜，在半夜起来，抓住城门的门扇和两个门框，把它们和门闩一起拆下来，扛在肩上，抬到 希伯仑 前面的山顶上。
JUDG|16|4|这事以后， 参孙 在 梭烈谷 爱上了一个女子，名叫 大利拉 。
JUDG|16|5|非利士 人的领袖上去，到那女子那里，对她说：“请你哄骗 参孙 ，探出他为何有这么大的力气，以及我们要用什么方法才能胜他，将他捆绑制伏。我们就每人给你一千一百块银子。”
JUDG|16|6|大利拉 对 参孙 说：“请你告诉我，你为何有这么大的力气，要用什么方法才能捆绑制伏你。”
JUDG|16|7|参孙 对她说：“若用七条未干的新绳子捆绑我，我就像平常人一样软弱。”
JUDG|16|8|于是 非利士 人的领袖拿了七条未干的新绳子来，交给她，她就用绳子捆绑 参孙 。
JUDG|16|9|当时，埋伏的人正在她的内室等着。她对 参孙 说：“ 参孙 ， 非利士 人来捉你了！” 参孙 就挣断绳子，绳子如遇到火的麻线断裂一样。这样，人还是不知道他的力量从哪里来。
JUDG|16|10|大利拉 对 参孙 说：“看哪，你欺骗我，对我说谎。现在请你告诉我，要用什么方法才能捆绑你。”
JUDG|16|11|参孙 对她说：“若用未曾用过的新绳子捆绑我，我就像平常人一样软弱。”
JUDG|16|12|大利拉 就用新绳子捆绑他，对他说：“ 参孙 ， 非利士 人来捉你了！”当时，埋伏的人在内室等着。 参孙 挣断手臂上的绳子，如挣断一条线一样。
JUDG|16|13|大利拉 对 参孙 说：“你到现在还是欺骗我，对我说谎。请你告诉我，要用什么方法才能捆绑你。” 参孙 对她说：“只要用织布的线将我头上的七条发绺编织起来就可以了”。
JUDG|16|14|于是 大利拉 用梭子将他的发绺钉住，对他说：“ 参孙 ， 非利士 人来捉你了！” 参孙 从睡中醒来，将织布机上的梭子和织布的线一齐都拔出来了。
JUDG|16|15|大利拉 对 参孙 说：“你既不与我同心，怎么能说‘我爱你’呢？你这三次欺骗我，不告诉我，你为什么有这么大的力气。”
JUDG|16|16|大利拉 天天用话催逼他，纠缠他，他就心里烦得要死，
JUDG|16|17|终于把心中的一切都告诉她。 参孙 对她说：“从来没有人用剃刀剃我的头，因为我一出母胎就归给上帝作拿细耳人。若有人剃了我的头发，我的力气就会离开我，我就像平常人一样软弱。”
JUDG|16|18|大利拉 见他说出了心中的一切，就派人去召 非利士 人的领袖，说：“请再上来一次，因为他已经说出了心中的一切。”于是 非利士 人的领袖手里拿着银子，上到她那里。
JUDG|16|19|大利拉 哄 参孙 睡在她的膝上，叫一个人来剃掉 参孙 头上的七条发绺。于是 大利拉 开始制伏 参孙 ，他的力气就离开他了。
JUDG|16|20|大利拉 说：“ 参孙 ， 非利士 人来捉你了！” 参孙 从睡中醒来，说：“我要像前几次一样脱身而去。”他却不知道耶和华已经离开他了。
JUDG|16|21|非利士 人逮住他，挖了他的眼睛，带他下到 迦萨 ，用铜链锁住他，叫他在监狱里推磨。
JUDG|16|22|然而他的头发被剃以后，又开始长起来了。
JUDG|16|23|非利士 人的领袖聚集，要向他们的神明 大衮 献大祭，并且庆祝，说：“我们的神明把我们的仇敌 参孙 交在我们手中了。”
JUDG|16|24|众人看见 参孙 ，就赞美他们的神明说：“我们的神明把那毁坏我们的地、杀害我们许多人的仇敌交在我们手中了。”
JUDG|16|25|他们心里高兴的时候，就说：“叫 参孙 来，逗我们欢乐。”于是他们把 参孙 从监狱里提出来，在他们面前戏耍。他们叫他站在两根柱子中间。
JUDG|16|26|参孙 对牵他手的童仆说：“让我摸摸支撑这庙宇的柱子，我要靠一靠。”
JUDG|16|27|那时庙宇内充满男女， 非利士 人的众领袖也都在那里，屋顶上约有三千男女观看 参孙 逗他们欢乐。
JUDG|16|28|参孙 求告耶和华说：“主耶和华啊，求你眷念我。上帝啊，就这一次，求你赐给我力量，使我向 非利士 人报那挖我双眼的仇。”
JUDG|16|29|参孙 抱住中间支撑庙宇的两根柱子，左手抱一根，右手抱一根。
JUDG|16|30|然后他说：“让我与 非利士 人一起死吧！”他尽力弯腰，庙宇就倒塌了，压住领袖和庙宇内的众人。这样， 参孙 死的时候所杀的人比活着所杀的还多。
JUDG|16|31|他的兄弟和他父亲的全家都下去收他的尸首，抬上去，葬在 琐拉 和 以实陶 中间、他父亲 玛挪亚 的坟墓里。 参孙 作 以色列 的士师二十年。
JUDG|17|1|以法莲 山区有一个人，名叫 米迦 。
JUDG|17|2|他对母亲说：“你的一千一百块银子被人拿走了，为此你发咒起誓，也说给我听。看哪，银子在我这里，是我拿的。”他母亲说：“愿我儿蒙耶和华赐福！”
JUDG|17|3|米迦 把这一千一百块银子还他母亲。他母亲说：“我把这银子分别为圣，亲手献给耶和华，为我儿子造一尊雕刻的像，以及一尊铸成的像。现在我把银子交给你。”
JUDG|17|4|米迦 把银子还他母亲，他母亲把二百块银子交给银匠，去造一尊雕刻的像，以及一尊铸成的像，安置在 米迦 的房子里。
JUDG|17|5|米迦 这个人有了神堂，又造了以弗得和家中的神像，派他的一个儿子作祭司。
JUDG|17|6|那时， 以色列 中没有王，各人照自己眼中看为对的去做。
JUDG|17|7|犹大 的 伯利恒 有一个年轻人，是 犹大 族的人。他是 利未 人，寄居在那里。
JUDG|17|8|这人离开 犹大 的 伯利恒城 ，要找一个可住的地方。他来到 以法莲 山区 米迦 的家，还要往前走。
JUDG|17|9|米迦 对他说：“你从哪里来？”他说：“我从 犹大 的 伯利恒 来。我是 利未 人，要找一个可住的地方。”
JUDG|17|10|米迦 说：“你就住在我这里吧！我以你为父为祭司，每年给你十块银子和一套衣服，以及生活所需的食物。” 利未 人就来了。
JUDG|17|11|利未 人愿意和这人同住；他待这年轻人如自己的儿子一样。
JUDG|17|12|米迦 授这年轻的 利未 人祭司的职任，他就住在 米迦 的家里。
JUDG|17|13|米迦 说：“现在我知道耶和华必恩待我，因为我有 利未 人作我的祭司。”
JUDG|18|1|那时， 以色列 中没有王。 但 支派的人还在觅地居住，因为直到那日，他们还没有在 以色列 支派中抽签得地为业。
JUDG|18|2|但 人从 琐拉 和 以实陶 派本族中的五个勇士，去窥探侦察那地，对他们说：“你们去侦察那地。”他们来到 以法莲 山区 米迦 的家中，就在那里住宿。
JUDG|18|3|他们临近 米迦 的家，听出那年轻的 利未 人的口音，就绕到那里，对他说：“谁领你到这里来？你在这里做什么？你在这里得了什么？”
JUDG|18|4|他对他们说：“ 米迦 如此如此待我，他雇用我，我就作了他的祭司。”
JUDG|18|5|他们对他说：“请你求问上帝，使我们知道所走的道路是否通达。”
JUDG|18|6|祭司对他们说：“你们平平安安去吧，你们所行的道路是在耶和华面前的。”
JUDG|18|7|五人就走了，来到 拉亿 ，见那里的人安居，像 西顿 人的生活一样安宁无虑，那地无人羞辱他们，无人夺取侵略。他们离 西顿 人很远，与世无争 。
JUDG|18|8|五人回到 琐拉 和 以实陶 他们的弟兄那里。他们的弟兄对他们说：“你们怎么了？”
JUDG|18|9|他们说：“起来，我们上去攻打他们吧！我们已经窥探了那地，看哪，那地非常好。你们还要待在这里吗？不要再迟延了，立刻出发去得那地为业吧！
JUDG|18|10|你们去，必来到安居的百姓和两边辽阔的地。上帝已将那地方交在你们手中了；那里不缺地上的任何东西。”
JUDG|18|11|于是 但 族的六百人，各带兵器，从 琐拉 和 以实陶 出发，
JUDG|18|12|上到 犹大 的 基列．耶琳 ，在那里安营。因此那地方名叫 玛哈尼．但 ，直到今日。看哪，它在 基列．耶琳 的西边。
JUDG|18|13|他们从那里往 以法莲 山区去，来到 米迦 的家。
JUDG|18|14|先前窥探 拉亿 地的五个人对他们的弟兄说：“你们知道吗？这些屋子里有以弗得和家中的神像，以及一尊雕刻的像与一尊铸成的像。现在你们要知道该怎么做。”
JUDG|18|15|五人转身，进入 米迦 的家，来到那年轻 利未 人的房间，向他问安。
JUDG|18|16|六百 但 人各带兵器，站在门口。
JUDG|18|17|那窥探这地的五个人上前去，进入里面，拿走雕刻的像、以弗得、家中的神像，以及铸成的像。祭司和带兵器的六百人一同站在门口。
JUDG|18|18|当五个人进入 米迦 的家，拿走雕刻的像、以弗得、家中的神像，以及铸成的像，祭司对他们说：“你们做什么呢？”
JUDG|18|19|他们对他说：“不要作声，用手捂口，跟我们去吧！我们必以你为父为祭司。你作一家的祭司好呢？还是作 以色列 一支派一族的祭司好呢？”
JUDG|18|20|祭司心里欢喜，拿着以弗得和家中的神像，以及雕刻的像，跟这些百姓走了。
JUDG|18|21|他们转身离开那里，把孩子、牲畜、财物安排在前头。
JUDG|18|22|他们离了 米迦 的家已远， 米迦 家附近的邻居被召来，追赶 但 人。
JUDG|18|23|他们呼叫 但 人， 但 人回头对 米迦 说：“你召集这许多人来做什么呢？”
JUDG|18|24|米迦 说：“你们把我所造的神像，还有祭司，都带走了，我还有什么呢？你怎么还对我说‘你在做什么’呢？”
JUDG|18|25|但 人对 米迦 说：“你不要让我们再听见你的声音，恐怕这群恼怒成性的人会攻击你们，你和你的全家就会丧命。”
JUDG|18|26|但 人仍走他们的路。 米迦 见他们的势力比自己强，就转身回家去了。
JUDG|18|27|但 人把 米迦 造的神像和他的祭司带走，来到 拉亿 安宁无虑的百姓那里，用刀杀了他们，放火烧了那城。
JUDG|18|28|没有人来搭救，因为这城离 西顿 很远，他们又与世无争；这城在靠近 伯．利合 的平原。 但 人建造这城，在那里居住，
JUDG|18|29|并照着他们祖先 以色列 之子 但 的名字，给这城起名叫 但 。原先这城名叫 拉亿 。
JUDG|18|30|但 人为自己设立了那雕刻的像。 摩西 的孙子， 革舜 的儿子 约拿单 和他的子孙作 但 支派的祭司，直到那地遭掳掠的日子。
JUDG|18|31|上帝的家在 示罗 多少日子， 但 人为自己设立 米迦 所雕刻的像也在 但 多少日子。
JUDG|19|1|当 以色列 中没有王的时候，有一个 利未 人寄居 以法莲 山区的边界，他娶了一个 犹大伯利恒 的女子为妾。
JUDG|19|2|这妾对丈夫生气 ，离开丈夫，回到 犹大伯利恒 的父家，在那里住了四个月。
JUDG|19|3|她的丈夫起来，带着一个仆人、两匹驴跟着她去，要用好话劝她回来。女子就带丈夫进到父亲家里。女子的父亲看见了他，就欢欢喜喜地迎接他。
JUDG|19|4|这岳父，就是女子的父亲，留他住了三天。他们在那里吃喝，住宿。
JUDG|19|5|第四日，他们清早起来， 利未 人起身要走，女子的父亲对女婿说：“先吃点东西，加添心力，然后你们才走。”
JUDG|19|6|于是二人坐下，一同吃喝。女子的父亲对那人说：“请你答应再住一夜，使你的心舒畅。”
JUDG|19|7|那人起身要走，他岳父挽留他，他就留下，在那里又住了一夜。
JUDG|19|8|第五日，他清早起来要走，女子的父亲说：“来，请加添心力，留到太阳偏西吧。”于是二人一同再吃。
JUDG|19|9|那人同他的妾和仆人起身要走，但他岳父，就是女子的父亲，对他说：“看哪，太阳下山，天快晚了，你们再住一夜吧。看哪，太阳偏西了，就在这里住宿，使你的心舒畅，明天你们一早起来上路，回你的帐棚去。”
JUDG|19|10|那人不愿再住一夜，就备上两匹驴，带着他的妾起身走了，来到 耶布斯 的对面， 耶布斯 就是 耶路撒冷 。
JUDG|19|11|将近 耶布斯 的时候，太阳快下山了，仆人对主人说：“来吧，我们进这 耶布斯 人的城，在这里住宿。”
JUDG|19|12|主人对他说：“我们不可进入外邦人的城，那不是 以色列 人的地方，我们越过这里到 基比亚 去吧。”
JUDG|19|13|他又对仆人说：“来，让我们到 基比亚 或 拉玛 的一个地方住宿。”
JUDG|19|14|于是他们越过那里往前走，将到 便雅悯 的 基比亚 的时候，太阳已经下山了。
JUDG|19|15|他们进入 基比亚 要在那里住宿。他来坐在城里的广场上，但没有人接待他们到家里住宿。
JUDG|19|16|看哪，晚上有一个老人从田间做工回来。他是 以法莲 山区的人，寄居在 基比亚 ；那地方的人是 便雅悯 人。
JUDG|19|17|老人举目看见那过路的人在城里的广场上，就说：“你从哪里来？要到哪里去？”
JUDG|19|18|他对他说：“我们从 犹大 的 伯利恒 过来，要到 以法莲 山区的边界去。我是那里的人，去了 犹大 的 伯利恒 ，现在要到耶和华的家去，却没有人接待我到他的家。
JUDG|19|19|其实我有饲料草料可以喂驴，我和你的使女，以及与我们在一起的仆人都有饼有酒，什么都不缺。”
JUDG|19|20|老人说：“愿你平安！你所需用的我都会给你们，只是不可在广场上过夜。”
JUDG|19|21|于是老人领他到家里，喂上驴。他们洗了脚，就吃喝起来。
JUDG|19|22|他们心里欢乐的时候，看哪，城中的无赖围住房子，连连叩门，对老人，这家的主人说：“把那进你家的人带出来，我们要与他交合。”
JUDG|19|23|这家的主人出来对他们说：“弟兄们，不要做这样的恶事。这人既然进了我的家，你们就不要做这样可耻的事。
JUDG|19|24|看哪，我有个女儿还是处女，还有这人的妾，我把她们领出来任由你们污辱她们，就照你们看为好的对待她们吧！但对这人你们不要做这样可耻的事。”
JUDG|19|25|那些人却不肯听从他。那人抓住他的妾，把她拉出去给他们。他们强奸了她，整夜凌辱她，直到早晨，天色快亮才放她走。
JUDG|19|26|到了早晨，妇人回来，仆倒在留她主人住宿的那人的家门前，直到天亮。
JUDG|19|27|早晨，她的主人起来开了门，出去要上路。看哪，那妇人，他的妾倒在屋子门前，双手搭在门槛上。
JUDG|19|28|他对妇人说：“起来，我们走吧！”妇人却没有回应。那人就将她驮在驴上，起身回自己的地方去了。
JUDG|19|29|到了家里，他拿刀，抓住他的妾，把她的尸身切成十二块，分送到 以色列 全境。
JUDG|19|30|凡看见的人都说：“自从 以色列 人离开 埃及 地上来，直到今日，像这样的事还没有发生过，也没有见过。大家应当想一想，商讨一下再说。”
JUDG|20|1|于是 以色列 众人从 但 到 别是巴 ，以及从 基列 地出来，如同一人，聚集在 米斯巴 耶和华那里。
JUDG|20|2|以色列 各支派中众百姓的领袖，都站在上帝百姓的会中。拿刀的步兵共有四十万。
JUDG|20|3|便雅悯 人听见 以色列 人上了 米斯巴 。 以色列 人说：“请说，这恶事是怎么发生的呢？”
JUDG|20|4|那 利未 人，就是被害妇人的丈夫，回答说：“我和我的妾来到 便雅悯 的 基比亚 住宿。
JUDG|20|5|基比亚 人夜间起来攻击我，包围我住的屋子。他们想要杀我，并把我的妾污辱致死。
JUDG|20|6|我把我的妾切成块，分送到 以色列 得为业的全地，因为 基比亚 人在 以色列 中做了邪恶可耻的事。
JUDG|20|7|看哪，你们大家， 以色列 人哪，在此提出你们的建议和对策吧！”
JUDG|20|8|众百姓都起来如同一人，说：“我们谁也不回自己的帐棚，谁也不回自己的家去！
JUDG|20|9|现在，我们要这样对付 基比亚 ，照所抽的签去攻打他们。
JUDG|20|10|我们要在 以色列 各支派中，一百人选十人，一千人选一百人，一万人选一千人，为那到 便雅悯 的 迦巴 去的士兵运粮；因为 基比亚 在 以色列 中行了可耻的事。”
JUDG|20|11|于是 以色列 众人彼此联合如同一人，聚集攻击那城。
JUDG|20|12|以色列 众支派派人去，问 便雅悯 支派的各家说：“你们中间怎么做了这样的恶事呢？
JUDG|20|13|现在你们要把 基比亚 的那些无赖交出来，我们好处死他们，从 以色列 中除掉这恶。” 便雅悯 人却不肯听从他们弟兄 以色列 人的话。
JUDG|20|14|便雅悯 人从各城聚集到 基比亚 ，出来要与 以色列 人打仗。
JUDG|20|15|那日， 便雅悯 人从各城里征召了拿刀的士兵，共有二万六千，另外还从 基比亚 居民中征召七百个精兵。
JUDG|20|16|全军中有特选的七百个精兵，都是惯用左手的，个个能用机弦甩石，毫发不差。
JUDG|20|17|以色列 人，除了 便雅悯 之外，共征召了四十万拿刀的，个个都是战士。
JUDG|20|18|以色列 人起来，上到 伯特利 去求问上帝说：“我们中间谁当首先上去与 便雅悯 人争战呢？”耶和华说：“ 犹大 先上去。”
JUDG|20|19|以色列 人早晨起来，对着 基比亚 安营。
JUDG|20|20|以色列 人出来与 便雅悯 人打仗， 以色列 人在 基比亚 对着他们摆阵。
JUDG|20|21|便雅悯 人从 基比亚 出来，当日把 以色列 中二万二千人杀倒在地。
JUDG|20|22|以色列 人的士兵鼓起勇气，在第一日摆阵的地方又摆阵。
JUDG|20|23|因 以色列 人上去，在耶和华面前哀哭，直到晚上。他们求问耶和华说：“我可以再出兵与我弟兄 便雅悯 人打仗吗？”耶和华说：“可以上去攻打他们。”
JUDG|20|24|第二日， 以色列 人就上前攻击 便雅悯 人。
JUDG|20|25|便雅悯 人也在第二日从 基比亚 出来与他们交战，又把 以色列 人一万八千个拿刀的士兵杀倒在地。
JUDG|20|26|以色列 众人和全体士兵上到 伯特利 ，坐在耶和华面前哭泣。那日，他们禁食直到晚上，又在耶和华面前献燔祭和平安祭。
JUDG|20|27|以色列 人去求问耶和华；那时，上帝的约柜在那里。
JUDG|20|28|那时， 亚伦 的孙子， 以利亚撒 的儿子 非尼哈 侍立在约柜前。他们说：“我可以再出去与我弟兄 便雅悯 人打仗吗？还是停战呢？”耶和华说：“你们可以上去，因为明日我必把他交在你手中。”
JUDG|20|29|以色列 在 基比亚 的四围设下埋伏。
JUDG|20|30|第三日， 以色列 人又上去攻击 便雅悯 人，在 基比亚 前摆阵，与前两次一样。
JUDG|20|31|便雅悯 人也出来迎敌，就被引诱出城外。在田间的两条路上，一条通往 伯特利 ，一条通往 基比亚 ，他们像前两次一样，动手杀了约三十个 以色列 人。
JUDG|20|32|便雅悯 人说：“他们仍像以前一样败在我们面前。”但 以色列 人说：“让我们逃跑，引诱他们离开城到路上来。”
JUDG|20|33|以色列 众人都起来，在 巴力．他玛 摆阵， 以色列 的伏兵从 马利．迦巴 埋伏的地方冲上前去。
JUDG|20|34|全 以色列 中的一万精兵来到 基比亚 前，战争十分激烈。 便雅悯 人却不知道灾祸临近了。
JUDG|20|35|耶和华在 以色列 面前击打 便雅悯 。那日， 以色列 人歼灭二万五千一百个 便雅悯 人，都是拿刀的士兵。
JUDG|20|36|便雅悯 人看到自己战败了。 以色列 人因为信任在 基比亚 前所设的伏兵，就在 便雅悯 人面前假装撤退。
JUDG|20|37|伏兵迅速闯进 基比亚 ；他们继续前进，用刀杀死全城的人。
JUDG|20|38|以色列 人预先与伏兵约定在城内放火，以上腾的烟为信号。
JUDG|20|39|以色列 人从阵上撤退， 便雅悯 人动手杀死 以色列 人，约有三十个，就说：“他们仍像以前一样败在我们面前。”
JUDG|20|40|当烟如柱一般从城中上腾的时候， 便雅悯 人回头，看哪，全城已经浓烟冲天了。
JUDG|20|41|以色列 人又转身回来， 便雅悯 人就很惊惶，因为看见灾祸临到自己了。
JUDG|20|42|他们在 以色列 人面前转身往旷野逃跑，战况对他们不利，那从城里出来的也去夹攻，杀灭他们。
JUDG|20|43|以色列 人围攻 便雅悯 人，追赶他们，在他们歇脚之处，直到向日出方向的 基比亚 的对面，践踏他们。
JUDG|20|44|便雅悯 人倒下的有一万八千名，这些全都是勇士。
JUDG|20|45|其余的人转身往旷野逃跑，到 临门岩 去。 以色列 人在路上杀了五千人，如拾穗一样，紧追他们直到 基顿 ，又杀了二千人。
JUDG|20|46|那日 便雅悯 人倒下的有二万五千名，这些全都是拿刀的勇士。
JUDG|20|47|有六百人转身往旷野逃跑，到了 临门岩 ，在 临门岩 住了四个月。
JUDG|20|48|以色列 人又转回去攻击 便雅悯 人，凡经过的各城，其中的人和牲畜都用刀杀了，又放火烧了所经过的一切城镇。
JUDG|21|1|以色列 人在 米斯巴 曾起誓说：“我们中谁都不把女儿嫁给 便雅悯 人。”
JUDG|21|2|以色列 人来到 伯特利 ，坐在那里直到晚上，在上帝面前放声大哭，
JUDG|21|3|说：“耶和华－ 以色列 的上帝啊，为何 以色列 中会发生这样的事，使 以色列 今日缺了一个支派呢？”
JUDG|21|4|次日，百姓清早起来，在那里筑了一座坛，献燔祭和平安祭。
JUDG|21|5|以色列 人说：“ 以色列 各支派中，谁没有同会众一起上到耶和华那里呢？”因为 以色列 人曾起重誓说：“凡不上 米斯巴 到耶和华那里的，必被处死。”
JUDG|21|6|以色列 人怜悯他们的弟兄 便雅悯 ，说：“如今 以色列 中断绝一个支派了。
JUDG|21|7|我们既然向耶和华起誓说，必不把我们的女儿嫁给 便雅悯 人，现在我们该怎么办，使他们剩下的人可以娶妻呢？”
JUDG|21|8|他们又说：“ 以色列 支派中谁没有上 米斯巴 到耶和华那里呢？”看哪， 基列 的 雅比 没有一人进营到会众那里，
JUDG|21|9|百姓被数点的时候，看哪， 基列 的 雅比 居民没有一人在那里。
JUDG|21|10|会众就派一万二千名大勇士，吩咐他们说：“你们去用刀把 基列 的 雅比 居民连妇女带孩子都杀了。
JUDG|21|11|这是你们当做的事：要把所有男人和曾与男人同房共寝的女人全都杀了。”
JUDG|21|12|他们在 基列 的 雅比 居民中，找到四百个未曾与男人同房共寝的处女，就带她们到 迦南 地的 示罗 营里。
JUDG|21|13|全会众派人到 临门岩 的 便雅悯 人那里，与他们讲和。
JUDG|21|14|当时 便雅悯 人回来了， 以色列 人就把所留下， 基列 的 雅比 活着的女子嫁给他们，可是还是不够。
JUDG|21|15|百姓怜悯 便雅悯 人，因为耶和华使 以色列 支派中有一个缺口。
JUDG|21|16|会众中的长老说：“ 便雅悯 中的女子既然都除灭了，我们该怎么办，使剩下的人可以娶妻呢？”
JUDG|21|17|他们又说：“ 便雅悯 逃脱的人应当有地业，免得 以色列 中的一个支派被涂去。
JUDG|21|18|只是我们不能把自己的女儿嫁给他们。”因为 以色列 人曾起誓说：“把女儿嫁给 便雅悯 人的必受诅咒。”
JUDG|21|19|他们又说：“看哪，一年一度耶和华的节期正在 示罗 举行。” 示罗 位于 利波拿 的南边， 伯特利 的北边，从 伯特利 往 示剑 大路的东边。
JUDG|21|20|他们吩咐 便雅悯 人说：“你们去，躲在葡萄园中，
JUDG|21|21|观看；看哪，若 示罗 的女子出来跳舞，你们就从葡萄园出来，各人从 示罗 的女子中抢一个为妻，然后到 便雅悯 地去。
JUDG|21|22|他们的父亲或兄弟若来与我们争论，我们就对他们说：‘请看我们的情面恩待这些人吧！因为我们在战争的时候没有给他们任何人留下女子为妻。这次也不是你们给他们的，若是你们给的，就算有罪了。’”
JUDG|21|23|于是 便雅悯 人就照样做了，按照他们的人数，把从跳舞女子中抢来的娶为妻子，带回自己的地业，重建城镇，居住在其中。
JUDG|21|24|那时 以色列 人离开那里，各自回到自己的支派、宗族；他们从那里起行，各自回到自己的地业去了。
JUDG|21|25|那时， 以色列 中没有王，各人照自己眼中看为对的去做。
