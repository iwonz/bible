2SAM|1|1|По смерти Саула, когда Давид возвратился от поражения Амаликитян и пробыл в Секелаге два дня,
2SAM|1|2|вот, на третий день приходит человек из стана Саулова; одежда на нем разодрана и прах на голове его. Придя к Давиду, он пал на землю и поклонился [ему].
2SAM|1|3|И сказал ему Давид: откуда ты пришел? И сказал тот: я убежал из стана Израильского.
2SAM|1|4|И сказал ему Давид: что произошло? расскажи мне. И тот сказал: народ побежал со сражения, и множество из народа пало и умерло, и умерли и Саул и сын его Ионафан.
2SAM|1|5|И сказал Давид отроку, рассказывавшему ему: как ты знаешь, что Саул и сын его Ионафан умерли?
2SAM|1|6|И сказал отрок, рассказывавший ему: я случайно пришел на гору Гелвуйскую, и вот, Саул пал на свое копье, колесницы же и всадники настигали его.
2SAM|1|7|Тогда он оглянулся назад и, увидев меня, позвал меня.
2SAM|1|8|И я сказал: вот я. Он сказал мне: кто ты? И я сказал ему: я – Амаликитянин.
2SAM|1|9|Тогда он сказал мне: подойди ко мне и убей меня, ибо тоска смертная объяла меня, душа моя все еще во мне.
2SAM|1|10|И я подошел к нему и убил его, ибо знал, что он не будет жив после своего падения; и взял я венец, бывший на голове его, и запястье, бывшее на руке его, и принес их к господину моему сюда.
2SAM|1|11|Тогда схватил Давид одежды свои и разодрал их, также и все люди, бывшие с ним.
2SAM|1|12|и рыдали и плакали, и постились до вечера о Сауле и о сыне его Ионафане, и о народе Господнем и о доме Израилевом, что пали они от меча.
2SAM|1|13|И сказал Давид отроку, рассказывавшему ему: откуда ты? И сказал он: я – сын пришельца Амаликитянина.
2SAM|1|14|Тогда Давид сказал ему: как не побоялся ты поднять руку, чтобы убить помазанника Господня?
2SAM|1|15|И призвал Давид одного из отроков и сказал ему: подойди, убей его.
2SAM|1|16|И [тот] убил его, и он умер. И сказал к нему Давид: кровь твоя на голове твоей, ибо твои уста свидетельствовали на тебя, когда ты говорил: я убил помазанника Господня.
2SAM|1|17|И оплакал Давид Саула и сына его Ионафана сею плачевною песнью,
2SAM|1|18|и повелел научить сынов Иудиных луку, как написано в книге Праведного, и сказал:
2SAM|1|19|краса твоя, о Израиль, поражена на высотах твоих! как пали сильные!
2SAM|1|20|Не рассказывайте в Гефе, не возвещайте на улицах Аскалона, чтобы не радовались дочери Филистимлян, чтобы не торжествовали дочери необрезанных.
2SAM|1|21|Горы Гелвуйские! да [не сойдет] ни роса, ни дождь на вас, и да не будет [на вас] полей с плодами, ибо там повержен щит сильных, щит Саула, как бы не был он помазан елеем.
2SAM|1|22|Без крови раненых, без тука сильных лук Ионафана не возвращался назад, и меч Саула не возвращался даром.
2SAM|1|23|Саул и Ионафан, любезные и согласные в жизни своей, не разлучились и в смерти своей; быстрее орлов, сильнее львов [они были].
2SAM|1|24|Дочери Израильские! плачьте о Сауле, который одевал вас в багряницу с украшениями и доставлял на одежды ваши золотые уборы.
2SAM|1|25|Как пали сильные на брани! Сражен Ионафан на высотах твоих.
2SAM|1|26|Скорблю о тебе, брат мой Ионафан; ты был очень дорог для меня; любовь твоя была для меня превыше любви женской.
2SAM|1|27|Как пали сильные, погибло оружие бранное!
2SAM|2|1|После сего Давид вопросил Господа, говоря: идти ли мне в какой–либо из городов Иудиных? И сказал ему Господь: иди. И сказал Давид: куда идти? И сказал Он: в Хеврон.
2SAM|2|2|И пошел туда Давид и обе жены его, Ахиноама Изреелитянка и Авигея, [бывшая] жена Навала, Кармилитянка.
2SAM|2|3|И людей, бывших с ним, привел Давид, каждого с семейством его, и поселились в городе Хевроне.
2SAM|2|4|И пришли мужи Иудины и помазали там Давида на царство над домом Иудиным. И донесли Давиду, что жители Иависа Галаадского погребли Саула.
2SAM|2|5|И отправил Давид послов к жителям Иависа Галаадского, сказать им: благословенны вы у Господа за то, что оказали эту милость господину своему Саулу, и погребли его.
2SAM|2|6|и ныне да воздаст вам Господь милостью и истиною; и я сделаю вам благодеяние за то, что вы это сделали;
2SAM|2|7|ныне да укрепятся руки ваши, и будьте мужественны; ибо господин ваш Саул умер, а меня помазал дом Иудин царем над собою.
2SAM|2|8|Но Авенир, сын Ниров, начальник войска Саулова, взял Иевосфея, сына Саулова, и привел его в Маханаим,
2SAM|2|9|и воцарил его над Галаадом, и Ашуром, и Изреелем, и Ефремом, и Вениамином, и над всем Израилем.
2SAM|2|10|Сорок лет было Иевосфею, сыну Саулову, когда он воцарился над Израилем, и царствовал два года. Только дом Иудин остался с Давидом.
2SAM|2|11|Всего времени, в которое Давид царствовал в Хевроне над домом Иудиным, было семь лет и шесть месяцев.
2SAM|2|12|И вышел Авенир, сын Ниров, и слуги Иевосфея, сына Саулова, из Маханаима в Гаваон.
2SAM|2|13|Вышел и Иоав, сын Саруи, со слугами Давида, и встретились у Гаваонского пруда, и засели те на одной стороне пруда, а эти на другой стороне пруда.
2SAM|2|14|И сказал Авенир Иоаву: пусть встанут юноши и поиграют пред нами. И сказал Иоав: пусть встанут.
2SAM|2|15|И встали и пошли числом двенадцать Вениамитян со стороны Иевосфея, сына Саулова, и двенадцать из слуг Давидовых.
2SAM|2|16|Они схватили друг друга за голову, [вонзили] меч один другому в бок и пали вместе. И было названо это место Хелкаф–Хаццурим, что в Гаваоне.
2SAM|2|17|И произошло в тот день жесточайшее сражение, и Авенир с людьми Израильскими был поражен слугами Давида.
2SAM|2|18|И были там три сына Саруи: Иоав, и Авесса, и Асаил. Асаил же был легок на ноги, как серна в поле.
2SAM|2|19|И погнался Асаил за Авениром и преследовал его, не уклоняясь ни направо, ни налево от следов Авенира.
2SAM|2|20|И оглянулся Авенир назад и сказал: ты ли это, Асаил? Тот сказал: я.
2SAM|2|21|И сказал ему Авенир: уклонись направо или налево, и выбери себе одного из отроков и возьми себе его вооружение. Но Асаил не захотел отстать от него.
2SAM|2|22|И повторил Авенир еще, говоря Асаилу: отстань от меня, чтоб я не поверг тебя на землю; тогда с каким лицем явлюсь я к Иоаву, брату твоему?
2SAM|2|23|Но тот не захотел отстать. Тогда Авенир, поворотив копье, поразил его в живот; копье прошло насквозь его, и он упал там же и умер на месте. Все проходившие чрез то место, где пал и умер Асаил, останавливались.
2SAM|2|24|И преследовали Иоав и Авесса Авенира. Солнце уже зашло, когда они пришли к холму Амма, что против Гиаха, на дороге к пустыне Гаваонской.
2SAM|2|25|И собрались Вениамитяне вокруг Авенира и составили одно ополчение, и стали на вершине одного холма.
2SAM|2|26|И воззвал Авенир к Иоаву, и сказал: вечно ли будет пожирать меч? Или ты не знаешь, что последствия будут горестные? И доколе ты не скажешь людям, чтобы они перестали преследовать братьев своих?
2SAM|2|27|И сказал Иоав: жив Бог! если бы ты не говорил иначе, то еще утром перестали бы люди преследовать братьев своих.
2SAM|2|28|И затрубил Иоав трубою, и остановился весь народ, и не преследовали более Израильтян; сражение прекратилось.
2SAM|2|29|Авенир же и люди его шли равниною всю ту ночь и перешли Иордан, и прошли весь Битрон, и пришли в Маханаим.
2SAM|2|30|И возвратился Иоав от преследования Авенира и собрал весь народ, и недоставало из слуг Давидовых девятнадцати человек кроме Асаила.
2SAM|2|31|Слуги же Давидовы поразили Вениамитян и людей Авенировых; пало их триста шестьдесят человек.
2SAM|2|32|И взяли Асаила и похоронили его во гробе отца его, что в Вифлееме. Иоав же с людьми своими шел всю ночь и на рассвете прибыл в Хеврон.
2SAM|3|1|И была продолжительная распря между домом Сауловым и домом Давидовым. Давид все более и более усиливался, а дом Саулов более и более ослабевал.
2SAM|3|2|И родились у Давида сыновей в Хевроне. Первенец его был Амнон от Ахиноамы Изреелитянки,
2SAM|3|3|а второй [сын] его – Далуиа от Авигеи, [бывшей] жены Навала, Кармилитянки; третий – Авессалом, сын Маахи, дочери Фалмая, царя Гессурского;
2SAM|3|4|четвертый – Адония, сын Аггифы; пятый – Сафатия, сын Авиталы;
2SAM|3|5|шестой – Иефераам от Эглы, жены Давидовой. Они родились у Давида в Хевроне.
2SAM|3|6|Когда была распря между домом Саула и домом Давида, то Авенир поддерживал дом Саула.
2SAM|3|7|У Саула была наложница, по имени Рицпа, дочь Айя. И сказал [Иевосфей] Авениру: зачем ты вошел к наложнице отца моего?
2SAM|3|8|Авенир же сильно разгневался на слова Иевосфея и сказал: разве я – собачья голова? Я против Иуды оказал ныне милость дому Саула, отца твоего, братьям его и друзьям его, и не предал тебя в руки Давида, а ты взыскиваешь ныне на мне грех из–за женщины.
2SAM|3|9|То и то пусть сделает Бог Авениру и еще больше сделает ему! Как клялся Господь Давиду, так и сделаю ему:
2SAM|3|10|отниму царство от дома Саулова и поставлю престол Давида над Израилем и над Иудою, от Дана до Вирсавии.
2SAM|3|11|И не мог Иевосфей возразить Авениру, ибо боялся его.
2SAM|3|12|И послал Авенир от себя послов к Давиду, сказать: чья эта земля? И еще сказать: заключи союз со мною, и рука моя будет с тобою, чтобы обратить к тебе весь народ Израильский.
2SAM|3|13|И сказал [Давид]: хорошо, я заключу союз с тобою, только прошу тебя об одном, именно – ты не увидишь лица моего, если не приведешь с собою Мелхолы, дочери Саула, когда придешь увидеться со мною.
2SAM|3|14|И отправил Давид послов к Иевосфею, сыну Саулову, сказать: отдай жену мою Мелхолу, которую я получил за сто краеобрезаний Филистимских.
2SAM|3|15|И послал Иевосфей и взял ее от мужа, от Фалтия, сына Лаишева.
2SAM|3|16|Пошел с нею и муж ее и с плачем провожал ее до Бахурима; но Авенир сказал ему: ступай назад. И он возвратился.
2SAM|3|17|И обратился Авенир к старейшинам Израильским, говоря: и вчера и третьего дня вы желали, чтобы Давид был царем над вами,
2SAM|3|18|теперь сделайте [это], ибо Господь сказал Давиду: "рукою раба Моего Давида Я спасу народ Мой Израиля от руки Филистимлян и от руки всех врагов его".
2SAM|3|19|То же говорил Авенир и Вениамитянам. И пошел Авенир в Хеврон, чтобы пересказать Давиду все, чего желали Израиль и весь дом Вениаминов.
2SAM|3|20|И пришел Авенир к Давиду в Хеврон и с ним двадцать человек, и сделал Давид пир для Авенира и людей, бывших с ним.
2SAM|3|21|И сказал Авенир Давиду: я встану и пойду и соберу к господину моему царю весь народ Израильский, и они вступят в завет с тобою, и будешь царствовать над всеми, как желает душа твоя. И отпустил Давид Авенира, и он ушел с миром.
2SAM|3|22|И вот, слуги Давидовы с Иоавом пришли из похода и принесли с собою много добычи; но Авенира уже не было с Давидом в Хевроне, ибо [Давид] отпустил его, и он ушел с миром.
2SAM|3|23|Когда Иоав и все войско, ходившее с ним, пришли, то Иоаву рассказали: приходил Авенир, сын Ниров, к царю, и тот отпустил его, и он ушел с миром.
2SAM|3|24|И пришел Иоав к царю и сказал: что ты сделал? Вот, приходил к тебе Авенир; зачем ты отпустил его, и он ушел?
2SAM|3|25|Ты знаешь Авенира, сына Нирова: он приходил обмануть тебя, узнать выход твой и вход твой и разведать все, что ты делаешь.
2SAM|3|26|И вышел Иоав от Давида и послал гонцов вслед за Авениром; и возвратили они его от колодезя Сира, без ведома Давида.
2SAM|3|27|Когда Авенир возвратился в Хеврон, то Иоав отвел его внутрь ворот, как будто для того, чтобы поговорить с ним тайно, и там поразил его в живот. И умер [Авенир] за кровь Асаила, брата Иоавова.
2SAM|3|28|И услышал после Давид [об этом] и сказал: невинен я и царство мое вовек пред Господом в крови Авенира, сына Нирова;
2SAM|3|29|пусть падет она на голову Иоава и на весь дом отца его; пусть никогда не остается дом Иоава без семеноточивого, или прокаженного, или опирающегося на посох, или падающего от меча, или нуждающегося в хлебе.
2SAM|3|30|Иоав же и брат его Авесса убили Авенира за то, что он умертвил брата их Асаила в сражении у Гаваона.
2SAM|3|31|И сказал Давид Иоаву и всем людям, бывшим с ним: раздерите одежды ваши и оденьтесь во вретища и плачьте над Авениром. И царь Давид шел за гробом [его].
2SAM|3|32|Когда погребали Авенира в Хевроне, то царь громко плакал над гробом Авенира; плакал и весь народ.
2SAM|3|33|И оплакал царь Авенира, говоря: смертью ли подлого умирать Авениру?
2SAM|3|34|Руки твои не были связаны, и ноги твои не в оковах, и ты пал, как падают от разбойников. И весь народ стал еще более плакать над ним.
2SAM|3|35|И пришел весь народ предложить Давиду хлеба, когда еще продолжался день; но Давид поклялся, говоря: то и то пусть сделает со мною Бог и еще больше сделает, если я до захождения солнца вкушу хлеба или чего–нибудь.
2SAM|3|36|И весь народ узнал это, и понравилось ему это, как и все, что делал царь, нравилось всему народу.
2SAM|3|37|И узнал весь народ и весь Израиль в тот день, что не от царя произошло умерщвление Авенира, сына Нирова.
2SAM|3|38|И сказал царь слугам своим: знаете ли, что вождь и великий муж пал в этот день в Израиле?
2SAM|3|39|Я теперь еще слаб, хотя и помазан на царство, а эти люди, сыновья Саруи, сильнее меня; пусть же воздаст Господь делающему злое по злобе его!
2SAM|4|1|И услышал [Иевосфей], сын Саулов, что умер Авенир в Хевроне, и опустились руки его, и весь Израиль смутился.
2SAM|4|2|У [Иевосфея], сына Саулова, два было предводителя войска; имя одного – Баана и имя другого – Рихав, сыновья Реммона Беерофянина, из потомков Вениаминовых, ибо и Беероф причислялся к Вениамину.
2SAM|4|3|И убежали Беерофяне в Гиффаим и остались там пришельцами до сего дня.
2SAM|4|4|У Ионафана, сына Саулова, был сын хромой. Пять лет было ему, когда пришло известие о Сауле и Ионафане из Изрееля, и нянька, взяв его, побежала. И когда она бежала поспешно, то он упал, и сделался хромым. Имя его Мемфивосфей.
2SAM|4|5|И пошли сыны Реммона Беерофянина, Рихав и Баана, и пришли в самый жар дня к дому Иевосфея; а он спал на постели в полдень.
2SAM|4|6|Рихав и Баана, брат его, вошли внутрь дома, [как бы] для того, чтобы взять пшеницы; и поразили его в живот и убежали.
2SAM|4|7|Когда они вошли в дом, [Иевосфей] лежал на постели своей, в спальной комнате своей; и они поразили его, и умертвили его, и отрубили голову его, и взяли голову его с собою, и шли пустынною дорогою всю ночь;
2SAM|4|8|и принесли голову Иевосфея к Давиду в Хеврон и сказали царю: вот голова Иевосфея, сына Саула, врага твоего, который искал души твоей; ныне Господь отмстил за господина моего царя Саулу и потомству его.
2SAM|4|9|И отвечал Давид Рихаву и Баане, брату его, сыновьям Реммона Беерофянина, и сказал им: жив Господь, избавивший душу мою от всякой скорби!
2SAM|4|10|если того, кто принес мне известие, сказав: "вот, умер Саул", и кто считал себя радостным вестником, я схватил и убил его в Секелаге, вместо того, чтобы дать ему награду,
2SAM|4|11|то теперь, когда негодные люди убили человека невинного в его доме на постели его, неужели я не взыщу крови его от руки вашей и не истреблю вас с земли?
2SAM|4|12|И приказал Давид слугам, и убили их, и отрубили им руки и ноги, и повесили их над прудом в Хевроне. А голову Иевосфея взяли и погребли во гробе Авенира, в Хевроне.
2SAM|5|1|И пришли все колена Израилевы к Давиду в Хеврон и сказали: вот, мы – кости твои и плоть твоя;
2SAM|5|2|еще вчера и третьего дня, когда Саул царствовал над нами, ты выводил и вводил Израиля; и сказал Господь тебе: "ты будешь пасти народ Мой Израиля и ты будешь вождем Израиля".
2SAM|5|3|И пришли все старейшины Израиля к царю в Хеврон, и заключил с ними царь Давид завет в Хевроне пред Господом; и помазали Давида в царя над Израилем.
2SAM|5|4|Тридцать лет было Давиду, когда он воцарился; царствовал сорок лет.
2SAM|5|5|В Хевроне царствовал над Иудою семь лет и шесть месяцев, и в Иерусалиме царствовал тридцать три года над всем Израилем и Иудою.
2SAM|5|6|И пошел царь и люди его на Иерусалим против Иевусеев, жителей той страны; но они говорили Давиду: "ты не войдешь сюда; тебя отгонят слепые и хромые", – это значило: "не войдет сюда Давид".
2SAM|5|7|Но Давид взял крепость Сион: это – город Давидов.
2SAM|5|8|И сказал Давид в тот день: всякий, убивая Иевусеев, пусть поражает копьем и хромых и слепых, ненавидящих душу Давида. Посему и говорится: слепой и хромой не войдет в дом [Господень].
2SAM|5|9|И поселился Давид в крепости, и назвал ее городом Давидовым, и обстроил кругом от Милло и внутри.
2SAM|5|10|И преуспевал Давид и возвышался, и Господь Бог Саваоф [был] с ним.
2SAM|5|11|И прислал Хирам, царь Тирский, послов к Давиду и кедровые деревья и плотников и каменщиков, и они построили дом Давиду.
2SAM|5|12|И уразумел Давид, что Господь утвердил его царем над Израилем и что возвысил царство его ради народа Своего Израиля.
2SAM|5|13|И взял Давид еще наложниц и жен из Иерусалима, после того, как пришел из Хеврона.
2SAM|5|14|И родились еще у Давида сыновья и дочери. И вот имена родившихся у него в Иерусалиме: Самус, и Совав, и Нафан, и Соломон,
2SAM|5|15|и Евеар, и Елисуа, и Нафек, и Иафиа,
2SAM|5|16|и Елисама, и Елидае, и Елифалеф.
2SAM|5|17|Когда Филистимляне услышали, что Давида помазали на царство над Израилем, то поднялись все Филистимляне искать Давида. И услышал Давид и пошел в крепость.
2SAM|5|18|А Филистимляне пришли и расположились в долине Рефаим.
2SAM|5|19|И вопросил Давид Господа, говоря: идти ли мне против Филистимлян? предашь ли их в руки мои? И сказал Господь Давиду: иди, ибо Я предам Филистимлян в руки твои.
2SAM|5|20|И пошел Давид в Ваал–Перацим и поразил их там, и сказал Давид: Господь разнес врагов моих предо мною, как разносит вода. Посему и месту тому дано имя Ваал–Перацим.
2SAM|5|21|И оставили там [Филистимляне] истуканов своих, а Давид с людьми своими взял их.
2SAM|5|22|И пришли опять Филистимляне и расположились в долине Рефаим.
2SAM|5|23|И вопросил Давид Господа, И Он отвечал ему: не выходи навстречу им, а зайди им с тылу и иди к ним со стороны тутовой рощи;
2SAM|5|24|и когда услышишь шум как бы идущего по вершинам тутовых дерев, то двинься, ибо тогда пошел Господь пред тобою, чтобы поразить войско Филистимское.
2SAM|5|25|И сделал Давид, как повелел ему Господь, и поразил Филистимлян от Гаваи до Газера.
2SAM|6|1|И собрал снова Давид всех отборных [людей] из Израиля, тридцать тысяч.
2SAM|6|2|И встал и пошел Давид и весь народ, бывший с ним из Ваала Иудина, чтобы перенести оттуда ковчег Божий, на котором нарицается имя Господа Саваофа, сидящего на херувимах.
2SAM|6|3|И поставили ковчег Божий на новую колесницу и вывезли его из дома Аминадава, что на холме. Сыновья же Аминадава, Оза и Ахио, вели новую колесницу.
2SAM|6|4|И повезли ее с ковчегом Божиим из дома Аминадава, что на холме; и Ахио шел пред ковчегом.
2SAM|6|5|А Давид и все сыны Израилевы играли пред Господом на всяких музыкальных орудиях из кипарисового дерева, и на цитрах, и на псалтирях, и на тимпанах, и на систрах, и на кимвалах.
2SAM|6|6|И когда дошли до гумна Нахонова, Оза простер руку свою к ковчегу Божию и взялся за него, ибо волы наклонили его.
2SAM|6|7|Но Господь прогневался на Озу, и поразил его Бог там же за дерзновение, и умер он там у ковчега Божия.
2SAM|6|8|И опечалился Давид, что Господь поразил Озу. Место сие и доныне называется: "поражение Озы".
2SAM|6|9|И устрашился Давид в тот день Господа и сказал: как войти ко мне ковчегу Господню?
2SAM|6|10|И не захотел Давид везти ковчег Господень к себе, в город Давидов, а обратил его в дом Аведдара Гефянина.
2SAM|6|11|И оставался ковчег Господень в доме Аведдара Гефянина три месяца, и благословил Господь Аведдара и весь дом его.
2SAM|6|12|Когда донесли царю Давиду, говоря: "Господь благословил дом Аведдара и все, что было у него, ради ковчега Божия", то пошел Давид и с торжеством перенес ковчег Божий из дома Аведдара в город Давидов.
2SAM|6|13|И когда несшие ковчег Господень проходили по шести шагов, он приносил в жертву тельца и овна.
2SAM|6|14|Давид скакал из всей силы пред Господом; одет же был Давид в льняной ефод.
2SAM|6|15|Так Давид и весь дом Израилев несли ковчег Господень с восклицаниями и трубными звуками.
2SAM|6|16|Когда входил ковчег Господень в город Давидов, Мелхола, дочь Саула, смотрела в окно и, увидев царя Давида, скачущего и пляшущего пред Господом, уничижила его в сердце своем.
2SAM|6|17|И принесли ковчег Господень и поставили его на своем месте посреди скинии, которую устроил для него Давид; и принес Давид всесожжения пред Господом и жертвы мирные.
2SAM|6|18|Когда Давид окончил приношение всесожжений и жертв мирных, то благословил он народ именем Господа Саваофа;
2SAM|6|19|и роздал всему народу, всему множеству Израильтян, как мужчинам, так и женщинам, по одному хлебу и по куску жареного мяса и по одной лепешке каждому. И пошел весь народ, каждый в дом свой.
2SAM|6|20|Когда Давид возвратился, чтобы благословить дом свой, то Мелхола, дочь Саула, вышла к нему на встречу и сказала: как отличился сегодня царь Израилев, обнажившись сегодня пред глазами рабынь рабов своих, как обнажается какой–нибудь пустой человек!
2SAM|6|21|И сказал Давид Мелхоле: пред Господом, Который предпочел меня отцу твоему и всему дому его, утвердив меня вождем народа Господня, Израиля; пред Господом играть и плясать буду;
2SAM|6|22|и я еще больше уничижусь, и сделаюсь еще ничтожнее в глазах моих, и пред служанками, о которых ты говоришь, я буду славен.
2SAM|6|23|И у Мелхолы, дочери Сауловой, не было детей до дня смерти ее.
2SAM|7|1|Когда царь жил в доме своем, и Господь успокоил его от всех окрестных врагов его,
2SAM|7|2|тогда сказал царь пророку Нафану: вот, я живу в доме кедровом, а ковчег Божий находится под шатром.
2SAM|7|3|И сказал Нафан царю: все, что у тебя на сердце, иди, делай; ибо Господь с тобою.
2SAM|7|4|Но в ту же ночь было слово Господа к Нафану:
2SAM|7|5|пойди, скажи рабу Моему Давиду: так говорит Господь: ты ли построишь Мне дом для Моего обитания,
2SAM|7|6|когда Я не жил в доме с того времени, как вывел сынов Израилевых из Египта, и до сего дня, но переходил в шатре и в скинии?
2SAM|7|7|Где Я ни ходил со всеми сынами Израиля, говорил ли Я хотя слово какому–либо из колен, которому Я назначил пасти народ Мой Израиля: "почему не построите Мне кедрового дома"?
2SAM|7|8|И теперь так скажи рабу Моему Давиду: так говорит Господь Саваоф: Я взял тебя от стада овец, чтобы ты был вождем народа Моего, Израиля;
2SAM|7|9|и был с тобою везде, куда ни ходил ты, и истребил всех врагов твоих пред лицем твоим, и сделал имя твое великим, как имя великих на земле.
2SAM|7|10|И Я устрою место для народа Моего, для Израиля, и укореню его, и будет он спокойно жить на месте своем, и не будет тревожиться больше, и люди нечестивые не станут более теснить его, как прежде,
2SAM|7|11|с того времени, как Я поставил судей над народом Моим, Израилем; и Я успокою тебя от всех врагов твоих. И Господь возвещает тебе, что Он устроит тебе дом.
2SAM|7|12|Когда же исполнятся дни твои, и ты почиешь с отцами твоими, то Я восставлю после тебя семя твое, которое произойдет из чресл твоих, и упрочу царство его.
2SAM|7|13|Он построит дом имени Моему, и Я утвержу престол царства его на веки.
2SAM|7|14|Я буду ему отцом, и он будет Мне сыном; и если он согрешит, Я накажу его жезлом мужей и ударами сынов человеческих;
2SAM|7|15|но милости Моей не отниму от него, как Я отнял от Саула, которого Я отверг пред лицем твоим.
2SAM|7|16|И будет непоколебим дом твой и царство твое на веки пред лицем Моим, и престол твой устоит во веки.
2SAM|7|17|Все эти слова и все это видение Нафан пересказал Давиду.
2SAM|7|18|И пошел царь Давид, и предстал пред лицем Господа, и сказал: кто я, Господи, Господи, и что такое дом мой, что Ты меня так возвеличил!
2SAM|7|19|И этого еще мало показалось в очах Твоих, Господи мой, Господи; но Ты возвестил еще о доме раба Твоего вдаль. Это уже по–человечески. Господи мой, Господи!
2SAM|7|20|Что еще может сказать Тебе Давид? Ты знаешь раба Твоего, Господи мой, Господи!
2SAM|7|21|Ради слова Твоего и по сердцу Твоему Ты делаешь это, открывая все это великое рабу Твоему.
2SAM|7|22|По всему велик Ты, Господи мой, Господи! ибо нет подобного Тебе и нет Бога, кроме Тебя, по всему, что слышали мы своими ушами.
2SAM|7|23|И кто подобен народу Твоему, Израилю, единственному народу на земле, для которого приходил Бог, чтобы приобрести [его] Себе в народ и прославить Свое имя [и] совершить великое и страшное пред народом Твоим, который Ты приобрел Себе от Египтян, изгнав народы и богов их?
2SAM|7|24|И Ты укрепил за Собою народ Твой, Израиля, как собственный народ, на веки, и Ты, Господи, сделался его Богом.
2SAM|7|25|И ныне, Господи Боже, утверди на веки слово, которое изрек Ты о рабе Твоем и о доме его, и исполни то, что Ты изрек.
2SAM|7|26|И да возвеличится имя Твое во веки, чтобы говорили: "Господь Саваоф – Бог над Израилем". И дом раба Твоего Давида да будет тверд пред лицем Твоим.
2SAM|7|27|Так как ты, Господи Саваоф, Боже Израилев, открыл рабу Твоему, говоря: "устрою тебе дом", то раб Твой уготовал сердце свое, чтобы молиться Тебе такою молитвою.
2SAM|7|28|Итак, Господи мой, Господи! Ты Бог, и слова Твои непреложны, и Ты возвестил рабу Твоему такое благо!
2SAM|7|29|И ныне начни и благослови дом раба Твоего, чтоб он был вечно пред лицем Твоим, ибо Ты, Господи мой, Господи, возвестил это, и благословением Твоим соделается дом раба Твоего благословенным во веки.
2SAM|8|1|После сего Давид поразил Филистимлян и смирил их, и взял Давид Мефег–Гаамма из рук Филистимлян.
2SAM|8|2|И поразил Моавитян и смерил их веревкою, положив их на землю; и отмерил две веревки на умерщвление, а одну веревку на оставление в живых. И сделались Моавитяне у Давида рабами, платящими дань.
2SAM|8|3|И поразил Давид Адраазара, сына Реховова, царя Сувского, когда тот шел, чтоб восстановить свое владычество при реке [Евфрате];
2SAM|8|4|и взял Давид у него тысячу семьсот всадников и двадцать тысяч человек пеших, и подрезал Давид жилы у всех коней колесничных, оставив [себе] из них для ста колесниц.
2SAM|8|5|И пришли Сирийцы Дамасские на помощь к Адраазару, царю Сувскому; но Давид поразил двадцать две тысячи человек Сирийцев.
2SAM|8|6|И поставил Давид охранные войска в Сирии Дамасской, и стали Сирийцы у Давида рабами, платящими дань. И хранил Господь Давида везде, куда он ни ходил.
2SAM|8|7|И взял Давид золотые щиты, которые были у рабов Адраазара, и принес их в Иерусалим.
2SAM|8|8|А в Бефе и Берофе, городах Адраазаровых, взял царь Давид весьма много меди.
2SAM|8|9|И услышал Фой, царь Имафа, что Давид поразил все войско Адраазарово,
2SAM|8|10|и послал Фой Иорама, сына своего, к царю Давиду, приветствовать его и благодарить его за то, что он воевал с Адраазаром и поразил его; ибо Адраазар вел войны с Фоем. В руках же [Иорама] были сосуды серебряные, золотые и медные.
2SAM|8|11|Их также посвятил царь Давид Господу, вместе с серебром и золотом, которое посвятил из [отнятого] у всех покоренных им народов:
2SAM|8|12|у Сирийцев, и Моавитян, и Аммонитян, и Филистимлян, и Амаликитян, и из отнятого у Адраазара, сына Реховова, царя Сувского.
2SAM|8|13|И сделал Давид себе имя, возвращаясь с поражения восемнадцати тысяч Сирийцев в долине Соленой.
2SAM|8|14|И поставил он охранные войска в Идумее; во всей Идумее поставил охранные войска, и все Идумеяне были рабами Давиду. И хранил Господь Давида везде, куда он ни ходил.
2SAM|8|15|И царствовал Давид над всем Израилем, и творил Давид суд и правду над всем народом своим.
2SAM|8|16|Иоав же, сын Саруи, [был начальником] войска; и Иосафат, сын Ахилуда, – дееписателем;
2SAM|8|17|Садок, сын Ахитува, и Ахимелех, сын Авиафара, – священниками, Сераия – писцом;
2SAM|8|18|и Ванея, сын Иодая – [начальником] над Хелефеями и Фелефеями, и сыновья Давида – первыми при дворе.
2SAM|9|1|И сказал Давид: не остался ли еще кто–нибудь из дома Саулова? я оказал бы ему милость ради Ионафана.
2SAM|9|2|В доме Саула был раб, по имени Сива; и позвали его к Давиду, и сказал ему царь: ты ли Сива? И тот сказал: я, раб твой.
2SAM|9|3|И сказал царь: нет ли еще кого–нибудь из дома Саулова? я оказал бы ему милость Божию. И сказал Сива царю: есть сын Ионафана, хромой ногами.
2SAM|9|4|И сказал ему царь: где он? И сказал Сива царю: вот, он в доме Махира, сына Аммиэлова, в Лодеваре.
2SAM|9|5|И послал царь Давид, и взяли его из дома Махира, сына Аммиэлова, из Лодевара.
2SAM|9|6|И пришел Мемфивосфей, сын Ионафана, сына Саулова, к Давиду, и пал на лице свое, и поклонился. И сказал Давид: Мемфивосфей! И сказал тот: вот раб твой.
2SAM|9|7|И сказал ему Давид: не бойся; я окажу тебе милость ради отца твоего Ионафана и возвращу тебе все поля Саула, отца твоего, и ты всегда будешь есть хлеб за моим столом.
2SAM|9|8|И поклонился [Мемфивосфей] и сказал: что такое раб твой, что ты призрел на такого мертвого пса, как я?
2SAM|9|9|И призвал царь Сиву, слугу Саула, и сказал ему: все, что принадлежало Саулу и всему дому его, я отдаю сыну господина твоего;
2SAM|9|10|итак обрабатывай для него землю ты и сыновья твои и рабы твои, и доставляй [плоды ее], чтобы у сына господина твоего был хлеб для пропитания; Мемфивосфей же, сын господина твоего, всегда будет есть за моим столом. У Сивы было пятнадцать сыновей и двадцать рабов.
2SAM|9|11|И сказал Сива царю: все, что приказывает господин мой царь рабу своему, исполнит раб твой. Мемфивосфей ел за столом [Давида], как один из сыновей царя.
2SAM|9|12|У Мемфивосфея был малолетний сын, по имени Миха. Все живущие в доме Сивы были рабами Мемфивосфея.
2SAM|9|13|И жил Мемфивосфей в Иерусалиме, ибо он ел всегда за царским столом. Он был хром на обе ноги.
2SAM|10|1|Спустя несколько времени умер царь Аммонитский, и воцарился вместо него сын его Аннон.
2SAM|10|2|И сказал Давид: окажу я милость Аннону, сыну Наасову, за благодеяние, которое оказал мне отец его. И послал Давид слуг своих утешить Аннона об отце его. И пришли слуги Давидовы в землю Аммонитскую.
2SAM|10|3|Но князья Аммонитские сказали Аннону, господину своему: неужели ты думаешь, что Давид из уважения к отцу твоему прислал к тебе утешителей? не для того ли, чтобы осмотреть город и высмотреть в нем и [после] разрушить его, прислал Давид слуг своих к тебе?
2SAM|10|4|И взял Аннон слуг Давидовых, и обрил каждому из них половину бороды, и обрезал одежды их наполовину, до чресл, и отпустил их.
2SAM|10|5|Когда донесли об этом Давиду, то он послал к ним навстречу, так как они были очень обесчещены. И велел царь сказать им: оставайтесь в Иерихоне, пока отрастут бороды ваши, и [тогда] возвратитесь.
2SAM|10|6|И увидели Аммонитяне, что они сделались ненавистными для Давида; и послали Аммонитяне нанять Сирийцев из Беф–Рехова и Сирийцев Сувы двадцать тысяч пеших, у царя Маахи тысячу человек и из Истова двенадцать тысяч человек.
2SAM|10|7|Когда услышал об этом Давид, то послал Иоава со всем войском храбрых.
2SAM|10|8|И вышли Аммонитяне и расположились к сражению у ворот, а Сирийцы Сувы и Рехова, и Истова, и Маахи, [стали] отдельно в поле.
2SAM|10|9|И увидел Иоав, что неприятельское войско было поставлено против него и спереди и сзади, и избрал [воинов] из всех отборных в Израиле, и выстроил их против Сирийцев;
2SAM|10|10|остальную же часть людей поручил Авессе, брату своему, чтоб он выстроил их против Аммонитян.
2SAM|10|11|И сказал [Иоав]: если Сирийцы будут одолевать меня, ты поможешь мне; а если Аммонитяне тебя будут одолевать, я приду к тебе на помощь;
2SAM|10|12|будь мужествен, и будем стоять твердо за народ наш и за города Бога нашего, а Господь сделает, что Ему угодно.
2SAM|10|13|И вступил Иоав в народ, который [был] у него, в сражение с Сирийцами, и они побежали от него.
2SAM|10|14|Аммонитяне же, увидев, что Сирийцы бегут, побежали от Авессы и ушли в город. И возвратился Иоав от Аммонитян и пришел в Иерусалим.
2SAM|10|15|Сирийцы, видя, что они поражены Израильтянами, собрались вместе.
2SAM|10|16|И послал Адраазар и призвал Сирийцев, которые за рекою, и пришли они к Еламу; а Совак, военачальник Адраазаров, предводительствовал ими.
2SAM|10|17|Когда донесли [об этом] Давиду, то он собрал всех Израильтян, и перешел Иордан и пришел к Еламу. Сирийцы выстроились против Давида и сразились с ним.
2SAM|10|18|И побежали Сирийцы от Израильтян. Давид истребил у Сирийцев семьсот колесниц и сорок тысяч всадников; поразил и военачальника Совака, который там и умер.
2SAM|10|19|Когда все цари покорные Адраазару увидели, что они поражены Израильтянами, то заключили мир с Израильтянами и покорились им. А Сирийцы боялись более помогать Аммонитянам.
2SAM|11|1|Через год, в то время, когда выходят цари [в походы], Давид послал Иоава и слуг своих с ним и всех Израильтян; и они поразили Аммонитян и осадили Равву; Давид же оставался в Иерусалиме.
2SAM|11|2|Однажды под вечер Давид, встав с постели, прогуливался на кровле царского дома и увидел с кровли купающуюся женщину; а та женщина была очень красива.
2SAM|11|3|И послал Давид разведать, кто эта женщина? И сказали ему: это Вирсавия, дочь Елиама, жена Урии Хеттеянина.
2SAM|11|4|Давид послал слуг взять ее; и она пришла к нему, и он спал с нею. Когда же она очистилась от нечистоты своей, возвратилась в дом свой.
2SAM|11|5|Женщина эта сделалась беременною и послала известить Давида, говоря: я беременна.
2SAM|11|6|И послал Давид [сказать] Иоаву: пришли ко мне Урию Хеттеянина. И послал Иоав Урию к Давиду.
2SAM|11|7|И пришел к нему Урия, и расспросил [его] Давид о положении Иоава и о положении народа, и о ходе войны.
2SAM|11|8|И сказал Давид Урии: иди домой и омой ноги свои. И вышел Урия из дома царского, а вслед за ним понесли и царское кушанье.
2SAM|11|9|Но Урия спал у ворот царского дома со всеми слугами своего господина, и не пошел в свой дом.
2SAM|11|10|И донесли Давиду, говоря: не пошел Урия в дом свой. И сказал Давид Урии: вот, ты пришел с дороги; отчего же не пошел ты в дом свой?
2SAM|11|11|И сказал Урия Давиду: ковчег и Израиль и Иуда находятся в шатрах, и господин мой Иоав и рабы господина моего пребывают в поле, а я вошел бы в дом свой и есть и пить и спать со своею женою! Клянусь твоею жизнью и жизнью души твоей, этого я не сделаю.
2SAM|11|12|И сказал Давид Урии: останься здесь и на этот день, а завтра я отпущу тебя. И остался Урия в Иерусалиме на этот день до завтра.
2SAM|11|13|И пригласил его Давид, и ел [Урия] пред ним и пил, и напоил его [Давид]. Но вечером [Урия] пошел спать на постель свою с рабами господина своего, а в свой дом не пошел.
2SAM|11|14|Поутру Давид написал письмо к Иоаву и послал [его] с Уриею.
2SAM|11|15|В письме он написал так: поставьте Урию там, где [будет] самое сильное сражение, и отступите от него, чтоб он был поражен и умер.
2SAM|11|16|Посему, когда Иоав осаждал город, то поставил он Урию на таком месте, о котором знал, что там храбрые люди.
2SAM|11|17|И вышли люди из города и сразились с Иоавом, и пало несколько из народа, из слуг Давидовых; был убит также и Урия Хеттеянин.
2SAM|11|18|И послал Иоав донести Давиду о всем ходе сражения.
2SAM|11|19|И приказал посланному, говоря: когда ты расскажешь царю о всем ходе сражения
2SAM|11|20|и увидишь, что царь разгневается, и скажет тебе: "зачем вы так близко подходили к городу сражаться? разве вы не знали, что со стены будут бросать на вас?
2SAM|11|21|кто убил Авимелеха, сына Иероваалова? не женщина ли бросила на него со стены обломок жернова, и он умер в Тевеце? Зачем же вы близко подходили к стене?" тогда ты скажи: и раб твой Урия Хеттеянин также умер.
2SAM|11|22|И пошел [посланный], и пришел, и рассказал Давиду обо всем, для чего послал его Иоав, обо всем ходе сражения.
2SAM|11|23|Тогда посланный сказал Давиду: одолевали нас те люди и вышли к нам в поле, и мы преследовали их до входа в ворота;
2SAM|11|24|тогда стреляли стрелки со стены на рабов твоих, и умерли [некоторые] из рабов царя; умер также и раб твой Урия Хеттеянин.
2SAM|11|25|Тогда сказал Давид посланному: так скажи Иоаву: "пусть не смущает тебя это дело, ибо меч поядает иногда того, иногда сего; усиль войну твою против города и разрушь его". Так ободри его.
2SAM|11|26|И услышала жена Урии, что умер Урия, муж ее, и плакала по муже своем.
2SAM|11|27|Когда кончилось время плача, Давид послал, и взял ее в дом свой, и она сделалась его женою и родила ему сына. И было это дело, которое сделал Давид, зло в очах Господа.
2SAM|12|1|И послал Господь Нафана к Давиду, и тот пришел к нему и сказал ему: в одном городе были два человека, один богатый, а другой бедный;
2SAM|12|2|у богатого было очень много мелкого и крупного скота,
2SAM|12|3|а у бедного ничего, кроме одной овечки, которую он купил маленькую и выкормил, и она выросла у него вместе с детьми его; от хлеба его она ела, и из его чаши пила, и на груди у него спала, и была для него, как дочь;
2SAM|12|4|и пришел к богатому человеку странник, и тот пожалел взять из своих овец или волов, чтобы приготовить [обед] для странника, который пришел к нему, а взял овечку бедняка и приготовил ее для человека, который пришел к нему.
2SAM|12|5|Сильно разгневался Давид на этого человека и сказал Нафану: жив Господь! достоин смерти человек, сделавший это;
2SAM|12|6|и за овечку он должен заплатить вчетверо, за то, что он сделал это, и за то, что не имел сострадания.
2SAM|12|7|И сказал Нафан Давиду: ты – тот человек. Так говорит Господь Бог Израилев: Я помазал тебя в царя над Израилем и Я избавил тебя от руки Саула,
2SAM|12|8|и дал тебе дом господина твоего и жен господина твоего на лоно твое, и дал тебе дом Израилев и Иудин, и, если этого [для тебя] мало, прибавил бы тебе еще больше;
2SAM|12|9|зачем же ты пренебрег слово Господа, сделав злое пред очами Его? Урию Хеттеянина ты поразил мечом; жену его взял себе в жену, а его ты убил мечом Аммонитян;
2SAM|12|10|итак не отступит меч от дома твоего во веки, за то, что ты пренебрег Меня и взял жену Урии Хеттеянина, чтоб она была тебе женою.
2SAM|12|11|Так говорит Господь: вот, Я воздвигну на тебя зло из дома твоего, и возьму жен твоих пред глазами твоими, и отдам ближнему твоему, и будет он спать с женами твоими пред этим солнцем;
2SAM|12|12|ты сделал тайно, а Я сделаю это пред всем Израилем и пред солнцем.
2SAM|12|13|И сказал Давид Нафану: согрешил я пред Господом. И сказал Нафан Давиду: и Господь снял [с тебя] грех твой; ты не умрешь;
2SAM|12|14|но как ты этим делом подал повод врагам Господа хулить Его, то умрет родившийся у тебя сын.
2SAM|12|15|И пошел Нафан в дом свой. И поразил Господь дитя, которое родила жена Урии Давиду, и оно заболело.
2SAM|12|16|И молился Давид Богу о младенце, и постился Давид, и, уединившись провел ночь, лежа на земле.
2SAM|12|17|И вошли к нему старейшины дома его, чтобы поднять его с земли; но он не хотел, и не ел с ними хлеба.
2SAM|12|18|На седьмой день дитя умерло, и слуги Давидовы боялись донести ему, что умер младенец; ибо, говорили они, когда дитя было еще живо, и мы уговаривали его, и он не слушал голоса нашего, как же мы скажем ему: "умерло дитя"? Он сделает что–нибудь худое.
2SAM|12|19|И увидел Давид, что слуги его перешептываются между собою, и понял Давид, что дитя умерло, и спросил Давид слуг своих: умерло дитя? И сказали: умерло.
2SAM|12|20|Тогда Давид встал с земли и умылся, и помазался, и переменил одежды свои, и пошел в дом Господень, и молился. Возвратившись домой, потребовал, чтобы подали ему хлеба, и он ел.
2SAM|12|21|И сказали ему слуги его: что значит, что ты так поступаешь: когда дитя было еще живо, ты постился и плакал; а когда дитя умерло, ты встал и ел хлеб?
2SAM|12|22|И сказал Давид: доколе дитя было живо, я постился и плакал, ибо думал: кто знает, не помилует ли меня Господь, и дитя останется живо?
2SAM|12|23|А теперь оно умерло; зачем же мне поститься? Разве я могу возвратить его? Я пойду к нему, а оно не возвратится ко мне.
2SAM|12|24|И утешил Давид Вирсавию, жену свою, и вошел к ней и спал с нею; и она родила сына, и нарекла ему имя: Соломон. И Господь возлюбил его
2SAM|12|25|и послал пророка Нафана, и он нарек ему имя: Иедидиа по слову Господа.
2SAM|12|26|Иоав воевал против Раввы Аммонитской и взял [почти] царственный город.
2SAM|12|27|И послал Иоав к Давиду сказать ему: я нападал на Равву и овладел водою города;
2SAM|12|28|теперь собери остальной народ и подступи к городу и возьми его; ибо, если я возьму его, то мое имя будет наречено ему.
2SAM|12|29|И собрал Давид весь народ и пошел к Равве, и воевал против нее и взял ее.
2SAM|12|30|И взял Давид венец царя их с головы его, – а в нем было золота талант и драгоценный камень, – и возложил его Давид на свою голову, и добычи из города вынес очень много.
2SAM|12|31|А народ, бывший в нем, он вывел и положил их под пилы, под железные молотилки, под железные топоры, и бросил их в обжигательные печи. Так он поступил со всеми городами Аммонитскими. И возвратился после того Давид и весь народ в Иерусалим.
2SAM|13|1|И было после того: у Авессалома, сына Давидова, [была] сестра красивая, по имени Фамарь, и полюбил ее Амнон, сын Давида.
2SAM|13|2|И скорбел Амнон до того, что заболел из–за Фамари, сестры своей; ибо она была девица, и Амнону казалось трудным что–нибудь сделать с нею.
2SAM|13|3|Но у Амнона был друг, по имени Ионадав, сын Самая, брата Давидова; и Ионадав был человек очень хитрый.
2SAM|13|4|И он сказал ему: отчего ты так худеешь с каждым днем, сын царев, – не откроешь ли мне? И сказал ему Амнон: Фамарь, сестру Авессалома, брата моего, люблю я.
2SAM|13|5|И сказал ему Ионадав: ложись в постель твою, и притворись больным; и когда отец твой придет навестить тебя: скажи ему: пусть придет Фамарь, сестра моя, и подкрепит меня пищею, приготовив кушанье при моих глазах, чтоб я видел, и ел из рук ее.
2SAM|13|6|И лег Амнон и притворился больным, и пришел царь навестить его; и сказал Амнон царю: пусть придет Фамарь, сестра моя, и испечет при моих глазах лепешку, или две, и я поем из рук ее.
2SAM|13|7|И послал Давид к Фамари в дом сказать: пойди в дом Амнона, брата твоего, и приготовь ему кушанье.
2SAM|13|8|И пошла она в дом брата своего Амнона; а он лежит. И взяла она муки и замесила, и изготовила пред глазами его и испекла лепешки,
2SAM|13|9|и взяла сковороду и выложила пред ним; но он не хотел есть. И сказал Амнон: пусть все выйдут от меня. И вышли от него все люди,
2SAM|13|10|и сказал Амнон Фамари: отнеси кушанье во внутреннюю комнату, и я поем из рук твоих. И взяла Фамарь лепешки, которые приготовила, и отнесла Амнону, брату своему, во внутреннюю комнату.
2SAM|13|11|И когда она поставила пред ним, чтоб он ел, то он схватил ее, и сказал ей: иди, ложись со мною, сестра моя.
2SAM|13|12|Но она сказала: нет, брат мой, не бесчести меня, ибо не делается так в Израиле; не делай этого безумия.
2SAM|13|13|И я, куда пойду я с моим бесчестием? И ты, ты будешь одним из безумных в Израиле. Ты поговори с царем; он не откажет отдать меня тебе.
2SAM|13|14|Но он не хотел слушать слов ее, и преодолел ее, и изнасиловал ее, и лежал с нею.
2SAM|13|15|Потом возненавидел ее Амнон величайшею ненавистью, так что ненависть, какою он возненавидел ее, была сильнее любви, какую имел к ней; и сказал ей Амнон: встань, уйди.
2SAM|13|16|И [Фамарь] сказала ему: нет, прогнать меня – это зло больше первого, которое ты сделал со мною. Но он не хотел слушать ее.
2SAM|13|17|И позвал отрока своего, который служил ему, и сказал: прогони эту от меня вон и запри дверь за нею.
2SAM|13|18|На ней была разноцветная одежда, ибо такие верхние одежды носили царские дочери–девицы. И вывел ее слуга вон и запер за нею дверь.
2SAM|13|19|И посыпала Фамарь пеплом голову свою, и разодрала разноцветную одежду, которую имела на себе, и положила руки свои на голову свою, и так шла и вопила.
2SAM|13|20|И сказал ей Авессалом, брат ее: не Амнон ли, брат твой, был с тобою? – но теперь молчи, сестра моя; он – брат твой; не сокрушайся сердцем твоим об этом деле. И жила Фамарь в одиночестве в доме Авессалома, брата своего.
2SAM|13|21|И услышал царь Давид обо всем этом, и сильно разгневался.
2SAM|13|22|Авессалом же не говорил с Амноном ни худого, ни хорошего; ибо возненавидел Авессалом Амнона за то, что он обесчестил Фамарь, сестру его.
2SAM|13|23|Чрез два года было стрижение [овец] у Авессалома в Ваал – Гацоре, что у Ефрема, и позвал Авессалом всех сыновей царских.
2SAM|13|24|И пришел Авессалом к царю и сказал: вот, ныне стрижение [овец] у раба твоего; пусть пойдет царь и слуги его с рабом твоим.
2SAM|13|25|Но царь сказал Авессалому: нет, сын мой, мы не пойдем все, чтобы не быть тебе в тягость. И сильно упрашивал его [Авессалом]; но он не захотел идти, и благословил его.
2SAM|13|26|И сказал ему Авессалом: по крайней мере пусть пойдет с нами Амнон, брат мой. И сказал ему царь: зачем ему идти с тобою?
2SAM|13|27|Но Авессалом упросил его, и он отпустил с ним Амнона и всех царских сыновей.
2SAM|13|28|Авессалом же приказал отрокам своим, сказав: смотрите, как только развеселится сердце Амнона от вина, и я скажу вам: "поразите Амнона", тогда убейте его, не бойтесь; это я приказываю вам, будьте смелы и мужественны.
2SAM|13|29|И поступили отроки Авессалома с Амноном, как приказал Авессалом. Тогда встали все царские сыновья, сели каждый на мула своего и убежали.
2SAM|13|30|Когда они были еще на пути, дошел слух до Давида, что Авессалом умертвил всех царских сыновей, и не осталось ни одного из них.
2SAM|13|31|И встал царь, и разодрал одежды свои, и повергся на землю, и все слуги его, предстоящие ему, разодрали одежды свои.
2SAM|13|32|Но Ионадав, сын Самая, брата Давидова, сказал: пусть не думает господин мой, что всех отроков, царских сыновей, умертвили; один только Амнон умер, ибо у Авессалома был этот замысел с того дня, как [Амнон] обесчестил сестру его;
2SAM|13|33|итак пусть господин мой, царь, не тревожится мыслью о том, будто умерли все царские сыновья: умер один только Амнон.
2SAM|13|34|И убежал Авессалом. И поднял отрок, стоявший на страже, глаза свои, и увидел: вот, много народа идет по дороге по скату горы.
2SAM|13|35|Тогда Ионадав сказал царю: это идут царские сыновья; как говорил раб твой, так и есть.
2SAM|13|36|И едва только сказал он это, вот пришли царские сыновья, и подняли вопль и плакали. И сам царь и все слуги его плакали очень великим плачем.
2SAM|13|37|Авессалом же убежал и пошел к Фалмаю, сыну Емиуда, царю Гессурскому. И плакал Давид о сыне своем во все дни.
2SAM|13|38|Авессалом убежал и пришел в Гессур и пробыл там три года.
2SAM|13|39|И не стал царь Давид преследовать Авессалома; ибо утешился о смерти Амнона.
2SAM|14|1|И заметил Иоав, сын Саруи, что сердце царя обратилось к Авессалому.
2SAM|14|2|И послал Иоав в Фекою, и взял оттуда умную женщину и сказал ей: притворись плачущею и надень печальную одежду, и не мажься елеем, и представься женщиною, много дней плакавшею по умершем;
2SAM|14|3|и пойди к царю и скажи ему так и так. И вложил Иоав в уста ее, что сказать.
2SAM|14|4|И вошла женщина Фекоитянка к царю и пала лицем своим на землю, и поклонилась и сказала: помоги, царь!
2SAM|14|5|И сказал ей царь: что тебе? И сказала она: я вдова, муж мой умер;
2SAM|14|6|и у рабы твоей [было] два сына; они поссорились в поле, и некому было разнять их, и поразил один другого и умертвил его.
2SAM|14|7|И вот, восстало все родство на рабу твою, и говорят: "отдай убийцу брата своего; мы убьем его за душу брата его, которую он погубил, и истребим даже наследника". И так они погасят остальную искру мою, чтобы не оставить мужу моему имени и потомства на лице земли.
2SAM|14|8|И сказал царь женщине: иди спокойно домой, я дам приказание о тебе.
2SAM|14|9|Но женщина Фекоитянка сказала царю: на мне, господин мой царь, да будет вина и на доме отца моего, царь же и престол его неповинен.
2SAM|14|10|И сказал царь: того, кто будет против тебя, приведи ко мне, и он более не тронет тебя.
2SAM|14|11|Она сказала: помяни, царь, Господа Бога твоего, чтобы не умножились мстители за кровь и не погубили сына моего. И сказал [царь]: жив Господь! не падет и волос сына твоего на землю.
2SAM|14|12|И сказала женщина: позволь рабе твоей сказать [еще] слово господину моему царю.
2SAM|14|13|Он сказал: говори. И сказала женщина: почему ты так мыслишь против народа Божия? Царь, произнеся это слово, обвинил себя самого, потому что не возвращает изгнанника своего.
2SAM|14|14|Мы умрем и [будем] как вода, вылитая на землю, которую нельзя собрать; но Бог не желает погубить душу и помышляет, как бы не отвергнуть от Себя и отверженного.
2SAM|14|15|И теперь я пришла сказать царю, господину моему, эти слова, потому что народ пугает меня; и раба твоя сказала: поговорю я с царем, не сделает ли он по слову рабы своей;
2SAM|14|16|верно царь выслушает и избавит рабу свою от руки людей, [хотящих] истребить меня вместе с сыном моим из наследия Божия.
2SAM|14|17|И сказала раба твоя: да будет слово господина моего царя в утешение мне, ибо господин мой царь, как Ангел Божий, и может выслушать и доброе и худое. И Господь Бог твой будет с тобою.
2SAM|14|18|И отвечал царь и сказал женщине: не скрой от меня, о чем я спрошу тебя. И сказала женщина: говори, господин мой царь.
2SAM|14|19|И сказал царь: не рука ли Иоава во всем этом с тобою? И отвечала женщина и сказала: да живет душа твоя, господин мой царь; ни направо, ни налево нельзя уклониться от того, что сказал господин мой, царь; точно, раб твой Иоав приказал мне, и он вложил в уста рабы твоей все эти слова;
2SAM|14|20|чтобы притчею дать делу такой вид, раб твой Иоав научил меня; но господин мой мудр, как мудр Ангел Божий, чтобы знать все, что на земле.
2SAM|14|21|И сказал царь Иоаву: вот, я сделал [по слову твоему]; пойди же, возврати отрока Авессалома.
2SAM|14|22|Тогда Иоав пал лицем на землю и поклонился, и благословил царя и сказал: теперь знает раб твой, что обрел благоволение пред очами твоими, господин мой царь, так как царь сделал по слову раба своего.
2SAM|14|23|И встал Иоав, и пошел в Гессур, и привел Авессалома в Иерусалим.
2SAM|14|24|И сказал царь: пусть он возвратится в дом свой, а лица моего не видит. И пошел Авессалом в свой дом, а лица царского не видал.
2SAM|14|25|Не было во всем Израиле мужчины столь красивого, как Авессалом, и столько хвалимого, как он; от подошвы ног до верха головы его не было у него недостатка.
2SAM|14|26|Когда он стриг голову свою, – а он стриг ее каждый год, потому что она отягощала его, – то волоса с головы его весили двести сиклей по весу царскому.
2SAM|14|27|И родились у Авессалома три сына и одна дочь, по имени Фамарь; она была женщина красивая.
2SAM|14|28|И оставался Авессалом в Иерусалиме два года, а лица царского не видал.
2SAM|14|29|И послал Авессалом за Иоавом, чтобы послать его к царю, но тот не захотел придти к нему. Послал и в другой раз; но тот не захотел придти.
2SAM|14|30|И сказал [Авессалом] слугам своим: видите участок поля Иоава подле моего, и у него там ячмень; пойдите, выжгите его огнем. И выжгли слуги Авессалома тот участок поля огнем.
2SAM|14|31|И встал Иоав, и пришел к Авессалому в дом, и сказал ему: зачем слуги твои выжгли мой участок огнем?
2SAM|14|32|И сказал Авессалом Иоаву: вот, я посылал за тобою, говоря: приди сюда, и я пошлю тебя к царю сказать: зачем я пришел из Гессура? Лучше было бы мне оставаться там. Я хочу увидеть лице царя. Если же я виноват, то убей меня.
2SAM|14|33|И пошел Иоав к царю и пересказал ему [это]. И позвал [царь] Авессалома; он пришел к царю, и пал лицем своим на землю пред царем; и поцеловал царь Авессалома.
2SAM|15|1|После сего Авессалом завел у себя колесницы и лошадей и пятьдесят скороходов.
2SAM|15|2|И вставал Авессалом рано утром, и становился при дороге у ворот, и когда кто–нибудь, имея тяжбу, шел к царю на суд, то Авессалом подзывал его к себе и спрашивал: из какого города ты? И когда тот отвечал: из такого–то колена Израилева раб твой,
2SAM|15|3|тогда говорил ему Авессалом: вот, дело твое доброе и справедливое, но у царя некому выслушать тебя.
2SAM|15|4|И говорил Авессалом: о, если бы меня поставили судьею в этой земле! ко мне приходил бы всякий, кто имеет спор и тяжбу, и я судил бы его по правде.
2SAM|15|5|И когда подходил кто–нибудь поклониться ему, то он простирал руку свою и обнимал его и целовал его.
2SAM|15|6|Так поступал Авессалом со всяким Израильтянином, приходившим на суд к царю, и вкрадывался Авессалом в сердце Израильтян.
2SAM|15|7|По прошествии сорока лет [царствования Давида], Авессалом сказал царю: пойду я и исполню обет мой, который я дал Господу, в Хевроне;
2SAM|15|8|ибо я, раб твой, живя в Гессуре в Сирии, дал обет: если Господь возвратит меня в Иерусалим, то я принесу жертву Господу.
2SAM|15|9|И сказал ему царь: иди с миром. И встал он и пошел в Хеврон.
2SAM|15|10|И разослал Авессалом лазутчиков во все колена Израилевы, сказав: когда вы услышите звук трубы, то говорите: Авессалом воцарился в Хевроне.
2SAM|15|11|С Авессаломом пошли из Иерусалима двести человек, которые были приглашены им, и пошли по простоте своей, не зная, в чем дело.
2SAM|15|12|Во время жертвоприношения Авессалом послал и призвал Ахитофела Гилонянина, советника Давидова, из его города Гило. И составился сильный заговор, и народ стекался и умножался около Авессалома.
2SAM|15|13|И пришел вестник к Давиду и сказал: сердце Израильтян уклонилось на сторону Авессалома.
2SAM|15|14|И сказал Давид всем слугам своим, которые были при нем в Иерусалиме: встаньте, убежим, ибо не будет нам спасения от Авессалома; спешите, чтобы нам уйти, чтоб он не застиг и не захватил нас, и не навел на нас беды и не истребил города мечом.
2SAM|15|15|И сказали слуги царские царю: во всем, что угодно господину нашему царю, мы – рабы твои.
2SAM|15|16|И вышел царь и весь дом его за ним пешком. Оставил же царь десять жен, наложниц [своих], для хранения дома.
2SAM|15|17|И вышел царь и весь народ пешие, и остановились у Беф–Мерхата.
2SAM|15|18|И все слуги его шли по сторонам его, и все Хелефеи, и все Фелефеи, и все Гефяне до шестисот человек, пришедшие вместе с ним из Гефа, шли впереди царя.
2SAM|15|19|И сказал царь Еффею Гефянину: зачем и ты идешь с нами? Возвратись и оставайся с тем царем; ибо ты – чужеземец и пришел сюда из своего места;
2SAM|15|20|вчера ты пришел, а сегодня я заставлю тебя идти с нами? Я иду, куда случится; возвратись и возврати братьев своих с собою; милость и истину [с тобою]!
2SAM|15|21|И отвечал Еффей царю и сказал: жив Господь, и да живет господин мой царь: где бы ни был господин мой царь, в жизни ли, в смерти ли, там будет и раб твой.
2SAM|15|22|И сказал Давид Еффею: итак иди и ходи со мною. И пошел Еффей Гефянин и все люди его и все дети, бывшие с ним.
2SAM|15|23|И плакала вся земля громким голосом. И весь народ переходил, и царь перешел поток Кедрон; и пошел весь народ по дороге к пустыне.
2SAM|15|24|Вот и Садок, и все левиты с ним несли ковчег завета Божия из Вефары и поставили ковчег Божий; Авиафар же стоял на возвышении, доколе весь народ не вышел из города.
2SAM|15|25|И сказал царь Садоку: возврати ковчег Божий в город. Если я обрету милость пред очами Господа, то Он возвратит меня и даст мне видеть его и жилище его.
2SAM|15|26|А если Он скажет так: "нет Моего благоволения к тебе", то вот я; пусть творит со мною, что Ему благоугодно.
2SAM|15|27|И сказал царь Садоку священнику: видишь ли, – возвратись в город с миром, и Ахимаас, сын твой, и Ионафан, сын Авиафара, оба сына ваши с вами;
2SAM|15|28|видите ли, я помедлю на равнине в пустыне, доколе не придет известие от вас ко мне.
2SAM|15|29|И возвратили Садок и Авиафар ковчег Божий в Иерусалим, и остались там.
2SAM|15|30|А Давид пошел на гору Елеонскую, шел и плакал; голова у него была покрыта; он шел босой, и все люди, бывшие с ним, покрыли каждый голову свою, шли и плакали.
2SAM|15|31|Донесли Давиду и сказали: и Ахитофел в числе заговорщиков с Авессаломом. И сказал Давид: Господи! разрушь совет Ахитофела.
2SAM|15|32|Когда Давид взошел на вершину горы, где он поклонялся Богу, вот навстречу ему идет Хусий Архитянин, друг Давидов; одежда на нем была разодрана, и прах на голове его.
2SAM|15|33|И сказал ему Давид: если ты пойдешь со мною, то будешь мне в тягость;
2SAM|15|34|но если возвратишься в город и скажешь Авессалому: "царь, я раб твой; доселе я был рабом отца твоего, а теперь я – твой раб": то ты расстроишь для меня совет Ахитофела.
2SAM|15|35|Вот, там с тобою Садок и Авиафар священники, и всякое слово, какое услышишь из дома царя, пересказывай Садоку и Авиафару священникам.
2SAM|15|36|Там с ними и два сына их, Ахимаас, сын Садока, и Ионафан, сын Авиафара; чрез них посылайте ко мне всякое известие, какое услышите.
2SAM|15|37|И пришел Хусий, друг Давида, в город; Авессалом же вступал тогда в Иерусалим.
2SAM|16|1|Когда Давид немного сошел с вершины горы, вот встречается ему Сива, слуга Мемфивосфея, с парою навьюченных ослов, и на них двести хлебов, сто связок изюму, сто связок смокв и мех с вином.
2SAM|16|2|И сказал царь Сиве: для чего это у тебя? И отвечал Сива: ослы для дома царского, для езды, а хлеб и плоды для пищи отрокам, а вино для питья ослабевшим в пустыне.
2SAM|16|3|И сказал царь: где сын господина твоего? И отвечал Сива царю: вот, он остался в Иерусалиме и говорит: теперь–то дом Израилев возвратит мне царство отца моего.
2SAM|16|4|И сказал царь Сиве: вот тебе все, что у Мемфивосфея. И отвечал Сива, поклонившись: да обрету милость в глазах господина моего царя!
2SAM|16|5|Когда дошел царь Давид до Бахурима, вот вышел оттуда человек из рода дома Саулова, по имени Семей, сын Геры; он шел и злословил,
2SAM|16|6|и бросал камнями на Давида и на всех рабов царя Давида; все же люди и все храбрые были по правую и по левую сторону [царя].
2SAM|16|7|Так говорил Семей, злословя его: уходи, уходи, убийца и беззаконник!
2SAM|16|8|Господь обратил на тебя всю кровь дома Саулова, вместо которого ты воцарился, и предал Господь царство в руки Авессалома, сына твоего; и вот, ты в беде, ибо ты – кровопийца.
2SAM|16|9|И сказал Авесса, сын Саруин, царю: зачем злословит этот мертвый пес господина моего царя? пойду я и сниму с него голову.
2SAM|16|10|И сказал царь: что мне и вам, сыны Саруины? пусть он злословит, ибо Господь повелел ему злословить Давида. Кто же может сказать: зачем ты так делаешь?
2SAM|16|11|И сказал Давид Авессе и всем слугам своим: вот, если мой сын, который вышел из чресл моих, ищет души моей, тем больше сын Вениамитянина; оставьте его, пусть злословит, ибо Господь повелел ему;
2SAM|16|12|может быть, Господь призрит на уничижение мое, и воздаст мне Господь благостью за теперешнее его злословие.
2SAM|16|13|И шел Давид и люди его [своим] путем, а Семей шел по окраине горы, со стороны его, шел и злословил, и бросал камнями на сторону его и пылью.
2SAM|16|14|И пришел царь и весь народ, бывший с ним, утомленный, и отдыхал там.
2SAM|16|15|Авессалом же и весь народ Израильский пришли в Иерусалим, и Ахитофел с ним.
2SAM|16|16|Когда Хусий Архитянин, друг Давидов, пришел к Авессалому, то сказал Хусий Авессалому: да живет царь, да живет царь!
2SAM|16|17|И сказал Авессалом Хусию: таково–то усердие твое к твоему другу! отчего ты не пошел с другом твоим?
2SAM|16|18|И сказал Хусий Авессалому: нет, кого избрал Господь и этот народ и весь Израиль, с тем и я, и с ним останусь.
2SAM|16|19|И притом кому я буду служить? Не сыну ли его? Как служил я отцу твоему, так буду служить и тебе.
2SAM|16|20|И сказал Авессалом Ахитофелу: дайте совет, что нам делать.
2SAM|16|21|И сказал Ахитофел Авессалому: войди к наложницам отца твоего, которых он оставил охранять дом свой; и услышат все Израильтяне, что ты сделался ненавистным для отца твоего, и укрепятся руки всех, которые с тобою.
2SAM|16|22|И поставили для Авессалома палатку на кровле, и вошел Авессалом к наложницам отца своего пред глазами всего Израиля.
2SAM|16|23|Советы же Ахитофела, которые он давал, в то время [считались], как если бы кто спрашивал наставления у Бога. Таков был всякий совет Ахитофела как для Давида, так и для Авессалома.
2SAM|17|1|И сказал Ахитофел Авессалому: выберу я двенадцать тысяч человек и встану и пойду в погоню за Давидом в эту ночь;
2SAM|17|2|и нападу на него, когда он будет утомлен и с опущенными руками, и приведу его в страх; и все люди, которые с ним, разбегутся; и я убью одного царя
2SAM|17|3|и всех людей обращу к тебе; и когда не будет одного, душу которого ты ищешь, тогда весь народ будет в мире.
2SAM|17|4|И понравилось это слово Авессалому и всем старейшинам Израилевым.
2SAM|17|5|И сказал Авессалом: позовите Хусия Архитянина; послушаем, что он скажет.
2SAM|17|6|И пришел Хусий к Авессалому, и сказал ему Авессалом, говоря: вот что говорит Ахитофел; сделать ли по его словам? а если нет, то говори ты.
2SAM|17|7|И сказал Хусий Авессалому: нехорош на этот раз совет, который дал Ахитофел.
2SAM|17|8|И продолжал Хусий: ты знаешь твоего отца и людей его; они храбры и сильно раздражены, как медведица в поле, у которой отняли детей, и отец твой – человек воинственный; он не остановится ночевать с народом.
2SAM|17|9|Вот, теперь он скрывается в какой–нибудь пещере, или в другом месте, и если кто падет при первом нападении на них, и услышат и скажут: "было поражение людей, последовавших за Авессаломом",
2SAM|17|10|тогда и самый храбрый, у которого сердце, как сердце львиное, упадет духом; ибо всему Израилю известно, как храбр отец твой и мужественны те, которые с ним.
2SAM|17|11|Посему я советую: пусть соберется к тебе весь Израиль, от Дана до Вирсавии, во множестве, как песок при море, и ты сам пойдешь посреди его;
2SAM|17|12|и тогда мы пойдем против него, в каком бы месте он ни находился, и нападем на него, как падает роса на землю; и не останется у него ни одного человека из всех, которые с ним;
2SAM|17|13|а если он войдет в какой–либо город, то весь Израиль принесет к тому городу веревки, и мы стащим его в реку, так что не останется ни одного камешка.
2SAM|17|14|И сказал Авессалом и весь Израиль: совет Хусия Архитянина лучше совета Ахитофелова. Так Господь судил разрушить лучший совет Ахитофела, чтобы навести Господу бедствие на Авессалома.
2SAM|17|15|И сказал Хусий Садоку и Авиафару священникам: так и так советовал Ахитофел Авессалому и старейшинам Израилевым, а так и так посоветовал я.
2SAM|17|16|И теперь пошлите поскорее и скажите Давиду так: не оставайся в эту ночь на равнине в пустыне, но поскорее перейди, чтобы не погибнуть царю и всем людям, которые с ним.
2SAM|17|17|Ионафан и Ахимаас стояли у источника Рогель. И пошла служанка и рассказала им, а они пошли и известили царя Давида; ибо они не могли показаться в городе.
2SAM|17|18|И увидел их отрок и донес Авессалому; но они оба скоро ушли и пришли в Бахурим, в дом одного человека, у которого на дворе был колодезь, и спустились туда.
2SAM|17|19|А женщина взяла и растянула над устьем колодезя покрывало и насыпала на него крупы, так что не было ничего заметно.
2SAM|17|20|И пришли рабы Авессалома к женщине в дом, и сказали: где Ахимаас и Ионафан? И сказала им женщина: они перешли вброд реку. И искали они, и не нашли, и возвратились в Иерусалим.
2SAM|17|21|Когда они ушли, те вышли из колодезя, пошли и известили царя Давида и сказали Давиду: встаньте и поскорее перейдите воду; ибо так и так советовал о вас Ахитофел.
2SAM|17|22|И встал Давид и все люди, бывшие с ним, и перешли Иордан; к рассвету не осталось ни одного, который не перешел бы Иордана.
2SAM|17|23|И увидел Ахитофел, что не исполнен совет его, и оседлал осла, и собрался, и пошел в дом свой, в город свой, и сделал завещание дому своему, и удавился, и умер, и был погребен в гробе отца своего.
2SAM|17|24|И пришел Давид в Маханаим, а Авессалом перешел Иордан, сам и весь Израиль с ним.
2SAM|17|25|Авессалом поставил Амессая, вместо Иоава, над войском. Амессай был сын одного человека, по имени Иефера из Изрееля, который вошел к Авигее, дочери Нааса, сестре Саруи, матери Иоава.
2SAM|17|26|И Израиль с Авессаломом расположился станом в земле Галаадской.
2SAM|17|27|Когда Давид пришел в Маханаим, то Сови, сын Нааса, из Раввы Аммонитской, и Махир, сын Аммиила, из Лодавара, и Верзеллий Галаадитянин из Роглима,
2SAM|17|28|принесли постелей, блюд и глиняных сосудов, и пшеницы, и ячменя, и муки, и пшена, и бобов, и чечевицы, и жареных зерен,
2SAM|17|29|и меду, и масла, и овец, и сыра коровьего, принесли Давиду и людям, бывшим с ним, в пищу; ибо говорили они: народ голоден и утомлен и терпел жажду в пустыне.
2SAM|18|1|И осмотрел Давид людей, бывших с ним, и поставил над ними тысяченачальников и сотников.
2SAM|18|2|И отправил Давид людей – третью часть под предводительством Иоава, третью часть под предводительством Авессы, сына Саруина, брата Иоава, третью часть под предводительством Еффея Гефянина. И сказал царь людям: я сам пойду с вами.
2SAM|18|3|Но люди отвечали ему: не ходи; ибо, если мы и побежим, то не обратят внимания на это; если и умрет половина из нас, также не обратят внимания; а ты один то же, что нас десять тысяч; итак для нас лучше, чтобы ты помогал нам из города.
2SAM|18|4|И сказал им царь: что угодно в глазах ваших, то и сделаю. И стал царь у ворот, и весь народ выходил по сотням и по тысячам.
2SAM|18|5|И приказал царь Иоаву и Авессе и Еффею, говоря: сберегите мне отрока Авессалома. И все люди слышали, как приказывал царь всем начальникам об Авессаломе.
2SAM|18|6|И вышли люди в поле навстречу Израильтянам, и было сражение в лесу Ефремовом.
2SAM|18|7|И был поражен народ Израильский рабами Давида; было там поражение великое в тот день, – поражены двадцать тысяч [человек].
2SAM|18|8|Сражение распространилось по всей той стране, и лес погубил народа больше, чем сколько истребил меч, в тот день.
2SAM|18|9|И встретился Авессалом с рабами Давидовыми; он был на муле. Когда мул вбежал с ним под ветви большого дуба, то [Авессалом] запутался волосами своими в ветвях дуба и повис между небом и землею, а мул, бывший под ним, убежал.
2SAM|18|10|И увидел это некто и донес Иоаву, говоря: вот, я видел Авессалома висящим на дубе.
2SAM|18|11|И сказал Иоав человеку, донесшему об этом: вот, ты видел; зачем же ты не поверг его там на землю? я дал бы тебе десять сиклей серебра и один пояс.
2SAM|18|12|И отвечал тот Иоаву: если бы положили на руки мои и тысячу сиклей серебра, и тогда я не поднял бы руки на царского сына; ибо вслух нас царь приказывал тебе и Авессе и Еффею, говоря: "сберегите мне отрока Авессалома";
2SAM|18|13|и если бы я поступил иначе с опасностью жизни моей, то это не скрылось бы от царя, и ты же восстал бы против меня.
2SAM|18|14|Иоав сказал: нечего мне медлить с тобою. И взял в руки три стрелы и вонзил их в сердце Авессалома, который был еще жив на дубе.
2SAM|18|15|И окружили Авессалома десять отроков, оруженосцев Иоава, и поразили и умертвили его.
2SAM|18|16|И затрубил Иоав трубою, и возвратились люди из погони за Израилем, ибо Иоав щадил народ.
2SAM|18|17|И взяли Авессалома, и бросили его в лесу в глубокую яму, и наметали над ним огромную кучу камней. И все Израильтяне разбежались, каждый в шатер свой.
2SAM|18|18|Авессалом еще при жизни своей взял и поставил себе памятник в царской долине; ибо сказал он: нет у меня сына, чтобы сохранилась память имени моего. И назвал памятник своим именем. И называется он "памятник Авессалома" до сего дня.
2SAM|18|19|Ахимаас, сын Садоков, сказал Иоаву: побегу я, извещу царя, что Господь судом Своим избавил его от рук врагов его.
2SAM|18|20|Но Иоав сказал ему: не будешь ты сегодня добрым вестником; известишь в другой день, а не сегодня, ибо умер сын царя.
2SAM|18|21|И сказал Иоав Хусию: пойди, донеси царю, что видел ты. И поклонился Хусий Иоаву и побежал.
2SAM|18|22|Но Ахимаас, сын Садоков, настаивал и говорил Иоаву: что бы ни было, но и я побегу за Хусием. Иоав же отвечал: зачем бежать тебе, сын мой? не принесешь ты доброй вести.
2SAM|18|23|[И сказал Ахимаас]: пусть так, но я побегу. И сказал ему [Иоав]: беги. И побежал Ахимаас по прямой дороге и опередил Хусия.
2SAM|18|24|Давид тогда сидел между двумя воротами. И сторож взошел на кровлю ворот к стене и, подняв глаза, увидел: вот, бежит один человек.
2SAM|18|25|И закричал сторож и известил царя. И сказал царь: если один, то весть в устах его. А тот подходил все ближе и ближе.
2SAM|18|26|Сторож увидел и другого бегущего человека; и закричал сторож привратнику: вот, еще бежит один человек. Царь сказал: и это – вестник.
2SAM|18|27|Сторож сказал: я вижу походку первого, похожую на походку Ахимааса, сына Садокова. И сказал царь: это человек хороший и идет с хорошею вестью.
2SAM|18|28|И воскликнул Ахимаас и сказал царю: мир. И поклонился царю лицем своим до земли и сказал: благословен Господь Бог твой, предавший людей, которые подняли руки свои на господина моего царя!
2SAM|18|29|И сказал царь: благополучен ли отрок Авессалом? И сказал Ахимаас: я видел большое волнение, когда раб царев Иоав посылал раба твоего; но я не знаю, что [там] было.
2SAM|18|30|И сказал царь: отойди, стань здесь. Он отошел и стал.
2SAM|18|31|Вот, пришел и Хусий. И сказал Хусий: добрая весть господину моему царю! Господь явил тебе ныне правду в избавлении от руки всех восставших против тебя.
2SAM|18|32|И сказал царь Хусию: благополучен ли отрок Авессалом? И сказал Хусий: да будет с врагами господина моего царя и со всеми, злоумышляющими против тебя то же, что постигло отрока!
2SAM|19|1|И смутился царь, и пошел в горницу над воротами, и плакал, и когда шел, говорил так: сын мой Авессалом! сын мой, сын мой Авессалом! о, кто дал бы мне умереть вместо тебя, Авессалом, сын мой, сын мой!
2SAM|19|2|И сказали Иоаву: вот, царь плачет и рыдает об Авессаломе.
2SAM|19|3|И обратилась победа того дня в плач для всего народа; ибо народ услышал в тот день и говорил, что царь скорбит о своем сыне.
2SAM|19|4|И входил тогда народ в город украдкою, как крадутся люди стыдящиеся, которые во время сражения обратились в бегство.
2SAM|19|5|А царь закрыл лице свое и громко взывал: сын мой Авессалом! Авессалом, сын мой, сын мой!
2SAM|19|6|И пришел Иоав к царю в дом и сказал: ты в стыд привел сегодня всех слуг твоих, спасших ныне жизнь твою и жизнь сыновей и дочерей твоих, и жизнь жен и жизнь наложниц твоих;
2SAM|19|7|ты любишь ненавидящих тебя и ненавидишь любящих тебя, ибо ты показал сегодня, что ничто для тебя и вожди и слуги; сегодня я узнал, что если бы Авессалом остался жив, а мы все умерли, то тебе было бы приятнее;
2SAM|19|8|итак встань, выйди и поговори к сердцу рабов твоих, ибо клянусь Господом, что, если ты не выйдешь, в эту ночь не останется у тебя ни одного человека; и это будет для тебя хуже всех бедствий, какие находили на тебя от юности твоей доныне.
2SAM|19|9|И встал царь и сел у ворот, а всему народу возвестили, что царь сидит у ворот. И пришел весь народ пред лице царя; Израильтяне же разбежались по своим шатрам.
2SAM|19|10|И весь народ во всех коленах Израилевых спорил и говорил: царь избавил нас от рук врагов наших и освободил нас от рук Филистимлян, а теперь сам бежал из земли сей, от Авессалома.
2SAM|19|11|Но Авессалом, которого мы помазали [в царя] над нами, умер на войне; почему же теперь вы медлите возвратить царя?
2SAM|19|12|И царь Давид послал сказать священникам Садоку и Авиафару: скажите старейшинам Иудиным: зачем хотите вы быть последними, чтобы возвратить царя в дом его, тогда как слова всего Израиля дошли до царя в дом его?
2SAM|19|13|Вы братья мои, кости мои и плоть моя – вы; зачем хотите вы быть последними в возвращении царя в дом его?
2SAM|19|14|И Амессаю скажите: не кость ли моя и плоть моя – ты? Пусть то и то сделает со мною Бог и еще больше сделает, если ты не будешь военачальником при мне, вместо Иоава, навсегда!
2SAM|19|15|И склонил он сердце всех Иудеев, как одного человека; и послали они к царю [сказать]: возвратись ты и все слуги твои.
2SAM|19|16|И возвратился царь, и пришел к Иордану, а Иудеи пришли в Галгал, чтобы встретить царя и перевезти царя чрез Иордан.
2SAM|19|17|И поспешил Семей, сын Геры, Вениамитянин из Бахурима, и пошел с Иудеями навстречу царю Давиду,
2SAM|19|18|и тысяча человек из Вениамитян с ним, и Сива, слуга дома Саулова, с пятнадцатью сыновьями своими и двадцатью рабами своими; и перешли они Иордан пред лицем царя.
2SAM|19|19|Когда переправили судно, чтобы перевезти дом царя и послужить ему, тогда Семей, сын Геры, пал пред царем, как только он перешел Иордан,
2SAM|19|20|и сказал царю: не поставь мне, господин мой, в преступление, и не помяни того, чем согрешил раб твой в тот день, когда господин мой царь выходил из Иерусалима, и не держи [того], царь, на сердце своем;
2SAM|19|21|ибо знает раб твой, что согрешил, и вот, ныне я пришел первый из всего дома Иосифова, чтобы выйти навстречу господину моему царю.
2SAM|19|22|И отвечал Авесса, сын Саруин, и сказал: неужели Семей не умрет за то, что злословил помазанника Господня?
2SAM|19|23|И сказал Давид: что мне и вам, сыны Саруины, что вы делаетесь ныне мне наветниками? Ныне ли умерщвлять кого–либо в Израиле? Не вижу ли я, что ныне я – царь над Израилем?
2SAM|19|24|И сказал царь Семею: ты не умрешь. И поклялся ему царь.
2SAM|19|25|И Мемфивосфей, сын [Ионафана, сына] Саулова, вышел навстречу царю. Он не омывал ног своих, не заботился о бороде своей и не мыл одежд своих с того дня, как вышел царь, до дня, когда он возвратился с миром.
2SAM|19|26|Когда он вышел из Иерусалима навстречу царю, царь сказал ему: почему ты, Мемфивосфей, не пошел со мною?
2SAM|19|27|Тот отвечал: господин мой царь! слуга мой обманул меня; ибо я, раб твой, говорил: "оседлаю себе осла и сяду на нем и поеду с царем", так как раб твой хром.
2SAM|19|28|А он оклеветал раба твоего пред господином моим царем. Но господин мой царь, как Ангел Божий; делай, что тебе угодно;
2SAM|19|29|хотя весь дом отца моего был повинен смерти пред господином моим царем, но ты посадил раба твоего между ядущими за столом твоим; какое же имею я право жаловаться еще пред царем?
2SAM|19|30|И сказал ему царь: к чему ты говоришь все это? я сказал, чтобы ты и Сива разделили [между собою] поля.
2SAM|19|31|Но Мемфивосфей отвечал царю: пусть он возьмет даже все, после того как господин мой царь, с миром возвратился в дом свой.
2SAM|19|32|И Верзеллий Галаадитянин пришел из Роглима и перешел с царем Иордан, чтобы проводить его за Иордан.
2SAM|19|33|Верзеллий же был очень стар, лет восьмидесяти. Он продовольствовал царя в пребывание его в Маханаиме, потому что был человек богатый.
2SAM|19|34|И сказал царь Верзеллию: иди со мною, и я буду продовольствовать тебя в Иерусалиме.
2SAM|19|35|Но Верзеллий отвечал царю: долго ли мне осталось жить, чтоб идти с царем в Иерусалим?
2SAM|19|36|Мне теперь восемьдесят лет; различу ли хорошее от худого? Узнает ли раб твой вкус в том, что буду есть, и в том, что буду пить? И буду ли в состоянии слышать голос певцов и певиц? Зачем же рабу твоему быть в тягость господину моему царю?
2SAM|19|37|Еще немного пройдет раб твой с царем за Иордан; за что же царю награждать меня такою милостью?
2SAM|19|38|Позволь рабу твоему возвратиться, чтобы умереть в своем городе, около гроба отца моего и матери моей. Но вот, раб твой, [сын мой] Кимгам пусть пойдет с господином моим, царем, и поступи с ним, как тебе угодно.
2SAM|19|39|И сказал царь: пусть идет со мною Кимгам, и я сделаю для него, что тебе угодно; и все, чего бы ни пожелал ты от меня, я сделаю для тебя.
2SAM|19|40|И перешел весь народ Иордан, и царь [также]. И поцеловал царь Верзеллия и благословил его, и он возвратился в место свое.
2SAM|19|41|И отправился царь в Галгал, отправился с ним и Кимгам; и весь народ Иудейский провожал царя, и половина народа Израильского.
2SAM|19|42|И вот, все Израильтяне пришли к царю и сказали царю: зачем братья наши, мужи Иудины, похитили тебя и проводили царя в дом его и всех людей Давида с ним через Иордан?
2SAM|19|43|И отвечали все мужи Иудины Израильтянам: затем, что царь ближний нам; и из–за чего сердиться вам на это? Разве мы что–нибудь съели у царя, или получили от него подарки?
2SAM|19|44|И отвечали Израильтяне мужам Иудиным и сказали: мы десять частей у царя, также и у Давида мы более, нежели вы; зачем же вы унизили нас? Не нам ли принадлежало первое слово о том, чтобы возвратить нашего царя? Но слово мужей Иудиных было сильнее, нежели слово Израильтян.
2SAM|20|1|Там случайно находился один негодный человек, по имени Савей, сын Бихри, Вениамитянин; он затрубил трубою и сказал: нет нам части в Давиде, и нет нам доли в сыне Иессеевом; все по шатрам своим, Израильтяне!
2SAM|20|2|И отделились все Израильтяне от Давида [и пошли] за Савеем, сыном Бихри; Иудеи же остались на стороне царя своего, от Иордана до Иерусалима.
2SAM|20|3|И пришел Давид в свой дом в Иерусалиме, и взял царь десять жен наложниц, которых он оставлял стеречь дом, и поместил их в особый дом под надзор, и содержал их, но не ходил к ним. И содержались они там до дня смерти своей, живя как вдовы.
2SAM|20|4|И сказал Давид Амессаю: созови ко мне Иудеев в течение трех дней и сам явись сюда.
2SAM|20|5|И пошел Амессай созвать Иудеев, но промедлил более назначенного ему времени.
2SAM|20|6|Тогда Давид сказал Авессе: теперь наделает нам зла Савей, сын Бихри, больше нежели Авессалом; возьми ты слуг господина твоего и преследуй его, чтобы он не нашел себе укрепленных городов и не скрылся от глаз наших.
2SAM|20|7|И вышли за ним люди Иоавовы, и Хелефеи и Фелефеи, и все храбрые пошли из Иерусалима преследовать Савея, сына Бихри.
2SAM|20|8|И когда они были близ большого камня, что у Гаваона, то встретился с ними Амессай. Иоав был одет в воинское одеяние свое и препоясан мечом, который висел при бедре в ножнах и который легко выходил из них и входил.
2SAM|20|9|И сказал Иоав Амессаю: здоров ли ты, брат мой? И взял Иоав правою рукою Амессая за бороду, чтобы поцеловать его.
2SAM|20|10|Амессай же не остерегся меча, бывшего в руке Иоава, и тот поразил его им в живот, так что выпали внутренности его на землю, и не повторил ему [удара], и он умер. Иоав и Авесса, брат его, погнались за Савеем, сыном Бихри.
2SAM|20|11|Один из отроков Иоавовых стоял над [Амессаем] и говорил: тот, кто предан Иоаву и кто за Давида, [пусть идет] за Иоавом!
2SAM|20|12|Амессай же лежал в крови среди дороги; и тот человек, увидев, что весь народ останавливается над ним, стащил Амессая с дороги в поле и набросил на него одежду, так как он видел, что всякий проходящий останавливался над ним.
2SAM|20|13|Но когда он был стащен с дороги, то весь народ Израильский пошел вслед за Иоавом преследовать Савея, сына Бихри.
2SAM|20|14|А он прошел чрез все колена Израильские до Авела–Беф–Мааха и чрез весь Берим; и [жители] собирались и шли за ним.
2SAM|20|15|И пришли и осадили его в Авеле–Беф–Маахе; и насыпали вал пред городом и подступили к стене, и все люди, бывшие с Иоавом, старались разрушить стену.
2SAM|20|16|[Тогда] одна умная женщина закричала со стены города: послушайте, послушайте, скажите Иоаву, чтоб он подошел сюда, и я поговорю с ним.
2SAM|20|17|И подошел к ней Иоав, и сказала женщина: ты ли Иоав? И сказал: я. Она сказала: послушай слов рабы твоей. И сказал он: слушаю.
2SAM|20|18|Она сказала: прежде говаривали: "кто хочет спросить, спроси в Авеле"; и так решали дело.
2SAM|20|19|Я из мирных, верных [городов] Израиля; а ты хочешь уничтожить город, и [притом] мать [городов] в Израиле; для чего тебе разрушать наследие Господне?
2SAM|20|20|И отвечал Иоав и сказал: да не будет этого от меня, чтобы я уничтожил или разрушил!
2SAM|20|21|Это не так; но человек с горы Ефремовой, по имени Савей, сын Бихри, поднял руку свою на царя Давида; выдайте мне его одного, и я отступлю от города. И сказала женщина Иоаву: вот, голова его [будет] тебе брошена со стены.
2SAM|20|22|И пошла женщина по всему народу со своим умным словом; и отсекли голову Савею, сыну Бихри, и бросили Иоаву. Тогда [Иоав] затрубил трубою, и разошлись от города все [люди] по своим шатрам; Иоав же возвратился в Иерусалим к царю.
2SAM|20|23|И был Иоав [поставлен] над всем войском Израильским, а Ванея, сын Иодаев, – над Хелефеями и над Фелефеями;
2SAM|20|24|Адорам – над сбором податей; Иосафат, сын Ахилуда – дееписателем;
2SAM|20|25|Суса – писцом; Садок и Авиафар – священниками;
2SAM|20|26|также и Ира Иаритянин был священником у Давида.
2SAM|21|1|Был голод на земле во дни Давида три года, год за годом. И вопросил Давид Господа. И сказал Господь: это ради Саула и кровожадного дома его, за то, что он умертвил Гаваонитян.
2SAM|21|2|Тогда царь призвал Гаваонитян и говорил с ними. Гаваонитяне были не из сынов Израилевых, но из остатков Аморреев; Израильтяне же дали им клятву, но Саул хотел истребить их по ревности своей о потомках Израиля и Иуды.
2SAM|21|3|И сказал Давид Гаваонитянам: что мне сделать для вас, и чем примирить вас, чтобы вы благословили наследие Господне?
2SAM|21|4|И сказали ему Гаваонитяне: не нужно нам ни серебра, ни золота от Саула, или от дома его, и не нужно нам, чтоб умертвили кого в Израиле. Он сказал: чего же вы хотите? я сделаю для вас.
2SAM|21|5|И сказали они царю: того человека, который губил нас и хотел истребить нас, чтобы не было нас ни в одном из пределов Израилевых, –
2SAM|21|6|из его потомков выдай нам семь человек, и мы повесим их пред Господом в Гиве Саула, избранного Господом. И сказал царь: я выдам.
2SAM|21|7|Но пощадил царь Мемфивосфея, сына Ионафана, сына Саулова, ради клятвы именем Господним, которая была между ними, между Давидом и Ионафаном, сыном Сауловым.
2SAM|21|8|И взял царь двух сыновей Рицпы, дочери Айя, которая родила Саулу Армона и Мемфивосфея, и пять сыновей Мелхолы, дочери Сауловой, которых она родила Адриэлу, сыну Верзеллия из Мехолы,
2SAM|21|9|и отдал их в руки Гаваонитян, и они повесили их на горе пред Господом. И погибли все семь вместе; они умерщвлены в первые дни жатвы, в начале жатвы ячменя.
2SAM|21|10|Тогда Рицпа, дочь Айя, взяла вретище и разостлала его себе на той горе [и сидела] от начала жатвы до того времени, пока не полились на них воды Божии с неба, и не допускала касаться их птицам небесным днем и зверям полевым ночью.
2SAM|21|11|И донесли Давиду, что сделала Рицпа, дочь Айя, наложница Саула.
2SAM|21|12|И пошел Давид и взял кости Саула и кости Ионафана, сына его, у жителей Иависа Галаадского, которые тайно взяли их с площади Беф–Сана, где они были повешены Филистимлянами, когда убили Филистимляне Саула на Гелвуе.
2SAM|21|13|И перенес он оттуда кости Саула и кости Ионафана, сына его; и собрали кости повешенных.
2SAM|21|14|И похоронили кости Саула и Ионафана, сына его, в земле Вениаминовой, в Цела, во гробе Киса, отца его. И сделали все, что повелел царь, и умилостивился Бог над страною после того.
2SAM|21|15|И открылась снова война между Филистимлянами и Израильтянами. И вышел Давид и слуги его с ним, и воевали с Филистимлянами; и Давид утомился.
2SAM|21|16|Тогда Иесвий, один из потомков Рефаимов, у которого копье было весом в триста сиклей меди и который опоясан был новым мечом, хотел поразить Давида.
2SAM|21|17|Но ему помог Авесса, сын Саруин, и поразил Филистимлянина и умертвил его. Тогда люди Давидовы поклялись, говоря: не выйдешь ты больше с нами на войну, чтобы не угас светильник Израиля.
2SAM|21|18|Потом была снова война с Филистимлянами в Гобе; тогда Совохай Хушатянин убил Сафута, одного из потомков Рефаимов.
2SAM|21|19|Было и другое сражение в Гобе; тогда убил Елханан, сын Ягаре–Оргима Вифлеемского, Голиафа Гефянина, у которого древко копья было, как навой у ткачей.
2SAM|21|20|Было еще сражение в Гефе; и был [там] один человек рослый, имевший по шести пальцев на руках и на ногах, всего двадцать четыре, также из потомков Рефаимов,
2SAM|21|21|и он поносил Израильтян; но его убил Ионафан, сын Сафая, брата Давидова.
2SAM|21|22|Эти четыре были из рода Рефаимов в Гефе, и они пали от руки Давида и слуг его.
2SAM|22|1|И воспел Давид песнь Господу в день, когда Господь избавил его от руки всех врагов его и от руки Саула, и сказал:
2SAM|22|2|Господь – твердыня моя и крепость моя и избавитель мой.
2SAM|22|3|Бог мой – скала моя; на Него я уповаю; щит мой, рог спасения моего, ограждение мое и убежище мое; Спаситель мой, от бед Ты избавил меня!
2SAM|22|4|Призову Господа достопоклоняемого и от врагов моих спасусь.
2SAM|22|5|Объяли меня волны смерти, и потоки беззакония устрашили меня;
2SAM|22|6|цепи ада облегли меня, и сети смерти опутали меня.
2SAM|22|7|Но в тесноте моей я призвал Господа и к Богу моему воззвал, и Он услышал из чертога Своего голос мой, и вопль мой [дошел] до слуха Его.
2SAM|22|8|Потряслась, всколебалась земля, дрогнули и подвиглись основания небес, ибо разгневался [на них Господь].
2SAM|22|9|Поднялся дым от гнева Его и из уст Его огонь поядающий; горящие угли сыпались от Него.
2SAM|22|10|Наклонил Он небеса и сошел; и мрак под ногами Его;
2SAM|22|11|и воссел на Херувимов, и полетел, и понесся на крыльях ветра;
2SAM|22|12|и мраком покрыл Себя, как сению, сгустив воды облаков небесных;
2SAM|22|13|от блистания пред Ним разгорались угли огненные.
2SAM|22|14|Возгремел с небес Господь, и Всевышний дал глас Свой;
2SAM|22|15|пустил стрелы и рассеял их; [блеснул] молниею и истребил их.
2SAM|22|16|И открылись источники моря, обнажились основания вселенной от грозного гласа Господа, от дуновения духа гнева Его.
2SAM|22|17|Простер Он [руку] с высоты и взял меня, и извлек меня из вод многих;
2SAM|22|18|избавил меня от врага моего сильного, от ненавидящих меня, которые были сильнее меня.
2SAM|22|19|Они восстали на меня в день бедствия моего; но Господь был опорою для меня
2SAM|22|20|и вывел меня на пространное место, избавил меня, ибо Он благоволит ко мне.
2SAM|22|21|Воздал мне Господь по правде моей, по чистоте рук моих вознаградил меня.
2SAM|22|22|Ибо я хранил пути Господа и не был нечестивым пред Богом моим,
2SAM|22|23|ибо все заповеди Его предо мною, и от уставов Его я не отступал,
2SAM|22|24|и был непорочен пред Ним, и остерегался, чтобы не согрешить мне.
2SAM|22|25|И воздал мне Господь по правде моей, по чистоте моей пред очами Его.
2SAM|22|26|С милостивым Ты поступаешь милостиво, с мужем искренним – искренно,
2SAM|22|27|с чистым – чисто, а с лукавым – по лукавству его.
2SAM|22|28|Людей угнетенных Ты спасаешь и взором Своим унижаешь надменных.
2SAM|22|29|Ты, Господи, светильник мой; Господь просвещает тьму мою.
2SAM|22|30|С Тобою я поражаю войско; с Богом моим восхожу на стену.
2SAM|22|31|Бог! – непорочен путь Его, чисто слово Господа, щит Он для всех, надеющихся на Него.
2SAM|22|32|Ибо кто Бог, кроме Господа, и кто защита, кроме Бога нашего?
2SAM|22|33|Бог препоясует меня силою, устрояет мне верный путь;
2SAM|22|34|делает ноги мои, как оленьи, и на высотах поставляет меня;
2SAM|22|35|научает руки мои брани и мышцы мои напрягает, как медный лук.
2SAM|22|36|Ты даешь мне щит спасения Твоего, и милость Твоя возвеличивает меня.
2SAM|22|37|Ты расширяешь шаг мой подо мною, и не колеблются ноги мои.
2SAM|22|38|Я гоняюсь за врагами моими и истребляю их, и не возвращаюсь, доколе не уничтожу их;
2SAM|22|39|и истребляю их и поражаю их, и не встают и падают под ноги мои.
2SAM|22|40|Ты препоясываешь меня силою для войны и низлагаешь предо мною восстающих на меня;
2SAM|22|41|Ты обращаешь ко мне тыл врагов моих, и я истребляю ненавидящих меня.
2SAM|22|42|Они взывают, но нет спасающего, – ко Господу, но Он не внемлет им.
2SAM|22|43|Я рассеваю их, как прах земной, как грязь уличную мну их и топчу их.
2SAM|22|44|Ты избавил меня от мятежа народа моего; Ты сохранил меня, чтоб быть мне главою над иноплеменниками; народ, которого я не знал, служит мне.
2SAM|22|45|Иноплеменники ласкательствуют предо мною; по слуху [обо мне] повинуются мне.
2SAM|22|46|Иноплеменники бледнеют и трепещут в укреплениях своих.
2SAM|22|47|Жив Господь и благословен защитник мой! Да будет превознесен Бог, убежище спасения моего,
2SAM|22|48|Бог, мстящий за меня и покоряющий мне народы
2SAM|22|49|и избавляющий меня от врагов моих! Над восстающими против меня Ты возвысил меня; от человека жестокого Ты избавил меня.
2SAM|22|50|За то я буду славить Тебя, Господи, между иноплеменниками и буду петь имени Твоему,
2SAM|22|51|величественно спасающий царя Своего и творящий милость помазаннику Своему Давиду и потомству его во веки!
2SAM|23|1|Вот последние слова Давида, изречение Давида, сына Иессеева, изречение мужа, поставленного высоко, помазанника Бога Иаковлева и сладкого певца Израилева:
2SAM|23|2|Дух Господень говорит во мне, и слово Его на языке у меня.
2SAM|23|3|Сказал Бог Израилев, говорил о мне скала Израилева: владычествующий над людьми будет праведен, владычествуя в страхе Божием.
2SAM|23|4|И как на рассвете утра, при восходе солнца на безоблачном небе, от сияния после дождя вырастает трава из земли,
2SAM|23|5|не так ли дом мой у Бога? Ибо завет вечный положил Он со мною, твердый и непреложный. Не так ли исходит от Него все спасение мое и все хотение мое?
2SAM|23|6|А нечестивые будут, как выброшенное терние, которого не берут рукою;
2SAM|23|7|но кто касается его, вооружается железом или деревом копья, и огнем сожигают его на месте.
2SAM|23|8|Вот имена храбрых у Давида: Исбосеф Ахаманитянин, главный из трех; он поднял копье свое на восемьсот человек и поразил их в один раз.
2SAM|23|9|По нем Елеазар, сын Додо, сына Ахохи, из трех храбрых, бывших с Давидом, когда они порицанием вызывали Филистимлян, собравшихся на войну;
2SAM|23|10|израильтяне вышли против них, и он стал и поражал Филистимлян до того, что рука его утомилась и прилипла к мечу. И даровал Господь в тот день великую победу, и народ последовал за ним для того только, чтоб обирать [убитых].
2SAM|23|11|За ним Шамма, сын Аге, Гараритянин. Когда Филистимляне собрались в Фирию, где было поле, засеянное чечевицею, и народ побежал от Филистимлян,
2SAM|23|12|то он стал среди поля и сберег его и поразил Филистимлян. И даровал тогда Господь великую победу.
2SAM|23|13|Трое сих главных из тридцати вождей пошли и вошли во время жатвы к Давиду в пещеру Одоллам, когда толпы Филистимлян стояли в долине Рефаимов.
2SAM|23|14|Давид был тогда в укрепленном месте, а отряд Филистимлян – в Вифлееме.
2SAM|23|15|И захотел Давид пить, и сказал: кто напоит меня водою из колодезя Вифлеемского, что у ворот?
2SAM|23|16|Тогда трое этих храбрых пробились сквозь стан Филистимский и почерпнули воды из колодезя Вифлеемского, что у ворот, и взяли и принесли Давиду. Но он не захотел пить ее и вылил ее во славу Господа,
2SAM|23|17|и сказал: сохрани меня Господь, чтоб я сделал это! не кровь ли это людей, ходивших с опасностью собственной жизни? И не захотел пить ее. Вот что сделали эти трое храбрых!
2SAM|23|18|И Авесса, брат Иоава, сын Саруин, был главным из трех; он убил копьем своим триста человек и был в славе у тех троих.
2SAM|23|19|Из трех он был знатнейшим и был начальником, но с теми тремя не равнялся.
2SAM|23|20|Ванея, сын Иодая, мужа храброго, великий по делам, из Кавцеила; он поразил двух сыновей Ариила Моавитского; он же сошел и убил льва во рве в снежное время;
2SAM|23|21|он же убил одного Египтянина человека видного; в руке Египтянина было копье, а он пошел к нему с палкою и отнял копье из руки Египтянина, и убил его собственным его копьем:
2SAM|23|22|вот что сделал Ванея, сын Иодаев, и он был в славе у трех храбрых;
2SAM|23|23|он был знатнее тридцати, но с теми тремя не равнялся. И поставил его Давид ближайшим исполнителем своих приказаний.
2SAM|23|24|Асаил, брат Иоава – в числе тридцати; Елханан, сын Додо, из Вифлеема,
2SAM|23|25|Шамма Хародитянин, Елика Хародитянин,
2SAM|23|26|Херец Палтитянин, Ира, сын Икеша, Фекоитянин,
2SAM|23|27|Евиезер Анафофянин, Мебуннай Хушатянин,
2SAM|23|28|Цалмон Ахохитянин, Магарай Нетофафянин,
2SAM|23|29|Хелев, сын Бааны, Нетофафянин, Иттай, сын Рибая, из Гивы сынов Вениаминовых,
2SAM|23|30|Ванея Пирафонянин, Иддай из Нахле–Гааша,
2SAM|23|31|Ави–Албон Арбатитянин, Азмавет Бархюмитянин,
2SAM|23|32|Елияхба Шаалбонянин; из сыновей Яшена – Ионафан,
2SAM|23|33|Шама Гараритянин, Ахиам, сын Шарара, Араритянин,
2SAM|23|34|Елифелет, сын Ахасбая, сына Магахати, Елиам, сын Ахитофела, Гилонянин,
2SAM|23|35|Хецрай Кармилитянин, Паарай Арбитянин,
2SAM|23|36|Игал, сын Нафана, из Цобы, Бани Гадитянин,
2SAM|23|37|Целек Аммонитянин, Нахарай Беротянин, оруженосец Иоава, сына Саруи,
2SAM|23|38|Ира Итритянин, Гареб Итритянин,
2SAM|23|39|Урия Хеттеянин. Всех тридцать семь.
2SAM|24|1|Гнев Господень опять возгорелся на Израильтян, и возбудил он в них Давида сказать: пойди, исчисли Израиля и Иуду.
2SAM|24|2|И сказал царь Иоаву военачальнику, который был при нем: пройди по всем коленам Израилевым от Дана до Вирсавии, и исчислите народ, чтобы мне знать число народа.
2SAM|24|3|И сказал Иоав царю: Господь Бог твой да умножит столько народа, сколько есть, и еще во сто раз столько, а очи господина моего царя да увидят [это]; но для чего господин мой царь желает этого дела?
2SAM|24|4|Но слово царя Иоаву и военачальникам превозмогло; и пошел Иоав с военачальниками от царя считать народ Израильский.
2SAM|24|5|И перешли они Иордан и остановились в Ароере, на правой стороне города, который среди долины Гадовой, к Иазеру;
2SAM|24|6|и пришли в Галаад и в землю Тахтим–Ходши; и пришли в Дан–Яан и обошли Сидон;
2SAM|24|7|и пришли к укреплению Тира и во все города Хивеян и Хананеян и вышли на юг Иудеи в Вирсавию;
2SAM|24|8|и обошли всю землю и пришли чрез девять месяцев и двадцать дней в Иерусалим.
2SAM|24|9|И подал Иоав список народной переписи царю; и оказалось, что Израильтян было восемьсот тысяч мужей сильных, способных к войне, а Иудеян пятьсот тысяч.
2SAM|24|10|И вздрогнуло сердце Давидово после того, как он сосчитал народ. И сказал Давид Господу: тяжко согрешил я, поступив так; и ныне молю Тебя, Господи, прости грех раба Твоего, ибо крайне неразумно поступил я.
2SAM|24|11|Когда Давид встал на другой день утром, то было слово Господа к Гаду пророку, прозорливцу Давида:
2SAM|24|12|пойди и скажи Давиду: так говорит Господь: три [наказания] предлагаю Я тебе; выбери себе одно из них, которое совершилось бы над тобою.
2SAM|24|13|И пришел Гад к Давиду, и возвестил ему, и сказал ему: избирай себе, быть ли голоду в стране твоей семь лет, или чтобы ты три месяца бегал от неприятелей твоих, и они преследовали тебя, или чтобы в продолжение трех дней была моровая язва в стране твоей? теперь рассуди и реши, что мне отвечать Пославшему меня.
2SAM|24|14|И сказал Давид Гаду: тяжело мне очень; но пусть впаду я в руки Господа, ибо велико милосердие Его; только бы в руки человеческие не впасть мне.
2SAM|24|15|И послал Господь язву на Израильтян от утра до назначенного времени; и умерло из народа, от Дана до Вирсавии, семьдесят тысяч человек.
2SAM|24|16|И простер Ангел руку свою на Иерусалим, чтобы опустошить его; но Господь пожалел о бедствии и сказал Ангелу, поражавшему народ: довольно, теперь опусти руку твою. Ангел же Господень был тогда у гумна Орны Иевусеянина.
2SAM|24|17|И сказал Давид Господу, когда увидел Ангела, поражавшего народ, говоря: вот, я согрешил, я поступил беззаконно; а эти овцы, что сделали они? пусть же рука Твоя обратится на меня и на дом отца моего.
2SAM|24|18|И пришел в тот день Гад к Давиду и сказал: иди, поставь жертвенник Господу на гумне Орны Иевусеянина.
2SAM|24|19|И пошел Давид по слову Гада, как повелел Господь.
2SAM|24|20|И взглянул Орна и увидел царя и слуг его, шедших к нему, и вышел Орна и поклонился царю лицем своим до земли.
2SAM|24|21|И сказал Орна: зачем пришел господин мой царь к рабу своему? И сказал Давид: купить у тебя гумно для устроения жертвенника Господу, чтобы прекратилось поражение народа.
2SAM|24|22|И сказал Орна Давиду: пусть возьмет и вознесет [в жертву] господин мой, царь, что ему угодно. Вот волы для всесожжения и повозки и упряжь воловья на дрова.
2SAM|24|23|Все это, царь, Орна отдает царю. Еще сказал Орна царю: Господь Бог твой да будет милостив к тебе!
2SAM|24|24|Но царь сказал Орне: нет, я заплачу тебе, что стоит, и не вознесу Господу Богу моему жертвы, [взятой] даром. И купил Давид гумно и волов за пятьдесят сиклей серебра.
2SAM|24|25|И соорудил там Давид жертвенник Господу и принес всесожжения и мирные жертвы. И умилостивился Господь над страною, и прекратилось поражение Израильтян.
