1KGS|1|1|et rex David senuerat habebatque aetatis plurimos dies cumque operiretur vestibus non calefiebat
1KGS|1|2|dixerunt ergo ei servi sui quaeramus domino nostro regi adulescentulam virginem et stet coram rege et foveat eum dormiatque in sinu tuo et calefaciat dominum nostrum regem
1KGS|1|3|quaesierunt igitur adulescentulam speciosam in omnibus finibus Israhel et invenerunt Abisag Sunamitin et adduxerunt eam ad regem
1KGS|1|4|erat autem puella pulchra nimis dormiebatque cum rege et ministrabat ei rex vero non cognovit eam
1KGS|1|5|Adonias autem filius Aggith elevabatur dicens ego regnabo fecitque sibi currum et equites et quinquaginta viros qui ante eum currerent
1KGS|1|6|nec corripuit eum pater suus aliquando dicens quare hoc fecisti erat autem et ipse pulcher valde secundus natu post Absalom
1KGS|1|7|et sermo ei cum Ioab filio Sarviae et cum Abiathar sacerdote qui adiuvabant partes Adoniae
1KGS|1|8|Sadoc vero sacerdos et Banaias filius Ioiadae et Nathan propheta et Semei et Rhei et robur exercitus David non erat cum Adonia
1KGS|1|9|immolatis ergo Adonias arietibus et vitulis et universis pinguibus iuxta lapidem Zoheleth qui erat vicinus fonti Rogel vocavit universos fratres suos filios regis et omnes viros Iuda servos regis
1KGS|1|10|Nathan autem prophetam et Banaiam et robustos quosque et Salomonem fratrem suum non vocavit
1KGS|1|11|dixit itaque Nathan ad Bethsabee matrem Salomonis num audisti quod regnaverit Adonias filius Aggith et dominus noster David hoc ignorat
1KGS|1|12|nunc ergo veni accipe a me consilium et salva animam tuam filiique tui Salomonis
1KGS|1|13|vade et ingredere ad regem David et dic ei nonne tu domine mi rex iurasti mihi ancillae tuae dicens quod Salomon filius tuus regnabit post me et ipse sedebit in solio meo quare ergo regnavit Adonias
1KGS|1|14|et adhuc ibi te loquente cum rege ego veniam post te et conplebo sermones tuos
1KGS|1|15|ingressa est itaque Bethsabee ad regem in cubiculo rex autem senuerat nimis et Abisag Sunamitis ministrabat ei
1KGS|1|16|inclinavit se Bethsabee et adoravit regem ad quam rex quid tibi inquit vis
1KGS|1|17|quae respondens ait domine mi tu iurasti per Dominum Deum tuum ancillae tuae Salomon filius tuus regnabit post me et ipse sedebit in solio meo
1KGS|1|18|et ecce nunc Adonias regnavit te domine mi rex ignorante
1KGS|1|19|mactavit boves et pinguia quaeque et arietes plurimos et vocavit omnes filios regis Abiathar quoque sacerdotem et Ioab principem militiae Salomonem autem servum tuum non vocavit
1KGS|1|20|verumtamen domine mi rex in te oculi respiciunt totius Israhel ut indices eis qui sedere debeat in solio tuo domine mi rex post te
1KGS|1|21|eritque cum dormierit dominus meus rex cum patribus suis erimus ego et filius meus Salomon peccatores
1KGS|1|22|adhuc illa loquente cum rege Nathan prophetes venit
1KGS|1|23|et nuntiaverunt regi dicentes adest Nathan propheta cumque introisset ante conspectum regis et adorasset eum pronus in terram
1KGS|1|24|dixit Nathan domine mi rex tu dixisti Adonias regnet post me et ipse sedeat super thronum meum
1KGS|1|25|quia descendit hodie et immolavit boves et pinguia et arietes plurimos et vocavit universos filios regis et principes exercitus Abiathar quoque sacerdotem illisque vescentibus et bibentibus coram eo et dicentibus vivat rex Adonias
1KGS|1|26|me servum tuum et Sadoc sacerdotem et Banaiam filium Ioiadae et Salomonem famulum tuum non vocavit
1KGS|1|27|numquid a domino meo rege exivit hoc verbum et mihi non indicasti servo tuo qui sessurus esset super thronum domini mei regis post eum
1KGS|1|28|et respondit rex David dicens vocate ad me Bethsabee quae cum fuisset ingressa coram rege et stetisset ante eum
1KGS|1|29|iuravit rex et ait vivit Dominus qui eruit animam meam de omni angustia
1KGS|1|30|quia sicut iuravi tibi per Dominum Deum Israhel dicens Salomon filius tuus regnabit post me et ipse sedebit super solium meum pro me sic faciam hodie
1KGS|1|31|submissoque Bethsabee in terram vultu adoravit regem dicens vivat dominus meus rex David in aeternum
1KGS|1|32|dixit quoque rex David vocate mihi Sadoc sacerdotem et Nathan propheten et Banaiam filium Ioiadae qui cum ingressi fuissent coram rege
1KGS|1|33|dixit ad eos tollite vobiscum servos domini vestri et inponite Salomonem filium meum super mulam meam et ducite eum in Gion
1KGS|1|34|et unguat eum ibi Sadoc sacerdos et Nathan propheta in regem super Israhel et canetis bucina atque dicetis vivat rex Salomon
1KGS|1|35|et ascendetis post eum et veniet et sedebit super solium meum et ipse regnabit pro me illique praecipiam ut sit dux super Israhel et super Iudam
1KGS|1|36|et respondit Banaias filius Ioiadae regi dicens amen sic loquatur Dominus Deus domini mei regis
1KGS|1|37|quomodo fuit Dominus cum domino meo rege sic sit cum Salomone et sublimius faciat solium eius a solio domini mei regis David
1KGS|1|38|descendit ergo Sadoc sacerdos et Nathan propheta et Banaias filius Ioiadae et Cherethi et Felethi et inposuerunt Salomonem super mulam regis David et adduxerunt eum in Gion
1KGS|1|39|sumpsitque Sadoc sacerdos cornu olei de tabernaculo et unxit Salomonem et cecinerunt bucina et dixit omnis populus vivat rex Salomon
1KGS|1|40|et ascendit universa multitudo post eum et populus canentium tibiis et laetantium gaudio magno et insonuit terra ad clamorem eorum
1KGS|1|41|audivit autem Adonias et omnes qui invitati fuerant ab eo iamque convivium finitum erat sed et Ioab audita voce tubae ait quid sibi vult clamor civitatis tumultuantis
1KGS|1|42|adhuc illo loquente Ionathan filius Abiathar sacerdotis venit cui dixit Adonias ingredere quia vir fortis es et bona nuntians
1KGS|1|43|responditque Ionathan Adoniae nequaquam dominus enim noster rex David regem constituit Salomonem
1KGS|1|44|misitque cum eo Sadoc sacerdotem et Nathan prophetam et Banaiam filium Ioiadae et Cherethi et Felethi et inposuerunt eum super mulam regis
1KGS|1|45|unxeruntque eum Sadoc sacerdos et Nathan propheta regem in Gion et ascenderunt inde laetantes et insonuit civitas haec est vox quam audistis
1KGS|1|46|sed et Salomon sedit super solio regni
1KGS|1|47|et ingressi servi regis benedixerunt domino nostro regi David dicentes amplificet Deus nomen Salomonis super nomen tuum et magnificet thronum eius super thronum tuum et adoravit rex in lectulo suo
1KGS|1|48|insuper et haec locutus est benedictus Dominus Deus Israhel qui dedit hodie sedentem in solio meo videntibus oculis meis
1KGS|1|49|territi sunt ergo et surrexerunt omnes qui invitati fuerant ab Adonia et ivit unusquisque in viam suam
1KGS|1|50|Adonias autem timens Salomonem surrexit et abiit tenuitque cornu altaris
1KGS|1|51|et nuntiaverunt Salomoni dicentes ecce Adonias timens regem Salomonem tenuit cornu altaris dicens iuret mihi hodie rex Salomon quod non interficiat servum suum gladio
1KGS|1|52|dixitque Salomon si fuerit vir bonus non cadet ne unus quidem capillus eius in terram sin autem malum inventum fuerit in eo morietur
1KGS|1|53|misit ergo rex Salomon et eduxit eum ab altari et ingressus adoravit regem Salomonem dixitque ei Salomon vade in domum tuam
1KGS|2|1|adpropinquaverant autem dies David ut moreretur praecepitque Salomoni filio suo dicens
1KGS|2|2|ego ingredior viam universae terrae confortare et esto vir
1KGS|2|3|et observa custodias Domini Dei tui ut ambules in viis eius et custodias caerimonias eius et praecepta eius et iudicia et testimonia sicut scriptum est in lege Mosi ut intellegas universa quae facis et quocumque te verteris
1KGS|2|4|ut confirmet Dominus sermones suos quos locutus est de me dicens si custodierint filii tui viam suam et ambulaverint coram me in veritate in omni corde suo et in omni anima sua non auferetur tibi vir de solio Israhel
1KGS|2|5|tu quoque nosti quae fecerit mihi Ioab filius Sarviae quae fecerit duobus principibus exercitus Israhel Abner filio Ner et Amasa filio Iether quos occidit et effudit sanguinem belli in pace et posuit cruorem proelii in balteo suo qui erat circa lumbos eius et in calciamento suo quod erat in pedibus eius
1KGS|2|6|facies ergo iuxta sapientiam tuam et non deduces canitiem eius pacifice ad inferos
1KGS|2|7|sed et filiis Berzellai Galaaditis reddes gratiam eruntque comedentes in mensa tua occurrerunt enim mihi quando fugiebam a facie Absalom fratris tui
1KGS|2|8|habes quoque apud te Semei filium Gera filii Iemini de Baurim qui maledixit mihi maledictione pessima quando ibam ad Castra sed quia descendit mihi in occursum cum transirem Iordanem et iuravi ei per Dominum dicens non te interficiam gladio
1KGS|2|9|tu noli pati esse eum innoxium vir autem sapiens es et scies quae facias ei deducesque canos eius cum sanguine ad infernum
1KGS|2|10|dormivit igitur David cum patribus suis et sepultus est in civitate David
1KGS|2|11|dies autem quibus regnavit David super Israhel quadraginta anni sunt in Hebron regnavit septem annis in Hierusalem triginta tribus
1KGS|2|12|Salomon autem sedit super thronum David patris sui et firmatum est regnum eius nimis
1KGS|2|13|et ingressus est Adonias filius Aggith ad Bethsabee matrem Salomonis quae dixit ei pacificusne ingressus tuus qui respondit pacificus
1KGS|2|14|addiditque sermo mihi est ad te cui ait loquere et ille
1KGS|2|15|tu inquit nosti quia meum erat regnum et me proposuerat omnis Israhel sibi in regem sed translatum est regnum et factum est fratris mei a Domino enim constitutum est ei
1KGS|2|16|nunc ergo petitionem unam deprecor a te ne confundas faciem meam quae dixit ad eum loquere
1KGS|2|17|et ille ait precor ut dicas Salomoni regi neque enim negare tibi quicquam potest ut det mihi Abisag Sunamitin uxorem
1KGS|2|18|et ait Bethsabee bene ego loquar pro te regi
1KGS|2|19|venit ergo Bethsabee ad regem Salomonem ut loqueretur ei pro Adonia et surrexit rex in occursum eius adoravitque eam et sedit super thronum suum positus quoque est thronus matri regis quae sedit ad dexteram eius
1KGS|2|20|dixitque ei petitionem unam parvulam ego deprecor a te ne confundas faciem meam dixit ei rex pete mater mi neque enim fas est ut avertam faciem tuam
1KGS|2|21|quae ait detur Abisag Sunamitis Adoniae fratri tuo uxor
1KGS|2|22|responditque rex Salomon et dixit matri suae quare postulas Abisag Sunamitin Adoniae postula ei et regnum ipse est enim frater meus maior me et habet Abiathar sacerdotem et Ioab filium Sarviae
1KGS|2|23|iuravit itaque rex Salomon per Dominum dicens haec faciat mihi Deus et haec addat quia contra animam suam locutus est Adonias verbum hoc
1KGS|2|24|et nunc vivit Dominus qui firmavit me et conlocavit super solium David patris mei et qui fecit mihi domum sicut locutus est quia hodie occidetur Adonias
1KGS|2|25|misitque rex Salomon per manum Banaiae filii Ioiadae qui interfecit eum et mortuus est
1KGS|2|26|Abiathar quoque sacerdoti dixit rex vade in Anathot ad agrum tuum es quidem vir mortis sed hodie te non interficiam quia portasti arcam Domini Dei coram David patre meo et sustinuisti laborem in omnibus in quibus laboravit pater meus
1KGS|2|27|eiecit ergo Salomon Abiathar ut non esset sacerdos Domini ut impleretur sermo Domini quem locutus est super domum Heli in Silo
1KGS|2|28|venit autem nuntius ad Ioab quod Ioab declinasset post Adoniam et post Absalom non declinasset fugit ergo Ioab in tabernaculum Domini et adprehendit cornu altaris
1KGS|2|29|nuntiatumque est regi Salomoni quod fugisset Ioab in tabernaculum Domini et esset iuxta altare misitque Salomon Banaiam filium Ioiadae dicens vade interfice eum
1KGS|2|30|venit Banaias ad tabernaculum Domini et dixit ei haec dicit rex egredere qui ait non egrediar sed hic moriar renuntiavit Banaias regi sermonem dicens haec locutus est Ioab et haec respondit mihi
1KGS|2|31|dixitque ei rex fac sicut locutus est et interfice eum et sepeli et amovebis sanguinem innocentem qui effusus est a Ioab a me et a domo patris mei
1KGS|2|32|et reddat Dominus sanguinem eius super caput eius quia interfecit duos viros iustos melioresque se et occidit eos gladio patre meo David ignorante Abner filium Ner principem militiae Israhel et Amasa filium Iether principem exercitus Iuda
1KGS|2|33|et revertetur sanguis illorum in caput Ioab et in caput seminis eius in sempiternum David autem et semini eius et domui et throno illius sit pax usque in aeternum a Domino
1KGS|2|34|ascendit itaque Banaias filius Ioiadae et adgressus eum interfecit sepultusque est in domo sua in deserto
1KGS|2|35|et constituit rex Banaiam filium Ioiadae pro eo super exercitum et Sadoc sacerdotem posuit pro Abiathar
1KGS|2|36|misit quoque rex et vocavit Semei dixitque ei aedifica tibi domum in Hierusalem et habita ibi et non egredieris inde huc atque illuc
1KGS|2|37|quacumque autem die egressus fueris et transieris torrentem Cedron scito te interficiendum sanguis tuus erit super caput tuum
1KGS|2|38|dixitque Semei regi bonus sermo sicut locutus est dominus meus rex sic faciet servus tuus habitavit itaque Semei in Hierusalem diebus multis
1KGS|2|39|factum est autem post annos tres ut fugerent servi Semei ad Achis filium Maacha regem Geth nuntiatumque est Semei quod servi eius essent in Geth
1KGS|2|40|et surrexit Semei et stravit asinum suum ivitque in Geth ad Achis ad requirendos servos suos et adduxit eos de Geth
1KGS|2|41|nuntiatum est autem Salomoni quod isset Semei in Geth de Hierusalem et redisset
1KGS|2|42|et mittens vocavit eum dixitque illi nonne testificatus sum tibi per Dominum et praedixi tibi quacumque die egressus ieris huc et illuc scito te esse moriturum et respondisti mihi bonus sermo audivi
1KGS|2|43|quare ergo non custodisti iusiurandum Domini et praeceptum quod praeceperam tibi
1KGS|2|44|dixitque rex ad Semei tu nosti omne malum cuius tibi conscium est cor tuum quod fecisti David patri meo reddidit Dominus malitiam tuam in caput tuum
1KGS|2|45|et rex Salomon benedictus et thronus David erit stabilis coram Domino usque in sempiternum
1KGS|2|46|iussit itaque rex Banaiae filio Ioiadae qui egressus percussit eum et mortuus est
1KGS|3|1|confirmatum est igitur regnum in manu Salomonis et adfinitate coniunctus est Pharaoni regi Aegypti accepit namque filiam eius et adduxit in civitatem David donec conpleret aedificans domum suam et domum Domini et murum Hierusalem per circuitum
1KGS|3|2|et tamen populus immolabat in excelsis non enim aedificatum erat templum nomini Domini usque in die illo
1KGS|3|3|dilexit autem Salomon Dominum ambulans in praeceptis David patris sui excepto quod in excelsis immolabat et accendebat thymiama
1KGS|3|4|abiit itaque in Gabaon ut immolaret ibi illud quippe erat excelsum maximum mille hostias in holocaustum obtulit Salomon super altare illud in Gabaon
1KGS|3|5|apparuit Dominus Salomoni per somnium nocte dicens postula quod vis ut dem tibi
1KGS|3|6|et ait Salomon tu fecisti cum servo tuo David patre meo misericordiam magnam sicut ambulavit in conspectu tuo in veritate et iustitia et recto corde tecum custodisti ei misericordiam tuam grandem et dedisti ei filium sedentem super thronum eius sicut et hodie
1KGS|3|7|et nunc Domine Deus tu regnare fecisti servum tuum pro David patre meo ego autem sum puer parvus et ignorans egressum et introitum meum
1KGS|3|8|et servus tuus in medio est populi quem elegisti populi infiniti qui numerari et supputari non potest prae multitudine
1KGS|3|9|dabis ergo servo tuo cor docile ut iudicare possit populum tuum et discernere inter malum et bonum quis enim potest iudicare populum istum populum tuum hunc multum
1KGS|3|10|placuit ergo sermo coram Domino quod Salomon rem huiuscemodi postulasset
1KGS|3|11|et dixit Deus Salomoni quia postulasti verbum hoc et non petisti tibi dies multos nec divitias aut animam inimicorum tuorum sed postulasti tibi sapientiam ad discernendum iudicium
1KGS|3|12|ecce feci tibi secundum sermones tuos et dedi tibi cor sapiens et intellegens in tantum ut nullus ante te similis tui fuerit nec post te surrecturus sit
1KGS|3|13|sed et haec quae non postulasti dedi tibi divitias scilicet et gloriam ut nemo fuerit similis tui in regibus cunctis retro diebus
1KGS|3|14|si autem ambulaveris in viis meis et custodieris praecepta mea et mandata mea sicut ambulavit pater tuus longos faciam dies tuos
1KGS|3|15|igitur evigilavit Salomon et intellexit quod esset somnium cumque venisset Hierusalem stetit coram arca foederis Domini et obtulit holocausta et fecit victimas pacificas et grande convivium universis famulis suis
1KGS|3|16|tunc venerunt duae mulieres meretrices ad regem steteruntque coram eo
1KGS|3|17|quarum una ait obsecro mi domine ego et mulier haec habitabamus in domo una et peperi apud eam in cubiculo
1KGS|3|18|tertia vero die postquam ego peperi peperit et haec et eramus simul nullusque alius in domo nobiscum exceptis nobis duabus
1KGS|3|19|mortuus est autem filius mulieris huius nocte dormiens quippe oppressit eum
1KGS|3|20|et consurgens intempesta nocte silentio tulit filium meum de latere meo ancillae tuae dormientis et conlocavit in sinu suo suum autem filium qui erat mortuus posuit in sinu meo
1KGS|3|21|cumque surrexissem mane ut darem lac filio meo apparuit mortuus quem diligentius intuens clara luce deprehendi non esse meum quem genueram
1KGS|3|22|responditque altera mulier non est ita sed filius tuus mortuus est meus autem vivit e contrario illa dicebat mentiris filius quippe meus vivit et filius tuus mortuus est atque in hunc modum contendebant coram rege
1KGS|3|23|tunc rex ait haec dicit filius meus vivit et filius tuus mortuus est et ista respondit non sed filius tuus mortuus est et filius meus vivit
1KGS|3|24|dixit ergo rex adferte mihi gladium cumque adtulissent gladium coram rege
1KGS|3|25|dividite inquit infantem vivum in duas partes et date dimidiam partem uni et dimidiam partem alteri
1KGS|3|26|dixit autem mulier cuius filius erat vivus ad regem commota sunt quippe viscera eius super filio suo obsecro domine date illi infantem vivum et nolite interficere eum contra illa dicebat nec mihi nec tibi sit dividatur
1KGS|3|27|respondens rex ait date huic infantem vivum et non occidatur haec est mater eius
1KGS|3|28|audivit itaque omnis Israhel iudicium quod iudicasset rex et timuerunt regem videntes sapientiam Dei esse in eo ad faciendum iudicium
1KGS|4|1|erat autem rex Salomon regnans super omnem Israhel
1KGS|4|2|et hii principes quos habebat Azarias filius Sadoc sacerdos
1KGS|4|3|Helioreph et Ahia filii Sesa scribae Iosaphat filius Ahilud a commentariis
1KGS|4|4|Banaias filius Ioiadae super exercitum Sadoc autem et Abiathar sacerdotes
1KGS|4|5|Azarias filius Nathan super eos qui adsistebant regi Zabud filius Nathan sacerdos amicus regis
1KGS|4|6|et Ahisar praepositus domus et Adoniram filius Abda super tributa
1KGS|4|7|habebat autem Salomon duodecim praefectos super omnem Israhel qui praebebant annonam regi et domui eius per singulos enim menses in anno singuli necessaria ministrabant
1KGS|4|8|et haec nomina eorum Benhur in monte Ephraim
1KGS|4|9|Bendecar in Macces et in Salebbim et in Bethsemes et Helon Bethanan
1KGS|4|10|Benesed in Araboth ipsius erat Soccho et omnis terra Epher
1KGS|4|11|Benabinadab cuius omnis Nepthad Dor Tapheth filiam Salomonis habebat uxorem
1KGS|4|12|Bana filius Ahilud regebat Thanac et Mageddo et universam Bethsan quae est iuxta Sarthana subter Hiezrahel a Bethsan usque Abelmeula e regione Iecmaan
1KGS|4|13|Bengaber in Ramoth Galaad habebat Avothiair filii Manasse in Galaad ipse praeerat in omni regione Argob quae est in Basan sexaginta civitatibus magnis atque muratis quae habebant seras aereas
1KGS|4|14|Ahinadab filius Addo praeerat in Manaim
1KGS|4|15|Ahimaas in Nepthali sed et ipse habebat Basmath filiam Salomonis in coniugio
1KGS|4|16|Baana filius Usi in Aser et in Balod
1KGS|4|17|Iosaphat filius Pharue in Isachar
1KGS|4|18|Semei filius Hela in Beniamin
1KGS|4|19|Gaber filius Uri in terra Galaad in terra Seon regis Amorrei et Og regis Basan super omnia quae erant in illa terra
1KGS|4|20|Iuda et Israhel innumerabiles sicut harena maris in multitudine comedentes et bibentes atque laetantes
1KGS|4|21|Salomon autem erat in dicione sua habens omnia regna sicut a flumine terrae Philisthim usque ad terminum Aegypti offerentium sibi munera et servientium ei cunctis diebus vitae eius
1KGS|4|22|erat autem cibus Salomonis per dies singulos triginta chori similae et sexaginta chori farinae
1KGS|4|23|decem boves pingues et viginti boves pascuales et centum arietes excepta venatione cervorum caprearum atque bubalorum et avium altilium
1KGS|4|24|ipse enim obtinebat omnem regionem quae erat trans flumen quasi a Thapsa usque Gazam et cunctos reges illarum regionum et habebat pacem ex omni parte in circuitu
1KGS|4|25|habitabatque Iudas et Israhel absque timore ullo unusquisque sub vite sua et sub ficu sua a Dan usque Bersabee cunctis diebus Salomonis
1KGS|4|26|et habebat Salomon quadraginta milia praesepia equorum currulium et duodecim milia equestrium
1KGS|4|27|nutriebantque eos supradicti regis praefecti sed et necessaria mensae regis Salomonis cum ingenti cura praebebant in tempore suo
1KGS|4|28|hordeum quoque et paleas equorum et iumentorum deferebant in locum ubi erat rex iuxta constitutum sibi
1KGS|4|29|dedit quoque Deus sapientiam Salomoni et prudentiam multam nimis et latitudinem cordis quasi harenam quae est in litore maris
1KGS|4|30|et praecedebat sapientia Salomonis sapientiam omnium Orientalium et Aegyptiorum
1KGS|4|31|et erat sapientior cunctis hominibus sapientior Aethan Ezraita et Heman et Chalcal et Dorda filiis Maol et erat nominatus in universis gentibus per circuitum
1KGS|4|32|locutus est quoque Salomon tria milia parabolas et fuerunt carmina eius quinque et mille
1KGS|4|33|et disputavit super lignis a cedro quae est in Libano usque ad hysopum quae egreditur de pariete et disseruit de iumentis et volucribus et reptilibus et piscibus
1KGS|4|34|et veniebant de cunctis populis ad audiendam sapientiam Salomonis et ab universis regibus terrae qui audiebant sapientiam eius
1KGS|5|1|misit quoque Hiram rex Tyri servos suos ad Salomonem audivit enim quod ipsum unxissent regem pro patre eius quia amicus fuerat Hiram David omni tempore
1KGS|5|2|misit autem et Salomon ad Hiram dicens
1KGS|5|3|tu scis voluntatem David patris mei et quia non potuerit aedificare domum nomini Domini Dei sui propter bella inminentia per circuitum donec daret Dominus eos sub vestigio pedum eius
1KGS|5|4|nunc autem requiem dedit Deus meus mihi per circuitum non est Satan neque occursus malus
1KGS|5|5|quam ob rem cogito aedificare templum nomini Domini Dei mei sicut locutus est Dominus David patri meo dicens filius tuus quem dabo pro te super solium tuum ipse aedificabit domum nomini meo
1KGS|5|6|praecipe igitur ut praecidant mihi cedros de Libano et servi mei sint cum servis tuis mercedem autem servorum tuorum dabo tibi quamcumque praeceperis scis enim quoniam non est in populo meo vir qui noverit ligna caedere sicut Sidonii
1KGS|5|7|cum ergo audisset Hiram verba Salomonis laetatus est valde et ait benedictus Dominus hodie qui dedit David filium sapientissimum super populum hunc plurimum
1KGS|5|8|et misit Hiram ad Salomonem dicens audivi quaecumque mandasti mihi ego faciam omnem voluntatem tuam in lignis cedrinis et abiegnis
1KGS|5|9|servi mei deponent ea de Libano ad mare et ego conponam ea in ratibus in mari usque ad locum quem significaveris mihi et adplicabo ea ibi et tu tolles ea praebebisque necessaria mihi ut detur cibus domui meae
1KGS|5|10|itaque Hiram dabat Salomoni ligna cedrina et ligna abiegna iuxta omnem voluntatem eius
1KGS|5|11|Salomon autem praebebat Hiram viginti milia chororum tritici in cibum domui eius et viginti choros purissimi olei haec tribuebat Salomon Hiram per annos singulos
1KGS|5|12|dedit quoque Dominus sapientiam Salomoni sicut locutus est ei et erat pax inter Hiram et Salomonem et percusserunt foedus ambo
1KGS|5|13|legitque rex Salomon operas de omni Israhel et erat indictio triginta milia virorum
1KGS|5|14|mittebatque eos in Libanum decem milia per menses singulos vicissim ita ut duobus mensibus essent in domibus suis et Adoniram erat super huiuscemodi indictione
1KGS|5|15|fuerunt itaque Salomoni septuaginta milia eorum qui onera portabant et octoginta milia latomorum in monte
1KGS|5|16|absque praepositis qui praeerant singulis operibus numero trium milium et trecentorum praecipientium populo et his qui faciebant opus
1KGS|5|17|praecepitque rex ut tollerent lapides grandes lapides pretiosos in fundamentum templi et quadrarent eos
1KGS|5|18|quos dolaverunt cementarii Salomonis et cementarii Hiram porro Biblii praeparaverunt ligna et lapides ad aedificandam domum
1KGS|6|1|factum est igitur quadringentesimo et octogesimo anno egressionis filiorum Israhel de terra Aegypti in anno quarto mense zio ipse est mensis secundus regis Salomonis super Israhel aedificare coepit domum Domino
1KGS|6|2|domus autem quam aedificabat rex Salomon Domino habebat sexaginta cubitos in longitudine et viginti cubitos in latitudine et triginta cubitos in altitudine
1KGS|6|3|et porticus erat ante templum viginti cubitorum longitudinis iuxta mensuram latitudinis templi et habebat decem cubitos latitudinis ante faciem templi
1KGS|6|4|fecitque in templo fenestras obliquas
1KGS|6|5|et aedificavit super parietem templi tabulata per gyrum in parietibus domus per circuitum templi et oraculi et fecit latera in circuitu
1KGS|6|6|tabulatum quod subter erat quinque cubitos habebat latitudinis et medium tabulatum sex cubitorum latitudinis et tertium tabulatum septem habens cubitos latitudinis trabes autem posuit in domo per circuitum forinsecus ut non hererent muris templi
1KGS|6|7|domus autem cum aedificaretur lapidibus dedolatis atque perfectis aedificata est et malleus et securis et omne ferramentum non sunt audita in domo cum aedificaretur
1KGS|6|8|ostium lateris medii in parte erat domus dexterae et per cocleam ascendebant in medium cenaculum et a medio in tertium
1KGS|6|9|et aedificavit domum et consummavit eam texit quoque domum laquearibus cedrinis
1KGS|6|10|et aedificavit tabulatum super omnem domum quinque cubitis altitudinis et operuit domum lignis cedrinis
1KGS|6|11|et factus est sermo Domini ad Salomonem dicens
1KGS|6|12|domus haec quam aedificas si ambulaveris in praeceptis meis et iudicia mea feceris et custodieris omnia mandata mea gradiens per ea firmabo sermonem meum tibi quem locutus sum ad David patrem tuum
1KGS|6|13|et habitabo in medio filiorum Israhel et non derelinquam populum meum Israhel
1KGS|6|14|igitur aedificavit Salomon domum et consummavit eam
1KGS|6|15|et aedificavit parietes domus intrinsecus tabulatis cedrinis a pavimento domus usque ad summitatem parietum et usque ad laquearia operuit lignis intrinsecus et texit pavimentum domus tabulis abiegnis
1KGS|6|16|aedificavitque viginti cubitorum ad posteriorem partem templi tabulata cedrina a pavimento usque ad superiora et fecit interiorem domum oraculi in sanctum sanctorum
1KGS|6|17|porro quadraginta cubitorum erat ipsum templum pro foribus oraculi
1KGS|6|18|et cedro omnis domus intrinsecus vestiebatur habens tornaturas suas et iuncturas fabrefactas et celaturas eminentes omnia cedrinis tabulis vestiebantur nec omnino lapis apparere poterat in pariete
1KGS|6|19|oraculum autem in medio domus in interiori parte fecerat ut poneret ibi arcam foederis Domini
1KGS|6|20|porro oraculum habebat viginti cubitos longitudinis et viginti cubitos latitudinis et viginti cubitos altitudinis et operuit illud atque vestivit auro purissimo sed et altare vestivit cedro
1KGS|6|21|domum quoque ante oraculum operuit auro purissimo et adfixit lamminas clavis aureis
1KGS|6|22|nihilque erat in templo quod non auro tegeretur sed et totum altare oraculi texit auro
1KGS|6|23|et fecit in oraculo duo cherubin de lignis olivarum decem cubitorum altitudinis
1KGS|6|24|quinque cubitorum ala cherub una et quinque cubitorum ala cherub altera id est decem cubitos habentes a summitate alae usque ad alae alterius summitatem
1KGS|6|25|decem quoque cubitorum erat cherub secundus mensura pari et opus unum erat in duobus cherubin
1KGS|6|26|id est altitudinem habebat unus cherub decem cubitorum et similiter cherub secundus
1KGS|6|27|posuitque cherubin in medio templi interioris extendebant autem alas suas cherubin et tangebat ala una parietem et ala cherub secundi tangebat parietem alterum alae autem alterae in media parte templi se invicem contingebant
1KGS|6|28|texit quoque cherubin auro
1KGS|6|29|et omnes parietes templi per circuitum scalpsit variis celaturis et torno et fecit in eis cherubin et palmas et picturas varias quasi prominentes de pariete et egredientes
1KGS|6|30|sed et pavimentum domus texit auro intrinsecus et extrinsecus
1KGS|6|31|et in ingressu oraculi fecit ostiola de lignis olivarum postesque angulorum quinque
1KGS|6|32|et duo ostia de lignis olivarum et scalpsit in eis picturam cherubin et palmarum species et anaglyfa valde prominentia et texit ea auro et operuit tam cherubin quam palmas et cetera auro
1KGS|6|33|fecitque in introitum templi postes de lignis olivarum quadrangulatos
1KGS|6|34|et duo ostia de lignis abiegnis altrinsecus et utrumque ostium duplex erat et se invicem tenens aperiebatur
1KGS|6|35|et scalpsit cherubin et palmas et celaturas valde eminentes operuitque omnia lamminis aureis opere quadro ad regulam
1KGS|6|36|et aedificavit atrium interius tribus ordinibus lapidum politorum et uno ordine lignorum cedri
1KGS|6|37|anno quarto fundata est domus Domini in mense zio
1KGS|6|38|et in anno undecimo mense bul ipse est mensis octavus perfecta est domus in omni opere suo et in universis utensilibus aedificavitque eam annis septem
1KGS|7|1|domum autem suam aedificavit Salomon tredecim annis et ad perfectum usque perduxit
1KGS|7|2|aedificavit quoque domum saltus Libani centum cubitorum longitudinis et quinquaginta cubitorum latitudinis et triginta cubitorum altitudinis et quattuor deambulacra inter columnas cedrinas ligna quippe cedrina exciderat in columnas
1KGS|7|3|et tabulatis cedrinis vestivit totam cameram quae quadraginta quinque columnis sustentabatur unus autem ordo habebat columnas quindecim
1KGS|7|4|contra se invicem positas
1KGS|7|5|et e regione se respicientes aequali spatio inter columnas et super columnas quadrangulata ligna in cunctis aequalia
1KGS|7|6|et porticum columnarum fecit quinquaginta cubitorum longitudinis et triginta cubitorum latitudinis et alteram porticum in facie maioris porticus et columnas et epistylia super columnas
1KGS|7|7|porticum quoque solii in qua tribunal est fecit et texit lignis cedrinis a pavimento usque ad summitatem
1KGS|7|8|et domuncula in qua sedetur ad iudicandum erat in media porticu simili opere domum quoque fecit filiae Pharaonis quam uxorem duxerat Salomon tali opere quali et hanc porticum
1KGS|7|9|omnia lapidibus pretiosis qui ad normam quandam atque mensuram tam intrinsecus quam extrinsecus serrati erant a fundamento usque ad summitatem parietum et intrinsecus usque ad atrium maius
1KGS|7|10|fundamenta autem de lapidibus pretiosis lapidibus magnis decem sive octo cubitorum
1KGS|7|11|et desuper lapides pretiosi aequalis mensurae secti erant similiterque de cedro
1KGS|7|12|et atrium maius rotundum trium ordinum de lapidibus sectis et unius ordinis dolata cedro necnon et in atrio domus Domini interiori et in porticu domus
1KGS|7|13|misit quoque rex Salomon et tulit Hiram de Tyro
1KGS|7|14|filium mulieris viduae de tribu Nepthali patre Tyrio artificem aerarium et plenum sapientia et intellegentia et doctrina ad faciendum omne opus ex aere qui cum venisset ad regem Salomonem fecit omne opus eius
1KGS|7|15|et finxit duas columnas aereas decem et octo cubitorum altitudinis columnam unam et linea duodecim cubitorum ambiebat columnam utramque
1KGS|7|16|duo quoque capitella fecit quae ponerentur super capita columnarum fusili aere quinque cubitorum altitudinis capitellum unum et quinque cubitorum altitudinis capitellum alterum
1KGS|7|17|et quasi in modum retis et catenarum sibi invicem miro opere contextarum utrumque capitellum columnarum fusile erat septena versuum retiacula in capitello uno et septena retiacula in capitello altero
1KGS|7|18|et perfecit columnas et duos ordines per circuitum retiaculorum singulorum ut tegerent capitella quae erant super summitatem malogranatorum eodem modo fecit et capitello secundo
1KGS|7|19|capitella autem quae erant super capita columnarum quasi opere lilii fabricata erant in porticu quattuor cubitorum
1KGS|7|20|et rursum alia capitella in summitate columnarum desuper iuxta mensuram columnae contra retiacula malogranatorum autem ducenti ordines erant in circuitu capitelli secundi
1KGS|7|21|et statuit duas columnas in porticum templi cumque statuisset columnam dexteram vocavit eam nomine Iachin similiter erexit columnam secundam et vocavit nomen eius Booz
1KGS|7|22|et super capita columnarum opus in modum lilii posuit perfectumque est opus columnarum
1KGS|7|23|fecit quoque mare fusile decem cubitorum a labio usque ad labium rotundum in circuitu quinque cubitorum altitudo eius et resticula triginta cubitorum cingebat illud per circuitum
1KGS|7|24|et scalptura subter labium circumibat illud decem cubitis ambiens mare duo ordines scalpturarum histriatarum erant fusiles
1KGS|7|25|et stabat super duodecim boves e quibus tres respiciebant ad aquilonem et tres ad occidentem et tres ad meridiem et tres ad orientem et mare super eos desuper erat quorum posteriora universa intrinsecus latitabant
1KGS|7|26|grossitudo autem luteris trium unciarum erat labiumque eius quasi labium calicis et folium repandi lilii duo milia batos capiebat
1KGS|7|27|et fecit bases decem aereas quattuor cubitorum longitudinis bases singulas et quattuor cubitorum latitudinis et trium cubitorum altitudinis
1KGS|7|28|et ipsum opus basium interrasile erat et scalpturae inter iuncturas
1KGS|7|29|et inter coronulas et plectas leones et boves et cherubin et in iuncturis similiter desuper et subter leones et boves quasi lora ex aere dependentia
1KGS|7|30|et quattuor rotae per bases singulas et axes aerei et per quattuor partes quasi umeruli subter luterem fusiles contra se invicem respectantes
1KGS|7|31|os quoque luteris intrinsecus erat in capitis summitate et quod forinsecus apparebat unius cubiti erat totum rotundum pariterque habebat unum cubitum et dimidium in angulis autem columnarum variae celaturae erant et media intercolumnia quadrata non rotunda
1KGS|7|32|quattuor quoque rotae quae per quattuor angulos basis erant coherebant subter basi una rota habebat altitudinis cubitum et semis
1KGS|7|33|tales autem rotae erant quales solent in curru fieri et axes earum et radii et canti et modioli omnia fusilia
1KGS|7|34|nam et umeruli illi quattuor per singulos angulos basis unius ex ipsa basi fusiles et coniuncti erant
1KGS|7|35|in summitate autem basis erat quaedam rotunditas dimidii cubiti ita fabrefacta ut luter desuper possit inponi habens celaturas suas et scalpturas varias ex semet ipso
1KGS|7|36|scalpsit quoque in tabulatis illis quae erant ex aere et in angulis cherubin et leones et palmas quasi in similitudinem stantis hominis ut non celata sed adposita per circuitum viderentur
1KGS|7|37|in hunc modum fecit decem bases fusura una et mensura scalpturaque consimili
1KGS|7|38|fecit quoque decem luteres aereos quadraginta batos capiebat luter unus eratque quattuor cubitorum singulosque luteres per singulas id est decem bases posuit
1KGS|7|39|et constituit decem bases quinque ad dexteram partem templi et quinque ad sinistram mare autem posuit ad dexteram partem templi contra orientem ad meridiem
1KGS|7|40|fecit ergo Hiram lebetas et scutras et amulas et perfecit omne opus regis Salomonis in templo Domini
1KGS|7|41|columnas duas et funiculos capitulorum super capitella columnarum duos et retiacula duo ut operirent duos funiculos qui erant super capita columnarum
1KGS|7|42|et malogranata quadringenta in duobus retiaculis duos versus malogranatorum in retiaculis singulis ad operiendos funiculos capitellorum qui erant super capita columnarum
1KGS|7|43|et bases decem et luteres decem super bases
1KGS|7|44|et mare unum et boves duodecim subter mare
1KGS|7|45|et lebetas et scutras et amulas omnia vasa quae fecit Hiram regi Salomoni in domo Domini de aurichalco erant
1KGS|7|46|in campestri regione Iordanis fudit ea rex in argillosa terra inter Socchoth et Sarthan
1KGS|7|47|et posuit Salomon omnia vasa propter multitudinem autem nimiam non erat pondus aeris
1KGS|7|48|fecitque Salomon omnia vasa in domo Domini altare aureum et mensam super quam ponerentur panes propositionis auream
1KGS|7|49|et candelabra aurea quinque ad dexteram et quinque ad sinistram contra oraculum ex auro primo et quasi lilii flores et lucernas desuper aureas et forcipes aureos
1KGS|7|50|et hydrias et fuscinulas et fialas et mortariola et turibula de auro purissimo et cardines ostiorum domus interioris sancti sanctorum et ostiorum domus templi ex auro erant
1KGS|7|51|et perfecit omne opus quod faciebat Salomon in domo Domini et intulit quae sanctificaverat David pater suus argentum et aurum et vasa reposuitque in thesauris domus Domini
1KGS|8|1|tunc congregavit omnes maiores natu Israhel cum principibus tribuum et duces familiarum filiorum Israhel ad regem Salomonem in Hierusalem ut deferrent arcam foederis Domini de civitate David id est de Sion
1KGS|8|2|convenitque ad regem Salomonem universus Israhel in mense hethanim in sollemni die ipse est mensis septimus
1KGS|8|3|veneruntque cuncti senes ex Israhel et tulerunt sacerdotes arcam
1KGS|8|4|et portaverunt arcam Domini et tabernaculum foederis et omnia vasa sanctuarii quae erant in tabernaculo et ferebant ea sacerdotes et Levitae
1KGS|8|5|rex autem Salomon et omnis multitudo Israhel quae convenerat ad eum gradiebatur cum illo ante arcam et immolabant oves et boves absque aestimatione et numero
1KGS|8|6|et intulerunt sacerdotes arcam foederis Domini in locum suum in oraculum templi in sanctum sanctorum subter alas cherubin
1KGS|8|7|siquidem cherubin expandebant alas super locum arcae et protegebant arcam et vectes eius desuper
1KGS|8|8|cumque eminerent vectes et apparerent summitates eorum foris sanctuarium ante oraculum non apparebant ultra extrinsecus qui et fuerunt ibi usque in praesentem diem
1KGS|8|9|in arca autem non est aliud nisi duae tabulae lapideae quas posuerat in ea Moses in Horeb quando pepigit foedus Dominus cum filiis Israhel cum egrederentur de terra Aegypti
1KGS|8|10|factum est autem cum exissent sacerdotes de sanctuario nebula implevit domum Domini
1KGS|8|11|et non poterant sacerdotes stare et ministrare propter nebulam impleverat enim gloria Domini domum Domini
1KGS|8|12|tunc ait Salomon Dominus dixit ut habitaret in nebula
1KGS|8|13|aedificans aedificavi domum in habitaculum tuum firmissimum solium tuum in sempiternum
1KGS|8|14|convertitque rex faciem suam et benedixit omni ecclesiae Israhel omnis enim ecclesia Israhel stabat
1KGS|8|15|et ait benedictus Dominus Deus Israhel qui locutus est ore suo ad David patrem meum et in manibus eius perfecit dicens
1KGS|8|16|a die qua eduxi populum meum Israhel de Aegypto non elegi civitatem de universis tribubus Israhel ut aedificaretur domus et esset nomen meum ibi sed elegi David ut esset super populum meum Israhel
1KGS|8|17|voluitque David pater meus aedificare domum nomini Domini Dei Israhel
1KGS|8|18|et ait Dominus ad David patrem meum quod cogitasti in corde tuo aedificare domum nomini meo bene fecisti hoc ipsum mente tractans
1KGS|8|19|verumtamen tu non aedificabis domum sed filius tuus qui egredietur de renibus tuis ipse aedificabit domum nomini meo
1KGS|8|20|confirmavit Dominus sermonem suum quem locutus est stetique pro David patre meo et sedi super thronum Israhel sicut locutus est Dominus et aedificavi domum nomini Domini Dei Israhel
1KGS|8|21|et constitui ibi locum arcae in qua foedus est Domini quod percussit cum patribus nostris quando egressi sunt de terra Aegypti
1KGS|8|22|stetit autem Salomon ante altare Domini in conspectu ecclesiae Israhel et expandit manus suas in caelum
1KGS|8|23|et ait Domine Deus Israhel non est similis tui Deus in caelo desuper et super terra deorsum qui custodis pactum et misericordiam servis tuis qui ambulant coram te in toto corde suo
1KGS|8|24|qui custodisti servo tuo David patri meo quae locutus es ei ore locutus es et manibus perfecisti ut et haec dies probat
1KGS|8|25|nunc igitur Domine Deus Israhel conserva famulo tuo David patri meo quae locutus es ei dicens non auferetur de te vir coram me qui sedeat super thronum Israhel ita tamen si custodierint filii tui viam suam ut ambulent coram me sicut tu ambulasti in conspectu meo
1KGS|8|26|et nunc Deus Israhel firmentur verba tua quae locutus es servo tuo David patri meo
1KGS|8|27|ergone putandum est quod vere Deus habitet super terram si enim caelum et caeli caelorum te capere non possunt quanto magis domus haec quam aedificavi
1KGS|8|28|sed respice ad orationem servi tui et ad preces eius Domine Deus meus audi hymnum et orationem quam servus tuus orat coram te hodie
1KGS|8|29|ut sint oculi tui aperti super domum hanc nocte et die super domum de qua dixisti erit nomen meum ibi ut exaudias orationem qua orat te servus tuus in loco isto
1KGS|8|30|ut exaudias deprecationem servi tui et populi tui Israhel quodcumque oraverint in loco isto et exaudies in loco habitaculi tui in caelo et cum exaudieris propitius eris
1KGS|8|31|si peccaverit homo in proximum suum et habuerit aliquod iuramentum quo teneatur adstrictus et venerit propter iuramentum coram altari tuo in domum tuam
1KGS|8|32|tu exaudies in caelo et facies et iudicabis servos tuos condemnans impium et reddens viam suam super caput eius iustificansque iustum et retribuens ei secundum iustitiam suam
1KGS|8|33|si fugerit populus tuus Israhel inimicos suos quia peccaturus est tibi et agentes paenitentiam et confitentes nomini tuo venerint et oraverint et deprecati te fuerint in domo hac
1KGS|8|34|exaudi in caelo et dimitte peccatum populi tui Israhel et reduces eos in terram quam dedisti patribus eorum
1KGS|8|35|si clausum fuerit caelum et non pluerit propter peccata eorum et orantes in loco isto paenitentiam egerint nomini tuo et a peccatis suis conversi fuerint propter adflictionem suam
1KGS|8|36|exaudi eos in caelo et dimitte peccata servorum tuorum et populi tui Israhel et ostende eis viam bonam per quam ambulent et da pluviam super terram tuam quam dedisti populo tuo in possessionem
1KGS|8|37|fames si oborta fuerit in terra aut pestilentia aut corruptus aer aurugo lucusta rubigo et adflixerit eum et inimicus eius portas obsidens omnis plaga universa infirmitas
1KGS|8|38|cuncta devotatio et inprecatio quae acciderit omni homini de populo tuo Israhel si quis cognoverit plagam cordis sui et expanderit manus suas in domo hac
1KGS|8|39|tu audies in caelo in loco habitationis tuae et repropitiaberis et facies ut des unicuique secundum omnes vias suas sicut videris cor eius quia tu nosti solus cor omnium filiorum hominum
1KGS|8|40|ut timeant te cunctis diebus quibus vivunt super faciem terrae quam dedisti patribus nostris
1KGS|8|41|insuper et alienigena qui non est de populo tuo Israhel cum venerit de terra longinqua propter nomen tuum audietur enim nomen tuum magnum et manus tua fortis et brachium tuum
1KGS|8|42|extentum ubique cum venerit ergo et oraverit in loco hoc
1KGS|8|43|tu exaudies in caelo in firmamento habitaculi tui et facies omnia pro quibus invocaverit te alienigena ut discant universi populi terrarum nomen tuum timere sicut populus tuus Israhel et probent quia nomen tuum invocatum est super domum hanc quam aedificavi
1KGS|8|44|si egressus fuerit populus tuus ad bellum contra inimicos suos per viam quocumque miseris eos orabunt te contra viam civitatis quam elegisti et contra domum quam aedificavi nomini tuo
1KGS|8|45|et exaudies in caelo orationem eorum et preces eorum et facies iudicium eorum
1KGS|8|46|quod si peccaverint tibi non est enim homo qui non peccet et iratus tradideris eos inimicis suis et capti ducti fuerint in terram inimicorum longe vel prope
1KGS|8|47|et egerint paenitentiam in corde suo in loco captivitatis et conversi deprecati te fuerint in captivitate sua dicentes peccavimus inique egimus impie gessimus
1KGS|8|48|et reversi fuerint ad te in universo corde suo et tota anima sua in terra inimicorum suorum ad quam captivi ducti sunt et oraverint te contra viam terrae suae quam dedisti patribus eorum et civitatis quam elegisti et templi quod aedificavi nomini tuo
1KGS|8|49|exaudies in caelo in firmamento solii tui orationem eorum et preces et facies iudicium eorum
1KGS|8|50|et propitiaberis populo tuo qui peccavit tibi et omnibus iniquitatibus eorum quibus praevaricati sunt in te et dabis misericordiam coram eis qui eos captivos habuerint ut misereantur eis
1KGS|8|51|populus enim tuus est et hereditas tua quos eduxisti de terra Aegypti de medio fornacis ferreae
1KGS|8|52|ut sint oculi tui aperti ad deprecationem servi tui et populi tui Israhel et exaudias eos in universis pro quibus invocaverint te
1KGS|8|53|tu enim separasti eos tibi in hereditatem de universis populis terrae sicut locutus es per Mosen servum tuum quando eduxisti patres nostros de Aegypto Domine Deus
1KGS|8|54|factum est autem cum conplesset Salomon orans Dominum omnem orationem et deprecationem hanc surrexit de conspectu altaris Domini utrumque enim genu in terram fixerat et manus expanderat ad caelum
1KGS|8|55|stetit ergo et benedixit omni ecclesiae Israhel voce magna dicens
1KGS|8|56|benedictus Dominus qui dedit requiem populo suo Israhel iuxta omnia quae locutus est non cecidit ne unus quidem sermo ex omnibus bonis quae locutus est per Mosen servum suum
1KGS|8|57|sit Dominus Deus noster nobiscum sicut fuit cum patribus nostris non derelinquens nos neque proiciens
1KGS|8|58|sed inclinet corda nostra ad se ut ambulemus in universis viis eius et custodiamus mandata eius et caerimonias et iudicia quaecumque mandavit patribus nostris
1KGS|8|59|et sint sermones mei isti quibus deprecatus sum coram Domino adpropinquantes Domino Deo nostro die et nocte ut faciat iudicium servo suo et populo suo Israhel per singulos dies
1KGS|8|60|et sciant omnes populi terrae quia Dominus ipse est Deus et non est ultra absque eo
1KGS|8|61|sit quoque cor nostrum perfectum cum Domino Deo nostro ut ambulemus in decretis eius et custodiamus mandata eius sicut et hodie
1KGS|8|62|igitur rex et omnis Israhel cum eo immolabant victimas coram Domino
1KGS|8|63|mactavitque Salomon hostias pacificas quas immolavit Domino boum viginti duo milia ovium centum viginti milia et dedicaverunt templum Domini rex et filii Israhel
1KGS|8|64|in die illa sanctificavit rex medium atrii quod erat ante domum Domini fecit quippe ibi holocaustum et sacrificium et adipem pacificorum quia altare aereum quod erat coram Domino minus erat et capere non poterat holocausta et sacrificium et adipem pacificorum
1KGS|8|65|fecit ergo Salomon in tempore illo festivitatem celebrem et omnis Israhel cum eo multitudo magna ab introitu Emath usque ad rivum Aegypti coram Domino Deo nostro septem diebus et septem diebus id est quattuordecim diebus
1KGS|8|66|et in die octava dimisit populos qui benedicentes regi profecti sunt in tabernacula sua laetantes et alacri corde super omnibus bonis quae fecerat Dominus David servo suo et Israhel populo suo
1KGS|9|1|factum est autem cum perfecisset Salomon aedificium domus Domini et aedificium regis et omne quod optaverat et voluerat facere
1KGS|9|2|apparuit Dominus ei secundo sicut apparuerat ei in Gabaon
1KGS|9|3|dixitque Dominus ad eum exaudivi orationem tuam et deprecationem tuam qua deprecatus es coram me sanctificavi domum hanc quam aedificasti ut ponerem nomen meum ibi in sempiternum et erunt oculi mei et cor meum ibi cunctis diebus
1KGS|9|4|tu quoque si ambulaveris coram me sicut ambulavit pater tuus in simplicitate cordis et in aequitate et feceris omnia quae praecepi tibi et legitima mea et iudicia mea servaveris
1KGS|9|5|ponam thronum regni tui super Israhel in sempiternum sicut locutus sum David patri tuo dicens non auferetur de genere tuo vir de solio Israhel
1KGS|9|6|si autem aversione aversi fueritis vos et filii vestri non sequentes me nec custodientes mandata mea et caerimonias quas proposui vobis sed abieritis et colueritis deos alienos et adoraveritis eos
1KGS|9|7|auferam Israhel de superficie terrae quam dedi eis et templum quod sanctificavi nomini meo proiciam a conspectu meo eritque Israhel in proverbium et in fabulam cunctis populis
1KGS|9|8|et domus haec erit in exemplum omnis qui transierit per eam stupebit et sibilabit et dicet quare fecit Dominus sic terrae huic et domui huic
1KGS|9|9|et respondebunt quia dereliquerunt Dominum Deum suum qui eduxit patres eorum de terra Aegypti et secuti sunt deos alienos et adoraverunt eos et coluerunt idcirco induxit Dominus super eos omne malum hoc
1KGS|9|10|expletis autem annis viginti postquam aedificaverat Salomon duas domos id est domum Domini et domum regis
1KGS|9|11|Hiram rege Tyri praebente Salomoni ligna cedrina et abiegna et aurum iuxta omne quod opus habuerat tunc dedit Salomon Hiram viginti oppida in terra Galileae
1KGS|9|12|egressusque est Hiram de Tyro ut videret oppida quae dederat ei Salomon et non placuerunt ei
1KGS|9|13|et ait haecine sunt civitates quas dedisti mihi frater et appellavit eas terram Chabul usque in diem hanc
1KGS|9|14|misit quoque Hiram ad regem centum viginti talenta auri
1KGS|9|15|haec est summa expensarum quam obtulit rex Salomon ad aedificandam domum Domini et domum suam et Mello et murum Hierusalem et Eser et Mageddo et Gazer
1KGS|9|16|Pharao rex Aegypti ascendit et cepit Gazer succenditque eam igni et Chananeum qui habitabat in civitate interfecit et dedit eam in dote filiae suae uxori Salomonis
1KGS|9|17|aedificavit ergo Salomon Gazer et Bethoron inferiorem
1KGS|9|18|et Baalath et Palmyram in terra solitudinis
1KGS|9|19|et omnes vicos qui ad se pertinebant et erant absque muro munivit et civitates curruum et civitates equitum et quodcumque ei placuit ut aedificaret in Hierusalem et in Libano et in omni terra potestatis suae
1KGS|9|20|universum populum qui remanserat de Amorreis et Hettheis et Ferezeis et Eveis et Iebuseis qui non sunt de filiis Israhel
1KGS|9|21|horum filios qui remanserant in terra quos scilicet non potuerant filii Israhel exterminare fecit Salomon tributarios usque ad diem hanc
1KGS|9|22|de filiis autem Israhel non constituit Salomon servire quemquam sed erant viri bellatores et ministri eius et principes et duces et praefecti curruum et equorum
1KGS|9|23|erant autem principes super omnia opera Salomonis praepositi quingenti quinquaginta qui habebant subiectum populum et statutis operibus imperabant
1KGS|9|24|filia autem Pharaonis ascendit de civitate David in domum suam quam aedificaverat ei tunc aedificavit Mello
1KGS|9|25|offerebat quoque Salomon tribus vicibus per annos singulos holocausta et pacificas victimas super altare quod aedificaverat Domino et adolebat thymiama coram Domino perfectumque est templum
1KGS|9|26|classem quoque fecit rex Salomon in Asiongaber quae est iuxta Ahilam in litore maris Rubri in terra Idumea
1KGS|9|27|misitque Hiram in classe illa servos suos viros nauticos et gnaros maris cum servis Salomonis
1KGS|9|28|qui cum venissent in Ophir sumptum inde aurum quadringentorum viginti talentorum detulerunt ad regem Salomonem
1KGS|10|1|sed et regina Saba audita fama Salomonis in nomine Domini venit temptare eum in enigmatibus
1KGS|10|2|et ingressa Hierusalem multo comitatu et divitiis camelis portantibus aromata et aurum infinitum nimis et gemmas pretiosas venit ad Salomonem et locuta est ei universa quae habebat in corde suo
1KGS|10|3|et docuit eam Salomon omnia verba quae proposuerat non fuit sermo qui regem posset latere et non responderet ei
1KGS|10|4|videns autem regina Saba omnem sapientiam Salomonis et domum quam aedificaverat
1KGS|10|5|et cibos mensae eius et habitacula servorum et ordinem ministrantium vestesque eorum et pincernas et holocausta quae offerebat in domo Domini non habebat ultra spiritum
1KGS|10|6|dixitque ad regem verus est sermo quem audivi in terra mea
1KGS|10|7|super sermonibus tuis et super sapientia tua et non credebam narrantibus mihi donec ipsa veni et vidi oculis meis et probavi quod media pars mihi nuntiata non fuerit maior est sapientia et opera tua quam rumor quem audivi
1KGS|10|8|beati viri tui et beati servi tui hii qui stant coram te semper et audiunt sapientiam tuam
1KGS|10|9|sit Dominus Deus tuus benedictus cui placuisti et posuit te super thronum Israhel eo quod dilexerit Dominus Israhel in sempiternum et constituit te regem ut faceres iudicium et iustitiam
1KGS|10|10|dedit ergo regi centum viginti talenta auri et aromata multa nimis et gemmas pretiosas non sunt adlata ultra aromata tam multa quam ea quae dedit regina Saba regi Salomoni
1KGS|10|11|sed et classis Hiram quae portabat aurum de Ophir adtulit ex Ophir ligna thyina multa nimis et gemmas pretiosas
1KGS|10|12|fecitque rex de lignis thyinis fulchra domus Domini et domus regiae et citharas lyrasque cantoribus non sunt adlata huiuscemodi ligna thyina neque visa usque in praesentem diem
1KGS|10|13|rex autem Salomon dedit reginae Saba omnia quae voluit et petivit ab eo exceptis his quae ultro obtulerat ei munere regio quae reversa est et abiit in terram suam cum servis suis
1KGS|10|14|erat autem pondus auri quod adferebatur Salomoni per annos singulos sescentorum sexaginta sex talentorum auri
1KGS|10|15|excepto eo quod offerebant viri qui super vectigalia erant et negotiatores universique scruta vendentes et omnes reges Arabiae ducesque terrae
1KGS|10|16|fecit quoque rex Salomon ducenta scuta de auro puro sescentos auri siclos dedit in lamminas scuti unius
1KGS|10|17|et trecentas peltas ex auro probato trecentae minae auri unam peltam vestiebant posuitque ea rex in domo silvae Libani
1KGS|10|18|fecit etiam rex Salomon thronum de ebore grandem et vestivit eum auro fulvo nimis
1KGS|10|19|qui habebat sex gradus et summitas throni rotunda erat in parte posteriori et duae manus hinc atque inde tenentes sedile et duo leones stabant iuxta manus singulas
1KGS|10|20|et duodecim leunculi stantes super sex gradus hinc atque inde non est factum tale opus in universis regnis
1KGS|10|21|sed et omnia vasa de quibus potabat rex Salomon erant aurea et universa supellex domus saltus Libani de auro purissimo non erat argentum nec alicuius pretii putabatur in diebus Salomonis
1KGS|10|22|quia classis regis per mare cum classe Hiram semel per tres annos ibat in Tharsis deferens inde aurum et argentum dentes elefantorum et simias et pavos
1KGS|10|23|magnificatus est ergo rex Salomon super omnes reges terrae divitiis et sapientia
1KGS|10|24|et universa terra desiderabat vultum Salomonis ut audiret sapientiam eius quam dederat Deus in corde eius
1KGS|10|25|et singuli deferebant ei munera vasa argentea et aurea vestes et arma bellica aromata quoque et equos et mulos per annos singulos
1KGS|10|26|congregavitque Salomon currus et equites et facti sunt ei mille quadringenti currus et duodecim milia equitum et disposuit eos per civitates munitas et cum rege in Hierusalem
1KGS|10|27|fecitque ut tanta esset abundantia argenti in Hierusalem quanta lapidum et cedrorum praebuit multitudinem quasi sycomoros quae nascuntur in campestribus
1KGS|10|28|et educebantur equi Salomoni de Aegypto et de Coa negotiatores enim regis emebant de Coa et statuto pretio perducebant
1KGS|10|29|egrediebatur autem quadriga ex Aegypto sescentis siclis argenti et equus centum quinquaginta atque in hunc modum cuncti reges Hettheorum et Syriae equos venundabant
1KGS|11|1|rex autem Salomon amavit mulieres alienigenas multas filiam quoque Pharaonis et Moabitidas et Ammanitidas Idumeas et Sidonias et Chettheas
1KGS|11|2|de gentibus super quibus dixit Dominus filiis Israhel non ingrediemini ad eas neque de illis ingredientur ad vestras certissimo enim avertent corda vestra ut sequamini deos earum his itaque copulatus est Salomon ardentissimo amore
1KGS|11|3|fueruntque ei uxores quasi reginae septingentae et concubinae trecentae et averterunt mulieres cor eius
1KGS|11|4|cumque iam esset senex depravatum est per mulieres cor eius ut sequeretur deos alienos nec erat cor eius perfectum cum Domino Deo suo sicut cor David patris eius
1KGS|11|5|sed colebat Salomon Astharthen deam Sidoniorum et Moloch idolum Ammanitarum
1KGS|11|6|fecitque Salomon quod non placuerat coram Domino et non adimplevit ut sequeretur Dominum sicut pater eius
1KGS|11|7|tunc aedificavit Salomon fanum Chamos idolo Moab in monte qui est contra Hierusalem et Moloch idolo filiorum Ammon
1KGS|11|8|atque in hunc modum fecit universis uxoribus suis alienigenis quae adolebant tura et immolabant diis suis
1KGS|11|9|igitur iratus est Dominus Salomoni quod aversa esset mens eius a Domino Deo Israhel qui apparuerat ei secundo
1KGS|11|10|et praeceperat de verbo hoc ne sequeretur deos alienos et non custodivit quae mandavit ei Dominus
1KGS|11|11|dixit itaque Dominus Salomoni quia habuisti hoc apud te et non custodisti pactum meum et praecepta mea quae mandavi tibi disrumpens scindam regnum tuum et dabo illud servo tuo
1KGS|11|12|verumtamen in diebus tuis non faciam propter David patrem tuum de manu filii tui scindam illud
1KGS|11|13|nec totum regnum auferam sed tribum unam dabo filio tuo propter David servum meum et Hierusalem quam elegi
1KGS|11|14|suscitavit autem Dominus adversarium Salomoni Adad Idumeum de semine regio qui erat in Edom
1KGS|11|15|cum enim esset David in Idumea et ascendisset Ioab princeps militiae ad sepeliendos eos qui fuerant interfecti et occidisset omne masculinum in Idumea
1KGS|11|16|sex enim mensibus ibi moratus est Ioab et omnis Israhel donec interimerent omne masculinum in Idumea
1KGS|11|17|fugit Adad ipse et viri idumei de servis patris eius cum eo ut ingrederetur Aegyptum erat autem Adad puer parvulus
1KGS|11|18|cumque surrexissent de Madian venerunt in Pharan tuleruntque secum viros de Pharan et introierunt Aegyptum ad Pharaonem regem Aegypti qui dedit ei domum et cibos constituit et terram delegavit
1KGS|11|19|et invenit Adad gratiam coram Pharao valde in tantum ut daret ei uxorem sororem uxoris suae germanam Tafnes reginae
1KGS|11|20|genuitque ei soror Tafnes Genebath filium et nutrivit eum Tafnes in domo Pharaonis eratque Genebath habitans apud Pharaonem cum filiis eius
1KGS|11|21|cumque audisset Adad in Aegypto dormisse David cum patribus suis et mortuum esse Ioab principem militiae dixit Pharaoni dimitte me ut vadam in terram meam
1KGS|11|22|dixitque ei Pharao qua enim re apud me indiges ut quaeras ire ad terram tuam at ille respondit nulla sed obsecro ut dimittas me
1KGS|11|23|suscitavit quoque ei Deus adversarium Razon filium Heliada qui fugerat Adadezer regem Soba dominum suum
1KGS|11|24|et congregavit contra eum viros et factus est princeps latronum cum interficeret eos David abieruntque Damascum et habitaverunt ibi et constituerunt eum regem in Damasco
1KGS|11|25|eratque adversarius Israhel cunctis diebus Salomonis et hoc est malum Adad et odium contra Israhel regnavitque in Syria
1KGS|11|26|Hieroboam quoque filius Nabath Ephratheus de Sareda cuius mater erat nomine Sarva mulier vidua servus Salomonis levavit manum contra regem
1KGS|11|27|et haec causa rebellionis adversus eum quia Salomon aedificavit Mello et coaequavit voraginem civitatis David patris sui
1KGS|11|28|erat autem Hieroboam vir fortis et potens vidensque Salomon adulescentem bonae indolis et industrium constituerat eum praefectum super tributa universae domus Ioseph
1KGS|11|29|factum est igitur in tempore illo ut Hieroboam egrederetur de Hierusalem et inveniret eum Ahias Silonites propheta in via opertus pallio novo erant autem duo tantum in agro
1KGS|11|30|adprehendensque Ahia pallium suum novum quo opertus erat scidit in duodecim partes
1KGS|11|31|et ait ad Hieroboam tolle tibi decem scissuras haec enim dicit Dominus Deus Israhel ecce ego scindam regnum de manu Salomonis et dabo tibi decem tribus
1KGS|11|32|porro una tribus remanebit ei propter servum meum David et Hierusalem civitatem quam elegi ex omnibus tribubus Israhel
1KGS|11|33|eo quod dereliquerint me et adoraverint Astharoth deam Sidoniorum et Chamos deum Moab et Melchom deum filiorum Ammon et non ambulaverint in viis meis ut facerent iustitiam coram me et praecepta mea et iudicia sicut David pater eius
1KGS|11|34|nec auferam omne regnum de manu eius sed ducem ponam eum cunctis diebus vitae suae propter David servum meum quem elegi qui custodivit mandata mea et praecepta mea
1KGS|11|35|auferam autem regnum de manu filii eius et dabo tibi decem tribus
1KGS|11|36|filio autem eius dabo tribum unam ut remaneat lucerna David servo meo cunctis diebus coram me in Hierusalem civitatem quam elegi ut esset nomen meum ibi
1KGS|11|37|te autem adsumam et regnabis super omnia quae desiderat anima tua erisque rex super Israhel
1KGS|11|38|si igitur audieris omnia quae praecepero tibi et ambulaveris in viis meis et feceris quod rectum est coram me custodiens mandata mea et praecepta mea sicut fecit David servus meus ero tecum et aedificabo tibi domum fidelem quomodo aedificavi David et tradam tibi Israhel
1KGS|11|39|et adfligam semen David super hoc verumtamen non cunctis diebus
1KGS|11|40|voluit ergo Salomon interficere Hieroboam qui surrexit et aufugit in Aegyptum ad Susac regem Aegypti et fuit in Aegypto usque ad mortem Salomonis
1KGS|11|41|reliquum autem verborum Salomonis et omnia quae fecit et sapientia eius ecce universa scripta sunt in libro verborum Salomonis
1KGS|11|42|dies autem quos regnavit Salomon in Hierusalem super omnem Israhel quadraginta anni sunt
1KGS|11|43|dormivitque Salomon cum patribus suis et sepultus est in civitate David patris sui regnavitque Roboam filius eius pro eo
1KGS|12|1|venit autem Roboam in Sychem illuc enim congregatus erat omnis Israhel ad constituendum eum regem
1KGS|12|2|at Hieroboam filius Nabath cum adhuc esset in Aegypto profugus a facie regis Salomonis audita morte eius reversus est de Aegypto
1KGS|12|3|miseruntque et vocaverunt eum venit ergo Hieroboam et omnis multitudo Israhel et locuti sunt ad Roboam dicentes
1KGS|12|4|pater tuus durissimum iugum inposuit nobis tu itaque nunc inminue paululum de imperio patris tui durissimo et de iugo gravissimo quod inposuit nobis et serviemus tibi
1KGS|12|5|qui ait eis ite usque ad tertium diem et revertimini ad me cumque abisset populus
1KGS|12|6|iniit consilium rex Roboam cum senibus qui adsistebant coram Salomone patre eius dum adviveret et ait quod mihi datis consilium ut respondeam populo
1KGS|12|7|qui dixerunt ei si hodie oboedieris populo huic et servieris et petitioni eorum cesseris locutusque fueris ad eos verba lenia erunt tibi servi cunctis diebus
1KGS|12|8|qui dereliquit consilium senum quod dederant ei et adhibuit adulescentes qui nutriti fuerant cum eo et adsistebant illi
1KGS|12|9|dixitque ad eos quod mihi datis consilium ut respondeam populo huic qui dixerunt mihi levius fac iugum quod inposuit pater tuus super nos
1KGS|12|10|et dixerunt ei iuvenes qui nutriti fuerant cum eo sic loquere populo huic qui locuti sunt ad te dicentes pater tuus adgravavit iugum nostrum tu releva nos sic loqueris ad eos minimus digitus meus grossior est dorso patris mei
1KGS|12|11|et nunc pater meus posuit super vos iugum grave ego autem addam super iugum vestrum pater meus cecidit vos flagellis ego autem caedam scorpionibus
1KGS|12|12|venit ergo Hieroboam et omnis populus ad Roboam die tertia sicut locutus fuerat rex dicens revertimini ad me die tertia
1KGS|12|13|responditque rex populo dura derelicto consilio seniorum quod ei dederant
1KGS|12|14|et locutus est eis secundum consilium iuvenum dicens pater meus adgravavit iugum vestrum ego autem addam iugo vestro pater meus cecidit vos flagellis et ego caedam scorpionibus
1KGS|12|15|et non adquievit rex populo quoniam aversatus eum fuerat Dominus ut suscitaret verbum suum quod locutus fuerat in manu Ahiae Silonitae ad Hieroboam filium Nabath
1KGS|12|16|videns itaque populus quod noluisset eos audire rex respondit ei dicens quae nobis pars in David vel quae hereditas in filio Isai in tabernacula tua Israhel nunc vide domum tuam David et abiit Israhel in tabernacula sua
1KGS|12|17|super filios autem Israhel quicumque habitabant in civitatibus Iuda regnavit Roboam
1KGS|12|18|misit igitur rex Roboam Aduram qui erat super tributum et lapidavit eum omnis Israhel et mortuus est porro rex Roboam festinus ascendit currum et fugit in Hierusalem
1KGS|12|19|recessitque Israhel a domo David usque in praesentem diem
1KGS|12|20|factum est autem cum audisset omnis Israhel quod reversus esset Hieroboam miserunt et vocaverunt eum congregato coetu et constituerunt regem super omnem Israhel nec secutus est quisquam domum David praeter tribum Iuda solam
1KGS|12|21|venit autem Roboam Hierusalem et congregavit universam domum Iuda et tribum Beniamin centum octoginta milia electorum virorum et bellatorum ut pugnaret contra domum Israhel et reduceret regnum Roboam filio Salomonis
1KGS|12|22|factus est vero sermo Domini ad Semeiam virum Dei dicens
1KGS|12|23|loquere ad Roboam filium Salomonis regem Iuda et ad omnem domum Iuda et Beniamin et reliquos de populo dicens
1KGS|12|24|haec dicit Dominus non ascendetis nec bellabitis contra fratres vestros filios Israhel revertatur vir in domum suam a me enim factum est verbum hoc audierunt sermonem Domini et reversi sunt de itinere sicut eis praeceperat Dominus
1KGS|12|25|aedificavit autem Hieroboam Sychem in monte Ephraim et habitavit ibi et egressus inde aedificavit Phanuhel
1KGS|12|26|dixitque Hieroboam in corde suo nunc revertetur regnum ad domum David
1KGS|12|27|si ascenderit populus iste ut faciat sacrificia in domo Domini in Hierusalem et convertetur cor populi huius ad dominum suum Roboam regem Iuda interficientque me et revertentur ad eum
1KGS|12|28|et excogitato consilio fecit duos vitulos aureos et dixit eis nolite ultra ascendere Hierusalem ecce dii tui Israhel qui eduxerunt te de terra Aegypti
1KGS|12|29|posuitque unum in Bethel et alterum in Dan
1KGS|12|30|et factum est verbum hoc in peccatum ibat enim populus ad adorandum vitulum usque in Dan
1KGS|12|31|et fecit fana in excelsis et sacerdotes de extremis populi qui non erant de filiis Levi
1KGS|12|32|constituitque diem sollemnem in mense octavo quintadecima die mensis in similitudinem sollemnitatis quae celebratur in Iuda et ascendens altare similiter fecit in Bethel ut immolaret vitulis quos fabricatus erat constituitque in Bethel sacerdotes excelsorum quae fecerat
1KGS|12|33|et ascendit super altare quod extruxerat in Bethel quintadecima die mensis octavi quem finxerat de corde suo et fecit sollemnitatem filiis Israhel et ascendit super altare ut adoleret incensum
1KGS|13|1|et ecce vir Dei venit de Iuda in sermone Domini in Bethel Hieroboam stante super altare et tus iaciente
1KGS|13|2|et exclamavit contra altare in sermone Domini et ait altare altare haec dicit Dominus ecce filius nascetur domui David Iosias nomine et immolabit super te sacerdotes excelsorum qui nunc in te tura succendunt et ossa hominum incendet super te
1KGS|13|3|deditque in die illa signum dicens hoc erit signum quod locutus est Dominus ecce altare scinditur et effunditur cinis qui in eo est
1KGS|13|4|cumque audisset rex sermonem hominis Dei quem inclamaverat contra altare in Bethel extendit manum suam de altari dicens adprehendite eum et exaruit manus eius quam extenderat contra eum nec valuit retrahere eam ad se
1KGS|13|5|altare quoque scissum est et effusus cinis de altari iuxta signum quod praedixerat vir Dei in sermone Domini
1KGS|13|6|et ait rex ad virum Dei deprecare faciem Domini Dei tui et ora pro me ut restituatur manus mea mihi oravit vir Dei faciem Domini et reversa est manus regis ad eum et facta est sicut prius fuerat
1KGS|13|7|locutus est autem rex ad virum Dei veni mecum domum ut prandeas et dabo tibi munera
1KGS|13|8|responditque vir Dei ad regem si dederis mihi mediam partem domus tuae non veniam tecum nec comedam panem neque bibam aquam in loco isto
1KGS|13|9|sic enim mandatum est mihi in sermone Domini praecipientis non comedes panem neque bibes aquam nec reverteris per viam qua venisti
1KGS|13|10|abiit ergo per aliam viam et non est reversus per iter quo venerat in Bethel
1KGS|13|11|prophetes autem quidam senex habitabat in Bethel ad quem venit filius suus et narravit ei omnia opera quae fecerat vir Dei illa die in Bethel et verba quae locutus fuerat ad regem et narraverunt patri suo
1KGS|13|12|et dixit eis pater eorum per quam viam abiit ostenderunt ei filii sui viam per quam abierat vir Dei qui venerat de Iuda
1KGS|13|13|et ait filiis suis sternite mihi asinum qui cum stravissent ascendit
1KGS|13|14|et abiit post virum Dei et invenit eum sedentem subtus terebinthum et ait illi tune es vir Dei qui venisti de Iuda respondit ille ego sum
1KGS|13|15|dixit ad eum veni mecum domum ut comedas panem
1KGS|13|16|qui ait non possum reverti neque venire tecum nec comedam panem nec bibam aquam in loco isto
1KGS|13|17|quia locutus est Dominus ad me in sermone Domini dicens non comedes panem et non bibes ibi aquam nec reverteris per viam qua ieris
1KGS|13|18|qui ait illi et ego propheta sum similis tui et angelus locutus est mihi in sermone Domini dicens reduc eum tecum in domum tuam et comedat panem et bibat aquam fefellit eum
1KGS|13|19|et reduxit secum comedit ergo panem in domo eius et bibit aquam
1KGS|13|20|cumque sederent ad mensam factus est sermo Domini ad prophetam qui reduxerat eum
1KGS|13|21|et exclamavit ad virum Dei qui venerat de Iuda dicens haec dicit Dominus quia inoboediens fuisti ori Domini et non custodisti mandatum quod praecepit tibi Dominus Deus tuus
1KGS|13|22|et reversus es et comedisti panem et bibisti aquam in loco in quo praecepit tibi ne comederes panem neque biberes aquam non inferetur cadaver tuum in sepulchrum patrum tuorum
1KGS|13|23|cumque comedisset et bibisset stravit asinum prophetae quem reduxerat
1KGS|13|24|qui cum abisset invenit eum leo in via et occidit et erat cadaver eius proiectum in itinere asinus autem stabat iuxta illum et leo stabat iuxta cadaver
1KGS|13|25|et ecce viri transeuntes viderunt cadaver proiectum in via et leonem stantem iuxta cadaver et venerunt et divulgaverunt in civitate in qua prophetes senex ille habitabat
1KGS|13|26|quod cum audisset propheta ille qui reduxerat eum de via ait vir Dei est qui inoboediens fuit ori Domini et tradidit eum Dominus leoni et confregit eum et occidit iuxta verbum Domini quod locutus est ei
1KGS|13|27|dixitque ad filios suos sternite mihi asinum qui cum stravissent
1KGS|13|28|et ille abisset invenit cadaver eius proiectum in via et asinum et leonem stantes iuxta cadaver non comedit leo de cadavere nec laesit asinum
1KGS|13|29|tulit ergo prophetes cadaver viri Dei et posuit illud super asinum et reversus intulit in civitatem prophetae senis ut plangerent eum
1KGS|13|30|et posuit cadaver eius in sepulchro suo et planxerunt eum heu frater
1KGS|13|31|cumque planxissent eum dixit ad filios suos cum mortuus fuero sepelite me in sepulchro in quo vir Dei sepultus est iuxta ossa eius ponite ossa mea
1KGS|13|32|profecto enim veniet sermo quem praedixit in sermone Domini contra altare quod est in Bethel et contra omnia fana excelsorum quae sunt in urbibus Samariae
1KGS|13|33|post verba haec non est reversus Hieroboam de via sua pessima sed e contrario fecit de novissimis populi sacerdotes excelsorum quicumque volebat implebat manum suam et fiebat sacerdos excelsorum
1KGS|13|34|et propter hanc causam peccavit domus Hieroboam et eversa est et deleta de superficie terrae
1KGS|14|1|in tempore illo aegrotavit Abia filius Hieroboam
1KGS|14|2|dixitque Hieroboam uxori suae surge et commuta habitum ne cognoscaris quod sis uxor Hieroboam et vade in Silo ubi est Ahia propheta qui locutus est mihi quod regnaturus essem super populum hunc
1KGS|14|3|tolle quoque in manu tua decem panes et crustula et vas mellis et vade ad illum ipse indicabit tibi quid eventurum sit huic puero
1KGS|14|4|fecit ut dixerat uxor Hieroboam et consurgens abiit in Silo et venit in domum Ahia at ille non poterat videre quia caligaverant oculi eius prae senectute
1KGS|14|5|dixit autem Dominus ad Ahiam ecce uxor Hieroboam ingreditur ut consulat te super filio suo qui aegrotat haec et haec loqueris ei cum ergo illa intraret et dissimularet se esse quae erat
1KGS|14|6|audivit Ahias sonitum pedum eius introeuntis per ostium et ait ingredere uxor Hieroboam quare aliam esse te simulas ego autem missus sum ad te durus nuntius
1KGS|14|7|vade et dic Hieroboam haec dicit Dominus Deus Israhel quia exaltavi te de medio populi et dedi te ducem super populum meum Israhel
1KGS|14|8|et scidi regnum domus David et dedi illud tibi et non fuisti sicut servus meus David qui custodivit mandata mea et secutus est me in toto corde suo faciens quod placitum esset in conspectu meo
1KGS|14|9|sed operatus es male super omnes qui fuerunt ante te et fecisti tibi deos alienos et conflatiles ut me ad iracundiam provocares me autem proiecisti post corpus tuum
1KGS|14|10|idcirco ecce ego inducam mala super domum Hieroboam et percutiam de Hieroboam mingentem ad parietem et clausum et novissimum in Israhel et mundabo reliquias domus Hieroboam sicut mundari solet fimus usque ad purum
1KGS|14|11|qui mortui fuerint de Hieroboam in civitate comedent eos canes qui autem mortui fuerint in agro vorabunt eos aves caeli quia Dominus locutus est
1KGS|14|12|tu igitur surge et vade in domum tuam et in ipso introitu pedum tuorum in urbem morietur puer
1KGS|14|13|et planget eum omnis Israhel et sepeliet iste enim solus infertur de Hieroboam in sepulchrum quia inventus est super eo sermo bonus ad Dominum Deum Israhel in domo Hieroboam
1KGS|14|14|constituet autem sibi Dominus regem super Israhel qui percutiat domum Hieroboam in hac die et in hoc tempore
1KGS|14|15|et percutiet Dominus Israhel sicut moveri solet harundo in aqua et evellet Israhel de terra bona hac quam dedit patribus eorum et ventilabit eos trans Flumen quia fecerunt sibi lucos ut inritarent Dominum
1KGS|14|16|et tradet Dominus Israhel propter peccata Hieroboam qui peccavit et peccare fecit Israhel
1KGS|14|17|surrexit itaque uxor Hieroboam et abiit et venit in Thersa cumque illa ingrederetur limen domus puer mortuus est
1KGS|14|18|et sepelierunt eum et planxit illum omnis Israhel iuxta sermonem Domini quem locutus est in manu servi sui Ahiae prophetae
1KGS|14|19|reliqua autem verborum Hieroboam quomodo pugnaverit et quomodo regnaverit ecce scripta sunt in libro verborum dierum regum Israhel
1KGS|14|20|dies autem quibus regnavit Hieroboam viginti duo anni sunt et dormivit cum patribus suis regnavitque Nadab filius eius pro eo
1KGS|14|21|porro Roboam filius Salomonis regnavit in Iuda quadraginta et unius anni erat Roboam cum regnare coepisset et decem et septem annis regnavit in Hierusalem civitatem quam elegit Dominus ut poneret nomen suum ibi ex omnibus tribubus Israhel nomen autem matris eius Naama Ammanites
1KGS|14|22|et fecit Iudas malum coram Domino et inritaverunt eum super omnibus quae fecerant patres eorum in peccatis suis quae peccaverant
1KGS|14|23|aedificaverunt enim et ipsi sibi aras et statuas et lucos super omnem collem excelsum et subter omnem arborem frondosam
1KGS|14|24|sed et effeminati fuerunt in terra feceruntque omnes abominationes gentium quas adtrivit Dominus ante faciem filiorum Israhel
1KGS|14|25|in quinto autem anno regni Roboam ascendit Sesac rex Aegypti in Hierusalem
1KGS|14|26|et tulit thesauros domus Domini et thesauros regios et universa diripuit scuta quoque aurea quae fecerat Salomon
1KGS|14|27|pro quibus fecit rex Roboam scuta aerea et tradidit ea in manu ducum scutariorum et eorum qui excubabant ante ostium domus regis
1KGS|14|28|cumque ingrederetur rex in domum Domini portabant ea qui praeeundi habebant officium et postea reportabant ad armamentarium scutariorum
1KGS|14|29|reliqua autem sermonum Roboam et omnium quae fecit ecce scripta sunt in libro verborum dierum regum Iuda
1KGS|14|30|fuitque bellum inter Roboam et Hieroboam cunctis diebus
1KGS|14|31|dormivit itaque Roboam cum patribus suis et sepultus est cum eis in civitate David nomen autem matris eius Naama Ammanites et regnavit Abiam filius eius pro eo
1KGS|15|1|igitur in octavodecimo anno regni Hieroboam filii Nabath regnavit Abiam super Iudam
1KGS|15|2|tribus annis regnavit in Hierusalem nomen matris eius Maacha filia Absalom
1KGS|15|3|ambulavitque in omnibus peccatis patris sui quae fecerat ante eum nec erat cor eius perfectum cum Domino Deo suo sicut cor David patris eius
1KGS|15|4|sed propter David dedit ei Dominus Deus suus lucernam in Hierusalem ut suscitaret filium eius post eum et staret Hierusalem
1KGS|15|5|eo quod fecisset David rectum in oculis Domini et non declinasset ab omnibus quae praeceperat ei cunctis diebus vitae suae excepto sermone Uriae Hetthei
1KGS|15|6|attamen bellum fuit inter Roboam et inter Hieroboam omni tempore vitae eius
1KGS|15|7|reliqua autem sermonum Abiam et omnia quae fecit nonne haec scripta sunt in libro verborum dierum regum Iuda fuitque proelium inter Abiam et inter Hieroboam
1KGS|15|8|et dormivit Abiam cum patribus suis et sepelierunt eum in civitate David regnavitque Asa filius eius pro eo
1KGS|15|9|in anno ergo vicesimo Hieroboam regis Israhel regnavit Asa rex Iuda
1KGS|15|10|et quadraginta uno anno regnavit in Hierusalem nomen matris eius Maacha filia Absalom
1KGS|15|11|et fecit Asa rectum ante conspectum Domini sicut David pater eius
1KGS|15|12|et abstulit effeminatos de terra purgavitque universas sordes idolorum quae fecerant patres eius
1KGS|15|13|insuper et Maacham matrem suam amovit ne esset princeps in sacris Priapi et in luco eius quem consecraverat subvertitque specum eius et confregit simulacrum turpissimum et conbusit in torrente Cedron
1KGS|15|14|excelsa autem non abstulit verumtamen cor Asa perfectum erat cum Deo cunctis diebus suis
1KGS|15|15|et intulit ea quae sanctificaverat pater suus et voverat in domum Domini argentum et aurum et vasa
1KGS|15|16|bellum autem erat inter Asa et Baasa regem Israhel cunctis diebus eorum
1KGS|15|17|ascendit quoque Baasa rex Israhel in Iudam et aedificavit Rama ut non possit quispiam egredi vel ingredi de parte Asa regis Iudae
1KGS|15|18|tollens itaque Asa omne argentum et aurum quod remanserat in thesauris domus Domini et in thesauris domus regiae dedit illud in manu servorum suorum et misit ad Benadad filium Tabremmon filii Ezion regem Syriae qui habitabat in Damasco dicens
1KGS|15|19|foedus est inter me et te et inter patrem meum et patrem tuum ideo misi tibi munera argentum et aurum et peto ut venias et irritum facias foedus quod habes cum Baasa rege Israhel et recedat a me
1KGS|15|20|adquiescens Benadad regi Asa misit principes exercitus sui in civitates Israhel et percusserunt Ahion et Dan et Abel domum Maacha et universam Cenneroth omnem scilicet terram Nepthalim
1KGS|15|21|quod cum audisset Baasa intermisit aedificare Rama et reversus est in Thersa
1KGS|15|22|rex autem Asa nuntium misit in omnem Iudam nemo sit excusatus et tulerunt lapides Rama et ligna eius quibus aedificaverat Baasa et extruxit de eis rex Asa Gaba Beniamin et Maspha
1KGS|15|23|reliqua autem omnium sermonum Asa et universae fortitudines eius et cuncta quae fecit et civitates quas extruxit nonne haec scripta sunt in libro verborum dierum regum Iuda verumtamen in tempore senectutis suae doluit pedes
1KGS|15|24|et dormivit cum patribus suis et sepultus est cum eis in civitate David patris sui regnavitque Iosaphat filius eius pro eo
1KGS|15|25|Nadab vero filius Hieroboam regnavit super Israhel anno secundo Asa regis Iuda regnavitque super Israhel duobus annis
1KGS|15|26|et fecit quod malum est in conspectu Domini et ambulavit in viis patris sui et in peccatis eius quibus peccare fecit Israhel
1KGS|15|27|insidiatus est autem ei Baasa filius Ahia de domo Isachar et percussit eum in Gebbethon quae est urbs Philisthinorum siquidem Nadab et omnis Israhel obsidebant Gebbethon
1KGS|15|28|interfecit igitur illum Baasa in anno tertio Asa regis Iuda et regnavit pro eo
1KGS|15|29|cumque regnasset percussit omnem domum Hieroboam non dimisit ne unam quidem animam de semine eius donec deleret eum iuxta verbum Domini quod locutus fuerat in manu servi sui Ahiae Silonitis
1KGS|15|30|propter peccata Hieroboam quae peccaverat et quibus peccare fecerat Israhel et propter delictum quo inritaverat Dominum Deum Israhel
1KGS|15|31|reliqua autem sermonum Nadab et omnia quae operatus est nonne haec scripta sunt in libro verborum dierum regum Israhel
1KGS|15|32|fuitque bellum inter Asa et Baasa regem Israhel cunctis diebus eorum
1KGS|15|33|anno tertio Asa regis Iuda regnavit Baasa filius Ahia super omnem Israhel in Thersa viginti quattuor annis
1KGS|15|34|et fecit malum coram Domino ambulavitque in via Hieroboam et in peccatis eius quibus peccare fecit Israhel
1KGS|16|1|factus est autem sermo Domini ad Hieu filium Anani contra Baasa dicens
1KGS|16|2|pro eo quod exaltavi te de pulvere et posui ducem super populum meum Israhel tu autem ambulasti in via Hieroboam et peccare fecisti populum meum Israhel ut me inritares in peccatis eorum
1KGS|16|3|ecce ego demetam posteriora Baasa et posteriora domus eius et faciam domum tuam sicut domum Hieroboam filii Nabath
1KGS|16|4|qui mortuus fuerit de Baasa in civitate comedent eum canes et qui mortuus fuerit ex eo in regione comedent eum volucres caeli
1KGS|16|5|reliqua autem sermonum Baasa et quaecumque fecit et proelia eius nonne haec scripta sunt in libro verborum dierum regum Israhel
1KGS|16|6|dormivit ergo Baasa cum patribus suis sepultusque est in Thersa et regnavit Hela filius eius pro eo
1KGS|16|7|cum autem in manu Hieu filii Anani prophetae verbum Domini factum esset contra Baasa et contra domum eius et contra omne malum quod fecerat coram Domino ad inritandum eum in operibus manuum suarum ut fieret sicut domus Hieroboam ob hanc causam occidit eum
1KGS|16|8|anno vicesimo sexto Asa regis Iuda regnavit Hela filius Baasa super Israhel in Thersa duobus annis
1KGS|16|9|et rebellavit contra eum servus suus Zamri dux mediae partis equitum erat autem Hela in Thersa bibens et temulentus in domo Arsa praefecti Thersa
1KGS|16|10|inruens ergo Zamri percussit et occidit eum anno vicesimo septimo Asa regis Iuda et regnavit pro eo
1KGS|16|11|cumque regnasset et sedisset super solium eius percussit omnem domum Baasa et non dereliquit ex eo mingentem ad parietem et propinquos et amicos eius
1KGS|16|12|delevitque Zamri omnem domum Baasa iuxta verbum Domini quod locutus fuerat ad Baasa in manu Hieu prophetae
1KGS|16|13|propter universa peccata Baasa et peccata Hela filii eius qui peccaverunt et peccare fecerunt Israhel provocantes Dominum Deum Israhel in vanitatibus suis
1KGS|16|14|reliqua autem sermonum Hela et omnia quae fecit nonne haec scripta sunt in libro verborum dierum regum Israhel
1KGS|16|15|anno vicesimo et septimo Asa regis Iuda regnavit Zamri septem diebus in Thersa porro exercitus obsidebat Gebbethon urbem Philisthinorum
1KGS|16|16|cumque audisset rebellasse Zamri et occidisse regem fecit sibi regem omnis Israhel Amri qui erat princeps militiae super Israhel in die illa in castris
1KGS|16|17|ascendit ergo Amri et omnis Israhel cum eo de Gebbethon et obsidebant Thersa
1KGS|16|18|videns autem Zamri quod expugnanda esset civitas ingressus est palatium et succendit secum domum regiam et mortuus est
1KGS|16|19|in peccatis suis quae peccaverat faciens malum coram Domino et ambulans in via Hieroboam et in peccato eius quo fecit peccare Israhel
1KGS|16|20|reliqua autem sermonum Zamri et insidiarum eius et tyrannidis nonne haec scripta sunt in libro verborum dierum regum Israhel
1KGS|16|21|tunc divisus est populus Israhel in duas partes media pars populi sequebatur Thebni filium Gineth ut constitueret eum regem et media pars Amri
1KGS|16|22|praevaluit autem populus qui erat cum Amri populo qui sequebatur Thebni filium Gineth mortuusque est Thebni et regnavit Amri
1KGS|16|23|anno tricesimo primo Asa regis Iuda regnavit Amri super Israhel duodecim annis in Thersa regnavit sex annis
1KGS|16|24|emitque montem Samariae a Somer duobus talentis argenti et aedificavit eam et vocavit nomen civitatis quam extruxerat nomine Somer domini montis Samariae
1KGS|16|25|fecit autem Amri malum in conspectu Domini et operatus est nequiter super omnes qui fuerant ante eum
1KGS|16|26|ambulavitque in omni via Hieroboam filii Nabath et in peccatis eius quibus peccare fecerat Israhel ut inritaret Dominum Deum Israhel in vanitatibus suis
1KGS|16|27|reliqua autem sermonum Amri et proelia eius quae gessit nonne haec scripta sunt in libro verborum dierum regum Israhel
1KGS|16|28|et dormivit Amri cum patribus suis et sepultus est in Samaria regnavitque Ahab filius eius pro eo
1KGS|16|29|Ahab vero filius Amri regnavit super Israhel anno tricesimo octavo Asa regis Iuda et regnavit Ahab filius Amri super Israhel in Samaria viginti et duobus annis
1KGS|16|30|et fecit Ahab filius Amri malum in conspectu Domini super omnes qui fuerunt ante eum
1KGS|16|31|nec suffecit ei ut ambularet in peccatis Hieroboam filii Nabath insuper duxit uxorem Hiezabel filiam Ethbaal regis Sidoniorum et abiit et servivit Baal et adoravit eum
1KGS|16|32|et posuit aram Baal in templo Baal quod aedificaverat in Samaria
1KGS|16|33|et plantavit lucum et addidit Ahab in opere suo inritans Dominum Deum Israhel super omnes reges Israhel qui fuerant ante eum
1KGS|16|34|in diebus eius aedificavit Ahiel de Bethel Hiericho in Abiram primitivo suo fundavit eam et in Segub novissimo suo posuit portas eius iuxta verbum Domini quod locutus fuerat in manu Iosue filii Nun
1KGS|17|1|et dixit Helias Thesbites de habitatoribus Galaad ad Ahab vivit Dominus Deus Israhel in cuius conspectu sto si erit annis his ros et pluvia nisi iuxta oris mei verba
1KGS|17|2|et factum est verbum Domini ad eum dicens
1KGS|17|3|recede hinc et vade contra orientem et abscondere in torrente Charith qui est contra Iordanem
1KGS|17|4|et ibi de torrente bibes corvisque praecepi ut pascant te ibi
1KGS|17|5|abiit ergo et fecit iuxta verbum Domini cumque abisset sedit in torrente Charith qui est contra Iordanem
1KGS|17|6|corvi quoque deferebant panem et carnes mane similiter panem et carnes vesperi et bibebat de torrente
1KGS|17|7|post dies autem siccatus est torrens non enim pluerat super terram
1KGS|17|8|factus est igitur sermo Domini ad eum dicens
1KGS|17|9|surge et vade in Sareptha Sidoniorum et manebis ibi praecepi enim ibi mulieri viduae ut pascat te
1KGS|17|10|surrexit et abiit Sareptham cumque venisset ad portam civitatis apparuit ei mulier vidua colligens ligna et vocavit eam dixitque da mihi paululum aquae in vase ut bibam
1KGS|17|11|cumque illa pergeret ut adferret clamavit post tergum eius dicens adfer mihi obsecro et buccellam panis in manu tua
1KGS|17|12|quae respondit vivit Dominus Deus tuus quia non habeo panem nisi quantum pugillus capere potest farinae in hydria et paululum olei in lecytho en colligo duo ligna ut ingrediar et faciam illud mihi et filio meo ut comedamus et moriamur
1KGS|17|13|ad quam Helias ait noli timere sed vade et fac sicut dixisti verumtamen mihi primum fac de ipsa farinula subcinericium panem parvulum et adfer ad me tibi autem et filio tuo facies postea
1KGS|17|14|haec autem dicit Dominus Deus Israhel hydria farinae non deficiet nec lecythus olei minuetur usque ad diem in qua daturus est Dominus pluviam super faciem terrae
1KGS|17|15|quae abiit et fecit iuxta verbum Heliae et comedit ipse et illa et domus eius et ex illa die
1KGS|17|16|hydria farinae non defecit et lecythus olei non est inminutus iuxta verbum Domini quod locutus fuerat in manu Heliae
1KGS|17|17|factum est autem post verba haec aegrotavit filius mulieris matris familiae et erat languor fortis nimis ita ut non remaneret in eo halitus
1KGS|17|18|dixit ergo ad Heliam quid mihi et tibi vir Dei ingressus es ad me ut rememorarentur iniquitates meae et interficeres filium meum
1KGS|17|19|et ait ad eam da mihi filium tuum tulitque eum de sinu illius et portavit in cenaculum ubi ipse manebat et posuit super lectulum suum
1KGS|17|20|et clamavit ad Dominum et dixit Domine Deus meus etiamne viduam apud quam ego utcumque sustentor adflixisti ut interficeres filium eius
1KGS|17|21|et expandit se atque mensus est super puerum tribus vicibus clamavitque ad Dominum et ait Domine Deus meus revertatur oro anima pueri huius in viscera eius
1KGS|17|22|exaudivit Dominus vocem Heliae et reversa est anima pueri intra eum et revixit
1KGS|17|23|tulitque Helias puerum et deposuit eum de cenaculo in inferiorem domum et tradidit matri suae et ait illi en vivit filius tuus
1KGS|17|24|dixitque mulier ad Heliam nunc in isto cognovi quoniam vir Dei es tu et verbum Domini in ore tuo verum est
1KGS|18|1|post dies multos verbum Domini factum est ad Heliam in anno tertio dicens vade et ostende te Ahab ut dem pluviam super faciem terrae
1KGS|18|2|ivit ergo Helias ut ostenderet se Ahab erat autem fames vehemens in Samaria
1KGS|18|3|vocavitque Ahab Abdiam dispensatorem domus suae Abdias autem timebat Dominum valde
1KGS|18|4|nam cum interficeret Hiezabel prophetas Domini tulit ille centum prophetas et abscondit eos quinquagenos in speluncis et pavit eos pane et aqua
1KGS|18|5|dixit ergo Ahab ad Abdiam vade in terram ad universos fontes aquarum et in cunctas valles si forte invenire possimus herbam et salvare equos et mulos et non penitus iumenta intereant
1KGS|18|6|diviseruntque sibi regiones ut circuirent eas Ahab ibat per viam unam et Abdias per viam alteram seorsum
1KGS|18|7|cumque esset Abdias in via Helias occurrit ei qui cum cognovisset eum cecidit super faciem suam et ait num tu es domine mi Helias
1KGS|18|8|cui ille respondit ego vade dic domino tuo adest Helias
1KGS|18|9|et ille quid peccavi inquit quoniam trades me servum tuum in manu Ahab ut interficiat me
1KGS|18|10|vivit Dominus Deus tuus non est gens aut regnum quo non miserit dominus meus te requirens et respondentibus cunctis non est hic adiuravit regna singula et gentes eo quod minime repperireris
1KGS|18|11|et nunc dicis mihi vade et dic domino tuo adest Helias
1KGS|18|12|cumque recessero a te spiritus Domini asportabit te in locum quem ego ignoro ingressus nuntiabo Ahab et non inveniet te et interficiet me servus autem tuus timet Dominum ab infantia sua
1KGS|18|13|numquid non indicatum est tibi domino meo quid fecerim cum interficeret Hiezabel prophetas Domini quod absconderim de prophetis Domini centum viros quinquagenos et quinquagenos in speluncis et paverim eos pane et aqua
1KGS|18|14|et nunc tu dicis vade et dic domino tuo adest Helias ut interficiat me
1KGS|18|15|dixit Helias vivit Dominus exercituum ante cuius vultum sto quia hodie apparebo ei
1KGS|18|16|abiit ergo Abdias in occursum Ahab et indicavit ei venitque Ahab in occursum Heliae
1KGS|18|17|et cum vidisset eum ait tune es ille qui conturbas Israhel
1KGS|18|18|et ille ait non turbavi Israhel sed tu et domus patris tui qui dereliquistis mandata Domini et secuti estis Baalim
1KGS|18|19|verumtamen nunc mitte et congrega ad me universum Israhel in monte Carmeli et prophetas Baal quadringentos quinquaginta prophetasque lucorum quadringentos qui comedunt de mensa Hiezabel
1KGS|18|20|misit Ahab ad omnes filios Israhel et congregavit prophetas in monte Carmeli
1KGS|18|21|accedens autem Helias ad omnem populum ait usquequo claudicatis in duas partes si Dominus est Deus sequimini eum si autem Baal sequimini illum et non respondit ei populus verbum
1KGS|18|22|et ait rursum Helias ad populum ego remansi propheta Domini solus prophetae autem Baal quadringenti et quinquaginta viri sunt
1KGS|18|23|dentur nobis duo boves et illi eligant bovem unum et in frusta caedentes ponant super ligna ignem autem non subponant et ego faciam bovem alterum et inponam super ligna ignemque non subponam
1KGS|18|24|invocate nomina deorum vestrorum et ego invocabo nomen Domini et deus qui exaudierit per ignem ipse sit Deus respondens omnis populus ait optima propositio
1KGS|18|25|dixit ergo Helias prophetis Baal eligite vobis bovem unum et facite primi quia vos plures estis et invocate nomina deorum vestrorum ignemque non subponatis
1KGS|18|26|qui cum tulissent bovem quem dederat eis fecerunt et invocabant nomen Baal de mane usque ad meridiem dicentes Baal exaudi nos et non erat vox nec qui responderet transiliebantque altare quod fecerant
1KGS|18|27|cumque esset iam meridies inludebat eis Helias dicens clamate voce maiore deus enim est et forsitan loquitur aut in diversorio est aut in itinere aut certe dormit ut excitetur
1KGS|18|28|clamabant ergo voce magna et incidebant se iuxta ritum suum cultris et lanceolis donec perfunderentur sanguine
1KGS|18|29|postquam autem transiit meridies et illis prophetantibus venerat tempus quo sacrificium offerri solet nec audiebatur vox neque aliquis respondebat nec adtendebat orantes
1KGS|18|30|dixit Helias omni populo venite ad me et accedente ad se populo curavit altare Domini quod destructum fuerat
1KGS|18|31|et tulit duodecim lapides iuxta numerum tribuum filiorum Iacob ad quem factus est sermo Domini dicens Israhel erit nomen tuum
1KGS|18|32|et aedificavit lapidibus altare in nomine Domini fecitque aquaeductum quasi per duas aratiunculas in circuitu altaris
1KGS|18|33|et conposuit ligna divisitque per membra bovem et posuit super ligna
1KGS|18|34|et ait implete quattuor hydrias aqua et fundite super holocaustum et super ligna rursumque dixit etiam secundo hoc facite qui cum fecissent et secundo ait etiam tertio id ipsum facite feceruntque et tertio
1KGS|18|35|et currebant aquae circa altare et fossa aquaeductus repleta est
1KGS|18|36|cumque iam tempus esset ut offerretur holocaustum accedens Helias propheta ait Domine Deus Abraham Isaac et Israhel hodie ostende quia tu es Deus Israhel et ego servus tuus et iuxta praeceptum tuum feci omnia verba haec
1KGS|18|37|exaudi me Domine exaudi me ut discat populus iste quia tu es Dominus Deus et tu convertisti cor eorum iterum
1KGS|18|38|cecidit autem ignis Domini et voravit holocaustum et ligna et lapides pulverem quoque et aquam quae erat in aquaeductu lambens
1KGS|18|39|quod cum vidisset omnis populus cecidit in faciem suam et ait Dominus ipse est Deus Dominus ipse est Deus
1KGS|18|40|dixitque Helias ad eos adprehendite prophetas Baal et ne unus quidem fugiat ex eis quos cum conprehendissent duxit eos Helias ad torrentem Cison et interfecit eos ibi
1KGS|18|41|et ait Helias ad Ahab ascende comede et bibe quia sonus multae pluviae est
1KGS|18|42|ascendit Ahab ut comederet et biberet Helias autem ascendit in vertice Carmeli et pronus in terram posuit faciem inter genua sua
1KGS|18|43|et dixit ad puerum suum ascende et prospice contra mare qui cum ascendisset et contemplatus esset ait non est quicquam et rursum ait illi revertere septem vicibus
1KGS|18|44|in septima autem vice ecce nubicula parva quasi vestigium hominis ascendebat de mari qui ait ascende et dic Ahab iunge et descende ne occupet te pluvia
1KGS|18|45|cumque se verterent huc atque illuc ecce caeli contenebrati sunt et nubes et ventus et facta est pluvia grandis ascendens itaque Ahab abiit in Hiezrahel
1KGS|18|46|et manus Domini facta est super Heliam accinctisque lumbis currebat ante Ahab donec veniret in Hiezrahel
1KGS|19|1|nuntiavit autem Ahab Hiezabel omnia quae fecerat Helias et quomodo occidisset universos prophetas gladio
1KGS|19|2|misitque Hiezabel nuntium ad Heliam dicens haec mihi faciant dii et haec addant nisi hac hora cras posuero animam tuam sicut animam unius ex illis
1KGS|19|3|timuit ergo Helias et surgens abiit quocumque eum ferebat voluntas venitque in Bersabee Iuda et dimisit ibi puerum suum
1KGS|19|4|et perrexit in desertum via unius diei cumque venisset et sederet subter unam iuniperum petivit animae suae ut moreretur et ait sufficit mihi Domine tolle animam meam neque enim melior sum quam patres mei
1KGS|19|5|proiecitque se et obdormivit in umbra iuniperi et ecce angelus tetigit eum et dixit illi surge comede
1KGS|19|6|respexit et ecce ad caput suum subcinericius panis et vas aquae comedit ergo et bibit et rursum obdormivit
1KGS|19|7|reversusque est angelus Domini secundo et tetigit eum dixitque illi surge comede grandis enim tibi restat via
1KGS|19|8|qui cum surrexisset comedit et bibit et ambulavit in fortitudine cibi illius quadraginta diebus et quadraginta noctibus usque ad montem Dei Horeb
1KGS|19|9|cumque venisset illuc mansit in spelunca et ecce sermo Domini ad eum dixitque illi quid hic agis Helia
1KGS|19|10|at ille respondit zelo zelatus sum pro Domino Deo exercituum quia dereliquerunt pactum Domini filii Israhel altaria tua destruxerunt et prophetas tuos occiderunt gladio et derelictus sum ego solus et quaerunt animam meam ut auferant eam
1KGS|19|11|et ait ei egredere et sta in monte coram Domino et ecce Dominus transit et spiritus grandis et fortis subvertens montes et conterens petras ante Dominum non in spiritu Dominus et post spiritum commotio non in commotione Dominus
1KGS|19|12|et post commotionem ignis non in igne Dominus et post ignem sibilus aurae tenuis
1KGS|19|13|quod cum audisset Helias operuit vultum suum pallio et egressus stetit in ostio speluncae et ecce vox ad eum dicens quid agis hic Helia
1KGS|19|14|et ille respondit zelo zelatus sum pro Domino Deo exercituum quia dereliquerunt pactum tuum filii Israhel altaria tua destruxerunt et prophetas tuos occiderunt gladio et derelictus sum ego solus et quaerunt animam meam ut auferant eam
1KGS|19|15|et ait Dominus ad eum vade et revertere in viam tuam per desertum in Damascum cumque perveneris ungues Azahel regem super Syriam
1KGS|19|16|et Hieu filium Namsi ungues regem super Israhel Heliseum autem filium Saphat qui est de Abelmaula ungues prophetam pro te
1KGS|19|17|et erit quicumque fugerit gladium Azahel occidet eum Hieu et qui fugerit gladium Hieu interficiet eum Heliseus
1KGS|19|18|et derelinquam mihi in Israhel septem milia universorum genua quae non sunt incurvata Baal et omne os quod non adoravit eum osculans manum
1KGS|19|19|profectus ergo inde repperit Heliseum filium Saphat arantem duodecim iugis boum et ipse in duodecim arantibus unus erat cumque venisset Helias ad eum misit pallium suum super illum
1KGS|19|20|qui statim relictis bubus cucurrit post Heliam et ait osculer oro te patrem meum et matrem meam et sic sequar te dixitque ei vade et revertere quod enim meum erat feci tibi
1KGS|19|21|reversus autem ab eo tulit par boum et mactavit illud et in aratro boum coxit carnes et dedit populo et comederunt consurgensque abiit et secutus est Heliam et ministrabat ei
1KGS|20|1|porro Benadad rex Syriae congregavit omnem exercitum suum et triginta et duos reges secum et equos et currus et ascendens pugnabat contra Samariam et obsidebat eam
1KGS|20|2|mittensque nuntios ad Ahab regem Israhel in civitatem
1KGS|20|3|ait haec dicit Benadad argentum tuum et aurum tuum meum est et uxores tuae et filii tui optimi mei sunt
1KGS|20|4|responditque rex Israhel iuxta verbum tuum domine mi rex tuus sum ego et omnia mea
1KGS|20|5|revertentesque nuntii dixerunt haec dicit Benadad qui misit nos ad te argentum tuum et aurum tuum et uxores tuas et filios tuos dabis mihi
1KGS|20|6|cras igitur hac eadem hora mittam servos meos ad te et scrutabuntur domum tuam et domum servorum tuorum et omne quod eis placuerit ponent in manibus suis et auferent
1KGS|20|7|vocavit autem rex Israhel omnes seniores terrae et ait animadvertite et videte quoniam insidietur nobis misit enim ad me pro uxoribus meis et filiis et pro argento et auro et non abnui
1KGS|20|8|dixeruntque omnes maiores natu et universus populus ad eum non audias neque adquiescas illi
1KGS|20|9|respondit itaque nuntiis Benadad dicite domino meo regi omnia propter quae misisti ad me servum tuum initio faciam hanc autem rem facere non possum
1KGS|20|10|reversique nuntii rettulerunt ei qui remisit et ait haec faciant mihi dii et haec addant si suffecerit pulvis Samariae pugillis omnis populi qui sequitur me
1KGS|20|11|et respondens rex Israhel ait dicite ei ne glorietur accinctus aeque ut discinctus
1KGS|20|12|factum est autem cum audisset verbum istud bibebat ipse et reges in umbraculis et ait servis suis circumdate civitatem et circumdederunt eam
1KGS|20|13|et ecce propheta unus accedens ad Ahab regem Israhel ait haec dicit Dominus certe vidisti omnem multitudinem hanc nimiam ecce ego tradam eam in manu tua hodie ut scias quia ego sum Dominus
1KGS|20|14|et ait Ahab per quem dixitque ei haec dicit Dominus per pedisequos principum provinciarum et ait quis incipiet proeliari et ille dixit tu
1KGS|20|15|recensuit ergo pueros principum provinciarum et repperit numerum ducentorum triginta duum et post eos recensuit populum omnes filios Israhel septem milia
1KGS|20|16|et egressi sunt meridie Benadad autem bibebat temulentus in umbraculo suo et reges triginta duo cum eo qui ad auxilium eius venerant
1KGS|20|17|egressi sunt autem pueri principum provinciarum in prima fronte misit itaque Benadad qui nuntiaverunt ei dicentes viri egressi sunt de Samaria
1KGS|20|18|at ille sive ait pro pace veniunt adprehendite eos vivos sive ut proelientur vivos eos capite
1KGS|20|19|egressi sunt ergo pueri principum provinciarum ac reliquus exercitus sequebatur
1KGS|20|20|et percussit unusquisque virum qui contra se venerat fugeruntque Syri et persecutus est eos Israhel fugit quoque Benadad rex Syriae in equo cum equitibus
1KGS|20|21|necnon et egressus rex Israhel percussit equos et currus et percussit Syriam plaga magna
1KGS|20|22|accedens autem propheta ad regem Israhel dixit ei vade et confortare et scito et vide quid facias sequenti enim anno rex Syriae ascendet contra te
1KGS|20|23|servi vero regis Syriae dixerunt ei dii montium sunt dii eorum ideo superaverunt nos sed melius est ut pugnemus contra eos in campestribus et obtinebimus eos
1KGS|20|24|tu ergo verbum hoc fac amove reges singulos ab exercitu suo et pone principes pro eis
1KGS|20|25|et instaura numerum militum qui ceciderunt de tuis et equos secundum equos pristinos et currus secundum currus quos ante habuisti et pugnabimus contra eos in campestribus et videbis quod obtinebimus eos credidit consilio eorum et fecit ita
1KGS|20|26|igitur postquam annus transierat recensuit Benadad Syros et ascendit in Afec ut pugnaret contra Israhel
1KGS|20|27|porro filii Israhel recensiti sunt et acceptis cibariis profecti ex adverso castraque metati contra eos quasi duo parvi greges caprarum Syri autem repleverunt terram
1KGS|20|28|et accedens unus vir Dei dixit ad regem Israhel haec dicit Dominus quia dixerunt Syri deus montium est Dominus et non est deus vallium dabo omnem multitudinem grandem hanc in manu tua et scietis quia ego Dominus
1KGS|20|29|dirigebant septem diebus ex adverso hii atque illi acies septima autem die commissum est bellum percusseruntque filii Israhel de Syris centum milia peditum in die una
1KGS|20|30|fugerunt autem qui remanserant in Afec in civitatem et cecidit murus super viginti septem milia hominum qui remanserant porro Benadad fugiens ingressus est civitatem in cubiculum quod erat intra cubiculum
1KGS|20|31|dixeruntque ei servi sui ecce audivimus quod reges domus Israhel clementes sint ponamus itaque saccos in lumbis nostris et funiculos in capitibus nostris et egrediamur ad regem Israhel forsitan salvabit animas nostras
1KGS|20|32|accinxerunt saccis lumbos suos et posuerunt funes in capitibus veneruntque ad regem Israhel et dixerunt servus tuus Benadad dicit vivat oro te anima mea et ille ait si adhuc vivit frater meus est
1KGS|20|33|quod acceperunt viri pro omine et festinantes rapuerunt verbum ex ore eius atque dixerunt frater tuus Benadad et dixit eis ite et adducite eum egressus est ergo ad eum Benadad et levavit eum in currum suum
1KGS|20|34|qui dixit ei civitates quas tulit pater meus a patre tuo reddam et plateas fac tibi in Damasco sicut fecit pater meus in Samaria et ego foederatus recedam a te pepigit ergo foedus et dimisit eum
1KGS|20|35|tunc vir quidam de filiis prophetarum dixit ad socium suum in sermone Domini percute me at ille noluit percutere
1KGS|20|36|cui ait quia noluisti audire vocem Domini ecce recedes a me et percutiet te leo cumque paululum recessisset ab eo invenit eum leo atque percussit
1KGS|20|37|sed et alterum conveniens virum dixit ad eum percute me qui percussit eum et vulneravit
1KGS|20|38|abiit ergo propheta et occurrit regi in via et mutavit aspersione pulveris os et oculos suos
1KGS|20|39|cumque rex transiret clamavit ad regem et ait servus tuus egressus est ad proeliandum comminus cumque fugisset vir unus adduxit eum quidam ad me et ait custodi virum istum qui si lapsus fuerit erit anima tua pro anima eius aut talentum argenti adpendes
1KGS|20|40|dum autem ego turbatus huc illucque me verterem subito non conparuit et ait rex Israhel ad eum hoc est iudicium tuum quod ipse decrevisti
1KGS|20|41|at ille statim abstersit pulverem de facie sua et cognovit eum rex Israhel quod esset de prophetis
1KGS|20|42|qui ait ad eum haec dicit Dominus quia dimisisti virum dignum morte de manu tua erit anima tua pro anima eius et populus tuus pro populo eius
1KGS|20|43|reversus est igitur rex Israhel in domum suam audire contemnens et furibundus venit Samariam
1KGS|21|1|post verba autem haec vinea erat Naboth Hiezrahelitae qui erat in Hiezrahel iuxta palatium Ahab regis Samariae
1KGS|21|2|locutus est ergo Ahab ad Naboth dicens da mihi vineam tuam ut faciam mihi hortum holerum quia vicina est et prope domum meam daboque tibi pro ea vineam meliorem aut si tibi commodius putas argenti pretium quanto digna est
1KGS|21|3|cui respondit Naboth propitius mihi sit Dominus ne dem hereditatem patrum meorum tibi
1KGS|21|4|venit ergo Ahab in domum suam indignans et frendens super verbo quod locutus fuerat ad eum Naboth Hiezrahelites dicens non do tibi hereditatem patrum meorum et proiciens se in lectulum suum avertit faciem ad parietem et non comedit panem
1KGS|21|5|ingressa est autem ad eum Hiezabel uxor sua dixitque ei quid est hoc unde anima tua contristata est et quare non comedis panem
1KGS|21|6|qui respondit ei locutus sum Naboth Hiezrahelitae et dixi ei da mihi vineam tuam accepta pecunia aut si tibi placet dabo tibi vineam pro ea et ille ait non do tibi vineam meam
1KGS|21|7|dixit ergo ad eum Hiezabel uxor eius grandis auctoritatis es et bene regis regnum Israhel surge et comede panem et aequo esto animo ego dabo tibi vineam Naboth Hiezrahelitae
1KGS|21|8|scripsit itaque litteras ex nomine Ahab et signavit eas anulo eius et misit ad maiores natu et ad optimates qui erant in civitate eius et habitabant cum Naboth
1KGS|21|9|litterarum autem erat ista sententia praedicate ieiunium et sedere facite Naboth inter primos populi
1KGS|21|10|et submittite duos viros filios Belial contra eum et falsum testimonium dicant benedixit Deum et regem et educite eum et lapidate sicque moriatur
1KGS|21|11|fecerunt ergo cives eius maiores natu et optimates qui habitabant cum eo in urbe sicut praeceperat eis Hiezabel et sicut scriptum erat in litteris quas miserat ad eos
1KGS|21|12|praedicaverunt ieiunium et sedere fecerunt Naboth inter primos populi
1KGS|21|13|et adductis duobus viris filiis diaboli fecerunt eos sedere contra eum at illi scilicet ut viri diabolici dixerunt contra eum testimonium coram multitudine benedixit Naboth Deo et regi quam ob rem eduxerunt eum extra civitatem et lapidibus interfecerunt
1KGS|21|14|miseruntque ad Hiezabel dicentes lapidatus est Naboth et mortuus est
1KGS|21|15|factum est autem cum audisset Hiezabel lapidatum Naboth et mortuum locuta est ad Ahab surge posside vineam Naboth Hiezrahelitae qui noluit tibi adquiescere et dare eam accepta pecunia non enim vivit Naboth sed mortuus est
1KGS|21|16|quod cum audisset Ahab mortuum videlicet Naboth surrexit et descendebat in vineam Naboth Hiezrahelitae ut possideret eam
1KGS|21|17|factus est igitur sermo Domini ad Heliam Thesbiten dicens
1KGS|21|18|surge et descende in occursum Ahab regis Israhel qui est in Samaria ecce ad vineam Naboth descendit ut possideat eam
1KGS|21|19|et loqueris ad eum dicens haec dicit Dominus occidisti insuper et possedisti et post haec addes haec dicit Dominus in loco hoc in quo linxerunt canes sanguinem Naboth lambent tuum quoque sanguinem
1KGS|21|20|et ait Ahab ad Heliam num invenisti me inimice mee qui dixit inveni eo quod venundatus sis ut faceres malum in conspectu Domini
1KGS|21|21|ecce ego inducam super te malum et demetam posteriora tua et interficiam de Ahab mingentem ad parietem et clausum et ultimum in Israhel
1KGS|21|22|et dabo domum tuam sicut domum Hieroboam filii Nabath et sicut domum Baasa filii Ahia quia egisti ut me ad iracundiam provocares et peccare fecisti Israhel
1KGS|21|23|sed et de Hiezabel locutus est Dominus dicens canes comedent Hiezabel in agro Hiezrahel
1KGS|21|24|si mortuus fuerit Ahab in civitate comedent eum canes si autem mortuus fuerit in agro comedent eum volucres caeli
1KGS|21|25|igitur non fuit alter talis ut Ahab qui venundatus est ut faceret malum in conspectu Domini concitavit enim eum Hiezabel uxor sua
1KGS|21|26|et abominabilis effectus est in tantum ut sequeretur idola quae fecerant Amorrei quos consumpsit Dominus a facie filiorum Israhel
1KGS|21|27|itaque cum audisset Ahab sermones istos scidit vestem suam et operuit cilicio carnem suam ieiunavitque et dormivit in sacco et ambulabat dimisso capite
1KGS|21|28|factus est autem sermo Domini ad Heliam Thesbiten dicens
1KGS|21|29|nonne vidisti humiliatum Ahab coram me quia igitur humiliatus est mei causa non inducam malum in diebus eius sed in diebus filii sui inferam malum domui eius
1KGS|22|1|transierunt igitur tres anni absque bello inter Syriam et Israhel
1KGS|22|2|in anno autem tertio descendit Iosaphat rex Iuda ad regem Israhel
1KGS|22|3|dixitque rex Israhel ad servos suos ignoratis quod nostra sit Ramoth Galaad et neglegimus tollere eam de manu regis Syriae
1KGS|22|4|et ait ad Iosaphat veniesne mecum ad proeliandum in Ramoth Galaad
1KGS|22|5|dixitque Iosaphat ad regem Israhel sicut ego sum ita et tu populus meus et populus tuus unum sunt et equites mei et equites tui dixitque Iosaphat ad regem Israhel quaere oro te hodie sermonem Domini
1KGS|22|6|congregavit ergo rex Israhel prophetas quadringentos circiter viros et ait ad eos ire debeo in Ramoth Galaad ad bellandum an quiescere qui responderunt ascende et dabit Dominus in manu regis
1KGS|22|7|dixit autem Iosaphat non est hic propheta Domini quispiam ut interrogemus per eum
1KGS|22|8|et ait rex Israhel ad Iosaphat remansit vir unus per quem possimus interrogare Dominum sed ego odi eum quia non prophetat mihi bonum sed malum Micheas filius Hiemla cui Iosaphat ait ne loquaris ita rex
1KGS|22|9|vocavit ergo rex Israhel eunuchum quendam et dixit ei festina adducere Micheam filium Hiemla
1KGS|22|10|rex autem Israhel et Iosaphat rex Iuda sedebat unusquisque in solio suo vestiti cultu regio in area iuxta ostium portae Samariae et universi prophetae prophetabant in conspectu eorum
1KGS|22|11|fecit quoque sibi Sedecias filius Chanaan cornua ferrea et ait haec dicit Dominus his ventilabis Syriam donec deleas eam
1KGS|22|12|omnesque prophetae similiter prophetabant dicentes ascende in Ramoth Galaad et vade prospere et tradet Dominus in manu regis
1KGS|22|13|nuntius vero qui ierat ut vocaret Micheam locutus est ad eum dicens ecce sermones prophetarum ore uno bona regi praedicant sit ergo et sermo tuus similis eorum et loquere bona
1KGS|22|14|cui Micheas ait vivit Dominus quia quodcumque dixerit mihi Dominus hoc loquar
1KGS|22|15|venit itaque ad regem et ait illi rex Michea ire debemus in Ramoth Galaad ad proeliandum an cessare cui ille respondit ascende et vade prospere et tradet Dominus in manu regis
1KGS|22|16|dixit autem rex ad eum iterum atque iterum adiuro te ut non loquaris mihi nisi quod verum est in nomine Domini
1KGS|22|17|et ille ait vidi cunctum Israhel dispersum in montibus quasi oves non habentes pastorem et ait Dominus non habent dominum isti revertatur unusquisque in domum suam in pace
1KGS|22|18|dixit ergo rex Israhel ad Iosaphat numquid non dixi tibi quia non prophetat mihi bonum sed semper malum
1KGS|22|19|ille vero addens ait propterea audi sermonem Domini vidi Dominum sedentem super solium suum et omnem exercitum caeli adsistentem ei a dextris et a sinistris
1KGS|22|20|et ait Dominus quis decipiet Ahab regem Israhel ut ascendat et cadat in Ramoth Galaad et dixit unus verba huiuscemodi et alius aliter
1KGS|22|21|egressus est autem spiritus et stetit coram Domino et ait ego decipiam illum cui locutus est Dominus in quo
1KGS|22|22|et ille ait egrediar et ero spiritus mendax in ore omnium prophetarum eius et dixit Dominus decipies et praevalebis egredere et fac ita
1KGS|22|23|nunc igitur ecce dedit Dominus spiritum mendacii in ore omnium prophetarum tuorum qui hic sunt et Dominus locutus est contra te malum
1KGS|22|24|accessit autem Sedecias filius Chanaan et percussit Micheam in maxillam et dixit mene ergo dimisit spiritus Domini et locutus est tibi
1KGS|22|25|et ait Micheas visurus es in die illa quando ingredieris cubiculum intra cubiculum ut abscondaris
1KGS|22|26|et ait rex Israhel tollite Micheam et maneat apud Amon principem civitatis et apud Ioas filium Ammelech
1KGS|22|27|et dicite eis haec dicit rex mittite virum istum in carcerem et sustentate eum pane tribulationis et aqua angustiae donec revertar in pace
1KGS|22|28|dixitque Micheas si reversus fueris in pace non est locutus Dominus in me et ait audite populi omnes
1KGS|22|29|ascendit itaque rex Israhel et Iosaphat rex Iuda in Ramoth Galaad
1KGS|22|30|dixitque rex Israhel ad Iosaphat sume arma et ingredere proelium et induere vestibus tuis porro rex Israhel mutavit habitum et ingressus est bellum
1KGS|22|31|rex autem Syriae praeceperat principibus curruum triginta duobus dicens non pugnabitis contra minorem et maiorem quempiam nisi contra regem Israhel solum
1KGS|22|32|cum ergo vidissent principes curruum Iosaphat suspicati sunt quod ipse esset rex Israhel et impetu facto pugnabant contra eum et exclamavit Iosaphat
1KGS|22|33|intellexeruntque principes curruum quod non esset rex Israhel et cessaverunt ab eo
1KGS|22|34|unus autem quidam tetendit arcum in incertum sagittam dirigens et casu percussit regem Israhel inter pulmonem et stomachum at ille dixit aurigae suo verte manum tuam et eice me de exercitu quia graviter vulneratus sum
1KGS|22|35|commissum est ergo proelium in die illa et rex Israhel stabat in curru suo contra Syros et mortuus est vesperi fluebat autem sanguis plagae in sinum currus
1KGS|22|36|et praeco personuit in universo exercitu antequam sol occumberet dicens unusquisque revertatur in civitatem et in terram suam
1KGS|22|37|mortuus est autem rex et perlatus est Samariam sepelieruntque regem in Samaria
1KGS|22|38|et laverunt currum in piscina Samariae et linxerunt canes sanguinem eius et habenas laverunt iuxta verbum Domini quod locutus fuerat
1KGS|22|39|reliqua vero sermonum Ahab et universa quae fecit et domus eburneae quam aedificavit cunctarumque urbium quas extruxit nonne scripta sunt haec in libro verborum dierum regum Israhel
1KGS|22|40|dormivit ergo Ahab cum patribus suis et regnavit Ohozias filius eius pro eo
1KGS|22|41|Iosaphat filius Asa regnare coeperat super Iudam anno quarto Ahab regis Israhel
1KGS|22|42|triginta quinque annorum erat cum regnare coepisset et viginti et quinque annos regnavit in Hierusalem nomen matris eius Azuba filia Salai
1KGS|22|43|et ambulavit in omni via Asa patris sui et non declinavit ex ea fecitque quod rectum est in conspectu Domini
1KGS|22|44|verumtamen excelsa non abstulit adhuc enim populus sacrificabat et adolebat incensum in excelsis
1KGS|22|45|pacemque habuit Iosaphat cum rege Israhel
1KGS|22|46|reliqua autem verborum Iosaphat et opera eius quae gessit et proelia nonne haec scripta sunt in libro verborum dierum regum Iuda
1KGS|22|47|sed et reliquias effeminatorum qui remanserant in diebus Asa patris eius abstulit de terra
1KGS|22|48|nec erat tunc rex constitutus in Edom
1KGS|22|49|rex vero Iosaphat fecerat classes in mari quae navigarent in Ophir propter aurum et ire non potuerunt quia confractae sunt in Asiongaber
1KGS|22|50|tunc ait Ohozias filius Ahab ad Iosaphat vadant servi mei cum servis tuis in navibus et noluit Iosaphat
1KGS|22|51|dormivitque cum patribus suis et sepultus est cum eis in civitate David patris sui regnavitque Ioram filius eius pro eo
1KGS|22|52|Ohozias autem filius Ahab regnare coeperat super Israhel in Samaria anno septimodecimo Iosaphat regis Iuda regnavitque super Israhel duobus annis
1KGS|22|53|et fecit malum in conspectu Domini et ambulavit in via patris sui et matris suae et in via Hieroboam filii Nabath qui peccare fecit Israhel
1KGS|22|54|servivit quoque Baal et adoravit eum et inritavit Dominum Deum Israhel iuxta omnia quae fecerat pater eius
