LUKE|1|1|Many have undertaken to draw up an account of the things that have been fulfilled among us,
LUKE|1|2|just as they were handed down to us by those who from the first were eyewitnesses and servants of the word.
LUKE|1|3|Therefore, since I myself have carefully investigated everything from the beginning, it seemed good also to me to write an orderly account for you, most excellent Theophilus,
LUKE|1|4|so that you may know the certainty of the things you have been taught.
LUKE|1|5|In the time of Herod king of Judea there was a priest named Zechariah, who belonged to the priestly division of Abijah; his wife Elizabeth was also a descendant of Aaron.
LUKE|1|6|Both of them were upright in the sight of God, observing all the Lord's commandments and regulations blamelessly.
LUKE|1|7|But they had no children, because Elizabeth was barren; and they were both well along in years.
LUKE|1|8|Once when Zechariah's division was on duty and he was serving as priest before God,
LUKE|1|9|he was chosen by lot, according to the custom of the priesthood, to go into the temple of the Lord and burn incense.
LUKE|1|10|And when the time for the burning of incense came, all the assembled worshipers were praying outside.
LUKE|1|11|Then an angel of the Lord appeared to him, standing at the right side of the altar of incense.
LUKE|1|12|When Zechariah saw him, he was startled and was gripped with fear.
LUKE|1|13|But the angel said to him: "Do not be afraid, Zechariah; your prayer has been heard. Your wife Elizabeth will bear you a son, and you are to give him the name John.
LUKE|1|14|He will be a joy and delight to you, and many will rejoice because of his birth,
LUKE|1|15|for he will be great in the sight of the Lord. He is never to take wine or other fermented drink, and he will be filled with the Holy Spirit even from birth.
LUKE|1|16|Many of the people of Israel will he bring back to the Lord their God.
LUKE|1|17|And he will go on before the Lord, in the spirit and power of Elijah, to turn the hearts of the fathers to their children and the disobedient to the wisdom of the righteous--to make ready a people prepared for the Lord."
LUKE|1|18|Zechariah asked the angel, "How can I be sure of this? I am an old man and my wife is well along in years."
LUKE|1|19|The angel answered, "I am Gabriel. I stand in the presence of God, and I have been sent to speak to you and to tell you this good news.
LUKE|1|20|And now you will be silent and not able to speak until the day this happens, because you did not believe my words, which will come true at their proper time."
LUKE|1|21|Meanwhile, the people were waiting for Zechariah and wondering why he stayed so long in the temple.
LUKE|1|22|When he came out, he could not speak to them. They realized he had seen a vision in the temple, for he kept making signs to them but remained unable to speak.
LUKE|1|23|When his time of service was completed, he returned home.
LUKE|1|24|After this his wife Elizabeth became pregnant and for five months remained in seclusion.
LUKE|1|25|"The Lord has done this for me," she said. "In these days he has shown his favor and taken away my disgrace among the people."
LUKE|1|26|In the sixth month, God sent the angel Gabriel to Nazareth, a town in Galilee,
LUKE|1|27|to a virgin pledged to be married to a man named Joseph, a descendant of David. The virgin's name was Mary.
LUKE|1|28|The angel went to her and said, "Greetings, you who are highly favored! The Lord is with you."
LUKE|1|29|Mary was greatly troubled at his words and wondered what kind of greeting this might be.
LUKE|1|30|But the angel said to her, "Do not be afraid, Mary, you have found favor with God.
LUKE|1|31|You will be with child and give birth to a son, and you are to give him the name Jesus.
LUKE|1|32|He will be great and will be called the Son of the Most High. The Lord God will give him the throne of his father David,
LUKE|1|33|and he will reign over the house of Jacob forever; his kingdom will never end."
LUKE|1|34|"How will this be," Mary asked the angel, "since I am a virgin?"
LUKE|1|35|The angel answered, "The Holy Spirit will come upon you, and the power of the Most High will overshadow you. So the holy one to be born will be called the Son of God.
LUKE|1|36|Even Elizabeth your relative is going to have a child in her old age, and she who was said to be barren is in her sixth month.
LUKE|1|37|For nothing is impossible with God."
LUKE|1|38|"I am the Lord's servant," Mary answered. "May it be to me as you have said." Then the angel left her.
LUKE|1|39|At that time Mary got ready and hurried to a town in the hill country of Judea,
LUKE|1|40|where she entered Zechariah's home and greeted Elizabeth.
LUKE|1|41|When Elizabeth heard Mary's greeting, the baby leaped in her womb, and Elizabeth was filled with the Holy Spirit.
LUKE|1|42|In a loud voice she exclaimed: "Blessed are you among women, and blessed is the child you will bear!
LUKE|1|43|But why am I so favored, that the mother of my Lord should come to me?
LUKE|1|44|As soon as the sound of your greeting reached my ears, the baby in my womb leaped for joy.
LUKE|1|45|Blessed is she who has believed that what the Lord has said to her will be accomplished!"
LUKE|1|46|And Mary said: "My soul glorifies the Lord
LUKE|1|47|and my spirit rejoices in God my Savior,
LUKE|1|48|for he has been mindful of the humble state of his servant. From now on all generations will call me blessed,
LUKE|1|49|for the Mighty One has done great things for me--holy is his name.
LUKE|1|50|His mercy extends to those who fear him, from generation to generation.
LUKE|1|51|He has performed mighty deeds with his arm; he has scattered those who are proud in their inmost thoughts.
LUKE|1|52|He has brought down rulers from their thrones but has lifted up the humble.
LUKE|1|53|He has filled the hungry with good things but has sent the rich away empty.
LUKE|1|54|He has helped his servant Israel, remembering to be merciful
LUKE|1|55|to Abraham and his descendants forever, even as he said to our fathers."
LUKE|1|56|Mary stayed with Elizabeth for about three months and then returned home.
LUKE|1|57|When it was time for Elizabeth to have her baby, she gave birth to a son.
LUKE|1|58|Her neighbors and relatives heard that the Lord had shown her great mercy, and they shared her joy.
LUKE|1|59|On the eighth day they came to circumcise the child, and they were going to name him after his father Zechariah,
LUKE|1|60|but his mother spoke up and said, "No! He is to be called John."
LUKE|1|61|They said to her, "There is no one among your relatives who has that name."
LUKE|1|62|Then they made signs to his father, to find out what he would like to name the child.
LUKE|1|63|He asked for a writing tablet, and to everyone's astonishment he wrote, "His name is John."
LUKE|1|64|Immediately his mouth was opened and his tongue was loosed, and he began to speak, praising God.
LUKE|1|65|The neighbors were all filled with awe, and throughout the hill country of Judea people were talking about all these things.
LUKE|1|66|Everyone who heard this wondered about it, asking, "What then is this child going to be?" For the Lord's hand was with him.
LUKE|1|67|His father Zechariah was filled with the Holy Spirit and prophesied:
LUKE|1|68|"Praise be to the Lord, the God of Israel, because he has come and has redeemed his people.
LUKE|1|69|He has raised up a horn of salvation for us in the house of his servant David
LUKE|1|70|(as he said through his holy prophets of long ago),
LUKE|1|71|salvation from our enemies and from the hand of all who hate us--
LUKE|1|72|to show mercy to our fathers and to remember his holy covenant,
LUKE|1|73|the oath he swore to our father Abraham:
LUKE|1|74|to rescue us from the hand of our enemies, and to enable us to serve him without fear
LUKE|1|75|in holiness and righteousness before him all our days.
LUKE|1|76|And you, my child, will be called a prophet of the Most High; for you will go on before the Lord to prepare the way for him,
LUKE|1|77|to give his people the knowledge of salvation through the forgiveness of their sins,
LUKE|1|78|because of the tender mercy of our God, by which the rising sun will come to us from heaven
LUKE|1|79|to shine on those living in darkness and in the shadow of death, to guide our feet into the path of peace."
LUKE|1|80|And the child grew and became strong in spirit; and he lived in the desert until he appeared publicly to Israel.
LUKE|2|1|In those days Caesar Augustus issued a decree that a census should be taken of the entire Roman world.
LUKE|2|2|(This was the first census that took place while Quirinius was governor of Syria.)
LUKE|2|3|And everyone went to his own town to register.
LUKE|2|4|So Joseph also went up from the town of Nazareth in Galilee to Judea, to Bethlehem the town of David, because he belonged to the house and line of David.
LUKE|2|5|He went there to register with Mary, who was pledged to be married to him and was expecting a child.
LUKE|2|6|While they were there, the time came for the baby to be born,
LUKE|2|7|and she gave birth to her firstborn, a son. She wrapped him in cloths and placed him in a manger, because there was no room for them in the inn.
LUKE|2|8|And there were shepherds living out in the fields nearby, keeping watch over their flocks at night.
LUKE|2|9|An angel of the Lord appeared to them, and the glory of the Lord shone around them, and they were terrified.
LUKE|2|10|But the angel said to them, "Do not be afraid. I bring you good news of great joy that will be for all the people.
LUKE|2|11|Today in the town of David a Savior has been born to you; he is Christ the Lord.
LUKE|2|12|This will be a sign to you: You will find a baby wrapped in cloths and lying in a manger."
LUKE|2|13|Suddenly a great company of the heavenly host appeared with the angel, praising God and saying,
LUKE|2|14|"Glory to God in the highest, and on earth peace to men on whom his favor rests."
LUKE|2|15|When the angels had left them and gone into heaven, the shepherds said to one another, "Let's go to Bethlehem and see this thing that has happened, which the Lord has told us about."
LUKE|2|16|So they hurried off and found Mary and Joseph, and the baby, who was lying in the manger.
LUKE|2|17|When they had seen him, they spread the word concerning what had been told them about this child,
LUKE|2|18|and all who heard it were amazed at what the shepherds said to them.
LUKE|2|19|But Mary treasured up all these things and pondered them in her heart.
LUKE|2|20|The shepherds returned, glorifying and praising God for all the things they had heard and seen, which were just as they had been told.
LUKE|2|21|On the eighth day, when it was time to circumcise him, he was named Jesus, the name the angel had given him before he had been conceived.
LUKE|2|22|When the time of their purification according to the Law of Moses had been completed, Joseph and Mary took him to Jerusalem to present him to the Lord
LUKE|2|23|(as it is written in the Law of the Lord, "Every firstborn male is to be consecrated to the Lord" ),
LUKE|2|24|and to offer a sacrifice in keeping with what is said in the Law of the Lord: "a pair of doves or two young pigeons."
LUKE|2|25|Now there was a man in Jerusalem called Simeon, who was righteous and devout. He was waiting for the consolation of Israel, and the Holy Spirit was upon him.
LUKE|2|26|It had been revealed to him by the Holy Spirit that he would not die before he had seen the Lord's Christ.
LUKE|2|27|Moved by the Spirit, he went into the temple courts. When the parents brought in the child Jesus to do for him what the custom of the Law required,
LUKE|2|28|Simeon took him in his arms and praised God, saying:
LUKE|2|29|"Sovereign Lord, as you have promised, you now dismiss your servant in peace.
LUKE|2|30|For my eyes have seen your salvation,
LUKE|2|31|which you have prepared in the sight of all people,
LUKE|2|32|a light for revelation to the Gentiles and for glory to your people Israel."
LUKE|2|33|The child's father and mother marveled at what was said about him.
LUKE|2|34|Then Simeon blessed them and said to Mary, his mother: "This child is destined to cause the falling and rising of many in Israel, and to be a sign that will be spoken against,
LUKE|2|35|so that the thoughts of many hearts will be revealed. And a sword will pierce your own soul too."
LUKE|2|36|There was also a prophetess, Anna, the daughter of Phanuel, of the tribe of Asher. She was very old; she had lived with her husband seven years after her marriage,
LUKE|2|37|and then was a widow until she was eighty-four. She never left the temple but worshiped night and day, fasting and praying.
LUKE|2|38|Coming up to them at that very moment, she gave thanks to God and spoke about the child to all who were looking forward to the redemption of Jerusalem.
LUKE|2|39|When Joseph and Mary had done everything required by the Law of the Lord, they returned to Galilee to their own town of Nazareth.
LUKE|2|40|And the child grew and became strong; he was filled with wisdom, and the grace of God was upon him.
LUKE|2|41|Every year his parents went to Jerusalem for the Feast of the Passover.
LUKE|2|42|When he was twelve years old, they went up to the Feast, according to the custom.
LUKE|2|43|After the Feast was over, while his parents were returning home, the boy Jesus stayed behind in Jerusalem, but they were unaware of it.
LUKE|2|44|Thinking he was in their company, they traveled on for a day. Then they began looking for him among their relatives and friends.
LUKE|2|45|When they did not find him, they went back to Jerusalem to look for him.
LUKE|2|46|After three days they found him in the temple courts, sitting among the teachers, listening to them and asking them questions.
LUKE|2|47|Everyone who heard him was amazed at his understanding and his answers.
LUKE|2|48|When his parents saw him, they were astonished. His mother said to him, "Son, why have you treated us like this? Your father and I have been anxiously searching for you."
LUKE|2|49|"Why were you searching for me?" he asked. "Didn't you know I had to be in my Father's house?"
LUKE|2|50|But they did not understand what he was saying to them.
LUKE|2|51|Then he went down to Nazareth with them and was obedient to them. But his mother treasured all these things in her heart.
LUKE|2|52|And Jesus grew in wisdom and stature, and in favor with God and men.
LUKE|3|1|In the fifteenth year of the reign of Tiberius Caesar--when Pontius Pilate was governor of Judea, Herod tetrarch of Galilee, his brother Philip tetrarch of Iturea and Traconitis, and Lysanias tetrarch of Abilene--
LUKE|3|2|during the high priesthood of Annas and Caiaphas, the word of God came to John son of Zechariah in the desert.
LUKE|3|3|He went into all the country around the Jordan, preaching a baptism of repentance for the forgiveness of sins.
LUKE|3|4|As is written in the book of the words of Isaiah the prophet: "A voice of one calling in the desert, 'Prepare the way for the Lord, make straight paths for him.
LUKE|3|5|Every valley shall be filled in, every mountain and hill made low. The crooked roads shall become straight, the rough ways smooth.
LUKE|3|6|And all mankind will see God's salvation.'"
LUKE|3|7|John said to the crowds coming out to be baptized by him, "You brood of vipers! Who warned you to flee from the coming wrath?
LUKE|3|8|Produce fruit in keeping with repentance. And do not begin to say to yourselves, 'We have Abraham as our father.' For I tell you that out of these stones God can raise up children for Abraham.
LUKE|3|9|The ax is already at the root of the trees, and every tree that does not produce good fruit will be cut down and thrown into the fire."
LUKE|3|10|"What should we do then?" the crowd asked.
LUKE|3|11|John answered, "The man with two tunics should share with him who has none, and the one who has food should do the same."
LUKE|3|12|Tax collectors also came to be baptized. "Teacher," they asked, "what should we do?"
LUKE|3|13|"Don't collect any more than you are required to," he told
LUKE|3|14|them. Then some soldiers asked him, "And what should we do?" He replied, "Don't extort money and don't accuse people falsely--be content with your pay."
LUKE|3|15|The people were waiting expectantly and were all wondering in their hearts if John might possibly be the Christ.
LUKE|3|16|John answered them all, "I baptize you with water. But one more powerful than I will come, the thongs of whose sandals I am not worthy to untie. He will baptize you with the Holy Spirit and with fire.
LUKE|3|17|His winnowing fork is in his hand to clear his threshing floor and to gather the wheat into his barn, but he will burn up the chaff with unquenchable fire."
LUKE|3|18|And with many other words John exhorted the people and preached the good news to them.
LUKE|3|19|But when John rebuked Herod the tetrarch because of Herodias, his brother's wife, and all the other evil things he had done,
LUKE|3|20|Herod added this to them all: He locked John up in prison.
LUKE|3|21|When all the people were being baptized, Jesus was baptized too. And as he was praying, heaven was opened
LUKE|3|22|and the Holy Spirit descended on him in bodily form like a dove. And a voice came from heaven: "You are my Son, whom I love; with you I am well pleased."
LUKE|3|23|Now Jesus himself was about thirty years old when he began his ministry. He was the son, so it was thought, of Joseph,
LUKE|3|24|the son of Heli, the son of Matthat, the son of Levi, the son of Melki, the son of Jannai, the son of Joseph,
LUKE|3|25|the son of Mattathias, the son of Amos, the son of Nahum, the son of Esli,
LUKE|3|26|the son of Naggai, the son of Maath, the son of Mattathias, the son of Semein, the son of Josech, the son of Joda,
LUKE|3|27|the son of Joanan, the son of Rhesa, the son of Zerubbabel, the son of Shealtiel,
LUKE|3|28|the son of Neri, the son of Melki, the son of Addi, the son of Cosam, the son of Elmadam, the son of Er,
LUKE|3|29|the son of Joshua, the son of Eliezer, the son of Jorim, the son of Matthat,
LUKE|3|30|the son of Levi, the son of Simeon, the son of Judah, the son of Joseph, the son of Jonam, the son of Eliakim,
LUKE|3|31|the son of Melea, the son of Menna, the son of Mattatha, the son of Nathan,
LUKE|3|32|the son of David, the son of Jesse, the son of Obed, the son of Boaz, the son of Salmon, the son of Nahshon,
LUKE|3|33|the son of Amminadab, the son of Ram, the son of Hezron, the son of Perez,
LUKE|3|34|the son of Judah, the son of Jacob, the son of Isaac, the son of Abraham, the son of Terah, the son of Nahor,
LUKE|3|35|the son of Serug, the son of Reu, the son of Peleg, the son of Eber,
LUKE|3|36|the son of Shelah, the son of Cainan, the son of Arphaxad, the son of Shem, the son of Noah, the son of Lamech,
LUKE|3|37|the son of Methuselah, the son of Enoch, the son of Jared, the son of Mahalalel,
LUKE|3|38|the son of Kenan, the son of Enosh, the son of Seth, the son of Adam, the son of God.
LUKE|4|1|Jesus, full of the Holy Spirit, returned from the Jordan and was led by the Spirit in the desert,
LUKE|4|2|where for forty days he was tempted by the devil. He ate nothing during those days, and at the end of them he was hungry.
LUKE|4|3|The devil said to him, "If you are the Son of God, tell this stone to become bread."
LUKE|4|4|Jesus answered, "It is written: 'Man does not live on bread alone.'"
LUKE|4|5|The devil led him up to a high place and showed him in an instant all the kingdoms of the world.
LUKE|4|6|And he said to him, "I will give you all their authority and splendor, for it has been given to me, and I can give it to anyone I want to.
LUKE|4|7|So if you worship me, it will all be yours."
LUKE|4|8|Jesus answered, "It is written: 'Worship the Lord your God and serve him only.'"
LUKE|4|9|The devil led him to Jerusalem and had him stand on the highest point of the temple. "If you are the Son of God," he said, "throw yourself down from here.
LUKE|4|10|For it is written: "'He will command his angels concerning you to guard you carefully;
LUKE|4|11|they will lift you up in their hands, so that you will not strike your foot against a stone.'"
LUKE|4|12|Jesus answered, "It says: 'Do not put the Lord your God to the test.'"
LUKE|4|13|When the devil had finished all this tempting, he left him until an opportune time.
LUKE|4|14|Jesus returned to Galilee in the power of the Spirit, and news about him spread through the whole countryside.
LUKE|4|15|He taught in their synagogues, and everyone praised him.
LUKE|4|16|He went to Nazareth, where he had been brought up, and on the Sabbath day he went into the synagogue, as was his custom. And he stood up to read.
LUKE|4|17|The scroll of the prophet Isaiah was handed to him. Unrolling it, he found the place where it is written:
LUKE|4|18|"The Spirit of the Lord is on me, because he has anointed me to preach good news to the poor. He has sent me to proclaim freedom for the prisoners and recovery of sight for the blind, to release the oppressed,
LUKE|4|19|to proclaim the year of the Lord's favor."
LUKE|4|20|Then he rolled up the scroll, gave it back to the attendant and sat down. The eyes of everyone in the synagogue were fastened on him,
LUKE|4|21|and he began by saying to them, "Today this scripture is fulfilled in your hearing."
LUKE|4|22|All spoke well of him and were amazed at the gracious words that came from his lips. "Isn't this Joseph's son?" they asked.
LUKE|4|23|Jesus said to them, "Surely you will quote this proverb to me: 'Physician, heal yourself! Do here in your hometown what we have heard that you did in Capernaum.'"
LUKE|4|24|"I tell you the truth," he continued, "no prophet is accepted in his hometown.
LUKE|4|25|I assure you that there were many widows in Israel in Elijah's time, when the sky was shut for three and a half years and there was a severe famine throughout the land.
LUKE|4|26|Yet Elijah was not sent to any of them, but to a widow in Zarephath in the region of Sidon.
LUKE|4|27|And there were many in Israel with leprosy in the time of Elisha the prophet, yet not one of them was cleansed--only Naaman the Syrian."
LUKE|4|28|All the people in the synagogue were furious when they heard this.
LUKE|4|29|They got up, drove him out of the town, and took him to the brow of the hill on which the town was built, in order to throw him down the cliff.
LUKE|4|30|But he walked right through the crowd and went on his way.
LUKE|4|31|Then he went down to Capernaum, a town in Galilee, and on the Sabbath began to teach the people.
LUKE|4|32|They were amazed at his teaching, because his message had authority.
LUKE|4|33|In the synagogue there was a man possessed by a demon, an evil spirit. He cried out at the top of his voice,
LUKE|4|34|"Ha! What do you want with us, Jesus of Nazareth? Have you come to destroy us? I know who you are--the Holy One of God!"
LUKE|4|35|"Be quiet!" Jesus said sternly. "Come out of him!" Then the demon threw the man down before them all and came out without injuring him.
LUKE|4|36|All the people were amazed and said to each other, "What is this teaching? With authority and power he gives orders to evil spirits and they come out!"
LUKE|4|37|And the news about him spread throughout the surrounding area.
LUKE|4|38|Jesus left the synagogue and went to the home of Simon. Now Simon's mother-in-law was suffering from a high fever, and they asked Jesus to help her.
LUKE|4|39|So he bent over her and rebuked the fever, and it left her. She got up at once and began to wait on them.
LUKE|4|40|When the sun was setting, the people brought to Jesus all who had various kinds of sickness, and laying his hands on each one, he healed them.
LUKE|4|41|Moreover, demons came out of many people, shouting, "You are the Son of God!" But he rebuked them and would not allow them to speak, because they knew he was the Christ.
LUKE|4|42|At daybreak Jesus went out to a solitary place. The people were looking for him and when they came to where he was, they tried to keep him from leaving them.
LUKE|4|43|But he said, "I must preach the good news of the kingdom of God to the other towns also, because that is why I was sent."
LUKE|4|44|And he kept on preaching in the synagogues of Judea.
LUKE|5|1|One day as Jesus was standing by the Lake of Gennesaret, with the people crowding around him and listening to the word of God,
LUKE|5|2|he saw at the water's edge two boats, left there by the fishermen, who were washing their nets.
LUKE|5|3|He got into one of the boats, the one belonging to Simon, and asked him to put out a little from shore. Then he sat down and taught the people from the boat.
LUKE|5|4|When he had finished speaking, he said to Simon, "Put out into deep water, and let down the nets for a catch."
LUKE|5|5|Simon answered, "Master, we've worked hard all night and haven't caught anything. But because you say so, I will let down the nets."
LUKE|5|6|When they had done so, they caught such a large number of fish that their nets began to break.
LUKE|5|7|So they signaled their partners in the other boat to come and help them, and they came and filled both boats so full that they began to sink.
LUKE|5|8|When Simon Peter saw this, he fell at Jesus' knees and said, "Go away from me, Lord; I am a sinful man!"
LUKE|5|9|For he and all his companions were astonished at the catch of fish they had taken,
LUKE|5|10|and so were James and John, the sons of Zebedee, Simon's partners.
LUKE|5|11|Then Jesus said to Simon, "Don't be afraid; from now on you will catch men." So they pulled their boats up on shore, left everything and followed him.
LUKE|5|12|While Jesus was in one of the towns, a man came along who was covered with leprosy. When he saw Jesus, he fell with his face to the ground and begged him, "Lord, if you are willing, you can make me clean."
LUKE|5|13|Jesus reached out his hand and touched the man. "I am willing," he said. "Be clean!" And immediately the leprosy left him.
LUKE|5|14|Then Jesus ordered him, "Don't tell anyone, but go, show yourself to the priest and offer the sacrifices that Moses commanded for your cleansing, as a testimony to them."
LUKE|5|15|Yet the news about him spread all the more, so that crowds of people came to hear him and to be healed of their sicknesses.
LUKE|5|16|But Jesus often withdrew to lonely places and prayed.
LUKE|5|17|One day as he was teaching, Pharisees and teachers of the law, who had come from every village of Galilee and from Judea and Jerusalem, were sitting there. And the power of the Lord was present for him to heal the sick.
LUKE|5|18|Some men came carrying a paralytic on a mat and tried to take him into the house to lay him before Jesus.
LUKE|5|19|When they could not find a way to do this because of the crowd, they went up on the roof and lowered him on his mat through the tiles into the middle of the crowd, right in front of Jesus.
LUKE|5|20|When Jesus saw their faith, he said, "Friend, your sins are forgiven."
LUKE|5|21|The Pharisees and the teachers of the law began thinking to themselves, "Who is this fellow who speaks blasphemy? Who can forgive sins but God alone?"
LUKE|5|22|Jesus knew what they were thinking and asked, "Why are you thinking these things in your hearts?
LUKE|5|23|Which is easier: to say, 'Your sins are forgiven,' or to say, 'Get up and walk'?
LUKE|5|24|But that you may know that the Son of Man has authority on earth to forgive sins...." He said to the paralyzed man, "I tell you, get up, take your mat and go home."
LUKE|5|25|Immediately he stood up in front of them, took what he had been lying on and went home praising God.
LUKE|5|26|Everyone was amazed and gave praise to God. They were filled with awe and said, "We have seen remarkable things today."
LUKE|5|27|After this, Jesus went out and saw a tax collector by the name of Levi sitting at his tax booth. "Follow me," Jesus said to him,
LUKE|5|28|and Levi got up, left everything and followed him.
LUKE|5|29|Then Levi held a great banquet for Jesus at his house, and a large crowd of tax collectors and others were eating with them.
LUKE|5|30|But the Pharisees and the teachers of the law who belonged to their sect complained to his disciples, "Why do you eat and drink with tax collectors and 'sinners'?"
LUKE|5|31|Jesus answered them, "It is not the healthy who need a doctor, but the sick.
LUKE|5|32|I have not come to call the righteous, but sinners to repentance."
LUKE|5|33|They said to him, "John's disciples often fast and pray, and so do the disciples of the Pharisees, but yours go on eating and drinking."
LUKE|5|34|Jesus answered, "Can you make the guests of the bridegroom fast while he is with them?
LUKE|5|35|But the time will come when the bridegroom will be taken from them; in those days they will fast."
LUKE|5|36|He told them this parable: "No one tears a patch from a new garment and sews it on an old one. If he does, he will have torn the new garment, and the patch from the new will not match the old.
LUKE|5|37|And no one pours new wine into old wineskins. If he does, the new wine will burst the skins, the wine will run out and the wineskins will be ruined.
LUKE|5|38|No, new wine must be poured into new wineskins.
LUKE|5|39|And no one after drinking old wine wants the new, for he says, 'The old is better.'"
LUKE|6|1|One Sabbath Jesus was going through the grainfields, and his disciples began to pick some heads of grain, rub them in their hands and eat the kernels.
LUKE|6|2|Some of the Pharisees asked, "Why are you doing what is unlawful on the Sabbath?"
LUKE|6|3|Jesus answered them, "Have you never read what David did when he and his companions were hungry?
LUKE|6|4|He entered the house of God, and taking the consecrated bread, he ate what is lawful only for priests to eat. And he also gave some to his companions."
LUKE|6|5|Then Jesus said to them, "The Son of Man is Lord of the Sabbath."
LUKE|6|6|On another Sabbath he went into the synagogue and was teaching, and a man was there whose right hand was shriveled.
LUKE|6|7|The Pharisees and the teachers of the law were looking for a reason to accuse Jesus, so they watched him closely to see if he would heal on the Sabbath.
LUKE|6|8|But Jesus knew what they were thinking and said to the man with the shriveled hand, "Get up and stand in front of everyone." So he got up and stood there.
LUKE|6|9|Then Jesus said to them, "I ask you, which is lawful on the Sabbath: to do good or to do evil, to save life or to destroy it?"
LUKE|6|10|He looked around at them all, and then said to the man, "Stretch out your hand." He did so, and his hand was completely restored.
LUKE|6|11|But they were furious and began to discuss with one another what they might do to Jesus.
LUKE|6|12|One of those days Jesus went out to a mountainside to pray, and spent the night praying to God.
LUKE|6|13|When morning came, he called his disciples to him and chose twelve of them, whom he also designated apostles:
LUKE|6|14|Simon (whom he named Peter), his brother Andrew, James, John, Philip, Bartholomew,
LUKE|6|15|Matthew, Thomas, James son of Alphaeus, Simon who was called the Zealot,
LUKE|6|16|Judas son of James, and Judas Iscariot, who became a traitor.
LUKE|6|17|He went down with them and stood on a level place. A large crowd of his disciples was there and a great number of people from all over Judea, from Jerusalem, and from the coast of Tyre and Sidon,
LUKE|6|18|who had come to hear him and to be healed of their diseases. Those troubled by evil spirits were cured,
LUKE|6|19|and the people all tried to touch him, because power was coming from him and healing them all.
LUKE|6|20|Looking at his disciples, he said: "Blessed are you who are poor, for yours is the kingdom of God.
LUKE|6|21|Blessed are you who hunger now, for you will be satisfied. Blessed are you who weep now, for you will laugh.
LUKE|6|22|Blessed are you when men hate you, when they exclude you and insult you and reject your name as evil, because of the Son of Man.
LUKE|6|23|"Rejoice in that day and leap for joy, because great is your reward in heaven. For that is how their fathers treated the prophets.
LUKE|6|24|"But woe to you who are rich, for you have already received your comfort.
LUKE|6|25|Woe to you who are well fed now, for you will go hungry. Woe to you who laugh now, for you will mourn and weep.
LUKE|6|26|Woe to you when all men speak well of you, for that is how their fathers treated the false prophets.
LUKE|6|27|"But I tell you who hear me: Love your enemies, do good to those who hate you,
LUKE|6|28|bless those who curse you, pray for those who mistreat you.
LUKE|6|29|If someone strikes you on one cheek, turn to him the other also. If someone takes your cloak, do not stop him from taking your tunic.
LUKE|6|30|Give to everyone who asks you, and if anyone takes what belongs to you, do not demand it back.
LUKE|6|31|Do to others as you would have them do to you.
LUKE|6|32|"If you love those who love you, what credit is that to you? Even 'sinners' love those who love them.
LUKE|6|33|And if you do good to those who are good to you, what credit is that to you? Even 'sinners' do that.
LUKE|6|34|And if you lend to those from whom you expect repayment, what credit is that to you? Even 'sinners' lend to 'sinners,' expecting to be repaid in full.
LUKE|6|35|But love your enemies, do good to them, and lend to them without expecting to get anything back. Then your reward will be great, and you will be sons of the Most High, because he is kind to the ungrateful and wicked.
LUKE|6|36|Be merciful, just as your Father is merciful.
LUKE|6|37|"Do not judge, and you will not be judged. Do not condemn, and you will not be condemned. Forgive, and you will be forgiven.
LUKE|6|38|Give, and it will be given to you. A good measure, pressed down, shaken together and running over, will be poured into your lap. For with the measure you use, it will be measured to you."
LUKE|6|39|He also told them this parable: "Can a blind man lead a blind man? Will they not both fall into a pit?
LUKE|6|40|A student is not above his teacher, but everyone who is fully trained will be like his teacher.
LUKE|6|41|"Why do you look at the speck of sawdust in your brother's eye and pay no attention to the plank in your own eye?
LUKE|6|42|How can you say to your brother, 'Brother, let me take the speck out of your eye,' when you yourself fail to see the plank in your own eye? You hypocrite, first take the plank out of your eye, and then you will see clearly to remove the speck from your brother's eye.
LUKE|6|43|"No good tree bears bad fruit, nor does a bad tree bear good fruit.
LUKE|6|44|Each tree is recognized by its own fruit. People do not pick figs from thornbushes, or grapes from briers.
LUKE|6|45|The good man brings good things out of the good stored up in his heart, and the evil man brings evil things out of the evil stored up in his heart. For out of the overflow of his heart his mouth speaks.
LUKE|6|46|"Why do you call me, 'Lord, Lord,' and do not do what I say?
LUKE|6|47|I will show you what he is like who comes to me and hears my words and puts them into practice.
LUKE|6|48|He is like a man building a house, who dug down deep and laid the foundation on rock. When a flood came, the torrent struck that house but could not shake it, because it was well built.
LUKE|6|49|But the one who hears my words and does not put them into practice is like a man who built a house on the ground without a foundation. The moment the torrent struck that house, it collapsed and its destruction was complete."
LUKE|7|1|When Jesus had finished saying all this in the hearing of the people, he entered Capernaum.
LUKE|7|2|There a centurion's servant, whom his master valued highly, was sick and about to die.
LUKE|7|3|The centurion heard of Jesus and sent some elders of the Jews to him, asking him to come and heal his servant.
LUKE|7|4|When they came to Jesus, they pleaded earnestly with him, "This man deserves to have you do this,
LUKE|7|5|because he loves our nation and has built our synagogue."
LUKE|7|6|So Jesus went with them. He was not far from the house when the centurion sent friends to say to him: "Lord, don't trouble yourself, for I do not deserve to have you come under my roof.
LUKE|7|7|That is why I did not even consider myself worthy to come to you. But say the word, and my servant will be healed.
LUKE|7|8|For I myself am a man under authority, with soldiers under me. I tell this one, 'Go,' and he goes; and that one, 'Come,' and he comes. I say to my servant, 'Do this,' and he does it."
LUKE|7|9|When Jesus heard this, he was amazed at him, and turning to the crowd following him, he said, "I tell you, I have not found such great faith even in Israel."
LUKE|7|10|Then the men who had been sent returned to the house and found the servant well.
LUKE|7|11|Soon afterward, Jesus went to a town called Nain, and his disciples and a large crowd went along with him.
LUKE|7|12|As he approached the town gate, a dead person was being carried out--the only son of his mother, and she was a widow. And a large crowd from the town was with her.
LUKE|7|13|When the Lord saw her, his heart went out to her and he said, "Don't cry."
LUKE|7|14|Then he went up and touched the coffin, and those carrying it stood still. He said, "Young man, I say to you, get up!"
LUKE|7|15|The dead man sat up and began to talk, and Jesus gave him back to his mother.
LUKE|7|16|They were all filled with awe and praised God. "A great prophet has appeared among us," they said. "God has come to help his people."
LUKE|7|17|This news about Jesus spread throughout Judea and the surrounding country.
LUKE|7|18|John's disciples told him about all these things. Calling two of them,
LUKE|7|19|he sent them to the Lord to ask, "Are you the one who was to come, or should we expect someone else?"
LUKE|7|20|When the men came to Jesus, they said, "John the Baptist sent us to you to ask, 'Are you the one who was to come, or should we expect someone else?'"
LUKE|7|21|At that very time Jesus cured many who had diseases, sicknesses and evil spirits, and gave sight to many who were blind.
LUKE|7|22|So he replied to the messengers, "Go back and report to John what you have seen and heard: The blind receive sight, the lame walk, those who have leprosy are cured, the deaf hear, the dead are raised, and the good news is preached to the poor.
LUKE|7|23|Blessed is the man who does not fall away on account of me."
LUKE|7|24|After John's messengers left, Jesus began to speak to the crowd about John: "What did you go out into the desert to see? A reed swayed by the wind?
LUKE|7|25|If not, what did you go out to see? A man dressed in fine clothes? No, those who wear expensive clothes and indulge in luxury are in palaces.
LUKE|7|26|But what did you go out to see? A prophet? Yes, I tell you, and more than a prophet.
LUKE|7|27|This is the one about whom it is written: "'I will send my messenger ahead of you, who will prepare your way before you.'
LUKE|7|28|I tell you, among those born of women there is no one greater than John; yet the one who is least in the kingdom of God is greater than he."
LUKE|7|29|(All the people, even the tax collectors, when they heard Jesus' words, acknowledged that God's way was right, because they had been baptized by John.
LUKE|7|30|But the Pharisees and experts in the law rejected God's purpose for themselves, because they had not been baptized by John.)
LUKE|7|31|"To what, then, can I compare the people of this generation? What are they like?
LUKE|7|32|They are like children sitting in the marketplace and calling out to each other: "'We played the flute for you, and you did not dance; we sang a dirge, and you did not cry.'
LUKE|7|33|For John the Baptist came neither eating bread nor drinking wine, and you say, 'He has a demon.'
LUKE|7|34|The Son of Man came eating and drinking, and you say, 'Here is a glutton and a drunkard, a friend of tax collectors and "sinners."'
LUKE|7|35|But wisdom is proved right by all her children."
LUKE|7|36|Now one of the Pharisees invited Jesus to have dinner with him, so he went to the Pharisee's house and reclined at the table.
LUKE|7|37|When a woman who had lived a sinful life in that town learned that Jesus was eating at the Pharisee's house, she brought an alabaster jar of perfume,
LUKE|7|38|and as she stood behind him at his feet weeping, she began to wet his feet with her tears. Then she wiped them with her hair, kissed them and poured perfume on them.
LUKE|7|39|When the Pharisee who had invited him saw this, he said to himself, "If this man were a prophet, he would know who is touching him and what kind of woman she is--that she is a sinner."
LUKE|7|40|Jesus answered him, "Simon, I have something to tell you.Tell me, teacher," he said.
LUKE|7|41|"Two men owed money to a certain moneylender. One owed him five hundred denarii, and the other fifty.
LUKE|7|42|Neither of them had the money to pay him back, so he canceled the debts of both. Now which of them will love him more?"
LUKE|7|43|Simon replied, "I suppose the one who had the bigger debt canceled.You have judged correctly," Jesus said.
LUKE|7|44|Then he turned toward the woman and said to Simon, "Do you see this woman? I came into your house. You did not give me any water for my feet, but she wet my feet with her tears and wiped them with her hair.
LUKE|7|45|You did not give me a kiss, but this woman, from the time I entered, has not stopped kissing my feet.
LUKE|7|46|You did not put oil on my head, but she has poured perfume on my feet.
LUKE|7|47|Therefore, I tell you, her many sins have been forgiven--for she loved much. But he who has been forgiven little loves little."
LUKE|7|48|Then Jesus said to her, "Your sins are forgiven."
LUKE|7|49|The other guests began to say among themselves, "Who is this who even forgives sins?"
LUKE|7|50|Jesus said to the woman, "Your faith has saved you; go in peace."
LUKE|8|1|After this, Jesus traveled about from one town and village to another, proclaiming the good news of the kingdom of God. The Twelve were with him,
LUKE|8|2|and also some women who had been cured of evil spirits and diseases: Mary (called Magdalene) from whom seven demons had come out;
LUKE|8|3|Joanna the wife of Cuza, the manager of Herod's household; Susanna; and many others. These women were helping to support them out of their own means.
LUKE|8|4|While a large crowd was gathering and people were coming to Jesus from town after town, he told this parable:
LUKE|8|5|"A farmer went out to sow his seed. As he was scattering the seed, some fell along the path; it was trampled on, and the birds of the air ate it up.
LUKE|8|6|Some fell on rock, and when it came up, the plants withered because they had no moisture.
LUKE|8|7|Other seed fell among thorns, which grew up with it and choked the plants.
LUKE|8|8|Still other seed fell on good soil. It came up and yielded a crop, a hundred times more than was sown." When he said this, he called out, "He who has ears to hear, let him hear."
LUKE|8|9|His disciples asked him what this parable meant.
LUKE|8|10|He said, "The knowledge of the secrets of the kingdom of God has been given to you, but to others I speak in parables, so that, "'though seeing, they may not see; though hearing, they may not understand.'
LUKE|8|11|"This is the meaning of the parable: The seed is the word of God.
LUKE|8|12|Those along the path are the ones who hear, and then the devil comes and takes away the word from their hearts, so that they may not believe and be saved.
LUKE|8|13|Those on the rock are the ones who receive the word with joy when they hear it, but they have no root. They believe for a while, but in the time of testing they fall away.
LUKE|8|14|The seed that fell among thorns stands for those who hear, but as they go on their way they are choked by life's worries, riches and pleasures, and they do not mature.
LUKE|8|15|But the seed on good soil stands for those with a noble and good heart, who hear the word, retain it, and by persevering produce a crop.
LUKE|8|16|"No one lights a lamp and hides it in a jar or puts it under a bed. Instead, he puts it on a stand, so that those who come in can see the light.
LUKE|8|17|For there is nothing hidden that will not be disclosed, and nothing concealed that will not be known or brought out into the open.
LUKE|8|18|Therefore consider carefully how you listen. Whoever has will be given more; whoever does not have, even what he thinks he has will be taken from him."
LUKE|8|19|Now Jesus' mother and brothers came to see him, but they were not able to get near him because of the crowd.
LUKE|8|20|Someone told him, "Your mother and brothers are standing outside, wanting to see you."
LUKE|8|21|He replied, "My mother and brothers are those who hear God's word and put it into practice."
LUKE|8|22|One day Jesus said to his disciples, "Let's go over to the other side of the lake." So they got into a boat and set out.
LUKE|8|23|As they sailed, he fell asleep. A squall came down on the lake, so that the boat was being swamped, and they were in great danger.
LUKE|8|24|The disciples went and woke him, saying, "Master, Master, we're going to drown!"
LUKE|8|25|He got up and rebuked the wind and the raging waters; the storm subsided, and all was calm. "Where is your faith?" he asked his disciples. In fear and amazement they asked one another, "Who is this? He commands even the winds and the water, and they obey him."
LUKE|8|26|They sailed to the region of the Gerasenes, which is across the lake from Galilee.
LUKE|8|27|When Jesus stepped ashore, he was met by a demon-possessed man from the town. For a long time this man had not worn clothes or lived in a house, but had lived in the tombs.
LUKE|8|28|When he saw Jesus, he cried out and fell at his feet, shouting at the top of his voice, "What do you want with me, Jesus, Son of the Most High God? I beg you, don't torture me!"
LUKE|8|29|For Jesus had commanded the evil spirit to come out of the man. Many times it had seized him, and though he was chained hand and foot and kept under guard, he had broken his chains and had been driven by the demon into solitary places.
LUKE|8|30|Jesus asked him, "What is your name?"
LUKE|8|31|"Legion," he replied, because many demons had gone into him. And they begged him repeatedly not to order them to go into the Abyss.
LUKE|8|32|A large herd of pigs was feeding there on the hillside. The demons begged Jesus to let them go into them, and he gave them permission.
LUKE|8|33|When the demons came out of the man, they went into the pigs, and the herd rushed down the steep bank into the lake and was drowned.
LUKE|8|34|When those tending the pigs saw what had happened, they ran off and reported this in the town and countryside,
LUKE|8|35|and the people went out to see what had happened. When they came to Jesus, they found the man from whom the demons had gone out, sitting at Jesus' feet, dressed and in his right mind; and they were afraid.
LUKE|8|36|Those who had seen it told the people how the demon-possessed man had been cured.
LUKE|8|37|Then all the people of the region of the Gerasenes asked Jesus to leave them, because they were overcome with fear. So he got into the boat and left.
LUKE|8|38|The man from whom the demons had gone out begged to go with him, but Jesus sent him away, saying,
LUKE|8|39|"Return home and tell how much God has done for you." So the man went away and told all over town how much Jesus had done for him.
LUKE|8|40|Now when Jesus returned, a crowd welcomed him, for they were all expecting him.
LUKE|8|41|Then a man named Jairus, a ruler of the synagogue, came and fell at Jesus' feet, pleading with him to come to his house
LUKE|8|42|because his only daughter, a girl of about twelve, was dying.
LUKE|8|43|As Jesus was on his way, the crowds almost crushed him. And a woman was there who had been subject to bleeding for twelve years, but no one could heal her.
LUKE|8|44|She came up behind him and touched the edge of his cloak, and immediately her bleeding stopped.
LUKE|8|45|"Who touched me?" Jesus asked. When they all denied it, Peter said, "Master, the people are crowding and pressing against you."
LUKE|8|46|But Jesus said, "Someone touched me; I know that power has gone out from me."
LUKE|8|47|Then the woman, seeing that she could not go unnoticed, came trembling and fell at his feet. In the presence of all the people, she told why she had touched him and how she had been instantly healed.
LUKE|8|48|Then he said to her, "Daughter, your faith has healed you. Go in peace."
LUKE|8|49|While Jesus was still speaking, someone came from the house of Jairus, the synagogue ruler. "Your daughter is dead," he said. "Don't bother the teacher any more."
LUKE|8|50|Hearing this, Jesus said to Jairus, "Don't be afraid; just believe, and she will be healed."
LUKE|8|51|When he arrived at the house of Jairus, he did not let anyone go in with him except Peter, John and James, and the child's father and mother.
LUKE|8|52|Meanwhile, all the people were wailing and mourning for her. "Stop wailing," Jesus said. "She is not dead but asleep."
LUKE|8|53|They laughed at him, knowing that she was dead.
LUKE|8|54|But he took her by the hand and said, "My child, get up!"
LUKE|8|55|Her spirit returned, and at once she stood up. Then Jesus told them to give her something to eat.
LUKE|8|56|Her parents were astonished, but he ordered them not to tell anyone what had happened.
LUKE|9|1|When Jesus had called the Twelve together, he gave them power and authority to drive out all demons and to cure diseases,
LUKE|9|2|and he sent them out to preach the kingdom of God and to heal the sick.
LUKE|9|3|He told them: "Take nothing for the journey--no staff, no bag, no bread, no money, no extra tunic.
LUKE|9|4|Whatever house you enter, stay there until you leave that town.
LUKE|9|5|If people do not welcome you, shake the dust off your feet when you leave their town, as a testimony against them."
LUKE|9|6|So they set out and went from village to village, preaching the gospel and healing people everywhere.
LUKE|9|7|Now Herod the tetrarch heard about all that was going on. And he was perplexed, because some were saying that John had been raised from the dead,
LUKE|9|8|others that Elijah had appeared, and still others that one of the prophets of long ago had come back to life.
LUKE|9|9|But Herod said, "I beheaded John. Who, then, is this I hear such things about?" And he tried to see him.
LUKE|9|10|When the apostles returned, they reported to Jesus what they had done. Then he took them with him and they withdrew by themselves to a town called Bethsaida,
LUKE|9|11|but the crowds learned about it and followed him. He welcomed them and spoke to them about the kingdom of God, and healed those who needed healing.
LUKE|9|12|Late in the afternoon the Twelve came to him and said, "Send the crowd away so they can go to the surrounding villages and countryside and find food and lodging, because we are in a remote place here."
LUKE|9|13|He replied, "You give them something to eat."
LUKE|9|14|They answered, "We have only five loaves of bread and two fish--unless we go and buy food for all this crowd." (About five thousand men were there.)
LUKE|9|15|But he said to his disciples, "Have them sit down in groups of about fifty each." The disciples did so, and everybody sat down.
LUKE|9|16|Taking the five loaves and the two fish and looking up to heaven, he gave thanks and broke them. Then he gave them to the disciples to set before the people.
LUKE|9|17|They all ate and were satisfied, and the disciples picked up twelve basketfuls of broken pieces that were left over.
LUKE|9|18|Once when Jesus was praying in private and his disciples were with him, he asked them, "Who do the crowds say I am?"
LUKE|9|19|They replied, "Some say John the Baptist; others say Elijah; and still others, that one of the prophets of long ago has come back to life."
LUKE|9|20|"But what about you?" he asked. "Who do you say I am?" Peter answered, "The Christ of God."
LUKE|9|21|Jesus strictly warned them not to tell this to anyone.
LUKE|9|22|And he said, "The Son of Man must suffer many things and be rejected by the elders, chief priests and teachers of the law, and he must be killed and on the third day be raised to life."
LUKE|9|23|Then he said to them all: "If anyone would come after me, he must deny himself and take up his cross daily and follow me.
LUKE|9|24|For whoever wants to save his life will lose it, but whoever loses his life for me will save it.
LUKE|9|25|What good is it for a man to gain the whole world, and yet lose or forfeit his very self?
LUKE|9|26|If anyone is ashamed of me and my words, the Son of Man will be ashamed of him when he comes in his glory and in the glory of the Father and of the holy angels.
LUKE|9|27|I tell you the truth, some who are standing here will not taste death before they see the kingdom of God."
LUKE|9|28|About eight days after Jesus said this, he took Peter, John and James with him and went up onto a mountain to pray.
LUKE|9|29|As he was praying, the appearance of his face changed, and his clothes became as bright as a flash of lightning.
LUKE|9|30|Two men, Moses and Elijah,
LUKE|9|31|appeared in glorious splendor, talking with Jesus. They spoke about his departure, which he was about to bring to fulfillment at Jerusalem.
LUKE|9|32|Peter and his companions were very sleepy, but when they became fully awake, they saw his glory and the two men standing with him.
LUKE|9|33|As the men were leaving Jesus, Peter said to him, "Master, it is good for us to be here. Let us put up three shelters--one for you, one for Moses and one for Elijah." (He did not know what he was saying.)
LUKE|9|34|While he was speaking, a cloud appeared and enveloped them, and they were afraid as they entered the cloud.
LUKE|9|35|A voice came from the cloud, saying, "This is my Son, whom I have chosen; listen to him."
LUKE|9|36|When the voice had spoken, they found that Jesus was alone. The disciples kept this to themselves, and told no one at that time what they had seen.
LUKE|9|37|The next day, when they came down from the mountain, a large crowd met him.
LUKE|9|38|A man in the crowd called out, "Teacher, I beg you to look at my son, for he is my only child.
LUKE|9|39|A spirit seizes him and he suddenly screams; it throws him into convulsions so that he foams at the mouth. It scarcely ever leaves him and is destroying him.
LUKE|9|40|I begged your disciples to drive it out, but they could not."
LUKE|9|41|"O unbelieving and perverse generation," Jesus replied, "how long shall I stay with you and put up with you? Bring your son here."
LUKE|9|42|Even while the boy was coming, the demon threw him to the ground in a convulsion. But Jesus rebuked the evil spirit, healed the boy and gave him back to his father.
LUKE|9|43|And they were all amazed at the greatness of God.
LUKE|9|44|While everyone was marveling at all that Jesus did, he said to his disciples, "Listen carefully to what I am about to tell you: The Son of Man is going to be betrayed into the hands of men."
LUKE|9|45|But they did not understand what this meant. It was hidden from them, so that they did not grasp it, and they were afraid to ask him about it.
LUKE|9|46|An argument started among the disciples as to which of them would be the greatest.
LUKE|9|47|Jesus, knowing their thoughts, took a little child and had him stand beside him.
LUKE|9|48|Then he said to them, "Whoever welcomes this little child in my name welcomes me; and whoever welcomes me welcomes the one who sent me. For he who is least among you all--he is the greatest."
LUKE|9|49|"Master," said John, "we saw a man driving out demons in your name and we tried to stop him, because he is not one of us."
LUKE|9|50|"Do not stop him," Jesus said, "for whoever is not against you is for you."
LUKE|9|51|As the time approached for him to be taken up to heaven, Jesus resolutely set out for Jerusalem.
LUKE|9|52|And he sent messengers on ahead, who went into a Samaritan village to get things ready for him;
LUKE|9|53|but the people there did not welcome him, because he was heading for Jerusalem.
LUKE|9|54|When the disciples James and John saw this, they asked, "Lord, do you want us to call fire down from heaven to destroy them?"
LUKE|9|55|But Jesus turned and rebuked them,
LUKE|9|56|and they went to another village.
LUKE|9|57|As they were walking along the road, a man said to him, "I will follow you wherever you go."
LUKE|9|58|Jesus replied, "Foxes have holes and birds of the air have nests, but the Son of Man has no place to lay his head."
LUKE|9|59|He said to another man, "Follow me." But the man replied, "Lord, first let me go and bury my father."
LUKE|9|60|Jesus said to him, "Let the dead bury their own dead, but you go and proclaim the kingdom of God."
LUKE|9|61|Still another said, "I will follow you, Lord; but first let me go back and say good bye to my family."
LUKE|9|62|Jesus replied, "No one who puts his hand to the plow and looks back is fit for service in the kingdom of God."
LUKE|10|1|After this the Lord appointed seventy-two others and sent them two by two ahead of him to every town and place where he was about to go.
LUKE|10|2|He told them, "The harvest is plentiful, but the workers are few. Ask the Lord of the harvest, therefore, to send out workers into his harvest field.
LUKE|10|3|Go! I am sending you out like lambs among wolves.
LUKE|10|4|Do not take a purse or bag or sandals; and do not greet anyone on the road.
LUKE|10|5|"When you enter a house, first say, 'Peace to this house.'
LUKE|10|6|If a man of peace is there, your peace will rest on him; if not, it will return to you.
LUKE|10|7|Stay in that house, eating and drinking whatever they give you, for the worker deserves his wages. Do not move around from house to house.
LUKE|10|8|"When you enter a town and are welcomed, eat what is set before you.
LUKE|10|9|Heal the sick who are there and tell them, 'The kingdom of God is near you.'
LUKE|10|10|But when you enter a town and are not welcomed, go into its streets and say,
LUKE|10|11|'Even the dust of your town that sticks to our feet we wipe off against you. Yet be sure of this: The kingdom of God is near.'
LUKE|10|12|I tell you, it will be more bearable on that day for Sodom than for that town.
LUKE|10|13|"Woe to you, Korazin! Woe to you, Bethsaida! For if the miracles that were performed in you had been performed in Tyre and Sidon, they would have repented long ago, sitting in sackcloth and ashes.
LUKE|10|14|But it will be more bearable for Tyre and Sidon at the judgment than for you.
LUKE|10|15|And you, Capernaum, will you be lifted up to the skies? No, you will go down to the depths.
LUKE|10|16|"He who listens to you listens to me; he who rejects you rejects me; but he who rejects me rejects him who sent me."
LUKE|10|17|The seventy-two returned with joy and said, "Lord, even the demons submit to us in your name."
LUKE|10|18|He replied, "I saw Satan fall like lightning from heaven.
LUKE|10|19|I have given you authority to trample on snakes and scorpions and to overcome all the power of the enemy; nothing will harm you.
LUKE|10|20|However, do not rejoice that the spirits submit to you, but rejoice that your names are written in heaven."
LUKE|10|21|At that time Jesus, full of joy through the Holy Spirit, said, "I praise you, Father, Lord of heaven and earth, because you have hidden these things from the wise and learned, and revealed them to little children. Yes, Father, for this was your good pleasure.
LUKE|10|22|"All things have been committed to me by my Father. No one knows who the Son is except the Father, and no one knows who the Father is except the Son and those to whom the Son chooses to reveal him."
LUKE|10|23|Then he turned to his disciples and said privately, "Blessed are the eyes that see what you see.
LUKE|10|24|For I tell you that many prophets and kings wanted to see what you see but did not see it, and to hear what you hear but did not hear it."
LUKE|10|25|On one occasion an expert in the law stood up to test Jesus. "Teacher," he asked, "what must I do to inherit eternal life?"
LUKE|10|26|"What is written in the Law?" he replied. "How do you read it?"
LUKE|10|27|He answered: "'Love the Lord your God with all your heart and with all your soul and with all your strength and with all your mind'; and, 'Love your neighbor as yourself.'"
LUKE|10|28|"You have answered correctly," Jesus replied. "Do this and you will live."
LUKE|10|29|But he wanted to justify himself, so he asked Jesus, "And who is my neighbor?"
LUKE|10|30|In reply Jesus said: "A man was going down from Jerusalem to Jericho, when he fell into the hands of robbers. They stripped him of his clothes, beat him and went away, leaving him half dead.
LUKE|10|31|A priest happened to be going down the same road, and when he saw the man, he passed by on the other side.
LUKE|10|32|So too, a Levite, when he came to the place and saw him, passed by on the other side.
LUKE|10|33|But a Samaritan, as he traveled, came where the man was; and when he saw him, he took pity on him.
LUKE|10|34|He went to him and bandaged his wounds, pouring on oil and wine. Then he put the man on his own donkey, took him to an inn and took care of him.
LUKE|10|35|The next day he took out two silver coins and gave them to the innkeeper. 'Look after him,' he said, 'and when I return, I will reimburse you for any extra expense you may have.'
LUKE|10|36|"Which of these three do you think was a neighbor to the man who fell into the hands of robbers?"
LUKE|10|37|The expert in the law replied, "The one who had mercy on him." Jesus told him, "Go and do likewise."
LUKE|10|38|As Jesus and his disciples were on their way, he came to a village where a woman named Martha opened her home to him.
LUKE|10|39|She had a sister called Mary, who sat at the Lord's feet listening to what he said.
LUKE|10|40|But Martha was distracted by all the preparations that had to be made. She came to him and asked, "Lord, don't you care that my sister has left me to do the work by myself? Tell her to help me!"
LUKE|10|41|"Martha, Martha," the Lord answered, "you are worried and upset about many things,
LUKE|10|42|but only one thing is needed. Mary has chosen what is better, and it will not be taken away from her."
LUKE|11|1|One day Jesus was praying in a certain place. When he finished, one of his disciples said to him, "Lord, teach us to pray, just as John taught his disciples."
LUKE|11|2|He said to them, "When you pray, say: "'Father, hallowed be your name, your kingdom come.
LUKE|11|3|Give us each day our daily bread.
LUKE|11|4|Forgive us our sins, for we also forgive everyone who sins against us. And lead us not into temptation. '"
LUKE|11|5|Then he said to them, "Suppose one of you has a friend, and he goes to him at midnight and says, 'Friend, lend me three loaves of bread,
LUKE|11|6|because a friend of mine on a journey has come to me, and I have nothing to set before him.'
LUKE|11|7|"Then the one inside answers, 'Don't bother me. The door is already locked, and my children are with me in bed. I can't get up and give you anything.'
LUKE|11|8|I tell you, though he will not get up and give him the bread because he is his friend, yet because of the man's boldness he will get up and give him as much as he needs.
LUKE|11|9|"So I say to you: Ask and it will be given to you; seek and you will find; knock and the door will be opened to you.
LUKE|11|10|For everyone who asks receives; he who seeks finds; and to him who knocks, the door will be opened.
LUKE|11|11|"Which of you fathers, if your son asks for a fish, will give him a snake instead?
LUKE|11|12|Or if he asks for an egg, will give him a scorpion?
LUKE|11|13|If you then, though you are evil, know how to give good gifts to your children, how much more will your Father in heaven give the Holy Spirit to those who ask him!"
LUKE|11|14|Jesus was driving out a demon that was mute. When the demon left, the man who had been mute spoke, and the crowd was amazed.
LUKE|11|15|But some of them said, "By Beelzebub, the prince of demons, he is driving out demons."
LUKE|11|16|Others tested him by asking for a sign from heaven.
LUKE|11|17|Jesus knew their thoughts and said to them: "Any kingdom divided against itself will be ruined, and a house divided against itself will fall.
LUKE|11|18|If Satan is divided against himself, how can his kingdom stand? I say this because you claim that I drive out demons by Beelzebub.
LUKE|11|19|Now if I drive out demons by Beelzebub, by whom do your followers drive them out? So then, they will be your judges.
LUKE|11|20|But if I drive out demons by the finger of God, then the kingdom of God has come to you.
LUKE|11|21|"When a strong man, fully armed, guards his own house, his possessions are safe.
LUKE|11|22|But when someone stronger attacks and overpowers him, he takes away the armor in which the man trusted and divides up the spoils.
LUKE|11|23|"He who is not with me is against me, and he who does not gather with me, scatters.
LUKE|11|24|"When an evil spirit comes out of a man, it goes through arid places seeking rest and does not find it. Then it says, 'I will return to the house I left.'
LUKE|11|25|When it arrives, it finds the house swept clean and put in order.
LUKE|11|26|Then it goes and takes seven other spirits more wicked than itself, and they go in and live there. And the final condition of that man is worse than the first."
LUKE|11|27|As Jesus was saying these things, a woman in the crowd called out, "Blessed is the mother who gave you birth and nursed you."
LUKE|11|28|He replied, "Blessed rather are those who hear the word of God and obey it."
LUKE|11|29|As the crowds increased, Jesus said, "This is a wicked generation. It asks for a miraculous sign, but none will be given it except the sign of Jonah.
LUKE|11|30|For as Jonah was a sign to the Ninevites, so also will the Son of Man be to this generation.
LUKE|11|31|The Queen of the South will rise at the judgment with the men of this generation and condemn them; for she came from the ends of the earth to listen to Solomon's wisdom, and now one greater than Solomon is here.
LUKE|11|32|The men of Nineveh will stand up at the judgment with this generation and condemn it; for they repented at the preaching of Jonah, and now one greater than Jonah is here.
LUKE|11|33|"No one lights a lamp and puts it in a place where it will be hidden, or under a bowl. Instead he puts it on its stand, so that those who come in may see the light.
LUKE|11|34|Your eye is the lamp of your body. When your eyes are good, your whole body also is full of light. But when they are bad, your body also is full of darkness.
LUKE|11|35|See to it, then, that the light within you is not darkness.
LUKE|11|36|Therefore, if your whole body is full of light, and no part of it dark, it will be completely lighted, as when the light of a lamp shines on you."
LUKE|11|37|When Jesus had finished speaking, a Pharisee invited him to eat with him; so he went in and reclined at the table.
LUKE|11|38|But the Pharisee, noticing that Jesus did not first wash before the meal, was surprised.
LUKE|11|39|Then the Lord said to him, "Now then, you Pharisees clean the outside of the cup and dish, but inside you are full of greed and wickedness.
LUKE|11|40|You foolish people! Did not the one who made the outside make the inside also?
LUKE|11|41|But give what is inside the dish to the poor, and everything will be clean for you.
LUKE|11|42|"Woe to you Pharisees, because you give God a tenth of your mint, rue and all other kinds of garden herbs, but you neglect justice and the love of God. You should have practiced the latter without leaving the former undone.
LUKE|11|43|"Woe to you Pharisees, because you love the most important seats in the synagogues and greetings in the marketplaces.
LUKE|11|44|"Woe to you, because you are like unmarked graves, which men walk over without knowing it."
LUKE|11|45|One of the experts in the law answered him, "Teacher, when you say these things, you insult us also."
LUKE|11|46|Jesus replied, "And you experts in the law, woe to you, because you load people down with burdens they can hardly carry, and you yourselves will not lift one finger to help them.
LUKE|11|47|"Woe to you, because you build tombs for the prophets, and it was your forefathers who killed them.
LUKE|11|48|So you testify that you approve of what your forefathers did; they killed the prophets, and you build their tombs.
LUKE|11|49|Because of this, God in his wisdom said, 'I will send them prophets and apostles, some of whom they will kill and others they will persecute.'
LUKE|11|50|Therefore this generation will be held responsible for the blood of all the prophets that has been shed since the beginning of the world,
LUKE|11|51|from the blood of Abel to the blood of Zechariah, who was killed between the altar and the sanctuary. Yes, I tell you, this generation will be held responsible for it all.
LUKE|11|52|"Woe to you experts in the law, because you have taken away the key to knowledge. You yourselves have not entered, and you have hindered those who were entering."
LUKE|11|53|When Jesus left there, the Pharisees and the teachers of the law began to oppose him fiercely and to besiege him with questions,
LUKE|11|54|waiting to catch him in something he might say.
LUKE|12|1|Meanwhile, when a crowd of many thousands had gathered, so that they were trampling on one another, Jesus began to speak first to his disciples, saying: "Be on your guard against the yeast of the Pharisees, which is hypocrisy.
LUKE|12|2|There is nothing concealed that will not be disclosed, or hidden that will not be made known.
LUKE|12|3|What you have said in the dark will be heard in the daylight, and what you have whispered in the ear in the inner rooms will be proclaimed from the roofs.
LUKE|12|4|"I tell you, my friends, do not be afraid of those who kill the body and after that can do no more.
LUKE|12|5|But I will show you whom you should fear: Fear him who, after the killing of the body, has power to throw you into hell. Yes, I tell you, fear him.
LUKE|12|6|Are not five sparrows sold for two pennies? Yet not one of them is forgotten by God.
LUKE|12|7|Indeed, the very hairs of your head are all numbered. Don't be afraid; you are worth more than many sparrows.
LUKE|12|8|"I tell you, whoever acknowledges me before men, the Son of Man will also acknowledge him before the angels of God.
LUKE|12|9|But he who disowns me before men will be disowned before the angels of God.
LUKE|12|10|And everyone who speaks a word against the Son of Man will be forgiven, but anyone who blasphemes against the Holy Spirit will not be forgiven.
LUKE|12|11|"When you are brought before synagogues, rulers and authorities, do not worry about how you will defend yourselves or what you will say,
LUKE|12|12|for the Holy Spirit will teach you at that time what you should say."
LUKE|12|13|Someone in the crowd said to him, "Teacher, tell my brother to divide the inheritance with me."
LUKE|12|14|Jesus replied, "Man, who appointed me a judge or an arbiter between you?"
LUKE|12|15|Then he said to them, "Watch out! Be on your guard against all kinds of greed; a man's life does not consist in the abundance of his possessions."
LUKE|12|16|And he told them this parable: "The ground of a certain rich man produced a good crop.
LUKE|12|17|He thought to himself, 'What shall I do? I have no place to store my crops.'
LUKE|12|18|"Then he said, 'This is what I'll do. I will tear down my barns and build bigger ones, and there I will store all my grain and my goods.
LUKE|12|19|And I'll say to myself, "You have plenty of good things laid up for many years. Take life easy; eat, drink and be merry."'
LUKE|12|20|"But God said to him, 'You fool! This very night your life will be demanded from you. Then who will get what you have prepared for yourself?'
LUKE|12|21|"This is how it will be with anyone who stores up things for himself but is not rich toward God."
LUKE|12|22|Then Jesus said to his disciples: "Therefore I tell you, do not worry about your life, what you will eat; or about your body, what you will wear.
LUKE|12|23|Life is more than food, and the body more than clothes.
LUKE|12|24|Consider the ravens: They do not sow or reap, they have no storeroom or barn; yet God feeds them. And how much more valuable you are than birds!
LUKE|12|25|Who of you by worrying can add a single hour to his life?
LUKE|12|26|Since you cannot do this very little thing, why do you worry about the rest?
LUKE|12|27|"Consider how the lilies grow. They do not labor or spin. Yet I tell you, not even Solomon in all his splendor was dressed like one of these.
LUKE|12|28|If that is how God clothes the grass of the field, which is here today, and tomorrow is thrown into the fire, how much more will he clothe you, O you of little faith!
LUKE|12|29|And do not set your heart on what you will eat or drink; do not worry about it.
LUKE|12|30|For the pagan world runs after all such things, and your Father knows that you need them.
LUKE|12|31|But seek his kingdom, and these things will be given to you as well.
LUKE|12|32|"Do not be afraid, little flock, for your Father has been pleased to give you the kingdom.
LUKE|12|33|Sell your possessions and give to the poor. Provide purses for yourselves that will not wear out, a treasure in heaven that will not be exhausted, where no thief comes near and no moth destroys.
LUKE|12|34|For where your treasure is, there your heart will be also.
LUKE|12|35|"Be dressed ready for service and keep your lamps burning,
LUKE|12|36|like men waiting for their master to return from a wedding banquet, so that when he comes and knocks they can immediately open the door for him.
LUKE|12|37|It will be good for those servants whose master finds them watching when he comes. I tell you the truth, he will dress himself to serve, will have them recline at the table and will come and wait on them.
LUKE|12|38|It will be good for those servants whose master finds them ready, even if he comes in the second or third watch of the night.
LUKE|12|39|But understand this: If the owner of the house had known at what hour the thief was coming, he would not have let his house be broken into.
LUKE|12|40|You also must be ready, because the Son of Man will come at an hour when you do not expect him."
LUKE|12|41|Peter asked, "Lord, are you telling this parable to us, or to everyone?"
LUKE|12|42|The Lord answered, "Who then is the faithful and wise manager, whom the master puts in charge of his servants to give them their food allowance at the proper time?
LUKE|12|43|It will be good for that servant whom the master finds doing so when he returns.
LUKE|12|44|I tell you the truth, he will put him in charge of all his possessions.
LUKE|12|45|But suppose the servant says to himself, 'My master is taking a long time in coming,' and he then begins to beat the menservants and maidservants and to eat and drink and get drunk.
LUKE|12|46|The master of that servant will come on a day when he does not expect him and at an hour he is not aware of. He will cut him to pieces and assign him a place with the unbelievers.
LUKE|12|47|"That servant who knows his master's will and does not get ready or does not do what his master wants will be beaten with many blows.
LUKE|12|48|But the one who does not know and does things deserving punishment will be beaten with few blows. From everyone who has been given much, much will be demanded; and from the one who has been entrusted with much, much more will be asked.
LUKE|12|49|"I have come to bring fire on the earth, and how I wish it were already kindled!
LUKE|12|50|But I have a baptism to undergo, and how distressed I am until it is completed!
LUKE|12|51|Do you think I came to bring peace on earth? No, I tell you, but division.
LUKE|12|52|From now on there will be five in one family divided against each other, three against two and two against three.
LUKE|12|53|They will be divided, father against son and son against father, mother against daughter and daughter against mother, mother-in-law against daughter-in-law and daughter-in-law against mother-in-law."
LUKE|12|54|He said to the crowd: "When you see a cloud rising in the west, immediately you say, 'It's going to rain,' and it does.
LUKE|12|55|And when the south wind blows, you say, 'It's going to be hot,' and it is.
LUKE|12|56|Hypocrites! You know how to interpret the appearance of the earth and the sky. How is it that you don't know how to interpret this present time?
LUKE|12|57|"Why don't you judge for yourselves what is right?
LUKE|12|58|As you are going with your adversary to the magistrate, try hard to be reconciled to him on the way, or he may drag you off to the judge, and the judge turn you over to the officer, and the officer throw you into prison.
LUKE|12|59|I tell you, you will not get out until you have paid the last penny. "
LUKE|13|1|Now there were some present at that time who told Jesus about the Galileans whose blood Pilate had mixed with their sacrifices.
LUKE|13|2|Jesus answered, "Do you think that these Galileans were worse sinners than all the other Galileans because they suffered this way?
LUKE|13|3|I tell you, no! But unless you repent, you too will all perish.
LUKE|13|4|Or those eighteen who died when the tower in Siloam fell on them--do you think they were more guilty than all the others living in Jerusalem?
LUKE|13|5|I tell you, no! But unless you repent, you too will all perish."
LUKE|13|6|Then he told this parable: "A man had a fig tree, planted in his vineyard, and he went to look for fruit on it, but did not find any.
LUKE|13|7|So he said to the man who took care of the vineyard, 'For three years now I've been coming to look for fruit on this fig tree and haven't found any. Cut it down! Why should it use up the soil?'
LUKE|13|8|"'Sir,' the man replied, 'leave it alone for one more year, and I'll dig around it and fertilize it.
LUKE|13|9|If it bears fruit next year, fine! If not, then cut it down.'"
LUKE|13|10|On a Sabbath Jesus was teaching in one of the synagogues,
LUKE|13|11|and a woman was there who had been crippled by a spirit for eighteen years. She was bent over and could not straighten up at all.
LUKE|13|12|When Jesus saw her, he called her forward and said to her, "Woman, you are set free from your infirmity."
LUKE|13|13|Then he put his hands on her, and immediately she straightened up and praised God.
LUKE|13|14|Indignant because Jesus had healed on the Sabbath, the synagogue ruler said to the people, "There are six days for work. So come and be healed on those days, not on the Sabbath."
LUKE|13|15|The Lord answered him, "You hypocrites! Doesn't each of you on the Sabbath untie his ox or donkey from the stall and lead it out to give it water?
LUKE|13|16|Then should not this woman, a daughter of Abraham, whom Satan has kept bound for eighteen long years, be set free on the Sabbath day from what bound her?"
LUKE|13|17|When he said this, all his opponents were humiliated, but the people were delighted with all the wonderful things he was doing.
LUKE|13|18|Then Jesus asked, "What is the kingdom of God like? What shall I compare it to?
LUKE|13|19|It is like a mustard seed, which a man took and planted in his garden. It grew and became a tree, and the birds of the air perched in its branches."
LUKE|13|20|Again he asked, "What shall I compare the kingdom of God to?
LUKE|13|21|It is like yeast that a woman took and mixed into a large amount of flour until it worked all through the dough."
LUKE|13|22|Then Jesus went through the towns and villages, teaching as he made his way to Jerusalem.
LUKE|13|23|Someone asked him, "Lord, are only a few people going to be saved?"
LUKE|13|24|He said to them, "Make every effort to enter through the narrow door, because many, I tell you, will try to enter and will not be able to.
LUKE|13|25|Once the owner of the house gets up and closes the door, you will stand outside knocking and pleading, 'Sir, open the door for us.'"But he will answer, 'I don't know you or where you come from.'
LUKE|13|26|"Then you will say, 'We ate and drank with you, and you taught in our streets.'
LUKE|13|27|"But he will reply, 'I don't know you or where you come from. Away from me, all you evildoers!'
LUKE|13|28|"There will be weeping there, and gnashing of teeth, when you see Abraham, Isaac and Jacob and all the prophets in the kingdom of God, but you yourselves thrown out.
LUKE|13|29|People will come from east and west and north and south, and will take their places at the feast in the kingdom of God.
LUKE|13|30|Indeed there are those who are last who will be first, and first who will be last."
LUKE|13|31|At that time some Pharisees came to Jesus and said to him, "Leave this place and go somewhere else. Herod wants to kill you."
LUKE|13|32|He replied, "Go tell that fox, 'I will drive out demons and heal people today and tomorrow, and on the third day I will reach my goal.'
LUKE|13|33|In any case, I must keep going today and tomorrow and the next day--for surely no prophet can die outside Jerusalem!
LUKE|13|34|"O Jerusalem, Jerusalem, you who kill the prophets and stone those sent to you, how often I have longed to gather your children together, as a hen gathers her chicks under her wings, but you were not willing!
LUKE|13|35|Look, your house is left to you desolate. I tell you, you will not see me again until you say, 'Blessed is he who comes in the name of the Lord.'"
LUKE|14|1|One Sabbath, when Jesus went to eat in the house of a prominent Pharisee, he was being carefully watched.
LUKE|14|2|There in front of him was a man suffering from dropsy.
LUKE|14|3|Jesus asked the Pharisees and experts in the law, "Is it lawful to heal on the Sabbath or not?"
LUKE|14|4|But they remained silent. So taking hold of the man, he healed him and sent him away.
LUKE|14|5|Then he asked them, "If one of you has a son or an ox that falls into a well on the Sabbath day, will you not immediately pull him out?"
LUKE|14|6|And they had nothing to say.
LUKE|14|7|When he noticed how the guests picked the places of honor at the table, he told them this parable:
LUKE|14|8|"When someone invites you to a wedding feast, do not take the place of honor, for a person more distinguished than you may have been invited.
LUKE|14|9|If so, the host who invited both of you will come and say to you, 'Give this man your seat.' Then, humiliated, you will have to take the least important place.
LUKE|14|10|But when you are invited, take the lowest place, so that when your host comes, he will say to you, 'Friend, move up to a better place.' Then you will be honored in the presence of all your fellow guests.
LUKE|14|11|For everyone who exalts himself will be humbled, and he who humbles himself will be exalted."
LUKE|14|12|Then Jesus said to his host, "When you give a luncheon or dinner, do not invite your friends, your brothers or relatives, or your rich neighbors; if you do, they may invite you back and so you will be repaid.
LUKE|14|13|But when you give a banquet, invite the poor, the crippled, the lame, the blind,
LUKE|14|14|and you will be blessed. Although they cannot repay you, you will be repaid at the resurrection of the righteous."
LUKE|14|15|When one of those at the table with him heard this, he said to Jesus, "Blessed is the man who will eat at the feast in the kingdom of God."
LUKE|14|16|Jesus replied: "A certain man was preparing a great banquet and invited many guests.
LUKE|14|17|At the time of the banquet he sent his servant to tell those who had been invited, 'Come, for everything is now ready.'
LUKE|14|18|"But they all alike began to make excuses. The first said, 'I have just bought a field, and I must go and see it. Please excuse me.'
LUKE|14|19|"Another said, 'I have just bought five yoke of oxen, and I'm on my way to try them out. Please excuse me.'
LUKE|14|20|"Still another said, 'I just got married, so I can't come.'
LUKE|14|21|"The servant came back and reported this to his master. Then the owner of the house became angry and ordered his servant, 'Go out quickly into the streets and alleys of the town and bring in the poor, the crippled, the blind and the lame.'
LUKE|14|22|"'Sir,' the servant said, 'what you ordered has been done, but there is still room.'
LUKE|14|23|"Then the master told his servant, 'Go out to the roads and country lanes and make them come in, so that my house will be full.
LUKE|14|24|I tell you, not one of those men who were invited will get a taste of my banquet.'"
LUKE|14|25|Large crowds were traveling with Jesus, and turning to them he said:
LUKE|14|26|"If anyone comes to me and does not hate his father and mother, his wife and children, his brothers and sisters--yes, even his own life--he cannot be my disciple.
LUKE|14|27|And anyone who does not carry his cross and follow me cannot be my disciple.
LUKE|14|28|"Suppose one of you wants to build a tower. Will he not first sit down and estimate the cost to see if he has enough money to complete it?
LUKE|14|29|For if he lays the foundation and is not able to finish it, everyone who sees it will ridicule him,
LUKE|14|30|saying, 'This fellow began to build and was not able to finish.'
LUKE|14|31|"Or suppose a king is about to go to war against another king. Will he not first sit down and consider whether he is able with ten thousand men to oppose the one coming against him with twenty thousand?
LUKE|14|32|If he is not able, he will send a delegation while the other is still a long way off and will ask for terms of peace.
LUKE|14|33|In the same way, any of you who does not give up everything he has cannot be my disciple.
LUKE|14|34|"Salt is good, but if it loses its saltiness, how can it be made salty again?
LUKE|14|35|It is fit neither for the soil nor for the manure pile; it is thrown out. "He who has ears to hear, let him hear."
LUKE|15|1|Now the tax collectors and "sinners" were all gathering around to hear him.
LUKE|15|2|But the Pharisees and the teachers of the law muttered, "This man welcomes sinners and eats with them."
LUKE|15|3|Then Jesus told them this parable:
LUKE|15|4|"Suppose one of you has a hundred sheep and loses one of them. Does he not leave the ninety-nine in the open country and go after the lost sheep until he finds it?
LUKE|15|5|And when he finds it, he joyfully puts it on his shoulders
LUKE|15|6|and goes home. Then he calls his friends and neighbors together and says, 'Rejoice with me; I have found my lost sheep.'
LUKE|15|7|I tell you that in the same way there will be more rejoicing in heaven over one sinner who repents than over ninety-nine righteous persons who do not need to repent.
LUKE|15|8|"Or suppose a woman has ten silver coins and loses one. Does she not light a lamp, sweep the house and search carefully until she finds it?
LUKE|15|9|And when she finds it, she calls her friends and neighbors together and says, 'Rejoice with me; I have found my lost coin.'
LUKE|15|10|In the same way, I tell you, there is rejoicing in the presence of the angels of God over one sinner who repents."
LUKE|15|11|Jesus continued: "There was a man who had two sons.
LUKE|15|12|The younger one said to his father, 'Father, give me my share of the estate.' So he divided his property between them.
LUKE|15|13|"Not long after that, the younger son got together all he had, set off for a distant country and there squandered his wealth in wild living.
LUKE|15|14|After he had spent everything, there was a severe famine in that whole country, and he began to be in need.
LUKE|15|15|So he went and hired himself out to a citizen of that country, who sent him to his fields to feed pigs.
LUKE|15|16|He longed to fill his stomach with the pods that the pigs were eating, but no one gave him anything.
LUKE|15|17|"When he came to his senses, he said, 'How many of my father's hired men have food to spare, and here I am starving to death!
LUKE|15|18|I will set out and go back to my father and say to him: Father, I have sinned against heaven and against you.
LUKE|15|19|I am no longer worthy to be called your son; make me like one of your hired men.'
LUKE|15|20|So he got up and went to his father. "But while he was still a long way off, his father saw him and was filled with compassion for him; he ran to his son, threw his arms around him and kissed him.
LUKE|15|21|"The son said to him, 'Father, I have sinned against heaven and against you. I am no longer worthy to be called your son. '
LUKE|15|22|"But the father said to his servants, 'Quick! Bring the best robe and put it on him. Put a ring on his finger and sandals on his feet.
LUKE|15|23|Bring the fattened calf and kill it. Let's have a feast and celebrate.
LUKE|15|24|For this son of mine was dead and is alive again; he was lost and is found.' So they began to celebrate.
LUKE|15|25|"Meanwhile, the older son was in the field. When he came near the house, he heard music and dancing.
LUKE|15|26|So he called one of the servants and asked him what was going on.
LUKE|15|27|'Your brother has come,' he replied, 'and your father has killed the fattened calf because he has him back safe and sound.'
LUKE|15|28|"The older brother became angry and refused to go in. So his father went out and pleaded with him.
LUKE|15|29|But he answered his father, 'Look! All these years I've been slaving for you and never disobeyed your orders. Yet you never gave me even a young goat so I could celebrate with my friends.
LUKE|15|30|But when this son of yours who has squandered your property with prostitutes comes home, you kill the fattened calf for him!'
LUKE|15|31|"'My son,' the father said, 'you are always with me, and everything I have is yours.
LUKE|15|32|But we had to celebrate and be glad, because this brother of yours was dead and is alive again; he was lost and is found.'"
LUKE|16|1|Jesus told his disciples: "There was a rich man whose manager was accused of wasting his possessions.
LUKE|16|2|So he called him in and asked him, 'What is this I hear about you? Give an account of your management, because you cannot be manager any longer.'
LUKE|16|3|"The manager said to himself, 'What shall I do now? My master is taking away my job. I'm not strong enough to dig, and I'm ashamed to beg--
LUKE|16|4|I know what I'll do so that, when I lose my job here, people will welcome me into their houses.'
LUKE|16|5|"So he called in each one of his master's debtors. He asked the first, 'How much do you owe my master?'
LUKE|16|6|"'Eight hundred gallons of olive oil,' he replied. "The manager told him, 'Take your bill, sit down quickly, and make it four hundred.'
LUKE|16|7|"Then he asked the second, 'And how much do you owe?'"'A thousand bushels of wheat,' he replied. "He told him, 'Take your bill and make it eight hundred.'
LUKE|16|8|"The master commended the dishonest manager because he had acted shrewdly. For the people of this world are more shrewd in dealing with their own kind than are the people of the light.
LUKE|16|9|I tell you, use worldly wealth to gain friends for yourselves, so that when it is gone, you will be welcomed into eternal dwellings.
LUKE|16|10|"Whoever can be trusted with very little can also be trusted with much, and whoever is dishonest with very little will also be dishonest with much.
LUKE|16|11|So if you have not been trustworthy in handling worldly wealth, who will trust you with true riches?
LUKE|16|12|And if you have not been trustworthy with someone else's property, who will give you property of your own?
LUKE|16|13|"No servant can serve two masters. Either he will hate the one and love the other, or he will be devoted to the one and despise the other. You cannot serve both God and Money."
LUKE|16|14|The Pharisees, who loved money, heard all this and were sneering at Jesus.
LUKE|16|15|He said to them, "You are the ones who justify yourselves in the eyes of men, but God knows your hearts. What is highly valued among men is detestable in God's sight.
LUKE|16|16|"The Law and the Prophets were proclaimed until John. Since that time, the good news of the kingdom of God is being preached, and everyone is forcing his way into it.
LUKE|16|17|It is easier for heaven and earth to disappear than for the least stroke of a pen to drop out of the Law.
LUKE|16|18|"Anyone who divorces his wife and marries another woman commits adultery, and the man who marries a divorced woman commits adultery.
LUKE|16|19|"There was a rich man who was dressed in purple and fine linen and lived in luxury every day.
LUKE|16|20|At his gate was laid a beggar named Lazarus, covered with sores
LUKE|16|21|and longing to eat what fell from the rich man's table. Even the dogs came and licked his sores.
LUKE|16|22|"The time came when the beggar died and the angels carried him to Abraham's side. The rich man also died and was buried.
LUKE|16|23|In hell, where he was in torment, he looked up and saw Abraham far away, with Lazarus by his side.
LUKE|16|24|So he called to him, 'Father Abraham, have pity on me and send Lazarus to dip the tip of his finger in water and cool my tongue, because I am in agony in this fire.'
LUKE|16|25|"But Abraham replied, 'Son, remember that in your lifetime you received your good things, while Lazarus received bad things, but now he is comforted here and you are in agony.
LUKE|16|26|And besides all this, between us and you a great chasm has been fixed, so that those who want to go from here to you cannot, nor can anyone cross over from there to us.'
LUKE|16|27|"He answered, 'Then I beg you, father, send Lazarus to my father's house,
LUKE|16|28|for I have five brothers. Let him warn them, so that they will not also come to this place of torment.'
LUKE|16|29|"Abraham replied, 'They have Moses and the Prophets; let them listen to them.'
LUKE|16|30|"'No, father Abraham,' he said, 'but if someone from the dead goes to them, they will repent.'
LUKE|16|31|"He said to him, 'If they do not listen to Moses and the Prophets, they will not be convinced even if someone rises from the dead.'"
LUKE|17|1|Jesus said to his disciples: "Things that cause people to sin are bound to come, but woe to that person through whom they come.
LUKE|17|2|It would be better for him to be thrown into the sea with a millstone tied around his neck than for him to cause one of these little ones to sin.
LUKE|17|3|So watch yourselves. "If your brother sins, rebuke him, and if he repents, forgive him.
LUKE|17|4|If he sins against you seven times in a day, and seven times comes back to you and says, 'I repent,' forgive him."
LUKE|17|5|The apostles said to the Lord, "Increase our faith!"
LUKE|17|6|He replied, "If you have faith as small as a mustard seed, you can say to this mulberry tree, 'Be uprooted and planted in the sea,' and it will obey you.
LUKE|17|7|"Suppose one of you had a servant plowing or looking after the sheep. Would he say to the servant when he comes in from the field, 'Come along now and sit down to eat'?
LUKE|17|8|Would he not rather say, 'Prepare my supper, get yourself ready and wait on me while I eat and drink; after that you may eat and drink'?
LUKE|17|9|Would he thank the servant because he did what he was told to do?
LUKE|17|10|So you also, when you have done everything you were told to do, should say, 'We are unworthy servants; we have only done our duty.'"
LUKE|17|11|Now on his way to Jerusalem, Jesus traveled along the border between Samaria and Galilee.
LUKE|17|12|As he was going into a village, ten men who had leprosy met him. They stood at a distance
LUKE|17|13|and called out in a loud voice, "Jesus, Master, have pity on us!"
LUKE|17|14|When he saw them, he said, "Go, show yourselves to the priests." And as they went, they were cleansed.
LUKE|17|15|One of them, when he saw he was healed, came back, praising God in a loud voice.
LUKE|17|16|He threw himself at Jesus' feet and thanked him--and he was a Samaritan.
LUKE|17|17|Jesus asked, "Were not all ten cleansed? Where are the other nine?
LUKE|17|18|Was no one found to return and give praise to God except this foreigner?"
LUKE|17|19|Then he said to him, "Rise and go; your faith has made you well."
LUKE|17|20|Once, having been asked by the Pharisees when the kingdom of God would come, Jesus replied, "The kingdom of God does not come with your careful observation,
LUKE|17|21|nor will people say, 'Here it is,' or 'There it is,' because the kingdom of God is within you."
LUKE|17|22|Then he said to his disciples, "The time is coming when you will long to see one of the days of the Son of Man, but you will not see it.
LUKE|17|23|Men will tell you, 'There he is!' or 'Here he is!' Do not go running off after them.
LUKE|17|24|For the Son of Man in his day will be like the lightning, which flashes and lights up the sky from one end to the other.
LUKE|17|25|But first he must suffer many things and be rejected by this generation.
LUKE|17|26|"Just as it was in the days of Noah, so also will it be in the days of the Son of Man.
LUKE|17|27|People were eating, drinking, marrying and being given in marriage up to the day Noah entered the ark. Then the flood came and destroyed them all.
LUKE|17|28|"It was the same in the days of Lot. People were eating and drinking, buying and selling, planting and building.
LUKE|17|29|But the day Lot left Sodom, fire and sulfur rained down from heaven and destroyed them all.
LUKE|17|30|"It will be just like this on the day the Son of Man is revealed.
LUKE|17|31|On that day no one who is on the roof of his house, with his goods inside, should go down to get them. Likewise, no one in the field should go back for anything.
LUKE|17|32|Remember Lot's wife!
LUKE|17|33|Whoever tries to keep his life will lose it, and whoever loses his life will preserve it.
LUKE|17|34|I tell you, on that night two people will be in one bed; one will be taken and the other left.
LUKE|17|35|Two women will be grinding grain together; one will be taken and the other left."
LUKE|17|36|See Footnote
LUKE|17|37|"Where, Lord?" they asked. He replied, "Where there is a dead body, there the vultures will gather."
LUKE|18|1|Then Jesus told his disciples a parable to show them that they should always pray and not give up.
LUKE|18|2|He said: "In a certain town there was a judge who neither feared God nor cared about men.
LUKE|18|3|And there was a widow in that town who kept coming to him with the plea, 'Grant me justice against my adversary.'
LUKE|18|4|"For some time he refused. But finally he said to himself, 'Even though I don't fear God or care about men,
LUKE|18|5|yet because this widow keeps bothering me, I will see that she gets justice, so that she won't eventually wear me out with her coming!'"
LUKE|18|6|And the Lord said, "Listen to what the unjust judge says.
LUKE|18|7|And will not God bring about justice for his chosen ones, who cry out to him day and night? Will he keep putting them off?
LUKE|18|8|I tell you, he will see that they get justice, and quickly. However, when the Son of Man comes, will he find faith on the earth?"
LUKE|18|9|To some who were confident of their own righteousness and looked down on everybody else, Jesus told this parable:
LUKE|18|10|"Two men went up to the temple to pray, one a Pharisee and the other a tax collector.
LUKE|18|11|The Pharisee stood up and prayed about himself: 'God, I thank you that I am not like other men--robbers, evildoers, adulterers--or even like this tax collector.
LUKE|18|12|I fast twice a week and give a tenth of all I get.'
LUKE|18|13|"But the tax collector stood at a distance. He would not even look up to heaven, but beat his breast and said, 'God, have mercy on me, a sinner.'
LUKE|18|14|"I tell you that this man, rather than the other, went home justified before God. For everyone who exalts himself will be humbled, and he who humbles himself will be exalted."
LUKE|18|15|People were also bringing babies to Jesus to have him touch them. When the disciples saw this, they rebuked them.
LUKE|18|16|But Jesus called the children to him and said, "Let the little children come to me, and do not hinder them, for the kingdom of God belongs to such as these.
LUKE|18|17|I tell you the truth, anyone who will not receive the kingdom of God like a little child will never enter it."
LUKE|18|18|A certain ruler asked him, "Good teacher, what must I do to inherit eternal life?"
LUKE|18|19|"Why do you call me good?" Jesus answered. "No one is good--except God alone.
LUKE|18|20|You know the commandments: 'Do not commit adultery, do not murder, do not steal, do not give false testimony, honor your father and mother.'"
LUKE|18|21|"All these I have kept since I was a boy," he said.
LUKE|18|22|When Jesus heard this, he said to him, "You still lack one thing. Sell everything you have and give to the poor, and you will have treasure in heaven. Then come, follow me."
LUKE|18|23|When he heard this, he became very sad, because he was a man of great wealth.
LUKE|18|24|Jesus looked at him and said, "How hard it is for the rich to enter the kingdom of God!
LUKE|18|25|Indeed, it is easier for a camel to go through the eye of a needle than for a rich man to enter the kingdom of God."
LUKE|18|26|Those who heard this asked, "Who then can be saved?"
LUKE|18|27|Jesus replied, "What is impossible with men is possible with God."
LUKE|18|28|Peter said to him, "We have left all we had to follow you!"
LUKE|18|29|"I tell you the truth," Jesus said to them, "no one who has left home or wife or brothers or parents or children for the sake of the kingdom of God
LUKE|18|30|will fail to receive many times as much in this age and, in the age to come, eternal life."
LUKE|18|31|Jesus took the Twelve aside and told them, "We are going up to Jerusalem, and everything that is written by the prophets about the Son of Man will be fulfilled.
LUKE|18|32|He will be handed over to the Gentiles. They will mock him, insult him, spit on him, flog him and kill him.
LUKE|18|33|On the third day he will rise again."
LUKE|18|34|The disciples did not understand any of this. Its meaning was hidden from them, and they did not know what he was talking about.
LUKE|18|35|As Jesus approached Jericho, a blind man was sitting by the roadside begging.
LUKE|18|36|When he heard the crowd going by, he asked what was happening.
LUKE|18|37|They told him, "Jesus of Nazareth is passing by."
LUKE|18|38|He called out, "Jesus, Son of David, have mercy on me!"
LUKE|18|39|Those who led the way rebuked him and told him to be quiet, but he shouted all the more, "Son of David, have mercy on me!"
LUKE|18|40|Jesus stopped and ordered the man to be brought to him. When he came near, Jesus asked him,
LUKE|18|41|"What do you want me to do for you?Lord, I want to see," he replied.
LUKE|18|42|Jesus said to him, "Receive your sight; your faith has healed you."
LUKE|18|43|Immediately he received his sight and followed Jesus, praising God. When all the people saw it, they also praised God.
LUKE|19|1|Jesus entered Jericho and was passing through.
LUKE|19|2|A man was there by the name of Zacchaeus; he was a chief tax collector and was wealthy.
LUKE|19|3|He wanted to see who Jesus was, but being a short man he could not, because of the crowd.
LUKE|19|4|So he ran ahead and climbed a sycamore-fig tree to see him, since Jesus was coming that way.
LUKE|19|5|When Jesus reached the spot, he looked up and said to him, "Zacchaeus, come down immediately. I must stay at your house today."
LUKE|19|6|So he came down at once and welcomed him gladly.
LUKE|19|7|All the people saw this and began to mutter, "He has gone to be the guest of a 'sinner.'"
LUKE|19|8|But Zacchaeus stood up and said to the Lord, "Look, Lord! Here and now I give half of my possessions to the poor, and if I have cheated anybody out of anything, I will pay back four times the amount."
LUKE|19|9|Jesus said to him, "Today salvation has come to this house, because this man, too, is a son of Abraham.
LUKE|19|10|For the Son of Man came to seek and to save what was lost."
LUKE|19|11|While they were listening to this, he went on to tell them a parable, because he was near Jerusalem and the people thought that the kingdom of God was going to appear at once.
LUKE|19|12|He said: "A man of noble birth went to a distant country to have himself appointed king and then to return.
LUKE|19|13|So he called ten of his servants and gave them ten minas. 'Put this money to work,' he said, 'until I come back.'
LUKE|19|14|"But his subjects hated him and sent a delegation after him to say, 'We don't want this man to be our king.'
LUKE|19|15|"He was made king, however, and returned home. Then he sent for the servants to whom he had given the money, in order to find out what they had gained with it.
LUKE|19|16|"The first one came and said, 'Sir, your mina has earned ten more.'
LUKE|19|17|"'Well done, my good servant!' his master replied. 'Because you have been trustworthy in a very small matter, take charge of ten cities.'
LUKE|19|18|"The second came and said, 'Sir, your mina has earned five more.'
LUKE|19|19|"His master answered, 'You take charge of five cities.'
LUKE|19|20|"Then another servant came and said, 'Sir, here is your mina; I have kept it laid away in a piece of cloth.
LUKE|19|21|I was afraid of you, because you are a hard man. You take out what you did not put in and reap what you did not sow.'
LUKE|19|22|"His master replied, 'I will judge you by your own words, you wicked servant! You knew, did you, that I am a hard man, taking out what I did not put in, and reaping what I did not sow?
LUKE|19|23|Why then didn't you put my money on deposit, so that when I came back, I could have collected it with interest?'
LUKE|19|24|"Then he said to those standing by, 'Take his mina away from him and give it to the one who has ten minas.'
LUKE|19|25|"'Sir,' they said, 'he already has ten!'
LUKE|19|26|"He replied, 'I tell you that to everyone who has, more will be given, but as for the one who has nothing, even what he has will be taken away.
LUKE|19|27|But those enemies of mine who did not want me to be king over them--bring them here and kill them in front of me.'"
LUKE|19|28|After Jesus had said this, he went on ahead, going up to Jerusalem.
LUKE|19|29|As he approached Bethphage and Bethany at the hill called the Mount of Olives, he sent two of his disciples, saying to them,
LUKE|19|30|"Go to the village ahead of you, and as you enter it, you will find a colt tied there, which no one has ever ridden. Untie it and bring it here.
LUKE|19|31|If anyone asks you, 'Why are you untying it?' tell him, 'The Lord needs it.'"
LUKE|19|32|Those who were sent ahead went and found it just as he had told them.
LUKE|19|33|As they were untying the colt, its owners asked them, "Why are you untying the colt?"
LUKE|19|34|They replied, "The Lord needs it."
LUKE|19|35|They brought it to Jesus, threw their cloaks on the colt and put Jesus on it.
LUKE|19|36|As he went along, people spread their cloaks on the road.
LUKE|19|37|When he came near the place where the road goes down the Mount of Olives, the whole crowd of disciples began joyfully to praise God in loud voices for all the miracles they had seen:
LUKE|19|38|"Blessed is the king who comes in the name of the Lord!Peace in heaven and glory in the highest!"
LUKE|19|39|Some of the Pharisees in the crowd said to Jesus, "Teacher, rebuke your disciples!"
LUKE|19|40|"I tell you," he replied, "if they keep quiet, the stones will cry out."
LUKE|19|41|As he approached Jerusalem and saw the city, he wept over it
LUKE|19|42|and said, "If you, even you, had only known on this day what would bring you peace--but now it is hidden from your eyes.
LUKE|19|43|The days will come upon you when your enemies will build an embankment against you and encircle you and hem you in on every side.
LUKE|19|44|They will dash you to the ground, you and the children within your walls. They will not leave one stone on another, because you did not recognize the time of God's coming to you."
LUKE|19|45|Then he entered the temple area and began driving out those who were selling.
LUKE|19|46|"It is written," he said to them, "'My house will be a house of prayer'; but you have made it 'a den of robbers.'"
LUKE|19|47|Every day he was teaching at the temple. But the chief priests, the teachers of the law and the leaders among the people were trying to kill him.
LUKE|19|48|Yet they could not find any way to do it, because all the people hung on his words.
LUKE|20|1|One day as he was teaching the people in the temple courts and preaching the gospel, the chief priests and the teachers of the law, together with the elders, came up to him.
LUKE|20|2|"Tell us by what authority you are doing these things," they said. "Who gave you this authority?"
LUKE|20|3|He replied, "I will also ask you a question. Tell me,
LUKE|20|4|John's baptism--was it from heaven, or from men?"
LUKE|20|5|They discussed it among themselves and said, "If we say, 'From heaven,' he will ask, 'Why didn't you believe him?'
LUKE|20|6|But if we say, 'From men,' all the people will stone us, because they are persuaded that John was a prophet."
LUKE|20|7|So they answered, "We don't know where it was from."
LUKE|20|8|Jesus said, "Neither will I tell you by what authority I am doing these things."
LUKE|20|9|He went on to tell the people this parable: "A man planted a vineyard, rented it to some farmers and went away for a long time.
LUKE|20|10|At harvest time he sent a servant to the tenants so they would give him some of the fruit of the vineyard. But the tenants beat him and sent him away empty-handed.
LUKE|20|11|He sent another servant, but that one also they beat and treated shamefully and sent away empty-handed.
LUKE|20|12|He sent still a third, and they wounded him and threw him out.
LUKE|20|13|"Then the owner of the vineyard said, 'What shall I do? I will send my son, whom I love; perhaps they will respect him.'
LUKE|20|14|"But when the tenants saw him, they talked the matter over. 'This is the heir,' they said. 'Let's kill him, and the inheritance will be ours.'
LUKE|20|15|So they threw him out of the vineyard and killed him.
LUKE|20|16|"What then will the owner of the vineyard do to them? He will come and kill those tenants and give the vineyard to others." When the people heard this, they said, "May this never be!"
LUKE|20|17|Jesus looked directly at them and asked, "Then what is the meaning of that which is written: "'The stone the builders rejected has become the capstone '?
LUKE|20|18|Everyone who falls on that stone will be broken to pieces, but he on whom it falls will be crushed."
LUKE|20|19|The teachers of the law and the chief priests looked for a way to arrest him immediately, because they knew he had spoken this parable against them. But they were afraid of the people.
LUKE|20|20|Keeping a close watch on him, they sent spies, who pretended to be honest. They hoped to catch Jesus in something he said so that they might hand him over to the power and authority of the governor.
LUKE|20|21|So the spies questioned him: "Teacher, we know that you speak and teach what is right, and that you do not show partiality but teach the way of God in accordance with the truth.
LUKE|20|22|Is it right for us to pay taxes to Caesar or not?"
LUKE|20|23|He saw through their duplicity and said to them,
LUKE|20|24|"Show me a denarius. Whose portrait and inscription are on it?"
LUKE|20|25|"Caesar's," they replied. He said to them, "Then give to Caesar what is Caesar's, and to God what is God's."
LUKE|20|26|They were unable to trap him in what he had said there in public. And astonished by his answer, they became silent.
LUKE|20|27|Some of the Sadducees, who say there is no resurrection, came to Jesus with a question.
LUKE|20|28|"Teacher," they said, "Moses wrote for us that if a man's brother dies and leaves a wife but no children, the man must marry the widow and have children for his brother.
LUKE|20|29|Now there were seven brothers. The first one married a woman and died childless.
LUKE|20|30|The second
LUKE|20|31|and then the third married her, and in the same way the seven died, leaving no children.
LUKE|20|32|Finally, the woman died too.
LUKE|20|33|Now then, at the resurrection whose wife will she be, since the seven were married to her?"
LUKE|20|34|Jesus replied, "The people of this age marry and are given in marriage.
LUKE|20|35|But those who are considered worthy of taking part in that age and in the resurrection from the dead will neither marry nor be given in marriage,
LUKE|20|36|and they can no longer die; for they are like the angels. They are God's children, since they are children of the resurrection.
LUKE|20|37|But in the account of the bush, even Moses showed that the dead rise, for he calls the Lord 'the God of Abraham, and the God of Isaac, and the God of Jacob.'
LUKE|20|38|He is not the God of the dead, but of the living, for to him all are alive."
LUKE|20|39|Some of the teachers of the law responded, "Well said, teacher!"
LUKE|20|40|And no one dared to ask him any more questions.
LUKE|20|41|Then Jesus said to them, "How is it that they say the Christ is the Son of David?
LUKE|20|42|David himself declares in the Book of Psalms: "'The Lord said to my Lord: "Sit at my right hand
LUKE|20|43|until I make your enemies a footstool for your feet."'
LUKE|20|44|David calls him 'Lord.' How then can he be his son?"
LUKE|20|45|While all the people were listening, Jesus said to his disciples,
LUKE|20|46|"Beware of the teachers of the law. They like to walk around in flowing robes and love to be greeted in the marketplaces and have the most important seats in the synagogues and the places of honor at banquets.
LUKE|20|47|They devour widows' houses and for a show make lengthy prayers. Such men will be punished most severely."
LUKE|21|1|As he looked up, Jesus saw the rich putting their gifts into the temple treasury.
LUKE|21|2|He also saw a poor widow put in two very small copper coins.
LUKE|21|3|"I tell you the truth," he said, "this poor widow has put in more than all the others.
LUKE|21|4|All these people gave their gifts out of their wealth; but she out of her poverty put in all she had to live on."
LUKE|21|5|Some of his disciples were remarking about how the temple was adorned with beautiful stones and with gifts dedicated to God. But Jesus said,
LUKE|21|6|"As for what you see here, the time will come when not one stone will be left on another; every one of them will be thrown down."
LUKE|21|7|"Teacher," they asked, "when will these things happen? And what will be the sign that they are about to take place?"
LUKE|21|8|He replied: "Watch out that you are not deceived. For many will come in my name, claiming, 'I am he,' and, 'The time is near.' Do not follow them.
LUKE|21|9|When you hear of wars and revolutions, do not be frightened. These things must happen first, but the end will not come right away."
LUKE|21|10|Then he said to them: "Nation will rise against nation, and kingdom against kingdom.
LUKE|21|11|There will be great earthquakes, famines and pestilences in various places, and fearful events and great signs from heaven.
LUKE|21|12|"But before all this, they will lay hands on you and persecute you. They will deliver you to synagogues and prisons, and you will be brought before kings and governors, and all on account of my name.
LUKE|21|13|This will result in your being witnesses to them.
LUKE|21|14|But make up your mind not to worry beforehand how you will defend yourselves.
LUKE|21|15|For I will give you words and wisdom that none of your adversaries will be able to resist or contradict.
LUKE|21|16|You will be betrayed even by parents, brothers, relatives and friends, and they will put some of you to death.
LUKE|21|17|All men will hate you because of me.
LUKE|21|18|But not a hair of your head will perish.
LUKE|21|19|By standing firm you will gain life.
LUKE|21|20|"When you see Jerusalem being surrounded by armies, you will know that its desolation is near.
LUKE|21|21|Then let those who are in Judea flee to the mountains, let those in the city get out, and let those in the country not enter the city.
LUKE|21|22|For this is the time of punishment in fulfillment of all that has been written.
LUKE|21|23|How dreadful it will be in those days for pregnant women and nursing mothers! There will be great distress in the land and wrath against this people.
LUKE|21|24|They will fall by the sword and will be taken as prisoners to all the nations. Jerusalem will be trampled on by the Gentiles until the times of the Gentiles are fulfilled.
LUKE|21|25|"There will be signs in the sun, moon and stars. On the earth, nations will be in anguish and perplexity at the roaring and tossing of the sea.
LUKE|21|26|Men will faint from terror, apprehensive of what is coming on the world, for the heavenly bodies will be shaken.
LUKE|21|27|At that time they will see the Son of Man coming in a cloud with power and great glory.
LUKE|21|28|When these things begin to take place, stand up and lift up your heads, because your redemption is drawing near."
LUKE|21|29|He told them this parable: "Look at the fig tree and all the trees.
LUKE|21|30|When they sprout leaves, you can see for yourselves and know that summer is near.
LUKE|21|31|Even so, when you see these things happening, you know that the kingdom of God is near.
LUKE|21|32|"I tell you the truth, this generation will certainly not pass away until all these things have happened.
LUKE|21|33|Heaven and earth will pass away, but my words will never pass away.
LUKE|21|34|"Be careful, or your hearts will be weighed down with dissipation, drunkenness and the anxieties of life, and that day will close on you unexpectedly like a trap.
LUKE|21|35|For it will come upon all those who live on the face of the whole earth.
LUKE|21|36|Be always on the watch, and pray that you may be able to escape all that is about to happen, and that you may be able to stand before the Son of Man."
LUKE|21|37|Each day Jesus was teaching at the temple, and each evening he went out to spend the night on the hill called the Mount of Olives,
LUKE|21|38|and all the people came early in the morning to hear him at the temple.
LUKE|22|1|Now the Feast of Unleavened Bread, called the Passover, was approaching,
LUKE|22|2|and the chief priests and the teachers of the law were looking for some way to get rid of Jesus, for they were afraid of the people.
LUKE|22|3|Then Satan entered Judas, called Iscariot, one of the Twelve.
LUKE|22|4|And Judas went to the chief priests and the officers of the temple guard and discussed with them how he might betray Jesus.
LUKE|22|5|They were delighted and agreed to give him money.
LUKE|22|6|He consented, and watched for an opportunity to hand Jesus over to them when no crowd was present.
LUKE|22|7|Then came the day of Unleavened Bread on which the Passover lamb had to be sacrificed.
LUKE|22|8|Jesus sent Peter and John, saying, "Go and make preparations for us to eat the Passover."
LUKE|22|9|"Where do you want us to prepare for it?" they asked.
LUKE|22|10|He replied, "As you enter the city, a man carrying a jar of water will meet you. Follow him to the house that he enters,
LUKE|22|11|and say to the owner of the house, 'The Teacher asks: Where is the guest room, where I may eat the Passover with my disciples?'
LUKE|22|12|He will show you a large upper room, all furnished. Make preparations there."
LUKE|22|13|They left and found things just as Jesus had told them. So they prepared the Passover.
LUKE|22|14|When the hour came, Jesus and his apostles reclined at the table.
LUKE|22|15|And he said to them, "I have eagerly desired to eat this Passover with you before I suffer.
LUKE|22|16|For I tell you, I will not eat it again until it finds fulfillment in the kingdom of God."
LUKE|22|17|After taking the cup, he gave thanks and said, "Take this and divide it among you.
LUKE|22|18|For I tell you I will not drink again of the fruit of the vine until the kingdom of God comes."
LUKE|22|19|And he took bread, gave thanks and broke it, and gave it to them, saying, "This is my body given for you; do this in remembrance of me."
LUKE|22|20|In the same way, after the supper he took the cup, saying, "This cup is the new covenant in my blood, which is poured out for you.
LUKE|22|21|But the hand of him who is going to betray me is with mine on the table.
LUKE|22|22|The Son of Man will go as it has been decreed, but woe to that man who betrays him."
LUKE|22|23|They began to question among themselves which of them it might be who would do this.
LUKE|22|24|Also a dispute arose among them as to which of them was considered to be greatest.
LUKE|22|25|Jesus said to them, "The kings of the Gentiles lord it over them; and those who exercise authority over them call themselves Benefactors.
LUKE|22|26|But you are not to be like that. Instead, the greatest among you should be like the youngest, and the one who rules like the one who serves.
LUKE|22|27|For who is greater, the one who is at the table or the one who serves? Is it not the one who is at the table? But I am among you as one who serves.
LUKE|22|28|You are those who have stood by me in my trials.
LUKE|22|29|And I confer on you a kingdom, just as my Father conferred one on me,
LUKE|22|30|so that you may eat and drink at my table in my kingdom and sit on thrones, judging the twelve tribes of Israel.
LUKE|22|31|"Simon, Simon, Satan has asked to sift you as wheat.
LUKE|22|32|But I have prayed for you, Simon, that your faith may not fail. And when you have turned back, strengthen your brothers."
LUKE|22|33|But he replied, "Lord, I am ready to go with you to prison and to death."
LUKE|22|34|Jesus answered, "I tell you, Peter, before the rooster crows today, you will deny three times that you know me."
LUKE|22|35|Then Jesus asked them, "When I sent you without purse, bag or sandals, did you lack anything?Nothing," they answered.
LUKE|22|36|He said to them, "But now if you have a purse, take it, and also a bag; and if you don't have a sword, sell your cloak and buy one.
LUKE|22|37|It is written: 'And he was numbered with the transgressors'; and I tell you that this must be fulfilled in me. Yes, what is written about me is reaching its fulfillment."
LUKE|22|38|The disciples said, "See, Lord, here are two swords.That is enough," he replied.
LUKE|22|39|Jesus went out as usual to the Mount of Olives, and his disciples followed him.
LUKE|22|40|On reaching the place, he said to them, "Pray that you will not fall into temptation."
LUKE|22|41|He withdrew about a stone's throw beyond them, knelt down and prayed,
LUKE|22|42|"Father, if you are willing, take this cup from me; yet not my will, but yours be done."
LUKE|22|43|An angel from heaven appeared to him and strengthened him.
LUKE|22|44|And being in anguish, he prayed more earnestly, and his sweat was like drops of blood falling to the ground.
LUKE|22|45|When he rose from prayer and went back to the disciples, he found them asleep, exhausted from sorrow.
LUKE|22|46|"Why are you sleeping?" he asked them. "Get up and pray so that you will not fall into temptation."
LUKE|22|47|While he was still speaking a crowd came up, and the man who was called Judas, one of the Twelve, was leading them. He approached Jesus to kiss him,
LUKE|22|48|but Jesus asked him, "Judas, are you betraying the Son of Man with a kiss?"
LUKE|22|49|When Jesus' followers saw what was going to happen, they said, "Lord, should we strike with our swords?"
LUKE|22|50|And one of them struck the servant of the high priest, cutting off his right ear.
LUKE|22|51|But Jesus answered, "No more of this!" And he touched the man's ear and healed him.
LUKE|22|52|Then Jesus said to the chief priests, the officers of the temple guard, and the elders, who had come for him, "Am I leading a rebellion, that you have come with swords and clubs?
LUKE|22|53|Every day I was with you in the temple courts, and you did not lay a hand on me. But this is your hour--when darkness reigns."
LUKE|22|54|Then seizing him, they led him away and took him into the house of the high priest. Peter followed at a distance.
LUKE|22|55|But when they had kindled a fire in the middle of the courtyard and had sat down together, Peter sat down with them.
LUKE|22|56|A servant girl saw him seated there in the firelight. She looked closely at him and said, "This man was with him."
LUKE|22|57|But he denied it. "Woman, I don't know him," he said.
LUKE|22|58|A little later someone else saw him and said, "You also are one of them.Man, I am not!" Peter replied.
LUKE|22|59|About an hour later another asserted, "Certainly this fellow was with him, for he is a Galilean."
LUKE|22|60|Peter replied, "Man, I don't know what you're talking about!" Just as he was speaking, the rooster crowed.
LUKE|22|61|The Lord turned and looked straight at Peter. Then Peter remembered the word the Lord had spoken to him: "Before the rooster crows today, you will disown me three times."
LUKE|22|62|And he went outside and wept bitterly.
LUKE|22|63|The men who were guarding Jesus began mocking and beating him.
LUKE|22|64|They blindfolded him and demanded, "Prophesy! Who hit you?"
LUKE|22|65|And they said many other insulting things to him.
LUKE|22|66|At daybreak the council of the elders of the people, both the chief priests and teachers of the law, met together, and Jesus was led before them.
LUKE|22|67|"If you are the Christ, "they said, "tell us."
LUKE|22|68|Jesus answered, "If I tell you, you will not believe me, and if I asked you, you would not answer.
LUKE|22|69|But from now on, the Son of Man will be seated at the right hand of the mighty God."
LUKE|22|70|They all asked, "Are you then the Son of God?" He replied, "You are right in saying I am."
LUKE|22|71|Then they said, "Why do we need any more testimony? We have heard it from his own lips."
LUKE|23|1|Then the whole assembly rose and led him off to Pilate.
LUKE|23|2|And they began to accuse him, saying, "We have found this man subverting our nation. He opposes payment of taxes to Caesar and claims to be Christ, a king."
LUKE|23|3|So Pilate asked Jesus, "Are you the king of the Jews?Yes, it is as you say," Jesus replied.
LUKE|23|4|Then Pilate announced to the chief priests and the crowd, "I find no basis for a charge against this man."
LUKE|23|5|But they insisted, "He stirs up the people all over Judea by his teaching. He started in Galilee and has come all the way here."
LUKE|23|6|On hearing this, Pilate asked if the man was a Galilean.
LUKE|23|7|When he learned that Jesus was under Herod's jurisdiction, he sent him to Herod, who was also in Jerusalem at that time.
LUKE|23|8|When Herod saw Jesus, he was greatly pleased, because for a long time he had been wanting to see him. From what he had heard about him, he hoped to see him perform some miracle.
LUKE|23|9|He plied him with many questions, but Jesus gave him no answer.
LUKE|23|10|The chief priests and the teachers of the law were standing there, vehemently accusing him.
LUKE|23|11|Then Herod and his soldiers ridiculed and mocked him. Dressing him in an elegant robe, they sent him back to Pilate.
LUKE|23|12|That day Herod and Pilate became friends--before this they had been enemies.
LUKE|23|13|Pilate called together the chief priests, the rulers and the people,
LUKE|23|14|and said to them, "You brought me this man as one who was inciting the people to rebellion. I have examined him in your presence and have found no basis for your charges against him.
LUKE|23|15|Neither has Herod, for he sent him back to us; as you can see, he has done nothing to deserve death.
LUKE|23|16|Therefore, I will punish him and then release him."
LUKE|23|17|See Footnote
LUKE|23|18|With one voice they cried out, "Away with this man! Release Barabbas to us!"
LUKE|23|19|(Barabbas had been thrown into prison for an insurrection in the city, and for murder.)
LUKE|23|20|Wanting to release Jesus, Pilate appealed to them again.
LUKE|23|21|But they kept shouting, "Crucify him! Crucify him!"
LUKE|23|22|For the third time he spoke to them: "Why? What crime has this man committed? I have found in him no grounds for the death penalty. Therefore I will have him punished and then release him."
LUKE|23|23|But with loud shouts they insistently demanded that he be crucified, and their shouts prevailed.
LUKE|23|24|So Pilate decided to grant their demand.
LUKE|23|25|He released the man who had been thrown into prison for insurrection and murder, the one they asked for, and surrendered Jesus to their will.
LUKE|23|26|As they led him away, they seized Simon from Cyrene, who was on his way in from the country, and put the cross on him and made him carry it behind Jesus.
LUKE|23|27|A large number of people followed him, including women who mourned and wailed for him.
LUKE|23|28|Jesus turned and said to them, "Daughters of Jerusalem, do not weep for me; weep for yourselves and for your children.
LUKE|23|29|For the time will come when you will say, 'Blessed are the barren women, the wombs that never bore and the breasts that never nursed!'
LUKE|23|30|Then "'they will say to the mountains, "Fall on us!" and to the hills, "Cover us!"'
LUKE|23|31|For if men do these things when the tree is green, what will happen when it is dry?"
LUKE|23|32|Two other men, both criminals, were also led out with him to be executed.
LUKE|23|33|When they came to the place called the Skull, there they crucified him, along with the criminals--one on his right, the other on his left.
LUKE|23|34|Jesus said, "Father, forgive them, for they do not know what they are doing." And they divided up his clothes by casting lots.
LUKE|23|35|The people stood watching, and the rulers even sneered at him. They said, "He saved others; let him save himself if he is the Christ of God, the Chosen One."
LUKE|23|36|The soldiers also came up and mocked him. They offered him wine vinegar
LUKE|23|37|and said, "If you are the king of the Jews, save yourself."
LUKE|23|38|There was a written notice above him, which read:|sc THIS IS THE KING OF THE JEWS.
LUKE|23|39|One of the criminals who hung there hurled insults at him: "Aren't you the Christ? Save yourself and us!"
LUKE|23|40|But the other criminal rebuked him. "Don't you fear God," he said, "since you are under the same sentence?
LUKE|23|41|We are punished justly, for we are getting what our deeds deserve. But this man has done nothing wrong."
LUKE|23|42|Then he said, "Jesus, remember me when you come into your kingdom. "
LUKE|23|43|Jesus answered him, "I tell you the truth, today you will be with me in paradise."
LUKE|23|44|It was now about the sixth hour, and darkness came over the whole land until the ninth hour,
LUKE|23|45|for the sun stopped shining. And the curtain of the temple was torn in two.
LUKE|23|46|Jesus called out with a loud voice, "Father, into your hands I commit my spirit." When he had said this, he breathed his last.
LUKE|23|47|The centurion, seeing what had happened, praised God and said, "Surely this was a righteous man."
LUKE|23|48|When all the people who had gathered to witness this sight saw what took place, they beat their breasts and went away.
LUKE|23|49|But all those who knew him, including the women who had followed him from Galilee, stood at a distance, watching these things.
LUKE|23|50|Now there was a man named Joseph, a member of the Council, a good and upright man,
LUKE|23|51|who had not consented to their decision and action. He came from the Judean town of Arimathea and he was waiting for the kingdom of God.
LUKE|23|52|Going to Pilate, he asked for Jesus' body.
LUKE|23|53|Then he took it down, wrapped it in linen cloth and placed it in a tomb cut in the rock, one in which no one had yet been laid.
LUKE|23|54|It was Preparation Day, and the Sabbath was about to begin.
LUKE|23|55|The women who had come with Jesus from Galilee followed Joseph and saw the tomb and how his body was laid in it.
LUKE|23|56|Then they went home and prepared spices and perfumes. But they rested on the Sabbath in obedience to the commandment.
LUKE|24|1|On the first day of the week, very early in the morning, the women took the spices they had prepared and went to the tomb.
LUKE|24|2|They found the stone rolled away from the tomb,
LUKE|24|3|but when they entered, they did not find the body of the Lord Jesus.
LUKE|24|4|While they were wondering about this, suddenly two men in clothes that gleamed like lightning stood beside them.
LUKE|24|5|In their fright the women bowed down with their faces to the ground, but the men said to them, "Why do you look for the living among the dead?
LUKE|24|6|He is not here; he has risen! Remember how he told you, while he was still with you in Galilee:
LUKE|24|7|'The Son of Man must be delivered into the hands of sinful men, be crucified and on the third day be raised again.'"
LUKE|24|8|Then they remembered his words.
LUKE|24|9|When they came back from the tomb, they told all these things to the Eleven and to all the others.
LUKE|24|10|It was Mary Magdalene, Joanna, Mary the mother of James, and the others with them who told this to the apostles.
LUKE|24|11|But they did not believe the women, because their words seemed to them like nonsense.
LUKE|24|12|Peter, however, got up and ran to the tomb. Bending over, he saw the strips of linen lying by themselves, and he went away, wondering to himself what had happened.
LUKE|24|13|Now that same day two of them were going to a village called Emmaus, about seven miles from Jerusalem.
LUKE|24|14|They were talking with each other about everything that had happened.
LUKE|24|15|As they talked and discussed these things with each other, Jesus himself came up and walked along with them;
LUKE|24|16|but they were kept from recognizing him.
LUKE|24|17|He asked them, "What are you discussing together as you walk along?"
LUKE|24|18|They stood still, their faces downcast. One of them, named Cleopas, asked him, "Are you only a visitor to Jerusalem and do not know the things that have happened there in these days?"
LUKE|24|19|"What things?" he asked.
LUKE|24|20|"About Jesus of Nazareth," they replied. "He was a prophet, powerful in word and deed before God and all the people. The chief priests and our rulers handed him over to be sentenced to death, and they crucified him;
LUKE|24|21|but we had hoped that he was the one who was going to redeem Israel. And what is more, it is the third day since all this took place.
LUKE|24|22|In addition, some of our women amazed us. They went to the tomb early this morning
LUKE|24|23|but didn't find his body. They came and told us that they had seen a vision of angels, who said he was alive.
LUKE|24|24|Then some of our companions went to the tomb and found it just as the women had said, but him they did not see."
LUKE|24|25|He said to them, "How foolish you are, and how slow of heart to believe all that the prophets have spoken!
LUKE|24|26|Did not the Christ have to suffer these things and then enter his glory?"
LUKE|24|27|And beginning with Moses and all the Prophets, he explained to them what was said in all the Scriptures concerning himself.
LUKE|24|28|As they approached the village to which they were going, Jesus acted as if he were going farther.
LUKE|24|29|But they urged him strongly, "Stay with us, for it is nearly evening; the day is almost over." So he went in to stay with them.
LUKE|24|30|When he was at the table with them, he took bread, gave thanks, broke it and began to give it to them.
LUKE|24|31|Then their eyes were opened and they recognized him, and he disappeared from their sight.
LUKE|24|32|They asked each other, "Were not our hearts burning within us while he talked with us on the road and opened the Scriptures to us?"
LUKE|24|33|They got up and returned at once to Jerusalem. There they found the Eleven and those with them, assembled together
LUKE|24|34|and saying, "It is true! The Lord has risen and has appeared to Simon."
LUKE|24|35|Then the two told what had happened on the way, and how Jesus was recognized by them when he broke the bread.
LUKE|24|36|While they were still talking about this, Jesus himself stood among them and said to them, "Peace be with you."
LUKE|24|37|They were startled and frightened, thinking they saw a ghost.
LUKE|24|38|He said to them, "Why are you troubled, and why do doubts rise in your minds?
LUKE|24|39|Look at my hands and my feet. It is I myself! Touch me and see; a ghost does not have flesh and bones, as you see I have."
LUKE|24|40|When he had said this, he showed them his hands and feet.
LUKE|24|41|And while they still did not believe it because of joy and amazement, he asked them, "Do you have anything here to eat?"
LUKE|24|42|They gave him a piece of broiled fish,
LUKE|24|43|and he took it and ate it in their presence.
LUKE|24|44|He said to them, "This is what I told you while I was still with you: Everything must be fulfilled that is written about me in the Law of Moses, the Prophets and the Psalms."
LUKE|24|45|Then he opened their minds so they could understand the Scriptures.
LUKE|24|46|He told them, "This is what is written: The Christ will suffer and rise from the dead on the third day,
LUKE|24|47|and repentance and forgiveness of sins will be preached in his name to all nations, beginning at Jerusalem.
LUKE|24|48|You are witnesses of these things.
LUKE|24|49|I am going to send you what my Father has promised; but stay in the city until you have been clothed with power from on high."
LUKE|24|50|When he had led them out to the vicinity of Bethany, he lifted up his hands and blessed them.
LUKE|24|51|While he was blessing them, he left them and was taken up into heaven.
LUKE|24|52|Then they worshiped him and returned to Jerusalem with great joy.
LUKE|24|53|And they stayed continually at the temple, praising God.
