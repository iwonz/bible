PHIL|1|1|Павел и Тимофей, рабы Иисуса Христа, всем святым во Христе Иисусе, находящимся в Филиппах, с епископами и диаконами:
PHIL|1|2|благодать вам и мир от Бога Отца нашего и Господа Иисуса Христа.
PHIL|1|3|Благодарю Бога моего при всяком воспоминании о вас,
PHIL|1|4|всегда во всякой молитве моей за всех вас принося с радостью молитву мою,
PHIL|1|5|за ваше участие в благовествовании от первого дня даже доныне,
PHIL|1|6|будучи уверен в том, что начавший в вас доброе дело будет совершать его даже до дня Иисуса Христа,
PHIL|1|7|как и должно мне помышлять о всех вас, потому что я имею вас в сердце в узах моих, при защищении и утверждении благовествования, вас всех, как соучастников моих в благодати.
PHIL|1|8|Бог – свидетель, что я люблю всех вас любовью Иисуса Христа;
PHIL|1|9|и молюсь о том, чтобы любовь ваша еще более и более возрастала в познании и всяком чувстве,
PHIL|1|10|чтобы, познавая лучшее, вы были чисты и непреткновенны в день Христов,
PHIL|1|11|исполнены плодов праведности Иисусом Христом, в славу и похвалу Божию.
PHIL|1|12|Желаю, братия, чтобы вы знали, что обстоятельства мои послужили к большему успеху благовествования,
PHIL|1|13|так что узы мои о Христе сделались известными всей претории и всем прочим,
PHIL|1|14|и большая часть из братьев в Господе, ободрившись узами моими, начали с большею смелостью, безбоязненно проповедывать слово Божие.
PHIL|1|15|Некоторые, правда, по зависти и любопрению, а другие с добрым расположением проповедуют Христа.
PHIL|1|16|Одни по любопрению проповедуют Христа не чисто, думая увеличить тяжесть уз моих;
PHIL|1|17|а другие – из любви, зная, что я поставлен защищать благовествование.
PHIL|1|18|Но что до того? Как бы ни проповедали Христа, притворно или искренно, я и тому радуюсь и буду радоваться,
PHIL|1|19|ибо знаю, что это послужит мне во спасение по вашей молитве и содействием Духа Иисуса Христа,
PHIL|1|20|при уверенности и надежде моей, что я ни в чем посрамлен не буду, но при всяком дерзновении, и ныне, как и всегда, возвеличится Христос в теле моем, жизнью ли то, или смертью.
PHIL|1|21|Ибо для меня жизнь – Христос, и смерть – приобретение.
PHIL|1|22|Если же жизнь во плоти [доставляет] плод моему делу, то не знаю, что избрать.
PHIL|1|23|Влечет меня то и другое: имею желание разрешиться и быть со Христом, потому что это несравненно лучше;
PHIL|1|24|а оставаться во плоти нужнее для вас.
PHIL|1|25|И я верно знаю, что останусь и пребуду со всеми вами для вашего успеха и радости в вере,
PHIL|1|26|дабы похвала ваша во Христе Иисусе умножилась через меня, при моем вторичном к вам пришествии.
PHIL|1|27|Только живите достойно благовествования Христова, чтобы мне, приду ли я и увижу вас, или не приду, слышать о вас, что вы стоите в одном духе, подвизаясь единодушно за веру Евангельскую,
PHIL|1|28|и не страшитесь ни в чем противников: это для них есть предзнаменование погибели, а для вас – спасения. И сие от Бога,
PHIL|1|29|потому что вам дано ради Христа не только веровать в Него, но и страдать за Него
PHIL|1|30|таким же подвигом, какой вы видели во мне и ныне слышите о мне.
PHIL|2|1|Итак, если [есть] какое утешение во Христе, если [есть] какая отрада любви, если [есть] какое общение духа, если [есть] какое милосердие и сострадательность,
PHIL|2|2|то дополните мою радость: имейте одни мысли, имейте ту же любовь, будьте единодушны и единомысленны;
PHIL|2|3|ничего [не делайте] по любопрению или по тщеславию, но по смиренномудрию почитайте один другого высшим себя.
PHIL|2|4|Не о себе [только] каждый заботься, но каждый и о других.
PHIL|2|5|Ибо в вас должны быть те же чувствования, какие и во Христе Иисусе:
PHIL|2|6|Он, будучи образом Божиим, не почитал хищением быть равным Богу;
PHIL|2|7|но уничижил Себя Самого, приняв образ раба, сделавшись подобным человекам и по виду став как человек;
PHIL|2|8|смирил Себя, быв послушным даже до смерти, и смерти крестной.
PHIL|2|9|Посему и Бог превознес Его и дал Ему имя выше всякого имени,
PHIL|2|10|дабы пред именем Иисуса преклонилось всякое колено небесных, земных и преисподних,
PHIL|2|11|и всякий язык исповедал, что Господь Иисус Христос в славу Бога Отца.
PHIL|2|12|Итак, возлюбленные мои, как вы всегда были послушны, не только в присутствии моем, но гораздо более ныне во время отсутствия моего, со страхом и трепетом совершайте свое спасение,
PHIL|2|13|потому что Бог производит в вас и хотение и действие по [Своему] благоволению.
PHIL|2|14|Все делайте без ропота и сомнения,
PHIL|2|15|чтобы вам быть неукоризненными и чистыми, чадами Божиими непорочными среди строптивого и развращенного рода, в котором вы сияете, как светила в мире,
PHIL|2|16|содержа слово жизни, к похвале моей в день Христов, что я не тщетно подвизался и не тщетно трудился.
PHIL|2|17|Но если я и соделываюсь жертвою за жертву и служение веры вашей, то радуюсь и сорадуюсь всем вам.
PHIL|2|18|О сем самом и вы радуйтесь и сорадуйтесь мне.
PHIL|2|19|Надеюсь же в Господе Иисусе вскоре послать к вам Тимофея, дабы и я, узнав о ваших обстоятельствах, утешился духом.
PHIL|2|20|Ибо я не имею никого равно усердного, кто бы столь искренно заботился о вас,
PHIL|2|21|потому что все ищут своего, а не того, что [угодно] Иисусу Христу.
PHIL|2|22|А его верность вам известна, потому что он, как сын отцу, служил мне в благовествовании.
PHIL|2|23|Итак я надеюсь послать его тотчас же, как скоро узнаю, что будет со мною.
PHIL|2|24|Я уверен в Господе, что и сам скоро приду к вам.
PHIL|2|25|Впрочем я почел нужным послать к вам Епафродита, брата и сотрудника и сподвижника моего, а вашего посланника и служителя в нужде моей,
PHIL|2|26|потому что он сильно желал видеть всех вас и тяжко скорбел о том, что до вас дошел слух о его болезни.
PHIL|2|27|Ибо он был болен при смерти; но Бог помиловал его, и не его только, но и меня, чтобы не прибавилась мне печаль к печали.
PHIL|2|28|Посему я скорее послал его, чтобы вы, увидев его снова, возрадовались, и я был менее печален.
PHIL|2|29|Примите же его в Господе со всякою радостью, и таких имейте в уважении,
PHIL|2|30|ибо он за дело Христово был близок к смерти, подвергая опасности жизнь, дабы восполнить недостаток ваших услуг мне.
PHIL|3|1|Впрочем, братия мои, радуйтесь о Господе. Писать вам о том же для меня не тягостно, а для вас назидательно.
PHIL|3|2|Берегитесь псов, берегитесь злых делателей, берегитесь обрезания,
PHIL|3|3|потому что обрезание – мы, служащие Богу духом и хвалящиеся Христом Иисусом, и не на плоть надеющиеся,
PHIL|3|4|хотя я могу надеяться и на плоть. Если кто другой думает надеяться на плоть, то более я,
PHIL|3|5|обрезанный в восьмой день, из рода Израилева, колена Вениаминова, Еврей от Евреев, по учению фарисей,
PHIL|3|6|по ревности – гонитель Церкви Божией, по правде законной – непорочный.
PHIL|3|7|Но что для меня было преимуществом, то ради Христа я почел тщетою.
PHIL|3|8|Да и все почитаю тщетою ради превосходства познания Христа Иисуса, Господа моего: для Него я от всего отказался, и все почитаю за сор, чтобы приобрести Христа
PHIL|3|9|и найтись в Нем не со своею праведностью, которая от закона, но с тою, которая через веру во Христа, с праведностью от Бога по вере;
PHIL|3|10|чтобы познать Его, и силу воскресения Его, и участие в страданиях Его, сообразуясь смерти Его,
PHIL|3|11|чтобы достигнуть воскресения мертвых.
PHIL|3|12|[Говорю так] не потому, чтобы я уже достиг, или усовершился; но стремлюсь, не достигну ли я, как достиг меня Христос Иисус.
PHIL|3|13|Братия, я не почитаю себя достигшим; а только, забывая заднее и простираясь вперед,
PHIL|3|14|стремлюсь к цели, к почести вышнего звания Божия во Христе Иисусе.
PHIL|3|15|Итак, кто из нас совершен, так должен мыслить; если же вы о чем иначе мыслите, то и это Бог вам откроет.
PHIL|3|16|Впрочем, до чего мы достигли, так и должны мыслить и по тому правилу жить.
PHIL|3|17|Подражайте, братия, мне и смотрите на тех, которые поступают по образу, какой имеете в нас.
PHIL|3|18|Ибо многие, о которых я часто говорил вам, а теперь даже со слезами говорю, поступают как враги креста Христова.
PHIL|3|19|Их конец – погибель, их бог – чрево, и слава их – в сраме, они мыслят о земном.
PHIL|3|20|Наше же жительство – на небесах, откуда мы ожидаем и Спасителя, Господа нашего Иисуса Христа,
PHIL|3|21|Который уничиженное тело наше преобразит так, что оно будет сообразно славному телу Его, силою, [которою] Он действует и покоряет Себе все.
PHIL|4|1|Итак, братия мои возлюбленные и вожделенные, радость и венец мой, стойте так в Господе, возлюбленные.
PHIL|4|2|Умоляю Еводию, умоляю Синтихию мыслить то же о Господе.
PHIL|4|3|Ей, прошу и тебя, искренний сотрудник, помогай им, подвизавшимся в благовествовании вместе со мною и с Климентом и с прочими сотрудниками моими, которых имена – в книге жизни.
PHIL|4|4|Радуйтесь всегда в Господе; и еще говорю: радуйтесь.
PHIL|4|5|Кротость ваша да будет известна всем человекам. Господь близко.
PHIL|4|6|Не заботьтесь ни о чем, но всегда в молитве и прошении с благодарением открывайте свои желания пред Богом,
PHIL|4|7|и мир Божий, который превыше всякого ума, соблюдет сердца ваши и помышления ваши во Христе Иисусе.
PHIL|4|8|Наконец, братия мои, что только истинно, что честно, что справедливо, что чисто, что любезно, что достославно, что только добродетель и похвала, о том помышляйте.
PHIL|4|9|Чему вы научились, что приняли и слышали и видели во мне, то исполняйте, – и Бог мира будет с вами.
PHIL|4|10|Я весьма возрадовался в Господе, что вы уже вновь начали заботиться о мне; вы и прежде заботились, но вам не благоприятствовали обстоятельства.
PHIL|4|11|Говорю это не потому, что нуждаюсь, ибо я научился быть довольным тем, что у меня есть.
PHIL|4|12|Умею жить и в скудости, умею жить и в изобилии; научился всему и во всем, насыщаться и терпеть голод, быть и в обилии и в недостатке.
PHIL|4|13|Все могу в укрепляющем меня Иисусе Христе.
PHIL|4|14|Впрочем вы хорошо поступили, приняв участие в моей скорби.
PHIL|4|15|Вы знаете, Филиппийцы, что в начале благовествования, когда я вышел из Македонии, ни одна церковь не оказала мне участия подаянием и принятием, кроме вас одних;
PHIL|4|16|вы и в Фессалонику и раз и два присылали мне на нужду.
PHIL|4|17|[Говорю это] не потому, чтобы я искал даяния; но ищу плода, умножающегося в пользу вашу.
PHIL|4|18|Я получил все, и избыточествую; я доволен, получив от Епафродита посланное вами, [как] благовонное курение, жертву приятную, благоугодную Богу.
PHIL|4|19|Бог мой да восполнит всякую нужду вашу, по богатству Своему в славе, Христом Иисусом.
PHIL|4|20|Богу же и Отцу нашему слава во веки веков! Аминь.
PHIL|4|21|Приветствуйте всякого святого во Христе Иисусе. Приветствуют вас находящиеся со мною братия.
PHIL|4|22|Приветствуют вас все святые, а наипаче из кесарева дома.
PHIL|4|23|Благодать Господа нашего Иисуса Христа со всеми вами. Аминь.
