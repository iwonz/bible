REV|1|1|Apocalypsis Iesu Christi, quam dedit illi Deus palam facere ser vis suis, quae oportet fieri cito, et significavit mittens per angelum suum servo suo Ioanni,
REV|1|2|qui testificatus est verbum Dei et testimonium Iesu Christi, quaecumque vidit.
REV|1|3|Beatus, qui legit et qui audiunt verba prophetiae et servant ea, quae in ea scripta sunt; tempus enim prope est.
REV|1|4|Ioannes septem ecclesiis, quae sunt in Asia: Gratia vobis et pax ab eo, qui est et qui erat et qui venturus est, et a septem spiritibus, qui in conspectu throni eius sunt,
REV|1|5|et ab Iesu Christo, qui est testis fidelis, primogenitus mortuorum et princeps regum terrae.Ei, qui diligit nos et solvit nos a peccatis nostris in sanguine suo
REV|1|6|et fecit nos regnum, sacerdotes Deo et Patri suo, ipsi gloria et imperium in saecula saeculorum. Amen.
REV|1|7|Ecce venit cum nubibus, et videbit eum omnis oculus et qui eum pupugerunt, et plangent se super eum omnes tribus terrae. Etiam, amen.
REV|1|8|Ego sum Alpha et Omega, dicit Dominus Deus, qui est et qui erat et qui venturus est, Omnipotens.
REV|1|9|Ego Ioannes, frater vester et particeps in tribulatione et regno et patientia in Iesu, fui in insula, quae appellatur Patmos, propter verbum Dei et testimonium Iesu.
REV|1|10|Fui in spiritu in dominica die et audivi post me vocem magnam tamquam tubae
REV|1|11|dicentis: " Quod vides, scribe in libro et mitte septem ecclesiis: Ephesum et Smyrnam et Pergamum et Thyatiram et Sardis et Philadelphiam et Laodiciam ".
REV|1|12|Et conversus sum, ut viderem vocem, quae loquebatur mecum; et conversus vidi septem candelabra aurea
REV|1|13|et in medio candelabrorum quasi Filium hominis, vestitum podere et praecinctum ad mamillas zonam auream;
REV|1|14|caput autem eius et capilli erant candidi tamquam lana alba, tamquam nix, et oculi eius velut flamma ignis,
REV|1|15|et pedes eius similes orichalco sicut in camino ardenti, et vox illius tamquam vox aquarum multarum,
REV|1|16|et habebat in dextera manu sua stellas septem, et de ore eius gladius anceps acutus exibat, et facies eius sicut sol lucet in virtute sua.
REV|1|17|Et cum vidissem eum, cecidi ad pedes eius tamquam mortuus; et posuit dexteram suam super me dicens: " Noli timere! Ego sum primus et novissimus,
REV|1|18|et vivens et fui mortuus et ecce sum vivens in saecula saeculorum et habeo claves mortis et inferni.
REV|1|19|Scribe ergo, quae vidisti et quae sunt et quae oportet fieri post haec.
REV|1|20|Mysterium septem stellarum, quas vidisti ad dexteram meam, et septem candelabra aurea: septem stellae, angeli sunt septem ecclesiarum; et candelabra septem, septem ecclesiae sunt.
REV|2|1|Angelo ecclesiae, quae est Ephesi, scribe:Haec dicit, qui tenet septem stellas in dextera sua, qui ambulat in medio septem candelabrorum aureorum:
REV|2|2|Scio opera tua et laborem et patientiam tuam, et quia non potes sustinere malos et tentasti eos, qui se dicunt apostolos et non sunt, et invenisti eos mendaces;
REV|2|3|et patientiam habes et sustinuisti propter nomen meum et non defecisti.
REV|2|4|Sed habeo adversus te quod caritatem tuam primam reliquisti.
REV|2|5|Memor esto itaque unde excideris, et age paenitentiam et prima opera fac; sin autem, venio tibi et movebo candelabrum tuum de loco suo, nisi paenitentiam egeris.
REV|2|6|Sed hoc habes, quia odisti facta Nicolaitarum, quae et ego odi.
REV|2|7|Qui habet aurem, audiat quid Spiritus dicat ecclesiis. Vincenti dabo ei edere de ligno vitae, quod est in paradiso Dei.
REV|2|8|Et angelo ecclesiae, quae est Smyrnae, scribe:Haec dicit Primus et Novissimus, qui fuit mortuus et vixit:
REV|2|9|Scio tribulationem tuam et paupertatem tuam - sed dives es - et blasphemiam ab his, qui se dicunt Iudaeos esse et non sunt, sed sunt synagoga Satanae.
REV|2|10|Nihil horum timeas, quae passurus es. Ecce missurus est Diabolus ex vobis in carcerem, ut tentemini, et habebitis tribulationem diebus decem. Esto fidelis usque ad mortem, et dabo tibi coronam vitae.
REV|2|11|Qui habet aurem, audiat quid Spiritus dicat ecclesiis. Qui vicerit, non laedetur a morte secunda.
REV|2|12|Et angelo ecclesiae, quae est Pergami, scribe:Haec dicit, qui habet romphaeam ancipitem acutam:
REV|2|13|Scio, ubi habitas, ubi thronus est Satanae, et tenes nomen meum et non negasti fidem meam et in diebus Antipas, testis meus fidelis, qui occisus est apud vos, ubi Satanas habitat.
REV|2|14|Sed habeo adversus te pauca, quia habes illic tenentes doctrinam Balaam, qui docebat Balac mittere scandalum coram filiis Israel, edere idolothyta et fornicari;
REV|2|15|ita habes et tu tenentes doctrinam Nicolaitarum similiter.
REV|2|16|Ergo paenitentiam age; si quo minus, venio tibi cito et pugnabo cum illis in gladio oris mei.
REV|2|17|Qui habet aurem, audiat quid Spiritus dicat ecclesiis. Vincenti dabo ei de manna abscondito et dabo illi calculum candidum, et in calculo nomen novum scriptum, quod nemo scit, nisi qui accipit.
REV|2|18|Et angelo ecclesiae, quae est Thyatirae, scribe: Haec dicit Filius Dei, qui habet oculos ut flammam ignis, et pedes eius similes orichalco:
REV|2|19|Novi opera tua et caritatem et fidem et ministerium et patientiam tuam et opera tua novissima plura prioribus.
REV|2|20|Sed habeo adversus te, quia permittis mulierem Iezabel, quae se dicit prophetissam, et docet et seducit servos meos fornicari et manducare idolothyta.
REV|2|21|Et dedi illi tempus, ut paenitentiam ageret, et non vult paeniteri a fornicatione sua.
REV|2|22|Ecce mitto eam in lectum et, qui moechantur cum ea, in tribulationem magnam, nisi paenitentiam egerint ab operibus eius.
REV|2|23|Et filios eius interficiam in morte, et scient omnes ecclesiae quia ego sum scrutans renes et corda, et dabo unicuique vestrum secundum opera vestra.
REV|2|24|Vobis autem dico ceteris, qui Thyatirae estis, quicumque non habent doctrinam hanc, qui non cognoverunt altitudines Satanae, quemadmodum dicunt, non mittam super vos aliud pondus;
REV|2|25|tamen id quod habetis, tenete, donec veniam.
REV|2|26|Et, qui vicerit et qui custodierit usque in finem opera mea, dabo illi potestatem super gentes,
REV|2|27|et reget illas in virga ferrea,tamquam vasa fictilia confringentur,
REV|2|28|sicut et ego accepi a Patre meo, et dabo illi stellam matutinam.
REV|2|29|Qui habet aurem, audiat quid Spiritus dicat ecclesiis.
REV|3|1|Et angelo ecclesiae, quae est Sardis, scribe:Haec dicit, qui habet septem spiritus Dei et septem stellas: Scio opera tua, quia nomen habes quod vivas, et mortuus es.
REV|3|2|Esto vigilans et confirma cetera, quae moritura erant, non enim invenio opera tua plena coram Deo meo;
REV|3|3|in mente ergo habe qualiter acceperis et audieris, et serva et paenitentiam age. Si ergo non vigilaveris, veniam tamquam fur, et nescies qua hora veniam ad te.
REV|3|4|Sed habes pauca nomina in Sardis, qui non inquinaverunt vestimenta sua et ambulabunt mecum in albis, quia digni sunt.
REV|3|5|Qui vicerit, sic vestietur vestimentis albis, et non delebo nomen eius de libro vitae et confitebor nomen eius coram Patre meo et coram angelis eius.
REV|3|6|Qui habet aurem, audiat quid Spiritus dicat ecclesiis.
REV|3|7|Et angelo ecclesiae, quae est Philadelphiae, scribe:Haec dicit Sanctus, Verus, qui habet clavem David, qui aperit, et nemo claudet; et claudit, et nemo aperit:
REV|3|8|Scio opera tua - ecce dedi coram te ostium apertum, quod nemo potest claudere - quia modicam habes virtutem, et servasti verbum meum et non negasti nomen meum.
REV|3|9|Ecce dabo de synagoga Satanae, qui dicunt se Iudaeos esse et non sunt, sed mentiuntur; ecce faciam illos, ut veniant et adorent ante pedes tuos et scient quia ego dilexi te.
REV|3|10|Quoniam servasti verbum patientiae meae, et ego te servabo ab hora tentationis, quae ventura est super orbem universum tentare habitantes in terra.
REV|3|11|Venio cito; tene quod habes, ut nemo accipiat coronam tuam.
REV|3|12|Qui vicerit, faciam illum columnam in templo Dei mei, et foras non egredietur amplius; et scribam super eum nomen Dei mei et nomen civitatis Dei mei, novae Ierusalem, quae descendit de caelo a Deo meo, et nomen meum novum.
REV|3|13|Qui habet aurem, audiat quid Spiritus dicat ecclesiis.
REV|3|14|Et angelo ecclesiae, quae est Laodiciae, scribe:Haec dicit Amen, testis fidelis et verus, principium creaturae Dei:
REV|3|15|Scio opera tua, quia neque frigidus es neque calidus. Utinam frigidus esses aut calidus!
REV|3|16|Sic quia tepidus es et nec calidus nec frigidus, incipiam te evomere ex ore meo.
REV|3|17|Quia dicis: "Dives sum et locupletatus et nullius egeo", et nescis quia tu es miser et miserabilis et pauper et caecus et nudus,
REV|3|18|suadeo tibi emere a me aurum igne probatum, ut locuples fias et vestimentis albis induaris, et non appareat confusio nuditatis tuae, et collyrium ad inunguendum oculos tuos, ut videas.
REV|3|19|Ego, quos amo, arguo et castigo. Aemulare ergo et paenitentiam age.
REV|3|20|Ecce sto ad ostium et pulso. Si quis audierit vocem meam et aperuerit ianuam, introibo ad illum et cenabo cum illo, et ipse mecum.
REV|3|21|Qui vicerit, dabo ei sedere mecum in throno meo, sicut et ego vici et sedi cum Patre meo in throno eius.
REV|3|22|Qui habet aurem, audiat quid Spiritus dicat ecclesiis ".
REV|4|1|Post haec vidi: et ecce ostium apertum in caelo, et vox prima, quam audivi, tamquam tubae loquentis mecum dicens: " Ascende huc, et ostendam tibi, quae oportet fieri post haec ".
REV|4|2|Statim fui in spiritu: et ecce thronus positus erat in caelo; et supra thronum sedens;
REV|4|3|et, qui sedebat, similis erat aspectu lapidi iaspidi et sardino; et iris erat in circuitu throni, aspectu similis smaragdo.
REV|4|4|Et in circuitu throni, viginti quattuor thronos, et super thronos viginti quattuor seniores sedentes, circumamictos vestimentis albis, et super capita eorum coronas aureas.
REV|4|5|Et de throno procedunt fulgura et voces et tonitrua; et septem lampades ignis ardentes ante thronum, quae sunt septem spiritus Dei;
REV|4|6|et in conspectu throni tamquam mare vitreum simile crystallo. Et in medio throni et in circuitu throni quattuor animalia, plena oculis ante et retro:
REV|4|7|et animal primum simile leoni, et secundum animal simile vitulo, et tertium animal habens faciem quasi hominis, et quartum animal simile aquilae volanti.
REV|4|8|Et quattuor animalia singula eorum habebant alas senas, in circuitu et intus plenae sunt oculis; et requiem non habent die et nocte dicentia: " Sanctus, sanctus, sanctus Dominus, Deus omnipotens, qui erat et qui est et qui venturus est! ".
REV|4|9|Et cum darent illa animalia gloriam et honorem et gratiarum actionem sedenti super thronum, viventi in saecula saeculorum,
REV|4|10|procidebant viginti quattuor seniores ante sedentem in throno et adorabant viventem in saecula saeculorum et mittebant coronas suas ante thronum dicentes:
REV|4|11|" Dignus es, Domine et Deus noster,accipere gloriam et honorem et virtutem,quia tu creasti omnia,et propter voluntatem tuam erant et creata sunt ".
REV|5|1|Et vidi in dextera sedentis super thronum librum scriptum intus et foris, signatum sigillis septem.
REV|5|2|Et vidi angelum fortem praedicantem voce magna: " Quis est dignus aperire librum et solvere signacula eius? ".
REV|5|3|Et nemo poterat in caelo neque in terra neque subtus terram aperire librum neque respicere illum.
REV|5|4|Et ego flebam multum, quoniam nemo dignus inventus est aperire librum nec respicere eum.
REV|5|5|Et unus de senioribus dicit mihi: " Ne fleveris; ecce vicit leo de tribu Iudae, radix David, aperire librum et septem signacula eius ".
REV|5|6|Et vidi in medio throni et quattuor animalium et in medio seniorum Agnum stantem tamquam occisum, habentem cornua septem et oculos septem, qui sunt septem spiritus Dei missi in omnem terram.
REV|5|7|Et venit et accepit de dextera sedentis in throno.
REV|5|8|Et cum accepisset librum, quattuor animalia et viginti quattuor seniores ceciderunt coram Agno, habentes singuli citharas et phialas aureas plenas incensorum, quae sunt orationes sanctorum.
REV|5|9|Et cantant novum canticum dicentes: Dignus es accipere librumet aperire signacula eius,quoniam occisus es et redemisti Deo in sanguine tuoex omni tribu et lingua et populo et natione;
REV|5|10|et fecisti eos Deo nostro regnum et sacerdotes,et regnabunt super terram ".
REV|5|11|Et vidi et audivi vocem angelorum multorum in circuitu throni et animalium et seniorum, et erat numerus eorum myriades myriadum et milia milium,
REV|5|12|dicentium voce magna: Dignus est Agnus, qui occisus est, accipere virtutem et divitias et sapientiamet fortitudinem et honorem et gloriam et benedictionem ".
REV|5|13|Et omnem creaturam, quae in caelo est et super terram et sub terra et super mare et quae in eis omnia, audivi dicentes: "Sedenti super thronum et Agno benedictio et honor et gloria et potestas in saecula saeculorum ".
REV|5|14|Et quattuor animalia dicebant: " Amen "; et seniores ceciderunt et adoraverunt.
REV|6|1|Et vidi, cum aperuisset Agnus unum de septem sigillis, et audi vi unum de quattuor animalibus dicens tamquam voce tonitrui: " Veni ".
REV|6|2|Et vidi: et ecce equus albus; et, qui sedebat super illum, habebat arcum, et data est ei corona, et exivit vincens et ut vinceret.
REV|6|3|Et cum aperuisset sigillum secundum, audivi secundum animal dicens: " Veni ".
REV|6|4|Et exivit alius equus rufus; et, qui sedebat super illum, datum est ei, ut sumeret pacem de terra, et ut invicem se interficiant; et datus est illi gladius magnus.
REV|6|5|Et cum aperuisset sigillum tertium, audivi tertium animal dicens: " Veni. Et vidi: et ecce equus niger; et, qui sedebat super eum, habebat stateram in manu sua.
REV|6|6|Et audivi tamquam vocem in medio quattuor animalium dicentem: " Bilibris tritici denario, et tres bilibres hordei denario; et oleum et vinum ne laeseris ".
REV|6|7|Et cum aperuisset sigillum quartum, audivi vocem quarti animalis dicentis: " Veni ".
REV|6|8|Et vidi: et ecce equus pallidus; et, qui sedebat desuper, nomen illi Mors, et Infernus sequebatur eum; et data est illis potestas super quartam partem terrae interficere gladio et fame et morte et a bestiis terrae.
REV|6|9|Et cum aperuisset quintum sigillum, vidi subtus altare animas interfectorum propter verbum Dei et propter testimonium, quod habebant.
REV|6|10|Et clamaverunt voce magna dicentes: " Usquequo, Domine, sanctus et verus, non iudicas et vindicas sanguinem nostrum de his, qui habitant in terra? ".
REV|6|11|Et datae sunt illis singulae stolae albae; et dictum est illis, ut requiescant tempus adhuc modicum, donec impleantur et conservi eorum et fratres eorum, qui interficiendi sunt sicut et illi.
REV|6|12|Et vidi, cum aperuisset sigillum sextum, et terraemotus factus est magnus, et sol factus est niger tamquam saccus cilicinus, et luna tota facta est sicut sanguis,
REV|6|13|et stellae caeli ceciderunt in terram, sicut ficus mittit grossos suos, cum vento magno movetur,
REV|6|14|et caelum recessit sicut liber involutus, et omnis mons et insula de locis suis motae sunt.
REV|6|15|Et reges terrae et magnates et tribuni et divites et fortes et omnis servus et liber absconderunt se in speluncis et in petris montium;
REV|6|16|et dicunt montibus et petris: " Cadite super nos et abscondite nos a facie sedentis super thronum et ab ira Agni,
REV|6|17|quoniam venit dies magnus irae ipsorum, et quis poterit stare? ".
REV|7|1|Post haec vidi quattuor angelos stantes super quattuor angulos terrae tenentes quattuor ventos terrae, ne flaret ventus super terram neque super mare neque in ullam arborem.
REV|7|2|Et vidi alterum angelum ascendentem ab ortu solis, habentem sigillum Dei vivi; et clamavit voce magna quattuor angelis, quibus datum est nocere terrae et mari,
REV|7|3|dicens: " Nolite nocere terrae neque mari neque arboribus, quoadusque signemus servos Dei nostri in frontibus eorum ".
REV|7|4|Et audivi numerum signatorum, centum quadraginta quattuor milia signati ex omni tribu filiorum Israel:
REV|7|5|ex tribu Iudae duodecim milia signati, ex tribu Ruben duodecim milia, ex tribu Gad duodecim milia,
REV|7|6|ex tribu Aser duodecim milia, ex tribu Nephthali duodecim milia, ex tribu Manasse duodecim milia,
REV|7|7|ex tribu Simeon duodecim milia, ex tribu Levi duodecim milia, ex tribu Issachar duodecim milia,
REV|7|8|ex tribu Zabulon duodecim milia, ex tribu Ioseph duodecim milia, ex tribu Beniamin duodecim milia signati.
REV|7|9|Post haec vidi: et ecce turba magna, quam dinumerare nemo poterat, ex omnibus gentibus et tribubus et populis et linguis stantes ante thronum et in conspectu Agni, amicti stolis albis, et palmae in manibus eorum;
REV|7|10|et clamant voce magna dicentes: " Salus Deo nostro, qui sedet super thronum, et Agno ".
REV|7|11|Et omnes angeli stabant in circuitu throni et seniorum et quattuor animalium, et ceciderunt in conspectu throni in facies suas et adoraverunt Deum
REV|7|12|dicentes: Amen! Benedictio et gloria et sapientia et gratiarum actio et honor et virtus et fortitudo Deo nostro in saecula saeculorum. Amen ".
REV|7|13|Et respondit unus de senioribus dicens mihi: " Hi, qui amicti sunt stolis albis, qui sunt et unde venerunt? ".
REV|7|14|Et dixi illi: " Domine mi, tu scis ". Et dixit mihi: " Hi sunt qui veniunt de tribulatione magna et laverunt stolas suas et dealbaverunt eas in sanguine Agni.
REV|7|15|Ideo sunt ante thronum Dei et serviunt ei die ac nocte in templo eius; et, qui sedet in throno, habitabit super illos.
REV|7|16|Non esurient amplius neque sitient amplius, neque cadet super illos sol neque ullus aestus,
REV|7|17|quoniam Agnus, qui in medio throni est, pascet illos et deducet eos ad vitae fontes aquarum, et absterget Deus omnem lacrimam ex oculis eorum ".
REV|8|1|Et cum aperuisset sigillum septimum, factum est silentium in caelo quasi media hora.
REV|8|2|Et vidi septem angelos, qui stant in conspectu Dei, et datae sunt illis septem tubae.
REV|8|3|Et alius angelus venit et stetit ante altare habens turibulum aureum, et data sunt illi incensa multa, ut daret orationibus sanctorum omnium super altare aureum, quod est ante thronum.
REV|8|4|Et ascendit fumus incensorum de orationibus sanctorum de manu angeli coram Deo.
REV|8|5|Et accepit angelus turibulum et implevit illud de igne altaris et misit in terram; et facta sunt tonitrua et voces et fulgura et terraemotus.
REV|8|6|Et septem angeli, qui habebant septem tubas, paraverunt se, ut tuba canerent.
REV|8|7|Et primus tuba cecinit. Et facta est grando et ignis mixta in sanguine, et missum est in terram: et tertia pars terrae combusta est, et tertia pars arborum combusta est, et omne fenum viride combustum est.
REV|8|8|Et secundus angelus tuba cecinit. Et tamquam mons magnus igne ardens missus est in mare: et facta est tertia pars maris sanguis,
REV|8|9|et mortua est tertia pars creaturarum, quae in mari sunt, quae habent animas, et tertia pars navium interiit.
REV|8|10|Et tertius angelus tuba cecinit. Et cecidit de caelo stella magna ardens tamquam facula et cecidit super tertiam partem fluminum et super fontes aquarum.
REV|8|11|Et nomen stellae dicitur Absinthius. Et facta est tertia pars aquarum in absinthium, et multi hominum mortui sunt de aquis, quia amarae factae sunt.
REV|8|12|Et quartus angelus tuba cecinit. Et percussa est tertia pars solis et tertia pars lunae et tertia pars stellarum, ut obscuraretur tertia pars eorum, et diei non luceret pars tertia, et nox similiter.
REV|8|13|Et vidi et audivi unam aquilam volantem per medium caelum dicentem voce magna: " Vae, vae, vae habitantibus in terra de ceteris vocibus tubae trium angelorum, qui tuba canituri sunt!".
REV|9|1|Et quintus angelus tuba cecinit. Et vidi stellam de caelo cecidis se in terram, et data est illi clavis putei abyssi.
REV|9|2|Et aperuit puteum abyssi, et ascendit fumus ex puteo sicut fumus fornacis magnae; et obscuratus est sol et aer de fumo putei.
REV|9|3|Et de fumo exierunt locustae in terram, et data est illis potestas, sicut habent potestatem scorpiones terrae.
REV|9|4|Et dictum est illis, ne laederent fenum terrae neque omne viride neque omnem arborem, nisi tantum homines, qui non habent signum Dei in frontibus.
REV|9|5|Et datum est illis, ne occiderent eos, sed ut cruciarentur mensibus quinque; et cruciatus eorum ut cruciatus scorpii, cum percutit hominem.
REV|9|6|Et in diebus illis quaerent homines mortem et non invenient eam; et desiderabunt mori, et fugit mors ab ipsis.
REV|9|7|Et similitudines locustarum similes equis paratis in proelium, et super capita earum tamquam coronae similes auro, et facies earum sicut facies hominum;
REV|9|8|et habebant capillos sicut capillos mulierum, et dentes earum sicut leonum erant,
REV|9|9|et habebant loricas sicut loricas ferreas, et vox alarum earum sicut vox curruum equorum multorum currentium in bellum.
REV|9|10|Et habent caudas similes scorpionibus et aculeos, et in caudis earum potestas earum nocere hominibus mensibus quinque.
REV|9|11|Habent super se regem angelum abyssi, cui nomen Hebraice Abaddon et Graece nomen habet Apollyon.
REV|9|12|Vae unum abiit. Ecce veniunt adhuc duo vae post haec.
REV|9|13|Et sextus angelus tuba cecinit. Et audivi vocem unam ex cornibus altaris aurei, quod est ante Deum,
REV|9|14|dicentem sexto angelo, qui habebat tubam: " Solve quattuor angelos, qui alligati sunt super flumen magnum Euphraten ".
REV|9|15|Et soluti sunt quattuor angeli, qui parati erant in horam et diem et mensem et annum, ut occiderent tertiam partem hominum.
REV|9|16|Et numerus equestris exercitus vicies milies dena milia; audivi numerum eorum.
REV|9|17|Et ita vidi equos in visione et, qui sedebant super eos, habentes loricas igneas et hyacinthinas et sulphureas; et capita equorum erant tamquam capita leonum, et de ore ipsorum procedit ignis et fumus et sulphur.
REV|9|18|Ab his tribus plagis occisa est tertia pars hominum, de igne et fumo et sulphure, quod procedebat ex ore ipsorum.
REV|9|19|Potestas enim equorum in ore eorum est et in caudis eorum; nam caudae illorum similes serpentibus habentes capita, et in his nocent.
REV|9|20|Et ceteri homines, qui non sunt occisi in his plagis neque paenitentiam egerunt de operibus manuum suarum, ut non adorarent daemonia et simulacra aurea et argentea et aerea et lapidea et lignea, quae neque videre possunt neque audire neque ambulare,
REV|9|21|et non egerunt paenitentiam ab homicidiis suis neque a veneficiis suis neque a fornicatione sua neque a furtis suis.
REV|10|1|Et vidi alium angelum for tem descendentem de caelo amictum nube, et iris super caput, et facies eius erat ut sol, et pedes eius tamquam columnae ignis;
REV|10|2|et habebat in manu sua libellum apertum. Et posuit pedem suum dexterum supra mare, sinistrum autem super terram,
REV|10|3|et clamavit voce magna, quemadmodum cum leo rugit. Et cum clamasset, locuta sunt septem tonitrua voces suas.
REV|10|4|Et cum locuta fuissent septem tonitrua, scripturus eram; et audivi vocem de caelo dicentem: " Signa, quae locuta sunt septem tonitrua, et noli ea scribere ".
REV|10|5|Et angelus, quem vidi stantem supra mare et supra terram, levavit manum suam dexteram ad caelum
REV|10|6|et iuravit per Viventem in saecula saeculorum, qui creavit caelum et ea, quae in illo sunt, et terram et ea, quae in ea sunt, et mare et ea, quae in eo sunt: " Tempus amplius non erit,
REV|10|7|sed in diebus vocis septimi angeli, cum coeperit tuba canere, et consummatum est mysterium Dei, sicut evangelizavit servis suis prophetis.
REV|10|8|Et vox, quam audivi de caelo, iterum loquentem mecum et dicentem: " Vade, accipe librum apertum de manu angeli stantis supra mare et supra terram ".
REV|10|9|Et abii ad angelum dicens ei, ut daret mihi libellum. Et dicit mihi: " Accipe et devora illum; et faciet amaricare ventrem tuum, sed in ore tuo erit dulcis tamquam mel ".
REV|10|10|Et accepi libellum de manu angeli et devoravi eum, et erat in ore meo tamquam mel dulcis; et cum devorassem eum, amaricatus est venter meus.
REV|10|11|Et dicunt mihi: " Oportet te iterum prophetare super populis et gentibus et linguis et regibus multis ".
REV|11|1|Et datus est mihi calamus similis virgae dicens: " Surge et metire templum Dei et altare et adorantes in eo.
REV|11|2|Atrium autem, quod est foris templum, eice foras et ne metiaris illud, quoniam datum est gentibus, et civitatem sanctam calcabunt mensibus quadraginta duobus.
REV|11|3|Et dabo duobus testibus meis, et prophetabunt diebus mille ducentis sexaginta amicti saccis ".
REV|11|4|Hi sunt duae olivae et duo candelabra in conspectu Domini terrae stantes.
REV|11|5|Et si quis eis vult nocere, ignis exit de ore illorum et devorat inimicos eorum; et si quis voluerit eos laedere, sic oportet eum occidi.
REV|11|6|Hi habent potestatem claudendi caelum, ne pluat pluvia diebus prophetiae ipsorum; et potestatem habent super aquas convertendi eas in sanguinem et percutere terram omni plaga, quotienscumque voluerint.
REV|11|7|Et cum finierint testimonium suum, bestia, quae ascendit de abysso, faciet adversus illos bellum et vincet eos et occidet illos.
REV|11|8|Et corpus eorum in platea civitatis magnae, quae vocatur spiritaliter Sodoma et Aegyptus, ubi et Dominus eorum crucifixus est;
REV|11|9|et vident de populis et tribubus et linguis et gentibus corpus eorum per tres dies et dimidium, et corpora eorum non sinunt poni in monumento.
REV|11|10|Et inhabitantes terram gaudent super illis et iucundantur et munera mittent invicem, quoniam hi duo prophetae cruciaverunt eos, qui inhabitant super terram.
REV|11|11|Et post dies tres et dimidium spiritus vitae a Deo intravit in eos, et steterunt super pedes suos; et timor magnus cecidit super eos, qui videbant eos.
REV|11|12|Et audierunt vocem magnam de caelo dicentem illis: " Ascendite huc "; et ascenderunt in caelum in nube, et viderunt illos inimici eorum.
REV|11|13|Et in illa hora factus est terraemotus magnus, et decima pars civitatis cecidit, et occisi sunt in terraemotu nomina hominum septem milia, et reliqui in timorem sunt missi et dederunt gloriam Deo caeli.
REV|11|14|Vae secundum abiit; ecce vae tertium venit cito.
REV|11|15|Et septimus angelus tuba cecinit, et factae sunt voces magnae in caelo dicentes: " Factum est regnum huius mundi Domini nostri et Christi eius, et regnabit in saecula saeculorum ".
REV|11|16|Et viginti quattuor seniores, qui in conspectu Dei sedent in thronis suis, ceciderunt super facies suas et adoraverunt Deum
REV|11|17|dicentes: Gratias agimus tibi,Domine, Deus omnipotens,qui es et qui eras,quia accepisti virtutem tuam magnam et regnasti.
REV|11|18|Et iratae sunt gentes,et advenit ira tua, et tempus mortuorum iudicariet reddere mercedem servis tuis prophetis et sanctiset timentibus nomen tuum, pusillis et magnis,et exterminare eos, qui exterminant terram ".
REV|11|19|Et apertum est templum Dei in caelo, et visa est arca testamenti eius in templo eius; et facta sunt fulgura et voces et terraemotus et grando magna.
REV|12|1|Et signum magnum appa ruit in caelo: mulier amicta sole, et luna sub pedibus eius, et super caput eius corona stellarum duodecim;
REV|12|2|et in utero habens, et clamat parturiens et cruciatur, ut pariat.
REV|12|3|Et visum est aliud signum in caelo: et ecce draco rufus magnus, habens capita septem et cornua decem, et super capita sua septem diademata;
REV|12|4|et cauda eius trahit tertiam partem stellarum caeli et misit eas in terram. Et draco stetit ante mulierem, quae erat paritura, ut, cum peperisset, filium eius devoraret.
REV|12|5|Et peperit filium, masculum, qui recturus est omnes gentes in virga ferrea; et raptus est filius eius ad Deum et ad thronum eius.
REV|12|6|Et mulier fugit in desertum, ubi habet locum paratum a Deo, ut ibi pascant illam diebus mille ducentis sexaginta.
REV|12|7|Et factum est proelium in caelo, Michael et angeli eius, ut proeliarentur cum dracone. Et draco pugnavit et angeli eius,
REV|12|8|et non valuit, neque locus inventus est eorum amplius in caelo.
REV|12|9|Et proiectus est draco ille magnus, serpens antiquus, qui vocatur Diabolus et Satanas, qui seducit universum orbem; proiectus est in terram, et angeli eius cum illo proiecti sunt.
REV|12|10|Et audivi vocem magnam in caelo dicentem: Nunc facta est salus et virtus et regnum Dei nostriet potestas Christi eius,quia proiectus est accusator fratrum nostrorum,qui accusabat illos ante conspectum Dei nostri die ac nocte.
REV|12|11|Et ipsi vicerunt illum propter sanguinem Agniet propter verbum testimonii sui;et non dilexerunt animam suamusque ad mortem.
REV|12|12|Propterea laetamini, caeliet qui habitatis in eis.Vae terrae et mari, quia descendit Diabolus ad vos habens iram magnam, sciens quod modicum tempus habet! ".
REV|12|13|Et postquam vidit draco quod proiectus est in terram, persecutus est mulierem, quae peperit masculum.
REV|12|14|Et datae sunt mulieri duae alae aquilae magnae, ut volaret in desertum in locum suum, ubi alitur per tempus et tempora et dimidium temporis a facie serpentis.
REV|12|15|Et misit serpens ex ore suo post mulierem aquam tamquam flumen, ut eam faceret trahi a flumine.
REV|12|16|Et adiuvit terra mulierem, et aperuit terra os suum et absorbuit flumen, quod misit draco de ore suo.
REV|12|17|Et iratus est draco in mulierem et abiit facere proelium cum reliquis de semine eius, qui custodiunt mandata Dei et habent testimonium Iesu.
REV|12|18|Et stetit super arenam maris.
REV|13|1|Et vidi de mari bestiam ascendentem, habentem cor nua decem et capita septem, et super cornua eius decem diademata, et super capita eius nomina blasphemiae.
REV|13|2|Et bestia, quam vidi, similis erat pardo, et pedes eius sicut ursi, et os eius sicut os leonis. Et dedit illi draco virtutem suam et thronum suum et potestatem magnam.
REV|13|3|Et unum de capitibus suis quasi occisum in mortem, et plaga mortis eius curata est.Et admirata est universa terra post bestiam,
REV|13|4|et adoraverunt draconem, quia dedit potestatem bestiae, et adoraverunt bestiam dicentes: " Quis similis bestiae, et quis potest pugnare cum ea?.
REV|13|5|Et datum est ei os loquens magna et blasphemias, et data est illi potestas facere menses quadraginta duos.
REV|13|6|Et aperuit os suum in blasphemias ad Deum, blasphemare nomen eius et tabernaculum eius, eos, qui in caelo habitant.
REV|13|7|Et datum est illi bellum facere cum sanctis et vincere illos, et data est ei potestas super omnem tribum et populum et linguam et gentem.
REV|13|8|Et adorabunt eum omnes, qui inhabitant terram, cuiuscumque non est scriptum nomen in libro vitae Agni, qui occisus est, ab origine mundi.
REV|13|9|Si quis habet aurem, audiat:
REV|13|10|Si quis in captivitatem,in captivitatem vadit;si quis in gladio debet occidi,oportet eum in gladio occidi.Hic est patientia et fides sanctorum.
REV|13|11|Et vidi aliam bestiam ascendentem de terra, et habebat cornua duo similia agni, et loquebatur sicut draco.
REV|13|12|Et potestatem prioris bestiae omnem facit in conspectu eius. Et facit terram et inhabitantes in ea adorare bestiam primam, cuius curata est plaga mortis.
REV|13|13|Et facit signa magna, ut etiam ignem faciat de caelo descendere in terram in conspectu hominum.
REV|13|14|Et seducit habitantes terram propter signa, quae data sunt illi facere in conspectu bestiae, dicens habitantibus in terra, ut faciant imaginem bestiae, quae habet plagam gladii et vixit.
REV|13|15|Et datum est illi, ut daret spiritum imagini bestiae, ut et loquatur imago bestiae; et faciat, ut quicumque non adoraverint imaginem bestiae, occidantur.
REV|13|16|Et facit omnes pusillos et magnos et divites et pauperes et liberos et servos accipere characterem in dextera manu sua aut in frontibus suis,
REV|13|17|et ne quis possit emere aut vendere, nisi qui habet characterem, nomen bestiae aut numerum nominis eius.
REV|13|18|Hic sapientia est: qui habet intellectum, computet numerum bestiae; numerus enim hominis est: et numerus eius est sescenti sexaginta sex.
REV|14|1|Et vidi: et ecce Agnus stans supra montem Sion, et cum illo centum quadraginta quattuor milia, habentes nomen eius et nomen Patris eius scriptum in frontibus suis.
REV|14|2|Et audivi vocem de caelo tamquam vocem aquarum multarum et tamquam vocem tonitrui magni; et vox, quam audivi, sicut citharoedorum citharizantium in citharis suis.
REV|14|3|Et cantant quasi canticum novum ante thronum et ante quattuor animalia et seniores. Et nemo poterat discere canticum, nisi illa centum quadraginta quattuor milia, qui empti sunt de terra.
REV|14|4|Hi sunt qui cum mulieribus non sunt coinquinati, virgines enim sunt. Hi qui sequuntur Agnum, quocumque abierit. Hi empti sunt ex hominibus primitiae Deo et Agno;
REV|14|5|et in ore ipsorum non est inventum mendacium: sine macula sunt.
REV|14|6|Et vidi alterum angelum volantem per medium caelum, habentem evangelium aeternum, ut evangelizaret super sedentes in terra et super omnem gentem et tribum et linguam et populum;
REV|14|7|dicens magna voce: " Timete Deum et date illi gloriam, quia venit hora iudicii eius; et adorate eum, qui fecit caelum et terram et mare et fontes aquarum ".
REV|14|8|Et alius angelus secutus est dicens: " Cecidit, cecidit Babylon illa magna, quae a vino irae fornicationis suae potionavit omnes gentes! ".
REV|14|9|Et alius angelus tertius secutus est illos dicens voce magna: " Si quis adoraverit bestiam et imaginem eius et acceperit characterem in fronte sua aut in manu sua,
REV|14|10|et hic bibet de vino irae Dei, quod mixtum est mero in calice irae ipsius, et cruciabitur igne et sulphure in conspectu angelorum sanctorum et ante conspectum Agni.
REV|14|11|Et fumus tormentorum eorum in saecula saeculorum ascendit, nec habent requiem die ac nocte, qui adoraverunt bestiam et imaginem eius, et si quis acceperit characterem nominis eius ".
REV|14|12|Hic patientia sanctorum est, qui custodiunt mandata Dei et fidem Iesu.
REV|14|13|Et audivi vocem de caelo dicentem: " Scribe: Beati mortui, qui in Domino moriuntur amodo. Etiam, dicit Spiritus, ut requiescant a laboribus suis; opera enim illorum sequuntur illos ".
REV|14|14|Et vidi: et ecce nubem candidam, et supra nubem sedentem quasi Filium hominis, habentem super caput suum coronam auream et in manu sua falcem acutam.
REV|14|15|Et alter angelus exivit de templo clamans voce magna ad sedentem super nubem: " Mitte falcem tuam et mete, quia venit hora, ut metatur, quoniam aruit messis terrae ".
REV|14|16|Et misit, qui sedebat supra nubem, falcem suam in terram, et messa est terra.
REV|14|17|Et alius angelus exivit de templo, quod est in caelo, habens et ipse falcem acutam.
REV|14|18|Et alius angelus de altari, habens potestatem supra ignem, et clamavit voce magna ad eum, qui habebat falcem acutam, dicens: " Mitte falcem tuam acutam et vindemia botros vineae terrae, quoniam maturae sunt uvae eius ".
REV|14|19|Et misit angelus falcem suam in terram et vindemiavit vineam terrae et misit in lacum irae Dei magnum.
REV|14|20|Et calcatus est lacus extra civitatem, et exivit sanguis de lacu usque ad frenos equorum per stadia mille sescenta.
REV|15|1|Et vidi aliud signum in caelo magnum et mirabile: angelos septem habentes plagas septem novissimas, quoniam in illis consummata est ira Dei.
REV|15|2|Et vidi tamquam mare vitreum mixtum igne; et eos, qui vicerunt bestiam et imaginem illius et numerum nominis eius, stantes supra mare vitreum, habentes citharas Dei.
REV|15|3|Et cantant canticum Moysis servi Dei et canticum Agni dicentes: Magna et mirabilia opera tua,Domine, Deus omnipotens;iustae et verae viae tuae,Rex gentium!
REV|15|4|Quis non timebit, Domine,et glorificabit nomen tuum?Quia solus Sanctus,quoniam omnes gentes venientet adorabunt in conspectu tuo,quoniam iudicia tua manifestata sunt ".
REV|15|5|Et post haec vidi: et apertum est templum tabernaculi testimonii in caelo,
REV|15|6|et exierunt septem angeli habentes septem plagas de templo, vestiti lino mundo candido et praecincti circa pectora zonis aureis.
REV|15|7|Et unum ex quattuor animalibus dedit septem angelis septem phialas aureas plenas iracundiae Dei viventis in saecula saeculorum.
REV|15|8|Et impletum est templum fumo de gloria Dei et de virtute eius; et nemo poterat introire in templum, donec consummarentur septem plagae septem angelorum.
REV|16|1|Et audivi vocem magnam de templo dicentem septem an gelis: " Ite et effundite septem phialas irae Dei in terram ".
REV|16|2|Et abiit primus et effudit phialam suam in terram; et factum est vulnus saevum ac pessimum in homines, qui habebant characterem bestiae, et eos, qui adorabant imaginem eius.
REV|16|3|Et secundus effudit phialam suam in mare; et factus est sanguis tamquam mortui, et omnis anima vivens mortua est, quae est in mari.
REV|16|4|Et tertius effudit phialam suam in flumina et in fontes aquarum; et factus est sanguis.
REV|16|5|Et audivi angelum aquarum dicentem: " Iustus es, qui es et qui eras, Sanctus, quia haec iudicasti;
REV|16|6|quia sanguinem sanctorum et prophetarum fuderunt, et sanguinem eis dedisti bibere: digni sunt! ".
REV|16|7|Et audivi altare dicens: " Etiam, Domine, Deus omnipotens, vera et iusta iudicia tua! ".
REV|16|8|Et quartus effudit phialam suam in solem; et datum est illi aestu afficere homines in igne.
REV|16|9|Et aestuaverunt homines aestu magno; et blasphemaverunt nomen Dei habentis potestatem super has plagas et non egerunt paenitentiam, ut darent illi gloriam.
REV|16|10|Et quintus effudit phialam suam super thronum bestiae; et factum est regnum eius tenebrosum, et commanducaverunt linguas suas prae dolore
REV|16|11|et blasphemaverunt Deum caeli prae doloribus suis et vulneribus suis et non egerunt paenitentiam ex operibus suis.
REV|16|12|Et sextus effudit phialam suam super flumen illud magnum Euphraten; et exsiccata est aqua eius, ut praepararetur via regibus, qui sunt ab ortu solis.
REV|16|13|Et vidi de ore draconis et de ore bestiae et de ore pseudoprophetae spiritus tres immundos velut ranas;
REV|16|14|sunt enim spiritus daemoniorum facientes signa, qui procedunt ad reges universi orbis congregare illos in proelium diei magni Dei omnipotentis.
REV|16|15|Ecce venio sicut fur. Beatus, qui vigilat et custodit vestimenta sua, ne nudus ambulet, et videant turpitudinem eius.
REV|16|16|Et congregavit illos in locum, qui vocatur Hebraice Harmagedon.
REV|16|17|Et septimus effudit phialam suam in aerem; et exivit vox magna de templo a throno dicens: " Factum est! ".
REV|16|18|Et facta sunt fulgura et voces et tonitrua, et terraemotus factus est magnus, qualis numquam fuit, ex quo homo fuit super terram, talis terraemotus sic magnus.
REV|16|19|Et facta est civitas magna in tres partes, et civitates gentium ceciderunt. Et Babylon magna venit in memoriam ante Deum dare ei calicem vini indignationis irae eius.
REV|16|20|Et omnis insula fugit, et montes non sunt inventi.
REV|16|21|Et grando magna sicut talentum descendit de caelo in homines; et blasphemaverunt homines Deum propter plagam grandinis, quoniam magna est plaga eius nimis.
REV|17|1|Et venit unus de septem angelis, qui habebant septem phialas, et locutus est mecum dicens: " Veni, ostendam tibi damnationem meretricis magnae, quae sedet super aquas multas,
REV|17|2|cum qua fornicati sunt reges terrae, et inebriati sunt, qui inhabitant terram, de vino prostitutionis eius ".
REV|17|3|Et abstulit me in desertum in spiritu. Et vidi mulierem sedentem super bestiam coccineam, plenam nominibus blasphemiae, habentem capita septem et cornua decem.
REV|17|4|Et mulier erat circumdata purpura et coccino, et inaurata auro et lapide pretioso et margaritis, habens poculum aureum in manu sua plenum abominationibus et immunditiis fornicationis eius;
REV|17|5|et in fronte eius nomen scriptum, mysterium: " Babylon magna, mater fornicationum et abominationum terrae ".
REV|17|6|Et vidi mulierem ebriam de sanguine sanctorum et de sanguine martyrum Iesu. Et miratus sum, cum vidissem illam, admiratione magna.
REV|17|7|Et dixit mihi angelus. " Quare miraris? Ego tibi dicam mysterium mulieris et bestiae, quae portat eam, quae habet capita septem et decem cornua:
REV|17|8|bestia, quam vidisti, fuit et non est, et ascensura est de abysso et in interitum ibit. Et mirabuntur inhabitantes terram, quorum non sunt scripta nomina in libro vitae a constitutione mundi, videntes bestiam, quia erat et non est et aderit.
REV|17|9|Hic est sensus, qui habet sapientiam. Septem capita, septem montes sunt, super quos mulier sedet. Et reges septem sunt:
REV|17|10|quinque ceciderunt, unus est, alius nondum venit; et, cum venerit, oportet illum breve tempus manere.
REV|17|11|Et bestia, quae erat et non est, et is octavus est et de septem est et in interitum vadit.
REV|17|12|Et decem cornua, quae vidisti, decem reges sunt, qui regnum nondum acceperunt, sed potestatem tamquam reges una hora accipiunt cum bestia.
REV|17|13|Hi unum consilium habent et virtutem et potestatem suam bestiae tradunt.
REV|17|14|Hi cum Agno pugnabunt; et Agnus vincet illos, quoniam Dominus dominorum est et Rex regum, et qui cum illo sunt vocati et electi et fideles ".
REV|17|15|Et dicit mihi: " Aquae, quas vidisti, ubi meretrix sedet, populi et turbae sunt et gentes et linguae.
REV|17|16|Et decem cornua, quae vidisti, et bestia, hi odient fornicariam et desolatam facient illam et nudam, et carnes eius manducabunt et ipsam igne concremabunt;
REV|17|17|Deus enim dedit in corda eorum, ut faciant, quod illi placitum est, et faciant unum consilium et dent regnum suum bestiae, donec consummentur verba Dei.
REV|17|18|Et mulier, quam vidisti, est civitas magna, quae habet regnum super reges terrae ".
REV|18|1|Post haec vidi alium ange lum descendentem de caelo, habentem potestatem magnam; et terra illuminata est a claritate eius.
REV|18|2|Et clamavit in forti voce dicens: " Cecidit, cecidit Babylon magna et facta est habitatio daemoniorum et custodia omnis spiritus immundi et custodia omnis bestiae immundae et odibilis;
REV|18|3|quia de vino irae fornicationis eius biberunt omnes gentes, et reges terrae cum illa fornicati sunt, et mercatores terrae de virtute deliciarum eius divites facti sunt! ".
REV|18|4|Et audivi aliam vocem de caelo dicentem: " Exite de illa, populus meus, ut ne comparticipes sitis peccatorum eius et de plagis eius non accipiatis,
REV|18|5|quoniam pervenerunt peccata eius usque ad caelum, et recordatus est Deus iniquitatum eius.
REV|18|6|Reddite illi, sicut et ipsa reddidit, et duplicate duplicia secundum opera eius; in poculo, quo miscuit, miscete illi duplum.
REV|18|7|Quantum glorificavit se et in deliciis fuit, tantum date illi tormentum et luctum. Quia in corde suo dicit: "Sedeo regina et vidua non sum et luctum non videbo",
REV|18|8|ideo in una die venient plagae eius, mors et luctus et fames, et igne comburetur, quia fortis est Dominus Deus, qui iudicavit illam ".
REV|18|9|Et flebunt et plangent se super illam reges terrae, qui cum illa fornicati sunt et in deliciis vixerunt, cum viderint fumum incendii eius,
REV|18|10|longe stantes propter timorem tormentorum eius, dicentes: " Vae, vae, civitas illa magna, Babylon, civitas illa fortis, quoniam una hora venit iudicium tuum! ".
REV|18|11|Et negotiatores terrae flent et lugent super illam, quoniam mercem eorum nemo emit amplius:
REV|18|12|mercem auri et argenti et lapidis pretiosi et margaritarum, et byssi et purpurae et serici et cocci, et omne lignum thyinum et omnia vasa eboris et omnia vasa de ligno pretiosissimo et aeramento et ferro et marmore,
REV|18|13|et cinnamomum et amomum et odoramenta et unguenta et tus, et vinum et oleum et similam et triticum, et iumenta et oves et equorum et raedarum, et mancipiorum et animas hominum.
REV|18|14|Et fructus tui, desiderium animae, discesserunt a te, et omnia pinguia et clara perierunt a te, et amplius illa iam non invenient.
REV|18|15|Mercatores horum, qui divites facti sunt ab ea, longe stabunt propter timorem tormentorum eius flentes ac lugentes,
REV|18|16|dicentes: " Vae, vae, civitas illa magna, quae amicta erat byssino et purpura et cocco, et deaurata auro et lapide pretioso et margarita,
REV|18|17|quoniam una hora desolatae sunt tantae divitiae! ".Et omnis gubernator et omnis, qui in locum navigat, et nautae et, quotquot maria operantur, longe steterunt
REV|18|18|et clamabant, videntes fumum incendii eius, dicentes: " Quae similis civitati huic magnae? ".
REV|18|19|Et miserunt pulverem super capita sua et clamabant, flentes et lugentes, dicentes: " Vae, vae, civitas illa magna, in qua divites facti sunt omnes, qui habent naves in mari, de opibus eius, quoniam una hora desolata est!
REV|18|20|Exsulta super eam, caelum, et sancti et apostoli et prophetae, quoniam iudicavit Deus iudicium vestrum de illa! ".
REV|18|21|Et sustulit unus angelus fortis lapidem quasi molarem magnum et misit in mare dicens: "Impetu sic mittetur Babylon magna illa civitas et ultra iam non invenietur.
REV|18|22|Et vox citharoedorum et musicorum et tibia canentium et tuba non audietur in te amplius, et omnis artifex omnis artis non invenietur in te amplius, et vox molae non audietur in te amplius,
REV|18|23|et lux lucernae non lucebit tibi amplius, et vox sponsi et sponsae non audietur in te amplius; quia mercatores tui erant magnates terrae, quia in veneficiis tuis erraverunt omnes gentes,
REV|18|24|et in ea sanguis prophetarum et sanctorum inventus est et omnium, qui interfecti sunt in terra! ".
REV|19|1|Post haec audivi quasi vo cem magnam turbae multae in caelo dicentium: Alleluia!Salus et gloria et virtus Deo nostro,
REV|19|2|quia vera et iusta iudicia eius;quia iudicavit de meretrice magna, quae corrupit terram in prostitutione sua, et vindicavit sanguinem servorum suorum de manibus eius! ".
REV|19|3|Et iterum dixerunt: " Alleluia! Et fumus eius ascendit in saecula saeculorum! ".
REV|19|4|Et ceciderunt seniores viginti quattuor et quattuor animalia et adoraverunt Deum sedentem super thronum dicentes: " Amen. Alleluia ".
REV|19|5|Et vox de throno exivit dicens: Laudem dicite Deo nostro, omnes servi eiuset qui timetis eum, pusilli et magni! ".
REV|19|6|Et audivi quasi vocem turbae magnae et sicut vocem aquarum multarum et sicut vocem tonitruum magnorum dicentium: Alleluia,quoniam regnavit Dominus, Deus noster omnipotens.
REV|19|7|Gaudeamus et exsultemus et demus gloriam ei,quia venerunt nuptiae Agni,et uxor eius praeparavit se.
REV|19|8|Et datum est illi, ut cooperiat se byssino splendenti mundo: byssinum enim iustificationes sunt sanctorum ".
REV|19|9|Et dicit mihi: " Scribe: Beati, qui ad cenam nuptiarum Agni vocati sunt!. Et dicit mihi: " Haec verba Dei vera sunt ".
REV|19|10|Et cecidi ante pedes eius, ut adorarem eum. Et dicit mihi: " Vide, ne feceris! Conservus tuus sum et fratrum tuorum habentium testimonium Iesu. Deum adora. Testimonium enim Iesu est spiritus prophetiae ".
REV|19|11|Et vidi caelum apertum: et ecce equus albus; et, qui sedebat super eum, vocabatur Fidelis et Verax, et in iustitia iudicat et pugnat.
REV|19|12|Oculi autem eius sicut flamma ignis, et in capite eius diademata multa, habens nomen scriptum, quod nemo novit nisi ipse;
REV|19|13|et vestitus veste aspersa sanguine, et vocatur nomen eius Verbum Dei.
REV|19|14|Et exercitus, qui sunt in caelo, sequebantur eum in equis albis, vestiti byssino albo mundo.
REV|19|15|Et de ore ipsius procedit gladius acutus, ut in ipso percutiat gentes, et ipse reget eos in virga ferrea; et ipse calcat torcular vini furoris irae Dei omnipotentis.
REV|19|16|Et habet super vestimentum et super femur suum nomen scriptum: Rex regum et Dominus dominorum.
REV|19|17|Et vidi unum angelum stantem in sole, et clamavit voce magna dicens omnibus avibus, quae volabant per medium caeli: "Venite, congregamini ad cenam magnam Dei,
REV|19|18|ut manducetis carnes regum et carnes tribunorum et carnes fortium et carnes equorum et sedentium in ipsis et carnes omnium liberorum ac servorum et pusillorum ac magnorum ".
REV|19|19|Et vidi bestiam et reges terrae et exercitus eorum congregatos ad faciendum proelium cum illo, qui sedebat super equum, et cum exercitu eius.
REV|19|20|Et apprehensa est bestia et cum illa pseudopropheta, qui fecit signa coram ipsa, quibus seduxit eos, qui acceperunt characterem bestiae et qui adorant imaginem eius; vivi missi sunt hi duo in stagnum ignis ardentis sulphure.
REV|19|21|Et ceteri occisi sunt in gladio sedentis super equum, qui procedit de ore ipsius, et omnes aves saturatae sunt carnibus eorum.
REV|20|1|Et vidi angelum descen dentem de caelo habentem clavem abyssi et catenam magnam in manu sua.
REV|20|2|Et apprehendit draconem, serpentem antiquum, qui est Diabolus et Satanas, et ligavit eum per annos mille;
REV|20|3|et misit eum in abyssum et clausit et signavit super illum, ut non seducat amplius gentes, donec consummentur mille anni; post haec oportet illum solvi modico tempore.
REV|20|4|Et vidi thronos, et sederunt super eos, et iudicium datum est illis; et animas decollatorum propter testimonium Iesu et propter verbum Dei, et qui non adoraverunt bestiam neque imaginem eius nec acceperunt characterem in frontibus et in manibus suis; et vixerunt et regnaverunt cum Christo mille annis.
REV|20|5|Ceteri mortuorum non vixerunt, donec consummentur mille anni. Haec est resurrectio prima.
REV|20|6|Beatus et sanctus, qui habet partem in resurrectione prima! In his secunda mors non habet potestatem, sed erunt sacerdotes Dei et Christi et regnabunt cum illo mille annis.
REV|20|7|Et cum consummati fuerint mille anni, solvetur Satanas de carcere suo
REV|20|8|et exibit seducere gentes, quae sunt in quattuor angulis terrae, Gog et Magog; congregare eos in proelium, quorum numerus est sicut arena maris.
REV|20|9|Et ascenderunt super latitudinem terrae et circumierunt castra sanctorum et civitatem dilectam. Et descendit ignis de caelo et devoravit eos;
REV|20|10|et Diabolus, qui seducebat eos, missus est in stagnum ignis et sulphuris, ubi et bestia et pseudopropheta, et cruciabuntur die ac nocte in saecula saeculorum.
REV|20|11|Et vidi thronum magnum candidum et sedentem super eum, a cuius aspectu fugit terra et caelum, et locus non est inventus eis.
REV|20|12|Et vidi mortuos, magnos et pusillos, stantes in conspectu throni; et libri aperti sunt. Et alius liber apertus est, qui est vitae; et iudicati sunt mortui ex his, quae scripta erant in libris, secundum opera ipsorum.
REV|20|13|Et dedit mare mortuos, qui in eo erant, et mors et infernus dederunt mortuos, qui in ipsis erant; et iudicati sunt singuli secundum opera ipsorum.
REV|20|14|Et mors et infernus missi sunt in stagnum ignis. Haec mors secunda est, stagnum ignis.
REV|20|15|Et si quis non est inventus in libro vitae scriptus, missus est in stagnum ignis.
REV|21|1|Et vidi caelum novum et ter ram novam; primum enim caelum et prima terra abierunt, et mare iam non est.
REV|21|2|Et civitatem sanctam Ierusalem novam vidi descendentem de caelo a Deo, paratam sicut sponsam ornatam viro suo.
REV|21|3|Et audivi vocem magnam de throno dicentem: "Ecce tabernaculum Dei cum hominibus! Et habitabit cum eis, et ipsi populi eius erunt, et ipse Deus cum eis erit eorum Deus;
REV|21|4|et absterget omnem lacrimam ab oculis eorum, et mors ultra non erit, neque luctus neque clamor neque dolor erit ultra, quia prima abierunt ".
REV|21|5|Et dixit, qui sedebat super throno: " Ecce nova facio omnia ". Et dicit: Scribe: Haec verba fidelia sunt et vera ".
REV|21|6|Et dixit mihi: " Facta sunt! Ego sum Alpha et Omega, principium et finis. Ego sitienti dabo de fonte aquae vivae gratis.
REV|21|7|Qui vicerit, hereditabit haec, et ero illi Deus, et ille erit mihi filius.
REV|21|8|Timidis autem et incredulis et exsecratis et homicidis et fornicatoribus et veneficis et idololatris et omnibus mendacibus, pars illorum erit in stagno ardenti igne et sulphure, quod est mors secunda ".
REV|21|9|Et venit unus de septem angelis habentibus septem phialas plenas septem plagis novissimis et locutus est mecum dicens: " Veni, ostendam tibi sponsam uxorem Agni ".
REV|21|10|Et sustulit me in spiritu super montem magnum et altum et ostendit mihi civitatem sanctam Ierusalem descendentem de caelo a Deo,
REV|21|11|habentem claritatem Dei; lumen eius simile lapidi pretiosissimo, tamquam lapidi iaspidi, in modum crystalli;
REV|21|12|et habebat murum magnum et altum et habebat portas duodecim et super portas angelos duodecim et nomina inscripta, quae sunt duodecim tribuum filiorum Israel.
REV|21|13|Ab oriente portae tres, et ab aquilone portae tres, et ab austro portae tres, et ab occasu portae tres;
REV|21|14|et murus civitatis habens fundamenta duodecim, et super ipsis duodecim nomina duodecim apostolorum Agni.
REV|21|15|Et, qui loquebatur mecum, habebat mensuram arundinem auream, ut metiretur civitatem et portas eius et murum eius.
REV|21|16|Et civitas in quadro posita est, et longitudo eius tanta est quanta et latitudo. Et mensus est civitatem arundine per stadia duodecim milia; longitudo et latitudo et altitudo eius aequales sunt.
REV|21|17|Et mensus est murum eius centum quadraginta quattuor cubitorum, mensura hominis, quae est angeli.
REV|21|18|Et erat structura muri eius ex iaspide, ipsa vero civitas aurum mundum simile vitro mundo.
REV|21|19|Fundamenta muri civitatis omni lapide pretioso ornata: fundamentum primum iaspis, secundus sapphirus, tertius chalcedonius, quartus smaragdus,
REV|21|20|quintus sardonyx, sextus sardinus, septimus chrysolithus, octavus beryllus, nonus topazius, decimus chrysoprasus, undecimus hyacinthus, duodecimus amethystus.
REV|21|21|Et duodecim portae duodecim margaritae sunt, et singulae portae erant ex singulis margaritis. Et platea civitatis aurum mundum tamquam vitrum perlucidum.
REV|21|22|Et templum non vidi in ea: Dominus enim, Deus omnipotens, templum illius est, et Agnus.
REV|21|23|Et civitas non eget sole neque luna, ut luceant ei, nam claritas Dei illuminavit eam, et lucerna eius est Agnus.
REV|21|24|Et ambulabunt gentes per lumen eius, et reges terrae afferunt gloriam suam in illam;
REV|21|25|et portae eius non claudentur per diem, nox enim non erit illic;
REV|21|26|et afferent gloriam et divitias gentium in illam.
REV|21|27|Nec intrabit in ea aliquid coinquinatum et faciens abominationem et mendacium, nisi qui scripti sunt in libro vitae Agni.
REV|22|1|Et ostendit mihi fluvium aquae vitae splendidum tamquam crystallum, procedentem de throno Dei et Agni.
REV|22|2|In medio plateae eius et fluminis ex utraque parte lignum vitae afferens fructus duodecim, per menses singulos reddens fructum suum; et folia ligni ad sanitatem gentium.
REV|22|3|Et omne maledictum non erit amplius. Et thronus Dei et Agni in illa erit; et servi eius servient illi
REV|22|4|et videbunt faciem eius, et nomen eius in frontibus eorum.
REV|22|5|Et nox ultra non erit, et non egent lumine lucernae neque lumine solis, quoniam Dominus Deus illuminabit super illos, et regnabunt in saecula saeculorum.
REV|22|6|Et dixit mihi: " Haec verba fidelissima et vera sunt, et Dominus, Deus spirituum prophetarum, misit angelum suum ostendere servis suis, quae oportet fieri cito.
REV|22|7|Et ecce venio velociter. Beatus, qui servat verba prophetiae libri huius.
REV|22|8|Et ego Ioannes, qui audivi et vidi haec. Et postquam audissem et vidissem, cecidi, ut adorarem ante pedes angeli, qui mihi haec ostendebat.
REV|22|9|Et dicit mihi: " Vide, ne feceris. Conservus tuus sum et fratrum tuorum prophetarum et eorum, qui servant verba libri huius; Deum adora! ".
REV|22|10|Et dicit mihi: " Ne signaveris verba prophetiae libri huius; tempus enim prope est!
REV|22|11|Qui nocet, noceat adhuc; et, qui sordidus est, sordescat adhuc; et iustus iustitiam faciat adhuc; et sanctus sanctificetur adhuc.
REV|22|12|Ecce venio cito, et merces mea mecum est, reddere unicuique sicut opus eius est.
REV|22|13|Ego Alpha et Omega, primus et novissimus, principium et finis.
REV|22|14|Beati, qui lavant stolas suas, ut sit potestas eorum super lignum vitae, et per portas intrent in civitatem.
REV|22|15|Foris canes et venefici et impudici et homicidae et idolis servientes et omnis, qui amat et facit mendacium!
REV|22|16|Ego Iesus misi angelum meum testificari vobis haec super ecclesiis. Ego sum radix et genus David, stella splendida matutina ".
REV|22|17|Et Spiritus et sponsa dicunt: " Veni! ". Et, qui audit, dicat: " Veni!. Et, qui sitit, veniat; qui vult, accipiat aquam vitae gratis.
REV|22|18|Contestor ego omni audienti verba prophetiae libri huius: Si quis apposuerit ad haec, apponet Deus super illum plagas scriptas in libro isto;
REV|22|19|et si quis abstulerit de verbis libri prophetiae huius, auferet Deus partem eius de ligno vitae et de civitate sancta, de his, quae scripta sunt in libro isto.
REV|22|20|Dicit, qui testimonium perhibet istorum: " Etiam, venio cito ". Amen. Veni, Domine Iesu! ".
REV|22|21|Gratia Domini Iesu cum omnibus.
