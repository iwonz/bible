MATT|1|1|The book of the generation of Jesus Christ, the son of David, the son of Abraham.
MATT|1|2|Abraham begat Isaac; and Isaac begat Jacob; and Jacob begat Judas and his brethren;
MATT|1|3|And Judas begat Phares and Zara of Thamar; and Phares begat Esrom; and Esrom begat Aram;
MATT|1|4|And Aram begat Aminadab; and Aminadab begat Naasson; and Naasson begat Salmon;
MATT|1|5|And Salmon begat Booz of Rachab; and Booz begat Obed of Ruth; and Obed begat Jesse;
MATT|1|6|And Jesse begat David the king; and David the king begat Solomon of her that had been the wife of Urias;
MATT|1|7|And Solomon begat Roboam; and Roboam begat Abia; and Abia begat Asa;
MATT|1|8|And Asa begat Josaphat; and Josaphat begat Joram; and Joram begat Ozias;
MATT|1|9|And Ozias begat Joatham; and Joatham begat Achaz; and Achaz begat Ezekias;
MATT|1|10|And Ezekias begat Manasses; and Manasses begat Amon; and Amon begat Josias;
MATT|1|11|And Josias begat Jechonias and his brethren, about the time they were carried away to Babylon:
MATT|1|12|And after they were brought to Babylon, Jechonias begat Salathiel; and Salathiel begat Zorobabel;
MATT|1|13|And Zorobabel begat Abiud; and Abiud begat Eliakim; and Eliakim begat Azor;
MATT|1|14|And Azor begat Sadoc; and Sadoc begat Achim; and Achim begat Eliud;
MATT|1|15|And Eliud begat Eleazar; and Eleazar begat Matthan; and Matthan begat Jacob;
MATT|1|16|And Jacob begat Joseph the husband of Mary, of whom was born Jesus, who is called Christ.
MATT|1|17|So all the generations from Abraham to David are fourteen generations; and from David until the carrying away into Babylon are fourteen generations; and from the carrying away into Babylon unto Christ are fourteen generations.
MATT|1|18|Now the birth of Jesus Christ was on this wise: When as his mother Mary was espoused to Joseph, before they came together, she was found with child of the Holy Ghost.
MATT|1|19|Then Joseph her husband, being a just man, and not willing to make her a publick example, was minded to put her away privily.
MATT|1|20|But while he thought on these things, behold, the angel of the LORD appeared unto him in a dream, saying, Joseph, thou son of David, fear not to take unto thee Mary thy wife: for that which is conceived in her is of the Holy Ghost.
MATT|1|21|And she shall bring forth a son, and thou shalt call his name JESUS: for he shall save his people from their sins.
MATT|1|22|Now all this was done, that it might be fulfilled which was spoken of the Lord by the prophet, saying,
MATT|1|23|Behold, a virgin shall be with child, and shall bring forth a son, and they shall call his name Emmanuel, which being interpreted is, God with us.
MATT|1|24|Then Joseph being raised from sleep did as the angel of the Lord had bidden him, and took unto him his wife:
MATT|1|25|And knew her not till she had brought forth her firstborn son: and he called his name JESUS.
MATT|2|1|Now when Jesus was born in Bethlehem of Judaea in the days of Herod the king, behold, there came wise men from the east to Jerusalem,
MATT|2|2|Saying, Where is he that is born King of the Jews? for we have seen his star in the east, and are come to worship him.
MATT|2|3|When Herod the king had heard these things, he was troubled, and all Jerusalem with him.
MATT|2|4|And when he had gathered all the chief priests and scribes of the people together, he demanded of them where Christ should be born.
MATT|2|5|And they said unto him, In Bethlehem of Judaea: for thus it is written by the prophet,
MATT|2|6|And thou Bethlehem, in the land of Juda, art not the least among the princes of Juda: for out of thee shall come a Governor, that shall rule my people Israel.
MATT|2|7|Then Herod, when he had privily called the wise men, enquired of them diligently what time the star appeared.
MATT|2|8|And he sent them to Bethlehem, and said, Go and search diligently for the young child; and when ye have found him, bring me word again, that I may come and worship him also.
MATT|2|9|When they had heard the king, they departed; and, lo, the star, which they saw in the east, went before them, till it came and stood over where the young child was.
MATT|2|10|When they saw the star, they rejoiced with exceeding great joy.
MATT|2|11|And when they were come into the house, they saw the young child with Mary his mother, and fell down, and worshipped him: and when they had opened their treasures, they presented unto him gifts; gold, and frankincense and myrrh.
MATT|2|12|And being warned of God in a dream that they should not return to Herod, they departed into their own country another way.
MATT|2|13|And when they were departed, behold, the angel of the Lord appeareth to Joseph in a dream, saying, Arise, and take the young child and his mother, and flee into Egypt, and be thou there until I bring thee word: for Herod will seek the young child to destroy him.
MATT|2|14|When he arose, he took the young child and his mother by night, and departed into Egypt:
MATT|2|15|And was there until the death of Herod: that it might be fulfilled which was spoken of the Lord by the prophet, saying, Out of Egypt have I called my son.
MATT|2|16|Then Herod, when he saw that he was mocked of the wise men, was exceeding wroth, and sent forth, and slew all the children that were in Bethlehem, and in all the coasts thereof, from two years old and under, according to the time which he had diligently enquired of the wise men.
MATT|2|17|Then was fulfilled that which was spoken by Jeremy the prophet, saying,
MATT|2|18|In Rama was there a voice heard, lamentation, and weeping, and great mourning, Rachel weeping for her children, and would not be comforted, because they are not.
MATT|2|19|But when Herod was dead, behold, an angel of the Lord appeareth in a dream to Joseph in Egypt,
MATT|2|20|Saying, Arise, and take the young child and his mother, and go into the land of Israel: for they are dead which sought the young child's life.
MATT|2|21|And he arose, and took the young child and his mother, and came into the land of Israel.
MATT|2|22|But when he heard that Archelaus did reign in Judaea in the room of his father Herod, he was afraid to go thither: notwithstanding, being warned of God in a dream, he turned aside into the parts of Galilee:
MATT|2|23|And he came and dwelt in a city called Nazareth: that it might be fulfilled which was spoken by the prophets, He shall be called a Nazarene.
MATT|3|1|In those days came John the Baptist, preaching in the wilderness of Judaea,
MATT|3|2|And saying, Repent ye: for the kingdom of heaven is at hand.
MATT|3|3|For this is he that was spoken of by the prophet Esaias, saying, The voice of one crying in the wilderness, Prepare ye the way of the Lord, make his paths straight.
MATT|3|4|And the same John had his raiment of camel's hair, and a leathern girdle about his loins; and his meat was locusts and wild honey.
MATT|3|5|Then went out to him Jerusalem, and all Judaea, and all the region round about Jordan,
MATT|3|6|And were baptized of him in Jordan, confessing their sins.
MATT|3|7|But when he saw many of the Pharisees and Sadducees come to his baptism, he said unto them, O generation of vipers, who hath warned you to flee from the wrath to come?
MATT|3|8|Bring forth therefore fruits meet for repentance:
MATT|3|9|And think not to say within yourselves, We have Abraham to our father: for I say unto you, that God is able of these stones to raise up children unto Abraham.
MATT|3|10|And now also the axe is laid unto the root of the trees: therefore every tree which bringeth not forth good fruit is hewn down, and cast into the fire.
MATT|3|11|I indeed baptize you with water unto repentance: but he that cometh after me is mightier than I, whose shoes I am not worthy to bear: he shall baptize you with the Holy Ghost, and with fire:
MATT|3|12|Whose fan is in his hand, and he will throughly purge his floor, and gather his wheat into the garner; but he will burn up the chaff with unquenchable fire.
MATT|3|13|Then cometh Jesus from Galilee to Jordan unto John, to be baptized of him.
MATT|3|14|But John forbad him, saying, I have need to be baptized of thee, and comest thou to me?
MATT|3|15|And Jesus answering said unto him, Suffer it to be so now: for thus it becometh us to fulfil all righteousness. Then he suffered him.
MATT|3|16|And Jesus, when he was baptized, went up straightway out of the water: and, lo, the heavens were opened unto him, and he saw the Spirit of God descending like a dove, and lighting upon him:
MATT|3|17|And lo a voice from heaven, saying, This is my beloved Son, in whom I am well pleased.
MATT|4|1|Then was Jesus led up of the spirit into the wilderness to be tempted of the devil.
MATT|4|2|And when he had fasted forty days and forty nights, he was afterward an hungred.
MATT|4|3|And when the tempter came to him, he said, If thou be the Son of God, command that these stones be made bread.
MATT|4|4|But he answered and said, It is written, Man shall not live by bread alone, but by every word that proceedeth out of the mouth of God.
MATT|4|5|Then the devil taketh him up into the holy city, and setteth him on a pinnacle of the temple,
MATT|4|6|And saith unto him, If thou be the Son of God, cast thyself down: for it is written, He shall give his angels charge concerning thee: and in their hands they shall bear thee up, lest at any time thou dash thy foot against a stone.
MATT|4|7|Jesus said unto him, It is written again, Thou shalt not tempt the Lord thy God.
MATT|4|8|Again, the devil taketh him up into an exceeding high mountain, and sheweth him all the kingdoms of the world, and the glory of them;
MATT|4|9|And saith unto him, All these things will I give thee, if thou wilt fall down and worship me.
MATT|4|10|Then saith Jesus unto him, Get thee hence, Satan: for it is written, Thou shalt worship the Lord thy God, and him only shalt thou serve.
MATT|4|11|Then the devil leaveth him, and, behold, angels came and ministered unto him.
MATT|4|12|Now when Jesus had heard that John was cast into prison, he departed into Galilee;
MATT|4|13|And leaving Nazareth, he came and dwelt in Capernaum, which is upon the sea coast, in the borders of Zabulon and Nephthalim:
MATT|4|14|That it might be fulfilled which was spoken by Esaias the prophet, saying,
MATT|4|15|The land of Zabulon, and the land of Nephthalim, by the way of the sea, beyond Jordan, Galilee of the Gentiles;
MATT|4|16|The people which sat in darkness saw great light; and to them which sat in the region and shadow of death light is sprung up.
MATT|4|17|From that time Jesus began to preach, and to say, Repent: for the kingdom of heaven is at hand.
MATT|4|18|And Jesus, walking by the sea of Galilee, saw two brethren, Simon called Peter, and Andrew his brother, casting a net into the sea: for they were fishers.
MATT|4|19|And he saith unto them, Follow me, and I will make you fishers of men.
MATT|4|20|And they straightway left their nets, and followed him.
MATT|4|21|And going on from thence, he saw other two brethren, James the son of Zebedee, and John his brother, in a ship with Zebedee their father, mending their nets; and he called them.
MATT|4|22|And they immediately left the ship and their father, and followed him.
MATT|4|23|And Jesus went about all Galilee, teaching in their synagogues, and preaching the gospel of the kingdom, and healing all manner of sickness and all manner of disease among the people.
MATT|4|24|And his fame went throughout all Syria: and they brought unto him all sick people that were taken with divers diseases and torments, and those which were possessed with devils, and those which were lunatick, and those that had the palsy; and he healed them.
MATT|4|25|And there followed him great multitudes of people from Galilee, and from Decapolis, and from Jerusalem, and from Judaea, and from beyond Jordan.
MATT|5|1|And seeing the multitudes, he went up into a mountain: and when he was set, his disciples came unto him:
MATT|5|2|And he opened his mouth, and taught them, saying,
MATT|5|3|Blessed are the poor in spirit: for theirs is the kingdom of heaven.
MATT|5|4|Blessed are they that mourn: for they shall be comforted.
MATT|5|5|Blessed are the meek: for they shall inherit the earth.
MATT|5|6|Blessed are they which do hunger and thirst after righteousness: for they shall be filled.
MATT|5|7|Blessed are the merciful: for they shall obtain mercy.
MATT|5|8|Blessed are the pure in heart: for they shall see God.
MATT|5|9|Blessed are the peacemakers: for they shall be called the children of God.
MATT|5|10|Blessed are they which are persecuted for righteousness' sake: for theirs is the kingdom of heaven.
MATT|5|11|Blessed are ye, when men shall revile you, and persecute you, and shall say all manner of evil against you falsely, for my sake.
MATT|5|12|Rejoice, and be exceeding glad: for great is your reward in heaven: for so persecuted they the prophets which were before you.
MATT|5|13|Ye are the salt of the earth: but if the salt have lost his savour, wherewith shall it be salted? it is thenceforth good for nothing, but to be cast out, and to be trodden under foot of men.
MATT|5|14|Ye are the light of the world. A city that is set on an hill cannot be hid.
MATT|5|15|Neither do men light a candle, and put it under a bushel, but on a candlestick; and it giveth light unto all that are in the house.
MATT|5|16|Let your light so shine before men, that they may see your good works, and glorify your Father which is in heaven.
MATT|5|17|Think not that I am come to destroy the law, or the prophets: I am not come to destroy, but to fulfil.
MATT|5|18|For verily I say unto you, Till heaven and earth pass, one jot or one tittle shall in no wise pass from the law, till all be fulfilled.
MATT|5|19|Whosoever therefore shall break one of these least commandments, and shall teach men so, he shall be called the least in the kingdom of heaven: but whosoever shall do and teach them, the same shall be called great in the kingdom of heaven.
MATT|5|20|For I say unto you, That except your righteousness shall exceed the righteousness of the scribes and Pharisees, ye shall in no case enter into the kingdom of heaven.
MATT|5|21|Ye have heard that it was said of them of old time, Thou shalt not kill; and whosoever shall kill shall be in danger of the judgment:
MATT|5|22|But I say unto you, That whosoever is angry with his brother without a cause shall be in danger of the judgment: and whosoever shall say to his brother, Raca, shall be in danger of the council: but whosoever shall say, Thou fool, shall be in danger of hell fire.
MATT|5|23|Therefore if thou bring thy gift to the altar, and there rememberest that thy brother hath ought against thee;
MATT|5|24|Leave there thy gift before the altar, and go thy way; first be reconciled to thy brother, and then come and offer thy gift.
MATT|5|25|Agree with thine adversary quickly, whiles thou art in the way with him; lest at any time the adversary deliver thee to the judge, and the judge deliver thee to the officer, and thou be cast into prison.
MATT|5|26|Verily I say unto thee, Thou shalt by no means come out thence, till thou hast paid the uttermost farthing.
MATT|5|27|Ye have heard that it was said by them of old time, Thou shalt not commit adultery:
MATT|5|28|But I say unto you, That whosoever looketh on a woman to lust after her hath committed adultery with her already in his heart.
MATT|5|29|And if thy right eye offend thee, pluck it out, and cast it from thee: for it is profitable for thee that one of thy members should perish, and not that thy whole body should be cast into hell.
MATT|5|30|And if thy right hand offend thee, cut it off, and cast it from thee: for it is profitable for thee that one of thy members should perish, and not that thy whole body should be cast into hell.
MATT|5|31|It hath been said, Whosoever shall put away his wife, let him give her a writing of divorcement:
MATT|5|32|But I say unto you, That whosoever shall put away his wife, saving for the cause of fornication, causeth her to commit adultery: and whosoever shall marry her that is divorced committeth adultery.
MATT|5|33|Again, ye have heard that it hath been said by them of old time, Thou shalt not forswear thyself, but shalt perform unto the Lord thine oaths:
MATT|5|34|But I say unto you, Swear not at all; neither by heaven; for it is God's throne:
MATT|5|35|Nor by the earth; for it is his footstool: neither by Jerusalem; for it is the city of the great King.
MATT|5|36|Neither shalt thou swear by thy head, because thou canst not make one hair white or black.
MATT|5|37|But let your communication be, Yea, yea; Nay, nay: for whatsoever is more than these cometh of evil.
MATT|5|38|Ye have heard that it hath been said, An eye for an eye, and a tooth for a tooth:
MATT|5|39|But I say unto you, That ye resist not evil: but whosoever shall smite thee on thy right cheek, turn to him the other also.
MATT|5|40|And if any man will sue thee at the law, and take away thy coat, let him have thy cloak also.
MATT|5|41|And whosoever shall compel thee to go a mile, go with him twain.
MATT|5|42|Give to him that asketh thee, and from him that would borrow of thee turn not thou away.
MATT|5|43|Ye have heard that it hath been said, Thou shalt love thy neighbour, and hate thine enemy.
MATT|5|44|But I say unto you, Love your enemies, bless them that curse you, do good to them that hate you, and pray for them which despitefully use you, and persecute you;
MATT|5|45|That ye may be the children of your Father which is in heaven: for he maketh his sun to rise on the evil and on the good, and sendeth rain on the just and on the unjust.
MATT|5|46|For if ye love them which love you, what reward have ye? do not even the publicans the same?
MATT|5|47|And if ye salute your brethren only, what do ye more than others? do not even the publicans so?
MATT|5|48|Be ye therefore perfect, even as your Father which is in heaven is perfect.
MATT|6|1|Take heed that ye do not your alms before men, to be seen of them: otherwise ye have no reward of your Father which is in heaven.
MATT|6|2|Therefore when thou doest thine alms, do not sound a trumpet before thee, as the hypocrites do in the synagogues and in the streets, that they may have glory of men. Verily I say unto you, They have their reward.
MATT|6|3|But when thou doest alms, let not thy left hand know what thy right hand doeth:
MATT|6|4|That thine alms may be in secret: and thy Father which seeth in secret himself shall reward thee openly.
MATT|6|5|And when thou prayest, thou shalt not be as the hypocrites are: for they love to pray standing in the synagogues and in the corners of the streets, that they may be seen of men. Verily I say unto you, They have their reward.
MATT|6|6|But thou, when thou prayest, enter into thy closet, and when thou hast shut thy door, pray to thy Father which is in secret; and thy Father which seeth in secret shall reward thee openly.
MATT|6|7|But when ye pray, use not vain repetitions, as the heathen do: for they think that they shall be heard for their much speaking.
MATT|6|8|Be not ye therefore like unto them: for your Father knoweth what things ye have need of, before ye ask him.
MATT|6|9|After this manner therefore pray ye: Our Father which art in heaven, Hallowed be thy name.
MATT|6|10|Thy kingdom come, Thy will be done in earth, as it is in heaven.
MATT|6|11|Give us this day our daily bread.
MATT|6|12|And forgive us our debts, as we forgive our debtors.
MATT|6|13|And lead us not into temptation, but deliver us from evil: For thine is the kingdom, and the power, and the glory, for ever. Amen.
MATT|6|14|For if ye forgive men their trespasses, your heavenly Father will also forgive you:
MATT|6|15|But if ye forgive not men their trespasses, neither will your Father forgive your trespasses.
MATT|6|16|Moreover when ye fast, be not, as the hypocrites, of a sad countenance: for they disfigure their faces, that they may appear unto men to fast. Verily I say unto you, They have their reward.
MATT|6|17|But thou, when thou fastest, anoint thine head, and wash thy face;
MATT|6|18|That thou appear not unto men to fast, but unto thy Father which is in secret: and thy Father, which seeth in secret, shall reward thee openly.
MATT|6|19|Lay not up for yourselves treasures upon earth, where moth and rust doth corrupt, and where thieves break through and steal:
MATT|6|20|But lay up for yourselves treasures in heaven, where neither moth nor rust doth corrupt, and where thieves do not break through nor steal:
MATT|6|21|For where your treasure is, there will your heart be also.
MATT|6|22|The light of the body is the eye: if therefore thine eye be single, thy whole body shall be full of light.
MATT|6|23|But if thine eye be evil, thy whole body shall be full of darkness. If therefore the light that is in thee be darkness, how great is that darkness!
MATT|6|24|No man can serve two masters: for either he will hate the one, and love the other; or else he will hold to the one, and despise the other. Ye cannot serve God and mammon.
MATT|6|25|Therefore I say unto you, Take no thought for your life, what ye shall eat, or what ye shall drink; nor yet for your body, what ye shall put on. Is not the life more than meat, and the body than raiment?
MATT|6|26|Behold the fowls of the air: for they sow not, neither do they reap, nor gather into barns; yet your heavenly Father feedeth them. Are ye not much better than they?
MATT|6|27|Which of you by taking thought can add one cubit unto his stature?
MATT|6|28|And why take ye thought for raiment? Consider the lilies of the field, how they grow; they toil not, neither do they spin:
MATT|6|29|And yet I say unto you, That even Solomon in all his glory was not arrayed like one of these.
MATT|6|30|Wherefore, if God so clothe the grass of the field, which to day is, and to morrow is cast into the oven, shall he not much more clothe you, O ye of little faith?
MATT|6|31|Therefore take no thought, saying, What shall we eat? or, What shall we drink? or, Wherewithal shall we be clothed?
MATT|6|32|(For after all these things do the Gentiles seek:) for your heavenly Father knoweth that ye have need of all these things.
MATT|6|33|But seek ye first the kingdom of God, and his righteousness; and all these things shall be added unto you.
MATT|6|34|Take therefore no thought for the morrow: for the morrow shall take thought for the things of itself. Sufficient unto the day is the evil thereof.
MATT|7|1|Judge not, that ye be not judged.
MATT|7|2|For with what judgment ye judge, ye shall be judged: and with what measure ye mete, it shall be measured to you again.
MATT|7|3|And why beholdest thou the mote that is in thy brother's eye, but considerest not the beam that is in thine own eye?
MATT|7|4|Or how wilt thou say to thy brother, Let me pull out the mote out of thine eye; and, behold, a beam is in thine own eye?
MATT|7|5|Thou hypocrite, first cast out the beam out of thine own eye; and then shalt thou see clearly to cast out the mote out of thy brother's eye.
MATT|7|6|Give not that which is holy unto the dogs, neither cast ye your pearls before swine, lest they trample them under their feet, and turn again and rend you.
MATT|7|7|Ask, and it shall be given you; seek, and ye shall find; knock, and it shall be opened unto you:
MATT|7|8|For every one that asketh receiveth; and he that seeketh findeth; and to him that knocketh it shall be opened.
MATT|7|9|Or what man is there of you, whom if his son ask bread, will he give him a stone?
MATT|7|10|Or if he ask a fish, will he give him a serpent?
MATT|7|11|If ye then, being evil, know how to give good gifts unto your children, how much more shall your Father which is in heaven give good things to them that ask him?
MATT|7|12|Therefore all things whatsoever ye would that men should do to you, do ye even so to them: for this is the law and the prophets.
MATT|7|13|Enter ye in at the strait gate: for wide is the gate, and broad is the way, that leadeth to destruction, and many there be which go in thereat:
MATT|7|14|Because strait is the gate, and narrow is the way, which leadeth unto life, and few there be that find it.
MATT|7|15|Beware of false prophets, which come to you in sheep's clothing, but inwardly they are ravening wolves.
MATT|7|16|Ye shall know them by their fruits. Do men gather grapes of thorns, or figs of thistles?
MATT|7|17|Even so every good tree bringeth forth good fruit; but a corrupt tree bringeth forth evil fruit.
MATT|7|18|A good tree cannot bring forth evil fruit, neither can a corrupt tree bring forth good fruit.
MATT|7|19|Every tree that bringeth not forth good fruit is hewn down, and cast into the fire.
MATT|7|20|Wherefore by their fruits ye shall know them.
MATT|7|21|Not every one that saith unto me, Lord, Lord, shall enter into the kingdom of heaven; but he that doeth the will of my Father which is in heaven.
MATT|7|22|Many will say to me in that day, Lord, Lord, have we not prophesied in thy name? and in thy name have cast out devils? and in thy name done many wonderful works?
MATT|7|23|And then will I profess unto them, I never knew you: depart from me, ye that work iniquity.
MATT|7|24|Therefore whosoever heareth these sayings of mine, and doeth them, I will liken him unto a wise man, which built his house upon a rock:
MATT|7|25|And the rain descended, and the floods came, and the winds blew, and beat upon that house; and it fell not: for it was founded upon a rock.
MATT|7|26|And every one that heareth these sayings of mine, and doeth them not, shall be likened unto a foolish man, which built his house upon the sand:
MATT|7|27|And the rain descended, and the floods came, and the winds blew, and beat upon that house; and it fell: and great was the fall of it.
MATT|7|28|And it came to pass, when Jesus had ended these sayings, the people were astonished at his doctrine:
MATT|7|29|For he taught them as one having authority, and not as the scribes.
MATT|8|1|When he was come down from the mountain, great multitudes followed him.
MATT|8|2|And, behold, there came a leper and worshipped him, saying, Lord, if thou wilt, thou canst make me clean.
MATT|8|3|And Jesus put forth his hand, and touched him, saying, I will; be thou clean. And immediately his leprosy was cleansed.
MATT|8|4|And Jesus saith unto him, See thou tell no man; but go thy way, shew thyself to the priest, and offer the gift that Moses commanded, for a testimony unto them.
MATT|8|5|And when Jesus was entered into Capernaum, there came unto him a centurion, beseeching him,
MATT|8|6|And saying, Lord, my servant lieth at home sick of the palsy, grievously tormented.
MATT|8|7|And Jesus saith unto him, I will come and heal him.
MATT|8|8|The centurion answered and said, Lord, I am not worthy that thou shouldest come under my roof: but speak the word only, and my servant shall be healed.
MATT|8|9|For I am a man under authority, having soldiers under me: and I say to this man, Go, and he goeth; and to another, Come, and he cometh; and to my servant, Do this, and he doeth it.
MATT|8|10|When Jesus heard it, he marvelled, and said to them that followed, Verily I say unto you, I have not found so great faith, no, not in Israel.
MATT|8|11|And I say unto you, That many shall come from the east and west, and shall sit down with Abraham, and Isaac, and Jacob, in the kingdom of heaven.
MATT|8|12|But the children of the kingdom shall be cast out into outer darkness: there shall be weeping and gnashing of teeth.
MATT|8|13|And Jesus said unto the centurion, Go thy way; and as thou hast believed, so be it done unto thee. And his servant was healed in the selfsame hour.
MATT|8|14|And when Jesus was come into Peter's house, he saw his wife's mother laid, and sick of a fever.
MATT|8|15|And he touched her hand, and the fever left her: and she arose, and ministered unto them.
MATT|8|16|When the even was come, they brought unto him many that were possessed with devils: and he cast out the spirits with his word, and healed all that were sick:
MATT|8|17|That it might be fulfilled which was spoken by Esaias the prophet, saying, Himself took our infirmities, and bare our sicknesses.
MATT|8|18|Now when Jesus saw great multitudes about him, he gave commandment to depart unto the other side.
MATT|8|19|And a certain scribe came, and said unto him, Master, I will follow thee whithersoever thou goest.
MATT|8|20|And Jesus saith unto him, The foxes have holes, and the birds of the air have nests; but the Son of man hath not where to lay his head.
MATT|8|21|And another of his disciples said unto him, Lord, suffer me first to go and bury my father.
MATT|8|22|But Jesus said unto him, Follow me; and let the dead bury their dead.
MATT|8|23|And when he was entered into a ship, his disciples followed him.
MATT|8|24|And, behold, there arose a great tempest in the sea, insomuch that the ship was covered with the waves: but he was asleep.
MATT|8|25|And his disciples came to him, and awoke him, saying, Lord, save us: we perish.
MATT|8|26|And he saith unto them, Why are ye fearful, O ye of little faith? Then he arose, and rebuked the winds and the sea; and there was a great calm.
MATT|8|27|But the men marvelled, saying, What manner of man is this, that even the winds and the sea obey him!
MATT|8|28|And when he was come to the other side into the country of the Gergesenes, there met him two possessed with devils, coming out of the tombs, exceeding fierce, so that no man might pass by that way.
MATT|8|29|And, behold, they cried out, saying, What have we to do with thee, Jesus, thou Son of God? art thou come hither to torment us before the time?
MATT|8|30|And there was a good way off from them an herd of many swine feeding.
MATT|8|31|So the devils besought him, saying, If thou cast us out, suffer us to go away into the herd of swine.
MATT|8|32|And he said unto them, Go. And when they were come out, they went into the herd of swine: and, behold, the whole herd of swine ran violently down a steep place into the sea, and perished in the waters.
MATT|8|33|And they that kept them fled, and went their ways into the city, and told every thing, and what was befallen to the possessed of the devils.
MATT|8|34|And, behold, the whole city came out to meet Jesus: and when they saw him, they besought him that he would depart out of their coasts.
MATT|9|1|And he entered into a ship, and passed over, and came into his own city.
MATT|9|2|And, behold, they brought to him a man sick of the palsy, lying on a bed: and Jesus seeing their faith said unto the sick of the palsy; Son, be of good cheer; thy sins be forgiven thee.
MATT|9|3|And, behold, certain of the scribes said within themselves, This man blasphemeth.
MATT|9|4|And Jesus knowing their thoughts said, Wherefore think ye evil in your hearts?
MATT|9|5|For whether is easier, to say, Thy sins be forgiven thee; or to say, Arise, and walk?
MATT|9|6|But that ye may know that the Son of man hath power on earth to forgive sins, (then saith he to the sick of the palsy,) Arise, take up thy bed, and go unto thine house.
MATT|9|7|And he arose, and departed to his house.
MATT|9|8|But when the multitudes saw it, they marvelled, and glorified God, which had given such power unto men.
MATT|9|9|And as Jesus passed forth from thence, he saw a man, named Matthew, sitting at the receipt of custom: and he saith unto him, Follow me. And he arose, and followed him.
MATT|9|10|And it came to pass, as Jesus sat at meat in the house, behold, many publicans and sinners came and sat down with him and his disciples.
MATT|9|11|And when the Pharisees saw it, they said unto his disciples, Why eateth your Master with publicans and sinners?
MATT|9|12|But when Jesus heard that, he said unto them, They that be whole need not a physician, but they that are sick.
MATT|9|13|But go ye and learn what that meaneth, I will have mercy, and not sacrifice: for I am not come to call the righteous, but sinners to repentance.
MATT|9|14|Then came to him the disciples of John, saying, Why do we and the Pharisees fast oft, but thy disciples fast not?
MATT|9|15|And Jesus said unto them, Can the children of the bridechamber mourn, as long as the bridegroom is with them? but the days will come, when the bridegroom shall be taken from them, and then shall they fast.
MATT|9|16|No man putteth a piece of new cloth unto an old garment, for that which is put in to fill it up taketh from the garment, and the rent is made worse.
MATT|9|17|Neither do men put new wine into old bottles: else the bottles break, and the wine runneth out, and the bottles perish: but they put new wine into new bottles, and both are preserved.
MATT|9|18|While he spake these things unto them, behold, there came a certain ruler, and worshipped him, saying, My daughter is even now dead: but come and lay thy hand upon her, and she shall live.
MATT|9|19|And Jesus arose, and followed him, and so did his disciples.
MATT|9|20|And, behold, a woman, which was diseased with an issue of blood twelve years, came behind him, and touched the hem of his garment:
MATT|9|21|For she said within herself, If I may but touch his garment, I shall be whole.
MATT|9|22|But Jesus turned him about, and when he saw her, he said, Daughter, be of good comfort; thy faith hath made thee whole. And the woman was made whole from that hour.
MATT|9|23|And when Jesus came into the ruler's house, and saw the minstrels and the people making a noise,
MATT|9|24|He said unto them, Give place: for the maid is not dead, but sleepeth. And they laughed him to scorn.
MATT|9|25|But when the people were put forth, he went in, and took her by the hand, and the maid arose.
MATT|9|26|And the fame hereof went abroad into all that land.
MATT|9|27|And when Jesus departed thence, two blind men followed him, crying, and saying, Thou son of David, have mercy on us.
MATT|9|28|And when he was come into the house, the blind men came to him: and Jesus saith unto them, Believe ye that I am able to do this? They said unto him, Yea, Lord.
MATT|9|29|Then touched he their eyes, saying, According to your faith be it unto you.
MATT|9|30|And their eyes were opened; and Jesus straitly charged them, saying, See that no man know it.
MATT|9|31|But they, when they were departed, spread abroad his fame in all that country.
MATT|9|32|As they went out, behold, they brought to him a dumb man possessed with a devil.
MATT|9|33|And when the devil was cast out, the dumb spake: and the multitudes marvelled, saying, It was never so seen in Israel.
MATT|9|34|But the Pharisees said, He casteth out devils through the prince of the devils.
MATT|9|35|And Jesus went about all the cities and villages, teaching in their synagogues, and preaching the gospel of the kingdom, and healing every sickness and every disease among the people.
MATT|9|36|But when he saw the multitudes, he was moved with compassion on them, because they fainted, and were scattered abroad, as sheep having no shepherd.
MATT|9|37|Then saith he unto his disciples, The harvest truly is plenteous, but the labourers are few;
MATT|9|38|Pray ye therefore the Lord of the harvest, that he will send forth labourers into his harvest.
MATT|10|1|And when he had called unto him his twelve disciples, he gave them power against unclean spirits, to cast them out, and to heal all manner of sickness and all manner of disease.
MATT|10|2|Now the names of the twelve apostles are these; The first, Simon, who is called Peter, and Andrew his brother; James the son of Zebedee, and John his brother;
MATT|10|3|Philip, and Bartholomew; Thomas, and Matthew the publican; James the son of Alphaeus, and Lebbaeus, whose surname was Thaddaeus;
MATT|10|4|Simon the Canaanite, and Judas Iscariot, who also betrayed him.
MATT|10|5|These twelve Jesus sent forth, and commanded them, saying, Go not into the way of the Gentiles, and into any city of the Samaritans enter ye not:
MATT|10|6|But go rather to the lost sheep of the house of Israel.
MATT|10|7|And as ye go, preach, saying, The kingdom of heaven is at hand.
MATT|10|8|Heal the sick, cleanse the lepers, raise the dead, cast out devils: freely ye have received, freely give.
MATT|10|9|Provide neither gold, nor silver, nor brass in your purses,
MATT|10|10|Nor scrip for your journey, neither two coats, neither shoes, nor yet staves: for the workman is worthy of his meat.
MATT|10|11|And into whatsoever city or town ye shall enter, enquire who in it is worthy; and there abide till ye go thence.
MATT|10|12|And when ye come into an house, salute it.
MATT|10|13|And if the house be worthy, let your peace come upon it: but if it be not worthy, let your peace return to you.
MATT|10|14|And whosoever shall not receive you, nor hear your words, when ye depart out of that house or city, shake off the dust of your feet.
MATT|10|15|Verily I say unto you, It shall be more tolerable for the land of Sodom and Gomorrha in the day of judgment, than for that city.
MATT|10|16|Behold, I send you forth as sheep in the midst of wolves: be ye therefore wise as serpents, and harmless as doves.
MATT|10|17|But beware of men: for they will deliver you up to the councils, and they will scourge you in their synagogues;
MATT|10|18|And ye shall be brought before governors and kings for my sake, for a testimony against them and the Gentiles.
MATT|10|19|But when they deliver you up, take no thought how or what ye shall speak: for it shall be given you in that same hour what ye shall speak.
MATT|10|20|For it is not ye that speak, but the Spirit of your Father which speaketh in you.
MATT|10|21|And the brother shall deliver up the brother to death, and the father the child: and the children shall rise up against their parents, and cause them to be put to death.
MATT|10|22|And ye shall be hated of all men for my name's sake: but he that endureth to the end shall be saved.
MATT|10|23|But when they persecute you in this city, flee ye into another: for verily I say unto you, Ye shall not have gone over the cities of Israel, till the Son of man be come.
MATT|10|24|The disciple is not above his master, nor the servant above his lord.
MATT|10|25|It is enough for the disciple that he be as his master, and the servant as his lord. If they have called the master of the house Beelzebub, how much more shall they call them of his household?
MATT|10|26|Fear them not therefore: for there is nothing covered, that shall not be revealed; and hid, that shall not be known.
MATT|10|27|What I tell you in darkness, that speak ye in light: and what ye hear in the ear, that preach ye upon the housetops.
MATT|10|28|And fear not them which kill the body, but are not able to kill the soul: but rather fear him which is able to destroy both soul and body in hell.
MATT|10|29|Are not two sparrows sold for a farthing? and one of them shall not fall on the ground without your Father.
MATT|10|30|But the very hairs of your head are all numbered.
MATT|10|31|Fear ye not therefore, ye are of more value than many sparrows.
MATT|10|32|Whosoever therefore shall confess me before men, him will I confess also before my Father which is in heaven.
MATT|10|33|But whosoever shall deny me before men, him will I also deny before my Father which is in heaven.
MATT|10|34|Think not that I am come to send peace on earth: I came not to send peace, but a sword.
MATT|10|35|For I am come to set a man at variance against his father, and the daughter against her mother, and the daughter in law against her mother in law.
MATT|10|36|And a man's foes shall be they of his own household.
MATT|10|37|He that loveth father or mother more than me is not worthy of me: and he that loveth son or daughter more than me is not worthy of me.
MATT|10|38|And he that taketh not his cross, and followeth after me, is not worthy of me.
MATT|10|39|He that findeth his life shall lose it: and he that loseth his life for my sake shall find it.
MATT|10|40|He that receiveth you receiveth me, and he that receiveth me receiveth him that sent me.
MATT|10|41|He that receiveth a prophet in the name of a prophet shall receive a prophet's reward; and he that receiveth a righteous man in the name of a righteous man shall receive a righteous man's reward.
MATT|10|42|And whosoever shall give to drink unto one of these little ones a cup of cold water only in the name of a disciple, verily I say unto you, he shall in no wise lose his reward.
MATT|11|1|And it came to pass, when Jesus had made an end of commanding his twelve disciples, he departed thence to teach and to preach in their cities.
MATT|11|2|Now when John had heard in the prison the works of Christ, he sent two of his disciples,
MATT|11|3|And said unto him, Art thou he that should come, or do we look for another?
MATT|11|4|Jesus answered and said unto them, Go and shew John again those things which ye do hear and see:
MATT|11|5|The blind receive their sight, and the lame walk, the lepers are cleansed, and the deaf hear, the dead are raised up, and the poor have the gospel preached to them.
MATT|11|6|And blessed is he, whosoever shall not be offended in me.
MATT|11|7|And as they departed, Jesus began to say unto the multitudes concerning John, What went ye out into the wilderness to see? A reed shaken with the wind?
MATT|11|8|But what went ye out for to see? A man clothed in soft raiment? behold, they that wear soft clothing are in kings' houses.
MATT|11|9|But what went ye out for to see? A prophet? yea, I say unto you, and more than a prophet.
MATT|11|10|For this is he, of whom it is written, Behold, I send my messenger before thy face, which shall prepare thy way before thee.
MATT|11|11|Verily I say unto you, Among them that are born of women there hath not risen a greater than John the Baptist: notwithstanding he that is least in the kingdom of heaven is greater than he.
MATT|11|12|And from the days of John the Baptist until now the kingdom of heaven suffereth violence, and the violent take it by force.
MATT|11|13|For all the prophets and the law prophesied until John.
MATT|11|14|And if ye will receive it, this is Elias, which was for to come.
MATT|11|15|He that hath ears to hear, let him hear.
MATT|11|16|But whereunto shall I liken this generation? It is like unto children sitting in the markets, and calling unto their fellows,
MATT|11|17|And saying, We have piped unto you, and ye have not danced; we have mourned unto you, and ye have not lamented.
MATT|11|18|For John came neither eating nor drinking, and they say, He hath a devil.
MATT|11|19|The Son of man came eating and drinking, and they say, Behold a man gluttonous, and a winebibber, a friend of publicans and sinners. But wisdom is justified of her children.
MATT|11|20|Then began he to upbraid the cities wherein most of his mighty works were done, because they repented not:
MATT|11|21|Woe unto thee, Chorazin! woe unto thee, Bethsaida! for if the mighty works, which were done in you, had been done in Tyre and Sidon, they would have repented long ago in sackcloth and ashes.
MATT|11|22|But I say unto you, It shall be more tolerable for Tyre and Sidon at the day of judgment, than for you.
MATT|11|23|And thou, Capernaum, which art exalted unto heaven, shalt be brought down to hell: for if the mighty works, which have been done in thee, had been done in Sodom, it would have remained until this day.
MATT|11|24|But I say unto you, That it shall be more tolerable for the land of Sodom in the day of judgment, than for thee.
MATT|11|25|At that time Jesus answered and said, I thank thee, O Father, Lord of heaven and earth, because thou hast hid these things from the wise and prudent, and hast revealed them unto babes.
MATT|11|26|Even so, Father: for so it seemed good in thy sight.
MATT|11|27|All things are delivered unto me of my Father: and no man knoweth the Son, but the Father; neither knoweth any man the Father, save the Son, and he to whomsoever the Son will reveal him.
MATT|11|28|Come unto me, all ye that labour and are heavy laden, and I will give you rest.
MATT|11|29|Take my yoke upon you, and learn of me; for I am meek and lowly in heart: and ye shall find rest unto your souls.
MATT|11|30|For my yoke is easy, and my burden is light.
MATT|12|1|At that time Jesus went on the sabbath day through the corn; and his disciples were an hungred, and began to pluck the ears of corn and to eat.
MATT|12|2|But when the Pharisees saw it, they said unto him, Behold, thy disciples do that which is not lawful to do upon the sabbath day.
MATT|12|3|But he said unto them, Have ye not read what David did, when he was an hungred, and they that were with him;
MATT|12|4|How he entered into the house of God, and did eat the shewbread, which was not lawful for him to eat, neither for them which were with him, but only for the priests?
MATT|12|5|Or have ye not read in the law, how that on the sabbath days the priests in the temple profane the sabbath, and are blameless?
MATT|12|6|But I say unto you, That in this place is one greater than the temple.
MATT|12|7|But if ye had known what this meaneth, I will have mercy, and not sacrifice, ye would not have condemned the guiltless.
MATT|12|8|For the Son of man is Lord even of the sabbath day.
MATT|12|9|And when he was departed thence, he went into their synagogue:
MATT|12|10|And, behold, there was a man which had his hand withered. And they asked him, saying, Is it lawful to heal on the sabbath days? that they might accuse him.
MATT|12|11|And he said unto them, What man shall there be among you, that shall have one sheep, and if it fall into a pit on the sabbath day, will he not lay hold on it, and lift it out?
MATT|12|12|How much then is a man better than a sheep? Wherefore it is lawful to do well on the sabbath days.
MATT|12|13|Then saith he to the man, Stretch forth thine hand. And he stretched it forth; and it was restored whole, like as the other.
MATT|12|14|Then the Pharisees went out, and held a council against him, how they might destroy him.
MATT|12|15|But when Jesus knew it, he withdrew himself from thence: and great multitudes followed him, and he healed them all;
MATT|12|16|And charged them that they should not make him known:
MATT|12|17|That it might be fulfilled which was spoken by Esaias the prophet, saying,
MATT|12|18|Behold my servant, whom I have chosen; my beloved, in whom my soul is well pleased: I will put my spirit upon him, and he shall shew judgment to the Gentiles.
MATT|12|19|He shall not strive, nor cry; neither shall any man hear his voice in the streets.
MATT|12|20|A bruised reed shall he not break, and smoking flax shall he not quench, till he send forth judgment unto victory.
MATT|12|21|And in his name shall the Gentiles trust.
MATT|12|22|Then was brought unto him one possessed with a devil, blind, and dumb: and he healed him, insomuch that the blind and dumb both spake and saw.
MATT|12|23|And all the people were amazed, and said, Is not this the son of David?
MATT|12|24|But when the Pharisees heard it, they said, This fellow doth not cast out devils, but by Beelzebub the prince of the devils.
MATT|12|25|And Jesus knew their thoughts, and said unto them, Every kingdom divided against itself is brought to desolation; and every city or house divided against itself shall not stand:
MATT|12|26|And if Satan cast out Satan, he is divided against himself; how shall then his kingdom stand?
MATT|12|27|And if I by Beelzebub cast out devils, by whom do your children cast them out? therefore they shall be your judges.
MATT|12|28|But if I cast out devils by the Spirit of God, then the kingdom of God is come unto you.
MATT|12|29|Or else how can one enter into a strong man's house, and spoil his goods, except he first bind the strong man? and then he will spoil his house.
MATT|12|30|He that is not with me is against me; and he that gathereth not with me scattereth abroad.
MATT|12|31|Wherefore I say unto you, All manner of sin and blasphemy shall be forgiven unto men: but the blasphemy against the Holy Ghost shall not be forgiven unto men.
MATT|12|32|And whosoever speaketh a word against the Son of man, it shall be forgiven him: but whosoever speaketh against the Holy Ghost, it shall not be forgiven him, neither in this world, neither in the world to come.
MATT|12|33|Either make the tree good, and his fruit good; or else make the tree corrupt, and his fruit corrupt: for the tree is known by his fruit.
MATT|12|34|O generation of vipers, how can ye, being evil, speak good things? for out of the abundance of the heart the mouth speaketh.
MATT|12|35|A good man out of the good treasure of the heart bringeth forth good things: and an evil man out of the evil treasure bringeth forth evil things.
MATT|12|36|But I say unto you, That every idle word that men shall speak, they shall give account thereof in the day of judgment.
MATT|12|37|For by thy words thou shalt be justified, and by thy words thou shalt be condemned.
MATT|12|38|Then certain of the scribes and of the Pharisees answered, saying, Master, we would see a sign from thee.
MATT|12|39|But he answered and said unto them, An evil and adulterous generation seeketh after a sign; and there shall no sign be given to it, but the sign of the prophet Jonas:
MATT|12|40|For as Jonas was three days and three nights in the whale's belly; so shall the Son of man be three days and three nights in the heart of the earth.
MATT|12|41|The men of Nineveh shall rise in judgment with this generation, and shall condemn it: because they repented at the preaching of Jonas; and, behold, a greater than Jonas is here.
MATT|12|42|The queen of the south shall rise up in the judgment with this generation, and shall condemn it: for she came from the uttermost parts of the earth to hear the wisdom of Solomon; and, behold, a greater than Solomon is here.
MATT|12|43|When the unclean spirit is gone out of a man, he walketh through dry places, seeking rest, and findeth none.
MATT|12|44|Then he saith, I will return into my house from whence I came out; and when he is come, he findeth it empty, swept, and garnished.
MATT|12|45|Then goeth he, and taketh with himself seven other spirits more wicked than himself, and they enter in and dwell there: and the last state of that man is worse than the first. Even so shall it be also unto this wicked generation.
MATT|12|46|While he yet talked to the people, behold, his mother and his brethren stood without, desiring to speak with him.
MATT|12|47|Then one said unto him, Behold, thy mother and thy brethren stand without, desiring to speak with thee.
MATT|12|48|But he answered and said unto him that told him, Who is my mother? and who are my brethren?
MATT|12|49|And he stretched forth his hand toward his disciples, and said, Behold my mother and my brethren!
MATT|12|50|For whosoever shall do the will of my Father which is in heaven, the same is my brother, and sister, and mother.
MATT|13|1|The same day went Jesus out of the house, and sat by the sea side.
MATT|13|2|And great multitudes were gathered together unto him, so that he went into a ship, and sat; and the whole multitude stood on the shore.
MATT|13|3|And he spake many things unto them in parables, saying, Behold, a sower went forth to sow;
MATT|13|4|And when he sowed, some seeds fell by the way side, and the fowls came and devoured them up:
MATT|13|5|Some fell upon stony places, where they had not much earth: and forthwith they sprung up, because they had no deepness of earth:
MATT|13|6|And when the sun was up, they were scorched; and because they had no root, they withered away.
MATT|13|7|And some fell among thorns; and the thorns sprung up, and choked them:
MATT|13|8|But other fell into good ground, and brought forth fruit, some an hundredfold, some sixtyfold, some thirtyfold.
MATT|13|9|Who hath ears to hear, let him hear.
MATT|13|10|And the disciples came, and said unto him, Why speakest thou unto them in parables?
MATT|13|11|He answered and said unto them, Because it is given unto you to know the mysteries of the kingdom of heaven, but to them it is not given.
MATT|13|12|For whosoever hath, to him shall be given, and he shall have more abundance: but whosoever hath not, from him shall be taken away even that he hath.
MATT|13|13|Therefore speak I to them in parables: because they seeing see not; and hearing they hear not, neither do they understand.
MATT|13|14|And in them is fulfilled the prophecy of Esaias, which saith, By hearing ye shall hear, and shall not understand; and seeing ye shall see, and shall not perceive:
MATT|13|15|For this people's heart is waxed gross, and their ears are dull of hearing, and their eyes they have closed; lest at any time they should see with their eyes and hear with their ears, and should understand with their heart, and should be converted, and I should heal them.
MATT|13|16|But blessed are your eyes, for they see: and your ears, for they hear.
MATT|13|17|For verily I say unto you, That many prophets and righteous men have desired to see those things which ye see, and have not seen them; and to hear those things which ye hear, and have not heard them.
MATT|13|18|Hear ye therefore the parable of the sower.
MATT|13|19|When any one heareth the word of the kingdom, and understandeth it not, then cometh the wicked one, and catcheth away that which was sown in his heart. This is he which received seed by the way side.
MATT|13|20|But he that received the seed into stony places, the same is he that heareth the word, and anon with joy receiveth it;
MATT|13|21|Yet hath he not root in himself, but dureth for a while: for when tribulation or persecution ariseth because of the word, by and by he is offended.
MATT|13|22|He also that received seed among the thorns is he that heareth the word; and the care of this world, and the deceitfulness of riches, choke the word, and he becometh unfruitful.
MATT|13|23|But he that received seed into the good ground is he that heareth the word, and understandeth it; which also beareth fruit, and bringeth forth, some an hundredfold, some sixty, some thirty.
MATT|13|24|Another parable put he forth unto them, saying, The kingdom of heaven is likened unto a man which sowed good seed in his field:
MATT|13|25|But while men slept, his enemy came and sowed tares among the wheat, and went his way.
MATT|13|26|But when the blade was sprung up, and brought forth fruit, then appeared the tares also.
MATT|13|27|So the servants of the householder came and said unto him, Sir, didst not thou sow good seed in thy field? from whence then hath it tares?
MATT|13|28|He said unto them, An enemy hath done this. The servants said unto him, Wilt thou then that we go and gather them up?
MATT|13|29|But he said, Nay; lest while ye gather up the tares, ye root up also the wheat with them.
MATT|13|30|Let both grow together until the harvest: and in the time of harvest I will say to the reapers, Gather ye together first the tares, and bind them in bundles to burn them: but gather the wheat into my barn.
MATT|13|31|Another parable put he forth unto them, saying, The kingdom of heaven is like to a grain of mustard seed, which a man took, and sowed in his field:
MATT|13|32|Which indeed is the least of all seeds: but when it is grown, it is the greatest among herbs, and becometh a tree, so that the birds of the air come and lodge in the branches thereof.
MATT|13|33|Another parable spake he unto them; The kingdom of heaven is like unto leaven, which a woman took, and hid in three measures of meal, till the whole was leavened.
MATT|13|34|All these things spake Jesus unto the multitude in parables; and without a parable spake he not unto them:
MATT|13|35|That it might be fulfilled which was spoken by the prophet, saying, I will open my mouth in parables; I will utter things which have been kept secret from the foundation of the world.
MATT|13|36|Then Jesus sent the multitude away, and went into the house: and his disciples came unto him, saying, Declare unto us the parable of the tares of the field.
MATT|13|37|He answered and said unto them, He that soweth the good seed is the Son of man;
MATT|13|38|The field is the world; the good seed are the children of the kingdom; but the tares are the children of the wicked one;
MATT|13|39|The enemy that sowed them is the devil; the harvest is the end of the world; and the reapers are the angels.
MATT|13|40|As therefore the tares are gathered and burned in the fire; so shall it be in the end of this world.
MATT|13|41|The Son of man shall send forth his angels, and they shall gather out of his kingdom all things that offend, and them which do iniquity;
MATT|13|42|And shall cast them into a furnace of fire: there shall be wailing and gnashing of teeth.
MATT|13|43|Then shall the righteous shine forth as the sun in the kingdom of their Father. Who hath ears to hear, let him hear.
MATT|13|44|Again, the kingdom of heaven is like unto treasure hid in a field; the which when a man hath found, he hideth, and for joy thereof goeth and selleth all that he hath, and buyeth that field.
MATT|13|45|Again, the kingdom of heaven is like unto a merchant man, seeking goodly pearls:
MATT|13|46|Who, when he had found one pearl of great price, went and sold all that he had, and bought it.
MATT|13|47|Again, the kingdom of heaven is like unto a net, that was cast into the sea, and gathered of every kind:
MATT|13|48|Which, when it was full, they drew to shore, and sat down, and gathered the good into vessels, but cast the bad away.
MATT|13|49|So shall it be at the end of the world: the angels shall come forth, and sever the wicked from among the just,
MATT|13|50|And shall cast them into the furnace of fire: there shall be wailing and gnashing of teeth.
MATT|13|51|Jesus saith unto them, Have ye understood all these things? They say unto him, Yea, Lord.
MATT|13|52|Then said he unto them, Therefore every scribe which is instructed unto the kingdom of heaven is like unto a man that is an householder, which bringeth forth out of his treasure things new and old.
MATT|13|53|And it came to pass, that when Jesus had finished these parables, he departed thence.
MATT|13|54|And when he was come into his own country, he taught them in their synagogue, insomuch that they were astonished, and said, Whence hath this man this wisdom, and these mighty works?
MATT|13|55|Is not this the carpenter's son? is not his mother called Mary? and his brethren, James, and Joses, and Simon, and Judas?
MATT|13|56|And his sisters, are they not all with us? Whence then hath this man all these things?
MATT|13|57|And they were offended in him. But Jesus said unto them, A prophet is not without honour, save in his own country, and in his own house.
MATT|13|58|And he did not many mighty works there because of their unbelief.
MATT|14|1|At that time Herod the tetrarch heard of the fame of Jesus,
MATT|14|2|And said unto his servants, This is John the Baptist; he is risen from the dead; and therefore mighty works do shew forth themselves in him.
MATT|14|3|For Herod had laid hold on John, and bound him, and put him in prison for Herodias' sake, his brother Philip's wife.
MATT|14|4|For John said unto him, It is not lawful for thee to have her.
MATT|14|5|And when he would have put him to death, he feared the multitude, because they counted him as a prophet.
MATT|14|6|But when Herod's birthday was kept, the daughter of Herodias danced before them, and pleased Herod.
MATT|14|7|Whereupon he promised with an oath to give her whatsoever she would ask.
MATT|14|8|And she, being before instructed of her mother, said, Give me here John Baptist's head in a charger.
MATT|14|9|And the king was sorry: nevertheless for the oath's sake, and them which sat with him at meat, he commanded it to be given her.
MATT|14|10|And he sent, and beheaded John in the prison.
MATT|14|11|And his head was brought in a charger, and given to the damsel: and she brought it to her mother.
MATT|14|12|And his disciples came, and took up the body, and buried it, and went and told Jesus.
MATT|14|13|When Jesus heard of it, he departed thence by ship into a desert place apart: and when the people had heard thereof, they followed him on foot out of the cities.
MATT|14|14|And Jesus went forth, and saw a great multitude, and was moved with compassion toward them, and he healed their sick.
MATT|14|15|And when it was evening, his disciples came to him, saying, This is a desert place, and the time is now past; send the multitude away, that they may go into the villages, and buy themselves victuals.
MATT|14|16|But Jesus said unto them, They need not depart; give ye them to eat.
MATT|14|17|And they say unto him, We have here but five loaves, and two fishes.
MATT|14|18|He said, Bring them hither to me.
MATT|14|19|And he commanded the multitude to sit down on the grass, and took the five loaves, and the two fishes, and looking up to heaven, he blessed, and brake, and gave the loaves to his disciples, and the disciples to the multitude.
MATT|14|20|And they did all eat, and were filled: and they took up of the fragments that remained twelve baskets full.
MATT|14|21|And they that had eaten were about five thousand men, beside women and children.
MATT|14|22|And straightway Jesus constrained his disciples to get into a ship, and to go before him unto the other side, while he sent the multitudes away.
MATT|14|23|And when he had sent the multitudes away, he went up into a mountain apart to pray: and when the evening was come, he was there alone.
MATT|14|24|But the ship was now in the midst of the sea, tossed with waves: for the wind was contrary.
MATT|14|25|And in the fourth watch of the night Jesus went unto them, walking on the sea.
MATT|14|26|And when the disciples saw him walking on the sea, they were troubled, saying, It is a spirit; and they cried out for fear.
MATT|14|27|But straightway Jesus spake unto them, saying, Be of good cheer; it is I; be not afraid.
MATT|14|28|And Peter answered him and said, Lord, if it be thou, bid me come unto thee on the water.
MATT|14|29|And he said, Come. And when Peter was come down out of the ship, he walked on the water, to go to Jesus.
MATT|14|30|But when he saw the wind boisterous, he was afraid; and beginning to sink, he cried, saying, Lord, save me.
MATT|14|31|And immediately Jesus stretched forth his hand, and caught him, and said unto him, O thou of little faith, wherefore didst thou doubt?
MATT|14|32|And when they were come into the ship, the wind ceased.
MATT|14|33|Then they that were in the ship came and worshipped him, saying, Of a truth thou art the Son of God.
MATT|14|34|And when they were gone over, they came into the land of Gennesaret.
MATT|14|35|And when the men of that place had knowledge of him, they sent out into all that country round about, and brought unto him all that were diseased;
MATT|14|36|And besought him that they might only touch the hem of his garment: and as many as touched were made perfectly whole.
MATT|15|1|Then came to Jesus scribes and Pharisees, which were of Jerusalem, saying,
MATT|15|2|Why do thy disciples transgress the tradition of the elders? for they wash not their hands when they eat bread.
MATT|15|3|But he answered and said unto them, Why do ye also transgress the commandment of God by your tradition?
MATT|15|4|For God commanded, saying, Honour thy father and mother: and, He that curseth father or mother, let him die the death.
MATT|15|5|But ye say, Whosoever shall say to his father or his mother, It is a gift, by whatsoever thou mightest be profited by me;
MATT|15|6|And honour not his father or his mother, he shall be free. Thus have ye made the commandment of God of none effect by your tradition.
MATT|15|7|Ye hypocrites, well did Esaias prophesy of you, saying,
MATT|15|8|This people draweth nigh unto me with their mouth, and honoureth me with their lips; but their heart is far from me.
MATT|15|9|But in vain they do worship me, teaching for doctrines the commandments of men.
MATT|15|10|And he called the multitude, and said unto them, Hear, and understand:
MATT|15|11|Not that which goeth into the mouth defileth a man; but that which cometh out of the mouth, this defileth a man.
MATT|15|12|Then came his disciples, and said unto him, Knowest thou that the Pharisees were offended, after they heard this saying?
MATT|15|13|But he answered and said, Every plant, which my heavenly Father hath not planted, shall be rooted up.
MATT|15|14|Let them alone: they be blind leaders of the blind. And if the blind lead the blind, both shall fall into the ditch.
MATT|15|15|Then answered Peter and said unto him, Declare unto us this parable.
MATT|15|16|And Jesus said, Are ye also yet without understanding?
MATT|15|17|Do not ye yet understand, that whatsoever entereth in at the mouth goeth into the belly, and is cast out into the draught?
MATT|15|18|But those things which proceed out of the mouth come forth from the heart; and they defile the man.
MATT|15|19|For out of the heart proceed evil thoughts, murders, adulteries, fornications, thefts, false witness, blasphemies:
MATT|15|20|These are the things which defile a man: but to eat with unwashen hands defileth not a man.
MATT|15|21|Then Jesus went thence, and departed into the coasts of Tyre and Sidon.
MATT|15|22|And, behold, a woman of Canaan came out of the same coasts, and cried unto him, saying, Have mercy on me, O Lord, thou son of David; my daughter is grievously vexed with a devil.
MATT|15|23|But he answered her not a word. And his disciples came and besought him, saying, Send her away; for she crieth after us.
MATT|15|24|But he answered and said, I am not sent but unto the lost sheep of the house of Israel.
MATT|15|25|Then came she and worshipped him, saying, Lord, help me.
MATT|15|26|But he answered and said, It is not meet to take the children's bread, and to cast it to dogs.
MATT|15|27|And she said, Truth, Lord: yet the dogs eat of the crumbs which fall from their masters' table.
MATT|15|28|Then Jesus answered and said unto her, O woman, great is thy faith: be it unto thee even as thou wilt. And her daughter was made whole from that very hour.
MATT|15|29|And Jesus departed from thence, and came nigh unto the sea of Galilee; and went up into a mountain, and sat down there.
MATT|15|30|And great multitudes came unto him, having with them those that were lame, blind, dumb, maimed, and many others, and cast them down at Jesus' feet; and he healed them:
MATT|15|31|Insomuch that the multitude wondered, when they saw the dumb to speak, the maimed to be whole, the lame to walk, and the blind to see: and they glorified the God of Israel.
MATT|15|32|Then Jesus called his disciples unto him, and said, I have compassion on the multitude, because they continue with me now three days, and have nothing to eat: and I will not send them away fasting, lest they faint in the way.
MATT|15|33|And his disciples say unto him, Whence should we have so much bread in the wilderness, as to fill so great a multitude?
MATT|15|34|And Jesus saith unto them, How many loaves have ye? And they said, Seven, and a few little fishes.
MATT|15|35|And he commanded the multitude to sit down on the ground.
MATT|15|36|And he took the seven loaves and the fishes, and gave thanks, and brake them, and gave to his disciples, and the disciples to the multitude.
MATT|15|37|And they did all eat, and were filled: and they took up of the broken meat that was left seven baskets full.
MATT|15|38|And they that did eat were four thousand men, beside women and children.
MATT|15|39|And he sent away the multitude, and took ship, and came into the coasts of Magdala.
MATT|16|1|The Pharisees also with the Sadducees came, and tempting desired him that he would shew them a sign from heaven.
MATT|16|2|He answered and said unto them, When it is evening, ye say, It will be fair weather: for the sky is red.
MATT|16|3|And in the morning, It will be foul weather to day: for the sky is red and lowering. O ye hypocrites, ye can discern the face of the sky; but can ye not discern the signs of the times?
MATT|16|4|A wicked and adulterous generation seeketh after a sign; and there shall no sign be given unto it, but the sign of the prophet Jonas. And he left them, and departed.
MATT|16|5|And when his disciples were come to the other side, they had forgotten to take bread.
MATT|16|6|Then Jesus said unto them, Take heed and beware of the leaven of the Pharisees and of the Sadducees.
MATT|16|7|And they reasoned among themselves, saying, It is because we have taken no bread.
MATT|16|8|Which when Jesus perceived, he said unto them, O ye of little faith, why reason ye among yourselves, because ye have brought no bread?
MATT|16|9|Do ye not yet understand, neither remember the five loaves of the five thousand, and how many baskets ye took up?
MATT|16|10|Neither the seven loaves of the four thousand, and how many baskets ye took up?
MATT|16|11|How is it that ye do not understand that I spake it not to you concerning bread, that ye should beware of the leaven of the Pharisees and of the Sadducees?
MATT|16|12|Then understood they how that he bade them not beware of the leaven of bread, but of the doctrine of the Pharisees and of the Sadducees.
MATT|16|13|When Jesus came into the coasts of Caesarea Philippi, he asked his disciples, saying, Whom do men say that I the Son of man am?
MATT|16|14|And they said, Some say that thou art John the Baptist: some, Elias; and others, Jeremias, or one of the prophets.
MATT|16|15|He saith unto them, But whom say ye that I am?
MATT|16|16|And Simon Peter answered and said, Thou art the Christ, the Son of the living God.
MATT|16|17|And Jesus answered and said unto him, Blessed art thou, Simon Barjona: for flesh and blood hath not revealed it unto thee, but my Father which is in heaven.
MATT|16|18|And I say also unto thee, That thou art Peter, and upon this rock I will build my church; and the gates of hell shall not prevail against it.
MATT|16|19|And I will give unto thee the keys of the kingdom of heaven: and whatsoever thou shalt bind on earth shall be bound in heaven: and whatsoever thou shalt loose on earth shall be loosed in heaven.
MATT|16|20|Then charged he his disciples that they should tell no man that he was Jesus the Christ.
MATT|16|21|From that time forth began Jesus to shew unto his disciples, how that he must go unto Jerusalem, and suffer many things of the elders and chief priests and scribes, and be killed, and be raised again the third day.
MATT|16|22|Then Peter took him, and began to rebuke him, saying, Be it far from thee, Lord: this shall not be unto thee.
MATT|16|23|But he turned, and said unto Peter, Get thee behind me, Satan: thou art an offence unto me: for thou savourest not the things that be of God, but those that be of men.
MATT|16|24|Then said Jesus unto his disciples, If any man will come after me, let him deny himself, and take up his cross, and follow me.
MATT|16|25|For whosoever will save his life shall lose it: and whosoever will lose his life for my sake shall find it.
MATT|16|26|For what is a man profited, if he shall gain the whole world, and lose his own soul? or what shall a man give in exchange for his soul?
MATT|16|27|For the Son of man shall come in the glory of his Father with his angels; and then he shall reward every man according to his works.
MATT|16|28|Verily I say unto you, There be some standing here, which shall not taste of death, till they see the Son of man coming in his kingdom.
MATT|17|1|And after six days Jesus taketh Peter, James, and John his brother, and bringeth them up into an high mountain apart,
MATT|17|2|And was transfigured before them: and his face did shine as the sun, and his raiment was white as the light.
MATT|17|3|And, behold, there appeared unto them Moses and Elias talking with him.
MATT|17|4|Then answered Peter, and said unto Jesus, Lord, it is good for us to be here: if thou wilt, let us make here three tabernacles; one for thee, and one for Moses, and one for Elias.
MATT|17|5|While he yet spake, behold, a bright cloud overshadowed them: and behold a voice out of the cloud, which said, This is my beloved Son, in whom I am well pleased; hear ye him.
MATT|17|6|And when the disciples heard it, they fell on their face, and were sore afraid.
MATT|17|7|And Jesus came and touched them, and said, Arise, and be not afraid.
MATT|17|8|And when they had lifted up their eyes, they saw no man, save Jesus only.
MATT|17|9|And as they came down from the mountain, Jesus charged them, saying, Tell the vision to no man, until the Son of man be risen again from the dead.
MATT|17|10|And his disciples asked him, saying, Why then say the scribes that Elias must first come?
MATT|17|11|And Jesus answered and said unto them, Elias truly shall first come, and restore all things.
MATT|17|12|But I say unto you, That Elias is come already, and they knew him not, but have done unto him whatsoever they listed. Likewise shall also the Son of man suffer of them.
MATT|17|13|Then the disciples understood that he spake unto them of John the Baptist.
MATT|17|14|And when they were come to the multitude, there came to him a certain man, kneeling down to him, and saying,
MATT|17|15|Lord, have mercy on my son: for he is lunatick, and sore vexed: for ofttimes he falleth into the fire, and oft into the water.
MATT|17|16|And I brought him to thy disciples, and they could not cure him.
MATT|17|17|Then Jesus answered and said, O faithless and perverse generation, how long shall I be with you? how long shall I suffer you? bring him hither to me.
MATT|17|18|And Jesus rebuked the devil; and he departed out of him: and the child was cured from that very hour.
MATT|17|19|Then came the disciples to Jesus apart, and said, Why could not we cast him out?
MATT|17|20|And Jesus said unto them, Because of your unbelief: for verily I say unto you, If ye have faith as a grain of mustard seed, ye shall say unto this mountain, Remove hence to yonder place; and it shall remove; and nothing shall be impossible unto you.
MATT|17|21|Howbeit this kind goeth not out but by prayer and fasting.
MATT|17|22|And while they abode in Galilee, Jesus said unto them, The Son of man shall be betrayed into the hands of men:
MATT|17|23|And they shall kill him, and the third day he shall be raised again. And they were exceeding sorry.
MATT|17|24|And when they were come to Capernaum, they that received tribute money came to Peter, and said, Doth not your master pay tribute?
MATT|17|25|He saith, Yes. And when he was come into the house, Jesus prevented him, saying, What thinkest thou, Simon? of whom do the kings of the earth take custom or tribute? of their own children, or of strangers?
MATT|17|26|Peter saith unto him, Of strangers. Jesus saith unto him, Then are the children free.
MATT|17|27|Notwithstanding, lest we should offend them, go thou to the sea, and cast an hook, and take up the fish that first cometh up; and when thou hast opened his mouth, thou shalt find a piece of money: that take, and give unto them for me and thee.
MATT|18|1|At the same time came the disciples unto Jesus, saying, Who is the greatest in the kingdom of heaven?
MATT|18|2|And Jesus called a little child unto him, and set him in the midst of them,
MATT|18|3|And said, Verily I say unto you, Except ye be converted, and become as little children, ye shall not enter into the kingdom of heaven.
MATT|18|4|Whosoever therefore shall humble himself as this little child, the same is greatest in the kingdom of heaven.
MATT|18|5|And whoso shall receive one such little child in my name receiveth me.
MATT|18|6|But whoso shall offend one of these little ones which believe in me, it were better for him that a millstone were hanged about his neck, and that he were drowned in the depth of the sea.
MATT|18|7|Woe unto the world because of offences! for it must needs be that offences come; but woe to that man by whom the offence cometh!
MATT|18|8|Wherefore if thy hand or thy foot offend thee, cut them off, and cast them from thee: it is better for thee to enter into life halt or maimed, rather than having two hands or two feet to be cast into everlasting fire.
MATT|18|9|And if thine eye offend thee, pluck it out, and cast it from thee: it is better for thee to enter into life with one eye, rather than having two eyes to be cast into hell fire.
MATT|18|10|Take heed that ye despise not one of these little ones; for I say unto you, That in heaven their angels do always behold the face of my Father which is in heaven.
MATT|18|11|For the Son of man is come to save that which was lost.
MATT|18|12|How think ye? if a man have an hundred sheep, and one of them be gone astray, doth he not leave the ninety and nine, and goeth into the mountains, and seeketh that which is gone astray?
MATT|18|13|And if so be that he find it, verily I say unto you, he rejoiceth more of that sheep, than of the ninety and nine which went not astray.
MATT|18|14|Even so it is not the will of your Father which is in heaven, that one of these little ones should perish.
MATT|18|15|Moreover if thy brother shall trespass against thee, go and tell him his fault between thee and him alone: if he shall hear thee, thou hast gained thy brother.
MATT|18|16|But if he will not hear thee, then take with thee one or two more, that in the mouth of two or three witnesses every word may be established.
MATT|18|17|And if he shall neglect to hear them, tell it unto the church: but if he neglect to hear the church, let him be unto thee as an heathen man and a publican.
MATT|18|18|Verily I say unto you, Whatsoever ye shall bind on earth shall be bound in heaven: and whatsoever ye shall loose on earth shall be loosed in heaven.
MATT|18|19|Again I say unto you, That if two of you shall agree on earth as touching any thing that they shall ask, it shall be done for them of my Father which is in heaven.
MATT|18|20|For where two or three are gathered together in my name, there am I in the midst of them.
MATT|18|21|Then came Peter to him, and said, Lord, how oft shall my brother sin against me, and I forgive him? till seven times?
MATT|18|22|Jesus saith unto him, I say not unto thee, Until seven times: but, Until seventy times seven.
MATT|18|23|Therefore is the kingdom of heaven likened unto a certain king, which would take account of his servants.
MATT|18|24|And when he had begun to reckon, one was brought unto him, which owed him ten thousand talents.
MATT|18|25|But forasmuch as he had not to pay, his lord commanded him to be sold, and his wife, and children, and all that he had, and payment to be made.
MATT|18|26|The servant therefore fell down, and worshipped him, saying, Lord, have patience with me, and I will pay thee all.
MATT|18|27|Then the lord of that servant was moved with compassion, and loosed him, and forgave him the debt.
MATT|18|28|But the same servant went out, and found one of his fellowservants, which owed him an hundred pence: and he laid hands on him, and took him by the throat, saying, Pay me that thou owest.
MATT|18|29|And his fellowservant fell down at his feet, and besought him, saying, Have patience with me, and I will pay thee all.
MATT|18|30|And he would not: but went and cast him into prison, till he should pay the debt.
MATT|18|31|So when his fellowservants saw what was done, they were very sorry, and came and told unto their lord all that was done.
MATT|18|32|Then his lord, after that he had called him, said unto him, O thou wicked servant, I forgave thee all that debt, because thou desiredst me:
MATT|18|33|Shouldest not thou also have had compassion on thy fellowservant, even as I had pity on thee?
MATT|18|34|And his lord was wroth, and delivered him to the tormentors, till he should pay all that was due unto him.
MATT|18|35|So likewise shall my heavenly Father do also unto you, if ye from your hearts forgive not every one his brother their trespasses.
MATT|19|1|And it came to pass, that when Jesus had finished these sayings, he departed from Galilee, and came into the coasts of Judaea beyond Jordan;
MATT|19|2|And great multitudes followed him; and he healed them there.
MATT|19|3|The Pharisees also came unto him, tempting him, and saying unto him, Is it lawful for a man to put away his wife for every cause?
MATT|19|4|And he answered and said unto them, Have ye not read, that he which made them at the beginning made them male and female,
MATT|19|5|And said, For this cause shall a man leave father and mother, and shall cleave to his wife: and they twain shall be one flesh?
MATT|19|6|Wherefore they are no more twain, but one flesh. What therefore God hath joined together, let not man put asunder.
MATT|19|7|They say unto him, Why did Moses then command to give a writing of divorcement, and to put her away?
MATT|19|8|He saith unto them, Moses because of the hardness of your hearts suffered you to put away your wives: but from the beginning it was not so.
MATT|19|9|And I say unto you, Whosoever shall put away his wife, except it be for fornication, and shall marry another, committeth adultery: and whoso marrieth her which is put away doth commit adultery.
MATT|19|10|His disciples say unto him, If the case of the man be so with his wife, it is not good to marry.
MATT|19|11|But he said unto them, All men cannot receive this saying, save they to whom it is given.
MATT|19|12|For there are some eunuchs, which were so born from their mother's womb: and there are some eunuchs, which were made eunuchs of men: and there be eunuchs, which have made themselves eunuchs for the kingdom of heaven's sake. He that is able to receive it, let him receive it.
MATT|19|13|Then were there brought unto him little children, that he should put his hands on them, and pray: and the disciples rebuked them.
MATT|19|14|But Jesus said, Suffer little children, and forbid them not, to come unto me: for of such is the kingdom of heaven.
MATT|19|15|And he laid his hands on them, and departed thence.
MATT|19|16|And, behold, one came and said unto him, Good Master, what good thing shall I do, that I may have eternal life?
MATT|19|17|And he said unto him, Why callest thou me good? there is none good but one, that is, God: but if thou wilt enter into life, keep the commandments.
MATT|19|18|He saith unto him, Which? Jesus said, Thou shalt do no murder, Thou shalt not commit adultery, Thou shalt not steal, Thou shalt not bear false witness,
MATT|19|19|Honour thy father and thy mother: and, Thou shalt love thy neighbour as thyself.
MATT|19|20|The young man saith unto him, All these things have I kept from my youth up: what lack I yet?
MATT|19|21|Jesus said unto him, If thou wilt be perfect, go and sell that thou hast, and give to the poor, and thou shalt have treasure in heaven: and come and follow me.
MATT|19|22|But when the young man heard that saying, he went away sorrowful: for he had great possessions.
MATT|19|23|Then said Jesus unto his disciples, Verily I say unto you, That a rich man shall hardly enter into the kingdom of heaven.
MATT|19|24|And again I say unto you, It is easier for a camel to go through the eye of a needle, than for a rich man to enter into the kingdom of God.
MATT|19|25|When his disciples heard it, they were exceedingly amazed, saying, Who then can be saved?
MATT|19|26|But Jesus beheld them, and said unto them, With men this is impossible; but with God all things are possible.
MATT|19|27|Then answered Peter and said unto him, Behold, we have forsaken all, and followed thee; what shall we have therefore?
MATT|19|28|And Jesus said unto them, Verily I say unto you, That ye which have followed me, in the regeneration when the Son of man shall sit in the throne of his glory, ye also shall sit upon twelve thrones, judging the twelve tribes of Israel.
MATT|19|29|And every one that hath forsaken houses, or brethren, or sisters, or father, or mother, or wife, or children, or lands, for my name's sake, shall receive an hundredfold, and shall inherit everlasting life.
MATT|19|30|But many that are first shall be last; and the last shall be first.
MATT|20|1|For the kingdom of heaven is like unto a man that is an householder, which went out early in the morning to hire labourers into his vineyard.
MATT|20|2|And when he had agreed with the labourers for a penny a day, he sent them into his vineyard.
MATT|20|3|And he went out about the third hour, and saw others standing idle in the marketplace,
MATT|20|4|And said unto them; Go ye also into the vineyard, and whatsoever is right I will give you. And they went their way.
MATT|20|5|Again he went out about the sixth and ninth hour, and did likewise.
MATT|20|6|And about the eleventh hour he went out, and found others standing idle, and saith unto them, Why stand ye here all the day idle?
MATT|20|7|They say unto him, Because no man hath hired us. He saith unto them, Go ye also into the vineyard; and whatsoever is right, that shall ye receive.
MATT|20|8|So when even was come, the lord of the vineyard saith unto his steward, Call the labourers, and give them their hire, beginning from the last unto the first.
MATT|20|9|And when they came that were hired about the eleventh hour, they received every man a penny.
MATT|20|10|But when the first came, they supposed that they should have received more; and they likewise received every man a penny.
MATT|20|11|And when they had received it, they murmured against the goodman of the house,
MATT|20|12|Saying, These last have wrought but one hour, and thou hast made them equal unto us, which have borne the burden and heat of the day.
MATT|20|13|But he answered one of them, and said, Friend, I do thee no wrong: didst not thou agree with me for a penny?
MATT|20|14|Take that thine is, and go thy way: I will give unto this last, even as unto thee.
MATT|20|15|Is it not lawful for me to do what I will with mine own? Is thine eye evil, because I am good?
MATT|20|16|So the last shall be first, and the first last: for many be called, but few chosen.
MATT|20|17|And Jesus going up to Jerusalem took the twelve disciples apart in the way, and said unto them,
MATT|20|18|Behold, we go up to Jerusalem; and the Son of man shall be betrayed unto the chief priests and unto the scribes, and they shall condemn him to death,
MATT|20|19|And shall deliver him to the Gentiles to mock, and to scourge, and to crucify him: and the third day he shall rise again.
MATT|20|20|Then came to him the mother of Zebedees children with her sons, worshipping him, and desiring a certain thing of him.
MATT|20|21|And he said unto her, What wilt thou? She saith unto him, Grant that these my two sons may sit, the one on thy right hand, and the other on the left, in thy kingdom.
MATT|20|22|But Jesus answered and said, Ye know not what ye ask. Are ye able to drink of the cup that I shall drink of, and to be baptized with the baptism that I am baptized with? They say unto him, We are able.
MATT|20|23|And he saith unto them, Ye shall drink indeed of my cup, and be baptized with the baptism that I am baptized with: but to sit on my right hand, and on my left, is not mine to give, but it shall be given to them for whom it is prepared of my Father.
MATT|20|24|And when the ten heard it, they were moved with indignation against the two brethren.
MATT|20|25|But Jesus called them unto him, and said, Ye know that the princes of the Gentiles exercise dominion over them, and they that are great exercise authority upon them.
MATT|20|26|But it shall not be so among you: but whosoever will be great among you, let him be your minister;
MATT|20|27|And whosoever will be chief among you, let him be your servant:
MATT|20|28|Even as the Son of man came not to be ministered unto, but to minister, and to give his life a ransom for many.
MATT|20|29|And as they departed from Jericho, a great multitude followed him.
MATT|20|30|And, behold, two blind men sitting by the way side, when they heard that Jesus passed by, cried out, saying, Have mercy on us, O Lord, thou son of David.
MATT|20|31|And the multitude rebuked them, because they should hold their peace: but they cried the more, saying, Have mercy on us, O Lord, thou son of David.
MATT|20|32|And Jesus stood still, and called them, and said, What will ye that I shall do unto you?
MATT|20|33|They say unto him, Lord, that our eyes may be opened.
MATT|20|34|So Jesus had compassion on them, and touched their eyes: and immediately their eyes received sight, and they followed him.
MATT|21|1|And when they drew nigh unto Jerusalem, and were come to Bethphage, unto the mount of Olives, then sent Jesus two disciples,
MATT|21|2|Saying unto them, Go into the village over against you, and straightway ye shall find an ass tied, and a colt with her: loose them, and bring them unto me.
MATT|21|3|And if any man say ought unto you, ye shall say, The Lord hath need of them; and straightway he will send them.
MATT|21|4|All this was done, that it might be fulfilled which was spoken by the prophet, saying,
MATT|21|5|Tell ye the daughter of Sion, Behold, thy King cometh unto thee, meek, and sitting upon an ass, and a colt the foal of an ass.
MATT|21|6|And the disciples went, and did as Jesus commanded them,
MATT|21|7|And brought the ass, and the colt, and put on them their clothes, and they set him thereon.
MATT|21|8|And a very great multitude spread their garments in the way; others cut down branches from the trees, and strawed them in the way.
MATT|21|9|And the multitudes that went before, and that followed, cried, saying, Hosanna to the son of David: Blessed is he that cometh in the name of the Lord; Hosanna in the highest.
MATT|21|10|And when he was come into Jerusalem, all the city was moved, saying, Who is this?
MATT|21|11|And the multitude said, This is Jesus the prophet of Nazareth of Galilee.
MATT|21|12|And Jesus went into the temple of God, and cast out all them that sold and bought in the temple, and overthrew the tables of the moneychangers, and the seats of them that sold doves,
MATT|21|13|And said unto them, It is written, My house shall be called the house of prayer; but ye have made it a den of thieves.
MATT|21|14|And the blind and the lame came to him in the temple; and he healed them.
MATT|21|15|And when the chief priests and scribes saw the wonderful things that he did, and the children crying in the temple, and saying, Hosanna to the son of David; they were sore displeased,
MATT|21|16|And said unto him, Hearest thou what these say? And Jesus saith unto them, Yea; have ye never read, Out of the mouth of babes and sucklings thou hast perfected praise?
MATT|21|17|And he left them, and went out of the city into Bethany; and he lodged there.
MATT|21|18|Now in the morning as he returned into the city, he hungered.
MATT|21|19|And when he saw a fig tree in the way, he came to it, and found nothing thereon, but leaves only, and said unto it, Let no fruit grow on thee henceforward for ever. And presently the fig tree withered away.
MATT|21|20|And when the disciples saw it, they marvelled, saying, How soon is the fig tree withered away!
MATT|21|21|Jesus answered and said unto them, Verily I say unto you, If ye have faith, and doubt not, ye shall not only do this which is done to the fig tree, but also if ye shall say unto this mountain, Be thou removed, and be thou cast into the sea; it shall be done.
MATT|21|22|And all things, whatsoever ye shall ask in prayer, believing, ye shall receive.
MATT|21|23|And when he was come into the temple, the chief priests and the elders of the people came unto him as he was teaching, and said, By what authority doest thou these things? and who gave thee this authority?
MATT|21|24|And Jesus answered and said unto them, I also will ask you one thing, which if ye tell me, I in like wise will tell you by what authority I do these things.
MATT|21|25|The baptism of John, whence was it? from heaven, or of men? And they reasoned with themselves, saying, If we shall say, From heaven; he will say unto us, Why did ye not then believe him?
MATT|21|26|But if we shall say, Of men; we fear the people; for all hold John as a prophet.
MATT|21|27|And they answered Jesus, and said, We cannot tell. And he said unto them, Neither tell I you by what authority I do these things.
MATT|21|28|But what think ye? A certain man had two sons; and he came to the first, and said, Son, go work to day in my vineyard.
MATT|21|29|He answered and said, I will not: but afterward he repented, and went.
MATT|21|30|And he came to the second, and said likewise. And he answered and said, I go, sir: and went not.
MATT|21|31|Whether of them twain did the will of his father? They say unto him, The first. Jesus saith unto them, Verily I say unto you, That the publicans and the harlots go into the kingdom of God before you.
MATT|21|32|For John came unto you in the way of righteousness, and ye believed him not: but the publicans and the harlots believed him: and ye, when ye had seen it, repented not afterward, that ye might believe him.
MATT|21|33|Hear another parable: There was a certain householder, which planted a vineyard, and hedged it round about, and digged a winepress in it, and built a tower, and let it out to husbandmen, and went into a far country:
MATT|21|34|And when the time of the fruit drew near, he sent his servants to the husbandmen, that they might receive the fruits of it.
MATT|21|35|And the husbandmen took his servants, and beat one, and killed another, and stoned another.
MATT|21|36|Again, he sent other servants more than the first: and they did unto them likewise.
MATT|21|37|But last of all he sent unto them his son, saying, They will reverence my son.
MATT|21|38|But when the husbandmen saw the son, they said among themselves, This is the heir; come, let us kill him, and let us seize on his inheritance.
MATT|21|39|And they caught him, and cast him out of the vineyard, and slew him.
MATT|21|40|When the lord therefore of the vineyard cometh, what will he do unto those husbandmen?
MATT|21|41|They say unto him, He will miserably destroy those wicked men, and will let out his vineyard unto other husbandmen, which shall render him the fruits in their seasons.
MATT|21|42|Jesus saith unto them, Did ye never read in the scriptures, The stone which the builders rejected, the same is become the head of the corner: this is the Lord's doing, and it is marvellous in our eyes?
MATT|21|43|Therefore say I unto you, The kingdom of God shall be taken from you, and given to a nation bringing forth the fruits thereof.
MATT|21|44|And whosoever shall fall on this stone shall be broken: but on whomsoever it shall fall, it will grind him to powder.
MATT|21|45|And when the chief priests and Pharisees had heard his parables, they perceived that he spake of them.
MATT|21|46|But when they sought to lay hands on him, they feared the multitude, because they took him for a prophet.
MATT|22|1|And Jesus answered and spake unto them again by parables, and said,
MATT|22|2|The kingdom of heaven is like unto a certain king, which made a marriage for his son,
MATT|22|3|And sent forth his servants to call them that were bidden to the wedding: and they would not come.
MATT|22|4|Again, he sent forth other servants, saying, Tell them which are bidden, Behold, I have prepared my dinner: my oxen and my fatlings are killed, and all things are ready: come unto the marriage.
MATT|22|5|But they made light of it, and went their ways, one to his farm, another to his merchandise:
MATT|22|6|And the remnant took his servants, and entreated them spitefully, and slew them.
MATT|22|7|But when the king heard thereof, he was wroth: and he sent forth his armies, and destroyed those murderers, and burned up their city.
MATT|22|8|Then saith he to his servants, The wedding is ready, but they which were bidden were not worthy.
MATT|22|9|Go ye therefore into the highways, and as many as ye shall find, bid to the marriage.
MATT|22|10|So those servants went out into the highways, and gathered together all as many as they found, both bad and good: and the wedding was furnished with guests.
MATT|22|11|And when the king came in to see the guests, he saw there a man which had not on a wedding garment:
MATT|22|12|And he saith unto him, Friend, how camest thou in hither not having a wedding garment? And he was speechless.
MATT|22|13|Then said the king to the servants, Bind him hand and foot, and take him away, and cast him into outer darkness, there shall be weeping and gnashing of teeth.
MATT|22|14|For many are called, but few are chosen.
MATT|22|15|Then went the Pharisees, and took counsel how they might entangle him in his talk.
MATT|22|16|And they sent out unto him their disciples with the Herodians, saying, Master, we know that thou art true, and teachest the way of God in truth, neither carest thou for any man: for thou regardest not the person of men.
MATT|22|17|Tell us therefore, What thinkest thou? Is it lawful to give tribute unto Caesar, or not?
MATT|22|18|But Jesus perceived their wickedness, and said, Why tempt ye me, ye hypocrites?
MATT|22|19|Shew me the tribute money. And they brought unto him a penny.
MATT|22|20|And he saith unto them, Whose is this image and superscription?
MATT|22|21|They say unto him, Caesar's. Then saith he unto them, Render therefore unto Caesar the things which are Caesar's; and unto God the things that are God's.
MATT|22|22|When they had heard these words, they marvelled, and left him, and went their way.
MATT|22|23|The same day came to him the Sadducees, which say that there is no resurrection, and asked him,
MATT|22|24|Saying, Master, Moses said, If a man die, having no children, his brother shall marry his wife, and raise up seed unto his brother.
MATT|22|25|Now there were with us seven brethren: and the first, when he had married a wife, deceased, and, having no issue, left his wife unto his brother:
MATT|22|26|Likewise the second also, and the third, unto the seventh.
MATT|22|27|And last of all the woman died also.
MATT|22|28|Therefore in the resurrection whose wife shall she be of the seven? for they all had her.
MATT|22|29|Jesus answered and said unto them, Ye do err, not knowing the scriptures, nor the power of God.
MATT|22|30|For in the resurrection they neither marry, nor are given in marriage, but are as the angels of God in heaven.
MATT|22|31|But as touching the resurrection of the dead, have ye not read that which was spoken unto you by God, saying,
MATT|22|32|I am the God of Abraham, and the God of Isaac, and the God of Jacob? God is not the God of the dead, but of the living.
MATT|22|33|And when the multitude heard this, they were astonished at his doctrine.
MATT|22|34|But when the Pharisees had heard that he had put the Sadducees to silence, they were gathered together.
MATT|22|35|Then one of them, which was a lawyer, asked him a question, tempting him, and saying,
MATT|22|36|Master, which is the great commandment in the law?
MATT|22|37|Jesus said unto him, Thou shalt love the Lord thy God with all thy heart, and with all thy soul, and with all thy mind.
MATT|22|38|This is the first and great commandment.
MATT|22|39|And the second is like unto it, Thou shalt love thy neighbour as thyself.
MATT|22|40|On these two commandments hang all the law and the prophets.
MATT|22|41|While the Pharisees were gathered together, Jesus asked them,
MATT|22|42|Saying, What think ye of Christ? whose son is he? They say unto him, The son of David.
MATT|22|43|He saith unto them, How then doth David in spirit call him Lord, saying,
MATT|22|44|The LORD said unto my Lord, Sit thou on my right hand, till I make thine enemies thy footstool?
MATT|22|45|If David then call him Lord, how is he his son?
MATT|22|46|And no man was able to answer him a word, neither durst any man from that day forth ask him any more questions.
MATT|23|1|Then spake Jesus to the multitude, and to his disciples,
MATT|23|2|Saying The scribes and the Pharisees sit in Moses' seat:
MATT|23|3|All therefore whatsoever they bid you observe, that observe and do; but do not ye after their works: for they say, and do not.
MATT|23|4|For they bind heavy burdens and grievous to be borne, and lay them on men's shoulders; but they themselves will not move them with one of their fingers.
MATT|23|5|But all their works they do for to be seen of men: they make broad their phylacteries, and enlarge the borders of their garments,
MATT|23|6|And love the uppermost rooms at feasts, and the chief seats in the synagogues,
MATT|23|7|And greetings in the markets, and to be called of men, Rabbi, Rabbi.
MATT|23|8|But be not ye called Rabbi: for one is your Master, even Christ; and all ye are brethren.
MATT|23|9|And call no man your father upon the earth: for one is your Father, which is in heaven.
MATT|23|10|Neither be ye called masters: for one is your Master, even Christ.
MATT|23|11|But he that is greatest among you shall be your servant.
MATT|23|12|And whosoever shall exalt himself shall be abased; and he that shall humble himself shall be exalted.
MATT|23|13|But woe unto you, scribes and Pharisees, hypocrites! for ye shut up the kingdom of heaven against men: for ye neither go in yourselves, neither suffer ye them that are entering to go in.
MATT|23|14|Woe unto you, scribes and Pharisees, hypocrites! for ye devour widows' houses, and for a pretence make long prayer: therefore ye shall receive the greater damnation.
MATT|23|15|Woe unto you, scribes and Pharisees, hypocrites! for ye compass sea and land to make one proselyte, and when he is made, ye make him twofold more the child of hell than yourselves.
MATT|23|16|Woe unto you, ye blind guides, which say, Whosoever shall swear by the temple, it is nothing; but whosoever shall swear by the gold of the temple, he is a debtor!
MATT|23|17|Ye fools and blind: for whether is greater, the gold, or the temple that sanctifieth the gold?
MATT|23|18|And, Whosoever shall swear by the altar, it is nothing; but whosoever sweareth by the gift that is upon it, he is guilty.
MATT|23|19|Ye fools and blind: for whether is greater, the gift, or the altar that sanctifieth the gift?
MATT|23|20|Whoso therefore shall swear by the altar, sweareth by it, and by all things thereon.
MATT|23|21|And whoso shall swear by the temple, sweareth by it, and by him that dwelleth therein.
MATT|23|22|And he that shall swear by heaven, sweareth by the throne of God, and by him that sitteth thereon.
MATT|23|23|Woe unto you, scribes and Pharisees, hypocrites! for ye pay tithe of mint and anise and cummin, and have omitted the weightier matters of the law, judgment, mercy, and faith: these ought ye to have done, and not to leave the other undone.
MATT|23|24|Ye blind guides, which strain at a gnat, and swallow a camel.
MATT|23|25|Woe unto you, scribes and Pharisees, hypocrites! for ye make clean the outside of the cup and of the platter, but within they are full of extortion and excess.
MATT|23|26|Thou blind Pharisee, cleanse first that which is within the cup and platter, that the outside of them may be clean also.
MATT|23|27|Woe unto you, scribes and Pharisees, hypocrites! for ye are like unto whited sepulchres, which indeed appear beautiful outward, but are within full of dead men's bones, and of all uncleanness.
MATT|23|28|Even so ye also outwardly appear righteous unto men, but within ye are full of hypocrisy and iniquity.
MATT|23|29|Woe unto you, scribes and Pharisees, hypocrites! because ye build the tombs of the prophets, and garnish the sepulchres of the righteous,
MATT|23|30|And say, If we had been in the days of our fathers, we would not have been partakers with them in the blood of the prophets.
MATT|23|31|Wherefore ye be witnesses unto yourselves, that ye are the children of them which killed the prophets.
MATT|23|32|Fill ye up then the measure of your fathers.
MATT|23|33|Ye serpents, ye generation of vipers, how can ye escape the damnation of hell?
MATT|23|34|Wherefore, behold, I send unto you prophets, and wise men, and scribes: and some of them ye shall kill and crucify; and some of them shall ye scourge in your synagogues, and persecute them from city to city:
MATT|23|35|That upon you may come all the righteous blood shed upon the earth, from the blood of righteous Abel unto the blood of Zacharias son of Barachias, whom ye slew between the temple and the altar.
MATT|23|36|Verily I say unto you, All these things shall come upon this generation.
MATT|23|37|O Jerusalem, Jerusalem, thou that killest the prophets, and stonest them which are sent unto thee, how often would I have gathered thy children together, even as a hen gathereth her chickens under her wings, and ye would not!
MATT|23|38|Behold, your house is left unto you desolate.
MATT|23|39|For I say unto you, Ye shall not see me henceforth, till ye shall say, Blessed is he that cometh in the name of the Lord.
MATT|24|1|And Jesus went out, and departed from the temple: and his disciples came to him for to shew him the buildings of the temple.
MATT|24|2|And Jesus said unto them, See ye not all these things? verily I say unto you, There shall not be left here one stone upon another, that shall not be thrown down.
MATT|24|3|And as he sat upon the mount of Olives, the disciples came unto him privately, saying, Tell us, when shall these things be? and what shall be the sign of thy coming, and of the end of the world?
MATT|24|4|And Jesus answered and said unto them, Take heed that no man deceive you.
MATT|24|5|For many shall come in my name, saying, I am Christ; and shall deceive many.
MATT|24|6|And ye shall hear of wars and rumours of wars: see that ye be not troubled: for all these things must come to pass, but the end is not yet.
MATT|24|7|For nation shall rise against nation, and kingdom against kingdom: and there shall be famines, and pestilences, and earthquakes, in divers places.
MATT|24|8|All these are the beginning of sorrows.
MATT|24|9|Then shall they deliver you up to be afflicted, and shall kill you: and ye shall be hated of all nations for my name's sake.
MATT|24|10|And then shall many be offended, and shall betray one another, and shall hate one another.
MATT|24|11|And many false prophets shall rise, and shall deceive many.
MATT|24|12|And because iniquity shall abound, the love of many shall wax cold.
MATT|24|13|But he that shall endure unto the end, the same shall be saved.
MATT|24|14|And this gospel of the kingdom shall be preached in all the world for a witness unto all nations; and then shall the end come.
MATT|24|15|When ye therefore shall see the abomination of desolation, spoken of by Daniel the prophet, stand in the holy place, (whoso readeth, let him understand:)
MATT|24|16|Then let them which be in Judaea flee into the mountains:
MATT|24|17|Let him which is on the housetop not come down to take any thing out of his house:
MATT|24|18|Neither let him which is in the field return back to take his clothes.
MATT|24|19|And woe unto them that are with child, and to them that give suck in those days!
MATT|24|20|But pray ye that your flight be not in the winter, neither on the sabbath day:
MATT|24|21|For then shall be great tribulation, such as was not since the beginning of the world to this time, no, nor ever shall be.
MATT|24|22|And except those days should be shortened, there should no flesh be saved: but for the elect's sake those days shall be shortened.
MATT|24|23|Then if any man shall say unto you, Lo, here is Christ, or there; believe it not.
MATT|24|24|For there shall arise false Christs, and false prophets, and shall shew great signs and wonders; insomuch that, if it were possible, they shall deceive the very elect.
MATT|24|25|Behold, I have told you before.
MATT|24|26|Wherefore if they shall say unto you, Behold, he is in the desert; go not forth: behold, he is in the secret chambers; believe it not.
MATT|24|27|For as the lightning cometh out of the east, and shineth even unto the west; so shall also the coming of the Son of man be.
MATT|24|28|For wheresoever the carcase is, there will the eagles be gathered together.
MATT|24|29|Immediately after the tribulation of those days shall the sun be darkened, and the moon shall not give her light, and the stars shall fall from heaven, and the powers of the heavens shall be shaken:
MATT|24|30|And then shall appear the sign of the Son of man in heaven: and then shall all the tribes of the earth mourn, and they shall see the Son of man coming in the clouds of heaven with power and great glory.
MATT|24|31|And he shall send his angels with a great sound of a trumpet, and they shall gather together his elect from the four winds, from one end of heaven to the other.
MATT|24|32|Now learn a parable of the fig tree; When his branch is yet tender, and putteth forth leaves, ye know that summer is nigh:
MATT|24|33|So likewise ye, when ye shall see all these things, know that it is near, even at the doors.
MATT|24|34|Verily I say unto you, This generation shall not pass, till all these things be fulfilled.
MATT|24|35|Heaven and earth shall pass away, but my words shall not pass away.
MATT|24|36|But of that day and hour knoweth no man, no, not the angels of heaven, but my Father only.
MATT|24|37|But as the days of Noe were, so shall also the coming of the Son of man be.
MATT|24|38|For as in the days that were before the flood they were eating and drinking, marrying and giving in marriage, until the day that Noe entered into the ark,
MATT|24|39|And knew not until the flood came, and took them all away; so shall also the coming of the Son of man be.
MATT|24|40|Then shall two be in the field; the one shall be taken, and the other left.
MATT|24|41|Two women shall be grinding at the mill; the one shall be taken, and the other left.
MATT|24|42|Watch therefore: for ye know not what hour your Lord doth come.
MATT|24|43|But know this, that if the goodman of the house had known in what watch the thief would come, he would have watched, and would not have suffered his house to be broken up.
MATT|24|44|Therefore be ye also ready: for in such an hour as ye think not the Son of man cometh.
MATT|24|45|Who then is a faithful and wise servant, whom his lord hath made ruler over his household, to give them meat in due season?
MATT|24|46|Blessed is that servant, whom his lord when he cometh shall find so doing.
MATT|24|47|Verily I say unto you, That he shall make him ruler over all his goods.
MATT|24|48|But and if that evil servant shall say in his heart, My lord delayeth his coming;
MATT|24|49|And shall begin to smite his fellowservants, and to eat and drink with the drunken;
MATT|24|50|The lord of that servant shall come in a day when he looketh not for him, and in an hour that he is not aware of,
MATT|24|51|And shall cut him asunder, and appoint him his portion with the hypocrites: there shall be weeping and gnashing of teeth.
MATT|25|1|Then shall the kingdom of heaven be likened unto ten virgins, which took their lamps, and went forth to meet the bridegroom.
MATT|25|2|And five of them were wise, and five were foolish.
MATT|25|3|They that were foolish took their lamps, and took no oil with them:
MATT|25|4|But the wise took oil in their vessels with their lamps.
MATT|25|5|While the bridegroom tarried, they all slumbered and slept.
MATT|25|6|And at midnight there was a cry made, Behold, the bridegroom cometh; go ye out to meet him.
MATT|25|7|Then all those virgins arose, and trimmed their lamps.
MATT|25|8|And the foolish said unto the wise, Give us of your oil; for our lamps are gone out.
MATT|25|9|But the wise answered, saying, Not so; lest there be not enough for us and you: but go ye rather to them that sell, and buy for yourselves.
MATT|25|10|And while they went to buy, the bridegroom came; and they that were ready went in with him to the marriage: and the door was shut.
MATT|25|11|Afterward came also the other virgins, saying, Lord, Lord, open to us.
MATT|25|12|But he answered and said, Verily I say unto you, I know you not.
MATT|25|13|Watch therefore, for ye know neither the day nor the hour wherein the Son of man cometh.
MATT|25|14|For the kingdom of heaven is as a man travelling into a far country, who called his own servants, and delivered unto them his goods.
MATT|25|15|And unto one he gave five talents, to another two, and to another one; to every man according to his several ability; and straightway took his journey.
MATT|25|16|Then he that had received the five talents went and traded with the same, and made them other five talents.
MATT|25|17|And likewise he that had received two, he also gained other two.
MATT|25|18|But he that had received one went and digged in the earth, and hid his lord's money.
MATT|25|19|After a long time the lord of those servants cometh, and reckoneth with them.
MATT|25|20|And so he that had received five talents came and brought other five talents, saying, Lord, thou deliveredst unto me five talents: behold, I have gained beside them five talents more.
MATT|25|21|His lord said unto him, Well done, thou good and faithful servant: thou hast been faithful over a few things, I will make thee ruler over many things: enter thou into the joy of thy lord.
MATT|25|22|He also that had received two talents came and said, Lord, thou deliveredst unto me two talents: behold, I have gained two other talents beside them.
MATT|25|23|His lord said unto him, Well done, good and faithful servant; thou hast been faithful over a few things, I will make thee ruler over many things: enter thou into the joy of thy lord.
MATT|25|24|Then he which had received the one talent came and said, Lord, I knew thee that thou art an hard man, reaping where thou hast not sown, and gathering where thou hast not strawed:
MATT|25|25|And I was afraid, and went and hid thy talent in the earth: lo, there thou hast that is thine.
MATT|25|26|His lord answered and said unto him, Thou wicked and slothful servant, thou knewest that I reap where I sowed not, and gather where I have not strawed:
MATT|25|27|Thou oughtest therefore to have put my money to the exchangers, and then at my coming I should have received mine own with usury.
MATT|25|28|Take therefore the talent from him, and give it unto him which hath ten talents.
MATT|25|29|For unto every one that hath shall be given, and he shall have abundance: but from him that hath not shall be taken away even that which he hath.
MATT|25|30|And cast ye the unprofitable servant into outer darkness: there shall be weeping and gnashing of teeth.
MATT|25|31|When the Son of man shall come in his glory, and all the holy angels with him, then shall he sit upon the throne of his glory:
MATT|25|32|And before him shall be gathered all nations: and he shall separate them one from another, as a shepherd divideth his sheep from the goats:
MATT|25|33|And he shall set the sheep on his right hand, but the goats on the left.
MATT|25|34|Then shall the King say unto them on his right hand, Come, ye blessed of my Father, inherit the kingdom prepared for you from the foundation of the world:
MATT|25|35|For I was an hungred, and ye gave me meat: I was thirsty, and ye gave me drink: I was a stranger, and ye took me in:
MATT|25|36|Naked, and ye clothed me: I was sick, and ye visited me: I was in prison, and ye came unto me.
MATT|25|37|Then shall the righteous answer him, saying, Lord, when saw we thee an hungred, and fed thee? or thirsty, and gave thee drink?
MATT|25|38|When saw we thee a stranger, and took thee in? or naked, and clothed thee?
MATT|25|39|Or when saw we thee sick, or in prison, and came unto thee?
MATT|25|40|And the King shall answer and say unto them, Verily I say unto you, Inasmuch as ye have done it unto one of the least of these my brethren, ye have done it unto me.
MATT|25|41|Then shall he say also unto them on the left hand, Depart from me, ye cursed, into everlasting fire, prepared for the devil and his angels:
MATT|25|42|For I was an hungred, and ye gave me no meat: I was thirsty, and ye gave me no drink:
MATT|25|43|I was a stranger, and ye took me not in: naked, and ye clothed me not: sick, and in prison, and ye visited me not.
MATT|25|44|Then shall they also answer him, saying, Lord, when saw we thee an hungred, or athirst, or a stranger, or naked, or sick, or in prison, and did not minister unto thee?
MATT|25|45|Then shall he answer them, saying, Verily I say unto you, Inasmuch as ye did it not to one of the least of these, ye did it not to me.
MATT|25|46|And these shall go away into everlasting punishment: but the righteous into life eternal.
MATT|26|1|And it came to pass, when Jesus had finished all these sayings, he said unto his disciples,
MATT|26|2|Ye know that after two days is the feast of the passover, and the Son of man is betrayed to be crucified.
MATT|26|3|Then assembled together the chief priests, and the scribes, and the elders of the people, unto the palace of the high priest, who was called Caiaphas,
MATT|26|4|And consulted that they might take Jesus by subtilty, and kill him.
MATT|26|5|But they said, Not on the feast day, lest there be an uproar among the people.
MATT|26|6|Now when Jesus was in Bethany, in the house of Simon the leper,
MATT|26|7|There came unto him a woman having an alabaster box of very precious ointment, and poured it on his head, as he sat at meat.
MATT|26|8|But when his disciples saw it, they had indignation, saying, To what purpose is this waste?
MATT|26|9|For this ointment might have been sold for much, and given to the poor.
MATT|26|10|When Jesus understood it, he said unto them, Why trouble ye the woman? for she hath wrought a good work upon me.
MATT|26|11|For ye have the poor always with you; but me ye have not always.
MATT|26|12|For in that she hath poured this ointment on my body, she did it for my burial.
MATT|26|13|Verily I say unto you, Wheresoever this gospel shall be preached in the whole world, there shall also this, that this woman hath done, be told for a memorial of her.
MATT|26|14|Then one of the twelve, called Judas Iscariot, went unto the chief priests,
MATT|26|15|And said unto them, What will ye give me, and I will deliver him unto you? And they covenanted with him for thirty pieces of silver.
MATT|26|16|And from that time he sought opportunity to betray him.
MATT|26|17|Now the first day of the feast of unleavened bread the disciples came to Jesus, saying unto him, Where wilt thou that we prepare for thee to eat the passover?
MATT|26|18|And he said, Go into the city to such a man, and say unto him, The Master saith, My time is at hand; I will keep the passover at thy house with my disciples.
MATT|26|19|And the disciples did as Jesus had appointed them; and they made ready the passover.
MATT|26|20|Now when the even was come, he sat down with the twelve.
MATT|26|21|And as they did eat, he said, Verily I say unto you, that one of you shall betray me.
MATT|26|22|And they were exceeding sorrowful, and began every one of them to say unto him, Lord, is it I?
MATT|26|23|And he answered and said, He that dippeth his hand with me in the dish, the same shall betray me.
MATT|26|24|The Son of man goeth as it is written of him: but woe unto that man by whom the Son of man is betrayed! it had been good for that man if he had not been born.
MATT|26|25|Then Judas, which betrayed him, answered and said, Master, is it I? He said unto him, Thou hast said.
MATT|26|26|And as they were eating, Jesus took bread, and blessed it, and brake it, and gave it to the disciples, and said, Take, eat; this is my body.
MATT|26|27|And he took the cup, and gave thanks, and gave it to them, saying, Drink ye all of it;
MATT|26|28|For this is my blood of the new testament, which is shed for many for the remission of sins.
MATT|26|29|But I say unto you, I will not drink henceforth of this fruit of the vine, until that day when I drink it new with you in my Father's kingdom.
MATT|26|30|And when they had sung an hymn, they went out into the mount of Olives.
MATT|26|31|Then saith Jesus unto them, All ye shall be offended because of me this night: for it is written, I will smite the shepherd, and the sheep of the flock shall be scattered abroad.
MATT|26|32|But after I am risen again, I will go before you into Galilee.
MATT|26|33|Peter answered and said unto him, Though all men shall be offended because of thee, yet will I never be offended.
MATT|26|34|Jesus said unto him, Verily I say unto thee, That this night, before the cock crow, thou shalt deny me thrice.
MATT|26|35|Peter said unto him, Though I should die with thee, yet will I not deny thee. Likewise also said all the disciples.
MATT|26|36|Then cometh Jesus with them unto a place called Gethsemane, and saith unto the disciples, Sit ye here, while I go and pray yonder.
MATT|26|37|And he took with him Peter and the two sons of Zebedee, and began to be sorrowful and very heavy.
MATT|26|38|Then saith he unto them, My soul is exceeding sorrowful, even unto death: tarry ye here, and watch with me.
MATT|26|39|And he went a little farther, and fell on his face, and prayed, saying, O my Father, if it be possible, let this cup pass from me: nevertheless not as I will, but as thou wilt.
MATT|26|40|And he cometh unto the disciples, and findeth them asleep, and saith unto Peter, What, could ye not watch with me one hour?
MATT|26|41|Watch and pray, that ye enter not into temptation: the spirit indeed is willing, but the flesh is weak.
MATT|26|42|He went away again the second time, and prayed, saying, O my Father, if this cup may not pass away from me, except I drink it, thy will be done.
MATT|26|43|And he came and found them asleep again: for their eyes were heavy.
MATT|26|44|And he left them, and went away again, and prayed the third time, saying the same words.
MATT|26|45|Then cometh he to his disciples, and saith unto them, Sleep on now, and take your rest: behold, the hour is at hand, and the Son of man is betrayed into the hands of sinners.
MATT|26|46|Rise, let us be going: behold, he is at hand that doth betray me.
MATT|26|47|And while he yet spake, lo, Judas, one of the twelve, came, and with him a great multitude with swords and staves, from the chief priests and elders of the people.
MATT|26|48|Now he that betrayed him gave them a sign, saying, Whomsoever I shall kiss, that same is he: hold him fast.
MATT|26|49|And forthwith he came to Jesus, and said, Hail, master; and kissed him.
MATT|26|50|And Jesus said unto him, Friend, wherefore art thou come? Then came they, and laid hands on Jesus and took him.
MATT|26|51|And, behold, one of them which were with Jesus stretched out his hand, and drew his sword, and struck a servant of the high priest's, and smote off his ear.
MATT|26|52|Then said Jesus unto him, Put up again thy sword into his place: for all they that take the sword shall perish with the sword.
MATT|26|53|Thinkest thou that I cannot now pray to my Father, and he shall presently give me more than twelve legions of angels?
MATT|26|54|But how then shall the scriptures be fulfilled, that thus it must be?
MATT|26|55|In that same hour said Jesus to the multitudes, Are ye come out as against a thief with swords and staves for to take me? I sat daily with you teaching in the temple, and ye laid no hold on me.
MATT|26|56|But all this was done, that the scriptures of the prophets might be fulfilled. Then all the disciples forsook him, and fled.
MATT|26|57|And they that had laid hold on Jesus led him away to Caiaphas the high priest, where the scribes and the elders were assembled.
MATT|26|58|But Peter followed him afar off unto the high priest's palace, and went in, and sat with the servants, to see the end.
MATT|26|59|Now the chief priests, and elders, and all the council, sought false witness against Jesus, to put him to death;
MATT|26|60|But found none: yea, though many false witnesses came, yet found they none. At the last came two false witnesses,
MATT|26|61|And said, This fellow said, I am able to destroy the temple of God, and to build it in three days.
MATT|26|62|And the high priest arose, and said unto him, Answerest thou nothing? what is it which these witness against thee?
MATT|26|63|But Jesus held his peace, And the high priest answered and said unto him, I adjure thee by the living God, that thou tell us whether thou be the Christ, the Son of God.
MATT|26|64|Jesus saith unto him, Thou hast said: nevertheless I say unto you, Hereafter shall ye see the Son of man sitting on the right hand of power, and coming in the clouds of heaven.
MATT|26|65|Then the high priest rent his clothes, saying, He hath spoken blasphemy; what further need have we of witnesses? behold, now ye have heard his blasphemy.
MATT|26|66|What think ye? They answered and said, He is guilty of death.
MATT|26|67|Then did they spit in his face, and buffeted him; and others smote him with the palms of their hands,
MATT|26|68|Saying, Prophesy unto us, thou Christ, Who is he that smote thee?
MATT|26|69|Now Peter sat without in the palace: and a damsel came unto him, saying, Thou also wast with Jesus of Galilee.
MATT|26|70|But he denied before them all, saying, I know not what thou sayest.
MATT|26|71|And when he was gone out into the porch, another maid saw him, and said unto them that were there, This fellow was also with Jesus of Nazareth.
MATT|26|72|And again he denied with an oath, I do not know the man.
MATT|26|73|And after a while came unto him they that stood by, and said to Peter, Surely thou also art one of them; for thy speech bewrayeth thee.
MATT|26|74|Then began he to curse and to swear, saying, I know not the man. And immediately the cock crew.
MATT|26|75|And Peter remembered the word of Jesus, which said unto him, Before the cock crow, thou shalt deny me thrice. And he went out, and wept bitterly.
MATT|27|1|When the morning was come, all the chief priests and elders of the people took counsel against Jesus to put him to death:
MATT|27|2|And when they had bound him, they led him away, and delivered him to Pontius Pilate the governor.
MATT|27|3|Then Judas, which had betrayed him, when he saw that he was condemned, repented himself, and brought again the thirty pieces of silver to the chief priests and elders,
MATT|27|4|Saying, I have sinned in that I have betrayed the innocent blood. And they said, What is that to us? see thou to that.
MATT|27|5|And he cast down the pieces of silver in the temple, and departed, and went and hanged himself.
MATT|27|6|And the chief priests took the silver pieces, and said, It is not lawful for to put them into the treasury, because it is the price of blood.
MATT|27|7|And they took counsel, and bought with them the potter's field, to bury strangers in.
MATT|27|8|Wherefore that field was called, The field of blood, unto this day.
MATT|27|9|Then was fulfilled that which was spoken by Jeremy the prophet, saying, And they took the thirty pieces of silver, the price of him that was valued, whom they of the children of Israel did value;
MATT|27|10|And gave them for the potter's field, as the Lord appointed me.
MATT|27|11|And Jesus stood before the governor: and the governor asked him, saying, Art thou the King of the Jews? And Jesus said unto him, Thou sayest.
MATT|27|12|And when he was accused of the chief priests and elders, he answered nothing.
MATT|27|13|Then said Pilate unto him, Hearest thou not how many things they witness against thee?
MATT|27|14|And he answered him to never a word; insomuch that the governor marvelled greatly.
MATT|27|15|Now at that feast the governor was wont to release unto the people a prisoner, whom they would.
MATT|27|16|And they had then a notable prisoner, called Barabbas.
MATT|27|17|Therefore when they were gathered together, Pilate said unto them, Whom will ye that I release unto you? Barabbas, or Jesus which is called Christ?
MATT|27|18|For he knew that for envy they had delivered him.
MATT|27|19|When he was set down on the judgment seat, his wife sent unto him, saying, Have thou nothing to do with that just man: for I have suffered many things this day in a dream because of him.
MATT|27|20|But the chief priests and elders persuaded the multitude that they should ask Barabbas, and destroy Jesus.
MATT|27|21|The governor answered and said unto them, Whether of the twain will ye that I release unto you? They said, Barabbas.
MATT|27|22|Pilate saith unto them, What shall I do then with Jesus which is called Christ? They all say unto him, Let him be crucified.
MATT|27|23|And the governor said, Why, what evil hath he done? But they cried out the more, saying, Let him be crucified.
MATT|27|24|When Pilate saw that he could prevail nothing, but that rather a tumult was made, he took water, and washed his hands before the multitude, saying, I am innocent of the blood of this just person: see ye to it.
MATT|27|25|Then answered all the people, and said, His blood be on us, and on our children.
MATT|27|26|Then released he Barabbas unto them: and when he had scourged Jesus, he delivered him to be crucified.
MATT|27|27|Then the soldiers of the governor took Jesus into the common hall, and gathered unto him the whole band of soldiers.
MATT|27|28|And they stripped him, and put on him a scarlet robe.
MATT|27|29|And when they had platted a crown of thorns, they put it upon his head, and a reed in his right hand: and they bowed the knee before him, and mocked him, saying, Hail, King of the Jews!
MATT|27|30|And they spit upon him, and took the reed, and smote him on the head.
MATT|27|31|And after that they had mocked him, they took the robe off from him, and put his own raiment on him, and led him away to crucify him.
MATT|27|32|And as they came out, they found a man of Cyrene, Simon by name: him they compelled to bear his cross.
MATT|27|33|And when they were come unto a place called Golgotha, that is to say, a place of a skull,
MATT|27|34|They gave him vinegar to drink mingled with gall: and when he had tasted thereof, he would not drink.
MATT|27|35|And they crucified him, and parted his garments, casting lots: that it might be fulfilled which was spoken by the prophet, They parted my garments among them, and upon my vesture did they cast lots.
MATT|27|36|And sitting down they watched him there;
MATT|27|37|And set up over his head his accusation written, THIS IS JESUS THE KING OF THE JEWS.
MATT|27|38|Then were there two thieves crucified with him, one on the right hand, and another on the left.
MATT|27|39|And they that passed by reviled him, wagging their heads,
MATT|27|40|And saying, Thou that destroyest the temple, and buildest it in three days, save thyself. If thou be the Son of God, come down from the cross.
MATT|27|41|Likewise also the chief priests mocking him, with the scribes and elders, said,
MATT|27|42|He saved others; himself he cannot save. If he be the King of Israel, let him now come down from the cross, and we will believe him.
MATT|27|43|He trusted in God; let him deliver him now, if he will have him: for he said, I am the Son of God.
MATT|27|44|The thieves also, which were crucified with him, cast the same in his teeth.
MATT|27|45|Now from the sixth hour there was darkness over all the land unto the ninth hour.
MATT|27|46|And about the ninth hour Jesus cried with a loud voice, saying, Eli, Eli, lama sabachthani? that is to say, My God, my God, why hast thou forsaken me?
MATT|27|47|Some of them that stood there, when they heard that, said, This man calleth for Elias.
MATT|27|48|And straightway one of them ran, and took a spunge, and filled it with vinegar, and put it on a reed, and gave him to drink.
MATT|27|49|The rest said, Let be, let us see whether Elias will come to save him.
MATT|27|50|Jesus, when he had cried again with a loud voice, yielded up the ghost.
MATT|27|51|And, behold, the veil of the temple was rent in twain from the top to the bottom; and the earth did quake, and the rocks rent;
MATT|27|52|And the graves were opened; and many bodies of the saints which slept arose,
MATT|27|53|And came out of the graves after his resurrection, and went into the holy city, and appeared unto many.
MATT|27|54|Now when the centurion, and they that were with him, watching Jesus, saw the earthquake, and those things that were done, they feared greatly, saying, Truly this was the Son of God.
MATT|27|55|And many women were there beholding afar off, which followed Jesus from Galilee, ministering unto him:
MATT|27|56|Among which was Mary Magdalene, and Mary the mother of James and Joses, and the mother of Zebedees children.
MATT|27|57|When the even was come, there came a rich man of Arimathaea, named Joseph, who also himself was Jesus' disciple:
MATT|27|58|He went to Pilate, and begged the body of Jesus. Then Pilate commanded the body to be delivered.
MATT|27|59|And when Joseph had taken the body, he wrapped it in a clean linen cloth,
MATT|27|60|And laid it in his own new tomb, which he had hewn out in the rock: and he rolled a great stone to the door of the sepulchre, and departed.
MATT|27|61|And there was Mary Magdalene, and the other Mary, sitting over against the sepulchre.
MATT|27|62|Now the next day, that followed the day of the preparation, the chief priests and Pharisees came together unto Pilate,
MATT|27|63|Saying, Sir, we remember that that deceiver said, while he was yet alive, After three days I will rise again.
MATT|27|64|Command therefore that the sepulchre be made sure until the third day, lest his disciples come by night, and steal him away, and say unto the people, He is risen from the dead: so the last error shall be worse than the first.
MATT|27|65|Pilate said unto them, Ye have a watch: go your way, make it as sure as ye can.
MATT|27|66|So they went, and made the sepulchre sure, sealing the stone, and setting a watch.
MATT|28|1|In the end of the sabbath, as it began to dawn toward the first day of the week, came Mary Magdalene and the other Mary to see the sepulchre.
MATT|28|2|And, behold, there was a great earthquake: for the angel of the Lord descended from heaven, and came and rolled back the stone from the door, and sat upon it.
MATT|28|3|His countenance was like lightning, and his raiment white as snow:
MATT|28|4|And for fear of him the keepers did shake, and became as dead men.
MATT|28|5|And the angel answered and said unto the women, Fear not ye: for I know that ye seek Jesus, which was crucified.
MATT|28|6|He is not here: for he is risen, as he said. Come, see the place where the Lord lay.
MATT|28|7|And go quickly, and tell his disciples that he is risen from the dead; and, behold, he goeth before you into Galilee; there shall ye see him: lo, I have told you.
MATT|28|8|And they departed quickly from the sepulchre with fear and great joy; and did run to bring his disciples word.
MATT|28|9|And as they went to tell his disciples, behold, Jesus met them, saying, All hail. And they came and held him by the feet, and worshipped him.
MATT|28|10|Then said Jesus unto them, Be not afraid: go tell my brethren that they go into Galilee, and there shall they see me.
MATT|28|11|Now when they were going, behold, some of the watch came into the city, and shewed unto the chief priests all the things that were done.
MATT|28|12|And when they were assembled with the elders, and had taken counsel, they gave large money unto the soldiers,
MATT|28|13|Saying, Say ye, His disciples came by night, and stole him away while we slept.
MATT|28|14|And if this come to the governor's ears, we will persuade him, and secure you.
MATT|28|15|So they took the money, and did as they were taught: and this saying is commonly reported among the Jews until this day.
MATT|28|16|Then the eleven disciples went away into Galilee, into a mountain where Jesus had appointed them.
MATT|28|17|And when they saw him, they worshipped him: but some doubted.
MATT|28|18|And Jesus came and spake unto them, saying, All power is given unto me in heaven and in earth.
MATT|28|19|Go ye therefore, and teach all nations, baptizing them in the name of the Father, and of the Son, and of the Holy Ghost:
MATT|28|20|Teaching them to observe all things whatsoever I have commanded you: and, lo, I am with you alway, even unto the end of the world. Amen.
