NEH|1|1|Слова Неемії, Гахаліїного сина: І сталося в місяці кіслеві двадцятого року, і був я в замку Шушан.
NEH|1|2|І прийшов Ханані, один із братів моїх, він та люди з Юдеї. І запитався я їх про юдеїв, що врятувалися, що позостали від полону, та про Єрусалим.
NEH|1|3|А вони сказали мені: Позосталі, що лишилися з полону, там в окрузі, живуть у великій біді та в ганьбі, а мур Єрусалиму поруйнований, а брами його попалені огнем...
NEH|1|4|І сталося, як почув я ці слова, сів я та й плакав, і був у жалобі кілька днів, і постив, і молився перед лицем Небесного Бога.
NEH|1|5|І сказав я: Молю Тебе, Господи, Боже Небесний, Боже великий та грізний, що дотримуєш заповіта та милість для тих, хто любить Тебе та дотримуєш заповіді Свої,
NEH|1|6|нехай же буде ухо Твоє чутке, а очі Твої відкриті, щоб прислухуватися до молитви раба Твого, якою я молюся сьогодні перед Твоїм лицем день та ніч за Ізраїлевих синів, Твоїх рабів, і сповідаюся в гріхах Ізраїлевих синів, якими грішили ми проти Тебе, і я і дім батька мого грішили!
NEH|1|7|Ми сильно провинилися перед Тобою, і не дотримували заповідей, і уставів, і прав, які наказав Ти Мойсеєві, рабові Своєму.
NEH|1|8|Пам'ятай же те слово, що Ти наказав був Мойсеєві, Своєму рабові, говорячи: як ви спроневіритеся, Я розпорошу вас поміж народами!
NEH|1|9|Та коли навернетеся до Мене, і будете дотримувати заповіді Мої й виконувати їх, то якщо будуть ваші вигнанці на краю небес, то й звідти позбираю їх, і приведу до того місця, яке Я вибрав, щоб там перебувало Ім'я Моє!
NEH|1|10|А вони раби Твої та народ Твій, якого Ти викупив Своєю великою силою та міцною Своєю рукою.
NEH|1|11|Молю Тебе, Господи, нехай же буде ухо Твоє чутке до молитви Твойого раба та до молитви Твоїх рабів, що прагнуть боятися Ймення Твого! І дай же сьогодні успіху Своєму рабові, і дай знайти милосердя перед оцим мужем! А я був чашником царевим.
NEH|2|1|І сталося в місяці нісані, двадцятого року царя Артаксеркса, було раз вино перед ним. І взяв я те вино й дав цареві. І я, здавалося, не був сумний перед ним.
NEH|2|2|Та сказав мені цар: Чому обличчя твоє сумне, чи ти не хворий? Це не інше що, як тільки сум серця... І я вельми сильно злякався!
NEH|2|3|І сказав я до царя: Нехай цар живе навіки! Чому не буде сумне обличчя моє, коли місто дому гробів батьків моїх поруйноване, а брами його попалені огнем!...
NEH|2|4|І сказав мені цар: Чого ж ти просиш? І я помолився до Небесного Бога,
NEH|2|5|і сказав цареві: Якщо це цареві вгодне, і якщо раб твій уподобаний перед обличчям твоїм, то пошли мене до Юдеї, до міста гробів батьків моїх, і я відбудую його!
NEH|2|6|І сказав мені цар (а цариця сиділа при ньому): Скільки часу буде дорога твоя, і коли ти повернешся? І сподобалось це цареві, і він послав мене, а я призначив йому час.
NEH|2|7|І сказав я цареві: Якщо це цареві вгодне, нехай дадуть мені листи до намісників Заріччя, щоб провадили мене, аж поки не прийду до Юдеї,
NEH|2|8|і листа до Асафа, дозорця царевого лісу, щоб дав мені дерева на брусся для замкових брам, що належать до Божого дому, і для міського муру, і для дому, що до нього ввійду. І дав мені цар в міру того, як добра була Божа рука надо мною.
NEH|2|9|І прибув я до намісників Заріччя, і дав їм цареві листи. А цар послав зо мною зверхників війська та верхівців.
NEH|2|10|І почув про це хоронянин Санваллат та раб аммонітянин Товія, і було їм прикро, дуже прикро, що прийшов чоловік клопотатися про добро для Ізраїлевих синів.
NEH|2|11|І прийшов я до Єрусалиму, і був там три дні.
NEH|2|12|І встав я вночі, я та трохи людей зо мною, і не розповів я нікому, що Бог мій дав до мого серця зробити для Єрусалиму. А худоби не було зо мною, окрім тієї худоби, що я нею їздив.
NEH|2|13|І вийшов я Долинною брамою вночі, і пішов до джерела Таннін, і до брами Смітникової. І я докладно оглянув мури Єрусалиму, що були поруйновані, а брами його були попалені огнем.
NEH|2|14|І перейшов я до Джерельної брами та до царського ставу, та там не було місця для переходу худоби, що була підо мною.
NEH|2|15|І йшов я долиною вночі, і докладно оглядав мура. Потім я вернувся, і ввійшов Долинною брамою, і вернувся.
NEH|2|16|А заступники не знали, куди я пішов та що я роблю, а юдеям, і священикам, і шляхті, і заступникам, і решті тих, що робили працю, я доти нічого не розповідав.
NEH|2|17|І сказав я до них: Ви бачите біду, що ми в ній, що Єрусалим зруйнований, а брами його попалені огнем. Ідіть, і збудуйте мура Єрусалиму, і вже не будемо ми ганьбою!...
NEH|2|18|І розповів я їм про руку Бога мого, що вона добра до мене, а також слова царя, які сказав він мені. І сказали вони: Станемо й збудуємо! І зміцнили вони руки свої на добре діло.
NEH|2|19|І почув це хоронянин Санваллат та аммонітянин раб Товія, і араб Ґешем, і сміялися з нас, і погорджували нами й говорили: Що це за річ, яку ви робите? Чи проти царя ви бунтуєтесь?
NEH|2|20|А я їм відповів і сказав до них: Небесний Бог Він дасть нам успіх, а ми, Його раби, станемо й збудуємо! А вам нема ані частки, ані права, ані пам'ятки в Єрусалимі!
NEH|3|1|І встав Еліяшів, первосвященик, та брати його священики, і збудували Овечу браму. Вони освятили її, і повставляли її двері, й аж до башти Меа освятили її, аж до башти Ханан'їла.
NEH|3|2|А поруч нього будували єрихоняни, а поруч них будував Заккур, син Імріїв.
NEH|3|3|А браму Рибну збудували сини Сенаїні, і вони покрили її бруссями, і повставляли двері її, замки її та засуви її.
NEH|3|4|А поруч них направляв Меремот, син Урії, Коцового сина, а поруч них направляв Мешуллам, син Берехії, Мешав'їлового сина, а поруч них направляв Садок, Баанин син.
NEH|3|5|А поруч них направляли текояни, але їхні вельможі не схилили своєї шиї в службу свого Господа.
NEH|3|6|А браму Стару направляли Йояда, син Пасеахів, та Мешуллам, син Бесодеїн, вони покривали бруссями, і вставляли двері її, і замки її та засуви її.
NEH|3|7|А поруч них направляв ґів'онеянин Мелатія та меронотеянин Ядон, люди Ґів'ону та Міцпи, що належали до володіння намісника Заріччя.
NEH|3|8|Поруч нього направляв Уззіїл, син Хархаїн, з золотарів, а поруч нього направляв Хананія, син Раккахімів, і вони відновили Єрусалима аж до Широкого муру.
NEH|3|9|А поруч нього направляв Рефая, син Хурів, зверхник половини єрусалимської округи.
NEH|3|10|А поруч нього направляв Єдая, син Харумафів, а то навпроти дому свого, а при його руці направляв Хаттуш, син Хашавнеїн.
NEH|3|11|Другу міру направляв Малкійя, син Харімів, та Хашшув, син Пахат-Моавів, та башту Печей.
NEH|3|12|А поруч нього направляв Шаллум, син Лохеша, зверхник половини єрусалимської округи, він та дочка його.
NEH|3|13|Браму Долинну направляв Ханун та мешканці Заноаху, вони збудували її, і повставляли двері її, замки її та засуви її, і тисячу ліктів у мурі аж до Смітникової брами.
NEH|3|14|А Смітникову браму направив Малкійя, син Рехавів, зверхник бет-керемської округи, він збудував її, і повставляв її двері, замки її та засуви її.
NEH|3|15|А Джерельну браму направив Шаллум, син Кол-Хезеїв, зверхник округи Міцпи, він збудував її, і покрив її, і повставляв її двері, замки її та засуви її, і направив мура ставу Шелах до царського садка, і аж до ступенів, що спускаються з Давидового Міста.
NEH|3|16|За ним направляв Неемія, син Азбуків, зверхник половини бетцурської округи аж до місця навпроти Давидових гробів і аж до зробленого ставу, і аж до дому Лицарів.
NEH|3|17|За ним направляли Левити: Рехум, син Баніїв, поруч нього направляв зверхник половини округи Кеїла, для своєї округи.
NEH|3|18|За ним направляли їхні брати: Баввай, син Хенададів, зверхник половини округи Кеїла.
NEH|3|19|І направляв поруч нього Езер, син Єшуїн, зверхник округи, міру другу, від місця навпроти виходу до зброярні наріжника.
NEH|3|20|За ним ревно направляв Барух, Заббаїв син, міру другу, від наріжника аж до входу до дому первосвященика Еліяшіва.
NEH|3|21|За ним направляв Меремот, син Урійї, сина Коцового, міру другу, від входу до Еліяшівового дому й аж до кінця Еліяшівового дому.
NEH|3|22|А за ним направляли священики, люди йорданської округи.
NEH|3|23|За ним направляв Веніямин, син Хашшувів, навпроти свого дому; за ним направляв Азарія, син Маасеї, сина Ананіїного, при своєму домі.
NEH|3|24|За ним направляв Біннуй, син Хенададів, міру другу, від Азаріїного дому аж до наріжника й аж до рогу.
NEH|3|25|Палал, син Узаїв, від місця навпроти наріжника та в горішній башті, що виходить із царського дому, що при в'язничному подвір'ї. За ним Педая, син Пар'ошів.
NEH|3|26|А підданці храму сиділи в Офелі аж до місця навпроти Водної брами на схід та навпроти виступаючої башти.
NEH|3|27|За ним направляли техояни, міру другу, від місця навпроти великої виступаючої башти й аж до офельського муру.
NEH|3|28|З-над Кінської брами направляли священики, кожен навпроти дому свого.
NEH|3|29|За ними направляв Садок, син Іммерів, навпроти свого дому, а за ним направляв Шемая, син Шеханіїн, сторож Східньої брами.
NEH|3|30|За ним направляв Хананія, син Шелеміїн, та Ханун, шостий син Цалафів, міру другу; за ним направляв Мешуллам, син Берехіїн, навпроти своєї кімнати.
NEH|3|31|За ним направляв Малкійя, син золотаря, аж до дому храмових підданців та крамарів, навпроти брами Міфкад і аж до наріжної горниці.
NEH|3|32|А між наріжною горницею до Овечої брами направляли золотарі та крамарі.
NEH|4|1|(3-33) І сталося, як почув Санваллат, що ми будуємо того мура, то він запалився гнівом, і дуже розгнівався, і сміявся з юдеїв.
NEH|4|2|(3-34) І говорив він перед своїми братами та самарійським військом і сказав: Що це роблять ці мізерні юдеї? Чи їм це позоставлять? Чи будуть вони приносити жертву? Чи закінчать цього дня? Чи оживлять вони ці каміння з куп пороху, а вони ж попалені?
NEH|4|3|(3-35) А аммонітянин Товійя був при ньому й сказав: Та й що вони будують? Якщо вийде лисиця, то вона зробить дірку в їхній камінній стіні!...
NEH|4|4|(3-36) Почуй, Боже наш, що ми стали погордою, і поверни їхню ганьбу на голову їхню, і дай їх на здобич у край полону!
NEH|4|5|(3-37) І не закрий їхньої провини, а їхній гріх нехай не буде стертий з-перед лиця Твого, бо вони образили будівничих!
NEH|4|6|(3-38) І збудували ми того мура, і був пов'язаний увесь той мур аж до половини його. А серце народу було, щоб далі робити!
NEH|4|7|(4-1) І сталося, як почув Санваллат, і Товійя, і араби, і аммонітяни, і ашдодяни, що направляється єрусалимський мур, що виломи в стіні стали затарасовуватися, то дуже запалилися гнівом.
NEH|4|8|(4-2) І змовилися вони всі разом, щоб іти воювати з Єрусалимом, та щоб учинити йому замішання.
NEH|4|9|(4-3) І ми молилися до нашого Бога, і поставили проти них сторожу вдень та вночі, перед ними.
NEH|4|10|(4-4) І сказав Юда: Ослабла сила носія, а звалищ багато, і ми не зможемо далі будувати мура!...
NEH|4|11|(4-5) А наші ненависники говорили: Вони не знатимуть і не побачать, як ми прийдемо до середини їх, і позабиваємо їх, та й спинимо працю!
NEH|4|12|(4-6) І сталося, як приходили ті юдеяни, що сиділи при них, то говорили нам про це разів десять, зо всіх місць, де вони пробували.
NEH|4|13|(4-7) Тоді поставив я сторожу здолу того місця за муром у печерах. І поставив я народ за їхніми родами, з їхніми мечами, їхніми ратищами та їхніми луками.
NEH|4|14|(4-8) І розглянув я це, і встав і сказав я до шляхетних, і до заступників, і до решти народу: Не бійтеся перед ними! Згадайте Господа великого та грізного, і воюйте за ваших братів, ваших синів, дочок ваших, жінок ваших та за доми ваші!
NEH|4|15|(4-9) І сталося, як почули наші вороги, що нам те відоме, то Господь зламав їхній задум, і всі ми вернулися до муру, кожен до праці своєї.
NEH|4|16|(4-10) І було від того дня, що половина моїх юнаків робили працю, а половина їх міцно тримала списи, щити, і луки та панцері, а зверхники стояли позад Юдиного дому.
NEH|4|17|(4-11) Будівничі працювали на мурі, а носії наладовували тягар, вони однією рукою робили працю, а однією міцно тримали списа...
NEH|4|18|(4-12) А в кожного будівничого його меч був прив'язаний на стегнах його, і так вони будували, а біля мене був сурмач.
NEH|4|19|(4-13) І сказав я до шляхетних, до заступників та до решти народу: Праця велика й простора, а ми повідділювані на мурі, далеко один від одного.
NEH|4|20|(4-14) Тому то в місце, де почуєте голос сурми, туди негайно збирайтеся до нас. Бог наш буде воювати для нас!
NEH|4|21|(4-15) І так ми робили працю, і половина їх міцно тримала списи від сходу ранньої зорі аж до появлення зір.
NEH|4|22|(4-16) Також того часу сказав я до народу: Кожен з юнаком своїм нехай ночують у середині Єрусалиму, і будуть вони для нас уночі сторожею, а вдень на працю.
NEH|4|23|(4-17) І ні я, ані брати мої, ані юнаки мої, ані сторожі, що були за мною, ми не здіймали своєї одежі, кожен мав свою зброю при своєму стегні.
NEH|5|1|І був великий крик народу та їхніх жінок на своїх братів юдеїв.
NEH|5|2|І були такі, що говорили: Ми даємо в заставу синів своїх та дочок своїх, і беремо збіжжя, і їмо й живемо!
NEH|5|3|І були такі, що говорили: Ми заставляємо поля свої, і виноградники свої, і доми свої, і беремо збіжжя в цьому голоді!
NEH|5|4|І були такі, що говорили: Ми позичаємо срібло на податок царський за наші поля та наші виноградники.
NEH|5|5|А наше ж тіло таке, як тіло наших братів, наші сини як їхні сини. А ось ми тиснемо наших синів та наших дочок за рабів, і є з наших дочок утискувані. Ми не в силі робити, а поля наші та виноградники наші належать іншим...
NEH|5|6|І сильно запалав у мені гнів, коли я почув їхній крик та ці слова!
NEH|5|7|А моє серце дало мені раду, і я сперечався з шляхетними та з заступниками та й сказав їм: Ви заставою тиснете один одного! І скликав я на них великі збори.
NEH|5|8|І сказав я до них: Ми викуповуємо своїх братів юдеїв, проданих поганам, за нашою спромогою, а ви будете продавати своїх братів, і вони продаються нам? І мовчали вони, і не знаходили слова...
NEH|5|9|І сказав я: Не добра це річ, що ви робите! Чи ж не в боязні нашого Бога ви маєте ходити, через ганьбу від тих поганів, наших ворогів?
NEH|5|10|Також і я, брати мої та юнаки мої були позикодавцями срібла та збіжжя. Опустімо ж ми оцей борг!
NEH|5|11|Верніть їм зараз їхні поля, їхні виноградники, їхні оливки, й їхні доми та відсоток срібла, і збіжжя, виноградний сік та нову оливу, що ви дали їм у заставу за них!
NEH|5|12|І вони сказали: Повернемо, і не будемо жадати від них! Зробимо так, як ти говориш! І покликав я священиків, і заприсягнув їх зробити за цим словом.
NEH|5|13|Витрусив я й свою пазуху та й сказав: Нехай отак витрусить Бог кожного чоловіка, хто не сповнить цього слова, з дому його та з труду його, і нехай буде такий витрушений та порожній! І сказали всі збори: Амінь! І славили вони Господа, і народ зробив за цим словом.
NEH|5|14|Також від дня, коли цар наказав мені бути їхнім намісником в Юдиному краї від року двадцятого й аж до року тридцять другого царя Артаксеркса, дванадцять літ не їв намісничого хліба ані я, ані брати мої.
NEH|5|15|А намісники попередні, що були передо мною, чинили тяжке над народом, і брали від них хлібом та вином одного дня сорок шеклів срібла; також їхні слуги панували над народом. А я не робив так через страх Божий.
NEH|5|16|також у праці того муру я підтримував, і поля не купували ми, а всі мої слуги були зібрані там над працею.
NEH|5|17|А за столом моїм були юдеї та заступники, сто й п'ятдесят чоловіка, та й ті, хто приходив до нас із народів, що навколо нас.
NEH|5|18|А що готовилося на один день, було: віл один, худоби дрібної шестеро вибраних, і птиця готувалася в мене, а за десять день виходило багато всякого вина. А при тому я не жадав намісничого хліба, бо та робота направи мурів була тяжка на тому народі.
NEH|5|19|Запам'ятай же мені, Боже мій, на добре все те, що я робив для цього народу!
NEH|6|1|І сталося, коли почув Санваллат, і Товійя, і араб Ґешем та решта наших ворогів, що я збудував мура, і що не позосталося в ньому вилому, але до цього часу дверей у брамах я не повставляв,
NEH|6|2|то послав Санваллат та Ґешем до мене, говорячи: Приходь, і вмовимося разом у Кефірімі в долині Оно! А вони замишляли зробити мені зло...
NEH|6|3|І послав я до них послів, говорячи: Я роблю велику працю, і не можу прийти. Нащо буде перервана ця праця, як кину її та піду до вас?
NEH|6|4|І посилали до мене так само чотири рази, а я відповідав їм так само.
NEH|6|5|І так само Санваллат п'ятий раз прислав до мене слугу свого, а в руці його був відкритий лист.
NEH|6|6|А в ньому написане: Чується серед народів, і Ґашму говорить: Ти та юдеї замишляєте відділитися, тому то ти будуєш того мура, і хочеш бути їм за царя, за тими словами.
NEH|6|7|Та й пророків ти понаставляв, щоб викрикували про тебе в Єрусалимі, говорячи: Цар в Юді! А тепер цар почує оці речі. Отож, приходь, і порадьмося разом!
NEH|6|8|І послав я до нього, говорячи: Не було таких речей, про які ти говориш, бо з серця свого ти їх повимишляв!...
NEH|6|9|Бо всі вони лякали нас, говорячи: Нехай ослабнуть їхні руки з цієї праці, і не буде вона зроблена! Та тепер, о Боже, зміцни мої руки!
NEH|6|10|І я ввійшов до дому Шемаї, сина Делаї, Мегетав'їлового сина, а він був задержаний. І він сказав: Умовмося піти до Божого дому, до середини храму, і замкнемо храмові двері, бо прийдуть забити тебе, власне вночі прийдуть забити тебе...
NEH|6|11|Та я відказав: Чи такий чоловік, як я, має втікати? І хто є такий, як я, що ввійде до храму й буде жити? Не ввійду!
NEH|6|12|І пізнав я, що то не Бог послав його, коли він говорив на мене те пророцтво, а то Товійя та Санваллат підкупили його...
NEH|6|13|Бо він був підкуплений, щоб я боявся, і зробив так, і згрішив. Це було для них на злий поговір, щоб образити мене.
NEH|6|14|Запам'ятай же, Боже мій, Товійї та Санваллатові за цими вчинками його, а також пророчиці Ноадії та решті пророків, що страхали мене!
NEH|6|15|І був закінчений мур двадцятого й п'ятого дня місяця елула, за п'ятдесят і два дні.
NEH|6|16|І сталося, як почули про це всі наші вороги, та побачили всі народи, що були навколо нас, то вони впали в очах своїх та й пізнали, що ця праця була зроблена від нашого Бога!
NEH|6|17|Тими днями також шляхетні юдеї писали багато своїх листів, що йшли до Товійї, а Товійїні приходили до них.
NEH|6|18|Бо багато-хто в Юдеї були заприсяженими приятелями йому, бо він був зять Шеханії, Арахового сина, а син його Єгоханан узяв дочку Мешуллама, Берехіїного сина.
NEH|6|19|І говорили передо мною добре про нього, а слова мої передавали йому. Товійя посилав листи, щоб настрахати мене.
NEH|7|1|І сталося, як був збудований мур, то повставляв я двері, і були понаставлювані придверні, співаки та Левити.
NEH|7|2|І призначив я над Єрусалимом свого брата Ханані та зверхника твердині Хананію, бо він був чоловік правдивий, і Бога боявся більше від багатьох інших.
NEH|7|3|І сказав я до них: Нехай не відчиняються єрусалимські брами аж до спеки сонця. І поки вони самі стоять, нехай позамикають двері, і так тримайте. І поставити варти з єрусалимських мешканців, кожного на його сторожі, і кожного навпроти його дому!
NEH|7|4|А місто було широко-просторе й велике, та народу в ньому мало, і доми не були побудовані.
NEH|7|5|І поклав мені Бог мій на серце моє зібрати шляхетних, і заступників та народ, щоб переписати. І знайшов я книжку перепису тих, хто прийшов перше, а в ній я знайшов написане таке:
NEH|7|6|Оце виходьки з округи, що прийшли з полону вигнання, яких вигнав був Навуходоносор, цар вавилонський, і вони повернулися до Єрусалиму та до Юдеї, кожен до міста свого,
NEH|7|7|ті, що прийшли були з Зоровавелем, Ісусом, Неемією, Азарією, Раамією, Нахаманієм, Мордехаєм, Білшаном, Місперетом, Біґваєм, Нехумом, Бааною. Число людей Ізраїлевого народу:
NEH|7|8|синів Пар'ошових дві тисячі сто й сімдесят і два,
NEH|7|9|синів Шеватіїних три сотні і сімдесят і два,
NEH|7|10|синів Арахових шість сотень п'ятдесят і два,
NEH|7|11|синів Пахат-Моавових, із синів Ісусових та Йоавових дві тисячі й вісім сотень вісімнадцять,
NEH|7|12|синів Еламових тисяча двісті п'ятдесят і чотири,
NEH|7|13|синів Заттуєвих вісім сотень сорок і п'ять,
NEH|7|14|синів Заккаєвих сім сотень і шістдесят,
NEH|7|15|синів Біннуєвих шість сотень сорок і вісім,
NEH|7|16|синів Беваєвих шість сотень двадцять і вісім,
NEH|7|17|синів Азґадових дві тисячі три сотні двадцять і два,
NEH|7|18|синів Адонікамових шість сотень шістдесят і сім,
NEH|7|19|синів Біґваєвих дві тисячі шістдесят і сім,
NEH|7|20|синів Адінових шість сотень п'ятдесят і п'ять,
NEH|7|21|синів Атерових, з синів Хізкійїних дев'ятдесят і вісім,
NEH|7|22|синів Хашумових три сотні двадцять і вісім,
NEH|7|23|синів Бецаєвих три сотні двадцять і чотири,
NEH|7|24|синів Харіфових сто дванадцять,
NEH|7|25|синів Ґів'онових дев'ятдесят і п'ять,
NEH|7|26|людей з Віфлеєму та Нетофи сто вісімдесят і вісім,
NEH|7|27|людей з Анототу сто двадцять і вісім,
NEH|7|28|людей з Бет-Азмавету сорок і два,
NEH|7|29|людей з Кір'ят-Єаріму, Кефіри та Беероту сім сотень сорок і три,
NEH|7|30|людей з Рами та Ґави шість сотень двадцять і один,
NEH|7|31|людей з Міхмасу сто двадцять і два,
NEH|7|32|людей з Бет-Елу та Аю сто двадцять і три,
NEH|7|33|людей з Нево Другого п'ятдесят і два,
NEH|7|34|виходьків з Еламу Другого тисяча двісті п'ятдесят і чотири,
NEH|7|35|виходьків з Харіму три сотні й двадцять,
NEH|7|36|виходьків з Єрихону три сотні сорок і п'ять,
NEH|7|37|виходьків з Лоду, Хадіду й Оно сім сотень і двадцять і один,
NEH|7|38|виходьків з Сенаї три тисячі дев'ять сотень і тридцять.
NEH|7|39|Священиків: синів Єдаїних з Ісусового дому дев'ять сотень сімдесят і три,
NEH|7|40|синів Іммерових тисяча п'ятдесят і два,
NEH|7|41|синів Пашхурових тисяча двісті сорок і сім,
NEH|7|42|синів Харімових тисяча сімнадцять.
NEH|7|43|Левитів: синів Ісусових з Кадміїлового дому, з Годевиних синів сімдесят і чотири.
NEH|7|44|Співаків: синів Асафових сто сорок і вісім.
NEH|7|45|Придверних: синів Шаллумових, синів Атерових, синів Талмонових, синів Аккувових, синів Хатітиних, синів Шоваєвих сто тридцять і вісім.
NEH|7|46|Храмових підданців: сини Ціхині, сини Хасуфині, сини Таббаотові,
NEH|7|47|сини Керосові, сини Сіїні, сини Падонові,
NEH|7|48|сини Леванині, сини Хаґавині, сини Салмаєві,
NEH|7|49|сини Хананові, сини Ґідделові, сини Ґахарові,
NEH|7|50|сини Реаїні, сини Рецінові, сини Некодині,
NEH|7|51|сини Ґаззамові, сини Уззині, сини Пасеахові,
NEH|7|52|сини Бесаєві, сини Меунімові, сини Нефішесінові,
NEH|7|53|сини Бакбутові, сини Хакуфині, сини Хархурові,
NEH|7|54|сини Бацлітові, сини Мехидині, сини Харшині,
NEH|7|55|сини Баркосові, сини Сісерині, сини Темахові,
NEH|7|56|сини Неціяхові, сини Хатіфині.
NEH|7|57|Синів Соломонових рабів: сини Сотаєві, сини Соферетові, сини Перідині,
NEH|7|58|сини Яалині, сини Дарконові, сини Ґідделові,
NEH|7|59|сини Шефатіїні, сини Хаттілові, сини Похерет-Гаццеваїмові, сини Амонові,
NEH|7|60|усього цих храмових підданців та синів Соломонових рабів три сотні дев'ятдесят і два.
NEH|7|61|А оце ті, що прийшли з Тел-Мелаху, з Тел-Харші, Керув-Аддону та Іммеру, та не могли довести роду батьків своїх та свого насіння, чи вони з Ізраїля:
NEH|7|62|синів Делаїних, синів Товійїних, синів Некодиних шість сотень сорок і два.
NEH|7|63|А з священиків: сини Ховаїні, сини Коцові, сини Барзіллая, що взяв жінку з дочок ґілеадянина Барзіллая, і став зватися їхнім ім'ям.
NEH|7|64|Вони шукали запису свого родоводу, але він не знайшовся, і були вони вилучені зо священства,
NEH|7|65|а намісник сказав їм, щоб вони не їли зо Святого Святих, аж поки не стане священик до уріму та тумміму.
NEH|7|66|Усього збору разом сорок дві тисячі триста й шістдесят,
NEH|7|67|окрім їхніх рабів та їхніх невільниць, цих було сім тисяч триста тридцять і сім; а в них співаків та співачок двісті й сорок і п'ять.
NEH|7|68|Їхніх коней було сім сотень тридцять і шість, їхніх мулів двісті сорок і п'ять,
NEH|7|69|верблюдів чотири сотні тридцять і п'ять, ослів шість тисяч і сім сотень і двадцять.
NEH|7|70|А частина голів батьківських родів дали на працю: намісник дав до скарбниці: золота тисячу дарейків, кропильниць п'ятдесят, священичих шат п'ятсот і тридцять.
NEH|7|71|А з голів батьківських родів дали до скарбниці на працю: золота двадцять тисяч дарейків, а срібла дві тисячі й двісті мін.
NEH|7|72|А що дала решта народу: золота двадцять тисяч дарейків, а срібла дві тисячі мін, а священичих шат шістдесят і сім.
NEH|7|73|І осілися священики, і Левити, і придверні, і співаки, і дехто з народу, і храмові підданці, і ввесь Ізраїль по своїх містах. Як настав сьомий місяць, то Ізраїлеві сини були по своїх містах.
NEH|8|1|І зібрався ввесь народ, як один чоловік, на майдан, що перед Водною брамою, і сказали учителеві Ездрі принести книги Мойсеєвого Закону, що наказав був Господь Ізраїлеві.
NEH|8|2|І приніс священик Ездра Закона перед збори з чоловіків та аж до жінок, і всіх, хто розумів чуте, першого дня сьомого місяця.
NEH|8|3|І читав він у нім на майдані, що перед Водною брамою, від світанку аж до полудня, перед чоловіками й жінками та тими, хто розуміє, а уші всього народу були звернені до книги Закону.
NEH|8|4|І стояв учитель Ездра на дерев'яному підвищенні, що зробили для цієї справи, а при ньому стояв Маттітія, і Шема, і Аная, і Урійя, і Хілкійя, і Маасея на правиці його, а на лівиці його: Педая, і Мішаїл, і Малкійя, і Хашум, і Хашбаддана, Захарій, Мешуллам.
NEH|8|5|І розгорнув Ездра цю книгу на очах усього народу, бо він був вище від усього народу, а коли він розгорнув, увесь народ устав.
NEH|8|6|І поблагословив Ездра Господа, Бога великого, а ввесь народ відповів: Амінь, Амінь! з піднесенням своїх рук. І всі схилялися, і вклонялися Господеві обличчям до землі!
NEH|8|7|А Ісус, і Бані, і Шеревея, Ямін, Аккув, Шаббетай, Годійя, Маасея, Келіта, Азарія, Йозавад, Ханан, Пелая та Левити пояснювали народові Закона, а народ був на своєму місці.
NEH|8|8|І читали в книзі, у Божому Законі виразно, і вияснювали значення, і робили зрозумілим читане.
NEH|8|9|І сказав намісник Неемія, і священик учитель Ездра й Левити, що вияснювали народові, до всього народу: День цей святий він для Господа, Бога вашого, не будьте в жалобі й не плачте! Бо плакав увесь народ, як почув слова Закону...
NEH|8|10|І сказав він до них: Ідіть, їжте сите та пийте солодке, і посилайте частки тому, в кого нема наготовленого. Бо святий цей день для нашого Господа, і не сумуйте, бо радість у Господі це ваша сила!
NEH|8|11|І Левити потішали ввесь народ, говорячи: Мовчіть, бо цей день святий, і не сумуйте!
NEH|8|12|І пішов увесь народ їсти та пити, і посилати частки та чинити велику радість, бо розумів ті слова, що розповіли йому.
NEH|8|13|А другого дня зібралися голови батьківських родів усього народу, священики та Левити, до вчителя Ездри, щоб він виясняв їм слова Закону.
NEH|8|14|І знайшли написане в Законі, що наказав був Господь через Мойсея, щоб Ізраїлеві сини сиділи в кучках у свято сьомого місяця,
NEH|8|15|і щоб розголосили й оголосили по всіх своїх містах та в Єрусалимі, говорячи: Вийдіть на гору, і понаносьте галуззя оливкового, і галуззя дерева оливкового, і галуззя миртового, і галуззя пальмового, і галуззя густолистого дерева, щоб поробити кучки, як написано.
NEH|8|16|І вийшов народ, і поназношували, і поробили собі кучки кожен на даху своїм, і в подвір'ях своїх, і в подвір'ях Божого дому, і на майдані Водної брами, і на майдані брами Єфремової.
NEH|8|17|І поробила кучки вся громада, що вернулася з полону, і сиділа в кучках, бо не робили так Ізраїлеві сини від днів Ісуса, Навинового сина, аж до дня цього. І була дуже велика радість!
NEH|8|18|І читали в книзі Божого Закону щоденно, від першого дня аж до дня останнього. І справляли свято сім день; а восьмого дня віддання, за уставом.
NEH|9|1|А двадцятого й четвертого дня того місяця зібралися Ізраїлеві сини в пості та в веретищах, а на них порох.
NEH|9|2|А Ізраїлеве насіння відділилося від усіх чужинців, і поставали й визнавали гріхи свої та провини своїх батьків.
NEH|9|3|І стали на місті своїм, і чверть дня читали з книги Закону Господа, Бога свого, а чверть сповідалися і вклонялися Господеві, Богові своєму.
NEH|9|4|І стали не левитському підвищенні Ісус, і Бані, Кадміїл, Шеванія, Бунні, Шеревея, Бані, Кенані, і кликали сильним голосом до Господа, Бога свого.
NEH|9|5|І сказали Левити: Ісус, і Кадміїл, Бані, Хашавнея, Шеревея, Годійя, Шеванія, Петахія: Устаньте, поблагословіть Господа, Бога свого, від віку аж до віку! І нехай благословляють Ім'я слави Твоєї, і нехай воно буде звеличене над усяке благословення та славу!
NEH|9|6|Ти Господь єдиний! Ти вчинив небо, небеса небес, і все їхнє військо, землю та все, що на ній, моря та все, що в них, і Ти оживляєш їх усіх, а небесне військо Тобі вклоняється!
NEH|9|7|Ти то Господь, Бог, що вибрав Аврама, і вивів його з халдейського Уру, і дав йому ім'я Авраам.
NEH|9|8|І Ти знайшов серце його вірним перед лицем Своїм, і склав був із ним заповіта, щоб дати Край хананеян, хіттеян, амореян, періззеян, євусеян, ґірґасеян, щоб дати насінню його. І Ти виконав слова Свої, бо Ти праведний!
NEH|9|9|І побачив Ти біду наших батьків ув Єгипті, а їхній зойк Ти почув над Червоним морем.
NEH|9|10|І дав Ти знаки та чуда на фараоні та на всіх його рабах, і на всім народі краю його, бо пізнав Ти, що вони гордо поводилися з ними, і зробив Ти Собі Ім'я, як видно цього дня.
NEH|9|11|І море Ти розсік перед ними, і вони перейшли серед моря по суходолу, а тих, хто гнався за ними, Ти кинув до глибин, як камінь до бурхливої води.
NEH|9|12|І Ти провадив їх стовпом хмари вдень, а стовпом огню вночі, щоб освітлювати їм ту дорогу, якою мали йти.
NEH|9|13|І Ти зійшов був на гору Сінай, і говорив з ними з небес, і дав їм справедливі права та правдиві закони, устави та заповіді добрі.
NEH|9|14|І святу Свою суботу Ти вказав їм, а заповіді, й устави та право наказав Ти їм через раба Свого Мойсея.
NEH|9|15|І хліб із небес дав Ти був їм на їхній голод, і воду зо скелі Ти вивів був їм на їхню спрагу. І Ти сказав їм, щоб ішли посісти Край, який Ти присягнув дати їм.
NEH|9|16|Та вони й наші батьки були вперті, і робили твердою свою шию, і не слухали Твоїх заповідей.
NEH|9|17|І відмовлялися вони слухати, і не пам'ятали чуд Твоїх, які Ти чинив був із ними, і стали твердошиї, і настановили собі голову, щоб вернутися до своєї неволі в непослуху. Та Ти Бог, що прощаєш, Ти ласкавий та милосердний, довготерпеливий та багатомилостивий, і Ти не покинув їх!
NEH|9|18|Хоч вони зробили були собі литого тельця та сказали: Оце бог твій, що вивів тебе з Єгипту, і робили великі образи,
NEH|9|19|та Ти в великім Своїм милосерді не залишив їх у пустині, стовп хмари не відходив від них удень, щоб вести їх дорогою, а стовп огню вночі, щоб освітлювати їм дорогу, якою мали йти.
NEH|9|20|І Духа Свого доброго Ти давав, щоб зробити їх мудрими, і манни Своєї не стримував від їхніх уст, і воду Ти їм давав на їхнє прагнення.
NEH|9|21|І сорок літ живив Ти їх у пустині. Не було недостатку ні в чому, одежі їхні не дерлися, а ноги їхні не пухли.
NEH|9|22|І дав Ти їм царства та народи, які призначив на поділ, і вони посіли край Сигона, і край царя хешбонського, і край Оґа, царя башанського.
NEH|9|23|А їхніх синів Ти помножив, як зорі небесні, і ввів їх до Краю, що про нього казав Ти їхнім батькам, щоб ішли посісти.
NEH|9|24|І ввійшли сини, і посіли той Край, і Ти впокорив перед ними мешканців того Краю ханаанеян, і дав у їхню руку їх та царів їхніх, та народи того Краю, щоб чинити з ними за своєю волею.
NEH|9|25|І поздобували вони міста укріплені, та землю ситу, і посіли доми, повні всякого добра, повитесувані в скелях водозбори, виноградники, і оливки, і багато овочевих дерев. І вони їли й наситилися, і поставали товсті, і насолоджувалися Твоїм великим добром.
NEH|9|26|І стали вони неслухняні, і побунтувалися проти Тебе, і кинули Закона Твого геть за свою спину, і позабивали пророків Твоїх, що свідчили між ними, щоб навернути їх до Тебе. І чинили вони великі образи.
NEH|9|27|І дав Ти їх у руку їхніх ворогів, а ті утискали їх. А в часі горя свого вони кликали до Тебе, а Ти з неба чув, і за Своїм великим милосердям давав їм спасителів, і вони спасали їх з руки їхніх ворогів.
NEH|9|28|Та коли був їм мир, вони знову чинили зло перед лицем Твоїм, і Ти давав їх у руку їхніх ворогів, і ті панували над ними. І вони знову кликали до Тебе, а Ти з неба їх вислуховував, і спасав їх за милосердям Своїм довгий час.
NEH|9|29|І свідчив Ти проти них, щоб навернути їх до Закону Твого, та вони чинили лихе, і не слухалися заповідей Твоїх, і грішили проти Твоїх прав, які коли б людина чинила, то жила б ними, і ставало рамено їх неслухняне, а шию свою робили твердою, і не слухалися.
NEH|9|30|І зволікав Ти їм довгі роки, і свідчив проти них Своїм Духом через Своїх пророків, та вони не слухали того, і Ти дав їх у руку народів цих країв.
NEH|9|31|І через велике Своє милосердя Ти не вигубив і не покинув їх, бо Ти Бог ласкавий та милосердний!
NEH|9|32|А тепер, Боже наш, Боже великий, сильний та страшний, що бережеш заповіта та милість, нехай не буде малою перед лицем Твоїм уся та мука, що спіткала нас, наших царів, наших зверхників, і священиків наших, і пророків наших, і батьків наших, і ввесь Твій народ від днів асирійських царів аж до цього дня!
NEH|9|33|А ти справедливий у всьому, що приходить на нас, бо Ти правду робив, а ми були несправедливі.
NEH|9|34|А наші царі, наші зверхники, наші священики та наші батьки не виконували Закона Твого, і не слухалися заповідей Твоїх та свідоцтв Твоїх, що Ти свідчив проти них.
NEH|9|35|І вони в царстві своїм та в великім добрі Твоїм, яке Ти їм давав, і в тому просторому та ситому Краї, що Ти дав перед ними, не служили Тобі, і не відвернулися від своїх злих чинів.
NEH|9|36|Ось ми сьогодні раби, а цей Край, що Ти дав його нашим батькам, щоб їсти плід його та добро його, ось ми раби в ньому!
NEH|9|37|І він множить свій урожай для царів, яких Ти дав над нами за наші гріхи, і вони панують над нашими тілами та над нашою худобою за своїм уподобанням, і ми в великому утискові!
NEH|9|38|(10-1) Через те все ми складаємо певну умову, і підписуємо, а печатки кладуть наші зверхники, наші Левити, наші священики.
NEH|10|1|(10-2) А між тих, що поклали печатки, були: намісник Неемія, син Хахаліїн, і Цідкійя,
NEH|10|2|(10-3) Серая, Азарія, Єремія,
NEH|10|3|(10-4) Пашхур, Амарія, Малкійя,
NEH|10|4|(10-5) Хаттуш, Шеванія, Маллух,
NEH|10|5|(10-6) Харім, Меремот, Овадія,
NEH|10|6|(10-7) Даніїл, Ґіннетон, Барух,
NEH|10|7|(10-8) Мешуллам, Авійя, Мійямін,
NEH|10|8|(10-9) Маазія, Білґай, Шемая, оце священики.
NEH|10|9|(10-10) А Левити: Ісус, син Азаніїн, Біннуй, з Хенададових синів, Кадміїл.
NEH|10|10|(10-11) А їхні брати: Шеванія, Годійя, Келіта, Пелая, Ханан,
NEH|10|11|(10-12) Міха, Рехов, Хашавія,
NEH|10|12|(10-13) Заккур, Шеревія, Шеванія,
NEH|10|13|(10-14) Годійя, Бані, Беніну.
NEH|10|14|(10-15) Голови народу: Пар'ош, Пахат-Моав, Елам, Затту, Бані,
NEH|10|15|(10-16) Бунні, Аз'дад, Бевай,
NEH|10|16|(10-17) Адонійя, Біґвай, Адін,
NEH|10|17|(10-18) Атер, Хізкійя, Аззур,
NEH|10|18|(10-19) Годійя, Хашум, Бецай,
NEH|10|19|(10-20) Харіф, Анатот, Невай,
NEH|10|20|(10-21) Маґпіяш, Мешуллам, Хезір,
NEH|10|21|(10-22) Мешезав'їл, Садок, Яддуя,
NEH|10|22|(10-23) Пелатія, Ханан, Аная,
NEH|10|23|(10-24) Осія, Хананія, Хашшув,
NEH|10|24|(10-25) Галлохеш, Пілха, Шовек,
NEH|10|25|(10-26) Рехум, Хашавна, Маасея,
NEH|10|26|(10-27) і Ахійя, Ханан, Анан,
NEH|10|27|(10-28) Маллух, Харім, Баана.
NEH|10|28|(10-29) І решта народу, священики, Левити, придверні, співаки, храмові підданці, і кожен, відділений від народів краю до Божого Закону, їхні жінки, їхні сини, та їхні дочки, кожен знаючий та розуміючий,
NEH|10|29|(10-30) зміцняють присягу при браттях своїх, при своїх шляхетних, і вступили в клятву та присягу, щоб ходити в Божому Законі, що був даний через Мойсея, Божого раба, і щоб дотримуватися, і щоб виконувати всі заповіді Господа, нашого Бога, і права Його, і постанови Його,
NEH|10|30|(10-31) і що не дамо наших синів народам Краю, а їхніх дочок не візьмемо для наших синів.
NEH|10|31|(10-32) А від народів цього Краю, що спроваджують товари та всяке збіжжя в день суботній на продаж, не візьмемо від них у суботу та в святі дні, і сьомого року понехаємо землю та всякого роду борги.
NEH|10|32|(10-33) І поставили ми собі за обов'язок, щоб давати нам третину шекля в рік на службу дому нашого Бога,
NEH|10|33|(10-34) на хліб показний, і на постійний дар, і на постійне цілопалення, на суботи, на молодики, на свята, і на освячені речі, і на жертви за гріх на окуплення за Ізраїля, і на всяку працю дому нашого Бога.
NEH|10|34|(10-35) І кинули ми жеребки про пожертву дров, священики, Левити та народ, щоб приносити до дому нашого Бога, за домом наших батьків, на означені часи рік-річно, щоб палити на жертівнику Господа, нашого Бога, як написано в Законі,
NEH|10|35|(10-36) і щоб приносити первоплоди нашої землі та первоплоди всякого плоду зо всякого дерева рік-річно до Господнього дому,
NEH|10|36|(10-37) і первороджених синів наших та нашої худоби, як написано в Законі, і первороджених худоби нашої великої та худоби нашої дрібної, щоб приносити до дому нашого Бога до священиків, що служать у домі нашого Бога,
NEH|10|37|(10-38) і первопочаток наших діж, і наші приношення, і плід усякого дерева, молоде вино та оливу спровадимо священикам до кімнат дому нашого Бога, а десятину нашої землі Левитам. А вони, Левити, будуть збирати десятину по всіх містах нашої роботи.
NEH|10|38|(10-39) І буде священик, син Ааронів, із Левитами, коли Левити будуть збирати десятину, і Левити віднесуть десятину від десятини до дому нашого Бога до комір, до скарбниці.
NEH|10|39|(10-40) Бо до комір будуть зносити сини Ізраїлеві та сини Левитів приношення збіжжя, молодого вина та оливи, і там є речі святині, служачі священики, і придверні, і співаки. І ми не опустимо дому нашого Бога!
NEH|11|1|І сиділи зверхники народу в Єрусалимі, а решта народу кинули жеребки, щоб привести одного з десяти сидіти в Єрусалимі, місті святому, а дев'ять частин зостаються по інших містах.
NEH|11|2|І поблагословив народ усіх тих людей, що пожертвувалися сидіти в Єрусалимі.
NEH|11|3|А оце голови округи, що сиділи в Єрусалимі, а по Юдиних містах сиділи, кожен у своїй посілості, по своїх містах, Ізраїль, священики, і Левити, і храмові підданці, і сини Соломонових рабів.
NEH|11|4|А в Єрусалимі сиділи оці з синів Юдиних та з синів Веніяминових. Із синів Юдиних: Атая, син Уззійї, сина Захарія, сина Амарії, сина Шефатії, сина Магаліїла, із синів Перецових.
NEH|11|5|І Маасея, син Баруха, сина Кол-Хозе, сина Хазаї, сина Адаї, сина Йояріва, сина Захарія, сина Шілоні.
NEH|11|6|Усіх синів Перецових, що сиділи в Єрусалимі, було чотири сотні шістдесят і вісім хоробрих людей.
NEH|11|7|А оце Веніяминові сини: Саллу, син Мешуллама, сина Йоеда, сина Педаї, сина Кадаї, сина Маасеї, сина Ітіїла, сина Ісаї.
NEH|11|8|А по ньому: Ґаббай, Саллай, дев'ять сотень двадцять і вісім.
NEH|11|9|А Йоїл, син Зіхрі, був провідником над ними, а Юда, син Сенуїн, другий над містом.
NEH|11|10|Із священиків: Єдая, син Йоярів, Яхін,
NEH|11|11|Серая, син Хілкійї, сина Мешуллама, сина Садока, сина Мерайота, сина Ахітува, начальник у Божому домі.
NEH|11|12|А їхніх братів, що робили службу для Божого дому, вісім сотень і двадцять і два. І Адая, син Єрохама, сина Пелалії, сина Амці, сина Захарія, сина Пашхура, сина Малкійї,
NEH|11|13|а їхніх братів, голів батьківських родів, двісті сорок і два. І Амашсай, син Азаріїла, сина Ахезая, сина Мешіллемота, сина Іммера,
NEH|11|14|а їхніх братів, хоробрих вояків, сто двадцять і вісім, а провідник над ними Завдіїл, син Ґедоліма.
NEH|11|15|А з Левитів: Шемая, син Хашшува, сина Азрікама, сина Хашавії, сина Бунні.
NEH|11|16|А Шаббетай та Йозавад були над зовнішньою службою для Божого дому, з голів Левитів.
NEH|11|17|А Матанія, син Міхи, сина Завді, сина Асафового, був головою, що починав славословити при молитві, і Бакбукія, другий з братів його, і Авда, син Шаммуї, сина Ґалала, сина Єдутунового.
NEH|11|18|Усіх Левитів у святому місті було двісті вісімдесят і чотири.
NEH|11|19|А придверні: Аккув, Талмон та їхні брати, що сторожили при брамах, сто сімдесят і два.
NEH|11|20|А решта Ізраїля, священики, Левити були по всіх Юдиних містах, кожен у наділі своїм.
NEH|11|21|А храмові підданці сиділи в Офелі, а Ціха та Ґішпа були над підданцями.
NEH|11|22|А провідником Левитів в Єрусалимі був Уззі, син Бані, сина Хашавії, сина Маттанії, сина Міхи, з Асафових синів, співаків при службі Божого дому,
NEH|11|23|бо був царів наказ про них та певна оплата на співаків про кожен день.
NEH|11|24|А Петахія, син Мешезав'їла, із синів Зераха, сина Юдиного, був при руці царя для всіх справ народу.
NEH|11|25|А по дворах на полях своїх з Юдиних синів сиділи: в Кір'ят-Арбі та залежних її містах, і в Дівоні та залежних його містах, і в Єкавцеїлі та залежних його містах,
NEH|11|26|і в Єшуї, і в Моладі, і в Бет-Пелеті,
NEH|11|27|і в Хасар-Шуалі, і в Беер-Шеві та залежних його містах,
NEH|11|28|і в Ціклаґу, і в Мехоні та в залежних її містах,
NEH|11|29|і в Ен-Ріммоні, і в Цор'ї, і в Ярмуті,
NEH|11|30|Заноаху, Адулламі та дворах її, в Лахішу та полях його, в Азці та залежних її містах. І таборували вони від Беер-Шеви аж до долини Гінном.
NEH|11|31|А Веніяминові сини, починаючи від Ґеви, заселили оці міста: Міхмаш, і Айя, і Бет-Ел та залежні його міста,
NEH|11|32|Анатот, Нов, Ананія,
NEH|11|33|Хацор, Рама, Ґіттаїм,
NEH|11|34|Хадід, Цевоїм, Неваллат,
NEH|11|35|Лод і Оно, долина Харашім.
NEH|11|36|А з Левитів Юдині відділи жили в краю Веніямина.
NEH|12|1|А оце священики та Левити, що прийшли з Зоровавелем, сином Шеалтіїловим, та з Ісусом: Серая, Їрмея, Ездра,
NEH|12|2|Амарія, Маллух, Хаттуш,
NEH|12|3|Шеханія, Рехум, Меремот,
NEH|12|4|Іддо, Ґіннетой, Авійя,
NEH|12|5|Мійямін, Маадія, Білґа,
NEH|12|6|Шемая, і Йоярів, Єдая,
NEH|12|7|Саллу, Амок, Хілкійя, Єдая. Це голови священиків та брати їхні за днів Ісуса.
NEH|12|8|А Левити: Ісус, Біннуй, Кадміїл, Шеревея, Юда, Матанія, головний над славослов'ям він та брати його.
NEH|12|9|І Бакбукія та Унні, їхні брати, були навпроти них на сторожі.
NEH|12|10|А Ісус породив Йоякима, а Йояким породив Ел'яшіва, а Ел'яшів породив Йояду,
NEH|12|11|а Йояда породив Йонатана, а Йонатан породив Яддуя.
NEH|12|12|А за Йоякимових днів були священики, голови батьківських родів: з роду Сераїного Мерая, з Їрмеїного Хананія,
NEH|12|13|з Ездриного Мешуллам, з Амаріїного Єгоханан,
NEH|12|14|з Меліхового Йонатан, з Шеваніїного Йосип,
NEH|12|15|з Харімового Адна, з Мерайотового Хелкай,
NEH|12|16|з Іддового Захарій, з Ґіннетонового Мешуллам,
NEH|12|17|з Авійїного Зіхрі, з Мін'ямінового та з Моадеїного Пілтай,
NEH|12|18|з Білґиного Шаммуя, з Шемаїного Йонатан,
NEH|12|19|а з Йоярівового Маттенай, з Єдаїного Уззі,
NEH|12|20|з Саллаєвого Каллай, з Амокового Евер,
NEH|12|21|з Хілкійїного Хашавія, з Єдаїного Натанаїл.
NEH|12|22|Левити, голови батьківських родів, були записані за днів Ел'яшіва, Йояди, і Йоханана, і Яддуя, а священики за царювання Дарія перського.
NEH|12|23|Сини Левія, голови батьківських родів, записані в Книгу Хронік, і аж до днів Йоханана, сина Ел'яшівового.
NEH|12|24|А голови Левитів: Хашавія, Шеревія, і Ісус, син Кадміїлів, та брати їхні були навпроти них, щоб хвалити та славити за наказом Давида, Божого чоловіка, черга за чергою.
NEH|12|25|Матанія, і Бакбукія, Овадія, Мешуллам, Талмон, Аккув, придверні, сторожа в брамних складах.
NEH|12|26|Вони були за днів Йоякима, сина Ісуса, сина Йоцадакового, та за днів намісника Неемії та священика вчителя Ездри.
NEH|12|27|А в свято освячення єрусалимського муру шукали Левитів по всіх їхніх місцях, щоб привести їх до Єрусалиму справити свято освячення та радости з похвалами, із піснею, цимбалами, арфами та з цитрами.
NEH|12|28|І позбиралися сини співаків та з округи навколо Єрусалиму та з осель нетофатян,
NEH|12|29|і з Бет-Гаґґілґала, і з піль Ґеви та Азмавету, бо співаки побудували собі двори навколо Єрусалиму.
NEH|12|30|І очистилися священики та Левити, і вони очистили народ, і брами та мур.
NEH|12|31|І повводив я Юдиних зверхників на мур, і поставив два великі збори славословників та походи, з них один пішов праворуч по муру до Смітникової брами.
NEH|12|32|А за ними йшов Гошая та половина Юдиних зверхників,
NEH|12|33|і Азарія, Ездра, і Мешуллам,
NEH|12|34|Юда, і Веніямин, Шемая, і Ірмея.
NEH|12|35|А з священичих синів із сурмами: Захарій, син Йонатана, сина Шемаї, сина Маттанії, сина Міхаї, сина Заккура, сина Асафового,
NEH|12|36|а брати його: Шемая, і Азаріїл, Мілай, Ґілалай, Маай, Натанаїл, і Юда, Ханані з музичними знаряддями Давида, Божого чоловіка, а вчитель Ездра перед ними.
NEH|12|37|А при Джерельній брамі, навпроти них, вони йшли ступенями Давидового Міста, входом на стіну над Давидовим домом і аж до Водної брами на схід.
NEH|12|38|А другий збір славословників ішов ліворуч, а за ним я та половина народу, зверху по муру вище башти Печей та аж до Широкого муру,
NEH|12|39|і від Єфремової брами та до брами Старої, і до брами Рибної, і башти Ханан'їла, і башти Меа, і аж до брами Овечої, і спинилися біля брами Ув'язнення.
NEH|12|40|І стали обидва збори славословників біля Божого дому, і я, і половина заступників зо мною,
NEH|12|41|і священики: Ел'яким, Маасея, Мін'ямин, Міхая, Елйоенай, Захарій, Хананія з сурмами,
NEH|12|42|і Маасея, і Шемая, і Елеазар, і Уззі, і Єгоханан, і Малкійя, і Елам, і Езер. І співаки співали, а Їзрахія був провідником.
NEH|12|43|І вони приносили того дня великі жертви та раділи, бо Бог порадував їх великою радістю. І раділи також жінки та діти, і аж далеко чута була радість Єрусалиму!
NEH|12|44|І того дня були попризначувані люди над коморами для скарбів, для приношень, для первоплодів та для десятин, щоб зносити в них з міських піль законні частки священикам та Левитам, бо радість Юдеї була дивитися на священиків та на Левитів, що стояли!
NEH|12|45|І вони стерегли постанови свого Бога, і постанови про очищення, і були співаками та придверними за наказом Давида та сина його Соломона.
NEH|12|46|Бо віддавна, за днів Давида та Асафа, були голови співаків та пісні хвали й збори славословників для Бога.
NEH|12|47|І ввесь Ізраїль за днів Зоровавеля та за днів Неемії давав частки співацькі та придверничі, щодня належне, і освячував це Левитам, а Левити освячували Аароновим синам.
NEH|13|1|Того дня читане було з Мойсеєвої книги вголос народу, і було знайдене написане в ній, що Аммонітянин та Моавітянин не ввійде до Божої громади, і так буде аж навіки,
NEH|13|2|бо вони не стріли були Ізраїлевих синів хлібом та водою, і найняли були на нього Валаама проклясти його, та Бог наш обернув те прокляття на благословення.
NEH|13|3|І сталося, як почули вони Закон, то відділили від Ізраїля все чуже.
NEH|13|4|А перед тим священик Ел'яшів, призначений до комори дому нашого Бога, близький Товійїн,
NEH|13|5|то зробив йому велику комору, а туди давали колись жертву хлібну, ладан, і посуд, і десятину збіжжя, молоде вино та оливу, призначені заповіддю для Левитів, і співаків, і придверних, і священичі принесення.
NEH|13|6|А за ввесь цей час не був я в Єрусалимі, бо в тридцять другому році Артаксеркса, царя вавилонського, я прийшов був до царя, та по певному часі випросився я від царя.
NEH|13|7|І прийшов я до Єрусалиму, і розглянувся в тому злі, що зробив Єл'яшів Товійї, роблячи йому комору на подвір'ях Божого дому.
NEH|13|8|І було мені дуже зле, й я всі домашні Товійїні речі повикидав геть із комори.
NEH|13|9|І я сказав, і очистили комори, а я вернув туди посуд Божого дому, хлібну жертву та ладан.
NEH|13|10|І довідався я, що левитські частки не давалися, а вони повтікали кожен на поле своє, ті Левити та співаки, що робили свою працю.
NEH|13|11|І докоряв я заступникам та й сказав: Чого опущений дім Божий? І зібрав я їх, і поставив їх на їхніх місцях.
NEH|13|12|І вся Юдея приносила десятину збіжжя, і молодого вина, і оливи до скарбниць.
NEH|13|13|І настановив я над скарбницями священика Шелемію й книжника Садока та Педаю з Левитів, а на їхню руку Ханана, сина Заккура, сина Маттаніїного, бо вони були уважані за вірних. І на них покладено ділити частки для їхніх братів.
NEH|13|14|Пам'ятай же мене, Боже, за це, і не зітри моїх добродійств, які я зробив у Божому домі та в сторожах!
NEH|13|15|Тими днями бачив я в Юдеї таких, що топтали в суботу чавила, і носили снопи, і нав'ючували на ослів вино, виноград, і фіґі, і всілякий тягар, і везли до Єрусалиму суботнього дня. І я при свідках остеріг їх того дня, коли вони продавали живність.
NEH|13|16|А тиряни мешкали в ньому, і постачали рибу й усе на продаж, і продавали в суботу Юдиним синам та в Єрусалимі.
NEH|13|17|І докоряв я Юдиним шляхетним та й сказав їм: Що це за річ, яку ви робите, і безчестите суботній день?
NEH|13|18|Чи ж не так робили ваші батьки, а наш Бог спровадив усе це зло на нас та на це місто? А ви побільшуєте жар гніву на Ізраїля зневажанням суботи.
NEH|13|19|І бувало, як падала вечерова тінь на єрусалимські брами перед суботою, то я наказував, і були замикувані брами. І звелів я, щоб не відчиняли їх, а тільки аж по суботі. А біля брам я поставив слуг своїх, щоб тягар не входив суботнього дня!
NEH|13|20|І ночували крамарі та продавці всього продажного раз і два поза Єрусалимом.
NEH|13|21|І остеріг я їх при свідках та й сказав їм: Чого ви ночуєте навпроти муру? Якщо ви повторите це, я простягну руку на вас! Від того часу вони не приходили в суботу.
NEH|13|22|І сказав я Левитам, щоб вони очистилися й приходили стерегти брами, щоб освятити суботній день. Також це запам'ятай мені, Боже мій, і змилуйся надо мною за великістю милости Твоєї!
NEH|13|23|Тими днями бачив я також юдеїв, що брали собі за жінок ашдодянок, аммонітянок, моавітянок.
NEH|13|24|А їхні сини говорили наполовину по-ашдодському, і не вміли говорити по-юдейському, а говорили мовою того чи того народу.
NEH|13|25|І докоряв я їм, і проклинав їх, і бив декого з них, і рвав їм волосся, і заприсягав їх Богом, кажучи: Не давайте ваших дочок їхнім синам, і не беріть їхніх дочок для ваших синів та для вас.
NEH|13|26|Чи ж не цим згрішив був Соломон, Ізраїлів цар, а між багатьма народами не було такого царя, як він, і був уподобаний Богові своєму, і Бог настановив його царем над усім Ізраїлем, і його ввели в гріх ті чужі жінки?
NEH|13|27|І тому чи ж чуте було таке, щоб чинити все це велике лихо на спроневірення проти нашого Бога, щоб брати чужих жінок?
NEH|13|28|А один із синів Йояди, сина Ел'яшіва, великого священика, був зятем хоронянина Санваллата, і я вигнав його від себе!
NEH|13|29|Запам'ятай же їм, Боже мій, за сплямлення священства та заповіту священичого та левитського!
NEH|13|30|І очистив я їх від усього чужого, і встановив черги для священиків та для Левитів, кожного в службі їх,
NEH|13|31|і для пожертви дров в означених часах, і для первоплодів. Запам'ятай же мене, боже мій, на добро!
