JOB|1|1|Vir erat in terra Us nomine Iob, et erat vir ille simplex et rectus ac timens Deum et recedens a malo.
JOB|1|2|Natique sunt ei septem filii et tres filiae.
JOB|1|3|Et fuit possessio eius septem milia ovium et tria milia camelorum, quingenta quoque iuga boum et quingentae asinae ac familia multa nimis; eratque vir ille magnus inter omnes Orientales.
JOB|1|4|Et ibant filii eius et faciebant convivium per domos unusquisque in die suo; et mittentes vocabant tres sorores suas, ut comederent et biberent cum eis.
JOB|1|5|Cumque in orbem transissent dies convivii, mittebat ad eos Iob et sanctificabat illos; consurgensque diluculo offerebat holocausta pro singulis. Dicebat enim: " Ne forte peccaverint filii mei et benedixerint Deo in cordibus suis ". Sic faciebat Iob cunctis diebus.
JOB|1|6|Quadam autem die, cum venissent filii Dei, ut assisterent coram Domino, affuit inter eos etiam Satan.
JOB|1|7|Cui dixit Dominus: " Unde venis? ". Qui respondens ait: " Circuivi terram et perambulavi eam ".
JOB|1|8|Dixitque Dominus ad eum: " Numquid considerasti servum meum Iob, quod non sit ei similis in terra, homo simplex et rectus ac timens Deum et recedens a malo? ".
JOB|1|9|Cui respondens Satan ait: " Numquid Iob frustra timet Deum?
JOB|1|10|Nonne tu vallasti eum ac domum eius universamque substantiam per circuitum, operibus manuum eius benedixisti, et possessio eius crevit in terra?
JOB|1|11|Sed extende paululum manum tuam et tange cuncta, quae possidet, nisi in faciem benedixerit tibi ".
JOB|1|12|Dixit ergo Dominus ad Satan: " Ecce, universa, quae habet, in manu tua sunt; tantum in eum ne extendas manum tuam ". Egressusque est Satan a facie Domini.
JOB|1|13|Cum autem quadam die filii et filiae eius comederent et biberent vinum in domo fratris sui primogeniti,
JOB|1|14|nuntius venit ad Iob, qui diceret: " Boves arabant, et asinae pascebantur iuxta eos;
JOB|1|15|et irruerunt Sabaei tuleruntque eos et pueros percusserunt gladio, et evasi ego solus, ut nuntiarem tibi ".
JOB|1|16|Cumque adhuc ille loqueretur, venit alter et dixit: " Ignis Dei cecidit e caelo et ussit oves puerosque consumpsit, et effugi ego solus, ut nuntiarem tibi ".
JOB|1|17|Sed et illo adhuc loquente, venit alius et dixit: " Chaldaei fecerunt tres turmas et invaserunt camelos et tulerunt eos necnon et pueros percusserunt gladio, et ego fugi solus, ut nuntiarem tibi ".
JOB|1|18|Adhuc loquebatur ille, et ecce alius intravit et dixit: " Filiis tuis et filiabus vescentibus et bibentibus vinum in domo fratris sui primogeniti,
JOB|1|19|repente ventus vehemens irruit a regione deserti et concussit quattuor angulos domus; quae corruens oppressit liberos tuos, et mortui sunt, et effugi ego solus, ut nuntiarem tibi ".
JOB|1|20|Tunc surrexit Iob et scidit vestimenta sua et, tonso capite, corruens in terram adoravit
JOB|1|21|et dixit: Nudus egressus sum de utero matris meaeet nudus revertar illuc.Dominus dedit, Dominus abstulit; sicut Domino placuit, ita factum est:sit nomen Domini benedictum ".
JOB|1|22|In omnibus his non peccavit Iob labiis suis neque stultum quid contra Deum locutus est.
JOB|2|1|Factum est autem, cum quadam die venissent filii Dei, ut starent coram Domino, venit quoque Satan inter eos, ut staret in conspectu eius.
JOB|2|2|Dixit Dominus ad Satan: " Unde venis? ". Qui respondens ait: " Circuivi terram et perambulavi eam ".
JOB|2|3|Et dixit Dominus ad Satan: " Numquid considerasti servum meum Iob, quod non sit ei similis in terra, vir simplex et rectus ac timens Deum et recedens a malo et adhuc retinens innocentiam? Tu autem commovisti me adversus eum, ut affligerem eum frustra ".
JOB|2|4|Cui respondens Satan ait: " Pellem pro pelle et cuncta, quae habet, homo dabit pro anima sua.
JOB|2|5|Alioquin mitte manum tuam et tange os eius et carnem; et tunc videbis, si in faciem benedicet tibi ".
JOB|2|6|Dixit ergo Dominus ad Satan: " Ecce, in manu tua est; verumtamen animam illius serva ".
JOB|2|7|Egressus igitur Satan a facie Domini, percussit Iob ulcere pessimo a planta pedis usque ad verticem eius.
JOB|2|8|Qui testa saniem radebat, sedens in sterquilinio.
JOB|2|9|Dixit autem illi uxor sua: Adhuctu permanes in simplicitate tua?Benedic Deo et morere ".
JOB|2|10|Qui ait ad illam: Quasi una de stultis mulieribuslocuta es!Si bona suscepimus de manu Dei,mala quare non suscipiamus? ".In omnibus his non peccavit Iob labiis suis.
JOB|2|11|Igitur, audientes tres amici Iob omne malum, quod accidisset ei, venerunt singuli de loco suo, Eliphaz Themanites et Baldad Suhites et Sophar Naamathites. Condixerant enim, ut pariter venientes visitarent eum et consolarentur.
JOB|2|12|Cumque elevassent procul oculos suos, non cognoverunt eum et exclamantes ploraverunt; scissisque vestibus, sparserunt pulverem super caput suum in caelum.
JOB|2|13|Et sederunt cum eo in terra septem diebus et septem noctibus, et nemo loquebatur ei verbum; videbant enim dolorem esse vehementem.
JOB|3|1|Post haec aperuit Iob os suum et maledixit diei suo
JOB|3|2|et locutus est:
JOB|3|3|" Pereat dies, in qua natus sum,et nox, in qua dictum est: "Conceptus est homo".
JOB|3|4|Dies ille vertatur in tenebras;non requirat eum Deus desuper,et non illustretur lumine.
JOB|3|5|Obscurent eum tenebrae et umbra mortis;occupet eum caligo,et involvatur amaritudine.
JOB|3|6|Noctem illam tenebrosus turbo possideat;non computetur in diebus anninec numeretur in mensibus.
JOB|3|7|Sit nox illa solitaria nec laude digna;
JOB|3|8|maledicant ei, qui maledicunt diei,qui parati sunt suscitare Leviathan.
JOB|3|9|Obtenebrentur stellae crepusculi eius;exspectet lucem, et non sit,nec videat palpebras aurorae,
JOB|3|10|quia non conclusit ostia ventris, qui portavit me,nec abstulit mala ab oculis meis.
JOB|3|11|Quare non in vulva mortuus sum?Egressus ex utero non statim perii?
JOB|3|12|Quare exceptus genibus?Cur lactatus uberibus?
JOB|3|13|Nunc enim dormiens sileremet somno meo requiescerem
JOB|3|14|cum regibus et consulibus terrae,qui aedificant sibi solitudines,
JOB|3|15|aut cum principibus, qui possident aurumet replent domos suas argento.
JOB|3|16|Aut sicut abortivum absconditum non subsisterem,vel qui concepti non viderunt lucem.
JOB|3|17|Ibi impii cessaverunt a tumultu,et ibi requieverunt fessi robore.
JOB|3|18|Et quondam vincti pariter sine molestianon audierunt vocem exactoris.
JOB|3|19|Parvus et magnus ibi sunt,et servus liber a domino suo.
JOB|3|20|Quare misero data est lux,et vita his, qui in amaritudine animae sunt?
JOB|3|21|Qui exspectant mortem, et non venit,et effodiunt quaerentes illam magis quam thesauros;
JOB|3|22|gaudentque vehementeret laetantur sepulcro.
JOB|3|23|Viro, cuius abscondita est via,et circumdedit eum Deus tenebris.
JOB|3|24|Antequam comedam, suspiro,et quasi inundantes aquae sic rugitus meus.
JOB|3|25|Quia timor, quem timebam, evenit mihi,et, quod verebar, accidit.
JOB|3|26|Non dissimulavi, non silui, non quievi,et venit super me indignatio ".
JOB|4|1|Respondens autem Eliphaz Themanites dixit:
JOB|4|2|" Si coeperimus loqui tibi, forsitan moleste accipies;sed conceptum sermonem tenere quis poterit?
JOB|4|3|Ecce, docuisti multoset manus lassas roborasti;
JOB|4|4|vacillantes confirmaverunt sermones tui,et genua trementia confortasti.
JOB|4|5|Nunc autem venit super te plaga, et defecisti;tetigit te, et conturbatus es.
JOB|4|6|Nonne timor tuus est fiducia tua,spes tua est perfectio viarum tuarum?
JOB|4|7|Recordare, obsecro te, quis umquam innocens periit,aut quando recti deleti sunt?
JOB|4|8|quin potius vidi eos, qui operantur iniquitatemet seminant dolores et metunt eos,
JOB|4|9|flante Deo perisse,et spiritu irae eius esse consumptos.
JOB|4|10|Rugitus leonis et vox leaenaeet dentes catulorum leonum contriti sunt.
JOB|4|11|Leo periit, eo quod non haberet praedam,et catuli leonis dissipati sunt.
JOB|4|12|Porro ad me furtive verbum delatum est,et suscepit auris mea sussurrum eius.
JOB|4|13|In horrore visionis nocturnae,quando solet sopor occupare homines,
JOB|4|14|pavor tenuit me et tremor,et omnia ossa mea perterrita sunt.
JOB|4|15|Et cum spiritus, me praesente, transiret,inhorruerunt pili carnis meae.
JOB|4|16|Stetit quidam, cuius non agnoscebam vultum,imago coram oculis meis,et vocem quasi aurae lenis audivi:
JOB|4|17|"Numquid homo Dei comparatione iustificabitur,aut factore suo purior erit vir?".
JOB|4|18|Ecce, in servis suis fiduciam non habetet in angelis suis reperit pravitatem.
JOB|4|19|Quanto magis hi, qui habitant domos luteas,quorum fundamentum est in pulvere.Consumentur velut tinea!
JOB|4|20|De mane usque ad vesperam succidenturet, quia nullus intellegit, in aeternum peribunt.
JOB|4|21|Nonne evulsum est reliquum eorum ab eis?Morientur, et non in sapientia.
JOB|5|1|Voca ergo, si est qui tibi re spondeat!Ad quem sanctorum converteris?
JOB|5|2|Vere stultum interficit iracundia,et fatuum occidit invidia.
JOB|5|3|Ego vidi stultum firma radiceet maledixi sedi eius statim.
JOB|5|4|Longe fient filii eius a saluteet conterentur in porta, et non erit qui eruat.
JOB|5|5|Cuius messem famelicus comedet,et ipsum rapiet armatus, et bibent sitientes divitias eius.
JOB|5|6|Quia non egreditur ex pulvere nequitia,et de humo non oritur dolor.
JOB|5|7|Sed homo generat laborem,et aves elevant volatum.
JOB|5|8|Quam ob rem ego deprecabor Dominumet ad Deum ponam eloquium meum,
JOB|5|9|qui facit magna et inscrutabiliaet mirabilia absque numero;
JOB|5|10|qui dat pluviam super faciem terraeet irrigat aquis rura;
JOB|5|11|qui ponit humiles in sublimeet maerentes erigit sospitate;
JOB|5|12|qui dissipat cogitationes malignorum,ne possint implere manus eorum, quod coeperant;
JOB|5|13|qui apprehendit sapientes in astutia eorumet consilium pravorum dissipat.
JOB|5|14|Per diem incurrent tenebraset, quasi in nocte, sic palpabunt in meridie.
JOB|5|15|Porro salvum faciet egenum a gladio oris eorumet de manu violenti pauperem;
JOB|5|16|et erit egeno spes,iniquitas autem contrahet os suum.
JOB|5|17|Beatus homo, qui corripitur a Deo;increpationem ergo Omnipotentis ne reprobes.
JOB|5|18|Quia ipse vulnerat et medetur,percutit, et manus eius sanabunt.
JOB|5|19|In sex tribulationibus liberabit te,et in septem non tanget te malum.
JOB|5|20|In fame eruet te de morteet in bello de manu gladii.
JOB|5|21|A flagello linguae absconderiset non timebis vastationem, cum venerit.
JOB|5|22|In vastitate et fame ridebiset bestias terrae non formidabis.
JOB|5|23|Sed cum lapidibus campi pactum tuum,et bestiae terrae pacificae erunt tibi.
JOB|5|24|Et scies quod pacem habeat tabernaculum tuum,et visitans habitationem tuam non falleris.
JOB|5|25|Scies quoque quoniam multiplex erit semen tuum,et progenies tua quasi herba terrae.
JOB|5|26|Ingredieris in abundantia sepulcrum,sicut infertur acervus tritici in tempore suo.
JOB|5|27|Ecce hoc, ut investigavimus, ita est;oboedi illi et tu sapias tibi ".
JOB|6|1|Respondens autem Iob dixit:
JOB|6|2|" Utinam appenderetur aegritu do mea,et calamitatem meam assumerent in statera!
JOB|6|3|Nunc vero arena maris haec gravior apparet,inde verbis meis haesito.
JOB|6|4|Quia sagittae Omnipotentis in me sunt,quarum venenum ebibit spiritus meus;et terrores Dei militant contra me.
JOB|6|5|Numquid rugiet onager, cum habuerit herbam?Aut mugiet bos, cum ante praesepe plenum steterit?
JOB|6|6|Aut poterit comedi insulsum, quod non est sale conditum?Aut poterit gustari herba insulsa?
JOB|6|7|Quae prius nolebat tangere anima mea,nunc prae angustia cibi mei sunt.
JOB|6|8|Quis det, ut veniat petitio mea,et, quod exspecto, tribuat mihi Deus?
JOB|6|9|Utinam Deus me conterat;solvat manum suam et succidat me!
JOB|6|10|Et haec mihi sit consolatio,et exsultabo vel in pavore, qui non parcat,nec celabo sermones Sancti.
JOB|6|11|Quae est enim fortitudo mea, ut sustineam?Aut quis finis meus, ut patienter agam?
JOB|6|12|Num fortitudo lapidum, fortitudo mea?Num caro mea aenea est?
JOB|6|13|An non est auxilium mihi in me,et virtus quoque remota est a me?
JOB|6|14|Qui tollit ab amico suo misericordiam,timorem Omnipotentis derelinquit.
JOB|6|15|Fratres mei mentiti sunt mesicut alveus torrentium, qui evanescunt
JOB|6|16|nigrescentes glacie,cum ingruit super eos nix.
JOB|6|17|Tempore, quo diffluunt, arescuntet, ut incaluerit, solvuntur de loco suo.
JOB|6|18|Deflectunt viatorum turmae de viis suis,ascendentes per desertum pereunt.
JOB|6|19|Commeatus Thema consideraverunt,viatores Saba speraverunt in eis.
JOB|6|20|Confusi sunt, quia speraverunt;venerunt eo usque, et pudore cooperti sunt.
JOB|6|21|Ita nunc vos facti estis mihi;videntes plagam meam, timetis.
JOB|6|22|Numquid dixi: Afferte mihiet de substantia vestra donate mihi?
JOB|6|23|vel: Liberate me de manu hostiset de manu robustorum eruite me?
JOB|6|24|Docete me, et ego tacebo,et, si quid forte ignoravi, instruite me.
JOB|6|25|Quare detraxistis sermonibus veritatis,cum e vobis nullus sit, qui possit arguere me?
JOB|6|26|Ad increpandum tantum eloquia concinnatis,sed in ventum verba desperati.
JOB|6|27|Super pupillum irruitiset subvertere nitimini amicum vestrum.
JOB|6|28|Nunc, quaeso, convertimini ad me,et in faciem vestram non mentiar.
JOB|6|29|Revertite! Nulla erit improbitas.Revertite! Adhuc praesens adest iustitia mea.
JOB|6|30|Estne in lingua mea improbitas?An palatum meum non discernit nequitiam?
JOB|7|1|Nonne militia est vita hominis super terram,et sicut dies mercennarii dies eius?
JOB|7|2|Sicut servus desiderat umbram,et sicut mercennarius praestolatur mercedem suam,
JOB|7|3|sic et ego habui menses vacuoset noctes laboriosas enumeravi mihi.
JOB|7|4|Si dormiero, dicam: Quando consurgam?Et rursum exspectabo vesperamet replebor doloribus usque crepusculum.
JOB|7|5|Induta est caro mea putredine et sordibus pulveris;cutis mea scinditur et diffluit.
JOB|7|6|Dies mei velocius transierunt quam navicula texentiset consumpti sunt deficiente filo.
JOB|7|7|Memento quia ventus est vita mea,et non revertetur oculus meus, ut videat bona.
JOB|7|8|Nec aspiciet me visus hominis;oculi tui in me, et non subsistam.
JOB|7|9|Sicut consumitur nubes et pertransit,sic, qui descenderit ad inferos, non ascendet
JOB|7|10|nec revertetur ultra in domum suam,neque cognoscet eum amplius locus eius.
JOB|7|11|Quapropter et ego non parcam ori meo;loquar in tribulatione spiritus mei, confabulabor cum amaritudine animae meae.
JOB|7|12|Numquid mare ego sum aut cetus,quia posuisti super me custodiam?
JOB|7|13|Si dixero: Consolabitur me lectulus meus,et assumet stratum meum querelam meam,
JOB|7|14|terrebis me per somniaet per visiones horrore concuties.
JOB|7|15|Quam ob rem eligit suspendium anima mea,et mortem ossa mea.
JOB|7|16|Desperavi; nequaquam ultra iam vivam.Parce mihi, nihil enim sunt dies mei.
JOB|7|17|Quid est homo, quia magnificas eum?Aut quid apponis erga eum cor tuum?
JOB|7|18|Visitas eum diluculoet singulis momentis probas illum.
JOB|7|19|Usquequo non avertes oculos a me?Nec dimittis me, ut glutiam salivam meam?
JOB|7|20|Peccavi; quid faciam tibi,o custos hominum?Quare posuisti me contrarium tibi, et factus sum mihimetipsi gravis?
JOB|7|21|Cur non tollis peccatum meumet quare non aufers iniquitatem meam?Ecce, nunc in pulvere dormiam;et, si mane me quaesieris, non subsistam! ".
JOB|8|1|Respondens autem Baldad Suhites dixit:
JOB|8|2|" Usquequo loqueris talia,et spiritus vehemens sermones oris tui?
JOB|8|3|Numquid Deus supplantat iudicium,aut Omnipotens subvertit, quod iustum est?
JOB|8|4|Et si filii tui peccaverunt ei,et dimisit eos in manu iniquitatis suae,
JOB|8|5|tu tamen, si diluculo consurrexeris ad Deumet Omnipotentem fueris deprecatus,
JOB|8|6|si mundus et rectus incesseris,statim evigilabit ad teet pacatum reddet habitaculum iustitiae tuae;
JOB|8|7|in tantum ut, si priora tua fuerint parva,et novissima tua multiplicentur nimis.
JOB|8|8|Interroga enim generationem pristinamet diligenter investiga patrum memoriam.
JOB|8|9|Hesterni quippe sumus et ignoramus,quoniam sicut umbra dies nostri sunt super terram.
JOB|8|10|Nonne ipsi docebunt te, loquentur tibiet de corde suo proferent eloquia?
JOB|8|11|Numquid virere potest scirpus absque umore,aut crescere carectum sine aqua?
JOB|8|12|Cum adhuc sit in flore, nec carpatur manu,ante omnes herbas arescit.
JOB|8|13|Sic viae omnium, qui obliviscuntur Deum,et spes impii peribit.
JOB|8|14|Cuius spes filum tenue,et sicut tela aranearum fiducia eius.
JOB|8|15|Innitetur super domum suam et non stabit;fulciet eam et non consurget.
JOB|8|16|Umectus videtur, antequam veniat sol,et in horto suo germen eius egredietur.
JOB|8|17|Super acervum petrarum radices eius densabuntur,et inter lapides commorabitur.
JOB|8|18|Si absorbuerit eum de loco suo,negabit eum et dicet: "Non novi te".
JOB|8|19|Haec est enim laetitia viae eius,ut rursum de terra alii germinentur.
JOB|8|20|Deus non proiciet simplicemnec porriget manum malignis,
JOB|8|21|donec impleatur risu os tuum,et labia tua iubilo.
JOB|8|22|Qui oderunt te, induentur confusione,et tabernaculum impiorum non subsistet ".
JOB|9|1|Et respondens Iob ait:
JOB|9|2|" Vere scio quod ita sit,et quomodo iustificabitur homo compositus Deo?
JOB|9|3|Si voluerit contendere cum eo,non poterit ei respondere unum pro mille.
JOB|9|4|Sapiens corde est et fortis robore;quis restitit ei, et pacem habuit?
JOB|9|5|Qui transtulit montes, et nescierunt hi, quos subvertit in furore suo.
JOB|9|6|Qui commovet terram de loco suo,et columnae eius concutiuntur.
JOB|9|7|Qui praecipit soli, et non oritur,et stellas claudit quasi sub signaculo.
JOB|9|8|Qui extendit caelos soluset graditur super fluctus maris.
JOB|9|9|Qui facit Arcturum et Orionaet Hyadas et interiora austri.
JOB|9|10|Qui facit magna et incomprehensibiliaet mirabilia, quorum non est numerus.
JOB|9|11|Si venerit ad me, non videbo eum;si abierit, non intellegam.
JOB|9|12|Si repente arripiet, quis eum impediet?Vel quis dicere potest: "Quid facis?".
JOB|9|13|Deus non retinet iram suam,et sub eo curvantur auxilia Rahab.
JOB|9|14|Quantus ergo sum ego, ut respondeam eiet loquar delectis verbis cum eo?
JOB|9|15|Quia, etiamsi iustus essem, non responderem,sed meum iudicem deprecarer;
JOB|9|16|et, cum invocantem exaudierit me,non credam quod audierit vocem meam.
JOB|9|17|In turbine enim conteret meet multiplicabit vulnera mea etiam sine causa.
JOB|9|18|Non concedit requiescere spiritum meumet implet me amaritudinibus.
JOB|9|19|Si fortitudo quaeritur, robustissimus est;si iudicium, quis eum arcesserit?
JOB|9|20|Si iustificare me voluero, os meum condemnabit me;si innocentem ostendero, pravum me comprobabit.
JOB|9|21|Etiamsi simplex fuero, hoc ipsum ignorabit anima mea,et contemnam vitam meam.
JOB|9|22|Unum est, quod locutus sum:Et innocentem et impium ipse consumit.
JOB|9|23|Si subito flagellum occidat,de afflictione innocentium ridebit.
JOB|9|24|Terra data est in manus impii,vultum iudicum eius operit;quod si non ille est, quis ergo est?
JOB|9|25|Dies mei velociores fuerunt cursore:fugerunt et non viderunt bonum;
JOB|9|26|pertransierunt quasi naves arundineae,sicut aquila volans ad escam.
JOB|9|27|Cum dixero: Obliviscar maerorem meum,commutabo faciem meam et hilaris fiam,
JOB|9|28|vereor omnes dolores meos,sciens quod non iustificaveris me.
JOB|9|29|Si autem et sic impius sum,quare frustra laboravi?
JOB|9|30|Si lotus fuero quasi aquis nivis,et lixivo mundavero manus meas,
JOB|9|31|tamen sordibus intinges me,et abominabuntur me vestimenta mea.
JOB|9|32|Neque enim viro, qui similis mei est, respondebo;nec vir, quocum in iudicio contendam.
JOB|9|33|Non est qui utrumque valeat arguereet ponere manum suam in ambobus.
JOB|9|34|Auferat a me virgam suam,et pavor eius non me terreat.
JOB|9|35|Loquar et non timebo eum;quia sic non mecum ipse sum.
JOB|10|1|Taedet animam meam vitae meae;dimittam adversum me eloquium meum,loquar in amaritudine animae meae.
JOB|10|2|Dicam Deo: Noli me condemnare,indica mihi cur me ita iudices.
JOB|10|3|Numquid bonum tibi videtur, si opprimas meet calumnieris me, opus manuum tuarum,et super consilium impiorum arrideas?
JOB|10|4|Numquid oculi carnei tibi sunt,aut, sicut videt homo, et tu videbis?
JOB|10|5|Numquid sicut dies hominis dies tui,et anni tui sicut humana sunt tempora,
JOB|10|6|ut quaeras iniquitatem meamet peccatum meum scruteris,
JOB|10|7|cum scias quia nihil impium fecerim,et sit nemo, qui de manu tua possit eruere?
JOB|10|8|Manus tuae fecerunt meet plasmaverunt me totum in circuitu;et sic repente praecipitas me?
JOB|10|9|Memento, quaeso, quod sicut lutum feceris meet in pulverem reduces me.
JOB|10|10|Nonne sicut lac mulsisti meet sicut caseum me coagulasti?
JOB|10|11|Pelle et carnibus vestisti me;ossibus et nervis compegisti me.
JOB|10|12|Vitam et misericordiam tribuisti mihi,et visitatio tua custodivit spiritum meum.
JOB|10|13|Licet haec celes in corde tuo,tamen scio haec in animo tuo versari.
JOB|10|14|Si peccaverim, observas meet ab iniquitate mea mundum me esse non pateris.
JOB|10|15|Et si impius fuero, vae mihi est;et si iustus, non levabo caput,saturatus afflictione et miseria.
JOB|10|16|Si superbia extollar, quasi catulum leonis capies meet iterum mirabilem te exhibebis in me.
JOB|10|17|Instauras testes tuos contra meet multiplicas iram tuam adversum me,et poenae militant in me.
JOB|10|18|Quare de vulva eduxisti me?Qui utinam consumptus essem, ne oculus me videret!
JOB|10|19|Fuissem quasi non essem,de utero translatus ad tumulum.
JOB|10|20|Numquid non paucitas dierum meorum finietur brevi?Dimitte ergo me, ut refrigerem paululum dolorem meum,
JOB|10|21|antequam vadam, et non revertar,ad terram tenebrarum et umbrae mortis,
JOB|10|22|terram caliginis et tenebrarum,ubi umbra mortis et nullus ordo,sed sempiternus horror inhabitat ".
JOB|11|1|Respondens autem Sophar Naamathites dixit:
JOB|11|2|" Numquid illi, qui multa loquitur, non et respondetur?Aut vir verbosus iustificabitur?
JOB|11|3|Vaniloquium tuum viros tacere faciet,et, cum ceteros irriseris, a nullo confutaberis?
JOB|11|4|Dixisti enim: "Purus est sermo meus,et mundus sum in conspectu tuo".
JOB|11|5|Atque utinam Deus ipse loqueretur tecumet aperiret labia sua tibi,
JOB|11|6|ut ostenderet tibi secreta sapientiaeet arcana consilia eius,et intellegeres quod multo minora quaerat a te,quam meretur iniquitas tua.
JOB|11|7|Forsitan vestigia Dei comprehendeset usque ad perfectum Omnipotentem reperies?
JOB|11|8|Excelsior caelo est, et quid facies?Profundior inferno, et quid cognosces?
JOB|11|9|Longior terra mensura eiuset latior mari.
JOB|11|10|Si subverterit vel concluserit et coarctaverit,quis contradicet ei?
JOB|11|11|Ipse enim novit hominum vanitatem;et videns iniquitatem nonne considerat?
JOB|11|12|Sed et vir vacuus cordatus fit,et homo tamquam pullum onagri nascitur.
JOB|11|13|Tu autem, si cor tuum firmaveriset expanderis ad eum manus tuas,
JOB|11|14|si iniquitatem, quae est in manu tua, abstuleris a te,et non manserit in tabernaculo tuo iniustitia,
JOB|11|15|tunc levare poteris faciem tuam absque maculaet eris stabilis et non timebis.
JOB|11|16|Miseriae quoque oblivisceriset quasi aquarum, quae praeterierunt, recordaberis.
JOB|11|17|Et quasi meridianus fulgor consurget tibi ad vesperam,et, cum te caligine tectum putaveris, orieris ut lucifer.
JOB|11|18|Et habebis fiduciam, proposita tibi spe,et defossus securus dormies.
JOB|11|19|Requiesces, et non erit qui te exterreat;et deprecabuntur faciem tuam plurimi.
JOB|11|20|Oculi autem impiorum deficient,et effugium peribit ab eis;et spes illorum exhalatio animae ".
JOB|12|1|Respondens autem Iob dixit:
JOB|12|2|" Ergo vos estis soli homines,et vobiscum morietur sapientia.
JOB|12|3|Et mihi est cor sicut et vobis,nec inferior vestri sum;quis enim haec, quae nostis, ignorat?
JOB|12|4|Qui deridetur ab amico suo sicut ego,invocabit Deum, et exaudiet eum; deridetur enim iusti integritas.
JOB|12|5|Lampas contempta apud cogitationes eorum, qui securi sunt,parata iis, qui vacillant pede.
JOB|12|6|Tranquilla sunt tabernacula praedonumet secura iis, qui provocant Deum, iis, qui Deum tenent manu sua.
JOB|12|7|Nimirum interroga iumenta, et docebunt te,et volatilia caeli, et indicabunt tibi.
JOB|12|8|Loquere terrae, et docebit te;et narrabunt pisces maris.
JOB|12|9|Quis ignorat in omnibus hisquod manus Domini hoc fecerit?
JOB|12|10|In cuius manu anima omnis viventiset spiritus universae carnis hominis.
JOB|12|11|Nonne auris verba diiudicat,et palatum cibum sibi gustat?
JOB|12|12|In senibus est sapientia,et in longaevis prudentia.
JOB|12|13|Apud ipsum est sapientia et fortitudo;ipse habet consilium et intellegentiam.
JOB|12|14|Si destruxerit, nemo est, qui aedificet;si incluserit hominem, nullus est, qui aperiat.
JOB|12|15|Si continuerit aquas, arescent;et, si emiserit eas, subvertent terram.
JOB|12|16|Apud ipsum est fortitudo et sapientia;ipse novit et decipientem et eum qui decipitur.
JOB|12|17|Inducit consiliarios spoliatoset iudices in stuporem.
JOB|12|18|Balteum regum dissolvitet praecingit fune renes eorum.
JOB|12|19|Inducit sacerdotes spoliatoset optimates supplantat,
JOB|12|20|commutans labium veraciumet doctrinam senum auferens.
JOB|12|21|Effundit despectionem super principeset cingulum fortium relaxat.
JOB|12|22|Qui revelat profunda de tenebriset producit in lucem umbram mortis.
JOB|12|23|Qui multiplicat gentes et perdit easet subversas in integrum restituit.
JOB|12|24|Qui immutat cor principum populi terrae et decipit eoset errare eos faciet per invium desertum.
JOB|12|25|Palpabunt quasi in tenebris et non in luce,et errare eos faciet quasi ebrios.
JOB|13|1|Ecce, omnia haec vidit oculus meus,et audivit auris mea, et intellexi singula.
JOB|13|2|Secundum scientiam vestram, et ego novi;nec inferior vestri sum.
JOB|13|3|Sed tamen ad Omnipotentem loquaret disputare cum Deo cupio;
JOB|13|4|vos autem ostendam fabricatores mendacii,medicos vanos vos omnes.
JOB|13|5|Atque utinam taceretis,ut sit vobis in sapientiam!
JOB|13|6|Audite ergo correptionem meamet contentiones labiorum meorum attendite.
JOB|13|7|Numquid pro Deo profertis mendaciumet pro illo loquimini dolos?
JOB|13|8|Numquid faciem eius accipitiset pro Deo in iudicio contendere nitimini?
JOB|13|9|Aut bonum est quod vos excutiat?Aut, ut illuditur homini, illudetis ei?
JOB|13|10|Ipse vos arguet,cum in abscondito faciem accipitis.
JOB|13|11|Nonne maiestas eius turbabit vos,et terror eius irruet super vos?
JOB|13|12|Sententiae vestrae sunt proverbia cineris;thoraces lutei thoraces vestri.
JOB|13|13|Tacete paulisper, ut loquar ipse,et transeat super me quodcumque.
JOB|13|14|Quare sumam carnes meas dentibus meiset animam meam ponam in manibus meis?
JOB|13|15|Etiamsi occiderit me, in ipso sperabo; verumtamen vias meas in conspectu eius arguam.
JOB|13|16|Et hoc erit salus mea:non enim veniet in conspectu eius omnis impius.
JOB|13|17|Audite sermonem meumet explicationem meam percipite auribus vestris.
JOB|13|18|Ecce iudicium paravi;scio quod iustus inveniar.
JOB|13|19|Quis est qui contendat mecum?Tunc enim tacebo et consummabor.
JOB|13|20|Duo tantum ne facias mihi,et tunc a facie tua non abscondar:
JOB|13|21|Manum tuam longe fac a me,et formido tua non me terreat.
JOB|13|22|Voca me, et ego respondebo tibi;aut ipse loquar, et tu respondebis mihi.
JOB|13|23|Quantas habeo iniquitates et peccata?Scelera mea et delicta ostende mihi.
JOB|13|24|Cur faciem tuam abscondiset arbitraris me inimicum tuum?
JOB|13|25|Contra folium, quod vento rapitur, dure agiset stipulam siccam persequeris.
JOB|13|26|Scribis enim contra me amaritudineset occupatum me vis peccatis adulescentiae meae.
JOB|13|27|Posuisti in nervo pedem meumet observasti omnes semitas measet vestigia pedum meorum considerasti.
JOB|13|28|Qui quasi uter consumendus sum,et quasi vestimentum, quod comeditur a tinea.
JOB|14|1|Homo natus de muliere,brevi vivens tempore, commotione satiatur.
JOB|14|2|Qui quasi flos egreditur et arescitet fugit velut umbra et non permanet.
JOB|14|3|Et dignum ducis super huiuscemodi aperire oculos tuoset adducere eum tecum in iudicium?
JOB|14|4|Quis potest facere mundum de immundo?Ne unus quidem!
JOB|14|5|Si statuti dies hominis sunt,et numerus mensium eius apud te est,et constituti sunt termini eius, quos non praeteribit,
JOB|14|6|averte oculos tuos ab eo, ut quiescat,donec solvat, sicut mercennarius, dies suos.
JOB|14|7|Nam lignum habet spem;si praecisum fuerit, rursum virescet,et rami eius non deficient.
JOB|14|8|Si senuerit in terra radix eius,et in pulvere emortuus fuerit truncus illius,
JOB|14|9|ad odorem aquae germinabitet faciet comam quasi novellae.
JOB|14|10|Homo vero cum mortuus fuerit et debilitatur,exspirat homo et, ubi, quaeso, est?
JOB|14|11|Recedent aquae de mari,et fluvius vacuefactus arescet;
JOB|14|12|sic homo, cum dormierit, non resurget:donec atteratur caelum, non evigilabitnec consurget de somno suo.
JOB|14|13|Quis mihi hoc tribuat, ut in inferno seponas meet abscondas me, donec pertranseat furor tuus,et constituas mihi tempus, in quo recorderis mei?
JOB|14|14|Putasne mortuus homo rursum vivat?Cunctis diebus, quibus nunc milito,exspectarem, donec veniat immutatio mea.
JOB|14|15|Vocares me, et ego responderem tibi;opus manuum tuarum requireres.
JOB|14|16|Tu quidem nunc gressus meos dinumerares,sed parceres peccatis meis.
JOB|14|17|Signares quasi in sacculo delicta mea,sed dealbares iniquitatem meam.
JOB|14|18|Mons cadens decidit,et saxum transfertur de loco suo;
JOB|14|19|lapides excavant aquae,et alluvione terra inundatur:et spem hominis perdes.
JOB|14|20|Praevales adversus eum, et in perpetuum transiet;immutas faciem eius et emittis eum.
JOB|14|21|Sive nobiles fuerint filii eius, non novit;sive ignobiles, non intellegit.
JOB|14|22|Attamen caro eius, dum vivet, dolet,et anima illius super semetipso luget ".
JOB|15|1|Respondens autem Eliphaz Themanites dixit:
JOB|15|2|" Numquid sapiens respondebit sapientia ventosaet implebit vento urente stomachum suum?
JOB|15|3|Arguens verbis, quae nihil prosunt,et sententiis, quae nihil iuvant?
JOB|15|4|Tu autem pietatem dissolviset detrahis meditationi coram Deo.
JOB|15|5|Docet enim iniquitas tua os tuum,et assumis linguam callidorum.
JOB|15|6|Condemnabit te os tuum et non ego,et labia tua respondebunt tibi.
JOB|15|7|Numquid primus homo tu natus eset ante colles formatus?
JOB|15|8|Numquid consilium Dei audistiet tibi attrahis sapientiam?
JOB|15|9|Quid nosti, quod nos ignoremus?Quid intellegis, quod nos nesciamus?
JOB|15|10|Et senes et antiqui sunt inter nos,multo vetustiores quam pater tuus.
JOB|15|11|Numquid parum tibi sunt consolationes Dei?Et verbum lene tecum factum?
JOB|15|12|Quid te elevat cor tuum,et cur attonitos habes oculos?
JOB|15|13|Quid vertis contra Deum spiritum tuumet profers de ore tuo huiuscemodi sermones?
JOB|15|14|Quid est homo, ut immaculatus sit,et ut iustus appareat natus de muliere?
JOB|15|15|Ecce, sanctis suis non fidit,et caeli non sunt mundi in conspectu eius;
JOB|15|16|quanto magis abominabilis et corruptus homo,qui bibit quasi aquam iniquitatem.
JOB|15|17|Ostendam tibi, audi me;quod vidi, narrabo tibi,
JOB|15|18|quod sapientes confitentur,et non celaverunt eos patres eorum:
JOB|15|19|quibus solis data est terra,et non transivit alienus per eos.
JOB|15|20|Cunctis diebus suis impius cruciatur,et numerus annorum incertus est tyranno.
JOB|15|21|Sonitus terroris semper in auribus illius,quasi, cum pax sit, vastator irruat in eum.
JOB|15|22|Non credit quod reverti possit de tenebris,cum sit destinatus gladio.
JOB|15|23|Cum se moverit ad quaerendum panem: "Ubinam?",novit quod paratus sit in manu eius tenebrarum dies.
JOB|15|24|Terrebit eum tribulatio et angustia,vallabit eum sicut regem, qui praeparatur ad proelium.
JOB|15|25|Tetendit enim adversus Deum manum suam,et contra Omnipotentem roboratus est.
JOB|15|26|Cucurrit adversus eum erecto collo,spisso scuto armatus.
JOB|15|27|Operuit faciem eius crassitudo,et de lateribus eius arvina dependet.
JOB|15|28|Habitavit in civitatibus desolatiset in domibus desertis, quae in tumulos sunt redactae.
JOB|15|29|Non ditabitur, nec perseverabit substantia eius;nec mittet in terra radicem suam.
JOB|15|30|Non recedet de tenebris;ramos eius arefaciet flamma,et auferet ventus florem eius.
JOB|15|31|Ne credat vanitati errore deceptus,quia vanitas erit remuneratio eius.
JOB|15|32|Antequam dies eius impleantur, abscindentur,et ramus eius non virescet.
JOB|15|33|Laedetur quasi vinea in primo flore botrus eius,et quasi oliva proiciens florem suum.
JOB|15|34|Cangregatio enim impii sterilis,et ignis devorabit tabernacula eorum, qui munera libenter accipiunt.
JOB|15|35|Concepit dolorem et peperit iniquitatem,et venter eius praeparat dolos.
JOB|16|1|Respondens autem Iob dixit:
JOB|16|2|" Audivi frequenter talia!onsolatores molesti omnes vos estis.
JOB|16|3|Numquid habebunt finem verba ventosa,aut quid te exacerbat, ut respondeas?
JOB|16|4|Poteram et ego similia vestri loqui,si esset anima vestra pro anima mea!Concinnarem super vos sermoneset moverem caput meum super vos.
JOB|16|5|Roborarem vos ore meoet motum labiorum meorum non cohiberem.
JOB|16|6|Si locutus fuero, non quiescet dolor meuset, si tacuero, non recedet a me;
JOB|16|7|nunc autem defatigavit me dolor meus,et tu vastasti omnem coetum meum.
JOB|16|8|Rugae meae testimonium dicunt contra me;et suscitatur falsiloquus adversus faciem meam contradicens mihi,
JOB|16|9|Ira eius discerpsit me et adversata est mihi,et infremuit contra me dentibus suis.Hostis meus acuit oculos suos in me.
JOB|16|10|Aperuerunt super me ora suaet exprobrantes percusserunt maxillam meam,simul conferti contra me.
JOB|16|11|Concludit me Deus apud iniquumet manibus impiorum me tradit.
JOB|16|12|Ego, ille quondam tranquillus, repente contritus sum.Tenuit cervicem meam, confregit meet posuit me sibi quasi in signum.
JOB|16|13|Circumdedit me lanceis suis,scidit lumbos meos, non pepercitet effudit in terra iecur meum.
JOB|16|14|Dirupit me rumpens et diruens,irruit in me quasi gigas.
JOB|16|15|Saccum consui super cutem meamet dimisi in terram cornu meum.
JOB|16|16|Facies mea rubuit a fletu,et palpebrae meae caligaverunt;
JOB|16|17|attamen absque iniquitate manus meae,cum haberem mundas preces.
JOB|16|18|Terra, ne operias sanguinem meum,neque inveniat in te locum latendi clamor meus.
JOB|16|19|Ecce enim in caelo testis meus,et conscius meus in excelsis.
JOB|16|20|Interpretes mei sunt cogitationes meae:ad Deum stillat oculus meus.
JOB|16|21|Atque utinam sic iudicaretur vir cum Deo,sicut iudicatur filius hominis cum collega suo.
JOB|16|22|Ecce enim breves anni transeunt,et semitam, per quam non revertar, ambulo.
JOB|17|1|Spiritus meus attenuatus est,dies mei exstincti,et solum mihi superest sepulcrum.
JOB|17|2|Nonne irrisiones circumdant me,et in amaritudinibus moratur oculus meus?
JOB|17|3|Pone pignus pro me iuxta te;et quis umquam spondens percutiet manum meam?
JOB|17|4|Cor eorum longe fecisti a disciplina;propterea non exaltabuntur.
JOB|17|5|Praedam pollicetur sociis,sed oculi filiorum eius deficient.
JOB|17|6|Posuit me quasi in proverbium vulgiet conspuendum in faciem.
JOB|17|7|Caligavit ab indignatione oculus meus,et membra mea quasi in umbram redacta sunt.
JOB|17|8|Stupebunt iusti super hoc,et innocens contra impium excitabitur.
JOB|17|9|Et tenebit iustus viam suam,et mundus manibus addet fortitudinem.
JOB|17|10|Igitur omnes vos convertimini et venite,et non inveniam in vobis ullum sapientem.
JOB|17|11|Dies mei transierunt, cogitationes meae dissipatae suntet desideria cordis mei.
JOB|17|12|Noctem verterunt in diem;et rursum post tenebras properat lux.
JOB|17|13|Si sustinuero, infernus domus mea est;et in tenebris stravi lectulum meum.
JOB|17|14|Putredini dixi: Pater meus es!;Mater mea et soror mea! vermibus.
JOB|17|15|Ubi est ergo nunc praestolatio mea,et patientiam meam quis considerat?
JOB|17|16|In profundissimum infernum descendent omnia mea;simul in pulvere erit requies mihi? ".
JOB|18|1|Respondens autem Baldad Suhites dixit:
JOB|18|2|" Usque ad quem finem verba iactabitis?Intellegite prius, et sic loquamur.
JOB|18|3|Quare reputati sumus ut iumentaet sorduimus coram vobis?
JOB|18|4|Qui perdis animam tuam in furore tuo,numquid propter te derelinquetur terra,et transferentur rupes de loco suo?
JOB|18|5|Etenim lux impii exstinguetur,nec splendebit flamma ignis eius.
JOB|18|6|Lux obtenebrescet in tabernaculo illius,et lucerna, quae super eum est, exstinguetur.
JOB|18|7|Arctabuntur gressus virtutis eius,et praecipitabit eum consilium suum.
JOB|18|8|Immissi sunt in rete pedes eius,et in reticulo ambulat.
JOB|18|9|Tenet plantam illius laqueus,et firmatur super eum tendiculum.
JOB|18|10|Abscondita est in terra pedica eius,et decipula illius super semitam.
JOB|18|11|Undique terrent eum formidineset involvunt pedes eius.
JOB|18|12|Attenuatur fame robur eius,et pernicies parata costis illius.
JOB|18|13|Devorat partes cutis eius,consumat membra illius primogenitus mortis.
JOB|18|14|Avellitur de tabernaculo suo fiducia eius,et urges eum ad regem formidinum.
JOB|18|15|Habitas in tabernaculo, quod iam non est ei;aspergitur in habitatione eius sulphur.
JOB|18|16|Deorsum radices eius siccantur,sursum autem atteruntur rami eius.
JOB|18|17|Memoria illius periit de terra,et non celebrabitur nomen eius in plateis.
JOB|18|18|Expellent eum de luce in tenebraset de orbe transferent eum.
JOB|18|19|Non erit semen eius neque progenies in populo suo,nec ullae reliquiae in commoratione eius.
JOB|18|20|In die eius stupebunt novissimi,et primos invadet horror.
JOB|18|21|Haec sunt ergo tabernacula iniqui;et iste locus eius, qui ignorat Deum ".
JOB|19|1|Respondens autem Iob dixit:
JOB|19|2|" Usquequo affligitis ani mam meamet atteritis me sermonibus?
JOB|19|3|En decies obiurgatis meet non erubescitis opprimentes me.
JOB|19|4|Nempe, etsi erravi,mecum erit error meus.
JOB|19|5|Si vos contra me erigiminiet arguitis me opprobriis meis,
JOB|19|6|saltem nunc intellegite quia Deus non aequo iudicio afflixerit meet rete suo me cinxerit.
JOB|19|7|Etsi clamo: Vim patior!, non exaudior;si vociferor, non est qui iudicet.
JOB|19|8|Semitam meam circumsaepsit, et transire non possum;et in calle meo tenebras posuit.
JOB|19|9|Spoliavit me gloria meaet abstulit coronam de capite meo.
JOB|19|10|Destruxit me undique, et pereo,et evellit quasi arborem spem meam.
JOB|19|11|Iratus est contra me furor eius,et sic me habuit quasi hostem suum.
JOB|19|12|Simul venerunt turmae eiuset fecerunt sibi viam adversus meet obsederunt in gyro tabernaculum meum.
JOB|19|13|Fratres meos longe fecit a me,et noti mei quasi alieni recesserunt a me.
JOB|19|14|Dereliquerunt me propinqui mei,et, qui me noverant, obliti sunt mei.
JOB|19|15|Inquilini domus meae et ancillae meae sicut alienum habuerunt me,et quasi peregrinus fui in oculis eorum.
JOB|19|16|Servum meum vocavi, et non respondit;ore proprio deprecabar illum.
JOB|19|17|Halitum meum exhorruit uxor mea,et fetui filiis uteri mei.
JOB|19|18|Vel infantes despiciebant meet, cum surgerem, detrahebant mihi.
JOB|19|19|Abominati sunt me quondam consiliarii mei;et, quem maxime diligebam, aversatus est me.
JOB|19|20|Pelli meae, consumptis carnibus, adhaesit os meum,et evanuit cutis mea circa dentes meos.
JOB|19|21|Miseremini mei, miseremini mei, saltem vos, amici mei,quia manus Domini tetigit me.
JOB|19|22|Quare persequimini me sicut Deuset carnibus meis non saturamini?
JOB|19|23|Quis mihi tribuat, ut scribantur sermones mei?Quis mihi det, ut exarentur in libro
JOB|19|24|stilo ferreo et plumbeo,in aeternum sculpantur in silice?
JOB|19|25|Scio enim quod redemptor meus vivitet in novissimo super pulvere stabit;
JOB|19|26|et post pellem meam hanc, quam abstraxerunt,et de carne mea videbo Deum.
JOB|19|27|Quem visurus sum ego ipse,et oculi mei conspecturi sunt, et non alienum.Consumpti sunt renes mei in sinu meo.
JOB|19|28|Si ergo nunc dicitis: "Quomodo persequemur eumet radicem verbi inveniemus contra eum?",
JOB|19|29|timete a facie gladii,quoniam ultor iniquitatum gladius est;et scitote esse iudicium ".
JOB|20|1|Respondens autem Sophar Naamathites dixit:
JOB|20|2|" Idcirco cogitationes meae reducunt me,eo quod intellectus effulsit in me.
JOB|20|3|Doctrinam, qua me arguis, audiam,at spiritus intellegentiae meae respondebit mihi.
JOB|20|4|Scisne hoc a principio,ex quo positus est homo super terram,
JOB|20|5|quod exsultatio iniquorum brevis sit,et gaudium impiorum ad instar puncti?
JOB|20|6|si ascenderit usque ad caelum superbia eius,et caput eius nubes tetigerit,
JOB|20|7|quasi sterquilinium in finem perdetur,et, qui eum viderant, dicent: "Ubi est?".
JOB|20|8|Velut somnium avolans non invenietur,transiet sicut visio nocturna.
JOB|20|9|Oculus, qui eum viderat, non videbit,neque ultra intuebitur eum locus suus.
JOB|20|10|Filii eius satagent complacere pauperibus,et manus illius reddent ei possessionem suam.
JOB|20|11|Ossa eius, quae implebantur adulescentia,cum eo in pulvere dormient.
JOB|20|12|Cum enim dulce fuerit in ore eius malum,abscondet illud sub lingua sua.
JOB|20|13|Parcet illi et non derelinquet illudet celabit in gutture suo.
JOB|20|14|Panis eius in visceribus illiusvertetur in fel aspidum intrinsecus.
JOB|20|15|Divitias, quas devoravit, evomet,et de ventre illius extrahet eas Deus.
JOB|20|16|Venenum aspidum sugebat,et occidet eum lingua viperae.
JOB|20|17|Non videat rivulos olei,torrentes mellis et butyri.
JOB|20|18|Restituet quaestum suum nec deglutiet,de opibus venditionum non laetabitur.
JOB|20|19|Quoniam confringens deseruit pauperes,domum rapuit et non aedificavit eam.
JOB|20|20|Nec est satiatus venter eius;et cum desideriis suis evadere non potuit.
JOB|20|21|Non fuerunt reliquiae de cibo eius,et propterea nihil permanebit de bonis eius.
JOB|20|22|Cum satiatus fuerit, arctabitur;et omnis dolor irruet super eum.
JOB|20|23|Impleat ventrem suum:emittet Deus in eum iram furoris suiet pluet super illum bellum suum.
JOB|20|24|Fugiet arma ferreaet irruet in arcum aereum.
JOB|20|25|Sagitta transverberabit corpus eius,et fulgur iecur eius;vadent et venient super eum horribilia.
JOB|20|26|Omnes tenebrae absconditae sunt in occultis eius,devorabit eum ignis, qui non succenditur;affligetur relictus in tabernaculo suo.
JOB|20|27|Revelabunt caeli iniquitatem eius,et terra consurget adversus eum.
JOB|20|28|Auferetur germen domus illius,detrahetur in die furoris Dei.
JOB|20|29|Haec est pars hominis impii a Deo,et hereditas verborum eius a Domino ".
JOB|21|1|Respondens autem Iob dixit:
JOB|21|2|" Audite, quaeso, sermonesmeos,et sint haec consolationes vestrae.
JOB|21|3|Sustinete me, et ego loquar;et post verba mea ridebitis.
JOB|21|4|Numquid contra hominem disputatio mea est,ut merito non debeam impatiens fieri?
JOB|21|5|Attendite me et obstupesciteet superponite digitum ori vestro.
JOB|21|6|Et ego, quando recordatus fuero, pertimesco,et concutit carnem meam tremor.
JOB|21|7|Quare ergo impii vivunt,senuerunt confortatique sunt divitiis?
JOB|21|8|Semen eorum permanet coram eis,et progenies eorum in conspectu eorum.
JOB|21|9|Domus eorum securae sunt et pacatae,et non est virga Dei super illos.
JOB|21|10|Bos eorum concepit et non abortivit,vacca peperit et non est privata fetu suo.
JOB|21|11|Egrediuntur quasi greges parvuli eorum,et infantes eorum exsultant lusibus.
JOB|21|12|Tenent tympanum et citharamet gaudent ad sonitum organi.
JOB|21|13|Ducunt in bonis dies suoset in puncto ad inferna descendunt.
JOB|21|14|Qui dixerant Deo: "Recede a nobis!Scientiam viarum tuarum nolumus.
JOB|21|15|Quis est Omnipotens, ut serviamus ei,et quid nobis prodest, si oraverimus illum?".
JOB|21|16|Sint in manu eorum bona sua;consilium vero impiorum longe sit a me.
JOB|21|17|Quam saepe lucerna impiorum exstinguitur,et superveniet eis pernicies,et dolores dividet in furore suo?
JOB|21|18|Erunt sicut paleae ante faciem venti,et sicut favilla, quam turbo dispergit.
JOB|21|19|"Servabitne Deus filiis iniquitatem eius?".Retribuat illi, ut sciat.
JOB|21|20|Videbunt oculi eius interfectionem suam,et de furore Omnipotentis bibet.
JOB|21|21|Quid enim ad eum pertinet de domo sua post se,et si numerus mensium eius recidetur?
JOB|21|22|Numquid Deum docebit quispiam scientiam,qui excelsos iudicat?
JOB|21|23|Iste moritur robustus et sanus,dives et felix;
JOB|21|24|viscera eius plena sunt adipe,et medullis ossa illius irrigantur.
JOB|21|25|Alius vero moritur in amaritudine animaeabsque ullis opibus;
JOB|21|26|et tamen simul in pulvere dormient,et vermes operient eos.
JOB|21|27|Certe novi cogitationes vestraset sententias contra me iniquas.
JOB|21|28|Dicitis enim: "Ubi est domus principis,et ubi tabernacula impiorum?".
JOB|21|29|Nonne interrogastis quemlibet de viatoribuset signa eorum non agnovistis?
JOB|21|30|Quia in diem perditionis servatur maluset ad diem furoris abducetur.
JOB|21|31|Quis arguet coram eo viam eius,et, quae fecit, quis reddet illi?
JOB|21|32|Ipse ad sepulcra ducetur,et super tumulum vigilabunt.
JOB|21|33|Dulces erunt ei glebae vallis,et post se omnem hominem trahetet ante se innumerabiles.
JOB|21|34|Quomodo igitur consolamini me frustra,et responsionis vestrae restat perfidia? ".
JOB|22|1|Respondens autem Eliphaz Themanites dixit:
JOB|22|2|" Numquid Deo prodesse potest homo,cum vix intellegens sibi ipse proderit?
JOB|22|3|Quid prodest Omnipotenti, si iustus fueris,aut quid ei confers, si immaculatam feceris viam tuam?
JOB|22|4|Numquid pro tua pietate arguet teet veniet tecum in iudicium?
JOB|22|5|Et non propter malitiam tuam plurimamet infinitas iniquitates tuas?
JOB|22|6|Sumpsisti enim pignori fratres tuos sine causaet nudos spoliasti vestibus.
JOB|22|7|Aquam lasso non dedistiet esurienti cohibuisti panem.
JOB|22|8|Numquid viro forti brachio erit terra,et acceptus sedebit in ea?
JOB|22|9|Viduas dimisisti vacuaset lacertos pupillorum comminuisti.
JOB|22|10|Propterea circumdatus es laqueis,et conturbat te subita formido.
JOB|22|11|Vel tenebras non vides,et impetus aquarum opprimit te.
JOB|22|12|"Nonne Deus excelsior caelo?Et inspice stellarum verticem: quam sublimis!".
JOB|22|13|Et dicis: "Quid enim novit Deuset quasi per caliginem iudicat?
JOB|22|14|Nubes latibulum eius, nec nostra considerat;et circa orbem caeli perambulat".
JOB|22|15|Numquid semitam saeculorum custodire cupis,quam calcaverunt viri iniqui?
JOB|22|16|Qui sublati ante tempus suum,et fluvius subvertit fundamentum eorum.
JOB|22|17|Qui dicebant Deo: "Recede a nobis!"et "Quid faciet Omnipotens nobis?".
JOB|22|18|Cum ille implesset domos eorum bonis,quorum sententia procul erat ab eo.
JOB|22|19|Videbunt iusti et laetabuntur,et innocens subsannabit eos:
JOB|22|20|"Vere succisus est status eorum,et reliquias eorum devoravit ignis".
JOB|22|21|Acquiesce igitur ei, et habeto pacem;et per haec habebis fructus optimos.
JOB|22|22|Suscipe ex ore illius legemet pone sermones eius in corde tuo.
JOB|22|23|Si reversus fueris ad Omnipotentem, aedificaberiset longe facies iniquitatem a tabernaculo tuo.
JOB|22|24|Comparabis tamquam terram aurumet tamquam glaream torrentis Ophir.
JOB|22|25|Eritque Omnipotens metallum tuum,et argentum coacervabitur tibi.
JOB|22|26|Tunc super Omnipotentem deliciis afflueset elevabis ad Deum faciem tuam.
JOB|22|27|Supplex rogabis eum, et exaudiet te,et vota tua reddes.
JOB|22|28|Decernes rem, et veniet tibi,et in viis tuis splendebit lumen.
JOB|22|29|Quia humiliat eum, qui loquitur superba,et demissus oculis ipse salvabitur.
JOB|22|30|Eripiet innocentem,eripietur autem in munditia manuum suarum ".
JOB|23|1|Respondens autem Iob ait:
JOB|23|2|" Nunc quoque in amaritu tudine est querela mea,et manus eius aggravata est super gemitum meum.
JOB|23|3|Quis mihi tribuat, ut cognoscam et inveniam illumet veniam usque ad solium eius?
JOB|23|4|Ponam coram eo iudiciumet os meum replebo increpationibus,
JOB|23|5|ut sciam verba, quae mihi respondeat,et intellegam quid loquatur mihi.
JOB|23|6|Num multa fortitudine contendet mecum?Non! Ipse tantum audiat!
JOB|23|7|Tunc iustus disceptabit cum illo,et ego evaderem in perpetuo a iudice meo.
JOB|23|8|Si ad orientem iero, non apparet;si ad occidentem, non intellegam eum.
JOB|23|9|Si ad sinistram pergam, non apprehendam eum;si me vertam ad dexteram, non videbo illum.
JOB|23|10|Ipse vero scit viam meam,et, si probaverit me, quasi aurum egrediar.
JOB|23|11|Vestigia eius secutus est pes meus,viam eius custodivi et non declinavi ex ea.
JOB|23|12|A mandatis labiorum eius non recessiet in sinu meo abscondi verba oris eius.
JOB|23|13|Ipse enim solus est, et quis repellet eum?Et anima eius, quodcumque voluit, hoc fecit.
JOB|23|14|Cum expleverit in me voluntatem suam,et alia multa similia praesto sunt ei;
JOB|23|15|et idcirco a facie eius turbatus sumet considerans eum timore sollicitor.
JOB|23|16|Deus mollivit cor meum,et Omnipotens conturbavit me.
JOB|23|17|Non enim perii propter imminentes tenebras,nec faciem meam operuit caligo.
JOB|24|1|Cur ab Omnipotente non sunt abscondita tempora,qui autem noverunt eum, ignorant dies illius?
JOB|24|2|Alii terminos transtulerunt,diripuerunt greges et paverunt eos.
JOB|24|3|Asinum pupillorum abegeruntet abstulerunt pro pignore bovem viduae.
JOB|24|4|Subverterunt pauperum viam,et simul se occultare coacti sunt mansueti terrae.
JOB|24|5|Alii, quasi onagri in deserto,egrediuntur ad opus suum:vigilantes ad praedamin terra arida ad panem liberis.
JOB|24|6|Agrum non suum demetuntet vineam peccatoris vindemiant.
JOB|24|7|Nudi pernoctant sine indumento,nec est eis operimentum in frigore.
JOB|24|8|Imbre montium riganturet non habentes refugium adhaerent rupibus.
JOB|24|9|Abripuerunt pupillum ab ubereet pauperem pignori sumpserunt;
JOB|24|10|nudi et incedentes absque vestituet esurientes portant spicas.
JOB|24|11|Inter muros oleum expresseruntet calcatis torcularibus sitiunt.
JOB|24|12|De civitatibus morientes ingemuerunt,et anima vulneratorum clamavit,et Deus non ponit aurem ad precem.
JOB|24|13|Ipsi fuerunt rebelles lumini,nescierunt vias eiusnec morati sunt in semitis eius.
JOB|24|14|Mane primo consurgit homicida,interficit egenum et pauperem;per noctem vero erit quasi fur.
JOB|24|15|Oculus adulteri observat caliginemdicens: "Non me videbit oculus";et operiet vultum suum.
JOB|24|16|Perfodit in tenebris domos, interdiu sese abdideruntet ignoraverunt lucem.
JOB|24|17|Si subito apparuerit aurora, arbitrantur umbram mortis,nam sunt assueti terroribus umbrae mortis.
JOB|24|18|"Levis est super faciem aquae;maledicta est pars eius in terra,nec est qui se dirigat ad vineas eius.
JOB|24|19|Siccitas et calor abstulerunt aquas nivium,et inferi eos, qui peccaverunt.
JOB|24|20|Sinus matris obliviscatur eius,dulcedo illius vermes fiant;non sit in recordatione,sed conteratur quasi lignum iniquitas.
JOB|24|21|Male egit cum sterili, quae non parit,et viduae bene non fecit.
JOB|24|22|Detraxit fortes in fortitudine suaet, cum steterit, ille non credet vitae suae.
JOB|24|23|Dedit ei locum securitatis, quo sustentetur;oculi autem eius sunt in viis illius.
JOB|24|24|Elevati sunt ad modicum et non subsistent,et humiliabuntur sicut omnia et auferenturet sicut summitates spicarum conterentur".
JOB|24|25|Quod si non est ita, quis me potest arguere esse mentitumet ponere in nihilum verba mea? ".
JOB|25|1|Respondens autem Baldad Suhites dixit:
JOB|25|2|" Potestas et terror apud eum est,qui facit pacem in sublimibus suis.
JOB|25|3|Numquid est numerus militum eius?Et super quem non surget lumen illius?
JOB|25|4|Numquid iustificari potest homo comparatus Deo,aut apparere mundus natus de muliere?
JOB|25|5|Ecce luna etiam non splendet,et stellae non sunt mundae in conspectu eius;
JOB|25|6|quanto magis homo putredo,et filius hominis vermis ".
JOB|26|1|Respondens autem Iob dixit:
JOB|26|2|" Quomodo adiuvisti imbecillem?Et sustentas brachium eius, qui non est fortis?
JOB|26|3|Quod dedisti illi consilium, qui non habet sapientiam?Et prudentiam tuam ostendisti plurimam!
JOB|26|4|Quem docere voluisti?Et cuius est spiritus, qui egreditur ex te?
JOB|26|5|Ecce umbrae gemunt sub aquis,et qui habitant cum eis.
JOB|26|6|Nudus est infernus coram illo,et nullum est operimentum Perditioni.
JOB|26|7|Qui extendit aquilonem super vacuumet appendit terram super nihilum.
JOB|26|8|Qui ligat aquas in nubibus suis,ut non erumpant pariter deorsum.
JOB|26|9|Qui operit faciem solii suiexpandens super illud nebulam suam.
JOB|26|10|Terminum circumdedit aquis,usque dum finiantur lux et tenebrae.
JOB|26|11|Columnae caeli contremiscuntet pavent ab increpatione eius.
JOB|26|12|In fortitudine sua terruit mareet prudentia sua percussit Rahab.
JOB|26|13|Spiritus eius serenavit caelos,et manus eius confodit colubrum fugientem.
JOB|26|14|Ecce haec sunt termini viarum eius;et, cum vix parvam stillam sermonis eius audierimus,quis poterit tonitruum magnitudinis illius intueri? ".
JOB|27|1|Addidit quoque Iob assu mens parabolam suam et dixit:
JOB|27|2|" Vivit Deus, qui abstulit ius meum, et Omnipotens, qui ad amaritudinem adduxit animam meam,
JOB|27|3|quia, donec superest halitus in me,et spiritus Dei in naribus meis,
JOB|27|4|non loquentur labia mea iniquitatem,nec lingua mea meditabitur mendacium!
JOB|27|5|Absit a me, ut iustos vos esse iudicem;donec exspirem, non recedam ab innocentia mea.
JOB|27|6|Iustificationem meam, quam coepi tenere, non deseram,neque enim reprehendit me cor meum in omni vita mea.
JOB|27|7|Sit ut impius inimicus meus,et adversarius meus quasi iniquus.
JOB|27|8|Quae est enim spes impii, cum secet,cum rapiat Deus animam eius?
JOB|27|9|Numquid Deus audiet clamorem eius,cum venerit super eum angustia?
JOB|27|10|Aut poterit in Omnipotente delectariet invocare Deum omni tempore?
JOB|27|11|Docebo vos manum Dei,quae Omnipotens habeat, nec abscondam.
JOB|27|12|Ecce vos omnes observastis,et quid sine causa vana loquimini?
JOB|27|13|Haec est pars hominis impii apud Deum,et hereditas violentorum, quam ab Omnipotente suscipient.
JOB|27|14|Si multiplicati fuerint filii eius, in gladio erunt,et nepotes eius non saturabuntur pane.
JOB|27|15|Qui reliqui fuerint ex eo, sepelientur in interitu,et viduae illius non plorabunt.
JOB|27|16|Si comportaverit quasi terram argentumet sicut lutum praeparaverit vestimenta,
JOB|27|17|praeparabit quidem, sed iustus vestietur illis,et argentum innocens dividet.
JOB|27|18|Aedificavit sicut aranea domum suam,et sicut custos fecit umbraculum.
JOB|27|19|Dives, cum dormierit, nihil secum auferet;aperiet oculos suos et nihil inveniet.
JOB|27|20|Apprehendet eum quasi aqua inopia,nocte opprimet eum tempestas.
JOB|27|21|Tollet eum ventus urens et auferet,et velut turbo rapiet eum de loco suo.
JOB|27|22|Et mittet super eum et non parcet;de manu eius fugiens fugiet.
JOB|27|23|Complodet super eum manus suaset sibilabit eum de loco suo.
JOB|28|1|Habet argentum venarum principiaet auro locus est, in quo conflatur.
JOB|28|2|Ferrum de terra tollitur,et lapis solutus calore in aes vertitur.
JOB|28|3|Terminum posuit tenebriset universorum finem ipse scrutatur,lapidem quoque caliginis et umbrae.
JOB|28|4|Aperuit cuniculos gens peregrina,ipsique obliti sunt pedes,penduli haerent plus quam vir nutans.
JOB|28|5|Terra, de qua oriebatur panis,in profundo subversa est sicut per ignem.
JOB|28|6|Locus sapphiri lapides eius,et glebae illius aurum.
JOB|28|7|Semitam ignoravit avis rapax,nec intuitus est eam oculus vulturis.
JOB|28|8|Non calcaverunt eam filii superbiae,nec pertransivit per eam leaena.
JOB|28|9|Ad silicem extendit manum suam,subvertit a radicibus montes.
JOB|28|10|In petris canales excidit,et omne pretiosum vidit oculus eius.
JOB|28|11|Profunda quoque fluviorum scrutatus estet abscondita in lucem produxit.
JOB|28|12|Sapientia vero ubi invenitur?Et quis est locus intellegentiae?
JOB|28|13|Nescit homo structuram eius,nec invenitur in terra viventium.
JOB|28|14|Abyssus dicit: "Non est in me";et mare loquitur: "Non est mecum".
JOB|28|15|Non dabitur aurum obryzum pro ea,nec appendetur argentum in commutatione eius.
JOB|28|16|Non appendetur auro Ophirnec lapidi sardonycho pretiosissimo vel sapphiro.
JOB|28|17|Non adaequabitur ei aurum vel vitrum,nec commutabuntur pro ea vasa auri.
JOB|28|18|Corallia et crystallum non memorabuntur comparatione eius;et possessio sapientiae potior margaritis.
JOB|28|19|Non adaequabitur ei topazius de Aethiopianec auro mundissimo componetur.
JOB|28|20|Unde ergo sapientia venit,et quis est locus intellegentiae?
JOB|28|21|Abscondita est ab oculis omnium viventium,volucres quoque caeli latet.
JOB|28|22|Perditio et mors dixerunt:Auribus nostris audivimus famam eius".
JOB|28|23|Deus intellegit viam eius,et ipse novit locum illius.
JOB|28|24|Ipse enim fines mundi intueturet omnia, quae sub caelo sunt, respicit.
JOB|28|25|Qui fecit ventis ponduset aquas appendit in mensura,
JOB|28|26|quando ponebat pluviis legemet viam procellis sonantibus,
JOB|28|27|tunc vidit illam et enarravitet praeparavit et investigavit.
JOB|28|28|Et dixit homini: "Ecce timor Domini, ipsa est sapientia;et recedere a malo intellegentia" ".
JOB|29|1|Addidit quoque Iob assumens parabolam suam et di xit:
JOB|29|2|" Quis mihi tribuat, ut sim iuxta menses pristinos,secundum dies, quibus Deus custodiebat me?
JOB|29|3|Quando splendebat lucerna eius super caput meum,et ad lumen eius ambulabam in tenebris.
JOB|29|4|Sicut fui in diebus adulescentiae meae,quando familiaris Deus erat in tabernaculo meo,
JOB|29|5|quando erat Omnipotens mecum,et in circuitu meo pueri mei,
JOB|29|6|quando lavabam pedes meos lacte,et petra fundebat mihi rivos olei.
JOB|29|7|Quando procedebam ad portam civitatiset in platea parabam cathedram mihi,
JOB|29|8|videbant me iuvenes et abscondebantur,et senes assurgentes stabant.
JOB|29|9|Principes cessabant loquiet digitum superponebant ori suo.
JOB|29|10|Vocem suam cohibebant duces,et lingua eorum palato suo adhaerebat.
JOB|29|11|Auris audiens beatificabat me,et oculus videns testimonium reddebat mihi,
JOB|29|12|eo quod liberassem pauperem vociferantemet pupillum, cui non esset adiutor.
JOB|29|13|Benedictio perituri super me veniebat,et cor viduae iubilare feci.
JOB|29|14|Iustitia indutus sum et vestivi me,sicut vestimento et diademate, iudicio meo.
JOB|29|15|Oculus fui caecoet pes claudo;
JOB|29|16|pater eram pauperumet causam viri ignoti diligentissime investigabam.
JOB|29|17|Conterebam molas iniquiet de dentibus illius auferebam praedam.
JOB|29|18|Dicebamque: In nidulo meo moriaret sicut palma multiplicabo dies.
JOB|29|19|Radix mea aperta est secus aquas,et ros morabitur in ramis meis.
JOB|29|20|Gloria mea semper innovabitur,et arcus meus in manu mea instaurabitur.
JOB|29|21|Qui me audiebant, blandiebanturet intenti tacebant ad consilium meum.
JOB|29|22|Verbis meis addere nihil audebant,et super illos stillabat eloquium meum.
JOB|29|23|Exspectabant me sicut pluviamet os suum aperiebant quasi ad imbrem serotinum.
JOB|29|24|Si quando ridebam ad eos, non credebant,et lux vultus mei non cadebat in terram.
JOB|29|25|Si voluissem ire ad eos, sedebam primus;cumque sederem quasi rex, circumstante exercitu,eram tamen maerentium consolator.
JOB|30|1|Nunc autem derident meiuniores tempore,quorum non dignabar patresponere cum canibus gregis mei;
JOB|30|2|quorum virtus manuum mihi erat pro nihilo,et robur iuvenile perierat totum.
JOB|30|3|Egestate et fame steriles, qui rodebant in solitudine,serotino tempore fiebant turbo et vastatio;
JOB|30|4|et mandebant herbas et arborum frutices,et radix iuniperorum erat cibus eorum.
JOB|30|5|De medio eiciebantur,clamabant contra eos tamquam fures;
JOB|30|6|ad ripas habitabant torrentiumet in cavernis terrae et petrarum;
JOB|30|7|inter frutices rudebant,sub sentibus se congerebant;
JOB|30|8|filii stultorum et ignobiliumet de terra penitus exturbati.
JOB|30|9|Nunc in eorum canticum versus sumet factus sum eis in proverbium.
JOB|30|10|Abominantur me et longe fugiunt a meet faciem meam conspuere non verentur.
JOB|30|11|Pharetram enim suam aperuit et afflixit meet frenum in os meum immisit.
JOB|30|12|Ad dexteram progenies surrexerunt;pedes meos subverteruntet complanaverunt contra me semitas ruinae.
JOB|30|13|Dissipaverunt itinera mea,insidiati sunt mihi et praevaluerunt,et non fuit qui ferret auxilium.
JOB|30|14|Quasi rupto muro et aperto irruerunt super meet sub ruinis devoluti sunt.
JOB|30|15|Versi sunt contra me in terrores,persequitur quasi ventus principatum meum,et velut nubes pertransiit salus mea.
JOB|30|16|Nunc autem in memetipso effunditur anima mea;et possident me dies afflictionis.
JOB|30|17|Nocte os meum perforatur doloribus;et, qui me comedunt, non dormiunt.
JOB|30|18|In multitudine roboris tenent vestimentum meumet quasi capitio tunicae succinxerunt me.
JOB|30|19|Proiecit me in lutum,et assimilatus sum favillae et cineri.
JOB|30|20|Clamo ad te, et non exaudis me;sto, et non respicis me.
JOB|30|21|Mutatus es mihi in crudelemet in duritia manus tuae adversaris mihi.
JOB|30|22|Elevasti meet quasi super ventum ponens dissolvisti me.
JOB|30|23|Scio quia morti trades me,ubi constituta est domus omni viventi.
JOB|30|24|Verumtamen non ad ruinam mittit manum;et in exitio eius erit salvatio.
JOB|30|25|An non flebam quondam super eo, qui afflictus erat,et compatiebatur anima mea pauperi?
JOB|30|26|Exspectabam bona, et venerunt mihi mala;praestolabar lucem, et eruperunt tenebrae.
JOB|30|27|Interiora mea efferbuerunt absque ulla requie;praevenerunt me dies afflictionis.
JOB|30|28|Taetro vultu incedebam sine consolatione,consurgens in turba clamabam.
JOB|30|29|Frater fui draconumet socius struthionum.
JOB|30|30|Cutis mea denigrata est super me,et ossa mea aruerunt prae caumate.
JOB|30|31|Versa est in luctum cithara mea,et organum meum in vocem flentium.
JOB|31|1|Pepigi foedus cum oculis meisut ne cogitarem quidem de virgine.
JOB|31|2|Quae enim pars mea apud Deum desuper,et quae hereditas apud Omnipotentem in excelsis?
JOB|31|3|Numquid non perditio est iniquo,et alienatio operantibus iniustitiam?
JOB|31|4|Nonne ipse considerat vias measet cunctos gressus meos dinumerat?
JOB|31|5|Si ambulavi in vanitate,et festinavit in dolo pes meus,
JOB|31|6|appendat me in statera iustaet sciat Deus integritatem meam.
JOB|31|7|Si declinavit gressus meus de via,et si secutum est oculos meos cor meum,et si manibus meis adhaesit macula,
JOB|31|8|seram, et alius comedat,et progenies mea eradicetur.
JOB|31|9|Si deceptum est cor meum super muliere,et si ad ostium amici mei insidiatus sum,
JOB|31|10|molat pro alio uxor mea,et super illam incurventur alii.
JOB|31|11|Hoc enim nefas estet iniquitas iudicialis;
JOB|31|12|ignis est usque ad perditionem devoranset omnia eradicans genimina.
JOB|31|13|Si contempsi subire iudicium cum servo meo et ancilla mea,cum disceptarent adversum me,
JOB|31|14|quid enim faciam, cum surrexerit ad iudicandum Deus;et, cum quaesierit, quid respondebo illi?
JOB|31|15|Numquid non in ventre fecit me,qui et illum operatus est,et formavit me in visceribus unus?
JOB|31|16|Si negavi, quod volebant, pauperibuset oculos viduae languescere feci;
JOB|31|17|si comedi buccellam meam solus,et non comedit pupillus ex ea,
JOB|31|18|quia ab infantia mea educavi eum ut pateret de ventre matris meae direxi eam;
JOB|31|19|si despexi pereuntem, eo quod non habuerit indumentum,et absque operimento pauperem;
JOB|31|20|si non benedixerunt mihi latera eius,et de velleribus ovium mearum calefactus est;
JOB|31|21|si levavi super pupillum manum meam,cum viderem in porta adiutorium mihi,
JOB|31|22|umerus meus a iunctura sua cadat,et brachium meum cum ossibus lacertorum confringatur,
JOB|31|23|quia timor super me calamitas a Deo,et contra maiestatem eius nihil valerem!
JOB|31|24|Si putavi aurum securitatem meamet obryzo dixi: Fiducia mea!;
JOB|31|25|si laetatus sum super multis divitiis meis,et quia plurima repperit manus mea;
JOB|31|26|si vidi solem, cum fulgeret,et lunam incedentem clare,
JOB|31|27|et decepit me in abscondito cor meum,et osculatus sum manum meam ore meo,
JOB|31|28|quae est iniquitas iudicialis,eo quod negassem Deum desuper;
JOB|31|29|si gavisus sum ad ruinam eius, qui me oderat,et exsultavi quod invenisset eum malum,
JOB|31|30|cum non dederim ad peccandum guttur meum,ut expeterem maledicens animam eius;
JOB|31|31|si non dixerunt viri tabernaculi mei: "Quis det, qui de carnibus eius non saturatus sit?";
JOB|31|32|foris non mansit peregrinus,ostium meum viatori patuit;
JOB|31|33|si abscondi quasi homo peccatum meumet celavi in sinu meo iniquitatem meam;
JOB|31|34|si expavi ad multitudinem nimiam,et despectio propinquorum terruit me,et magis tacui nec egressus sum ostium.
JOB|31|35|Quis mihi tribuat auditorem?Ecce signum meum! Omnipotens respondeat mihi!Ecce liber, quem scripsit vir litis meae,
JOB|31|36|ut in umero meo portem illumet alligem illum quasi coronam mihi.
JOB|31|37|Numerum graduum meorum pronuntiabo illiet quasi principem adibo eum.
JOB|31|38|Si adversum me terra mea clamat,et cum ipsa sulci eius deflent;
JOB|31|39|si fructus eius comedi absque pecuniaet animam agricolarum eius afflixi,
JOB|31|40|pro frumento oriatur mihi tribulus,et pro hordeo herba foetida! ".Finita sunt verba Iob.
JOB|32|1|Omiserunt autem tres viri isti respondere Iob, eo quod iustus sibi videretur.
JOB|32|2|Et iratus indignatusque est Eliu filius Barachel Buzites de cognatione Ram; iratus est autem adversum Iob, eo quod iustum se esse diceret coram Deo.
JOB|32|3|Porro adversum amicos eius indignatus est, eo quod non invenissent responsionem, sed tantummodo condemnassent Iob.
JOB|32|4|Igitur Eliu exspectavit Iob loquentem, eo quod seniores essent, qui loquebantur;
JOB|32|5|cum autem vidisset Eliu quod tres respondere non potuissent, iratus est vehementer.
JOB|32|6|Respondensque Eliu filius Barachel Buzites dixit: Iunior sum tempore,vos autem antiquiores;idcirco veritus sum et timuivobis indicare meam sententiam.
JOB|32|7|Dixi: Aetas loquetur,et annorum multitudo docebit sapientiam.
JOB|32|8|Sed, ut video, spiritus est in hominibus,et inspiratio Omnipotentis dat intellegentiam.
JOB|32|9|Non sunt longaevi sapientes,nec senes intellegunt iudicium.
JOB|32|10|Ideo dicam: Audite me,ostendam vobis etiam ego meam sapientiam.
JOB|32|11|Exspectavi enim sermones vestros,intendi aurem in prudentiam vestram, donec investigaretis,
JOB|32|12|et ut vos intellegerem nitebar.Sed, ut video, non est qui possit arguere Iobet respondere ex vobis sermonibus eius.
JOB|32|13|Ne forte dicatis: "Invenimus sapientiam;Deus proiecit eum, non homo".
JOB|32|14|Non parabo mihi verba,et ego non secundum sermones vestros respondebo illi.
JOB|32|15|Extimuerunt nec responderunt ultra;abstuleruntque a se eloquia.
JOB|32|16|Quoniam igitur exspectavi, et non sunt locuti,steterunt, nec ultra responderunt,
JOB|32|17|respondebo et ego partem meamet ostendam scientiam meam.
JOB|32|18|Plenus sum enim sermonibus,et coarctat me spiritus pectoris mei;
JOB|32|19|en venter meus quasi mustum absque spiraculo,quod lagunculas novas disrumpit.
JOB|32|20|Loquar et respirabo paululum,aperiam labia mea et respondebo.
JOB|32|21|Non accipiam personam viriet nulli homini blandiar.
JOB|32|22|Nescio enim blandiri,quia in brevi tolleret me Factor meus.
JOB|33|1|Audi igitur, Iob, eloquia meaet omnes sermones meos ausculta.
JOB|33|2|Ecce aperui os meum,loquatur lingua mea in faucibus meis.
JOB|33|3|Ex recto corde sermones mei sunt,et sententiam puram labia mea loquentur.
JOB|33|4|Spiritus Dei fecit me,et spiraculum Omnipotentis vivificavit me.
JOB|33|5|Si potes, responde mihi,praepara te coram me et consiste.
JOB|33|6|Ecce ego sicut tu coram Deo sumet de eodem luto abscissus sum et ego.
JOB|33|7|Verumtamen terror meus non te terreat,et onus meum non sit tibi grave.
JOB|33|8|Dixisti ergo in auribus meis,et vocem verborum tuorum audivi:
JOB|33|9|"Mundus sum ego et absque delicto;immaculatus, et non est iniquitas in me.
JOB|33|10|Quia querelas in me repperit,ideo arbitratus est me inimicum sibi;
JOB|33|11|posuit in nervo pedes meos,custodivit omnes semitas meas".
JOB|33|12|Hoc est ergo, in quo non es iustificatus, respondebo tibi,quia maior est Deus homine.
JOB|33|13|Quare adversus eum contendis,quod non ad omnia verba responderit tibi?
JOB|33|14|Semel loquitur Deus,et secundo idipsum non repetit.
JOB|33|15|Per somnium in visione nocturna,quando irruit sopor super homines,et dormiunt in lectulo,
JOB|33|16|tunc aperit aures virorumet in visionibus terret eos,
JOB|33|17|ut avertat hominem ab his, quae facit,et liberet eum de superbia,
JOB|33|18|eruens animam eius a foveaet vitam illius, ut non transeat canalem mortis.
JOB|33|19|Increpat quoque per dolorem in lectulo,et tremitus ossium eius continuus.
JOB|33|20|Abominabilis ei fit in vita sua panis,et animae illius cibus ante desiderabilis.
JOB|33|21|Tabescet caro eius in conspectu,et ossa, quae non videbantur, nudabuntur.
JOB|33|22|Appropinquavit corruptioni foveae,et vita illius mortiferis sedibus.
JOB|33|23|Si fuerit apud eum angelus, unus de milibus interpres,ut annuntiet homini aequitatem,
JOB|33|24|miserebitur eius et dicet:Libera eum, ut non descendat in foveam;inveni, in quo ei propitier".
JOB|33|25|Revirescet caro eius plus quam in iuventute,revertetur ad dies adulescentiae suae.
JOB|33|26|Deprecabitur Deum, et placabilis ei erit;et videbit faciem eius in iubilo,et reddet homini iustitiam suam.
JOB|33|27|Canit ad homines et dicit: "Peccavi et iustitiam pervertiet non debui satisfacere.
JOB|33|28|Liberavit animam suam, ne pergeret in foveam,sed vivens lucem videret".
JOB|33|29|Ecce haec omnia operatur Deusduobus, tribus vicibus cum homine,
JOB|33|30|ut revocet animas eorum a foveaet illuminet luce viventium.
JOB|33|31|Attende, Iob, et audi meet tace, dum ego loquor.
JOB|33|32|Si autem habes quod loquaris, responde mihi; loquere, volo enim te apparere iustum.
JOB|33|33|Quod si non habes, audi me;tace, et docebo te sapientiam ".
JOB|34|1|Pronuntians itaque Eliu etiam haec locutus est:
JOB|34|2|" Audite, sapientes, verba mea;et eruditi, auscultate me.
JOB|34|3|Auris enim verba probat,et guttur escas gustu diiudicat.
JOB|34|4|Iudicium eligamus nobiset inter nos videamus quid sit melius.
JOB|34|5|Quia dixit Iob: "Iustus sum,et Deus avertit iudicium meum;
JOB|34|6|in iudicando enim me mendacium est,violenta sagitta mea absque ullo peccato".
JOB|34|7|Quis est vir, ut est Iob,qui bibit subsannationem quasi aquam,
JOB|34|8|qui graditur una cum operantibus iniquitatemet ambulat cum viris impiis?
JOB|34|9|Dixit enim: "Non prodest viro,etiamsi cum Deo familiariter agit".
JOB|34|10|Ideo, viri cordati, audite me:Absit a Deo impietas, et ab Omnipotente iniquitas.
JOB|34|11|Opus enim hominis reddet eiet iuxta vias singulorum restituet eis.
JOB|34|12|Vere enim Deus non operatur malum,nec Omnipotens subvertet iudicium.
JOB|34|13|Quis commisit ei terram suam,aut quis posuit totum orbem?
JOB|34|14|Si direxerit ad se cor suum,spiritum illius et halitum ad se trahat,
JOB|34|15|deficiet omnis caro simul,et homo in cinerem revertetur.
JOB|34|16|Si habes ergo intellectum, audi hocet ausculta vocem eloquii mei:
JOB|34|17|Numquid, qui non amat iudicium, reget imperio?Num iustum magnum condemnabis,
JOB|34|18|qui dicet regi: "Nequam!",qui vocabit duces: "Impios!",
JOB|34|19|qui non accipit personas principumnec cognovit opulentum,cum disceptaret contra pauperem?Opus enim manuum eius sunt universi.
JOB|34|20|Subito morientur; et in media nocteturbabuntur populi et pertransibunt,et auferent violentum absque conatu.
JOB|34|21|Oculi enim eius super vias hominum,et omnes gressus eorum considerat.
JOB|34|22|Non sunt tenebrae, et non est umbra mortis,ut abscondantur ibi, qui operantur iniquitatem.
JOB|34|23|Nec enim ultra homini ponit conveniendi locum,ut veniat ad Deum in iudicium.
JOB|34|24|Conteret potentes sine inquisitioneet stare faciet alios pro eis.
JOB|34|25|Novit enim opera eorumet idcirco inducet noctem, et conterentur.
JOB|34|26|Quasi impios percussit eosin loco videntium,
JOB|34|27|qui quasi de industria recesserunt ab eoet omnes vias eius intellegere noluerunt,
JOB|34|28|cum induceret ad se clamorem egeni et audiret vocem pauperum.
JOB|34|29|Ipse enim si quieverit, quis est qui condemnet?Et si absconderit vultum, quis est qui contempletur eum,super gentem et super homines simul?
JOB|34|30|Ne regnet homo impius,ne sint laquei populo.
JOB|34|31|Si enim dixit quispiam Deo:Ferre debui! Iam non perverse agam.
JOB|34|32|Dum videam, tu doce me;si iniquitatem operatus sum, ultra non addam".
JOB|34|33|Numquid pro te Deus satisfaciet,quia respuisti?Tu enim eliges, et non ego;et si quid nosti melius, loquere.
JOB|34|34|Viri intellegentes loquentur mihi,et vir sapiens, qui audiet me:
JOB|34|35|"Iob autem non in sapientia locutus est,et verba illius non sonant disciplinam".
JOB|34|36|Utique, probetur Iob usque ad finemde responsionibus hominum iniquitatis.
JOB|34|37|Quia addit super peccata sua delictum,inter nos plaudit manibuset multiplicat sermones suos contra Deum ".
JOB|35|1|Igitur Eliu haec rursum locutus est:
JOB|35|2|" Numquid aequa tibi videtur tua cogitatio,ut diceres: "Iustificatio mea coram Deo"?
JOB|35|3|Dixisti enim: "Quid ad te?Vel quid tibi proderit, si ego peccavero?".
JOB|35|4|Itaque ego respondebo sermonibus tuiset amicis tuis tecum.
JOB|35|5|Suspice caelum et intuereet contemplare nubes quod altiores te sint.
JOB|35|6|Si peccaveris, quid facies ei?Et si multiplicatae fuerint iniquitates tuae, quid facies contra eum?
JOB|35|7|Porro si iuste egeris, quid donabis ei?Aut quid de manu tua accipiet?
JOB|35|8|Homini, qui similis tui est, nocebit impietas tua,et filium hominis adiuvabit iustitia tua.
JOB|35|9|Propter multitudinem oppressorum clamabuntet eiulabunt propter vim brachii tyrannorum,
JOB|35|10|sed nemo dixit: "Ubi est Deus, qui fecit me,qui dedit carmina in nocte,
JOB|35|11|qui docet nos super iumenta terraeet super volucres caeli erudit nos?".
JOB|35|12|Ibi clamabunt, et non exaudiet,propter superbiam malorum.
JOB|35|13|Etiam, frustra: non audiet Deus,et Omnipotens non intuebitur.
JOB|35|14|Omnino cum dixeris: "Non considerat",iudicium est coram illo, et exspectas eum.
JOB|35|15|Et nunc cum dicis: "Ira eius poenas non infert,nec ulciscitur scelus valde",
JOB|35|16|Iob frustra aperit os suumet absque scientia verba multiplicat ".
JOB|36|1|Addens quoque Eliu haec locutus est:
JOB|36|2|" Sustine me paululum, et indicabo tibi:adhuc enim habeo quod pro Deo loquar.
JOB|36|3|Repetam scientiam meam a longeet Factori meo tribuam iustitiam.
JOB|36|4|Vere enim absque mendacio sermones mei,et perfectus scientia adest tecum.
JOB|36|5|Deus potens est; non abicit,potens virtute cordis.
JOB|36|6|Non vivere faciet impium,sed iudicium pauperibus tribuit.
JOB|36|7|Non auferet a iusto oculos suoset reges in solio collocat in perpetuum,et illi eriguntur.
JOB|36|8|Et si fuerint vincti compedibuset vinciantur funibus paupertatis,
JOB|36|9|indicabit eis opera eorumet scelera eorum, quia violenti fuerunt.
JOB|36|10|Revelabit quoque aurem eorum, ut corripiat,et loquetur, ut revertantur ab iniquitate.
JOB|36|11|Si audierint et observaverint,complebunt dies suos in bonoet annos suos in deliciis.
JOB|36|12|Si autem non audierint, transibunt per canalem mortiset consumentur in stultitia.
JOB|36|13|Impii corde sibi reponent iram Deineque clamabunt, cum vincti fuerint.
JOB|36|14|Morietur in iuventute anima eorum,et vita eorum in adulescentia.
JOB|36|15|Eripiet de angustia sua pauperemet revelabit in tribulatione aurem eius.
JOB|36|16|Igitur salvabit te de ore angusto,amplitudo et non angustiae erunt sub te;requies autem mensae tuae erit plena pinguedine.
JOB|36|17|Causa tua quasi impii iudicata est,causam iudiciumque tenebunt.
JOB|36|18|Cave, ne te seducat abundantia,nec multitudo donorum inclinet te.
JOB|36|19|Nonne proferetur clamor tuus nisi in angustia?Et omnes conatus roboris?
JOB|36|20|Ne inhies nocti,ut ascendat turba pro eis.
JOB|36|21|Cave, ne declines ad iniquitatem;propter hoc enim expertus es miseriam.
JOB|36|22|Ecce, Deus excelsus in fortitudine sua.Quis ei similis doctor?
JOB|36|23|Quis poterit scrutari vias eius,aut quis potest ei dicere: "Operatus es iniquitatem"?
JOB|36|24|Memento, ut magnifices opus eius,de quo cecinerunt viri.
JOB|36|25|Omnes homines vident eum,unusquisque intuetur procul.
JOB|36|26|Ecce, Deus magnus vincens scientiam nostram;numerus annorum eius inaestimabilis.
JOB|36|27|Qui aufert stillas pluviaeet effundit imbres ad instar fluminis,
JOB|36|28|quos nubes effundunt,stillantes super homines multos.
JOB|36|29|Profecto quis intellegit dilatationem nubium,strepitum tabernaculi eius?
JOB|36|30|Ecce extendit circum se lumen suumet fundamenta maris texit.
JOB|36|31|Per haec enim iudicat populoset dat escas copiose.
JOB|36|32|In manibus abscondit lucemet praecipit ei, ut percutiat.
JOB|36|33|Fragor eius de eo annuntiat,zelans ira contra iniquitatem.
JOB|37|1|Super hoc expavit cor meumet emotum est de loco suo.
JOB|37|2|Audite fremitum vocis eiuset murmur de ore illius procedens.
JOB|37|3|Subter omnes caelos ipsum revolvit,et lumen illius super terminos terrae.
JOB|37|4|Post eum rugiet sonitus,tonabit voce magnitudinis suae;et non retardabit, cum audita fuerit vox eius.
JOB|37|5|Tonabit Deus in voce sua mirabiliter,qui facit magna et inscrutabilia.
JOB|37|6|Qui praecipit nivi, ut descendat in terram,et hiemis pluviis et imbri, ut roborentur.
JOB|37|7|Qui in manu omnium hominum signat,ut noverint singuli opera sua.
JOB|37|8|Ingredietur bestia latibulumet in antro suo morabitur.
JOB|37|9|Ab interioribus egredietur tempestas,et ab Arcturo frigus.
JOB|37|10|Flante Deo, datur gelu,et expansio aquarum solidatur.
JOB|37|11|Fulgur proicitur a nube,et nubes spargunt lumen suum;
JOB|37|12|quae lustrant per circuitum,quocumque eas voluntas gubernantis duxerit,ad omne, quod praeceperit illis super faciem orbis terrarum,
JOB|37|13|sive in castigatione terrae suae,sive in misericordia eas iusserit inveniri.
JOB|37|14|Ausculta haec, Iob;sta et considera mirabilia Dei.
JOB|37|15|Numquid scis quando praeceperit Deus,ut ostenderent lucem nubes eius?
JOB|37|16|Numquid nosti semitas nubium magnaset mirabilia perfecti scientia?
JOB|37|17|Nonne vestimenta tua calida sunt,cum quieverit terra austro?
JOB|37|18|Tu forsitan cum eo expandisti caelos,qui solidissimi, quasi aere, fusi sunt?
JOB|37|19|Ostende nobis quid dicamus illi;nos disponere verba nescimus propter tenebras.
JOB|37|20|Quis narrabit ei, quae loquor?Et, si locutus fuerit, homo deglutietur.
JOB|37|21|At nunc non vident lucem:aer offuscatus est nubibus,sed ventus transiens fugabit eas.
JOB|37|22|Ab aquilone splendor auri venit;et circa Deum terribilis maiestas.
JOB|37|23|Omnipotentem attingere non possumus: magnus fortitudine;et iudicium et multam iustitiam deprimere non potest.
JOB|37|24|Ideo timebunt eum homines,non contemplabitur omnes, qui sibi videntur corde sapientes ".
JOB|38|1|Respondens autem Dominus Iob de turbine dixit:
JOB|38|2|" Quis est iste obscurans consiliumsermonibus imperitis?
JOB|38|3|Accinge sicut vir lumbos tuos;interrogabo te, et edoce me.
JOB|38|4|Ubi eras, quando ponebam fundamenta terrae?Indica mihi, si habes intellegentiam.
JOB|38|5|Quis posuit mensuras eius, si nosti?Vel quis tetendit super eam lineam?
JOB|38|6|Super quo bases illius solidatae sunt?Aut quis demisit lapidem angularem eius,
JOB|38|7|cum clamarent simul astra matutina,et iubilarent omnes filii Dei?
JOB|38|8|Quis conclusit ostiis mare,quando erumpebat quasi de visceribus procedens,
JOB|38|9|cum ponerem nubem vestimentum eiuset caligine illud quasi fascia obvolverem?
JOB|38|10|Definivi illud terminis meiset posui vectem et ostia
JOB|38|11|et dixi: Usque huc venies et non procedes ampliuset hic confringes tumentes fluctus tuos.
JOB|38|12|Numquid in diebus tuis praecepisti diluculoet assignasti aurorae locum suum,
JOB|38|13|et, cum extrema terrae teneres,excussi sunt impii ex ea?
JOB|38|14|Vertetur in lutum signatumet stabit sicut vestimentum.
JOB|38|15|Cohibetur ab impiis lux sua,et brachium excelsum confringetur.
JOB|38|16|Numquid ingressus es scaturigines mariset in novissimis abyssi deambulasti?
JOB|38|17|Numquid apertae sunt tibi portae mortis,et ostia tenebrosa vidisti?
JOB|38|18|Numquid considerasti latitudinem terrae?Indica mihi, si nosti omnia:
JOB|38|19|In qua via lux habitet,et tenebrarum quis locus sit;
JOB|38|20|ut ducas unumquodque ad terminos suoset intellegas semitas domus eius?
JOB|38|21|Novisti, nam tunc natus eras,et numerus dierum tuorum multus!
JOB|38|22|Numquid ingressus es thesauros nivisaut thesauros grandinis aspexisti,
JOB|38|23|quae praeparavi in tempus angustiae,in diem pugnae et belli?
JOB|38|24|Per quam viam spargitur lux,diffunditur ventus urens super terram?
JOB|38|25|Quis dedit vehementissimo imbri cursumet viam fulmini tonanti,
JOB|38|26|ut plueret super terram absque homine,in deserto, ubi nullus mortalium commoratur,
JOB|38|27|ut impleret inviam et desolatamet produceret herbas in terra arida?
JOB|38|28|Quis est pluviae pater,vel quis genuit stillas roris?
JOB|38|29|De cuius sinu egressa est glacies,et pruinam de caelo quis genuit?
JOB|38|30|In similitudinem lapidis aquae durantur,et superficies abyssi constringitur.
JOB|38|31|Numquid coniungere valebis nexus stellarum Pleiadumaut funiculum Arcturi poteris solvere?
JOB|38|32|Numquid produces Coronam in tempore suoet Ursam cum filiis ducis tu?
JOB|38|33|Numquid nosti leges caeliet pones scripturam eius in terra?
JOB|38|34|Numquid elevabis in nebula vocem tuam,et impetus aquarum operiet te?
JOB|38|35|Numquid mittes fulgura, et ibuntet dicent tibi: "Adsumus!"?
JOB|38|36|Quis posuit in visceribus ibis sapientiam,vel quis dedit gallo intellegentiam?
JOB|38|37|Quis recensebit nubes in sapientia,et utres caeli quis declinabit,
JOB|38|38|quando funditur pulvis in solidum,et glebae compinguntur?
JOB|38|39|Numquid capies leaenae praedamet animam catulorum eius implebis,
JOB|38|40|quando cubant in antriset in specubus insidiantur?
JOB|38|41|Quis praeparat corvo escam suam,quando pulli eius clamant ad Deum vagantes,eo quod non habeant cibos?
JOB|39|1|Numquid nosti tempus partus ibicum in petrisvel parturientes cervas observasti?
JOB|39|2|Dinumerasti menses conceptus earumet scisti tempus partus earum?
JOB|39|3|Incurvantur ad fetum et pariuntet fetus suos emittunt.
JOB|39|4|Impinguantur filii earum et adolescunt in campo,egrediuntur et non revertuntur ad eas.
JOB|39|5|Quis dimisit onagrum liberum,et vincula ipsius quis solvit?
JOB|39|6|Cui dedi in solitudine domumet tabernacula eius in terra salsuginis.
JOB|39|7|Contemnit multitudinem civitatis,clamorem exactoris non audit.
JOB|39|8|Explorat montes pascuae suaeet virentia quaeque perquirit.
JOB|39|9|Numquid volet taurus ferus servire tibiaut morabitur ad praesepe tuum?
JOB|39|10|Numquid alligabis taurum ferum ad arandum loro tuo,aut confringet glebas vallium post te?
JOB|39|11|Numquid fiduciam habebis in magna fortitudine eiuset derelinques ei labores tuos?
JOB|39|12|Numquid credes illi quod revertaturet sementem in aream tuam congreget?
JOB|39|13|Ala struthionis laeta est,penna vero ciconiae et avolat.
JOB|39|14|Quando derelinquit ova sua in terra,in pulvere calefiunt.
JOB|39|15|Obliviscitur quod pes conculcet ea,aut bestia agri conterat.
JOB|39|16|Duratur ad filios suos quasi non sint sui;frustra laborans nullo timore anxiatur.
JOB|39|17|Privavit enim eam Deus sapientianec dedit illi intellegentiam.
JOB|39|18|Cum tempus fuerit, in altum alas erigit,deridet equum et ascensorem eius.
JOB|39|19|Numquid praebebis equo fortitudinemaut circumdabis collo eius iubam?
JOB|39|20|Numquid suscitabis eum quasi locustas?Gloria hinnitus eius terror;
JOB|39|21|vallem ungula fodit, exsultat audacter,in occursum pergit armatis.
JOB|39|22|Contemnit pavorem nec territurneque cedit gladio.
JOB|39|23|Super ipsum sonabit pharetra,micat hasta et acinaces.
JOB|39|24|Fervens et fremens sorbet terramnec consistet, cum tubae sonaverit clangor.
JOB|39|25|Ubi audierit bucinam, dicit: "Uah!".Procul odoratur bellum,exhortationem ducum et ululatum exercitus.
JOB|39|26|Numquid per sapientiam tuam plumescit accipiter,expandens alas suas ad austrum?
JOB|39|27|Numquid ad praeceptum tuum elevabitur aquilaet in arduis ponet nidum suum?
JOB|39|28|In petris manetet in praeruptis silicibus commoraturatque in culmine et arce.
JOB|39|29|Inde contemplatur escam,et de longe oculi eius prospiciunt.
JOB|39|30|Pulli eius lambent sanguinem;et, ubicumque cadaver fuerit, statim adest ".
JOB|40|1|Et respondens Dominus locutus est ad Iob:
JOB|40|2|" Numquid contendit cum Omnipotente reprehensor?Qui arguit Deum, debet respondere ad ea ".
JOB|40|3|Respondens autem Iob Domino dixit:
JOB|40|4|" Ecce leviter locutus sum, quid respondebo tibi?Manum meam ponam super os meum.
JOB|40|5|Unum locutus sum, quod non repetam,et alterum, quibus ultra non addam ".
JOB|40|6|Respondens autem Dominus Iob de turbine dixit:
JOB|40|7|" Accinge sicut vir lumbos tuos;interrogabo te, et edoce me.
JOB|40|8|Numquid irritum facies iudicium meumet condemnabis me, ut tu iustificeris?
JOB|40|9|Et si habes brachium sicut Deuset si voce simili tonas?
JOB|40|10|Circumda tibi decorem et sublimitatem;gloria et decore induere.
JOB|40|11|Effunde vehementiam furoris tuiet respiciens omnem arrogantem humilia.
JOB|40|12|Respice cunctos superbos et confunde eoset contere impios in loco suo.
JOB|40|13|Absconde eos in pulvere simulet facies eorum claude in fovea;
JOB|40|14|et ego confiteborquod salvare te possit dextera tua.
JOB|40|15|Ecce Behemoth, quem feci tecum;fenum quasi bos comedit.
JOB|40|16|Fortitudo eius in lumbis eius,et virtus illius in umbilico ventris eius.
JOB|40|17|Stringit caudam suam quasi cedrum,nervi femorum eius perplexi sunt.
JOB|40|18|Ossa eius velut fistulae aeris,cartilago illius quasi laminae ferreae.
JOB|40|19|Ipse est principium viarum Dei;qui fecit eum, applicabit gladium eius.
JOB|40|20|Huic montes tributum ferunt,omnes bestiae agri ludunt ibi.
JOB|40|21|Sub lotis silvestribus dormit,in secreto calami et in locis umentibus;
JOB|40|22|loti silvestres umbra eum protegunt,circumdant eum salices torrentis.
JOB|40|23|Si fluvius intumescat, non tremit;securus est, si prorumpat fluctus ad os eius.
JOB|40|24|In oculis eius quis capiet eumet in sudibus perforabit nares eius?
JOB|40|25|An extrahere poteris Leviathan hamoet fune ligabis linguam eius?
JOB|40|26|Numquid pones iuncum in naribus eiusaut spina perforabis maxillam eius?
JOB|40|27|Numquid multiplicabit ad te precesaut loquetur tibi mollia?
JOB|40|28|Numquid feriet tecum pactum,et accipies eum servum sempiternum?
JOB|40|29|Numquid illudes ei quasi aviaut ligabis eum pro puellis tuis?
JOB|40|30|Speculabuntur super eum socii,divident illum negotiatores?
JOB|40|31|Numquid implebis telis pellem eiuset iaculo hamato piscium caput illius?
JOB|40|32|Pone super eum manum tuam;memento belli nec ultra addas.
JOB|41|1|Ecce spes eius frustrabitur eum,et aspectu eius praecipitabitur.
JOB|41|2|Nemo tam audax, ut suscitet eum.Quis enim resistere potest vultui eius?
JOB|41|3|Quis eum aggressus est et salvus fuit?Sub omni caelo quisnam?
JOB|41|4|Non tacebo super membra eiuset eloquar robur et gratiam struis.
JOB|41|5|Quis revelabit faciem indumenti eius,et duplicia mandibulae eius quis intrabit?
JOB|41|6|Portas vultus eius quis aperiet?Per gyrum dentium eius formido.
JOB|41|7|Corpus illius quasi scuta fusilia,compactum sigillo siliceo:
JOB|41|8|unum uni coniungitur,et ne spiraculum quidem incedit per ea;
JOB|41|9|unum alteri adhaeret,et tenentes se nequaquam separantur.
JOB|41|10|Sternutatio eius favillae ignis,et oculi eius ut palpebrae diluculi.
JOB|41|11|De ore eius lampades procedunt,sicut scintillae ignis emittuntur.
JOB|41|12|De naribus eius procedit fumus,sicut ollae succensae atque ferventis.
JOB|41|13|Halitus eius prunas ardere facit,et flamma de ore eius egreditur.
JOB|41|14|In collo eius morabitur fortitudo,et faciem eius praecedit angor.
JOB|41|15|Palearia eius cohaerentia sibicompressa non moventur.
JOB|41|16|Cor eius induratur tamquam lapiset duratur quasi mola inferior.
JOB|41|17|Cum surrexerit, tremunt forteset ab undis retrorsum convertuntur.
JOB|41|18|Qui impegerit in eum, gladius eius non stabitnec hasta neque pilum neque thorax;
JOB|41|19|reputat enim quasi paleas ferrumet quasi lignum putridum aes.
JOB|41|20|Non fugat eum vir sagittarius,in stipulam versi sunt ei lapides fundae.
JOB|41|21|Quasi stipulam aestimat fustemet deridet vibrantem acinacem.
JOB|41|22|Sub ipso acumina testae,et sternit tribula super lutum.
JOB|41|23|Fervescere facit quasi ollam profundumet mare ponit quasi vas unguentarium.
JOB|41|24|Post se illuminat semitam,aestimatur abyssus quasi canescens.
JOB|41|25|Non est super terram potestas, quae comparetur ei,qui factus est, ut nullum timeret.
JOB|41|26|Omne sublime videt:ipse est rex super universos filios superbiae ".
JOB|42|1|Respondens autem Iob Domino dixit:
JOB|42|2|" Scio quia omnia potes,et nulla te latet cogitatio.
JOB|42|3|Quis est iste, qui celat consiliumabsque scientia?Ideo insipienter locutus sumet mirabilia, quae excederent scientiam meam.
JOB|42|4|Audi, et ego loquar;interrogabo te, et responde mihi.
JOB|42|5|Auditu auris audivi te;nunc autem oculus meus videt te.
JOB|42|6|Idcirco ipse me reprehendoet ago paenitentiam in favilla et cinere ".
JOB|42|7|Postquam autem locutus est Dominus verba haec ad Iob, dixit ad Eliphaz Themanitem: " Iratus est furor meus in te et in duos amicos tuos, quoniam non estis locuti coram me rectum sicut servus meus Iob.
JOB|42|8|Sumite ergo vobis septem tauros et septem arietes et ite ad servum meum Iob et offerte holocaustum pro vobis; Iob autem servus meus orabit pro vobis. Faciem eius suscipiam, ut non vobis imputetur stultitia; neque enim locuti estis ad me recta sicut servus meus Iob ".
JOB|42|9|Abierunt ergo Eliphaz Themanites et Baldad Suhites et Sophar Naamathites et fecerunt, sicut locutus fuerat Dominus ad eos, et suscepit Dominus faciem Iob.
JOB|42|10|Dominus vertit sortem Iob, cum oraret ille pro amicis suis; et addidit Dominus omnia, quaecumque fuerant Iob, duplicia.
JOB|42|11|Venerunt autem ad eum omnes fratres sui et universae sorores suae et cuncti, qui noverant eum prius; et comederunt cum eo panem in domo eius et moverunt super eum caput et consolati sunt eum super omni malo, quod intulerat Dominus super eum; et dederunt ei unusquisque argenteum unum et inaurem auream unam.
JOB|42|12|Dominus autem benedixit novissimis Iob magis quam principio eius; et facta sunt ei quattuordecim milia ovium et sex milia camelorum et mille iuga boum et mille asinae.
JOB|42|13|Et fuerunt ei septem filii et tres filiae;
JOB|42|14|et vocavit nomen unius Columbam et nomen secundae Cassiam et nomen tertiae Cornustibii.
JOB|42|15|Non sunt autem inventae mulieres speciosae sicut filiae Iob in universa terra; deditque eis pater suus hereditatem inter fratres earum.
JOB|42|16|Vixit autem Iob post haec centum quadraginta annis et vidit filios suos et filios filiorum suorum usque ad quartam generationem; et mortuus est senex et plenus dierum.
