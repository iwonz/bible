PHIL|1|1|Paul and Timothy, servants of Christ Jesus, To all the saints in Christ Jesus who are at Philippi, with the overseers and deacons:
PHIL|1|2|Grace to you and peace from God our Father and the Lord Jesus Christ.
PHIL|1|3|I thank my God in all my remembrance of you,
PHIL|1|4|always in every prayer of mine for you all making my prayer with joy,
PHIL|1|5|because of your partnership in the gospel from the first day until now.
PHIL|1|6|And I am sure of this, that he who began a good work in you will bring it to completion at the day of Jesus Christ.
PHIL|1|7|It is right for me to feel this way about you all, because I hold you in my heart, for you are all partakers with me of grace, both in my imprisonment and in the defense and confirmation of the gospel.
PHIL|1|8|For God is my witness, how I yearn for you all with the affection of Christ Jesus.
PHIL|1|9|And it is my prayer that your love may abound more and more, with knowledge and all discernment,
PHIL|1|10|so that you may approve what is excellent, and so be pure and blameless for the day of Christ,
PHIL|1|11|filled with the fruit of righteousness that comes through Jesus Christ, to the glory and praise of God.
PHIL|1|12|I want you to know, brothers, that what has happened to me has really served to advance the gospel,
PHIL|1|13|so that it has become known throughout the whole imperial guard and to all the rest that my imprisonment is for Christ.
PHIL|1|14|And most of the brothers, having become confident in the Lord by my imprisonment, are much more bold to speak the word without fear.
PHIL|1|15|Some indeed preach Christ from envy and rivalry, but others from good will.
PHIL|1|16|The latter do it out of love, knowing that I am put here for the defense of the gospel.
PHIL|1|17|The former proclaim Christ out of rivalry, not sincerely but thinking to afflict me in my imprisonment.
PHIL|1|18|What then? Only that in every way, whether in pretense or in truth, Christ is proclaimed, and in that I rejoice. Yes, and I will rejoice,
PHIL|1|19|for I know that through your prayers and the help of the Spirit of Jesus Christ this will turn out for my deliverance,
PHIL|1|20|as it is my eager expectation and hope that I will not be at all ashamed, but that with full courage now as always Christ will be honored in my body, whether by life or by death.
PHIL|1|21|For to me to live is Christ, and to die is gain.
PHIL|1|22|If I am to live in the flesh, that means fruitful labor for me. Yet which I shall choose I cannot tell.
PHIL|1|23|I am hard pressed between the two. My desire is to depart and be with Christ, for that is far better.
PHIL|1|24|But to remain in the flesh is more necessary on your account.
PHIL|1|25|Convinced of this, I know that I will remain and continue with you all, for your progress and joy in the faith,
PHIL|1|26|so that in me you may have ample cause to glory in Christ Jesus, because of my coming to you again.
PHIL|1|27|Only let your manner of life be worthy of the gospel of Christ, so that whether I come and see you or am absent, I may hear of you that you are standing firm in one spirit, with one mind striving side by side for the faith of the gospel,
PHIL|1|28|and not frightened in anything by your opponents. This is a clear sign to them of their destruction, but of your salvation, and that from God.
PHIL|1|29|For it has been granted to you that for the sake of Christ you should not only believe in him but also suffer for his sake,
PHIL|1|30|engaged in the same conflict that you saw I had and now hear that I still have.
PHIL|2|1|So if there is any encouragement in Christ, any comfort from love, any participation in the Spirit, any affection and sympathy,
PHIL|2|2|complete my joy by being of the same mind, having the same love, being in full accord and of one mind.
PHIL|2|3|Do nothing from rivalry or conceit, but in humility count others more significant than yourselves.
PHIL|2|4|Let each of you look not only to his own interests, but also to the interests of others.
PHIL|2|5|Have this mind among yourselves, which is yours in Christ Jesus,
PHIL|2|6|who, though he was in the form of God, did not count equality with God a thing to be grasped,
PHIL|2|7|but made himself nothing, taking the form of a servant, being born in the likeness of men. And being found in human form,
PHIL|2|8|he humbled himself by becoming obedient to the point of death, even death on a cross.
PHIL|2|9|Therefore God has highly exalted him and bestowed on him the name that is above every name,
PHIL|2|10|so that at the name of Jesus every knee should bow, in heaven and on earth and under the earth,
PHIL|2|11|and every tongue confess that Jesus Christ is Lord, to the glory of God the Father.
PHIL|2|12|Therefore, my beloved, as you have always obeyed, so now, not only as in my presence but much more in my absence, work out your own salvation with fear and trembling,
PHIL|2|13|for it is God who works in you, both to will and to work for his good pleasure.
PHIL|2|14|Do all things without grumbling or questioning,
PHIL|2|15|that you may be blameless and innocent, children of God without blemish in the midst of a crooked and twisted generation, among whom you shine as lights in the world,
PHIL|2|16|holding fast to the word of life, so that in the day of Christ I may be proud that I did not run in vain or labor in vain.
PHIL|2|17|Even if I am to be poured out as a drink offering upon the sacrificial offering of your faith, I am glad and rejoice with you all.
PHIL|2|18|Likewise you also should be glad and rejoice with me.
PHIL|2|19|I hope in the Lord Jesus to send Timothy to you soon, so that I too may be cheered by news of you.
PHIL|2|20|For I have no one like him, who will be genuinely concerned for your welfare.
PHIL|2|21|They all seek their own interests, not those of Jesus Christ.
PHIL|2|22|But you know Timothy's proven worth, how as a son with a father he has served with me in the gospel.
PHIL|2|23|I hope therefore to send him just as soon as I see how it will go with me,
PHIL|2|24|and I trust in the Lord that shortly I myself will come also.
PHIL|2|25|I have thought it necessary to send to you Epaphroditus my brother and fellow worker and fellow soldier, and your messenger and minister to my need,
PHIL|2|26|for he has been longing for you all and has been distressed because you heard that he was ill.
PHIL|2|27|Indeed he was ill, near to death. But God had mercy on him, and not only on him but on me also, lest I should have sorrow upon sorrow.
PHIL|2|28|I am the more eager to send him, therefore, that you may rejoice at seeing him again, and that I may be less anxious.
PHIL|2|29|So receive him in the Lord with all joy, and honor such men,
PHIL|2|30|for he nearly died for the work of Christ, risking his life to complete what was lacking in your service to me.
PHIL|3|1|Finally, my brothers, rejoice in the Lord. To write the same things to you is no trouble to me and is safe for you.
PHIL|3|2|Look out for the dogs, look out for the evildoers, look out for those who mutilate the flesh.
PHIL|3|3|For we are the real circumcision, who worship by the Spirit of God and glory in Christ Jesus and put no confidence in the flesh-
PHIL|3|4|though I myself have reason for confidence in the flesh also. If anyone else thinks he has reason for confidence in the flesh, I have more:
PHIL|3|5|circumcised on the eighth day, of the people of Israel, of the tribe of Benjamin, a Hebrew of Hebrews; as to the law, a Pharisee;
PHIL|3|6|as to zeal, a persecutor of the church; as to righteousness, under the law blameless.
PHIL|3|7|But whatever gain I had, I counted as loss for the sake of Christ.
PHIL|3|8|Indeed, I count everything as loss because of the surpassing worth of knowing Christ Jesus my Lord. For his sake I have suffered the loss of all things and count them as rubbish, in order that I may gain Christ
PHIL|3|9|and be found in him, not having a righteousness of my own that comes from the law, but that which comes through faith in Christ, the righteousness from God that depends on faith-
PHIL|3|10|that I may know him and the power of his resurrection, and may share his sufferings, becoming like him in his death,
PHIL|3|11|that by any means possible I may attain the resurrection from the dead.
PHIL|3|12|Not that I have already obtained this or am already perfect, but I press on to make it my own, because Christ Jesus has made me his own.
PHIL|3|13|Brothers, I do not consider that I have made it my own. But one thing I do: forgetting what lies behind and straining forward to what lies ahead,
PHIL|3|14|I press on toward the goal for the prize of the upward call of God in Christ Jesus.
PHIL|3|15|Let those of us who are mature think this way, and if in anything you think otherwise, God will reveal that also to you.
PHIL|3|16|Only let us hold true to what we have attained.
PHIL|3|17|Brothers, join in imitating me, and keep your eyes on those who walk according to the example you have in us.
PHIL|3|18|For many, of whom I have often told you and now tell you even with tears, walk as enemies of the cross of Christ.
PHIL|3|19|Their end is destruction, their god is their belly, and they glory in their shame, with minds set on earthly things.
PHIL|3|20|But our citizenship is in heaven, and from it we await a Savior, the Lord Jesus Christ,
PHIL|3|21|who will transform our lowly body to be like his glorious body, by the power that enables him even to subject all things to himself.
PHIL|4|1|Therefore, my brothers, whom I love and long for, my joy and crown, stand firm thus in the Lord, my beloved.
PHIL|4|2|I entreat Euodia and I entreat Syntyche to agree in the Lord.
PHIL|4|3|Yes, I ask you also, true companion, help these women, who have labored side by side with me in the gospel together with Clement and the rest of my fellow workers, whose names are in the book of life.
PHIL|4|4|Rejoice in the Lord always; again I will say, Rejoice.
PHIL|4|5|Let your reasonableness be known to everyone. The Lord is at hand;
PHIL|4|6|do not be anxious about anything, but in everything by prayer and supplication with thanksgiving let your requests be made known to God.
PHIL|4|7|And the peace of God, which surpasses all understanding, will guard your hearts and your minds in Christ Jesus.
PHIL|4|8|Finally, brothers, whatever is true, whatever is honorable, whatever is just, whatever is pure, whatever is lovely, whatever is commendable, if there is any excellence, if there is anything worthy of praise, think about these things.
PHIL|4|9|What you have learned and received and heard and seen in me- practice these things, and the God of peace will be with you.
PHIL|4|10|I rejoiced in the Lord greatly that now at length you have revived your concern for me. You were indeed concerned for me, but you had no opportunity.
PHIL|4|11|Not that I am speaking of being in need, for I have learned in whatever situation I am to be content.
PHIL|4|12|I know how to be brought low, and I know how to abound. In any and every circumstance, I have learned the secret of facing plenty and hunger, abundance and need.
PHIL|4|13|I can do all things through him who strengthens me.
PHIL|4|14|Yet it was kind of you to share my trouble.
PHIL|4|15|And you Philippians yourselves know that in the beginning of the gospel, when I left Macedonia, no church entered into partnership with me in giving and receiving, except you only.
PHIL|4|16|Even in Thessalonica you sent me help for my needs once and again.
PHIL|4|17|Not that I seek the gift, but I seek the fruit that increases to your credit.
PHIL|4|18|I have received full payment, and more. I am well supplied, having received from Epaphroditus the gifts you sent, a fragrant offering, a sacrifice acceptable and pleasing to God.
PHIL|4|19|And my God will supply every need of yours according to his riches in glory in Christ Jesus.
PHIL|4|20|To our God and Father be glory forever and ever. Amen.
PHIL|4|21|Greet every saint in Christ Jesus. The brothers who are with me greet you.
PHIL|4|22|All the saints greet you, especially those of Caesar's household.
PHIL|4|23|The grace of the Lord Jesus Christ be with your spirit.
