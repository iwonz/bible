GAL|1|1|Paul, an apostle, (not of men, neither by man, but by Jesus Christ, and God the Father, who raised him from the dead;)
GAL|1|2|And all the brethren which are with me, unto the churches of Galatia:
GAL|1|3|Grace be to you and peace from God the Father, and from our Lord Jesus Christ,
GAL|1|4|Who gave himself for our sins, that he might deliver us from this present evil world, according to the will of God and our Father:
GAL|1|5|To whom be glory for ever and ever. Amen.
GAL|1|6|I marvel that ye are so soon removed from him that called you into the grace of Christ unto another gospel:
GAL|1|7|Which is not another; but there be some that trouble you, and would pervert the gospel of Christ.
GAL|1|8|But though we, or an angel from heaven, preach any other gospel unto you than that which we have preached unto you, let him be accursed.
GAL|1|9|As we said before, so say I now again, if any man preach any other gospel unto you than that ye have received, let him be accursed.
GAL|1|10|For do I now persuade men, or God? or do I seek to please men? for if I yet pleased men, I should not be the servant of Christ.
GAL|1|11|But I certify you, brethren, that the gospel which was preached of me is not after man.
GAL|1|12|For I neither received it of man, neither was I taught it, but by the revelation of Jesus Christ.
GAL|1|13|For ye have heard of my conversation in time past in the Jews' religion, how that beyond measure I persecuted the church of God, and wasted it:
GAL|1|14|And profited in the Jews' religion above many my equals in mine own nation, being more exceedingly zealous of the traditions of my fathers.
GAL|1|15|But when it pleased God, who separated me from my mother's womb, and called me by his grace,
GAL|1|16|To reveal his Son in me, that I might preach him among the heathen; immediately I conferred not with flesh and blood:
GAL|1|17|Neither went I up to Jerusalem to them which were apostles before me; but I went into Arabia, and returned again unto Damascus.
GAL|1|18|Then after three years I went up to Jerusalem to see Peter, and abode with him fifteen days.
GAL|1|19|But other of the apostles saw I none, save James the Lord's brother.
GAL|1|20|Now the things which I write unto you, behold, before God, I lie not.
GAL|1|21|Afterwards I came into the regions of Syria and Cilicia;
GAL|1|22|And was unknown by face unto the churches of Judaea which were in Christ:
GAL|1|23|But they had heard only, That he which persecuted us in times past now preacheth the faith which once he destroyed.
GAL|1|24|And they glorified God in me.
GAL|2|1|Then fourteen years after I went up again to Jerusalem with Barnabas, and took Titus with me also.
GAL|2|2|And I went up by revelation, and communicated unto them that gospel which I preach among the Gentiles, but privately to them which were of reputation, lest by any means I should run, or had run, in vain.
GAL|2|3|But neither Titus, who was with me, being a Greek, was compelled to be circumcised:
GAL|2|4|And that because of false brethren unawares brought in, who came in privily to spy out our liberty which we have in Christ Jesus, that they might bring us into bondage:
GAL|2|5|To whom we gave place by subjection, no, not for an hour; that the truth of the gospel might continue with you.
GAL|2|6|But of these who seemed to be somewhat, (whatsoever they were, it maketh no matter to me: God accepteth no man's person:) for they who seemed to be somewhat in conference added nothing to me:
GAL|2|7|But contrariwise, when they saw that the gospel of the uncircumcision was committed unto me, as the gospel of the circumcision was unto Peter;
GAL|2|8|(For he that wrought effectually in Peter to the apostleship of the circumcision, the same was mighty in me toward the Gentiles:)
GAL|2|9|And when James, Cephas, and John, who seemed to be pillars, perceived the grace that was given unto me, they gave to me and Barnabas the right hands of fellowship; that we should go unto the heathen, and they unto the circumcision.
GAL|2|10|Only they would that we should remember the poor; the same which I also was forward to do.
GAL|2|11|But when Peter was come to Antioch, I withstood him to the face, because he was to be blamed.
GAL|2|12|For before that certain came from James, he did eat with the Gentiles: but when they were come, he withdrew and separated himself, fearing them which were of the circumcision.
GAL|2|13|And the other Jews dissembled likewise with him; insomuch that Barnabas also was carried away with their dissimulation.
GAL|2|14|But when I saw that they walked not uprightly according to the truth of the gospel, I said unto Peter before them all, If thou, being a Jew, livest after the manner of Gentiles, and not as do the Jews, why compellest thou the Gentiles to live as do the Jews?
GAL|2|15|We who are Jews by nature, and not sinners of the Gentiles,
GAL|2|16|Knowing that a man is not justified by the works of the law, but by the faith of Jesus Christ, even we have believed in Jesus Christ, that we might be justified by the faith of Christ, and not by the works of the law: for by the works of the law shall no flesh be justified.
GAL|2|17|But if, while we seek to be justified by Christ, we ourselves also are found sinners, is therefore Christ the minister of sin? God forbid.
GAL|2|18|For if I build again the things which I destroyed, I make myself a transgressor.
GAL|2|19|For I through the law am dead to the law, that I might live unto God.
GAL|2|20|I am crucified with Christ: neverthless I live; yet not I, but Christ liveth in me: and the life which I now live in the flesh I live by the faith of the Son of God, who loved me, and gave himself for me.
GAL|2|21|I do not frustrate the grace of God: for if righteousness come by the law, then Christ is dead in vain.
GAL|3|1|O foolish Galatians, who hath bewitched you, that ye should not obey the truth, before whose eyes Jesus Christ hath been evidently set forth, crucified among you?
GAL|3|2|This only would I learn of you, Received ye the Spirit by the works of the law, or by the hearing of faith?
GAL|3|3|Are ye so foolish? having begun in the Spirit, are ye now made perfect by the flesh?
GAL|3|4|Have ye suffered so many things in vain? if it be yet in vain.
GAL|3|5|He therefore that ministereth to you the Spirit, and worketh miracles among you, doeth he it by the works of the law, or by the hearing of faith?
GAL|3|6|Even as Abraham believed God, and it was accounted to him for righteousness.
GAL|3|7|Know ye therefore that they which are of faith, the same are the children of Abraham.
GAL|3|8|And the scripture, foreseeing that God would justify the heathen through faith, preached before the gospel unto Abraham, saying, In thee shall all nations be blessed.
GAL|3|9|So then they which be of faith are blessed with faithful Abraham.
GAL|3|10|For as many as are of the works of the law are under the curse: for it is written, Cursed is every one that continueth not in all things which are written in the book of the law to do them.
GAL|3|11|But that no man is justified by the law in the sight of God, it is evident: for, The just shall live by faith.
GAL|3|12|And the law is not of faith: but, The man that doeth them shall live in them.
GAL|3|13|Christ hath redeemed us from the curse of the law, being made a curse for us: for it is written, Cursed is every one that hangeth on a tree:
GAL|3|14|That the blessing of Abraham might come on the Gentiles through Jesus Christ; that we might receive the promise of the Spirit through faith.
GAL|3|15|Brethren, I speak after the manner of men; Though it be but a man's covenant, yet if it be confirmed, no man disannulleth, or addeth thereto.
GAL|3|16|Now to Abraham and his seed were the promises made. He saith not, And to seeds, as of many; but as of one, And to thy seed, which is Christ.
GAL|3|17|And this I say, that the covenant, that was confirmed before of God in Christ, the law, which was four hundred and thirty years after, cannot disannul, that it should make the promise of none effect.
GAL|3|18|For if the inheritance be of the law, it is no more of promise: but God gave it to Abraham by promise.
GAL|3|19|Wherefore then serveth the law? It was added because of transgressions, till the seed should come to whom the promise was made; and it was ordained by angels in the hand of a mediator.
GAL|3|20|Now a mediator is not a mediator of one, but God is one.
GAL|3|21|Is the law then against the promises of God? God forbid: for if there had been a law given which could have given life, verily righteousness should have been by the law.
GAL|3|22|But the scripture hath concluded all under sin, that the promise by faith of Jesus Christ might be given to them that believe.
GAL|3|23|But before faith came, we were kept under the law, shut up unto the faith which should afterwards be revealed.
GAL|3|24|Wherefore the law was our schoolmaster to bring us unto Christ, that we might be justified by faith.
GAL|3|25|But after that faith is come, we are no longer under a schoolmaster.
GAL|3|26|For ye are all the children of God by faith in Christ Jesus.
GAL|3|27|For as many of you as have been baptized into Christ have put on Christ.
GAL|3|28|There is neither Jew nor Greek, there is neither bond nor free, there is neither male nor female: for ye are all one in Christ Jesus.
GAL|3|29|And if ye be Christ's, then are ye Abraham's seed, and heirs according to the promise.
GAL|4|1|Now I say, That the heir, as long as he is a child, differeth nothing from a servant, though he be lord of all;
GAL|4|2|But is under tutors and governors until the time appointed of the father.
GAL|4|3|Even so we, when we were children, were in bondage under the elements of the world:
GAL|4|4|But when the fulness of the time was come, God sent forth his Son, made of a woman, made under the law,
GAL|4|5|To redeem them that were under the law, that we might receive the adoption of sons.
GAL|4|6|And because ye are sons, God hath sent forth the Spirit of his Son into your hearts, crying, Abba, Father.
GAL|4|7|Wherefore thou art no more a servant, but a son; and if a son, then an heir of God through Christ.
GAL|4|8|Howbeit then, when ye knew not God, ye did service unto them which by nature are no gods.
GAL|4|9|But now, after that ye have known God, or rather are known of God, how turn ye again to the weak and beggarly elements, whereunto ye desire again to be in bondage?
GAL|4|10|Ye observe days, and months, and times, and years.
GAL|4|11|I am afraid of you, lest I have bestowed upon you labour in vain.
GAL|4|12|Brethren, I beseech you, be as I am; for I am as ye are: ye have not injured me at all.
GAL|4|13|Ye know how through infirmity of the flesh I preached the gospel unto you at the first.
GAL|4|14|And my temptation which was in my flesh ye despised not, nor rejected; but received me as an angel of God, even as Christ Jesus.
GAL|4|15|Where is then the blessedness ye spake of? for I bear you record, that, if it had been possible, ye would have plucked out your own eyes, and have given them to me.
GAL|4|16|Am I therefore become your enemy, because I tell you the truth?
GAL|4|17|They zealously affect you, but not well; yea, they would exclude you, that ye might affect them.
GAL|4|18|But it is good to be zealously affected always in a good thing, and not only when I am present with you.
GAL|4|19|My little children, of whom I travail in birth again until Christ be formed in you,
GAL|4|20|I desire to be present with you now, and to change my voice; for I stand in doubt of you.
GAL|4|21|Tell me, ye that desire to be under the law, do ye not hear the law?
GAL|4|22|For it is written, that Abraham had two sons, the one by a bondmaid, the other by a freewoman.
GAL|4|23|But he who was of the bondwoman was born after the flesh; but he of the freewoman was by promise.
GAL|4|24|Which things are an allegory: for these are the two covenants; the one from the mount Sinai, which gendereth to bondage, which is Agar.
GAL|4|25|For this Agar is mount Sinai in Arabia, and answereth to Jerusalem which now is, and is in bondage with her children.
GAL|4|26|But Jerusalem which is above is free, which is the mother of us all.
GAL|4|27|For it is written, Rejoice, thou barren that bearest not; break forth and cry, thou that travailest not: for the desolate hath many more children than she which hath an husband.
GAL|4|28|Now we, brethren, as Isaac was, are the children of promise.
GAL|4|29|But as then he that was born after the flesh persecuted him that was born after the Spirit, even so it is now.
GAL|4|30|Nevertheless what saith the scripture? Cast out the bondwoman and her son: for the son of the bondwoman shall not be heir with the son of the freewoman.
GAL|4|31|So then, brethren, we are not children of the bondwoman, but of the free.
GAL|5|1|Stand fast therefore in the liberty wherewith Christ hath made us free, and be not entangled again with the yoke of bondage.
GAL|5|2|Behold, I Paul say unto you, that if ye be circumcised, Christ shall profit you nothing.
GAL|5|3|For I testify again to every man that is circumcised, that he is a debtor to do the whole law.
GAL|5|4|Christ is become of no effect unto you, whosoever of you are justified by the law; ye are fallen from grace.
GAL|5|5|For we through the Spirit wait for the hope of righteousness by faith.
GAL|5|6|For in Jesus Christ neither circumcision availeth any thing, nor uncircumcision; but faith which worketh by love.
GAL|5|7|Ye did run well; who did hinder you that ye should not obey the truth?
GAL|5|8|This persuasion cometh not of him that calleth you.
GAL|5|9|A little leaven leaveneth the whole lump.
GAL|5|10|I have confidence in you through the Lord, that ye will be none otherwise minded: but he that troubleth you shall bear his judgment, whosoever he be.
GAL|5|11|And I, brethren, if I yet preach circumcision, why do I yet suffer persecution? then is the offence of the cross ceased.
GAL|5|12|I would they were even cut off which trouble you.
GAL|5|13|For, brethren, ye have been called unto liberty; only use not liberty for an occasion to the flesh, but by love serve one another.
GAL|5|14|For all the law is fulfilled in one word, even in this; Thou shalt love thy neighbour as thyself.
GAL|5|15|But if ye bite and devour one another, take heed that ye be not consumed one of another.
GAL|5|16|This I say then, Walk in the Spirit, and ye shall not fulfil the lust of the flesh.
GAL|5|17|For the flesh lusteth against the Spirit, and the Spirit against the flesh: and these are contrary the one to the other: so that ye cannot do the things that ye would.
GAL|5|18|But if ye be led of the Spirit, ye are not under the law.
GAL|5|19|Now the works of the flesh are manifest, which are these; Adultery, fornication, uncleanness, lasciviousness,
GAL|5|20|Idolatry, witchcraft, hatred, variance, emulations, wrath, strife, seditions, heresies,
GAL|5|21|Envyings, murders, drunkenness, revellings, and such like: of the which I tell you before, as I have also told you in time past, that they which do such things shall not inherit the kingdom of God.
GAL|5|22|But the fruit of the Spirit is love, joy, peace, longsuffering, gentleness, goodness, faith,
GAL|5|23|Meekness, temperance: against such there is no law.
GAL|5|24|And they that are Christ's have crucified the flesh with the affections and lusts.
GAL|5|25|If we live in the Spirit, let us also walk in the Spirit.
GAL|5|26|Let us not be desirous of vain glory, provoking one another, envying one another.
GAL|6|1|Brethren, if a man be overtaken in a fault, ye which are spiritual, restore such an one in the spirit of meekness; considering thyself, lest thou also be tempted.
GAL|6|2|Bear ye one another's burdens, and so fulfil the law of Christ.
GAL|6|3|For if a man think himself to be something, when he is nothing, he deceiveth himself.
GAL|6|4|But let every man prove his own work, and then shall he have rejoicing in himself alone, and not in another.
GAL|6|5|For every man shall bear his own burden.
GAL|6|6|Let him that is taught in the word communicate unto him that teacheth in all good things.
GAL|6|7|Be not deceived; God is not mocked: for whatsoever a man soweth, that shall he also reap.
GAL|6|8|For he that soweth to his flesh shall of the flesh reap corruption; but he that soweth to the Spirit shall of the Spirit reap life everlasting.
GAL|6|9|And let us not be weary in well doing: for in due season we shall reap, if we faint not.
GAL|6|10|As we have therefore opportunity, let us do good unto all men, especially unto them who are of the household of faith.
GAL|6|11|Ye see how large a letter I have written unto you with mine own hand.
GAL|6|12|As many as desire to make a fair shew in the flesh, they constrain you to be circumcised; only lest they should suffer persecution for the cross of Christ.
GAL|6|13|For neither they themselves who are circumcised keep the law; but desire to have you circumcised, that they may glory in your flesh.
GAL|6|14|But God forbid that I should glory, save in the cross of our Lord Jesus Christ, by whom the world is crucified unto me, and I unto the world.
GAL|6|15|For in Christ Jesus neither circumcision availeth any thing, nor uncircumcision, but a new creature.
GAL|6|16|And as many as walk according to this rule, peace be on them, and mercy, and upon the Israel of God.
GAL|6|17|From henceforth let no man trouble me: for I bear in my body the marks of the Lord Jesus.
GAL|6|18|Brethren, the grace of our Lord Jesus Christ be with your spirit. Amen.
