2COR|1|1|奉上帝旨意作基督耶稣使徒的 保罗 和弟兄 提摩太 ，写信给在 哥林多 上帝的教会和全 亚该亚 的众圣徒。
2COR|1|2|愿恩惠、平安 从我们的父上帝和主耶稣基督归给你们！
2COR|1|3|愿颂赞归于上帝—我们主耶稣基督的父；他是发慈悲的父，赐各样安慰的上帝。
2COR|1|4|我们在一切患难中，他安慰我们，使我们能用上帝所赐的安慰去安慰那些遭各样患难的人。
2COR|1|5|正如我们跟基督同受许多苦楚，我们也靠基督得许多安慰。
2COR|1|6|如果我们受患难，那是为使你们得安慰，得拯救；如果我们得安慰，那也是为使你们得安慰，这安慰能使你们忍受我们所受同样的苦楚。
2COR|1|7|我们为你们所存的盼望是确定的，因为知道你们分担了我们的痛苦，也要分享我们的安慰。
2COR|1|8|弟兄们，我们不要你们不知道，我们从前在 亚细亚 遭遇苦难，因受到无法忍受的压力，甚至连活命的指望都没有了。
2COR|1|9|自己心里也断定是必死无疑，这是要使我们不依靠自己，只依靠使死人复活的上帝。
2COR|1|10|他曾救我们脱离那极大的死亡，他要继续救我们，而且我们指望他将来还要救我们。
2COR|1|11|你们也要一同用祈祷来帮助我们，好使许多人为我们感恩，因着他们许多的祷告，我们获得了恩赐。
2COR|1|12|我们所夸的是：我们在世为人，特别是跟你们的关系，是凭着上帝所赐的坦率和真诚，不是靠人的聪明，而是靠上帝的恩惠；这是我们的良心可以作证的。
2COR|1|13|我们现在写给你们的话，无非是你们所能诵读、所能明白的，我也盼望你们真能彻底明白。
2COR|1|14|你们已经有几分认识我们，在我们主耶稣 的日子，你们会以我们为荣，正像我们也以你们为荣。
2COR|1|15|既然我这样深信，早就有意先到你们那里去，让你们得加倍的益处。
2COR|1|16|我要路过你们那里往 马其顿 去，再从 马其顿 回到你们那里，让你们给我送行往 犹太 去。
2COR|1|17|我有此意，难道是反覆不定吗？难道我的意愿是从私欲起的，以致我忽是忽非吗？
2COR|1|18|我指着信实的上帝说，我们向你们所传的道并非又是又非的。
2COR|1|19|因为，我、 西拉 和 提摩太 在你们中间传上帝的儿子耶稣基督，从没有“又是又非”的；在他只有一个“是”。
2COR|1|20|上帝的应许，不论有多少，在基督都是“是”的。所以，我们藉着他说“阿们”，使上帝因我们得荣耀。
2COR|1|21|那在基督里坚固我们和你们，并且膏抹我们的，就是上帝。
2COR|1|22|他在我们身上盖了印，并赐圣灵在我们心里作凭据。
2COR|1|23|我指着我的性命求告上帝作证，我没有再往 哥林多 去是为了要宽容你们。
2COR|1|24|我们并不是要控制你们的信心，而是要作你们的同工，让你们得快乐，因为你们在信仰上已经站得稳了。
2COR|2|1|我自己定了主意，下次不再带着悲伤到你们那里去。
2COR|2|2|我若使你们悲伤，除了因我而使他悲伤的那人以外，谁能使我喜乐呢？
2COR|2|3|我曾把这事写给你们，免得我到的时候，那该令我喜乐的人反倒令我悲伤。我也深信，你们众人都以我的喜乐为自己的喜乐。
2COR|2|4|我先前忧心忡忡、眼泪汪汪地给你们写了信，并非要使你们悲伤，而是要你们知道我格外疼爱你们。
2COR|2|5|如果有人使人悲伤，他不但使我悲伤，也是使你们众人有些悲伤。我说有些，恐怕说得太重了。
2COR|2|6|这样的人受了大多数人的责备也就够了，
2COR|2|7|倒不如赦免他，安慰他，免得他过分悲伤，甚至受不了啦！
2COR|2|8|所以，我劝你们，要向他肯定你们的爱心。
2COR|2|9|为此，我先前也写信给你们，正是要考验你们，看你们是否在一切事上都顺从我。
2COR|2|10|你们赦免谁，我也赦免谁。我若有所赦免，是在基督面前为你们的缘故赦免的，
2COR|2|11|免得撒但趁着机会胜过我们，因我们并非不知道他的诡计。
2COR|2|12|我从前为基督的福音到了 特罗亚 ，主给我开了门。
2COR|2|13|那时，因为没有遇见我的弟兄 提多 ，我心里不安，就辞别那里的人，往 马其顿 去了。
2COR|2|14|感谢上帝！他常率领我们在基督里得胜，并藉着我们在各处显扬那因认识基督而有的香气。
2COR|2|15|因为无论在得救的人或在灭亡的人当中，我们都是基督馨香之气，是献给上帝的。
2COR|2|16|对灭亡的人，这是死而又死的气味；对得救的人，这是生而又生的气味。这些事谁能当得起呢？
2COR|2|17|我们不像许多人，把上帝的道当商品贩卖，而是由于真诚，而是受命于上帝，在上帝面前凭着基督讲道。
2COR|3|1|难道我们又开始推荐自己吗？难道我们像某些人那样要用人的推荐信介绍给你们，或用你们的推荐信给人吗？
2COR|3|2|你们就是我们的推荐信，写在我们心里，被众人所知道、所诵读的，
2COR|3|3|而你们显明自己是基督的书信，藉着我们写成的。不是用墨写的，而是用永生上帝的灵写的；不是写在石版上，而是写在心版上的。
2COR|3|4|我们藉着基督才对上帝有这样的信心。
2COR|3|5|并不是我们凭自己配做什么事，我们之所以配做是出于上帝；
2COR|3|6|他使我们能配作新约的执事，不是文字上的约，而是圣灵的约；因为文字使人死，圣灵能使人活。
2COR|3|7|那用字刻在石头上属死的事奉尚且有荣光，以致 以色列 人因 摩西 脸上那逐渐褪色的荣光不能定睛看他的脸，
2COR|3|8|那属圣灵的事奉不是更有荣光吗？
2COR|3|9|若是那使人定罪的事奉有荣光，那使人称义的事奉的荣光就越发大了。
2COR|3|10|那从前有荣光的，因这更大的荣光，就算不得有荣光了；
2COR|3|11|若是那逐渐褪色的有荣光，这长存的就更有荣光了。
2COR|3|12|既然我们有这样的盼望，就大有胆量，
2COR|3|13|不像 摩西 将面纱蒙在脸上，使 以色列 人不能定睛看到那逐渐褪色的荣光的结局。
2COR|3|14|但他们的心地刚硬，直到今日诵读旧约的时候，这同样的面纱还没有揭去；因为这面纱在基督里才被废去。
2COR|3|15|然而直到今日，每逢诵读 摩西 书的时候，面纱还在他们心上。
2COR|3|16|但他们的心何时归向主，面纱就何时除去。
2COR|3|17|主就是那灵；主的灵在哪里，哪里就有自由。
2COR|3|18|既然我们众人以揭去面纱的脸得以看见 主的荣光，好像从镜子里返照，就变成了与主有同样的形像，荣上加荣，如同从主的灵 变成的。
2COR|4|1|所以，既然我们蒙怜悯受了这事奉的责任，就不丧胆，
2COR|4|2|反而把那些暗昧可耻的事弃绝了，不行诡诈，不曲解上帝的道，只将真理显扬出来，好在上帝面前把自己推荐给各人的良心。
2COR|4|3|即使我们的福音被遮蔽，那只是对灭亡的人遮蔽。
2COR|4|4|这些不信的人被这世界的神明弄瞎了心眼，使他们看不见基督荣耀的福音。基督本是上帝的像。
2COR|4|5|我们不是传自己，而是传耶稣基督为主，并且自己因耶稣作你们的仆人。
2COR|4|6|那吩咐光从黑暗里照出来的上帝已经照在我们心里，使我们知道上帝荣耀的光显在耶稣基督的脸上。
2COR|4|7|我们有这宝贝放在瓦器里，为要显明这莫大的能力是出于上帝，不是出于我们。
2COR|4|8|我们处处受困，却不被捆住；内心困扰，却没有绝望；
2COR|4|9|遭受迫害，却不被撇弃；击倒在地，却不致灭亡。
2COR|4|10|我们身上常带着耶稣的死，使耶稣的生也在我们身上显明。
2COR|4|11|因为我们这活着的人常为耶稣被置于死地，使耶稣的生命在我们这必死的人身上显明出来。
2COR|4|12|这样看来，死是在我们身上运作，生却在你们身上运作。
2COR|4|13|但我们既然有从同一位灵而来的信心，正如经上记着：“我信，故我说话”，我们也信，所以也说话；
2COR|4|14|因为知道，那使主耶稣复活的也必使我们与耶稣一同复活，并且使我们与你们一起站在他面前。
2COR|4|15|凡事都是为了你们，好使恩惠既藉着更多的人而加增，感恩也格外显多，好归荣耀给上帝。
2COR|4|16|所以，我们不丧胆。虽然我们外在的人日渐朽坏，内在的人却日日更新。
2COR|4|17|我们这短暂而轻微的苦楚要为我们成就极重、无比、永远的荣耀。
2COR|4|18|因为我们不是顾念看得见的，而是顾念看不见的；原来看得见的是暂时的，看不见的才是永远的。
2COR|5|1|因为我们知道，我们这地上的帐篷若拆毁了，我们将有上帝所造的居所，不是人手所造的，而是在天上永存的。
2COR|5|2|我们在这帐篷里叹息，渴望得到那从天上来的居所，好像穿上衣服；
2COR|5|3|倘若脱下也 不至于赤身了。
2COR|5|4|其实，我们在这帐篷里的人劳苦叹息，并不是愿意脱下地上的帐篷，而是愿意穿上天上的居所，好使这必死的被生命吞灭了。
2COR|5|5|那为我们安排这事的是上帝，他赐给我们圣灵作凭据 。
2COR|5|6|所以，我们总是勇敢的，并且知道，只要我们住在这身体内就是离开了主。
2COR|5|7|因为我们行事为人是凭着信心，不是凭着眼见。
2COR|5|8|我们勇敢，更情愿离开身体，与主同住。
2COR|5|9|所以，无论是住在身内或住在身外，我们都立了志向要得主的喜悦。
2COR|5|10|因为我们众人必须站在基督审判台前受审，为使各人按着本身所行的，或善或恶受报。
2COR|5|11|既然我们知道主是可畏的，就劝导人；但是上帝是认识我们的，我盼望你们的良心也认识我们。
2COR|5|12|我们不是向你们再推荐自己，而是要让你们有夸耀我们的机会，使你们好面对那凭外貌、不凭内心夸耀的人。
2COR|5|13|如果我们癫狂，是为上帝；如果我们清醒，是为你们。
2COR|5|14|原来基督的爱激励我们；因我们这样断定，一人既替众人死了，众人就都死了。
2COR|5|15|并且他替众人死，是叫那些活着的人不再为自己活，乃为替他们死而复活的主活。
2COR|5|16|所以，从今以后，我们不再按照人的看法来认识人，纵使我们曾经按照人的看法认识基督，如今却不再这样认识他了。
2COR|5|17|所以，若有人在基督里，他就是新造的人：旧事已过，都变成新的了。
2COR|5|18|一切都是出于上帝；他藉着基督使我们与他和好，又将劝人与他和好的使命赐给我们。
2COR|5|19|这就是：上帝在基督里使世人与自己和好，不将他们的过犯归到他们身上，并且将这和好的信息托付了我们。
2COR|5|20|所以，我们作基督的特使，就好像上帝藉我们劝你们一般。我们替基督求你们，与上帝和好吧！
2COR|5|21|上帝使那无罪 的，替我们成为罪，好使我们在他里面成为上帝的义。
2COR|6|1|我们与上帝同工的也劝你们，不可白受他的恩典；
2COR|6|2|因为他说： “在悦纳的时候，我应允了你； 在拯救的日子，我帮助了你。” 看哪，现在正是悦纳的时候！看哪，现在正是拯救的日子！
2COR|6|3|我们不在任何事上妨碍任何人，免得这使命被人毁谤；
2COR|6|4|反倒在各样的事上表明自己是上帝的用人：就如在持久的忍耐、患难、困苦、灾难、
2COR|6|5|鞭打、监禁、动乱、劳碌、失眠、饥饿、
2COR|6|6|廉洁、知识、坚忍、恩慈、圣灵的感化、无伪的爱心、
2COR|6|7|真实的言语、上帝的大能、藉着仁义的兵器在左在右、
2COR|6|8|荣誉或羞辱、恶名或美名。我们似乎是诱惑人的，却是诚实的；
2COR|6|9|似乎不为人所知，却是人所共知；似乎是死了，却是活着；似乎受惩罚，却没有被处死；
2COR|6|10|似乎忧愁，却常有喜乐；似乎贫穷，却使许多人富足；似乎一无所有，却样样都有。
2COR|6|11|哥林多 人哪，我们对你们，口是诚实的，心是宽宏的。
2COR|6|12|你们的狭窄不是由于我们，而是由于你们自己的心肠狭窄。
2COR|6|13|你们也要照样用宽宏的心报答我；我这话正像对自己的孩子说的。
2COR|6|14|你们不要和不信的人同负一轭。义和不义有什么相关？光明和黑暗有什么相连？
2COR|6|15|基督和 彼列 有什么相和？信主的和不信主的有什么相干？
2COR|6|16|上帝的殿和偶像有什么相同？因为我们是永生上帝的殿，就如上帝曾说： “我要在他们中间居住来往； 我要作他们的上帝， 他们要作我的子民。”
2COR|6|17|所以主说： “你们务要从他们中间出来， 跟他们分别； 不要沾不洁净的东西， 我就收纳你们。
2COR|6|18|我要作你们的父， 你们要作我的儿女。 这是全能的主说的。”
2COR|7|1|所以，亲爱的，既然我们有这样的应许，就当洁净自己，除去身体和灵魂一切的污秽，藉着敬畏上帝，得以成圣。
2COR|7|2|宽宏大量地接纳我们吧！我们未曾亏负谁，未曾败坏谁，未曾占谁的便宜。
2COR|7|3|我说这话，不是要定你们的罪，我已经说过，你们常在我们心里，我们情愿与你们同生共死。
2COR|7|4|我对你们很是放心，多多夸耀你们；我满有安慰，在我们一切患难中格外喜乐。
2COR|7|5|我们从前到了 马其顿 的时候，身体没有丝毫安宁，反而到处遭患难，外有纷争，内有惧怕。
2COR|7|6|但那安慰灰心之人的上帝藉着 提多 来安慰了我们；
2COR|7|7|不但藉着他来，也藉着他从你们所得的安慰安慰了我们，因为他把你们的思念，你们的哀恸，你们对我的热忱，都告诉了我，使我更加欢喜。
2COR|7|8|即使我先前那封信使你们忧愁，后来我曾懊悔，如今却不懊悔；因为我知道，那封信使你们忧愁，不过是暂时的。
2COR|7|9|如今我欢喜，不是因你们曾忧愁，而是因忧愁导致你们的悔改。你们依着上帝的意思忧愁，凡事就不至于因我们受亏损了。
2COR|7|10|因为依着上帝的意思而忧愁，就生出没有懊悔的悔改来，以致得救；但世俗的忧愁叫人死。
2COR|7|11|你看，你们依着上帝的意思而忧愁，这在你们当中产生了何等的殷勤、甚至辩白、甚至愤慨、甚至恐惧、甚至渴望、甚至热忱、甚至责罚。在这一切事上，你们都表明自己是无可指责的。
2COR|7|12|所以，虽然我从前写信给你们，却不是为那亏负人的，也不是为那受人亏负的，而是要在上帝面前把你们顾念我们的热忱表现出来。
2COR|7|13|因此，我们得了安慰。 在我们所得的安慰之外，又因你们众人使 提多 心里畅快喜乐，我们就更加欢喜了。
2COR|7|14|我若对 提多 夸奖过你们什么，也不觉得惭愧，因为我对 提多 夸奖你们的话是真的，正如我对你们所说的话也向来都是真的。
2COR|7|15|提多 一想起你们众人的顺服，怎样恐惧战兢地接待他，他爱你们的心就越发热切了。
2COR|7|16|我如今欢喜，因为我在一切事上对你们有信心。
2COR|8|1|弟兄们，我们要把上帝赐给 马其顿 众教会的恩惠告诉你们：
2COR|8|2|他们在患难中受大考验的时候，仍然满有喜乐，在极度贫穷中还格外显出他们乐捐的慷慨。
2COR|8|3|我可以证明，他们是按着能力，而且超过了能力来捐助，主动
2COR|8|4|再三恳求我们，准他们在这供给圣徒的善事上有份；
2COR|8|5|并且他们所做的，不但照我们所期望的，更照上帝的旨意先把自己献给主，又给了我们。
2COR|8|6|因此，我们劝 提多 ，既然在你们中间开始这慈善的事，就当把它办成。
2COR|8|7|既然你们在信心、口才、知识、万分的热忱，以及我们对你们 的爱心上，都胜人一等，那么，当在这慈善的事上也要胜人一等。
2COR|8|8|我说这话，并不是命令你们，而是藉着别人的热忱来考验你们爱心的真诚。
2COR|8|9|你们知道我们主耶稣基督的恩典：他本是富足，却为你们成了贫穷，好使你们因他的贫穷而成为富足。
2COR|8|10|我在这事上把我的意见告诉你们，是对你们有益，因为你们开始办这事，而且起此心意已经有一年了。
2COR|8|11|如今就当办成这事，既然有愿做的心，也当照你们所有的去办成。
2COR|8|12|因为人只要有愿做的心，必照他所有的蒙悦纳，并不是照他所没有的。
2COR|8|13|我不是要别人轻松，你们受累，而是要均匀：
2COR|8|14|就是要你们现在的富余补他们的不足，使他们的富余将来也可以补你们的不足，这就均匀了。
2COR|8|15|如经上所记： 多收的没有余， 少收的也没有缺。
2COR|8|16|感谢上帝，把我对你们的热忱同样放在 提多 心里。
2COR|8|17|他固然听了我的劝告，但自己更加热心，自愿往你们那里去。
2COR|8|18|我们还差遣一位弟兄和他同去，这人在传福音的事上得了众教会的称赞；
2COR|8|19|不但这样，他也被众教会选派跟我们同行，把所交托我们的这捐款送到了，为的是荣耀主，也表明我们的好意。
2COR|8|20|我们这样做，免得有人因我们收的捐款多而挑剔我们。
2COR|8|21|我们留心做好事，不但在主面前，就是在人面前也是这样。
2COR|8|22|我们又差遣一位弟兄同去。这人的热忱，我们在许多事上屡次考验过，现在他因为深深信任你们，就更加热心了。
2COR|8|23|至于 提多 ，他是我的伙伴，为服事你们作我的同工。至于那两位弟兄，他们是众教会的使者，是基督的荣耀。
2COR|8|24|所以，你们务要在众教会面前向他们显明你们的爱心和我所夸奖你们的凭据。
2COR|9|1|关于供给圣徒的事，我本来不必写信给你们；
2COR|9|2|因为我知道你们的好意，常对 马其顿 人夸奖你们，说 亚该亚 人预备好已经有一年了。你们的热心感动了许多人。
2COR|9|3|但我差遣那几位弟兄去，要使你们照我的话预备妥当，免得我们在这事上夸奖你们的话落了空。
2COR|9|4|万一有 马其顿 人与我同去，见你们没有预备好，就使我们所确信的反成了羞愧；你们的羞愧更不用说了。
2COR|9|5|因此，我想必须鼓励那几位弟兄先到你们那里去，把从前所应许的捐款预备妥当，好显出你们所捐的是出于乐意，不是出于勉强。
2COR|9|6|还有一点：“少种的少收；多种的多收。”
2COR|9|7|各人要随心所愿，不要为难，不要勉强，因为上帝爱乐捐的人。
2COR|9|8|上帝能将各样的恩惠多多加给你们，使你们凡事常常充足，能多做各样善事。
2COR|9|9|如经上所记： “他施舍，周济贫穷； 他的义行存到永远。”
2COR|9|10|那赐种子给撒种的，赐粮食给人吃的，必多多加给你们种地的种子，又增添你们仁义的果子。
2COR|9|11|你们必凡事富足，能多多施舍，使人藉着我们而生感谢上帝的心。
2COR|9|12|因为办这供给的事，不但补圣徒的缺乏，而且使许多人对上帝充满更多的感谢。
2COR|9|13|他们从这供给的事上得了凭据，知道你们宣认基督，顺服他的福音，慷慨捐助给他们和众人，把荣耀归给上帝。
2COR|9|14|他们也因上帝极大的恩赐显在你们身上而切切想念你们，为你们祈祷。
2COR|9|15|感谢上帝，因他有说不尽的恩赐！
2COR|10|1|我－ 保罗 与你们见面的时候是温和的，不在你们那里的时候向你们是勇敢的，如今亲自藉着基督的温柔和慈祥劝你们。
2COR|10|2|有人认为我们是凭着血气行事，我认为必须敢于对付这等人；我但求在那里的时候，不必这样勇敢。
2COR|10|3|我们虽然在血气中行事，却不凭着血气争战。
2COR|10|4|因为我们争战的兵器本不是属血气的，而是凭着上帝的能力，能够攻破坚固的营垒。我们攻破各样的计谋，
2COR|10|5|和各样拦阻人认识上帝的高垒，又夺回人心来顺服基督。
2COR|10|6|我已经预备好了，等你们完全顺服的时候来惩罚所有不顺服的人。
2COR|10|7|你们只看事情的外表。倘若有人自信是属基督的，他要再想想，他属基督，我们也属基督。
2COR|10|8|主赐给我们权柄，是要造就你们，并不是要拆毁你们；我就是为这权柄稍微夸口也不觉得惭愧。
2COR|10|9|我说这话，免得你们以为我写信是要恐吓你们。
2COR|10|10|因为有人说：“他信上的语气既严厉又强硬，他本人却软弱无能，言语粗俗。”
2COR|10|11|这等人当明白，我们不在那里时信上怎么说，见面时也必怎么做。
2COR|10|12|因为我们不敢将自己和某些自我推荐的人并列相比；他们用自己度量自己，用自己比较自己，是不明智的。
2COR|10|13|我们不愿意过分夸口，但是我们只在上帝划定的界限内夸口。这界限甚至扩展到你们那里。
2COR|10|14|我们扩展到你们那里时并没有越过了自己的界限，其实我们是首先到你们那里传基督福音的。
2COR|10|15|我们不靠别人所劳碌的过分夸口；我们只希望你们信心增长的时候，所划定给我们的范围也能够因着你们更加扩展，
2COR|10|16|使福音得以传到你们以外的地方，而不在别人的范围之内，以别人所成就的事夸口。
2COR|10|17|但“要夸耀的，该夸耀主”。
2COR|10|18|因为蒙悦纳的，不是自我称许的，而是主所称许的。
2COR|11|1|但愿你们容忍我小小的愚蠢；请你们务必容忍我。
2COR|11|2|我以上帝嫉妒的爱来爱你们，因为我曾把你们许配给一个丈夫，要把你们如同贞洁的童女献给基督。
2COR|11|3|我只怕你们的心偏邪了，失去那向基督所献诚恳贞洁 的心，就像蛇用诡诈诱惑了 夏娃 一样。
2COR|11|4|假如有人来，传另一个耶稣，不是我们所传过的；或者你们另受一个灵，不是你们所受过的圣灵；或者接纳另一个福音，不是你们所接纳过的；你们居然容忍了！
2COR|11|5|但我想，我一点也不在那些超级使徒以下。
2COR|11|6|虽然我不擅长说话，我的知识却不如此。这点我们已经在每一方面各样事上向你们表明了。
2COR|11|7|我贬低自己，为了使你们高升，因为我白白地传上帝的福音给你们，难道这算是我犯了错吗？
2COR|11|8|我剥夺了别的教会，向他们取了报酬来效劳你们。
2COR|11|9|我在你们那里有缺乏的时候，并没有连累你们一个人，因为我所缺乏的，那些从 马其顿 来的弟兄都补足了。我向来凡事谨慎，将来也必谨慎，总不要连累你们。
2COR|11|10|既有基督的真诚在我里面，在 亚该亚 一带地方就没有人能阻止我这样自夸。
2COR|11|11|为什么呢？是因我不爱你们吗？上帝知道，我爱你们！
2COR|11|12|我现在所做的，将来还要做，为要断绝那些寻机会之人的机会，不让他们在所夸耀的事上被人认为与我们一样。
2COR|11|13|那样的人是假使徒，行事诡诈，装作基督的使徒。
2COR|11|14|这也不足为奇，因为连撒但也装作光明的天使。
2COR|11|15|所以，他的差役若装作公义的差役也没有什么大不了。他们的结局必然跟他们的行为相符。
2COR|11|16|我再说，谁都不可把我看作愚蠢的；即使你们把我当作愚蠢人，那么，也让我稍微夸夸口吧。
2COR|11|17|我说的话不是奉主的权柄说的，而是像愚蠢人具有自信地放胆夸口。
2COR|11|18|既然有好些人凭着血气在夸口，我也要夸口了。
2COR|11|19|你们是聪明人，竟能甘心容忍愚蠢人！
2COR|11|20|假若有人奴役你们，或侵吞你们，或压榨你们，或侮辱你们，或打你们的脸，你们居然都能容忍。
2COR|11|21|说来惭愧，在这方面好像我们是太软弱了。 然而，我说句蠢话，人在什么事上敢夸口，我也敢夸口。
2COR|11|22|他们是 希伯来 人吗？我也是。他们是 以色列 人吗？我也是。他们是 亚伯拉罕 的后裔吗？我也是。
2COR|11|23|他们是基督的用人吗？我说句狂话，我更是。我比他们忍受更多劳苦，坐过更多次监牢，受过无数次的鞭打，常常冒死。
2COR|11|24|我被 犹太 人鞭打五次，每次四十减去一下；
2COR|11|25|被棍打了三次，被石头打了一次，遭海难三次，一昼一夜在深海里挣扎。
2COR|11|26|我又屡次行远路，遭江河的危险，盗贼的危险，同族人的危险，外族人的危险，城里的危险，旷野的危险，海中的危险，假弟兄的危险。
2COR|11|27|我劳碌困苦，常常失眠，又饥又渴，忍饥耐寒，赤身露体。
2COR|11|28|除了这些外表的事以外，我还有为众教会操心的事天天压在我身上。
2COR|11|29|有谁软弱，我不软弱呢？有谁跌倒，我不焦急呢？
2COR|11|30|我若必须夸口，就夸我软弱的事好了。
2COR|11|31|那永远可称颂之主耶稣的父上帝知道我不说谎。
2COR|11|32|在 大马士革 的 亚哩达 王手下的提督把守 大马士革城 ，要捉拿我，
2COR|11|33|我被人用筐子从城墙上的窗口缒下，逃脱了他的手。
2COR|12|1|虽然自夸无益，我还是不得不夸。我现在要提到主的异象和启示。
2COR|12|2|我认识一个在基督里的人，他在十四年前被提到第三层天上去；或在身内，我不知道，或在身外，我也不知道，只有上帝知道。
2COR|12|3|我认识的这样的一个人—或在身内，或在身外，我都不知道，只有上帝知道—
2COR|12|4|他被提到乐园里，听见隐秘的言语，是人不可说的。
2COR|12|5|为这人，我要夸口；但是为我自己，除了我的软弱以外，我并不夸口。
2COR|12|6|就是我愿意夸口也不算狂，因为我会说实话；只是我绝口不谈，恐怕有人把我看得太高了，过于他在我身上所看见所听见的；
2COR|12|7|又恐怕我因所得的启示太高深，就过于高抬自己，所以 有一根刺加在我身上，就是撒但的差役来折磨我，免得我过于高抬自己。
2COR|12|8|为了这事，我曾三次求主使这根刺离开我。
2COR|12|9|他对我说：“我的恩典是够你用的，因为我的能力是在人的软弱上显得完全。”所以，我更喜欢夸耀自己的软弱，好使基督的能力覆庇我。
2COR|12|10|为基督的缘故，我以软弱、凌辱、艰难、迫害、困苦为可喜乐的事；因为我什么时候软弱，什么时候就刚强了。
2COR|12|11|我成了愚蠢人，是被你们逼出来的，因为我本该被你们赞许才是。虽然我算不了什么，却没有一件事在那些超级使徒以下。
2COR|12|12|我在你们中间，用百般的忍耐，藉着神迹、奇事、异能显出使徒的凭据来。
2COR|12|13|除了我不曾连累你们这一件事，你们还有什么事不及别的教会呢？这不公平之处，请你们饶恕我吧。
2COR|12|14|如今，我准备第三次到你们那里去。我仍不会连累你们，因为我所求的是你们，不是你们的财物。儿女不该为父母积财，父母该为儿女积财。
2COR|12|15|我也甘心乐意为你们的灵魂费财费力。难道我越爱你们，就越少得你们的爱吗？
2COR|12|16|罢了，我自己并没有连累你们，你们却有人说，我施诡诈，用心计牢笼你们。
2COR|12|17|我所差遣到你们那里去的人，我何曾藉着他们中的任何人占过你们的便宜呢？
2COR|12|18|我劝 提多 到你们那里去，又差遣那位弟兄与他同去， 提多 占过你们的便宜吗？我们的行事为人不是同一心灵 吗？不是同一步伐吗？
2COR|12|19|你们一直认为我们是在你们面前为自己辩护吗？其实，我们本是在基督里当着上帝面前说话。亲爱的，一切的事都是为了造就你们。
2COR|12|20|我怕我再来的时候，见你们不合我所期望的，而你们见我也不合你们所期望的。我怕有纷争、嫉妒、愤怒、自私、毁谤、谗言、狂傲、动乱的事。
2COR|12|21|我怕我再来的时候，我的上帝使我在你们面前蒙羞，并且又因许多人从前犯罪，行污秽、淫乱、放荡的事，不肯悔改而悲伤。
2COR|13|1|这是我第三次要到你们那里去。“任何指控都要凭两个或三个证人的口述才能成立”。
2COR|13|2|对那些犯了罪的人和其余所有的人，正如我第二次见你们的时候曾说过，现在不在你们那里再次说：“我若再来，必不宽容。”
2COR|13|3|因为你们想求证基督是否藉着我说话。基督对你们并不是软弱的，而是在你们里面大有能力的。
2COR|13|4|他因软弱被钉在十字架上，却因上帝的大能仍然活着。我们在他里面也成为软弱的，但对你们，我们将因上帝的大能而与他一同活着。
2COR|13|5|你们总要省察自己是否在信仰中生活；你们要考验自己。除非你们经不起考验，你们自己岂不应该知道有耶稣基督在你们里面吗？
2COR|13|6|我希望你们知道，我们并不是经不起考验的人。
2COR|13|7|我们祈求上帝使你们不做任何恶事；这不是要显明我们是经得起考验的，而是要你们行事端正，即使我们似乎经不起考验也没有关系。
2COR|13|8|我们不能做任何对抗真理的事，只能维护真理。
2COR|13|9|当我们软弱而你们刚强时，我们也欢喜。我们所祈求的是：你们能成为完全人。
2COR|13|10|所以，我不在你们那里的时候，把这些话写给你们，好使我见你们的时候不用照主所给我的权柄严厉地待你们；这权柄原是为造就人，而不是为摧毁人。
2COR|13|11|末了，弟兄们，愿你们喜乐。要追求完全；要接受鼓励；要同心合意；要彼此和睦。如此，慈爱和平的上帝必与你们同在。
2COR|13|12|你们要用圣洁的吻彼此问安。众圣徒都向你们问安。
2COR|13|13|愿主耶稣基督的恩惠、上帝的慈爱、圣灵的感动常与你们众人同在！
