OBAD|1|1|visio Abdiae haec dicit Dominus Deus ad Edom auditum audivimus a Domino et legatum ad gentes misit surgite et consurgamus adversum eum in proelium
OBAD|1|2|ecce parvulum te dedi in gentibus contemptibilis tu es valde
OBAD|1|3|superbia cordis tui extulit te habitantem in scissuris petrae exaltantem solium suum qui dicit in corde suo quis detrahet me in terram
OBAD|1|4|si exaltatus fueris ut aquila et si inter sidera posueris nidum tuum inde detraham te dicit Dominus
OBAD|1|5|si fures introissent ad te si latrones per noctem quomodo conticuisses nonne furati essent sufficientia sibi si vindemiatores introissent ad te numquid saltim racemos reliquissent tibi
OBAD|1|6|quomodo scrutati sunt Esau investigaverunt abscondita eius
OBAD|1|7|usque ad terminum emiserunt te omnes viri foederis tui inluserunt tibi invaluerunt adversum te viri pacis tuae qui comedunt tecum ponent insidias subter te non est prudentia in eo
OBAD|1|8|numquid non in die illa dicit Dominus perdam sapientes de Idumea et prudentiam de monte Esau
OBAD|1|9|et timebunt fortes tui a meridie ut intereat vir de monte Esau
OBAD|1|10|propter interfectionem et propter iniquitatem in fratrem tuum Iacob operiet te confusio et peribis in aeternum
OBAD|1|11|in die cum stares adversus quando capiebant alieni exercitum eius et extranei ingrediebantur portas eius et super Hierusalem mittebant sortem tu quoque eras quasi unus ex eis
OBAD|1|12|et non despicies in die fratris tui in die peregrinationis eius et non laetaberis super filios Iuda in die perditionis eorum et non magnificabis os tuum in die angustiae
OBAD|1|13|neque ingredieris portam populi mei in die ruinae eorum neque despicies et tu in malis eius in die vastitatis illius et non emitteris adversum exercitum eius in die vastitatis illius
OBAD|1|14|neque stabis in exitibus ut interficias eos qui fugerint et non concludes reliquos eius in die tribulationis
OBAD|1|15|quoniam iuxta est dies Domini super omnes gentes sicut fecisti fiet tibi retributionem tuam convertet in caput tuum
OBAD|1|16|quomodo enim bibisti super montem sanctum meum bibent omnes gentes iugiter et bibent et absorbent et erunt quasi non sint
OBAD|1|17|et in monte Sion erit salvatio et erit sanctus et possidebit domus Iacob eos qui se possederant
OBAD|1|18|et erit domus Iacob ignis et domus Ioseph flamma et domus Esau stipula et succendentur in eis et devorabunt eos et non erunt reliquiae domus Esau quia Dominus locutus est
OBAD|1|19|et hereditabunt hii qui ad austrum montem Esau et qui in campestribus Philisthim et possidebunt regionem Ephraim et regionem Samariae et Beniamin possidebit Galaad
OBAD|1|20|et transmigratio exercitus huius filiorum Israhel omnia Chananeorum usque ad Saraptham et transmigratio Hierusalem quae in Bosforo est possidebit civitates austri
OBAD|1|21|et ascendent salvatores in montem Sion iudicare montem Esau et erit Domino regnum
