JOEL|1|1|Слово Господне, которое было к Иоилю, сыну Вафуила.
JOEL|1|2|Слушайте это, старцы, и внимайте, все жители земли сей: бывало ли такое во дни ваши, или во дни отцов ваших?
JOEL|1|3|Передайте об этом детям вашим; а дети ваши пусть скажут своим детям, а их дети следующему роду:
JOEL|1|4|оставшееся от гусеницы ела саранча, оставшееся от саранчи ели черви, а оставшееся от червей доели жуки.
JOEL|1|5|Пробудитесь, пьяницы, и плачьте и рыдайте, все пьющие вино, о виноградном соке, ибо он отнят от уст ваших!
JOEL|1|6|Ибо пришел на землю Мою народ сильный и бесчисленный; зубы у него – зубы львиные, и челюсти у него – как у львицы.
JOEL|1|7|Опустошил он виноградную лозу Мою, и смоковницу Мою обломал, ободрал ее догола, и бросил; сделались белыми ветви ее.
JOEL|1|8|Рыдай, как молодая жена, препоясавшись [вретищем], о муже юности своей!
JOEL|1|9|Прекратилось хлебное приношение и возлияние в доме Господнем; плачут священники, служители Господни.
JOEL|1|10|Опустошено поле, сетует земля; ибо истреблен хлеб, высох виноградный сок, завяла маслина.
JOEL|1|11|Краснейте от стыда, земледельцы, рыдайте, виноградари, о пшенице и ячмене, потому что погибла жатва в поле,
JOEL|1|12|засохла виноградная лоза и смоковница завяла; гранатовое дерево, пальма и яблоня, все дерева в поле посохли; потому и веселье у сынов человеческих исчезло.
JOEL|1|13|Препояшьтесь [вретищем] и плачьте, священники! рыдайте, служители алтаря! войдите, ночуйте во вретищах, служители Бога моего! ибо не стало в доме Бога вашего хлебного приношения и возлияния.
JOEL|1|14|Назначьте пост, объявите торжественное собрание, созовите старцев и всех жителей страны сей в дом Господа Бога вашего, и взывайте к Господу.
JOEL|1|15|О, какой день! ибо день Господень близок; как опустошение от Всемогущего придет он.
JOEL|1|16|Не пред нашими ли глазами отнимается пища, от дома Бога нашего – веселье и радость?
JOEL|1|17|Истлели зерна под глыбами своими, опустели житницы, разрушены кладовые, ибо не стало хлеба.
JOEL|1|18|Как стонет скот! уныло ходят стада волов, ибо нет для них пажити; томятся и стада овец.
JOEL|1|19|К Тебе, Господи, взываю; ибо огонь пожрал злачные пастбища пустыни, и пламя попалило все дерева в поле.
JOEL|1|20|Даже и животные на поле взывают к Тебе, потому что иссохли потоки вод, и огонь истребил пастбища пустыни.
JOEL|2|1|Трубите трубою на Сионе и бейте тревогу на святой горе Моей; да трепещут все жители земли, ибо наступает день Господень, ибо он близок –
JOEL|2|2|день тьмы и мрака, день облачный и туманный: как утренняя заря распространяется по горам народ многочисленный и сильный, какого не бывало от века и после того не будет в роды родов.
JOEL|2|3|Перед ним пожирает огонь, а за ним палит пламя; перед ним земля как сад Едемский, а позади него будет опустошенная степь, и никому не будет спасения от него.
JOEL|2|4|Вид его как вид коней, и скачут они как всадники;
JOEL|2|5|скачут по вершинам гор как бы со стуком колесниц, как бы с треском огненного пламени, пожирающего солому, как сильный народ, выстроенный к битве.
JOEL|2|6|При виде его затрепещут народы, у всех лица побледнеют.
JOEL|2|7|Как борцы бегут они и как храбрые воины влезают на стену, и каждый идет своею дорогою, и не сбивается с путей своих.
JOEL|2|8|Не давят друг друга, каждый идет своею стезею, и падают на копья, но остаются невредимы.
JOEL|2|9|Бегают по городу, поднимаются на стены, влезают на дома, входят в окна, как вор.
JOEL|2|10|Перед ними потрясется земля, поколеблется небо; солнце и луна помрачатся, и звезды потеряют свой свет.
JOEL|2|11|И Господь даст глас Свой пред воинством Своим, ибо весьма многочисленно полчище Его и могуществен исполнитель слова Его; ибо велик день Господень и весьма страшен, и кто выдержит его?
JOEL|2|12|Но и ныне еще говорит Господь: обратитесь ко Мне всем сердцем своим в посте, плаче и рыдании.
JOEL|2|13|Раздирайте сердца ваши, а не одежды ваши, и обратитесь к Господу Богу вашему; ибо Он благ и милосерд, долготерпелив и многомилостив и сожалеет о бедствии.
JOEL|2|14|Кто знает, не сжалится ли Он, и не оставит ли благословения, хлебного приношения и возлияния Господу Богу вашему?
JOEL|2|15|Вострубите трубою на Сионе, назначьте пост и объявите торжественное собрание.
JOEL|2|16|Соберите народ, созовите собрание, пригласите старцев, соберите отроков и грудных младенцев; пусть выйдет жених из чертога своего и невеста из своей горницы.
JOEL|2|17|Между притвором и жертвенником да плачут священники, служители Господни, и говорят: "пощади, Господи, народ Твой, не предай наследия Твоего на поругание, чтобы не издевались над ним народы; для чего будут говорить между народами: где Бог их?"
JOEL|2|18|И тогда возревнует Господь о земле Своей, и пощадит народ Свой.
JOEL|2|19|И ответит Господь, и скажет народу Своему: вот, Я пошлю вам хлеб и вино и елей, и будете насыщаться ими, и более не отдам вас на поругание народам.
JOEL|2|20|И пришедшего от севера удалю от вас, и изгоню в землю безводную и пустую, переднее полчище его – в море восточное, а заднее – в море западное, и пойдет от него зловоние, и поднимется от него смрад, так как он много наделал [зла].
JOEL|2|21|Не бойся, земля: радуйся и веселись, ибо Господь велик, чтобы совершить это.
JOEL|2|22|Не бойтесь, животные, ибо пастбища пустыни произрастят траву, дерево принесет плод свой, смоковница и виноградная лоза окажут свою силу.
JOEL|2|23|И вы, чада Сиона, радуйтесь и веселитесь о Господе Боге вашем; ибо Он даст вам дождь в меру и будет ниспосылать вам дождь, дождь ранний и поздний, как прежде.
JOEL|2|24|И наполнятся гумна хлебом, и переполнятся подточилия виноградным соком и елеем.
JOEL|2|25|И воздам вам за те годы, которые пожирали саранча, черви, жуки и гусеница, великое войско Мое, которое послал Я на вас.
JOEL|2|26|И до сытости будете есть и насыщаться и славить имя Господа Бога вашего, Который дивное соделал с вами, и не посрамится народ Мой во веки.
JOEL|2|27|И узнаете, что Я посреди Израиля, и Я – Господь Бог ваш, и нет другого, и Мой народ не посрамится вовеки.
JOEL|2|28|И будет после того, излию от Духа Моего на всякую плоть, и будут пророчествовать сыны ваши и дочери ваши; старцам вашим будут сниться сны, и юноши ваши будут видеть видения.
JOEL|2|29|И также на рабов и на рабынь в те дни излию от Духа Моего.
JOEL|2|30|И покажу знамения на небе и на земле: кровь и огонь и столпы дыма.
JOEL|2|31|Солнце превратится во тьму и луна – в кровь, прежде нежели наступит день Господень, великий и страшный.
JOEL|2|32|И будет: всякий, кто призовет имя Господне, спасется; ибо на горе Сионе и в Иерусалиме будет спасение, как сказал Господь, и у остальных, которых призовет Господь.
JOEL|3|1|Ибо вот, в те дни и в то самое время, когда Я возвращу плен Иуды и Иерусалима,
JOEL|3|2|Я соберу все народы, и приведу их в долину Иосафата, и там произведу над ними суд за народ Мой и за наследие Мое, Израиля, который они рассеяли между народами, и землю Мою разделили.
JOEL|3|3|И о народе Моем они бросали жребий, и отдавали отрока за блудницу, и продавали отроковицу за вино, и пили.
JOEL|3|4|И что вы Мне, Тир и Сидон и все округи Филистимские? Хотите ли воздать Мне возмездие? хотите ли воздать Мне? Легко и скоро Я обращу возмездие ваше на головы ваши,
JOEL|3|5|потому что вы взяли серебро Мое и золото Мое, и наилучшие драгоценности Мои внесли в капища ваши,
JOEL|3|6|и сынов Иуды и сынов Иерусалима продавали сынам Еллинов, чтобы удалить их от пределов их.
JOEL|3|7|Вот, Я подниму их из того места, куда вы продали их, и обращу мзду вашу на голову вашу.
JOEL|3|8|И предам сыновей ваших и дочерей ваших в руки сынов Иуды, и они продадут их Савеям, народу отдаленному; так Господь сказал.
JOEL|3|9|Провозгласите об этом между народами, приготовьтесь к войне, возбудите храбрых; пусть выступят, поднимутся все ратоборцы.
JOEL|3|10|Перекуйте орала ваши на мечи и серпы ваши на копья; слабый пусть говорит: "я силен".
JOEL|3|11|Спешите и сходитесь, все народы окрестные, и соберитесь; туда, Господи, веди Твоих героев.
JOEL|3|12|Пусть воспрянут народы и низойдут в долину Иосафата; ибо там Я воссяду, чтобы судить все народы отовсюду.
JOEL|3|13|Пустите в дело серпы, ибо жатва созрела; идите, спуститесь, ибо точило полно и подточилия переливаются, потому что злоба их велика.
JOEL|3|14|Толпы, толпы в долине суда! ибо близок день Господень к долине суда!
JOEL|3|15|Солнце и луна померкнут и звезды потеряют блеск свой.
JOEL|3|16|И возгремит Господь с Сиона, и даст глас Свой из Иерусалима; содрогнутся небо и земля; но Господь будет защитою для народа Своего и обороною для сынов Израилевых.
JOEL|3|17|Тогда узнаете, что Я Господь Бог ваш, обитающий на Сионе, на святой горе Моей; и будет Иерусалим святынею, и не будут уже иноплеменники проходить через него.
JOEL|3|18|И будет в тот день: горы будут капать вином и холмы потекут молоком, и все русла Иудейские наполнятся водою, а из дома Господня выйдет источник, и будет напоять долину Ситтим.
JOEL|3|19|Египет сделается пустынею и Едом будет пустою степью – за то, что они притесняли сынов Иудиных и проливали невинную кровь в земле их.
JOEL|3|20|А Иуда будет жить вечно и Иерусалим – в роды родов.
JOEL|3|21|Я смою кровь их, которую не смыл еще, и Господь будет обитать на Сионе.
