MARK|1|1|上帝的儿子 ，耶稣基督福音的起头。
MARK|1|2|正如 以赛亚 先知书上记着： “看哪，我要差遣我的使者在你面前， 他要为你预备道路。
MARK|1|3|在旷野有声音呼喊着： 预备主的道， 修直他的路。”
MARK|1|4|照这话，施洗 约翰 来到旷野 ，宣讲悔改的洗礼，使罪得赦。
MARK|1|5|犹太 全地和全 耶路撒冷 的人都出去，到 约翰 那里，承认他们的罪，在 约旦河 里受他的洗。
MARK|1|6|约翰 穿骆驼毛的衣服，腰束皮带，吃的是蝗虫和野蜜。
MARK|1|7|他宣讲，说：“有一位在我以后来的，能力比我更大，我就是弯腰给他解鞋带也不配。
MARK|1|8|我用水给你们施洗，他却要用圣灵给你们施洗。”
MARK|1|9|那时，耶稣从 加利利 的 拿撒勒 来，在 约旦河 里受了 约翰 的洗。
MARK|1|10|他从水里一上来，就看见天裂开了，圣灵仿佛鸽子降在他身上。
MARK|1|11|又有声音从天上来，说：“你是我的爱子，我喜爱你。”
MARK|1|12|圣灵立刻把耶稣催促到旷野里去。
MARK|1|13|他在旷野四十天，受撒但的试探，并与野兽同在一起，且有天使来伺候他。
MARK|1|14|约翰 下监以后，耶稣来到 加利利 ，宣讲上帝的福音，
MARK|1|15|说：“日期满了，上帝的国近了。你们要悔改，信福音！”
MARK|1|16|耶稣沿着 加利利 的海边走，看见 西门 和 西门 的弟弟 安得烈 在海上撒网；他们本是打鱼的。
MARK|1|17|耶稣对他们说：“来跟从我，我要叫你们得人如得鱼一样。”
MARK|1|18|他们立刻舍了网，跟从他。
MARK|1|19|耶稣稍往前走，又见 西庇太 的儿子 雅各 和他弟弟 约翰 在船上补网。
MARK|1|20|耶稣随即呼召他们，他们就把父亲 西庇太 和雇工留在船上，跟从了耶稣。
MARK|1|21|他们到了 迦百农 ，耶稣就在安息日进了会堂教导人。
MARK|1|22|他们对他的教导感到很惊奇，因为他教导他们正像有权柄的人，不像文士。
MARK|1|23|当时，会堂里有一个污灵附身的人，他在喊叫，
MARK|1|24|说：“ 拿撒勒 人耶稣，你为什么干扰我们？你来消灭我们吗？我知道你是谁，你是上帝的圣者。”
MARK|1|25|耶稣斥责他说：“不要作声，从这人身上出来吧！”
MARK|1|26|污灵使那人抽了一阵风，大声喊叫，就出来了。
MARK|1|27|众人都惊讶，以致彼此对问：“这是什么事？是个新的教导啊！他用权柄命令污灵，连污灵也听从了他。”
MARK|1|28|于是耶稣的名声立刻传遍了全 加利利 周围地区。
MARK|1|29|他们一出会堂，就同 雅各 和 约翰 进了 西门 和 安得烈 的家。
MARK|1|30|西门 的岳母正发烧躺着，就有人告诉耶稣。
MARK|1|31|耶稣进前拉着她的手，扶她起来，烧就退了，于是她服事他们。
MARK|1|32|傍晚日落的时候，有人带着一切害病的和被鬼附的，来到耶稣跟前。
MARK|1|33|全城的人都聚集在门前。
MARK|1|34|耶稣治好了许多害各样病的人，又赶出许多鬼，不许鬼说话，因为鬼认识他。
MARK|1|35|次日早晨，天未亮的时候，耶稣起来，到旷野地方去，在那里祷告。
MARK|1|36|西门 和同伴出去找他，
MARK|1|37|找到了就对他说：“众人都在找你！”
MARK|1|38|耶稣对他们说：“让我们往别处去，到邻近的乡村，我也好在那里传道，因为我是为这事出来的。”
MARK|1|39|于是他走遍全 加利利 ，在他们的会堂传道，并且赶鬼。
MARK|1|40|有一个痲疯病人来求耶稣，向他跪下 ，说：“你若肯，你能使我洁净。”
MARK|1|41|耶稣动了慈心，就伸手摸他，说：“我肯，你洁净了吧！”
MARK|1|42|痲疯病立刻离开他，他就洁净了。
MARK|1|43|耶稣严严地叮嘱他，立刻打发他走，
MARK|1|44|对他说：“你要注意，千万不可告诉任何人，只要去，让祭司为你检查，又因为你已经洁净，献上 摩西 所吩咐的祭物，作为证据给众人看。”
MARK|1|45|那人出去，倒说许多的话，把这件事传扬开了，使耶稣不能再公开进城，只好留在外边旷野地方，人从各处都到他跟前来。
MARK|2|1|过了些日子，耶稣又进了 迦百农 。人听说他在屋里，
MARK|2|2|于是许多人聚集，甚至连门前都没有空地；耶稣就对他们讲道。
MARK|2|3|有人带着一个瘫子来见耶稣，是由四个人抬来的；
MARK|2|4|因为人多，无法抬到耶稣跟前，就把他所在那房子的屋顶拆了，既拆通了，就把瘫子连所躺卧的褥子都缒下去。
MARK|2|5|耶稣见他们的信心，就对瘫子说：“孩子，你的罪赦了。”
MARK|2|6|有几个文士坐在那里，心里议论，说：
MARK|2|7|“这个人为什么这样说呢？他说亵渎的话了。除了上帝一位之外，谁能赦罪呢？”
MARK|2|8|耶稣心中立刻知道他们心里这样议论，就说：“你们心里为什么这样议论呢？
MARK|2|9|对瘫子说‘你的罪赦了’，或说‘起来！拿你的褥子行走’，哪一样容易呢？
MARK|2|10|但要让你们知道，人子在地上有赦罪的权柄。”就对瘫子说：
MARK|2|11|“我吩咐你，起来！拿你的褥子回家去吧。”
MARK|2|12|那人就起来，立刻拿着褥子，当着众人面前出去了，以致众人都惊奇，归荣耀给上帝，说：“我们从来没有见过这样的事！”
MARK|2|13|耶稣又到海边去，众人都到他跟前来，他就教导他们。
MARK|2|14|耶稣往前走，看见 亚勒腓 的儿子 利未 在税关坐着，就对他说：“来跟从我！”他就起来跟从耶稣。
MARK|2|15|耶稣在 利未 家里坐席的时候，有好些税吏和罪人与耶稣和他的门徒一同坐席，因为有很多人也跟随耶稣。
MARK|2|16|法利赛人中的文士 看见耶稣与罪人和税吏一同吃饭，就对他的门徒说：“他与税吏和罪人一同吃饭吗？”
MARK|2|17|耶稣听见，就对他们说：“健康的人用不着医生，有病的人才用得着。我不是来召义人，而是召罪人。”
MARK|2|18|那时， 约翰 的门徒和法利赛人都禁食。他们来问耶稣说：“ 约翰 的门徒和法利赛人的门徒禁食，你的门徒却不禁食，这是为什么呢？”
MARK|2|19|耶稣对他们说：“新郎和宾客在一起的时候，宾客怎么能禁食呢？只要新郎和他们在一起，他们不能禁食。
MARK|2|20|但日子将到，新郎要被带走，那日他们就要禁食了。
MARK|2|21|“没有人把新布缝在旧衣服上，若是这样，所补上的新布会撕破旧衣服，裂口就更大了。
MARK|2|22|也没有人把新酒装在旧皮袋里，若是这样，酒会胀破皮袋，酒和皮袋都糟蹋了 。相反地，新酒要装在新皮袋里 。”
MARK|2|23|有一个安息日，耶稣从麦田经过。他的门徒走路的时候，摘起麦穗来。
MARK|2|24|法利赛人对耶稣说：“看哪！他们为什么做安息日不合法的事呢？”
MARK|2|25|耶稣对他们说：“ 大卫 和跟从他的人饥饿需要食物时所做的事，你们没有念过吗？
MARK|2|26|他在 亚比亚他 作大祭司的时候，怎么进了上帝的居所，吃了供饼，又给跟从他的人吃呢？这饼除了祭司以外，人都不可以吃。”
MARK|2|27|他又对他们说：“安息日是为人设立的，人不是为安息日设立的。
MARK|2|28|所以，人子也是安息日的主。”
MARK|3|1|耶稣又进了会堂，在那里有一个人，他的一只手萎缩了。
MARK|3|2|众人为了要控告耶稣，就窥探他会不会在安息日医治那人。
MARK|3|3|耶稣对那手萎缩了的人说：“起来站在当中！”
MARK|3|4|他又问众人：“在安息日行善行恶，救命害命，哪样是合法的呢？”他们都不作声。
MARK|3|5|耶稣怒目环视他们，因他们的心刚硬而忧伤，就对那人说：“伸出手来！”他把手一伸，手就复原了。
MARK|3|6|法利赛人出去，立刻同 希律 一党的人商议怎样除掉耶稣。
MARK|3|7|耶稣和门徒退到海边去，有许多人从 加利利 跟随他。还有许多人听见他所做的事，就从 犹太 、 耶路撒冷 、 以土买 、 约旦河 的东边，以及 推罗 和 西顿 的附近地方来到他那里。
MARK|3|8|
MARK|3|9|因为人多，他吩咐门徒为他预备一只小船，免得众人拥挤他。
MARK|3|10|他治好了许多人，所以凡有疾病的，都挤着要摸他。
MARK|3|11|每当污灵看见他，就俯伏在他面前，喊着说：“你是上帝的儿子。”
MARK|3|12|耶稣再三嘱咐他们不要把他宣扬出去。
MARK|3|13|耶稣上了山，把自己所要的人召来，他们就来到他那里。
MARK|3|14|于是他设立十二个人，又称他们为使徒 ，要他们常和自己同在，也要差他们去传道，
MARK|3|15|并给他们权柄赶鬼。
MARK|3|16|他设立的十二个人 有 西门 －耶稣又给他起名叫 彼得 ，
MARK|3|17|还有 西庇太 的儿子 雅各 和 雅各 的弟弟 约翰 —耶稣又给他们起名叫 半尼其 ，就是雷的儿子—
MARK|3|18|又有 安得烈 、 腓力 、 巴多罗买 、 马太 、 多马 、 亚勒腓 的儿子 雅各 、 达太 和激进党的 西门 ，
MARK|3|19|还有出卖耶稣的 加略 人 犹大 。
MARK|3|20|耶稣进了屋子，众人又聚集，甚至他连饭也顾不得吃。
MARK|3|21|耶稣的家人听见，就出来要拉住他，因为他们说他癫狂了。
MARK|3|22|从 耶路撒冷 下来的文士说：“他是被 别西卜 附身的”，又说：“他是靠着鬼王赶鬼的。”
MARK|3|23|耶稣叫他们来，用比喻对他们说：“撒但怎能赶出撒但呢？
MARK|3|24|一国若自相纷争，那国就立不住；
MARK|3|25|一家若自相纷争，那家就立不住。
MARK|3|26|撒但若自相攻打纷争，他就立不住，必定灭亡。
MARK|3|27|没有人能进壮士家里，抢夺他的东西；除非先绑住那壮士，否则无法抢夺他的家。
MARK|3|28|我实在告诉你们，世人一切的罪和一切亵渎的话都可以得到赦免；
MARK|3|29|凡亵渎圣灵的，却永不得赦免，而要担当永远的罪。”
MARK|3|30|因为他们说：“他是被污灵附身的。”
MARK|3|31|那时，耶稣的母亲和他兄弟来，站在外边，打发人去叫他。
MARK|3|32|有许多人在耶稣周围坐着，他们就告诉他说：“看哪！你母亲、你兄弟和你姊妹 在外边找你。”
MARK|3|33|耶稣回答他们：“谁是我的母亲？谁是我的兄弟？”
MARK|3|34|就环视那周围坐着的人，说：“看哪，我的母亲，我的兄弟！
MARK|3|35|凡遵行上帝旨意的人就是我的兄弟姊妹和母亲。”
MARK|4|1|耶稣又在海边教导人。有一大群人到他那里聚集，他只好上船坐下。船在海里，众人都靠近海，站在岸上。
MARK|4|2|耶稣就用许多比喻教导他们。在教导的时候，他对他们说：
MARK|4|3|“你们听啊，有一个撒种的出去撒种。
MARK|4|4|他撒的时候，有的落在路旁，飞鸟来把它吃掉了。
MARK|4|5|有的落在土浅的石头地上，因为土不深，很快就长出苗来，
MARK|4|6|太阳出来一晒，因为没有根就枯干了。
MARK|4|7|有的落在荆棘里，荆棘长起来，把它挤住了，就结不出果实。
MARK|4|8|又有的落在好土里，就发芽长大，结出果实，有三十倍的，有六十倍的，有一百倍的。”
MARK|4|9|耶稣又说：“有耳可听的，就应当听！”
MARK|4|10|耶稣独自一人的时候，跟随他的人和十二使徒问他这些比喻的意思。
MARK|4|11|耶稣对他们说：“上帝国的奥秘只让你们知道，若是对外人讲，凡事就用比喻，
MARK|4|12|要 他们看了又看，却看不清， 听了又听，却不明白， 免得他们回转过来，获得赦免。”
MARK|4|13|耶稣又对他们说：“你们不明白这比喻吗？这样怎能明白一切的比喻呢？
MARK|4|14|撒种的人所撒的就是道。
MARK|4|15|那撒在路旁的种子，就是人听了道，撒但立刻来，把撒在他们心里的道夺了去。
MARK|4|16|那撒在石头地上的，就是人听了道，立刻欢喜领受，
MARK|4|17|因心里没有根，不过是暂时的，一旦为道遭受患难或迫害，立刻就跌倒。
MARK|4|18|还有那撒在荆棘里的，就是人听了道，
MARK|4|19|后来有世上的忧虑、钱财的迷惑，和别样的私欲进来，把道挤住了，结不出果实。
MARK|4|20|那撒在好土里的，就是人听了道，领受了，并且结了果实，有三十倍的，有六十倍的，有一百倍的。”
MARK|4|21|耶稣又对他们说：“人拿灯来，难道是要放在斗底下，床底下，而不放在灯台上吗？
MARK|4|22|因为掩藏的事没有不显出来的，隐瞒的事也没有不露出来的。
MARK|4|23|有耳可听的，就应当听！”
MARK|4|24|他又说：“你们要留心所听的。你们用什么量器来量，也将要用什么来量给你们，并且要多给你们。
MARK|4|25|因为有的，还要给他；没有的，连他所有的也要夺去。”
MARK|4|26|耶稣又说：“上帝的国如同人把种子撒在地上，
MARK|4|27|黑夜睡觉，白日起来，这种子就发芽生长，那人却不知道如何会这样。
MARK|4|28|土地自然而然地出产五谷，先发苗，后长穗，然后穗上结成饱满的谷子。
MARK|4|29|五谷熟了，就用镰刀去割，因为收成的时候到了。”
MARK|4|30|耶稣又说：“我们可用什么来比拟上帝的国呢？可用什么比喻来说明呢？
MARK|4|31|它像一粒芥菜种，种在地里的时候，虽比地上所有的种子都小，
MARK|4|32|但种下去以后，它长起来，比各样的菜都大，又长出大枝，以致天上的飞鸟可以在它的荫下筑巢。”
MARK|4|33|耶稣用许多这样的比喻，照他们所能听的，对他们讲道；
MARK|4|34|若不用比喻，他就不对他们讲，但私下没有人的时候，就把一切的道讲给门徒听。
MARK|4|35|那天晚上，耶稣对门徒说：“我们渡到对岸去吧。”
MARK|4|36|门徒离开众人，耶稣已在船上，他们就请他一同去；也有别的船和他同行。
MARK|4|37|忽然狂风大作，波浪打入船内，以致船灌满了水。
MARK|4|38|耶稣在船尾上，枕着枕头睡觉。门徒叫醒他，说：“老师！我们快没命了，你不管吗？”
MARK|4|39|耶稣醒了，斥责那风，向海说：“住了吧！静了吧！”风就止住，大大平静了。
MARK|4|40|耶稣对他们说：“为什么胆怯？你们还没有信心吗？”
MARK|4|41|他们就非常惧怕，彼此说：“这到底是谁？连风和海都听从他。”
MARK|5|1|他们渡到海的对岸，到 格拉森 人 的地区。
MARK|5|2|耶稣一下船，就有一个污灵附身的人从坟墓迎着他走来。
MARK|5|3|那人常住在坟墓里，没有人能捆住他，就是用铁链也不能；
MARK|5|4|因为人屡次用脚镣和铁链捆锁他，铁链被他挣断，脚镣也被他弄碎了，总没有人能制伏他。
MARK|5|5|他昼夜常在坟墓里和山中喊叫，又用石头打自己。
MARK|5|6|他远远看见耶稣，就跑过来拜他，
MARK|5|7|大声呼叫说：“至高上帝的儿子耶稣，你为什么干扰我？我指着上帝恳求你，不要叫我受苦！”
MARK|5|8|这是因耶稣曾吩咐他说：“污灵啊，从这人身上出来！”
MARK|5|9|耶稣问他：“你叫什么名字？”他说：“我名叫 群 ，因为我们数目众多。”
MARK|5|10|他就再三求耶稣不要叫他们离开那地方。
MARK|5|11|在山坡那里，有一大群猪正在吃食；
MARK|5|12|污灵就央求耶稣，说：“求你打发我们进入猪群，好附着它们。”
MARK|5|13|耶稣准了他们，污灵就出来，进入猪里，那群猪就闯下山崖，投进海里，淹死了。猪的数目约有二千。
MARK|5|14|放猪的逃跑了，去告诉城里和乡下的人。众人就来，要看发生了什么事。
MARK|5|15|他们来到耶稣那里，看见那被鬼附的人，就是曾被群鬼所附的，坐着，穿着衣服，神智清醒，他们就害怕。
MARK|5|16|看见这事的人把被鬼附的人所遇见的，和那群猪的事，都告诉了众人，
MARK|5|17|众人就央求耶稣离开他们的地区。
MARK|5|18|耶稣上船的时候，那曾被鬼附的人恳求要和耶稣在一起。
MARK|5|19|耶稣不许，却对他说：“你回家去，到你的亲友那里，将主为你所做多么大的事和他怎样怜悯你，都告诉他们。”
MARK|5|20|那人就走了，开始在 低加坡里 传扬耶稣为他做了多么大的事，众人就都惊讶。
MARK|5|21|耶稣又坐船 渡到对岸，有一大群人聚集到他身边；他正在海边。
MARK|5|22|有一个会堂主管，名叫 叶鲁 ，也来了，一见到耶稣，就俯伏在他脚前，
MARK|5|23|再三求他，说：“我的小女儿快要死了，求你去为她按手，使她痊愈，可以活下去。”
MARK|5|24|耶稣就和他同去。 有一大群人跟随他，拥挤着他。
MARK|5|25|有一个女人，患了经血不止的病有十二年，
MARK|5|26|在好多医生手里受了许多苦，又花尽了她所有的，一点也不见好，反而更重了。
MARK|5|27|她听见耶稣的事，就夹在众人中间，从后面来摸耶稣的衣裳，
MARK|5|28|因她想：“我只摸到他的衣裳，就会痊愈。”
MARK|5|29|于是她的流血立刻止住，她觉得身上的疾病好了。
MARK|5|30|耶稣顿时心里觉得有能力从自己身上出去，就在众人中间转过来，说：“谁摸我的衣裳？”
MARK|5|31|门徒对他说：“你看众人拥挤着你，还说‘谁摸我’呢？”
MARK|5|32|耶稣周围观看，要见做这事的女人。
MARK|5|33|那女人知道在自己身上所成的事，就恐惧战兢，来俯伏在耶稣跟前，将实情全告诉他。
MARK|5|34|耶稣对她说：“女儿，你的信救了你，平安地回去吧！你的疾病痊愈了。”
MARK|5|35|耶稣还在说话的时候，有人从会堂主管的家里来，说：“你的女儿死了，何必还劳驾老师呢？”
MARK|5|36|耶稣不理会他们所说的话，就对会堂主管说：“不要怕，只要信！”
MARK|5|37|于是他带着 彼得 、 雅各 和 雅各 的弟弟 约翰 同去，不许别人跟着他。
MARK|5|38|他们来到会堂主管的家里，耶稣看到一片吵闹，并有人大声哭泣哀号，
MARK|5|39|就进到里面，对他们说：“为什么大吵大哭呢？孩子不是死了，是睡着了。”
MARK|5|40|他们就嘲笑耶稣。耶稣把他们都赶出去，带着孩子的父母和跟随的人进了孩子所在的地方，
MARK|5|41|就拉着孩子的手，对她说：“大利大，古米！”翻出来就是说：“女孩，我吩咐你，起来！”
MARK|5|42|那女孩子立刻起来走动—她已经十二岁了；他们就非常惊奇。
MARK|5|43|耶稣切切地嘱咐他们，不要让人知道这事，又吩咐给她东西吃。
MARK|6|1|耶稣离开那里，来到自己的家乡；门徒也跟从他。
MARK|6|2|到了安息日，他在会堂里教导人。众人听见，就很惊奇，说：“这人哪来这本事呢？所赐给他的是什么智慧？他手所做的是何等的异能呢？
MARK|6|3|这不是那木匠吗？不是 马利亚 的儿子 雅各 、 约西 、 犹大 、 西门 的长兄吗？他姊妹们不也是在我们这里吗？”他们就厌弃他。
MARK|6|4|耶稣对他们说：“先知除了在本乡、本族和自己的家之外，没有不被尊敬的。”
MARK|6|5|耶稣在那里不能行什么异能，不过为几个病人按手，治好他们。
MARK|6|6|他也诧异他们不信。 耶稣走遍周围乡村教导人。
MARK|6|7|他叫了十二个使徒来，差遣他们两个两个地出去，也赐给他们权柄制伏污灵，
MARK|6|8|并且吩咐他们：途中不要带食物和行囊，腰袋里也不要带钱，除了手杖以外，什么都不要带；
MARK|6|9|只要穿鞋子，也不要穿两件内衣。
MARK|6|10|他又对他们说：“你们无论到何处，进哪家，就住在哪里，直到离开那地方。
MARK|6|11|若有什么地方的人不接待你们，不听你们，你们离开那里的时候，要跺掉你们脚上的尘土，证明他们的不是。”
MARK|6|12|使徒就出去传道，叫人悔改，
MARK|6|13|又赶出许多鬼，用油抹了许多病人，治好他们。
MARK|6|14|耶稣的名声传开了， 希律 王也听见。有人说：“施洗的 约翰 从死人中复活了，因此才有这些异能在他里面运行。”
MARK|6|15|但别人说：“他是 以利亚 。”又有人说：“是先知，正如先知中的一位。”
MARK|6|16|希律 听见却说：“是我所斩的 约翰 ，他复活了。”
MARK|6|17|原来， 希律 为他兄弟 腓力 的妻子 希罗底 的缘故，派人去抓了 约翰 ，把他绑了在监狱里，因为 希律 已经娶了那妇人。
MARK|6|18|约翰 曾对 希律 说：“你占有你兄弟的妻子是不合法的。”
MARK|6|19|于是 希罗底 怀恨他，想要杀他，只是不能。
MARK|6|20|因为 希律 怕 约翰 ，知道他是义人，是圣人，所以就保护他，虽然听了他的讲论十分困惑 ，仍然乐意听他。
MARK|6|21|有一天，恰巧是 希律 的生日， 希律 摆设宴席，请了大臣、千夫长和 加利利 的领袖。
MARK|6|22|他的女儿 希罗底 进来跳舞，使 希律 和同席的人都很高兴。王就对女孩说：“无论你要什么，向我求，我都会给你”；
MARK|6|23|又对她多次 起誓说：“无论你向我求什么，就是我国家的一半，我也会给你。”
MARK|6|24|她就出去对她母亲说：“我该求什么呢？”她母亲说：“施洗 约翰 的头。”
MARK|6|25|她就急忙进去见王，求他说：“我愿王立刻把施洗 约翰 的头放在盘子里给我。”
MARK|6|26|王就很忧愁，然而因他所发的誓，又因同席的人，不愿食言，
MARK|6|27|就立刻派一个卫兵，吩咐拿 约翰 的头来。卫兵就去，在监狱里斩了 约翰 ，
MARK|6|28|把头放在盘子里，拿来给那女孩，她就给她母亲。
MARK|6|29|约翰 的门徒听到了，就来把他的尸体领去，放在坟墓里。
MARK|6|30|使徒们聚集到耶稣那里，把一切所做的事、所传的道全告诉他。
MARK|6|31|他就说：“你们来，同我私下到荒野的地方去歇一歇。”这是因为来往的人多，他们连吃饭的时间也没有。
MARK|6|32|他们就坐船，私下往荒野的地方去。
MARK|6|33|众人看见他们走了，有许多认识他们的，就从各城步行，一同跑到那里，比他们先赶到了。
MARK|6|34|耶稣出来，见有一大群的人，就怜悯他们，因为他们如同羊没有牧人一般，于是开始教导他们许多事。
MARK|6|35|天已经很晚，门徒进前来，说：“这地方偏僻，而且天已经很晚了，
MARK|6|36|请叫众人散去，他们好往四面的乡镇村庄去，自己买些东西吃。”
MARK|6|37|耶稣回答他们说：“你们给他们吃吧！”门徒对他说：“我们要拿两百个银币去买饼给他们吃吗？”
MARK|6|38|耶稣说：“你们有多少饼？去看看。”他们知道后就说：“有五个，还有两条鱼。”
MARK|6|39|耶稣吩咐他们，叫众人一组一组地坐在青草地上。
MARK|6|40|众人就一群一群地坐下，有一百的，有五十的。
MARK|6|41|耶稣拿着这五个饼和两条鱼，望着天祝福，擘开饼，递给门徒，摆在众人面前，也把那两条鱼分给众人。
MARK|6|42|他们都吃，并且吃饱了。
MARK|6|43|门徒把饼和鱼的碎屑收拾起来，装满了十二个篮子。
MARK|6|44|吃饼的男人共有五千。
MARK|6|45|耶稣随即催门徒上船，先渡到对岸，到 伯赛大 去，等他叫众人散去。
MARK|6|46|他辞别了他们，就往山上去祷告。
MARK|6|47|到了晚上，船在海中，耶稣独自在岸上。
MARK|6|48|他看见门徒因风不顺，摇橹很苦。天快亮的时候，他在海面上走，往他们那里去，想要超过他们。
MARK|6|49|但门徒看见他在海面上走，以为是鬼怪，就喊叫起来；
MARK|6|50|因为他们都看见了他，甚为惊慌。耶稣连忙对他们说：“放心！是我，不要怕！”
MARK|6|51|于是他到他们那里，一上船，风就停了；他们心里十分惊奇。
MARK|6|52|这是因为他们不明白那分饼的事，心里还是愚顽。
MARK|6|53|他们渡过了海，在 革尼撒勒 靠岸，泊了船，
MARK|6|54|他们一下来，众人立刻认出是耶稣，
MARK|6|55|就跑遍那整个地区，听到他在哪里，就把有病的人用褥子抬到哪里。
MARK|6|56|耶稣所到的地方，或村中、或城里、或乡间，他们都把病人放在街市上，求耶稣让他们摸一摸他的衣裳繸子，摸着的人就都好了。
MARK|7|1|有法利赛人和几个从 耶路撒冷 来的文士聚集到耶稣那里。
MARK|7|2|他们曾看见他的门徒中有人用不洁净的手，就是没有洗的手吃饭。
MARK|7|3|法利赛人和所有的 犹太 人都拘守古人的传统，若不按规矩洗手就不吃饭；
MARK|7|4|从市场来，若不洗净也不吃饭；他们还拘守好些别的规矩，如洗杯、罐、铜器、床铺 等。
MARK|7|5|法利赛人和文士问他说：“你的门徒为什么不照古人的传统，竟然用不洁净的手吃饭呢？”
MARK|7|6|耶稣对他们说：“ 以赛亚 指着你们假冒为善的人所预言的说得好。如经上所记： ‘这百姓用嘴唇尊敬我， 他们的心却远离我。
MARK|7|7|他们把人的规条当作教义教导人； 他们拜我也是枉然。’
MARK|7|8|你们是离弃上帝的诫命，拘守人的传统。”
MARK|7|9|耶稣又说：“你们诚然是废弃上帝的诫命，为要守自己的传统。
MARK|7|10|摩西 说：‘当孝敬父母’；又说：‘咒骂父母的，必须处死。’
MARK|7|11|你们倒说：‘人若对父母说：我所当供奉你的已经作了各耳板’（各耳板就是奉献的意思），
MARK|7|12|你们就容许他不必再奉养父母。
MARK|7|13|这就是你们藉着继承传统，废了上帝的话。你们还做许多这样的事。”
MARK|7|14|耶稣又叫众人来，对他们说：“你们都要听我的话，也要明白。
MARK|7|15|从外面进去的不能玷污人，惟有从里面出来的才玷污人。 ”
MARK|7|16|
MARK|7|17|耶稣离开众人，进了屋子，门徒就问他这比喻的意思。
MARK|7|18|耶稣对他们说：“你们也是这样不明白吗？难道你们不了解，凡从外面进去的不能玷污人吗？
MARK|7|19|因为不是进入他的心，而是进入他的肚子，又排入厕所。”（这是说，各样的食物都是洁净的。）
MARK|7|20|耶稣又说：“从人里面出来的，那才玷污人；
MARK|7|21|因为从人心里发出种种恶念，如淫乱、偷盗、凶杀、
MARK|7|22|奸淫、贪婪、邪恶、诡诈、淫荡、嫉妒、毁谤、骄傲、狂妄。
MARK|7|23|这一切的恶都是从里面出来，且能玷污人。”
MARK|7|24|耶稣从那里起身，往 推罗 境内去，进了一家，他不愿意人知道，却隐藏不住。
MARK|7|25|立刻有一个妇人，她的小女儿被污灵附着，一听见耶稣的事，就来俯伏在他脚前。
MARK|7|26|这妇人是 希腊 人，属 叙利亚 的 腓尼基 族。她求耶稣从她女儿身上赶出那鬼。
MARK|7|27|耶稣对她说：“让孩子们先吃饱，拿孩子的饼丢给小狗吃是不妥的。”
MARK|7|28|妇人回答：“主啊，桌子底下的小狗也吃小孩子的碎屑呀！”
MARK|7|29|耶稣对她说：“凭着这句话，你回去吧，鬼已经离开你的女儿了。”
MARK|7|30|她就回家去，见小孩子躺在床上，鬼已经出去了。
MARK|7|31|耶稣又离开了 推罗 地区，经过 西顿 ，就从 低加坡里 境内来到 加利利海 。
MARK|7|32|有人带着一个耳聋舌结的人来见耶稣，求他为他按手。
MARK|7|33|耶稣领他离开众人，到一边去，就用指头探他的耳朵，吐唾沫抹他的舌头，
MARK|7|34|望天叹息，对他说：“以法大！”就是说“开了吧！”
MARK|7|35|他的耳朵立刻 开了，舌结也解了，他说话也清楚了。
MARK|7|36|耶稣嘱咐他们不要告诉人；但他越嘱咐，他们越发传扬。
MARK|7|37|众人分外惊奇，说：“他所做的事样样都好，他甚至使聋子听见，哑巴说话。”
MARK|8|1|那时，又有一大群人聚集，没有什么吃的。耶稣叫门徒来，说：
MARK|8|2|“我怜悯这群人，因为他们同我在这里已经三天，没有吃的东西了。
MARK|8|3|我若叫他们饿着回家，他们会在路上饿昏，因为其中有从远处来的。”
MARK|8|4|门徒回答：“在这野地，从哪里能得饼使这些人吃饱呢？”
MARK|8|5|耶稣问他们：“你们有多少饼？”他们说：“七个。”
MARK|8|6|他吩咐众人坐在地上，就拿着这七个饼祝谢了，擘开，递给门徒，叫他们摆开，门徒就摆在众人面前。
MARK|8|7|他们还有几条小鱼；耶稣祝谢了，就吩咐也摆在众人面前。
MARK|8|8|他们都吃，并且吃饱了，收拾剩下的碎屑，有七筐子。
MARK|8|9|人数约有四千。耶稣打发他们走了，
MARK|8|10|随即同门徒上船，来到 大玛努他 境内。
MARK|8|11|法利赛人出来盘问耶稣，要求他从天上显个神迹给他们看，想要试探他。
MARK|8|12|耶稣心里深深叹息，说：“这世代为什么求神迹呢？我实在告诉你们，没有神迹给这世代看。”
MARK|8|13|他就离开他们，又上船往海的对岸去了。
MARK|8|14|门徒忘了带饼，在船上除了一个饼，没有别的食物。
MARK|8|15|耶稣嘱咐他们说：“你们要谨慎，要防备法利赛人的酵和 希律 的酵。”
MARK|8|16|他们彼此议论说：“这是因为我们没有饼吧。”
MARK|8|17|耶稣知道了，就说：“你们为什么因为没有饼就议论呢？你们还不领悟，还不明白吗？你们的心还是愚顽吗？
MARK|8|18|你们有眼睛，看不见吗？有耳朵，听不到吗？也不记得吗？
MARK|8|19|我擘开那五个饼分给五千人，你们收拾的碎屑装满了多少个篮子呢？”他们说：“十二个。”
MARK|8|20|“又擘开那七个饼分给四千人，你们收拾的碎屑装满了多少个筐子呢？”他们说：“七个。”
MARK|8|21|耶稣说：“你们还不明白吗？”
MARK|8|22|他们来到 伯赛大 ，有人带一个盲人来，求耶稣摸他。
MARK|8|23|耶稣拉着盲人的手，领他到村外，就吐唾沫在他眼睛上，为他按手，问他：“你看见什么？”
MARK|8|24|他抬头一看，说：“我看见人，他们好像树木，并且行走。”
MARK|8|25|随后耶稣又按手在他眼睛上，他定睛一看，就复原了，样样都看得清楚了。
MARK|8|26|耶稣打发他回家，说：“连这村子你也不要进去。”
MARK|8|27|耶稣和门徒出去，往 凯撒利亚．腓立比 附近的村庄去。在路上，他问门徒：“人们说我是谁？”
MARK|8|28|他们对他说：“是施洗的 约翰 ；有人说是 以利亚 ；又有人说是先知中的一位。”
MARK|8|29|他又问他们：“你们说我是谁？” 彼得 回答他：“你是基督。”
MARK|8|30|于是耶稣切切地嘱咐他们不可对任何人说起他。
MARK|8|31|从此，他教导他们说：“人子必须受许多的苦，被长老、祭司长和文士弃绝，并且被杀，三天后复活。”
MARK|8|32|耶稣明白地说了这话， 彼得 就拉着他，责备他。
MARK|8|33|耶稣转过来看着门徒，斥责 彼得 说：“撒但，退到我后边去！因为你不体会上帝的心意，而是体会人的意思。”
MARK|8|34|于是他叫众人和门徒来，对他们说：“若有人要跟从我，就当舍己，背起自己的十字架来跟从我。
MARK|8|35|因为凡要救自己生命的，必丧失生命；凡为我和福音丧失生命的，必救自己的生命。
MARK|8|36|人就是赚得全世界，赔上自己的生命，有什么益处呢？
MARK|8|37|人还能拿什么换生命呢？
MARK|8|38|凡在这淫乱罪恶的世代，把我和我的道当作可耻的，人子在他父的荣耀里与圣天使一同来临的时候，也要把那人当作可耻的。”
MARK|9|1|耶稣又对他们说：“我实在告诉你们，站在这里的，有人在没经历死亡以前，必定看见上帝的国带着能力临到。”
MARK|9|2|过了六天，耶稣带着 彼得 、 雅各 、 约翰 ，领他们悄悄地上了高山。他在他们面前变了形像，
MARK|9|3|衣服放光，极其洁白，地上漂布的人没有一个能漂得那样白。
MARK|9|4|有 以利亚 和 摩西 向他们显现，并且与耶稣说话。
MARK|9|5|彼得 对耶稣说：“拉比 ，我们在这里真好！我们来搭三座棚，一座为你，一座为 摩西 ，一座为 以利亚 。”
MARK|9|6|彼得 不知道说什么才好，因为他们很害怕。
MARK|9|7|有一朵云彩来遮盖他们，又有声音从云彩里出来，说：“这是我的爱子，你们要听从他！”
MARK|9|8|门徒连忙向周围观看，不再看见任何人，只见耶稣同他们在一起。
MARK|9|9|下山的时候，耶稣嘱咐他们说：“人子还没有从死人中复活，你们不要把所看到的告诉人。”
MARK|9|10|门徒将这话存记在心，彼此议论“从死人中复活”是什么意思。
MARK|9|11|他们就问耶稣：“文士为什么说 以利亚 必须先来？”
MARK|9|12|耶稣说：“ 以利亚 的确先来复兴万事。经上不是指着人子说，他要受许多的苦和被人轻慢吗？
MARK|9|13|我告诉你们， 以利亚 已经来了，他们任意待他，正如经上指着他说的。”
MARK|9|14|他们到了门徒那里，看见有一大群人围着他们，又有文士和他们辩论。
MARK|9|15|众人一见耶稣，都很惊奇，就跑上去向他问安。
MARK|9|16|耶稣问他们：“你们和他们辩论什么？”
MARK|9|17|众人中的一个回答：“老师，我带了我的儿子到你这里来，他被哑巴的灵附着。
MARK|9|18|无论在哪里，那灵拿住他，把他摔倒，他就口吐白沫，牙关紧锁，身体僵硬。我请过你的门徒把那灵赶出去，他们却不能。”
MARK|9|19|耶稣回答：“唉！这不信的世代啊，我和你们在一起要到几时呢？我忍耐你们要到几时呢？把他带到我这里！”
MARK|9|20|他们就带了他来。那灵一见耶稣，就使他重重地抽风，倒在地上，翻来覆去，口吐白沫。
MARK|9|21|耶稣问他父亲：“他得这病有多久了呢？”父亲说：“从小的时候。
MARK|9|22|那灵屡次把他扔在火里、水里，要治死他。你若能做什么，求你怜悯我们，帮助我们。”
MARK|9|23|耶稣对他说：“‘你若能’，在信的人，凡事都能。”
MARK|9|24|孩子的父亲立刻喊着说：“我信；求你帮助我的不信！”
MARK|9|25|耶稣看见众人都跑上来，就斥责那污灵说：“你这聋哑的灵，我命令你从他里头出来，再不要进去！”
MARK|9|26|那灵大喊一声，使孩子猛烈地抽了一阵风，就出来了。孩子好像死了一般，以致众人多半说：“他死了。”
MARK|9|27|但耶稣拉着他的手，扶他起来，他就站起来了。
MARK|9|28|耶稣进了屋子，门徒就私下问他：“我们为什么不能赶出那灵呢？”
MARK|9|29|耶稣对他们说：“非用祷告 ，这一类的邪灵总赶不出来。”
MARK|9|30|他们离开那地方，经过 加利利 ；耶稣不愿意人知道，
MARK|9|31|因为他正教导门徒说：“人子将要被交在人手里，他们要杀害他；被杀以后，三天后他要复活。”
MARK|9|32|门徒却不明白这话，又不敢问他。
MARK|9|33|他们来到 迦百农 。耶稣在屋里问门徒说：“你们在路上议论的是什么？”
MARK|9|34|门徒不作声，因为他们在路上彼此争论谁最大。
MARK|9|35|耶稣坐下，叫十二个使徒来，说：“若有人愿意为首，他要作众人之后，作众人的用人。”
MARK|9|36|于是耶稣领一个小孩过来，让他站在门徒当中，又抱起他来，对他们说：
MARK|9|37|“凡为我的名接纳一个像这小孩子的，就是接纳我；凡接纳我的，不是接纳我，而是接纳那差我来的。”
MARK|9|38|约翰 对耶稣说：“老师，我们看见一个人奉你的名赶鬼，我们就阻止他，因为他不跟从我们。”
MARK|9|39|耶稣说：“不要阻止他，因为没有人奉我的名行异能，反倒轻易毁谤我。
MARK|9|40|不抵挡我们的，就是帮助我们的。
MARK|9|41|凡因你们是属基督，给你们一杯水喝的，我实在告诉你们，他一定会得到赏赐。”
MARK|9|42|“凡使这些信我的小子 中的一个跌倒的，倒不如把大磨石拴在这人的颈项上，扔在海里。
MARK|9|43|如果你一只手使你跌倒，就把它砍下来；你缺一只手进入永生，比有两只手落到地狱，入那不灭的火里去还好。
MARK|9|44|
MARK|9|45|如果你一只脚使你跌倒，就把它砍下来；你瘸腿进入永生，比有两只脚被扔进地狱里还好。
MARK|9|46|
MARK|9|47|如果你一只眼使你跌倒，就去掉它；你只有一只眼进入上帝的国，比有两只眼被扔进地狱里还好。
MARK|9|48|在那里，虫是不死的，火是不灭的。
MARK|9|49|因为每个人必被火像盐一般腌起来。
MARK|9|50|盐本是好的，若失了咸味，你们怎能用它调味呢？你们中间要有盐，彼此和睦。”
MARK|10|1|耶稣从那里起身，来到 犹太 的境内， 约旦河 的东边。众人又聚集到他那里，他又照常教导他们。
MARK|10|2|有法利赛人来问他说：“男人休妻合不合法？”意思是要试探他。
MARK|10|3|耶稣回答他们说：“ 摩西 吩咐你们的是什么？”
MARK|10|4|他们说：“ 摩西 准许写了休书就可以休妻。”
MARK|10|5|耶稣对他们说：“ 摩西 因为你们的心硬，所以写这诫命给你们。
MARK|10|6|但从起初创造的时候，上帝造人是造男造女。
MARK|10|7|因此，人要离开他的父母，与妻子结合 ，
MARK|10|8|二人成为一体。既然如此，夫妻不再是两个人，而是一体的了。
MARK|10|9|所以，上帝配合的，人不可分开。”
MARK|10|10|他们到了屋里，门徒又问他这事。
MARK|10|11|耶稣对他们说：“凡休妻另娶的，就是犯奸淫，辜负他的妻子；
MARK|10|12|妻子若离弃丈夫另嫁，也是犯奸淫了。”
MARK|10|13|有人带着小孩子来见耶稣，要他摸他们，门徒就责备那些人。
MARK|10|14|耶稣看见就很生气，对门徒说：“让小孩到我这里来，不要阻止他们，因为在上帝国的正是这样的人。
MARK|10|15|我实在告诉你们，凡要接受上帝国的，若不像小孩子，绝不能进去。”
MARK|10|16|于是他抱着小孩子，给他们按手，为他们祝福。
MARK|10|17|耶稣刚上路的时候，有一个人跑来，跪在他面前，问他：“善良的老师，我该做什么事才能承受永生？”
MARK|10|18|耶稣对他说：“你为什么称我是善良的？除了上帝一位之外，再没有善良的。
MARK|10|19|诫命你是知道的：‘不可杀人；不可奸淫；不可偷盗；不可作假见证；不可亏负人；当孝敬父母。’”
MARK|10|20|他对耶稣说：“老师，这一切我从小都遵守了。”
MARK|10|21|耶稣看着他，就爱他，对他说：“你还缺少一件：去变卖你所有的，分给穷人，就必有财宝在天上；然后来跟从我。”
MARK|10|22|他听见这话，脸就变了色，忧忧愁愁地走了，因为他的产业很多。
MARK|10|23|耶稣看了看周围，对门徒说：“有钱财的人进上帝的国是何等的难哪！”
MARK|10|24|门徒对他的话非常惊奇。耶稣又对他们说：“孩子们， 要进上帝的国是何等的难哪！
MARK|10|25|骆驼穿过针眼比财主进上帝的国还容易呢！”
MARK|10|26|门徒就更为惊讶，彼此对问：“这样，谁能得救呢？”
MARK|10|27|耶稣看着他们，说：“在人不能，在上帝却不然，因为在上帝凡事都能。”
MARK|10|28|彼得 就对他说：“看哪，我们已经撇下一切跟从你了。”
MARK|10|29|耶稣说：“我实在告诉你们，凡为我和福音撇下房屋，或是兄弟、姊妹、父亲、母亲、儿女、田地，
MARK|10|30|没有不在今世得百倍的，就是房屋、兄弟、姊妹、母亲、儿女、田地，并且要受迫害，在来世得永生。
MARK|10|31|然而，有许多在前的，将要在后；在后的，将要在前。”
MARK|10|32|他们行路上 耶路撒冷 去。耶稣在前头走，他们很惊讶，跟从的人也害怕。耶稣又叫十二使徒来，把自己将要遭遇的事告诉他们，
MARK|10|33|说：“看哪，我们上 耶路撒冷 去，人子将被交给祭司长和文士；他们要定他死罪，又交给外邦人。
MARK|10|34|他们要戏弄他，向他吐唾沫，鞭打他，杀害他；三天后，他要复活。”
MARK|10|35|西庇太 的儿子 雅各 和 约翰 进前来，对耶稣说：“老师，我们无论求你什么，愿你为我们做。”
MARK|10|36|耶稣对他们说：“要我为你们做什么？”
MARK|10|37|他们对他说：“在你的荣耀里，请赐我们一个坐在你右边，一个坐在你左边。”
MARK|10|38|耶稣对他们说：“你们不知道所求的是什么。我所喝的杯，你们能喝吗？我所受的洗，你们能受吗？”
MARK|10|39|他们对他说：“我们能。”耶稣对他们说：“我所喝的杯，你们要喝；我所受的洗，你们也要受。
MARK|10|40|可是坐在我的左右，不是我可以赐的，而是为谁预备就赐给谁。”
MARK|10|41|其余十个门徒听见，就对 雅各 和 约翰 很生气。
MARK|10|42|耶稣叫了他们来，对他们说：“你们知道，外邦人有君王作主治理他们，有大臣操权管辖他们。
MARK|10|43|但是在你们中间，不可这样。你们中间谁愿为大，就要作你们的用人；
MARK|10|44|在你们中间谁愿为首，就要作众人的仆人。
MARK|10|45|因为人子来，并不是要受人的服事，乃是要服事人，并且要舍命作多人的赎价。”
MARK|10|46|他们到了 耶利哥 。耶稣同门徒并许多人离开 耶利哥 的时候，有一个讨饭的盲人，是 底买 的儿子 巴底买 ，坐在路旁。
MARK|10|47|他听见是 拿撒勒 的耶稣，就喊了起来，说：“ 大卫 之子耶稣啊，可怜我吧！”
MARK|10|48|有许多人责备他，不许他作声，他却越发喊着：“ 大卫 之子啊，可怜我吧！”
MARK|10|49|耶稣就站住，说：“叫他过来。”他们就叫那盲人，对他说：“放心，起来！他在叫你啦。”
MARK|10|50|盲人就丢下衣服，跳起来，走到耶稣那里。
MARK|10|51|耶稣回答他说：“你要我为你做什么？”盲人对他说：“拉波尼 ，我要能看见。”
MARK|10|52|耶稣对他说：“你去吧！你的信救了你。”盲人立刻看得见，就在路上跟随耶稣。
MARK|11|1|耶稣和门徒快到 耶路撒冷 ，来到 伯法其 和 伯大尼 ，在 橄榄山 那里。耶稣打发两个门徒，
MARK|11|2|对他们说：“你们往对面村子里去，一进去的时候会看见一匹驴驹拴在那里，是从来没有人骑过的，把它解开，牵来。
MARK|11|3|若有人对你们说：‘为什么做这事？’你们就说：‘主要用它，但会立刻把它牵回到这里来。’”
MARK|11|4|他们去了，看见一匹驴驹拴在门外街道上，就把它解开。
MARK|11|5|在那里站着的人，有几个说：“你们解开驴驹做什么？”
MARK|11|6|门徒照着耶稣的话说，那些人就任凭他们牵去了。
MARK|11|7|他们把驴驹牵到耶稣那里，把自己的衣服搭在上面，耶稣就骑上。
MARK|11|8|有许多人把衣服铺在路上，还有人把田间的树枝砍下来铺上。
MARK|11|9|前呼后拥的人都喊着说： “和散那 ！ 奉主名来的是应当称颂的！
MARK|11|10|那将要来的我祖 大卫 之国是应当称颂的！ 至高无上的，和散那！”
MARK|11|11|耶稣到了 耶路撒冷 ，进入圣殿，看了周围的一切。天色已晚，他就和十二使徒出城，往 伯大尼 去。
MARK|11|12|第二天，他们从 伯大尼 出来，耶稣饿了。
MARK|11|13|他远远地看见一棵无花果树，树上有叶子，就过去，看是不是在树上可以找到什么。他到了树下，竟找不到什么，只有叶子，因为不是无花果的季节。
MARK|11|14|耶稣就对树说：“从今以后，永没有人吃你的果子。”他的门徒都听到了。
MARK|11|15|他们来到 耶路撒冷 。耶稣一进圣殿，就赶出在圣殿里做买卖的人，推倒兑换银钱之人的桌子和卖鸽子之人的凳子；
MARK|11|16|也不许人拿着器具从圣殿里经过。
MARK|11|17|他教导他们说：“经上不是记着： ‘我的殿要称为万国祷告的殿吗？ 你们倒使它成为贼窝了。’”
MARK|11|18|祭司长和文士听见这话，就想法子要除掉耶稣，却又怕他，因为众人都对他的教导感到惊奇。
MARK|11|19|每天晚上，他们 都到城外去。
MARK|11|20|早晨，他们从那里经过，看见无花果树连根都枯干了。
MARK|11|21|彼得 想起耶稣的话来，就对他说：“拉比，你看！你所诅咒的无花果树已经枯干了。”
MARK|11|22|耶稣回答：“你们对上帝要有信心。
MARK|11|23|我实在告诉你们，无论何人对这座山说：‘离开此地，投在海里！’他心里若不疑惑，只信所说的必成，就为他实现。
MARK|11|24|所以我告诉你们，凡你们祷告祈求的，无论是什么，只要信你们已经得着了，就为你们实现。
MARK|11|25|你们站着祷告的时候，若想起有人得罪你们，就该饶恕他，好让你们在天上的父也饶恕你们的过犯。 ”
MARK|11|26|
MARK|11|27|他们又来到 耶路撒冷 。耶稣在圣殿里行走的时候，祭司长、文士和长老进前来，
MARK|11|28|问他说：“你仗着什么权柄做这些事？给你权柄做这些事的是谁呢？”
MARK|11|29|耶稣对他们说：“我要问你们一句话，你们回答我，我就告诉你们我仗着什么权柄做这些事。
MARK|11|30|约翰 的洗礼是从天上来的，还是从人间来的呢？你们回答我吧。”
MARK|11|31|他们彼此商议说：“我们若说‘从天上来的’，他会说：‘这样，你们为什么不信他呢？’
MARK|11|32|但若说‘从人间来的’，却又怕众人，因为大家认为 约翰 确是先知。”
MARK|11|33|于是他们回答耶稣：“我们不知道。”耶稣说：“我也不告诉你们，我仗着什么权柄做这些事。”
MARK|12|1|耶稣就用比喻对他们说：“有人开垦了一个葡萄园，四周围上篱笆，挖了一个榨酒池，盖了一座守望楼，租给园户，就出外远行去了。
MARK|12|2|到了时候，他打发一个仆人到园户那里，要向他们收葡萄园的果子。
MARK|12|3|他们拿住他，打了他，叫他空手回去。
MARK|12|4|园主再打发一个仆人到他们那里。他们打伤他的头，并且侮辱他。
MARK|12|5|园主又打发一个仆人去，他们就杀了他。以后又打发好些仆人去，有的被他们打了，有的被他们杀了。
MARK|12|6|园主还有一位，是他的爱子，最后又打发他去，说：‘他们会尊敬我的儿子。’
MARK|12|7|那些园户却彼此说：‘这是承受产业的。来，我们杀了他，产业就归我们了！’
MARK|12|8|于是他们拿住他，杀了他，把他扔出葡萄园。
MARK|12|9|这样，葡萄园主要怎么做呢？他要来除灭那些园户，将葡萄园转给别人。
MARK|12|10|‘匠人所丢弃的石头 已作了房角的头块石头。 这是主所做的， 在我们眼中看为奇妙。’ 这经文你们没有念过吗？”
MARK|12|11|
MARK|12|12|他们看出这比喻是指着他们说的，就想要捉拿他，但是惧怕众人，于是离开他走了。
MARK|12|13|后来，他们打发几个法利赛人和 希律 党人到耶稣那里，要用他自己的话陷害他。
MARK|12|14|他们来了，就对他说：“老师，我们知道你是诚实的，无论谁你都一视同仁；因为你不看人的面子，而是诚诚实实传上帝的道。纳税给凯撒合不合法？
MARK|12|15|我们该不该纳？”耶稣知道他们的虚伪，就对他们说：“你们为什么试探我？拿一个银币来给我看。”
MARK|12|16|他们就拿了来。耶稣问他们：“这像和这名号是谁的？”他们对他说：“是凯撒的。”
MARK|12|17|耶稣对他们说：“凯撒的归凯撒；上帝的归上帝。”他们对他非常惊讶。
MARK|12|18|撒都该人来见耶稣。他们说没有复活这回事，于是问耶稣：
MARK|12|19|“老师， 摩西 为我们写下这话：‘某人的哥哥若死了，撇下妻子，没有孩子，他该娶哥哥的妻子，为哥哥生子立后。’
MARK|12|20|那么，有兄弟七人，第一个娶了妻，死了，没有留下孩子。
MARK|12|21|第二个娶了她，也死了，没有留下孩子。第三个也是这样。
MARK|12|22|那七个人都没有留下孩子。最后，那妇人也死了。
MARK|12|23|在复活的时候， 她是哪一个的妻子呢？因为他们七个人都娶过她。”
MARK|12|24|耶稣说：“你们错了，不正是因为不明白圣经，也不知道上帝的大能吗？
MARK|12|25|当人从死人中复活后，也不娶也不嫁，而是像天上的天使一样。
MARK|12|26|论到死人复活，你们没有念过 摩西 书中《荆棘篇》上所记载的吗？上帝对 摩西 说：‘我是 亚伯拉罕 的上帝， 以撒 的上帝， 雅各 的上帝。’
MARK|12|27|上帝不是死人的上帝，而是活人的上帝。你们是大错了。”
MARK|12|28|有一个文士来，听见他们的辩论，知道耶稣回答得好，就问他说：“诫命中哪一条是第一呢？”
MARK|12|29|耶稣回答：“第一是：‘ 以色列 啊，你要听，主—我们的上帝是独一的主。
MARK|12|30|你要尽心、尽性、尽意、尽力爱主—你的上帝。’
MARK|12|31|第二是：‘要爱邻 如己。’再没有比这两条诫命更大的了。”
MARK|12|32|那文士对耶稣说：“好，老师，你说得对，上帝是一位，除了他以外，再没有别的了；
MARK|12|33|并且尽心、尽智、尽力爱他，又爱邻如己，要比一切燔祭和祭祀好得多。”
MARK|12|34|耶稣见他回答得有智慧，就对他说：“你离上帝的国不远了。”从此以后，没有人敢再问他什么。
MARK|12|35|耶稣在圣殿里教导人，问他们说：“文士怎么说基督是 大卫 的后裔呢？
MARK|12|36|大卫 被圣灵感动，说： ‘主对我主说： 你坐在我的右边， 等我把你的仇敌放在你脚下 。’
MARK|12|37|大卫 亲自称他为主，他怎么又是 大卫 的后裔呢？”一大群的人都喜欢听他。
MARK|12|38|他在教导的时候，说：“你们要防备文士。他们好穿长袍走来走去，喜欢人们在街市上向他们问安，
MARK|12|39|又喜爱会堂里的高位，宴席上的首座。
MARK|12|40|他们侵吞寡妇的家产，假意作很长的祷告。这些人要受更重的惩罚！”
MARK|12|41|耶稣面向圣殿银库坐着，看众人怎样把钱投入银库。有好些财主投了许多钱。
MARK|12|42|有一个穷寡妇来，投了两个小文钱 ，就是一个大文钱 。
MARK|12|43|耶稣叫门徒来，对他们说：“我实在告诉你们，这穷寡妇投入银库里的比众人所投的更多。
MARK|12|44|因为，众人都是拿有余的捐献，但这寡妇，虽然自己不足，却把她一生所有的全都投进去了。”
MARK|13|1|耶稣从圣殿里出来的时候，有一个门徒对他说：“老师，请看，这是多么了不起的石头！多么了不起的建筑！”
MARK|13|2|耶稣对他说：“你看见这些宏伟的建筑吗？这里将没有一块石头会留在另一块石头上而不被拆毁的。”
MARK|13|3|耶稣在 橄榄山 上，面向圣殿坐着； 彼得 、 雅各 、 约翰 和 安得烈 私下问他说：
MARK|13|4|“请告诉我们，什么时候有这些事呢？这一切事将成的时候有什么预兆呢？”
MARK|13|5|耶稣说：“你们要谨慎，免得有人迷惑你们。
MARK|13|6|将有好些人冒我的名来，说‘我是基督’，并且要迷惑许多人。
MARK|13|7|当你们听见打仗和打仗的风声，不要惊慌；这些事必须发生，但这还不是终结。
MARK|13|8|民要攻打民，国要攻打国，多处必有地震、饥荒。这都是灾难 的起头。
MARK|13|9|但你们自己要谨慎；因为有人要把你们交给议会，并且你们在会堂里要受鞭打，又为我的缘故站在统治者和君王面前，对他们作见证。
MARK|13|10|然而，福音必须先传给万民。
MARK|13|11|有人把你们解送去受审的时候，不要事先担心说什么；到那时候，赐给你们什么话，你们就说什么；因为说话的不是你们，而是圣灵。
MARK|13|12|兄弟要把兄弟、父亲要把儿女置于死地；儿女要起来与父母为敌，害死他们；
MARK|13|13|而且你们要为我的名被众人憎恨。但坚忍到底的终必得救。”
MARK|13|14|“当你们看见那‘施行毁灭的亵渎者’站在不当站的地方（读这经的人要会意），那时，在 犹太 的，应当逃到山上；
MARK|13|15|在屋顶上的，不要下来，也不要进家里去拿东西；
MARK|13|16|在田里的，不要回去取衣裳。
MARK|13|17|在那些日子，怀孕的和奶孩子的就苦了。
MARK|13|18|你们要祈求，叫这事不在冬天发生。
MARK|13|19|因为，在那些日子必有灾难，自从上帝创造万物直到如今，从没有这样的灾难，将来也不会有。
MARK|13|20|若不是主减少那些日子，凡血肉之躯的，就没有一个能得救；但是为了他所拣选的选民，他将那些日子减少了。
MARK|13|21|那时，若有人对你们说：‘看哪，基督在这里！看哪，在那里！’你们不要信。
MARK|13|22|因为假基督和假先知将要起来，显神迹奇事，如果可能，连选民也迷惑了。
MARK|13|23|你们要谨慎！凡事我都预先告诉你们了。”
MARK|13|24|“在那些日子、那灾难以后， 太阳要变黑，月亮也不放光，
MARK|13|25|众星要从天上坠落， 天上的万象都要震动。
MARK|13|26|那时，他们要看见人子带着大能力和荣耀驾云来临。
MARK|13|27|他要差遣天使，从四方，从地极直到天边，召集他的选民。”
MARK|13|28|“你们要从无花果树学习功课：当树枝发芽长叶的时候，你们就知道夏天近了。
MARK|13|29|同样，当你们看见这些事发生，就知道那时候近了，就在门口了。
MARK|13|30|我实在告诉你们，这世代还没有过去，这一切都要发生。
MARK|13|31|天地要废去，我的话却绝不废去。”
MARK|13|32|“但那日子，那时辰，没有人知道，连天上的天使也不知道，子也不知道，惟有父知道。
MARK|13|33|你们要谨慎，要警醒 ，因为你们不知道那时刻几时来到。
MARK|13|34|这事正如一个人离家远行，授权给仆人们，分派各人的工作，又吩咐看门的警醒。
MARK|13|35|所以，你们要警醒，因为你们不知道这家的主人什么时候来，是晚上，或半夜，或鸡叫时，或早晨，
MARK|13|36|免得他忽然来到，看见你们睡着了。
MARK|13|37|我对你们所说的话，也是对众人说的：要警醒！”
MARK|14|1|过两天是逾越节，又是除酵节，祭司长和文士在想法子怎样设计捉拿耶稣，把他杀掉。
MARK|14|2|他们说：“不可在过节的日子，恐怕百姓生乱。”
MARK|14|3|耶稣在 伯大尼 痲疯病人 西门 家里坐席的时候，有一个女人拿着一玉瓶极贵的纯哪哒 香膏来，打破玉瓶，把膏浇在耶稣的头上。
MARK|14|4|有几个人心中很不高兴，说：“何必这样浪费香膏呢？
MARK|14|5|这香膏可以卖三百多个银币周济穷人。”他们就对那女人生气。
MARK|14|6|耶稣说：“由她吧！为什么难为她呢？她在我身上做的是一件美事。
MARK|14|7|因为常有穷人和你们在一起，要向他们行善，随时都可以，但是你们不常有我。
MARK|14|8|她所做的是尽她所能的；她是为了我的安葬，把香膏预先浇在我身上。
MARK|14|9|我实在告诉你们，普天之下，无论在什么地方传这福音，都要述说这女人所做的，来记念她。”
MARK|14|10|十二使徒中有一个 加略 人 犹大 ，去见祭司长，要把耶稣交给他们。
MARK|14|11|他们听见就很高兴，又应许给他银子；他就想怎样找机会把耶稣交给他们。
MARK|14|12|除酵节的第一天，就是宰逾越节羔羊的那一天，门徒对耶稣说：“你要我们到哪里去预备你吃逾越节的宴席呢？”
MARK|14|13|耶稣就打发两个门徒，对他们说：“你们进城去，会有人拿着一罐水迎面而来，你们就跟着他。
MARK|14|14|无论他进哪一家，你们就对那家的主人说：‘老师问：我的客房在哪里？我和我的门徒要在那里吃逾越节的宴席。’
MARK|14|15|他会带你们看一间摆设齐全、准备妥当的楼上大厅，你们就在那里为我们预备。”
MARK|14|16|门徒出去，进了城，所看到的正如耶稣所说的。他们就预备了逾越节的宴席。
MARK|14|17|到了晚上，耶稣和十二使徒都来了。
MARK|14|18|他们坐席，正吃的时候，耶稣说：“我实在告诉你们，你们中间有一个与我同吃的人要出卖我了。”
MARK|14|19|他们就忧愁起来，一个个地问他：“不是我吧？”
MARK|14|20|耶稣对他们说：“是十二人中的一个，就是同我蘸饼在盘子里的那个人。
MARK|14|21|人子要去了，正如经上所写有关他的；但出卖人子的人有祸了！那人没有出生倒好。”
MARK|14|22|他们吃的时候，耶稣拿起饼来，祝福了，就擘开，递给他们，说：“你们拿去，这是我的身体。”
MARK|14|23|他又拿起杯来，祝谢了，递给他们；他们都喝了。
MARK|14|24|耶稣对他们说：“这是我立约的血，为许多人流出来的。
MARK|14|25|我实在告诉你们，我不再喝这葡萄汁，直到我在上帝的国里喝新的那日子。”
MARK|14|26|他们唱了诗，就出来往 橄榄山 去。
MARK|14|27|耶稣对他们说：“你们都要跌倒，因为经上记着： ‘我要击打牧人， 羊就分散了。’，　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　
MARK|14|28|但我复活以后，要在你们之前往 加利利 去。”
MARK|14|29|彼得 说：“虽然众人跌倒，但我不会。”
MARK|14|30|耶稣对他说：“我实在告诉你，今天夜里，鸡叫两遍 以前，你要三次不认我。”
MARK|14|31|彼得 却极力地说：“我就是必须和你同死，也绝不会不认你。”所有的门徒 都是这样说。
MARK|14|32|他们来到一个地方，名叫 客西马尼 。耶稣对门徒说：“你们坐在这里，我去祷告。”
MARK|14|33|于是他带着 彼得 、 雅各 和 约翰 同去。他惊恐起来，极其难过，
MARK|14|34|对他们说：“我心里非常忧伤，几乎要死；你们留在这里，要警醒。”
MARK|14|35|他就稍往前走，俯伏在地，祷告说，如果可能，就叫那时候离开他。
MARK|14|36|他说：“阿爸，父啊！在你凡事都能；求你将这杯撤去。然而，不是照我所愿的，而是照你所愿的。”
MARK|14|37|耶稣回来，见他们睡着了，就对 彼得 说：“ 西门 ，你睡着了吗？不能警醒一小时吗？
MARK|14|38|总要警醒祷告，免得陷入试探。你们心灵固然愿意，肉体却软弱了。”
MARK|14|39|耶稣又去祷告，说的话跟先前一样。
MARK|14|40|他又来，见他们睡着了，因为他们的眼睛很困倦；他们也不知道怎么回答他。
MARK|14|41|他第三次来对他们说：“现在你们仍在睡觉安歇吗？够了，时候到了。看哪，人子被出卖在罪人手里了。
MARK|14|42|起来，我们走吧！看哪，那出卖我的人快来了。”
MARK|14|43|耶稣还在说话的时候，忽然十二使徒之一的 犹大 来了，还有一群人带着刀棒，从祭司长、文士和长老那里跟他同来。
MARK|14|44|那出卖耶稣的人曾给他们一个暗号，说：“我亲谁，谁就是。你们把他抓住，稳妥地带走。”
MARK|14|45|犹大 来了，随即到耶稣跟前，说：“拉比”，就跟他亲吻。
MARK|14|46|他们就下手抓住他。
MARK|14|47|旁边站着的人，有一个拔出刀来，把大祭司的仆人砍了一刀，削掉了他一只耳朵。
MARK|14|48|耶稣回应他们说：“你们带着刀棒出来拿我，如同拿强盗吗？
MARK|14|49|我天天教导人，同你们在殿里，你们并没有抓我。但这是要应验经上的话。”
MARK|14|50|门徒都离开他，逃走了。
MARK|14|51|有一个青年光着身子，只披一块麻布，跟随耶稣，众人就抓住他。
MARK|14|52|他却丢下麻布，赤身逃走了。
MARK|14|53|他们把耶稣带到大祭司那里，又有众祭司长、长老和文士都来一同聚集。
MARK|14|54|彼得 远远地跟着耶稣，直到进了大祭司的院子，和警卫一同坐在火边取暖。
MARK|14|55|祭司长和全议会寻找见证控告耶稣，要处死他，却找不到实据。
MARK|14|56|因为有好些人作假见证告他，他们的见证又各不相符。
MARK|14|57|又有几个人站起来，作假见证告他说：
MARK|14|58|“我们听见他说：‘我要拆毁这人手所造的殿，三日内另造一座不是人手所造的。’”
MARK|14|59|就是这样，他们的见证还是不相符。
MARK|14|60|大祭司起来站在中间，问耶稣说：“这些人作证告你的事，你什么都不回答吗？”
MARK|14|61|耶稣却不言语，一句也不回答。大祭司又问他：“你是不是基督，那当称颂者的儿子？”
MARK|14|62|耶稣说：“我是。 你们要看见人子 坐在那权能者的右边， 驾着天上的云来临。”
MARK|14|63|大祭司就撕裂衣服，说：“我们何必再要证人呢？
MARK|14|64|你们已经听见他这亵渎的话了。你们的决定如何？”他们都判定他该处死。
MARK|14|65|于是有人开始向他吐唾沫，又蒙着他的脸，用拳头打他，对他说：“你说预言吧！”警卫把他拉过来，打他耳光。
MARK|14|66|彼得 在下边院子里，大祭司的一个使女来了，
MARK|14|67|见 彼得 取暖，就看着他，说：“你素来也是同 拿撒勒 人耶稣一起的。”
MARK|14|68|彼得 却不承认，说：“我不知道，也不明白你说的是什么！”于是他出来，到了前院，鸡就叫了 。
MARK|14|69|那使女看见他，又对旁边站着的人说：“这个人也是他们一伙的。”
MARK|14|70|彼得 又不承认。过了不久，旁边站着的人又对 彼得 说：“你真是他们一伙的，因为你也是 加利利 人。”
MARK|14|71|彼得 就赌咒发誓说：“我不认得你们说的这个人。”
MARK|14|72|立刻，鸡叫了第二遍。 彼得 想起耶稣对他所说的话：“鸡叫两遍以前，你要三次不认我。”他就忍不住哭了。
MARK|15|1|一到早晨，众祭司长、长老、文士，和全议会的人大家商议，就把耶稣绑着，解去，交给 彼拉多 。
MARK|15|2|彼拉多 问他：“你是 犹太 人的王吗？”耶稣回答：“是你说的。”
MARK|15|3|祭司长们告他许多的事。
MARK|15|4|彼拉多 又问他：“你看，他们告你这么多的事，你什么都不回答吗？”
MARK|15|5|耶稣仍不回答，以致 彼拉多 觉得惊讶。
MARK|15|6|每逢这节期， 彼拉多 照众人所求的，释放一个囚犯给他们。
MARK|15|7|有一个人名叫 巴拉巴 ，和作乱的人监禁在一起。他们作乱的时候曾杀过人。
MARK|15|8|众人上去求 彼拉多 照常例给他们办理。
MARK|15|9|彼拉多 说：“你们要我释放 犹太 人的王给你们吗？”
MARK|15|10|他原知道祭司长们是因嫉妒才把耶稣解了来。
MARK|15|11|但是祭司长们煽动众人，宁可要他释放 巴拉巴 给他们。
MARK|15|12|彼拉多 又说：“那么，你们称为 犹太 人的王的 ，要 我怎么办他呢？”
MARK|15|13|他们又再喊着：“把他钉十字架！”
MARK|15|14|彼拉多 说：“为什么？他做了什么恶事呢？”他们更加喊着：“把他钉十字架！”
MARK|15|15|彼拉多 要讨好众人，就释放 巴拉巴 给他们，把耶稣鞭打后交给人钉十字架。
MARK|15|16|士兵把耶稣带进总督府的庭院里，叫齐了全营的兵。
MARK|15|17|他们给他穿上紫袍，又用荆棘编了冠冕给他戴上，
MARK|15|18|然后向他致敬，说：“万岁， 犹太 人的王！”
MARK|15|19|他们又拿一根芦苇秆打他的头，向他吐唾沫，屈膝拜他。
MARK|15|20|他们戏弄完了，就给他脱了紫袍，又穿上他自己的衣服，带他出去，要把他钉十字架。
MARK|15|21|有一个 古利奈 人 西门 ，就是 亚历山大 和 鲁孚 的父亲，从乡下来，经过那地方，他们就强迫他同去，好背耶稣的十字架。
MARK|15|22|他们带耶稣到了一个地方叫 各各他 （翻出来就是“髑髅地”），
MARK|15|23|拿没药调和的酒给耶稣，他却不受。
MARK|15|24|于是他们把他钉在十字架上，抽签分他的衣服，看谁得什么。
MARK|15|25|他们把他钉十字架的时候是上午九点钟。
MARK|15|26|罪状牌上写的是：“ 犹太 人的王。”
MARK|15|27|他们又把两个强盗和他同钉十字架，一个在右边，一个在左边。
MARK|15|28|
MARK|15|29|从那里经过的人讥笑他，摇着头，说：“哼！你这拆毁殿、三日又建造起来的，
MARK|15|30|救救你自己，从十字架上下来呀！”
MARK|15|31|众祭司长和文士也这样嘲笑他，彼此说：“他救了别人，不能救自己。
MARK|15|32|以色列 的王基督，现在从十字架上下来，好让我们看见就信了呀！”那和他同钉的人也讥讽他。
MARK|15|33|到了正午，全地都黑暗了，直到下午三点钟。
MARK|15|34|下午三点钟的时候，耶稣大声呼喊：“以罗伊！以罗伊！拉马撒巴各大尼？”（翻出来就是：我的上帝！我的上帝！为什么离弃我？）
MARK|15|35|旁边站着的人，有的听见就说：“看哪，他叫 以利亚 呢！”
MARK|15|36|有一个人跑去，把海绵蘸满了醋，绑在芦苇秆上，送给他喝，说：“且等着，看 以利亚 会不会来把他放下来。”
MARK|15|37|耶稣大喊一声，气就断了。
MARK|15|38|殿的幔子从上到下裂为两半。
MARK|15|39|对面站着的百夫长看见耶稣这样断气 ，就说：“这人真是上帝的儿子！”
MARK|15|40|还有些妇女远远地观看，其中有 抹大拉 的 马利亚 ，又有小 雅各 和 约西 的母亲 马利亚 ，并有 撒罗米 ，
MARK|15|41|就是耶稣在 加利利 的时候，跟随他、服事他的那些人，还有同耶稣上 耶路撒冷 的好些妇女。
MARK|15|42|到了晚上，因为这是预备日，就是安息日的前一日，
MARK|15|43|有 亚利马太 的 约瑟 前来，他是尊贵的议员，也是盼望着上帝国的，他放胆进去见 彼拉多 ，请求要耶稣的身体。
MARK|15|44|彼拉多 诧异耶稣已经死了，就叫百夫长来，问他耶稣是不是死了很久；
MARK|15|45|既从百夫长得知实情，就把耶稣的身体赐给 约瑟 。
MARK|15|46|约瑟 买了细麻布，把耶稣取下来，用细麻布裹好，安放在岩石中凿出来的墓穴里，又滚来一块石头挡住墓门。
MARK|15|47|抹大拉 的 马利亚 和 约西 的母亲 马利亚 都看见安放他的地方。
MARK|16|1|过了安息日， 抹大拉 的 马利亚 、 雅各 的母亲 马利亚 ，和 撒罗米 ，买了香料，要去膏耶稣的身体。
MARK|16|2|七日的第一日清早，太阳出来后，她们来到坟墓那里，
MARK|16|3|彼此说：“谁要替我们把石头从墓门滚开呢？”
MARK|16|4|她们抬头一看，看见石头已经滚开了，原来那石头很大。
MARK|16|5|她们进了坟墓，看见一个年轻人坐在右边，穿着白袍，就很惊奇。
MARK|16|6|那年轻人对她们说：“不要惊慌！你们寻找那钉十字架的 拿撒勒 人耶稣，他已经复活了，不在这里。来看安放他的地方。
MARK|16|7|你们去，对他的门徒和 彼得 说：‘他要比你们先到 加利利 去，在那里你们会看见他，正如他从前所告诉你们的。’”
MARK|16|8|于是她们出来，从坟墓那里逃走，又发抖又惊讶，什么也没有告诉人，因为她们害怕。 〔
MARK|16|9|凡耶稣所吩咐的，她们简洁地告诉 彼得 和他周围的人。这些事以后，耶稣亲自藉着他的门徒，从东到西，把那神圣、不朽、永远拯救的福音传出去。阿们！〕 〔 在七日的第一日清早，耶稣复活了，先向 抹大拉 的 马利亚 显现；耶稣曾从她身上赶出七个鬼。
MARK|16|10|她去告诉那向来跟随耶稣的人；那时他们正哀恸哭泣。
MARK|16|11|他们听见耶稣活了，被 马利亚 看见，可是不信。〕 〔
MARK|16|12|这些事以后，门徒中有两个人往乡下去；正走着的时候，耶稣以另一种形像向他们显现。
MARK|16|13|他们去告诉其余的门徒，那些门徒还是不信。〕 〔
MARK|16|14|后来十一使徒坐席的时候，耶稣向他们显现，责备他们不信，心里刚硬，因为他们不信那些在他复活以后看见他的人。
MARK|16|15|他又对他们说：“你们往普天下去，传福音给万民 听。
MARK|16|16|信而受洗的必然得救，不信的必被定罪。
MARK|16|17|信的人将有神迹随着他们：就是奉我的名赶鬼；说新方言；
MARK|16|18|手 能拿蛇；若喝了什么毒物，也不会受害；手按病人，病人就好了。”〕 〔
MARK|16|19|主耶稣 和他们说完了话以后，被接到天上，坐在上帝的右边。
MARK|16|20|门徒出去，到处传福音。主和他们同工，藉着伴随的神迹证实所传的道。 〕
