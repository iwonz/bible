DAN|1|1|В третий год царствования Иоакима, царя Иудейского, пришел Навуходоносор, царь Вавилонский, к Иерусалиму и осадил его.
DAN|1|2|И предал Господь в руку его Иоакима, царя Иудейского, и часть сосудов дома Божия, и он отправил их в землю Сеннаар, в дом бога своего, и внес эти сосуды в сокровищницу бога своего.
DAN|1|3|И сказал царь Асфеназу, начальнику евнухов своих, чтобы он из сынов Израилевых, из рода царского и княжеского, привел
DAN|1|4|отроков, у которых нет никакого телесного недостатка, красивых видом, и понятливых для всякой науки, и разумеющих науки, и смышленых и годных служить в чертогах царских, и чтобы научил их книгам и языку Халдейскому.
DAN|1|5|И назначил им царь ежедневную пищу с царского стола и вино, которое сам пил, и велел воспитывать их три года, по истечении которых они должны были предстать пред царя.
DAN|1|6|Между ними были из сынов Иудиных Даниил, Анания, Мисаил и Азария.
DAN|1|7|И переименовал их начальник евнухов – Даниила Валтасаром, Ананию Седрахом, Мисаила Мисахом и Азарию Авденаго.
DAN|1|8|Даниил положил в сердце своем не оскверняться яствами со стола царского и вином, какое пьет царь, и потому просил начальника евнухов о том, чтобы не оскверняться ему.
DAN|1|9|Бог даровал Даниилу милость и благорасположение начальника евнухов;
DAN|1|10|и начальник евнухов сказал Даниилу: боюсь я господина моего, царя, который сам назначил вам пищу и питье; если он увидит лица ваши худощавее, нежели у отроков, сверстников ваших, то вы сделаете голову мою виновною перед царем.
DAN|1|11|Тогда сказал Даниил Амелсару, которого начальник евнухов приставил к Даниилу, Анании, Мисаилу и Азарии:
DAN|1|12|сделай опыт над рабами твоими в течение десяти дней; пусть дают нам в пищу овощи и воду для питья;
DAN|1|13|и потом пусть явятся перед тобою лица наши и лица тех отроков, которые питаются царскою пищею, и затем поступай с рабами твоими, как увидишь.
DAN|1|14|Он послушался их в этом и испытывал их десять дней.
DAN|1|15|По истечении же десяти дней лица их оказались красивее, и телом они были полнее всех тех отроков, которые питались царскими яствами.
DAN|1|16|Тогда Амелсар брал их кушанье и вино для питья и давал им овощи.
DAN|1|17|И даровал Бог четырем сим отрокам знание и разумение всякой книги и мудрости, а Даниилу еще даровал разуметь и всякие видения и сны.
DAN|1|18|По окончании тех дней, когда царь приказал представить их, начальник евнухов представил их Навуходоносору.
DAN|1|19|И царь говорил с ними, и из всех [отроков] не нашлось подобных Даниилу, Анании, Мисаилу и Азарии, и стали они служить пред царем.
DAN|1|20|И во всяком деле мудрого уразумения, о чем ни спрашивал их царь, он находил их в десять раз выше всех тайноведцев и волхвов, какие были во всем царстве его.
DAN|1|21|И был там Даниил до первого года царя Кира.
DAN|2|1|Во второй год царствования Навуходоносора снились Навуходоносору сны, и возмутился дух его, и сон удалился от него.
DAN|2|2|И велел царь созвать тайноведцев, и гадателей, и чародеев, и Халдеев, чтобы они рассказали царю сновидения его. Они пришли, и стали перед царем.
DAN|2|3|И сказал им царь: сон снился мне, и тревожится дух мой; желаю знать этот сон.
DAN|2|4|И сказали Халдеи царю по–арамейски: царь! вовеки живи! скажи сон рабам твоим, и мы объясним значение его.
DAN|2|5|Отвечал царь и сказал Халдеям: слово отступило от меня; если вы не скажете мне сновидения и значения его, то в куски будете изрублены, и домы ваши обратятся в развалины.
DAN|2|6|Если же расскажете сон и значение его, то получите от меня дары, награду и великую почесть; итак скажите мне сон и значение его.
DAN|2|7|Они вторично отвечали и сказали: да скажет царь рабам своим сновидение, и мы объясним его значение.
DAN|2|8|Отвечал царь и сказал: верно знаю, что вы хотите выиграть время, потому что видите, что слово отступило от меня.
DAN|2|9|Так как вы не объявляете мне сновидения, то у вас один умысел: вы собираетесь сказать мне ложь и обман, пока минет время; итак расскажите мне сон, и тогда я узнаю, что вы можете объяснить мне и значение его.
DAN|2|10|Халдеи отвечали царю и сказали: нет на земле человека, который мог бы открыть это дело царю, и потому ни один царь, великий и могущественный, не требовал подобного ни от какого тайноведца, гадателя и Халдея.
DAN|2|11|Дело, которого царь требует, так трудно, что никто другой не может открыть его царю, кроме богов, которых обитание не с плотью.
DAN|2|12|Рассвирепел царь и сильно разгневался на это, и приказал истребить всех мудрецов Вавилонских.
DAN|2|13|Когда вышло это повеление, чтобы убивать мудрецов, искали Даниила и товарищей его, чтобы умертвить их.
DAN|2|14|Тогда Даниил обратился с советом и мудростью к Ариоху, начальнику царских телохранителей, который вышел убивать мудрецов Вавилонских;
DAN|2|15|и спросил Ариоха, сильного при царе: "почему такое грозное повеление от царя?" Тогда Ариох рассказал все дело Даниилу.
DAN|2|16|И Даниил вошел, и упросил царя дать ему время, и он представит царю толкование [сна].
DAN|2|17|Даниил пришел в дом свой, и рассказал дело Анании, Мисаилу и Азарии, товарищам своим,
DAN|2|18|чтобы они просили милости у Бога небесного об этой тайне, дабы Даниил и товарищи его не погибли с прочими мудрецами Вавилонскими.
DAN|2|19|И тогда открыта была тайна Даниилу в ночном видении, и Даниил благословил Бога небесного.
DAN|2|20|И сказал Даниил: да будет благословенно имя Господа от века и до века! ибо у Него мудрость и сила;
DAN|2|21|он изменяет времена и лета, низлагает царей и поставляет царей; дает мудрость мудрым и разумение разумным;
DAN|2|22|он открывает глубокое и сокровенное, знает, что во мраке, и свет обитает с Ним.
DAN|2|23|Славлю и величаю Тебя, Боже отцов моих, что Ты даровал мне мудрость и силу и открыл мне то, о чем мы молили Тебя; ибо Ты открыл нам дело царя.
DAN|2|24|После сего Даниил вошел к Ариоху, которому царь повелел умертвить мудрецов Вавилонских, пришел и сказал ему: не убивай мудрецов Вавилонских; введи меня к царю, и я открою значение [сна].
DAN|2|25|Тогда Ариох немедленно привел Даниила к царю и сказал ему: я нашел из пленных сынов Иудеи человека, который может открыть царю значение [сна].
DAN|2|26|Царь сказал Даниилу, который назван был Валтасаром: можешь ли ты сказать мне сон, который я видел, и значение его?
DAN|2|27|Даниил отвечал царю и сказал: тайны, о которой царь спрашивает, не могут открыть царю ни мудрецы, ни обаятели, ни тайноведцы, ни гадатели.
DAN|2|28|Но есть на небесах Бог, открывающий тайны; и Он открыл царю Навуходоносору, что будет в последние дни. Сон твой и видения главы твоей на ложе твоем были такие:
DAN|2|29|ты, царь, на ложе твоем думал о том, что будет после сего? и Открывающий тайны показал тебе то, что будет.
DAN|2|30|А мне тайна сия открыта не потому, чтобы я был мудрее всех живущих, но для того, чтобы открыто было царю разумение и чтобы ты узнал помышления сердца твоего.
DAN|2|31|Тебе, царь, было такое видение: вот, какой–то большой истукан; огромный был этот истукан, в чрезвычайном блеске стоял он пред тобою, и страшен был вид его.
DAN|2|32|У этого истукана голова была из чистого золота, грудь его и руки его – из серебра, чрево его и бедра его медные,
DAN|2|33|голени его железные, ноги его частью железные, частью глиняные.
DAN|2|34|Ты видел его, доколе камень не оторвался от горы без содействия рук, ударил в истукана, в железные и глиняные ноги его, и разбил их.
DAN|2|35|Тогда все вместе раздробилось: железо, глина, медь, серебро и золото сделались как прах на летних гумнах, и ветер унес их, и следа не осталось от них; а камень, разбивший истукана, сделался великою горою и наполнил всю землю.
DAN|2|36|Вот сон! Скажем пред царем и значение его.
DAN|2|37|Ты, царь, царь царей, которому Бог небесный даровал царство, власть, силу и славу,
DAN|2|38|и всех сынов человеческих, где бы они ни жили, зверей земных и птиц небесных Он отдал в твои руки и поставил тебя владыкою над всеми ими. Ты – это золотая голова!
DAN|2|39|После тебя восстанет другое царство, ниже твоего, и еще третье царство, медное, которое будет владычествовать над всею землею.
DAN|2|40|А четвертое царство будет крепко, как железо; ибо как железо разбивает и раздробляет все, так и оно, подобно всесокрушающему железу, будет раздроблять и сокрушать.
DAN|2|41|А что ты видел ноги и пальцы на ногах частью из глины горшечной, а частью из железа, то будет царство разделенное, и в нем останется несколько крепости железа, так как ты видел железо, смешанное с горшечною глиною.
DAN|2|42|И как персты ног были частью из железа, а частью из глины, так и царство будет частью крепкое, частью хрупкое.
DAN|2|43|А что ты видел железо, смешанное с глиною горшечною, это значит, что они смешаются через семя человеческое, но не сольются одно с другим, как железо не смешивается с глиною.
DAN|2|44|И во дни тех царств Бог небесный воздвигнет царство, которое вовеки не разрушится, и царство это не будет передано другому народу; оно сокрушит и разрушит все царства, а само будет стоять вечно,
DAN|2|45|так как ты видел, что камень отторгнут был от горы не руками и раздробил железо, медь, глину, серебро и золото. Великий Бог дал знать царю, что будет после сего. И верен этот сон, и точно истолкование его!
DAN|2|46|Тогда царь Навуходоносор пал на лице свое и поклонился Даниилу, и велел принести ему дары и благовонные курения.
DAN|2|47|И сказал царь Даниилу: истинно Бог ваш есть Бог богов и Владыка царей, открывающий тайны, когда ты мог открыть эту тайну!
DAN|2|48|Тогда возвысил царь Даниила и дал ему много больших подарков, и поставил его над всею областью Вавилонскою и главным начальником над всеми мудрецами Вавилонскими.
DAN|2|49|Но Даниил просил царя, и он поставил Седраха, Мисаха и Авденаго над делами страны Вавилонской, а Даниил остался при дворе царя.
DAN|3|1|Царь Навуходоносор сделал золотой истукан, вышиною в шестьдесят локтей, шириною в шесть локтей, поставил его на поле Деире, в области Вавилонской.
DAN|3|2|И послал царь Навуходоносор собрать сатрапов, наместников, воевод, верховных судей, казнохранителей, законоведцев, блюстителей суда и всех областных правителей, чтобы они пришли на торжественное открытие истукана, которого поставил царь Навуходоносор.
DAN|3|3|И собрались сатрапы, наместники, военачальники, верховные судьи, казнохранители, законоведцы, блюстители суда и все областные правители на открытие истукана, которого Навуходоносор царь поставил, и стали перед истуканом, которого воздвиг Навуходоносор.
DAN|3|4|Тогда глашатай громко воскликнул: объявляется вам, народы, племена и языки:
DAN|3|5|в то время, как услышите звук трубы, свирели, цитры, цевницы, гуслей и симфонии и всяких музыкальных орудий, падите и поклонитесь золотому истукану, которого поставил царь Навуходоносор.
DAN|3|6|А кто не падет и не поклонится, тотчас брошен будет в печь, раскаленную огнем.
DAN|3|7|Посему, когда все народы услышали звук трубы, свирели, цитры, цевницы, гуслей и всякого рода музыкальных орудий, то пали все народы, племена и языки, и поклонились золотому истукану, которого поставил Навуходоносор царь.
DAN|3|8|В это самое время приступили некоторые из Халдеев и донесли на Иудеев.
DAN|3|9|Они сказали царю Навуходоносору: царь, вовеки живи!
DAN|3|10|Ты, царь, дал повеление, чтобы каждый человек, который услышит звук трубы, свирели, цитры, цевницы, гуслей и симфонии и всякого рода музыкальных орудий, пал и поклонился золотому истукану;
DAN|3|11|а кто не падет и не поклонится, тот должен быть брошен в печь, раскаленную огнем.
DAN|3|12|Есть мужи Иудейские, которых ты поставил над делами страны Вавилонской: Седрах, Мисах и Авденаго; эти мужи не повинуются повелению твоему, царь, богам твоим не служат и золотому истукану, которого ты поставил, не поклоняются.
DAN|3|13|Тогда Навуходоносор во гневе и ярости повелел привести Седраха, Мисаха и Авденаго; и приведены были эти мужи к царю.
DAN|3|14|Навуходоносор сказал им: с умыслом ли вы, Седрах, Мисах и Авденаго, богам моим не служите, и золотому истукану, которого я поставил, не поклоняетесь?
DAN|3|15|Отныне, если вы готовы, как скоро услышите звук трубы, свирели, цитры, цевницы, гуслей, симфонии и всякого рода музыкальных орудий, падите и поклонитесь истукану, которого я сделал; если же не поклонитесь, то в тот же час брошены будете в печь, раскаленную огнем, и тогда какой Бог избавит вас от руки моей?
DAN|3|16|И отвечали Седрах, Мисах и Авденаго, и сказали царю Навуходоносору: нет нужды нам отвечать тебе на это.
DAN|3|17|Бог наш, Которому мы служим, силен спасти нас от печи, раскаленной огнем, и от руки твоей, царь, избавит.
DAN|3|18|Если же и не будет того, то да будет известно тебе, царь, что мы богам твоим служить не будем и золотому истукану, которого ты поставил, не поклонимся.
DAN|3|19|Тогда Навуходоносор исполнился ярости, и вид лица его изменился на Седраха, Мисаха и Авденаго, и он повелел разжечь печь в семь раз сильнее, нежели как обыкновенно разжигали ее,
DAN|3|20|и самым сильным мужам из войска своего приказал связать Седраха, Мисаха и Авденаго и бросить их в печь, раскаленную огнем.
DAN|3|21|Тогда мужи сии связаны были в исподнем и верхнем платье своем, в головных повязках и в прочих одеждах своих, и брошены в печь, раскаленную огнем.
DAN|3|22|И как повеление царя было строго, и печь раскалена была чрезвычайно, то пламя огня убило тех людей, которые бросали Седраха, Мисаха и Авденаго.
DAN|3|23|А сии три мужа, Седрах, Мисах и Авденаго, упали в раскаленную огнем печь связанные.
DAN|3|24|Навуходоносор царь изумился, и поспешно встал, и сказал вельможам своим: не троих ли мужей бросили мы в огонь связанными? Они в ответ сказали царю: истинно так, царь!
DAN|3|25|На это он сказал: вот, я вижу четырех мужей несвязанных, ходящих среди огня, и нет им вреда; и вид четвертого подобен сыну Божию.
DAN|3|26|Тогда подошел Навуходоносор к устью печи, раскаленной огнем, и сказал: Седрах, Мисах и Авденаго, рабы Бога Всевышнего! выйдите и подойдите! Тогда Седрах, Мисах и Авденаго вышли из среды огня.
DAN|3|27|И, собравшись, сатрапы, наместники, военачальники и советники царя усмотрели, что над телами мужей сих огонь не имел силы, и волосы на голове не опалены, и одежды их не изменились, и даже запаха огня не было от них.
DAN|3|28|Тогда Навуходоносор сказал: благословен Бог Седраха, Мисаха и Авденаго, Который послал Ангела Своего и избавил рабов Своих, которые надеялись на Него и не послушались царского повеления, и предали тела свои [огню], чтобы не служить и не поклоняться иному богу, кроме Бога своего!
DAN|3|29|И от меня дается повеление, чтобы из всякого народа, племени и языка кто произнесет хулу на Бога Седраха, Мисаха и Авденаго, был изрублен в куски, и дом его обращен в развалины, ибо нет иного бога, который мог бы так спасать.
DAN|3|30|Тогда царь возвысил Седраха, Мисаха и Авденаго в стране Вавилонской.
DAN|3|31|Навуходоносор царь всем народам, племенам и языкам, живущим
DAN|3|32|Знамения и чудеса, какие совершил надо мною Всевышний Бог, угодно мне возвестить вам.
DAN|3|33|Как велики знамения Его и как могущественны чудеса Его! Царство Его – царство вечное, и владычество Его – в роды и роды.
DAN|4|1|Я, Навуходоносор, спокоен был в доме моем и благоденствовал в чертогах моих.
DAN|4|2|Но я видел сон, который устрашил меня, и размышления на ложе моем и видения головы моей смутили меня.
DAN|4|3|И дано было мною повеление привести ко мне всех мудрецов Вавилонских, чтобы они сказали мне значение сна.
DAN|4|4|Тогда пришли тайноведцы, обаятели, Халдеи и гадатели; я рассказал им сон, но они не могли мне объяснить значения его.
DAN|4|5|Наконец вошел ко мне Даниил, которому имя было Валтасар, по имени бога моего, и в котором дух святаго Бога; ему рассказал я сон.
DAN|4|6|Валтасар, глава мудрецов! я знаю, что в тебе дух святаго Бога, и никакая тайна не затрудняет тебя; объясни мне видения сна моего, который я видел, и значение его.
DAN|4|7|Видения же головы моей на ложе моем были такие: я видел, вот, среди земли дерево весьма высокое.
DAN|4|8|Большое было это дерево и крепкое, и высота его достигала до неба, и оно видимо было до краев всей земли.
DAN|4|9|Листья его прекрасные, и плодов на нем множество, и пища на нем для всех; под ним находили тень полевые звери, и в ветвях его гнездились птицы небесные, и от него питалась всякая плоть.
DAN|4|10|И видел я в видениях головы моей на ложе моем, и вот, нисшел с небес Бодрствующий и Святый.
DAN|4|11|Воскликнув громко, Он сказал: "срубите это дерево, обрубите ветви его, стрясите листья с него и разбросайте плоды его; пусть удалятся звери из–под него и птицы с ветвей его;
DAN|4|12|но главный корень его оставьте в земле, и пусть он в узах железных и медных среди полевой травы орошается небесною росою, и с животными пусть будет часть его в траве земной.
DAN|4|13|Сердце человеческое отнимется от него и дастся ему сердце звериное, и пройдут над ним семь времен.
DAN|4|14|Повелением Бодрствующих это определено, и по приговору Святых назначено, дабы знали живущие, что Всевышний владычествует над царством человеческим, и дает его, кому хочет, и поставляет над ним уничиженного между людьми".
DAN|4|15|Такой сон видел я, царь Навуходоносор; а ты, Валтасар, скажи значение его, так как никто из мудрецов в моем царстве не мог объяснить его значения, а ты можешь, потому что дух святаго Бога в тебе.
DAN|4|16|Тогда Даниил, которому имя Валтасар, около часа пробыл в изумлении, и мысли его смущали его. Царь начал говорить и сказал: Валтасар! да не смущает тебя этот сон и значение его. Валтасар отвечал и сказал: господин мой! твоим бы ненавистникам этот сон, и врагам твоим значение его!
DAN|4|17|Дерево, которое ты видел, которое было большое и крепкое, высотою своею достигало до небес и видимо было по всей земле,
DAN|4|18|на котором листья были прекрасные и множество плодов и пропитание для всех, под которым обитали звери полевые и в ветвях которого гнездились птицы небесные,
DAN|4|19|это ты, царь, возвеличившийся и укрепившийся, и величие твое возросло и достигло до небес, и власть твоя – до краев земли.
DAN|4|20|А что царь видел Бодрствующего и Святаго, сходящего с небес, Который сказал: "срубите дерево и истребите его, только главный корень его оставьте в земле, и пусть он в узах железных и медных, среди полевой травы, орошается росою небесною, и с полевыми зверями пусть будет часть его, доколе не пройдут над ним семь времен", –
DAN|4|21|то вот значение этого, царь, и вот определение Всевышнего, которое постигнет господина моего, царя:
DAN|4|22|тебя отлучат от людей, и обитание твое будет с полевыми зверями; травою будут кормить тебя, как вола, росою небесною ты будешь орошаем, и семь времен пройдут над тобою, доколе познаешь, что Всевышний владычествует над царством человеческим и дает его, кому хочет.
DAN|4|23|А что повелено было оставить главный корень дерева, это значит, что царство твое останется при тебе, когда ты познаешь власть небесную.
DAN|4|24|Посему, царь, да будет благоугоден тебе совет мой: искупи грехи твои правдою и беззакония твои милосердием к бедным; вот чем может продлиться мир твой.
DAN|4|25|Все это сбылось над царем Навуходоносором.
DAN|4|26|По прошествии двенадцати месяцев, расхаживая по царским чертогам в Вавилоне,
DAN|4|27|царь сказал: это ли не величественный Вавилон, который построил я в дом царства силою моего могущества и в славу моего величия!
DAN|4|28|Еще речь сия была в устах царя, как был с неба голос: "тебе говорят, царь Навуходоносор: царство отошло от тебя!
DAN|4|29|И отлучат тебя от людей, и будет обитание твое с полевыми зверями; травою будут кормить тебя, как вола, и семь времен пройдут над тобою, доколе познаешь, что Всевышний владычествует над царством человеческим и дает его, кому хочет!"
DAN|4|30|Тотчас и исполнилось это слово над Навуходоносором, и отлучен он был от людей, ел траву, как вол, и орошалось тело его росою небесною, так что волосы у него выросли как у льва, и ногти у него – как у птицы.
DAN|4|31|По окончании же дней тех, я, Навуходоносор, возвел глаза мои к небу, и разум мой возвратился ко мне; и благословил я Всевышнего, восхвалил и прославил Присносущего, Которого владычество – владычество вечное, и Которого царство – в роды и роды.
DAN|4|32|И все, живущие на земле, ничего не значат; по воле Своей Он действует как в небесном воинстве, так и у живущих на земле; и нет никого, кто мог бы противиться руке Его и сказать Ему: "что Ты сделал?"
DAN|4|33|В то время возвратился ко мне разум мой, и к славе царства моего возвратились ко мне сановитость и прежний вид мой; тогда взыскали меня советники мои и вельможи мои, и я восстановлен на царство мое, и величие мое еще более возвысилось.
DAN|4|34|Ныне я, Навуходоносор, славлю, превозношу и величаю Царя Небесного, Которого все дела истинны и пути праведны, и Который силен смирить ходящих гордо.
DAN|5|1|Валтасар царь сделал большое пиршество для тысячи вельмож своих и перед глазами тысячи пил вино.
DAN|5|2|Вкусив вина, Валтасар приказал принести золотые и серебряные сосуды, которые Навуходоносор, отец его, вынес из храма Иерусалимского, чтобы пить из них царю, вельможам его, женам его и наложницам его.
DAN|5|3|Тогда принесли золотые сосуды, которые взяты были из святилища дома Божия в Иерусалиме; и пили из них царь и вельможи его, жены его и наложницы его.
DAN|5|4|Пили вино, и славили богов золотых и серебряных, медных, железных, деревянных и каменных.
DAN|5|5|В тот самый час вышли персты руки человеческой и писали против лампады на извести стены чертога царского, и царь видел кисть руки, которая писала.
DAN|5|6|Тогда царь изменился в лице своем; мысли его смутили его, связи чресл его ослабели, и колени его стали биться одно о другое.
DAN|5|7|Сильно закричал царь, чтобы привели обаятелей, Халдеев и гадателей. Царь начал говорить, и сказал мудрецам Вавилонским: кто прочитает это написанное и объяснит мне значение его, тот будет облечен в багряницу, и золотая цепь будет на шее у него, и третьим властелином будет в царстве.
DAN|5|8|И вошли все мудрецы царя, но не могли прочитать написанного и объяснить царю значения его.
DAN|5|9|Царь Валтасар чрезвычайно встревожился, и вид лица его изменился на нем, и вельможи его смутились.
DAN|5|10|Царица же, по поводу слов царя и вельмож его, вошла в палату пиршества; начала говорить царица и сказала: царь, вовеки живи! да не смущают тебя мысли твои, и да не изменяется вид лица твоего!
DAN|5|11|Есть в царстве твоем муж, в котором дух святаго Бога; во дни отца твоего найдены были в нем свет, разум и мудрость, подобная мудрости богов, и царь Навуходоносор, отец твой, поставил его главою тайноведцев, обаятелей, Халдеев и гадателей, – сам отец твой, царь,
DAN|5|12|потому что в нем, в Данииле, которого царь переименовал Валтасаром, оказались высокий дух, ведение и разум, способный изъяснять сны, толковать загадочное и разрешать узлы. Итак пусть призовут Даниила и он объяснит значение.
DAN|5|13|Тогда введен был Даниил пред царя, и царь начал речь и сказал Даниилу: ты ли Даниил, один из пленных сынов Иудейских, которых отец мой, царь, привел из Иудеи?
DAN|5|14|Я слышал о тебе, что дух Божий в тебе и свет, и разум, и высокая мудрость найдена в тебе.
DAN|5|15|Вот, приведены были ко мне мудрецы и обаятели, чтобы прочитать это написанное и объяснить мне значение его; но они не могли объяснить мне этого.
DAN|5|16|А о тебе я слышал, что ты можешь объяснять значение и разрешать узлы; итак, если можешь прочитать это написанное и объяснить мне значение его, то облечен будешь в багряницу, и золотая цепь будет на шее твоей, и третьим властелином будешь в царстве.
DAN|5|17|Тогда отвечал Даниил, и сказал царю: дары твои пусть останутся у тебя, и почести отдай другому; а написанное я прочитаю царю и значение объясню ему.
DAN|5|18|Царь! Всевышний Бог даровал отцу твоему Навуходоносору царство, величие, честь и славу.
DAN|5|19|Пред величием, которое Он дал ему, все народы, племена и языки трепетали и страшились его: кого хотел, он убивал, и кого хотел, оставлял в живых; кого хотел, возвышал, и кого хотел, унижал.
DAN|5|20|Но когда сердце его надмилось и дух его ожесточился до дерзости, он был свержен с царского престола своего и лишен славы своей,
DAN|5|21|и отлучен был от сынов человеческих, и сердце его уподобилось звериному, и жил он с дикими ослами; кормили его травою, как вола, и тело его орошаемо было небесною росою, доколе он познал, что над царством человеческим владычествует Всевышний Бог и поставляет над ним, кого хочет.
DAN|5|22|И ты, сын его Валтасар, не смирил сердца твоего, хотя знал все это,
DAN|5|23|но вознесся против Господа небес, и сосуды дома Его принесли к тебе, и ты и вельможи твои, жены твои и наложницы твои пили из них вино, и ты славил богов серебряных и золотых, медных, железных, деревянных и каменных, которые ни видят, ни слышат, ни разумеют; а Бога, в руке Которого дыхание твое и у Которого все пути твои, ты не прославил.
DAN|5|24|За это и послана от Него кисть руки, и начертано это писание.
DAN|5|25|И вот что начертано: мене, мене, текел, упарсин.
DAN|5|26|Вот и значение слов: мене – исчислил Бог царство твое и положил конец ему;
DAN|5|27|Текел – ты взвешен на весах и найден очень легким;
DAN|5|28|Перес – разделено царство твое и дано Мидянам и Персам.
DAN|5|29|Тогда по повелению Валтасара облекли Даниила в багряницу и возложили золотую цепь на шею его, и провозгласили его третьим властелином в царстве.
DAN|5|30|В ту же самую ночь Валтасар, царь Халдейский, был убит,
DAN|5|31|и Дарий Мидянин принял царство, будучи шестидесяти двух лет.
DAN|6|1|Угодно было Дарию поставить над царством сто двадцать сатрапов, чтобы они были во всем царстве,
DAN|6|2|а над ними трех князей, – из которых один был Даниил, – чтобы сатрапы давали им отчет и чтобы царю не было никакого обременения.
DAN|6|3|Даниил превосходил прочих князей и сатрапов, потому что в нем был высокий дух, и царь помышлял уже поставить его над всем царством.
DAN|6|4|Тогда князья и сатрапы начали искать предлога к обвинению Даниила по управлению царством; но никакого предлога и погрешностей не могли найти, потому что он был верен, и никакой погрешности или вины не оказывалось в нем.
DAN|6|5|И эти люди сказали: не найти нам предлога против Даниила, если мы не найдем его против него в законе Бога его.
DAN|6|6|Тогда эти князья и сатрапы приступили к царю и так сказали ему: царь Дарий! вовеки живи!
DAN|6|7|Все князья царства, наместники, сатрапы, советники и военачальники согласились между собою, чтобы сделано было царское постановление и издано повеление, чтобы, кто в течение тридцати дней будет просить какого–либо бога или человека, кроме тебя, царь, того бросить в львиный ров.
DAN|6|8|Итак утверди, царь, это определение и подпиши указ, чтобы он был неизменен, как закон Мидийский и Персидский, и чтобы он не был нарушен.
DAN|6|9|Царь Дарий подписал указ и это повеление.
DAN|6|10|Даниил же, узнав, что подписан такой указ, пошел в дом свой; окна же в горнице его были открыты против Иерусалима, и он три раза в день преклонял колени, и молился своему Богу, и славословил Его, как это делал он и прежде того.
DAN|6|11|Тогда эти люди подсмотрели и нашли Даниила молящегося и просящего милости пред Богом своим,
DAN|6|12|потом пришли и сказали царю о царском повелении: не ты ли подписал указ, чтобы всякого человека, который в течение тридцати дней будет просить какого–либо бога или человека, кроме тебя, царь, бросать в львиный ров? Царь отвечал и сказал: это слово твердо, как закон Мидян и Персов, не допускающий изменения.
DAN|6|13|Тогда отвечали они и сказали царю, что Даниил, который из пленных сынов Иудеи, не обращает внимания ни на тебя, царь, ни на указ, тобою подписанный, но три раза в день молится своими молитвами.
DAN|6|14|Царь, услышав это, сильно опечалился и положил в сердце своем спасти Даниила, и даже до захождения солнца усиленно старался избавить его.
DAN|6|15|Но те люди приступили к царю и сказали ему: знай, царь, что по закону Мидян и Персов никакое определение или постановление, утвержденное царем, не может быть изменено.
DAN|6|16|Тогда царь повелел, и привели Даниила, и бросили в ров львиный; при этом царь сказал Даниилу: Бог твой, Которому ты неизменно служишь, Он спасет тебя!
DAN|6|17|И принесен был камень и положен на отверстие рва, и царь запечатал его перстнем своим, и перстнем вельмож своих, чтобы ничто не переменилось в распоряжении о Данииле.
DAN|6|18|Затем царь пошел в свой дворец, лег спать без ужина, и даже не велел вносить к нему пищи, и сон бежал от него.
DAN|6|19|Поутру же царь встал на рассвете и поспешно пошел ко рву львиному,
DAN|6|20|и, подойдя ко рву, жалобным голосом кликнул Даниила, и сказал царь Даниилу: Даниил, раб Бога живаго! Бог твой, Которому ты неизменно служишь, мог ли спасти тебя от львов?
DAN|6|21|Тогда Даниил сказал царю: царь! вовеки живи!
DAN|6|22|Бог мой послал Ангела Своего и заградил пасть львам, и они не повредили мне, потому что я оказался пред Ним чист, да и перед тобою, царь, я не сделал преступления.
DAN|6|23|Тогда царь чрезвычайно возрадовался о нем и повелел поднять Даниила изо рва; и поднят был Даниил изо рва, и никакого повреждения не оказалось на нем, потому что он веровал в Бога своего.
DAN|6|24|И приказал царь, и приведены были те люди, которые обвиняли Даниила, и брошены в львиный ров, как они сами, так и дети их и жены их; и они не достигли до дна рва, как львы овладели ими и сокрушили все кости их.
DAN|6|25|После того царь Дарий написал всем народам, племенам и языкам, живущим по всей земле: "Мир вам да умножится!
DAN|6|26|Мною дается повеление, чтобы во всякой области царства моего трепетали и благоговели пред Богом Данииловым, потому что Он есть Бог живый и присносущий, и царство Его несокрушимо, и владычество Его бесконечно.
DAN|6|27|Он избавляет и спасает, и совершает чудеса и знамения на небе и на земле; Он избавил Даниила от силы львов".
DAN|6|28|И Даниил благоуспевал и в царствование Дария, и в царствование Кира Персидского.
DAN|7|1|В первый год Валтасара, царя Вавилонского, Даниил видел сон и пророческие видения головы своей на ложе своем. Тогда он записал этот сон, изложив сущность дела.
DAN|7|2|Начав речь, Даниил сказал: видел я в ночном видении моем, и вот, четыре ветра небесных боролись на великом море,
DAN|7|3|и четыре больших зверя вышли из моря, непохожие один на другого.
DAN|7|4|Первый – как лев, но у него крылья орлиные; я смотрел, доколе не вырваны были у него крылья, и он поднят был от земли, и стал на ноги, как человек, и сердце человеческое дано ему.
DAN|7|5|И вот еще зверь, второй, похожий на медведя, стоял с одной стороны, и три клыка во рту у него, между зубами его; ему сказано так: "встань, ешь мяса много!"
DAN|7|6|Затем видел я, вот еще зверь, как барс; на спине у него четыре птичьих крыла, и четыре головы были у зверя сего, и власть дана была ему.
DAN|7|7|После сего видел я в ночных видениях, и вот зверь четвертый, страшный и ужасный и весьма сильный; у него большие железные зубы; он пожирает и сокрушает, остатки же попирает ногами; он отличен был от всех прежних зверей, и десять рогов было у него.
DAN|7|8|Я смотрел на эти рога, и вот, вышел между ними еще небольшой рог, и три из прежних рогов с корнем исторгнуты были перед ним, и вот, в этом роге были глаза, как глаза человеческие, и уста, говорящие высокомерно.
DAN|7|9|Видел я, наконец, что поставлены были престолы, и воссел Ветхий днями; одеяние на Нем было бело, как снег, и волосы главы Его – как чистая волна; престол Его – как пламя огня, колеса Его – пылающий огонь.
DAN|7|10|Огненная река выходила и проходила пред Ним; тысячи тысяч служили Ему и тьмы тем предстояли пред Ним; судьи сели, и раскрылись книги.
DAN|7|11|Видел я тогда, что за изречение высокомерных слов, какие говорил рог, зверь был убит в глазах моих, и тело его сокрушено и предано на сожжение огню.
DAN|7|12|И у прочих зверей отнята власть их, и продолжение жизни дано им только на время и на срок.
DAN|7|13|Видел я в ночных видениях, вот, с облаками небесными шел как бы Сын человеческий, дошел до Ветхого днями и подведен был к Нему.
DAN|7|14|И Ему дана власть, слава и царство, чтобы все народы, племена и языки служили Ему; владычество Его – владычество вечное, которое не прейдет, и царство Его не разрушится.
DAN|7|15|Вострепетал дух мой во мне, Данииле, в теле моем, и видения головы моей смутили меня.
DAN|7|16|Я подошел к одному из предстоящих и спросил у него об истинном значении всего этого, и он стал говорить со мною, и объяснил мне смысл сказанного:
DAN|7|17|"эти большие звери, которых четыре, [означают], что четыре царя восстанут от земли.
DAN|7|18|Потом примут царство святые Всевышнего и будут владеть царством вовек и вовеки веков".
DAN|7|19|Тогда пожелал я точного объяснения о четвертом звере, который был отличен от всех и очень страшен, с зубами железными и когтями медными, пожирал и сокрушал, а остатки попирал ногами,
DAN|7|20|и о десяти рогах, которые были на голове у него, и о другом, вновь вышедшем, перед которым выпали три, о том самом роге, у которого были глаза и уста, говорящие высокомерно, и который по виду стал больше прочих.
DAN|7|21|Я видел, как этот рог вел брань со святыми и превозмогал их,
DAN|7|22|доколе не пришел Ветхий днями, и суд дан был святым Всевышнего, и наступило время, чтобы царством овладели святые.
DAN|7|23|Об этом он сказал: зверь четвертый – четвертое царство будет на земле, отличное от всех царств, которое будет пожирать всю землю, попирать и сокрушать ее.
DAN|7|24|А десять рогов значат, что из этого царства восстанут десять царей, и после них восстанет иной, отличный от прежних, и уничижит трех царей,
DAN|7|25|и против Всевышнего будет произносить слова и угнетать святых Всевышнего; даже возмечтает отменить у них [праздничные] времена и закон, и они преданы будут в руку его до времени и времен и полувремени.
DAN|7|26|Затем воссядут судьи и отнимут у него власть губить и истреблять до конца.
DAN|7|27|Царство же и власть и величие царственное во всей поднебесной дано будет народу святых Всевышнего, Которого царство – царство вечное, и все властители будут служить и повиноваться Ему.
DAN|7|28|Здесь конец слова. Меня, Даниила, сильно смущали размышления мои, и лице мое изменилось на мне; но слово я сохранил в сердце моем.
DAN|8|1|В третий год царствования Валтасара царя явилось мне, Даниилу, видение после того, которое явилось мне прежде.
DAN|8|2|И видел я в видении, и когда видел, я был в Сузах, престольном городе в области Еламской, и видел я в видении, – как бы я был у реки Улая.
DAN|8|3|Поднял я глаза мои и увидел: вот, один овен стоит у реки; у него два рога, и рога высокие, но один выше другого, и высший поднялся после.
DAN|8|4|Видел я, как этот овен бодал к западу и к северу и к югу, и никакой зверь не мог устоять против него, и никто не мог спасти от него; он делал, что хотел, и величался.
DAN|8|5|Я внимательно смотрел на это, и вот, с запада шел козел по лицу всей земли, не касаясь земли; у этого козла был видный рог между его глазами.
DAN|8|6|Он пошел на того овна, имеющего рога, которого я видел стоящим у реки, и бросился на него в сильной ярости своей.
DAN|8|7|И я видел, как он, приблизившись к овну, рассвирепел на него и поразил овна, и сломил у него оба рога; и недостало силы у овна устоять против него, и он поверг его на землю и растоптал его, и не было никого, кто мог бы спасти овна от него.
DAN|8|8|Тогда козел чрезвычайно возвеличился; но когда он усилился, то сломился большой рог, и на место его вышли четыре, обращенные на четыре ветра небесных.
DAN|8|9|От одного из них вышел небольшой рог, который чрезвычайно разросся к югу и к востоку и к прекрасной стране,
DAN|8|10|и вознесся до воинства небесного, и низринул на землю часть сего воинства и звезд, и попрал их,
DAN|8|11|и даже вознесся на Вождя воинства сего, и отнята была у Него ежедневная жертва, и поругано было место святыни Его.
DAN|8|12|И воинство предано вместе с ежедневною жертвою за нечестие, и он, повергая истину на землю, действовал и успевал.
DAN|8|13|И услышал я одного святого говорящего, и сказал этот святой кому–то, вопрошавшему: "на сколько времени простирается это видение о ежедневной жертве и об опустошительном нечестии, когда святыня и воинство будут попираемы?"
DAN|8|14|И сказал мне: "на две тысячи триста вечеров и утр; и тогда святилище очистится".
DAN|8|15|И было: когда я, Даниил, увидел это видение и искал значения его, вот, стал предо мною как облик мужа.
DAN|8|16|И услышал я от средины Улая голос человеческий, который воззвал и сказал: "Гавриил! объясни ему это видение!"
DAN|8|17|И он подошел к тому месту, где я стоял, и когда он пришел, я ужаснулся и пал на лице мое; и сказал он мне: "знай, сын человеческий, что видение относится к концу времени!"
DAN|8|18|И когда он говорил со мною, я без чувств лежал лицем моим на земле; но он прикоснулся ко мне и поставил меня на место мое,
DAN|8|19|и сказал: "вот, я открываю тебе, что будет в последние дни гнева; ибо это относится к концу определенного времени.
DAN|8|20|Овен, которого ты видел с двумя рогами, это цари Мидийский и Персидский.
DAN|8|21|А козел косматый – царь Греции, а большой рог, который между глазами его, это первый ее царь;
DAN|8|22|он сломился, и вместо него вышли другие четыре: это – четыре царства восстанут из этого народа, но не с его силою.
DAN|8|23|Под конец же царства их, когда отступники исполнят меру беззаконий своих, восстанет царь наглый и искусный в коварстве;
DAN|8|24|и укрепится сила его, хотя и не его силою, и он будет производить удивительные опустошения и успевать и действовать и губить сильных и народ святых,
DAN|8|25|и при уме его и коварство будет иметь успех в руке его, и сердцем своим он превознесется, и среди мира погубит многих, и против Владыки владык восстанет, но будет сокрушен – не рукою.
DAN|8|26|Видение же о вечере и утре, о котором сказано, истинно; но ты сокрой это видение, ибо оно относится к отдаленным временам".
DAN|8|27|И я, Даниил, изнемог, и болел несколько дней; потом встал и начал заниматься царскими делами; я изумлен был видением сим и не понимал его.
DAN|9|1|В первый год Дария, сына Ассуирова, из рода Мидийского, который поставлен был царем над царством Халдейским,
DAN|9|2|в первый год царствования его я, Даниил, сообразил по книгам число лет, о котором было слово Господне к Иеремии пророку, что семьдесят лет исполнятся над опустошением Иерусалима.
DAN|9|3|И обратил я лице мое к Господу Богу с молитвою и молением, в посте и вретище и пепле.
DAN|9|4|И молился я Господу Богу моему, и исповедывался и сказал: "Молю Тебя, Господи Боже великий и дивный, хранящий завет и милость любящим Тебя и соблюдающим повеления Твои!
DAN|9|5|Согрешили мы, поступали беззаконно, действовали нечестиво, упорствовали и отступили от заповедей Твоих и от постановлений Твоих;
DAN|9|6|и не слушали рабов Твоих, пророков, которые Твоим именем говорили царям нашим, и вельможам нашим, и отцам нашим, и всему народу страны.
DAN|9|7|У Тебя, Господи, правда, а у нас на лицах стыд, как день сей, у каждого Иудея, у жителей Иерусалима и у всего Израиля, у ближних и дальних, во всех странах, куда Ты изгнал их за отступление их, с каким они отступили от Тебя.
DAN|9|8|Господи! у нас на лицах стыд, у царей наших, у князей наших и у отцов наших, потому что мы согрешили пред Тобою.
DAN|9|9|А у Господа Бога нашего милосердие и прощение, ибо мы возмутились против Него
DAN|9|10|и не слушали гласа Господа Бога нашего, чтобы поступать по законам Его, которые Он дал нам через рабов Своих, пророков.
DAN|9|11|И весь Израиль преступил закон Твой и отвратился, чтобы не слушать гласа Твоего; и за то излились на нас проклятие и клятва, которые написаны в законе Моисея, раба Божия: ибо мы согрешили пред Ним.
DAN|9|12|И Он исполнил слова Свои, которые изрек на нас и на судей наших, судивших нас, наведя на нас великое бедствие, какого не бывало под небесами и какое совершилось над Иерусалимом.
DAN|9|13|Как написано в законе Моисея, так все это бедствие постигло нас; но мы не умоляли Господа Бога нашего, чтобы нам обратиться от беззаконий наших и уразуметь истину Твою.
DAN|9|14|Наблюдал Господь это бедствие и навел его на нас: ибо праведен Господь Бог наш во всех делах Своих, которые совершает, но мы не слушали гласа Его.
DAN|9|15|И ныне, Господи Боже наш, изведший народ Твой из земли Египетской рукою сильною и явивший славу Твою, как день сей! согрешили мы, поступали нечестиво.
DAN|9|16|Господи! по всей правде Твоей да отвратится гнев Твой и негодование Твое от града Твоего, Иерусалима, от святой горы Твоей; ибо за грехи наши и беззакония отцов наших Иерусалим и народ Твой в поругании у всех, окружающих нас.
DAN|9|17|И ныне услыши, Боже наш, молитву раба Твоего и моление его и воззри светлым лицем Твоим на опустошенное святилище Твое, ради Тебя, Господи.
DAN|9|18|Приклони, Боже мой, ухо Твое и услыши, открой очи Твои и воззри на опустошения наши и на город, на котором наречено имя Твое; ибо мы повергаем моления наши пред Тобою, уповая не на праведность нашу, но на Твое великое милосердие.
DAN|9|19|Господи! услыши; Господи! прости; Господи! внемли и соверши, не умедли ради Тебя Самого, Боже мой, ибо Твое имя наречено на городе Твоем и на народе Твоем".
DAN|9|20|И когда я еще говорил и молился, и исповедывал грехи мои и грехи народа моего, Израиля, и повергал мольбу мою пред Господом Богом моим о святой горе Бога моего;
DAN|9|21|когда я еще продолжал молитву, муж Гавриил, которого я видел прежде в видении, быстро прилетев, коснулся меня около времени вечерней жертвы
DAN|9|22|и вразумлял меня, говорил со мною и сказал: "Даниил! теперь я исшел, чтобы научить тебя разумению.
DAN|9|23|В начале моления твоего вышло слово, и я пришел возвестить [его] [тебе], ибо ты муж желаний; итак вникни в слово и уразумей видение.
DAN|9|24|Семьдесят седмин определены для народа твоего и святаго города твоего, чтобы покрыто было преступление, запечатаны были грехи и заглажены беззакония, и чтобы приведена была правда вечная, и запечатаны были видение и пророк, и помазан был Святый святых.
DAN|9|25|Итак знай и разумей: с того времени, как выйдет повеление о восстановлении Иерусалима, до Христа Владыки семь седмин и шестьдесят две седмины; и возвратится [народ] и обстроятся улицы и стены, но в трудные времена.
DAN|9|26|И по истечении шестидесяти двух седмин предан будет смерти Христос, и не будет; а город и святилище разрушены будут народом вождя, который придет, и конец его будет как от наводнения, и до конца войны будут опустошения.
DAN|9|27|И утвердит завет для многих одна седмина, а в половине седмины прекратится жертва и приношение, и на крыле [святилища] будет мерзость запустения, и окончательная предопределенная гибель постигнет опустошителя".
DAN|10|1|В третий год Кира, царя Персидского, было откровение Даниилу, который назывался именем Валтасара; и истинно было это откровение и великой силы. Он понял это откровение и уразумел это видение.
DAN|10|2|В эти дни я, Даниил, был в сетовании три седмицы дней.
DAN|10|3|Вкусного хлеба я не ел; мясо и вино не входило в уста мои, и мастями я не умащал себя до исполнения трех седмиц дней.
DAN|10|4|А в двадцать четвертый день первого месяца был я на берегу большой реки Тигра,
DAN|10|5|и поднял глаза мои, и увидел: вот один муж, облеченный в льняную одежду, и чресла его опоясаны золотом из Уфаза.
DAN|10|6|Тело его – как топаз, лице его – как вид молнии; очи его – как горящие светильники, руки его и ноги его по виду – как блестящая медь, и глас речей его – как голос множества людей.
DAN|10|7|И только один я, Даниил, видел это видение, а бывшие со мною люди не видели этого видения; но сильный страх напал на них и они убежали, чтобы скрыться.
DAN|10|8|И остался я один и смотрел на это великое видение, но во мне не осталось крепости, и вид лица моего чрезвычайно изменился, не стало во мне бодрости.
DAN|10|9|И услышал я глас слов его; и как только услышал глас слов его, в оцепенении пал я на лице мое и лежал лицем к земле.
DAN|10|10|Но вот, коснулась меня рука и поставила меня на колени мои и на длани рук моих.
DAN|10|11|И сказал он мне: "Даниил, муж желаний! вникни в слова, которые я скажу тебе, и стань прямо на ноги твои; ибо к тебе я послан ныне". Когда он сказал мне эти слова, я встал с трепетом.
DAN|10|12|Но он сказал мне: "не бойся, Даниил; с первого дня, как ты расположил сердце твое, чтобы достигнуть разумения и смирить тебя пред Богом твоим, слова твои услышаны, и я пришел бы по словам твоим.
DAN|10|13|Но князь царства Персидского стоял против меня двадцать один день; но вот, Михаил, один из первых князей, пришел помочь мне, и я остался там при царях Персидских.
DAN|10|14|А теперь я пришел возвестить тебе, что будет с народом твоим в последние времена, так как видение относится к отдаленным дням".
DAN|10|15|Когда он говорил мне такие слова, я припал лицем моим к земле и онемел.
DAN|10|16|Но вот, некто, по виду похожий на сынов человеческих, коснулся уст моих, и я открыл уста мои, стал говорить и сказал стоящему передо мною: "господин мой! от этого видения внутренности мои повернулись во мне, и не стало во мне силы.
DAN|10|17|И как может говорить раб такого господина моего с таким господином моим? ибо во мне нет силы, и дыхание замерло во мне".
DAN|10|18|Тогда снова прикоснулся ко мне тот человеческий облик и укрепил меня
DAN|10|19|и сказал: "не бойся, муж желаний! мир тебе; мужайся, мужайся!" И когда он говорил со мною, я укрепился и сказал: "говори, господин мой; ибо ты укрепил меня".
DAN|10|20|И он сказал: "знаешь ли, для чего я пришел к тебе? Теперь я возвращусь, чтобы бороться с князем Персидским; а когда я выйду, то вот, придет князь Греции.
DAN|10|21|Впрочем я возвещу тебе, что начертано в истинном писании; и нет никого, кто поддерживал бы меня в том, кроме Михаила, князя вашего.
DAN|11|1|Итак я с первого года Дария Мидянина стал ему подпорою и подкреплением.
DAN|11|2|Теперь возвещу тебе истину: вот, еще три царя восстанут в Персии; потом четвертый превзойдет всех великим богатством, и когда усилится богатством своим, то поднимет всех против царства Греческого.
DAN|11|3|И восстанет царь могущественный, который будет владычествовать с великою властью, и будет действовать по своей воле.
DAN|11|4|Но когда он восстанет, царство его разрушится и разделится по четырем ветрам небесным, и не к его потомкам перейдет, и не с тою властью, с какою он владычествовал; ибо раздробится царство его и достанется другим, кроме этих.
DAN|11|5|И усилится южный царь и один из князей его пересилит его и будет владычествовать, и велико будет владычество его.
DAN|11|6|Но через несколько лет они сблизятся, и дочь южного царя придет к царю северному, чтобы установить правильные отношения между ними; но она не удержит силы в руках своих, не устоит и род ее, но преданы будут как она, так и сопровождавшие ее, и рожденный ею, и помогавшие ей в те времена.
DAN|11|7|Но восстанет отрасль от корня ее, придет к войску и войдет в укрепления царя северного, и будет действовать в них, и усилится.
DAN|11|8|Даже и богов их, истуканы их с драгоценными сосудами их, серебряными и золотыми, увезет в плен в Египет и на несколько лет будет стоять выше царя северного.
DAN|11|9|Хотя этот и сделает нашествие на царство южного царя, но возвратится в свою землю.
DAN|11|10|Потом вооружатся сыновья его и соберут многочисленное войско, и один из них быстро пойдет, наводнит и пройдет, и потом, возвращаясь, будет сражаться с ним до укреплений его.
DAN|11|11|И раздражится южный царь, и выступит, сразится с ним, с царем северным, и выставит большое войско, и предано будет войско в руки его.
DAN|11|12|И ободрится войско, и сердце [царя] вознесется; он низложит многие тысячи, но от этого не будет сильнее.
DAN|11|13|Ибо царь северный возвратится и выставит войско больше прежнего, и через несколько лет быстро придет с огромным войском и большим богатством.
DAN|11|14|В те времена многие восстанут против южного царя, и мятежные из сынов твоего народа поднимутся, чтобы исполнилось видение, и падут.
DAN|11|15|И придет царь северный, устроит вал и овладеет укрепленным городом, и не устоят мышцы юга, ни отборное войско его; недостанет силы противостоять.
DAN|11|16|И кто выйдет к нему, будет действовать по воле его, и никто не устоит перед ним; и на славной земле поставит стан свой, и она пострадает от руки его.
DAN|11|17|И вознамерится войти со всеми силами царства своего, и праведные с ним, и совершит это; и дочь жен отдаст ему, на погибель ее, но этот замысел не состоится, и ему не будет пользы из того.
DAN|11|18|Потом обратит лице свое к островам и овладеет многими; но некий вождь прекратит нанесенный им позор и даже свой позор обратит на него.
DAN|11|19|Затем он обратит лице свое на крепости своей земли; но споткнется, падет и не станет его.
DAN|11|20|На место его восстанет некий, который пошлет сборщика податей, пройти по царству славы; но и он после немногих дней погибнет, и не от возмущения и не в сражении.
DAN|11|21|И восстанет на место его презренный, и не воздадут ему царских почестей, но он придет без шума и лестью овладеет царством.
DAN|11|22|И всепотопляющие полчища будут потоплены и сокрушены им, даже и сам вождь завета.
DAN|11|23|Ибо после того, как он вступит в союз с ним, он будет действовать обманом, и взойдет, и одержит верх с малым народом.
DAN|11|24|Он войдет в мирные и плодоносные страны, и совершит то, чего не делали отцы его и отцы отцов его; добычу, награбленное имущество и богатство будет расточать своим и на крепости будет иметь замыслы свои, но только до времени.
DAN|11|25|Потом возбудит силы свои и дух свой с многочисленным войском против царя южного, и южный царь выступит на войну с великим и еще более сильным войском, но не устоит, потому что будет против него коварство.
DAN|11|26|Даже участники трапезы его погубят его, и войско его разольется, и падет много убитых.
DAN|11|27|У обоих царей сих на сердце будет коварство, и за одним столом будут говорить ложь, но успеха не будет, потому что конец еще отложен до времени.
DAN|11|28|И отправится он в землю свою с великим богатством и враждебным намерением против святаго завета, и он исполнит его, и возвратится в свою землю.
DAN|11|29|В назначенное время опять пойдет он на юг; но последний [поход] не такой будет, как прежний,
DAN|11|30|ибо в одно время с ним придут корабли Киттимские; и он упадет духом, и возвратится, и озлобится на святый завет, и исполнит свое намерение, и опять войдет в соглашение с отступниками от святаго завета.
DAN|11|31|И поставлена будет им часть войска, которая осквернит святилище могущества, и прекратит ежедневную жертву, и поставит мерзость запустения.
DAN|11|32|Поступающих нечестиво против завета он привлечет к себе лестью; но люди, чтущие своего Бога, усилятся и будут действовать.
DAN|11|33|И разумные из народа вразумят многих, хотя будут несколько времени страдать от меча и огня, от плена и грабежа;
DAN|11|34|и во время страдания своего будут иметь некоторую помощь, и многие присоединятся к ним, но притворно.
DAN|11|35|Пострадают некоторые и из разумных для испытания их, очищения и для убеления к последнему времени; ибо есть еще время до срока.
DAN|11|36|И будет поступать царь тот по своему произволу, и вознесется и возвеличится выше всякого божества, и о Боге богов станет говорить хульное и будет иметь успех, доколе не совершится гнев: ибо, что предопределено, то исполнится.
DAN|11|37|И о богах отцов своих он не помыслит, и ни желания жен, ни даже божества никакого не уважит; ибо возвеличит себя выше всех.
DAN|11|38|Но богу крепостей на месте его будет он воздавать честь, и этого бога, которого не знали отцы его, он будет чествовать золотом и серебром, и дорогими камнями, и разными драгоценностями,
DAN|11|39|и устроит твердую крепость с чужим богом: которые признают его, тем увеличит почести и даст власть над многими, и землю раздаст в награду.
DAN|11|40|Под конец же времени сразится с ним царь южный, и царь северный устремится как буря на него с колесницами, всадниками и многочисленными кораблями, и нападет на области, наводнит их, и пройдет через них.
DAN|11|41|И войдет он в прекраснейшую из земель, и многие области пострадают и спасутся от руки его только Едом, Моав и большая часть сынов Аммоновых.
DAN|11|42|И прострет руку свою на разные страны; не спасется и земля Египетская.
DAN|11|43|И завладеет он сокровищами золота и серебра и разными драгоценностями Египта; Ливийцы и Ефиопляне последуют за ним.
DAN|11|44|Но слухи с востока и севера встревожат его, и выйдет он в величайшей ярости, чтобы истреблять и губить многих,
DAN|11|45|и раскинет он царские шатры свои между морем и горою преславного святилища; но придет к своему концу, и никто не поможет ему.
DAN|12|1|И восстанет в то время Михаил, князь великий, стоящий за сынов народа твоего; и наступит время тяжкое, какого не бывало с тех пор, как существуют люди, до сего времени; но спасутся в это время из народа твоего все, которые найдены будут записанными в книге.
DAN|12|2|И многие из спящих в прахе земли пробудятся, одни для жизни вечной, другие на вечное поругание и посрамление.
DAN|12|3|И разумные будут сиять, как светила на тверди, и обратившие многих к правде – как звезды, вовеки, навсегда.
DAN|12|4|А ты, Даниил, сокрой слова сии и запечатай книгу сию до последнего времени; многие прочитают ее, и умножится ведение".
DAN|12|5|Тогда я, Даниил, посмотрел, и вот, стоят двое других, один на этом берегу реки, другой на том берегу реки.
DAN|12|6|И [один] сказал мужу в льняной одежде, который стоял над водами реки: "когда будет конец этих чудных происшествий?"
DAN|12|7|И слышал я, как муж в льняной одежде, находившийся над водами реки, подняв правую и левую руку к небу, клялся Живущим вовеки, что к концу времени и времен и полувремени, и по совершенном низложении силы народа святого, все это совершится.
DAN|12|8|Я слышал это, но не понял, и потому сказал: "господин мой! что же после этого будет?"
DAN|12|9|И отвечал он: "иди, Даниил; ибо сокрыты и запечатаны слова сии до последнего времени.
DAN|12|10|Многие очистятся, убелятся и переплавлены будут [в искушении]; нечестивые же будут поступать нечестиво, и не уразумеет сего никто из нечестивых, а мудрые уразумеют.
DAN|12|11|Со времени прекращения ежедневной жертвы и поставления мерзости запустения пройдет тысяча двести девяносто дней.
DAN|12|12|Блажен, кто ожидает и достигнет тысячи трехсот тридцати пяти дней.
DAN|12|13|А ты иди к твоему концу и упокоишься, и восстанешь для получения твоего жребия в конце дней".
