ESTH|1|1|Now it came to pass in the days of Ahasuerus, (this is Ahasuerus which reigned, from India even unto Ethiopia, over an hundred and seven and twenty provinces:)
ESTH|1|2|That in those days, when the king Ahasuerus sat on the throne of his kingdom, which was in Shushan the palace,
ESTH|1|3|In the third year of his reign, he made a feast unto all his princes and his servants; the power of Persia and Media, the nobles and princes of the provinces, being before him:
ESTH|1|4|When he shewed the riches of his glorious kingdom and the honour of his excellent majesty many days, even an hundred and fourscore days.
ESTH|1|5|And when these days were expired, the king made a feast unto all the people that were present in Shushan the palace, both unto great and small, seven days, in the court of the garden of the king's palace;
ESTH|1|6|Where were white, green, and blue, hangings, fastened with cords of fine linen and purple to silver rings and pillars of marble: the beds were of gold and silver, upon a pavement of red, and blue, and white, and black, marble.
ESTH|1|7|And they gave them drink in vessels of gold, (the vessels being diverse one from another,) and royal wine in abundance, according to the state of the king.
ESTH|1|8|And the drinking was according to the law; none did compel: for so the king had appointed to all the officers of his house, that they should do according to every man's pleasure.
ESTH|1|9|Also Vashti the queen made a feast for the women in the royal house which belonged to king Ahasuerus.
ESTH|1|10|On the seventh day, when the heart of the king was merry with wine, he commanded Mehuman, Biztha, Harbona, Bigtha, and Abagtha, Zethar, and Carcas, the seven chamberlains that served in the presence of Ahasuerus the king,
ESTH|1|11|To bring Vashti the queen before the king with the crown royal, to shew the people and the princes her beauty: for she was fair to look on.
ESTH|1|12|But the queen Vashti refused to come at the king's commandment by his chamberlains: therefore was the king very wroth, and his anger burned in him.
ESTH|1|13|Then the king said to the wise men, which knew the times, (for so was the king's manner toward all that knew law and judgment:
ESTH|1|14|And the next unto him was Carshena, Shethar, Admatha, Tarshish, Meres, Marsena, and Memucan, the seven princes of Persia and Media, which saw the king's face, and which sat the first in the kingdom;)
ESTH|1|15|What shall we do unto the queen Vashti according to law, because she hath not performed the commandment of the king Ahasuerus by the chamberlains?
ESTH|1|16|And Memucan answered before the king and the princes, Vashti the queen hath not done wrong to the king only, but also to all the princes, and to all the people that are in all the provinces of the king Ahasuerus.
ESTH|1|17|For this deed of the queen shall come abroad unto all women, so that they shall despise their husbands in their eyes, when it shall be reported, The king Ahasuerus commanded Vashti the queen to be brought in before him, but she came not.
ESTH|1|18|Likewise shall the ladies of Persia and Media say this day unto all the king's princes, which have heard of the deed of the queen. Thus shall there arise too much contempt and wrath.
ESTH|1|19|If it please the king, let there go a royal commandment from him, and let it be written among the laws of the Persians and the Medes, that it be not altered, That Vashti come no more before king Ahasuerus; and let the king give her royal estate unto another that is better than she.
ESTH|1|20|And when the king's decree which he shall make shall be published throughout all his empire, (for it is great,) all the wives shall give to their husbands honour, both to great and small.
ESTH|1|21|And the saying pleased the king and the princes; and the king did according to the word of Memucan:
ESTH|1|22|For he sent letters into all the king's provinces, into every province according to the writing thereof, and to every people after their language, that every man should bear rule in his own house, and that it should be published according to the language of every people.
ESTH|2|1|After these things, when the wrath of king Ahasuerus was appeased, he remembered Vashti, and what she had done, and what was decreed against her.
ESTH|2|2|Then said the king's servants that ministered unto him, Let there be fair young virgins sought for the king:
ESTH|2|3|And let the king appoint officers in all the provinces of his kingdom, that they may gather together all the fair young virgins unto Shushan the palace, to the house of the women, unto the custody of Hege the king's chamberlain, keeper of the women; and let their things for purification be given them:
ESTH|2|4|And let the maiden which pleaseth the king be queen instead of Vashti. And the thing pleased the king; and he did so.
ESTH|2|5|Now in Shushan the palace there was a certain Jew, whose name was Mordecai, the son of Jair, the son of Shimei, the son of Kish, a Benjamite;
ESTH|2|6|Who had been carried away from Jerusalem with the captivity which had been carried away with Jeconiah king of Judah, whom Nebuchadnezzar the king of Babylon had carried away.
ESTH|2|7|And he brought up Hadassah, that is, Esther, his uncle's daughter: for she had neither father nor mother, and the maid was fair and beautiful; whom Mordecai, when her father and mother were dead, took for his own daughter.
ESTH|2|8|So it came to pass, when the king's commandment and his decree was heard, and when many maidens were gathered together unto Shushan the palace, to the custody of Hegai, that Esther was brought also unto the king's house, to the custody of Hegai, keeper of the women.
ESTH|2|9|And the maiden pleased him, and she obtained kindness of him; and he speedily gave her her things for purification, with such things as belonged to her, and seven maidens, which were meet to be given her, out of the king's house: and he preferred her and her maids unto the best place of the house of the women.
ESTH|2|10|Esther had not shewed her people nor her kindred: for Mordecai had charged her that she should not shew it.
ESTH|2|11|And Mordecai walked every day before the court of the women's house, to know how Esther did, and what should become of her.
ESTH|2|12|Now when every maid's turn was come to go in to king Ahasuerus, after that she had been twelve months, according to the manner of the women, (for so were the days of their purifications accomplished, to wit, six months with oil of myrrh, and six months with sweet odours, and with other things for the purifying of the women;)
ESTH|2|13|Then thus came every maiden unto the king; whatsoever she desired was given her to go with her out of the house of the women unto the king's house.
ESTH|2|14|In the evening she went, and on the morrow she returned into the second house of the women, to the custody of Shaashgaz, the king's chamberlain, which kept the concubines: she came in unto the king no more, except the king delighted in her, and that she were called by name.
ESTH|2|15|Now when the turn of Esther, the daughter of Abihail the uncle of Mordecai, who had taken her for his daughter, was come to go in unto the king, she required nothing but what Hegai the king's chamberlain, the keeper of the women, appointed. And Esther obtained favour in the sight of all them that looked upon her.
ESTH|2|16|So Esther was taken unto king Ahasuerus into his house royal in the tenth month, which is the month Tebeth, in the seventh year of his reign.
ESTH|2|17|And the king loved Esther above all the women, and she obtained grace and favour in his sight more than all the virgins; so that he set the royal crown upon her head, and made her queen instead of Vashti.
ESTH|2|18|Then the king made a great feast unto all his princes and his servants, even Esther's feast; and he made a release to the provinces, and gave gifts, according to the state of the king.
ESTH|2|19|And when the virgins were gathered together the second time, then Mordecai sat in the king's gate.
ESTH|2|20|Esther had not yet shewed her kindred nor her people; as Mordecai had charged her: for Esther did the commandment of Mordecai, like as when she was brought up with him.
ESTH|2|21|In those days, while Mordecai sat in the king's gate, two of the king's chamberlains, Bigthan and Teresh, of those which kept the door, were wroth, and sought to lay hands on the king Ahasuerus.
ESTH|2|22|And the thing was known to Mordecai, who told it unto Esther the queen; and Esther certified the king thereof in Mordecai's name.
ESTH|2|23|And when inquisition was made of the matter, it was found out; therefore they were both hanged on a tree: and it was written in the book of the chronicles before the king.
ESTH|3|1|After these things did king Ahasuerus promote Haman the son of Hammedatha the Agagite, and advanced him, and set his seat above all the princes that were with him.
ESTH|3|2|And all the king's servants, that were in the king's gate, bowed, and reverenced Haman: for the king had so commanded concerning him. But Mordecai bowed not, nor did him reverence.
ESTH|3|3|Then the king's servants, which were in the king's gate, said unto Mordecai, Why transgressest thou the king's commandment?
ESTH|3|4|Now it came to pass, when they spake daily unto him, and he hearkened not unto them, that they told Haman, to see whether Mordecai's matters would stand: for he had told them that he was a Jew.
ESTH|3|5|And when Haman saw that Mordecai bowed not, nor did him reverence, then was Haman full of wrath.
ESTH|3|6|And he thought scorn to lay hands on Mordecai alone; for they had shewed him the people of Mordecai: wherefore Haman sought to destroy all the Jews that were throughout the whole kingdom of Ahasuerus, even the people of Mordecai.
ESTH|3|7|In the first month, that is, the month Nisan, in the twelfth year of king Ahasuerus, they cast Pur, that is, the lot, before Haman from day to day, and from month to month, to the twelfth month, that is, the month Adar.
ESTH|3|8|And Haman said unto king Ahasuerus, There is a certain people scattered abroad and dispersed among the people in all the provinces of thy kingdom; and their laws are diverse from all people; neither keep they the king's laws: therefore it is not for the king's profit to suffer them.
ESTH|3|9|If it please the king, let it be written that they may be destroyed: and I will pay ten thousand talents of silver to the hands of those that have the charge of the business, to bring it into the king's treasuries.
ESTH|3|10|And the king took his ring from his hand, and gave it unto Haman the son of Hammedatha the Agagite, the Jews' enemy.
ESTH|3|11|And the king said unto Haman, The silver is given to thee, the people also, to do with them as it seemeth good to thee.
ESTH|3|12|Then were the king's scribes called on the thirteenth day of the first month, and there was written according to all that Haman had commanded unto the king's lieutenants, and to the governors that were over every province, and to the rulers of every people of every province according to the writing thereof, and to every people after their language; in the name of king Ahasuerus was it written, and sealed with the king's ring.
ESTH|3|13|And the letters were sent by posts into all the king's provinces, to destroy, to kill, and to cause to perish, all Jews, both young and old, little children and women, in one day, even upon the thirteenth day of the twelfth month, which is the month Adar, and to take the spoil of them for a prey.
ESTH|3|14|The copy of the writing for a commandment to be given in every province was published unto all people, that they should be ready against that day.
ESTH|3|15|The posts went out, being hastened by the king's commandment, and the decree was given in Shushan the palace. And the king and Haman sat down to drink; but the city Shushan was perplexed.
ESTH|4|1|When Mordecai perceived all that was done, Mordecai rent his clothes, and put on sackcloth with ashes, and went out into the midst of the city, and cried with a loud and a bitter cry;
ESTH|4|2|And came even before the king's gate: for none might enter into the king's gate clothed with sackcloth.
ESTH|4|3|And in every province, whithersoever the king's commandment and his decree came, there was great mourning among the Jews, and fasting, and weeping, and wailing; and many lay in sackcloth and ashes.
ESTH|4|4|So Esther's maids and her chamberlains came and told it her. Then was the queen exceedingly grieved; and she sent raiment to clothe Mordecai, and to take away his sackcloth from him: but he received it not.
ESTH|4|5|Then called Esther for Hatach, one of the king's chamberlains, whom he had appointed to attend upon her, and gave him a commandment to Mordecai, to know what it was, and why it was.
ESTH|4|6|So Hatach went forth to Mordecai unto the street of the city, which was before the king's gate.
ESTH|4|7|And Mordecai told him of all that had happened unto him, and of the sum of the money that Haman had promised to pay to the king's treasuries for the Jews, to destroy them.
ESTH|4|8|Also he gave him the copy of the writing of the decree that was given at Shushan to destroy them, to shew it unto Esther, and to declare it unto her, and to charge her that she should go in unto the king, to make supplication unto him, and to make request before him for her people.
ESTH|4|9|And Hatach came and told Esther the words of Mordecai.
ESTH|4|10|Again Esther spake unto Hatach, and gave him commandment unto Mordecai;
ESTH|4|11|All the king's servants, and the people of the king's provinces, do know, that whosoever, whether man or women, shall come unto the king into the inner court, who is not called, there is one law of his to put him to death, except such to whom the king shall hold out the golden sceptre, that he may live: but I have not been called to come in unto the king these thirty days.
ESTH|4|12|And they told to Mordecai Esther's words.
ESTH|4|13|Then Mordecai commanded to answer Esther, Think not with thyself that thou shalt escape in the king's house, more than all the Jews.
ESTH|4|14|For if thou altogether holdest thy peace at this time, then shall there enlargement and deliverance arise to the Jews from another place; but thou and thy father's house shall be destroyed: and who knoweth whether thou art come to the kingdom for such a time as this?
ESTH|4|15|Then Esther bade them return Mordecai this answer,
ESTH|4|16|Go, gather together all the Jews that are present in Shushan, and fast ye for me, and neither eat nor drink three days, night or day: I also and my maidens will fast likewise; and so will I go in unto the king, which is not according to the law: and if I perish, I perish.
ESTH|4|17|So Mordecai went his way, and did according to all that Esther had commanded him.
ESTH|5|1|Now it came to pass on the third day, that Esther put on her royal apparel, and stood in the inner court of the king's house, over against the king's house: and the king sat upon his royal throne in the royal house, over against the gate of the house.
ESTH|5|2|And it was so, when the king saw Esther the queen standing in the court, that she obtained favour in his sight: and the king held out to Esther the golden sceptre that was in his hand. So Esther drew near, and touched the top of the sceptre.
ESTH|5|3|Then said the king unto her, What wilt thou, queen Esther? and what is thy request? it shall be even given thee to the half of the kingdom.
ESTH|5|4|And Esther answered, If it seem good unto the king, let the king and Haman come this day unto the banquet that I have prepared for him.
ESTH|5|5|Then the king said, Cause Haman to make haste, that he may do as Esther hath said. So the king and Haman came to the banquet that Esther had prepared.
ESTH|5|6|And the king said unto Esther at the banquet of wine, What is thy petition? and it shall be granted thee: and what is thy request? even to the half of the kingdom it shall be performed.
ESTH|5|7|Then answered Esther, and said, My petition and my request is;
ESTH|5|8|If I have found favour in the sight of the king, and if it please the king to grant my petition, and to perform my request, let the king and Haman come to the banquet that I shall prepare for them, and I will do to morrow as the king hath said.
ESTH|5|9|Then went Haman forth that day joyful and with a glad heart: but when Haman saw Mordecai in the king's gate, that he stood not up, nor moved for him, he was full of indignation against Mordecai.
ESTH|5|10|Nevertheless Haman refrained himself: and when he came home, he sent and called for his friends, and Zeresh his wife.
ESTH|5|11|And Haman told them of the glory of his riches, and the multitude of his children, and all the things wherein the king had promoted him, and how he had advanced him above the princes and servants of the king.
ESTH|5|12|Haman said moreover, Yea, Esther the queen did let no man come in with the king unto the banquet that she had prepared but myself; and to morrow am I invited unto her also with the king.
ESTH|5|13|Yet all this availeth me nothing, so long as I see Mordecai the Jew sitting at the king's gate.
ESTH|5|14|Then said Zeresh his wife and all his friends unto him, Let a gallows be made of fifty cubits high, and to morrow speak thou unto the king that Mordecai may be hanged thereon: then go thou in merrily with the king unto the banquet. And the thing pleased Haman; and he caused the gallows to be made.
ESTH|6|1|On that night could not the king sleep, and he commanded to bring the book of records of the chronicles; and they were read before the king.
ESTH|6|2|And it was found written, that Mordecai had told of Bigthana and Teresh, two of the king's chamberlains, the keepers of the door, who sought to lay hand on the king Ahasuerus.
ESTH|6|3|And the king said, What honour and dignity hath been done to Mordecai for this? Then said the king's servants that ministered unto him, There is nothing done for him.
ESTH|6|4|And the king said, Who is in the court? Now Haman was come into the outward court of the king's house, to speak unto the king to hang Mordecai on the gallows that he had prepared for him.
ESTH|6|5|And the king's servants said unto him, Behold, Haman standeth in the court. And the king said, Let him come in.
ESTH|6|6|So Haman came in. And the king said unto him, What shall be done unto the man whom the king delighteth to honour? Now Haman thought in his heart, To whom would the king delight to do honour more than to myself?
ESTH|6|7|And Haman answered the king, For the man whom the king delighteth to honour,
ESTH|6|8|Let the royal apparel be brought which the king useth to wear, and the horse that the king rideth upon, and the crown royal which is set upon his head:
ESTH|6|9|And let this apparel and horse be delivered to the hand of one of the king's most noble princes, that they may array the man withal whom the king delighteth to honour, and bring him on horseback through the street of the city, and proclaim before him, Thus shall it be done to the man whom the king delighteth to honour.
ESTH|6|10|Then the king said to Haman, Make haste, and take the apparel and the horse, as thou hast said, and do even so to Mordecai the Jew, that sitteth at the king's gate: let nothing fail of all that thou hast spoken.
ESTH|6|11|Then took Haman the apparel and the horse, and arrayed Mordecai, and brought him on horseback through the street of the city, and proclaimed before him, Thus shall it be done unto the man whom the king delighteth to honour.
ESTH|6|12|And Mordecai came again to the king's gate. But Haman hasted to his house mourning, and having his head covered.
ESTH|6|13|And Haman told Zeresh his wife and all his friends every thing that had befallen him. Then said his wise men and Zeresh his wife unto him, If Mordecai be of the seed of the Jews, before whom thou hast begun to fall, thou shalt not prevail against him, but shalt surely fall before him.
ESTH|6|14|And while they were yet talking with him, came the king's chamberlains, and hasted to bring Haman unto the banquet that Esther had prepared.
ESTH|7|1|So the king and Haman came to banquet with Esther the queen.
ESTH|7|2|And the king said again unto Esther on the second day at the banquet of wine, What is thy petition, queen Esther? and it shall be granted thee: and what is thy request? and it shall be performed, even to the half of the kingdom.
ESTH|7|3|Then Esther the queen answered and said, If I have found favour in thy sight, O king, and if it please the king, let my life be given me at my petition, and my people at my request:
ESTH|7|4|For we are sold, I and my people, to be destroyed, to be slain, and to perish. But if we had been sold for bondmen and bondwomen, I had held my tongue, although the enemy could not countervail the king's damage.
ESTH|7|5|Then the king Ahasuerus answered and said unto Esther the queen, Who is he, and where is he, that durst presume in his heart to do so?
ESTH|7|6|And Esther said, The adversary and enemy is this wicked Haman. Then Haman was afraid before the king and the queen.
ESTH|7|7|And the king arising from the banquet of wine in his wrath went into the palace garden: and Haman stood up to make request for his life to Esther the queen; for he saw that there was evil determined against him by the king.
ESTH|7|8|Then the king returned out of the palace garden into the place of the banquet of wine; and Haman was fallen upon the bed whereon Esther was. Then said the king, Will he force the queen also before me in the house? As the word went out of king's mouth, they covered Haman's face.
ESTH|7|9|And Harbonah, one of the chamberlains, said before the king, Behold also, the gallows fifty cubits high, which Haman had made for Mordecai, who spoken good for the king, standeth in the house of Haman. Then the king said, Hang him thereon.
ESTH|7|10|So they hanged Haman on the gallows that he had prepared for Mordecai. Then was the king's wrath pacified.
ESTH|8|1|On that day did the king Ahasuerus give the house of Haman the Jews' enemy unto Esther the queen. And Mordecai came before the king; for Esther had told what he was unto her.
ESTH|8|2|And the king took off his ring, which he had taken from Haman, and gave it unto Mordecai. And Esther set Mordecai over the house of Haman.
ESTH|8|3|And Esther spake yet again before the king, and fell down at his feet, and besought him with tears to put away the mischief of Haman the Agagite, and his device that he had devised against the Jews.
ESTH|8|4|Then the king held out the golden sceptre toward Esther. So Esther arose, and stood before the king,
ESTH|8|5|And said, If it please the king, and if I have favour in his sight, and the thing seem right before the king, and I be pleasing in his eyes, let it be written to reverse the letters devised by Haman the son of Hammedatha the Agagite, which he wrote to destroy the Jews which are in all the king's provinces:
ESTH|8|6|For how can I endure to see the evil that shall come unto my people? or how can I endure to see the destruction of my kindred?
ESTH|8|7|Then the king Ahasuerus said unto Esther the queen and to Mordecai the Jew, Behold, I have given Esther the house of Haman, and him they have hanged upon the gallows, because he laid his hand upon the Jews.
ESTH|8|8|Write ye also for the Jews, as it liketh you, in the king's name, and seal it with the king's ring: for the writing which is written in the king's name, and sealed with the king's ring, may no man reverse.
ESTH|8|9|Then were the king's scribes called at that time in the third month, that is, the month Sivan, on the three and twentieth day thereof; and it was written according to all that Mordecai commanded unto the Jews, and to the lieutenants, and the deputies and rulers of the provinces which are from India unto Ethiopia, an hundred twenty and seven provinces, unto every province according to the writing thereof, and unto every people after their language, and to the Jews according to their writing, and according to their language.
ESTH|8|10|And he wrote in the king Ahasuerus' name, and sealed it with the king's ring, and sent letters by posts on horseback, and riders on mules, camels, and young dromedaries:
ESTH|8|11|Wherein the king granted the Jews which were in every city to gather themselves together, and to stand for their life, to destroy, to slay and to cause to perish, all the power of the people and province that would assault them, both little ones and women, and to take the spoil of them for a prey,
ESTH|8|12|Upon one day in all the provinces of king Ahasuerus, namely, upon the thirteenth day of the twelfth month, which is the month Adar.
ESTH|8|13|The copy of the writing for a commandment to be given in every province was published unto all people, and that the Jews should be ready against that day to avenge themselves on their enemies.
ESTH|8|14|So the posts that rode upon mules and camels went out, being hastened and pressed on by the king's commandment. And the decree was given at Shushan the palace.
ESTH|8|15|And Mordecai went out from the presence of the king in royal apparel of blue and white, and with a great crown of gold, and with a garment of fine linen and purple: and the city of Shushan rejoiced and was glad.
ESTH|8|16|The Jews had light, and gladness, and joy, and honour.
ESTH|8|17|And in every province, and in every city, whithersoever the king's commandment and his decree came, the Jews had joy and gladness, a feast and a good day. And many of the people of the land became Jews; for the fear of the Jews fell upon them.
ESTH|9|1|Now in the twelfth month, that is, the month Adar, on the thirteenth day of the same, when the king's commandment and his decree drew near to be put in execution, in the day that the enemies of the Jews hoped to have power over them, (though it was turned to the contrary, that the Jews had rule over them that hated them;)
ESTH|9|2|The Jews gathered themselves together in their cities throughout all the provinces of the king Ahasuerus, to lay hand on such as sought their hurt: and no man could withstand them; for the fear of them fell upon all people.
ESTH|9|3|And all the rulers of the provinces, and the lieutenants, and the deputies, and officers of the king, helped the Jews; because the fear of Mordecai fell upon them.
ESTH|9|4|For Mordecai was great in the king's house, and his fame went out throughout all the provinces: for this man Mordecai waxed greater and greater.
ESTH|9|5|Thus the Jews smote all their enemies with the stroke of the sword, and slaughter, and destruction, and did what they would unto those that hated them.
ESTH|9|6|And in Shushan the palace the Jews slew and destroyed five hundred men.
ESTH|9|7|And Parshandatha, and Dalphon, and Aspatha,
ESTH|9|8|And Poratha, and Adalia, and Aridatha,
ESTH|9|9|And Parmashta, and Arisai, and Aridai, and Vajezatha,
ESTH|9|10|The ten sons of Haman the son of Hammedatha, the enemy of the Jews, slew they; but on the spoil laid they not their hand.
ESTH|9|11|On that day the number of those that were slain in Shushan the palace was brought before the king.
ESTH|9|12|And the king said unto Esther the queen, The Jews have slain and destroyed five hundred men in Shushan the palace, and the ten sons of Haman; what have they done in the rest of the king's provinces? now what is thy petition? and it shall be granted thee: or what is thy request further? and it shall be done.
ESTH|9|13|Then said Esther, If it please the king, let it be granted to the Jews which are in Shushan to do to morrow also according unto this day's decree, and let Haman's ten sons be hanged upon the gallows.
ESTH|9|14|And the king commanded it so to be done: and the decree was given at Shushan; and they hanged Haman's ten sons.
ESTH|9|15|For the Jews that were in Shushan gathered themselves together on the fourteenth day also of the month Adar, and slew three hundred men at Shushan; but on the prey they laid not their hand.
ESTH|9|16|But the other Jews that were in the king's provinces gathered themselves together, and stood for their lives, and had rest from their enemies, and slew of their foes seventy and five thousand, but they laid not their hands on the prey,
ESTH|9|17|On the thirteenth day of the month Adar; and on the fourteenth day of the same rested they, and made it a day of feasting and gladness.
ESTH|9|18|But the Jews that were at Shushan assembled together on the thirteenth day thereof, and on the fourteenth thereof; and on the fifteenth day of the same they rested, and made it a day of feasting and gladness.
ESTH|9|19|Therefore the Jews of the villages, that dwelt in the unwalled towns, made the fourteenth day of the month Adar a day of gladness and feasting, and a good day, and of sending portions one to another.
ESTH|9|20|And Mordecai wrote these things, and sent letters unto all the Jews that were in all the provinces of the king Ahasuerus, both nigh and far,
ESTH|9|21|To stablish this among them, that they should keep the fourteenth day of the month Adar, and the fifteenth day of the same, yearly,
ESTH|9|22|As the days wherein the Jews rested from their enemies, and the month which was turned unto them from sorrow to joy, and from mourning into a good day: that they should make them days of feasting and joy, and of sending portions one to another, and gifts to the poor.
ESTH|9|23|And the Jews undertook to do as they had begun, and as Mordecai had written unto them;
ESTH|9|24|Because Haman the son of Hammedatha, the Agagite, the enemy of all the Jews, had devised against the Jews to destroy them, and had cast Pur, that is, the lot, to consume them, and to destroy them;
ESTH|9|25|But when Esther came before the king, he commanded by letters that his wicked device, which he devised against the Jews, should return upon his own head, and that he and his sons should be hanged on the gallows.
ESTH|9|26|Wherefore they called these days Purim after the name of Pur. Therefore for all the words of this letter, and of that which they had seen concerning this matter, and which had come unto them,
ESTH|9|27|The Jews ordained, and took upon them, and upon their seed, and upon all such as joined themselves unto them, so as it should not fail, that they would keep these two days according to their writing, and according to their appointed time every year;
ESTH|9|28|And that these days should be remembered and kept throughout every generation, every family, every province, and every city; and that these days of Purim should not fail from among the Jews, nor the memorial of them perish from their seed.
ESTH|9|29|Then Esther the queen, the daughter of Abihail, and Mordecai the Jew, wrote with all authority, to confirm this second letter of Purim.
ESTH|9|30|And he sent the letters unto all the Jews, to the hundred twenty and seven provinces of the kingdom of Ahasuerus, with words of peace and truth,
ESTH|9|31|To confirm these days of Purim in their times appointed, according as Mordecai the Jew and Esther the queen had enjoined them, and as they had decreed for themselves and for their seed, the matters of the fastings and their cry.
ESTH|9|32|And the decree of Esther confirmed these matters of Purim; and it was written in the book.
ESTH|10|1|And the king Ahasuerus laid a tribute upon the land, and upon the isles of the sea.
ESTH|10|2|And all the acts of his power and of his might, and the declaration of the greatness of Mordecai, whereunto the king advanced him, are they not written in the book of the chronicles of the kings of Media and Persia?
ESTH|10|3|For Mordecai the Jew was next unto king Ahasuerus, and great among the Jews, and accepted of the multitude of his brethren, seeking the wealth of his people, and speaking peace to all his seed.
