ROM|1|1|Paulus servus Christi Iesu vocatus apostolus segregatus in evangelium Dei
ROM|1|2|quod ante promiserat per prophetas suos in scripturis sanctis
ROM|1|3|de Filio suo qui factus est ex semine David secundum carnem
ROM|1|4|qui praedestinatus est Filius Dei in virtute secundum Spiritum sanctificationis ex resurrectione mortuorum Iesu Christi Domini nostri
ROM|1|5|per quem accepimus gratiam et apostolatum ad oboediendum fidei in omnibus gentibus pro nomine eius
ROM|1|6|in quibus estis et vos vocati Iesu Christi
ROM|1|7|omnibus qui sunt Romae dilectis Dei vocatis sanctis gratia vobis et pax a Deo Patre nostro et Domino Iesu Christo
ROM|1|8|primum quidem gratias ago Deo meo per Iesum Christum pro omnibus vobis quia fides vestra adnuntiatur in universo mundo
ROM|1|9|testis enim mihi est Deus cui servio in spiritu meo in evangelio Filii eius quod sine intermissione memoriam vestri facio
ROM|1|10|semper in orationibus meis obsecrans si quo modo tandem aliquando prosperum iter habeam in voluntate Dei veniendi ad vos
ROM|1|11|desidero enim videre vos ut aliquid inpertiar gratiae vobis spiritalis ad confirmandos vos
ROM|1|12|id est simul consolari in vobis per eam quae invicem est fidem vestram atque meam
ROM|1|13|nolo autem vos ignorare fratres quia saepe proposui venire ad vos et prohibitus sum usque adhuc ut aliquem fructum habeam et in vobis sicut et in ceteris gentibus
ROM|1|14|Graecis ac barbaris sapientibus et insipientibus debitor sum
ROM|1|15|ita quod in me promptum est et vobis qui Romae estis evangelizare
ROM|1|16|non enim erubesco evangelium virtus enim Dei est in salutem omni credenti Iudaeo primum et Graeco
ROM|1|17|iustitia enim Dei in eo revelatur ex fide in fidem sicut scriptum est iustus autem ex fide vivit
ROM|1|18|revelatur enim ira Dei de caelo super omnem impietatem et iniustitiam hominum eorum qui veritatem in iniustitiam detinent
ROM|1|19|quia quod notum est Dei manifestum est in illis Deus enim illis manifestavit
ROM|1|20|invisibilia enim ipsius a creatura mundi per ea quae facta sunt intellecta conspiciuntur sempiterna quoque eius virtus et divinitas ut sint inexcusabiles
ROM|1|21|quia cum cognovissent Deum non sicut Deum glorificaverunt aut gratias egerunt sed evanuerunt in cogitationibus suis et obscuratum est insipiens cor eorum
ROM|1|22|dicentes enim se esse sapientes stulti facti sunt
ROM|1|23|et mutaverunt gloriam incorruptibilis Dei in similitudinem imaginis corruptibilis hominis et volucrum et quadrupedum et serpentium
ROM|1|24|propter quod tradidit illos Deus in desideria cordis eorum in inmunditiam ut contumeliis adficiant corpora sua in semet ipsis
ROM|1|25|qui commutaverunt veritatem Dei in mendacio et coluerunt et servierunt creaturae potius quam creatori qui est benedictus in saecula amen
ROM|1|26|propterea tradidit illos Deus in passiones ignominiae nam feminae eorum inmutaverunt naturalem usum in eum usum qui est contra naturam
ROM|1|27|similiter autem et masculi relicto naturali usu feminae exarserunt in desideriis suis in invicem masculi in masculos turpitudinem operantes et mercedem quam oportuit erroris sui in semet ipsis recipientes
ROM|1|28|et sicut non probaverunt Deum habere in notitia tradidit eos Deus in reprobum sensum ut faciant quae non conveniunt
ROM|1|29|repletos omni iniquitate malitia fornicatione avaritia nequitia plenos invidia homicidio contentione dolo malignitate susurrones
ROM|1|30|detractores Deo odibiles contumeliosos superbos elatos inventores malorum parentibus non oboedientes
ROM|1|31|insipientes inconpositos sine affectione absque foedere sine misericordia
ROM|1|32|qui cum iustitiam Dei cognovissent non intellexerunt quoniam qui talia agunt digni sunt morte non solum ea faciunt sed et consentiunt facientibus
ROM|2|1|propter quod inexcusabilis es o homo omnis qui iudicas in quo enim iudicas alterum te ipsum condemnas eadem enim agis qui iudicas
ROM|2|2|scimus enim quoniam iudicium Dei est secundum veritatem in eos qui talia agunt
ROM|2|3|existimas autem hoc o homo qui iudicas eos qui talia agunt et facis ea quia tu effugies iudicium Dei
ROM|2|4|an divitias bonitatis eius et patientiae et longanimitatis contemnis ignorans quoniam benignitas Dei ad paenitentiam te adducit
ROM|2|5|secundum duritiam autem tuam et inpaenitens cor thesaurizas tibi iram in die irae et revelationis iusti iudicii Dei
ROM|2|6|qui reddet unicuique secundum opera eius
ROM|2|7|his quidem qui secundum patientiam boni operis gloriam et honorem et incorruptionem quaerentibus vitam aeternam
ROM|2|8|his autem qui ex contentione et qui non adquiescunt veritati credunt autem iniquitati ira et indignatio
ROM|2|9|tribulatio et angustia in omnem animam hominis operantis malum Iudaei primum et Graeci
ROM|2|10|gloria autem et honor et pax omni operanti bonum Iudaeo primum et Graeco
ROM|2|11|non est enim personarum acceptio apud Deum
ROM|2|12|quicumque enim sine lege peccaverunt sine lege et peribunt et quicumque in lege peccaverunt per legem iudicabuntur
ROM|2|13|non enim auditores legis iusti sunt apud Deum sed factores legis iustificabuntur
ROM|2|14|cum enim gentes quae legem non habent naturaliter quae legis sunt faciunt eiusmodi legem non habentes ipsi sibi sunt lex
ROM|2|15|qui ostendunt opus legis scriptum in cordibus suis testimonium reddente illis conscientia ipsorum et inter se invicem cogitationum accusantium aut etiam defendentium
ROM|2|16|in die cum iudicabit Deus occulta hominum secundum evangelium meum per Iesum Christum
ROM|2|17|si autem tu Iudaeus cognominaris et requiescis in lege et gloriaris in Deo
ROM|2|18|et nosti voluntatem et probas utiliora instructus per legem
ROM|2|19|confidis te ipsum ducem esse caecorum lumen eorum qui in tenebris sunt
ROM|2|20|eruditorem insipientium magistrum infantium habentem formam scientiae et veritatis in lege
ROM|2|21|qui ergo alium doces te ipsum non doces qui praedicas non furandum furaris
ROM|2|22|qui dicis non moechandum moecharis qui abominaris idola sacrilegium facis
ROM|2|23|qui in lege gloriaris per praevaricationem legis Deum inhonoras
ROM|2|24|nomen enim Dei per vos blasphematur inter gentes sicut scriptum est
ROM|2|25|circumcisio quidem prodest si legem observes si autem praevaricator legis sis circumcisio tua praeputium facta est
ROM|2|26|si igitur praeputium iustitias legis custodiat nonne praeputium illius in circumcisionem reputabitur
ROM|2|27|et iudicabit quod ex natura est praeputium legem consummans te qui per litteram et circumcisionem praevaricator legis es
ROM|2|28|non enim qui in manifesto Iudaeus est neque quae in manifesto in carne circumcisio
ROM|2|29|sed qui in abscondito Iudaeus et circumcisio cordis in spiritu non littera cuius laus non ex hominibus sed ex Deo est
ROM|3|1|quid ergo amplius est Iudaeo aut quae utilitas circumcisionis
ROM|3|2|multum per omnem modum primum quidem quia credita sunt illis eloquia Dei
ROM|3|3|quid enim si quidam illorum non crediderunt numquid incredulitas illorum fidem Dei evacuabit absit
ROM|3|4|est autem Deus verax omnis autem homo mendax sicut scriptum est ut iustificeris in sermonibus tuis et vincas cum iudicaris
ROM|3|5|si autem iniquitas nostra iustitiam Dei commendat quid dicemus numquid iniquus Deus qui infert iram secundum hominem dico
ROM|3|6|absit alioquin quomodo iudicabit Deus mundum
ROM|3|7|si enim veritas Dei in meo mendacio abundavit in gloriam ipsius quid adhuc et ego tamquam peccator iudicor
ROM|3|8|et non sicut blasphemamur et sicut aiunt nos quidam dicere faciamus mala ut veniant bona quorum damnatio iusta est
ROM|3|9|quid igitur praecellimus eos nequaquam causati enim sumus Iudaeos et Graecos omnes sub peccato esse
ROM|3|10|sicut scriptum est quia non est iustus quisquam
ROM|3|11|non est intellegens non est requirens Deum
ROM|3|12|omnes declinaverunt simul inutiles facti sunt non est qui faciat bonum non est usque ad unum
ROM|3|13|sepulchrum patens est guttur eorum linguis suis dolose agebant venenum aspidum sub labiis eorum
ROM|3|14|quorum os maledictione et amaritudine plenum est
ROM|3|15|veloces pedes eorum ad effundendum sanguinem
ROM|3|16|contritio et infelicitas in viis eorum
ROM|3|17|et viam pacis non cognoverunt
ROM|3|18|non est timor Dei ante oculos eorum
ROM|3|19|scimus autem quoniam quaecumque lex loquitur his qui in lege sunt loquitur ut omne os obstruatur et subditus fiat omnis mundus Deo
ROM|3|20|quia ex operibus legis non iustificabitur omnis caro coram illo per legem enim cognitio peccati
ROM|3|21|nunc autem sine lege iustitia Dei manifestata est testificata a lege et prophetis
ROM|3|22|iustitia autem Dei per fidem Iesu Christi super omnes qui credunt non enim est distinctio
ROM|3|23|omnes enim peccaverunt et egent gloriam Dei
ROM|3|24|iustificati gratis per gratiam ipsius per redemptionem quae est in Christo Iesu
ROM|3|25|quem proposuit Deus propitiationem per fidem in sanguine ipsius ad ostensionem iustitiae suae propter remissionem praecedentium delictorum
ROM|3|26|in sustentatione Dei ad ostensionem iustitiae eius in hoc tempore ut sit ipse iustus et iustificans eum qui ex fide est Iesu
ROM|3|27|ubi est ergo gloriatio exclusa est per quam legem factorum non sed per legem fidei
ROM|3|28|arbitramur enim iustificari hominem per fidem sine operibus legis
ROM|3|29|an Iudaeorum Deus tantum nonne et gentium immo et gentium
ROM|3|30|quoniam quidem unus Deus qui iustificabit circumcisionem ex fide et praeputium per fidem
ROM|3|31|legem ergo destruimus per fidem absit sed legem statuimus
ROM|4|1|quid ergo dicemus invenisse Abraham patrem nostrum secundum carnem
ROM|4|2|si enim Abraham ex operibus iustificatus est habet gloriam sed non apud Deum
ROM|4|3|quid enim scriptura dicit credidit Abraham Deo et reputatum est illi ad iustitiam
ROM|4|4|ei autem qui operatur merces non inputatur secundum gratiam sed secundum debitum
ROM|4|5|ei vero qui non operatur credenti autem in eum qui iustificat impium reputatur fides eius ad iustitiam
ROM|4|6|sicut et David dicit beatitudinem hominis cui Deus accepto fert iustitiam sine operibus
ROM|4|7|beati quorum remissae sunt iniquitates et quorum tecta sunt peccata
ROM|4|8|beatus vir cui non inputabit Dominus peccatum
ROM|4|9|beatitudo ergo haec in circumcisione an etiam in praeputio dicimus enim quia reputata est Abrahae fides ad iustitiam
ROM|4|10|quomodo ergo reputata est in circumcisione an in praeputio non in circumcisione sed in praeputio
ROM|4|11|et signum accepit circumcisionis signaculum iustitiae fidei quae est in praeputio ut sit pater omnium credentium per praeputium ut reputetur et illis ad iustitiam
ROM|4|12|et sit pater circumcisionis non his tantum qui sunt ex circumcisione sed et his qui sectantur vestigia quae est in praeputio fidei patris nostri Abrahae
ROM|4|13|non enim per legem promissio Abrahae aut semini eius ut heres esset mundi sed per iustitiam fidei
ROM|4|14|si enim qui ex lege heredes sunt exinanita est fides abolita est promissio
ROM|4|15|lex enim iram operatur ubi enim non est lex nec praevaricatio
ROM|4|16|ideo ex fide ut secundum gratiam ut firma sit promissio omni semini non ei qui ex lege est solum sed et ei qui ex fide est Abrahae qui est pater omnium nostrum
ROM|4|17|sicut scriptum est quia patrem multarum gentium posui te ante Deum cui credidit qui vivificat mortuos et vocat quae non sunt tamquam ea quae sunt
ROM|4|18|qui contra spem in spem credidit ut fieret pater multarum gentium secundum quod dictum est sic erit semen tuum
ROM|4|19|et non infirmatus fide consideravit corpus suum emortuum cum fere centum annorum esset et emortuam vulvam Sarrae
ROM|4|20|in repromissione etiam Dei non haesitavit diffidentia sed confortatus est fide dans gloriam Deo
ROM|4|21|plenissime sciens quia quaecumque promisit potens est et facere
ROM|4|22|ideo et reputatum est illi ad iustitiam
ROM|4|23|non est autem scriptum tantum propter ipsum quia reputatum est illi
ROM|4|24|sed et propter nos quibus reputabitur credentibus in eum qui suscitavit Iesum Dominum nostrum a mortuis
ROM|4|25|qui traditus est propter delicta nostra et resurrexit propter iustificationem nostram
ROM|5|1|iustificati igitur ex fide pacem habeamus ad Deum per Dominum nostrum Iesum Christum
ROM|5|2|per quem et accessum habemus fide in gratiam istam in qua stamus et gloriamur in spe gloriae filiorum Dei
ROM|5|3|non solum autem sed et gloriamur in tribulationibus scientes quod tribulatio patientiam operatur
ROM|5|4|patientia autem probationem probatio vero spem
ROM|5|5|spes autem non confundit quia caritas Dei diffusa est in cordibus nostris per Spiritum Sanctum qui datus est nobis
ROM|5|6|ut quid enim Christus cum adhuc infirmi essemus secundum tempus pro impiis mortuus est
ROM|5|7|vix enim pro iusto quis moritur nam pro bono forsitan quis et audeat mori
ROM|5|8|commendat autem suam caritatem Deus in nos quoniam cum adhuc peccatores essemus
ROM|5|9|Christus pro nobis mortuus est multo igitur magis iustificati nunc in sanguine ipsius salvi erimus ab ira per ipsum
ROM|5|10|si enim cum inimici essemus reconciliati sumus Deo per mortem Filii eius multo magis reconciliati salvi erimus in vita ipsius
ROM|5|11|non solum autem sed et gloriamur in Deo per Dominum nostrum Iesum Christum per quem nunc reconciliationem accepimus
ROM|5|12|propterea sicut per unum hominem in hunc mundum peccatum intravit et per peccatum mors et ita in omnes homines mors pertransiit in quo omnes peccaverunt
ROM|5|13|usque ad legem enim peccatum erat in mundo peccatum autem non inputatur cum lex non est
ROM|5|14|sed regnavit mors ab Adam usque ad Mosen etiam in eos qui non peccaverunt in similitudinem praevaricationis Adae qui est forma futuri
ROM|5|15|sed non sicut delictum ita et donum si enim unius delicto multi mortui sunt multo magis gratia Dei et donum in gratiam unius hominis Iesu Christi in plures abundavit
ROM|5|16|et non sicut per unum peccantem ita et donum nam iudicium ex uno in condemnationem gratia autem ex multis delictis in iustificationem
ROM|5|17|si enim in unius delicto mors regnavit per unum multo magis abundantiam gratiae et donationis et iustitiae accipientes in vita regnabunt per unum Iesum Christum
ROM|5|18|igitur sicut per unius delictum in omnes homines in condemnationem sic et per unius iustitiam in omnes homines in iustificationem vitae
ROM|5|19|sicut enim per inoboedientiam unius hominis peccatores constituti sunt multi ita et per unius oboeditionem iusti constituentur multi
ROM|5|20|lex autem subintravit ut abundaret delictum ubi autem abundavit delictum superabundavit gratia
ROM|5|21|ut sicut regnavit peccatum in morte ita et gratia regnet per iustitiam in vitam aeternam per Iesum Christum Dominum nostrum
ROM|6|1|quid ergo dicemus permanebimus in peccato ut gratia abundet
ROM|6|2|absit qui enim mortui sumus peccato quomodo adhuc vivemus in illo
ROM|6|3|an ignoratis quia quicumque baptizati sumus in Christo Iesu in morte ipsius baptizati sumus
ROM|6|4|consepulti enim sumus cum illo per baptismum in mortem ut quomodo surrexit Christus a mortuis per gloriam Patris ita et nos in novitate vitae ambulemus
ROM|6|5|si enim conplantati facti sumus similitudini mortis eius simul et resurrectionis erimus
ROM|6|6|hoc scientes quia vetus homo noster simul crucifixus est ut destruatur corpus peccati ut ultra non serviamus peccato
ROM|6|7|qui enim mortuus est iustificatus est a peccato
ROM|6|8|si autem mortui sumus cum Christo credimus quia simul etiam vivemus cum Christo
ROM|6|9|scientes quod Christus surgens ex mortuis iam non moritur mors illi ultra non dominabitur
ROM|6|10|quod enim mortuus est peccato mortuus est semel quod autem vivit vivit Deo
ROM|6|11|ita et vos existimate vos mortuos quidem esse peccato viventes autem Deo in Christo Iesu
ROM|6|12|non ergo regnet peccatum in vestro mortali corpore ut oboediatis concupiscentiis eius
ROM|6|13|sed neque exhibeatis membra vestra arma iniquitatis peccato sed exhibete vos Deo tamquam ex mortuis viventes et membra vestra arma iustitiae Deo
ROM|6|14|peccatum enim vobis non dominabitur non enim sub lege estis sed sub gratia
ROM|6|15|quid ergo peccavimus quoniam non sumus sub lege sed sub gratia absit
ROM|6|16|nescitis quoniam cui exhibetis vos servos ad oboediendum servi estis eius cui oboeditis sive peccati sive oboeditionis ad iustitiam
ROM|6|17|gratias autem Deo quod fuistis servi peccati oboedistis autem ex corde in eam formam doctrinae in qua traditi estis
ROM|6|18|liberati autem a peccato servi facti estis iustitiae
ROM|6|19|humanum dico propter infirmitatem carnis vestrae sicut enim exhibuistis membra vestra servire inmunditiae et iniquitati ad iniquitatem ita nunc exhibete membra vestra servire iustitiae in sanctificationem
ROM|6|20|cum enim servi essetis peccati liberi fuistis iustitiae
ROM|6|21|quem ergo fructum habuistis tunc in quibus nunc erubescitis nam finis illorum mors est
ROM|6|22|nunc vero liberati a peccato servi autem facti Deo habetis fructum vestrum in sanctificationem finem vero vitam aeternam
ROM|6|23|stipendia enim peccati mors gratia autem Dei vita aeterna in Christo Iesu Domino nostro
ROM|7|1|an ignoratis fratres scientibus enim legem loquor quia lex in homine dominatur quanto tempore vivit
ROM|7|2|nam quae sub viro est mulier vivente viro alligata est legi si autem mortuus fuerit vir soluta est a lege viri
ROM|7|3|igitur vivente viro vocabitur adultera si fuerit cum alio viro si autem mortuus fuerit vir eius liberata est a lege ut non sit adultera si fuerit cum alio viro
ROM|7|4|itaque fratres mei et vos mortificati estis legi per corpus Christi ut sitis alterius qui ex mortuis resurrexit ut fructificaremus Deo
ROM|7|5|cum enim essemus in carne passiones peccatorum quae per legem erant operabantur in membris nostris ut fructificarent morti
ROM|7|6|nunc autem soluti sumus a lege morientes in quo detinebamur ita ut serviamus in novitate spiritus et non in vetustate litterae
ROM|7|7|quid ergo dicemus lex peccatum est absit sed peccatum non cognovi nisi per legem nam concupiscentiam nesciebam nisi lex diceret non concupisces
ROM|7|8|occasione autem accepta peccatum per mandatum operatum est in me omnem concupiscentiam sine lege enim peccatum mortuum erat
ROM|7|9|ego autem vivebam sine lege aliquando sed cum venisset mandatum peccatum revixit
ROM|7|10|ego autem mortuus sum et inventum est mihi mandatum quod erat ad vitam hoc esse ad mortem
ROM|7|11|nam peccatum occasione accepta per mandatum seduxit me et per illud occidit
ROM|7|12|itaque lex quidem sancta et mandatum sanctum et iustum et bonum
ROM|7|13|quod ergo bonum est mihi factum est mors absit sed peccatum ut appareat peccatum per bonum mihi operatum est mortem ut fiat supra modum peccans peccatum per mandatum
ROM|7|14|scimus enim quod lex spiritalis est ego autem carnalis sum venundatus sub peccato
ROM|7|15|quod enim operor non intellego non enim quod volo hoc ago sed quod odi illud facio
ROM|7|16|si autem quod nolo illud facio consentio legi quoniam bona
ROM|7|17|nunc autem iam non ego operor illud sed quod habitat in me peccatum
ROM|7|18|scio enim quia non habitat in me hoc est in carne mea bonum nam velle adiacet mihi perficere autem bonum non invenio
ROM|7|19|non enim quod volo bonum hoc facio sed quod nolo malum hoc ago
ROM|7|20|si autem quod nolo illud facio non ego operor illud sed quod habitat in me peccatum
ROM|7|21|invenio igitur legem volenti mihi facere bonum quoniam mihi malum adiacet
ROM|7|22|condelector enim legi Dei secundum interiorem hominem
ROM|7|23|video autem aliam legem in membris meis repugnantem legi mentis meae et captivantem me in lege peccati quae est in membris meis
ROM|7|24|infelix ego homo quis me liberabit de corpore mortis huius
ROM|7|25|gratia Dei per Iesum Christum Dominum nostrum igitur ego ipse mente servio legi Dei carne autem legi peccati
ROM|8|1|nihil ergo nunc damnationis est his qui sunt in Christo Iesu qui non secundum carnem ambulant
ROM|8|2|lex enim Spiritus vitae in Christo Iesu liberavit me a lege peccati et mortis
ROM|8|3|nam quod inpossibile erat legis in quo infirmabatur per carnem Deus Filium suum mittens in similitudinem carnis peccati et de peccato damnavit peccatum in carne
ROM|8|4|ut iustificatio legis impleretur in nobis qui non secundum carnem ambulamus sed secundum Spiritum
ROM|8|5|qui enim secundum carnem sunt quae carnis sunt sapiunt qui vero secundum Spiritum quae sunt Spiritus sentiunt
ROM|8|6|nam prudentia carnis mors prudentia autem Spiritus vita et pax
ROM|8|7|quoniam sapientia carnis inimicitia est in Deum legi enim Dei non subicitur nec enim potest
ROM|8|8|qui autem in carne sunt Deo placere non possunt
ROM|8|9|vos autem in carne non estis sed in Spiritu si tamen Spiritus Dei habitat in vobis si quis autem Spiritum Christi non habet hic non est eius
ROM|8|10|si autem Christus in vobis est corpus quidem mortuum est propter peccatum spiritus vero vita propter iustificationem
ROM|8|11|quod si Spiritus eius qui suscitavit Iesum a mortuis habitat in vobis qui suscitavit Iesum Christum a mortuis vivificabit et mortalia corpora vestra propter inhabitantem Spiritum eius in vobis
ROM|8|12|ergo fratres debitores sumus non carni ut secundum carnem vivamus
ROM|8|13|si enim secundum carnem vixeritis moriemini si autem Spiritu facta carnis mortificatis vivetis
ROM|8|14|quicumque enim Spiritu Dei aguntur hii filii sunt Dei
ROM|8|15|non enim accepistis spiritum servitutis iterum in timore sed accepistis Spiritum adoptionis filiorum in quo clamamus Abba Pater
ROM|8|16|ipse Spiritus testimonium reddit spiritui nostro quod sumus filii Dei
ROM|8|17|si autem filii et heredes heredes quidem Dei coheredes autem Christi si tamen conpatimur ut et conglorificemur
ROM|8|18|existimo enim quod non sunt condignae passiones huius temporis ad futuram gloriam quae revelabitur in nobis
ROM|8|19|nam expectatio creaturae revelationem filiorum Dei expectat
ROM|8|20|vanitati enim creatura subiecta est non volens sed propter eum qui subiecit in spem
ROM|8|21|quia et ipsa creatura liberabitur a servitute corruptionis in libertatem gloriae filiorum Dei
ROM|8|22|scimus enim quod omnis creatura ingemescit et parturit usque adhuc
ROM|8|23|non solum autem illa sed et nos ipsi primitias Spiritus habentes et ipsi intra nos gemimus adoptionem filiorum expectantes redemptionem corporis nostri
ROM|8|24|spe enim salvi facti sumus spes autem quae videtur non est spes nam quod videt quis quid sperat
ROM|8|25|si autem quod non videmus speramus per patientiam expectamus
ROM|8|26|similiter autem et Spiritus adiuvat infirmitatem nostram nam quid oremus sicut oportet nescimus sed ipse Spiritus postulat pro nobis gemitibus inenarrabilibus
ROM|8|27|qui autem scrutatur corda scit quid desideret Spiritus quia secundum Deum postulat pro sanctis
ROM|8|28|scimus autem quoniam diligentibus Deum omnia cooperantur in bonum his qui secundum propositum vocati sunt sancti
ROM|8|29|nam quos praescivit et praedestinavit conformes fieri imaginis Filii eius ut sit ipse primogenitus in multis fratribus
ROM|8|30|quos autem praedestinavit hos et vocavit et quos vocavit hos et iustificavit quos autem iustificavit illos et glorificavit
ROM|8|31|quid ergo dicemus ad haec si Deus pro nobis quis contra nos
ROM|8|32|qui etiam Filio suo non pepercit sed pro nobis omnibus tradidit illum quomodo non etiam cum illo omnia nobis donabit
ROM|8|33|quis accusabit adversus electos Dei Deus qui iustificat
ROM|8|34|quis est qui condemnet Christus Iesus qui mortuus est immo qui resurrexit qui et est ad dexteram Dei qui etiam interpellat pro nobis
ROM|8|35|quis nos separabit a caritate Christi tribulatio an angustia an persecutio an fames an nuditas an periculum an gladius
ROM|8|36|sicut scriptum est quia propter te mortificamur tota die aestimati sumus ut oves occisionis
ROM|8|37|sed in his omnibus superamus propter eum qui dilexit nos
ROM|8|38|certus sum enim quia neque mors neque vita neque angeli neque principatus neque instantia neque futura neque fortitudines
ROM|8|39|neque altitudo neque profundum neque creatura alia poterit nos separare a caritate Dei quae est in Christo Iesu Domino nostro
ROM|9|1|veritatem dico in Christo non mentior testimonium mihi perhibente conscientia mea in Spiritu Sancto
ROM|9|2|quoniam tristitia est mihi magna et continuus dolor cordi meo
ROM|9|3|optabam enim ipse ego anathema esse a Christo pro fratribus meis qui sunt cognati mei secundum carnem
ROM|9|4|qui sunt Israhelitae quorum adoptio est filiorum et gloria et testamenta et legislatio et obsequium et promissa
ROM|9|5|quorum patres et ex quibus Christus secundum carnem qui est super omnia Deus benedictus in saecula amen
ROM|9|6|non autem quod exciderit verbum Dei non enim omnes qui ex Israhel hii sunt Israhel
ROM|9|7|neque quia semen sunt Abrahae omnes filii sed in Isaac vocabitur tibi semen
ROM|9|8|id est non qui filii carnis hii filii Dei sed qui filii sunt promissionis aestimantur in semine
ROM|9|9|promissionis enim verbum hoc est secundum hoc tempus veniam et erit Sarrae filius
ROM|9|10|non solum autem sed et Rebecca ex uno concubitum habens Isaac patre nostro
ROM|9|11|cum enim nondum nati fuissent aut aliquid egissent bonum aut malum ut secundum electionem propositum Dei maneret
ROM|9|12|non ex operibus sed ex vocante dictum est ei quia maior serviet minori
ROM|9|13|sicut scriptum est Iacob dilexi Esau autem odio habui
ROM|9|14|quid ergo dicemus numquid iniquitas apud Deum absit
ROM|9|15|Mosi enim dicit miserebor cuius misereor et misericordiam praestabo cuius miserebor
ROM|9|16|igitur non volentis neque currentis sed miserentis Dei
ROM|9|17|dicit enim scriptura Pharaoni quia in hoc ipsum excitavi te ut ostendam in te virtutem meam et ut adnuntietur nomen meum in universa terra
ROM|9|18|ergo cuius vult miseretur et quem vult indurat
ROM|9|19|dicis itaque mihi quid adhuc queritur voluntati enim eius quis resistit
ROM|9|20|o homo tu quis es qui respondeas Deo numquid dicit figmentum ei qui se finxit quid me fecisti sic
ROM|9|21|an non habet potestatem figulus luti ex eadem massa facere aliud quidem vas in honorem aliud vero in contumeliam
ROM|9|22|quod si volens Deus ostendere iram et notam facere potentiam suam sustinuit in multa patientia vasa irae aptata in interitum
ROM|9|23|ut ostenderet divitias gloriae suae in vasa misericordiae quae praeparavit in gloriam
ROM|9|24|quos et vocavit nos non solum ex Iudaeis sed etiam ex gentibus
ROM|9|25|sicut in Osee dicit vocabo non plebem meam plebem meam et non misericordiam consecutam misericordiam consecutam
ROM|9|26|et erit in loco ubi dictum est eis non plebs mea vos ibi vocabuntur filii Dei vivi
ROM|9|27|Esaias autem clamat pro Israhel si fuerit numerus filiorum Israhel tamquam harena maris reliquiae salvae fient
ROM|9|28|verbum enim consummans et brevians in aequitate quia verbum breviatum faciet Dominus super terram
ROM|9|29|et sicut praedixit Esaias nisi Dominus Sabaoth reliquisset nobis semen sicut Sodoma facti essemus et sicut Gomorra similes fuissemus
ROM|9|30|quid ergo dicemus quod gentes quae non sectabantur iustitiam adprehenderunt iustitiam iustitiam autem quae ex fide est
ROM|9|31|Israhel vero sectans legem iustitiae in legem iustitiae non pervenit
ROM|9|32|quare quia non ex fide sed quasi ex operibus offenderunt in lapidem offensionis
ROM|9|33|sicut scriptum est ecce pono in Sion lapidem offensionis et petram scandali et omnis qui credit in eum non confundetur
ROM|10|1|fratres voluntas quidem cordis mei et obsecratio ad Deum fit pro illis in salutem
ROM|10|2|testimonium enim perhibeo illis quod aemulationem Dei habent sed non secundum scientiam
ROM|10|3|ignorantes enim Dei iustitiam et suam quaerentes statuere iustitiae Dei non sunt subiecti
ROM|10|4|finis enim legis Christus ad iustitiam omni credenti
ROM|10|5|Moses enim scripsit quoniam iustitiam quae ex lege est qui fecerit homo vivet in ea
ROM|10|6|quae autem ex fide est iustitia sic dicit ne dixeris in corde tuo quis ascendit in caelum id est Christum deducere
ROM|10|7|aut quis descendit in abyssum hoc est Christum ex mortuis revocare
ROM|10|8|sed quid dicit prope est verbum in ore tuo et in corde tuo hoc est verbum fidei quod praedicamus
ROM|10|9|quia si confitearis in ore tuo Dominum Iesum et in corde tuo credideris quod Deus illum excitavit ex mortuis salvus eris
ROM|10|10|corde enim creditur ad iustitiam ore autem confessio fit in salutem
ROM|10|11|dicit enim scriptura omnis qui credit in illum non confundetur
ROM|10|12|non enim est distinctio Iudaei et Graeci nam idem Dominus omnium dives in omnes qui invocant illum
ROM|10|13|omnis enim quicumque invocaverit nomen Domini salvus erit
ROM|10|14|quomodo ergo invocabunt in quem non crediderunt aut quomodo credent ei quem non audierunt quomodo autem audient sine praedicante
ROM|10|15|quomodo vero praedicabunt nisi mittantur sicut scriptum est quam speciosi pedes evangelizantium pacem evangelizantium bona
ROM|10|16|sed non omnes oboedierunt evangelio Esaias enim dicit Domine quis credidit auditui nostro
ROM|10|17|ergo fides ex auditu auditus autem per verbum Christi
ROM|10|18|sed dico numquid non audierunt et quidem in omnem terram exiit sonus eorum et in fines orbis terrae verba eorum
ROM|10|19|sed dico numquid Israhel non cognovit primus Moses dicit ego ad aemulationem vos adducam in non gentem in gentem insipientem in iram vos mittam
ROM|10|20|Esaias autem audet et dicit inventus sum non quaerentibus me palam apparui his qui me non interrogabant
ROM|10|21|ad Israhel autem dicit tota die expandi manus meas ad populum non credentem et contradicentem
ROM|11|1|dico ergo numquid reppulit Deus populum suum absit nam et ego Israhelita sum ex semine Abraham tribu Beniamin
ROM|11|2|non reppulit Deus plebem suam quam praesciit an nescitis in Helia quid dicit scriptura quemadmodum interpellat Deum adversus Israhel
ROM|11|3|Domine prophetas tuos occiderunt altaria tua suffoderunt et ego relictus sum solus et quaerunt animam meam
ROM|11|4|sed quid dicit illi responsum divinum reliqui mihi septem milia virorum qui non curvaverunt genu Baal
ROM|11|5|sic ergo et in hoc tempore reliquiae secundum electionem gratiae factae sunt
ROM|11|6|si autem gratia non ex operibus alioquin gratia iam non est gratia
ROM|11|7|quid ergo quod quaerebat Israhel hoc non est consecutus electio autem consecuta est ceteri vero excaecati sunt
ROM|11|8|sicut scriptum est dedit illis Deus spiritum conpunctionis oculos ut non videant et aures ut non audiant usque in hodiernum diem
ROM|11|9|et David dicit fiat mensa eorum in laqueum et in captionem et in scandalum et in retributionem illis
ROM|11|10|obscurentur oculi eorum ne videant et dorsum illorum semper incurva
ROM|11|11|dico ergo numquid sic offenderunt ut caderent absit sed illorum delicto salus gentibus ut illos aemulentur
ROM|11|12|quod si delictum illorum divitiae sunt mundi et deminutio eorum divitiae gentium quanto magis plenitudo eorum
ROM|11|13|vobis enim dico gentibus quamdiu quidem ego sum gentium apostolus ministerium meum honorificabo
ROM|11|14|si quo modo ad aemulandum provocem carnem meam et salvos faciam aliquos ex illis
ROM|11|15|si enim amissio eorum reconciliatio est mundi quae adsumptio nisi vita ex mortuis
ROM|11|16|quod si delibatio sancta est et massa et si radix sancta et rami
ROM|11|17|quod si aliqui ex ramis fracti sunt tu autem cum oleaster esses insertus es in illis et socius radicis et pinguidinis olivae factus es
ROM|11|18|noli gloriari adversus ramos quod si gloriaris non tu radicem portas sed radix te
ROM|11|19|dices ergo fracti sunt rami ut ego inserar
ROM|11|20|bene propter incredulitatem fracti sunt tu autem fide stas noli altum sapere sed time
ROM|11|21|si enim Deus naturalibus ramis non pepercit ne forte nec tibi parcat
ROM|11|22|vide ergo bonitatem et severitatem Dei in eos quidem qui ceciderunt severitatem in te autem bonitatem Dei si permanseris in bonitate alioquin et tu excideris
ROM|11|23|sed et illi si non permanserint in incredulitate inserentur potens est enim Deus iterum inserere illos
ROM|11|24|nam si tu ex naturali excisus es oleastro et contra naturam insertus es in bonam olivam quanto magis hii secundum naturam inserentur suae olivae
ROM|11|25|nolo enim vos ignorare fratres mysterium hoc ut non sitis vobis ipsis sapientes quia caecitas ex parte contigit in Israhel donec plenitudo gentium intraret
ROM|11|26|et sic omnis Israhel salvus fieret sicut scriptum est veniet ex Sion qui eripiat avertet impietates ab Iacob
ROM|11|27|et hoc illis a me testamentum cum abstulero peccata eorum
ROM|11|28|secundum evangelium quidem inimici propter vos secundum electionem autem carissimi propter patres
ROM|11|29|sine paenitentia enim sunt dona et vocatio Dei
ROM|11|30|sicut enim aliquando et vos non credidistis Deo nunc autem misericordiam consecuti estis propter illorum incredulitatem
ROM|11|31|ita et isti nunc non crediderunt in vestram misericordiam ut et ipsi misericordiam consequantur
ROM|11|32|conclusit enim Deus omnia in incredulitatem ut omnium misereatur
ROM|11|33|o altitudo divitiarum sapientiae et scientiae Dei quam inconprehensibilia sunt iudicia eius et investigabiles viae eius
ROM|11|34|quis enim cognovit sensum Domini aut quis consiliarius eius fuit
ROM|11|35|aut quis prior dedit illi et retribuetur ei
ROM|11|36|quoniam ex ipso et per ipsum et in ipso omnia ipsi gloria in saecula amen
ROM|12|1|obsecro itaque vos fratres per misericordiam Dei ut exhibeatis corpora vestra hostiam viventem sanctam Deo placentem rationabile obsequium vestrum
ROM|12|2|et nolite conformari huic saeculo sed reformamini in novitate sensus vestri ut probetis quae sit voluntas Dei bona et placens et perfecta
ROM|12|3|dico enim per gratiam quae data est mihi omnibus qui sunt inter vos non plus sapere quam oportet sapere sed sapere ad sobrietatem unicuique sicut Deus divisit mensuram fidei
ROM|12|4|sicut enim in uno corpore multa membra habemus omnia autem membra non eundem actum habent
ROM|12|5|ita multi unum corpus sumus in Christo singuli autem alter alterius membra
ROM|12|6|habentes autem donationes secundum gratiam quae data est nobis differentes sive prophetiam secundum rationem fidei
ROM|12|7|sive ministerium in ministrando sive qui docet in doctrina
ROM|12|8|qui exhortatur in exhortando qui tribuit in simplicitate qui praeest in sollicitudine qui miseretur in hilaritate
ROM|12|9|dilectio sine simulatione odientes malum adherentes bono
ROM|12|10|caritatem fraternitatis invicem diligentes honore invicem praevenientes
ROM|12|11|sollicitudine non pigri spiritu ferventes Domino servientes
ROM|12|12|spe gaudentes in tribulatione patientes orationi instantes
ROM|12|13|necessitatibus sanctorum communicantes hospitalitatem sectantes
ROM|12|14|benedicite persequentibus benedicite et nolite maledicere
ROM|12|15|gaudere cum gaudentibus flere cum flentibus
ROM|12|16|id ipsum invicem sentientes non alta sapientes sed humilibus consentientes nolite esse prudentes apud vosmet ipsos
ROM|12|17|nulli malum pro malo reddentes providentes bona non tantum coram Deo sed etiam coram omnibus hominibus
ROM|12|18|si fieri potest quod ex vobis est cum omnibus hominibus pacem habentes
ROM|12|19|non vosmet ipsos defendentes carissimi sed date locum irae scriptum est enim mihi vindictam ego retribuam dicit Dominus
ROM|12|20|sed si esurierit inimicus tuus ciba illum si sitit potum da illi hoc enim faciens carbones ignis congeres super caput eius
ROM|12|21|noli vinci a malo sed vince in bono malum
ROM|13|1|omnis anima potestatibus sublimioribus subdita sit non est enim potestas nisi a Deo quae autem sunt a Deo ordinatae sunt
ROM|13|2|itaque qui resistit potestati Dei ordinationi resistit qui autem resistunt ipsi sibi damnationem adquirunt
ROM|13|3|nam principes non sunt timori boni operis sed mali vis autem non timere potestatem bonum fac et habebis laudem ex illa
ROM|13|4|Dei enim minister est tibi in bonum si autem male feceris time non enim sine causa gladium portat Dei enim minister est vindex in iram ei qui malum agit
ROM|13|5|ideo necessitate subditi estote non solum propter iram sed et propter conscientiam
ROM|13|6|ideo enim et tributa praestatis ministri enim Dei sunt in hoc ipsum servientes
ROM|13|7|reddite omnibus debita cui tributum tributum cui vectigal vectigal cui timorem timorem cui honorem honorem
ROM|13|8|nemini quicquam debeatis nisi ut invicem diligatis qui enim diligit proximum legem implevit
ROM|13|9|nam non adulterabis non occides non furaberis non concupisces et si quod est aliud mandatum in hoc verbo instauratur diliges proximum tuum tamquam te ipsum
ROM|13|10|dilectio proximo malum non operatur plenitudo ergo legis est dilectio
ROM|13|11|et hoc scientes tempus quia hora est iam nos de somno surgere nunc enim propior est nostra salus quam cum credidimus
ROM|13|12|nox praecessit dies autem adpropiavit abiciamus ergo opera tenebrarum et induamur arma lucis
ROM|13|13|sicut in die honeste ambulemus non in comesationibus et ebrietatibus non in cubilibus et inpudicitiis non in contentione et aemulatione
ROM|13|14|sed induite Dominum Iesum Christum et carnis curam ne feceritis in desideriis
ROM|14|1|infirmum autem in fide adsumite non in disceptationibus cogitationum
ROM|14|2|alius enim credit manducare omnia qui autem infirmus est holus manducat
ROM|14|3|is qui manducat non manducantem non spernat et qui non manducat manducantem non iudicet Deus enim illum adsumpsit
ROM|14|4|tu quis es qui iudices alienum servum suo domino stat aut cadit stabit autem potens est enim Deus statuere illum
ROM|14|5|nam alius iudicat diem plus inter diem alius iudicat omnem diem unusquisque in suo sensu abundet
ROM|14|6|qui sapit diem Domino sapit et qui manducat Domino manducat gratias enim agit Deo et qui non manducat Domino non manducat et gratias agit Deo
ROM|14|7|nemo enim nostrum sibi vivit et nemo sibi moritur
ROM|14|8|sive enim vivimus Domino vivimus sive morimur Domino morimur sive ergo vivimus sive morimur Domini sumus
ROM|14|9|in hoc enim Christus et mortuus est et revixit ut et mortuorum et vivorum dominetur
ROM|14|10|tu autem quid iudicas fratrem tuum aut tu quare spernis fratrem tuum omnes enim stabimus ante tribunal Dei
ROM|14|11|scriptum est enim vivo ego dicit Dominus quoniam mihi flectet omne genu et omnis lingua confitebitur Deo
ROM|14|12|itaque unusquisque nostrum pro se rationem reddet Deo
ROM|14|13|non ergo amplius invicem iudicemus sed hoc iudicate magis ne ponatis offendiculum fratri vel scandalum
ROM|14|14|scio et confido in Domino Iesu quia nihil commune per ipsum nisi ei qui existimat quid commune esse illi commune est
ROM|14|15|si enim propter cibum frater tuus contristatur iam non secundum caritatem ambulas noli cibo tuo illum perdere pro quo Christus mortuus est
ROM|14|16|non ergo blasphemetur bonum nostrum
ROM|14|17|non est regnum Dei esca et potus sed iustitia et pax et gaudium in Spiritu Sancto
ROM|14|18|qui enim in hoc servit Christo placet Deo et probatus est hominibus
ROM|14|19|itaque quae pacis sunt sectemur et quae aedificationis sunt in invicem
ROM|14|20|noli propter escam destruere opus Dei omnia quidem munda sunt sed malum est homini qui per offendiculum manducat
ROM|14|21|bonum est non manducare carnem et non bibere vinum neque in quo frater tuus offendit aut scandalizatur aut infirmatur
ROM|14|22|tu fidem habes penes temet ipsum habe coram Deo beatus qui non iudicat semet ipsum in eo quo probat
ROM|14|23|qui autem discernit si manducaverit damnatus est quia non ex fide omne autem quod non ex fide peccatum est
ROM|15|1|debemus autem nos firmiores inbecillitates infirmorum sustinere et non nobis placere
ROM|15|2|unusquisque vestrum proximo suo placeat in bonum ad aedificationem
ROM|15|3|etenim Christus non sibi placuit sed sicut scriptum est inproperia inproperantium tibi ceciderunt super me
ROM|15|4|quaecumque enim scripta sunt ad nostram doctrinam scripta sunt ut per patientiam et consolationem scripturarum spem habeamus
ROM|15|5|Deus autem patientiae et solacii det vobis id ipsum sapere in alterutrum secundum Iesum Christum
ROM|15|6|ut unianimes uno ore honorificetis Deum et Patrem Domini nostri Iesu Christi
ROM|15|7|propter quod suscipite invicem sicut et Christus suscepit vos in honorem Dei
ROM|15|8|dico enim Christum Iesum ministrum fuisse circumcisionis propter veritatem Dei ad confirmandas promissiones patrum
ROM|15|9|gentes autem super misericordiam honorare Deum sicut scriptum est propter hoc confitebor tibi in gentibus et nomini tuo cantabo
ROM|15|10|et iterum dicit laetamini gentes cum plebe eius
ROM|15|11|et iterum laudate omnes gentes Dominum et magnificate eum omnes populi
ROM|15|12|et rursus Esaias ait erit radix Iesse et qui exsurget regere gentes in eo gentes sperabunt
ROM|15|13|Deus autem spei repleat vos omni gaudio et pace in credendo ut abundetis in spe in virtute Spiritus Sancti
ROM|15|14|certus sum autem fratres mei et ego ipse de vobis quoniam et ipsi pleni estis dilectione repleti omni scientia ita ut possitis alterutrum monere
ROM|15|15|audacius autem scripsi vobis fratres ex parte tamquam in memoriam vos reducens propter gratiam quae data est mihi a Deo
ROM|15|16|ut sim minister Christi Iesu in gentibus sanctificans evangelium Dei ut fiat oblatio gentium accepta sanctificata in Spiritu Sancto
ROM|15|17|habeo igitur gloriam in Christo Iesu ad Deum
ROM|15|18|non enim audeo aliquid loqui eorum quae per me non effecit Christus in oboedientiam gentium verbo et factis
ROM|15|19|in virtute signorum et prodigiorum in virtute Spiritus Sancti ita ut ab Hierusalem per circuitum usque in Illyricum repleverim evangelium Christi
ROM|15|20|sic autem hoc praedicavi evangelium non ubi nominatus est Christus ne super alienum fundamentum aedificarem
ROM|15|21|sed sicut scriptum est quibus non est adnuntiatum de eo videbunt et qui non audierunt intellegent
ROM|15|22|propter quod et inpediebar plurimum venire ad vos
ROM|15|23|nunc vero ulterius locum non habens in his regionibus cupiditatem autem habens veniendi ad vos ex multis iam annis
ROM|15|24|cum in Hispaniam proficisci coepero spero quod praeteriens videam vos et a vobis deducar illuc si vobis primum ex parte fruitus fuero
ROM|15|25|nunc igitur proficiscar in Hierusalem ministrare sanctis
ROM|15|26|probaverunt enim Macedonia et Achaia conlationem aliquam facere in pauperes sanctorum qui sunt in Hierusalem
ROM|15|27|placuit enim eis et debitores sunt eorum nam si spiritalium eorum participes facti sunt gentiles debent et in carnalibus ministrare eis
ROM|15|28|hoc igitur cum consummavero et adsignavero eis fructum hunc proficiscar per vos in Hispaniam
ROM|15|29|scio autem quoniam veniens ad vos in abundantia benedictionis Christi veniam
ROM|15|30|obsecro igitur vos fratres per Dominum nostrum Iesum Christum et per caritatem Spiritus ut adiuvetis me in orationibus pro me ad Deum
ROM|15|31|ut liberer ab infidelibus qui sunt in Iudaea et obsequii mei oblatio accepta fiat in Hierosolyma sanctis
ROM|15|32|ut veniam ad vos in gaudio per voluntatem Dei et refrigerer vobiscum
ROM|15|33|Deus autem pacis sit cum omnibus vobis amen
ROM|16|1|commendo autem vobis Phoebem sororem nostram quae est in ministerio ecclesiae quae est Cenchris
ROM|16|2|ut eam suscipiatis in Domino digne sanctis et adsistatis ei in quocumque negotio vestri indiguerit etenim ipsa quoque adstitit multis et mihi ipsi
ROM|16|3|salutate Priscam et Aquilam adiutores meos in Christo Iesu
ROM|16|4|qui pro anima mea suas cervices subposuerunt quibus non solus ego gratias ago sed et cunctae ecclesiae gentium
ROM|16|5|et domesticam eorum ecclesiam salutate Ephaenetum dilectum mihi qui est primitivus Asiae in Christo
ROM|16|6|salutate Mariam quae multum laboravit in vobis
ROM|16|7|salutate Andronicum et Iuniam cognatos et concaptivos meos qui sunt nobiles in apostolis qui et ante me fuerunt in Christo
ROM|16|8|salutate Ampliatum dilectissimum mihi in Domino
ROM|16|9|salutate Urbanum adiutorem nostrum in Christo et Stachyn dilectum meum
ROM|16|10|salutate Apellen probum in Christo
ROM|16|11|salutate eos qui sunt ex Aristoboli salutate Herodionem cognatum meum salutate eos qui sunt ex Narcissi qui sunt in Domino
ROM|16|12|salutate Tryfenam et Tryfosam quae laborant in Domino salutate Persidam carissimam quae multum laboravit in Domino
ROM|16|13|salutate Rufum electum in Domino et matrem eius et meam
ROM|16|14|salutate Asyncritum Flegonta Hermen Patrobam Hermam et qui cum eis sunt fratres
ROM|16|15|salutate Filologum et Iuliam Nereum et sororem eius et Olympiadem et omnes qui cum eis sunt sanctos
ROM|16|16|salutate invicem in osculo sancto salutant vos omnes ecclesiae Christi
ROM|16|17|rogo autem vos fratres ut observetis eos qui dissensiones et offendicula praeter doctrinam quam vos didicistis faciunt et declinate ab illis
ROM|16|18|huiusmodi enim Christo Domino nostro non serviunt sed suo ventri et per dulces sermones et benedictiones seducunt corda innocentium
ROM|16|19|vestra enim oboedientia in omnem locum divulgata est gaudeo igitur in vobis sed volo vos sapientes esse in bono et simplices in malo
ROM|16|20|Deus autem pacis conteret Satanan sub pedibus vestris velociter gratia Domini nostri Iesu Christi vobiscum
ROM|16|21|salutat vos Timotheus adiutor meus et Lucius et Iason et Sosipater cognati mei
ROM|16|22|saluto vos ego Tertius qui scripsi epistulam in Domino
ROM|16|23|salutat vos Gaius hospes meus et universae ecclesiae salutat vos Erastus arcarius civitatis et Quartus frater
ROM|16|24|
ROM|16|25|ei autem qui potens est vos confirmare iuxta evangelium meum et praedicationem Iesu Christi secundum revelationem mysterii temporibus aeternis taciti
ROM|16|26|quod nunc patefactum est per scripturas prophetarum secundum praeceptum aeterni Dei ad oboeditionem fidei in cunctis gentibus cognito
ROM|16|27|solo sapienti Deo per Iesum Christum cui honor in saecula saeculorum amen
