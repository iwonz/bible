HAG|1|1|in anno secundo Darii regis in mense sexto in die una mensis factum est verbum Domini in manu Aggei prophetae ad Zorobabel filium Salathihel ducem Iuda et ad Iesum filium Iosedech sacerdotem magnum dicens
HAG|1|2|haec ait Dominus exercituum dicens populus iste dicit nondum venit tempus domus Domini aedificandae
HAG|1|3|et factum est verbum Domini in manu Aggei prophetae dicens
HAG|1|4|numquid tempus vobis est ut habitetis in domibus laqueatis et domus ista deserta
HAG|1|5|et nunc haec dicit Dominus exercituum ponite corda vestra super vias vestras
HAG|1|6|seminastis multum et intulistis parum comedistis et non estis satiati bibistis et non estis inebriati operuistis vos et non estis calefacti et qui mercedes congregavit misit eas in sacculum pertusum
HAG|1|7|haec dicit Dominus exercituum ponite corda vestra super vias vestras
HAG|1|8|ascendite in montem portate lignum et aedificate domum et acceptabilis mihi erit et glorificabor dicit Dominus
HAG|1|9|respexistis ad amplius et ecce factum est minus et intulistis in domum et exsuflavi illud quam ob causam dicit Dominus exercituum quia domus mea deserta est et vos festinatis unusquisque in domum suam
HAG|1|10|propter hoc super vos prohibiti sunt caeli ne darent rorem et terra prohibita est ne daret germen suum
HAG|1|11|et vocavi siccitatem super terram et super montes et super triticum et super vinum et super oleum et quaecumque profert humus et super homines et super iumenta et super omnem laborem manuum
HAG|1|12|et audivit Zorobabel filius Salathihel et Iesus filius Iosedech sacerdos magnus et omnes reliquiae populi vocem Dei sui et verba Aggei prophetae sicut misit eum Dominus Deus eorum ad ipsos et timuit populus a facie Domini
HAG|1|13|et dixit Aggeus nuntius Domini de nuntiis Domini populo dicens ego vobiscum dicit Dominus
HAG|1|14|et suscitavit Dominus spiritum Zorobabel filii Salathihel ducis Iuda et spiritum Iesu filii Iosedech sacerdotis magni et spiritum reliquorum de omni populo et ingressi sunt et faciebant opus in domo Domini exercituum Dei sui
HAG|2|1|in die vicesima et quarta mensis in sexto mense in anno secundo Darii regis
HAG|2|2|in septimo mense vicesima et prima mensis factum est verbum Domini in manu Aggei prophetae dicens
HAG|2|3|loquere ad Zorobabel filium Salathihel ducem Iuda et ad Iesum filium Iosedech sacerdotem magnum et ad reliquos populi dicens
HAG|2|4|quis in vobis est derelictus qui vidit domum istam in gloria sua prima et quid vos videtis hanc nunc numquid non ita est quasi non sit in oculis vestris
HAG|2|5|et nunc confortare Zorobabel dicit Dominus et confortare Iesu fili Iosedech sacerdos magne et confortare omnis popule terrae dicit Dominus exercituum et facite quoniam ego vobiscum sum dicit Dominus exercituum
HAG|2|6|verbum quod placui vobiscum cum egrederemini de terra Aegypti et spiritus meus erit in medio vestrum nolite timere
HAG|2|7|quia haec dicit Dominus exercituum adhuc unum modicum est et ego commovebo caelum et terram et mare et aridam
HAG|2|8|et movebo omnes gentes et veniet desideratus cunctis gentibus et implebo domum istam gloria dicit Dominus exercituum
HAG|2|9|meum est argentum et meum est aurum dicit Dominus exercituum
HAG|2|10|magna erit gloria domus istius novissimae plus quam primae dicit Dominus exercituum et in loco isto dabo pacem dicit Dominus exercituum
HAG|2|11|in vicesima et quarta noni mensis in anno secundo Darii factum est verbum Domini ad Aggeum prophetam dicens
HAG|2|12|haec dicit Dominus exercituum interroga sacerdotes legem dicens
HAG|2|13|si tulerit homo carnem sanctificatam in ora vestimenti sui et tetigerit de summitate eius panem aut pulmentum aut vinum aut oleum aut omnem cibum numquid sanctificabitur respondentes autem sacerdotes dixerunt non
HAG|2|14|et dixit Aggeus si tetigerit pollutus in anima ex omnibus his numquid contaminabitur et responderunt sacerdotes et dixerunt contaminabitur
HAG|2|15|et respondit Aggeus et dixit sic populus iste et sic gens ista ante faciem meam dicit Dominus et sic omne opus manuum eorum et omnia quae obtulerint ibi contaminata erunt
HAG|2|16|et nunc ponite corda vestra a die hac et supra antequam poneretur lapis super lapidem in templo Domini
HAG|2|17|cum accederetis ad acervum viginti modiorum et fierent decem intraretis ad torcular ut exprimeretis quinquaginta lagoenas et fiebant viginti
HAG|2|18|percussi vos vento urente et aurugine et grandine omnia opera manuum vestrarum et non fuit in vobis qui reverteretur ad me dicit Dominus
HAG|2|19|ponite corda vestra ex die ista et in futurum a die vicesima et quarta noni mensis a die qua fundamenta iacta sunt templi Domini ponite super cor vestrum
HAG|2|20|numquid iam semen in germine est et adhuc vinea et ficus et malogranatum et lignum olivae non floruit ex die ista benedicam
HAG|2|21|et factum est verbum Domini secundo ad Aggeum in vicesima et quarta mensis dicens
HAG|2|22|loquere ad Zorobabel ducem Iuda dicens ego movebo caelum pariter et terram
HAG|2|23|et subvertam solium regnorum et conteram fortitudinem regni gentium et subvertam quadrigam et ascensorem eius et descendent equi et ascensores eorum vir in gladio fratris sui
HAG|2|24|in die illo dicit Dominus exercituum adsumam te Zorobabel fili Salathihel serve meus dicit Dominus et ponam te quasi signaculum quia te elegi dicit Dominus exercituum
