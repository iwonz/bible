1COR|1|1|Paul called to be an apostle of Jesus Christ through the will of God, and Sosthenes our brother,
1COR|1|2|Unto the church of God which is at Corinth, to them that are sanctified in Christ Jesus, called to be saints, with all that in every place call upon the name of Jesus Christ our Lord, both their's and our's:
1COR|1|3|Grace be unto you, and peace, from God our Father, and from the Lord Jesus Christ.
1COR|1|4|I thank my God always on your behalf, for the grace of God which is given you by Jesus Christ;
1COR|1|5|That in every thing ye are enriched by him, in all utterance, and in all knowledge;
1COR|1|6|Even as the testimony of Christ was confirmed in you:
1COR|1|7|So that ye come behind in no gift; waiting for the coming of our Lord Jesus Christ:
1COR|1|8|Who shall also confirm you unto the end, that ye may be blameless in the day of our Lord Jesus Christ.
1COR|1|9|God is faithful, by whom ye were called unto the fellowship of his Son Jesus Christ our Lord.
1COR|1|10|Now I beseech you, brethren, by the name of our Lord Jesus Christ, that ye all speak the same thing, and that there be no divisions among you; but that ye be perfectly joined together in the same mind and in the same judgment.
1COR|1|11|For it hath been declared unto me of you, my brethren, by them which are of the house of Chloe, that there are contentions among you.
1COR|1|12|Now this I say, that every one of you saith, I am of Paul; and I of Apollos; and I of Cephas; and I of Christ.
1COR|1|13|Is Christ divided? was Paul crucified for you? or were ye baptized in the name of Paul?
1COR|1|14|I thank God that I baptized none of you, but Crispus and Gaius;
1COR|1|15|Lest any should say that I had baptized in mine own name.
1COR|1|16|And I baptized also the household of Stephanas: besides, I know not whether I baptized any other.
1COR|1|17|For Christ sent me not to baptize, but to preach the gospel: not with wisdom of words, lest the cross of Christ should be made of none effect.
1COR|1|18|For the preaching of the cross is to them that perish foolishness; but unto us which are saved it is the power of God.
1COR|1|19|For it is written, I will destroy the wisdom of the wise, and will bring to nothing the understanding of the prudent.
1COR|1|20|Where is the wise? where is the scribe? where is the disputer of this world? hath not God made foolish the wisdom of this world?
1COR|1|21|For after that in the wisdom of God the world by wisdom knew not God, it pleased God by the foolishness of preaching to save them that believe.
1COR|1|22|For the Jews require a sign, and the Greeks seek after wisdom:
1COR|1|23|But we preach Christ crucified, unto the Jews a stumblingblock, and unto the Greeks foolishness;
1COR|1|24|But unto them which are called, both Jews and Greeks, Christ the power of God, and the wisdom of God.
1COR|1|25|Because the foolishness of God is wiser than men; and the weakness of God is stronger than men.
1COR|1|26|For ye see your calling, brethren, how that not many wise men after the flesh, not many mighty, not many noble, are called:
1COR|1|27|But God hath chosen the foolish things of the world to confound the wise; and God hath chosen the weak things of the world to confound the things which are mighty;
1COR|1|28|And base things of the world, and things which are despised, hath God chosen, yea, and things which are not, to bring to nought things that are:
1COR|1|29|That no flesh should glory in his presence.
1COR|1|30|But of him are ye in Christ Jesus, who of God is made unto us wisdom, and righteousness, and sanctification, and redemption:
1COR|1|31|That, according as it is written, He that glorieth, let him glory in the Lord.
1COR|2|1|And I, brethren, when I came to you, came not with excellency of speech or of wisdom, declaring unto you the testimony of God.
1COR|2|2|For I determined not to know any thing among you, save Jesus Christ, and him crucified.
1COR|2|3|And I was with you in weakness, and in fear, and in much trembling.
1COR|2|4|And my speech and my preaching was not with enticing words of man's wisdom, but in demonstration of the Spirit and of power:
1COR|2|5|That your faith should not stand in the wisdom of men, but in the power of God.
1COR|2|6|Howbeit we speak wisdom among them that are perfect: yet not the wisdom of this world, nor of the princes of this world, that come to nought:
1COR|2|7|But we speak the wisdom of God in a mystery, even the hidden wisdom, which God ordained before the world unto our glory:
1COR|2|8|Which none of the princes of this world knew: for had they known it, they would not have crucified the Lord of glory.
1COR|2|9|But as it is written, Eye hath not seen, nor ear heard, neither have entered into the heart of man, the things which God hath prepared for them that love him.
1COR|2|10|But God hath revealed them unto us by his Spirit: for the Spirit searcheth all things, yea, the deep things of God.
1COR|2|11|For what man knoweth the things of a man, save the spirit of man which is in him? even so the things of God knoweth no man, but the Spirit of God.
1COR|2|12|Now we have received, not the spirit of the world, but the spirit which is of God; that we might know the things that are freely given to us of God.
1COR|2|13|Which things also we speak, not in the words which man's wisdom teacheth, but which the Holy Ghost teacheth; comparing spiritual things with spiritual.
1COR|2|14|But the natural man receiveth not the things of the Spirit of God: for they are foolishness unto him: neither can he know them, because they are spiritually discerned.
1COR|2|15|But he that is spiritual judgeth all things, yet he himself is judged of no man.
1COR|2|16|For who hath known the mind of the Lord, that he may instruct him? But we have the mind of Christ.
1COR|3|1|And I, brethren, could not speak unto you as unto spiritual, but as unto carnal, even as unto babes in Christ.
1COR|3|2|I have fed you with milk, and not with meat: for hitherto ye were not able to bear it, neither yet now are ye able.
1COR|3|3|For ye are yet carnal: for whereas there is among you envying, and strife, and divisions, are ye not carnal, and walk as men?
1COR|3|4|For while one saith, I am of Paul; and another, I am of Apollos; are ye not carnal?
1COR|3|5|Who then is Paul, and who is Apollos, but ministers by whom ye believed, even as the Lord gave to every man?
1COR|3|6|I have planted, Apollos watered; but God gave the increase.
1COR|3|7|So then neither is he that planteth any thing, neither he that watereth; but God that giveth the increase.
1COR|3|8|Now he that planteth and he that watereth are one: and every man shall receive his own reward according to his own labour.
1COR|3|9|For we are labourers together with God: ye are God's husbandry, ye are God's building.
1COR|3|10|According to the grace of God which is given unto me, as a wise masterbuilder, I have laid the foundation, and another buildeth thereon. But let every man take heed how he buildeth thereupon.
1COR|3|11|For other foundation can no man lay than that is laid, which is Jesus Christ.
1COR|3|12|Now if any man build upon this foundation gold, silver, precious stones, wood, hay, stubble;
1COR|3|13|Every man's work shall be made manifest: for the day shall declare it, because it shall be revealed by fire; and the fire shall try every man's work of what sort it is.
1COR|3|14|If any man's work abide which he hath built thereupon, he shall receive a reward.
1COR|3|15|If any man's work shall be burned, he shall suffer loss: but he himself shall be saved; yet so as by fire.
1COR|3|16|Know ye not that ye are the temple of God, and that the Spirit of God dwelleth in you?
1COR|3|17|If any man defile the temple of God, him shall God destroy; for the temple of God is holy, which temple ye are.
1COR|3|18|Let no man deceive himself. If any man among you seemeth to be wise in this world, let him become a fool, that he may be wise.
1COR|3|19|For the wisdom of this world is foolishness with God. For it is written, He taketh the wise in their own craftiness.
1COR|3|20|And again, The Lord knoweth the thoughts of the wise, that they are vain.
1COR|3|21|Therefore let no man glory in men. For all things are your's;
1COR|3|22|Whether Paul, or Apollos, or Cephas, or the world, or life, or death, or things present, or things to come; all are your's;
1COR|3|23|And ye are Christ's; and Christ is God's.
1COR|4|1|Let a man so account of us, as of the ministers of Christ, and stewards of the mysteries of God.
1COR|4|2|Moreover it is required in stewards, that a man be found faithful.
1COR|4|3|But with me it is a very small thing that I should be judged of you, or of man's judgment: yea, I judge not mine own self.
1COR|4|4|For I know nothing by myself; yet am I not hereby justified: but he that judgeth me is the Lord.
1COR|4|5|Therefore judge nothing before the time, until the Lord come, who both will bring to light the hidden things of darkness, and will make manifest the counsels of the hearts: and then shall every man have praise of God.
1COR|4|6|And these things, brethren, I have in a figure transferred to myself and to Apollos for your sakes; that ye might learn in us not to think of men above that which is written, that no one of you be puffed up for one against another.
1COR|4|7|For who maketh thee to differ from another? and what hast thou that thou didst not receive? now if thou didst receive it, why dost thou glory, as if thou hadst not received it?
1COR|4|8|Now ye are full, now ye are rich, ye have reigned as kings without us: and I would to God ye did reign, that we also might reign with you.
1COR|4|9|For I think that God hath set forth us the apostles last, as it were appointed to death: for we are made a spectacle unto the world, and to angels, and to men.
1COR|4|10|We are fools for Christ's sake, but ye are wise in Christ; we are weak, but ye are strong; ye are honourable, but we are despised.
1COR|4|11|Even unto this present hour we both hunger, and thirst, and are naked, and are buffeted, and have no certain dwellingplace;
1COR|4|12|And labour, working with our own hands: being reviled, we bless; being persecuted, we suffer it:
1COR|4|13|Being defamed, we intreat: we are made as the filth of the world, and are the offscouring of all things unto this day.
1COR|4|14|I write not these things to shame you, but as my beloved sons I warn you.
1COR|4|15|For though ye have ten thousand instructers in Christ, yet have ye not many fathers: for in Christ Jesus I have begotten you through the gospel.
1COR|4|16|Wherefore I beseech you, be ye followers of me.
1COR|4|17|For this cause have I sent unto you Timotheus, who is my beloved son, and faithful in the Lord, who shall bring you into remembrance of my ways which be in Christ, as I teach every where in every church.
1COR|4|18|Now some are puffed up, as though I would not come to you.
1COR|4|19|But I will come to you shortly, if the Lord will, and will know, not the speech of them which are puffed up, but the power.
1COR|4|20|For the kingdom of God is not in word, but in power.
1COR|4|21|What will ye? shall I come unto you with a rod, or in love, and in the spirit of meekness?
1COR|5|1|It is reported commonly that there is fornication among you, and such fornication as is not so much as named among the Gentiles, that one should have his father's wife.
1COR|5|2|And ye are puffed up, and have not rather mourned, that he that hath done this deed might be taken away from among you.
1COR|5|3|For I verily, as absent in body, but present in spirit, have judged already, as though I were present, concerning him that hath so done this deed,
1COR|5|4|In the name of our Lord Jesus Christ, when ye are gathered together, and my spirit, with the power of our Lord Jesus Christ,
1COR|5|5|To deliver such an one unto Satan for the destruction of the flesh, that the spirit may be saved in the day of the Lord Jesus.
1COR|5|6|Your glorying is not good. Know ye not that a little leaven leaveneth the whole lump?
1COR|5|7|Purge out therefore the old leaven, that ye may be a new lump, as ye are unleavened. For even Christ our passover is sacrificed for us:
1COR|5|8|Therefore let us keep the feast, not with old leaven, neither with the leaven of malice and wickedness; but with the unleavened bread of sincerity and truth.
1COR|5|9|I wrote unto you in an epistle not to company with fornicators:
1COR|5|10|Yet not altogether with the fornicators of this world, or with the covetous, or extortioners, or with idolaters; for then must ye needs go out of the world.
1COR|5|11|But now I have written unto you not to keep company, if any man that is called a brother be a fornicator, or covetous, or an idolater, or a railer, or a drunkard, or an extortioner; with such an one no not to eat.
1COR|5|12|For what have I to do to judge them also that are without? do not ye judge them that are within?
1COR|5|13|But them that are without God judgeth. Therefore put away from among yourselves that wicked person.
1COR|6|1|Dare any of you, having a matter against another, go to law before the unjust, and not before the saints?
1COR|6|2|Do ye not know that the saints shall judge the world? and if the world shall be judged by you, are ye unworthy to judge the smallest matters?
1COR|6|3|Know ye not that we shall judge angels? how much more things that pertain to this life?
1COR|6|4|If then ye have judgments of things pertaining to this life, set them to judge who are least esteemed in the church.
1COR|6|5|I speak to your shame. Is it so, that there is not a wise man among you? no, not one that shall be able to judge between his brethren?
1COR|6|6|But brother goeth to law with brother, and that before the unbelievers.
1COR|6|7|Now therefore there is utterly a fault among you, because ye go to law one with another. Why do ye not rather take wrong? why do ye not rather suffer yourselves to be defrauded?
1COR|6|8|Nay, ye do wrong, and defraud, and that your brethren.
1COR|6|9|Know ye not that the unrighteous shall not inherit the kingdom of God? Be not deceived: neither fornicators, nor idolaters, nor adulterers, nor effeminate, nor abusers of themselves with mankind,
1COR|6|10|Nor thieves, nor covetous, nor drunkards, nor revilers, nor extortioners, shall inherit the kingdom of God.
1COR|6|11|And such were some of you: but ye are washed, but ye are sanctified, but ye are justified in the name of the Lord Jesus, and by the Spirit of our God.
1COR|6|12|All things are lawful unto me, but all things are not expedient: all things are lawful for me, but I will not be brought under the power of any.
1COR|6|13|Meats for the belly, and the belly for meats: but God shall destroy both it and them. Now the body is not for fornication, but for the Lord; and the Lord for the body.
1COR|6|14|And God hath both raised up the Lord, and will also raise up us by his own power.
1COR|6|15|Know ye not that your bodies are the members of Christ? shall I then take the members of Christ, and make them the members of an harlot? God forbid.
1COR|6|16|What? know ye not that he which is joined to an harlot is one body? for two, saith he, shall be one flesh.
1COR|6|17|But he that is joined unto the Lord is one spirit.
1COR|6|18|Flee fornication. Every sin that a man doeth is without the body; but he that committeth fornication sinneth against his own body.
1COR|6|19|What? know ye not that your body is the temple of the Holy Ghost which is in you, which ye have of God, and ye are not your own?
1COR|6|20|For ye are bought with a price: therefore glorify God in your body, and in your spirit, which are God's.
1COR|7|1|Now concerning the things whereof ye wrote unto me: It is good for a man not to touch a woman.
1COR|7|2|Nevertheless, to avoid fornication, let every man have his own wife, and let every woman have her own husband.
1COR|7|3|Let the husband render unto the wife due benevolence: and likewise also the wife unto the husband.
1COR|7|4|The wife hath not power of her own body, but the husband: and likewise also the husband hath not power of his own body, but the wife.
1COR|7|5|Defraud ye not one the other, except it be with consent for a time, that ye may give yourselves to fasting and prayer; and come together again, that Satan tempt you not for your incontinency.
1COR|7|6|But I speak this by permission, and not of commandment.
1COR|7|7|For I would that all men were even as I myself. But every man hath his proper gift of God, one after this manner, and another after that.
1COR|7|8|I say therefore to the unmarried and widows, It is good for them if they abide even as I.
1COR|7|9|But if they cannot contain, let them marry: for it is better to marry than to burn.
1COR|7|10|And unto the married I command, yet not I, but the Lord, Let not the wife depart from her husband:
1COR|7|11|But and if she depart, let her remain unmarried or be reconciled to her husband: and let not the husband put away his wife.
1COR|7|12|But to the rest speak I, not the Lord: If any brother hath a wife that believeth not, and she be pleased to dwell with him, let him not put her away.
1COR|7|13|And the woman which hath an husband that believeth not, and if he be pleased to dwell with her, let her not leave him.
1COR|7|14|For the unbelieving husband is sanctified by the wife, and the unbelieving wife is sanctified by the husband: else were your children unclean; but now are they holy.
1COR|7|15|But if the unbelieving depart, let him depart. A brother or a sister is not under bondage in such cases: but God hath called us to peace.
1COR|7|16|For what knowest thou, O wife, whether thou shalt save thy husband? or how knowest thou, O man, whether thou shalt save thy wife?
1COR|7|17|But as God hath distributed to every man, as the Lord hath called every one, so let him walk. And so ordain I in all churches.
1COR|7|18|Is any man called being circumcised? let him not become uncircumcised. Is any called in uncircumcision? let him not be circumcised.
1COR|7|19|Circumcision is nothing, and uncircumcision is nothing, but the keeping of the commandments of God.
1COR|7|20|Let every man abide in the same calling wherein he was called.
1COR|7|21|Art thou called being a servant? care not for it: but if thou mayest be made free, use it rather.
1COR|7|22|For he that is called in the Lord, being a servant, is the Lord's freeman: likewise also he that is called, being free, is Christ's servant.
1COR|7|23|Ye are bought with a price; be not ye the servants of men.
1COR|7|24|Brethren, let every man, wherein he is called, therein abide with God.
1COR|7|25|Now concerning virgins I have no commandment of the Lord: yet I give my judgment, as one that hath obtained mercy of the Lord to be faithful.
1COR|7|26|I suppose therefore that this is good for the present distress, I say, that it is good for a man so to be.
1COR|7|27|Art thou bound unto a wife? seek not to be loosed. Art thou loosed from a wife? seek not a wife.
1COR|7|28|But and if thou marry, thou hast not sinned; and if a virgin marry, she hath not sinned. Nevertheless such shall have trouble in the flesh: but I spare you.
1COR|7|29|But this I say, brethren, the time is short: it remaineth, that both they that have wives be as though they had none;
1COR|7|30|And they that weep, as though they wept not; and they that rejoice, as though they rejoiced not; and they that buy, as though they possessed not;
1COR|7|31|And they that use this world, as not abusing it: for the fashion of this world passeth away.
1COR|7|32|But I would have you without carefulness. He that is unmarried careth for the things that belong to the Lord, how he may please the Lord:
1COR|7|33|But he that is married careth for the things that are of the world, how he may please his wife.
1COR|7|34|There is difference also between a wife and a virgin. The unmarried woman careth for the things of the Lord, that she may be holy both in body and in spirit: but she that is married careth for the things of the world, how she may please her husband.
1COR|7|35|And this I speak for your own profit; not that I may cast a snare upon you, but for that which is comely, and that ye may attend upon the Lord without distraction.
1COR|7|36|But if any man think that he behaveth himself uncomely toward his virgin, if she pass the flower of her age, and need so require, let him do what he will, he sinneth not: let them marry.
1COR|7|37|Nevertheless he that standeth stedfast in his heart, having no necessity, but hath power over his own will, and hath so decreed in his heart that he will keep his virgin, doeth well.
1COR|7|38|So then he that giveth her in marriage doeth well; but he that giveth her not in marriage doeth better.
1COR|7|39|The wife is bound by the law as long as her husband liveth; but if her husband be dead, she is at liberty to be married to whom she will; only in the Lord.
1COR|7|40|But she is happier if she so abide, after my judgment: and I think also that I have the Spirit of God.
1COR|8|1|Now as touching things offered unto idols, we know that we all have knowledge. Knowledge puffeth up, but charity edifieth.
1COR|8|2|And if any man think that he knoweth any thing, he knoweth nothing yet as he ought to know.
1COR|8|3|But if any man love God, the same is known of him.
1COR|8|4|As concerning therefore the eating of those things that are offered in sacrifice unto idols, we know that an idol is nothing in the world, and that there is none other God but one.
1COR|8|5|For though there be that are called gods, whether in heaven or in earth, (as there be gods many, and lords many,)
1COR|8|6|But to us there is but one God, the Father, of whom are all things, and we in him; and one Lord Jesus Christ, by whom are all things, and we by him.
1COR|8|7|Howbeit there is not in every man that knowledge: for some with conscience of the idol unto this hour eat it as a thing offered unto an idol; and their conscience being weak is defiled.
1COR|8|8|But meat commendeth us not to God: for neither, if we eat, are we the better; neither, if we eat not, are we the worse.
1COR|8|9|But take heed lest by any means this liberty of your's become a stumblingblock to them that are weak.
1COR|8|10|For if any man see thee which hast knowledge sit at meat in the idol's temple, shall not the conscience of him which is weak be emboldened to eat those things which are offered to idols;
1COR|8|11|And through thy knowledge shall the weak brother perish, for whom Christ died?
1COR|8|12|But when ye sin so against the brethren, and wound their weak conscience, ye sin against Christ.
1COR|8|13|Wherefore, if meat make my brother to offend, I will eat no flesh while the world standeth, lest I make my brother to offend.
1COR|9|1|Am I not an apostle? am I not free? have I not seen Jesus Christ our Lord? are not ye my work in the Lord?
1COR|9|2|If I be not an apostle unto others, yet doubtless I am to you: for the seal of mine apostleship are ye in the Lord.
1COR|9|3|Mine answer to them that do examine me is this,
1COR|9|4|Have we not power to eat and to drink?
1COR|9|5|Have we not power to lead about a sister, a wife, as well as other apostles, and as the brethren of the Lord, and Cephas?
1COR|9|6|Or I only and Barnabas, have not we power to forbear working?
1COR|9|7|Who goeth a warfare any time at his own charges? who planteth a vineyard, and eateth not of the fruit thereof? or who feedeth a flock, and eateth not of the milk of the flock?
1COR|9|8|Say I these things as a man? or saith not the law the same also?
1COR|9|9|For it is written in the law of Moses, Thou shalt not muzzle the mouth of the ox that treadeth out the corn. Doth God take care for oxen?
1COR|9|10|Or saith he it altogether for our sakes? For our sakes, no doubt, this is written: that he that ploweth should plow in hope; and that he that thresheth in hope should be partaker of his hope.
1COR|9|11|If we have sown unto you spiritual things, is it a great thing if we shall reap your carnal things?
1COR|9|12|If others be partakers of this power over you, are not we rather? Nevertheless we have not used this power; but suffer all things, lest we should hinder the gospel of Christ.
1COR|9|13|Do ye not know that they which minister about holy things live of the things of the temple? and they which wait at the altar are partakers with the altar?
1COR|9|14|Even so hath the Lord ordained that they which preach the gospel should live of the gospel.
1COR|9|15|But I have used none of these things: neither have I written these things, that it should be so done unto me: for it were better for me to die, than that any man should make my glorying void.
1COR|9|16|For though I preach the gospel, I have nothing to glory of: for necessity is laid upon me; yea, woe is unto me, if I preach not the gospel!
1COR|9|17|For if I do this thing willingly, I have a reward: but if against my will, a dispensation of the gospel is committed unto me.
1COR|9|18|What is my reward then? Verily that, when I preach the gospel, I may make the gospel of Christ without charge, that I abuse not my power in the gospel.
1COR|9|19|For though I be free from all men, yet have I made myself servant unto all, that I might gain the more.
1COR|9|20|And unto the Jews I became as a Jew, that I might gain the Jews; to them that are under the law, as under the law, that I might gain them that are under the law;
1COR|9|21|To them that are without law, as without law, (being not without law to God, but under the law to Christ,) that I might gain them that are without law.
1COR|9|22|To the weak became I as weak, that I might gain the weak: I am made all things to all men, that I might by all means save some.
1COR|9|23|And this I do for the gospel's sake, that I might be partaker thereof with you.
1COR|9|24|Know ye not that they which run in a race run all, but one receiveth the prize? So run, that ye may obtain.
1COR|9|25|And every man that striveth for the mastery is temperate in all things. Now they do it to obtain a corruptible crown; but we an incorruptible.
1COR|9|26|I therefore so run, not as uncertainly; so fight I, not as one that beateth the air:
1COR|9|27|But I keep under my body, and bring it into subjection: lest that by any means, when I have preached to others, I myself should be a castaway.
1COR|10|1|Moreover, brethren, I would not that ye should be ignorant, how that all our fathers were under the cloud, and all passed through the sea;
1COR|10|2|And were all baptized unto Moses in the cloud and in the sea;
1COR|10|3|And did all eat the same spiritual meat;
1COR|10|4|And did all drink the same spiritual drink: for they drank of that spiritual Rock that followed them: and that Rock was Christ.
1COR|10|5|But with many of them God was not well pleased: for they were overthrown in the wilderness.
1COR|10|6|Now these things were our examples, to the intent we should not lust after evil things, as they also lusted.
1COR|10|7|Neither be ye idolaters, as were some of them; as it is written, The people sat down to eat and drink, and rose up to play.
1COR|10|8|Neither let us commit fornication, as some of them committed, and fell in one day three and twenty thousand.
1COR|10|9|Neither let us tempt Christ, as some of them also tempted, and were destroyed of serpents.
1COR|10|10|Neither murmur ye, as some of them also murmured, and were destroyed of the destroyer.
1COR|10|11|Now all these things happened unto them for ensamples: and they are written for our admonition, upon whom the ends of the world are come.
1COR|10|12|Wherefore let him that thinketh he standeth take heed lest he fall.
1COR|10|13|There hath no temptation taken you but such as is common to man: but God is faithful, who will not suffer you to be tempted above that ye are able; but will with the temptation also make a way to escape, that ye may be able to bear it.
1COR|10|14|Wherefore, my dearly beloved, flee from idolatry.
1COR|10|15|I speak as to wise men; judge ye what I say.
1COR|10|16|The cup of blessing which we bless, is it not the communion of the blood of Christ? The bread which we break, is it not the communion of the body of Christ?
1COR|10|17|For we being many are one bread, and one body: for we are all partakers of that one bread.
1COR|10|18|Behold Israel after the flesh: are not they which eat of the sacrifices partakers of the altar?
1COR|10|19|What say I then? that the idol is any thing, or that which is offered in sacrifice to idols is any thing?
1COR|10|20|But I say, that the things which the Gentiles sacrifice, they sacrifice to devils, and not to God: and I would not that ye should have fellowship with devils.
1COR|10|21|Ye cannot drink the cup of the Lord, and the cup of devils: ye cannot be partakers of the Lord's table, and of the table of devils.
1COR|10|22|Do we provoke the Lord to jealousy? are we stronger than he?
1COR|10|23|All things are lawful for me, but all things are not expedient: all things are lawful for me, but all things edify not.
1COR|10|24|Let no man seek his own, but every man another's wealth.
1COR|10|25|Whatsoever is sold in the shambles, that eat, asking no question for conscience sake:
1COR|10|26|For the earth is the Lord's, and the fulness thereof.
1COR|10|27|If any of them that believe not bid you to a feast, and ye be disposed to go; whatsoever is set before you, eat, asking no question for conscience sake.
1COR|10|28|But if any man say unto you, This is offered in sacrifice unto idols, eat not for his sake that shewed it, and for conscience sake: for the earth is the Lord's, and the fulness thereof:
1COR|10|29|Conscience, I say, not thine own, but of the other: for why is my liberty judged of another man's conscience?
1COR|10|30|For if I by grace be a partaker, why am I evil spoken of for that for which I give thanks?
1COR|10|31|Whether therefore ye eat, or drink, or whatsoever ye do, do all to the glory of God.
1COR|10|32|Give none offence, neither to the Jews, nor to the Gentiles, nor to the church of God:
1COR|10|33|Even as I please all men in all things, not seeking mine own profit, but the profit of many, that they may be saved.
1COR|11|1|Be ye followers of me, even as I also am of Christ.
1COR|11|2|Now I praise you, brethren, that ye remember me in all things, and keep the ordinances, as I delivered them to you.
1COR|11|3|But I would have you know, that the head of every man is Christ; and the head of the woman is the man; and the head of Christ is God.
1COR|11|4|Every man praying or prophesying, having his head covered, dishonoureth his head.
1COR|11|5|But every woman that prayeth or prophesieth with her head uncovered dishonoureth her head: for that is even all one as if she were shaven.
1COR|11|6|For if the woman be not covered, let her also be shorn: but if it be a shame for a woman to be shorn or shaven, let her be covered.
1COR|11|7|For a man indeed ought not to cover his head, forasmuch as he is the image and glory of God: but the woman is the glory of the man.
1COR|11|8|For the man is not of the woman: but the woman of the man.
1COR|11|9|Neither was the man created for the woman; but the woman for the man.
1COR|11|10|For this cause ought the woman to have power on her head because of the angels.
1COR|11|11|Nevertheless neither is the man without the woman, neither the woman without the man, in the Lord.
1COR|11|12|For as the woman is of the man, even so is the man also by the woman; but all things of God.
1COR|11|13|Judge in yourselves: is it comely that a woman pray unto God uncovered?
1COR|11|14|Doth not even nature itself teach you, that, if a man have long hair, it is a shame unto him?
1COR|11|15|But if a woman have long hair, it is a glory to her: for her hair is given her for a covering.
1COR|11|16|But if any man seem to be contentious, we have no such custom, neither the churches of God.
1COR|11|17|Now in this that I declare unto you I praise you not, that ye come together not for the better, but for the worse.
1COR|11|18|For first of all, when ye come together in the church, I hear that there be divisions among you; and I partly believe it.
1COR|11|19|For there must be also heresies among you, that they which are approved may be made manifest among you.
1COR|11|20|When ye come together therefore into one place, this is not to eat the Lord's supper.
1COR|11|21|For in eating every one taketh before other his own supper: and one is hungry, and another is drunken.
1COR|11|22|What? have ye not houses to eat and to drink in? or despise ye the church of God, and shame them that have not? What shall I say to you? shall I praise you in this? I praise you not.
1COR|11|23|For I have received of the Lord that which also I delivered unto you, That the Lord Jesus the same night in which he was betrayed took bread:
1COR|11|24|And when he had given thanks, he brake it, and said, Take, eat: this is my body, which is broken for you: this do in remembrance of me.
1COR|11|25|After the same manner also he took the cup, when he had supped, saying, This cup is the new testament in my blood: this do ye, as oft as ye drink it, in remembrance of me.
1COR|11|26|For as often as ye eat this bread, and drink this cup, ye do shew the Lord's death till he come.
1COR|11|27|Wherefore whosoever shall eat this bread, and drink this cup of the Lord, unworthily, shall be guilty of the body and blood of the Lord.
1COR|11|28|But let a man examine himself, and so let him eat of that bread, and drink of that cup.
1COR|11|29|For he that eateth and drinketh unworthily, eateth and drinketh damnation to himself, not discerning the Lord's body.
1COR|11|30|For this cause many are weak and sickly among you, and many sleep.
1COR|11|31|For if we would judge ourselves, we should not be judged.
1COR|11|32|But when we are judged, we are chastened of the Lord, that we should not be condemned with the world.
1COR|11|33|Wherefore, my brethren, when ye come together to eat, tarry one for another.
1COR|11|34|And if any man hunger, let him eat at home; that ye come not together unto condemnation. And the rest will I set in order when I come.
1COR|12|1|Now concerning spiritual gifts, brethren, I would not have you ignorant.
1COR|12|2|Ye know that ye were Gentiles, carried away unto these dumb idols, even as ye were led.
1COR|12|3|Wherefore I give you to understand, that no man speaking by the Spirit of God calleth Jesus accursed: and that no man can say that Jesus is the Lord, but by the Holy Ghost.
1COR|12|4|Now there are diversities of gifts, but the same Spirit.
1COR|12|5|And there are differences of administrations, but the same Lord.
1COR|12|6|And there are diversities of operations, but it is the same God which worketh all in all.
1COR|12|7|But the manifestation of the Spirit is given to every man to profit withal.
1COR|12|8|For to one is given by the Spirit the word of wisdom; to another the word of knowledge by the same Spirit;
1COR|12|9|To another faith by the same Spirit; to another the gifts of healing by the same Spirit;
1COR|12|10|To another the working of miracles; to another prophecy; to another discerning of spirits; to another divers kinds of tongues; to another the interpretation of tongues:
1COR|12|11|But all these worketh that one and the selfsame Spirit, dividing to every man severally as he will.
1COR|12|12|For as the body is one, and hath many members, and all the members of that one body, being many, are one body: so also is Christ.
1COR|12|13|For by one Spirit are we all baptized into one body, whether we be Jews or Gentiles, whether we be bond or free; and have been all made to drink into one Spirit.
1COR|12|14|For the body is not one member, but many.
1COR|12|15|If the foot shall say, Because I am not the hand, I am not of the body; is it therefore not of the body?
1COR|12|16|And if the ear shall say, Because I am not the eye, I am not of the body; is it therefore not of the body?
1COR|12|17|If the whole body were an eye, where were the hearing? If the whole were hearing, where were the smelling?
1COR|12|18|But now hath God set the members every one of them in the body, as it hath pleased him.
1COR|12|19|And if they were all one member, where were the body?
1COR|12|20|But now are they many members, yet but one body.
1COR|12|21|And the eye cannot say unto the hand, I have no need of thee: nor again the head to the feet, I have no need of you.
1COR|12|22|Nay, much more those members of the body, which seem to be more feeble, are necessary:
1COR|12|23|And those members of the body, which we think to be less honourable, upon these we bestow more abundant honour; and our uncomely parts have more abundant comeliness.
1COR|12|24|For our comely parts have no need: but God hath tempered the body together, having given more abundant honour to that part which lacked.
1COR|12|25|That there should be no schism in the body; but that the members should have the same care one for another.
1COR|12|26|And whether one member suffer, all the members suffer with it; or one member be honoured, all the members rejoice with it.
1COR|12|27|Now ye are the body of Christ, and members in particular.
1COR|12|28|And God hath set some in the church, first apostles, secondarily prophets, thirdly teachers, after that miracles, then gifts of healings, helps, governments, diversities of tongues.
1COR|12|29|Are all apostles? are all prophets? are all teachers? are all workers of miracles?
1COR|12|30|Have all the gifts of healing? do all speak with tongues? do all interpret?
1COR|12|31|But covet earnestly the best gifts: and yet shew I unto you a more excellent way.
1COR|13|1|Though I speak with the tongues of men and of angels, and have not charity, I am become as sounding brass, or a tinkling cymbal.
1COR|13|2|And though I have the gift of prophecy, and understand all mysteries, and all knowledge; and though I have all faith, so that I could remove mountains, and have not charity, I am nothing.
1COR|13|3|And though I bestow all my goods to feed the poor, and though I give my body to be burned, and have not charity, it profiteth me nothing.
1COR|13|4|Charity suffereth long, and is kind; charity envieth not; charity vaunteth not itself, is not puffed up,
1COR|13|5|Doth not behave itself unseemly, seeketh not her own, is not easily provoked, thinketh no evil;
1COR|13|6|Rejoiceth not in iniquity, but rejoiceth in the truth;
1COR|13|7|Beareth all things, believeth all things, hopeth all things, endureth all things.
1COR|13|8|Charity never faileth: but whether there be prophecies, they shall fail; whether there be tongues, they shall cease; whether there be knowledge, it shall vanish away.
1COR|13|9|For we know in part, and we prophesy in part.
1COR|13|10|But when that which is perfect is come, then that which is in part shall be done away.
1COR|13|11|When I was a child, I spake as a child, I understood as a child, I thought as a child: but when I became a man, I put away childish things.
1COR|13|12|For now we see through a glass, darkly; but then face to face: now I know in part; but then shall I know even as also I am known.
1COR|13|13|And now abideth faith, hope, charity, these three; but the greatest of these is charity.
1COR|14|1|Follow after charity, and desire spiritual gifts, but rather that ye may prophesy.
1COR|14|2|For he that speaketh in an unknown tongue speaketh not unto men, but unto God: for no man understandeth him; howbeit in the spirit he speaketh mysteries.
1COR|14|3|But he that prophesieth speaketh unto men to edification, and exhortation, and comfort.
1COR|14|4|He that speaketh in an unknown tongue edifieth himself; but he that prophesieth edifieth the church.
1COR|14|5|I would that ye all spake with tongues but rather that ye prophesied: for greater is he that prophesieth than he that speaketh with tongues, except he interpret, that the church may receive edifying.
1COR|14|6|Now, brethren, if I come unto you speaking with tongues, what shall I profit you, except I shall speak to you either by revelation, or by knowledge, or by prophesying, or by doctrine?
1COR|14|7|And even things without life giving sound, whether pipe or harp, except they give a distinction in the sounds, how shall it be known what is piped or harped?
1COR|14|8|For if the trumpet give an uncertain sound, who shall prepare himself to the battle?
1COR|14|9|So likewise ye, except ye utter by the tongue words easy to be understood, how shall it be known what is spoken? for ye shall speak into the air.
1COR|14|10|There are, it may be, so many kinds of voices in the world, and none of them is without signification.
1COR|14|11|Therefore if I know not the meaning of the voice, I shall be unto him that speaketh a barbarian, and he that speaketh shall be a barbarian unto me.
1COR|14|12|Even so ye, forasmuch as ye are zealous of spiritual gifts, seek that ye may excel to the edifying of the church.
1COR|14|13|Wherefore let him that speaketh in an unknown tongue pray that he may interpret.
1COR|14|14|For if I pray in an unknown tongue, my spirit prayeth, but my understanding is unfruitful.
1COR|14|15|What is it then? I will pray with the spirit, and I will pray with the understanding also: I will sing with the spirit, and I will sing with the understanding also.
1COR|14|16|Else when thou shalt bless with the spirit, how shall he that occupieth the room of the unlearned say Amen at thy giving of thanks, seeing he understandeth not what thou sayest?
1COR|14|17|For thou verily givest thanks well, but the other is not edified.
1COR|14|18|I thank my God, I speak with tongues more than ye all:
1COR|14|19|Yet in the church I had rather speak five words with my understanding, that by my voice I might teach others also, than ten thousand words in an unknown tongue.
1COR|14|20|Brethren, be not children in understanding: howbeit in malice be ye children, but in understanding be men.
1COR|14|21|In the law it is written, With men of other tongues and other lips will I speak unto this people; and yet for all that will they not hear me, saith the Lord.
1COR|14|22|Wherefore tongues are for a sign, not to them that believe, but to them that believe not: but prophesying serveth not for them that believe not, but for them which believe.
1COR|14|23|If therefore the whole church be come together into one place, and all speak with tongues, and there come in those that are unlearned, or unbelievers, will they not say that ye are mad?
1COR|14|24|But if all prophesy, and there come in one that believeth not, or one unlearned, he is convinced of all, he is judged of all:
1COR|14|25|And thus are the secrets of his heart made manifest; and so falling down on his face he will worship God, and report that God is in you of a truth.
1COR|14|26|How is it then, brethren? when ye come together, every one of you hath a psalm, hath a doctrine, hath a tongue, hath a revelation, hath an interpretation. Let all things be done unto edifying.
1COR|14|27|If any man speak in an unknown tongue, let it be by two, or at the most by three, and that by course; and let one interpret.
1COR|14|28|But if there be no interpreter, let him keep silence in the church; and let him speak to himself, and to God.
1COR|14|29|Let the prophets speak two or three, and let the other judge.
1COR|14|30|If any thing be revealed to another that sitteth by, let the first hold his peace.
1COR|14|31|For ye may all prophesy one by one, that all may learn, and all may be comforted.
1COR|14|32|And the spirits of the prophets are subject to the prophets.
1COR|14|33|For God is not the author of confusion, but of peace, as in all churches of the saints.
1COR|14|34|Let your women keep silence in the churches: for it is not permitted unto them to speak; but they are commanded to be under obedience as also saith the law.
1COR|14|35|And if they will learn any thing, let them ask their husbands at home: for it is a shame for women to speak in the church.
1COR|14|36|What? came the word of God out from you? or came it unto you only?
1COR|14|37|If any man think himself to be a prophet, or spiritual, let him acknowledge that the things that I write unto you are the commandments of the Lord.
1COR|14|38|But if any man be ignorant, let him be ignorant.
1COR|14|39|Wherefore, brethren, covet to prophesy, and forbid not to speak with tongues.
1COR|14|40|Let all things be done decently and in order.
1COR|15|1|Moreover, brethren, I declare unto you the gospel which I preached unto you, which also ye have received, and wherein ye stand;
1COR|15|2|By which also ye are saved, if ye keep in memory what I preached unto you, unless ye have believed in vain.
1COR|15|3|For I delivered unto you first of all that which I also received, how that Christ died for our sins according to the scriptures;
1COR|15|4|And that he was buried, and that he rose again the third day according to the scriptures:
1COR|15|5|And that he was seen of Cephas, then of the twelve:
1COR|15|6|After that, he was seen of above five hundred brethren at once; of whom the greater part remain unto this present, but some are fallen asleep.
1COR|15|7|After that, he was seen of James; then of all the apostles.
1COR|15|8|And last of all he was seen of me also, as of one born out of due time.
1COR|15|9|For I am the least of the apostles, that am not meet to be called an apostle, because I persecuted the church of God.
1COR|15|10|But by the grace of God I am what I am: and his grace which was bestowed upon me was not in vain; but I laboured more abundantly than they all: yet not I, but the grace of God which was with me.
1COR|15|11|Therefore whether it were I or they, so we preach, and so ye believed.
1COR|15|12|Now if Christ be preached that he rose from the dead, how say some among you that there is no resurrection of the dead?
1COR|15|13|But if there be no resurrection of the dead, then is Christ not risen:
1COR|15|14|And if Christ be not risen, then is our preaching vain, and your faith is also vain.
1COR|15|15|Yea, and we are found false witnesses of God; because we have testified of God that he raised up Christ: whom he raised not up, if so be that the dead rise not.
1COR|15|16|For if the dead rise not, then is not Christ raised:
1COR|15|17|And if Christ be not raised, your faith is vain; ye are yet in your sins.
1COR|15|18|Then they also which are fallen asleep in Christ are perished.
1COR|15|19|If in this life only we have hope in Christ, we are of all men most miserable.
1COR|15|20|But now is Christ risen from the dead, and become the firstfruits of them that slept.
1COR|15|21|For since by man came death, by man came also the resurrection of the dead.
1COR|15|22|For as in Adam all die, even so in Christ shall all be made alive.
1COR|15|23|But every man in his own order: Christ the firstfruits; afterward they that are Christ's at his coming.
1COR|15|24|Then cometh the end, when he shall have delivered up the kingdom to God, even the Father; when he shall have put down all rule and all authority and power.
1COR|15|25|For he must reign, till he hath put all enemies under his feet.
1COR|15|26|The last enemy that shall be destroyed is death.
1COR|15|27|For he hath put all things under his feet. But when he saith all things are put under him, it is manifest that he is excepted, which did put all things under him.
1COR|15|28|And when all things shall be subdued unto him, then shall the Son also himself be subject unto him that put all things under him, that God may be all in all.
1COR|15|29|Else what shall they do which are baptized for the dead, if the dead rise not at all? why are they then baptized for the dead?
1COR|15|30|And why stand we in jeopardy every hour?
1COR|15|31|I protest by your rejoicing which I have in Christ Jesus our Lord, I die daily.
1COR|15|32|If after the manner of men I have fought with beasts at Ephesus, what advantageth it me, if the dead rise not? let us eat and drink; for to morrow we die.
1COR|15|33|Be not deceived: evil communications corrupt good manners.
1COR|15|34|Awake to righteousness, and sin not; for some have not the knowledge of God: I speak this to your shame.
1COR|15|35|But some man will say, How are the dead raised up? and with what body do they come?
1COR|15|36|Thou fool, that which thou sowest is not quickened, except it die:
1COR|15|37|And that which thou sowest, thou sowest not that body that shall be, but bare grain, it may chance of wheat, or of some other grain:
1COR|15|38|But God giveth it a body as it hath pleased him, and to every seed his own body.
1COR|15|39|All flesh is not the same flesh: but there is one kind of flesh of men, another flesh of beasts, another of fishes, and another of birds.
1COR|15|40|There are also celestial bodies, and bodies terrestrial: but the glory of the celestial is one, and the glory of the terrestrial is another.
1COR|15|41|There is one glory of the sun, and another glory of the moon, and another glory of the stars: for one star differeth from another star in glory.
1COR|15|42|So also is the resurrection of the dead. It is sown in corruption; it is raised in incorruption:
1COR|15|43|It is sown in dishonour; it is raised in glory: it is sown in weakness; it is raised in power:
1COR|15|44|It is sown a natural body; it is raised a spiritual body. There is a natural body, and there is a spiritual body.
1COR|15|45|And so it is written, The first man Adam was made a living soul; the last Adam was made a quickening spirit.
1COR|15|46|Howbeit that was not first which is spiritual, but that which is natural; and afterward that which is spiritual.
1COR|15|47|The first man is of the earth, earthy; the second man is the Lord from heaven.
1COR|15|48|As is the earthy, such are they also that are earthy: and as is the heavenly, such are they also that are heavenly.
1COR|15|49|And as we have borne the image of the earthy, we shall also bear the image of the heavenly.
1COR|15|50|Now this I say, brethren, that flesh and blood cannot inherit the kingdom of God; neither doth corruption inherit incorruption.
1COR|15|51|Behold, I shew you a mystery; We shall not all sleep, but we shall all be changed,
1COR|15|52|In a moment, in the twinkling of an eye, at the last trump: for the trumpet shall sound, and the dead shall be raised incorruptible, and we shall be changed.
1COR|15|53|For this corruptible must put on incorruption, and this mortal must put on immortality.
1COR|15|54|So when this corruptible shall have put on incorruption, and this mortal shall have put on immortality, then shall be brought to pass the saying that is written, Death is swallowed up in victory.
1COR|15|55|O death, where is thy sting? O grave, where is thy victory?
1COR|15|56|The sting of death is sin; and the strength of sin is the law.
1COR|15|57|But thanks be to God, which giveth us the victory through our Lord Jesus Christ.
1COR|15|58|Therefore, my beloved brethren, be ye stedfast, unmoveable, always abounding in the work of the Lord, forasmuch as ye know that your labour is not in vain in the Lord.
1COR|16|1|Now concerning the collection for the saints, as I have given order to the churches of Galatia, even so do ye.
1COR|16|2|Upon the first day of the week let every one of you lay by him in store, as God hath prospered him, that there be no gatherings when I come.
1COR|16|3|And when I come, whomsoever ye shall approve by your letters, them will I send to bring your liberality unto Jerusalem.
1COR|16|4|And if it be meet that I go also, they shall go with me.
1COR|16|5|Now I will come unto you, when I shall pass through Macedonia: for I do pass through Macedonia.
1COR|16|6|And it may be that I will abide, yea, and winter with you, that ye may bring me on my journey whithersoever I go.
1COR|16|7|For I will not see you now by the way; but I trust to tarry a while with you, if the Lord permit.
1COR|16|8|But I will tarry at Ephesus until Pentecost.
1COR|16|9|For a great door and effectual is opened unto me, and there are many adversaries.
1COR|16|10|Now if Timotheus come, see that he may be with you without fear: for he worketh the work of the Lord, as I also do.
1COR|16|11|Let no man therefore despise him: but conduct him forth in peace, that he may come unto me: for I look for him with the brethren.
1COR|16|12|As touching our brother Apollos, I greatly desired him to come unto you with the brethren: but his will was not at all to come at this time; but he will come when he shall have convenient time.
1COR|16|13|Watch ye, stand fast in the faith, quit you like men, be strong.
1COR|16|14|Let all your things be done with charity.
1COR|16|15|I beseech you, brethren, (ye know the house of Stephanas, that it is the firstfruits of Achaia, and that they have addicted themselves to the ministry of the saints,)
1COR|16|16|That ye submit yourselves unto such, and to every one that helpeth with us, and laboureth.
1COR|16|17|I am glad of the coming of Stephanas and Fortunatus and Achaicus: for that which was lacking on your part they have supplied.
1COR|16|18|For they have refreshed my spirit and your's: therefore acknowledge ye them that are such.
1COR|16|19|The churches of Asia salute you. Aquila and Priscilla salute you much in the Lord, with the church that is in their house.
1COR|16|20|All the brethren greet you. Greet ye one another with an holy kiss.
1COR|16|21|The salutation of me Paul with mine own hand.
1COR|16|22|If any man love not the Lord Jesus Christ, let him be Anathema Maranatha.
1COR|16|23|The grace of our Lord Jesus Christ be with you.
1COR|16|24|My love be with you all in Christ Jesus. Amen.
