EPH|1|1|Paul, an apostle of Jesus Christ by the will of God, to the saints which are at Ephesus, and to the faithful in Christ Jesus:
EPH|1|2|Grace be to you, and peace, from God our Father, and from the Lord Jesus Christ.
EPH|1|3|Blessed be the God and Father of our Lord Jesus Christ, who hath blessed us with all spiritual blessings in heavenly places in Christ:
EPH|1|4|According as he hath chosen us in him before the foundation of the world, that we should be holy and without blame before him in love:
EPH|1|5|Having predestinated us unto the adoption of children by Jesus Christ to himself, according to the good pleasure of his will,
EPH|1|6|To the praise of the glory of his grace, wherein he hath made us accepted in the beloved.
EPH|1|7|In whom we have redemption through his blood, the forgiveness of sins, according to the riches of his grace;
EPH|1|8|Wherein he hath abounded toward us in all wisdom and prudence;
EPH|1|9|Having made known unto us the mystery of his will, according to his good pleasure which he hath purposed in himself:
EPH|1|10|That in the dispensation of the fulness of times he might gather together in one all things in Christ, both which are in heaven, and which are on earth; even in him:
EPH|1|11|In whom also we have obtained an inheritance, being predestinated according to the purpose of him who worketh all things after the counsel of his own will:
EPH|1|12|That we should be to the praise of his glory, who first trusted in Christ.
EPH|1|13|In whom ye also trusted, after that ye heard the word of truth, the gospel of your salvation: in whom also after that ye believed, ye were sealed with that holy Spirit of promise,
EPH|1|14|Which is the earnest of our inheritance until the redemption of the purchased possession, unto the praise of his glory.
EPH|1|15|Wherefore I also, after I heard of your faith in the Lord Jesus, and love unto all the saints,
EPH|1|16|Cease not to give thanks for you, making mention of you in my prayers;
EPH|1|17|That the God of our Lord Jesus Christ, the Father of glory, may give unto you the spirit of wisdom and revelation in the knowledge of him:
EPH|1|18|The eyes of your understanding being enlightened; that ye may know what is the hope of his calling, and what the riches of the glory of his inheritance in the saints,
EPH|1|19|And what is the exceeding greatness of his power to us-ward who believe, according to the working of his mighty power,
EPH|1|20|Which he wrought in Christ, when he raised him from the dead, and set him at his own right hand in the heavenly places,
EPH|1|21|Far above all principality, and power, and might, and dominion, and every name that is named, not only in this world, but also in that which is to come:
EPH|1|22|And hath put all things under his feet, and gave him to be the head over all things to the church,
EPH|1|23|Which is his body, the fulness of him that filleth all in all.
EPH|2|1|And you hath he quickened, who were dead in trespasses and sins;
EPH|2|2|Wherein in time past ye walked according to the course of this world, according to the prince of the power of the air, the spirit that now worketh in the children of disobedience:
EPH|2|3|Among whom also we all had our conversation in times past in the lusts of our flesh, fulfilling the desires of the flesh and of the mind; and were by nature the children of wrath, even as others.
EPH|2|4|But God, who is rich in mercy, for his great love wherewith he loved us,
EPH|2|5|Even when we were dead in sins, hath quickened us together with Christ, (by grace ye are saved;)
EPH|2|6|And hath raised us up together, and made us sit together in heavenly places in Christ Jesus:
EPH|2|7|That in the ages to come he might shew the exceeding riches of his grace in his kindness toward us through Christ Jesus.
EPH|2|8|For by grace are ye saved through faith; and that not of yourselves: it is the gift of God:
EPH|2|9|Not of works, lest any man should boast.
EPH|2|10|For we are his workmanship, created in Christ Jesus unto good works, which God hath before ordained that we should walk in them.
EPH|2|11|Wherefore remember, that ye being in time past Gentiles in the flesh, who are called Uncircumcision by that which is called the Circumcision in the flesh made by hands;
EPH|2|12|That at that time ye were without Christ, being aliens from the commonwealth of Israel, and strangers from the covenants of promise, having no hope, and without God in the world:
EPH|2|13|But now in Christ Jesus ye who sometimes were far off are made nigh by the blood of Christ.
EPH|2|14|For he is our peace, who hath made both one, and hath broken down the middle wall of partition between us;
EPH|2|15|Having abolished in his flesh the enmity, even the law of commandments contained in ordinances; for to make in himself of twain one new man, so making peace;
EPH|2|16|And that he might reconcile both unto God in one body by the cross, having slain the enmity thereby:
EPH|2|17|And came and preached peace to you which were afar off, and to them that were nigh.
EPH|2|18|For through him we both have access by one Spirit unto the Father.
EPH|2|19|Now therefore ye are no more strangers and foreigners, but fellowcitizens with the saints, and of the household of God;
EPH|2|20|And are built upon the foundation of the apostles and prophets, Jesus Christ himself being the chief corner stone;
EPH|2|21|In whom all the building fitly framed together groweth unto an holy temple in the Lord:
EPH|2|22|In whom ye also are builded together for an habitation of God through the Spirit.
EPH|3|1|For this cause I Paul, the prisoner of Jesus Christ for you Gentiles,
EPH|3|2|If ye have heard of the dispensation of the grace of God which is given me to you-ward:
EPH|3|3|How that by revelation he made known unto me the mystery; (as I wrote afore in few words,
EPH|3|4|Whereby, when ye read, ye may understand my knowledge in the mystery of Christ)
EPH|3|5|Which in other ages was not made known unto the sons of men, as it is now revealed unto his holy apostles and prophets by the Spirit;
EPH|3|6|That the Gentiles should be fellowheirs, and of the same body, and partakers of his promise in Christ by the gospel:
EPH|3|7|Whereof I was made a minister, according to the gift of the grace of God given unto me by the effectual working of his power.
EPH|3|8|Unto me, who am less than the least of all saints, is this grace given, that I should preach among the Gentiles the unsearchable riches of Christ;
EPH|3|9|And to make all men see what is the fellowship of the mystery, which from the beginning of the world hath been hid in God, who created all things by Jesus Christ:
EPH|3|10|To the intent that now unto the principalities and powers in heavenly places might be known by the church the manifold wisdom of God,
EPH|3|11|According to the eternal purpose which he purposed in Christ Jesus our Lord:
EPH|3|12|In whom we have boldness and access with confidence by the faith of him.
EPH|3|13|Wherefore I desire that ye faint not at my tribulations for you, which is your glory.
EPH|3|14|For this cause I bow my knees unto the Father of our Lord Jesus Christ,
EPH|3|15|Of whom the whole family in heaven and earth is named,
EPH|3|16|That he would grant you, according to the riches of his glory, to be strengthened with might by his Spirit in the inner man;
EPH|3|17|That Christ may dwell in your hearts by faith; that ye, being rooted and grounded in love,
EPH|3|18|May be able to comprehend with all saints what is the breadth, and length, and depth, and height;
EPH|3|19|And to know the love of Christ, which passeth knowledge, that ye might be filled with all the fulness of God.
EPH|3|20|Now unto him that is able to do exceeding abundantly above all that we ask or think, according to the power that worketh in us,
EPH|3|21|Unto him be glory in the church by Christ Jesus throughout all ages, world without end. Amen.
EPH|4|1|I therefore, the prisoner of the Lord, beseech you that ye walk worthy of the vocation wherewith ye are called,
EPH|4|2|With all lowliness and meekness, with longsuffering, forbearing one another in love;
EPH|4|3|Endeavouring to keep the unity of the Spirit in the bond of peace.
EPH|4|4|There is one body, and one Spirit, even as ye are called in one hope of your calling;
EPH|4|5|One Lord, one faith, one baptism,
EPH|4|6|One God and Father of all, who is above all, and through all, and in you all.
EPH|4|7|But unto every one of us is given grace according to the measure of the gift of Christ.
EPH|4|8|Wherefore he saith, When he ascended up on high, he led captivity captive, and gave gifts unto men.
EPH|4|9|(Now that he ascended, what is it but that he also descended first into the lower parts of the earth?
EPH|4|10|He that descended is the same also that ascended up far above all heavens, that he might fill all things.)
EPH|4|11|And he gave some, apostles; and some, prophets; and some, evangelists; and some, pastors and teachers;
EPH|4|12|For the perfecting of the saints, for the work of the ministry, for the edifying of the body of Christ:
EPH|4|13|Till we all come in the unity of the faith, and of the knowledge of the Son of God, unto a perfect man, unto the measure of the stature of the fulness of Christ:
EPH|4|14|That we henceforth be no more children, tossed to and fro, and carried about with every wind of doctrine, by the sleight of men, and cunning craftiness, whereby they lie in wait to deceive;
EPH|4|15|But speaking the truth in love, may grow up into him in all things, which is the head, even Christ:
EPH|4|16|From whom the whole body fitly joined together and compacted by that which every joint supplieth, according to the effectual working in the measure of every part, maketh increase of the body unto the edifying of itself in love.
EPH|4|17|This I say therefore, and testify in the Lord, that ye henceforth walk not as other Gentiles walk, in the vanity of their mind,
EPH|4|18|Having the understanding darkened, being alienated from the life of God through the ignorance that is in them, because of the blindness of their heart:
EPH|4|19|Who being past feeling have given themselves over unto lasciviousness, to work all uncleanness with greediness.
EPH|4|20|But ye have not so learned Christ;
EPH|4|21|If so be that ye have heard him, and have been taught by him, as the truth is in Jesus:
EPH|4|22|That ye put off concerning the former conversation the old man, which is corrupt according to the deceitful lusts;
EPH|4|23|And be renewed in the spirit of your mind;
EPH|4|24|And that ye put on the new man, which after God is created in righteousness and true holiness.
EPH|4|25|Wherefore putting away lying, speak every man truth with his neighbour: for we are members one of another.
EPH|4|26|Be ye angry, and sin not: let not the sun go down upon your wrath:
EPH|4|27|Neither give place to the devil.
EPH|4|28|Let him that stole steal no more: but rather let him labour, working with his hands the thing which is good, that he may have to give to him that needeth.
EPH|4|29|Let no corrupt communication proceed out of your mouth, but that which is good to the use of edifying, that it may minister grace unto the hearers.
EPH|4|30|And grieve not the holy Spirit of God, whereby ye are sealed unto the day of redemption.
EPH|4|31|Let all bitterness, and wrath, and anger, and clamour, and evil speaking, be put away from you, with all malice:
EPH|4|32|And be ye kind one to another, tenderhearted, forgiving one another, even as God for Christ's sake hath forgiven you.
EPH|5|1|Be ye therefore followers of God, as dear children;
EPH|5|2|And walk in love, as Christ also hath loved us, and hath given himself for us an offering and a sacrifice to God for a sweetsmelling savour.
EPH|5|3|But fornication, and all uncleanness, or covetousness, let it not be once named among you, as becometh saints;
EPH|5|4|Neither filthiness, nor foolish talking, nor jesting, which are not convenient: but rather giving of thanks.
EPH|5|5|For this ye know, that no whoremonger, nor unclean person, nor covetous man, who is an idolater, hath any inheritance in the kingdom of Christ and of God.
EPH|5|6|Let no man deceive you with vain words: for because of these things cometh the wrath of God upon the children of disobedience.
EPH|5|7|Be not ye therefore partakers with them.
EPH|5|8|For ye were sometimes darkness, but now are ye light in the Lord: walk as children of light:
EPH|5|9|(For the fruit of the Spirit is in all goodness and righteousness and truth;)
EPH|5|10|Proving what is acceptable unto the Lord.
EPH|5|11|And have no fellowship with the unfruitful works of darkness, but rather reprove them.
EPH|5|12|For it is a shame even to speak of those things which are done of them in secret.
EPH|5|13|But all things that are reproved are made manifest by the light: for whatsoever doth make manifest is light.
EPH|5|14|Wherefore he saith, Awake thou that sleepest, and arise from the dead, and Christ shall give thee light.
EPH|5|15|See then that ye walk circumspectly, not as fools, but as wise,
EPH|5|16|Redeeming the time, because the days are evil.
EPH|5|17|Wherefore be ye not unwise, but understanding what the will of the Lord is.
EPH|5|18|And be not drunk with wine, wherein is excess; but be filled with the Spirit;
EPH|5|19|Speaking to yourselves in psalms and hymns and spiritual songs, singing and making melody in your heart to the Lord;
EPH|5|20|Giving thanks always for all things unto God and the Father in the name of our Lord Jesus Christ;
EPH|5|21|Submitting yourselves one to another in the fear of God.
EPH|5|22|Wives, submit yourselves unto your own husbands, as unto the Lord.
EPH|5|23|For the husband is the head of the wife, even as Christ is the head of the church: and he is the saviour of the body.
EPH|5|24|Therefore as the church is subject unto Christ, so let the wives be to their own husbands in every thing.
EPH|5|25|Husbands, love your wives, even as Christ also loved the church, and gave himself for it;
EPH|5|26|That he might sanctify and cleanse it with the washing of water by the word,
EPH|5|27|That he might present it to himself a glorious church, not having spot, or wrinkle, or any such thing; but that it should be holy and without blemish.
EPH|5|28|So ought men to love their wives as their own bodies. He that loveth his wife loveth himself.
EPH|5|29|For no man ever yet hated his own flesh; but nourisheth and cherisheth it, even as the Lord the church:
EPH|5|30|For we are members of his body, of his flesh, and of his bones.
EPH|5|31|For this cause shall a man leave his father and mother, and shall be joined unto his wife, and they two shall be one flesh.
EPH|5|32|This is a great mystery: but I speak concerning Christ and the church.
EPH|5|33|Nevertheless let every one of you in particular so love his wife even as himself; and the wife see that she reverence her husband.
EPH|6|1|Children, obey your parents in the Lord: for this is right.
EPH|6|2|Honour thy father and mother; which is the first commandment with promise;
EPH|6|3|That it may be well with thee, and thou mayest live long on the earth.
EPH|6|4|And, ye fathers, provoke not your children to wrath: but bring them up in the nurture and admonition of the Lord.
EPH|6|5|Servants, be obedient to them that are your masters according to the flesh, with fear and trembling, in singleness of your heart, as unto Christ;
EPH|6|6|Not with eyeservice, as menpleasers; but as the servants of Christ, doing the will of God from the heart;
EPH|6|7|With good will doing service, as to the Lord, and not to men:
EPH|6|8|Knowing that whatsoever good thing any man doeth, the same shall he receive of the Lord, whether he be bond or free.
EPH|6|9|And, ye masters, do the same things unto them, forbearing threatening: knowing that your Master also is in heaven; neither is there respect of persons with him.
EPH|6|10|Finally, my brethren, be strong in the Lord, and in the power of his might.
EPH|6|11|Put on the whole armour of God, that ye may be able to stand against the wiles of the devil.
EPH|6|12|For we wrestle not against flesh and blood, but against principalities, against powers, against the rulers of the darkness of this world, against spiritual wickedness in high places.
EPH|6|13|Wherefore take unto you the whole armour of God, that ye may be able to withstand in the evil day, and having done all, to stand.
EPH|6|14|Stand therefore, having your loins girt about with truth, and having on the breastplate of righteousness;
EPH|6|15|And your feet shod with the preparation of the gospel of peace;
EPH|6|16|Above all, taking the shield of faith, wherewith ye shall be able to quench all the fiery darts of the wicked.
EPH|6|17|And take the helmet of salvation, and the sword of the Spirit, which is the word of God:
EPH|6|18|Praying always with all prayer and supplication in the Spirit, and watching thereunto with all perseverance and supplication for all saints;
EPH|6|19|And for me, that utterance may be given unto me, that I may open my mouth boldly, to make known the mystery of the gospel,
EPH|6|20|For which I am an ambassador in bonds: that therein I may speak boldly, as I ought to speak.
EPH|6|21|But that ye also may know my affairs, and how I do, Tychicus, a beloved brother and faithful minister in the Lord, shall make known to you all things:
EPH|6|22|Whom I have sent unto you for the same purpose, that ye might know our affairs, and that he might comfort your hearts.
EPH|6|23|Peace be to the brethren, and love with faith, from God the Father and the Lord Jesus Christ.
EPH|6|24|Grace be with all them that love our Lord Jesus Christ in sincerity. Amen.
