1THESS|1|1|Paul, and Silvanus, and Timotheus, unto the church of the Thessalonians which is in God the Father and in the Lord Jesus Christ: Grace be unto you, and peace, from God our Father, and the Lord Jesus Christ.
1THESS|1|2|We give thanks to God always for you all, making mention of you in our prayers;
1THESS|1|3|Remembering without ceasing your work of faith, and labour of love, and patience of hope in our Lord Jesus Christ, in the sight of God and our Father;
1THESS|1|4|Knowing, brethren beloved, your election of God.
1THESS|1|5|For our gospel came not unto you in word only, but also in power, and in the Holy Ghost, and in much assurance; as ye know what manner of men we were among you for your sake.
1THESS|1|6|And ye became followers of us, and of the Lord, having received the word in much affliction, with joy of the Holy Ghost.
1THESS|1|7|So that ye were ensamples to all that believe in Macedonia and Achaia.
1THESS|1|8|For from you sounded out the word of the Lord not only in Macedonia and Achaia, but also in every place your faith to God-ward is spread abroad; so that we need not to speak any thing.
1THESS|1|9|For they themselves shew of us what manner of entering in we had unto you, and how ye turned to God from idols to serve the living and true God;
1THESS|1|10|And to wait for his Son from heaven, whom he raised from the dead, even Jesus, which delivered us from the wrath to come.
1THESS|2|1|For yourselves, brethren, know our entrance in unto you, that it was not in vain:
1THESS|2|2|But even after that we had suffered before, and were shamefully entreated, as ye know, at Philippi, we were bold in our God to speak unto you the gospel of God with much contention.
1THESS|2|3|For our exhortation was not of deceit, nor of uncleanness, nor in guile:
1THESS|2|4|But as we were allowed of God to be put in trust with the gospel, even so we speak; not as pleasing men, but God, which trieth our hearts.
1THESS|2|5|For neither at any time used we flattering words, as ye know, nor a cloke of covetousness; God is witness:
1THESS|2|6|Nor of men sought we glory, neither of you, nor yet of others, when we might have been burdensome, as the apostles of Christ.
1THESS|2|7|But we were gentle among you, even as a nurse cherisheth her children:
1THESS|2|8|So being affectionately desirous of you, we were willing to have imparted unto you, not the gospel of God only, but also our own souls, because ye were dear unto us.
1THESS|2|9|For ye remember, brethren, our labour and travail: for labouring night and day, because we would not be chargeable unto any of you, we preached unto you the gospel of God.
1THESS|2|10|Ye are witnesses, and God also, how holily and justly and unblameably we behaved ourselves among you that believe:
1THESS|2|11|As ye know how we exhorted and comforted and charged every one of you, as a father doth his children,
1THESS|2|12|That ye would walk worthy of God, who hath called you unto his kingdom and glory.
1THESS|2|13|For this cause also thank we God without ceasing, because, when ye received the word of God which ye heard of us, ye received it not as the word of men, but as it is in truth, the word of God, which effectually worketh also in you that believe.
1THESS|2|14|For ye, brethren, became followers of the churches of God which in Judaea are in Christ Jesus: for ye also have suffered like things of your own countrymen, even as they have of the Jews:
1THESS|2|15|Who both killed the Lord Jesus, and their own prophets, and have persecuted us; and they please not God, and are contrary to all men:
1THESS|2|16|Forbidding us to speak to the Gentiles that they might be saved, to fill up their sins alway: for the wrath is come upon them to the uttermost.
1THESS|2|17|But we, brethren, being taken from you for a short time in presence, not in heart, endeavoured the more abundantly to see your face with great desire.
1THESS|2|18|Wherefore we would have come unto you, even I Paul, once and again; but Satan hindered us.
1THESS|2|19|For what is our hope, or joy, or crown of rejoicing? Are not even ye in the presence of our Lord Jesus Christ at his coming?
1THESS|2|20|For ye are our glory and joy.
1THESS|3|1|Wherefore when we could no longer forbear, we thought it good to be left at Athens alone;
1THESS|3|2|And sent Timotheus, our brother, and minister of God, and our fellowlabourer in the gospel of Christ, to establish you, and to comfort you concerning your faith:
1THESS|3|3|That no man should be moved by these afflictions: for yourselves know that we are appointed thereunto.
1THESS|3|4|For verily, when we were with you, we told you before that we should suffer tribulation; even as it came to pass, and ye know.
1THESS|3|5|For this cause, when I could no longer forbear, I sent to know your faith, lest by some means the tempter have tempted you, and our labour be in vain.
1THESS|3|6|But now when Timotheus came from you unto us, and brought us good tidings of your faith and charity, and that ye have good remembrance of us always, desiring greatly to see us, as we also to see you:
1THESS|3|7|Therefore, brethren, we were comforted over you in all our affliction and distress by your faith:
1THESS|3|8|For now we live, if ye stand fast in the Lord.
1THESS|3|9|For what thanks can we render to God again for you, for all the joy wherewith we joy for your sakes before our God;
1THESS|3|10|Night and day praying exceedingly that we might see your face, and might perfect that which is lacking in your faith?
1THESS|3|11|Now God himself and our Father, and our Lord Jesus Christ, direct our way unto you.
1THESS|3|12|And the Lord make you to increase and abound in love one toward another, and toward all men, even as we do toward you:
1THESS|3|13|To the end he may stablish your hearts unblameable in holiness before God, even our Father, at the coming of our Lord Jesus Christ with all his saints.
1THESS|4|1|Furthermore then we beseech you, brethren, and exhort you by the Lord Jesus, that as ye have received of us how ye ought to walk and to please God, so ye would abound more and more.
1THESS|4|2|For ye know what commandments we gave you by the Lord Jesus.
1THESS|4|3|For this is the will of God, even your sanctification, that ye should abstain from fornication:
1THESS|4|4|That every one of you should know how to possess his vessel in sanctification and honour;
1THESS|4|5|Not in the lust of concupiscence, even as the Gentiles which know not God:
1THESS|4|6|That no man go beyond and defraud his brother in any matter: because that the Lord is the avenger of all such, as we also have forewarned you and testified.
1THESS|4|7|For God hath not called us unto uncleanness, but unto holiness.
1THESS|4|8|He therefore that despiseth, despiseth not man, but God, who hath also given unto us his holy Spirit.
1THESS|4|9|But as touching brotherly love ye need not that I write unto you: for ye yourselves are taught of God to love one another.
1THESS|4|10|And indeed ye do it toward all the brethren which are in all Macedonia: but we beseech you, brethren, that ye increase more and more;
1THESS|4|11|And that ye study to be quiet, and to do your own business, and to work with your own hands, as we commanded you;
1THESS|4|12|That ye may walk honestly toward them that are without, and that ye may have lack of nothing.
1THESS|4|13|But I would not have you to be ignorant, brethren, concerning them which are asleep, that ye sorrow not, even as others which have no hope.
1THESS|4|14|For if we believe that Jesus died and rose again, even so them also which sleep in Jesus will God bring with him.
1THESS|4|15|For this we say unto you by the word of the Lord, that we which are alive and remain unto the coming of the Lord shall not prevent them which are asleep.
1THESS|4|16|For the Lord himself shall descend from heaven with a shout, with the voice of the archangel, and with the trump of God: and the dead in Christ shall rise first:
1THESS|4|17|Then we which are alive and remain shall be caught up together with them in the clouds, to meet the Lord in the air: and so shall we ever be with the Lord.
1THESS|4|18|Wherefore comfort one another with these words.
1THESS|5|1|But of the times and the seasons, brethren, ye have no need that I write unto you.
1THESS|5|2|For yourselves know perfectly that the day of the Lord so cometh as a thief in the night.
1THESS|5|3|For when they shall say, Peace and safety; then sudden destruction cometh upon them, as travail upon a woman with child; and they shall not escape.
1THESS|5|4|But ye, brethren, are not in darkness, that that day should overtake you as a thief.
1THESS|5|5|Ye are all the children of light, and the children of the day: we are not of the night, nor of darkness.
1THESS|5|6|Therefore let us not sleep, as do others; but let us watch and be sober.
1THESS|5|7|For they that sleep sleep in the night; and they that be drunken are drunken in the night.
1THESS|5|8|But let us, who are of the day, be sober, putting on the breastplate of faith and love; and for an helmet, the hope of salvation.
1THESS|5|9|For God hath not appointed us to wrath, but to obtain salvation by our Lord Jesus Christ,
1THESS|5|10|Who died for us, that, whether we wake or sleep, we should live together with him.
1THESS|5|11|Wherefore comfort yourselves together, and edify one another, even as also ye do.
1THESS|5|12|And we beseech you, brethren, to know them which labour among you, and are over you in the Lord, and admonish you;
1THESS|5|13|And to esteem them very highly in love for their work's sake. And be at peace among yourselves.
1THESS|5|14|Now we exhort you, brethren, warn them that are unruly, comfort the feebleminded, support the weak, be patient toward all men.
1THESS|5|15|See that none render evil for evil unto any man; but ever follow that which is good, both among yourselves, and to all men.
1THESS|5|16|Rejoice evermore.
1THESS|5|17|Pray without ceasing.
1THESS|5|18|In every thing give thanks: for this is the will of God in Christ Jesus concerning you.
1THESS|5|19|Quench not the Spirit.
1THESS|5|20|Despise not prophesyings.
1THESS|5|21|Prove all things; hold fast that which is good.
1THESS|5|22|Abstain from all appearance of evil.
1THESS|5|23|And the very God of peace sanctify you wholly; and I pray God your whole spirit and soul and body be preserved blameless unto the coming of our Lord Jesus Christ.
1THESS|5|24|Faithful is he that calleth you, who also will do it.
1THESS|5|25|Brethren, pray for us.
1THESS|5|26|Greet all the brethren with an holy kiss.
1THESS|5|27|I charge you by the Lord that this epistle be read unto all the holy brethren.
1THESS|5|28|The grace of our Lord Jesus Christ be with you. Amen.
