HAB|1|1|The oracle that Habakkuk the prophet received.
HAB|1|2|How long, O LORD, must I call for help, but you do not listen? Or cry out to you, "Violence!" but you do not save?
HAB|1|3|Why do you make me look at injustice? Why do you tolerate wrong? Destruction and violence are before me; there is strife, and conflict abounds.
HAB|1|4|Therefore the law is paralyzed, and justice never prevails. The wicked hem in the righteous, so that justice is perverted.
HAB|1|5|"Look at the nations and watch- and be utterly amazed. For I am going to do something in your days that you would not believe, even if you were told.
HAB|1|6|I am raising up the Babylonians, that ruthless and impetuous people, who sweep across the whole earth to seize dwelling places not their own.
HAB|1|7|They are a feared and dreaded people; they are a law to themselves and promote their own honor.
HAB|1|8|Their horses are swifter than leopards, fiercer than wolves at dusk. Their cavalry gallops headlong; their horsemen come from afar. They fly like a vulture swooping to devour;
HAB|1|9|they all come bent on violence. Their hordes advance like a desert wind and gather prisoners like sand.
HAB|1|10|They deride kings and scoff at rulers. They laugh at all fortified cities; they build earthen ramps and capture them.
HAB|1|11|Then they sweep past like the wind and go on- guilty men, whose own strength is their god."
HAB|1|12|O LORD, are you not from everlasting? My God, my Holy One, we will not die. O LORD, you have appointed them to execute judgment; O Rock, you have ordained them to punish.
HAB|1|13|Your eyes are too pure to look on evil; you cannot tolerate wrong. Why then do you tolerate the treacherous? Why are you silent while the wicked swallow up those more righteous than themselves?
HAB|1|14|You have made men like fish in the sea, like sea creatures that have no ruler.
HAB|1|15|The wicked foe pulls all of them up with hooks, he catches them in his net, he gathers them up in his dragnet; and so he rejoices and is glad.
HAB|1|16|Therefore he sacrifices to his net and burns incense to his dragnet, for by his net he lives in luxury and enjoys the choicest food.
HAB|1|17|Is he to keep on emptying his net, destroying nations without mercy?
HAB|2|1|I will stand at my watch and station myself on the ramparts; I will look to see what he will say to me, and what answer I am to give to this complaint.
HAB|2|2|Then the LORD replied: "Write down the revelation and make it plain on tablets so that a herald may run with it.
HAB|2|3|For the revelation awaits an appointed time; it speaks of the end and will not prove false. Though it linger, wait for it; it will certainly come and will not delay.
HAB|2|4|"See, he is puffed up; his desires are not upright- but the righteous will live by his faith -
HAB|2|5|indeed, wine betrays him; he is arrogant and never at rest. Because he is as greedy as the grave and like death is never satisfied, he gathers to himself all the nations and takes captive all the peoples.
HAB|2|6|"Will not all of them taunt him with ridicule and scorn, saying, "'Woe to him who piles up stolen goods and makes himself wealthy by extortion! How long must this go on?'
HAB|2|7|Will not your debtors suddenly arise? Will they not wake up and make you tremble? Then you will become their victim.
HAB|2|8|Because you have plundered many nations, the peoples who are left will plunder you. For you have shed man's blood; you have destroyed lands and cities and everyone in them.
HAB|2|9|"Woe to him who builds his realm by unjust gain to set his nest on high, to escape the clutches of ruin!
HAB|2|10|You have plotted the ruin of many peoples, shaming your own house and forfeiting your life.
HAB|2|11|The stones of the wall will cry out, and the beams of the woodwork will echo it.
HAB|2|12|"Woe to him who builds a city with bloodshed and establishes a town by crime!
HAB|2|13|Has not the LORD Almighty determined that the people's labor is only fuel for the fire, that the nations exhaust themselves for nothing?
HAB|2|14|For the earth will be filled with the knowledge of the glory of the LORD, as the waters cover the sea.
HAB|2|15|"Woe to him who gives drink to his neighbors, pouring it from the wineskin till they are drunk, so that he can gaze on their naked bodies.
HAB|2|16|You will be filled with shame instead of glory. Now it is your turn! Drink and be exposed! The cup from the LORD's right hand is coming around to you, and disgrace will cover your glory.
HAB|2|17|The violence you have done to Lebanon will overwhelm you, and your destruction of animals will terrify you. For you have shed man's blood; you have destroyed lands and cities and everyone in them.
HAB|2|18|"Of what value is an idol, since a man has carved it? Or an image that teaches lies? For he who makes it trusts in his own creation; he makes idols that cannot speak.
HAB|2|19|Woe to him who says to wood, 'Come to life!' Or to lifeless stone, 'Wake up!' Can it give guidance? It is covered with gold and silver; there is no breath in it.
HAB|2|20|But the LORD is in his holy temple; let all the earth be silent before him."
HAB|3|1|A prayer of Habakkuk the prophet. On shigionoth.
HAB|3|2|LORD, I have heard of your fame; I stand in awe of your deeds, O LORD. Renew them in our day, in our time make them known; in wrath remember mercy.
HAB|3|3|God came from Teman, the Holy One from Mount Paran. Selah His glory covered the heavens and his praise filled the earth.
HAB|3|4|His splendor was like the sunrise; rays flashed from his hand, where his power was hidden.
HAB|3|5|Plague went before him; pestilence followed his steps.
HAB|3|6|He stood, and shook the earth; he looked, and made the nations tremble. The ancient mountains crumbled and the age-old hills collapsed. His ways are eternal.
HAB|3|7|I saw the tents of Cushan in distress, the dwellings of Midian in anguish.
HAB|3|8|Were you angry with the rivers, O LORD? Was your wrath against the streams? Did you rage against the sea when you rode with your horses and your victorious chariots?
HAB|3|9|You uncovered your bow, you called for many arrows. Selah You split the earth with rivers;
HAB|3|10|the mountains saw you and writhed. Torrents of water swept by; the deep roared and lifted its waves on high.
HAB|3|11|Sun and moon stood still in the heavens at the glint of your flying arrows, at the lightning of your flashing spear.
HAB|3|12|In wrath you strode through the earth and in anger you threshed the nations.
HAB|3|13|You came out to deliver your people, to save your anointed one. You crushed the leader of the land of wickedness, you stripped him from head to foot. Selah
HAB|3|14|With his own spear you pierced his head when his warriors stormed out to scatter us, gloating as though about to devour the wretched who were in hiding.
HAB|3|15|You trampled the sea with your horses, churning the great waters.
HAB|3|16|I heard and my heart pounded, my lips quivered at the sound; decay crept into my bones, and my legs trembled. Yet I will wait patiently for the day of calamity to come on the nation invading us.
HAB|3|17|Though the fig tree does not bud and there are no grapes on the vines, though the olive crop fails and the fields produce no food, though there are no sheep in the pen and no cattle in the stalls,
HAB|3|18|yet I will rejoice in the LORD, I will be joyful in God my Savior.
HAB|3|19|The Sovereign LORD is my strength; he makes my feet like the feet of a deer, he enables me to go on the heights. For the director of music. On my stringed instruments.
