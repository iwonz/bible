ZECH|1|1|In mense octavo, in anno se cundo Darii, factum est verbum Domini ad Zachariam filium Barachiae filii Addo prophetam dicens:
ZECH|1|2|" Iratus est Dominus super patres vestros iracundia.
ZECH|1|3|Et dices ad eos: Haec dicit Dominus exercituum: Convertimini ad me, ait Dominus exercituum; et convertar ad vos, dicit Dominus exercituum.
ZECH|1|4|Ne sitis sicut patres vestri, ad quos clamabant prophetae priores dicentes: Haec dicit Dominus exercituum: Convertimini de viis vestris malis et de cogitationibus vestris malis; et non audierunt neque attenderunt ad me, dicit Dominus.
ZECH|1|5|Patres vestri ubi sunt? Et prophetae numquid in sempiternum vivent?
ZECH|1|6|Verumtamen verba mea et praecepta mea, quae mandavi servis meis prophetis, numquid non attigerunt patres vestros? Et conversi sunt et dixerunt: "Sicut cogitavit Dominus exercituum facere nobis, secundum vias nostras et secundum adinventiones nostras fecit nobis" ".
ZECH|1|7|In die vicesima et quarta undecimi mensis, qui est mensis Sabath, in anno secundo Darii, factum est verbum Domini ad Zachariam filium Barachiae filii Addo prophetam dicens:
ZECH|1|8|" Vidi per noctem, et ecce vir sedens super equum rufum et ipse stabat inter myrteta, quae erant in profundo; et post eum equi rufi, fulvi et albi.
ZECH|1|9|Et dixi: "Quid sunt isti, domine mi?". Et dixit ad me angelus, qui loquebatur in me: "Ego ostendam tibi quid sint isti".
ZECH|1|10|Et respondit vir, qui stabat inter myrteta, et dixit: "Isti sunt quos misit Dominus, ut perambularent terram".
ZECH|1|11|Et responderunt angelo Domini, qui stabat inter myrteta, et dixerunt: Perambulavimus terram, et ecce omnis terra habitatur et quiescit".
ZECH|1|12|Et respondit angelus Domini et dixit: "Domine exercituum, usquequo tu non misereberis Ierusalem et urbium Iudae, quibus iratus es? Iste septuagesimus annus est!".
ZECH|1|13|Et respondit Dominus angelo, qui loquebatur in me verba bona, verba consolatoria.
ZECH|1|14|Et dixit ad me angelus, qui loquebatur in me: "Clama dicens: Haec dixit Dominus exercituum: Zelatus sum Ierusalem et Sion zelo magno,
ZECH|1|15|sed ira magna ego irascor super gentes opulentas, quia ego iratus sum parum, ipsi vero adiuverunt in malum.
ZECH|1|16|Propterea haec dicit Dominus: Revertar ad Ierusalem in misericordiis. Domus mea aedificabitur in ea, ait Dominus exercituum, et perpendiculum extendetur super Ierusalem.
ZECH|1|17|Adhuc clama dicens: Haec dicit Dominus exercituum: Adhuc affluent civitates meae bonis, et consolabitur adhuc Dominus Sion et eliget adhuc Ierusalem".
ZECH|2|1|Et levavi oculos meos et vidi, et ecce quattuor cornua;
ZECH|2|2|et dixi ad angelum, qui loquebatur in me: "Quid sunt haec?". Et dixit ad me: "Haec sunt cornua, quae ventilaverunt Iudam et Israel et Ierusalem".
ZECH|2|3|Et ostendit mihi Dominus quattuor fabros;
ZECH|2|4|et dixi: "Quid isti veniunt facere?". Qui respondit dicens: "Haec sunt cornua, quae ventilaverunt Iudam per singulos viros, ut nemo eorum levaret caput suum; et venerunt isti deterrere ea, ut deiciant cornua gentium, quae levaverunt cornu super terram Iudae, ut dispergerent eam".
ZECH|2|5|Et levavi oculos meos et vidi; et ecce vir, et in manu eius funiculus mensorum.
ZECH|2|6|Et dixi: "Quo tu vadis?". Et dixit ad me: "Ut metiar Ierusalem et videam, quanta sit latitudo eius et quanta longitudo eius".
ZECH|2|7|Et ecce angelus, qui loquebatur in me, egrediebatur, et angelus alius egrediebatur in occursum eius;
ZECH|2|8|et dixit ad eum: "Curre, loquere ad puerum istum dicens: Absque muris habitabitur Ierusalem prae multitudine hominum et iumentorum in medio eius.
ZECH|2|9|Et ego ero ei, ait Dominus, murus ignis in circuitu et in gloria ero in medio eius.
ZECH|2|10|Heu, heu! Fugite de terra aquilonis, dicit Dominus, quoniam in quattuor ventos caeli dispersi vos, dicit Dominus.
ZECH|2|11|Heu, Sion, fuge, quae habitas apud filiam Babylonis!
ZECH|2|12|Quia haec dicit Dominus exercituum, cuius gloria misit me ad gentes, quae spoliaverunt vos: Qui tetigerit vos, tangit pupillam oculi mei.
ZECH|2|13|Quia ecce ego levo manum meam super eos, et erunt praeda servorum suorum; et cognoscetis quia Dominus exercituum misit me.
ZECH|2|14|Iubila et laetare, filia Sion,quia ecce ego venioet habitabo in medio tui,ait Dominus.
ZECH|2|15|Et applicabuntur gentes multaead Dominum in die illaet erunt ei in populum.Et habitabo in medio tui,et scies quia Dominus exercituummisit me ad te.
ZECH|2|16|Et possidebit Dominus Iudampartem suam super terram sanctamet eliget adhuc Ierusalem.
ZECH|2|17|Sileat omnis caro a facie Domini,quia consurrexit de habitaculo sancto suo".
ZECH|3|1|Et ostendit mihi Iesua sacer dotem magnum stantem coram angelo Domini; et Satan stabat a dextris eius, ut adversaretur ei.
ZECH|3|2|Et dixit angelus Domini ad Satan: "Increpet Dominus in te, Satan! Et increpet Dominus in te, qui elegit Ierusalem! Numquid non iste torris est erutus de igne?".
ZECH|3|3|Et Iesua erat indutus vestibus sordidis et stabat ante faciem angeli.
ZECH|3|4|Qui respondit et ait ad eos, qui stabant coram se, dicens: "Auferte vestimenta sordida ab eo". Et dixit ad eum: "Ecce, abstuli a te iniquitatem tuam; induam te mutatoriis".
ZECH|3|5|Et dixit: "Ponite cidarim mundam super caput eius". Et posuerunt cidarim mundam super caput eius et induerunt eum vestibus; et angelus Domini stabat.
ZECH|3|6|Et contestabatur angelus Domini Iesua dicens:
ZECH|3|7|"Haec dicit Dominus exercituum: Si in viis meis ambulaveris et ministerium meum custodieris, tu quoque iudicabis domum meam et custodies atria mea; et dabo tibi accessum inter eos, qui nunc hic assistunt.
ZECH|3|8|Audi, Iesua sacerdos magne, tu et amici tui, qui sedent coram te, quia viri portendentes sunt: Ecce enim ego adduco servum meum Germen.
ZECH|3|9|Quia ecce lapis, quem dedi coram Iesua: super lapidem unum septem oculi sunt; ecce ego caelabo sculpturam eius, ait Dominus exercituum, et auferam iniquitatem terrae illius in die una.
ZECH|3|10|In die illa, oraculum Domini exercituum, vocabit vir amicum suum subter vitem et subter ficum".
ZECH|4|1|Et reversus est angelus, qui loquebatur in me, et excitavit me quasi virum, qui excitatur de somno suo.
ZECH|4|2|Et dixit ad me: "Quid tu vides?". Et dixi: "Vidi: et ecce candelabrum aureum totum, et ampulla super caput ipsius, et septem lucernae eius super illud, et septena infusoria lucernis, quae erant super caput eius.
ZECH|4|3|Et duae olivae super illud, una a dextris ampullae et una a sinistris eius".
ZECH|4|4|Et respondi et aio ad angelum, qui loquebatur in me, dicens: "Quid sunt haec, domine mi?".
ZECH|4|5|Et respondit angelus, qui loquebatur in me, et dixit ad me: "Numquid nescis quid sunt haec?". Et dixi: "Non, domine mi".
ZECH|4|6|Et respondit et ait ad me dicens: "Hoc est verbum Domini ad Zorobabel dicens: Non in exercitu nec in robore sed in spiritu meo, dicit Dominus exercituum.
ZECH|4|7|Quis tu, mons magne, coram Zorobabel? Eris in planum. Et educet lapidem primarium inter clamores: Quam venustus!
ZECH|4|8|Et factum est verbum Domini ad me dicens:
ZECH|4|9|Manus Zorobabel fundaverunt domum istam et manus eius perficient eam, et scietis quia Dominus exercituum misit me ad vos.
ZECH|4|10|Quis enim despexit diem initiorum parvorum? Et laetabuntur et videbunt lapidem stanneum in manu Zorobabel. Septem illae oculi sunt Domini, qui discurrunt in universa terra".
ZECH|4|11|Et respondi et dixi ad eum: "Quid sunt duae olivae istae ad dexteram candelabri et ad sinistram eius?".
ZECH|4|12|Et respondi secundo et dixi ad eum: "Quid sunt duo rami olivarum, qui duabus fistulis aureis effundunt ex se aurum?".
ZECH|4|13|Et ait ad me dicens: "Numquid nescis quid sunt haec?". Et dixi: "Non, domine mi".
ZECH|4|14|Et dixit: "Isti sunt duo filii olei, qui assistunt Dominatori universae terrae".
ZECH|5|1|Et conversus sum et levavi ocu los meos et vidi: et ecce volu men volans.
ZECH|5|2|Et dixit ad me: "Quid tu vides?". Et dixi: "Ego video volumen volans; longitudo eius viginti cubitorum et latitudo eius decem cubitorum".
ZECH|5|3|Et dixit ad me: "Haec est maledictio, quae egreditur super faciem omnis terrae; quia omnis fur hinc iuxta illud expurgatur, et omnis periurus illinc iuxta illud expurgatur.
ZECH|5|4|Educo illud, dicit Dominus exercituum, et veniet ad domum furis et ad domum iurantis in nomine meo mendaciter; et commorabitur in medio domus eius, et consumet eam et ligna eius et lapides eius".
ZECH|5|5|Et egressus est angelus, qui loquebatur in me, et dixit ad me: "Leva, quaeso, oculos tuos et vide. Quid est hoc, quod egreditur?".
ZECH|5|6|Et dixi: "Quidnam est?". Et ait: "Haec est epha egrediens". Et dixit: Hoc est peccatum eorum in universa terra".
ZECH|5|7|Et ecce operculum plumbi elevatum est, et ecce mulier una sedens in medio ephae.
ZECH|5|8|Et dixit: "Haec est impietas". Et proiecit eam in epham et misit massam plumbeam in os eius.
ZECH|5|9|Et levavi oculos meos et vidi: et ecce duae mulieres egredientes, et ventus in alis earum, et habebant alas quasi alas milvi; et levaverunt epham inter terram et caelum.
ZECH|5|10|Et dixi ad angelum, qui loquebatur in me: "Quo istae deferunt epham?".
ZECH|5|11|Et dixit ad me: "Ut aedificetur ei domus in terra Sennaar; et, postquam constructa fuerit, ponetur ibi super basem suam".
ZECH|6|1|Et rursus levavi oculos meos et vidi: et ecce quattuor quadrigae egredientes de medio duorum montium; et montes, montes aerei.
ZECH|6|2|In quadriga prima equi rufi, et in quadriga secunda equi nigri,
ZECH|6|3|et in quadriga tertia equi albi, et in quadriga quarta equi varii.
ZECH|6|4|Et respondi et dixi ad angelum, qui loquebatur in me: "Quid sunt haec, domine mi?".
ZECH|6|5|Et respondit angelus et ait ad me: "Isti sunt quattuor venti caeli, qui egrediuntur, postquam steterunt coram Dominatore omnis terrae".
ZECH|6|6|In qua erant equi nigri, egrediebantur in terram aquilonis, et albi egressi sunt post eos, et varii egressi sunt ad terram austri.
ZECH|6|7|Et equi fortes exierunt et quaerebant ire et discurrere per terram. Et dixit: "Ite, perambulate terram". Et perambulaverunt terram.
ZECH|6|8|Et vocavit me et locutus est ad me dicens: "Ecce, qui egrediuntur in terram aquilonis requiescere fecerunt spiritum meum in terra aquilonis".
ZECH|6|9|Et factum est verbum Domini ad me dicens:
ZECH|6|10|"Sume ab his, qui de captivitate sunt, ab Holdai et a Thobia et ab Iedaia, et venies tu in die illa et intrabis domum Iosiae filii Sophoniae, qui venerunt de Babylone.
ZECH|6|11|Et sumes argentum et aurum et facies coronam et pones in capite Iesua filii Iosedec, sacerdotis magni,
ZECH|6|12|et loqueris ad eum dicens: Haec ait Dominus exercituum dicens: Ecce vir, Germen nomen eius; et in loco suo aliquid germinabit et aedificabit templum Domini.
ZECH|6|13|Et ipse exstruet templum Domini; et ipse portabit gloriam et sedebit et dominabitur super solio suo; et erit sacerdos ad dexteram eius, et consilium pacis erit inter illos duos.
ZECH|6|14|Et corona erit Helem et Thobiae et Iedaiae et Hen filio Sophoniae memoriale in templo Domini.
ZECH|6|15|Et qui procul sunt, venient et aedificabunt in templo Domini; et scietis quia Dominus exercituum misit me ad vos. Erit autem hoc, si oboedieritis voci Domini Dei vestri" ".
ZECH|7|1|Et factum est in anno quarto Darii regis, factum est verbum Domini ad Zachariam in quarta mensis noni, qui est Casleu.
ZECH|7|2|Et Bethel miserat Sarasar et Regemmelech et viros, qui erant cum eo, ad deprecandam faciem Domini,
ZECH|7|3|ut dicerent sacerdotibus domus Domini exercituum et prophetis loquentes: Numquid flendum est mihi in quinto mense vel ieiunandum, sicut iam feci multis annis? ".
ZECH|7|4|Et factum est verbum Domini exercituum ad me dicens:
ZECH|7|5|" Loquere ad omnem populum terrae et ad sacerdotes dicens: Cum ieiunaretis et plangeretis in quinto et septimo mense per hos septuaginta annos, numquid revera ieiunastis mihi?
ZECH|7|6|Et cum comedistis et bibistis, numquid non vobis comedistis et vobismetipsis bibistis?
ZECH|7|7|Numquid non sunt verba, quae locutus est Dominus in manu prophetarum priorum, cum adhuc Ierusalem habitaretur et esset opulenta, ipsa et urbes in circuitu eius, et Nageb habitaretur simul cum Sephela? ".
ZECH|7|8|Et factum est verbum Domini ad Zachariam dicens:
ZECH|7|9|" Haec ait Dominus exercituum dicens: Iudicium verum iudicate et misericordiam et miserationes facite unusquisque cum fratre suo;
ZECH|7|10|et viduam et pupillum et advenam et pauperem nolite calumniari, et malum unusquisque contra fratrem suum nolite cogitare in corde vestro.
ZECH|7|11|Et noluerunt attendere; et opposuerunt dorsum rebelle et aures suas aggravaverunt, ne audirent.
ZECH|7|12|Et cor suum posuerunt adamantem, ne audirent legem et verba, quae misit Dominus exercituum in spiritu suo per manum prophetarum priorum, et facta est indignatio magna a Domino exercituum.
ZECH|7|13|Et factum est, sicut cum clamaret, et ipsi non audierunt, sic clamabunt, et non exaudiam, dicit Dominus exercituum.
ZECH|7|14|Et disperdam eos per omnes gentes, quas nesciunt; et terra desolata est post eos, ita ut non esset transiens et revertens. Et posuerunt terram desiderabilem in desertum ".
ZECH|8|1|Et factum est verbum Domini exercituum dicens:
ZECH|8|2|" Haec dicit Dominus exercituum:Zelatus sum Sion zelo magnoet ardore magno zelatus sum eam.
ZECH|8|3|Haec dicit Dominus: Reversus sum ad Sion et habitabo in medio Ierusalem; et vocabitur Ierusalem civitas Veritatis, et mons Domini exercituum mons Sanctitatis.
ZECH|8|4|Haec dicit Dominus exercituum: Adhuc sedebunt senes et anus in plateis Ierusalem et unusquisque cum baculo suo in manu sua prae multitudine dierum;
ZECH|8|5|et plateae civitatis complebuntur pueris et puellis ludentibus in plateis eius.
ZECH|8|6|Haec dicit Dominus exercituum: Si videbitur difficile in oculis reliquiarum populi huius in diebus illis, numquid etiam in oculis meis difficile erit?, dicit Dominus exercituum.
ZECH|8|7|Haec dicit Dominus exercituum:Ecce ego salvabo populum meum de terra orientiset de terra occasus solis:
ZECH|8|8|et adducam eos,et habitabunt in medio Ierusalem;et erunt mihi in populum,et ego ero eis in Deumin veritate et iustitia.
ZECH|8|9|Haec dicit Dominus exercituum: Confortentur manus vestrae, qui auditis in his diebus sermones istos per os prophetarum in die, qua fundata est domus Domini exercituum, ut templum aedificaretur.
ZECH|8|10|Siquidem ante dies istosmerces hominis non erat,nec merces iumenti erat,neque introeunti neque exeuntierat pax prae tribulatione;et dimisi omnes homines,unumquemque contra proximum suum.
ZECH|8|11|Nunc autem non iuxta dies priores ego sumreliquiis populi huius,dicit Dominus exercituum;
ZECH|8|12|sed semen pacis erit:vinea dabit fructum suum,et terra dabit proventum suum,et possidere faciamreliquias populi huiusuniversa haec.
ZECH|8|13|Et erit: sicut eratis maledictio in gentibus, domus Iudae et domus Israel, sic salvabo vos, et eritis benedictio. Nolite timere; confortentur manus vestrae.
ZECH|8|14|Quia haec dicit Dominus exercituum: Sicut cogitavi, ut affligerem vos, cum ad iracundiam provocassent patres vestri me, dicit Dominus exercituum,
ZECH|8|15|et non sum misertus, sic conversus cogitavi in diebus istis, ut benefaciam Ierusalem et domui Iudae; nolite timere.
ZECH|8|16|Haec sunt ergo, quae facietis: Loquimini veritatem unusquisque cum proximo suo et iudicium pacis iudicate in portis vestris,
ZECH|8|17|et unusquisque malum contra amicum suum ne cogitetis in cordibus vestris et iuramentum mendax ne diligatis: omnia enim haec sunt quae odi, dicit Dominus.
ZECH|8|18|Et factum est verbum Domini exercituum ad me dicens:
ZECH|8|19|" Haec dicit Dominus exercituum: Ieiunium quarti et ieiunium quinti et ieiunium septimi et ieiunium decimi erit domui Iudae in gaudium et laetitiam et in sollemnitates praeclaras; veritatem tantum et pacem diligite.
ZECH|8|20|Haec dicit Dominus exercituum: Adhuc venient populi et habitatores civitatum magnarum,
ZECH|8|21|et ibunt habitatores unius ad alteram dicentes: "Eamus, ut deprecemur faciem Domini et quaeramus Dominum exercituum; vadam etiam ego".
ZECH|8|22|Et venient populi multi et gentes robustae ad quaerendum Dominum exercituum in Ierusalem et deprecandam faciem Domini.
ZECH|8|23|Haec dicit Dominus exercituum: In diebus illis apprehendent decem homines ex omnibus linguis gentium, apprehendent fimbriam viri Iudaei dicentes: "Ibimus vobiscum; audivimus enim quoniam Deus vobiscum est" ".
ZECH|9|1|Oraculum. Verbum Domini in terra Ha drachet Damasci requiei eius,quia Domini est oculus Aramsicut omnes tribus Israel.
ZECH|9|2|Emath quoque in terminis eiuset Tyrus et Sidon, quae sapiens est valde.
ZECH|9|3|Et aedificavit Tyrus munitionem suamet coacervavit argentum quasi pulveremet aurum ut lutum platearum.
ZECH|9|4|Ecce Dominus possidebit eamet percutiet in mari fortitudinem eius;et haec igni devorabitur.
ZECH|9|5|Videbit Ascalon et timebit,et Gaza dolore torquetur nimis,et Accaron, quoniam confusa est spes eius;et peribit rex de Gaza,et Ascalon non habitabitur.
ZECH|9|6|Et habitabit spurius in Azoto,et disperdam superbiam Philisthim.
ZECH|9|7|Et auferam sanguinem eius de ore eiuset abominationes eius de medio dentium eius,et relinquetur etiam ipse Deo nostro,et erit quasi dux in Iuda,et Accaron quasi Iebusaeus.
ZECH|9|8|Et circumdabo domum meam ut praesidiumcontra euntes et revertentes;et non transibit super eos ultra exactor,quia nunc vidi in oculis meis.
ZECH|9|9|Exsulta satis, filia Sion;iubila, filia Ierusalem.Ecce rex tuus venit tibiiustus et salvator ipse,pauper et sedens super asinumet super pullum filium asinae.
ZECH|9|10|Et disperdam currum ex Ephraimet equum de Ierusalem;et confringetur arcus belli,et loquetur pacem gentibus.Et imperium eius a mari usque ad mareet a flumine usque ad fines terrae.
ZECH|9|11|Tu quoque: in sanguine testamenti tuiextraho vinctos tuos de lacu,in quo non est aqua.
ZECH|9|12|Convertimini ad munitionem,vincti spei;hodie quoque annuntians:Duplicia reddam tibi.
ZECH|9|13|Nam extendi mihi Iudam quasi arcum,implevi Ephraim;et suscitabo filios tuos, Sion,super filios tuos, Graecia,et ponam te quasi gladium fortium.
ZECH|9|14|Et Dominus super eos videbitur,et exibit ut fulgur iaculum eius;et Dominus Deus in tuba canetet vadet in procellis austri.
ZECH|9|15|Dominus exercituum proteget eos;et devorabunt et conculcabunt lapides fundaeet bibent, agitabuntur quasi vinoet replebuntur ut phialae et quasi cornua altaris.
ZECH|9|16|Et salvabit eos Dominus Deus eorumin die illaut gregem populi sui,quia lapides coronaefulgebunt super terram eius.
ZECH|9|17|Quid enim bonum eius est,et quid pulchrum eius!Frumentum succrescere facit iuvenes,et mustum virgines.
ZECH|10|1|Petite a Domino pluviamin tempore pluviae serotinae.Dominus facit fulguraet pluviam imbris dabit eis,singulis herbam in agro.
ZECH|10|2|Quia theraphim loquuntur inania,et divini vident mendacium,et somnia loquuntur vana,vane consolantur;idcirco migrant quasi grex,affliguntur, quia non est eis pastor.
ZECH|10|3|Super pastores iratus est furor meus,et super hircos visitabo:certe visitat Dominus exercituumgregem suum, domum Iudae,et faciet eos quasi equum gloriae suaein bello.
ZECH|10|4|Ex ipso angulus,ex ipso paxillus,ex ipso arcus proelii,ex ipso egredietur omnis exactor simul.
ZECH|10|5|Et erunt quasi fortesconculcantes lutum viarum in proelioet bellabunt, quia Dominus cum eis; et confundentur ascensores equorum.
ZECH|10|6|Et confortabo domum Iudaeet domum Ioseph salvaboet reducam eos, quia miserebor eorum;et erunt, sicut non proiecissem eos:ego enim Dominus Deus eorum et exaudiam eos.
ZECH|10|7|Et erunt quasi fortes Ephraim,et laetabitur cor eorum quasi a vino,et filii eorum videbunt et laetabuntur,et exsultabit cor eorum in Domino.
ZECH|10|8|Sibilabo eis et congregabo illos,quia redemi eos,et multi erunt, sicut multi ante fuerant.
ZECH|10|9|Et seminabo eos in populis,et de longe recordabuntur mei;et alent filios suos et revertentur.
ZECH|10|10|Et reducam eos de terra Aegyptiet de Assyria congregabo eoset ad terram Galaad et Libani adducam eos,et non invenietur eis locus.
ZECH|10|11|Et transibunt per mare angustiae,et percutiet in mari fluctus,et exiccabuntur omnia profunda fluminis;et humiliabitur superbia Assyriae,et sceptrum Aegypti recedet.
ZECH|10|12|Confortabo eos in Domino,et in nomine eius ambulabunt ",dicit Dominus.
ZECH|11|1|Aperi, Libane, portas tuas,et comedat ignis cedros tuas.
ZECH|11|2|Ulula, abies, quia cecidit cedrus,quoniam magnifici vastati sunt;ululate, quercus Basan,quoniam corruit saltus impervius.
ZECH|11|3|Vox ululatus pastorum,quia vastata est magnificentia eorum;vox rugitus leonum,quoniam vastata est superbia Iordanis.
ZECH|11|4|Haec dicit Dominus Deus meus: " Pasce pecora occisionis.
ZECH|11|5|Quae, qui emunt, occidunt et non dolent; et, qui vendunt ea, dicunt: Benedictus Dominus! Dives factus sum". Et pastores eorum non miserentur eorum.
ZECH|11|6|Et ego non miserebor ultra super habitantes terram, dicit Dominus; ecce ego tradam homines, unumquemque in manu proximi sui et in manu regis sui; et concident terram, et non eruam de manu eorum ".
ZECH|11|7|Et ego pavi pecus occisionis pro mercatoribus gregis. Et assumpsi mihi duas virgas: unam vocavi Gratiam et alteram vocavi Funiculum; et pavi gregem.
ZECH|11|8|Et succidi tres pastores in mense uno, et taeduit eorum animam meam; siquidem et animam eorum taeduit mei.
ZECH|11|9|Et dixi: " Non pascam vos. Quae moritura est, moriatur; et, quae succidenda est, succidatur; et reliquae devorent unaquaeque carnem proximae suae ".
ZECH|11|10|Et tuli virgam meam, quae vocabatur Gratia, et abscidi eam, ut irritum facerem foedus meum, quod percussi cum omnibus populis.
ZECH|11|11|Et irritum factum est in die illa; et cognoverunt mercatores gregis, qui observabant me, quia verbum Domini est.
ZECH|11|12|Et dixi ad eos: " Si bonum est in oculis vestris, afferte mercedem meam et, si non, quiescite ". Et appenderunt mercedem meam triginta siclos argenteos.
ZECH|11|13|Et dixit Dominus ad me: " Proice illud in thesaurum, decorum pretium, quo appretiatus sum ab eis ".Et tuli triginta siclos argenteos et proieci illos in domum Domini in thesaurum.
ZECH|11|14|Et praecidi virgam meam secundam, quae appellabatur Funiculus, ut dissolverem germanitatem inter Iudam et Israel.
ZECH|11|15|Et dixit Dominus ad me: Adhuc sume tibi vasa pastoris stulti;
ZECH|11|16|quia ecce ego suscitabo pastorem in terra,qui perituram ovem non visitabit,dispersam non quaeretet contritam non sanabitet stantem non sustinebitet carnes pinguium comedetet ungulas earum confringet.
ZECH|11|17|Vae stulto meo pastoriderelinquenti gregem!Gladius super brachium eiuset super oculum dextrum eius;brachium eius ariditate siccetur,et oculus dexter eius tenebrescens obscuretur ".
ZECH|12|1|Oraculum. Verbum Domini super Israel et super Iudam. Oraculum Domini, qui extendit caelum et fundat terram et fingit spiritum hominis in eo:
ZECH|12|2|" Ecce ego pono Ierusalem pateram crapulae omnibus populis in circuitu. Hoc erit in obsidione contra Ierusalem.
ZECH|12|3|Et erit: in die illa ponam Ierusalem lapidem portandum cunctis populis; omnes portantes eam concisione lacerabuntur, et colligentur adversus eam omnes gentes terrae.
ZECH|12|4|In die illa, dicit Dominus, percutiam omnem equum in stuporem et ascensorem eius in amentiam; et super domum Iudae aperiam oculos meos et omnem equum populorum percutiam caecitate.
ZECH|12|5|Et dicent duces Iudae in corde suo: "Robur habitantium Ierusalem est in Domino exercituum, Deo eorum".
ZECH|12|6|In die illa ponam duces Iudae sicut ollam ignis super ligna et sicut facem ignis super fenum; et devorabunt ad dexteram et ad sinistram omnes populos in circuitu, et habitabitur Ierusalem rursus in loco suo.
ZECH|12|7|Et salvabit Dominus prius tabernacula Iudae, ut non elevetur gloria domus David et gloria habitantium Ierusalem contra Iudam.
ZECH|12|8|In die illa proteget Dominus habitatores Ierusalem; et erit, qui offenderit ex eis in die illa quasi David, et domus David quasi Deus, sicut angelus Domini in conspectu eorum.
ZECH|12|9|Et erit: in die illa quaeram conterere omnes gentes, quae veniunt contra Ierusalem,
ZECH|12|10|et effundam super domum David et super habitatores Ierusalem spiritum gratiae et precum; et aspicient ad me. Quem confixerunt, plangent quasi planctu super unigenitum et dolebunt super eum, ut doleri solet super primogenitum.
ZECH|12|11|In die illa magnus erit planctus in Ierusalem sicut planctus Adadremmon in campo Mageddo;
ZECH|12|12|et planget terra, singulae familiae seorsum:familia domus David seorsumet mulieres eorum seorsum;familia domus Nathan seorsumet mulieres eorum seorsum;
ZECH|12|13|familia domus Levi seorsumet mulieres eorum seorsum;familia Semei seorsumet mulieres eorum seorsum;
ZECH|12|14|omnes reliquae familiae, singulae familiae seorsumet mulieres eorum seorsum.
ZECH|13|1|In die illa erit fons patens domui David et habitantibus Ierusalem pro peccatis et immunditia.
ZECH|13|2|Et erit in die illa, dicit Dominus exercituum, disperdam nomina idolorum de terra, et non memorabuntur ultra; et pseudoprophetas et spiritum immundum auferam de terra.
ZECH|13|3|Et erit: cum prophetaverit quispiam ultra, dicent ei pater eius et mater eius, qui genuerunt eum: "Non vives, quia mendacium locutus es in nomine Domini"; et configent eum pater eius et mater eius, qui genuerunt eum, cum prophetaverit.
ZECH|13|4|Et erit: in die illa confundentur prophetae, unusquisque ex visione sua, cum prophetaverit; nec operientur pallio saccino, ut mentiantur,
ZECH|13|5|sed dicet: "Non sum propheta; homo operans terram ego sum, quoniam terra est possessio mea ab adulescentia mea".
ZECH|13|6|Et dicetur ei: "Quid sunt plagae istae in medio manuum tuarum?". Et dicet: "His plagatus sum in domo eorum, qui diligebant me".
ZECH|13|7|Framea, suscitare super pastorem meumet super virum cohaerentem mihi,dicit Dominus exercituum.Percute pastorem, et dispergentur oves,et convertam manum meam contra parvulos.
ZECH|13|8|Et erit in omni terra,dicit Dominus:partes duae in ea dispergentur et deficient,et tertia pars relinquetur in ea;
ZECH|13|9|et ducam tertiam partem per ignemet purgabo eos, sicut purgatur argentum,et probabo eos, sicut probatur aurum:ipse vocabit nomen meum,et ego exaudiam eum.Dicam: Populus meus est ille;et ipse dicet: "Dominus est Deus meus".
ZECH|14|1|Ecce venit dies Domino, et dividentur spolia tua in me dio tui,
ZECH|14|2|et congregabo omnes gentes ad Ierusalem in proelium, et capietur civitas, et vastabuntur domus, et mulieres violabuntur; et egredietur media pars civitatis in captivitatem, et reliquum populi non auferetur ex urbe.
ZECH|14|3|Et egredietur Dominus et proeliabitur contra gentes illas, sicut proeliatus est in die certaminis.
ZECH|14|4|Et stabunt pedes eius in die illa super montem Olivarum, qui est contra Ierusalem ad orientem; et scindetur mons Olivarum ex media parte sui ad orientem et ad occidentem, praerupto grandi valde, et separabitur medium montis ad aquilonem et medium eius ad meridiem.
ZECH|14|5|Et fugietis ad vallem montium eorum, quoniam vallis montium pertinget usque ad Iasol; et fugietis, sicut fugistis a facie terraemotus in diebus Oziae regis Iudae, et veniet Dominus Deus meus, omnesque sancti cum eo.
ZECH|14|6|Erit: in die illa non erit lux sed frigus et gelu;
ZECH|14|7|et erit dies una, quae nota est Domino, non dies neque nox; et in tempore vesperi erit lux.
ZECH|14|8|Et erit: in die illa exibunt aquae vivae de Ierusalem, medium earum ad mare orientale, et medium earum ad mare occidentale: in aestate et in hieme erunt.
ZECH|14|9|Et erit Dominus rex super omnem terram: in die illa erit Dominus unus, et erit nomen eius unum.
ZECH|14|10|Et revertetur omnis terra in desertum, a Gabaa usque ad Remmon ad austrum Ierusalem, quae exaltabitur et habitabitur in loco suo, a porta Beniamin usque ad locum portae Prioris, et usque ad portam Angulorum, et a turre Hananeel usque ad Torcularia regis.
ZECH|14|11|Et habitabunt in ea, et anathema non erit amplius; sed habitabitur Ierusalem secura.
ZECH|14|12|Et haec erit plaga, qua percutiet Dominus omnes gentes, quae pugnaverunt adversus Ierusalem: tabescet caro uniuscuiusque stantis super pedes suos, et oculi eius contabescent in foraminibus suis, et lingua eius contabescet in ore suo.
ZECH|14|13|In die illa erit tumultus Domini magnus in eis, et apprehendet vir manum proximi sui, et elevabitur manus eius super manum proximi sui.
ZECH|14|14|Sed et Iudas pugnabit in Ierusalem, et congregabuntur divitiae omnium gentium in circuitu, aurum et argentum et vestes multae nimis.
ZECH|14|15|Et sic erit ruina equi, muli, cameli et asini et omnium iumentorum, quae fuerint in castris illis, sicut ruina haec.
ZECH|14|16|Et omnes, qui reliqui fuerint de universis gentibus, quae venerunt contra Ierusalem, ascendent ab anno in annum, ut adorent Regem, Dominum exercituum, et celebrent festivitatem Tabernaculorum.
ZECH|14|17|Et erit: qui non ascenderit de familiis terrae ad Ierusalem, ut adoret Regem, Dominum exercituum, non erit super eos imber.
ZECH|14|18|Quod et si familia Aegypti non ascenderit et non venerit, super eos erit plaga, qua percutit Dominus gentes, quae non ascenderint ad celebrandam festivitatem Tabernaculorum.
ZECH|14|19|Haec erit poena Aegypti, et haec poena omnium gentium, quae non ascenderint ad celebrandam festivitatem Tabernaculorum.
ZECH|14|20|In die illa erit super tintinnabula equorum; "Sanctum Domino"; et erunt lebetes in domo Domini quasi phialae coram altari.
ZECH|14|21|Et erit omnis lebes in Ierusalem et in Iuda sanctificatus Domino exercituum; et venient omnes immolantes et sument ex eis et coquent in eis, et non erit mercator ultra in domo Domini exercituum in die illo ".
