JUDE|1|1|Юда, раб Ісуса Христа, а брат Якова, покликаним, улюбленим у Бозі Отці та збереженим Ісусом Христом:
JUDE|1|2|милість вам, і мир, і любов хай примножиться!
JUDE|1|3|Улюблені, всяке дбання чинивши писати до вас про наше спільне спасіння, я признав за потрібне писати до вас, благаючи боротись за віру, раз дану святим.
JUDE|1|4|Бо крадькома повходили деякі люди, на цей осуд віддавна призначені, безбожні, що благодать нашого Бога обертають у розпусту, і відкидаються єдиного Владики і Господа нашого Ісуса Христа.
JUDE|1|5|А я хочу нагадати вам, що раз усе знаєте, що Господь визволив людей від землі єгипетської, а згодом вигубив тих, хто не вірував.
JUDE|1|6|І Анголів, що не зберегли початкового стану свого, але кинули житло своє, Він зберіг у вічних кайданах під темрявою на суд великого дня.
JUDE|1|7|Як Содом і Гоморра та міста коло них, що таким самим способом чинили перелюб та ходили за іншим тілом, понесли кару вічного огню, і поставлені в приклад,
JUDE|1|8|так само буде й цим сновидам, що опоганюють тіло, погорджують владами, зневажають слави.
JUDE|1|9|І сам Архангол Михаїл, коли сперечався з дияволом і говорив про Мойсеєве тіло, не наважився винести суду зневажливого, а сказав: Хай Господь докорить тобі!
JUDE|1|10|А ці зневажають, чого не знають; а що знають із природи, як німа звірина, то й у тому псуються.
JUDE|1|11|Горе їм, бо пішли вони дорогою Каїновою, і попали в обману Валаамової заплати, і загинули в бунті Корея!
JUDE|1|12|Вони скелі підводні на ваших вечерях любови, бо з вами без страху їдять та себе попасають; хмари безводні, що носяться вітром; осінні дерева безплідні, двічі померлі, викорінені;
JUDE|1|13|люті хвилі морські, що з піною викидають власний сором; зорі блудні, що для них морок темряви бережеться повік.
JUDE|1|14|Про них же звіщав був Енох, сьомий від Адама, і казав: Ось іде Господь зо Своїми десятками тисяч святих,
JUDE|1|15|щоб суд учинити над усіма, і винуватити всіх безбожних за всі вчинки безбожности їхньої, що безбожно накоїли, та за всі жорстокі слова, що їх говорили на Нього безбожні грішники.
JUDE|1|16|Це ремствувачі, незадоволені з долі своєї, що ходять у своїх пожадливостях, а уста їхні говорять чванливе; вони вихваляють особи для зиску!
JUDE|1|17|А ви, улюблені, згадуйте слова, що їх давніше казали апостоли Господа нашого Ісуса Христа,
JUDE|1|18|які вам говорили: За останнього часу будуть глузії, що ходитимуть за своїми пожадливостями та безбожністю.
JUDE|1|19|Це ті, хто відлучується від єдности, тілесні, що духа не мають.
JUDE|1|20|А ви, улюблені, будуйте себе найсвятішою вашою вірою, моліться Духом Святим,
JUDE|1|21|бережіть себе самих у Божій любові, і чекайте милости Господа нашого Ісуса Христа для вічного життя.
JUDE|1|22|І до одних, хто вагається, будьте милостиві,
JUDE|1|23|спасайте і виривайте з огню, а до інших будьте милосердні зо страхом, і ненавидьте навіть одежу, опоганену від тіла!
JUDE|1|24|А Тому, Хто може вас зберегти від упадку, і поставити перед Своєю славою непорочними в радості,
JUDE|1|25|Єдиному премудрому Богові, Спасителеві нашому через Ісуса Христа, Господа нашого, слава, могутність, сила та влада перше всього віку, і тепер, і на всі віки! Амінь.
