LEV|1|1|The LORD called to Moses and spoke to him from the Tent of Meeting. He said,
LEV|1|2|"Speak to the Israelites and say to them: 'When any of you brings an offering to the LORD, bring as your offering an animal from either the herd or the flock.
LEV|1|3|"'If the offering is a burnt offering from the herd, he is to offer a male without defect. He must present it at the entrance to the Tent of Meeting so that it will be acceptable to the LORD.
LEV|1|4|He is to lay his hand on the head of the burnt offering, and it will be accepted on his behalf to make atonement for him.
LEV|1|5|He is to slaughter the young bull before the LORD, and then Aaron's sons the priests shall bring the blood and sprinkle it against the altar on all sides at the entrance to the Tent of Meeting.
LEV|1|6|He is to skin the burnt offering and cut it into pieces.
LEV|1|7|The sons of Aaron the priest are to put fire on the altar and arrange wood on the fire.
LEV|1|8|Then Aaron's sons the priests shall arrange the pieces, including the head and the fat, on the burning wood that is on the altar.
LEV|1|9|He is to wash the inner parts and the legs with water, and the priest is to burn all of it on the altar. It is a burnt offering, an offering made by fire, an aroma pleasing to the LORD.
LEV|1|10|"'If the offering is a burnt offering from the flock, from either the sheep or the goats, he is to offer a male without defect.
LEV|1|11|He is to slaughter it at the north side of the altar before the LORD, and Aaron's sons the priests shall sprinkle its blood against the altar on all sides.
LEV|1|12|He is to cut it into pieces, and the priest shall arrange them, including the head and the fat, on the burning wood that is on the altar.
LEV|1|13|He is to wash the inner parts and the legs with water, and the priest is to bring all of it and burn it on the altar. It is a burnt offering, an offering made by fire, an aroma pleasing to the LORD.
LEV|1|14|"'If the offering to the LORD is a burnt offering of birds, he is to offer a dove or a young pigeon.
LEV|1|15|The priest shall bring it to the altar, wring off the head and burn it on the altar; its blood shall be drained out on the side of the altar.
LEV|1|16|He is to remove the crop with its contents and throw it to the east side of the altar, where the ashes are.
LEV|1|17|He shall tear it open by the wings, not severing it completely, and then the priest shall burn it on the wood that is on the fire on the altar. It is a burnt offering, an offering made by fire, an aroma pleasing to the LORD.
LEV|2|1|"'When someone brings a grain offering to the LORD, his offering is to be of fine flour. He is to pour oil on it, put incense on it
LEV|2|2|and take it to Aaron's sons the priests. The priest shall take a handful of the fine flour and oil, together with all the incense, and burn this as a memorial portion on the altar, an offering made by fire, an aroma pleasing to the LORD.
LEV|2|3|The rest of the grain offering belongs to Aaron and his sons; it is a most holy part of the offerings made to the LORD by fire.
LEV|2|4|"'If you bring a grain offering baked in an oven, it is to consist of fine flour: cakes made without yeast and mixed with oil, or wafers made without yeast and spread with oil.
LEV|2|5|If your grain offering is prepared on a griddle, it is to be made of fine flour mixed with oil, and without yeast.
LEV|2|6|Crumble it and pour oil on it; it is a grain offering.
LEV|2|7|If your grain offering is cooked in a pan, it is to be made of fine flour and oil.
LEV|2|8|Bring the grain offering made of these things to the LORD; present it to the priest, who shall take it to the altar.
LEV|2|9|He shall take out the memorial portion from the grain offering and burn it on the altar as an offering made by fire, an aroma pleasing to the LORD.
LEV|2|10|The rest of the grain offering belongs to Aaron and his sons; it is a most holy part of the offerings made to the LORD by fire.
LEV|2|11|"'Every grain offering you bring to the LORD must be made without yeast, for you are not to burn any yeast or honey in an offering made to the LORD by fire.
LEV|2|12|You may bring them to the LORD as an offering of the firstfruits, but they are not to be offered on the altar as a pleasing aroma.
LEV|2|13|Season all your grain offerings with salt. Do not leave the salt of the covenant of your God out of your grain offerings; add salt to all your offerings.
LEV|2|14|"'If you bring a grain offering of firstfruits to the LORD, offer crushed heads of new grain roasted in the fire.
LEV|2|15|Put oil and incense on it; it is a grain offering.
LEV|2|16|The priest shall burn the memorial portion of the crushed grain and the oil, together with all the incense, as an offering made to the LORD by fire.
LEV|3|1|"'If someone's offering is a fellowship offering, and he offers an animal from the herd, whether male or female, he is to present before the LORD an animal without defect.
LEV|3|2|He is to lay his hand on the head of his offering and slaughter it at the entrance to the Tent of Meeting. Then Aaron's sons the priests shall sprinkle the blood against the altar on all sides.
LEV|3|3|From the fellowship offering he is to bring a sacrifice made to the LORD by fire: all the fat that covers the inner parts or is connected to them,
LEV|3|4|both kidneys with the fat on them near the loins, and the covering of the liver, which he will remove with the kidneys.
LEV|3|5|Then Aaron's sons are to burn it on the altar on top of the burnt offering that is on the burning wood, as an offering made by fire, an aroma pleasing to the LORD.
LEV|3|6|"'If he offers an animal from the flock as a fellowship offering to the LORD, he is to offer a male or female without defect.
LEV|3|7|If he offers a lamb, he is to present it before the LORD.
LEV|3|8|He is to lay his hand on the head of his offering and slaughter it in front of the Tent of Meeting. Then Aaron's sons shall sprinkle its blood against the altar on all sides.
LEV|3|9|From the fellowship offering he is to bring a sacrifice made to the LORD by fire: its fat, the entire fat tail cut off close to the backbone, all the fat that covers the inner parts or is connected to them,
LEV|3|10|both kidneys with the fat on them near the loins, and the covering of the liver, which he will remove with the kidneys.
LEV|3|11|The priest shall burn them on the altar as food, an offering made to the LORD by fire.
LEV|3|12|"'If his offering is a goat, he is to present it before the LORD.
LEV|3|13|He is to lay his hand on its head and slaughter it in front of the Tent of Meeting. Then Aaron's sons shall sprinkle its blood against the altar on all sides.
LEV|3|14|From what he offers he is to make this offering to the LORD by fire: all the fat that covers the inner parts or is connected to them,
LEV|3|15|both kidneys with the fat on them near the loins, and the covering of the liver, which he will remove with the kidneys.
LEV|3|16|The priest shall burn them on the altar as food, an offering made by fire, a pleasing aroma. All the fat is the LORD's.
LEV|3|17|"'This is a lasting ordinance for the generations to come, wherever you live: You must not eat any fat or any blood.'"
LEV|4|1|The LORD said to Moses,
LEV|4|2|"Say to the Israelites: 'When anyone sins unintentionally and does what is forbidden in any of the LORD's commands-
LEV|4|3|"'If the anointed priest sins, bringing guilt on the people, he must bring to the LORD a young bull without defect as a sin offering for the sin he has committed.
LEV|4|4|He is to present the bull at the entrance to the Tent of Meeting before the LORD. He is to lay his hand on its head and slaughter it before the LORD.
LEV|4|5|Then the anointed priest shall take some of the bull's blood and carry it into the Tent of Meeting.
LEV|4|6|He is to dip his finger into the blood and sprinkle some of it seven times before the LORD, in front of the curtain of the sanctuary.
LEV|4|7|The priest shall then put some of the blood on the horns of the altar of fragrant incense that is before the LORD in the Tent of Meeting. The rest of the bull's blood he shall pour out at the base of the altar of burnt offering at the entrance to the Tent of Meeting.
LEV|4|8|He shall remove all the fat from the bull of the sin offering-the fat that covers the inner parts or is connected to them,
LEV|4|9|both kidneys with the fat on them near the loins, and the covering of the liver, which he will remove with the kidneys-
LEV|4|10|just as the fat is removed from the ox sacrificed as a fellowship offering. Then the priest shall burn them on the altar of burnt offering.
LEV|4|11|But the hide of the bull and all its flesh, as well as the head and legs, the inner parts and offal-
LEV|4|12|that is, all the rest of the bull-he must take outside the camp to a place ceremonially clean, where the ashes are thrown, and burn it in a wood fire on the ash heap.
LEV|4|13|"'If the whole Israelite community sins unintentionally and does what is forbidden in any of the LORD's commands, even though the community is unaware of the matter, they are guilty.
LEV|4|14|When they become aware of the sin they committed, the assembly must bring a young bull as a sin offering and present it before the Tent of Meeting.
LEV|4|15|The elders of the community are to lay their hands on the bull's head before the LORD, and the bull shall be slaughtered before the LORD.
LEV|4|16|Then the anointed priest is to take some of the bull's blood into the Tent of Meeting.
LEV|4|17|He shall dip his finger into the blood and sprinkle it before the LORD seven times in front of the curtain.
LEV|4|18|He is to put some of the blood on the horns of the altar that is before the LORD in the Tent of Meeting. The rest of the blood he shall pour out at the base of the altar of burnt offering at the entrance to the Tent of Meeting.
LEV|4|19|He shall remove all the fat from it and burn it on the altar,
LEV|4|20|and do with this bull just as he did with the bull for the sin offering. In this way the priest will make atonement for them, and they will be forgiven.
LEV|4|21|Then he shall take the bull outside the camp and burn it as he burned the first bull. This is the sin offering for the community.
LEV|4|22|"'When a leader sins unintentionally and does what is forbidden in any of the commands of the LORD his God, he is guilty.
LEV|4|23|When he is made aware of the sin he committed, he must bring as his offering a male goat without defect.
LEV|4|24|He is to lay his hand on the goat's head and slaughter it at the place where the burnt offering is slaughtered before the LORD. It is a sin offering.
LEV|4|25|Then the priest shall take some of the blood of the sin offering with his finger and put it on the horns of the altar of burnt offering and pour out the rest of the blood at the base of the altar.
LEV|4|26|He shall burn all the fat on the altar as he burned the fat of the fellowship offering. In this way the priest will make atonement for the man's sin, and he will be forgiven.
LEV|4|27|"'If a member of the community sins unintentionally and does what is forbidden in any of the LORD's commands, he is guilty.
LEV|4|28|When he is made aware of the sin he committed, he must bring as his offering for the sin he committed a female goat without defect.
LEV|4|29|He is to lay his hand on the head of the sin offering and slaughter it at the place of the burnt offering.
LEV|4|30|Then the priest is to take some of the blood with his finger and put it on the horns of the altar of burnt offering and pour out the rest of the blood at the base of the altar.
LEV|4|31|He shall remove all the fat, just as the fat is removed from the fellowship offering, and the priest shall burn it on the altar as an aroma pleasing to the LORD. In this way the priest will make atonement for him, and he will be forgiven.
LEV|4|32|"'If he brings a lamb as his sin offering, he is to bring a female without defect.
LEV|4|33|He is to lay his hand on its head and slaughter it for a sin offering at the place where the burnt offering is slaughtered.
LEV|4|34|Then the priest shall take some of the blood of the sin offering with his finger and put it on the horns of the altar of burnt offering and pour out the rest of the blood at the base of the altar.
LEV|4|35|He shall remove all the fat, just as the fat is removed from the lamb of the fellowship offering, and the priest shall burn it on the altar on top of the offerings made to the LORD by fire. In this way the priest will make atonement for him for the sin he has committed, and he will be forgiven.
LEV|5|1|"'If a person sins because he does not speak up when he hears a public charge to testify regarding something he has seen or learned about, he will be held responsible.
LEV|5|2|"'Or if a person touches anything ceremonially unclean-whether the carcasses of unclean wild animals or of unclean livestock or of unclean creatures that move along the ground-even though he is unaware of it, he has become unclean and is guilty.
LEV|5|3|"'Or if he touches human uncleanness-anything that would make him unclean-even though he is unaware of it, when he learns of it he will be guilty.
LEV|5|4|"'Or if a person thoughtlessly takes an oath to do anything, whether good or evil-in any matter one might carelessly swear about-even though he is unaware of it, in any case when he learns of it he will be guilty.
LEV|5|5|"'When anyone is guilty in any of these ways, he must confess in what way he has sinned
LEV|5|6|and, as a penalty for the sin he has committed, he must bring to the LORD a female lamb or goat from the flock as a sin offering; and the priest shall make atonement for him for his sin.
LEV|5|7|"'If he cannot afford a lamb, he is to bring two doves or two young pigeons to the LORD as a penalty for his sin-one for a sin offering and the other for a burnt offering.
LEV|5|8|He is to bring them to the priest, who shall first offer the one for the sin offering. He is to wring its head from its neck, not severing it completely,
LEV|5|9|and is to sprinkle some of the blood of the sin offering against the side of the altar; the rest of the blood must be drained out at the base of the altar. It is a sin offering.
LEV|5|10|The priest shall then offer the other as a burnt offering in the prescribed way and make atonement for him for the sin he has committed, and he will be forgiven.
LEV|5|11|"'If, however, he cannot afford two doves or two young pigeons, he is to bring as an offering for his sin a tenth of an ephah of fine flour for a sin offering. He must not put oil or incense on it, because it is a sin offering.
LEV|5|12|He is to bring it to the priest, who shall take a handful of it as a memorial portion and burn it on the altar on top of the offerings made to the LORD by fire. It is a sin offering.
LEV|5|13|In this way the priest will make atonement for him for any of these sins he has committed, and he will be forgiven. The rest of the offering will belong to the priest, as in the case of the grain offering.'"
LEV|5|14|The LORD said to Moses:
LEV|5|15|"When a person commits a violation and sins unintentionally in regard to any of the LORD's holy things, he is to bring to the LORD as a penalty a ram from the flock, one without defect and of the proper value in silver, according to the sanctuary shekel. It is a guilt offering.
LEV|5|16|He must make restitution for what he has failed to do in regard to the holy things, add a fifth of the value to that and give it all to the priest, who will make atonement for him with the ram as a guilt offering, and he will be forgiven.
LEV|5|17|"If a person sins and does what is forbidden in any of the LORD's commands, even though he does not know it, he is guilty and will be held responsible.
LEV|5|18|He is to bring to the priest as a guilt offering a ram from the flock, one without defect and of the proper value. In this way the priest will make atonement for him for the wrong he has committed unintentionally, and he will be forgiven.
LEV|5|19|It is a guilt offering; he has been guilty of wrongdoing against the LORD."
LEV|6|1|The LORD said to Moses:
LEV|6|2|"If anyone sins and is unfaithful to the LORD by deceiving his neighbor about something entrusted to him or left in his care or stolen, or if he cheats him,
LEV|6|3|or if he finds lost property and lies about it, or if he swears falsely, or if he commits any such sin that people may do-
LEV|6|4|when he thus sins and becomes guilty, he must return what he has stolen or taken by extortion, or what was entrusted to him, or the lost property he found,
LEV|6|5|or whatever it was he swore falsely about. He must make restitution in full, add a fifth of the value to it and give it all to the owner on the day he presents his guilt offering.
LEV|6|6|And as a penalty he must bring to the priest, that is, to the LORD, his guilt offering, a ram from the flock, one without defect and of the proper value.
LEV|6|7|In this way the priest will make atonement for him before the LORD, and he will be forgiven for any of these things he did that made him guilty."
LEV|6|8|The LORD said to Moses:
LEV|6|9|"Give Aaron and his sons this command: 'These are the regulations for the burnt offering: The burnt offering is to remain on the altar hearth throughout the night, till morning, and the fire must be kept burning on the altar.
LEV|6|10|The priest shall then put on his linen clothes, with linen undergarments next to his body, and shall remove the ashes of the burnt offering that the fire has consumed on the altar and place them beside the altar.
LEV|6|11|Then he is to take off these clothes and put on others, and carry the ashes outside the camp to a place that is ceremonially clean.
LEV|6|12|The fire on the altar must be kept burning; it must not go out. Every morning the priest is to add firewood and arrange the burnt offering on the fire and burn the fat of the fellowship offerings on it.
LEV|6|13|The fire must be kept burning on the altar continuously; it must not go out.
LEV|6|14|"'These are the regulations for the grain offering: Aaron's sons are to bring it before the LORD, in front of the altar.
LEV|6|15|The priest is to take a handful of fine flour and oil, together with all the incense on the grain offering, and burn the memorial portion on the altar as an aroma pleasing to the LORD.
LEV|6|16|Aaron and his sons shall eat the rest of it, but it is to be eaten without yeast in a holy place; they are to eat it in the courtyard of the Tent of Meeting.
LEV|6|17|It must not be baked with yeast; I have given it as their share of the offerings made to me by fire. Like the sin offering and the guilt offering, it is most holy.
LEV|6|18|Any male descendant of Aaron may eat it. It is his regular share of the offerings made to the LORD by fire for the generations to come. Whatever touches them will become holy. '"
LEV|6|19|The LORD also said to Moses,
LEV|6|20|"This is the offering Aaron and his sons are to bring to the LORD on the day he is anointed: a tenth of an ephah of fine flour as a regular grain offering, half of it in the morning and half in the evening.
LEV|6|21|Prepare it with oil on a griddle; bring it well-mixed and present the grain offering broken in pieces as an aroma pleasing to the LORD.
LEV|6|22|The son who is to succeed him as anointed priest shall prepare it. It is the LORD's regular share and is to be burned completely.
LEV|6|23|Every grain offering of a priest shall be burned completely; it must not be eaten."
LEV|6|24|The LORD said to Moses,
LEV|6|25|"Say to Aaron and his sons: 'These are the regulations for the sin offering: The sin offering is to be slaughtered before the LORD in the place the burnt offering is slaughtered; it is most holy.
LEV|6|26|The priest who offers it shall eat it; it is to be eaten in a holy place, in the courtyard of the Tent of Meeting.
LEV|6|27|Whatever touches any of the flesh will become holy, and if any of the blood is spattered on a garment, you must wash it in a holy place.
LEV|6|28|The clay pot the meat is cooked in must be broken; but if it is cooked in a bronze pot, the pot is to be scoured and rinsed with water.
LEV|6|29|Any male in a priest's family may eat it; it is most holy.
LEV|6|30|But any sin offering whose blood is brought into the Tent of Meeting to make atonement in the Holy Place must not be eaten; it must be burned.
LEV|7|1|"'These are the regulations for the guilt offering, which is most holy:
LEV|7|2|The guilt offering is to be slaughtered in the place where the burnt offering is slaughtered, and its blood is to be sprinkled against the altar on all sides.
LEV|7|3|All its fat shall be offered: the fat tail and the fat that covers the inner parts,
LEV|7|4|both kidneys with the fat on them near the loins, and the covering of the liver, which is to be removed with the kidneys.
LEV|7|5|The priest shall burn them on the altar as an offering made to the LORD by fire. It is a guilt offering.
LEV|7|6|Any male in a priest's family may eat it, but it must be eaten in a holy place; it is most holy.
LEV|7|7|"'The same law applies to both the sin offering and the guilt offering: They belong to the priest who makes atonement with them.
LEV|7|8|The priest who offers a burnt offering for anyone may keep its hide for himself.
LEV|7|9|Every grain offering baked in an oven or cooked in a pan or on a griddle belongs to the priest who offers it,
LEV|7|10|and every grain offering, whether mixed with oil or dry, belongs equally to all the sons of Aaron.
LEV|7|11|"'These are the regulations for the fellowship offering a person may present to the LORD:
LEV|7|12|"'If he offers it as an expression of thankfulness, then along with this thank offering he is to offer cakes of bread made without yeast and mixed with oil, wafers made without yeast and spread with oil, and cakes of fine flour well-kneaded and mixed with oil.
LEV|7|13|Along with his fellowship offering of thanksgiving he is to present an offering with cakes of bread made with yeast.
LEV|7|14|He is to bring one of each kind as an offering, a contribution to the LORD; it belongs to the priest who sprinkles the blood of the fellowship offerings.
LEV|7|15|The meat of his fellowship offering of thanksgiving must be eaten on the day it is offered; he must leave none of it till morning.
LEV|7|16|"'If, however, his offering is the result of a vow or is a freewill offering, the sacrifice shall be eaten on the day he offers it, but anything left over may be eaten on the next day.
LEV|7|17|Any meat of the sacrifice left over till the third day must be burned up.
LEV|7|18|If any meat of the fellowship offering is eaten on the third day, it will not be accepted. It will not be credited to the one who offered it, for it is impure; the person who eats any of it will be held responsible.
LEV|7|19|"'Meat that touches anything ceremonially unclean must not be eaten; it must be burned up. As for other meat, anyone ceremonially clean may eat it.
LEV|7|20|But if anyone who is unclean eats any meat of the fellowship offering belonging to the LORD, that person must be cut off from his people.
LEV|7|21|If anyone touches something unclean-whether human uncleanness or an unclean animal or any unclean, detestable thing-and then eats any of the meat of the fellowship offering belonging to the LORD, that person must be cut off from his people.'"
LEV|7|22|The LORD said to Moses,
LEV|7|23|"Say to the Israelites: 'Do not eat any of the fat of cattle, sheep or goats.
LEV|7|24|The fat of an animal found dead or torn by wild animals may be used for any other purpose, but you must not eat it.
LEV|7|25|Anyone who eats the fat of an animal from which an offering by fire may be made to the LORD must be cut off from his people.
LEV|7|26|And wherever you live, you must not eat the blood of any bird or animal.
LEV|7|27|If anyone eats blood, that person must be cut off from his people.'"
LEV|7|28|The LORD said to Moses,
LEV|7|29|"Say to the Israelites: 'Anyone who brings a fellowship offering to the LORD is to bring part of it as his sacrifice to the LORD.
LEV|7|30|With his own hands he is to bring the offering made to the LORD by fire; he is to bring the fat, together with the breast, and wave the breast before the LORD as a wave offering.
LEV|7|31|The priest shall burn the fat on the altar, but the breast belongs to Aaron and his sons.
LEV|7|32|You are to give the right thigh of your fellowship offerings to the priest as a contribution.
LEV|7|33|The son of Aaron who offers the blood and the fat of the fellowship offering shall have the right thigh as his share.
LEV|7|34|From the fellowship offerings of the Israelites, I have taken the breast that is waved and the thigh that is presented and have given them to Aaron the priest and his sons as their regular share from the Israelites.'"
LEV|7|35|This is the portion of the offerings made to the LORD by fire that were allotted to Aaron and his sons on the day they were presented to serve the LORD as priests.
LEV|7|36|On the day they were anointed, the LORD commanded that the Israelites give this to them as their regular share for the generations to come.
LEV|7|37|These, then, are the regulations for the burnt offering, the grain offering, the sin offering, the guilt offering, the ordination offering and the fellowship offering,
LEV|7|38|which the LORD gave Moses on Mount Sinai on the day he commanded the Israelites to bring their offerings to the LORD, in the Desert of Sinai.
LEV|8|1|The LORD said to Moses,
LEV|8|2|"Bring Aaron and his sons, their garments, the anointing oil, the bull for the sin offering, the two rams and the basket containing bread made without yeast,
LEV|8|3|and gather the entire assembly at the entrance to the Tent of Meeting."
LEV|8|4|Moses did as the LORD commanded him, and the assembly gathered at the entrance to the Tent of Meeting.
LEV|8|5|Moses said to the assembly, "This is what the LORD has commanded to be done."
LEV|8|6|Then Moses brought Aaron and his sons forward and washed them with water.
LEV|8|7|He put the tunic on Aaron, tied the sash around him, clothed him with the robe and put the ephod on him. He also tied the ephod to him by its skillfully woven waistband; so it was fastened on him.
LEV|8|8|He placed the breastpiece on him and put the Urim and Thummim in the breastpiece.
LEV|8|9|Then he placed the turban on Aaron's head and set the gold plate, the sacred diadem, on the front of it, as the LORD commanded Moses.
LEV|8|10|Then Moses took the anointing oil and anointed the tabernacle and everything in it, and so consecrated them.
LEV|8|11|He sprinkled some of the oil on the altar seven times, anointing the altar and all its utensils and the basin with its stand, to consecrate them.
LEV|8|12|He poured some of the anointing oil on Aaron's head and anointed him to consecrate him.
LEV|8|13|Then he brought Aaron's sons forward, put tunics on them, tied sashes around them and put headbands on them, as the LORD commanded Moses.
LEV|8|14|He then presented the bull for the sin offering, and Aaron and his sons laid their hands on its head.
LEV|8|15|Moses slaughtered the bull and took some of the blood, and with his finger he put it on all the horns of the altar to purify the altar. He poured out the rest of the blood at the base of the altar. So he consecrated it to make atonement for it.
LEV|8|16|Moses also took all the fat around the inner parts, the covering of the liver, and both kidneys and their fat, and burned it on the altar.
LEV|8|17|But the bull with its hide and its flesh and its offal he burned up outside the camp, as the LORD commanded Moses.
LEV|8|18|He then presented the ram for the burnt offering, and Aaron and his sons laid their hands on its head.
LEV|8|19|Then Moses slaughtered the ram and sprinkled the blood against the altar on all sides.
LEV|8|20|He cut the ram into pieces and burned the head, the pieces and the fat.
LEV|8|21|He washed the inner parts and the legs with water and burned the whole ram on the altar as a burnt offering, a pleasing aroma, an offering made to the LORD by fire, as the LORD commanded Moses.
LEV|8|22|He then presented the other ram, the ram for the ordination, and Aaron and his sons laid their hands on its head.
LEV|8|23|Moses slaughtered the ram and took some of its blood and put it on the lobe of Aaron's right ear, on the thumb of his right hand and on the big toe of his right foot.
LEV|8|24|Moses also brought Aaron's sons forward and put some of the blood on the lobes of their right ears, on the thumbs of their right hands and on the big toes of their right feet. Then he sprinkled blood against the altar on all sides.
LEV|8|25|He took the fat, the fat tail, all the fat around the inner parts, the covering of the liver, both kidneys and their fat and the right thigh.
LEV|8|26|Then from the basket of bread made without yeast, which was before the LORD, he took a cake of bread, and one made with oil, and a wafer; he put these on the fat portions and on the right thigh.
LEV|8|27|He put all these in the hands of Aaron and his sons and waved them before the LORD as a wave offering.
LEV|8|28|Then Moses took them from their hands and burned them on the altar on top of the burnt offering as an ordination offering, a pleasing aroma, an offering made to the LORD by fire.
LEV|8|29|He also took the breast-Moses' share of the ordination ram-and waved it before the LORD as a wave offering, as the LORD commanded Moses.
LEV|8|30|Then Moses took some of the anointing oil and some of the blood from the altar and sprinkled them on Aaron and his garments and on his sons and their garments. So he consecrated Aaron and his garments and his sons and their garments.
LEV|8|31|Moses then said to Aaron and his sons, "Cook the meat at the entrance to the Tent of Meeting and eat it there with the bread from the basket of ordination offerings, as I commanded, saying, 'Aaron and his sons are to eat it.'
LEV|8|32|Then burn up the rest of the meat and the bread.
LEV|8|33|Do not leave the entrance to the Tent of Meeting for seven days, until the days of your ordination are completed, for your ordination will last seven days.
LEV|8|34|What has been done today was commanded by the LORD to make atonement for you.
LEV|8|35|You must stay at the entrance to the Tent of Meeting day and night for seven days and do what the LORD requires, so you will not die; for that is what I have been commanded."
LEV|8|36|So Aaron and his sons did everything the LORD commanded through Moses.
LEV|9|1|On the eighth day Moses summoned Aaron and his sons and the elders of Israel.
LEV|9|2|He said to Aaron, "Take a bull calf for your sin offering and a ram for your burnt offering, both without defect, and present them before the LORD.
LEV|9|3|Then say to the Israelites: 'Take a male goat for a sin offering, a calf and a lamb-both a year old and without defect-for a burnt offering,
LEV|9|4|and an ox and a ram for a fellowship offering to sacrifice before the LORD, together with a grain offering mixed with oil. For today the LORD will appear to you.'"
LEV|9|5|They took the things Moses commanded to the front of the Tent of Meeting, and the entire assembly came near and stood before the LORD.
LEV|9|6|Then Moses said, "This is what the LORD has commanded you to do, so that the glory of the LORD may appear to you."
LEV|9|7|Moses said to Aaron, "Come to the altar and sacrifice your sin offering and your burnt offering and make atonement for yourself and the people; sacrifice the offering that is for the people and make atonement for them, as the LORD has commanded."
LEV|9|8|So Aaron came to the altar and slaughtered the calf as a sin offering for himself.
LEV|9|9|His sons brought the blood to him, and he dipped his finger into the blood and put it on the horns of the altar; the rest of the blood he poured out at the base of the altar.
LEV|9|10|On the altar he burned the fat, the kidneys and the covering of the liver from the sin offering, as the LORD commanded Moses;
LEV|9|11|the flesh and the hide he burned up outside the camp.
LEV|9|12|Then he slaughtered the burnt offering. His sons handed him the blood, and he sprinkled it against the altar on all sides.
LEV|9|13|They handed him the burnt offering piece by piece, including the head, and he burned them on the altar.
LEV|9|14|He washed the inner parts and the legs and burned them on top of the burnt offering on the altar.
LEV|9|15|Aaron then brought the offering that was for the people. He took the goat for the people's sin offering and slaughtered it and offered it for a sin offering as he did with the first one.
LEV|9|16|He brought the burnt offering and offered it in the prescribed way.
LEV|9|17|He also brought the grain offering, took a handful of it and burned it on the altar in addition to the morning's burnt offering.
LEV|9|18|He slaughtered the ox and the ram as the fellowship offering for the people. His sons handed him the blood, and he sprinkled it against the altar on all sides.
LEV|9|19|But the fat portions of the ox and the ram-the fat tail, the layer of fat, the kidneys and the covering of the liver-
LEV|9|20|these they laid on the breasts, and then Aaron burned the fat on the altar.
LEV|9|21|Aaron waved the breasts and the right thigh before the LORD as a wave offering, as Moses commanded.
LEV|9|22|Then Aaron lifted his hands toward the people and blessed them. And having sacrificed the sin offering, the burnt offering and the fellowship offering, he stepped down.
LEV|9|23|Moses and Aaron then went into the Tent of Meeting. When they came out, they blessed the people; and the glory of the LORD appeared to all the people.
LEV|9|24|Fire came out from the presence of the LORD and consumed the burnt offering and the fat portions on the altar. And when all the people saw it, they shouted for joy and fell facedown.
LEV|10|1|Aaron's sons Nadab and Abihu took their censers, put fire in them and added incense; and they offered unauthorized fire before the LORD, contrary to his command.
LEV|10|2|So fire came out from the presence of the LORD and consumed them, and they died before the LORD.
LEV|10|3|Moses then said to Aaron, "This is what the LORD spoke of when he said: "'Among those who approach me I will show myself holy; in the sight of all the people I will be honored.'" Aaron remained silent.
LEV|10|4|Moses summoned Mishael and Elzaphan, sons of Aaron's uncle Uzziel, and said to them, "Come here; carry your cousins outside the camp, away from the front of the sanctuary."
LEV|10|5|So they came and carried them, still in their tunics, outside the camp, as Moses ordered.
LEV|10|6|Then Moses said to Aaron and his sons Eleazar and Ithamar, "Do not let your hair become unkempt, and do not tear your clothes, or you will die and the LORD will be angry with the whole community. But your relatives, all the house of Israel, may mourn for those the LORD has destroyed by fire.
LEV|10|7|Do not leave the entrance to the Tent of Meeting or you will die, because the LORD's anointing oil is on you." So they did as Moses said.
LEV|10|8|Then the LORD said to Aaron,
LEV|10|9|"You and your sons are not to drink wine or other fermented drink whenever you go into the Tent of Meeting, or you will die. This is a lasting ordinance for the generations to come.
LEV|10|10|You must distinguish between the holy and the common, between the unclean and the clean,
LEV|10|11|and you must teach the Israelites all the decrees the LORD has given them through Moses."
LEV|10|12|Moses said to Aaron and his remaining sons, Eleazar and Ithamar, "Take the grain offering left over from the offerings made to the LORD by fire and eat it prepared without yeast beside the altar, for it is most holy.
LEV|10|13|Eat it in a holy place, because it is your share and your sons' share of the offerings made to the LORD by fire; for so I have been commanded.
LEV|10|14|But you and your sons and your daughters may eat the breast that was waved and the thigh that was presented. Eat them in a ceremonially clean place; they have been given to you and your children as your share of the Israelites' fellowship offerings.
LEV|10|15|The thigh that was presented and the breast that was waved must be brought with the fat portions of the offerings made by fire, to be waved before the LORD as a wave offering. This will be the regular share for you and your children, as the LORD has commanded."
LEV|10|16|When Moses inquired about the goat of the sin offering and found that it had been burned up, he was angry with Eleazar and Ithamar, Aaron's remaining sons, and asked,
LEV|10|17|"Why didn't you eat the sin offering in the sanctuary area? It is most holy; it was given to you to take away the guilt of the community by making atonement for them before the LORD.
LEV|10|18|Since its blood was not taken into the Holy Place, you should have eaten the goat in the sanctuary area, as I commanded."
LEV|10|19|Aaron replied to Moses, "Today they sacrificed their sin offering and their burnt offering before the LORD, but such things as this have happened to me. Would the LORD have been pleased if I had eaten the sin offering today?"
LEV|10|20|When Moses heard this, he was satisfied.
LEV|11|1|The LORD said to Moses and Aaron,
LEV|11|2|"Say to the Israelites: 'Of all the animals that live on land, these are the ones you may eat:
LEV|11|3|You may eat any animal that has a split hoof completely divided and that chews the cud.
LEV|11|4|"'There are some that only chew the cud or only have a split hoof, but you must not eat them. The camel, though it chews the cud, does not have a split hoof; it is ceremonially unclean for you.
LEV|11|5|The coney, though it chews the cud, does not have a split hoof; it is unclean for you.
LEV|11|6|The rabbit, though it chews the cud, does not have a split hoof; it is unclean for you.
LEV|11|7|And the pig, though it has a split hoof completely divided, does not chew the cud; it is unclean for you.
LEV|11|8|You must not eat their meat or touch their carcasses; they are unclean for you.
LEV|11|9|"'Of all the creatures living in the water of the seas and the streams, you may eat any that have fins and scales.
LEV|11|10|But all creatures in the seas or streams that do not have fins and scales-whether among all the swarming things or among all the other living creatures in the water-you are to detest.
LEV|11|11|And since you are to detest them, you must not eat their meat and you must detest their carcasses.
LEV|11|12|Anything living in the water that does not have fins and scales is to be detestable to you.
LEV|11|13|"'These are the birds you are to detest and not eat because they are detestable: the eagle, the vulture, the black vulture,
LEV|11|14|the red kite, any kind of black kite,
LEV|11|15|any kind of raven,
LEV|11|16|the horned owl, the screech owl, the gull, any kind of hawk,
LEV|11|17|the little owl, the cormorant, the great owl,
LEV|11|18|the white owl, the desert owl, the osprey,
LEV|11|19|the stork, any kind of heron, the hoopoe and the bat.
LEV|11|20|"'All flying insects that walk on all fours are to be detestable to you.
LEV|11|21|There are, however, some winged creatures that walk on all fours that you may eat: those that have jointed legs for hopping on the ground.
LEV|11|22|Of these you may eat any kind of locust, katydid, cricket or grasshopper.
LEV|11|23|But all other winged creatures that have four legs you are to detest.
LEV|11|24|"'You will make yourselves unclean by these; whoever touches their carcasses will be unclean till evening.
LEV|11|25|Whoever picks up one of their carcasses must wash his clothes, and he will be unclean till evening.
LEV|11|26|"'Every animal that has a split hoof not completely divided or that does not chew the cud is unclean for you; whoever touches the carcass of any of them will be unclean.
LEV|11|27|Of all the animals that walk on all fours, those that walk on their paws are unclean for you; whoever touches their carcasses will be unclean till evening.
LEV|11|28|Anyone who picks up their carcasses must wash his clothes, and he will be unclean till evening. They are unclean for you.
LEV|11|29|"'Of the animals that move about on the ground, these are unclean for you: the weasel, the rat, any kind of great lizard,
LEV|11|30|the gecko, the monitor lizard, the wall lizard, the skink and the chameleon.
LEV|11|31|Of all those that move along the ground, these are unclean for you. Whoever touches them when they are dead will be unclean till evening.
LEV|11|32|When one of them dies and falls on something, that article, whatever its use, will be unclean, whether it is made of wood, cloth, hide or sackcloth. Put it in water; it will be unclean till evening, and then it will be clean.
LEV|11|33|If one of them falls into a clay pot, everything in it will be unclean, and you must break the pot.
LEV|11|34|Any food that could be eaten but has water on it from such a pot is unclean, and any liquid that could be drunk from it is unclean.
LEV|11|35|Anything that one of their carcasses falls on becomes unclean; an oven or cooking pot must be broken up. They are unclean, and you are to regard them as unclean.
LEV|11|36|A spring, however, or a cistern for collecting water remains clean, but anyone who touches one of these carcasses is unclean.
LEV|11|37|If a carcass falls on any seeds that are to be planted, they remain clean.
LEV|11|38|But if water has been put on the seed and a carcass falls on it, it is unclean for you.
LEV|11|39|"'If an animal that you are allowed to eat dies, anyone who touches the carcass will be unclean till evening.
LEV|11|40|Anyone who eats some of the carcass must wash his clothes, and he will be unclean till evening. Anyone who picks up the carcass must wash his clothes, and he will be unclean till evening.
LEV|11|41|"'Every creature that moves about on the ground is detestable; it is not to be eaten.
LEV|11|42|You are not to eat any creature that moves about on the ground, whether it moves on its belly or walks on all fours or on many feet; it is detestable.
LEV|11|43|Do not defile yourselves by any of these creatures. Do not make yourselves unclean by means of them or be made unclean by them.
LEV|11|44|I am the LORD your God; consecrate yourselves and be holy, because I am holy. Do not make yourselves unclean by any creature that moves about on the ground.
LEV|11|45|I am the LORD who brought you up out of Egypt to be your God; therefore be holy, because I am holy.
LEV|11|46|"'These are the regulations concerning animals, birds, every living thing that moves in the water and every creature that moves about on the ground.
LEV|11|47|You must distinguish between the unclean and the clean, between living creatures that may be eaten and those that may not be eaten.'"
LEV|12|1|The LORD said to Moses,
LEV|12|2|"Say to the Israelites: 'A woman who becomes pregnant and gives birth to a son will be ceremonially unclean for seven days, just as she is unclean during her monthly period.
LEV|12|3|On the eighth day the boy is to be circumcised.
LEV|12|4|Then the woman must wait thirty-three days to be purified from her bleeding. She must not touch anything sacred or go to the sanctuary until the days of her purification are over.
LEV|12|5|If she gives birth to a daughter, for two weeks the woman will be unclean, as during her period. Then she must wait sixty-six days to be purified from her bleeding.
LEV|12|6|"'When the days of her purification for a son or daughter are over, she is to bring to the priest at the entrance to the Tent of Meeting a year-old lamb for a burnt offering and a young pigeon or a dove for a sin offering.
LEV|12|7|He shall offer them before the LORD to make atonement for her, and then she will be ceremonially clean from her flow of blood. "'These are the regulations for the woman who gives birth to a boy or a girl.
LEV|12|8|If she cannot afford a lamb, she is to bring two doves or two young pigeons, one for a burnt offering and the other for a sin offering. In this way the priest will make atonement for her, and she will be clean.'"
LEV|13|1|The LORD said to Moses and Aaron,
LEV|13|2|"When anyone has a swelling or a rash or a bright spot on his skin that may become an infectious skin disease, he must be brought to Aaron the priest or to one of his sons who is a priest.
LEV|13|3|The priest is to examine the sore on his skin, and if the hair in the sore has turned white and the sore appears to be more than skin deep, it is an infectious skin disease. When the priest examines him, he shall pronounce him ceremonially unclean.
LEV|13|4|If the spot on his skin is white but does not appear to be more than skin deep and the hair in it has not turned white, the priest is to put the infected person in isolation for seven days.
LEV|13|5|On the seventh day the priest is to examine him, and if he sees that the sore is unchanged and has not spread in the skin, he is to keep him in isolation another seven days.
LEV|13|6|On the seventh day the priest is to examine him again, and if the sore has faded and has not spread in the skin, the priest shall pronounce him clean; it is only a rash. The man must wash his clothes, and he will be clean.
LEV|13|7|But if the rash does spread in his skin after he has shown himself to the priest to be pronounced clean, he must appear before the priest again.
LEV|13|8|The priest is to examine him, and if the rash has spread in the skin, he shall pronounce him unclean; it is an infectious disease.
LEV|13|9|"When anyone has an infectious skin disease, he must be brought to the priest.
LEV|13|10|The priest is to examine him, and if there is a white swelling in the skin that has turned the hair white and if there is raw flesh in the swelling,
LEV|13|11|it is a chronic skin disease and the priest shall pronounce him unclean. He is not to put him in isolation, because he is already unclean.
LEV|13|12|"If the disease breaks out all over his skin and, so far as the priest can see, it covers all the skin of the infected person from head to foot,
LEV|13|13|the priest is to examine him, and if the disease has covered his whole body, he shall pronounce that person clean. Since it has all turned white, he is clean.
LEV|13|14|But whenever raw flesh appears on him, he will be unclean.
LEV|13|15|When the priest sees the raw flesh, he shall pronounce him unclean. The raw flesh is unclean; he has an infectious disease.
LEV|13|16|Should the raw flesh change and turn white, he must go to the priest.
LEV|13|17|The priest is to examine him, and if the sores have turned white, the priest shall pronounce the infected person clean; then he will be clean.
LEV|13|18|"When someone has a boil on his skin and it heals,
LEV|13|19|and in the place where the boil was, a white swelling or reddish-white spot appears, he must present himself to the priest.
LEV|13|20|The priest is to examine it, and if it appears to be more than skin deep and the hair in it has turned white, the priest shall pronounce him unclean. It is an infectious skin disease that has broken out where the boil was.
LEV|13|21|But if, when the priest examines it, there is no white hair in it and it is not more than skin deep and has faded, then the priest is to put him in isolation for seven days.
LEV|13|22|If it is spreading in the skin, the priest shall pronounce him unclean; it is infectious.
LEV|13|23|But if the spot is unchanged and has not spread, it is only a scar from the boil, and the priest shall pronounce him clean.
LEV|13|24|"When someone has a burn on his skin and a reddish-white or white spot appears in the raw flesh of the burn,
LEV|13|25|the priest is to examine the spot, and if the hair in it has turned white, and it appears to be more than skin deep, it is an infectious disease that has broken out in the burn. The priest shall pronounce him unclean; it is an infectious skin disease.
LEV|13|26|But if the priest examines it and there is no white hair in the spot and if it is not more than skin deep and has faded, then the priest is to put him in isolation for seven days.
LEV|13|27|On the seventh day the priest is to examine him, and if it is spreading in the skin, the priest shall pronounce him unclean; it is an infectious skin disease.
LEV|13|28|If, however, the spot is unchanged and has not spread in the skin but has faded, it is a swelling from the burn, and the priest shall pronounce him clean; it is only a scar from the burn.
LEV|13|29|"If a man or woman has a sore on the head or on the chin,
LEV|13|30|the priest is to examine the sore, and if it appears to be more than skin deep and the hair in it is yellow and thin, the priest shall pronounce that person unclean; it is an itch, an infectious disease of the head or chin.
LEV|13|31|But if, when the priest examines this kind of sore, it does not seem to be more than skin deep and there is no black hair in it, then the priest is to put the infected person in isolation for seven days.
LEV|13|32|On the seventh day the priest is to examine the sore, and if the itch has not spread and there is no yellow hair in it and it does not appear to be more than skin deep,
LEV|13|33|he must be shaved except for the diseased area, and the priest is to keep him in isolation another seven days.
LEV|13|34|On the seventh day the priest is to examine the itch, and if it has not spread in the skin and appears to be no more than skin deep, the priest shall pronounce him clean. He must wash his clothes, and he will be clean.
LEV|13|35|But if the itch does spread in the skin after he is pronounced clean,
LEV|13|36|the priest is to examine him, and if the itch has spread in the skin, the priest does not need to look for yellow hair; the person is unclean.
LEV|13|37|If, however, in his judgment it is unchanged and black hair has grown in it, the itch is healed. He is clean, and the priest shall pronounce him clean.
LEV|13|38|"When a man or woman has white spots on the skin,
LEV|13|39|the priest is to examine them, and if the spots are dull white, it is a harmless rash that has broken out on the skin; that person is clean.
LEV|13|40|"When a man has lost his hair and is bald, he is clean.
LEV|13|41|If he has lost his hair from the front of his scalp and has a bald forehead, he is clean.
LEV|13|42|But if he has a reddish-white sore on his bald head or forehead, it is an infectious disease breaking out on his head or forehead.
LEV|13|43|The priest is to examine him, and if the swollen sore on his head or forehead is reddish-white like an infectious skin disease,
LEV|13|44|the man is diseased and is unclean. The priest shall pronounce him unclean because of the sore on his head.
LEV|13|45|"The person with such an infectious disease must wear torn clothes, let his hair be unkempt, cover the lower part of his face and cry out, 'Unclean! Unclean!'
LEV|13|46|As long as he has the infection he remains unclean. He must live alone; he must live outside the camp.
LEV|13|47|"If any clothing is contaminated with mildew-any woolen or linen clothing,
LEV|13|48|any woven or knitted material of linen or wool, any leather or anything made of leather-
LEV|13|49|and if the contamination in the clothing, or leather, or woven or knitted material, or any leather article, is greenish or reddish, it is a spreading mildew and must be shown to the priest.
LEV|13|50|The priest is to examine the mildew and isolate the affected article for seven days.
LEV|13|51|On the seventh day he is to examine it, and if the mildew has spread in the clothing, or the woven or knitted material, or the leather, whatever its use, it is a destructive mildew; the article is unclean.
LEV|13|52|He must burn up the clothing, or the woven or knitted material of wool or linen, or any leather article that has the contamination in it, because the mildew is destructive; the article must be burned up.
LEV|13|53|"But if, when the priest examines it, the mildew has not spread in the clothing, or the woven or knitted material, or the leather article,
LEV|13|54|he shall order that the contaminated article be washed. Then he is to isolate it for another seven days.
LEV|13|55|After the affected article has been washed, the priest is to examine it, and if the mildew has not changed its appearance, even though it has not spread, it is unclean. Burn it with fire, whether the mildew has affected one side or the other.
LEV|13|56|If, when the priest examines it, the mildew has faded after the article has been washed, he is to tear the contaminated part out of the clothing, or the leather, or the woven or knitted material.
LEV|13|57|But if it reappears in the clothing, or in the woven or knitted material, or in the leather article, it is spreading, and whatever has the mildew must be burned with fire.
LEV|13|58|The clothing, or the woven or knitted material, or any leather article that has been washed and is rid of the mildew, must be washed again, and it will be clean."
LEV|13|59|These are the regulations concerning contamination by mildew in woolen or linen clothing, woven or knitted material, or any leather article, for pronouncing them clean or unclean.
LEV|14|1|The LORD said to Moses,
LEV|14|2|"These are the regulations for the diseased person at the time of his ceremonial cleansing, when he is brought to the priest:
LEV|14|3|The priest is to go outside the camp and examine him. If the person has been healed of his infectious skin disease,
LEV|14|4|the priest shall order that two live clean birds and some cedar wood, scarlet yarn and hyssop be brought for the one to be cleansed.
LEV|14|5|Then the priest shall order that one of the birds be killed over fresh water in a clay pot.
LEV|14|6|He is then to take the live bird and dip it, together with the cedar wood, the scarlet yarn and the hyssop, into the blood of the bird that was killed over the fresh water.
LEV|14|7|Seven times he shall sprinkle the one to be cleansed of the infectious disease and pronounce him clean. Then he is to release the live bird in the open fields.
LEV|14|8|"The person to be cleansed must wash his clothes, shave off all his hair and bathe with water; then he will be ceremonially clean. After this he may come into the camp, but he must stay outside his tent for seven days.
LEV|14|9|On the seventh day he must shave off all his hair; he must shave his head, his beard, his eyebrows and the rest of his hair. He must wash his clothes and bathe himself with water, and he will be clean.
LEV|14|10|"On the eighth day he must bring two male lambs and one ewe lamb a year old, each without defect, along with three-tenths of an ephah of fine flour mixed with oil for a grain offering, and one log of oil.
LEV|14|11|The priest who pronounces him clean shall present both the one to be cleansed and his offerings before the LORD at the entrance to the Tent of Meeting.
LEV|14|12|"Then the priest is to take one of the male lambs and offer it as a guilt offering, along with the log of oil; he shall wave them before the LORD as a wave offering.
LEV|14|13|He is to slaughter the lamb in the holy place where the sin offering and the burnt offering are slaughtered. Like the sin offering, the guilt offering belongs to the priest; it is most holy.
LEV|14|14|The priest is to take some of the blood of the guilt offering and put it on the lobe of the right ear of the one to be cleansed, on the thumb of his right hand and on the big toe of his right foot.
LEV|14|15|The priest shall then take some of the log of oil, pour it in the palm of his own left hand,
LEV|14|16|dip his right forefinger into the oil in his palm, and with his finger sprinkle some of it before the LORD seven times.
LEV|14|17|The priest is to put some of the oil remaining in his palm on the lobe of the right ear of the one to be cleansed, on the thumb of his right hand and on the big toe of his right foot, on top of the blood of the guilt offering.
LEV|14|18|The rest of the oil in his palm the priest shall put on the head of the one to be cleansed and make atonement for him before the LORD.
LEV|14|19|"Then the priest is to sacrifice the sin offering and make atonement for the one to be cleansed from his uncleanness. After that, the priest shall slaughter the burnt offering
LEV|14|20|and offer it on the altar, together with the grain offering, and make atonement for him, and he will be clean.
LEV|14|21|"If, however, he is poor and cannot afford these, he must take one male lamb as a guilt offering to be waved to make atonement for him, together with a tenth of an ephah of fine flour mixed with oil for a grain offering, a log of oil,
LEV|14|22|and two doves or two young pigeons, which he can afford, one for a sin offering and the other for a burnt offering.
LEV|14|23|"On the eighth day he must bring them for his cleansing to the priest at the entrance to the Tent of Meeting, before the LORD.
LEV|14|24|The priest is to take the lamb for the guilt offering, together with the log of oil, and wave them before the LORD as a wave offering.
LEV|14|25|He shall slaughter the lamb for the guilt offering and take some of its blood and put it on the lobe of the right ear of the one to be cleansed, on the thumb of his right hand and on the big toe of his right foot.
LEV|14|26|The priest is to pour some of the oil into the palm of his own left hand,
LEV|14|27|and with his right forefinger sprinkle some of the oil from his palm seven times before the LORD.
LEV|14|28|Some of the oil in his palm he is to put on the same places he put the blood of the guilt offering-on the lobe of the right ear of the one to be cleansed, on the thumb of his right hand and on the big toe of his right foot.
LEV|14|29|The rest of the oil in his palm the priest shall put on the head of the one to be cleansed, to make atonement for him before the LORD.
LEV|14|30|Then he shall sacrifice the doves or the young pigeons, which the person can afford,
LEV|14|31|one as a sin offering and the other as a burnt offering, together with the grain offering. In this way the priest will make atonement before the LORD on behalf of the one to be cleansed."
LEV|14|32|These are the regulations for anyone who has an infectious skin disease and who cannot afford the regular offerings for his cleansing.
LEV|14|33|The LORD said to Moses and Aaron,
LEV|14|34|"When you enter the land of Canaan, which I am giving you as your possession, and I put a spreading mildew in a house in that land,
LEV|14|35|the owner of the house must go and tell the priest, 'I have seen something that looks like mildew in my house.'
LEV|14|36|The priest is to order the house to be emptied before he goes in to examine the mildew, so that nothing in the house will be pronounced unclean. After this the priest is to go in and inspect the house.
LEV|14|37|He is to examine the mildew on the walls, and if it has greenish or reddish depressions that appear to be deeper than the surface of the wall,
LEV|14|38|the priest shall go out the doorway of the house and close it up for seven days.
LEV|14|39|On the seventh day the priest shall return to inspect the house. If the mildew has spread on the walls,
LEV|14|40|he is to order that the contaminated stones be torn out and thrown into an unclean place outside the town.
LEV|14|41|He must have all the inside walls of the house scraped and the material that is scraped off dumped into an unclean place outside the town.
LEV|14|42|Then they are to take other stones to replace these and take new clay and plaster the house.
LEV|14|43|"If the mildew reappears in the house after the stones have been torn out and the house scraped and plastered,
LEV|14|44|the priest is to go and examine it and, if the mildew has spread in the house, it is a destructive mildew; the house is unclean.
LEV|14|45|It must be torn down-its stones, timbers and all the plaster-and taken out of the town to an unclean place.
LEV|14|46|"Anyone who goes into the house while it is closed up will be unclean till evening.
LEV|14|47|Anyone who sleeps or eats in the house must wash his clothes.
LEV|14|48|"But if the priest comes to examine it and the mildew has not spread after the house has been plastered, he shall pronounce the house clean, because the mildew is gone.
LEV|14|49|To purify the house he is to take two birds and some cedar wood, scarlet yarn and hyssop.
LEV|14|50|He shall kill one of the birds over fresh water in a clay pot.
LEV|14|51|Then he is to take the cedar wood, the hyssop, the scarlet yarn and the live bird, dip them into the blood of the dead bird and the fresh water, and sprinkle the house seven times.
LEV|14|52|He shall purify the house with the bird's blood, the fresh water, the live bird, the cedar wood, the hyssop and the scarlet yarn.
LEV|14|53|Then he is to release the live bird in the open fields outside the town. In this way he will make atonement for the house, and it will be clean."
LEV|14|54|These are the regulations for any infectious skin disease, for an itch,
LEV|14|55|for mildew in clothing or in a house,
LEV|14|56|and for a swelling, a rash or a bright spot,
LEV|14|57|to determine when something is clean or unclean. These are the regulations for infectious skin diseases and mildew.
LEV|15|1|The LORD said to Moses and Aaron,
LEV|15|2|"Speak to the Israelites and say to them: 'When any man has a bodily discharge, the discharge is unclean.
LEV|15|3|Whether it continues flowing from his body or is blocked, it will make him unclean. This is how his discharge will bring about uncleanness:
LEV|15|4|"'Any bed the man with a discharge lies on will be unclean, and anything he sits on will be unclean.
LEV|15|5|Anyone who touches his bed must wash his clothes and bathe with water, and he will be unclean till evening.
LEV|15|6|Whoever sits on anything that the man with a discharge sat on must wash his clothes and bathe with water, and he will be unclean till evening.
LEV|15|7|"'Whoever touches the man who has a discharge must wash his clothes and bathe with water, and he will be unclean till evening.
LEV|15|8|"'If the man with the discharge spits on someone who is clean, that person must wash his clothes and bathe with water, and he will be unclean till evening.
LEV|15|9|"'Everything the man sits on when riding will be unclean,
LEV|15|10|and whoever touches any of the things that were under him will be unclean till evening; whoever picks up those things must wash his clothes and bathe with water, and he will be unclean till evening.
LEV|15|11|"'Anyone the man with a discharge touches without rinsing his hands with water must wash his clothes and bathe with water, and he will be unclean till evening.
LEV|15|12|"'A clay pot that the man touches must be broken, and any wooden article is to be rinsed with water.
LEV|15|13|"'When a man is cleansed from his discharge, he is to count off seven days for his ceremonial cleansing; he must wash his clothes and bathe himself with fresh water, and he will be clean.
LEV|15|14|On the eighth day he must take two doves or two young pigeons and come before the LORD to the entrance to the Tent of Meeting and give them to the priest.
LEV|15|15|The priest is to sacrifice them, the one for a sin offering and the other for a burnt offering. In this way he will make atonement before the LORD for the man because of his discharge.
LEV|15|16|"'When a man has an emission of semen, he must bathe his whole body with water, and he will be unclean till evening.
LEV|15|17|Any clothing or leather that has semen on it must be washed with water, and it will be unclean till evening.
LEV|15|18|When a man lies with a woman and there is an emission of semen, both must bathe with water, and they will be unclean till evening.
LEV|15|19|"'When a woman has her regular flow of blood, the impurity of her monthly period will last seven days, and anyone who touches her will be unclean till evening.
LEV|15|20|"'Anything she lies on during her period will be unclean, and anything she sits on will be unclean.
LEV|15|21|Whoever touches her bed must wash his clothes and bathe with water, and he will be unclean till evening.
LEV|15|22|Whoever touches anything she sits on must wash his clothes and bathe with water, and he will be unclean till evening.
LEV|15|23|Whether it is the bed or anything she was sitting on, when anyone touches it, he will be unclean till evening.
LEV|15|24|"'If a man lies with her and her monthly flow touches him, he will be unclean for seven days; any bed he lies on will be unclean.
LEV|15|25|"'When a woman has a discharge of blood for many days at a time other than her monthly period or has a discharge that continues beyond her period, she will be unclean as long as she has the discharge, just as in the days of her period.
LEV|15|26|Any bed she lies on while her discharge continues will be unclean, as is her bed during her monthly period, and anything she sits on will be unclean, as during her period.
LEV|15|27|Whoever touches them will be unclean; he must wash his clothes and bathe with water, and he will be unclean till evening.
LEV|15|28|"'When she is cleansed from her discharge, she must count off seven days, and after that she will be ceremonially clean.
LEV|15|29|On the eighth day she must take two doves or two young pigeons and bring them to the priest at the entrance to the Tent of Meeting.
LEV|15|30|The priest is to sacrifice one for a sin offering and the other for a burnt offering. In this way he will make atonement for her before the LORD for the uncleanness of her discharge.
LEV|15|31|"'You must keep the Israelites separate from things that make them unclean, so they will not die in their uncleanness for defiling my dwelling place, which is among them.'"
LEV|15|32|These are the regulations for a man with a discharge, for anyone made unclean by an emission of semen,
LEV|15|33|for a woman in her monthly period, for a man or a woman with a discharge, and for a man who lies with a woman who is ceremonially unclean.
LEV|16|1|The LORD spoke to Moses after the death of the two sons of Aaron who died when they approached the LORD.
LEV|16|2|The LORD said to Moses: "Tell your brother Aaron not to come whenever he chooses into the Most Holy Place behind the curtain in front of the atonement cover on the ark, or else he will die, because I appear in the cloud over the atonement cover.
LEV|16|3|"This is how Aaron is to enter the sanctuary area: with a young bull for a sin offering and a ram for a burnt offering.
LEV|16|4|He is to put on the sacred linen tunic, with linen undergarments next to his body; he is to tie the linen sash around him and put on the linen turban. These are sacred garments; so he must bathe himself with water before he puts them on.
LEV|16|5|From the Israelite community he is to take two male goats for a sin offering and a ram for a burnt offering.
LEV|16|6|"Aaron is to offer the bull for his own sin offering to make atonement for himself and his household.
LEV|16|7|Then he is to take the two goats and present them before the LORD at the entrance to the Tent of Meeting.
LEV|16|8|He is to cast lots for the two goats-one lot for the LORD and the other for the scapegoat.
LEV|16|9|Aaron shall bring the goat whose lot falls to the LORD and sacrifice it for a sin offering.
LEV|16|10|But the goat chosen by lot as the scapegoat shall be presented alive before the LORD to be used for making atonement by sending it into the desert as a scapegoat.
LEV|16|11|"Aaron shall bring the bull for his own sin offering to make atonement for himself and his household, and he is to slaughter the bull for his own sin offering.
LEV|16|12|He is to take a censer full of burning coals from the altar before the LORD and two handfuls of finely ground fragrant incense and take them behind the curtain.
LEV|16|13|He is to put the incense on the fire before the LORD, and the smoke of the incense will conceal the atonement cover above the Testimony, so that he will not die.
LEV|16|14|He is to take some of the bull's blood and with his finger sprinkle it on the front of the atonement cover; then he shall sprinkle some of it with his finger seven times before the atonement cover.
LEV|16|15|"He shall then slaughter the goat for the sin offering for the people and take its blood behind the curtain and do with it as he did with the bull's blood: He shall sprinkle it on the atonement cover and in front of it.
LEV|16|16|In this way he will make atonement for the Most Holy Place because of the uncleanness and rebellion of the Israelites, whatever their sins have been. He is to do the same for the Tent of Meeting, which is among them in the midst of their uncleanness.
LEV|16|17|No one is to be in the Tent of Meeting from the time Aaron goes in to make atonement in the Most Holy Place until he comes out, having made atonement for himself, his household and the whole community of Israel.
LEV|16|18|"Then he shall come out to the altar that is before the LORD and make atonement for it. He shall take some of the bull's blood and some of the goat's blood and put it on all the horns of the altar.
LEV|16|19|He shall sprinkle some of the blood on it with his finger seven times to cleanse it and to consecrate it from the uncleanness of the Israelites.
LEV|16|20|"When Aaron has finished making atonement for the Most Holy Place, the Tent of Meeting and the altar, he shall bring forward the live goat.
LEV|16|21|He is to lay both hands on the head of the live goat and confess over it all the wickedness and rebellion of the Israelites-all their sins-and put them on the goat's head. He shall send the goat away into the desert in the care of a man appointed for the task.
LEV|16|22|The goat will carry on itself all their sins to a solitary place; and the man shall release it in the desert.
LEV|16|23|"Then Aaron is to go into the Tent of Meeting and take off the linen garments he put on before he entered the Most Holy Place, and he is to leave them there.
LEV|16|24|He shall bathe himself with water in a holy place and put on his regular garments. Then he shall come out and sacrifice the burnt offering for himself and the burnt offering for the people, to make atonement for himself and for the people.
LEV|16|25|He shall also burn the fat of the sin offering on the altar.
LEV|16|26|"The man who releases the goat as a scapegoat must wash his clothes and bathe himself with water; afterward he may come into the camp.
LEV|16|27|The bull and the goat for the sin offerings, whose blood was brought into the Most Holy Place to make atonement, must be taken outside the camp; their hides, flesh and offal are to be burned up.
LEV|16|28|The man who burns them must wash his clothes and bathe himself with water; afterward he may come into the camp.
LEV|16|29|"This is to be a lasting ordinance for you: On the tenth day of the seventh month you must deny yourselves and not do any work-whether native-born or an alien living among you-
LEV|16|30|because on this day atonement will be made for you, to cleanse you. Then, before the LORD, you will be clean from all your sins.
LEV|16|31|It is a sabbath of rest, and you must deny yourselves; it is a lasting ordinance.
LEV|16|32|The priest who is anointed and ordained to succeed his father as high priest is to make atonement. He is to put on the sacred linen garments
LEV|16|33|and make atonement for the Most Holy Place, for the Tent of Meeting and the altar, and for the priests and all the people of the community.
LEV|16|34|"This is to be a lasting ordinance for you: Atonement is to be made once a year for all the sins of the Israelites." And it was done, as the LORD commanded Moses.
LEV|17|1|The LORD said to Moses,
LEV|17|2|"Speak to Aaron and his sons and to all the Israelites and say to them: 'This is what the LORD has commanded:
LEV|17|3|Any Israelite who sacrifices an ox, a lamb or a goat in the camp or outside of it
LEV|17|4|instead of bringing it to the entrance to the Tent of Meeting to present it as an offering to the LORD in front of the tabernacle of the LORD -that man shall be considered guilty of bloodshed; he has shed blood and must be cut off from his people.
LEV|17|5|This is so the Israelites will bring to the LORD the sacrifices they are now making in the open fields. They must bring them to the priest, that is, to the LORD, at the entrance to the Tent of Meeting and sacrifice them as fellowship offerings.
LEV|17|6|The priest is to sprinkle the blood against the altar of the LORD at the entrance to the Tent of Meeting and burn the fat as an aroma pleasing to the LORD.
LEV|17|7|They must no longer offer any of their sacrifices to the goat idols to whom they prostitute themselves. This is to be a lasting ordinance for them and for the generations to come.'
LEV|17|8|"Say to them: 'Any Israelite or any alien living among them who offers a burnt offering or sacrifice
LEV|17|9|and does not bring it to the entrance to the Tent of Meeting to sacrifice it to the LORD -that man must be cut off from his people.
LEV|17|10|"'Any Israelite or any alien living among them who eats any blood-I will set my face against that person who eats blood and will cut him off from his people.
LEV|17|11|For the life of a creature is in the blood, and I have given it to you to make atonement for yourselves on the altar; it is the blood that makes atonement for one's life.
LEV|17|12|Therefore I say to the Israelites, "None of you may eat blood, nor may an alien living among you eat blood."
LEV|17|13|"'Any Israelite or any alien living among you who hunts any animal or bird that may be eaten must drain out the blood and cover it with earth,
LEV|17|14|because the life of every creature is its blood. That is why I have said to the Israelites, "You must not eat the blood of any creature, because the life of every creature is its blood; anyone who eats it must be cut off."
LEV|17|15|"'Anyone, whether native-born or alien, who eats anything found dead or torn by wild animals must wash his clothes and bathe with water, and he will be ceremonially unclean till evening; then he will be clean.
LEV|17|16|But if he does not wash his clothes and bathe himself, he will be held responsible.'"
LEV|18|1|The LORD said to Moses,
LEV|18|2|"Speak to the Israelites and say to them: 'I am the LORD your God.
LEV|18|3|You must not do as they do in Egypt, where you used to live, and you must not do as they do in the land of Canaan, where I am bringing you. Do not follow their practices.
LEV|18|4|You must obey my laws and be careful to follow my decrees. I am the LORD your God.
LEV|18|5|Keep my decrees and laws, for the man who obeys them will live by them. I am the LORD.
LEV|18|6|"'No one is to approach any close relative to have sexual relations. I am the LORD.
LEV|18|7|"'Do not dishonor your father by having sexual relations with your mother. She is your mother; do not have relations with her.
LEV|18|8|"'Do not have sexual relations with your father's wife; that would dishonor your father.
LEV|18|9|"'Do not have sexual relations with your sister, either your father's daughter or your mother's daughter, whether she was born in the same home or elsewhere.
LEV|18|10|"'Do not have sexual relations with your son's daughter or your daughter's daughter; that would dishonor you.
LEV|18|11|"'Do not have sexual relations with the daughter of your father's wife, born to your father; she is your sister.
LEV|18|12|"'Do not have sexual relations with your father's sister; she is your father's close relative.
LEV|18|13|"'Do not have sexual relations with your mother's sister, because she is your mother's close relative.
LEV|18|14|"'Do not dishonor your father's brother by approaching his wife to have sexual relations; she is your aunt.
LEV|18|15|"'Do not have sexual relations with your daughter-in-law. She is your son's wife; do not have relations with her.
LEV|18|16|"'Do not have sexual relations with your brother's wife; that would dishonor your brother.
LEV|18|17|"'Do not have sexual relations with both a woman and her daughter. Do not have sexual relations with either her son's daughter or her daughter's daughter; they are her close relatives. That is wickedness.
LEV|18|18|"'Do not take your wife's sister as a rival wife and have sexual relations with her while your wife is living.
LEV|18|19|"'Do not approach a woman to have sexual relations during the uncleanness of her monthly period.
LEV|18|20|"'Do not have sexual relations with your neighbor's wife and defile yourself with her.
LEV|18|21|"'Do not give any of your children to be sacrificed to Molech, for you must not profane the name of your God. I am the LORD.
LEV|18|22|"'Do not lie with a man as one lies with a woman; that is detestable.
LEV|18|23|"'Do not have sexual relations with an animal and defile yourself with it. A woman must not present herself to an animal to have sexual relations with it; that is a perversion.
LEV|18|24|"'Do not defile yourselves in any of these ways, because this is how the nations that I am going to drive out before you became defiled.
LEV|18|25|Even the land was defiled; so I punished it for its sin, and the land vomited out its inhabitants.
LEV|18|26|But you must keep my decrees and my laws. The native-born and the aliens living among you must not do any of these detestable things,
LEV|18|27|for all these things were done by the people who lived in the land before you, and the land became defiled.
LEV|18|28|And if you defile the land, it will vomit you out as it vomited out the nations that were before you.
LEV|18|29|"'Everyone who does any of these detestable things-such persons must be cut off from their people.
LEV|18|30|Keep my requirements and do not follow any of the detestable customs that were practiced before you came and do not defile yourselves with them. I am the LORD your God.'"
LEV|19|1|The LORD said to Moses,
LEV|19|2|"Speak to the entire assembly of Israel and say to them: 'Be holy because I, the LORD your God, am holy.
LEV|19|3|"'Each of you must respect his mother and father, and you must observe my Sabbaths. I am the LORD your God.
LEV|19|4|"'Do not turn to idols or make gods of cast metal for yourselves. I am the LORD your God.
LEV|19|5|"'When you sacrifice a fellowship offering to the LORD, sacrifice it in such a way that it will be accepted on your behalf.
LEV|19|6|It shall be eaten on the day you sacrifice it or on the next day; anything left over until the third day must be burned up.
LEV|19|7|If any of it is eaten on the third day, it is impure and will not be accepted.
LEV|19|8|Whoever eats it will be held responsible because he has desecrated what is holy to the LORD; that person must be cut off from his people.
LEV|19|9|"'When you reap the harvest of your land, do not reap to the very edges of your field or gather the gleanings of your harvest.
LEV|19|10|Do not go over your vineyard a second time or pick up the grapes that have fallen. Leave them for the poor and the alien. I am the LORD your God.
LEV|19|11|"'Do not steal. "'Do not lie. "'Do not deceive one another.
LEV|19|12|"'Do not swear falsely by my name and so profane the name of your God. I am the LORD.
LEV|19|13|"'Do not defraud your neighbor or rob him. "'Do not hold back the wages of a hired man overnight.
LEV|19|14|"'Do not curse the deaf or put a stumbling block in front of the blind, but fear your God. I am the LORD.
LEV|19|15|"'Do not pervert justice; do not show partiality to the poor or favoritism to the great, but judge your neighbor fairly.
LEV|19|16|"'Do not go about spreading slander among your people. "'Do not do anything that endangers your neighbor's life. I am the LORD.
LEV|19|17|"'Do not hate your brother in your heart. Rebuke your neighbor frankly so you will not share in his guilt.
LEV|19|18|"'Do not seek revenge or bear a grudge against one of your people, but love your neighbor as yourself. I am the LORD.
LEV|19|19|"'Keep my decrees. "'Do not mate different kinds of animals. "'Do not plant your field with two kinds of seed. "'Do not wear clothing woven of two kinds of material.
LEV|19|20|"'If a man sleeps with a woman who is a slave girl promised to another man but who has not been ransomed or given her freedom, there must be due punishment. Yet they are not to be put to death, because she had not been freed.
LEV|19|21|The man, however, must bring a ram to the entrance to the Tent of Meeting for a guilt offering to the LORD.
LEV|19|22|With the ram of the guilt offering the priest is to make atonement for him before the LORD for the sin he has committed, and his sin will be forgiven.
LEV|19|23|"'When you enter the land and plant any kind of fruit tree, regard its fruit as forbidden. For three years you are to consider it forbidden; it must not be eaten.
LEV|19|24|In the fourth year all its fruit will be holy, an offering of praise to the LORD.
LEV|19|25|But in the fifth year you may eat its fruit. In this way your harvest will be increased. I am the LORD your God.
LEV|19|26|"'Do not eat any meat with the blood still in it. "'Do not practice divination or sorcery.
LEV|19|27|"'Do not cut the hair at the sides of your head or clip off the edges of your beard.
LEV|19|28|"'Do not cut your bodies for the dead or put tattoo marks on yourselves. I am the LORD.
LEV|19|29|"'Do not degrade your daughter by making her a prostitute, or the land will turn to prostitution and be filled with wickedness.
LEV|19|30|"'Observe my Sabbaths and have reverence for my sanctuary. I am the LORD.
LEV|19|31|"'Do not turn to mediums or seek out spiritists, for you will be defiled by them. I am the LORD your God.
LEV|19|32|"'Rise in the presence of the aged, show respect for the elderly and revere your God. I am the LORD.
LEV|19|33|"'When an alien lives with you in your land, do not mistreat him.
LEV|19|34|The alien living with you must be treated as one of your native-born. Love him as yourself, for you were aliens in Egypt. I am the LORD your God.
LEV|19|35|"'Do not use dishonest standards when measuring length, weight or quantity.
LEV|19|36|Use honest scales and honest weights, an honest ephah and an honest hin. I am the LORD your God, who brought you out of Egypt.
LEV|19|37|"'Keep all my decrees and all my laws and follow them. I am the LORD.'"
LEV|20|1|The LORD said to Moses,
LEV|20|2|"Say to the Israelites: 'Any Israelite or any alien living in Israel who gives any of his children to Molech must be put to death. The people of the community are to stone him.
LEV|20|3|I will set my face against that man and I will cut him off from his people; for by giving his children to Molech, he has defiled my sanctuary and profaned my holy name.
LEV|20|4|If the people of the community close their eyes when that man gives one of his children to Molech and they fail to put him to death,
LEV|20|5|I will set my face against that man and his family and will cut off from their people both him and all who follow him in prostituting themselves to Molech.
LEV|20|6|"'I will set my face against the person who turns to mediums and spiritists to prostitute himself by following them, and I will cut him off from his people.
LEV|20|7|"'Consecrate yourselves and be holy, because I am the LORD your God.
LEV|20|8|Keep my decrees and follow them. I am the LORD, who makes you holy.
LEV|20|9|"'If anyone curses his father or mother, he must be put to death. He has cursed his father or his mother, and his blood will be on his own head.
LEV|20|10|"'If a man commits adultery with another man's wife-with the wife of his neighbor-both the adulterer and the adulteress must be put to death.
LEV|20|11|"'If a man sleeps with his father's wife, he has dishonored his father. Both the man and the woman must be put to death; their blood will be on their own heads.
LEV|20|12|"'If a man sleeps with his daughter-in-law, both of them must be put to death. What they have done is a perversion; their blood will be on their own heads.
LEV|20|13|"'If a man lies with a man as one lies with a woman, both of them have done what is detestable. They must be put to death; their blood will be on their own heads.
LEV|20|14|"'If a man marries both a woman and her mother, it is wicked. Both he and they must be burned in the fire, so that no wickedness will be among you.
LEV|20|15|"'If a man has sexual relations with an animal, he must be put to death, and you must kill the animal.
LEV|20|16|"'If a woman approaches an animal to have sexual relations with it, kill both the woman and the animal. They must be put to death; their blood will be on their own heads.
LEV|20|17|"'If a man marries his sister, the daughter of either his father or his mother, and they have sexual relations, it is a disgrace. They must be cut off before the eyes of their people. He has dishonored his sister and will be held responsible.
LEV|20|18|"'If a man lies with a woman during her monthly period and has sexual relations with her, he has exposed the source of her flow, and she has also uncovered it. Both of them must be cut off from their people.
LEV|20|19|"'Do not have sexual relations with the sister of either your mother or your father, for that would dishonor a close relative; both of you would be held responsible.
LEV|20|20|"'If a man sleeps with his aunt, he has dishonored his uncle. They will be held responsible; they will die childless.
LEV|20|21|"'If a man marries his brother's wife, it is an act of impurity; he has dishonored his brother. They will be childless.
LEV|20|22|"'Keep all my decrees and laws and follow them, so that the land where I am bringing you to live may not vomit you out.
LEV|20|23|You must not live according to the customs of the nations I am going to drive out before you. Because they did all these things, I abhorred them.
LEV|20|24|But I said to you, "You will possess their land; I will give it to you as an inheritance, a land flowing with milk and honey." I am the LORD your God, who has set you apart from the nations.
LEV|20|25|"'You must therefore make a distinction between clean and unclean animals and between unclean and clean birds. Do not defile yourselves by any animal or bird or anything that moves along the ground-those which I have set apart as unclean for you.
LEV|20|26|You are to be holy to me because I, the LORD, am holy, and I have set you apart from the nations to be my own.
LEV|20|27|"'A man or woman who is a medium or spiritist among you must be put to death. You are to stone them; their blood will be on their own heads.'"
LEV|21|1|The LORD said to Moses, "Speak to the priests, the sons of Aaron, and say to them: 'A priest must not make himself ceremonially unclean for any of his people who die,
LEV|21|2|except for a close relative, such as his mother or father, his son or daughter, his brother,
LEV|21|3|or an unmarried sister who is dependent on him since she has no husband-for her he may make himself unclean.
LEV|21|4|He must not make himself unclean for people related to him by marriage, and so defile himself.
LEV|21|5|"'Priests must not shave their heads or shave off the edges of their beards or cut their bodies.
LEV|21|6|They must be holy to their God and must not profane the name of their God. Because they present the offerings made to the LORD by fire, the food of their God, they are to be holy.
LEV|21|7|"'They must not marry women defiled by prostitution or divorced from their husbands, because priests are holy to their God.
LEV|21|8|Regard them as holy, because they offer up the food of your God. Consider them holy, because I the LORD am holy-I who make you holy.
LEV|21|9|"'If a priest's daughter defiles herself by becoming a prostitute, she disgraces her father; she must be burned in the fire.
LEV|21|10|"'The high priest, the one among his brothers who has had the anointing oil poured on his head and who has been ordained to wear the priestly garments, must not let his hair become unkempt or tear his clothes.
LEV|21|11|He must not enter a place where there is a dead body. He must not make himself unclean, even for his father or mother,
LEV|21|12|nor leave the sanctuary of his God or desecrate it, because he has been dedicated by the anointing oil of his God. I am the LORD.
LEV|21|13|"'The woman he marries must be a virgin.
LEV|21|14|He must not marry a widow, a divorced woman, or a woman defiled by prostitution, but only a virgin from his own people,
LEV|21|15|so he will not defile his offspring among his people. I am the LORD, who makes him holy. '"
LEV|21|16|The LORD said to Moses,
LEV|21|17|"Say to Aaron: 'For the generations to come none of your descendants who has a defect may come near to offer the food of his God.
LEV|21|18|No man who has any defect may come near: no man who is blind or lame, disfigured or deformed;
LEV|21|19|no man with a crippled foot or hand,
LEV|21|20|or who is hunchbacked or dwarfed, or who has any eye defect, or who has festering or running sores or damaged testicles.
LEV|21|21|No descendant of Aaron the priest who has any defect is to come near to present the offerings made to the LORD by fire. He has a defect; he must not come near to offer the food of his God.
LEV|21|22|He may eat the most holy food of his God, as well as the holy food;
LEV|21|23|yet because of his defect, he must not go near the curtain or approach the altar, and so desecrate my sanctuary. I am the LORD, who makes them holy. '"
LEV|21|24|So Moses told this to Aaron and his sons and to all the Israelites.
LEV|22|1|The LORD said to Moses,
LEV|22|2|"Tell Aaron and his sons to treat with respect the sacred offerings the Israelites consecrate to me, so they will not profane my holy name. I am the LORD.
LEV|22|3|"Say to them: 'For the generations to come, if any of your descendants is ceremonially unclean and yet comes near the sacred offerings that the Israelites consecrate to the LORD, that person must be cut off from my presence. I am the LORD.
LEV|22|4|"'If a descendant of Aaron has an infectious skin disease or a bodily discharge, he may not eat the sacred offerings until he is cleansed. He will also be unclean if he touches something defiled by a corpse or by anyone who has an emission of semen,
LEV|22|5|or if he touches any crawling thing that makes him unclean, or any person who makes him unclean, whatever the uncleanness may be.
LEV|22|6|The one who touches any such thing will be unclean till evening. He must not eat any of the sacred offerings unless he has bathed himself with water.
LEV|22|7|When the sun goes down, he will be clean, and after that he may eat the sacred offerings, for they are his food.
LEV|22|8|He must not eat anything found dead or torn by wild animals, and so become unclean through it. I am the LORD.
LEV|22|9|"'The priests are to keep my requirements so that they do not become guilty and die for treating them with contempt. I am the LORD, who makes them holy.
LEV|22|10|"'No one outside a priest's family may eat the sacred offering, nor may the guest of a priest or his hired worker eat it.
LEV|22|11|But if a priest buys a slave with money, or if a slave is born in his household, that slave may eat his food.
LEV|22|12|If a priest's daughter marries anyone other than a priest, she may not eat any of the sacred contributions.
LEV|22|13|But if a priest's daughter becomes a widow or is divorced, yet has no children, and she returns to live in her father's house as in her youth, she may eat of her father's food. No unauthorized person, however, may eat any of it.
LEV|22|14|"'If anyone eats a sacred offering by mistake, he must make restitution to the priest for the offering and add a fifth of the value to it.
LEV|22|15|The priests must not desecrate the sacred offerings the Israelites present to the LORD
LEV|22|16|by allowing them to eat the sacred offerings and so bring upon them guilt requiring payment. I am the LORD, who makes them holy.'"
LEV|22|17|The LORD said to Moses,
LEV|22|18|"Speak to Aaron and his sons and to all the Israelites and say to them: 'If any of you-either an Israelite or an alien living in Israel-presents a gift for a burnt offering to the LORD, either to fulfill a vow or as a freewill offering,
LEV|22|19|you must present a male without defect from the cattle, sheep or goats in order that it may be accepted on your behalf.
LEV|22|20|Do not bring anything with a defect, because it will not be accepted on your behalf.
LEV|22|21|When anyone brings from the herd or flock a fellowship offering to the LORD to fulfill a special vow or as a freewill offering, it must be without defect or blemish to be acceptable.
LEV|22|22|Do not offer to the LORD the blind, the injured or the maimed, or anything with warts or festering or running sores. Do not place any of these on the altar as an offering made to the LORD by fire.
LEV|22|23|You may, however, present as a freewill offering an ox or a sheep that is deformed or stunted, but it will not be accepted in fulfillment of a vow.
LEV|22|24|You must not offer to the LORD an animal whose testicles are bruised, crushed, torn or cut. You must not do this in your own land,
LEV|22|25|and you must not accept such animals from the hand of a foreigner and offer them as the food of your God. They will not be accepted on your behalf, because they are deformed and have defects.'"
LEV|22|26|The LORD said to Moses,
LEV|22|27|"When a calf, a lamb or a goat is born, it is to remain with its mother for seven days. From the eighth day on, it will be acceptable as an offering made to the LORD by fire.
LEV|22|28|Do not slaughter a cow or a sheep and its young on the same day.
LEV|22|29|"When you sacrifice a thank offering to the LORD, sacrifice it in such a way that it will be accepted on your behalf.
LEV|22|30|It must be eaten that same day; leave none of it till morning. I am the LORD.
LEV|22|31|"Keep my commands and follow them. I am the LORD.
LEV|22|32|Do not profane my holy name. I must be acknowledged as holy by the Israelites. I am the LORD, who makes you holy
LEV|22|33|and who brought you out of Egypt to be your God. I am the LORD."
LEV|23|1|The LORD said to Moses,
LEV|23|2|"Speak to the Israelites and say to them: 'These are my appointed feasts, the appointed feasts of the LORD, which you are to proclaim as sacred assemblies.
LEV|23|3|"'There are six days when you may work, but the seventh day is a Sabbath of rest, a day of sacred assembly. You are not to do any work; wherever you live, it is a Sabbath to the LORD.
LEV|23|4|"'These are the LORD's appointed feasts, the sacred assemblies you are to proclaim at their appointed times:
LEV|23|5|The LORD's Passover begins at twilight on the fourteenth day of the first month.
LEV|23|6|On the fifteenth day of that month the LORD's Feast of Unleavened Bread begins; for seven days you must eat bread made without yeast.
LEV|23|7|On the first day hold a sacred assembly and do no regular work.
LEV|23|8|For seven days present an offering made to the LORD by fire. And on the seventh day hold a sacred assembly and do no regular work.'"
LEV|23|9|The LORD said to Moses,
LEV|23|10|"Speak to the Israelites and say to them: 'When you enter the land I am going to give you and you reap its harvest, bring to the priest a sheaf of the first grain you harvest.
LEV|23|11|He is to wave the sheaf before the LORD so it will be accepted on your behalf; the priest is to wave it on the day after the Sabbath.
LEV|23|12|On the day you wave the sheaf, you must sacrifice as a burnt offering to the LORD a lamb a year old without defect,
LEV|23|13|together with its grain offering of two-tenths of an ephah of fine flour mixed with oil-an offering made to the LORD by fire, a pleasing aroma-and its drink offering of a quarter of a hin of wine.
LEV|23|14|You must not eat any bread, or roasted or new grain, until the very day you bring this offering to your God. This is to be a lasting ordinance for the generations to come, wherever you live.
LEV|23|15|"'From the day after the Sabbath, the day you brought the sheaf of the wave offering, count off seven full weeks.
LEV|23|16|Count off fifty days up to the day after the seventh Sabbath, and then present an offering of new grain to the LORD.
LEV|23|17|From wherever you live, bring two loaves made of two-tenths of an ephah of fine flour, baked with yeast, as a wave offering of firstfruits to the LORD.
LEV|23|18|Present with this bread seven male lambs, each a year old and without defect, one young bull and two rams. They will be a burnt offering to the LORD, together with their grain offerings and drink offerings-an offering made by fire, an aroma pleasing to the LORD.
LEV|23|19|Then sacrifice one male goat for a sin offering and two lambs, each a year old, for a fellowship offering.
LEV|23|20|The priest is to wave the two lambs before the LORD as a wave offering, together with the bread of the firstfruits. They are a sacred offering to the LORD for the priest.
LEV|23|21|On that same day you are to proclaim a sacred assembly and do no regular work. This is to be a lasting ordinance for the generations to come, wherever you live.
LEV|23|22|"'When you reap the harvest of your land, do not reap to the very edges of your field or gather the gleanings of your harvest. Leave them for the poor and the alien. I am the LORD your God.'"
LEV|23|23|The LORD said to Moses,
LEV|23|24|"Say to the Israelites: 'On the first day of the seventh month you are to have a day of rest, a sacred assembly commemorated with trumpet blasts.
LEV|23|25|Do no regular work, but present an offering made to the LORD by fire.'"
LEV|23|26|The LORD said to Moses,
LEV|23|27|"The tenth day of this seventh month is the Day of Atonement. Hold a sacred assembly and deny yourselves, and present an offering made to the LORD by fire.
LEV|23|28|Do no work on that day, because it is the Day of Atonement, when atonement is made for you before the LORD your God.
LEV|23|29|Anyone who does not deny himself on that day must be cut off from his people.
LEV|23|30|I will destroy from among his people anyone who does any work on that day.
LEV|23|31|You shall do no work at all. This is to be a lasting ordinance for the generations to come, wherever you live.
LEV|23|32|It is a sabbath of rest for you, and you must deny yourselves. From the evening of the ninth day of the month until the following evening you are to observe your sabbath."
LEV|23|33|The LORD said to Moses,
LEV|23|34|"Say to the Israelites: 'On the fifteenth day of the seventh month the LORD's Feast of Tabernacles begins, and it lasts for seven days.
LEV|23|35|The first day is a sacred assembly; do no regular work.
LEV|23|36|For seven days present offerings made to the LORD by fire, and on the eighth day hold a sacred assembly and present an offering made to the LORD by fire. It is the closing assembly; do no regular work.
LEV|23|37|("'These are the LORD's appointed feasts, which you are to proclaim as sacred assemblies for bringing offerings made to the LORD by fire-the burnt offerings and grain offerings, sacrifices and drink offerings required for each day.
LEV|23|38|These offerings are in addition to those for the LORD's Sabbaths and in addition to your gifts and whatever you have vowed and all the freewill offerings you give to the LORD.)
LEV|23|39|"'So beginning with the fifteenth day of the seventh month, after you have gathered the crops of the land, celebrate the festival to the LORD for seven days; the first day is a day of rest, and the eighth day also is a day of rest.
LEV|23|40|On the first day you are to take choice fruit from the trees, and palm fronds, leafy branches and poplars, and rejoice before the LORD your God for seven days.
LEV|23|41|Celebrate this as a festival to the LORD for seven days each year. This is to be a lasting ordinance for the generations to come; celebrate it in the seventh month.
LEV|23|42|Live in booths for seven days: All native-born Israelites are to live in booths
LEV|23|43|so your descendants will know that I had the Israelites live in booths when I brought them out of Egypt. I am the LORD your God.'"
LEV|23|44|So Moses announced to the Israelites the appointed feasts of the LORD.
LEV|24|1|The LORD said to Moses,
LEV|24|2|"Command the Israelites to bring you clear oil of pressed olives for the light so that the lamps may be kept burning continually.
LEV|24|3|Outside the curtain of the Testimony in the Tent of Meeting, Aaron is to tend the lamps before the LORD from evening till morning, continually. This is to be a lasting ordinance for the generations to come.
LEV|24|4|The lamps on the pure gold lampstand before the LORD must be tended continually.
LEV|24|5|"Take fine flour and bake twelve loaves of bread, using two-tenths of an ephah for each loaf.
LEV|24|6|Set them in two rows, six in each row, on the table of pure gold before the LORD.
LEV|24|7|Along each row put some pure incense as a memorial portion to represent the bread and to be an offering made to the LORD by fire.
LEV|24|8|This bread is to be set out before the LORD regularly, Sabbath after Sabbath, on behalf of the Israelites, as a lasting covenant.
LEV|24|9|It belongs to Aaron and his sons, who are to eat it in a holy place, because it is a most holy part of their regular share of the offerings made to the LORD by fire." A Blasphemer Stoned
LEV|24|10|Now the son of an Israelite mother and an Egyptian father went out among the Israelites, and a fight broke out in the camp between him and an Israelite.
LEV|24|11|The son of the Israelite woman blasphemed the Name with a curse; so they brought him to Moses. (His mother's name was Shelomith, the daughter of Dibri the Danite.)
LEV|24|12|They put him in custody until the will of the LORD should be made clear to them.
LEV|24|13|Then the LORD said to Moses:
LEV|24|14|"Take the blasphemer outside the camp. All those who heard him are to lay their hands on his head, and the entire assembly is to stone him.
LEV|24|15|Say to the Israelites: 'If anyone curses his God, he will be held responsible;
LEV|24|16|anyone who blasphemes the name of the LORD must be put to death. The entire assembly must stone him. Whether an alien or native-born, when he blasphemes the Name, he must be put to death.
LEV|24|17|"'If anyone takes the life of a human being, he must be put to death.
LEV|24|18|Anyone who takes the life of someone's animal must make restitution-life for life.
LEV|24|19|If anyone injures his neighbor, whatever he has done must be done to him:
LEV|24|20|fracture for fracture, eye for eye, tooth for tooth. As he has injured the other, so he is to be injured.
LEV|24|21|Whoever kills an animal must make restitution, but whoever kills a man must be put to death.
LEV|24|22|You are to have the same law for the alien and the native-born. I am the LORD your God.'"
LEV|24|23|Then Moses spoke to the Israelites, and they took the blasphemer outside the camp and stoned him. The Israelites did as the LORD commanded Moses.
LEV|25|1|The LORD said to Moses on Mount Sinai,
LEV|25|2|"Speak to the Israelites and say to them: 'When you enter the land I am going to give you, the land itself must observe a sabbath to the LORD.
LEV|25|3|For six years sow your fields, and for six years prune your vineyards and gather their crops.
LEV|25|4|But in the seventh year the land is to have a sabbath of rest, a sabbath to the LORD. Do not sow your fields or prune your vineyards.
LEV|25|5|Do not reap what grows of itself or harvest the grapes of your untended vines. The land is to have a year of rest.
LEV|25|6|Whatever the land yields during the sabbath year will be food for you-for yourself, your manservant and maidservant, and the hired worker and temporary resident who live among you,
LEV|25|7|as well as for your livestock and the wild animals in your land. Whatever the land produces may be eaten.
LEV|25|8|"'Count off seven sabbaths of years-seven times seven years-so that the seven sabbaths of years amount to a period of forty-nine years.
LEV|25|9|Then have the trumpet sounded everywhere on the tenth day of the seventh month; on the Day of Atonement sound the trumpet throughout your land.
LEV|25|10|Consecrate the fiftieth year and proclaim liberty throughout the land to all its inhabitants. It shall be a jubilee for you; each one of you is to return to his family property and each to his own clan.
LEV|25|11|The fiftieth year shall be a jubilee for you; do not sow and do not reap what grows of itself or harvest the untended vines.
LEV|25|12|For it is a jubilee and is to be holy for you; eat only what is taken directly from the fields.
LEV|25|13|"'In this Year of Jubilee everyone is to return to his own property.
LEV|25|14|"'If you sell land to one of your countrymen or buy any from him, do not take advantage of each other.
LEV|25|15|You are to buy from your countryman on the basis of the number of years since the Jubilee. And he is to sell to you on the basis of the number of years left for harvesting crops.
LEV|25|16|When the years are many, you are to increase the price, and when the years are few, you are to decrease the price, because what he is really selling you is the number of crops.
LEV|25|17|Do not take advantage of each other, but fear your God. I am the LORD your God.
LEV|25|18|"'Follow my decrees and be careful to obey my laws, and you will live safely in the land.
LEV|25|19|Then the land will yield its fruit, and you will eat your fill and live there in safety.
LEV|25|20|You may ask, "What will we eat in the seventh year if we do not plant or harvest our crops?"
LEV|25|21|I will send you such a blessing in the sixth year that the land will yield enough for three years.
LEV|25|22|While you plant during the eighth year, you will eat from the old crop and will continue to eat from it until the harvest of the ninth year comes in.
LEV|25|23|"'The land must not be sold permanently, because the land is mine and you are but aliens and my tenants.
LEV|25|24|Throughout the country that you hold as a possession, you must provide for the redemption of the land.
LEV|25|25|"'If one of your countrymen becomes poor and sells some of his property, his nearest relative is to come and redeem what his countryman has sold.
LEV|25|26|If, however, a man has no one to redeem it for him but he himself prospers and acquires sufficient means to redeem it,
LEV|25|27|he is to determine the value for the years since he sold it and refund the balance to the man to whom he sold it; he can then go back to his own property.
LEV|25|28|But if he does not acquire the means to repay him, what he sold will remain in the possession of the buyer until the Year of Jubilee. It will be returned in the Jubilee, and he can then go back to his property.
LEV|25|29|"'If a man sells a house in a walled city, he retains the right of redemption a full year after its sale. During that time he may redeem it.
LEV|25|30|If it is not redeemed before a full year has passed, the house in the walled city shall belong permanently to the buyer and his descendants. It is not to be returned in the Jubilee.
LEV|25|31|But houses in villages without walls around them are to be considered as open country. They can be redeemed, and they are to be returned in the Jubilee.
LEV|25|32|"'The Levites always have the right to redeem their houses in the Levitical towns, which they possess.
LEV|25|33|So the property of the Levites is redeemable-that is, a house sold in any town they hold-and is to be returned in the Jubilee, because the houses in the towns of the Levites are their property among the Israelites.
LEV|25|34|But the pastureland belonging to their towns must not be sold; it is their permanent possession.
LEV|25|35|"'If one of your countrymen becomes poor and is unable to support himself among you, help him as you would an alien or a temporary resident, so he can continue to live among you.
LEV|25|36|Do not take interest of any kind from him, but fear your God, so that your countryman may continue to live among you.
LEV|25|37|You must not lend him money at interest or sell him food at a profit.
LEV|25|38|I am the LORD your God, who brought you out of Egypt to give you the land of Canaan and to be your God.
LEV|25|39|"'If one of your countrymen becomes poor among you and sells himself to you, do not make him work as a slave.
LEV|25|40|He is to be treated as a hired worker or a temporary resident among you; he is to work for you until the Year of Jubilee.
LEV|25|41|Then he and his children are to be released, and he will go back to his own clan and to the property of his forefathers.
LEV|25|42|Because the Israelites are my servants, whom I brought out of Egypt, they must not be sold as slaves.
LEV|25|43|Do not rule over them ruthlessly, but fear your God.
LEV|25|44|"'Your male and female slaves are to come from the nations around you; from them you may buy slaves.
LEV|25|45|You may also buy some of the temporary residents living among you and members of their clans born in your country, and they will become your property.
LEV|25|46|You can will them to your children as inherited property and can make them slaves for life, but you must not rule over your fellow Israelites ruthlessly.
LEV|25|47|"'If an alien or a temporary resident among you becomes rich and one of your countrymen becomes poor and sells himself to the alien living among you or to a member of the alien's clan,
LEV|25|48|he retains the right of redemption after he has sold himself. One of his relatives may redeem him:
LEV|25|49|An uncle or a cousin or any blood relative in his clan may redeem him. Or if he prospers, he may redeem himself.
LEV|25|50|He and his buyer are to count the time from the year he sold himself up to the Year of Jubilee. The price for his release is to be based on the rate paid to a hired man for that number of years.
LEV|25|51|If many years remain, he must pay for his redemption a larger share of the price paid for him.
LEV|25|52|If only a few years remain until the Year of Jubilee, he is to compute that and pay for his redemption accordingly.
LEV|25|53|He is to be treated as a man hired from year to year; you must see to it that his owner does not rule over him ruthlessly.
LEV|25|54|"'Even if he is not redeemed in any of these ways, he and his children are to be released in the Year of Jubilee,
LEV|25|55|for the Israelites belong to me as servants. They are my servants, whom I brought out of Egypt. I am the LORD your God.
LEV|26|1|"'Do not make idols or set up an image or a sacred stone for yourselves, and do not place a carved stone in your land to bow down before it. I am the LORD your God.
LEV|26|2|"'Observe my Sabbaths and have reverence for my sanctuary. I am the LORD.
LEV|26|3|"'If you follow my decrees and are careful to obey my commands,
LEV|26|4|I will send you rain in its season, and the ground will yield its crops and the trees of the field their fruit.
LEV|26|5|Your threshing will continue until grape harvest and the grape harvest will continue until planting, and you will eat all the food you want and live in safety in your land.
LEV|26|6|"'I will grant peace in the land, and you will lie down and no one will make you afraid. I will remove savage beasts from the land, and the sword will not pass through your country.
LEV|26|7|You will pursue your enemies, and they will fall by the sword before you.
LEV|26|8|Five of you will chase a hundred, and a hundred of you will chase ten thousand, and your enemies will fall by the sword before you.
LEV|26|9|"'I will look on you with favor and make you fruitful and increase your numbers, and I will keep my covenant with you.
LEV|26|10|You will still be eating last year's harvest when you will have to move it out to make room for the new.
LEV|26|11|I will put my dwelling place among you, and I will not abhor you.
LEV|26|12|I will walk among you and be your God, and you will be my people.
LEV|26|13|I am the LORD your God, who brought you out of Egypt so that you would no longer be slaves to the Egyptians; I broke the bars of your yoke and enabled you to walk with heads held high.
LEV|26|14|"'But if you will not listen to me and carry out all these commands,
LEV|26|15|and if you reject my decrees and abhor my laws and fail to carry out all my commands and so violate my covenant,
LEV|26|16|then I will do this to you: I will bring upon you sudden terror, wasting diseases and fever that will destroy your sight and drain away your life. You will plant seed in vain, because your enemies will eat it.
LEV|26|17|I will set my face against you so that you will be defeated by your enemies; those who hate you will rule over you, and you will flee even when no one is pursuing you.
LEV|26|18|"'If after all this you will not listen to me, I will punish you for your sins seven times over.
LEV|26|19|I will break down your stubborn pride and make the sky above you like iron and the ground beneath you like bronze.
LEV|26|20|Your strength will be spent in vain, because your soil will not yield its crops, nor will the trees of the land yield their fruit.
LEV|26|21|"'If you remain hostile toward me and refuse to listen to me, I will multiply your afflictions seven times over, as your sins deserve.
LEV|26|22|I will send wild animals against you, and they will rob you of your children, destroy your cattle and make you so few in number that your roads will be deserted.
LEV|26|23|"'If in spite of these things you do not accept my correction but continue to be hostile toward me,
LEV|26|24|I myself will be hostile toward you and will afflict you for your sins seven times over.
LEV|26|25|And I will bring the sword upon you to avenge the breaking of the covenant. When you withdraw into your cities, I will send a plague among you, and you will be given into enemy hands.
LEV|26|26|When I cut off your supply of bread, ten women will be able to bake your bread in one oven, and they will dole out the bread by weight. You will eat, but you will not be satisfied.
LEV|26|27|"'If in spite of this you still do not listen to me but continue to be hostile toward me,
LEV|26|28|then in my anger I will be hostile toward you, and I myself will punish you for your sins seven times over.
LEV|26|29|You will eat the flesh of your sons and the flesh of your daughters.
LEV|26|30|I will destroy your high places, cut down your incense altars and pile your dead bodies on the lifeless forms of your idols, and I will abhor you.
LEV|26|31|I will turn your cities into ruins and lay waste your sanctuaries, and I will take no delight in the pleasing aroma of your offerings.
LEV|26|32|I will lay waste the land, so that your enemies who live there will be appalled.
LEV|26|33|I will scatter you among the nations and will draw out my sword and pursue you. Your land will be laid waste, and your cities will lie in ruins.
LEV|26|34|Then the land will enjoy its sabbath years all the time that it lies desolate and you are in the country of your enemies; then the land will rest and enjoy its sabbaths.
LEV|26|35|All the time that it lies desolate, the land will have the rest it did not have during the sabbaths you lived in it.
LEV|26|36|"'As for those of you who are left, I will make their hearts so fearful in the lands of their enemies that the sound of a windblown leaf will put them to flight. They will run as though fleeing from the sword, and they will fall, even though no one is pursuing them.
LEV|26|37|They will stumble over one another as though fleeing from the sword, even though no one is pursuing them. So you will not be able to stand before your enemies.
LEV|26|38|You will perish among the nations; the land of your enemies will devour you.
LEV|26|39|Those of you who are left will waste away in the lands of their enemies because of their sins; also because of their fathers' sins they will waste away.
LEV|26|40|"'But if they will confess their sins and the sins of their fathers-their treachery against me and their hostility toward me,
LEV|26|41|which made me hostile toward them so that I sent them into the land of their enemies-then when their uncircumcised hearts are humbled and they pay for their sin,
LEV|26|42|I will remember my covenant with Jacob and my covenant with Isaac and my covenant with Abraham, and I will remember the land.
LEV|26|43|For the land will be deserted by them and will enjoy its sabbaths while it lies desolate without them. They will pay for their sins because they rejected my laws and abhorred my decrees.
LEV|26|44|Yet in spite of this, when they are in the land of their enemies, I will not reject them or abhor them so as to destroy them completely, breaking my covenant with them. I am the LORD their God.
LEV|26|45|But for their sake I will remember the covenant with their ancestors whom I brought out of Egypt in the sight of the nations to be their God. I am the LORD.'"
LEV|26|46|These are the decrees, the laws and the regulations that the LORD established on Mount Sinai between himself and the Israelites through Moses.
LEV|27|1|The LORD said to Moses,
LEV|27|2|"Speak to the Israelites and say to them: 'If anyone makes a special vow to dedicate persons to the LORD by giving equivalent values,
LEV|27|3|set the value of a male between the ages of twenty and sixty at fifty shekels of silver, according to the sanctuary shekel;
LEV|27|4|and if it is a female, set her value at thirty shekels.
LEV|27|5|If it is a person between the ages of five and twenty, set the value of a male at twenty shekels and of a female at ten shekels.
LEV|27|6|If it is a person between one month and five years, set the value of a male at five shekels of silver and that of a female at three shekels of silver.
LEV|27|7|If it is a person sixty years old or more, set the value of a male at fifteen shekels and of a female at ten shekels.
LEV|27|8|If anyone making the vow is too poor to pay the specified amount, he is to present the person to the priest, who will set the value for him according to what the man making the vow can afford.
LEV|27|9|"'If what he vowed is an animal that is acceptable as an offering to the LORD, such an animal given to the LORD becomes holy.
LEV|27|10|He must not exchange it or substitute a good one for a bad one, or a bad one for a good one; if he should substitute one animal for another, both it and the substitute become holy.
LEV|27|11|If what he vowed is a ceremonially unclean animal-one that is not acceptable as an offering to the LORD -the animal must be presented to the priest,
LEV|27|12|who will judge its quality as good or bad. Whatever value the priest then sets, that is what it will be.
LEV|27|13|If the owner wishes to redeem the animal, he must add a fifth to its value.
LEV|27|14|"'If a man dedicates his house as something holy to the LORD, the priest will judge its quality as good or bad. Whatever value the priest then sets, so it will remain.
LEV|27|15|If the man who dedicates his house redeems it, he must add a fifth to its value, and the house will again become his.
LEV|27|16|"'If a man dedicates to the LORD part of his family land, its value is to be set according to the amount of seed required for it-fifty shekels of silver to a homer of barley seed.
LEV|27|17|If he dedicates his field during the Year of Jubilee, the value that has been set remains.
LEV|27|18|But if he dedicates his field after the Jubilee, the priest will determine the value according to the number of years that remain until the next Year of Jubilee, and its set value will be reduced.
LEV|27|19|If the man who dedicates the field wishes to redeem it, he must add a fifth to its value, and the field will again become his.
LEV|27|20|If, however, he does not redeem the field, or if he has sold it to someone else, it can never be redeemed.
LEV|27|21|When the field is released in the Jubilee, it will become holy, like a field devoted to the LORD; it will become the property of the priests.
LEV|27|22|"'If a man dedicates to the LORD a field he has bought, which is not part of his family land,
LEV|27|23|the priest will determine its value up to the Year of Jubilee, and the man must pay its value on that day as something holy to the LORD.
LEV|27|24|In the Year of Jubilee the field will revert to the person from whom he bought it, the one whose land it was.
LEV|27|25|Every value is to be set according to the sanctuary shekel, twenty gerahs to the shekel.
LEV|27|26|"'No one, however, may dedicate the firstborn of an animal, since the firstborn already belongs to the LORD; whether an ox or a sheep, it is the LORD's.
LEV|27|27|If it is one of the unclean animals, he may buy it back at its set value, adding a fifth of the value to it. If he does not redeem it, it is to be sold at its set value.
LEV|27|28|"'But nothing that a man owns and devotes to the LORD -whether man or animal or family land-may be sold or redeemed; everything so devoted is most holy to the LORD.
LEV|27|29|"'No person devoted to destruction may be ransomed; he must be put to death.
LEV|27|30|"'A tithe of everything from the land, whether grain from the soil or fruit from the trees, belongs to the LORD; it is holy to the LORD.
LEV|27|31|If a man redeems any of his tithe, he must add a fifth of the value to it.
LEV|27|32|The entire tithe of the herd and flock-every tenth animal that passes under the shepherd's rod-will be holy to the LORD.
LEV|27|33|He must not pick out the good from the bad or make any substitution. If he does make a substitution, both the animal and its substitute become holy and cannot be redeemed.'"
LEV|27|34|These are the commands the LORD gave Moses on Mount Sinai for the Israelites.
