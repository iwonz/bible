1TIM|1|1|Павло, апостол Христа Ісуса, з волі Бога, Спасителя нашого й Христа Ісуса, надії нашої,
1TIM|1|2|до Тимофія, щирого сина за вірою: благодать, милість, мир від Бога Отця і Христа Ісуса, Господа нашого!
1TIM|1|3|Як я йшов у Македонію, я тебе вблагав був позостатися в Ефесі, щоб ти декому наказав не навчати іншої науки,
1TIM|1|4|і не звертати уваги на вигадки й на родоводи безкраї, що викликують більше сварки, ніж збудування Боже, що в вірі воно.
1TIM|1|5|Ціль же наказу любов від чистого серця, і доброго сумління, і нелукавої віри.
1TIM|1|6|Дехто в тім прогрішили були та вдалися в пустомовність,
1TIM|1|7|вони забажали бути вчителями Закону, та не розуміли ні того, що говорять, ні про що запевняють.
1TIM|1|8|А ми знаємо, що добрий Закон, коли хто законно вживає його,
1TIM|1|9|та відає те, що Закон не покладений для праведного, але для беззаконних та для неслухняних, нечестивих і грішників, безбожних та нечистих, для зневажників батька та зневажників матері, для душогубців,
1TIM|1|10|розпусників, мужоложників, розбійників, неправдомовців, кривоприсяжників, і для всього іншого, що противне здоровій науці,
1TIM|1|11|за славною Євангелією блаженного Бога, яка мені звірена.
1TIM|1|12|Я дяку складаю Тому, Хто зміцнив мене, Христу Ісусу, Господу нашому, що мене за вірного визнав і поставив на службу,
1TIM|1|13|мене, що давніше був богозневажник, і гнобитель, і напасник, але був помилуваний, бо я те чинив нетямучий у невірстві.
1TIM|1|14|І багато збільшилась у мені благодать Господа нашого з вірою та з любов'ю в Христі Ісусі.
1TIM|1|15|Вірне це слово, і гідне всякого прийняття, що Христос Ісус прийшов у світ спасти грішних, із яких перший то я.
1TIM|1|16|Але я тому був помилуваний, щоб Ісус Христос на першім мені показав усе довготерпіння, для прикладу тим, що мають увірувати в Нього на вічне життя.
1TIM|1|17|А Цареві віків, нетлінному, невидимому, єдиному Богові честь і слава на вічні віки. Амінь.
1TIM|1|18|Цього наказа я передаю тобі, сину мій Тимофіє, за тими пророцтвами, що про тебе давніше були, щоб ними провадив ти добру війну,
1TIM|1|19|маючи віру та добре сумління, якого дехто відкинулися та й розбилися в вірі.
1TIM|1|20|Серед них Гіменей та Олександер, яких я передав сатані, щоб навчились вони не зневажати Бога.
1TIM|2|1|Отже, перш над усе я благаю чинити молитви, благання, прохання, подяки за всіх людей,
1TIM|2|2|за царів та за всіх, хто при владі, щоб могли ми провадити тихе й мирне життя в усякій побожності та чистості.
1TIM|2|3|Бо це добре й приємне Спасителеві нашому Богові,
1TIM|2|4|що хоче, щоб усі люди спаслися, і прийшли до пізнання правди.
1TIM|2|5|Один бо є Бог, і один Посередник між Богом та людьми, людина Христос Ісус,
1TIM|2|6|що дав Самого Себе на викуп за всіх. Таке було свідоцтво часу свого,
1TIM|2|7|на що я поставлений був за проповідника та за апостола, правду кажу, не обманюю, за вчителя поганів у вірі та в правді.
1TIM|2|8|Отож, хочу я, щоб мужі чинили молитви на кожному місці, підіймаючи чисті руки без гніву та сумніву.
1TIM|2|9|Так само й жінки, у скромнім убранні, з соромливістю та невинністю, нехай прикрашають себе не плетінням волосся, не коштовними шатами,
1TIM|2|10|але добрими вчинками, як то личить жінкам, що присвячуються на побожність.
1TIM|2|11|Нехай жінка навчається мовчки в повній покорі.
1TIM|2|12|А жінці навчати я не дозволяю, ані панувати над мужем, але бути в мовчанні.
1TIM|2|13|Адам бо був створений перше, а Єва потому.
1TIM|2|14|І Адам не був зведений, але, зведена бувши, жінка попала в переступ.
1TIM|2|15|Та спасеться вона дітородженням, якщо пробуватиме в вірі й любові, та в посвяті з розвагою.
1TIM|3|1|Вірне це слово: коли хто єпископства хоче, доброго діла він прагне.
1TIM|3|2|А єпископ має бути бездоганний, муж однієї дружини, тверезий, невинний, чесний, гостинний до приходнів, здібний навчати,
1TIM|3|3|не п'яниця, не заводіяка, але тихий, несварливий, не сріблолюбець,
1TIM|3|4|щоб добре рядив власним домом, що має дітей у слухняності з повною чесністю,
1TIM|3|5|бо хто власним домом рядити не вміє, як він зможе пильнувати про Божу Церкву?
1TIM|3|6|не новонавернений, щоб він не запишався, і не впав у ворожий осуд.
1TIM|3|7|Треба, щоб мав він і добре засвідчення від чужинців, щоб не впасти в догану та в сітку диявольську.
1TIM|3|8|Так само диякони мають бути поважні, не двомовці, не багато віддані вину, не соромнозахланні,
1TIM|3|9|такі, що мають таємницю віри при чистім сумлінні.
1TIM|3|10|Отже, і вони нехай перш випробовуються, а потому хай служать, якщо будуть бездоганні.
1TIM|3|11|Так само жінки нехай будуть поважні, не обмовливі, тверезі та вірні в усьому.
1TIM|3|12|Диякони мусять бути мужі однієї дружини, що добре рядять дітьми й своїми домами.
1TIM|3|13|Бо хто добре виконує службу, той добрий ступінь набуває собі та велику відвагу в вірі через Христа Ісуса.
1TIM|3|14|Це пишу я тобі, і сподіваюсь до тебе прийти незабаром.
1TIM|3|15|А коли я спізнюся, то щоб знав ти, як треба поводитися в Божому домі, що ним є Церква Бога Живого, стовп і підвалина правди.
1TIM|3|16|Безсумнівно, велика це таємниця благочестя: Хто в тілі з'явився, Той оправданий Духом, Анголам показався, проповіданий був між народами, увірувано в Нього в світі, Він у славі вознісся!
1TIM|4|1|А Дух ясно говорить, що від віри відступляться дехто в останні часи, ті, хто слухає духів підступних і наук демонів,
1TIM|4|2|хто в лицемірстві говорить неправду, і спалив сумління своє,
1TIM|4|3|хто одружуватися забороняє, наказує стримуватися від їжі, яку Бог створив на поживу з подякою віруючим та тим, хто правду пізнав.
1TIM|4|4|Кожне бо Боже твориво добре, і ніщо не негідне, що приймаємо з подякою,
1TIM|4|5|воно бо освячується Божим Словом і молитвою.
1TIM|4|6|Як будеш оце подавати братам, то будеш ти добрий служитель Христа Ісуса, годований словами віри та доброї науки, що за нею слідом ти пішов.
1TIM|4|7|Цурайся нечистих та бабських байок, а вправляйся в благочесті.
1TIM|4|8|Бо вправа тілесна мало корисна, а благочестя корисне на все, бо має обітницю життя теперішнього та майбутнього.
1TIM|4|9|Вірне це слово, і гідне всякого прийняття!
1TIM|4|10|Бо на це ми й працюємо і зносимо ганьбу, що надію кладемо на Бога Живого, Який усім людям Спаситель, найбільше ж для вірних.
1TIM|4|11|Наказуй оце та навчай!
1TIM|4|12|Нехай молодим твоїм віком ніхто не гордує, але будь зразком для вірних у слові, у житті, у любові, у дусі, у вірі, у чистості!
1TIM|4|13|Поки прийду я, пильнуй читання, нагадування та науки!
1TIM|4|14|Не занедбуй благодатного дара в собі, що був даний тобі за пророцтвом із покладенням рук пресвітерів.
1TIM|4|15|Про це піклуйся, у цім пробувай, щоб успіх твій був явний для всіх!
1TIM|4|16|Уважай на самого себе та на науку, тримайся цього. Бо чинячи так, ти спасеш і самого себе, і тих, хто тебе слухає!
1TIM|5|1|Старшого не докоряй, але вмовляй, немов батька, а молодших як братів,
1TIM|5|2|старших жінок немов матірок, молодших як сестер, зо всякою чистістю.
1TIM|5|3|Шануй вдів, удів правдивих.
1TIM|5|4|А як має вдовиця яка дітей чи внучат, нехай учаться перше побожно шанувати родину свою, і віддячуватися батькам, бо це Богові вгодно.
1TIM|5|5|А вдовиця правдива й самотна надію складає на Бога, та перебуває день і ніч у молитвах і благаннях.
1TIM|5|6|А котра у розкошах живе, та живою померла.
1TIM|5|7|І це наказуй, щоб були непорочні.
1TIM|5|8|Коли ж хто про своїх, особливо ж про домашніх не дбає, той вирікся віри, і він гірший від невірного.
1TIM|5|9|А вдову вносити до списку не менше, як шістдесятлітню, що була за дружину одному чоловікові,
1TIM|5|10|засвідчену в добрих ділах, якщо дітей виховала, якщо подорожніх приймала, якщо ноги святим умивала, якщо помагала обездоленим, якщо всякий добрий учинок виконувала.
1TIM|5|11|Але вдів молодих не приймай, бо вони, розпалившися, хочуть, наперекір Христові, заміж виходити,
1TIM|5|12|через що мають осуд, бо від першої віри відкинулись.
1TIM|5|13|А разом із тим неробітні вони, бо вчаться ходити по домах, і не тільки неробітні, але й лепетливі, і занадто цікаві, і говорять, чого не годиться.
1TIM|5|14|Отож бо, я хочу, щоб молодші заміж виходили, родили дітей, домом рядили, не давали противникові ані жадного поводу для лихомовства.
1TIM|5|15|Бо вже дехто пішли слідом за сатаною.
1TIM|5|16|А коли має вдів який вірний, нехай їх утримує, а Церква нехай не обтяжується, щоб могла вона втримувати вдів правдивих.
1TIM|5|17|А пресвітери, які добре пильнують діла, нехай будуть наділені подвійною честю, а надто ті, хто працює у слові й науці.
1TIM|5|18|Бо каже Писання: Не в'яжи рота волові, що молотить, та: Вартий працівник своєї нагороди.
1TIM|5|19|Не приймай скарги проти пресвітера, хібащо при двох чи трьох свідках.
1TIM|5|20|А тих, хто грішить, картай перед усіма, щоб і інші страх мали.
1TIM|5|21|Заклинаю тебе перед Богом й Ісусом Христом та вибраними Анголами, щоб ти заховав це без лицемірства, нічого не роблячи з упередженням.
1TIM|5|22|Не рукополагай скоро нікого, і не приставай до чужих гріхів. Бережи себе чистим!
1TIM|5|23|Води більше не пий, але трохи вина заживай ради шлунка твого та частих недугів твоїх.
1TIM|5|24|У інших людей гріхи явні і йдуть перед ними на осуд, а за іншими йдуть слідкома.
1TIM|5|25|Явні так само й добрі діла, а ті, хто інакший, сховатись не можуть.
1TIM|6|1|Усі раби, які під ярмом, нехай уважають панів своїх гідними всякої чести, щоб не зневажалися Боже Ім'я та наука.
1TIM|6|2|А ті, хто має панів віруючих, не повинні недбати про них через те, що браття вони, але нехай служать їм тим більше, що вони віруючі та улюблені, що вони добродійства Божі приймають. Оцього навчай та нагадуй!
1TIM|6|3|А коли хто навчає інакше, і не приступає до здорових слів Господа нашого Ісуса Христа та до науки, що вона за правдивою вірою,
1TIM|6|4|той згордів, нічого не знає, але захворів на суперечки й змагання, що від них повстають заздрість, сварки, богозневаги, лукаві здогади,
1TIM|6|5|постійні сварні між людьми зіпсутого розуму й позбавлених правди, які думають, ніби благочестя то зиск. Цурайся таких!
1TIM|6|6|Великий же зиск то благочестя із задоволенням.
1TIM|6|7|Бо ми не принесли в світ нічого, то нічого не можемо й винести.
1TIM|6|8|А як маєм поживу та одяг, то ми задоволені будьмо з того.
1TIM|6|9|А ті, хто хоче багатіти, упадають у спокуси та в сітку, та в численні нерозумні й шкідливі пожадливості, що втручають людей на загладу й загибіль.
1TIM|6|10|Бо корень усього лихого то грошолюбство, якому віддавшись, дехто відбились від віри й поклали на себе великі страждання.
1TIM|6|11|Але ти, о Божа людино, утікай від такого, а женися за правдою, благочестям, вірою, любов'ю, терпеливістю, лагідністю!
1TIM|6|12|Змагай добрим змагом віри, ухопися за вічне життя, до якого й покликаний ти, і визнав був добре визнання перед свідками багатьома.
1TIM|6|13|Наказую перед Богом, що оживлює все, і перед Христом Ісусом, Який добре визнання засвідчив за Понтія Пилата,
1TIM|6|14|щоб додержав ти заповідь чистою та бездоганною аж до з'явлення Господа нашого Ісуса Христа,
1TIM|6|15|що його свого часу покаже блаженний і єдиний міцний, Цар над царями та Пан над панами,
1TIM|6|16|Єдиний, що має безсмертя, і живе в неприступному світлі, Якого не бачив ніхто із людей, ані бачити не може. Честь Йому й вічна влада, амінь!
1TIM|6|17|Наказуй багатим за віку теперішнього, щоб не неслися високо, і щоб надії не клали на багатство непевне, а на Бога Живого, що щедро дає нам усе на спожиток,
1TIM|6|18|щоб робили добро, багатилися в добрих ділах, були щедрі та пильні,
1TIM|6|19|щоб збирали собі скарб, як добру основу в майбутньому, щоб прийняти правдиве життя.
1TIM|6|20|О Тимофію, бережи передання, стережися марного базікання та суперечок знання, неправдиво названого так.
1TIM|6|21|Дехто віддався йому, та й від віри відпав. Благодать з тобою. Амінь.
