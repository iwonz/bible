1PET|1|1|耶稣基督的使徒 彼得 写信给那些被拣选，分散在 本都 、 加拉太 、 加帕多家 、 亚细亚 、 庇推尼 寄居的人，
1PET|1|2|就是照父上帝的预知，藉着圣灵得以成圣，以致顺服耶稣基督，又蒙他血所洒的人。愿恩惠、平安 多多地赐给你们！
1PET|1|3|愿颂赞归于我们主耶稣基督的父上帝！他曾照自己的大怜悯，藉着耶稣基督从死人中复活，重生了我们，使我们有活的盼望，
1PET|1|4|好得到不朽坏、不玷污、不衰残、为你们存留在天上的基业，
1PET|1|5|就是为你们这些藉着信、蒙上帝大能保守的人，能获得他所预备、到末世要显现的救恩。
1PET|1|6|虽然你们必须在百般试炼中暂时忧愁，你们要为此喜乐 ，
1PET|1|7|使你们的信心既被考验，就比那被火试炼仍然能坏的金子更显宝贵，可以在耶稣基督显现的时候得著称赞、荣耀、尊贵。
1PET|1|8|虽然你们没有见过他，却是爱他；如今虽看不见，你们却因信他而有说不出来、满有荣光的喜乐，
1PET|1|9|因为你们 得到信心的效果，就是灵魂的得救。
1PET|1|10|论到这救恩，那预先说你们要得恩典的众先知已经详细地搜索查考过，
1PET|1|11|查考在他们心里的基督的灵预先证明基督受苦难，后来得荣耀，是指什么时候，什么样的情况。
1PET|1|12|他们得了启示，知道他们所服事的不是自己，而是你们。那藉着从天上差来的圣灵传福音给你们的人，现在将这些事传给你们；这些事连天使也都切望察看呢！
1PET|1|13|所以，要准备 好你们的心，谨慎自守，专心盼望耶稣基督显现的时候带给你们的恩惠。
1PET|1|14|作为顺服的儿女，就不要效法从前蒙昧无知的时候那放纵私欲的样子。
1PET|1|15|但那召你们的既是圣洁，你们在一切所行的事上也要圣洁；
1PET|1|16|因为经上记着：“你们要成为圣，因为我是神圣的。”
1PET|1|17|既然你们称那不偏待人、按各人行为审判人的主为父 ，就当存敬畏的心，度你们在世寄居的日子。
1PET|1|18|你们知道，你们得以从你们祖先传下来虚妄的行为中救赎出来，不是靠着会朽坏的金银等物，
1PET|1|19|而是凭着基督的宝血，如同无瑕疵、无玷污的羔羊的血。
1PET|1|20|基督是上帝在创世以前所预知，而在这末世才为你们显现的。
1PET|1|21|你们也因着他而信那使他从死人中复活、又给他荣耀的上帝，好让你们的信心和盼望都在于上帝。
1PET|1|22|既然你们因顺从真理而洁净了自己的心灵，能真诚爱弟兄，就该以清洁的心 彼此切实相爱。
1PET|1|23|你们蒙了重生，不是由于会朽坏的种子，而是由于不会朽坏的种子，是藉着上帝永活常存的道。
1PET|1|24|因为 “凡血肉之躯的尽都如草， 他的一切荣美像草上的花； 草必枯干，花必凋谢，
1PET|1|25|惟有主的道永远常存。” 这话就是传给你们的福音。
1PET|2|1|所以，你们要除去一切的恶毒，一切诡诈、假善、嫉妒，和一切毁谤的话。
1PET|2|2|要爱慕那纯净的灵奶，像初生的婴孩爱慕奶一样，好使你们藉着它成长，以致得救，
1PET|2|3|因为你们已经尝过主恩的滋味。
1PET|2|4|要亲近主，他是活石，虽然被人所丢弃，却是上帝所拣选、所珍贵的。
1PET|2|5|你们作为活石，要被建造成属灵的殿，成为圣洁的祭司，藉着耶稣基督献上蒙上帝悦纳的属灵祭物。
1PET|2|6|因为经上说： “看哪，我把一块石头放在 锡安 — 一块蒙拣选、珍贵的房角石； 信靠他的人必不蒙羞。”
1PET|2|7|所以，这石头在你们信的人是珍贵的；在那不信的人却有话说： “匠人所丢弃的石头 已作了房角的头块石头。”
1PET|2|8|又说： “作了绊脚的石头， 使人跌倒的磐石。” 他们绊跌，因为不顺从这道，这也是预定的。
1PET|2|9|不过，你们是被拣选的一族，是君尊的祭司，是神圣的国度，是属上帝的子民，要使你们宣扬那召你们出黑暗入奇妙光明者的美德。
1PET|2|10|“你们从前不是子民， 现在却成了上帝的子民； 从前未曾蒙怜悯， 现在却蒙了怜悯。”
1PET|2|11|亲爱的，你们是客旅，是寄居的，我劝你们要禁戒肉体的情欲；这情欲是与灵魂争战的。
1PET|2|12|你们在外邦人中要品行端正，好让那些人，虽然毁谤你们是作恶的，会因看见你们的好行为而在鉴察 的日子归荣耀给上帝。
1PET|2|13|你们为主的缘故要顺服人的一切制度，或是在上的君王，
1PET|2|14|或是君王所派惩恶赏善的官员。
1PET|2|15|因为上帝的旨意原是要你们以行善来堵住糊涂无知人的口。
1PET|2|16|虽然你们是自由的，却不可藉着自由遮盖恶毒，总要作上帝的仆人。
1PET|2|17|务要尊重众人；要敬爱教中的弟兄姊妹；要敬畏上帝；要尊敬君王。
1PET|2|18|你们作奴仆的，凡事要存敬畏的心顺服主人；不但顺服善良温和的，就是乖僻的也要顺服。
1PET|2|19|倘若你们为使良心对得起上帝，忍受冤屈的痛苦，这是可赞许的。
1PET|2|20|你们若因犯罪受责打而忍耐，有什么可称赞的呢？但你们若因行善受苦而忍耐，这在上帝看来是可赞许的。
1PET|2|21|你们蒙召就是为此，因为基督也为你们受过苦，给你们留下榜样，为要使你们跟随他的脚踪。
1PET|2|22|“他并没有犯罪， 口里也没有诡诈。”
1PET|2|23|他被辱骂不还口，受害也不说威吓的话，只将自己交托给公义的审判者。
1PET|2|24|他被挂在木头上，亲身担当了我们的罪，使我们既然在罪上死，就得以在义上活。因他受的鞭伤，你们得了医治。
1PET|2|25|你们从前好像迷路的羊，如今却归回你们灵魂的牧人和监督了。
1PET|3|1|同样，你们作妻子的，要顺服自己的丈夫，这样，即使有不信从道理的丈夫，也会因妻子的品行，并非言语，而感化过来，
1PET|3|2|因为看见了你们敬虔纯洁的品行。
1PET|3|3|你们不要藉外表来妆饰自己，如编头发，戴金饰，穿美丽的衣裳等，
1PET|3|4|而要有蕴藏在人内心不衰退的美，以温柔娴静的心妆饰自己；这在上帝面前是极宝贵的。
1PET|3|5|因为古时仰赖上帝的圣洁妇人正是以此为妆饰，顺服自己的丈夫。
1PET|3|6|就如 撒拉 听从 亚伯拉罕 ，称他为主。你们只要行善，不怕任何恐吓，就成为 撒拉 的女儿了。
1PET|3|7|同样，你们作丈夫的，要按情理 跟妻子共同生活，体贴女性是比较软弱的器皿；要尊重她，因为她也与你一同承受生命之恩。这样，你们的祷告就不会受阻碍。
1PET|3|8|总而言之，你们都要同心，彼此体恤，相爱如弟兄，存怜悯和谦卑的心。
1PET|3|9|不要以恶报恶，以辱骂还辱骂，倒要祝福，因为你们正是为此蒙召的，好使你们承受福气。
1PET|3|10|因为经上说： “凡要爱惜生命、 享受好日子的人， 要禁止舌头不出恶言， 嘴唇不说诡诈的话。
1PET|3|11|也要弃恶行善， 寻求和睦，一心追求。
1PET|3|12|因为主的眼看顾义人， 他的耳听他们的祈祷； 但主向行恶的人变脸。”
1PET|3|13|你们若热心行善，有谁会害你们呢？
1PET|3|14|即使你们为义受苦，也是有福的。不要怕人的威吓，也不要惊慌；
1PET|3|15|只要心里奉主基督为圣，尊他为主。有人问你们心中盼望的理由，要随时准备答覆；
1PET|3|16|不过，要以温柔、敬畏的心回答。要存无亏的良心，使你们在何事上被毁谤，就在何事上使那些凌辱你们在基督里有好品行的人自觉羞愧。
1PET|3|17|上帝的旨意若是要你们因行善受苦，这总比因行恶受苦好。
1PET|3|18|因为基督也曾一次为罪受苦 ， 就是义的代替不义的， 为要引领你们 到上帝面前。 在肉体里，他被治死； 但在灵里，他复活了。
1PET|3|19|他藉这灵也曾去向那些在监狱里的灵传道，
1PET|3|20|就是那些从前在 挪亚 预备方舟、上帝容忍等待的时候不信从的人。当时进入方舟，藉着水得救的不多，只有八个人。
1PET|3|21|这水所预表的洗礼，现在藉着耶稣基督的复活拯救你们，不是除掉肉体的污秽，而是向上帝恳求有无亏的良心。
1PET|3|22|耶稣已经到天上去，在上帝的右边，众天使、有权柄的、有权能的都服从了他。
1PET|4|1|既然基督在肉身受苦，你们也该将这样的心志作为兵器，因为在肉身受过苦的已经与罪断绝了，
1PET|4|2|使你们从今以后不再随从人的情欲，只顺从上帝的旨意，在世度余下的光阴。
1PET|4|3|因为你们从前随从外邦人的心意，生活在淫荡、情欲、醉酒、荒宴、狂饮和可憎的偶像崇拜中，时候已经够了。
1PET|4|4|在这些事上，他们见你们不与他们同奔放荡无度的路就以为怪，毁谤你们。
1PET|4|5|他们必须在那位将要审判活人死人的主面前交账。
1PET|4|6|为此，死人也曾有福音传给他们，要使他们的肉体按着人受审判，他们的灵却靠上帝活着。
1PET|4|7|万物的结局近了。所以你们要谨慎自守，要警醒祷告。
1PET|4|8|最要紧的是彼此切实相爱，因为爱能遮掩许多的罪。
1PET|4|9|你们要互相款待，不发怨言。
1PET|4|10|人人要照自己所得的恩赐彼此服事，作上帝各种恩赐的好管家。
1PET|4|11|若有人讲道，他要按着上帝的圣言讲；若有人服事，他要按着上帝所赐的力量服事，好让上帝在凡事上因耶稣基督得荣耀。愿荣耀和权能都归给他，直到永永远远。阿们！
1PET|4|12|亲爱的，有火一般的考验临到你们，不要奇怪，似乎是遭遇非常的事；
1PET|4|13|倒要欢喜，因为你们是与基督一同受苦，使你们在他荣耀显现的时候也可以欢喜快乐。
1PET|4|14|你们若为基督的名受辱骂是有福的，因为荣耀的灵，就是上帝的灵，在你们身上。
1PET|4|15|你们中间，不可有人因为杀人、偷窃、作恶、好管闲事而受苦。
1PET|4|16|若有人因是基督徒而受苦，不要引以为耻，倒要因这名而归荣耀给上帝。
1PET|4|17|因为时候到了，审判要从上帝的家开始；若是先从我们开始，那么，不信从上帝福音的人将有何等的结局呢？
1PET|4|18|“若是义人还仅仅得救， 不虔敬和犯罪的人将有何地可站呢？”
1PET|4|19|所以，照上帝旨意受苦的人要一心为善，将自己的灵魂交给那信实的造物主。
1PET|5|1|所以，我这同作长老，作基督受苦的证人和分享将来所要显现的荣耀的人，勉励在你们中间的长老们：
1PET|5|2|务要牧养在你们当中上帝的群羊，按着上帝的旨意照顾他们 ，不是出于勉强，而是出于甘心；也不是因为贪财，而是出于乐意。
1PET|5|3|不要辖制所托付你们的群羊，而是要作他们的榜样。
1PET|5|4|到了大牧人显现的时候，你们必得到那永不衰残、荣耀的冠冕。
1PET|5|5|同样，你们年轻的，要顺服年长的。你们大家都要以谦卑当衣服穿上，彼此顺服，因为 “上帝抵挡骄傲的人， 但赐恩给谦卑的人。”
1PET|5|6|所以，你们要谦卑服在上帝大能的手下，这样，到了适当的时候，他必使你们升高。
1PET|5|7|你们要将一切的忧虑卸给上帝，因为他顾念你们。
1PET|5|8|务要谨慎，要警醒。因为你们的仇敌魔鬼，如同咆哮的狮子，走来走去，寻找可吞吃的人。
1PET|5|9|你们要用坚固的信心抵挡他，因为知道你们在世上的众弟兄也正在经历这样的苦难。
1PET|5|10|那赐一切恩典的上帝曾在基督 里召了你们，得享他永远的荣耀，在你们暂受苦难之后，必要亲自成全你们，坚固你们，赐力量给你们，建立你们 。
1PET|5|11|愿权能归给他，直到永永远远。阿们！
1PET|5|12|我简单地写了这信，托我所看为忠心的弟兄 西拉 交给你们，劝勉你们，又证明这恩是上帝真实的恩典；你们务要在这恩上站立得住。
1PET|5|13|在 巴比伦 与你们同蒙拣选的教会向你们问安。我儿子 马可 也向你们问安。
1PET|5|14|你们要用爱心彼此亲吻问安。愿平安 归给你们所有在基督里的人！
