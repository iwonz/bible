RUTH|1|1|In the days when the judges ruled there was a famine in the land, and a man of Bethlehem in Judah went to sojourn in the country of Moab, he and his wife and his two sons.
RUTH|1|2|The name of the man was Elimelech and the name of his wife Naomi, and the names of his two sons were Mahlon and Chilion. They were Ephrathites from Bethlehem in Judah. They went into the country of Moab and remained there.
RUTH|1|3|But Elimelech, the husband of Naomi, died, and she was left with her two sons.
RUTH|1|4|These took Moabite wives; the name of the one was Orpah and the name of the other Ruth. They lived there about ten years,
RUTH|1|5|and both Mahlon and Chilion died, so that the woman was left without her two sons and her husband.
RUTH|1|6|Then she arose with her daughters-in-law to return from the country of Moab, for she had heard in the fields of Moab that the LORD had visited his people and given them food.
RUTH|1|7|So she set out from the place where she was with her two daughters-in-law, and they went on the way to return to the land of Judah.
RUTH|1|8|But Naomi said to her two daughters-in-law, "Go, return each of you to her mother's house. May the LORD deal kindly with you, as you have dealt with the dead and with me.
RUTH|1|9|The LORD grant that you may find rest, each of you in the house of her husband!" Then she kissed them, and they lifted up their voices and wept.
RUTH|1|10|And they said to her, "No, we will return with you to your people."
RUTH|1|11|But Naomi said, "Turn back, my daughters; why will you go with me? Have I yet sons in my womb that they may become your husbands?
RUTH|1|12|Turn back, my daughters; go your way, for I am too old to have a husband. If I should say I have hope, even if I should have a husband this night and should bear sons,
RUTH|1|13|would you therefore wait till they were grown? Would you therefore refrain from marrying? No, my daughters, for it is exceedingly bitter to me for your sake that the hand of the LORD has gone out against me."
RUTH|1|14|Then they lifted up their voices and wept again. And Orpah kissed her mother-in-law, but Ruth clung to her.
RUTH|1|15|And she said, "See, your sister-in-law has gone back to her people and to her gods; return after your sister-in-law."
RUTH|1|16|But Ruth said, "Do not urge me to leave you or to return from following you. For where you go I will go, and where you lodge I will lodge. Your people shall be my people, and your God my God.
RUTH|1|17|Where you die I will die, and there will I be buried. May the LORD do so to me and more also if anything but death parts me from you."
RUTH|1|18|And when Naomi saw that she was determined to go with her, she said no more.
RUTH|1|19|So the two of them went on until they came to Bethlehem. And when they came to Bethlehem, the whole town was stirred because of them. And the women said, "Is this Naomi?"
RUTH|1|20|She said to them, "Do not call me Naomi; call me Mara, for the Almighty has dealt very bitterly with me.
RUTH|1|21|I went away full, and the LORD has brought me back empty. Why call me Naomi, when the LORD has testified against me and the Almighty has brought calamity upon me?"
RUTH|1|22|So Naomi returned, and Ruth the Moabite her daughter-in-law with her, who returned from the country of Moab. And they came to Bethlehem at the beginning of barley harvest.
RUTH|2|1|Now Naomi had a relative of her husband's, a worthy man of the clan of Elimelech, whose name was Boaz.
RUTH|2|2|And Ruth the Moabite said to Naomi, "Let me go to the field and glean among the ears of grain after him in whose sight I shall find favor." And she said to her, "Go, my daughter."
RUTH|2|3|So she set out and went and gleaned in the field after the reapers, and she happened to come to the part of the field belonging to Boaz, who was of the clan of Elimelech.
RUTH|2|4|And behold, Boaz came from Bethlehem. And he said to the reapers, "The LORD be with you!" And they answered, "The LORD bless you."
RUTH|2|5|Then Boaz said to his young man who was in charge of the reapers, "Whose young woman is this?"
RUTH|2|6|And the servant who was in charge of the reapers answered, "She is the young Moabite woman, who came back with Naomi from the country of Moab.
RUTH|2|7|She said, 'Please let me glean and gather among the sheaves after the reapers.' So she came, and she has continued from early morning until now, except for a short rest."
RUTH|2|8|Then Boaz said to Ruth, "Now, listen, my daughter, do not go to glean in another field or leave this one, but keep close to my young women.
RUTH|2|9|Let your eyes be on the field that they are reaping, and go after them. Have I not charged the young men not to touch you? And when you are thirsty, go to the vessels and drink what the young men have drawn."
RUTH|2|10|Then she fell on her face, bowing to the ground, and said to him, "Why have I found favor in your eyes, that you should take notice of me, since I am a foreigner?"
RUTH|2|11|But Boaz answered her, "All that you have done for your mother-in-law since the death of your husband has been fully told to me, and how you left your father and mother and your native land and came to a people that you did not know before.
RUTH|2|12|The LORD repay you for what you have done, and a full reward be given you by the LORD, the God of Israel, under whose wings you have come to take refuge!"
RUTH|2|13|Then she said, "I have found favor in your eyes, my lord, for you have comforted me and spoken kindly to your servant, though I am not one of your servants."
RUTH|2|14|And at mealtime Boaz said to her, "Come here and eat some bread and dip your morsel in the wine." So she sat beside the reapers, and he passed to her roasted grain. And she ate until she was satisfied, and she had some left over.
RUTH|2|15|When she rose to glean, Boaz instructed his young men, saying, "Let her glean even among the sheaves, and do not reproach her.
RUTH|2|16|And also pull out some from the bundles for her and leave it for her to glean, and do not rebuke her."
RUTH|2|17|So she gleaned in the field until evening. Then she beat out what she had gleaned, and it was about an ephah of barley.
RUTH|2|18|And she took it up and went into the city. Her mother-in-law saw what she had gleaned. She also brought out and gave her what food she had left over after being satisfied.
RUTH|2|19|And her mother-in-law said to her, "Where did you glean today? And where have you worked? Blessed be the man who took notice of you." So she told her mother-in-law with whom she had worked and said, "The man's name with whom I worked today is Boaz."
RUTH|2|20|And Naomi said to her daughter-in-law, "May he be blessed by the LORD, whose kindness has not forsaken the living or the dead!" Naomi also said to her, "The man is a close relative of ours, one of our redeemers."
RUTH|2|21|And Ruth the Moabite said, "Besides, he said to me, 'You shall keep close by my young men until they have finished all my harvest.'"
RUTH|2|22|And Naomi said to Ruth, her daughter-in-law, "It is good, my daughter, that you go out with his young women, lest in another field you be assaulted."
RUTH|2|23|So she kept close to the young women of Boaz, gleaning until the end of the barley and wheat harvests. And she lived with her mother-in-law.
RUTH|3|1|Then Naomi her mother-in-law said to her, "My daughter, should I not seek rest for you, that it may be well with you?
RUTH|3|2|Is not Boaz our relative, with whose young women you were? See, he is winnowing barley tonight at the threshing floor.
RUTH|3|3|Wash therefore and anoint yourself, and put on your cloak and go down to the threshing floor, but do not make yourself known to the man until he has finished eating and drinking.
RUTH|3|4|But when he lies down, observe the place where he lies. Then go and uncover his feet and lie down, and he will tell you what to do."
RUTH|3|5|And she replied, "All that you say I will do."
RUTH|3|6|So she went down to the threshing floor and did just as her mother-in-law had commanded her.
RUTH|3|7|And when Boaz had eaten and drunk, and his heart was merry, he went to lie down at the end of the heap of grain. Then she came softly and uncovered his feet and lay down.
RUTH|3|8|At midnight the man was startled and turned over, and behold, a woman lay at his feet!
RUTH|3|9|He said, "Who are you?" And she answered, "I am Ruth, your servant. Spread your wings over your servant, for you are a redeemer."
RUTH|3|10|And he said, "May you be blessed by the LORD, my daughter. You have made this last kindness greater than the first in that you have not gone after young men, whether poor or rich.
RUTH|3|11|And now, my daughter, do not fear. I will do for you all that you ask, for all my fellow townsmen know that you are a worthy woman.
RUTH|3|12|And now it is true that I am a redeemer. Yet there is a redeemer nearer than I.
RUTH|3|13|Remain tonight, and in the morning, if he will redeem you, good; let him do it. But if he is not willing to redeem you, then, as the LORD lives, I will redeem you. Lie down until the morning."
RUTH|3|14|So she lay at his feet until the morning, but arose before one could recognize another. And he said, "Let it not be known that the woman came to the threshing floor."
RUTH|3|15|And he said, "Bring the garment you are wearing and hold it out." So she held it, and he measured out six measures of barley and put it on her. Then she went into the city.
RUTH|3|16|And when she came to her mother-in-law, she said, "How did you fare, my daughter?" Then she told her all that the man had done for her,
RUTH|3|17|saying, "These six measures of barley he gave to me, for he said to me, 'You must not go back empty-handed to your mother-in-law.'"
RUTH|3|18|She replied, "Wait, my daughter, until you learn how the matter turns out, for the man will not rest but will settle the matter today."
RUTH|4|1|Now Boaz had gone up to the gate and sat down there. And behold, the redeemer, of whom Boaz had spoken, came by. So Boaz said, "Turn aside, friend; sit down here." And he turned aside and sat down.
RUTH|4|2|And he took ten men of the elders of the city and said, "Sit down here." So they sat down.
RUTH|4|3|Then he said to the redeemer, "Naomi, who has come back from the country of Moab, is selling the parcel of land that belonged to our relative Elimelech.
RUTH|4|4|So I thought I would tell you of it and say, 'Buy it in the presence of those sitting here and in the presence of the elders of my people.' If you will redeem it, redeem it. But if you will not, tell me, that I may know, for there is no one besides you to redeem it, and I come after you." And he said, "I will redeem it."
RUTH|4|5|Then Boaz said, "The day you buy the field from the hand of Naomi, you also acquire Ruth the Moabite, the widow of the dead, in order to perpetuate the name of the dead in his inheritance."
RUTH|4|6|Then the redeemer said, "I cannot redeem it for myself, lest I impair my own inheritance. Take my right of redemption yourself, for I cannot redeem it."
RUTH|4|7|Now this was the custom in former times in Israel concerning redeeming and exchanging: to confirm a transaction, the one drew off his sandal and gave it to the other, and this was the manner of attesting in Israel.
RUTH|4|8|So when the redeemer said to Boaz, "Buy it for yourself," he drew off his sandal.
RUTH|4|9|Then Boaz said to the elders and all the people, "You are witnesses this day that I have bought from the hand of Naomi all that belonged to Elimelech and all that belonged to Chilion and to Mahlon.
RUTH|4|10|Also Ruth the Moabite, the widow of Mahlon, I have bought to be my wife, to perpetuate the name of the dead in his inheritance, that the name of the dead may not be cut off from among his brothers and from the gate of his native place. You are witnesses this day."
RUTH|4|11|Then all the people who were at the gate and the elders said, "We are witnesses. May the LORD make the woman, who is coming into your house, like Rachel and Leah, who together built up the house of Israel. May you act worthily in Ephrathah and be renowned in Bethlehem,
RUTH|4|12|and may your house be like the house of Perez, whom Tamar bore to Judah, because of the offspring that the LORD will give you by this young woman."
RUTH|4|13|So Boaz took Ruth, and she became his wife. And he went in to her, and the LORD gave her conception, and she bore a son.
RUTH|4|14|Then the women said to Naomi, "Blessed be the LORD, who has not left you this day without a redeemer, and may his name be renowned in Israel!
RUTH|4|15|He shall be to you a restorer of life and a nourisher of your old age, for your daughter-in-law who loves you, who is more to you than seven sons, has given birth to him."
RUTH|4|16|Then Naomi took the child and laid him on her lap and became his nurse.
RUTH|4|17|And the women of the neighborhood gave him a name, saying, "A son has been born to Naomi." They named him Obed. He was the father of Jesse, the father of David.
RUTH|4|18|Now these are the generations of Perez: Perez fathered Hezron,
RUTH|4|19|Hezron fathered Ram, Ram fathered Amminadab,
RUTH|4|20|Amminadab fathered Nahshon, Nahshon fathered Salmon,
RUTH|4|21|Salmon fathered Boaz, Boaz fathered Obed,
RUTH|4|22|Obed fathered Jesse, and Jesse fathered David.
