LEV|1|1|耶和华从会幕中呼叫 摩西 ，吩咐他说：
LEV|1|2|“你要吩咐 以色列 人，对他们说：你们中间若有人要献供物给耶和华，可以从牛群羊群中献牲畜为供物。
LEV|1|3|“他的供物若以牛为燔祭，要献一头没有残疾的公牛，献在会幕的门口，他就可以在耶和华面前蒙悦纳。
LEV|1|4|他要按手在燔祭牲的头上，为自己赎罪，就蒙悦纳。
LEV|1|5|他要在耶和华面前宰公牛犊； 亚伦 子孙作祭司的要献上血，把血洒在会幕门口坛的周围。
LEV|1|6|他要剥去燔祭牲的皮，把燔祭牲切成块。
LEV|1|7|亚伦 祭司的子孙要在坛上生火，把柴摆在火上。
LEV|1|8|亚伦 子孙作祭司的要把肉块连头和脂肪，摆在坛上烧着火的柴上。
LEV|1|9|燔祭牲的内脏与小腿要用水洗净，祭司要把整只全烧在坛上，当作燔祭，是献给耶和华为馨香的火祭。
LEV|1|10|“人的供物若以绵羊或山羊为燔祭，要献一只没有残疾的公羊。
LEV|1|11|他要在坛的北边，在耶和华面前宰羊； 亚伦 子孙作祭司的要把血洒在坛的周围。
LEV|1|12|他要把燔祭牲切成块，祭司就要把肉块连头和脂肪，摆在坛上烧着火的柴上。
LEV|1|13|内脏与小腿要用水洗净，祭司要把整只献上，全烧在坛上。这是燔祭，是献给耶和华为馨香的火祭。
LEV|1|14|“人献给耶和华的供物若以鸟为燔祭，就要献斑鸠或雏鸽为他的供物。
LEV|1|15|祭司要把鸟拿到坛前，扭断它的头，把鸟烧在坛上，鸟的血要流在坛的旁边；
LEV|1|16|又要把鸟的嗉囊和里面的脏物 除掉，丢在坛东边倒灰的地方。
LEV|1|17|他要拿着鸟的两个翅膀，把鸟撕开，却不可撕断；祭司要把它摆在坛上烧着火的柴上焚烧。这是燔祭，是献给耶和华为馨香的火祭。”
LEV|2|1|“若有人献素祭为供物给耶和华，就要献细面为供物，把油浇在上面，加上乳香，
LEV|2|2|带到 亚伦 子孙作祭司的那里。祭司要从细面中取出满满的一把，又取些油和所有的乳香，把这些作为纪念的烧在坛上，是献给耶和华为馨香的火祭。
LEV|2|3|素祭所剩的要归给 亚伦 和他的子孙；在献给耶和华的火祭中，这是至圣的。
LEV|2|4|“若献炉中烤的素祭为供物，要用调了油的无酵细面饼，或抹了油的无酵薄饼。
LEV|2|5|若以铁盘上的素祭为供物，就要用调了油的无酵细面，
LEV|2|6|分成小块，浇上油；这是素祭。
LEV|2|7|若以煎锅煎的素祭为供物，就要用油与细面做成。
LEV|2|8|要把这样做成的素祭带到耶和华面前，拿给祭司，祭司要带到坛前。
LEV|2|9|祭司要从素祭中取出作为纪念的烧在坛上，是献给耶和华为馨香的火祭。
LEV|2|10|素祭所剩的要归给 亚伦 和他的子孙；在献给耶和华的火祭中，这是至圣的。
LEV|2|11|“凡献给耶和华的素祭都不可以有酵，因为你们不可把任何的酵或蜜烧了，当作火祭献给耶和华。
LEV|2|12|你们可以把这些献给耶和华当作初熟的供物，但是不可献在坛上作为馨香的祭。
LEV|2|13|凡献为素祭的供物都要用盐调和；在素祭中，不可缺少你与上帝立约的盐。一切的供物都要加盐献上。
LEV|2|14|“你若献初熟之物给耶和华为素祭，就要献在火中烘过的新麦穗，就是磨碎的新谷物，当作初熟之物的素祭。
LEV|2|15|你要加上油和乳香；这是素祭。
LEV|2|16|祭司要把供物中作为纪念的，就是一些磨碎的新谷物和一些油，以及所有的乳香，都焚烧，是献给耶和华的火祭。”
LEV|3|1|“人献平安祭为供物，若是从牛群中献，无论是公的母的，要用没有残疾的，献在耶和华面前。
LEV|3|2|他要按手在供物的头上，在会幕的门口宰了它。 亚伦 子孙作祭司的，要把血洒在坛的周围。
LEV|3|3|从平安祭中，他要把火祭献给耶和华，就是包着内脏的脂肪和内脏上所有的脂肪，
LEV|3|4|两个肾和肾上的脂肪，即靠近肾两旁的脂肪，以及肝上的网油，连同肾一起取下。
LEV|3|5|亚伦 的子孙要把这些摆在烧着火的柴上，烧在坛的燔祭上，是献给耶和华为馨香的火祭。
LEV|3|6|“人向耶和华献平安祭为供物，若是从羊群中献，无论是公的母的，要用没有残疾的。
LEV|3|7|若他献一只绵羊为供物，就要把它献在耶和华面前。
LEV|3|8|要按手在供物的头上，在会幕前宰了它。 亚伦 的子孙要把血洒在坛的周围。
LEV|3|9|从平安祭中，他要取脂肪当作火祭献给耶和华，就是靠近脊骨处取下的整条肥尾巴，包着内脏的脂肪和内脏上所有的脂肪，
LEV|3|10|两个肾和肾上的脂肪，即靠近肾两旁的脂肪，以及肝上的网油，连同肾一起取下。
LEV|3|11|祭司要把这些烧在坛上，是献给耶和华为食物的火祭。
LEV|3|12|“人的供物若是山羊，就要把它献在耶和华面前。
LEV|3|13|要按手在它的头上，在会幕前宰了它。 亚伦 的子孙要把血洒在坛的周围，
LEV|3|14|又要从供物中把火祭献给耶和华，就是包着内脏的脂肪和内脏上所有的脂肪，
LEV|3|15|两个肾和肾上的脂肪，即靠近肾两旁的脂肪，以及肝上的网油，连同肾一起取下。
LEV|3|16|祭司要把这些烧在坛上，作为馨香火祭的食物；所有的脂肪都是耶和华的。
LEV|3|17|在你们一切的住处，脂肪和血都不可吃，这要成为你们世世代代永远的定例。”
LEV|4|1|耶和华吩咐 摩西 说：
LEV|4|2|“你要吩咐 以色列 人说：若有人无意中犯罪，在任何事上犯了一条耶和华所吩咐的禁令，
LEV|4|3|或是受膏的祭司犯了罪，使百姓陷在罪里，他就当为自己所犯的罪，把没有残疾的公牛犊献给耶和华为赎罪祭。
LEV|4|4|他要把公牛牵到会幕的门口，在耶和华面前按手在牛的头上，把牛宰于耶和华面前。
LEV|4|5|受膏的祭司要取些公牛的血，带到会幕那里。
LEV|4|6|祭司要把手指蘸在血中，在耶和华面前对着圣所的幔子弹血七次，
LEV|4|7|又要把一些血抹在会幕内，耶和华面前香坛的四个翘角上，再把公牛其余的血全倒在会幕门口燔祭坛的底座上；
LEV|4|8|又要取出这头赎罪祭公牛所有的脂肪，就是包着内脏的脂肪和内脏上所有的脂肪，
LEV|4|9|两个肾和肾上的脂肪，即靠近肾两旁的脂肪，以及肝上的网油，连同肾一起取下，
LEV|4|10|正如从平安祭的牛身上所取的，祭司要把这些烧在燔祭坛上。
LEV|4|11|但公牛的皮和所有的肉，以及头、腿、内脏、粪，
LEV|4|12|就是全公牛，要搬到营外清洁的地方倒灰之处，放在柴上用火焚烧。
LEV|4|13|“ 以色列 全会众若犯了错，在任何事上犯了一条耶和华所吩咐的禁令，而有了罪，会众看不出这隐藏的事；
LEV|4|14|他们一知道犯了罪，就要献一头公牛犊为赎罪祭，牵它到会幕前。
LEV|4|15|会众的长老要在耶和华面前按手在公牛的头上，把牛宰于耶和华面前。
LEV|4|16|受膏的祭司要取些公牛的血，带到会幕那里。
LEV|4|17|祭司要用手指蘸一些血，在耶和华面前对着幔子弹七次，
LEV|4|18|又要把一些血抹在会幕内，耶和华面前坛的四个翘角上，再把其余的血全倒在会幕门口燔祭坛的底座上。
LEV|4|19|他要取出公牛所有的脂肪，烧在坛上。
LEV|4|20|他要处理这牛，正如处理那头赎罪祭的公牛一样，他要如此去做。祭司要为他们赎罪，他们就蒙赦免。
LEV|4|21|他要把牛搬到营外烧了，像烧前一头公牛一样；这是会众的赎罪祭。
LEV|4|22|“官长若犯罪，在任何事上无意中犯了一条耶和华－他的上帝所吩咐的禁令，而有了罪，
LEV|4|23|他一知道自己犯了罪，就要牵一只没有残疾的公山羊为供物。
LEV|4|24|他要按手在羊的头上，在耶和华面前宰燔祭牲的地方把它宰了；这是赎罪祭。
LEV|4|25|祭司要用手指蘸一些赎罪祭牲的血，抹在燔祭坛的四个翘角上，再把其余的血倒在燔祭坛的底座上。
LEV|4|26|祭牲所有的脂肪都要烧在坛上，正如平安祭的脂肪一样。祭司要为他的罪赎了他，他就蒙赦免。
LEV|4|27|“这地的百姓若有人无意中犯罪，在任何事上犯了一条耶和华所吩咐的禁令，而有了罪，
LEV|4|28|他一知道自己犯了罪，就要为所犯的罪牵一只没有残疾的母山羊为供物。
LEV|4|29|他要按手在赎罪祭牲的头上，在燔祭牲的地方把它宰了。
LEV|4|30|祭司要用手指蘸一些祭牲的血，抹在燔祭坛的四个翘角上，再把其余的血全倒在坛的底座上；
LEV|4|31|又要把祭牲所有的脂肪都取下，正如取平安祭牲的脂肪一样。祭司要把脂肪烧在坛上，在耶和华面前作为馨香的祭。祭司要为他赎罪，他就蒙赦免。
LEV|4|32|“人若牵一只绵羊为赎罪祭作供物，就要牵一只没有残疾的母羊。
LEV|4|33|他要按手在赎罪祭牲的头上，在宰燔祭牲的地方宰了它，作为赎罪祭。
LEV|4|34|祭司要用手指蘸一些赎罪祭牲的血，抹在燔祭坛的四个翘角上，再把其余的血全倒在坛的底座上；
LEV|4|35|又要把祭牲所有的脂肪都取下，正如取平安祭的羊的脂肪一样。祭司要按献给耶和华火祭的条例，把脂肪烧在坛上。祭司要为他所犯的罪赎了他，他就蒙赦免。”
LEV|5|1|“若有人犯了罪，就是听见了誓言，他本来可以作证，却不把所看见、所知道的说出来，必须担当他的罪孽。
LEV|5|2|若有人摸了任何不洁之物，无论是野兽的不洁尸体，家畜的不洁尸体，或是群聚动物的不洁尸体，他虽不察觉，也是不洁净，就有罪了。
LEV|5|3|或是他摸了人的不洁之物，就是任何使人成为不洁的不洁之物，他虽不察觉，但一知道，就有罪了。
LEV|5|4|若有人随口发誓，或出于恶意，或出于善意，这人无论在什么事上随意发誓，虽不察觉，但一知道，就在这其中的一件事上有罪了。
LEV|5|5|当他在这其中的一件事上有罪的时候，就要承认所犯的罪，
LEV|5|6|并要为所犯的罪，把他的赎愆祭牲，就是羊群中的一只母绵羊或母山羊，献给耶和华为赎罪祭，祭司要为他的罪赎了他。
LEV|5|7|“若他的力量不够献一只绵羊，就要为所犯的罪，把两只斑鸠或是两只雏鸽献给耶和华为赎愆祭：一只作赎罪祭，一只作燔祭。
LEV|5|8|他要把这些带到祭司那里，祭司就先把赎罪祭献上，从鸟的颈项上扭断它的头，但不把鸟撕断。
LEV|5|9|祭司要把一些赎罪祭牲的血弹在祭坛的边上，其余的血要倒在坛的底座上；这是赎罪祭。
LEV|5|10|他要依照条例献第二只鸟为燔祭。祭司要为他所犯的罪赎了他，他就蒙赦免。
LEV|5|11|“他的力量若不够献两只斑鸠或两只雏鸽，就要为所犯的罪把供物，就是十分之一伊法细面，献上为赎罪祭；不可加上油，也不可加上乳香，因为这是赎罪祭。
LEV|5|12|他要把细面带到祭司那里，祭司要取出满满的一把，作为纪念，按照献火祭给耶和华的条例把它烧在坛上；这是赎罪祭。
LEV|5|13|至于他在这几件事中所犯的任何罪，祭司要为他赎了，他就蒙赦免。剩下的都归给祭司，和素祭一样。”
LEV|5|14|耶和华吩咐 摩西 说：
LEV|5|15|“若有人在耶和华的圣物上无意中犯了罪，有了过犯，就要献羊群中一只没有残疾的公绵羊给耶和华为赎愆祭，或依圣所的舍客勒所估定的银子，作为赎愆祭。
LEV|5|16|他要为在圣物上的疏忽赔偿，另外加五分之一，把这些都交给祭司。祭司要用赎愆祭的公绵羊为他赎罪，他就蒙赦免。
LEV|5|17|“若有人犯罪，在任何事上犯了一条耶和华所吩咐的禁令，他虽不察觉，仍算有罪，必须担当自己的罪孽。
LEV|5|18|他要牵羊群中一只没有残疾的公绵羊，或照你所估定的价值，给祭司作赎愆祭。祭司要为他赎他因不知道而无意中所犯的罪，他就蒙赦免。
LEV|5|19|这是赎愆祭；因他确实得罪了耶和华。”
LEV|6|1|耶和华吩咐 摩西 说：
LEV|6|2|“若有人犯罪，得罪了耶和华，就是在邻舍寄托他的东西或抵押品上行诡诈，或抢夺，或欺压邻舍，
LEV|6|3|或是捡了失物行了诡诈，起了假誓，在人所做的任何事上犯了罪；
LEV|6|4|他既犯了罪，有了过犯，就要归还他所抢夺的，或是因欺压所得的，或是别人寄托他的，或是他所捡到的失物，
LEV|6|5|或是起假誓得来的任何东西，就要全数归还，另外再加五分之一。在查出他有罪的日子，就要立刻赔还给原主。
LEV|6|6|他要献羊群中一只没有残疾的公绵羊，给耶和华为赎愆祭，或照你所估定的价值，给祭司 作赎愆祭。
LEV|6|7|祭司要在耶和华面前为他赎罪；他无论做了什么事，以致有了罪，都必蒙赦免。”
LEV|6|8|耶和华吩咐 摩西 说：
LEV|6|9|“你要吩咐 亚伦 和他的子孙说，燔祭的条例是这样：燔祭要放在坛的底盘上，从晚上到天亮，坛上的火要不断地烧着。
LEV|6|10|祭司要穿上细麻布衣服，又要把细麻布裤子穿在身上，把在坛上烧剩的燔祭灰收起来，放在坛的旁边。
LEV|6|11|然后，他要脱去这衣服，穿上别的衣服，把灰拿到营外洁净之处。
LEV|6|12|坛上的火要不断地烧着，不可熄灭。每日早晨，祭司要在坛上烧柴，把燔祭摆在坛上，并烧平安祭牲的脂肪。
LEV|6|13|坛上的火要不断地烧着，不可熄灭。”
LEV|6|14|“素祭的条例是这样： 亚伦 的子孙要在坛前把这祭献在耶和华面前。
LEV|6|15|祭司要从素祭中的细面取出一把，再取些油和素祭上所有的乳香，把这些作为纪念的烧在坛上，是献给耶和华为馨香的祭。
LEV|6|16|亚伦 和他子孙要吃素祭剩下的；要在圣处吃这无酵饼，在会幕的院子里吃。
LEV|6|17|烤饼不可加酵。这是从献给我的火祭中归给他们的一份；如赎罪祭和赎愆祭一样，这份是至圣的。
LEV|6|18|亚伦 子孙中的男丁都要吃，因为这是你们世世代代从献给耶和华的火祭中，他们永远应得的份。凡摸这些祭物的都要成为圣。”
LEV|6|19|耶和华吩咐 摩西 说：
LEV|6|20|“这是 亚伦 受膏的日子，他和他的子孙所要献给耶和华的供物：十分之一伊法细面，如他们经常献的素祭，早晨一半，晚上一半。
LEV|6|21|要在铁盘上用油调和，调匀后，就拿去烤。素祭烤熟了要分成小块，作为献给耶和华馨香的祭。
LEV|6|22|亚伦 子孙中接续他受膏为祭司的，要把这素祭献上，全烧给耶和华。这是永远的定例。
LEV|6|23|祭司一切的素祭要全部烧了，不可以吃。”
LEV|6|24|耶和华吩咐 摩西 说：
LEV|6|25|“你要吩咐 亚伦 和他的子孙说，赎罪祭的条例是这样：要在耶和华面前宰燔祭牲的地方宰赎罪祭牲；这是至圣的。
LEV|6|26|献赎罪祭的祭司要吃这祭物；要在圣处，就是在会幕的院子里吃。
LEV|6|27|凡摸这祭肉的都要成为圣；这祭牲的血若溅在衣服上，你要在圣处洗净那溅到血的衣服 。
LEV|6|28|煮这祭物的瓦器要打碎；若祭物是在铜器里煮，要把这铜器擦净，用水冲洗。
LEV|6|29|祭司中所有的男丁都可以吃；这是至圣的。
LEV|6|30|若将任何赎罪祭的血带进会幕，为要在圣所赎罪，那肉就不可吃，要用火焚烧。”
LEV|7|1|“赎愆祭的条例是这样：这祭是至圣的。
LEV|7|2|人在哪里宰燔祭牲，也要在哪里宰赎愆祭牲；其血，祭司要洒在坛的周围。
LEV|7|3|祭司要献上它所有的脂肪，把肥尾巴和包着内脏的脂肪，
LEV|7|4|两个肾和肾上的脂肪，即靠近肾两旁的脂肪，以及肝上的网油，连同肾一起取下。
LEV|7|5|祭司要把这些烧在坛上，献给耶和华为火祭，作为赎愆祭。
LEV|7|6|祭司中所有的男丁都可以吃这祭物，要在圣处吃；这是至圣的。
LEV|7|7|赎罪祭怎样，赎愆祭也是怎样，都有一样的条例，用赎愆祭赎罪的祭司要得这祭物。
LEV|7|8|献燔祭的祭司，无论为谁献，所献燔祭牲的皮要归给那祭司，那是他的。
LEV|7|9|任何素祭，无论是在炉中烤的，用煎锅或铁盘做成的，都要归给献祭的祭司。
LEV|7|10|任何素祭，无论是用油调和的，是干的，都要归 亚伦 的子孙，大家均分。”
LEV|7|11|“献给耶和华平安祭的条例是这样：
LEV|7|12|若有人为感谢献祭，就要把用油调和的无酵饼、抹了油的无酵薄饼，和用油调匀细面做成的饼，与感谢祭一同献上。
LEV|7|13|要用有酵的饼，和那为感谢而献的平安祭，与供物一同献上。
LEV|7|14|他要从每一种供物中拿一个饼，献给耶和华为举祭，是要归给那洒平安祭牲血的祭司。
LEV|7|15|为感谢而献的平安祭的肉，要在献祭当天吃，一点也不可留到早晨。
LEV|7|16|若所献的是还愿祭或甘心祭，要在献祭当天吃，剩下的，第二天也可以吃。
LEV|7|17|第三天，所剩下的祭肉要用火焚烧。
LEV|7|18|第三天若吃平安祭的肉，必不蒙悦纳，所献的也不算为祭；这祭物是不洁净的，凡吃这祭物的，必担当自己的罪孽。
LEV|7|19|“沾了不洁净之物的肉就不可吃，要用火焚烧。至于其他的肉，凡洁净的人都可以吃这肉；
LEV|7|20|但不洁净的人若吃了献给耶和华平安祭的肉，这人必从民中剪除。
LEV|7|21|若有人摸了不洁之物，无论是人体的不洁净，或是不洁的牲畜，或是不洁的可憎之物 ，再吃了献给耶和华平安祭的肉，这人必从民中剪除。”
LEV|7|22|耶和华吩咐 摩西 说：
LEV|7|23|“你要吩咐 以色列 人说：牛、绵羊、山羊的脂肪，你们都不可吃。
LEV|7|24|自然死去的或被野兽撕裂的，那脂肪可以作别的用途，你们却万不可吃。
LEV|7|25|任何人吃了献给耶和华作火祭祭牲的脂肪，这人必从民中剪除。
LEV|7|26|在你们一切的住处，无论是鸟或兽的血，你们都不可吃。
LEV|7|27|无论谁吃了血，这人必从民中剪除。”
LEV|7|28|耶和华吩咐 摩西 说：
LEV|7|29|“你要吩咐 以色列 人说：献平安祭给耶和华的，要从他的平安祭中取些供物来献给耶和华。
LEV|7|30|他要亲手把献给耶和华的火祭带来，要把脂肪和胸带来，把胸在耶和华面前摇一摇，作为摇祭。
LEV|7|31|祭司要把脂肪烧在坛上，但胸要归给 亚伦 和他的子孙。
LEV|7|32|你们要从平安祭牲中把右腿作为举祭，送给祭司。
LEV|7|33|亚伦 子孙中献平安祭牲的血和脂肪的，要得这右腿，作为他当得的份。
LEV|7|34|因为我从 以色列 人的平安祭中，把这摇祭的胸和这举祭的腿给 亚伦 祭司和他子孙，作为他们在 以色列 人中永远当得的份。”
LEV|7|35|这是从耶和华的火祭中取出，作为 亚伦 和他子孙受膏的份，就是 摩西 叫他们前来，给耶和华供祭司职分的那一天开始的。
LEV|7|36|这是在 摩西 膏他们的日子，耶和华吩咐给他们的，作为他们在 以色列 人中世世代代永远当得的份。
LEV|7|37|这就是燔祭、素祭、赎罪祭、赎愆祭、圣职礼和平安祭的条例，
LEV|7|38|都是耶和华在 西奈山 上吩咐 摩西 的，也是他在 西奈 旷野吩咐 以色列 人献供物给耶和华的日子所说的。
LEV|8|1|耶和华吩咐 摩西 说：
LEV|8|2|“你领 亚伦 和他儿子前来，并将圣衣、膏油，与赎罪祭的一头公牛、两只公绵羊、一筐无酵饼都一同带来；
LEV|8|3|又要召集全会众到会幕的门口。”
LEV|8|4|摩西 就遵照耶和华的吩咐做了，于是会众聚集在会幕的门口。
LEV|8|5|摩西 对会众说：“这是耶和华所吩咐当做的事。”
LEV|8|6|摩西 领了 亚伦 和他儿子前来，用水洗他们。
LEV|8|7|他给 亚伦 穿上内袍，束上腰带，套上外袍，加上以弗得，再束上精致的带子，把以弗得系在他身上。
LEV|8|8|他又给 亚伦 戴上胸袋，把乌陵和土明放在胸袋内。
LEV|8|9|他把礼冠戴在 亚伦 的头上，礼冠前面安上金牌，成为圣冕，是照耶和华所吩咐 摩西 的。
LEV|8|10|摩西 用膏油抹帐幕和其中所有的，使它们成为圣。
LEV|8|11|他又用膏油在祭坛上弹了七次，抹了坛和坛的一切器皿，以及洗濯盆和盆座，使它们成为圣。
LEV|8|12|他把膏油倒在 亚伦 的头上膏他，使他成为圣。
LEV|8|13|摩西 带了 亚伦 的儿子来，给他们穿上内袍，束上腰带，裹上头巾，是照耶和华所吩咐 摩西 的。
LEV|8|14|他把赎罪祭的公牛牵来， 亚伦 和他儿子按手在赎罪祭公牛的头上，
LEV|8|15|就宰了公牛。 摩西 取了血，用指头抹在祭坛周围的四个翘角上，使坛洁净，再把其余的血倒在坛的底座上，使坛成为圣，为坛赎罪。
LEV|8|16|摩西 把内脏所有的脂肪和肝上的网油，以及两个肾与肾上的脂肪取出，都烧在坛上。
LEV|8|17|至于公牛，连皮带肉和粪，他都用火烧在营外，是照耶和华所吩咐 摩西 的。
LEV|8|18|他把燔祭的公绵羊牵来， 亚伦 和他儿子按手在羊的头上，
LEV|8|19|就宰了公羊。 摩西 把血洒在祭坛的周围，
LEV|8|20|把羊切成块，把头和肉块，以及脂肪拿去烧，
LEV|8|21|他用水洗了内脏和腿之后，就把全羊烧在坛上，作为馨香的燔祭，是献给耶和华的火祭，都是照耶和华所吩咐 摩西 的。
LEV|8|22|他又牵来第二只公绵羊，就是圣职礼的羊， 亚伦 和他儿子按手在羊的头上，
LEV|8|23|就宰了羊。 摩西 把一些血抹在 亚伦 的右耳垂上，右手的大拇指上和右脚的大脚趾上。
LEV|8|24|他领了 亚伦 的儿子来，把一些血抹在他们的右耳垂上，右手的大拇指上和右脚的大脚趾上。 摩西 把其余的血洒在坛的周围。
LEV|8|25|他把脂肪，肥尾巴、内脏所有的脂肪、肝上的网油、两个肾、肾上的脂肪，和右腿取下，
LEV|8|26|再从耶和华面前那装无酵饼的篮子中取一个无酵饼、一个油饼和一个薄饼，把这些放在脂肪和右腿上。
LEV|8|27|他把这一切放在 亚伦 和他儿子的手上，在耶和华面前摇一摇，作为摇祭。
LEV|8|28|摩西 从他们的手上把这些祭物拿来，放在坛的燔祭上烧，这就是圣职礼中献给耶和华馨香的火祭。
LEV|8|29|摩西 拿羊的胸，在耶和华面前摇一摇，作为摇祭，这是圣职礼的羊归给 摩西 的一份，是照耶和华所吩咐 摩西 的。
LEV|8|30|摩西 取些膏油和坛上的血，弹在 亚伦 和他的衣服上，以及他儿子和他们的衣服上，使 亚伦 和他的衣服，他儿子和他们的衣服都成为圣。
LEV|8|31|摩西 对 亚伦 和他儿子说：“你们要在会幕的门口把肉煮了，在那里吃这肉和圣职礼中篮子里的饼，按我所吩咐的说：‘这是 亚伦 和他儿子当吃的。’
LEV|8|32|剩下的肉和饼，你们要用火焚烧。
LEV|8|33|这七天，你们不可走出会幕的门口，直等到你们圣职礼的日子满了，因为授予你们圣职需要七天 。
LEV|8|34|今天所做的，都是耶和华吩咐要做的，好为你们赎罪。
LEV|8|35|这七天，你们要昼夜留在会幕门内，遵守耶和华所吩咐的，免得你们死亡，因为所吩咐我的就是这样。”
LEV|8|36|于是， 亚伦 和他的儿子就做了耶和华藉着 摩西 所吩咐的一切事。
LEV|9|1|到了第八天， 摩西 召 亚伦 和他儿子，以及 以色列 的众长老来，
LEV|9|2|对 亚伦 说：“你当取一头公牛犊作赎罪祭，一只公绵羊作燔祭，都要没有残疾的，献在耶和华面前。
LEV|9|3|你要对 以色列 人说：‘你们当取一只公山羊作赎罪祭，再取一头牛犊和一只小绵羊，都要一岁没有残疾的，作燔祭；
LEV|9|4|又当取一头公牛，一只公绵羊作平安祭，宰杀献在耶和华面前，再加上调油的素祭。因为今天耶和华要向你们显现。’”
LEV|9|5|于是，他们把 摩西 所吩咐的带到会幕前；全会众都近前来，站在耶和华面前。
LEV|9|6|摩西 说：“这是耶和华吩咐你们当做的事，耶和华的荣光要向你们显现。”
LEV|9|7|摩西 对 亚伦 说：“你靠近祭坛前，献你的赎罪祭和燔祭，为自己与百姓赎罪，再献上百姓的供物，为他们赎罪，都是照耶和华所吩咐的。”
LEV|9|8|于是， 亚伦 靠近坛前，宰了那头为自己赎罪的牛犊。
LEV|9|9|亚伦 的儿子把血递给他，他就把指头蘸在血中，抹在坛的四个翘角上，再把其余的血倒在坛的底座上。
LEV|9|10|他把赎罪祭的脂肪和肾，以及肝上的网油，烧在坛上，是照耶和华所吩咐 摩西 的。
LEV|9|11|他用火将肉和皮烧在营外。
LEV|9|12|亚伦 把燔祭牲宰了，他儿子把血递给他，他就把血洒在坛的周围。
LEV|9|13|他们又把燔祭一块一块地，连头递给他，他就烧在坛上。
LEV|9|14|他又洗了内脏和腿，放在坛的燔祭上烧。
LEV|9|15|然后，他奉上百姓的供物。他牵来给百姓作赎罪祭的公山羊，把它宰了，献为赎罪祭，和先前的一样。
LEV|9|16|他也奉上燔祭，按照条例献上。
LEV|9|17|除了早晨的燔祭以外，他又献上素祭，用手取了满满的一把，烧在坛上。
LEV|9|18|亚伦 宰了那给百姓作平安祭的公牛和公绵羊，他儿子把血递给他，他就把血洒在坛的周围；
LEV|9|19|他们把公牛和公绵羊的脂肪、肥尾巴，包着内脏的脂肪，肾和肝上的网油，都递给他。
LEV|9|20|他们把脂肪放在祭牲的胸上，他就把脂肪烧在坛上。
LEV|9|21|亚伦 把祭牲的胸和右腿在耶和华面前摇一摇，作为摇祭，是照 摩西 所吩咐的。
LEV|9|22|亚伦 向百姓举手，为他们祝福。他献了赎罪祭、燔祭、平安祭就下来了。
LEV|9|23|摩西 和 亚伦 进了会幕。他们出来，为百姓祝福；耶和华的荣光向全体百姓显现。
LEV|9|24|有火从耶和华面前出来，焚烧了坛上的燔祭和脂肪；全体百姓一看见，就都欢呼，脸伏于地。
LEV|10|1|亚伦 的儿子 拿答 和 亚比户 各拿着自己的香炉，把火放在炉里，加上香，在耶和华面前献上凡火，是耶和华没有吩咐他们的。
LEV|10|2|有火从耶和华面前出来，把他们吞灭，他们就死在耶和华面前。
LEV|10|3|于是， 摩西 对 亚伦 说：“这就是耶和华所吩咐的，说：‘我在那亲近我的人中要显为圣；在全体百姓面前，我要得着荣耀。’” 亚伦 就默默不言。
LEV|10|4|摩西 召 亚伦 的叔父 乌薛 的儿子 米沙利 和 以利撒反 前来，对他们说：“过来，把你们的亲属从圣所前抬到营外。”
LEV|10|5|于是，二人过来把尸体连袍子一起抬到营外，是照 摩西 所吩咐的。
LEV|10|6|摩西 对 亚伦 和他儿子 以利亚撒 和 以他玛 说：“不可蓬头散发，也不可撕裂衣服，免得你们死亡，免得耶和华向全会众发怒。但你们的弟兄 以色列 全家却要为耶和华发出的火哀哭。
LEV|10|7|你们也不可出会幕的门口，免得你们死亡，因为耶和华的膏油在你们身上。”他们就遵照 摩西 的话去做了。
LEV|10|8|耶和华吩咐 亚伦 说：
LEV|10|9|“你和你儿子进会幕的时候，清酒烈酒都不可喝，免得你们死亡，这要作你们世世代代永远的定例。
LEV|10|10|你们必须分辨圣的俗的，洁净的和不洁净的，
LEV|10|11|也要将耶和华藉 摩西 吩咐 以色列 人的一切律例教导他们。”
LEV|10|12|摩西 对 亚伦 和他剩下的儿子 以利亚撒 和 以他玛 说：“献给耶和华的火祭中所剩下的素祭，你们要拿来，在祭坛旁吃这无酵饼，因为它是至圣的。
LEV|10|13|你们要在圣处吃，因为在献给耶和华的火祭中，这是你和你儿子当得的份；所吩咐我的就是这样。
LEV|10|14|这摇祭的胸和这举祭的腿，你要在洁净的地方和你的儿女一同吃，因为这些是从 以色列 人的平安祭中归给你，作为你和你儿子当得的份。
LEV|10|15|他们要把举祭的腿、摇祭的胸和火祭的脂肪一同带来，在耶和华面前摇一摇，作为摇祭。这些要归给你和你儿子，作永远当得的份，都是照耶和华所吩咐的。”
LEV|10|16|那时， 摩西 急切地寻找那只赎罪祭的公山羊，看哪，它已经烧掉了。他向 亚伦 剩下的儿子 以利亚撒 和 以他玛 发怒，说：
LEV|10|17|“你们为何没有在圣所吃这赎罪祭呢？它是至圣的，是耶和华给你们的，为了除掉会众的罪孽，在耶和华面前为他们赎罪。
LEV|10|18|看哪，这祭牲的血没有拿到圣所里去！你们应当照我所吩咐的，在圣所里吃这祭肉。”
LEV|10|19|亚伦 对 摩西 说：“看哪，他们今天在耶和华面前献上赎罪祭和燔祭，但是我却遭遇这样的灾难。我若今天吃这赎罪祭，耶和华岂能看为美呢？”
LEV|10|20|摩西 听了，就看为美。
LEV|11|1|耶和华吩咐 摩西 和 亚伦 ，对他们说：
LEV|11|2|“你们要吩咐 以色列 人说，地上一切的走兽中可吃的动物是这些：
LEV|11|3|凡蹄分两瓣，分趾蹄而又反刍食物的走兽，你们都可以吃。
LEV|11|4|但那反刍或分蹄之中不可吃的是：骆驼，反刍却不分蹄，对你们是不洁净的；
LEV|11|5|石獾，反刍却不分蹄，对你们是不洁净的；
LEV|11|6|兔子，反刍却不分蹄，对你们是不洁净的；
LEV|11|7|猪，蹄分两瓣，分趾蹄却不反刍，对你们是不洁净的。
LEV|11|8|这些兽的肉，你们不可吃；它们的尸体，你们也不可摸，对你们都是不洁净的。
LEV|11|9|“水中可吃的是这些：凡在水里，无论是海或河，有鳍有鳞的，都可以吃。
LEV|11|10|凡在海里、河里和水里滋生的动物，就是在水里所有的动物，无鳍无鳞的，对你们是可憎的。
LEV|11|11|它们对你们都是可憎的。你们不可吃它们的肉；它们的尸体，也当以为可憎。
LEV|11|12|凡在水里无鳍无鳞的，对你们是可憎的。
LEV|11|13|“飞鸟中你们当以为可憎，不可吃且可憎的是：雕、狗头雕、红头雕，
LEV|11|14|鹞鹰、小鹰的类群，
LEV|11|15|所有乌鸦的类群，
LEV|11|16|鸵鸟、夜鹰、鱼鹰、鹰的类群，
LEV|11|17|鸮鸟、鸬鹚、猫头鹰，
LEV|11|18|角鸱、鹈鹕、秃雕，
LEV|11|19|鹳、鹭鸶的类群，戴鵀与蝙蝠。
LEV|11|20|“凡有翅膀却用四足爬行的群聚动物，对你们是可憎的。
LEV|11|21|只是有翅膀却用四足爬行的群聚动物中，足上有腿在地上跳的，你们还可以吃；
LEV|11|22|其中你们可以吃的有蝗虫的类群，蚂蚱的类群，蟋蟀的类群和蚱蜢的类群。
LEV|11|23|其余有翅膀有四足的群聚动物，对你们都是可憎的。
LEV|11|24|“这些都能使你们不洁净。凡摸它们尸体的，必不洁净到晚上。
LEV|11|25|任何人搬动了它们的尸体，要把衣服洗净，必不洁净到晚上。
LEV|11|26|凡蹄分两瓣却不分趾或不反刍食物的走兽，对你们是不洁净的；谁摸了它们就不洁净。
LEV|11|27|凡用脚掌行走，四足行走的动物，对你们是不洁净的；凡摸它们尸体的，必不洁净到晚上。
LEV|11|28|谁搬动了它们的尸体，要把衣服洗净，必不洁净到晚上。这些对你们是不洁净的。
LEV|11|29|“在地上成群的群聚动物中，对你们不洁净的是这些：鼬鼠、鼫鼠、蜥蜴的类群，
LEV|11|30|壁虎、龙子、守宫、蛇医、蝘蜓。
LEV|11|31|这些群聚动物对你们都是不洁净的。在它们死后，凡摸了它们尸体的，必不洁净到晚上。
LEV|11|32|其中死了的，若掉在任何东西上，这东西就不洁净，无论是木器、衣服、皮革、麻袋，或是任何工作需用的器皿，都要泡在水中，必不洁净到晚上，然后才是洁净的。
LEV|11|33|若有一点掉在瓦器里，里面的任何东西就不洁净了； 你们要把这瓦器打破。
LEV|11|34|其中一切可吃的食物，沾到那水的就不洁净；器皿里可喝的东西，也必不洁净。
LEV|11|35|它们的尸体，只要有一点掉在任何物件上，那物件就不洁净。无论是烤炉或炉灶，都要打碎；它们不洁净，而且对你们也不洁净。
LEV|11|36|但是水泉或池子，就是聚水的地方，仍是洁净的；凡摸这些尸体的才不洁净。
LEV|11|37|若它们的尸体有一点掉在要播的种子上，种子仍是洁净的；
LEV|11|38|若水已经浇在种子上，它们的尸体有一点掉在上面，这种子对你们就是不洁净的了。
LEV|11|39|“你们可吃的走兽中若有死了的，谁摸了它的尸体，就必不洁净到晚上。
LEV|11|40|人若吃了那已死的走兽，要把衣服洗净，必不洁净到晚上。人若搬动了那已死的牲畜，要把衣服洗净，必不洁净到晚上。
LEV|11|41|“凡在地上成群的群聚动物都是可憎的，都不可吃。
LEV|11|42|凡用肚子爬行或用四脚爬行，或是用多足的，地上一切群聚的动物，你们都不可吃，因为是可憎的。
LEV|11|43|你们不可因任何群聚的动物使自己成为可憎的，也不可因它们成为不洁净，染了污秽。
LEV|11|44|我是耶和华－你们的上帝。你们要使自己分别为圣，要成为圣，因为我是神圣的。你们不可因地上爬行的群聚动物使自己不洁净。
LEV|11|45|我是把你们从 埃及 地领出来的耶和华，要作你们的上帝。你们要成为圣，因为我是神圣的。”
LEV|11|46|这是牲畜、飞鸟、水中一切游动的生物和地上一切爬行的动物的条例，
LEV|11|47|为要使你们能分辨洁净的和不洁净的，可吃的和不可吃的动物。
LEV|12|1|耶和华吩咐 摩西 说：
LEV|12|2|“你要吩咐 以色列 人说：妇人若怀孕生男孩，就不洁净七天，像在月经污秽的期间不洁净一样。
LEV|12|3|第八天，要给婴孩行割礼。
LEV|12|4|妇人产后流血的洁净，要家居三十三天。她洁净的日子未满，不可摸圣物，也不可进入圣所。
LEV|12|5|她若生女孩，就不洁净两个七天，像经期中一样。她产后流血的洁净，要家居六十六天。
LEV|12|6|“洁净的日子满了，无论生儿子或女儿，她要把一只一岁的羔羊作燔祭，一只雏鸽或一只斑鸠作赎罪祭，带到会幕的门口交给祭司。
LEV|12|7|祭司要把这祭物献在耶和华面前，为她赎罪。这样，她就从流血中得洁净了。这是为生男或生女之妇人的条例。
LEV|12|8|妇人的能力若不足，无法献一只羔羊，她就要取两只斑鸠或两只雏鸽，一只为燔祭，一只为赎罪祭。祭司要为她赎罪，她就洁净了。”
LEV|13|1|耶和华吩咐 摩西 和 亚伦 说：
LEV|13|2|“人身上的皮肤若肿胀，或发疹，或有斑点，可能成为痲疯 的灾病，就要把他带到 亚伦 祭司或 亚伦 的一个作祭司的子孙那里。
LEV|13|3|祭司要检查他身上皮肤的患处，若患处的毛已经变白，灾病的现象深入身上皮肤内，这就是痲疯的灾病。祭司检查后，要宣布他为不洁净。
LEV|13|4|若这人身上的皮肤有白斑，看起来并没有深入皮肤内，其上的毛也没有变白，祭司就要将这病人隔离七天。
LEV|13|5|第七天，祭司要检查他，看哪，若灾病在祭司眼前止住了，没有在皮肤上扩散，要将他再隔离七天。
LEV|13|6|到了第七天，祭司要再检查他。看哪，若灾病减轻，没有在皮肤上扩散，祭司就要宣布他为洁净，因为他患的不过是疹子。那人要洗自己的衣服，就洁净了。
LEV|13|7|他给祭司检查宣布为洁净后，疹子若在皮肤上大大扩散，他就要再给祭司检查。
LEV|13|8|祭司要检查，看哪，疹子若在皮肤上扩散了，祭司就要宣布他为不洁净，是痲疯病。
LEV|13|9|“人若得了痲疯的灾病，就要把他带到祭司那里。
LEV|13|10|祭司要检查，看哪，若皮肤有白色肿块，使毛变白，肿块里有嫩的新长的肉，
LEV|13|11|这就是他身上皮肤慢性的痲疯病。祭司要宣布他为不洁净，不必将他隔离，因为他已是不洁净了。
LEV|13|12|若痲疯在皮肤四处扩散，长满在患灾病之人的皮肤上，据祭司察看，从头到脚无处不有，
LEV|13|13|祭司就要检查，看哪，若这病人全身已长满了痲疯，就要宣布他为洁净；他全身都变白了，他是洁净的。
LEV|13|14|但他身上一旦出现新长的肉，就不洁净了。
LEV|13|15|祭司一见新长的肉，就要宣布他为不洁净。新长的肉是不洁净的，这就是痲疯病。
LEV|13|16|新长的肉若变白了，他就要到祭司那里。
LEV|13|17|祭司要检查，看哪，患处若变白了，祭司就要宣布那患灾病的人为洁净，他就洁净了。
LEV|13|18|“人身上的皮肤 若长了疮，却已经好了，
LEV|13|19|在长疮之处又发肿变白，或是出现白中带红的斑点，就要给祭司检查。
LEV|13|20|祭司要检查，看哪，若灾病的现象已深入皮肤内，其上的毛也变白了，祭司就要宣布他为不洁净，有痲疯的灾病生在疮中。
LEV|13|21|祭司若检查，看哪，其上没有白毛，也没有深入皮肤内，而且灾病减轻，祭司就要将他隔离七天。
LEV|13|22|若在皮肤上大大扩散，祭司就要宣布他为不洁净，这是灾病。
LEV|13|23|斑点若留在原处，没有扩散，这就是疮的疤痕，祭司就要宣布他为洁净。
LEV|13|24|“人身上的皮肤若被火烧伤，伤口新长的肉有了斑点，无论是白中带红，或是全白，
LEV|13|25|祭司就要检查，看哪，斑点上的毛若变白了，现象又深入皮肤内，这就是痲疯长在烧伤处；祭司就要宣布他为不洁净，是痲疯的灾病。
LEV|13|26|若祭司检查，看哪，斑点上没有白毛，也没有深入皮肤内，而且灾病减轻，祭司就要将他隔离七天。
LEV|13|27|第七天，祭司要检查他。斑点若在皮肤上大大扩散，祭司就要宣布他为不洁净，是患了痲疯的灾病。
LEV|13|28|斑点若留在原处，没有在皮肤上扩散，并减轻了，它只是烧伤的肿块，祭司要宣布他为洁净，这不过是烧伤后的疤痕。
LEV|13|29|“无论男女，若在头上或下巴有灾病，
LEV|13|30|祭司就要检查这灾病，看哪，若灾病的现象深入皮肤内，其上有黄色的细毛，祭司就要宣布他为不洁净，这是疥疮，是头上或下巴的痲疯病。
LEV|13|31|祭司要检查这疥疮的灾病，看哪，现象若未深入皮肤内，其上也没有黑毛，祭司就要将长疥疮的人隔离七天。
LEV|13|32|第七天，祭司要检查这灾病，看哪，若疥疮没有扩散，其上没有黄色的毛，疥疮的现象也没有深入皮肤内，
LEV|13|33|那人就要剃去须发，但不可剃长疥疮之处。祭司要将那长疥疮的人，再隔离七天。
LEV|13|34|第七天，祭司要检查疥疮，看哪，疥疮若没有在皮肤上扩散，现象也未深入在皮肤内，祭司就要宣布他为洁净；那人要洗自己的衣服，就洁净了。
LEV|13|35|但他被宣布为洁净后，疥疮若在皮肤上大大扩散，
LEV|13|36|祭司就要检查他。看哪，疥疮若在皮肤上扩散，祭司就不必找黄色的毛，这人是不洁净了。
LEV|13|37|若疥疮在祭司眼前止住了，其上长了黑毛，疥疮就已痊愈了，那人是洁净的，祭司要宣布他为洁净。
LEV|13|38|“无论男女，身上的皮肤若有斑点，是白色的斑点，
LEV|13|39|祭司就要检查，看哪，若皮肤的斑点是暗白色的，这是皮肤长了斑；那人是洁净的。
LEV|13|40|“人的头发若掉了，变成秃头，他是洁净的。
LEV|13|41|他头顶的前面若掉了头发，以致顶门光秃，他是洁净的。
LEV|13|42|头秃处或顶门秃处，若有白中带红的灾病，这就是痲疯长在他的头秃处或顶门秃处。
LEV|13|43|祭司要检查他，看哪，若头秃处或顶门秃处的灾病肿块白中带红，像身上皮肤痲疯病的现象一样，
LEV|13|44|那人就是患了痲疯病，是不洁净的。祭司要宣布他为不洁净；他的灾病是生在头上。
LEV|13|45|“患有痲疯灾病的人，他的衣服要撕裂，也要蓬头散发，遮住上唇，喊着说：‘不洁净！不洁净！’
LEV|13|46|灾病还在他身上的时候，他就是不洁净的；既然不洁净，他就要独居，住在营外。”
LEV|13|47|“衣服若发霉 了，无论是羊毛衣服、麻布衣服，
LEV|13|48|无论是经线、纬线，是麻布的、羊毛的，是皮革，或是任何皮制的物件；
LEV|13|49|若是衣服、皮革、经线、纬线，或是任何皮制的物件呈现绿色或红色，这就是发霉，必须给祭司检查。
LEV|13|50|祭司要检查这霉，把发霉的物件隔离七天。
LEV|13|51|第七天，他要检查这霉。若霉在衣服上，无论是经线、纬线，或任何用途的皮制物件上扩散，这是侵蚀性的霉，是不洁净的。
LEV|13|52|发霉的衣服，无论在经线、纬线，羊毛的、麻布的，或是任何皮制物件，都要把它烧掉；因为这是侵蚀性的霉，必须用火焚烧。
LEV|13|53|祭司检查，看哪，霉若在衣服上，无论是经线、纬线，或在任何的皮制物件上没有扩散，
LEV|13|54|祭司就要吩咐人把发霉的物件洗了，再隔离七天。
LEV|13|55|洗过之后，祭司要检查，看哪，若那霉在他眼前没有变色，霉虽没有扩散，也是不洁净的。这是侵蚀性的灾病，无论是在正面或反面，都要用火焚烧那物件。
LEV|13|56|祭司若检查，看哪，那霉在洗过之后已经褪色，他就要从衣服，皮革，或经线、纬线，把发霉的部分撕去。
LEV|13|57|若霉再出现在衣服上，无论是经线、纬线、或在任何皮制物件上，这就是旧霉复发，必须用火将那发霉的物件焚烧。
LEV|13|58|洗过的衣服，或是经线，纬线，或是任何皮制的物件，若霉已经消失了，仍要再洗，这衣服就洁净了。”
LEV|13|59|这就是衣服发霉的条例。无论是羊毛衣服，麻布衣服，或是经线、纬线，或任何皮制的物件，都按照这条例宣布为洁净或不洁净。
LEV|14|1|耶和华吩咐 摩西 说：
LEV|14|2|“这是患痲疯病的人得洁净时的条例：要带他到祭司那里，
LEV|14|3|祭司要出到营外，检查那患痲疯病的人，看哪，他的痲疯灾病已经痊愈了，
LEV|14|4|祭司就要吩咐人为那求洁净的人带两只洁净的活鸟和香柏木、朱红色纱，以及牛膝草来。
LEV|14|5|祭司要吩咐用瓦器盛清水，把第一只鸟宰在上面。
LEV|14|6|至于那只活鸟，祭司要把它和香柏木、朱红色纱，以及牛膝草，一同蘸在宰于清水上的鸟血中。
LEV|14|7|他要向那从痲疯病中得洁净的人身上弹血七次，宣布他为洁净，然后把那活鸟在野地里放走。
LEV|14|8|求洁净的人要洗衣服，剃去所有的毛发，用水洗澡，他就洁净了。然后，他可以进营，不过仍要在自己的帐棚外居住七天。
LEV|14|9|到了第七天，他要剃所有的毛发，头发、胡须、眼睛的眉毛，他全身的毛都剃了；然后，他要洗衣服，用水洗身，才洁净了。
LEV|14|10|“第八天，他要取两只没有残疾的小公羊和一只没有残疾、一岁的小母羊，以及作为素祭的十分之三伊法调了油的细面和一罗革的油。
LEV|14|11|宣布洁净的祭司要将那求洁净的人，连同这些东西，安置在耶和华面前，会幕的门口。
LEV|14|12|祭司要取一只小公羊献为赎愆祭，又取一罗革的油，把它们在耶和华面前摇一摇，作为摇祭；
LEV|14|13|再把小公羊宰于圣处，就是宰赎罪祭牲和燔祭牲的地方。赎愆祭要归给祭司，与赎罪祭一样，是至圣的。
LEV|14|14|祭司要取一些赎愆祭牲的血，抹在求洁净的人的右耳垂上、右手的大拇指上和右脚的大脚趾上。
LEV|14|15|祭司要从那一罗革的油中，取一些倒在自己的左手掌里，
LEV|14|16|祭司要用右手指蘸在他左手掌的油里，在耶和华面前用手指弹七次。
LEV|14|17|祭司要把手掌里剩下的油抹在那求洁净的人的右耳垂上、右手的大拇指上和右脚的大脚趾上，在赎愆祭牲之血抹过的上面。
LEV|14|18|祭司手掌里剩下的油要抹在那求洁净的人的头上，祭司就在耶和华面前为他赎罪。
LEV|14|19|祭司要献赎罪祭，为那从不洁净中得洁净的人赎罪，然后要宰燔祭牲，
LEV|14|20|祭司要把燔祭和素祭献在坛上，祭司要为他赎罪，他就洁净了。
LEV|14|21|“他若贫穷，手头财力不及，就要取一只小公羊作赎愆祭，作摇祭为他赎罪。他也要把作为素祭的十分之一伊法调了油的细面，和一罗革的油，一同取来。
LEV|14|22|他又要照手头财力所及，取两只斑鸠或两只雏鸽，一只作赎罪祭，一只作燔祭。
LEV|14|23|第八天，为了使自己洁净，他要把这些祭物带到耶和华面前，在会幕的门口交给祭司。
LEV|14|24|祭司要把赎愆祭的羔羊和那一罗革的油一同在耶和华面前摇一摇，作为摇祭。
LEV|14|25|祭司要宰赎愆祭的羔羊，取一些赎愆祭牲的血，抹在那求洁净的人的右耳垂上、右手的大拇指上和右脚的大脚趾上。
LEV|14|26|祭司要把一些油倒在自己的左手掌里，
LEV|14|27|祭司要用右手指，把他左手掌里的油在耶和华面前弹七次。
LEV|14|28|祭司要把手掌里的油抹一些在那求洁净的人的右耳垂上、右手的大拇指上和右脚的大脚趾上，在赎愆祭牲之血抹过之处的上面。
LEV|14|29|祭司手掌里剩下的油要抹在那求洁净的人的头上，在耶和华面前为他赎罪。
LEV|14|30|那人又要照他手头财力所及，献上斑鸠中的一只或雏鸽中的一只，
LEV|14|31|照他手头财力所及，一只为赎罪祭，一只为燔祭，与素祭一同献上。祭司就在耶和华面前为他赎罪。
LEV|14|32|这是为患痲疯灾病，手头财力不及而求洁净的人所定的条例。”
LEV|14|33|耶和华吩咐 摩西 和 亚伦 说：
LEV|14|34|“你们到了我所赐给你们为业的 迦南 地，我若使你们所得为业之地的房屋发霉 ，
LEV|14|35|屋主就要去告诉祭司说：‘据我看，房屋似乎发霉了。’
LEV|14|36|祭司进去检查这霉之前，要吩咐把屋内的东西全部搬走，免得屋子里所有的东西成为不洁净。然后，祭司要进去检查房屋。
LEV|14|37|他要检查这霉，看哪，若屋子墙上的霉有发绿或发红凹入的斑纹，其现象深入墙内，
LEV|14|38|祭司就要出到屋子的门外，把屋子封锁七天。
LEV|14|39|第七天，祭司要再去检查，看哪，霉若在屋子的墙上扩散，
LEV|14|40|祭司要吩咐把发霉的石头挖出来，扔在城外不洁净之处。
LEV|14|41|他也要叫人刮屋内的四围，把刮出来的灰泥倒在城外不洁净之处。
LEV|14|42|他们要用别的石头取代挖出来的石头，用别的灰泥涂抹屋子。
LEV|14|43|“他挖出石头，刮了屋子，涂抹以后，霉若又在屋子里出现，
LEV|14|44|祭司就要进去检查，看哪，霉若在屋子里扩散，那就是有侵蚀性的霉在屋子里，是不洁净的。
LEV|14|45|他要拆毁屋子，把石头、木料和所有的灰泥都搬到城外不洁净之处。
LEV|14|46|屋子封锁的任何时候，进去的人必不洁净到晚上。
LEV|14|47|在屋子里躺卧的人必须把衣服洗净，在屋子里吃饭的人也必须把衣服洗净。
LEV|14|48|“屋子涂抹了之后，祭司若进去检查，看哪，霉没有在屋内扩散，就要宣布这房屋为洁净，因为霉已经消除了。
LEV|14|49|他要为洁净房屋取两只鸟和香柏木、朱红色纱，以及牛膝草，
LEV|14|50|用瓦器盛清水，把一只鸟宰在上面。
LEV|14|51|他要把香柏木、牛膝草、朱红色纱和那一只活鸟，都蘸在被宰的鸟血和清水中，用来弹屋子七次。
LEV|14|52|他要用鸟血、清水、活鸟、香柏木、牛膝草和朱红色纱洁净那房屋。
LEV|14|53|他要把活鸟在城外野地里放走。他要为房屋赎罪，房屋就洁净了。”
LEV|14|54|这条例是为痲疯灾病和疥疮，
LEV|14|55|衣服和房屋发霉，
LEV|14|56|以及皮肤肿胀、发疹、有斑点等，
LEV|14|57|用以分辨何时洁净，何时不洁净。这是痲疯病的条例。
LEV|15|1|耶和华吩咐 摩西 和 亚伦 说：
LEV|15|2|“你们要吩咐 以色列 人，对他们说：人若身体 患了漏症，他因这症就不洁净了。
LEV|15|3|这就是他因漏症而有的不洁净：无论是身体流出液体，或身体已经止住不再有液体，他都是不洁净的。
LEV|15|4|那患漏症的人所躺的床都不洁净，所坐的任何东西也不洁净。
LEV|15|5|凡摸他床的人，要洗衣服，用水洗澡，必不洁净到晚上。
LEV|15|6|人坐了漏症患者坐过的东西，他要洗衣服，用水洗澡，必不洁净到晚上。
LEV|15|7|人摸了漏症患者，他要洗衣服，用水洗澡，必不洁净到晚上。
LEV|15|8|若漏症患者吐唾沫在洁净的人身上，这人要洗衣服，用水洗澡，必不洁净到晚上。
LEV|15|9|漏症患者所骑的任何鞍子也不洁净。
LEV|15|10|凡摸了他坐过的任何东西，必不洁净到晚上；拿了这些东西的，要洗衣服，用水洗澡，必不洁净到晚上。
LEV|15|11|漏症患者若没有用水冲洗他的手，无论摸了谁，谁就要洗衣服，用水洗澡，必不洁净到晚上。
LEV|15|12|漏症患者所摸的瓦器必要打破；他所摸的一切木器必要用水冲洗。
LEV|15|13|“漏症患者的漏症痊愈了，就要为洁净自己计算七天，也要洗衣服，用清水洗身，就洁净了。
LEV|15|14|第八天，他要带两只斑鸠或两只雏鸽，来到耶和华面前，在会幕门口把鸟交给祭司。
LEV|15|15|祭司要献上一只为赎罪祭，一只为燔祭。祭司要因这人所患的漏症，在耶和华面前为他赎罪。
LEV|15|16|“人若遗精，他要用水洗全身，必不洁净到晚上。
LEV|15|17|无论是衣服或皮革，若沾染了精液，要用水洗净，必不洁净到晚上。
LEV|15|18|女人，若有男人与她同寝，沾染了精液，二人要用水洗澡，必不洁净到晚上。”
LEV|15|19|“女人月经期间，有血从体内流出，她必不洁净七天；凡摸她的，必不洁净到晚上。
LEV|15|20|在不洁净期间，女人所躺的东西都不洁净，所坐的任何东西也不洁净。
LEV|15|21|凡摸她床的，要洗衣服，用水洗澡，必不洁净到晚上；
LEV|15|22|凡摸她坐过的东西的，要洗衣服，用水洗澡，必不洁净到晚上；
LEV|15|23|不论是床，或她坐过的东西，人摸了，必不洁净到晚上。
LEV|15|24|男人若和这女人同寝，沾了她的不洁净，就不洁净七天，所躺的床也都不洁净。
LEV|15|25|“女人若在经期之外仍然流血多日，或是经期过长，她在流血的一切日子都不洁净，和她在经期的日子不洁净一样。
LEV|15|26|在流血的日子，她所躺的床、所坐的任何东西都不洁净，和在月经期间不洁净一样。
LEV|15|27|凡摸这些东西的，就不洁净；他要洗衣服，用水洗澡，必不洁净到晚上。
LEV|15|28|这女人的血漏若痊愈了，就要计算七天，然后才洁净。
LEV|15|29|第八天，她要取两只斑鸠或两只雏鸽，带到会幕门口祭司那里。
LEV|15|30|祭司要献一只为赎罪祭，一只为燔祭。祭司要因这女人血漏的不洁净，在耶和华面前为她赎罪。
LEV|15|31|“你们要使 以色列 人与他们的不洁净隔离，免得他们玷污我在他们中间的帐幕，因自己的不洁净死亡。”
LEV|15|32|这条例是为漏症患者或遗精而不洁净者，
LEV|15|33|女人经期的不洁，男女患漏症，以及男人与不洁净女人同寝而立的。
LEV|16|1|亚伦 的两个儿子靠近耶和华面前，死了。他们死后，耶和华吩咐 摩西 ；
LEV|16|2|耶和华对 摩西 说：“你要吩咐你哥哥 亚伦 ，不可随时进入圣所的幔子内、到柜盖 前，免得他死亡，因为我在柜盖上的云中显现。
LEV|16|3|亚伦 进圣所要带这些：一头公牛犊为赎罪祭，一只公绵羊为燔祭。
LEV|16|4|他要穿上细麻布圣内袍，把细麻布裤子穿在身上，腰束细麻布带子，头戴细麻布礼冠；这些都是圣服。他要用水洗身，然后穿上圣服。
LEV|16|5|他要从 以色列 会众中取两只公山羊为赎罪祭，一只公绵羊为燔祭。
LEV|16|6|“亚伦要把他自己赎罪祭的公牛献上，为自己和家人赎罪；
LEV|16|7|也要把两只公山羊牵到耶和华面前，安置在会幕的门口。
LEV|16|8|亚伦 要为那两只山羊抽签，一签归给耶和华，一签归给 阿撒泻勒 。
LEV|16|9|亚伦 要把那抽中归给耶和华的山羊牵来献为赎罪祭，
LEV|16|10|至于抽中归给 阿撒泻勒 的山羊，却要活着安放在耶和华面前，用以赎罪，然后送到旷野去，归给 阿撒泻勒 。
LEV|16|11|“ 亚伦 要把他自己赎罪祭的公牛献上，为自己和家人赎罪，他要宰作自己赎罪祭的公牛。
LEV|16|12|他要从耶和华面前的坛上取盛满火炭的香炉，再拿一捧捣细的香料，把这些都带入幔子内。
LEV|16|13|在耶和华面前，他要把香放在火上，使香的烟云遮着法柜上的盖子，免得他死亡。
LEV|16|14|他要取一些公牛的血，用手指弹在柜盖的前面，就是东面，又在柜盖的前面用手指弹血七次。
LEV|16|15|“他要宰那只为百姓作赎罪祭的公山羊，把羊的血带入幔子内，把血弹在柜盖的上面和前面，好像弹公牛的血一样。
LEV|16|16|因 以色列 人的不洁净和过犯，就是他们一切的罪，他要为圣所赎罪；因会幕在他们不洁净之中，他也要为会幕照样做。
LEV|16|17|他进圣所赎罪的时候，会幕里都不准有人，直等到他为自己和家人，以及 以色列 全会众赎了罪出来。
LEV|16|18|他出来后，要到耶和华面前的祭坛那里，为坛赎罪。他要取一些公牛的血和公山羊的血，抹在坛周围的四个翘角上。
LEV|16|19|他也要用手指把血弹在坛上七次，使坛从 以色列 人的不洁净中得以洁净，成为圣。”
LEV|16|20|“ 亚伦 为圣所和会幕，以及祭坛赎罪后，就要把那只活的公山羊牵来。
LEV|16|21|他的双手要按在活的山羊的头上，承认 以色列 人所有的罪孽过犯，就是他们一切的罪，把这些罪都归在羊的头上，再指派一个人把它送到旷野去。
LEV|16|22|这羊要担当他们一切的罪孽，带到无人之地；那人要把羊送到旷野去。
LEV|16|23|“ 亚伦 要进入会幕，把他进圣所时所穿的细麻布衣服脱下，放在那里，
LEV|16|24|又要在圣处用水洗身，穿上衣服出来，把自己的燔祭和百姓的燔祭献上，为自己和百姓赎罪。
LEV|16|25|赎罪祭牲的脂肪要烧在坛上。
LEV|16|26|那放走山羊归给 阿撒泻勒 的人要洗衣服，用水洗身，然后才可以回到营里。
LEV|16|27|作赎罪祭的公牛和作赎罪祭的公山羊的血被带入圣所赎罪之后，就要把这牛羊搬到营外，皮、肉、粪都用火焚烧。
LEV|16|28|焚烧的人要洗衣服，用水洗身，然后才可以回到营里。”
LEV|16|29|“这是你们永远的定例：每年七月初十，你们要刻苦己心；无论是本地人，是寄居在你们中间的外人，任何工都不可做。
LEV|16|30|因为这日要为你们赎罪，洁净你们，使你们脱离一切的罪，在耶和华面前得以洁净。
LEV|16|31|这日你们要守完全安息的安息日，刻苦己心；这是永远的定例。
LEV|16|32|那受膏接续他父亲担任圣职的祭司要赎罪，穿上细麻布衣服，就是圣衣，
LEV|16|33|为至圣所和会幕赎罪，为祭坛赎罪，并要为祭司和会众的全体百姓赎罪。
LEV|16|34|这要作你们永远的定例：因 以色列 人一切的罪，要一年一次为他们赎罪。”于是， 亚伦 照耶和华所吩咐 摩西 的做了 。
LEV|17|1|耶和华吩咐 摩西 说：
LEV|17|2|“你要吩咐 亚伦 和他儿子，以及 以色列 众人，对他们说，耶和华所吩咐的话是这样：
LEV|17|3|凡 以色列 家中的人宰公牛，或小绵羊，或山羊，无论是在营内或营外，
LEV|17|4|若不把牲畜牵到会幕门口耶和华的帐幕前，献给耶和华为供物，所流的血必归到那人身上。他既使血流出，就要从百姓中剪除。
LEV|17|5|这是为要使 以色列 人把他们在野地里所宰的祭牲带来，带到耶和华前，会幕门口祭司那里，宰杀这些祭牲，把它们献给耶和华为平安祭。
LEV|17|6|祭司要在会幕门口，把血洒在耶和华的祭坛上，把脂肪焚烧，献给耶和华为馨香的祭。
LEV|17|7|他们不可再宰杀祭牲献给他们行淫所随从的山羊鬼魔。这要作他们世世代代永远的定例。
LEV|17|8|“你要对他们说：凡 以色列 家中的任何人，或寄居在他们中间的外人献燔祭或祭物，
LEV|17|9|若不带到会幕门口献给耶和华，那人必从百姓中剪除。
LEV|17|10|“凡 以色列 家中的任何人，或寄居在他们中间的外人，吃任何的血，我必向那吃血的人变脸，把他从百姓中剪除。
LEV|17|11|因为动物的生命是在血中。我把这血赐给你们，可以在祭坛上为你们的生命赎罪；因为血就是生命，能够赎罪。
LEV|17|12|因此，我对 以色列 人说：你们都不可吃血；寄居在你们中间的外人也不可吃血。
LEV|17|13|凡 以色列 人，或寄居在他们中间的外人，猎取了可吃的飞禽走兽，必须把它的血放出来，用土掩盖。
LEV|17|14|“因一切动物的生命，它的血就是它的生命。所以我对 以色列 人说：无论什么动物的血，你们都不可吃，因为一切动物的生命就是它的血。凡吃血的必被剪除。
LEV|17|15|无论是本地人，是寄居的，若吃了自然死去或被野兽撕裂的动物，要洗衣服，用水洗澡，必不洁净到晚上，晚上就洁净了。
LEV|17|16|但他若不洗衣服，也不洗身，就要担当自己的罪孽。”
LEV|18|1|耶和华吩咐 摩西 说：
LEV|18|2|“你要吩咐 以色列 人，对他们说：我是耶和华－你们的上帝。
LEV|18|3|你们不可做你们从前住 埃及 地的人所做的，也不可做我要领你们去的 迦南 地的人所做的。你们不可照他们的习俗行。
LEV|18|4|你们要遵行我的典章，谨守我的律例，按此而行。我是耶和华－你们的上帝。
LEV|18|5|你们要谨守我的律例典章；遵行的人就必因此得生。我是耶和华。
LEV|18|6|“任何人都不可亲近骨肉之亲，露其下体。我是耶和华。
LEV|18|7|你父亲的下体，就是你母亲的下体，你不可露；她是你的母亲，不可露她的下体。
LEV|18|8|不可露你继母的下体，就是你父亲的下体。
LEV|18|9|你姊妹的下体，或是同父异母的，或是同母异父的，无论生在家或生在外的，都不可露她们的下体。
LEV|18|10|不可露你孙女或外孙女的下体，因为她们的下体就是你自己的下体。
LEV|18|11|你继母为你父亲所生的女儿是你的姊妹，不可露她的下体。
LEV|18|12|不可露你姑母的下体；她是你父亲的骨肉之亲。
LEV|18|13|不可露你姨母的下体；她是你母亲的骨肉之亲。
LEV|18|14|不可露你叔伯的下体，不可亲近他的妻子；她是你的叔母、伯母。
LEV|18|15|不可露你媳妇的下体，她是你儿子的妻，不可露她的下体。
LEV|18|16|不可露你兄弟妻子的下体，这是你兄弟的下体。
LEV|18|17|不可露妇人的下体，又露她女儿的下体，也不可娶她的孙女或外孙女，露她们的下体；她们是骨肉之亲 。这是邪恶的事。
LEV|18|18|你妻子还活着的时候，不可另娶她的姊妹与她作对，露她姊妹的下体。
LEV|18|19|“不可亲近经期中不洁净的女人，露她的下体。
LEV|18|20|不可跟邻舍的妻交合，因她玷污自己。
LEV|18|21|不可使你儿女经火献给 摩洛 ，也不可亵渎你上帝的名。我是耶和华。
LEV|18|22|不可跟男人同寝，像跟女人同寝；这是可憎恶的事。
LEV|18|23|不可跟兽交合，因它玷污自己。女人也不可站在兽前，与它交合；这是逆性的事。
LEV|18|24|“在这一切的事上，你们都不可玷污自己，因为我在你们面前所逐出的列国，在这一切的事上玷污了自己。
LEV|18|25|连地也玷污了，我惩罚那地的罪孽，地就吐出它的居民来。
LEV|18|26|但你们要遵守我的律例典章。这一切可憎恶的事，无论是本地人或寄居在你们中间的外人，都不可以做。
LEV|18|27|在你们之前居住那地的人做了这一切可憎恶的事，地就玷污了。
LEV|18|28|不要让地因你们玷污了它而把你们吐出来，像吐出在你们之前的国一样。
LEV|18|29|无论是谁，若做了这其中一件可憎恶的事，必从百姓中剪除。
LEV|18|30|你们要遵守我的吩咐，免得你们随从那些可憎的习俗，就是在你们之前的人所做的，玷污了自己。我是耶和华－你们的上帝。”
LEV|19|1|耶和华吩咐 摩西 说：
LEV|19|2|“你要吩咐 以色列 全会众，对他们说：你们要成为圣，因为我耶和华－你们的上帝是神圣的。
LEV|19|3|你们各人都当孝敬父母，也要守我的安息日。我是耶和华－你们的上帝。
LEV|19|4|你们不可转向虚无的神明，也不可为自己铸造神像。我是耶和华－你们的上帝。
LEV|19|5|“你们宰杀祭牲献平安祭给耶和华的时候，要献得使你们可蒙悦纳。
LEV|19|6|这祭物要在献的当天或第二天吃；若有剩到第三天的，就要用火焚烧。
LEV|19|7|第三天若再吃，这祭物是不洁净的，必不蒙悦纳。
LEV|19|8|吃的人必担当自己的罪孽，因为他亵渎了耶和华的圣物，这人必从百姓中剪除。
LEV|19|9|“你们在自己的地收割庄稼时，不可割尽田的角落，也不可拾取庄稼所掉落的。
LEV|19|10|不可摘尽葡萄园的葡萄，也不可拾取葡萄园中掉落的葡萄，要把它们留给穷人和寄居的。我是耶和华－你们的上帝。
LEV|19|11|“你们不可偷盗，不可欺骗，也不可彼此说谎。
LEV|19|12|不可指着我的名起假誓，亵渎你上帝的名。我是耶和华。
LEV|19|13|“不可欺压你的邻舍，也不可偷盗。雇工的工钱不可在你那里过夜，留到早晨。
LEV|19|14|不可咒骂聋子，也不可将绊脚石放在盲人面前。你要敬畏你的上帝。我是耶和华。
LEV|19|15|“你们审判的时候，不可不公正；不可偏护贫穷人，也不可看重有权势人的脸，总要公平审判你的邻舍。
LEV|19|16|不可在百姓中到处搬弄是非，不可陷害邻舍的性命 。我是耶和华。
LEV|19|17|“不可心里恨你的弟兄；要指摘你的邻舍，免得因他承担罪过。
LEV|19|18|不可报仇，也不可埋怨你本国的子民。你要爱邻如己。我是耶和华。
LEV|19|19|“你们要遵守我的律例。不可使你的牲畜与异类交配；不可在你的田地播下两样的种子；也不可穿两种原料做成的衣服。
LEV|19|20|“若有人与女子同寝交合，而她是婢女，许配了丈夫，尚未被赎或得自由，就要受到惩罚，却不可把他们处死，因为婢女还没有得自由。
LEV|19|21|男的要把赎愆祭，就是一只公绵羊牵到耶和华面前，会幕的门口。
LEV|19|22|祭司要用赎愆祭的羊在耶和华面前为他所犯的罪赎罪，他所犯的罪就必蒙赦免。
LEV|19|23|“你们到了 迦南 地，栽种各样的果树，就要把所结的果子当作不洁净的 ；三年之内，你们要把它视为不洁净，是不可吃的。
LEV|19|24|但第四年所结的果子全是圣的，用以赞美耶和华 。
LEV|19|25|第五年，你们就可以吃树上的果子，使树给你们结出更多的果子。我是耶和华－你们的上帝。
LEV|19|26|“你们不可吃带血的食物。不可占卜，也不可观星象。
LEV|19|27|头的周围 不可剃，胡须的周围不可损坏。
LEV|19|28|不可为死人割划自己的身体，也不可在身上刺花纹。我是耶和华。
LEV|19|29|“不可侮辱你的女儿，使她沦为娼妓，免得这地行淫乱，地就充满了邪恶。
LEV|19|30|你们要谨守我的安息日，敬畏我的圣所。我是耶和华。
LEV|19|31|“不可转向招魂的，也不可求问行巫术的，免得被他们玷污。我是耶和华－你们的上帝。
LEV|19|32|“在白发的人面前，你要站起来，要尊敬老人；要敬畏你的上帝，我是耶和华。
LEV|19|33|“若有外人寄居在你们的地上和你同住，不可欺负他。
LEV|19|34|寄居在你们那里的外人，你们要看他如本地人，并要爱他如己，因为你们在 埃及 地也作过寄居的。我是耶和华－你们的上帝。
LEV|19|35|“你们审判的时候，不可用不公正的度量衡。
LEV|19|36|你们要用公正的天平、公正的法码、公正的伊法和公正的欣。我是耶和华－你们的上帝，曾把你们从 埃及 地领出来。
LEV|19|37|你们要谨守我一切的律例典章，遵行它们。我是耶和华。”
LEV|20|1|耶和华吩咐 摩西 说：
LEV|20|2|“你要对 以色列 人说：凡 以色列 人，或是寄居在 以色列 的外人，把自己儿女献给 摩洛 的，必被处死；本地的百姓要用石头打死他。
LEV|20|3|我也要向那人变脸，把他从百姓中剪除，因为他把儿女献给 摩洛 ，玷污了我的圣所，亵渎了我的圣名。
LEV|20|4|那人把儿女献给 摩洛 ，本地的百姓若假装没看见，不把他处死，
LEV|20|5|我就要向这人和他的家人变脸，把他和所有跟随他与 摩洛 行淫的人都从百姓中剪除。
LEV|20|6|“人若转向招魂的和行巫术的，随从他们行淫，我就要向这人变脸，把他从百姓中剪除。
LEV|20|7|你们要使自己分别为圣，要成为圣，因为我是耶和华－你们的上帝。
LEV|20|8|你们要谨守我的律例，遵行它们；我是使你们分别为圣的耶和华。
LEV|20|9|凡咒骂父母的，必被处死；他咒骂了父母，他的血要归在他身上。
LEV|20|10|“凡与有夫之妇行奸淫，就是与邻舍的妻子行奸淫的，奸夫淫妇必被处死。
LEV|20|11|人若与继母同寝，就是露了父亲的下体，二人必被处死，血要归在他们身上。
LEV|20|12|人若与媳妇同寝，二人必被处死；他们行了乱伦的事，血要归在他们身上。
LEV|20|13|男人若跟男人同寝，像跟女人同寝，他们二人行了可憎恶的事，必被处死，血要归在他们身上。
LEV|20|14|人若娶妻，又娶妻子的母亲，这是邪恶的事；要把这三人用火焚烧，在你们中间除去这邪恶。
LEV|20|15|人若与兽交合，必被处死；你们也要杀死那兽。
LEV|20|16|女人若与兽亲近，与它交合，你要把那女人和兽杀死；他们必被处死，血要归在他们身上。
LEV|20|17|“人若娶自己的姊妹，或是同父异母的，或是同母异父的，彼此见了下体，这是可耻的事；他们必在自己百姓眼前被剪除。他露了姊妹的下体，必担当自己的罪孽。
LEV|20|18|若有人跟经期中的妇人同寝，露了她的下体，暴露妇人的血源，妇人也露了自己的血源，二人必从百姓中剪除。
LEV|20|19|不可露姨母或姑母的下体，因为这是露了骨肉之亲的下体，他们必担当自己的罪孽。
LEV|20|20|人若与叔伯之妻同寝，就露了他叔伯的下体，他们必担当自己的罪，必没有子女而死。
LEV|20|21|人若娶了自己兄弟的妻子，就露了他兄弟的下体，这是不洁净的事，他们必没有子女。
LEV|20|22|“你们要谨守我一切的律例典章，遵行它们，免得我领你们去住的那地把你们吐出来。
LEV|20|23|我在你们面前所逐出的国民，你们不可随从他们的风俗。因为他们行了这一切的事，所以我厌恶他们。
LEV|20|24|但我对你们说过，你们要承受他们的土地；我要把这流奶与蜜之地赐给你们，作为你们的产业。我是耶和华－你们的上帝，是把你们从万民中分别出来的。
LEV|20|25|你们要分辨洁净和不洁净的飞禽走兽；不可因我定为不洁净的飞禽走兽，或爬行在土地上的任何生物，使自己成为可憎恶的。
LEV|20|26|你们要归我为圣，因为－我耶和华是神圣的；我把你们从万民中分别出来，作我的子民。
LEV|20|27|“无论男女，是招魂的或行巫术的，他们必被处死。人要用石头打死他们，血要归在他们身上。”
LEV|21|1|耶和华对 摩西 说：“你要告诉 亚伦 子孙作祭司的，对他们说：祭司不可为自己百姓中的死人玷污自己，
LEV|21|2|除非是他的骨肉之亲，他的父母、儿女、兄弟、
LEV|21|3|或未出嫁还是处女的姊妹，因她是至亲，才可以玷污自己。
LEV|21|4|祭司既然在自己百姓中为首，就不可从俗玷污自己 。
LEV|21|5|“不可使头光秃，不可剃除胡须的边缘，也不可割划自己的身体。
LEV|21|6|他们要归上帝为圣，不可亵渎他们上帝的名，因为耶和华的火祭，就是上帝的食物，是他们献的，所以他们要成为圣。
LEV|21|7|“祭司不可娶妓女，或被玷污的女人为妻，也不可娶被休的妇人为妻，因为他是归上帝为圣的。
LEV|21|8|你要使祭司分别为圣，因为他献你上帝的食物。你要以他为圣，因为我是使你们分别为圣 的耶和华，是神圣的。
LEV|21|9|“祭司的女儿若行淫玷污自己，就侮辱了父亲，要用火将她焚烧。
LEV|21|10|“在弟兄中作大祭司的，头上倒了膏油，承接圣职，穿了圣衣，不可蓬头散发，也不可撕裂衣服；
LEV|21|11|不可挨近任何死尸，即使为了父母也不可玷污自己。
LEV|21|12|他不可出圣所，免得亵渎了上帝的圣所，因为在他身上有上帝的膏油为圣冕。我是耶和华。
LEV|21|13|他要娶处女为妻。
LEV|21|14|大祭司不可娶寡妇，被休的妇人，或被玷污的妓女为妻；他只可以娶自己百姓中的处女为妻。
LEV|21|15|他不可在自己百姓中侮辱他的儿女，因为我是使他分别为圣的耶和华。”
LEV|21|16|耶和华吩咐 摩西 说：
LEV|21|17|“你吩咐 亚伦 说：你世世代代的后裔，凡有残疾的都不可近前来献上帝的食物。
LEV|21|18|因为凡有残疾的，无论是失明的、瘸腿的、五官不正的、肢体之一过长的、
LEV|21|19|断脚的、断手的、
LEV|21|20|驼背的、侏儒的、有眼疾的、长癣的、长疥的，或是睾丸压伤的，都不可近前来。
LEV|21|21|亚伦 祭司的后裔，凡有残疾的都不可近前来献耶和华的火祭。他有残疾，不可近前来献上帝的食物。
LEV|21|22|上帝的食物，无论是圣的，或是至圣的，他都可以吃。
LEV|21|23|但他不可进到幔子前，也不可挨近祭坛前，因为他有残疾，免得他亵渎我的圣所。我是使他们分别为圣的耶和华。”
LEV|21|24|于是， 摩西 吩咐了 亚伦 和他的儿子，以及 以色列 众人。
LEV|22|1|耶和华吩咐 摩西 说：
LEV|22|2|“你要吩咐 亚伦 和他子孙说：你们要谨慎处理 以色列 人所分别为圣，归给我的圣物，免得亵渎我的圣名。我是耶和华。
LEV|22|3|你要对他们说：你们世世代代的后裔，凡不洁净，却挨近 以色列 人所分别为圣，归给耶和华的圣物，那人必从我面前剪除。我是耶和华。
LEV|22|4|亚伦 的后裔中，凡有痲疯病的，或患漏症的，都不可吃圣物，直等他洁净了。无论谁摸了那因尸体而不洁净的东西，或遗精的人，
LEV|22|5|或摸到任何使他不洁净的群聚动物或使他不洁净的人，无论那人有什么不洁净，
LEV|22|6|摸了这些的人必不洁净到晚上；若不用水洗身，就不可吃圣物。
LEV|22|7|日落的时候，他就洁净了，然后可以吃圣物，因为这是他的食物。
LEV|22|8|自然死去的或被野兽撕裂的，他不可吃，免得玷污自己。我是耶和华。
LEV|22|9|他们要遵守我的吩咐，免得因亵渎圣物 ，担当自己的罪而死。我是使他们分别为圣的耶和华。
LEV|22|10|“任何外人都不可吃圣物；寄居在祭司家的，或雇工，都不可吃圣物。
LEV|22|11|若是祭司用自己的银钱买来的人，就可以吃圣物；在他家出生的人也可以吃他的食物。
LEV|22|12|祭司的女儿若嫁给外人，就不可吃举祭的圣物。
LEV|22|13|但祭司的女儿若成为寡妇或被休，又没有后裔，她回到父家，好像年轻的时候，就可以吃她父亲的食物。只是任何外人都不可吃它。
LEV|22|14|若有人误吃了圣物，要把圣物加上五分之一交给祭司。
LEV|22|15|祭司不可亵渎 以色列 人献给耶和华的圣物，
LEV|22|16|免得他们因吃圣物而自取罪孽。我是使他们分别为圣的耶和华。”
LEV|22|17|耶和华吩咐 摩西 说：
LEV|22|18|“你要吩咐 亚伦 和他子孙，以及 以色列 众人，对他们说： 以色列 家中的人，或在 以色列 中寄居的 ，若要献供物给耶和华作燔祭，无论是为所许的愿或是甘心献的，
LEV|22|19|就要将一头公的，没有残疾的牛，或绵羊，或山羊献上，这样你们才蒙悦纳。
LEV|22|20|凡有残疾的，你们不可献上，因为这样你们必不蒙悦纳。
LEV|22|21|若有人从牛群或羊群中，将平安祭献给耶和华，无论是为还所许特别的愿，或是甘心献的，所献的必须是健康、无任何残疾的，才蒙悦纳。
LEV|22|22|凡瞎眼的、受伤的、断腿的、溃烂的、长癣的、长疥的，都不可献给耶和华，不可在坛上作为火祭献给耶和华。
LEV|22|23|无论是公牛或小绵羊，若一条腿太长或太短，只可作甘心祭献上；若用来还愿，就不蒙悦纳。
LEV|22|24|凡睾丸损伤，或压碎，或破裂，或阉割的，都不可献给耶和华；不可在你们的地上行这事。
LEV|22|25|从外人的手里得到任何这类的动物，也不可献上作你们上帝的食物；因为它们有缺陷，有残疾，它们必不为你们而蒙悦纳。”
LEV|22|26|耶和华吩咐 摩西 说：
LEV|22|27|“刚出生的公牛，或绵羊，或山羊，七天当跟着它的母亲；从第八天起，可以当供物作为耶和华的火祭，这是蒙悦纳的。
LEV|22|28|无论是牛或羊，不可在同一日宰它和它的小牛小羊。
LEV|22|29|你们宰杀祭牲献感谢祭给耶和华，要献得使你们可蒙悦纳；
LEV|22|30|要在当天吃，一点也不可留到早晨。我是耶和华。
LEV|22|31|“你们要谨守我的诫命，遵行它们。我是耶和华。
LEV|22|32|你们不可亵渎我的圣名；我在 以色列 人中要被尊为圣。我是使你们分别为圣的耶和华，
LEV|22|33|曾把你们从 埃及 地领出来，作你们的上帝。我是耶和华。”
LEV|23|1|耶和华吩咐 摩西 说：
LEV|23|2|“你要吩咐 以色列 人，对他们说：以下是我的节期，是你们要宣告为圣会的耶和华的节期。”
LEV|23|3|“六日要做工，第七日是完全安息的安息日，要有圣会；你们任何工都不可做。这是在你们一切的住处向耶和华当守的安息日。”
LEV|23|4|“以下是你们要按时宣告为圣会的耶和华的节期。”
LEV|23|5|“正月十四日黄昏的时候 ，是向耶和华守的逾越节。
LEV|23|6|这月的十五日是向耶和华守的除酵节；你们要吃无酵饼七日。
LEV|23|7|第一日要有圣会，任何劳动的工都不可做；
LEV|23|8|要将火祭献给耶和华七日。第七日要有圣会，任何劳动的工都不可做。”
LEV|23|9|耶和华吩咐 摩西 说：
LEV|23|10|“你要吩咐 以色列 人，对他们说：你们到了我赐给你们的地，收割庄稼的时候，要把初熟庄稼中的一捆拿来给祭司。
LEV|23|11|他要把这捆在耶和华面前摇一摇，使你们蒙悦纳。祭司要在安息日的次日把这捆摇一摇。
LEV|23|12|摇这捆的那一日，你们要献一只一岁没有残疾的小公绵羊，给耶和华作燔祭。
LEV|23|13|同献的素祭是十分之二伊法调了油的细面，作为献给耶和华馨香的火祭；同献的浇酒祭是四分之一欣酒。
LEV|23|14|无论是饼，是烘熟的谷物，是新穗子，你们都不可吃；直等到你们把这供物带来献给你们上帝的那一天，才可以吃。在你们一切的住处，这要成为你们世世代代永远的定例。”
LEV|23|15|“你们要从安息日的次日，就是献那捆庄稼为摇祭的那日起，计算足足的七个安息日。
LEV|23|16|到第七个安息日的次日，共计五十天，你们要将新的素祭献给耶和华。
LEV|23|17|要从你们的住处取十分之二伊法细面，加酵烤成两个摇祭的饼，作为初熟之物献给耶和华。
LEV|23|18|又要将七只一岁没有残疾的羔羊、一头公牛犊、两只公绵羊和饼一同奉上。这些要和素祭和浇酒祭一同作为燔祭献给耶和华，作馨香的火祭献给耶和华。
LEV|23|19|你们要献一只公山羊为赎罪祭，两只一岁的小公绵羊为平安祭。
LEV|23|20|祭司要把这些和初熟庄稼做成的饼，与两只小公绵羊一同在耶和华面前摇一摇，作为摇祭。这些献给耶和华的圣物是归给祭司的。
LEV|23|21|在这一日，你们要宣告圣会；任何劳动的工都不可做。在你们一切的住处，这要成为你们世世代代永远的定例。
LEV|23|22|“你们在自己的地收割庄稼时，不可割尽田的角落，也不可拾取庄稼所掉落的，要把它们留给穷人和寄居的。我是耶和华－你们的上帝。”
LEV|23|23|耶和华吩咐 摩西 说：
LEV|23|24|“你要吩咐 以色列 人说：七月初一，你们要守为完全安息的日子，要吹角作纪念，当有圣会。
LEV|23|25|任何劳动的工都不可做；要将火祭献给耶和华。”
LEV|23|26|耶和华吩咐 摩西 说：
LEV|23|27|“但是，七月初十是赎罪日；你们要守为圣会，刻苦己心，并要将火祭献给耶和华。
LEV|23|28|在这一日，任何工都不可做；因为这是赎罪日，要在耶和华－你们的上帝面前赎罪。
LEV|23|29|在这一日，凡不刻苦己心的，必从百姓中剪除。
LEV|23|30|凡在这一日做任何工的，我必将他从百姓中除灭。
LEV|23|31|任何工你们都不可做。在你们一切的住处，这要成为你们世世代代永远的定例。
LEV|23|32|你们要守这日为完全安息的安息日，刻苦己心；从这月初九晚上到次日晚上，你们要守为安息日。”
LEV|23|33|耶和华吩咐 摩西 说：
LEV|23|34|“你要吩咐 以色列 人说：这七月十五日是住棚节，要向耶和华守这节七日。
LEV|23|35|第一日当有圣会，任何劳动的工都不可做。
LEV|23|36|要将火祭献给耶和华七日。第八日当守圣会，并要献火祭给耶和华。这是严肃会，任何劳动的工都不可做。
LEV|23|37|“这是耶和华的节期，就是你们要宣告为圣会的节期；要将火祭，就是燔祭、素祭、祭物和浇酒祭，按照每日的规定献给耶和华。
LEV|23|38|除此之外，还有耶和华的安息日，你们献给耶和华的供物，一切的还愿祭，和一切的甘心祭。
LEV|23|39|“但是，从七月十五日起，你们收藏了地的出产之后，要守耶和华的节期七日。第一日为要完全安息，第八日也要完全安息。
LEV|23|40|第一日，你们要拿美好树上的果子、棕树枝、树叶茂密的枝条和河边的柳枝，在耶和华－你们的上帝面前欢乐七日。
LEV|23|41|每年你们要向耶和华守这节七日。你们在七月里所守的节，要成为世世代代永远的定例。
LEV|23|42|你们要住在棚里七日；凡 以色列 家出生的人都要住在棚里，
LEV|23|43|好叫你们世世代代知道，我领 以色列 人出 埃及 地的时候，曾使他们住在棚里。我是耶和华－你们的上帝。”
LEV|23|44|于是， 摩西 向 以色列 人颁布了耶和华的节期。
LEV|24|1|耶和华吩咐 摩西 说：
LEV|24|2|“你要吩咐 以色列 人，把那捣成的纯橄榄油拿来给你，用以点灯，使灯经常点着。
LEV|24|3|在会幕中法柜前的幔子外， 亚伦 从晚上到早晨要在耶和华面前照管这灯。这要成为你们世世代代永远的定例。
LEV|24|4|他要在耶和华面前经常照管纯金 灯台上的灯。”
LEV|24|5|“你要取细面，烤成十二个饼，每个用十分之二伊法。
LEV|24|6|要把饼排成两行 ，每行六个，供在耶和华面前的纯金桌子上。
LEV|24|7|再把纯乳香撒在每行饼上，作为纪念，是献给耶和华为食物的火祭。
LEV|24|8|每个安息日， 亚伦 要把饼不间断地供在耶和华面前。这是 以色列 人永远的约。
LEV|24|9|这饼要归给 亚伦 和他的子孙。他们要在圣处吃这饼，因为在献给耶和华的火祭中，这饼是至圣的，归给他作永远当得的份。”
LEV|24|10|有一个 以色列 妇人的儿子，他父亲是 埃及 人。有一日他出去，到 以色列 人中。这 以色列 妇人的儿子和一个 以色列 人在营里争吵。
LEV|24|11|以色列 妇人的儿子诅咒，亵渎了圣名。有人把他送到 摩西 那里。他的母亲名叫 示罗密 ，是 但 支派 底伯利 的女儿。
LEV|24|12|他们把这人收押在监里，等候耶和华指示的话。
LEV|24|13|耶和华吩咐 摩西 说：
LEV|24|14|“把那诅咒的人带到营外。凡听见的人都要把手放在他头上，全会众要用石头打死他。
LEV|24|15|你要吩咐 以色列 人说：凡诅咒上帝的，必要担当自己的罪。
LEV|24|16|亵渎耶和华名的，必被处死；全会众必须用石头打死他。无论是寄居的，是本地人，他亵渎圣名的时候必被处死。
LEV|24|17|“打死人的，必被处死；
LEV|24|18|打死牲畜的，必赔上牲畜，以命偿命。
LEV|24|19|人若伤害邻舍以致残疾，他怎样做，也要照样向他做：
LEV|24|20|以伤还伤，以眼还眼，以牙还牙。他怎样使人有残疾，也要照样向他做。
LEV|24|21|打死牲畜的，必赔上牲畜；打死人的，必被处死。
LEV|24|22|无论是寄居的，是本地人，都依照同一条例。我是耶和华－你们的上帝。”
LEV|24|23|于是， 摩西 吩咐 以色列 人，他们就把那诅咒的人带到营外，用石头打死。 以色列 人就照耶和华所吩咐 摩西 的做了。
LEV|25|1|耶和华在 西奈山 吩咐 摩西 说：
LEV|25|2|“你要吩咐 以色列 人，对他们说：你们到了我所赐你们那地的时候，地要休耕，向耶和华守安息。
LEV|25|3|你们六年要耕种田地，六年要修整葡萄园，收藏地的出产。
LEV|25|4|第七年，地要守完全安息的安息年，就是向耶和华守安息。你们不可耕种田地，也不可修整葡萄园。
LEV|25|5|不可收割自然生长的庄稼，也不可摘取没有修剪的葡萄树上的葡萄。这年，地要完全安息。
LEV|25|6|地在安息年所长出的，要给你和你的奴仆、使女、雇工，以及寄居在你那里的外人作食物。
LEV|25|7|所有的出产也要给你的牲畜和你地上的走兽作食物。”
LEV|25|8|“你要计算七个安息年，就是七个七年。这就成为你的七个安息年，一共四十九年。
LEV|25|9|七月初十，你要大声吹角；这是赎罪日，你要在全地吹角。
LEV|25|10|你们要以第五十年为圣年，在全地向所有的居民宣告自由。这是你们的禧年，各人的产业要归还自己，各人要归回自己的家。
LEV|25|11|第五十年要作为你们的禧年。你们不可耕种，不可收割自然生长的庄稼，也不可摘取没有修剪的葡萄树上的葡萄。
LEV|25|12|因为这是禧年，是你们的圣年；你们要吃地中自然生长的农作物。
LEV|25|13|“这禧年，你们各人的产业要归还自己。
LEV|25|14|无论你卖什么给邻舍，或从邻舍的手中买什么，彼此不可亏负。
LEV|25|15|你要按照禧年后的年数向邻舍买；他要按照可收成的年数卖给你；
LEV|25|16|年数越多，价钱就越高；年数越少，价钱就越低，因为他卖给你的是收成的数量。
LEV|25|17|你们彼此不可亏负，只要敬畏你的上帝，因为我是耶和华－你们的上帝。”
LEV|25|18|“你们要遵行我的律例，谨守我的典章，遵行它们，就可以在那地上安然居住。
LEV|25|19|地必出产果实，你们可以吃饱，在那地上安然居住。
LEV|25|20|你们若说：‘看哪，第七年我们不耕种，也不收藏农作物，我们吃什么呢？’
LEV|25|21|我必在第六年发令赐福给你们，地就长出三年的农作物来。
LEV|25|22|第八年你们要耕种，也要吃陈粮；等到第九年农作物收成的时候，你们还有陈粮吃。”
LEV|25|23|“地不可以卖断，因为地是我的；你们在我面前是客旅，是寄居的。
LEV|25|24|在你们所得为业的全地，要准许人有权将地赎回。
LEV|25|25|“你的弟兄若渐渐贫穷，卖了他的一些产业，他的至亲就要来把弟兄所卖的赎回。
LEV|25|26|若没有人能为他赎回，他的手头渐渐宽裕，能够赎回，
LEV|25|27|就要计算卖后的年数，把剩余年数的价钱归还给那买主，他的地业便归还自己。
LEV|25|28|若他手头的财力不够赎回，所卖的地就要留在买主的手里，直到禧年。到了禧年，地业要归还卖主。
LEV|25|29|“人若卖城墙内的住宅，卖了以后，一整年内他有权赎回；这是他可以赎回的期限。
LEV|25|30|若他在一整年内不赎回，这有墙之城的房屋就确定永归买主，直到世世代代；在禧年也不必归还。
LEV|25|31|但周围无城墙之村庄的房屋，要看为乡下的田地，可以赎回；到了禧年就要归还。
LEV|25|32|至于 利未 人所得为业的城镇， 利未 人可以随时赎回他们城镇中的房屋。
LEV|25|33|在所得为业的城镇， 利未 人若卖了房屋，又不赎回，到了禧年仍要归还原主，因为 利未 人城镇的房屋是他们在 以色列 人中的产业。
LEV|25|34|但是 利未 人各城郊外之地是不可卖的，因为这是他们永远的产业。”
LEV|25|35|“你的弟兄在你那里若渐渐贫穷，手头缺乏，你就要帮补他，使他与你一同生活，像外人和寄居的一样。
LEV|25|36|不可向他取利息，也不可向他索取高利；要敬畏你的上帝，使你的弟兄与你一同生活。
LEV|25|37|你不可为了利息借钱给他，也不可为了高利而借粮。
LEV|25|38|我是耶和华－你们的上帝，曾领你们从 埃及 地出来，为要把 迦南 地赐给你们，要作你们的上帝。
LEV|25|39|“你的弟兄在你那里若渐渐贫穷，将自己卖给你，你不可叫他像奴仆服事你。
LEV|25|40|他在你那里要像雇工和寄居的，服事你直到禧年。
LEV|25|41|他和他儿女要离开你，一同出去，归回自己的家，回到他祖宗的地业去。
LEV|25|42|因为他们是我的仆人，是我从 埃及 地领出来的。他们不可被卖为奴仆。
LEV|25|43|不可苛刻管辖他，只要敬畏你的上帝。
LEV|25|44|至于你所要的奴仆和使女，可以来自你们四围的列国，你们可以从他们中买奴仆和使女。
LEV|25|45|那些寄居在你们中间的外人和他们的家属，就是在你们地上所生的，你们可以从其中买人；他们要作你们的产业。
LEV|25|46|你们可以把他们遗留给你们后代的子孙，作为永远继承的产业；你们可以使他们作奴仆。至于你们的弟兄 以色列 人，你们彼此不可苛刻管辖。
LEV|25|47|“住在你那里的外人或寄居的，若手头渐渐宽裕，你的弟兄却渐渐贫穷，将自己卖给那外人或寄居的，或外人家族的一支，
LEV|25|48|卖了以后，有权把自己赎回。他弟兄中的一位可以把他赎回。
LEV|25|49|他的叔伯或叔伯的儿子可以赎他。他家族中的骨肉之亲也可以赎他。他自己若手头渐渐宽裕，也可以赎回自己。
LEV|25|50|他要跟买主计算，从卖自己的那年起，算到禧年；所卖的价钱要按照年数计算，就是雇工跟买主在一起的日子。
LEV|25|51|若剩余的年数多，就要按着年数从买价中偿还他的赎价。
LEV|25|52|若到禧年只剩下几年，就要按着年数跟买主计算，偿还他的赎价。
LEV|25|53|他和买主同住，要像按年雇用的工人，买主不可苛刻管辖他。
LEV|25|54|他若不这样被赎，到了禧年，仍要和他的儿女一同出去。
LEV|25|55|因为 以色列 人都是我的仆人，他们是我的仆人，是我领他们从 埃及 地出来的。我是耶和华－你们的上帝。”
LEV|26|1|“你们不可为自己造虚无的神明，不可竖立雕刻的偶像或柱像，也不可在你们的地上安放石像，向它跪拜，因为我是耶和华－你们的上帝。
LEV|26|2|你们要谨守我的安息日，敬畏我的圣所。我是耶和华。
LEV|26|3|“你们若遵行我的律例，谨守我的诫命，实行它们，
LEV|26|4|我必按时降雨给你们，使地长出农作物，田野的树结出果实。
LEV|26|5|你们打谷物要打到摘葡萄的时候，摘葡萄要摘到播种的时候。你们要吃粮食得饱足，在你们的地上安然居住。
LEV|26|6|我要赐平安在地上；你们躺卧，无人惊吓。我要使你们地上的恶兽消灭，刀剑必不穿越你们的地。
LEV|26|7|你们要追赶仇敌，他们必倒在你们刀下。
LEV|26|8|你们五个人要追赶一百人，一百人要追赶一万人；仇敌必在你们面前倒在刀下。
LEV|26|9|我要眷顾你们，使你们生养众多，也要与你们坚立我的约。
LEV|26|10|你们要吃储存的陈粮，又要为新粮清理陈粮。
LEV|26|11|我要在你们中间立我的帐幕，我的心也不厌恶你们。
LEV|26|12|我要行走在你们中间，作你们的上帝，你们要作我的子民。
LEV|26|13|我是耶和华－你们的上帝，曾将你们从 埃及 地领出来，使你们不再作 埃及 人的奴仆；我曾折断你们所负的轭，使你们挺身前行。”
LEV|26|14|“你们若不听从我，不遵行我这一切的诫命，
LEV|26|15|厌弃我的律例，心中厌恶我的典章，不遵行我一切的诫命，背弃了我的约，
LEV|26|16|我就要这样对待你们：我必使惊惶临到你们，使你们患痨病，害热病，以致眼睛失明，身体衰弱。你们要白白撒种，因为仇敌要吃尽你们所种的。
LEV|26|17|我要向你们变脸，使你们败在仇敌的面前。恨恶你们的必管辖你们；无人追赶，你们却要逃跑。
LEV|26|18|如果这样，你们还不听从我，我就要因你们的罪，加重七倍惩罚你们。
LEV|26|19|我必粉碎你们因势力而有的骄傲，又要使你们的天坚如铁，地硬如铜。
LEV|26|20|你们劳力却白费，因为你们的地没有出产，地上的树也不结果实。
LEV|26|21|“你们行事若与我作对，不肯听从我，我就要因你们的罪，加重七倍灾祸击打你们。
LEV|26|22|我要打发野地的走兽到你们中间，夺去你们的儿女，吞灭你们的牲畜，使你们人数减少，道路荒凉。
LEV|26|23|“如果这样，你们还不接受管教归向我，行事与我作对，
LEV|26|24|我就要行事与你们作对，因你们的罪，加重七倍击打你们。
LEV|26|25|我要使刀剑临到你们，报复你们的背约。你们若被赶入城中，我要降瘟疫在你们中间，把你们交在仇敌手中。
LEV|26|26|我要断绝你们粮食的供应 ，使十个女人用一个烤炉给你们烤饼，按配给的定量秤给你们。你们要吃，却吃不饱。
LEV|26|27|“如果这样，你们还不听从我，行事与我作对，
LEV|26|28|我就要向你们发烈怒，行事与你们作对，因你们的罪，加重七倍惩罚你们。
LEV|26|29|你们要吃你们儿子的肉，也要吃你们女儿的肉。
LEV|26|30|我要摧毁你们的丘坛，砍掉你们的香坛，把你们的尸首扔在你们偶像的残骸上。我的心也必厌恶你们，
LEV|26|31|使你们的城镇变成废墟，你们的众圣所变荒凉，我也不闻你们芬芳的香气。
LEV|26|32|我要使这地变荒凉，甚至占领这地的敌人都惊讶。
LEV|26|33|我要把你们驱散到列国中，也要拔刀追赶你们。你们的地要成为荒凉，你们的城镇要变成废墟。
LEV|26|34|“当你们在敌人之地的时候，你们的地要在一切荒凉的日子重享安息；在那时候，地要休息，重享安息。
LEV|26|35|地在一切荒凉的日子都要安息，这是你们住在其上的时候所不能得的安息。
LEV|26|36|至于你们幸存的人，我要使他们在敌人之地心中惊慌，甚至风吹落叶的声音也把他们吓跑。他们要逃避，像人逃避刀剑，虽无人追赶，却要跌倒。
LEV|26|37|虽然无人追赶，他们却要彼此绊倒，像逃避刀剑一样。你们在仇敌面前必站立不住。
LEV|26|38|你们要在列国中灭亡，敌人之地要吞灭你们，
LEV|26|39|你们幸存的人必因自己的罪孽在敌人之地衰残，也要因祖先的罪孽衰残。
LEV|26|40|“他们要承认自己的罪孽和祖先的罪孽，就是背叛我，行事与我作对的过犯。
LEV|26|41|我也行事与他们作对，把他们遣送到敌人之地。那时，他们未受割礼的心若肯谦卑，也服了罪孽的惩罚，
LEV|26|42|我就要记念我与 雅各 的约，记念我与 以撒 的约，与 亚伯拉罕 的约；我也要记念这地。
LEV|26|43|地被他们离弃，因他们不在而荒凉的时候，就要重享安息。他们服了罪孽的惩罚，因为他们厌弃我的典章，心中厌恶我的律例。
LEV|26|44|虽然如此，当他们在敌人之地时，我却不厌弃他们，不厌恶他们，将他们全然灭绝，也不背弃我与他们的约，因为我是耶和华－他们的上帝。
LEV|26|45|我要为他们的缘故记念我与他们祖先的约；我在列国眼前曾把他们的祖先从 埃及 地领出来，为要作他们的上帝。我是耶和华。”
LEV|26|46|这些律例、典章和法度是耶和华在 西奈山 上藉着 摩西 与 以色列 人立的。
LEV|27|1|耶和华吩咐 摩西 说：
LEV|27|2|“你要吩咐 以色列 人，对他们说：人向耶和华许特别的愿，要按照你所估一个人的价钱。
LEV|27|3|你所估的是：二十岁到六十岁男的，按照圣所的舍客勒，估价是五十舍客勒银子。
LEV|27|4|若是女的，估价是三十舍客勒。
LEV|27|5|五岁到二十岁男的，估价是二十舍客勒，女的十舍客勒。
LEV|27|6|一个月到五岁男的，估价是五舍客勒，女的三舍客勒。
LEV|27|7|六十岁以上男的，估价是十五舍客勒，女的十舍客勒。
LEV|27|8|他若贫穷，不能按照你的估价，就要把他带到祭司面前，让祭司为他估价；祭司要按许愿者手头财力所及估价。
LEV|27|9|“许愿要献给耶和华的供物若是牲畜，凡这类献给耶和华的都要成为圣。
LEV|27|10|不可更换，也不可用另一只取代，无论是好的换坏的，或是坏的换好的，都不可。若一定要以牲畜取代牲畜，所许的与所取代的都要成为圣。
LEV|27|11|若牲畜不洁净，不可献给耶和华为供物，就要把牲畜带到祭司面前。
LEV|27|12|祭司要估价；牲畜是好是坏，祭司怎样估定，就是你的估价。
LEV|27|13|许愿者若一定要把它赎回，就要在你的估价上加五分之一。
LEV|27|14|“人将房屋分别为圣，归给耶和华为圣，祭司就要估价。房屋是好是坏，祭司怎样估定，就要以他的估价为准。
LEV|27|15|将房屋分别为圣的人，若要赎回房屋，必须付你所估定的价钱，再加上五分之一，房屋才可以归还给他。
LEV|27|16|“人若将所继承的一块田地分别为圣，归给耶和华，就要按照这地撒种多少来估价；能撒一贺梅珥大麦种子的，是五十舍客勒银子。
LEV|27|17|他若从禧年起将地分别为圣，就要以你的估价为准。
LEV|27|18|倘若他在禧年以后将地分别为圣，祭司就要按照从那时到下一个禧年所剩的年数推算，从你的估价中减掉。
LEV|27|19|将地分别为圣的人若要把地赎回，必须付你所估定的价钱，再加上五分之一，地才可以归还给他。
LEV|27|20|他若不赎回那地，或是将地卖给别人，就不能再赎了。
LEV|27|21|到了禧年，那田地要从买主手中退还，归耶和华为圣，和永献的地一样，要归祭司为业。
LEV|27|22|若分别为圣归耶和华的田地不是继承的，而是买来的，
LEV|27|23|祭司就要依照你的估价，推算到禧年。当天，这人要将你所估的归给耶和华为圣。
LEV|27|24|到了禧年，那田地要退还给卖主，就是继承那地的原主。
LEV|27|25|凡你所估的价钱都要按照圣所的舍客勒：二十季拉是一舍客勒。
LEV|27|26|“头生的，就是牲畜中头生属耶和华的，人不可再将它分别为圣，无论是牛是羊都是耶和华的。
LEV|27|27|头生的牲畜若是不洁净的，就要按照所估定的价钱，再加上五分之一，把它赎回。若不赎回，就要按照你的估价把它卖了。
LEV|27|28|“但一切永献作当灭的，就是人从他所有永献给耶和华作当灭的，无论是人，是牲畜，是他继承的田地，都不可卖，也不可赎。凡永献作当灭的都归耶和华为至圣。
LEV|27|29|凡从人中永献作当灭的都不可赎，必被处死。
LEV|27|30|“地上所有的，无论是地上的种子，是树上的果子，十分之一是耶和华的，是归耶和华为圣的。
LEV|27|31|人若要赎回这十分之一，就要另加五分之一。
LEV|27|32|凡牛群羊群中的十分之一，就是一切从牧人杖下经过的，每第十只要归耶和华为圣。
LEV|27|33|不可追究是好是坏，也不可取代；若一定要取代，所取代的和本来当献的牲畜都要成为圣，不可赎回。”
LEV|27|34|这些是耶和华在 西奈山 为 以色列 人所吩咐 摩西 的命令。
