PROV|1|1|The proverbs of Solomon the son of David, king of Israel;
PROV|1|2|To know wisdom and instruction; to perceive the words of understanding;
PROV|1|3|To receive the instruction of wisdom, justice, and judgment, and equity;
PROV|1|4|To give subtilty to the simple, to the young man knowledge and discretion.
PROV|1|5|A wise man will hear, and will increase learning; and a man of understanding shall attain unto wise counsels:
PROV|1|6|To understand a proverb, and the interpretation; the words of the wise, and their dark sayings.
PROV|1|7|The fear of the LORD is the beginning of knowledge: but fools despise wisdom and instruction.
PROV|1|8|My son, hear the instruction of thy father, and forsake not the law of thy mother:
PROV|1|9|For they shall be an ornament of grace unto thy head, and chains about thy neck.
PROV|1|10|My son, if sinners entice thee, consent thou not.
PROV|1|11|If they say, Come with us, let us lay wait for blood, let us lurk privily for the innocent without cause:
PROV|1|12|Let us swallow them up alive as the grave; and whole, as those that go down into the pit:
PROV|1|13|We shall find all precious substance, we shall fill our houses with spoil:
PROV|1|14|Cast in thy lot among us; let us all have one purse:
PROV|1|15|My son, walk not thou in the way with them; refrain thy foot from their path:
PROV|1|16|For their feet run to evil, and make haste to shed blood.
PROV|1|17|Surely in vain the net is spread in the sight of any bird.
PROV|1|18|And they lay wait for their own blood; they lurk privily for their own lives.
PROV|1|19|So are the ways of every one that is greedy of gain; which taketh away the life of the owners thereof.
PROV|1|20|Wisdom crieth without; she uttereth her voice in the streets:
PROV|1|21|She crieth in the chief place of concourse, in the openings of the gates: in the city she uttereth her words, saying,
PROV|1|22|How long, ye simple ones, will ye love simplicity? and the scorners delight in their scorning, and fools hate knowledge?
PROV|1|23|Turn you at my reproof: behold, I will pour out my spirit unto you, I will make known my words unto you.
PROV|1|24|Because I have called, and ye refused; I have stretched out my hand, and no man regarded;
PROV|1|25|But ye have set at nought all my counsel, and would none of my reproof:
PROV|1|26|I also will laugh at your calamity; I will mock when your fear cometh;
PROV|1|27|When your fear cometh as desolation, and your destruction cometh as a whirlwind; when distress and anguish cometh upon you.
PROV|1|28|Then shall they call upon me, but I will not answer; they shall seek me early, but they shall not find me:
PROV|1|29|For that they hated knowledge, and did not choose the fear of the LORD:
PROV|1|30|They would none of my counsel: they despised all my reproof.
PROV|1|31|Therefore shall they eat of the fruit of their own way, and be filled with their own devices.
PROV|1|32|For the turning away of the simple shall slay them, and the prosperity of fools shall destroy them.
PROV|1|33|But whoso hearkeneth unto me shall dwell safely, and shall be quiet from fear of evil.
PROV|2|1|My son, if thou wilt receive my words, and hide my commandments with thee;
PROV|2|2|So that thou incline thine ear unto wisdom, and apply thine heart to understanding;
PROV|2|3|Yea, if thou criest after knowledge, and liftest up thy voice for understanding;
PROV|2|4|If thou seekest her as silver, and searchest for her as for hid treasures;
PROV|2|5|Then shalt thou understand the fear of the LORD, and find the knowledge of God.
PROV|2|6|For the LORD giveth wisdom: out of his mouth cometh knowledge and understanding.
PROV|2|7|He layeth up sound wisdom for the righteous: he is a buckler to them that walk uprightly.
PROV|2|8|He keepeth the paths of judgment, and preserveth the way of his saints.
PROV|2|9|Then shalt thou understand righteousness, and judgment, and equity; yea, every good path.
PROV|2|10|When wisdom entereth into thine heart, and knowledge is pleasant unto thy soul;
PROV|2|11|Discretion shall preserve thee, understanding shall keep thee:
PROV|2|12|To deliver thee from the way of the evil man, from the man that speaketh froward things;
PROV|2|13|Who leave the paths of uprightness, to walk in the ways of darkness;
PROV|2|14|Who rejoice to do evil, and delight in the frowardness of the wicked;
PROV|2|15|Whose ways are crooked, and they froward in their paths:
PROV|2|16|To deliver thee from the strange woman, even from the stranger which flattereth with her words;
PROV|2|17|Which forsaketh the guide of her youth, and forgetteth the covenant of her God.
PROV|2|18|For her house inclineth unto death, and her paths unto the dead.
PROV|2|19|None that go unto her return again, neither take they hold of the paths of life.
PROV|2|20|That thou mayest walk in the way of good men, and keep the paths of the righteous.
PROV|2|21|For the upright shall dwell in the land, and the perfect shall remain in it.
PROV|2|22|But the wicked shall be cut off from the earth, and the transgressors shall be rooted out of it.
PROV|3|1|My son, forget not my law; but let thine heart keep my commandments:
PROV|3|2|For length of days, and long life, and peace, shall they add to thee.
PROV|3|3|Let not mercy and truth forsake thee: bind them about thy neck; write them upon the table of thine heart:
PROV|3|4|So shalt thou find favour and good understanding in the sight of God and man.
PROV|3|5|Trust in the LORD with all thine heart; and lean not unto thine own understanding.
PROV|3|6|In all thy ways acknowledge him, and he shall direct thy paths.
PROV|3|7|Be not wise in thine own eyes: fear the LORD, and depart from evil.
PROV|3|8|It shall be health to thy navel, and marrow to thy bones.
PROV|3|9|Honour the LORD with thy substance, and with the firstfruits of all thine increase:
PROV|3|10|So shall thy barns be filled with plenty, and thy presses shall burst out with new wine.
PROV|3|11|My son, despise not the chastening of the LORD; neither be weary of his correction:
PROV|3|12|For whom the LORD loveth he correcteth; even as a father the son in whom he delighteth.
PROV|3|13|Happy is the man that findeth wisdom, and the man that getteth understanding.
PROV|3|14|For the merchandise of it is better than the merchandise of silver, and the gain thereof than fine gold.
PROV|3|15|She is more precious than rubies: and all the things thou canst desire are not to be compared unto her.
PROV|3|16|Length of days is in her right hand; and in her left hand riches and honour.
PROV|3|17|Her ways are ways of pleasantness, and all her paths are peace.
PROV|3|18|She is a tree of life to them that lay hold upon her: and happy is every one that retaineth her.
PROV|3|19|The LORD by wisdom hath founded the earth; by understanding hath he established the heavens.
PROV|3|20|By his knowledge the depths are broken up, and the clouds drop down the dew.
PROV|3|21|My son, let not them depart from thine eyes: keep sound wisdom and discretion:
PROV|3|22|So shall they be life unto thy soul, and grace to thy neck.
PROV|3|23|Then shalt thou walk in thy way safely, and thy foot shall not stumble.
PROV|3|24|When thou liest down, thou shalt not be afraid: yea, thou shalt lie down, and thy sleep shall be sweet.
PROV|3|25|Be not afraid of sudden fear, neither of the desolation of the wicked, when it cometh.
PROV|3|26|For the LORD shall be thy confidence, and shall keep thy foot from being taken.
PROV|3|27|Withhold not good from them to whom it is due, when it is in the power of thine hand to do it.
PROV|3|28|Say not unto thy neighbour, Go, and come again, and to morrow I will give; when thou hast it by thee.
PROV|3|29|Devise not evil against thy neighbour, seeing he dwelleth securely by thee.
PROV|3|30|Strive not with a man without cause, if he have done thee no harm.
PROV|3|31|Envy thou not the oppressor, and choose none of his ways.
PROV|3|32|For the froward is abomination to the LORD: but his secret is with the righteous.
PROV|3|33|The curse of the LORD is in the house of the wicked: but he blesseth the habitation of the just.
PROV|3|34|Surely he scorneth the scorners: but he giveth grace unto the lowly.
PROV|3|35|The wise shall inherit glory: but shame shall be the promotion of fools.
PROV|4|1|Hear, ye children, the instruction of a father, and attend to know understanding.
PROV|4|2|For I give you good doctrine, forsake ye not my law.
PROV|4|3|For I was my father's son, tender and only beloved in the sight of my mother.
PROV|4|4|He taught me also, and said unto me, Let thine heart retain my words: keep my commandments, and live.
PROV|4|5|Get wisdom, get understanding: forget it not; neither decline from the words of my mouth.
PROV|4|6|Forsake her not, and she shall preserve thee: love her, and she shall keep thee.
PROV|4|7|Wisdom is the principal thing; therefore get wisdom: and with all thy getting get understanding.
PROV|4|8|Exalt her, and she shall promote thee: she shall bring thee to honour, when thou dost embrace her.
PROV|4|9|She shall give to thine head an ornament of grace: a crown of glory shall she deliver to thee.
PROV|4|10|Hear, O my son, and receive my sayings; and the years of thy life shall be many.
PROV|4|11|I have taught thee in the way of wisdom; I have led thee in right paths.
PROV|4|12|When thou goest, thy steps shall not be straitened; and when thou runnest, thou shalt not stumble.
PROV|4|13|Take fast hold of instruction; let her not go: keep her; for she is thy life.
PROV|4|14|Enter not into the path of the wicked, and go not in the way of evil men.
PROV|4|15|Avoid it, pass not by it, turn from it, and pass away.
PROV|4|16|For they sleep not, except they have done mischief; and their sleep is taken away, unless they cause some to fall.
PROV|4|17|For they eat the bread of wickedness, and drink the wine of violence.
PROV|4|18|But the path of the just is as the shining light, that shineth more and more unto the perfect day.
PROV|4|19|The way of the wicked is as darkness: they know not at what they stumble.
PROV|4|20|My son, attend to my words; incline thine ear unto my sayings.
PROV|4|21|Let them not depart from thine eyes; keep them in the midst of thine heart.
PROV|4|22|For they are life unto those that find them, and health to all their flesh.
PROV|4|23|Keep thy heart with all diligence; for out of it are the issues of life.
PROV|4|24|Put away from thee a froward mouth, and perverse lips put far from thee.
PROV|4|25|Let thine eyes look right on, and let thine eyelids look straight before thee.
PROV|4|26|Ponder the path of thy feet, and let all thy ways be established.
PROV|4|27|Turn not to the right hand nor to the left: remove thy foot from evil.
PROV|5|1|My son, attend unto my wisdom, and bow thine ear to my understanding:
PROV|5|2|That thou mayest regard discretion, and that thy lips may keep knowledge.
PROV|5|3|For the lips of a strange woman drop as an honeycomb, and her mouth is smoother than oil:
PROV|5|4|But her end is bitter as wormwood, sharp as a two-edged sword.
PROV|5|5|Her feet go down to death; her steps take hold on hell.
PROV|5|6|Lest thou shouldest ponder the path of life, her ways are moveable, that thou canst not know them.
PROV|5|7|Hear me now therefore, O ye children, and depart not from the words of my mouth.
PROV|5|8|Remove thy way far from her, and come not nigh the door of her house:
PROV|5|9|Lest thou give thine honour unto others, and thy years unto the cruel:
PROV|5|10|Lest strangers be filled with thy wealth; and thy labours be in the house of a stranger;
PROV|5|11|And thou mourn at the last, when thy flesh and thy body are consumed,
PROV|5|12|And say, How have I hated instruction, and my heart despised reproof;
PROV|5|13|And have not obeyed the voice of my teachers, nor inclined mine ear to them that instructed me!
PROV|5|14|I was almost in all evil in the midst of the congregation and assembly.
PROV|5|15|Drink waters out of thine own cistern, and running waters out of thine own well.
PROV|5|16|Let thy fountains be dispersed abroad, and rivers of waters in the streets.
PROV|5|17|Let them be only thine own, and not strangers' with thee.
PROV|5|18|Let thy fountain be blessed: and rejoice with the wife of thy youth.
PROV|5|19|Let her be as the loving hind and pleasant roe; let her breasts satisfy thee at all times; and be thou ravished always with her love.
PROV|5|20|And why wilt thou, my son, be ravished with a strange woman, and embrace the bosom of a stranger?
PROV|5|21|For the ways of man are before the eyes of the LORD, and he pondereth all his goings.
PROV|5|22|His own iniquities shall take the wicked himself, and he shall be holden with the cords of his sins.
PROV|5|23|He shall die without instruction; and in the greatness of his folly he shall go astray.
PROV|6|1|My son, if thou be surety for thy friend, if thou hast stricken thy hand with a stranger,
PROV|6|2|Thou art snared with the words of thy mouth, thou art taken with the words of thy mouth.
PROV|6|3|Do this now, my son, and deliver thyself, when thou art come into the hand of thy friend; go, humble thyself, and make sure thy friend.
PROV|6|4|Give not sleep to thine eyes, nor slumber to thine eyelids.
PROV|6|5|Deliver thyself as a roe from the hand of the hunter, and as a bird from the hand of the fowler.
PROV|6|6|Go to the ant, thou sluggard; consider her ways, and be wise:
PROV|6|7|Which having no guide, overseer, or ruler,
PROV|6|8|Provideth her meat in the summer, and gathereth her food in the harvest.
PROV|6|9|How long wilt thou sleep, O sluggard? when wilt thou arise out of thy sleep?
PROV|6|10|Yet a little sleep, a little slumber, a little folding of the hands to sleep:
PROV|6|11|So shall thy poverty come as one that travelleth, and thy want as an armed man.
PROV|6|12|A naughty person, a wicked man, walketh with a froward mouth.
PROV|6|13|He winketh with his eyes, he speaketh with his feet, he teacheth with his fingers;
PROV|6|14|Frowardness is in his heart, he deviseth mischief continually; he soweth discord.
PROV|6|15|Therefore shall his calamity come suddenly; suddenly shall he be broken without remedy.
PROV|6|16|These six things doth the LORD hate: yea, seven are an abomination unto him:
PROV|6|17|A proud look, a lying tongue, and hands that shed innocent blood,
PROV|6|18|An heart that deviseth wicked imaginations, feet that be swift in running to mischief,
PROV|6|19|A false witness that speaketh lies, and he that soweth discord among brethren.
PROV|6|20|My son, keep thy father's commandment, and forsake not the law of thy mother:
PROV|6|21|Bind them continually upon thine heart, and tie them about thy neck.
PROV|6|22|When thou goest, it shall lead thee; when thou sleepest, it shall keep thee; and when thou awakest, it shall talk with thee.
PROV|6|23|For the commandment is a lamp; and the law is light; and reproofs of instruction are the way of life:
PROV|6|24|To keep thee from the evil woman, from the flattery of the tongue of a strange woman.
PROV|6|25|Lust not after her beauty in thine heart; neither let her take thee with her eyelids.
PROV|6|26|For by means of a whorish woman a man is brought to a piece of bread: and the adultress will hunt for the precious life.
PROV|6|27|Can a man take fire in his bosom, and his clothes not be burned?
PROV|6|28|Can one go upon hot coals, and his feet not be burned?
PROV|6|29|So he that goeth in to his neighbour's wife; whosoever toucheth her shall not be innocent.
PROV|6|30|Men do not despise a thief, if he steal to satisfy his soul when he is hungry;
PROV|6|31|But if he be found, he shall restore sevenfold; he shall give all the substance of his house.
PROV|6|32|But whoso committeth adultery with a woman lacketh understanding: he that doeth it destroyeth his own soul.
PROV|6|33|A wound and dishonour shall he get; and his reproach shall not be wiped away.
PROV|6|34|For jealousy is the rage of a man: therefore he will not spare in the day of vengeance.
PROV|6|35|He will not regard any ransom; neither will he rest content, though thou givest many gifts.
PROV|7|1|My son, keep my words, and lay up my commandments with thee.
PROV|7|2|Keep my commandments, and live; and my law as the apple of thine eye.
PROV|7|3|Bind them upon thy fingers, write them upon the table of thine heart.
PROV|7|4|Say unto wisdom, Thou art my sister; and call understanding thy kinswoman:
PROV|7|5|That they may keep thee from the strange woman, from the stranger which flattereth with her words.
PROV|7|6|For at the window of my house I looked through my casement,
PROV|7|7|And beheld among the simple ones, I discerned among the youths, a young man void of understanding,
PROV|7|8|Passing through the street near her corner; and he went the way to her house,
PROV|7|9|In the twilight, in the evening, in the black and dark night:
PROV|7|10|And, behold, there met him a woman with the attire of an harlot, and subtil of heart.
PROV|7|11|(She is loud and stubborn; her feet abide not in her house:
PROV|7|12|Now is she without, now in the streets, and lieth in wait at every corner.)
PROV|7|13|So she caught him, and kissed him, and with an impudent face said unto him,
PROV|7|14|I have peace offerings with me; this day have I payed my vows.
PROV|7|15|Therefore came I forth to meet thee, diligently to seek thy face, and I have found thee.
PROV|7|16|I have decked my bed with coverings of tapestry, with carved works, with fine linen of Egypt.
PROV|7|17|I have perfumed my bed with myrrh, aloes, and cinnamon.
PROV|7|18|Come, let us take our fill of love until the morning: let us solace ourselves with loves.
PROV|7|19|For the goodman is not at home, he is gone a long journey:
PROV|7|20|He hath taken a bag of money with him, and will come home at the day appointed.
PROV|7|21|With her much fair speech she caused him to yield, with the flattering of her lips she forced him.
PROV|7|22|He goeth after her straightway, as an ox goeth to the slaughter, or as a fool to the correction of the stocks;
PROV|7|23|Till a dart strike through his liver; as a bird hasteth to the snare, and knoweth not that it is for his life.
PROV|7|24|Hearken unto me now therefore, O ye children, and attend to the words of my mouth.
PROV|7|25|Let not thine heart decline to her ways, go not astray in her paths.
PROV|7|26|For she hath cast down many wounded: yea, many strong men have been slain by her.
PROV|7|27|Her house is the way to hell, going down to the chambers of death.
PROV|8|1|Doth not wisdom cry? and understanding put forth her voice?
PROV|8|2|She standeth in the top of high places, by the way in the places of the paths.
PROV|8|3|She crieth at the gates, at the entry of the city, at the coming in at the doors.
PROV|8|4|Unto you, O men, I call; and my voice is to the sons of man.
PROV|8|5|O ye simple, understand wisdom: and, ye fools, be ye of an understanding heart.
PROV|8|6|Hear; for I will speak of excellent things; and the opening of my lips shall be right things.
PROV|8|7|For my mouth shall speak truth; and wickedness is an abomination to my lips.
PROV|8|8|All the words of my mouth are in righteousness; there is nothing froward or perverse in them.
PROV|8|9|They are all plain to him that understandeth, and right to them that find knowledge.
PROV|8|10|Receive my instruction, and not silver; and knowledge rather than choice gold.
PROV|8|11|For wisdom is better than rubies; and all the things that may be desired are not to be compared to it.
PROV|8|12|I wisdom dwell with prudence, and find out knowledge of witty inventions.
PROV|8|13|The fear of the LORD is to hate evil: pride, and arrogancy, and the evil way, and the froward mouth, do I hate.
PROV|8|14|Counsel is mine, and sound wisdom: I am understanding; I have strength.
PROV|8|15|By me kings reign, and princes decree justice.
PROV|8|16|By me princes rule, and nobles, even all the judges of the earth.
PROV|8|17|I love them that love me; and those that seek me early shall find me.
PROV|8|18|Riches and honour are with me; yea, durable riches and righteousness.
PROV|8|19|My fruit is better than gold, yea, than fine gold; and my revenue than choice silver.
PROV|8|20|I lead in the way of righteousness, in the midst of the paths of judgment:
PROV|8|21|That I may cause those that love me to inherit substance; and I will fill their treasures.
PROV|8|22|The LORD possessed me in the beginning of his way, before his works of old.
PROV|8|23|I was set up from everlasting, from the beginning, or ever the earth was.
PROV|8|24|When there were no depths, I was brought forth; when there were no fountains abounding with water.
PROV|8|25|Before the mountains were settled, before the hills was I brought forth:
PROV|8|26|While as yet he had not made the earth, nor the fields, nor the highest part of the dust of the world.
PROV|8|27|When he prepared the heavens, I was there: when he set a compass upon the face of the depth:
PROV|8|28|When he established the clouds above: when he strengthened the fountains of the deep:
PROV|8|29|When he gave to the sea his decree, that the waters should not pass his commandment: when he appointed the foundations of the earth:
PROV|8|30|Then I was by him, as one brought up with him: and I was daily his delight, rejoicing always before him;
PROV|8|31|Rejoicing in the habitable part of his earth; and my delights were with the sons of men.
PROV|8|32|Now therefore hearken unto me, O ye children: for blessed are they that keep my ways.
PROV|8|33|Hear instruction, and be wise, and refuse it not.
PROV|8|34|Blessed is the man that heareth me, watching daily at my gates, waiting at the posts of my doors.
PROV|8|35|For whoso findeth me findeth life, and shall obtain favour of the LORD.
PROV|8|36|But he that sinneth against me wrongeth his own soul: all they that hate me love death.
PROV|9|1|Wisdom hath builded her house, she hath hewn out her seven pillars:
PROV|9|2|She hath killed her beasts; she hath mingled her wine; she hath also furnished her table.
PROV|9|3|She hath sent forth her maidens: she crieth upon the highest places of the city,
PROV|9|4|Whoso is simple, let him turn in hither: as for him that wanteth understanding, she saith to him,
PROV|9|5|Come, eat of my bread, and drink of the wine which I have mingled.
PROV|9|6|Forsake the foolish, and live; and go in the way of understanding.
PROV|9|7|He that reproveth a scorner getteth to himself shame: and he that rebuketh a wicked man getteth himself a blot.
PROV|9|8|Reprove not a scorner, lest he hate thee: rebuke a wise man, and he will love thee.
PROV|9|9|Give instruction to a wise man, and he will be yet wiser: teach a just man, and he will increase in learning.
PROV|9|10|The fear of the LORD is the beginning of wisdom: and the knowledge of the holy is understanding.
PROV|9|11|For by me thy days shall be multiplied, and the years of thy life shall be increased.
PROV|9|12|If thou be wise, thou shalt be wise for thyself: but if thou scornest, thou alone shalt bear it.
PROV|9|13|A foolish woman is clamorous: she is simple, and knoweth nothing.
PROV|9|14|For she sitteth at the door of her house, on a seat in the high places of the city,
PROV|9|15|To call passengers who go right on their ways:
PROV|9|16|Whoso is simple, let him turn in hither: and as for him that wanteth understanding, she saith to him,
PROV|9|17|Stolen waters are sweet, and bread eaten in secret is pleasant.
PROV|9|18|But he knoweth not that the dead are there; and that her guests are in the depths of hell.
PROV|10|1|The proverbs of Solomon. A wise son maketh a glad father: but a foolish son is the heaviness of his mother.
PROV|10|2|Treasures of wickedness profit nothing: but righteousness delivereth from death.
PROV|10|3|The LORD will not suffer the soul of the righteous to famish: but he casteth away the substance of the wicked.
PROV|10|4|He becometh poor that dealeth with a slack hand: but the hand of the diligent maketh rich.
PROV|10|5|He that gathereth in summer is a wise son: but he that sleepeth in harvest is a son that causeth shame.
PROV|10|6|Blessings are upon the head of the just: but violence covereth the mouth of the wicked.
PROV|10|7|The memory of the just is blessed: but the name of the wicked shall rot.
PROV|10|8|The wise in heart will receive commandments: but a prating fool shall fall.
PROV|10|9|He that walketh uprightly walketh surely: but he that perverteth his ways shall be known.
PROV|10|10|He that winketh with the eye causeth sorrow: but a prating fool shall fall.
PROV|10|11|The mouth of a righteous man is a well of life: but violence covereth the mouth of the wicked.
PROV|10|12|Hatred stirreth up strifes: but love covereth all sins.
PROV|10|13|In the lips of him that hath understanding wisdom is found: but a rod is for the back of him that is void of understanding.
PROV|10|14|Wise men lay up knowledge: but the mouth of the foolish is near destruction.
PROV|10|15|The rich man's wealth is his strong city: the destruction of the poor is their poverty.
PROV|10|16|The labour of the righteous tendeth to life: the fruit of the wicked to sin.
PROV|10|17|He is in the way of life that keepeth instruction: but he that refuseth reproof erreth.
PROV|10|18|He that hideth hatred with lying lips, and he that uttereth a slander, is a fool.
PROV|10|19|In the multitude of words there wanteth not sin: but he that refraineth his lips is wise.
PROV|10|20|The tongue of the just is as choice silver: the heart of the wicked is little worth.
PROV|10|21|The lips of the righteous feed many: but fools die for want of wisdom.
PROV|10|22|The blessing of the LORD, it maketh rich, and he addeth no sorrow with it.
PROV|10|23|It is as sport to a fool to do mischief: but a man of understanding hath wisdom.
PROV|10|24|The fear of the wicked, it shall come upon him: but the desire of the righteous shall be granted.
PROV|10|25|As the whirlwind passeth, so is the wicked no more: but the righteous is an everlasting foundation.
PROV|10|26|As vinegar to the teeth, and as smoke to the eyes, so is the sluggard to them that send him.
PROV|10|27|The fear of the LORD prolongeth days: but the years of the wicked shall be shortened.
PROV|10|28|The hope of the righteous shall be gladness: but the expectation of the wicked shall perish.
PROV|10|29|The way of the LORD is strength to the upright: but destruction shall be to the workers of iniquity.
PROV|10|30|The righteous shall never be removed: but the wicked shall not inhabit the earth.
PROV|10|31|The mouth of the just bringeth forth wisdom: but the froward tongue shall be cut out.
PROV|10|32|The lips of the righteous know what is acceptable: but the mouth of the wicked speaketh frowardness.
PROV|11|1|A false balance is abomination to the LORD: but a just weight is his delight.
PROV|11|2|When pride cometh, then cometh shame: but with the lowly is wisdom.
PROV|11|3|The integrity of the upright shall guide them: but the perverseness of transgressors shall destroy them.
PROV|11|4|Riches profit not in the day of wrath: but righteousness delivereth from death.
PROV|11|5|The righteousness of the perfect shall direct his way: but the wicked shall fall by his own wickedness.
PROV|11|6|The righteousness of the upright shall deliver them: but transgressors shall be taken in their own naughtiness.
PROV|11|7|When a wicked man dieth, his expectation shall perish: and the hope of unjust men perisheth.
PROV|11|8|The righteous is delivered out of trouble, and the wicked cometh in his stead.
PROV|11|9|An hypocrite with his mouth destroyeth his neighbour: but through knowledge shall the just be delivered.
PROV|11|10|When it goeth well with the righteous, the city rejoiceth: and when the wicked perish, there is shouting.
PROV|11|11|By the blessing of the upright the city is exalted: but it is overthrown by the mouth of the wicked.
PROV|11|12|He that is void of wisdom despiseth his neighbour: but a man of understanding holdeth his peace.
PROV|11|13|A talebearer revealeth secrets: but he that is of a faithful spirit concealeth the matter.
PROV|11|14|Where no counsel is, the people fall: but in the multitude of counsellors there is safety.
PROV|11|15|He that is surety for a stranger shall smart for it: and he that hateth suretiship is sure.
PROV|11|16|A gracious woman retaineth honour: and strong men retain riches.
PROV|11|17|The merciful man doeth good to his own soul: but he that is cruel troubleth his own flesh.
PROV|11|18|The wicked worketh a deceitful work: but to him that soweth righteousness shall be a sure reward.
PROV|11|19|As righteousness tendeth to life: so he that pursueth evil pursueth it to his own death.
PROV|11|20|They that are of a froward heart are abomination to the LORD: but such as are upright in their way are his delight.
PROV|11|21|Though hand join in hand, the wicked shall not be unpunished: but the seed of the righteous shall be delivered.
PROV|11|22|As a jewel of gold in a swine's snout, so is a fair woman which is without discretion.
PROV|11|23|The desire of the righteous is only good: but the expectation of the wicked is wrath.
PROV|11|24|There is that scattereth, and yet increaseth; and there is that withholdeth more than is meet, but it tendeth to poverty.
PROV|11|25|The liberal soul shall be made fat: and he that watereth shall be watered also himself.
PROV|11|26|He that withholdeth corn, the people shall curse him: but blessing shall be upon the head of him that selleth it.
PROV|11|27|He that diligently seeketh good procureth favour: but he that seeketh mischief, it shall come unto him.
PROV|11|28|He that trusteth in his riches shall fall; but the righteous shall flourish as a branch.
PROV|11|29|He that troubleth his own house shall inherit the wind: and the fool shall be servant to the wise of heart.
PROV|11|30|The fruit of the righteous is a tree of life; and he that winneth souls is wise.
PROV|11|31|Behold, the righteous shall be recompensed in the earth: much more the wicked and the sinner.
PROV|12|1|Whoso loveth instruction loveth knowledge: but he that hateth reproof is brutish.
PROV|12|2|A good man obtaineth favour of the LORD: but a man of wicked devices will he condemn.
PROV|12|3|A man shall not be established by wickedness: but the root of the righteous shall not be moved.
PROV|12|4|A virtuous woman is a crown to her husband: but she that maketh ashamed is as rottenness in his bones.
PROV|12|5|The thoughts of the righteous are right: but the counsels of the wicked are deceit.
PROV|12|6|The words of the wicked are to lie in wait for blood: but the mouth of the upright shall deliver them.
PROV|12|7|The wicked are overthrown, and are not: but the house of the righteous shall stand.
PROV|12|8|A man shall be commended according to his wisdom: but he that is of a perverse heart shall be despised.
PROV|12|9|He that is despised, and hath a servant, is better than he that honoureth himself, and lacketh bread.
PROV|12|10|A righteous man regardeth the life of his beast: but the tender mercies of the wicked are cruel.
PROV|12|11|He that tilleth his land shall be satisfied with bread: but he that followeth vain persons is void of understanding.
PROV|12|12|The wicked desireth the net of evil men: but the root of the righteous yieldeth fruit.
PROV|12|13|The wicked is snared by the transgression of his lips: but the just shall come out of trouble.
PROV|12|14|A man shall be satisfied with good by the fruit of his mouth: and the recompence of a man's hands shall be rendered unto him.
PROV|12|15|The way of a fool is right in his own eyes: but he that hearkeneth unto counsel is wise.
PROV|12|16|A fool's wrath is presently known: but a prudent man covereth shame.
PROV|12|17|He that speaketh truth sheweth forth righteousness: but a false witness deceit.
PROV|12|18|There is that speaketh like the piercings of a sword: but the tongue of the wise is health.
PROV|12|19|The lip of truth shall be established for ever: but a lying tongue is but for a moment.
PROV|12|20|Deceit is in the heart of them that imagine evil: but to the counsellors of peace is joy.
PROV|12|21|There shall no evil happen to the just: but the wicked shall be filled with mischief.
PROV|12|22|Lying lips are abomination to the LORD: but they that deal truly are his delight.
PROV|12|23|A prudent man concealeth knowledge: but the heart of fools proclaimeth foolishness.
PROV|12|24|The hand of the diligent shall bear rule: but the slothful shall be under tribute.
PROV|12|25|Heaviness in the heart of man maketh it stoop: but a good word maketh it glad.
PROV|12|26|The righteous is more excellent than his neighbour: but the way of the wicked seduceth them.
PROV|12|27|The slothful man roasteth not that which he took in hunting: but the substance of a diligent man is precious.
PROV|12|28|In the way of righteousness is life: and in the pathway thereof there is no death.
PROV|13|1|A wise son heareth his father's instruction: but a scorner heareth not rebuke.
PROV|13|2|A man shall eat good by the fruit of his mouth: but the soul of the transgressors shall eat violence.
PROV|13|3|He that keepeth his mouth keepeth his life: but he that openeth wide his lips shall have destruction.
PROV|13|4|The soul of the sluggard desireth, and hath nothing: but the soul of the diligent shall be made fat.
PROV|13|5|A righteous man hateth lying: but a wicked man is loathsome, and cometh to shame.
PROV|13|6|Righteousness keepeth him that is upright in the way: but wickedness overthroweth the sinner.
PROV|13|7|There is that maketh himself rich, yet hath nothing: there is that maketh himself poor, yet hath great riches.
PROV|13|8|The ransom of a man's life are his riches: but the poor heareth not rebuke.
PROV|13|9|The light of the righteous rejoiceth: but the lamp of the wicked shall be put out.
PROV|13|10|Only by pride cometh contention: but with the well advised is wisdom.
PROV|13|11|Wealth gotten by vanity shall be diminished: but he that gathereth by labour shall increase.
PROV|13|12|Hope deferred maketh the heart sick: but when the desire cometh, it is a tree of life.
PROV|13|13|Whoso despiseth the word shall be destroyed: but he that feareth the commandment shall be rewarded.
PROV|13|14|The law of the wise is a fountain of life, to depart from the snares of death.
PROV|13|15|Good understanding giveth favour: but the way of transgressors is hard.
PROV|13|16|Every prudent man dealeth with knowledge: but a fool layeth open his folly.
PROV|13|17|A wicked messenger falleth into mischief: but a faithful ambassador is health.
PROV|13|18|Poverty and shame shall be to him that refuseth instruction: but he that regardeth reproof shall be honoured.
PROV|13|19|The desire accomplished is sweet to the soul: but it is abomination to fools to depart from evil.
PROV|13|20|He that walketh with wise men shall be wise: but a companion of fools shall be destroyed.
PROV|13|21|Evil pursueth sinners: but to the righteous good shall be repayed.
PROV|13|22|A good man leaveth an inheritance to his children's children: and the wealth of the sinner is laid up for the just.
PROV|13|23|Much food is in the tillage of the poor: but there is that is destroyed for want of judgment.
PROV|13|24|He that spareth his rod hateth his son: but he that loveth him chasteneth him betimes.
PROV|13|25|The righteous eateth to the satisfying of his soul: but the belly of the wicked shall want.
PROV|14|1|Every wise woman buildeth her house: but the foolish plucketh it down with her hands.
PROV|14|2|He that walketh in his uprightness feareth the LORD: but he that is perverse in his ways despiseth him.
PROV|14|3|In the mouth of the foolish is a rod of pride: but the lips of the wise shall preserve them.
PROV|14|4|Where no oxen are, the crib is clean: but much increase is by the strength of the ox.
PROV|14|5|A faithful witness will not lie: but a false witness will utter lies.
PROV|14|6|A scorner seeketh wisdom, and findeth it not: but knowledge is easy unto him that understandeth.
PROV|14|7|Go from the presence of a foolish man, when thou perceivest not in him the lips of knowledge.
PROV|14|8|The wisdom of the prudent is to understand his way: but the folly of fools is deceit.
PROV|14|9|Fools make a mock at sin: but among the righteous there is favour.
PROV|14|10|The heart knoweth his own bitterness; and a stranger doth not intermeddle with his joy.
PROV|14|11|The house of the wicked shall be overthrown: but the tabernacle of the upright shall flourish.
PROV|14|12|There is a way which seemeth right unto a man, but the end thereof are the ways of death.
PROV|14|13|Even in laughter the heart is sorrowful; and the end of that mirth is heaviness.
PROV|14|14|The backslider in heart shall be filled with his own ways: and a good man shall be satisfied from himself.
PROV|14|15|The simple believeth every word: but the prudent man looketh well to his going.
PROV|14|16|A wise man feareth, and departeth from evil: but the fool rageth, and is confident.
PROV|14|17|He that is soon angry dealeth foolishly: and a man of wicked devices is hated.
PROV|14|18|The simple inherit folly: but the prudent are crowned with knowledge.
PROV|14|19|The evil bow before the good; and the wicked at the gates of the righteous.
PROV|14|20|The poor is hated even of his own neighbour: but the rich hath many friends.
PROV|14|21|He that despiseth his neighbour sinneth: but he that hath mercy on the poor, happy is he.
PROV|14|22|Do they not err that devise evil? but mercy and truth shall be to them that devise good.
PROV|14|23|In all labour there is profit: but the talk of the lips tendeth only to penury.
PROV|14|24|The crown of the wise is their riches: but the foolishness of fools is folly.
PROV|14|25|A true witness delivereth souls: but a deceitful witness speaketh lies.
PROV|14|26|In the fear of the LORD is strong confidence: and his children shall have a place of refuge.
PROV|14|27|The fear of the LORD is a fountain of life, to depart from the snares of death.
PROV|14|28|In the multitude of people is the king's honour: but in the want of people is the destruction of the prince.
PROV|14|29|He that is slow to wrath is of great understanding: but he that is hasty of spirit exalteth folly.
PROV|14|30|A sound heart is the life of the flesh: but envy the rottenness of the bones.
PROV|14|31|He that oppresseth the poor reproacheth his Maker: but he that honoureth him hath mercy on the poor.
PROV|14|32|The wicked is driven away in his wickedness: but the righteous hath hope in his death.
PROV|14|33|Wisdom resteth in the heart of him that hath understanding: but that which is in the midst of fools is made known.
PROV|14|34|Righteousness exalteth a nation: but sin is a reproach to any people.
PROV|14|35|The king's favour is toward a wise servant: but his wrath is against him that causeth shame.
PROV|15|1|A soft answer turneth away wrath: but grievous words stir up anger.
PROV|15|2|The tongue of the wise useth knowledge aright: but the mouth of fools poureth out foolishness.
PROV|15|3|The eyes of the LORD are in every place, beholding the evil and the good.
PROV|15|4|A wholesome tongue is a tree of life: but perverseness therein is a breach in the spirit.
PROV|15|5|A fool despiseth his father's instruction: but he that regardeth reproof is prudent.
PROV|15|6|In the house of the righteous is much treasure: but in the revenues of the wicked is trouble.
PROV|15|7|The lips of the wise disperse knowledge: but the heart of the foolish doeth not so.
PROV|15|8|The sacrifice of the wicked is an abomination to the LORD: but the prayer of the upright is his delight.
PROV|15|9|The way of the wicked is an abomination unto the LORD: but he loveth him that followeth after righteousness.
PROV|15|10|Correction is grievous unto him that forsaketh the way: and he that hateth reproof shall die.
PROV|15|11|Hell and destruction are before the LORD: how much more then the hearts of the children of men?
PROV|15|12|A scorner loveth not one that reproveth him: neither will he go unto the wise.
PROV|15|13|A merry heart maketh a cheerful countenance: but by sorrow of the heart the spirit is broken.
PROV|15|14|The heart of him that hath understanding seeketh knowledge: but the mouth of fools feedeth on foolishness.
PROV|15|15|All the days of the afflicted are evil: but he that is of a merry heart hath a continual feast.
PROV|15|16|Better is little with the fear of the LORD than great treasure and trouble therewith.
PROV|15|17|Better is a dinner of herbs where love is, than a stalled ox and hatred therewith.
PROV|15|18|A wrathful man stirreth up strife: but he that is slow to anger appeaseth strife.
PROV|15|19|The way of the slothful man is as an hedge of thorns: but the way of the righteous is made plain.
PROV|15|20|A wise son maketh a glad father: but a foolish man despiseth his mother.
PROV|15|21|Folly is joy to him that is destitute of wisdom: but a man of understanding walketh uprightly.
PROV|15|22|Without counsel purposes are disappointed: but in the multitude of counsellors they are established.
PROV|15|23|A man hath joy by the answer of his mouth: and a word spoken in due season, how good is it!
PROV|15|24|The way of life is above to the wise, that he may depart from hell beneath.
PROV|15|25|The LORD will destroy the house of the proud: but he will establish the border of the widow.
PROV|15|26|The thoughts of the wicked are an abomination to the LORD: but the words of the pure are pleasant words.
PROV|15|27|He that is greedy of gain troubleth his own house; but he that hateth gifts shall live.
PROV|15|28|The heart of the righteous studieth to answer: but the mouth of the wicked poureth out evil things.
PROV|15|29|The LORD is far from the wicked: but he heareth the prayer of the righteous.
PROV|15|30|The light of the eyes rejoiceth the heart: and a good report maketh the bones fat.
PROV|15|31|The ear that heareth the reproof of life abideth among the wise.
PROV|15|32|He that refuseth instruction despiseth his own soul: but he that heareth reproof getteth understanding.
PROV|15|33|The fear of the LORD is the instruction of wisdom; and before honour is humility.
PROV|16|1|The preparations of the heart in man, and the answer of the tongue, is from the LORD.
PROV|16|2|All the ways of a man are clean in his own eyes; but the LORD weigheth the spirits.
PROV|16|3|Commit thy works unto the LORD, and thy thoughts shall be established.
PROV|16|4|The LORD hath made all things for himself: yea, even the wicked for the day of evil.
PROV|16|5|Every one that is proud in heart is an abomination to the LORD: though hand join in hand, he shall not be unpunished.
PROV|16|6|By mercy and truth iniquity is purged: and by the fear of the LORD men depart from evil.
PROV|16|7|When a man's ways please the LORD, he maketh even his enemies to be at peace with him.
PROV|16|8|Better is a little with righteousness than great revenues without right.
PROV|16|9|A man's heart deviseth his way: but the LORD directeth his steps.
PROV|16|10|A divine sentence is in the lips of the king: his mouth transgresseth not in judgment.
PROV|16|11|A just weight and balance are the LORD's: all the weights of the bag are his work.
PROV|16|12|It is an abomination to kings to commit wickedness: for the throne is established by righteousness.
PROV|16|13|Righteous lips are the delight of kings; and they love him that speaketh right.
PROV|16|14|The wrath of a king is as messengers of death: but a wise man will pacify it.
PROV|16|15|In the light of the king's countenance is life; and his favour is as a cloud of the latter rain.
PROV|16|16|How much better is it to get wisdom than gold! and to get understanding rather to be chosen than silver!
PROV|16|17|The highway of the upright is to depart from evil: he that keepeth his way preserveth his soul.
PROV|16|18|Pride goeth before destruction, and an haughty spirit before a fall.
PROV|16|19|Better it is to be of an humble spirit with the lowly, than to divide the spoil with the proud.
PROV|16|20|He that handleth a matter wisely shall find good: and whoso trusteth in the LORD, happy is he.
PROV|16|21|The wise in heart shall be called prudent: and the sweetness of the lips increaseth learning.
PROV|16|22|Understanding is a wellspring of life unto him that hath it: but the instruction of fools is folly.
PROV|16|23|The heart of the wise teacheth his mouth, and addeth learning to his lips.
PROV|16|24|Pleasant words are as an honeycomb, sweet to the soul, and health to the bones.
PROV|16|25|There is a way that seemeth right unto a man, but the end thereof are the ways of death.
PROV|16|26|He that laboureth laboureth for himself; for his mouth craveth it of him.
PROV|16|27|An ungodly man diggeth up evil: and in his lips there is as a burning fire.
PROV|16|28|A froward man soweth strife: and a whisperer separateth chief friends.
PROV|16|29|A violent man enticeth his neighbour, and leadeth him into the way that is not good.
PROV|16|30|He shutteth his eyes to devise froward things: moving his lips he bringeth evil to pass.
PROV|16|31|The hoary head is a crown of glory, if it be found in the way of righteousness.
PROV|16|32|He that is slow to anger is better than the mighty; and he that ruleth his spirit than he that taketh a city.
PROV|16|33|The lot is cast into the lap; but the whole disposing thereof is of the LORD.
PROV|17|1|Better is a dry morsel, and quietness therewith, than an house full of sacrifices with strife.
PROV|17|2|A wise servant shall have rule over a son that causeth shame, and shall have part of the inheritance among the brethren.
PROV|17|3|The fining pot is for silver, and the furnace for gold: but the LORD trieth the hearts.
PROV|17|4|A wicked doer giveth heed to false lips; and a liar giveth ear to a naughty tongue.
PROV|17|5|Whoso mocketh the poor reproacheth his Maker: and he that is glad at calamities shall not be unpunished.
PROV|17|6|Children's children are the crown of old men; and the glory of children are their fathers.
PROV|17|7|Excellent speech becometh not a fool: much less do lying lips a prince.
PROV|17|8|A gift is as a precious stone in the eyes of him that hath it: whithersoever it turneth, it prospereth.
PROV|17|9|He that covereth a transgression seeketh love; but he that repeateth a matter separateth very friends.
PROV|17|10|A reproof entereth more into a wise man than an hundred stripes into a fool.
PROV|17|11|An evil man seeketh only rebellion: therefore a cruel messenger shall be sent against him.
PROV|17|12|Let a bear robbed of her whelps meet a man, rather than a fool in his folly.
PROV|17|13|Whoso rewardeth evil for good, evil shall not depart from his house.
PROV|17|14|The beginning of strife is as when one letteth out water: therefore leave off contention, before it be meddled with.
PROV|17|15|He that justifieth the wicked, and he that condemneth the just, even they both are abomination to the LORD.
PROV|17|16|Wherefore is there a price in the hand of a fool to get wisdom, seeing he hath no heart to it?
PROV|17|17|A friend loveth at all times, and a brother is born for adversity.
PROV|17|18|A man void of understanding striketh hands, and becometh surety in the presence of his friend.
PROV|17|19|He loveth transgression that loveth strife: and he that exalteth his gate seeketh destruction.
PROV|17|20|He that hath a froward heart findeth no good: and he that hath a perverse tongue falleth into mischief.
PROV|17|21|He that begetteth a fool doeth it to his sorrow: and the father of a fool hath no joy.
PROV|17|22|A merry heart doeth good like a medicine: but a broken spirit drieth the bones.
PROV|17|23|A wicked man taketh a gift out of the bosom to pervert the ways of judgment.
PROV|17|24|Wisdom is before him that hath understanding; but the eyes of a fool are in the ends of the earth.
PROV|17|25|A foolish son is a grief to his father, and bitterness to her that bare him.
PROV|17|26|Also to punish the just is not good, nor to strike princes for equity.
PROV|17|27|He that hath knowledge spareth his words: and a man of understanding is of an excellent spirit.
PROV|17|28|Even a fool, when he holdeth his peace, is counted wise: and he that shutteth his lips is esteemed a man of understanding.
PROV|18|1|Through desire a man, having separated himself, seeketh and intermeddleth with all wisdom.
PROV|18|2|A fool hath no delight in understanding, but that his heart may discover itself.
PROV|18|3|When the wicked cometh, then cometh also contempt, and with ignominy reproach.
PROV|18|4|The words of a man's mouth are as deep waters, and the wellspring of wisdom as a flowing brook.
PROV|18|5|It is not good to accept the person of the wicked, to overthrow the righteous in judgment.
PROV|18|6|A fool's lips enter into contention, and his mouth calleth for strokes.
PROV|18|7|A fool's mouth is his destruction, and his lips are the snare of his soul.
PROV|18|8|The words of a talebearer are as wounds, and they go down into the innermost parts of the belly.
PROV|18|9|He also that is slothful in his work is brother to him that is a great waster.
PROV|18|10|The name of the LORD is a strong tower: the righteous runneth into it, and is safe.
PROV|18|11|The rich man's wealth is his strong city, and as an high wall in his own conceit.
PROV|18|12|Before destruction the heart of man is haughty, and before honour is humility.
PROV|18|13|He that answereth a matter before he heareth it, it is folly and shame unto him.
PROV|18|14|The spirit of a man will sustain his infirmity; but a wounded spirit who can bear?
PROV|18|15|The heart of the prudent getteth knowledge; and the ear of the wise seeketh knowledge.
PROV|18|16|A man's gift maketh room for him, and bringeth him before great men.
PROV|18|17|He that is first in his own cause seemeth just; but his neighbour cometh and searcheth him.
PROV|18|18|The lot causeth contentions to cease, and parteth between the mighty.
PROV|18|19|A brother offended is harder to be won than a strong city: and their contentions are like the bars of a castle.
PROV|18|20|A man's belly shall be satisfied with the fruit of his mouth; and with the increase of his lips shall he be filled.
PROV|18|21|Death and life are in the power of the tongue: and they that love it shall eat the fruit thereof.
PROV|18|22|Whoso findeth a wife findeth a good thing, and obtaineth favour of the LORD.
PROV|18|23|The poor useth intreaties; but the rich answereth roughly.
PROV|18|24|A man that hath friends must shew himself friendly: and there is a friend that sticketh closer than a brother.
PROV|19|1|Better is the poor that walketh in his integrity, than he that is perverse in his lips, and is a fool.
PROV|19|2|Also, that the soul be without knowledge, it is not good; and he that hasteth with his feet sinneth.
PROV|19|3|The foolishness of man perverteth his way: and his heart fretteth against the LORD.
PROV|19|4|Wealth maketh many friends; but the poor is separated from his neighbour.
PROV|19|5|A false witness shall not be unpunished, and he that speaketh lies shall not escape.
PROV|19|6|Many will intreat the favour of the prince: and every man is a friend to him that giveth gifts.
PROV|19|7|All the brethren of the poor do hate him: how much more do his friends go far from him? he pursueth them with words, yet they are wanting to him.
PROV|19|8|He that getteth wisdom loveth his own soul: he that keepeth understanding shall find good.
PROV|19|9|A false witness shall not be unpunished, and he that speaketh lies shall perish.
PROV|19|10|Delight is not seemly for a fool; much less for a servant to have rule over princes.
PROV|19|11|The discretion of a man deferreth his anger; and it is his glory to pass over a transgression.
PROV|19|12|The king's wrath is as the roaring of a lion; but his favour is as dew upon the grass.
PROV|19|13|A foolish son is the calamity of his father: and the contentions of a wife are a continual dropping.
PROV|19|14|House and riches are the inheritance of fathers: and a prudent wife is from the LORD.
PROV|19|15|Slothfulness casteth into a deep sleep; and an idle soul shall suffer hunger.
PROV|19|16|He that keepeth the commandment keepeth his own soul; but he that despiseth his ways shall die.
PROV|19|17|He that hath pity upon the poor lendeth unto the LORD; and that which he hath given will he pay him again.
PROV|19|18|Chasten thy son while there is hope, and let not thy soul spare for his crying.
PROV|19|19|A man of great wrath shall suffer punishment: for if thou deliver him, yet thou must do it again.
PROV|19|20|Hear counsel, and receive instruction, that thou mayest be wise in thy latter end.
PROV|19|21|There are many devices in a man's heart; nevertheless the counsel of the LORD, that shall stand.
PROV|19|22|The desire of a man is his kindness: and a poor man is better than a liar.
PROV|19|23|The fear of the LORD tendeth to life: and he that hath it shall abide satisfied; he shall not be visited with evil.
PROV|19|24|A slothful man hideth his hand in his bosom, and will not so much as bring it to his mouth again.
PROV|19|25|Smite a scorner, and the simple will beware: and reprove one that hath understanding, and he will understand knowledge.
PROV|19|26|He that wasteth his father, and chaseth away his mother, is a son that causeth shame, and bringeth reproach.
PROV|19|27|Cease, my son, to hear the instruction that causeth to err from the words of knowledge.
PROV|19|28|An ungodly witness scorneth judgment: and the mouth of the wicked devoureth iniquity.
PROV|19|29|Judgments are prepared for scorners, and stripes for the back of fools.
PROV|20|1|Wine is a mocker, strong drink is raging: and whosoever is deceived thereby is not wise.
PROV|20|2|The fear of a king is as the roaring of a lion: whoso provoketh him to anger sinneth against his own soul.
PROV|20|3|It is an honour for a man to cease from strife: but every fool will be meddling.
PROV|20|4|The sluggard will not plow by reason of the cold; therefore shall he beg in harvest, and have nothing.
PROV|20|5|Counsel in the heart of man is like deep water; but a man of understanding will draw it out.
PROV|20|6|Most men will proclaim every one his own goodness: but a faithful man who can find?
PROV|20|7|The just man walketh in his integrity: his children are blessed after him.
PROV|20|8|A king that sitteth in the throne of judgment scattereth away all evil with his eyes.
PROV|20|9|Who can say, I have made my heart clean, I am pure from my sin?
PROV|20|10|Divers weights, and divers measures, both of them are alike abomination to the LORD.
PROV|20|11|Even a child is known by his doings, whether his work be pure, and whether it be right.
PROV|20|12|The hearing ear, and the seeing eye, the LORD hath made even both of them.
PROV|20|13|Love not sleep, lest thou come to poverty; open thine eyes, and thou shalt be satisfied with bread.
PROV|20|14|It is naught, it is naught, saith the buyer: but when he is gone his way, then he boasteth.
PROV|20|15|There is gold, and a multitude of rubies: but the lips of knowledge are a precious jewel.
PROV|20|16|Take his garment that is surety for a stranger: and take a pledge of him for a strange woman.
PROV|20|17|Bread of deceit is sweet to a man; but afterwards his mouth shall be filled with gravel.
PROV|20|18|Every purpose is established by counsel: and with good advice make war.
PROV|20|19|He that goeth about as a talebearer revealeth secrets: therefore meddle not with him that flattereth with his lips.
PROV|20|20|Whoso curseth his father or his mother, his lamp shall be put out in obscure darkness.
PROV|20|21|An inheritance may be gotten hastily at the beginning; but the end thereof shall not be blessed.
PROV|20|22|Say not thou, I will recompense evil; but wait on the LORD, and he shall save thee.
PROV|20|23|Divers weights are an abomination unto the LORD; and a false balance is not good.
PROV|20|24|Man's goings are of the LORD; how can a man then understand his own way?
PROV|20|25|It is a snare to the man who devoureth that which is holy, and after vows to make enquiry.
PROV|20|26|A wise king scattereth the wicked, and bringeth the wheel over them.
PROV|20|27|The spirit of man is the candle of the LORD, searching all the inward parts of the belly.
PROV|20|28|Mercy and truth preserve the king: and his throne is upholden by mercy.
PROV|20|29|The glory of young men is their strength: and the beauty of old men is the grey head.
PROV|20|30|The blueness of a wound cleanseth away evil: so do stripes the inward parts of the belly.
PROV|21|1|The king's heart is in the hand of the LORD, as the rivers of water: he turneth it whithersoever he will.
PROV|21|2|Every way of a man is right in his own eyes: but the LORD pondereth the hearts.
PROV|21|3|To do justice and judgment is more acceptable to the LORD than sacrifice.
PROV|21|4|An high look, and a proud heart, and the plowing of the wicked, is sin.
PROV|21|5|The thoughts of the diligent tend only to plenteousness; but of every one that is hasty only to want.
PROV|21|6|The getting of treasures by a lying tongue is a vanity tossed to and fro of them that seek death.
PROV|21|7|The robbery of the wicked shall destroy them; because they refuse to do judgment.
PROV|21|8|The way of man is froward and strange: but as for the pure, his work is right.
PROV|21|9|It is better to dwell in a corner of the housetop, than with a brawling woman in a wide house.
PROV|21|10|The soul of the wicked desireth evil: his neighbour findeth no favour in his eyes.
PROV|21|11|When the scorner is punished, the simple is made wise: and when the wise is instructed, he receiveth knowledge.
PROV|21|12|The righteous man wisely considereth the house of the wicked: but God overthroweth the wicked for their wickedness.
PROV|21|13|Whoso stoppeth his ears at the cry of the poor, he also shall cry himself, but shall not be heard.
PROV|21|14|A gift in secret pacifieth anger: and a reward in the bosom strong wrath.
PROV|21|15|It is joy to the just to do judgment: but destruction shall be to the workers of iniquity.
PROV|21|16|The man that wandereth out of the way of understanding shall remain in the congregation of the dead.
PROV|21|17|He that loveth pleasure shall be a poor man: he that loveth wine and oil shall not be rich.
PROV|21|18|The wicked shall be a ransom for the righteous, and the transgressor for the upright.
PROV|21|19|It is better to dwell in the wilderness, than with a contentious and an angry woman.
PROV|21|20|There is treasure to be desired and oil in the dwelling of the wise; but a foolish man spendeth it up.
PROV|21|21|He that followeth after righteousness and mercy findeth life, righteousness, and honour.
PROV|21|22|A wise man scaleth the city of the mighty, and casteth down the strength of the confidence thereof.
PROV|21|23|Whoso keepeth his mouth and his tongue keepeth his soul from troubles.
PROV|21|24|Proud and haughty scorner is his name, who dealeth in proud wrath.
PROV|21|25|The desire of the slothful killeth him; for his hands refuse to labour.
PROV|21|26|He coveteth greedily all the day long: but the righteous giveth and spareth not.
PROV|21|27|The sacrifice of the wicked is abomination: how much more, when he bringeth it with a wicked mind?
PROV|21|28|A false witness shall perish: but the man that heareth speaketh constantly.
PROV|21|29|A wicked man hardeneth his face: but as for the upright, he directeth his way.
PROV|21|30|There is no wisdom nor understanding nor counsel against the LORD.
PROV|21|31|The horse is prepared against the day of battle: but safety is of the LORD.
PROV|22|1|A GOOD name is rather to be chosen than great riches, and loving favour rather than silver and gold.
PROV|22|2|The rich and poor meet together: the LORD is the maker of them all.
PROV|22|3|A prudent man foreseeth the evil, and hideth himself: but the simple pass on, and are punished.
PROV|22|4|By humility and the fear of the LORD are riches, and honour, and life.
PROV|22|5|Thorns and snares are in the way of the froward: he that doth keep his soul shall be far from them.
PROV|22|6|Train up a child in the way he should go: and when he is old, he will not depart from it.
PROV|22|7|The rich ruleth over the poor, and the borrower is servant to the lender.
PROV|22|8|He that soweth iniquity shall reap vanity: and the rod of his anger shall fail.
PROV|22|9|He that hath a bountiful eye shall be blessed; for he giveth of his bread to the poor.
PROV|22|10|Cast out the scorner, and contention shall go out; yea, strife and reproach shall cease.
PROV|22|11|He that loveth pureness of heart, for the grace of his lips the king shall be his friend.
PROV|22|12|The eyes of the LORD preserve knowledge, and he overthroweth the words of the transgressor.
PROV|22|13|The slothful man saith, There is a lion without, I shall be slain in the streets.
PROV|22|14|The mouth of strange women is a deep pit: he that is abhorred of the LORD shall fall therein.
PROV|22|15|Foolishness is bound in the heart of a child; but the rod of correction shall drive it far from him.
PROV|22|16|He that oppresseth the poor to increase his riches, and he that giveth to the rich, shall surely come to want.
PROV|22|17|Bow down thine ear, and hear the words of the wise, and apply thine heart unto my knowledge.
PROV|22|18|For it is a pleasant thing if thou keep them within thee; they shall withal be fitted in thy lips.
PROV|22|19|That thy trust may be in the LORD, I have made known to thee this day, even to thee.
PROV|22|20|Have not I written to thee excellent things in counsels and knowledge,
PROV|22|21|That I might make thee know the certainty of the words of truth; that thou mightest answer the words of truth to them that send unto thee?
PROV|22|22|Rob not the poor, because he is poor: neither oppress the afflicted in the gate:
PROV|22|23|For the LORD will plead their cause, and spoil the soul of those that spoiled them.
PROV|22|24|Make no friendship with an angry man; and with a furious man thou shalt not go:
PROV|22|25|Lest thou learn his ways, and get a snare to thy soul.
PROV|22|26|Be not thou one of them that strike hands, or of them that are sureties for debts.
PROV|22|27|If thou hast nothing to pay, why should he take away thy bed from under thee?
PROV|22|28|Remove not the ancient landmark, which thy fathers have set.
PROV|22|29|Seest thou a man diligent in his business? he shall stand before kings; he shall not stand before mean men.
PROV|23|1|When thou sittest to eat with a ruler, consider diligently what is before thee:
PROV|23|2|And put a knife to thy throat, if thou be a man given to appetite.
PROV|23|3|Be not desirous of his dainties: for they are deceitful meat.
PROV|23|4|Labour not to be rich: cease from thine own wisdom.
PROV|23|5|Wilt thou set thine eyes upon that which is not? for riches certainly make themselves wings; they fly away as an eagle toward heaven.
PROV|23|6|Eat thou not the bread of him that hath an evil eye, neither desire thou his dainty meats:
PROV|23|7|For as he thinketh in his heart, so is he: Eat and drink, saith he to thee; but his heart is not with thee.
PROV|23|8|The morsel which thou hast eaten shalt thou vomit up, and lose thy sweet words.
PROV|23|9|Speak not in the ears of a fool: for he will despise the wisdom of thy words.
PROV|23|10|Remove not the old landmark; and enter not into the fields of the fatherless:
PROV|23|11|For their redeemer is mighty; he shall plead their cause with thee.
PROV|23|12|Apply thine heart unto instruction, and thine ears to the words of knowledge.
PROV|23|13|Withhold not correction from the child: for if thou beatest him with the rod, he shall not die.
PROV|23|14|Thou shalt beat him with the rod, and shalt deliver his soul from hell.
PROV|23|15|My son, if thine heart be wise, my heart shall rejoice, even mine.
PROV|23|16|Yea, my reins shall rejoice, when thy lips speak right things.
PROV|23|17|Let not thine heart envy sinners: but be thou in the fear of the LORD all the day long.
PROV|23|18|For surely there is an end; and thine expectation shall not be cut off.
PROV|23|19|Hear thou, my son, and be wise, and guide thine heart in the way.
PROV|23|20|Be not among winebibbers; among riotous eaters of flesh:
PROV|23|21|For the drunkard and the glutton shall come to poverty: and drowsiness shall clothe a man with rags.
PROV|23|22|Hearken unto thy father that begat thee, and despise not thy mother when she is old.
PROV|23|23|Buy the truth, and sell it not; also wisdom, and instruction, and understanding.
PROV|23|24|The father of the righteous shall greatly rejoice: and he that begetteth a wise child shall have joy of him.
PROV|23|25|Thy father and thy mother shall be glad, and she that bare thee shall rejoice.
PROV|23|26|My son, give me thine heart, and let thine eyes observe my ways.
PROV|23|27|For a whore is a deep ditch; and a strange woman is a narrow pit.
PROV|23|28|She also lieth in wait as for a prey, and increaseth the transgressors among men.
PROV|23|29|Who hath woe? who hath sorrow? who hath contentions? who hath babbling? who hath wounds without cause? who hath redness of eyes?
PROV|23|30|They that tarry long at the wine; they that go to seek mixed wine.
PROV|23|31|Look not thou upon the wine when it is red, when it giveth his colour in the cup, when it moveth itself aright.
PROV|23|32|At the last it biteth like a serpent, and stingeth like an adder.
PROV|23|33|Thine eyes shall behold strange women, and thine heart shall utter perverse things.
PROV|23|34|Yea, thou shalt be as he that lieth down in the midst of the sea, or as he that lieth upon the top of a mast.
PROV|23|35|They have stricken me, shalt thou say, and I was not sick; they have beaten me, and I felt it not: when shall I awake? I will seek it yet again.
PROV|24|1|Be not thou envious against evil men, neither desire to be with them.
PROV|24|2|For their heart studieth destruction, and their lips talk of mischief.
PROV|24|3|Through wisdom is an house builded; and by understanding it is established:
PROV|24|4|And by knowledge shall the chambers be filled with all precious and pleasant riches.
PROV|24|5|A wise man is strong; yea, a man of knowledge increaseth strength.
PROV|24|6|For by wise counsel thou shalt make thy war: and in multitude of counsellors there is safety.
PROV|24|7|Wisdom is too high for a fool: he openeth not his mouth in the gate.
PROV|24|8|He that deviseth to do evil shall be called a mischievous person.
PROV|24|9|The thought of foolishness is sin: and the scorner is an abomination to men.
PROV|24|10|If thou faint in the day of adversity, thy strength is small.
PROV|24|11|If thou forbear to deliver them that are drawn unto death, and those that are ready to be slain;
PROV|24|12|If thou sayest, Behold, we knew it not; doth not he that pondereth the heart consider it? and he that keepeth thy soul, doth not he know it? and shall not he render to every man according to his works?
PROV|24|13|My son, eat thou honey, because it is good; and the honeycomb, which is sweet to thy taste:
PROV|24|14|So shall the knowledge of wisdom be unto thy soul: when thou hast found it, then there shall be a reward, and thy expectation shall not be cut off.
PROV|24|15|Lay not wait, O wicked man, against the dwelling of the righteous; spoil not his resting place:
PROV|24|16|For a just man falleth seven times, and riseth up again: but the wicked shall fall into mischief.
PROV|24|17|Rejoice not when thine enemy falleth, and let not thine heart be glad when he stumbleth:
PROV|24|18|Lest the LORD see it, and it displease him, and he turn away his wrath from him.
PROV|24|19|Fret not thyself because of evil men, neither be thou envious at the wicked:
PROV|24|20|For there shall be no reward to the evil man; the candle of the wicked shall be put out.
PROV|24|21|My son, fear thou the LORD and the king: and meddle not with them that are given to change:
PROV|24|22|For their calamity shall rise suddenly; and who knoweth the ruin of them both?
PROV|24|23|These things also belong to the wise. It is not good to have respect of persons in judgment.
PROV|24|24|He that saith unto the wicked, Thou are righteous; him shall the people curse, nations shall abhor him:
PROV|24|25|But to them that rebuke him shall be delight, and a good blessing shall come upon them.
PROV|24|26|Every man shall kiss his lips that giveth a right answer.
PROV|24|27|Prepare thy work without, and make it fit for thyself in the field; and afterwards build thine house.
PROV|24|28|Be not a witness against thy neighbour without cause; and deceive not with thy lips.
PROV|24|29|Say not, I will do so to him as he hath done to me: I will render to the man according to his work.
PROV|24|30|I went by the field of the slothful, and by the vineyard of the man void of understanding;
PROV|24|31|And, lo, it was all grown over with thorns, and nettles had covered the face thereof, and the stone wall thereof was broken down.
PROV|24|32|Then I saw, and considered it well: I looked upon it, and received instruction.
PROV|24|33|Yet a little sleep, a little slumber, a little folding of the hands to sleep:
PROV|24|34|So shall thy poverty come as one that travelleth; and thy want as an armed man.
PROV|25|1|These are also proverbs of Solomon, which the men of Hezekiah king of Judah copied out.
PROV|25|2|It is the glory of God to conceal a thing: but the honour of kings is to search out a matter.
PROV|25|3|The heaven for height, and the earth for depth, and the heart of kings is unsearchable.
PROV|25|4|Take away the dross from the silver, and there shall come forth a vessel for the finer.
PROV|25|5|Take away the wicked from before the king, and his throne shall be established in righteousness.
PROV|25|6|Put not forth thyself in the presence of the king, and stand not in the place of great men:
PROV|25|7|For better it is that it be said unto thee, Come up hither; than that thou shouldest be put lower in the presence of the prince whom thine eyes have seen.
PROV|25|8|Go not forth hastily to strive, lest thou know not what to do in the end thereof, when thy neighbour hath put thee to shame.
PROV|25|9|Debate thy cause with thy neighbour himself; and discover not a secret to another:
PROV|25|10|Lest he that heareth it put thee to shame, and thine infamy turn not away.
PROV|25|11|A word fitly spoken is like apples of gold in pictures of silver.
PROV|25|12|As an earring of gold, and an ornament of fine gold, so is a wise reprover upon an obedient ear.
PROV|25|13|As the cold of snow in the time of harvest, so is a faithful messenger to them that send him: for he refresheth the soul of his masters.
PROV|25|14|Whoso boasteth himself of a false gift is like clouds and wind without rain.
PROV|25|15|By long forbearing is a prince persuaded, and a soft tongue breaketh the bone.
PROV|25|16|Hast thou found honey? eat so much as is sufficient for thee, lest thou be filled therewith, and vomit it.
PROV|25|17|Withdraw thy foot from thy neighbour's house; lest he be weary of thee, and so hate thee.
PROV|25|18|A man that beareth false witness against his neighbour is a maul, and a sword, and a sharp arrow.
PROV|25|19|Confidence in an unfaithful man in time of trouble is like a broken tooth, and a foot out of joint.
PROV|25|20|As he that taketh away a garment in cold weather, and as vinegar upon nitre, so is he that singeth songs to an heavy heart.
PROV|25|21|If thine enemy be hungry, give him bread to eat; and if he be thirsty, give him water to drink:
PROV|25|22|For thou shalt heap coals of fire upon his head, and the LORD shall reward thee.
PROV|25|23|The north wind driveth away rain: so doth an angry countenance a backbiting tongue.
PROV|25|24|It is better to dwell in the corner of the housetop, than with a brawling woman and in a wide house.
PROV|25|25|As cold waters to a thirsty soul, so is good news from a far country.
PROV|25|26|A righteous man falling down before the wicked is as a troubled fountain, and a corrupt spring.
PROV|25|27|It is not good to eat much honey: so for men to search their own glory is not glory.
PROV|25|28|He that hath no rule over his own spirit is like a city that is broken down, and without walls.
PROV|26|1|As snow in summer, and as rain in harvest, so honour is not seemly for a fool.
PROV|26|2|As the bird by wandering, as the swallow by flying, so the curse causeless shall not come.
PROV|26|3|A whip for the horse, a bridle for the ass, and a rod for the fool's back.
PROV|26|4|Answer not a fool according to his folly, lest thou also be like unto him.
PROV|26|5|Answer a fool according to his folly, lest he be wise in his own conceit.
PROV|26|6|He that sendeth a message by the hand of a fool cutteth off the feet, and drinketh damage.
PROV|26|7|The legs of the lame are not equal: so is a parable in the mouth of fools.
PROV|26|8|As he that bindeth a stone in a sling, so is he that giveth honour to a fool.
PROV|26|9|As a thorn goeth up into the hand of a drunkard, so is a parable in the mouths of fools.
PROV|26|10|The great God that formed all things both rewardeth the fool, and rewardeth transgressors.
PROV|26|11|As a dog returneth to his vomit, so a fool returneth to his folly.
PROV|26|12|Seest thou a man wise in his own conceit? there is more hope of a fool than of him.
PROV|26|13|The slothful man saith, There is a lion in the way; a lion is in the streets.
PROV|26|14|As the door turneth upon his hinges, so doth the slothful upon his bed.
PROV|26|15|The slothful hideth his hand in his bosom; it grieveth him to bring it again to his mouth.
PROV|26|16|The sluggard is wiser in his own conceit than seven men that can render a reason.
PROV|26|17|He that passeth by, and meddleth with strife belonging not to him, is like one that taketh a dog by the ears.
PROV|26|18|As a mad man who casteth firebrands, arrows, and death,
PROV|26|19|So is the man that deceiveth his neighbour, and saith, Am not I in sport?
PROV|26|20|Where no wood is, there the fire goeth out: so where there is no talebearer, the strife ceaseth.
PROV|26|21|As coals are to burning coals, and wood to fire; so is a contentious man to kindle strife.
PROV|26|22|The words of a talebearer are as wounds, and they go down into the innermost parts of the belly.
PROV|26|23|Burning lips and a wicked heart are like a potsherd covered with silver dross.
PROV|26|24|He that hateth dissembleth with his lips, and layeth up deceit within him;
PROV|26|25|When he speaketh fair, believe him not: for there are seven abominations in his heart.
PROV|26|26|Whose hatred is covered by deceit, his wickedness shall be shewed before the whole congregation.
PROV|26|27|Whoso diggeth a pit shall fall therein: and he that rolleth a stone, it will return upon him.
PROV|26|28|A lying tongue hateth those that are afflicted by it; and a flattering mouth worketh ruin.
PROV|27|1|Boast not thyself of to morrow; for thou knowest not what a day may bring forth.
PROV|27|2|Let another man praise thee, and not thine own mouth; a stranger, and not thine own lips.
PROV|27|3|A stone is heavy, and the sand weighty; but a fool's wrath is heavier than them both.
PROV|27|4|Wrath is cruel, and anger is outrageous; but who is able to stand before envy?
PROV|27|5|Open rebuke is better than secret love.
PROV|27|6|Faithful are the wounds of a friend; but the kisses of an enemy are deceitful.
PROV|27|7|The full soul loatheth an honeycomb; but to the hungry soul every bitter thing is sweet.
PROV|27|8|As a bird that wandereth from her nest, so is a man that wandereth from his place.
PROV|27|9|Ointment and perfume rejoice the heart: so doth the sweetness of a man's friend by hearty counsel.
PROV|27|10|Thine own friend, and thy father's friend, forsake not; neither go into thy brother's house in the day of thy calamity: for better is a neighbour that is near than a brother far off.
PROV|27|11|My son, be wise, and make my heart glad, that I may answer him that reproacheth me.
PROV|27|12|A prudent man foreseeth the evil, and hideth himself; but the simple pass on, and are punished.
PROV|27|13|Take his garment that is surety for a stranger, and take a pledge of him for a strange woman.
PROV|27|14|He that blesseth his friend with a loud voice, rising early in the morning, it shall be counted a curse to him.
PROV|27|15|A continual dropping in a very rainy day and a contentious woman are alike.
PROV|27|16|Whosoever hideth her hideth the wind, and the ointment of his right hand, which bewrayeth itself.
PROV|27|17|Iron sharpeneth iron; so a man sharpeneth the countenance of his friend.
PROV|27|18|Whoso keepeth the fig tree shall eat the fruit thereof: so he that waiteth on his master shall be honoured.
PROV|27|19|As in water face answereth to face, so the heart of man to man.
PROV|27|20|Hell and destruction are never full; so the eyes of man are never satisfied.
PROV|27|21|As the fining pot for silver, and the furnace for gold; so is a man to his praise.
PROV|27|22|Though thou shouldest bray a fool in a mortar among wheat with a pestle, yet will not his foolishness depart from him.
PROV|27|23|Be thou diligent to know the state of thy flocks, and look well to thy herds.
PROV|27|24|For riches are not for ever: and doth the crown endure to every generation?
PROV|27|25|The hay appeareth, and the tender grass sheweth itself, and herbs of the mountains are gathered.
PROV|27|26|The lambs are for thy clothing, and the goats are the price of the field.
PROV|27|27|And thou shalt have goats' milk enough for thy food, for the food of thy household, and for the maintenance for thy maidens.
PROV|28|1|The wicked flee when no man pursueth: but the righteous are bold as a lion.
PROV|28|2|For the transgression of a land many are the princes thereof: but by a man of understanding and knowledge the state thereof shall be prolonged.
PROV|28|3|A poor man that oppresseth the poor is like a sweeping rain which leaveth no food.
PROV|28|4|They that forsake the law praise the wicked: but such as keep the law contend with them.
PROV|28|5|Evil men understand not judgment: but they that seek the LORD understand all things.
PROV|28|6|Better is the poor that walketh in his uprightness, than he that is perverse in his ways, though he be rich.
PROV|28|7|Whoso keepeth the law is a wise son: but he that is a companion of riotous men shameth his father.
PROV|28|8|He that by usury and unjust gain increaseth his substance, he shall gather it for him that will pity the poor.
PROV|28|9|He that turneth away his ear from hearing the law, even his prayer shall be abomination.
PROV|28|10|Whoso causeth the righteous to go astray in an evil way, he shall fall himself into his own pit: but the upright shall have good things in possession.
PROV|28|11|The rich man is wise in his own conceit; but the poor that hath understanding searcheth him out.
PROV|28|12|When righteous men do rejoice, there is great glory: but when the wicked rise, a man is hidden.
PROV|28|13|He that covereth his sins shall not prosper: but whoso confesseth and forsaketh them shall have mercy.
PROV|28|14|Happy is the man that feareth alway: but he that hardeneth his heart shall fall into mischief.
PROV|28|15|As a roaring lion, and a ranging bear; so is a wicked ruler over the poor people.
PROV|28|16|The prince that wanteth understanding is also a great oppressor: but he that hateth covetousness shall prolong his days.
PROV|28|17|A man that doeth violence to the blood of any person shall flee to the pit; let no man stay him.
PROV|28|18|Whoso walketh uprightly shall be saved: but he that is perverse in his ways shall fall at once.
PROV|28|19|He that tilleth his land shall have plenty of bread: but he that followeth after vain persons shall have poverty enough.
PROV|28|20|A faithful man shall abound with blessings: but he that maketh haste to be rich shall not be innocent.
PROV|28|21|To have respect of persons is not good: for for a piece of bread that man will transgress.
PROV|28|22|He that hasteth to be rich hath an evil eye, and considereth not that poverty shall come upon him.
PROV|28|23|He that rebuketh a man afterwards shall find more favour than he that flattereth with the tongue.
PROV|28|24|Whoso robbeth his father or his mother, and saith, It is no transgression; the same is the companion of a destroyer.
PROV|28|25|He that is of a proud heart stirreth up strife: but he that putteth his trust in the LORD shall be made fat.
PROV|28|26|He that trusteth in his own heart is a fool: but whoso walketh wisely, he shall be delivered.
PROV|28|27|He that giveth unto the poor shall not lack: but he that hideth his eyes shall have many a curse.
PROV|28|28|When the wicked rise, men hide themselves: but when they perish, the righteous increase.
PROV|29|1|He, that being often reproved hardeneth his neck, shall suddenly be destroyed, and that without remedy.
PROV|29|2|When the righteous are in authority, the people rejoice: but when the wicked beareth rule, the people mourn.
PROV|29|3|Whoso loveth wisdom rejoiceth his father: but he that keepeth company with harlots spendeth his substance.
PROV|29|4|The king by judgment establisheth the land: but he that receiveth gifts overthroweth it.
PROV|29|5|A man that flattereth his neighbour spreadeth a net for his feet.
PROV|29|6|In the transgression of an evil man there is a snare: but the righteous doth sing and rejoice.
PROV|29|7|The righteous considereth the cause of the poor: but the wicked regardeth not to know it.
PROV|29|8|Scornful men bring a city into a snare: but wise men turn away wrath.
PROV|29|9|If a wise man contendeth with a foolish man, whether he rage or laugh, there is no rest.
PROV|29|10|The bloodthirsty hate the upright: but the just seek his soul.
PROV|29|11|A fool uttereth all his mind: but a wise man keepeth it in till afterwards.
PROV|29|12|If a ruler hearken to lies, all his servants are wicked.
PROV|29|13|The poor and the deceitful man meet together: the LORD lighteneth both their eyes.
PROV|29|14|The king that faithfully judgeth the poor, his throne shall be established for ever.
PROV|29|15|The rod and reproof give wisdom: but a child left to himself bringeth his mother to shame.
PROV|29|16|When the wicked are multiplied, transgression increaseth: but the righteous shall see their fall.
PROV|29|17|Correct thy son, and he shall give thee rest; yea, he shall give delight unto thy soul.
PROV|29|18|Where there is no vision, the people perish: but he that keepeth the law, happy is he.
PROV|29|19|A servant will not be corrected by words: for though he understand he will not answer.
PROV|29|20|Seest thou a man that is hasty in his words? there is more hope of a fool than of him.
PROV|29|21|He that delicately bringeth up his servant from a child shall have him become his son at the length.
PROV|29|22|An angry man stirreth up strife, and a furious man aboundeth in transgression.
PROV|29|23|A man's pride shall bring him low: but honour shall uphold the humble in spirit.
PROV|29|24|Whoso is partner with a thief hateth his own soul: he heareth cursing, and bewrayeth it not.
PROV|29|25|The fear of man bringeth a snare: but whoso putteth his trust in the LORD shall be safe.
PROV|29|26|Many seek the ruler's favour; but every man's judgment cometh from the LORD.
PROV|29|27|An unjust man is an abomination to the just: and he that is upright in the way is abomination to the wicked.
PROV|30|1|The words of Agur the son of Jakeh, even the prophecy: the man spake unto Ithiel, even unto Ithiel and Ucal,
PROV|30|2|Surely I am more brutish than any man, and have not the understanding of a man.
PROV|30|3|I neither learned wisdom, nor have the knowledge of the holy.
PROV|30|4|Who hath ascended up into heaven, or descended? who hath gathered the wind in his fists? who hath bound the waters in a garment? who hath established all the ends of the earth? what is his name, and what is his son's name, if thou canst tell?
PROV|30|5|Every word of God is pure: he is a shield unto them that put their trust in him.
PROV|30|6|Add thou not unto his words, lest he reprove thee, and thou be found a liar.
PROV|30|7|Two things have I required of thee; deny me them not before I die:
PROV|30|8|Remove far from me vanity and lies: give me neither poverty nor riches; feed me with food convenient for me:
PROV|30|9|Lest I be full, and deny thee, and say, Who is the LORD? or lest I be poor, and steal, and take the name of my God in vain.
PROV|30|10|Accuse not a servant unto his master, lest he curse thee, and thou be found guilty.
PROV|30|11|There is a generation that curseth their father, and doth not bless their mother.
PROV|30|12|There is a generation that are pure in their own eyes, and yet is not washed from their filthiness.
PROV|30|13|There is a generation, O how lofty are their eyes! and their eyelids are lifted up.
PROV|30|14|There is a generation, whose teeth are as swords, and their jaw teeth as knives, to devour the poor from off the earth, and the needy from among men.
PROV|30|15|The horseleach hath two daughters, crying, Give, give. There are three things that are never satisfied, yea, four things say not, It is enough:
PROV|30|16|The grave; and the barren womb; the earth that is not filled with water; and the fire that saith not, It is enough.
PROV|30|17|The eye that mocketh at his father, and despiseth to obey his mother, the ravens of the valley shall pick it out, and the young eagles shall eat it.
PROV|30|18|There be three things which are too wonderful for me, yea, four which I know not:
PROV|30|19|The way of an eagle in the air; the way of a serpent upon a rock; the way of a ship in the midst of the sea; and the way of a man with a maid.
PROV|30|20|Such is the way of an adulterous woman; she eateth, and wipeth her mouth, and saith, I have done no wickedness.
PROV|30|21|For three things the earth is disquieted, and for four which it cannot bear:
PROV|30|22|For a servant when he reigneth; and a fool when he is filled with meat;
PROV|30|23|For an odious woman when she is married; and an handmaid that is heir to her mistress.
PROV|30|24|There be four things which are little upon the earth, but they are exceeding wise:
PROV|30|25|The ants are a people not strong, yet they prepare their meat in the summer;
PROV|30|26|The conies are but a feeble folk, yet make they their houses in the rocks;
PROV|30|27|The locusts have no king, yet go they forth all of them by bands;
PROV|30|28|The spider taketh hold with her hands, and is in kings' palaces.
PROV|30|29|There be three things which go well, yea, four are comely in going:
PROV|30|30|A lion which is strongest among beasts, and turneth not away for any;
PROV|30|31|A greyhound; an he goat also; and a king, against whom there is no rising up.
PROV|30|32|If thou hast done foolishly in lifting up thyself, or if thou hast thought evil, lay thine hand upon thy mouth.
PROV|30|33|Surely the churning of milk bringeth forth butter, and the wringing of the nose bringeth forth blood: so the forcing of wrath bringeth forth strife.
PROV|31|1|The words of king Lemuel, the prophecy that his mother taught him.
PROV|31|2|What, my son? and what, the son of my womb? and what, the son of my vows?
PROV|31|3|Give not thy strength unto women, nor thy ways to that which destroyeth kings.
PROV|31|4|It is not for kings, O Lemuel, it is not for kings to drink wine; nor for princes strong drink:
PROV|31|5|Lest they drink, and forget the law, and pervert the judgment of any of the afflicted.
PROV|31|6|Give strong drink unto him that is ready to perish, and wine unto those that be of heavy hearts.
PROV|31|7|Let him drink, and forget his poverty, and remember his misery no more.
PROV|31|8|Open thy mouth for the dumb in the cause of all such as are appointed to destruction.
PROV|31|9|Open thy mouth, judge righteously, and plead the cause of the poor and needy.
PROV|31|10|Who can find a virtuous woman? for her price is far above rubies.
PROV|31|11|The heart of her husband doth safely trust in her, so that he shall have no need of spoil.
PROV|31|12|She will do him good and not evil all the days of her life.
PROV|31|13|She seeketh wool, and flax, and worketh willingly with her hands.
PROV|31|14|She is like the merchants' ships; she bringeth her food from afar.
PROV|31|15|She riseth also while it is yet night, and giveth meat to her household, and a portion to her maidens.
PROV|31|16|She considereth a field, and buyeth it: with the fruit of her hands she planteth a vineyard.
PROV|31|17|She girdeth her loins with strength, and strengtheneth her arms.
PROV|31|18|She perceiveth that her merchandise is good: her candle goeth not out by night.
PROV|31|19|She layeth her hands to the spindle, and her hands hold the distaff.
PROV|31|20|She stretcheth out her hand to the poor; yea, she reacheth forth her hands to the needy.
PROV|31|21|She is not afraid of the snow for her household: for all her household are clothed with scarlet.
PROV|31|22|She maketh herself coverings of tapestry; her clothing is silk and purple.
PROV|31|23|Her husband is known in the gates, when he sitteth among the elders of the land.
PROV|31|24|She maketh fine linen, and selleth it; and delivereth girdles unto the merchant.
PROV|31|25|Strength and honour are her clothing; and she shall rejoice in time to come.
PROV|31|26|She openeth her mouth with wisdom; and in her tongue is the law of kindness.
PROV|31|27|She looketh well to the ways of her household, and eateth not the bread of idleness.
PROV|31|28|Her children arise up, and call her blessed; her husband also, and he praiseth her.
PROV|31|29|Many daughters have done virtuously, but thou excellest them all.
PROV|31|30|Favour is deceitful, and beauty is vain: but a woman that feareth the LORD, she shall be praised.
PROV|31|31|Give her of the fruit of her hands; and let her own works praise her in the gates.
