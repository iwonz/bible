JOHN|1|1|In principio erat Verbum, et Verbum erat apud Deum, et Deus erat Verbum.
JOHN|1|2|Hoc erat in principio apud Deum.
JOHN|1|3|Omnia per ipsum facta sunt, et sine ipso factum est nihil, quod factum est;
JOHN|1|4|in ipso vita erat, et vita erat lux hominum,
JOHN|1|5|et lux in tenebris lucet, et tenebrae eam non comprehenderunt.
JOHN|1|6|Fuit homo missus a Deo, cui nomen erat Ioannes;
JOHN|1|7|hic venit in testimonium, ut testimonium perhiberet de lumine, ut omnes crederent per illum.
JOHN|1|8|Non erat ille lux, sed ut testimonium perhiberet de lumine.
JOHN|1|9|Erat lux vera, quae illuminat omnem hominem, veniens in mundum.
JOHN|1|10|In mundo erat, et mundus per ipsum factus est, et mundus eum non cognovit.
JOHN|1|11|In propria venit, et sui eum non receperunt.
JOHN|1|12|Quotquot autem acceperunt eum, dedit eis potestatem filios Dei fieri, his, qui credunt in nomine eius,
JOHN|1|13|qui non ex sanguinibus neque ex voluntate carnis neque ex voluntate viri, sed ex Deo nati sunt.
JOHN|1|14|Et Verbum caro factum est et habitavit in nobis; et vidimus gloriam eius, gloriam quasi Unigeniti a Patre, plenum gratiae et veritatis.
JOHN|1|15|Ioannes testimonium perhibet de ipso et clamat dicens: " Hic erat, quem dixi: Qui post me venturus est, ante me factus est, quia prior me erat ".
JOHN|1|16|Et de plenitudine eius nos omnes accepimus, et gratiam pro gratia;
JOHN|1|17|quia lex per Moysen data est, gratia et veritas per Iesum Christum facta est.
JOHN|1|18|Deum nemo vidit umquam; unigenitus Deus, qui est in sinum Patris, ipse enarravit.
JOHN|1|19|Et hoc est testimonium Ioannis, quando miserunt ad eum Iudaei ab Hierosolymis sacerdotes et Levitas, ut interrogarent eum: " Tu quis es? ".
JOHN|1|20|Et confessus est et non negavit; et confessus est: " Non sum ego Christus ".
JOHN|1|21|Et interrogaverunt eum: " Quid ergo? Elias es tu? ". Et dicit: " Non sum ". " Propheta es tu? ". Et respondit: " Non ".
JOHN|1|22|Dixerunt ergo ei: " Quis es? Ut responsum demus his, qui miserunt nos. Quid dicis de teipso? ".
JOHN|1|23|Ait: Ego vox clamantis in deserto:Dirigite viam Domini",sicut dixit Isaias propheta ".
JOHN|1|24|Et qui missi fuerant, erant ex pharisaeis;
JOHN|1|25|et interrogaverunt eum et dixerunt ei: " Quid ergo baptizas, si tu non es Christus neque Elias neque propheta? ".
JOHN|1|26|Respondit eis Ioannes dicens: " Ego baptizo in aqua; medius vestrum stat, quem vos non scitis,
JOHN|1|27|qui post me venturus est, cuius ego non sum dignus, ut solvam eius corrigiam calceamenti ".
JOHN|1|28|Haec in Bethania facta sunt trans Iordanem, ubi erat Ioannes baptizans.
JOHN|1|29|Altera die videt Iesum venientem ad se et ait: " Ecce agnus Dei, qui tollit peccatum mundi.
JOHN|1|30|Hic est, de quo dixi: Post me venit vir, qui ante me factus est, quia prior me erat.
JOHN|1|31|Et ego nesciebam eum, sed ut manifestetur Israel, propterea veni ego in aqua baptizans ".
JOHN|1|32|Et testimonium perhibuit Ioannes dicens: " Vidi Spiritum descendentem quasi columbam de caelo, et mansit super eum;
JOHN|1|33|et ego nesciebam eum, sed, qui misit me baptizare in aqua, ille mihi dixit: "Super quem videris Spiritum descendentem et manentem super eum, hic est qui baptizat in Spiritu Sancto".
JOHN|1|34|Et ego vidi et testimonium perhibui quia hic est Filius Dei ".
JOHN|1|35|Altera die iterum stabat Ioannes et ex discipulis eius duo,
JOHN|1|36|et respiciens Iesum ambulantem dicit: " Ecce agnus Dei ".
JOHN|1|37|Et audierunt eum duo discipuli loquentem et secuti sunt Iesum.
JOHN|1|38|Conversus autem Iesus et videns eos sequentes se dicit eis: " Quid quaeritis? ". Qui dixerunt ei: " Rabbi - quod dicitur interpretatum Magister - ubi manes? ".
JOHN|1|39|Dicit eis: " Venite et videbitis ". Venerunt ergo et viderunt, ubi maneret, et apud eum manserunt die illo; hora erat quasi decima.
JOHN|1|40|Erat Andreas, frater Simonis Petri, unus ex duobus, qui audierant ab Ioanne et secuti fuerant eum.
JOHN|1|41|Invenit hic primum fratrem suum Simonem et dicit ei: " Invenimus Messiam " - quod est interpretatum Christus C;
JOHN|1|42|adduxit eum ad Iesum. Intuitus eum Iesus dixit: " Tu es Simon filius Ioannis; tu vocaberis Cephas " - quod interpretatur Petrus C.
JOHN|1|43|In crastinum voluit exire in Galilaeam et invenit Philippum. Et dicit ei Iesus: " Sequere me ".
JOHN|1|44|Erat autem Philippus a Bethsaida, civitate Andreae et Petri.
JOHN|1|45|Invenit Philippus Nathanael et dicit ei: " Quem scripsit Moyses in Lege et Prophetae invenimus, Iesum filium Ioseph a Nazareth ".
JOHN|1|46|Et dixit ei Nathanael: " A Nazareth potest aliquid boni esse? ". Dicit ei Philippus: " Veni et vide ".
JOHN|1|47|Vidit Iesus Nathanael venientem ad se et dicit de eo: " Ecce vere Israelita, in quo dolus non est ".
JOHN|1|48|Dicit ei Nathanael: " Unde me nosti? ". Respondit Iesus et dixit ei: " Priusquam te Philippus vocaret, cum esses sub ficu, vidi te ".
JOHN|1|49|Respondit ei Nathanael: " Rabbi, tu es Filius Dei, tu rex es Israel! ".
JOHN|1|50|Respondit Iesus et dixit ei: " Quia dixi tibi: Vidi te sub ficu, credis? Maiora his videbis ".
JOHN|1|51|Et dicit ei: " Amen, amen dico vobis: Videbitis caelum apertum et angelos Dei ascendentes et descendentes supra Filium hominis ".
JOHN|2|1|Et die tertio nuptiae factae sunt in Cana Galilaeae, et erat mater Iesu ibi;
JOHN|2|2|vocatus est autem et Iesus et discipuli eius ad nuptias.
JOHN|2|3|Et deficiente vino, dicit mater Iesu ad eum: " Vinum non habent ".
JOHN|2|4|Et dicit ei Iesus: " Quid mihi et tibi, mulier? Nondum venit hora mea ".
JOHN|2|5|Dicit mater eius ministris: " Quodcumque dixerit vobis, facite ".
JOHN|2|6|Erant autem ibi lapideae hydriae sex positae secundum purificationem Iudaeorum, capientes singulae metretas binas vel ternas.
JOHN|2|7|Dicit eis Iesus: " Implete hydrias aqua ". Et impleverunt eas usque ad summum.
JOHN|2|8|Et dicit eis: " Haurite nunc et ferte architriclino ". Illi autem tulerunt.
JOHN|2|9|Ut autem gustavit architriclinus aquam vinum factam et non sciebat unde esset, ministri autem sciebant, qui haurierant aquam, vocat sponsum architriclinus
JOHN|2|10|et dicit ei: " Omnis homo primum bonum vinum ponit et, cum inebriati fuerint, id quod deterius est; tu servasti bonum vinum usque adhuc ".
JOHN|2|11|Hoc fecit initium signorum Iesus in Cana Galilaeae et manifestavit gloriam suam, et crediderunt in eum discipuli eius.
JOHN|2|12|Post hoc descendit Capharnaum ipse et mater eius et fratres eius et discipuli eius, et ibi manserunt non multis diebus.
JOHN|2|13|Et prope erat Pascha Iudaeorum, et ascendit Hierosolymam Iesus.
JOHN|2|14|Et invenit in templo vendentes boves et oves et columbas, et nummularios sedentes;
JOHN|2|15|et cum fecisset flagellum de funiculis, omnes eiecit de templo, oves quoque et boves, et nummulariorum effudit aes et mensas subvertit;
JOHN|2|16|et his, qui columbas vendebant, dixit: " Auferte ista hinc! Nolite facere domum Patris mei domum negotiationis ".
JOHN|2|17|Recordati sunt discipuli eius quia scriptum est: " Zelus domus tuae comedit me ".
JOHN|2|18|Responderunt ergo Iudaei et dixerunt ei: " Quod signum ostendis nobis, quia haec facis? ".
JOHN|2|19|Respondit Iesus et dixit eis: " Solvite templum hoc, et in tribus diebus excitabo illud ".
JOHN|2|20|Dixerunt ergo Iudaei: " Quadraginta et sex annis aedificatum est templum hoc, et tu tribus diebus excitabis illud? ".
JOHN|2|21|Ille autem dicebat de templo corporis sui.
JOHN|2|22|Cum ergo resurrexisset a mortuis, recordati sunt discipuli eius quia hoc dicebat, et crediderunt Scripturae et sermoni, quem dixit Iesus.
JOHN|2|23|Cum autem esset Hierosolymis in Pascha, in die festo, multi crediderunt in nomine eius, videntes signa eius, quae faciebat.
JOHN|2|24|Ipse autem Iesus non credebat semetipsum eis, eo quod ipse nosset omnes,
JOHN|2|25|et quia opus ei non erat, ut quis testimonium perhiberet de homine; ipse enim sciebat quid esset in homine.
JOHN|3|1|Erat autem homo ex pharisaeis, Nicodemus nomine, princeps Iudaeorum;
JOHN|3|2|hic venit ad eum nocte et dixit ei: " Rabbi, scimus quia a Deo venisti magister; nemo enim potest haec signa facere, quae tu facis, nisi fuerit Deus cum eo ".
JOHN|3|3|Respondit Iesus et dixit ei: " Amen, amen dico tibi: Nisi quis natus fuerit desuper, non potest videre regnum Dei ".
JOHN|3|4|Dicit ad eum Nicodemus: " Quomodo potest homo nasci, cum senex sit? Numquid potest in ventrem matris suae iterato introire et nasci? ".
JOHN|3|5|Respondit Iesus: " Amen, amen dico tibi: Nisi quis natus fuerit ex aqua et Spiritu, non potest introire in regnum Dei.
JOHN|3|6|Quod natum est ex carne, caro est; et, quod natum est ex Spiritu, spiritus est.
JOHN|3|7|Non mireris quia dixi tibi: Oportet vos nasci denuo.
JOHN|3|8|Spiritus, ubi vult, spirat, et vocem eius audis, sed non scis unde veniat et quo vadat; sic est omnis, qui natus est ex Spiritu ".
JOHN|3|9|Respondit Nicodemus et dixit ei: " Quomodo possunt haec fieri? ".
JOHN|3|10|Respondit Iesus et dixit ei: " Tu es magister Israel et haec ignoras?
JOHN|3|11|Amen, amen dico tibi: Quod scimus, loquimur et, quod vidimus, testamur; et testimonium nostrum non accipitis.
JOHN|3|12|Si terrena dixi vobis, et non creditis, quomodo, si dixero vobis caelestia, credetis?
JOHN|3|13|Et nemo ascendit in caelum, nisi qui descendit de caelo, Filius hominis.
JOHN|3|14|Et sicut Moyses exaltavit serpentem in deserto, ita exaltari oportet Filium hominis,
JOHN|3|15|ut omnis, qui credit, in ipso habeat vitam aeternam ".
JOHN|3|16|Sic enim dilexit Deus mundum, ut Filium suum unigenitum daret, ut omnis, qui credit in eum, non pereat, sed habeat vitam aeternam.
JOHN|3|17|Non enim misit Deus Filium in mundum, ut iudicet mundum, sed ut salvetur mundus per ipsum.
JOHN|3|18|Qui credit in eum, non iudicatur; qui autem non credit, iam iudicatus est, quia non credidit in nomen Unigeniti Filii Dei.
JOHN|3|19|Hoc est autem iudicium: Lux venit in mundum, et dilexerunt homines magis tenebras quam lucem; erant enim eorum mala opera.
JOHN|3|20|Omnis enim, qui mala agit, odit lucem et non venit ad lucem, ut non arguantur opera eius;
JOHN|3|21|qui autem facit veritatem, venit ad lucem, ut manifestentur eius opera, quia in Deo sunt facta.
JOHN|3|22|Post haec venit Iesus et discipuli eius in Iudaeam terram, et illic demorabatur cum eis et baptizabat.
JOHN|3|23|Erat autem et Ioannes baptizans in Enon iuxta Salim, quia aquae multae erant illic, et adveniebant et baptizabantur;
JOHN|3|24|nondum enim missus fuerat in carcerem Ioannes.
JOHN|3|25|Facta est ergo quaestio ex discipulis Ioannis cum Iudaeo de purificatione.
JOHN|3|26|Et venerunt ad Ioannem et dixerunt ei: " Rabbi, qui erat tecum trans Iordanem, cui tu testimonium perhibuisti, ecce hic baptizat, et omnes veniunt ad eum! ".
JOHN|3|27|Respondit Ioannes et dixit: " Non potest homo accipere quidquam, nisi fuerit ei datum de caelo.
JOHN|3|28|Ipsi vos mihi testimonium perhibetis, quod dixerim: Non sum ego Christus, sed: Missus sum ante illum.
JOHN|3|29|Qui habet sponsam, sponsus est; amicus autem sponsi, qui stat et audit eum, gaudio gaudet propter vocem sponsi. Hoc ergo gaudium meum impletum est.
JOHN|3|30|Illum oportet crescere, me autem minui ".
JOHN|3|31|Qui de sursum venit, supra omnes est; qui est de terra, de terra est et de terra loquitur. Qui de caelo venit, supra omnes est;
JOHN|3|32|et quod vidit et audivit, hoc testatur, et testimonium eius nemo accipit.
JOHN|3|33|Qui accipit eius testimonium, signavit quia Deus verax est.
JOHN|3|34|Quem enim misit Deus, verba Dei loquitur; non enim ad mensuram dat Spiritum.
JOHN|3|35|Pater diligit Filium et omnia dedit in manu eius.
JOHN|3|36|Qui credit in Filium, habet vitam aeternam; qui autem incredulus est Filio, non videbit vitam, sed ira Dei manet super eum.
JOHN|4|1|Ut ergo cognovit Iesus quia audierunt pharisaei quia Iesus plures discipulos facit et baptizat quam Ioannes
JOHN|4|2|- quamquam Iesus ipse non baptizaret sed discipuli eius -
JOHN|4|3|reliquit Iudaeam et abiit iterum in Galilaeam.
JOHN|4|4|Oportebat autem eum transire per Samariam.
JOHN|4|5|Venit ergo in civitatem Samariae, quae dicitur Sichar, iuxta praedium, quod dedit Iacob Ioseph filio suo;
JOHN|4|6|erat autem ibi fons Iacob. Iesus ergo fatigatus ex itinere sedebat sic super fontem; hora erat quasi sexta.
JOHN|4|7|Venit mulier de Samaria haurire aquam. Dicit ei Iesus: " Da mihi bibere;
JOHN|4|8|discipuli enim eius abierant in civitatem, ut cibos emerent.
JOHN|4|9|Dicit ergo ei mulier illa Samaritana: " Quomodo tu, Iudaeus cum sis, bibere a me poscis, quae sum mulier Samaritana? ". Non enim coutuntur Iudaei Samaritanis.
JOHN|4|10|Respondit Iesus et dixit ei: " Si scires donum Dei, et quis est, qui dicit tibi: "Da mihi bibere", tu forsitan petisses ab eo, et dedisset tibi aquam vivam ".
JOHN|4|11|Dicit ei mulier: " Domine, neque in quo haurias habes, et puteus altus est; unde ergo habes aquam vivam?
JOHN|4|12|Numquid tu maior es patre nostro Iacob, qui dedit nobis puteum, et ipse ex eo bibit et filii eius et pecora eius? ".
JOHN|4|13|Respondit Iesus et dixit ei: " Omnis, qui bibit ex aqua hac, sitiet iterum;
JOHN|4|14|qui autem biberit ex aqua, quam ego dabo ei, non sitiet in aeternum; sed aqua, quam dabo ei, fiet in eo fons aquae salientis in vitam aeternam.
JOHN|4|15|Dicit ad eum mulier: " Domine, da mihi hanc aquam, ut non sitiam neque veniam huc haurire ".
JOHN|4|16|Dicit ei: " Vade, voca virum tuum et veni huc ".
JOHN|4|17|Respondit mulier et dixit ei: " Non habeo virum ". Dicit ei Iesus: " Bene dixisti: "Non habeo virum";
JOHN|4|18|quinque enim viros habuisti, et nunc, quem habes, non est tuus vir. Hoc vere dixisti ".
JOHN|4|19|Dicit ei mulier: " Domine, video quia propheta es tu.
JOHN|4|20|Patres nostri in monte hoc adoraverunt, et vos dicitis quia in Hierosolymis est locus, ubi adorare oportet ".
JOHN|4|21|Dicit ei Iesus: " Crede mihi, mulier, quia venit hora, quando neque in monte hoc neque in Hierosolymis adorabitis Patrem.
JOHN|4|22|Vos adoratis, quod nescitis; nos adoramus, quod scimus, quia salus ex Iudaeis est.
JOHN|4|23|Sed venit hora, et nunc est, quando veri adoratores adorabunt Patrem in Spiritu et veritate; nam et Pater tales quaerit, qui adorent eum.
JOHN|4|24|Spiritus est Deus, et eos, qui adorant eum, in Spiritu et veritate oportet adorare ".
JOHN|4|25|Dicit ei mulier: " Scio quia Messias venit - qui dicitur Christus C; cum venerit ille, nobis annuntiabit omnia ".
JOHN|4|26|Dicit ei Iesus: " Ego sum, qui loquor tecum ".
JOHN|4|27|Et continuo venerunt discipuli eius et mirabantur quia cum muliere loquebatur; nemo tamen dixit: " Quid quaeris aut quid loqueris cum ea? ".
JOHN|4|28|Reliquit ergo hydriam suam mulier et abiit in civitatem et dicit illis hominibus:
JOHN|4|29|" Venite, videte hominem, qui dixit mihi omnia, quaecumque feci; numquid ipse est Christus? ".
JOHN|4|30|Exierunt de civitate et veniebant ad eum.
JOHN|4|31|Interea rogabant eum discipuli dicentes: " Rabbi, manduca ".
JOHN|4|32|Ille autem dixit eis: " Ego cibum habeo manducare, quem vos nescitis ".
JOHN|4|33|Dicebant ergo discipuli ad invicem: " Numquid aliquis attulit ei manducare? ".
JOHN|4|34|Dicit eis Iesus: " Meus cibus est, ut faciam voluntatem eius, qui misit me, et ut perficiam opus eius.
JOHN|4|35|Nonne vos dicitis: "Adhuc quattuor menses sunt, et messis venit"? Ecce dico vobis: Levate oculos vestros et videte regiones, quia albae sunt ad messem! Iam
JOHN|4|36|qui metit, mercedem accipit et congregat fructum in vitam aeternam, ut et qui seminat, simul gaudeat et qui metit.
JOHN|4|37|In hoc enim est verbum verum: Alius est qui seminat, et alius est qui metit.
JOHN|4|38|Ego misi vos metere, quod vos non laborastis; alii laboraverunt, et vos in laborem eorum introistis ".
JOHN|4|39|Ex civitate autem illa multi crediderunt in eum Samaritanorum propter verbum mulieris testimonium perhibentis: " Dixit mihi omnia, quaecumque feci! ".
JOHN|4|40|Cum venissent ergo ad illum Samaritani, rogaverunt eum, ut apud ipsos maneret; et mansit ibi duos dies.
JOHN|4|41|Et multo plures crediderunt propter sermonem eius;
JOHN|4|42|et mulieri dicebant: " Iam non propter tuam loquelam credimus; ipsi enim audivimus et scimus quia hic est vere Salvator mundi! ".
JOHN|4|43|Post duos autem dies exiit inde in Galilaeam;
JOHN|4|44|ipse enim Iesus testimonium perhibuit, quia propheta in sua patria honorem non habet.
JOHN|4|45|Cum ergo venisset in Galilaeam, exceperunt eum Galilaei, cum omnia vidissent, quae fecerat Hierosolymis in die festo; et ipsi enim venerant in diem festum.
JOHN|4|46|Venit ergo iterum in Cana Galilaeae, ubi fecit aquam vinum. Et erat quidam regius, cuius filius infirmabatur Capharnaum;
JOHN|4|47|hic, cum audisset quia Iesus advenerit a Iudaea in Galilaeam, abiit ad eum et rogabat, ut descenderet et sanaret filium eius; incipiebat enim mori.
JOHN|4|48|Dixit ergo Iesus ad eum: " Nisi signa et prodigia videritis, non credetis ".
JOHN|4|49|Dicit ad eum regius: " Domine, descende priusquam moriatur puer meus ".
JOHN|4|50|Dicit ei Iesus: " Vade. Filius tuus vivit ". Credidit homo sermoni, quem dixit ei Iesus, et ibat.
JOHN|4|51|Iam autem eo descendente, servi eius occurrerunt ei dicentes quia puer eius vivit.
JOHN|4|52|Interrogabat ergo horam ab eis, in qua melius habuerit. Dixerunt ergo ei: " Heri hora septima reliquit eum febris ".
JOHN|4|53|Cognovit ergo pater quia illa hora erat, in qua dixit ei Iesus: " Filius tuus vivit ", et credidit ipse et domus eius tota.
JOHN|4|54|Hoc iterum secundum signum fecit Iesus, cum venisset a Iudaea in Galilaeam.
JOHN|5|1|Post haec erat dies festus Iu daeorum, et ascendit Iesus Hie rosolymam.
JOHN|5|2|Est autem Hierosolymis, super Probatica, piscina, quae cognominatur HebraiceBethsatha, quinque porticus habens.
JOHN|5|3|In his iacebat multitudo languentium, caecorum, claudorum, aridorum.
JOHN|5|4|()
JOHN|5|5|Erat autem quidam homo ibi triginta et octo annos habens in infirmitate sua.
JOHN|5|6|Hunc cum vidisset Iesus iacentem, et cognovisset quia multum iam tempus habet, dicit ei: " Vis sanus fieri? ".
JOHN|5|7|Respondit ei languidus: " Domine, hominem non habeo, ut, cum turbata fuerit aqua, mittat me in piscinam; dum autem venio ego, alius ante me descendit ".
JOHN|5|8|Dicit ei Iesus: " Surge, tolle grabatum tuum et ambula ".
JOHN|5|9|Et statim sanus factus est homo et sustulit grabatum suum et ambulabat.Erat autem sabbatum in illo die.
JOHN|5|10|Dicebant ergo Iudaei illi, qui sanatus fuerat: " Sabbatum est, et non licet tibi tollere grabatum tuum ".
JOHN|5|11|Ille autem respondit eis: " Qui me fecit sanum, ille mihi dixit: "Tolle grabatum tuum et ambula" ".
JOHN|5|12|Interrogaverunt eum: " Quis est ille homo, qui dixit tibi: "Tolle et ambula"? ".
JOHN|5|13|Is autem, qui sanus fuerat effectus, nesciebat quis esset; Iesus enim declinavit a turba constituta in loco.
JOHN|5|14|Postea invenit eum Iesus in templo et dixit illi: " Ecce sanus factus es; iam noli peccare, ne deterius tibi aliquid contingat ".
JOHN|5|15|Abiit ille homo et nuntiavit Iudaeis quia Iesus esset, qui fecit eum sanum.
JOHN|5|16|Et propterea persequebantur Iudaei Iesum, quia haec faciebat in sabbato.
JOHN|5|17|Iesus autem respondit eis: " Pater meus usque modo operatur, et ego operor ".
JOHN|5|18|Propterea ergo magis quaerebant eum Iudaei interficere, quia non solum solvebat sabbatum, sed et Patrem suum dicebat Deum, aequalem se faciens Deo.
JOHN|5|19|Respondit itaque Iesus et dixit eis: " Amen, amen dico vobis: Non potest Filius a se facere quidquam, nisi quod viderit Patrem facientem; quaecumque enim ille faciat, haec et Filius similiter facit.
JOHN|5|20|Pater enim diligit Filium et omnia demonstrat ei, quae ipse facit, et maiora his demonstrabit ei opera, ut vos miremini.
JOHN|5|21|Sicut enim Pater suscitat mortuos et vivificat, sic et Filius, quos vult, vivificat.
JOHN|5|22|Neque enim Pater iudicat quemquam, sed iudicium omne dedit Filio,
JOHN|5|23|ut omnes honorificent Filium, sicut honorificant Patrem. Qui non honorificat Filium, non honorificat Patrem, qui misit illum.
JOHN|5|24|Amen, amen dico vobis: Qui verbum meum audit et credit ei, qui misit me, habet vitam aeternam et in iudicium non venit, sed transiit a morte in vitam.
JOHN|5|25|Amen, amen dico vobis: Venit hora, et nunc est, quando mortui audient vocem Filii Dei et, qui audierint, vivent.
JOHN|5|26|Sicut enim Pater habet vitam in semetipso, sic dedit et Filio vitam habere in semetipso;
JOHN|5|27|et potestatem dedit ei iudicium facere, quia Filius hominis est.
JOHN|5|28|Nolite mirari hoc, quia venit hora, in qua omnes, qui in monumentis sunt, audient vocem eius;
JOHN|5|29|et procedent, qui bona fecerunt, in resurrectionem vitae, qui vero mala egerunt, in resurrectionem iudicii.
JOHN|5|30|Non possum ego a meipso facere quidquam; sicut audio, iudico, et iudicium meum iustum est, quia non quaero voluntatem meam, sed voluntatem eius, qui misit me.
JOHN|5|31|Si ego testimonium perhibeo de meipso, testimonium meum non est verum;
JOHN|5|32|alius est, qui testimonium perhibet de me, et scio quia verum est testimonium, quod perhibet de me.
JOHN|5|33|Vos misistis ad Ioannem, et testimonium perhibuit veritati;
JOHN|5|34|ego autem non ab homine testimonium accipio, sed haec dico, ut vos salvi sitis.
JOHN|5|35|Ille erat lucerna ardens et lucens; vos autem voluistis exsultare ad horam in luce eius.
JOHN|5|36|Ego autem habeo testimonium maius Ioanne; opera enim, quae dedit mihi Pater, ut perficiam ea, ipsa opera, quae ego facio, testimonium perhibent de me, quia Pater me misit;
JOHN|5|37|et, qui misit me, Pater, ipse testimonium perhibuit de me. Neque vocem eius umquam audistis neque speciem eius vidistis;
JOHN|5|38|et verbum eius non habetis in vobis manens, quia, quem misit ille, huic vos non creditis.
JOHN|5|39|Scrutamini Scripturas, quia vos putatis in ipsis vitam aeternam habere; et illae sunt, quae testimonium perhibent de me.
JOHN|5|40|Et non vultis venire ad me, ut vitam habeatis.
JOHN|5|41|Gloriam ab hominibus non accipio,
JOHN|5|42|sed cognovi vos, quia dilectionem Dei non habetis in vobis.
JOHN|5|43|Ego veni in nomine Patris mei, et non accipitis me; si alius venerit in nomine suo, illum accipietis.
JOHN|5|44|Quomodo potestis vos credere, qui gloriam ab invicem accipitis, et gloriam, quae a solo est Deo, non quaeritis?
JOHN|5|45|Nolite putare quia ego accusaturus sim vos apud Patrem; est qui accuset vos: Moyses, in quo vos speratis.
JOHN|5|46|Si enim crederetis Moysi, crederetis forsitan et mihi; de me enim ille scripsit.
JOHN|5|47|Si autem illius litteris non creditis, quomodo meis verbis credetis? ".
JOHN|6|1|Post haec abiit Iesus trans mare Galilaeae, quod est Tiberiadis.
JOHN|6|2|Et sequebatur eum multitudo magna, quia videbant signa, quae faciebat super his, qui infirmabantur.
JOHN|6|3|Subiit autem in montem Iesus et ibi sedebat cum discipulis suis.
JOHN|6|4|Erat autem proximum Pascha, dies festus Iudaeorum.
JOHN|6|5|Cum sublevasset ergo oculos Iesus et vidisset quia multitudo magna venit ad eum, dicit ad Philippum: " Unde ememus panes, ut manducent hi? ".
JOHN|6|6|Hoc autem dicebat tentans eum; ipse enim sciebat quid esset facturus.
JOHN|6|7|Respondit ei Philippus: " Ducentorum denariorum panes non sufficiunt eis, ut unusquisque modicum quid accipiat! ".
JOHN|6|8|Dicit ei unus ex discipulis eius, Andreas frater Simonis Petri:
JOHN|6|9|" Est puer hic, qui habet quinque panes hordeaceos et duos pisces; sed haec quid sunt propter tantos? ".
JOHN|6|10|Dixit Iesus: " Facite homines discumbere ". Erat autem fenum multum in loco. Discubuerunt ergo viri numero quasi quinque milia.
JOHN|6|11|Accepit ergo panes Iesus et, cum gratias egisset, distribuit discumbentibus; similiter et ex piscibus, quantum volebant.
JOHN|6|12|Ut autem impleti sunt, dicit discipulis suis: " Colligite, quae superaverunt, fragmenta, ne quid pereat ".
JOHN|6|13|Collegerunt ergo et impleverunt duodecim cophinos fragmentorum ex quinque panibus hordeaceis, quae superfuerunt his, qui manducaverunt.
JOHN|6|14|Illi ergo homines, cum vidissent quod fecerat signum, dicebant: " Hic est vere propheta, qui venit in mundum! ".
JOHN|6|15|Iesus ergo, cum cognovisset quia venturi essent, ut raperent eum et facerent eum regem, secessit iterum in montem ipse solus.
JOHN|6|16|Ut autem sero factum est, descenderunt discipuli eius ad mare
JOHN|6|17|et, cum ascendissent navem, veniebant trans mare in Capharnaum. Et tenebrae iam factae erant, et nondum venerat ad eos Iesus.
JOHN|6|18|Mare autem, vento magno flante, exsurgebat.
JOHN|6|19|Cum remigassent ergo quasi stadia viginti quinque aut triginta, vident Iesum ambulantem super mare et proximum navi fieri, et timuerunt.
JOHN|6|20|Ille autem dicit eis: " Ego sum, nolite timere! ".
JOHN|6|21|Volebant ergo accipere eum in navem, et statim fuit navis ad terram, in quam ibant.
JOHN|6|22|Altera die turba, quae stabat trans mare, vidit quia navicula alia non erat ibi, nisi una, et quia non introisset cum discipulis suis Iesus in navem, sed soli discipuli eius abiissent;
JOHN|6|23|aliae supervenerunt naves a Tiberiade iuxta locum, ubi manducaverant panem, gratias agente Domino.
JOHN|6|24|Cum ergo vidisset turba quia Iesus non esset ibi neque discipuli eius, ascenderunt ipsi naviculas et venerunt Capharnaum quaerentes Iesum.
JOHN|6|25|Et cum invenissent eum trans mare, dixerunt ei: " Rabbi, quando huc venisti? ".
JOHN|6|26|Respondit eis Iesus et dixit: " Amen, amen dico vobis: Quaeritis me, non quia vidistis signa, sed quia manducastis ex panibus et saturati estis.
JOHN|6|27|Operamini non cibum, qui perit, sed cibum, qui permanet in vitam aeternam, quem Filius hominis vobis dabit; hunc enim Pater signavit Deus!.
JOHN|6|28|Dixerunt ergo ad eum: " Quid faciemus, ut operemur opera Dei? ".
JOHN|6|29|Respondit Iesus et dixit eis: " Hoc est opus Dei, ut credatis in eum, quem misit ille ".
JOHN|6|30|Dixerunt ergo ei: " Quod ergo tu facis signum, ut videamus et credamus tibi? Quid operaris?
JOHN|6|31|Patres nostri manna manducaverunt in deserto, sicut scriptum est: Panem de caelo dedit eis manducare" ".
JOHN|6|32|Dixit ergo eis Iesus: " Amen, amen dico vobis: Non Moyses dedit vobis panem de caelo, sed Pater meus dat vobis panem de caelo verum;
JOHN|6|33|panis enim Dei est, qui descendit de caelo et dat vitam mundo ".
JOHN|6|34|Dixerunt ergo ad eum: " Domine, semper da nobis panem hunc ".
JOHN|6|35|Dixit eis Iesus: " Ego sum panis vitae. Qui venit ad me, non esuriet; et, qui credit in me, non sitiet umquam.
JOHN|6|36|Sed dixi vobis, quia et vidistis me et non creditis.
JOHN|6|37|Omne, quod dat mihi Pater, ad me veniet; et eum, qui venit ad me, non eiciam foras,
JOHN|6|38|quia descendi de caelo, non ut faciam voluntatem meam sed voluntatem eius, qui misit me.
JOHN|6|39|Haec est autem voluntas eius, qui misit me, ut omne, quod dedit mihi, non perdam ex eo, sed resuscitem illud in novissimo die.
JOHN|6|40|Haec est enim voluntas Patris mei, ut omnis, qui videt Filium et credit in eum, habeat vitam aeternam; et resuscitabo ego eum in novissimo die ".
JOHN|6|41|Murmurabant ergo Iudaei de illo, quia dixisset: " Ego sum panis, qui de caelo descendi ",
JOHN|6|42|et dicebant: " Nonne hic est Iesus filius Ioseph, cuius nos novimus patrem et matrem? Quomodo dicit nunc: "De caelo descendi"? ".
JOHN|6|43|Respondit Iesus et dixit eis: " Nolite murmurare in invicem.
JOHN|6|44|Nemo potest venire ad me, nisi Pater, qui misit me, traxerit eum; et ego resuscitabo eum in novissimo die.
JOHN|6|45|Est scriptum in Prophetis: "Et erunt omnes docibiles Dei ". Omnis, qui audivit a Patre et didicit, venit ad me.
JOHN|6|46|Non quia Patrem vidit quisquam, nisi is qui est a Deo, hic vidit Patrem.
JOHN|6|47|Amen, amen dico vobis: Qui credit, habet vitam aeternam.
JOHN|6|48|Ego sum panis vitae.
JOHN|6|49|Patres vestri manducaverunt in deserto manna et mortui sunt.
JOHN|6|50|Hic est panis de caelo descendens, ut, si quis ex ipso manducaverit, non moriatur.
JOHN|6|51|Ego sum panis vivus, qui de caelo descendi. Si quis manducaverit ex hoc pane, vivet in aeternum; panis autem, quem ego dabo, caro mea est pro mundi vita ".
JOHN|6|52|Litigabant ergo Iudaei ad invicem dicentes: " Quomodo potest hic nobis carnem suam dare ad manducandum? ".
JOHN|6|53|Dixit ergo eis Iesus: " Amen, amen dico vobis: Nisi manducaveritis carnem Filii hominis et biberitis eius sanguinem, non habetis vitam in vobismetipsis.
JOHN|6|54|Qui manducat meam carnem et bibit meum sanguinem, habet vitam aeternam; et ego resuscitabo eum in novissimo die.
JOHN|6|55|Caro enim mea verus est cibus, et sanguis meus verus est potus.
JOHN|6|56|Qui manducat meam carnem et bibit meum sanguinem, in me manet, et ego in illo.
JOHN|6|57|Sicut misit me vivens Pater, et ego vivo propter Patrem; et, qui manducat me, et ipse vivet propter me.
JOHN|6|58|Hic est panis, qui de caelo descendit, non sicut manducaverunt patres et mortui sunt; qui manducat hunc panem, vivet in aeternum ".
JOHN|6|59|Haec dixit in synagoga docens in Capharnaum.
JOHN|6|60|Multi ergo audientes ex discipulis eius dixerunt: " Durus est hic sermo! Quis potest eum audire? ".
JOHN|6|61|Sciens autem Iesus apud semetipsum quia murmurarent de hoc discipuli eius, dixit eis: " Hoc vos scandalizat?
JOHN|6|62|Si ergo videritis Filium hominis ascendentem, ubi erat prius?
JOHN|6|63|Spiritus est, qui vivificat, caro non prodest quidquam; verba, quae ego locutus sum vobis, Spiritus sunt et vita sunt.
JOHN|6|64|Sed sunt quidam ex vobis, qui non credunt ". Sciebat enim ab initio Iesus, qui essent non credentes, et quis traditurus esset eum.
JOHN|6|65|Et dicebat: " Propterea dixi vobis: Nemo potest venire ad me, nisi fuerit ei datum a Patre ".
JOHN|6|66|Ex hoc multi discipulorum eius abierunt retro et iam non cum illo ambulabant.
JOHN|6|67|Dixit ergo Iesus ad Duodecim: " Numquid et vos vultis abire? ".
JOHN|6|68|Respondit ei Simon Petrus: " Domine, ad quem ibimus? Verba vitae aeternae habes;
JOHN|6|69|et nos credidimus et cognovimus quia tu es Sanctus Dei ".
JOHN|6|70|Respondit eis Iesus: " Nonne ego vos Duodecim elegi? Et ex vobis unus Diabolus est ".
JOHN|6|71|Dicebat autem Iudam Simonis Iscariotis; hic enim erat traditurus eum, cum esset unus ex Duodecim.
JOHN|7|1|Et post haec ambulabat Iesus in Galilaeam; non enim volebat in Iudaeam ambulare, quia quaerebant eum Iudaei interficere.
JOHN|7|2|Erat autem in proximo dies festus Iudaeorum, Scenopegia.
JOHN|7|3|Dixerunt ergo ad eum fratres eius: " Transi hinc et vade in Iudaeam, ut et discipuli tui videant opera tua, quae facis.
JOHN|7|4|Nemo quippe in occulto quid facit et quaerit ipse in palam esse. Si haec facis, manifesta teipsum mundo ".
JOHN|7|5|Neque enim fratres eius credebant in eum.
JOHN|7|6|Dicit ergo eis Iesus: " Tempus meum nondum adest, tempus autem vestrum semer est paratum.
JOHN|7|7|Non potest mundus odisse vos; me autem odit, quia ego testimonium perhibeo de illo, quia opera eius mala sunt.
JOHN|7|8|Vos ascendite ad diem festum; ego non ascendo ad diem festum istum, quia meum tempus nondum impletum est ".
JOHN|7|9|Haec autem cum dixisset, ipse mansit in Galilaea.
JOHN|7|10|Ut autem ascenderunt fratres eius ad diem festum, tunc et ipse ascendit, non manifeste sed quasi in occulto.
JOHN|7|11|Iudaei ergo quaerebant eum in die festo et dicebant: " Ubi est ille? ".
JOHN|7|12|Et murmur multus de eo erat in turba. Alii quidem dicebant: " Bonus est! "; alii autem dicebant: " Non, sed seducit turbam! ".
JOHN|7|13|Nemo tamen palam loquebatur de illo propter metum Iudaeorum.
JOHN|7|14|Iam autem die festo mediante, ascendit Iesus in templum et docebat.
JOHN|7|15|Mirabantur ergo Iudaei dicentes: " Quomodo hic litteras scit, cum non didicerit? ".
JOHN|7|16|Respondit ergo eis Iesus et dixit: " Mea doctrina non est mea sed eius, qui misit me.
JOHN|7|17|Si quis voluerit voluntatem eius facere, cognoscet de doctrina utrum ex Deo sit, an ego a meipso loquar.
JOHN|7|18|Qui a semetipso loquitur, gloriam propriam quaerit; qui autem quaerit gloriam eius, qui misit illum, hic verax est, et iniustitia in illo non est.
JOHN|7|19|Nonne Moyses dedit vobis legem? Et nemo ex vobis facit legem. Quid me quaeritis interficere? ".
JOHN|7|20|Respondit turba: " Daemonium habes! Quis te quaerit interficere? ".
JOHN|7|21|Respondit Iesus et dixit eis: " Unum opus feci, et omnes miramini.
JOHN|7|22|Propterea Moyses dedit vobis circumcisionem - non quia ex Moyse est sed ex patribus - et in sabbato circumciditis hominem.
JOHN|7|23|Si circumcisionem accipit homo in sabbato, ut non solvatur lex Moysis, mihi indignamini, quia totum hominem sanum feci in sabbato?
JOHN|7|24|Nolite iudicare secundum faciem, sed iustum iudicium iudicate ".
JOHN|7|25|Dicebant ergo quidam ex Hierosolymitis: " Nonne hic est, quem quaerunt interficere?
JOHN|7|26|Et ecce palam loquitur, et nihil ei dicunt. Numquid vere cognoverunt principes quia hic est Christus?
JOHN|7|27|Sed hunc scimus unde sit, Christus autem cum venerit, nemo scit unde sit ".
JOHN|7|28|Clamavit ergo docens in templo Iesus et dicens: " Et me scitis et unde sim scitis. Et a meipso non veni, sed est verus, qui misit me, quem vos non scitis.
JOHN|7|29|Ego scio eum, quia ab ipso sum, et ipse me misit ".
JOHN|7|30|Quaerebant ergo eum apprehendere, et nemo misit in illum manus, quia nondum venerat hora eius.
JOHN|7|31|De turba autem multi crediderunt in eum et dicebant: " Christus cum venerit, numquid plura signa faciet quam quae hic fecit? ".
JOHN|7|32|Audierunt pharisaei turbam murmurantem de illo haec et miserunt pontifices et pharisaei ministros, ut apprehenderent eum.
JOHN|7|33|Dixit ergo Iesus: " Adhuc modicum tempus vobiscum sum et vado ad eum, qui misit me.
JOHN|7|34|Quaeretis me et non invenietis; et ubi sum ego, vos non potestis venire.
JOHN|7|35|Dixerunt ergo Iudaei ad seipsos: " Quo hic iturus est, quia nos non inveniemus eum? Numquid in dispersionem Graecorum iturus est et docturus Graecos?
JOHN|7|36|Quis est hic sermo, quem dixit: "Quaeretis me et non invenietis" et: Ubi sum ego, vos non potestis venire"? ".
JOHN|7|37|In novissimo autem die magno festivitatis stabat Iesus et clamavit dicens: " Si quis sitit, veniat ad me et bibat,
JOHN|7|38|qui credit in me. Sicut dixit Scriptura, flumina de ventre eius fluent aquae vivae ".
JOHN|7|39|Hoc autem dixit de Spiritu, quem accepturi erant qui crediderant in eum. Nondum enim erat Spiritus, quia Iesus nondum fuerat glorificatus.
JOHN|7|40|Ex illa ergo turba, cum audissent hos sermones, dicebant: " Hic est vere propheta! ";
JOHN|7|41|alii dicebant: " Hic est Christus! "; quidam autem dicebant: " Numquid a Galilaea Christus venit?
JOHN|7|42|Nonne Scriptura dixit: "Ex semine David et de Bethlehem castello, ubi erat David, venit Christus"? ".
JOHN|7|43|Dissensio itaque facta est in turba propter eum.
JOHN|7|44|Quidam autem ex ipsis volebant apprehendere eum, sed nemo misit super illum manus.
JOHN|7|45|Venerunt ergo ministri ad pontifices et pharisaeos; et dixerunt eis illi: " Quare non adduxistis eum? ".
JOHN|7|46|Responderunt ministri: " Numquam sic locutus est homo ".
JOHN|7|47|Responderunt ergo eis pharisaei: " Numquid et vos seducti estis?
JOHN|7|48|Numquid aliquis ex principibus credidit in eum aut ex pharisaeis?
JOHN|7|49|Sed turba haec, quae non novit legem, maledicti sunt! ".
JOHN|7|50|Dicit Nicodemus ad eos, ille qui venit ad eum antea, qui unus erat ex ipsis:
JOHN|7|51|" Numquid lex nostra iudicat hominem, nisi audierit ab ipso prius et cognoverit quid faciat? ".
JOHN|7|52|Responderunt et dixerunt ei: " Numquid et tu ex Galilaea es? Scrutare et vide quia propheta a Galilaea non surgit! ".
JOHN|7|53|Et reversi sunt unusquisque in domum suam.
JOHN|8|1|Iesus autem perrexit in montem Oliveti.
JOHN|8|2|Diluculo autem iterum venit in templum, et omnis populus veniebat ad eum, et sedens docebat eos.
JOHN|8|3|Adducunt autem scribae et pharisaei mulierem in adulterio deprehensam et statuerunt eam in medio
JOHN|8|4|et dicunt ei: " Magister, haec mulier manifesto deprehensa est in adulterio.
JOHN|8|5|In lege autem Moyses mandavit nobis huiusmodi lapidare; tu ergo quid dicis? ".
JOHN|8|6|Hoc autem dicebant tentantes eum, ut possent accusare eum. Iesus autem inclinans se deorsum digito scribebat in terra.
JOHN|8|7|Cum autem perseverarent interrogantes eum, erexit se et dixit eis: " Qui sine peccato est vestrum, primus in illam lapidem mittat ";
JOHN|8|8|et iterum se inclinans scribebat in terra.
JOHN|8|9|Audientes autem unus post unum exibant, incipientes a senioribus, et remansit solus, et mulier in medio stans.
JOHN|8|10|Erigens autem se Iesus dixit ei: " Mulier, ubi sunt? Nemo te condemnavit? ".
JOHN|8|11|Quae dixit: " Nemo, Domine ". Dixit autem Iesus: " Nec ego te condemno; vade et amplius iam noli peccare ".
JOHN|8|12|Iterum ergo locutus est eis Iesus dicens: " Ego sum lux mundi; qui sequitur me, non ambulabit in tenebris, sed habebit lucem vitae ".
JOHN|8|13|Dixerunt ergo ei pharisaei: " Tu de teipso testimonium perhibes; testimonium tuum non est verum ".
JOHN|8|14|Respondit Iesus et dixit eis: " Et si ego testimonium perhibeo de meipso, verum est testimonium meum, quia scio unde veni et quo vado; vos autem nescitis unde venio aut quo vado.
JOHN|8|15|Vos secundum carnem iudicatis, ego non iudico quemquam.
JOHN|8|16|Et si iudico ego, iudicium meum verum est, quia solus non sum, sed ego et, qui me misit, Pater.
JOHN|8|17|Sed et in lege vestra scriptum est, quia duorum hominum testimonium verum est.
JOHN|8|18|Ego sum, qui testimonium perhibeo de meipso, et testimonium perhibet de me, qui misit me, Pater ".
JOHN|8|19|Dicebant ergo ei: " Ubi est Pater tuus? ". Respondit Iesus: " Neque me scitis neque Patrem meum; si me sciretis, forsitan et Patrem meum sciretis.
JOHN|8|20|Haec verba locutus est in gazophylacio docens in templo; et nemo apprehendit eum, quia necdum venerat hora eius.
JOHN|8|21|Dixit ergo iterum eis: " Ego vado, et quaeretis me et in peccato vestro moriemini! Quo ego vado, vos non potestis venire ".
JOHN|8|22|Dicebant ergo Iudaei: " Numquid interficiet semetipsum, quia dicit: Quo ego vado, vos non potestis venire"? ".
JOHN|8|23|Et dicebat eis: " Vos de deorsum estis, ego de supernis sum; vos de mundo hoc estis, ego non sum de hoc mundo.
JOHN|8|24|Dixi ergo vobis quia moriemini in peccatis vestris; si enim non credideritis quia ego sum, moriemini in peccatis vestris ".
JOHN|8|25|Dicebant ergo ei: " Tu quis es? ". Dixit eis Iesus: " In principio: id quod et loquor vobis!
JOHN|8|26|Multa habeo de vobis loqui et iudicare; sed, qui misit me, verax est, et ego, quae audivi ab eo, haec loquor ad mundum ".
JOHN|8|27|Non cognoverunt quia Patrem eis dicebat.
JOHN|8|28|Dixit ergo eis Iesus: " Cum exaltaveritis Filium hominis, tunc cognoscetis quia ego sum et a meipso facio nihil, sed, sicut docuit me Pater, haec loquor.
JOHN|8|29|Et qui me misit, mecum est; non reliquit me solum, quia ego, quae placita sunt ei, facio semper ".
JOHN|8|30|Haec illo loquente, multi crediderunt in eum.
JOHN|8|31|Dicebat ergo Iesus ad eos, qui crediderunt ei, Iudaeos: " Si vos manseritis in sermone meo, vere discipuli mei estis
JOHN|8|32|et cognoscetis veritatem, et veritas liberabit vos ".
JOHN|8|33|Responderunt ei: " Semen Abrahae sumus et nemini servivimus umquam! Quomodo tu dicis: "Liberi fietis"? ".
JOHN|8|34|Respondit eis Iesus: " Amen, amen dico vobis: Omnis, qui facit peccatum, servus est peccati.
JOHN|8|35|Servus autem non manet in domo in aeternum; filius manet in aeternum.
JOHN|8|36|Si ergo Filius vos liberaverit, vere liberi eritis.
JOHN|8|37|Scio quia semen Abrahae estis; sed quaeritis me interficere, quia sermo meus non capit in vobis.
JOHN|8|38|Ego, quae vidi apud Patrem, loquor; et vos ergo, quae audivistis a patre, facitis ".
JOHN|8|39|Responderunt et dixerunt ei: " Pater noster Abraham est ". Dicit eis Iesus: " Si filii Abrahae essetis, opera Abrahae faceretis.
JOHN|8|40|Nunc autem quaeritis me interficere, hominem, qui veritatem vobis locutus sum, quam audivi a Deo; hoc Abraham non fecit.
JOHN|8|41|Vos facitis opera patris vestri ". Dixerunt itaque ei: " Nos ex fornicatione non sumus nati; unum patrem habemus Deum! ".
JOHN|8|42|Dixit eis Iesus: " Si Deus pater vester esset, diligeretis me; ego enim ex Deo processi et veni; neque enim a meipso veni, sed ille me misit.
JOHN|8|43|Quare loquelam meam non cognoscitis? Quia non potestis audire sermonem meum.
JOHN|8|44|Vos ex patre Diabolo estis et desideria patris vestri vultis facere. Ille homicida erat ab initio et in veritate non stabat, quia non est veritas in eo. Cum loquitur mendacium, ex propriis loquitur, quia mendax est et pater eius.
JOHN|8|45|Ego autem quia veritatem dico, non creditis mihi.
JOHN|8|46|Quis ex vobis arguit me de peccato? Si veritatem dico, quare vos non creditis mihi?
JOHN|8|47|Qui est ex Deo, verba Dei audit; propterea vos non auditis, quia ex Deo non estis ".
JOHN|8|48|Responderunt Iudaei et dixerunt ei: " Nonne bene dicimus nos, quia Samaritanus es tu et daemonium habes? ".
JOHN|8|49|Respondit Iesus: " Ego daemonium non habeo, sed honorifico Patrem meum, et vos inhonoratis me.
JOHN|8|50|Ego autem non quaero gloriam meam; est qui quaerit et iudicat.
JOHN|8|51|Amen, amen dico vobis: Si quis sermonem meum servaverit, mortem non videbit in aeternum ".
JOHN|8|52|Dixerunt ergo ei Iudaei: " Nunc cognovimus quia daemonium habes. Abraham mortuus est et prophetae, et tu dicis: "Si quis sermonem meum servaverit, non gustabit mortem in aeternum".
JOHN|8|53|Numquid tu maior es patre nostro Abraham, qui mortuus est? Et prophetae mortui sunt! Quem teipsum facis? ".
JOHN|8|54|Respondit Iesus: " Si ego glorifico meipsum, gloria mea nihil est; est Pater meus, qui glorificat me, quem vos dicitis: "Deus noster est!",
JOHN|8|55|et non cognovistis eum. Ego autem novi eum. Et si dixero: Non scio eum, ero similis vobis, mendax; sed scio eum et sermonem eius servo.
JOHN|8|56|Abraham pater vester exsultavit, ut videret diem meum; et vidit et gavisus est ".
JOHN|8|57|Dixerunt ergo Iudaei ad eum: " Quinquaginta annos nondum habes et Abraham vidisti? ".
JOHN|8|58|Dixit eis Iesus: " Amen, amen dico vobis: Antequam Abraham fieret, ego sum ".
JOHN|8|59|Tulerunt ergo lapides, ut iacerent in eum; Iesus autem abscondit se et exivit de templo.
JOHN|9|1|Et praeteriens vidit hominem caecum a nativitate.
JOHN|9|2|Et interro gaverunt eum discipuli sui dicentes: " Rabbi, quis peccavit, hic aut parentes eius, ut caecus nasceretur? ".
JOHN|9|3|Respondit Iesus: " Neque hic peccavit neque parentes eius, sed ut manifestentur opera Dei in illo.
JOHN|9|4|Nos oportet operari opera eius, qui misit me, donec dies est; venit nox, quando nemo potest operari.
JOHN|9|5|Quamdiu in mundo sum, lux sum mundi ".
JOHN|9|6|Haec cum dixisset, exspuit in terram et fecit lutum ex sputo et linivit lutum super oculos eius
JOHN|9|7|et dixit ei: " Vade, lava in natatoria Siloae! " - quod interpretatur Missus C. Abiit ergo et lavit et venit videns.
JOHN|9|8|Itaque vicini et, qui videbant eum prius quia mendicus erat, dicebant: " Nonne hic est, qui sedebat et mendicabat? ";
JOHN|9|9|alii dicebant: " Hic est! "; alii dicebant: " Nequaquam, sed similis est eius! ". Ille dicebat: " Ego sum! ".
JOHN|9|10|Dicebant ergo ei: " Quomodo igitur aperti sunt oculi tibi? ".
JOHN|9|11|Respondit ille: " Homo, qui dicitur Iesus, lutum fecit et unxit oculos meos et dixit mihi: "Vade ad Siloam et lava! ". Abii ergo et lavi et vidi.
JOHN|9|12|Et dixerunt ei: " Ubi est ille? ". Ait: " Nescio ".
JOHN|9|13|Adducunt eum ad pharisaeos, qui caecus fuerat.
JOHN|9|14|Erat autem sabbatum, in qua die lutum fecit Iesus et aperuit oculos eius.
JOHN|9|15|Iterum ergo interrogabant et eum pharisaei quomodo vidisset. Ille autem dixit eis: " Lutum posuit super oculos meos, et lavi et video ".
JOHN|9|16|Dicebant ergo ex pharisaeis quidam: " Non est hic homo a Deo, quia sabbatum non custodit! "; alii autem dicebant: " Quomodo potest homo peccator haec signa facere? ". Et schisma erat in eis.
JOHN|9|17|Dicunt ergo caeco iterum: " Tu quid dicis de eo quia aperuit oculos tuos? ". Ille autem dixit: " Propheta est! ".
JOHN|9|18|Non crediderunt ergo Iudaei de illo quia caecus fuisset et vidisset, donec vocaverunt parentes eius, qui viderat.
JOHN|9|19|Et interrogaverunt eos dicentes: " Hic est filius vester, quem vos dicitis quia caecus natus est? Quomodo ergo nunc videt? ".
JOHN|9|20|Responderunt ergo parentes eius et dixerunt: " Scimus quia hic est filius noster et quia caecus natus est.
JOHN|9|21|Quomodo autem nunc videat nescimus, aut quis eius aperuit oculos nos nescimus; ipsum interrogate. Aetatem habet; ipse de se loquetur! ".
JOHN|9|22|Haec dixerunt parentes eius, quia timebant Iudaeos; iam enim conspiraverant Iudaei, ut, si quis eum confiteretur Christum, extra synagogam fieret.
JOHN|9|23|Propterea parentes eius dixerunt: " Aetatem habet; ipsum interrogate!.
JOHN|9|24|Vocaverunt ergo rursum hominem, qui fuerat caecus, et dixerunt ei: " Da gloriam Deo! Nos scimus quia hic homo peccator est ".
JOHN|9|25|Respondit ergo ille: " Si peccator est nescio; unum scio quia, caecus cum essem, modo video ".
JOHN|9|26|Dixerunt ergo illi: " Quid fecit tibi? Quomodo aperuit oculos tuos? ".
JOHN|9|27|Respondit eis: " Dixi vobis iam, et non audistis; quid iterum vultis audire? Numquid et vos vultis discipuli eius fieri? ".
JOHN|9|28|Et maledixerunt ei et dixerunt: " Tu discipulus illius es, nos autem Moysis discipuli sumus.
JOHN|9|29|Nos scimus quia Moysi locutus est Deus; hunc autem nescimus unde sit ".
JOHN|9|30|Respondit homo et dixit eis: " In hoc enim mirabile est, quia vos nescitis unde sit, et aperuit meos oculos!
JOHN|9|31|Scimus quia peccatores Deus non audit; sed, si quis Dei cultor est et voluntatem eius facit, hunc exaudit.
JOHN|9|32|A saeculo non est auditum quia aperuit quis oculos caeci nati;
JOHN|9|33|nisi esset hic a Deo, non poterat facere quidquam ".
JOHN|9|34|Responderunt et dixerunt ei: " In peccatis tu natus es totus et tu doces nos? ". Et eiecerunt eum foras.
JOHN|9|35|Audivit Iesus quia eiecerunt eum foras et, cum invenisset eum, dixit ei: " Tu credis in Filium hominis? ".
JOHN|9|36|Respondit ille et dixit: " Et quis est, Domine, ut credam in eum? ".
JOHN|9|37|Dixit ei Iesus: " Et vidisti eum; et, qui loquitur tecum, ipse est ".
JOHN|9|38|At ille ait: " Credo, Domine! "; et adoravit eum.
JOHN|9|39|Et dixit Iesus: " In iudicium ego in hunc mundum veni, ut, qui non vident, videant, et, qui vident, caeci fiant ".
JOHN|9|40|Audierunt haec ex pharisaeis, qui cum ipso erant, et dixerunt ei: " Numquid et nos caeci sumus? ".
JOHN|9|41|Dixit eis Iesus: " Si caeci essetis, non haberetis peccatum. Nunc vero dicitis: "Videmus!"; peccatum vestrum manet ".
JOHN|10|1|" Amen, amen dico vobis: Qui non intrat per ostium in ovile ovium, sed ascendit aliunde, ille fur est et latro;
JOHN|10|2|qui autem intrat per ostium, pastor est ovium.
JOHN|10|3|Huic ostiarius aperit, et oves vocem eius audiunt, et proprias oves vocat nominatim et educit eas.
JOHN|10|4|Cum proprias omnes emiserit, ante eas vadit, et oves illum sequuntur, quia sciunt vocem eius;
JOHN|10|5|alienum autem non sequentur, sed fugient ab eo, quia non noverunt vocem alienorum ".
JOHN|10|6|Hoc proverbium dixit eis Iesus; illi autem non cognoverunt quid esset, quod loquebatur eis.
JOHN|10|7|Dixit ergo iterum Iesus: " Amen, amen dico vobis: Ego sum ostium ovium.
JOHN|10|8|Omnes, quotquot venerunt ante me, fures sunt et latrones, sed non audierunt eos oves.
JOHN|10|9|Ego sum ostium; per me, si quis introierit, salvabitur et ingredietur et egredietur et pascua inveniet.
JOHN|10|10|Fur non venit, nisi ut furetur et mactet et perdat; ego veni, ut vitam habeant et abundantius habeant.
JOHN|10|11|Ego sum pastor bonus; bonus pastor animam suam ponit pro ovibus;
JOHN|10|12|mercennarius et, qui non est pastor, cuius non sunt oves propriae, videt lupum venientem et dimittit oves et fugit - et lupus rapit eas et dispergit -
JOHN|10|13|quia mercennarius est et non pertinet ad eum de ovibus.
JOHN|10|14|Ego sum pastor bonus et cognosco meas, et cognoscunt me meae,
JOHN|10|15|sicut cognoscit me Pater, et ego cognosco Patrem; et animam meam pono pro ovibus.
JOHN|10|16|Et alias oves habeo, quae non sunt ex hoc ovili, et illas oportet me adducere, et vocem meam audient et fient unus grex, unus pastor.
JOHN|10|17|Propterea me Pater diligit, quia ego pono animam meam, ut iterum sumam eam.
JOHN|10|18|Nemo tollit eam a me, sed ego pono eam a meipso. Potestatem habeo ponendi eam et potestatem habeo iterum sumendi eam. Hoc mandatum accepi a Patre meo ".
JOHN|10|19|Dissensio iterum facta est inter Iudaeos propter sermones hos.
JOHN|10|20|Dicebant autem multi ex ipsis: " Daemonium habet et insanit! Quid eum auditis? ".
JOHN|10|21|Alii dicebant: " Haec verba non sunt daemonium habentis! Numquid daemonium potest caecorum oculos aperire? ".
JOHN|10|22|Facta sunt tunc Encaenia in Hierosolymis. Hiems erat;
JOHN|10|23|et ambulabat Iesus in templo in porticu Salomonis.
JOHN|10|24|Circumdederunt ergo eum Iudaei et dicebant ei: " Quousque animam nostram tollis? Si tu es Christus, dic nobis palam! ".
JOHN|10|25|Respondit eis Iesus: " Dixi vobis, et non creditis; opera, quae ego facio in nomine Patris mei, haec testimonium perhibent de me.
JOHN|10|26|Sed vos non creditis, quia non estis ex ovibus meis.
JOHN|10|27|Oves meae vocem meam audiunt, et ego cognosco eas, et sequuntur me;
JOHN|10|28|et ego vitam aeternam do eis, et non peribunt in aeternum, et non rapiet eas quisquam de manu mea.
JOHN|10|29|Pater meus quod dedit mihi, maius omnibus est, et nemo potest rapere de manu Patris.
JOHN|10|30|Ego et Pater unum sumus ".
JOHN|10|31|Sustulerunt iterum lapides Iudaei, ut lapidarent eum.
JOHN|10|32|Respondit eis Iesus: " Multa opera bona ostendi vobis ex Patre; propter quod eorum opus me lapidatis? ".
JOHN|10|33|Responderunt ei Iudaei: " De bono opere non lapidamus te sed de blasphemia, et quia tu, homo cum sis, facis teipsum Deum ".
JOHN|10|34|Respondit eis Iesus: " Nonne scriptum est in lege vestra: "Ego dixi: Dii estis?".
JOHN|10|35|Si illos dixit deos, ad quos sermo Dei factus est, et non potest solvi Scriptura,
JOHN|10|36|quem Pater sanctificavit et misit in mundum, vos dicitis: Blasphemas!", quia dixi: Filius Dei sum?
JOHN|10|37|Si non facio opera Patris mei, nolite credere mihi;
JOHN|10|38|si autem facio, et si mihi non vultis credere, operibus credite, ut cognoscatis et sciatis quia in me est Pater, et ego in Patre ".
JOHN|10|39|Quaerebant ergo iterum eum prehendere; et exivit de manibus eorum.
JOHN|10|40|Et abiit iterum trans Iordanem in eum locum, ubi erat Ioannes baptizans primum, et mansit illic.
JOHN|10|41|Et multi venerunt ad eum et dicebant: " Ioannes quidem signum fecit nullum; omnia autem, quaecumque dixit Ioannes de hoc, vera erant ".
JOHN|10|42|Et multi crediderunt in eum illic.
JOHN|11|1|Erat autem quidam lan guens Lazarus a Bethania, de castello Mariae et Marthae sororis eius.
JOHN|11|2|Maria autem erat, quae unxit Dominum unguento et extersit pedes eius capillis suis, cuius frater Lazarus infirmabatur.
JOHN|11|3|Miserunt ergo sorores ad eum dicentes: " Domine, ecce, quem amas, infirmatur ".
JOHN|11|4|Audiens autem Iesus dixit: " Infirmitas haec non est ad mortem sed pro gloria Dei, ut glorificetur Filius Dei per eam ".
JOHN|11|5|Diligebat autem Iesus Martham et sororem eius et Lazarum.
JOHN|11|6|Ut ergo audivit quia infirmabatur, tunc quidem mansit in loco, in quo erat, duobus diebus;
JOHN|11|7|deinde post hoc dicit discipulis: " Eamus in Iudaeam iterum ".
JOHN|11|8|Dicunt ei discipuli: " Rabbi, nunc quaerebant te Iudaei lapidare, et iterum vadis illuc? ".
JOHN|11|9|Respondit Iesus: " Nonne duodecim horae sunt diei? Si quis ambulaverit in die, non offendit, quia lucem huius mundi videt;
JOHN|11|10|si quis autem ambulaverit in nocte, offendit, quia lux non est in eo ".
JOHN|11|11|Haec ait et post hoc dicit eis: " Lazarus amicus noster dormit, sed vado, ut a somno exsuscitem eum ".
JOHN|11|12|Dixerunt ergo ei discipuli: " Domine, si dormit, salvus erit ".
JOHN|11|13|Dixerat autem Iesus de morte eius, illi autem putaverunt quia de dormitione somni diceret.
JOHN|11|14|Tunc ergo dixit eis Iesus manifeste: " Lazarus mortuus est,
JOHN|11|15|et gaudeo propter vos, ut credatis, quoniam non eram ibi; sed eamus ad eum ".
JOHN|11|16|Dixit ergo Thomas, qui dicitur Didymus, ad condiscipulos: " Eamus et nos, ut moriamur cum eo! ".
JOHN|11|17|Venit itaque Iesus et invenit eum quattuor dies iam in monumento habentem.
JOHN|11|18|Erat autem Bethania iuxta Hierosolymam quasi stadiis quindecim.
JOHN|11|19|Multi autem ex Iudaeis venerant ad Martham et Mariam, ut consolarentur eas de fratre.
JOHN|11|20|Martha ergo ut audivit quia Iesus venit, occurrit illi; Maria autem domi sedebat.
JOHN|11|21|Dixit ergo Martha ad Iesum: " Domine, si fuisses hic, frater meus non esset mortuus!
JOHN|11|22|Sed et nunc scio quia, quaecumque poposceris a Deo, dabit tibi Deus ".
JOHN|11|23|Dicit illi Iesus: " Resurget frater tuus ".
JOHN|11|24|Dicit ei Martha: " Scio quia resurget in resurrectione in novissimo die.
JOHN|11|25|Dixit ei Iesus: " Ego sum resurrectio et vita. Qui credit in me, etsi mortuus fuerit, vivet;
JOHN|11|26|et omnis, qui vivit et credit in me, non morietur in aeternum. Credis hoc? ".
JOHN|11|27|Ait illi: " Utique, Domine; ego credidi quia tu es Christus Filius Dei, qui in mundum venisti ".
JOHN|11|28|Et cum haec dixisset, abiit et vocavit Mariam sororem suam silentio dicens: " Magister adest et vocat te ".
JOHN|11|29|Illa autem ut audivit, surrexit cito et venit ad eum;
JOHN|11|30|nondum enim venerat Iesus in castellum, sed erat adhuc in illo loco, ubi occurrerat ei Martha.
JOHN|11|31|Iudaei igitur, qui erant cum ea in domo et consolabantur eam, cum vidissent Mariam quia cito surrexit et exiit, secuti sunt eam putantes: " Vadit ad monumentum, ut ploret ibi ".
JOHN|11|32|Maria ergo, cum venisset ubi erat Iesus, videns eum cecidit ad pedes eius dicens ei: " Domine, si fuisses hic, non esset mortuus frater meus!.
JOHN|11|33|Iesus ergo, ut vidit eam plorantem et Iudaeos, qui venerant cum ea, plorantes, fremuit spiritu et turbavit seipsum
JOHN|11|34|et dixit: " Ubi posuistis eum? ". Dicunt ei: " Domine, veni et vide ".
JOHN|11|35|Lacrimatus est Iesus.
JOHN|11|36|Dicebant ergo Iudaei: " Ecce quomodo amabat eum! ".
JOHN|11|37|Quidam autem dixerunt ex ipsis: " Non poterat hic, qui aperuit oculos caeci, facere, ut et hic non moreretur? ".
JOHN|11|38|Iesus ergo rursum fremens in semetipso, venit ad monumentum; erat autem spelunca, et lapis superpositus erat ei.
JOHN|11|39|Ait Iesus: " Tollite lapidem! ". Dicit ei Martha, soror eius, qui mortuus fuerat: " Domine, iam foetet; quatriduanus enim est! ".
JOHN|11|40|Dicit ei Iesus: " Nonne dixi tibi quoniam, si credideris, videbis gloriam Dei? ".
JOHN|11|41|Tulerunt ergo lapidem. Iesus autem, elevatis sursum oculis, dixit: " Pater, gratias ago tibi quoniam audisti me.
JOHN|11|42|Ego autem sciebam quia semper me audis, sed propter populum, qui circumstat, dixi, ut credant quia tu me misisti ".
JOHN|11|43|Et haec cum dixisset, voce magna clamavit: " Lazare, veni foras! ".
JOHN|11|44|Prodiit, qui fuerat mortuus, ligatus pedes et manus institis; et facies illius sudario erat ligata. Dicit Iesus eis: " Solvite eum et sinite eum abire ".
JOHN|11|45|Multi ergo ex Iudaeis, qui venerant ad Mariam et viderant, quae fecit, crediderunt in eum;
JOHN|11|46|quidam autem ex ipsis abierunt ad pharisaeos et dixerunt eis, quae fecit Iesus.
JOHN|11|47|Collegerunt ergo pontifices et pharisaei concilium et dicebant: " Quid facimus, quia hic homo multa signa facit?
JOHN|11|48|Si dimittimus eum sic, omnes credent in eum, et venient Romani et tollent nostrum et locum et gentem! ".
JOHN|11|49|Unus autem ex ipsis, Caiphas, cum esset pontifex anni illius, dixit eis: " Vos nescitis quidquam
JOHN|11|50|nec cogitatis quia expedit vobis, ut unus moriatur homo pro populo, et non tota gens pereat! ".
JOHN|11|51|Hoc autem a semetipso non dixit; sed, cum esset pontifex anni illius, prophetavit quia Iesus moriturus erat pro gente
JOHN|11|52|et non tantum pro gente, sed et ut filios Dei, qui erant dispersi, congregaret in unum.
JOHN|11|53|Ab illo ergo die cogitaverunt, ut interficerent eum.
JOHN|11|54|Iesus ergo iam non in palam ambulabat apud Iudaeos, sed abiit inde in regionem iuxta desertum, in civitatem, quae dicitur Ephraim, et ibi morabatur cum discipulis.
JOHN|11|55|Proximum autem erat Pascha Iudaeorum, et ascenderunt multi Hierosolymam de regione ante Pascha, ut sanctificarent seipsos.
JOHN|11|56|Quaerebant ergo Iesum et colloquebantur ad invicem in templo stantes: " Quid videtur vobis? Numquid veniet ad diem festum? ".
JOHN|11|57|Dederant autem pontifices et pharisaei mandatum, ut, si quis cognoverit, ubi sit, indicet, ut apprehendant eum.
JOHN|12|1|Iesus ergo ante sex dies Paschae venit Bethaniam, ubi erat Lazarus, quem suscitavit a mortuis Iesus.
JOHN|12|2|Fecerunt ergo ei cenam ibi, et Martha ministrabat, Lazarus vero unus erat ex discumbentibus cum eo.
JOHN|12|3|Maria ergo accepit libram unguenti nardi puri, pretiosi, et unxit pedes Iesu et extersit capillis suis pedes eius; domus autem impleta est ex odore unguenti.
JOHN|12|4|Dicit autem Iudas Iscariotes, unus ex discipulis eius, qui erat eum traditurus:
JOHN|12|5|" Quare hoc unguentum non veniit trecentis denariis et datum est egenis?.
JOHN|12|6|Dixit autem hoc, non quia de egenis pertinebat ad eum, sed quia fur erat et, loculos habens, ea, quae mittebantur, portabat.
JOHN|12|7|Dixit ergo Iesus: " Sine illam, ut in diem sepulturae meae servet illud.
JOHN|12|8|Pauperes enim semper habetis vobiscum, me autem non semper habetis ".
JOHN|12|9|Cognovit ergo turba multa ex Iudaeis quia illic est, et venerunt non propter Iesum tantum, sed ut et Lazarum viderent, quem suscitavit a mortuis.
JOHN|12|10|Cogitaverunt autem principes sacerdotum, ut et Lazarum interficerent,
JOHN|12|11|quia multi propter illum abibant ex Iudaeis et credebant in Iesum.
JOHN|12|12|In crastinum turba multa, quae venerat ad diem festum, cum audissent quia venit Iesus Hierosolymam,
JOHN|12|13|acceperunt ramos palmarum et processerunt obviam ei et clamabant: Hosanna!Benedictus, qui venit in nomine Domini, et rex Israel! ".
JOHN|12|14|Invenit autem Iesus asellum et sedit super eum, sicut scriptum est:
JOHN|12|15|" Noli timere, filia Sion.Ecce rex tuus venitsedens super pullum asinae ".
JOHN|12|16|Haec non cognoverunt discipuli eius primum, sed quando glorificatus est Iesus, tunc recordati sunt quia haec erant scripta de eo, et haec fecerunt ei.
JOHN|12|17|Testimonium ergo perhibebat turba, quae erat cum eo, quando Lazarum vocavit de monumento et suscitavit eum a mortuis.
JOHN|12|18|Propterea et obviam venit ei turba, quia audierunt eum fecisse hoc signum.
JOHN|12|19|Pharisaei ergo dixerunt ad semetipsos: " Videtis quia nihil proficitis? Ecce mundus post eum abiit! ".
JOHN|12|20|Erant autem Graeci quidam ex his, qui ascenderant, ut adorarent in die festo;
JOHN|12|21|hi ergo accesserunt ad Philippum, qui erat a Bethsaida Galilaeae, et rogabant eum dicentes: " Domine, volumus Iesum videre ".
JOHN|12|22|Venit Philippus et dicit Andreae; venit Andreas et Philippus et dicunt Iesu.
JOHN|12|23|Iesus autem respondet eis dicens: " Venit hora, ut glorificetur Filius hominis.
JOHN|12|24|Amen, amen dico vobis: Nisi granum frumenti cadens in terram mortuum fuerit, ipsum solum manet; si autem mortuum fuerit, multum fructum affert.
JOHN|12|25|Qui amat animam suam, perdit eam; et, qui odit animam suam in hoc mundo, in vitam aeternam custodiet eam.
JOHN|12|26|Si quis mihi ministrat, me sequatur, et ubi sum ego, illic et minister meus erit; si quis mihi ministraverit, honorificabit eum Pater.
JOHN|12|27|Nunc anima mea turbata est. Et quid dicam? Pater, salvifica me ex hora hac? Sed propterea veni in horam hanc.
JOHN|12|28|Pater, glorifica tuum nomen! ". Venit ergo vox de caelo: " Et glorificavi et iterum glorificabo ".
JOHN|12|29|Turba ergo, quae stabat et audierat, dicebat tonitruum factum esse; alii dicebant: " Angelus ei locutus est ".
JOHN|12|30|Respondit Iesus et dixit: " Non propter me vox haec facta est sed propter vos.
JOHN|12|31|Nunc iudicium est huius mundi, nunc princeps huius mundi eicietur foras;
JOHN|12|32|et ego, si exaltatus fuero a terra, omnes traham ad meipsum ".
JOHN|12|33|Hoc autem dicebat significans, qua morte esset moriturus.
JOHN|12|34|Respondit ergo ei turba: " Nos audivimus ex Lege, quia Christus manet in aeternum; et quomodo tu dicis: "Oportet exaltari Filium hominis"? Quis est iste Filius hominis? ".
JOHN|12|35|Dixit ergo eis Iesus: " Adhuc modicum tempus lumen in vobis est. Ambulate, dum lucem habetis, ut non tenebrae vos comprehendant; et, qui ambulat in tenebris, nescit quo vadat.
JOHN|12|36|Dum lucem habetis, credite in lucem, ut filii lucis fiatis ". Haec locutus est Iesus et abiit et abscondit se ab eis.
JOHN|12|37|Cum autem tanta signa fecisset coram eis, non credebant in eum,
JOHN|12|38|ut sermo Isaiae prophetae impleretur, quem dixit: Domine, quis credidit auditui nostro,et brachium Domini cui revelatum est? ".
JOHN|12|39|Propterea non poterant credere, quia iterum dixit Isaias:
JOHN|12|40|" Excaecavit oculos eorumet induravit eorum cor,ut non videant oculiset intellegant corde et convertantur,et sanem eos ".
JOHN|12|41|Haec dixit Isaias, quia vidit gloriam eius et locutus est de eo.
JOHN|12|42|Verumtamen et ex principibus multi crediderunt in eum, sed propter pharisaeos non confitebantur, ut de synagoga non eicerentur;
JOHN|12|43|dilexerunt enim gloriam hominum magis quam gloriam Dei.
JOHN|12|44|Iesus autem clamavit et dixit: " Qui credit in me, non credit in me sed in eum, qui misit me;
JOHN|12|45|et, qui videt me, videt eum, qui misit me.
JOHN|12|46|Ego lux in mundum veni, ut omnis, qui credit in me, in tenebris non maneat.
JOHN|12|47|Et si quis audierit verba mea et non custodierit, ego non iudico eum; non enim veni, ut iudicem mundum, sed ut salvificem mundum.
JOHN|12|48|Qui spernit me et non accipit verba mea, habet, qui iudicet eum: sermo, quem locutus sum, ille iudicabit eum in novissimo die,
JOHN|12|49|quia ego ex meipso non sum locutus, sed, qui misit me, Pater, ipse mihi mandatum dedit quid dicam et quid loquar.
JOHN|12|50|Et scio quia mandatum eius vita aeterna est. Quae ergo ego loquor, sicut dixit mihi Pater, sic loquor ".
JOHN|13|1|Ante diem autem festum Pa schae, sciens Iesus quia venit eius hora, ut transeat ex hoc mundo ad Patrem, cum dilexisset suos, qui erant in mundo, in finem dilexit eos.
JOHN|13|2|Et in cena, cum Diabolus iam misisset in corde, ut traderet eum Iudas Simonis Iscariotis,
JOHN|13|3|sciens quia omnia dedit ei Pater in manus, et quia a Deo exivit et ad Deum vadit,
JOHN|13|4|surgit a cena et ponit vestimenta sua et, cum accepisset linteum, praecinxit se.
JOHN|13|5|Deinde mittit aquam in pelvem et coepit lavare pedes discipulorum et extergere linteo, quo erat praecinctus.
JOHN|13|6|Venit ergo ad Simonem Petrum. Dicit ei: " Domine, tu mihi lavas pedes?.
JOHN|13|7|Respondit Iesus et dixit ei: " Quod ego facio, tu nescis modo, scies autem postea ".
JOHN|13|8|Dicit ei Petrus: " Non lavabis mihi pedes in aeternum! ". Respondit Iesus ei: " Si non lavero te, non habes partem mecum ".
JOHN|13|9|Dicit ei Simon Petrus: " Domine, non tantum pedes meos sed et manus et caput! ".
JOHN|13|10|Dicit ei Iesus: " Qui lotus est, non indiget nisi ut pedes lavet, sed est mundus totus; et vos mundi estis sed non omnes ".
JOHN|13|11|Sciebat enim quisnam esset, qui traderet eum; propterea dixit: " Non estis mundi omnes ".
JOHN|13|12|Postquam ergo lavit pedes eorum et accepit vestimenta sua, cum recubuisset iterum, dixit eis: " Scitis quid fecerim vobis?
JOHN|13|13|Vos vocatis me: "Magister" et: "Domine", et bene dicitis; sum etenim.
JOHN|13|14|Si ergo ego lavi vestros pedes, Dominus et Magister, et vos debetis alter alterius lavare pedes.
JOHN|13|15|Exemplum enim dedi vobis, ut, quemadmodum ego feci vobis, et vos faciatis.
JOHN|13|16|Amen, amen dico vobis: Non est servus maior domino suo, neque apostolus maior eo, qui misit illum.
JOHN|13|17|Si haec scitis, beati estis, si facitis ea.
JOHN|13|18|Non de omnibus vobis dico, ego scio, quos elegerim, sed ut impleatur Scriptura: "Qui manducat meum panem, levavit contra me calcaneum suum".
JOHN|13|19|Amodo dico vobis priusquam fiat, ut credatis, cum factum fuerit, quia ego sum.
JOHN|13|20|Amen, amen dico vobis: Qui accipit, si quem misero, me accipit; qui autem me accipit, accipit eum, qui me misit ".
JOHN|13|21|Cum haec dixisset Iesus, turbatus est spiritu et protestatus est et dixit: " Amen, amen dico vobis: Unus ex vobis tradet me ".
JOHN|13|22|Aspiciebant ad invicem discipuli, haesitantes de quo diceret.
JOHN|13|23|Erat recumbens unus ex discipulis eius in sinu Iesu, quem diligebat Iesus.
JOHN|13|24|Innuit ergo huic Simon Petrus, ut interrogaret: " Quis est, de quo dicit? ".
JOHN|13|25|Cum ergo recumberet ille ita supra pectus Iesu, dicit ei: " Domine, quis est? ".
JOHN|13|26|Respondet Iesus: " Ille est, cui ego intinctam buccellam porrexero ". Cum ergo intinxisset buccellam, dat Iudae Simonis Iscariotis.
JOHN|13|27|Et post buccellam tunc introivit in illum Satanas. Dicit ergo ei Iesus: Quod facis, fac citius ".
JOHN|13|28|Hoc autem nemo scivit discumbentium ad quid dixerit ei;
JOHN|13|29|quidam enim putabant quia loculos habebat Iudas, quia dicit ei Iesus: " Eme ea, quae opus sunt nobis ad diem festum ", aut egenis ut aliquid daret.
JOHN|13|30|Cum ergo accepisset ille buccellam, exivit continuo; erat autem nox.
JOHN|13|31|Cum ergo exisset, dicit Iesus: " Nunc clarificatus est Filius hominis, et Deus clarificatus est in eo;
JOHN|13|32|si Deus clarificatus est in eo, et Deus clarificabit eum in semetipso et continuo clarificabit eum.
JOHN|13|33|Filioli, adhuc modicum vobiscum sum; quaeretis me, et sicut dixi Iudaeis: Quo ego vado, vos non potestis venire, et vobis dico modo.
JOHN|13|34|Mandatum novum do vobis, ut diligatis invicem; sicut dilexi vos, ut et vos diligatis invicem.
JOHN|13|35|In hoc cognoscent omnes quia mei discipuli estis: si dilectionem habueritis ad invicem ".
JOHN|13|36|Dicit ei Simon Petrus: " Domine, quo vadis? ". Respondit Iesus: " Quo vado, non potes me modo sequi, sequeris autem postea ".
JOHN|13|37|Dicit ei Petrus: " Domine, quare non possum te sequi modo? Animam meam pro te ponam ".
JOHN|13|38|Respondet Iesus: " Animam tuam pro me pones? Amen, amen dico tibi: Non cantabit gallus, donec me ter neges.
JOHN|14|1|Non turbetur cor vestrum. Creditis in Deum et in me credite.
JOHN|14|2|In domo Patris mei mansiones multae sunt; si quo minus, dixissem vobis, quia vado parare vobis locum?
JOHN|14|3|Et si abiero et praeparavero vobis locum, iterum venio et accipiam vos ad meipsum, ut, ubi sum ego, et vos sitis.
JOHN|14|4|Et quo ego vado, scitis viam ".
JOHN|14|5|Dicit ei Thomas: " Domine, nescimus quo vadis; quomodo possumus viam scire? ".
JOHN|14|6|Dicit ei Iesus: " Ego sum via et veritas et vita; nemo venit ad Patrem nisi per me.
JOHN|14|7|Si cognovistis me, et Patrem meum utique cognoscetis; et amodo cognoscitis eum et vidistis eum ".
JOHN|14|8|Dicit ei Philippus: " Domine, ostende nobis Patrem, et sufficit nobis ".
JOHN|14|9|Dicit ei Iesus: " Tanto tempore vobiscum sum, et non cognovisti me, Philippe? Qui vidit me, vidit Patrem. Quomodo tu dicis: "Ostende nobis Patrem"?
JOHN|14|10|Non credis quia ego in Patre, et Pater in me est? Verba, quae ego loquor vobis, a meipso non loquor; Pater autem in me manens facit opera sua.
JOHN|14|11|Credite mihi quia ego in Patre, et Pater in me est; alioquin propter opera ipsa credite.
JOHN|14|12|Amen, amen dico vobis: Qui credit in me, opera, quae ego facio, et ipse faciet et maiora horum faciet, quia ego ad Patrem vado.
JOHN|14|13|Et quodcumque petieritis in nomine meo, hoc faciam, ut glorificetur Pater in Filio;
JOHN|14|14|si quid petieritis me in nomine meo, ego faciam.
JOHN|14|15|Si diligitis me, mandata mea servabitis;
JOHN|14|16|et ego rogabo Patrem, et alium Paraclitum dabit vobis, ut maneat vobiscum in aeternum,
JOHN|14|17|Spiritum veritatis, quem mundus non potest accipere, quia non videt eum nec cognoscit. Vos cognoscitis eum, quia apud vos manet; et in vobis erit.
JOHN|14|18|Non relinquam vos orphanos; venio ad vos.
JOHN|14|19|Adhuc modicum, et mundus me iam non videt; vos autem videtis me, quia ego vivo et vos vivetis.
JOHN|14|20|In illo die vos cognoscetis quia ego sum in Patre meo, et vos in me, et ego in vobis.
JOHN|14|21|Qui habet mandata mea et servat ea, ille est, qui diligit me; qui autem diligit me, diligetur a Patre meo, et ego diligam eum et manifestabo ei meipsum ".
JOHN|14|22|Dicit ei Iudas, non ille Iscariotes: " Domine, et quid factum est, quia nobis manifestaturus es teipsum et non mundo? ".
JOHN|14|23|Respondit Iesus et dixit ei: " Si quis diligit me, sermonem meum servabit, et Pater meus diliget eum, et ad eum veniemus et mansionem apud eum faciemus;
JOHN|14|24|qui non diligit me, sermones meos non servat. Et sermo, quem auditis, non est meus, sed eius qui misit me, Patris.
JOHN|14|25|Haec locutus sum vobis apud vos manens.
JOHN|14|26|Paraclitus autem, Spiritus Sanctus, quem mittet Pater in nomine meo, ille vos docebit omnia et suggeret vobis omnia, quae dixi vobis.
JOHN|14|27|Pacem relinquo vobis, pacem meam do vobis; non quomodo mundus dat, ego do vobis. Non turbetur cor vestrum neque formidet.
JOHN|14|28|Audistis quia ego dixi vobis: Vado et venio ad vos. Si diligeretis me, gauderetis quia vado ad Patrem, quia Pater maior me est.
JOHN|14|29|Et nunc dixi vobis, priusquam fiat, ut, cum factum fuerit, credatis.
JOHN|14|30|Iam non multa loquar vobiscum, venit enim princeps mundi et in me non habet quidquam;
JOHN|14|31|sed, ut cognoscat mundus quia diligo Patrem, et sicut mandatum dedit mihi Pater, sic facio. Surgite, eamus hinc.
JOHN|15|1|Ego sum vitis vera, et Pater meus agricola est.
JOHN|15|2|Omnem palmitem in me non ferentem fructum tollit eum; et omnem, qui fert fructum, purgat eum, ut fructum plus afferat.
JOHN|15|3|Iam vos mundi estis propter sermonem, quem locutus sum vobis.
JOHN|15|4|Manete in me, et ego in vobis. Sicut palmes non potest ferre fructum a semetipso, nisi manserit in vite, sic nec vos, nisi in me manseritis.
JOHN|15|5|Ego sum vitis, vos palmites. Qui manet in me, et ego in eo, hic fert fructum multum, quia sine me nihil potestis facere.
JOHN|15|6|Si quis in me non manserit, missus est foras sicut palmes et aruit; et colligunt eos et in ignem mittunt, et ardent.
JOHN|15|7|Si manseritis in me, et verba mea in vobis manserint, quodcumque volueritis, petite, et fiet vobis.
JOHN|15|8|In hoc clarificatus est Pater meus, ut fructum multum afferatis et efficiamini mei discipuli.
JOHN|15|9|Sicut dilexit me Pater, et ego dilexi vos; manete in dilectione mea.
JOHN|15|10|Si praecepta mea servaveritis, manebitis in dilectione mea, sicut ego Patris mei praecepta servavi et maneo in eius dilectione.
JOHN|15|11|Haec locutus sum vobis, ut gaudium meum in vobis sit, et gaudium vestrum impleatur.
JOHN|15|12|Hoc est praeceptum meum, ut diligatis invicem, sicut dilexi vos;
JOHN|15|13|maiorem hac dilectionem nemo habet, ut animam suam quis ponat pro amicis suis.
JOHN|15|14|Vos amici mei estis, si feceritis, quae ego praecipio vobis.
JOHN|15|15|Iam non dico vos servos, quia servus nescit quid facit dominus eius; vos autem dixi amicos, quia omnia, quae audivi a Patre meo, nota feci vobis.
JOHN|15|16|Non vos me elegistis, sed ego elegi vos et posui vos, ut vos eatis et fructum afferatis, et fructus vester maneat, ut quodcumque petieritis Patrem in nomine meo, det vobis.
JOHN|15|17|Haec mando vobis, ut diligatis invicem.
JOHN|15|18|Si mundus vos odit, scitote quia me priorem vobis odio habuit.
JOHN|15|19|Si de mundo essetis, mundus, quod suum est, diligeret; quia vero de mundo non estis, sed ego elegi vos de mundo, propterea odit vos mundus.
JOHN|15|20|Mementote sermonis, quem ego dixi vobis: Non est servus maior domino suo. Si me persecuti sunt, et vos persequentur; si sermonem meum servaverunt, et vestrum servabunt.
JOHN|15|21|Sed haec omnia facient vobis propter nomen meum, quia nesciunt eum, qui misit me.
JOHN|15|22|Si non venissem et locutus fuissem eis, peccatum non haberent; nunc autem excusationem non habent de peccato suo.
JOHN|15|23|Qui me odit et Patrem meum odit.
JOHN|15|24|Si opera non fecissem in eis, quae nemo alius fecit, peccatum non haberent; nunc autem et viderunt et oderunt et me et Patrem meum.
JOHN|15|25|Sed ut impleatur sermo, qui in lege eorum scriptus est: "Odio me habuerunt gratis".
JOHN|15|26|Cum autem venerit Paraclitus, quem ego mittam vobis a Patre, Spiritum veritatis, qui a Patre procedit, ille testimonium perhibebit de me;
JOHN|15|27|sed et vos testimonium perhibetis, quia ab initio mecum estis.
JOHN|16|1|Haec locutus sum vobis, ut non scandalizemini.
JOHN|16|2|Absque synagogis facient vos; sed venit hora, ut omnis, qui interficit vos, arbitretur obsequium se praestare Deo.
JOHN|16|3|Et haec facient, quia non noverunt Patrem neque me.
JOHN|16|4|Sed haec locutus sum vobis, ut, cum venerit hora eorum, reminiscamini eorum, quia ego dixi vobis. Haec autem vobis ab initio non dixi, quia vobiscum eram.
JOHN|16|5|At nunc vado ad eum, qui me misit, et nemo ex vobis interrogat me: "Quo vadis?".
JOHN|16|6|Sed quia haec locutus sum vobis, tristitia implevit cor vestrum.
JOHN|16|7|Sed ego veritatem dico vobis: Expedit vobis, ut ego vadam. Si enim non abiero, Paraclitus non veniet ad vos; si autem abiero, mittam eum ad vos.
JOHN|16|8|Et cum venerit ille, arguet mundum de peccato et de iustitia et de iudicio:
JOHN|16|9|de peccato quidem, quia non credunt in me;
JOHN|16|10|de iustitia vero, quia ad Patrem vado, et iam non videtis me;
JOHN|16|11|de iudicio autem, quia princeps mundi huius iudicatus est.
JOHN|16|12|Adhuc multa habeo vobis dicere, sed non potestis portare modo.
JOHN|16|13|Cum autem venerit ille, Spiritus veritatis, deducet vos in omnem veritatem; non enim loquetur a semetipso, sed quaecumque audiet, loquetur et, quae ventura sunt, annuntiabit vobis.
JOHN|16|14|Ille me clarificabit, quia de meo accipiet et annuntiabit vobis.
JOHN|16|15|Omnia, quaecumque habet Pater, mea sunt; propterea dixi quia de meo accipit et annuntiabit vobis.
JOHN|16|16|Modicum, et iam non videtis me; et iterum modicum, et videbitis me ".
JOHN|16|17|Dixerunt ergo ex discipulis eius ad invicem: " Quid est hoc, quod dicit nobis: "Modicum, et non videtis me; et iterum modicum, et videbitis me" et: "Vado ad Patrem"? ".
JOHN|16|18|Dicebant ergo: " Quid est hoc, quod dicit: "Modicum"? Nescimus quid loquitur ".
JOHN|16|19|Cognovit Iesus quia volebant eum interrogare et dixit eis: " De hoc quaeritis inter vos, quia dixi: "Modicum, et non videtis me; et iterum modicum, et videbitis me"?
JOHN|16|20|Amen, amen dico vobis quia plorabitis et flebitis vos, mundus autem gaudebit; vos contristabimini, sed tristitia vestra vertetur in gaudium.
JOHN|16|21|Mulier, cum parit, tristitiam habet, quia venit hora eius; cum autem pepererit puerum, iam non meminit pressurae propter gaudium, quia natus est homo in mundum.
JOHN|16|22|Et vos igitur nunc quidem tristitiam habetis; iterum autem videbo vos, et gaudebit cor vestrum, et gaudium vestrum nemo tollit a vobis.
JOHN|16|23|Et in illo die me non rogabitis quidquam.Amen, amen dico vobis: Si quid petieritis Patrem in nomine meo, dabit vobis.
JOHN|16|24|Usque modo non petistis quidquam in nomine meo. Petite et accipietis, ut gaudium vestrum sit plenum.
JOHN|16|25|Haec in proverbiis locutus sum vobis; venit hora, cum iam non in proverbiis loquar vobis, sed palam de Patre annuntiabo vobis.
JOHN|16|26|Illo die in nomine meo petetis, et non dico vobis quia ego rogabo Patrem de vobis;
JOHN|16|27|ipse enim Pater amat vos, quia vos me amastis et credidistis quia ego a Deo exivi.
JOHN|16|28|Exivi a Patre et veni in mundum; iterum relinquo mundum et vado ad Patrem ".
JOHN|16|29|Dicunt discipuli eius: " Ecce nunc palam loqueris, et proverbium nullum dicis.
JOHN|16|30|Nunc scimus quia scis omnia, et non opus est tibi, ut quis te interroget; in hoc credimus quia a Deo existi ".
JOHN|16|31|Respondit eis Iesus: " Modo creditis?
JOHN|16|32|Ecce venit hora et iam venit, ut dispergamini unusquisque in propria et me solum relinquatis; et non sum solus, quia Pater mecum est.
JOHN|16|33|Haec locutus sum vobis, ut in me pacem habeatis; in mundo pressuram habetis, sed confidite, ego vici mundum ".
JOHN|17|1|Haec locutus est Iesus; et, sublevatis oculis suis in cae lum, dixit: " Pater, venit hora: clarifica Filium tuum, ut Filius clarificet te,
JOHN|17|2|sicut dedisti ei potestatem omnis carnis, ut omne, quod dedisti ei, det eis vitam aeternam.
JOHN|17|3|Haec est autem vita aeterna, ut cognoscant te solum verum Deum et, quem misisti, Iesum Christum.
JOHN|17|4|Ego te clarificavi super terram; opus consummavi, quod dedisti mihi, ut faciam;
JOHN|17|5|et nunc clarifica me tu, Pater, apud temetipsum claritate, quam habebam, priusquam mundus esset, apud te.
JOHN|17|6|Manifestavi nomen tuum hominibus, quos dedisti mihi de mundo. Tui erant, et mihi eos dedisti, et sermonem tuum servaverunt.
JOHN|17|7|Nunc cognoverunt quia omnia, quae dedisti mihi, abs te sunt,
JOHN|17|8|quia verba, quae dedisti mihi, dedi eis; et ipsi acceperunt et cognoverunt vere quia a te exivi et crediderunt quia tu me misisti.
JOHN|17|9|Ego pro eis rogo; non pro mundo rogo, sed pro his, quos dedisti mihi, quia tui sunt;
JOHN|17|10|et mea omnia tua sunt, et tua mea; et clarificatus sum in eis.
JOHN|17|11|Et iam non sum in mundo, et hi in mundo sunt, et ego ad te venio.Pater sancte, serva eos in nomine tuo, quod dedisti mihi, ut sint unum sicut nos.
JOHN|17|12|Cum essem cum eis, ego servabam eos in nomine tuo, quod dedisti mihi, et custodivi, et nemo ex his periit, nisi filius perditionis, ut Scriptura impleatur.
JOHN|17|13|Nunc autem ad te venio et haec loquor in mundo, ut habeant gaudium meum impletum in semetipsis.
JOHN|17|14|Ego dedi eis sermonem tuum, et mundus odio eos habuit, quia non sunt de mundo, sicut ego non sum de mundo.
JOHN|17|15|Non rogo, ut tollas eos de mundo, sed ut serves eos ex Malo.
JOHN|17|16|De mundo non sunt, sicut ego non sum de mundo.
JOHN|17|17|Sanctifica eos in veritate; sermo tuus veritas est.
JOHN|17|18|Sicut me misisti in mundum, et ego misi eos in mundum;
JOHN|17|19|et pro eis ego sanctifico meipsum, ut sint et ipsi sanctificati in veritate.
JOHN|17|20|Non pro his autem rogo tantum, sed et pro eis, qui credituri sunt per verbum eorum in me,
JOHN|17|21|ut omnes unum sint, sicut tu, Pater, in me et ego in te, ut et ipsi in nobis unum sint; ut mundus credat quia tu me misisti.
JOHN|17|22|Et ego claritatem, quam dedisti mihi, dedi illis, ut sint unum, sicut nos unum sumus;
JOHN|17|23|ego in eis, et tu in me, ut sint consummati in unum; ut cognoscat mundus, quia tu me misisti et dilexisti eos, sicut me dilexisti.
JOHN|17|24|Pater, quod dedisti mihi, volo, ut ubi ego sum, et illi sint mecum, ut videant claritatem meam, quam dedisti mihi, quia dilexisti me ante constitutionem mundi.
JOHN|17|25|Pater iuste, et mundus te non cognovit; ego autem te cognovi, et hi cognoverunt quia tu me misisti;
JOHN|17|26|et notum feci eis nomen tuum et notum faciam, ut dilectio, qua dilexisti me, in ipsis sit, et ego in ipsis ".
JOHN|18|1|Haec cum dixisset Iesus, egressus est cum discipulis suis trans torrentem Cedron, ubi erat hortus, in quem introivit ipse et discipuli eius.
JOHN|18|2|Sciebat autem et Iudas, qui tradebat eum, locum, quia frequenter Iesus convenerat illuc cum discipulis suis.
JOHN|18|3|Iudas ergo, cum accepisset cohortem et a pontificibus et pharisaeis ministros, venit illuc cum lanternis et facibus et armis.
JOHN|18|4|Iesus itaque sciens omnia, quae ventura erant super eum, processit et dicit eis: " Quem quaeritis? ".
JOHN|18|5|Responderunt ei: " Iesum Nazarenum ". Dicit eis: " Ego sum! ". Stabat autem et Iudas, qui tradebat eum, cum ipsis.
JOHN|18|6|Ut ergo dixit eis: " Ego sum! ", abierunt retrorsum et ceciderunt in terram.
JOHN|18|7|Iterum ergo eos interrogavit: " Quem quaeritis? ". Illi autem dixerunt: Iesum Nazarenum ".
JOHN|18|8|Respondit Iesus: " Dixi vobis: Ego sum! Si ergo me quaeritis, sinite hos abire ",
JOHN|18|9|ut impleretur sermo, quem dixit: " Quos dedisti mihi, non perdidi ex ipsis quemquam ".
JOHN|18|10|Simon ergo Petrus, habens gladium, eduxit eum et percussit pontificis servum et abscidit eius auriculam dextram. Erat autem nomen servo Malchus.
JOHN|18|11|Dixit ergo Iesus Petro: " Mitte gladium in vaginam; calicem, quem dedit mihi Pater, non bibam illum? ".
JOHN|18|12|Cohors ergo et tribunus et ministri Iudaeorum comprehenderunt Iesum et ligaverunt eum
JOHN|18|13|et adduxerunt ad Annam primum; erat enim socer Caiphae, qui erat pontifex anni illius.
JOHN|18|14|Erat autem Caiphas, qui consilium dederat Iudaeis: " Expedit unum hominem mori pro populo ".
JOHN|18|15|Sequebatur autem Iesum Simon Petrus et alius discipulus. Discipulus autem ille erat notus pontifici et introivit cum Iesu in atrium pontificis;
JOHN|18|16|Petrus autem stabat ad ostium foris. Exivit ergo discipulus alius, qui erat notus pontifici, et dixit ostiariae et introduxit Petrum.
JOHN|18|17|Dicit ergo Petro ancilla ostiaria: " Numquid et tu ex discipulis es hominis istius? ". Dicit ille: " Non sum! ".
JOHN|18|18|Stabant autem servi et ministri, qui prunas fecerant, quia frigus erat, et calefaciebant se; erat autem cum eis et Petrus stans et calefaciens se.
JOHN|18|19|Pontifex ergo interrogavit Iesum de discipulis suis et de doctrina eius.
JOHN|18|20|Respondit ei Iesus: " Ego palam locutus sum mundo; ego semper docui in synagoga et in templo, quo omnes Iudaei conveniunt, et in occulto locutus sum nihil.
JOHN|18|21|Quid me interrogas? Interroga eos, qui audierunt quid locutus sum ipsis; ecce hi sciunt, quae dixerim ego ".
JOHN|18|22|Haec autem cum dixisset, unus assistens ministrorum dedit alapam Iesu dicens: " Sic respondes pontifici? ".
JOHN|18|23|Respondit ei Iesus: " Si male locutus sum, testimonium perhibe de malo; si autem bene, quid me caedis? ".
JOHN|18|24|Misit ergo eum Annas ligatum ad Caipham pontificem.
JOHN|18|25|Erat autem Simon Petrus stans et calefaciens se. Dixerunt ergo ei: " Numquid et tu ex discipulis eius es? ". Negavit ille et dixit: " Non sum!.
JOHN|18|26|Dicit unus ex servis pontificis, cognatus eius, cuius abscidit Petrus auriculam: " Nonne ego te vidi in horto cum illo? ".
JOHN|18|27|Iterum ergo negavit Petrus; et statim gallus cantavit.
JOHN|18|28|Adducunt ergo Iesum a Caipha in praetorium. Erat autem mane. Et ipsi non introierunt in praetorium, ut non contaminarentur, sed manducarent Pascha.
JOHN|18|29|Exivit ergo Pilatus ad eos foras et dicit: " Quam accusationem affertis adversus hominem hunc? ".
JOHN|18|30|Responderunt et dixerunt ei: " Si non esset hic malefactor, non tibi tradidissemus eum ".
JOHN|18|31|Dixit ergo eis Pilatus: " Accipite eum vos et secundum legem vestram iudicate eum! ". Dixerunt ei Iudaei: " Nobis non licet interficere quemquam ",
JOHN|18|32|ut sermo Iesu impleretur, quem dixit, significans qua esset morte moriturus.
JOHN|18|33|Introivit ergo iterum in praetorium Pilatus et vocavit Iesum et dixit ei: " Tu es rex Iudaeorum? ".
JOHN|18|34|Respondit Iesus: " A temetipso tu hoc dicis, an alii tibi dixerunt de me? ".
JOHN|18|35|Respondit Pilatus: " Numquid ego Iudaeus sum? Gens tua et pontifices tradiderunt te mihi; quid fecisti? ".
JOHN|18|36|Respondit Iesus: " Regnum meum non est de mundo hoc; si ex hoc mundo esset regnum meum, ministri mei decertarent, ut non traderer Iudaeis; nunc autem meum regnum non est hinc ".
JOHN|18|37|Dixit itaque ei Pilatus: " Ergo rex es tu? ". Respondit Iesus: " Tu dicis quia rex sum. Ego in hoc natus sum et ad hoc veni in mundum, ut testimonium perhibeam veritati; omnis, qui est ex veritate, audit meam vocem ".
JOHN|18|38|Dicit ei Pilatus: " Quid est veritas? ". Et cum hoc dixisset, iterum exivit ad Iudaeos et dicit eis: " Ego nullam invenio in eo causam.
JOHN|18|39|Est autem consuetudo vobis, ut unum dimittam vobis in Pascha; vultis ergo dimittam vobis regem Iudaeorum? ".
JOHN|18|40|Clamaverunt ergo rursum dicentes: " Non hunc sed Barabbam! ". Erat autem Barabbas latro.
JOHN|19|1|Tunc ergo apprehendit Pi latus Iesum et flagellavit.
JOHN|19|2|Et milites, plectentes coronam de spinis, imposuerunt capiti eius et veste purpurea circumdederunt eum;
JOHN|19|3|et veniebant ad eum et dicebant: " Ave, rex Iudaeorum! ", et dabant ei alapas.
JOHN|19|4|Et exiit iterum Pilatus foras et dicit eis: " Ecce adduco vobis eum foras, ut cognoscatis quia in eo invenio causam nullam ".
JOHN|19|5|Exiit ergo Iesus foras, portans spineam coronam et purpureum vestimentum. Et dicit eis: " Ecce homo! ".
JOHN|19|6|Cum ergo vidissent eum pontifices et ministri, clamaverunt dicentes: " Crucifige, crucifige! ". Dicit eis Pilatus: " Accipite eum vos et crucifigite; ego enim non invenio in eo causam ".
JOHN|19|7|Responderunt ei Iudaei: " Nos legem habemus, et secundum legem debet mori, quia Filium Dei se fecit ".
JOHN|19|8|Cum ergo audisset Pilatus hunc sermonem, magis timuit
JOHN|19|9|et ingressus est praetorium iterum et dicit ad Iesum: " Unde es tu? ". Iesus autem responsum non dedit ei.
JOHN|19|10|Dicit ergo ei Pilatus: " Mihi non loqueris? Nescis quia potestatem habeo dimittere te et potestatem habeo crucifigere te? ".
JOHN|19|11|Respondit Iesus: " Non haberes potestatem adversum me ullam, nisi tibi esset datum desuper; propterea, qui tradidit me tibi, maius peccatum habet.
JOHN|19|12|Exinde quaerebat Pilatus dimittere eum; Iudaei autem clamabant dicentes: " Si hunc dimittis, non es amicus Caesaris! Omnis, qui se regem facit, contradicit Caesari ".
JOHN|19|13|Pilatus ergo, cum audisset hos sermones, adduxit foras Iesum et sedit pro tribunali in locum, qui dicitur Lithostrotos, Hebraice autem Gabbatha.
JOHN|19|14|Erat autem Parasceve Paschae, hora erat quasi sexta. Et dicit Iudaeis: Ecce rex vester! ".
JOHN|19|15|Clamaverunt ergo illi: " Tolle, tolle, crucifige eum! ". Dicit eis Pilatus: " Regem vestrum crucifigam? ". Responderunt pontifices: " Non habemus regem, nisi Caesarem ".
JOHN|19|16|Tunc ergo tradidit eis illum, ut crucifigeretur. Susceperunt ergo Iesum.
JOHN|19|17|Et baiulans sibi crucem exivit in eum, qui dicitur Calvariae locum, quod Hebraice dicitur Golgotha,
JOHN|19|18|ubi eum crucifixerunt et cum eo alios duos hinc et hinc, medium autem Iesum.
JOHN|19|19|Scripsit autem et titulum Pilatus et posuit super crucem; erat autem scriptum: " Iesus Nazarenus Rex Iudaeorum ".
JOHN|19|20|Hunc ergo titulum multi legerunt Iudaeorum, quia prope civitatem erat locus, ubi crucifixus est Iesus; et erat scriptum Hebraice, Latine, Graece.
JOHN|19|21|Dicebant ergo Pilato pontifices Iudaeorum: " Noli scribere: Rex Iudaeorum, sed: Ipse dixit: "Rex sum Iudaeorum" ".
JOHN|19|22|Respondit Pilatus: " Quod scripsi, scripsi! ".
JOHN|19|23|Milites ergo cum crucifixissent Iesum, acceperunt vestimenta eius et fecerunt quattuor partes, unicuique militi partem, et tunicam. Erat autem tunica inconsutilis, desuper contexta per totum.
JOHN|19|24|Dixerunt ergo ad invicem: " Non scindamus eam, sed sortiamur de illa,cuius sit ", ut Scriptura impleatur dicens: Partiti sunt vestimenta mea sibiet in vestem meam miserunt sortem ".Et milites quidem haec fecerunt.
JOHN|19|25|Stabant autem iuxta crucem Iesu mater eius et soror matris eius, Maria Cleopae, et Maria Magdalene.
JOHN|19|26|Cum vidisset ergo Iesus matrem et discipulum stantem, quem diligebat, dicit matri: " Mulier, ecce filius tuus ".
JOHN|19|27|Deinde dicit discipulo: " Ecce mater tua ". Et ex illa hora accepit eam discipulus in sua.
JOHN|19|28|Post hoc sciens Iesus quia iam omnia consummata sunt, ut consummaretur Scriptura, dicit: " Sitio ".
JOHN|19|29|Vas positum erat aceto plenum; spongiam ergo plenam aceto hyssopo circumponentes, obtulerunt ori eius.
JOHN|19|30|Cum ergo accepisset acetum, Iesus dixit: " Consummatum est! ". Et inclinato capite tradidit spiritum.
JOHN|19|31|Iudaei ergo, quoniam Parasceve erat, ut non remanerent in cruce corpora sabbato, erat enim magnus dies illius sabbati, rogaverunt Pilatum, ut frangerentur eorum crura, et tollerentur.
JOHN|19|32|Venerunt ergo milites et primi quidem fregerunt crura et alterius, qui crucifixus est cum eo;
JOHN|19|33|ad Iesum autem cum venissent, ut viderunt eum iam mortuum, non fregerunt eius crura,
JOHN|19|34|sed unus militum lancea latus eius aperuit, et continuo exivit sanguis et aqua.
JOHN|19|35|Et qui vidit, testimonium perhibuit, et verum est eius testimonium, et ille scit quia vera dicit, ut et vos credatis.
JOHN|19|36|Facta sunt enim haec, ut Scriptura impleatur: " Os non comminuetur eius,
JOHN|19|37|et iterum alia Scriptura dicit: " Videbunt in quem transfixerunt ".
JOHN|19|38|Post haec autem rogavit Pilatum Ioseph ab Arimathaea, qui erat discipulus Iesu, occultus autem propter metum Iudaeorum, ut tolleret corpus Iesu; et permisit Pilatus. Venit ergo et tulit corpus eius.
JOHN|19|39|Venit autem et Nicodemus, qui venerat ad eum nocte primum, ferens mixturam myrrhae et aloes quasi libras centum.
JOHN|19|40|Acceperunt ergo corpus Iesu et ligaverunt illud linteis cum aromatibus, sicut mos Iudaeis est sepelire.
JOHN|19|41|Erat autem in loco, ubi crucifixus est, hortus, et in horto monumentum novum, in quo nondum quisquam positus erat.
JOHN|19|42|Ibi ergo propter Parascevem Iudaeorum, quia iuxta erat monumentum, posuerunt Iesum.
JOHN|20|1|Prima autem sabbatorum Maria Magdalene venit ma ne, cum adhuc tenebrae essent, ad monumentum et videt lapidem sublatum a monumento.
JOHN|20|2|Currit ergo et venit ad Simonem Petrum et ad alium discipulum, quem amabat Iesus, et dicit eis: " Tulerunt Dominum de monumento, et nescimus, ubi posuerunt eum! ".
JOHN|20|3|Exiit ergo Petrus et ille alius discipulus, et veniebant ad monumentum.
JOHN|20|4|Currebant autem duo simul, et ille alius discipulus praecucurrit citius Petro et venit primus ad monumentum;
JOHN|20|5|et cum se inclinasset, videt posita linteamina, non tamen introivit.
JOHN|20|6|Venit ergo et Simon Petrus sequens eum et introivit in monumentum; et videt linteamina posita
JOHN|20|7|et sudarium, quod fuerat super caput eius, non cum linteaminibus positum, sed separatim involutum in unum locum.
JOHN|20|8|Tunc ergo introivit et alter discipulus, qui venerat primus ad monumentum, et vidit et credidit.
JOHN|20|9|Nondum enim sciebant Scripturam, quia oportet eum a mortuis resurgere.
JOHN|20|10|Abierunt ergo iterum ad semetipsos discipuli.
JOHN|20|11|Maria autem stabat ad monumentum foris plorans. Dum ergo fleret, inclinavit se in monumentum
JOHN|20|12|et videt duos angelos in albis sedentes, unum ad caput et unum ad pedes, ubi positum fuerat corpus Iesu.
JOHN|20|13|Et dicunt ei illi: " Mulier, quid ploras? ". Dicit eis: " Tulerunt Dominum meum, et nescio, ubi posuerunt eum ".
JOHN|20|14|Haec cum dixisset, conversa est retrorsum et videt Iesum stantem; et non sciebat quia Iesus est.
JOHN|20|15|Dicit ei Iesus: " Mulier, quid ploras? Quem quaeris? ". Illa, existimans quia hortulanus esset, dicit ei: " Domine, si tu sustulisti eum, dicito mihi, ubi posuisti eum, et ego eum tollam ".
JOHN|20|16|Dicit ei Iesus: " Maria! ". Conversa illa dicit ei Hebraice: " Rabbuni! - quod dicitur Magister C.
JOHN|20|17|Dicit ei Iesus: " Iam noli me tenere, nondum enim ascendi ad Patrem; vade autem ad fratres meos et dic eis: Ascendo ad Patrem meum et Patrem vestrum, et Deum meum et Deum vestrum ".
JOHN|20|18|Venit Maria Magdalene annuntians discipulis: " Vidi Dominum! ", et quia haec dixit ei.
JOHN|20|19|Cum esset ergo sero die illa prima sabbatorum, et fores essent clausae, ubi erant discipuli, propter metum Iudaeorum, venit Iesus et stetit in medio et dicit eis: " Pax vobis! ".
JOHN|20|20|Et hoc cum dixisset, ostendit eis manus et latus. Gavisi sunt ergo discipuli, viso Domino.
JOHN|20|21|Dixit ergo eis iterum: " Pax vobis! Sicut misit me Pater, et ego mitto vos ".
JOHN|20|22|Et cum hoc dixisset, insufflavit et dicit eis: " Accipite Spiritum Sanctum.
JOHN|20|23|Quorum remiseritis peccata, remissa sunt eis; quorum retinueritis, retenta sunt ".
JOHN|20|24|Thomas autem, unus ex Duodecim, qui dicitur Didymus, non erat cum eis, quando venit Iesus.
JOHN|20|25|Dicebant ergo ei alii discipuli: " Vidimus Dominum! ". Ille autem dixit eis: " Nisi videro in manibus eius signum clavorum et mittam digitum meum in signum clavorum et mittam manum meam in latus eius, non credam ".
JOHN|20|26|Et post dies octo iterum erant discipuli eius intus, et Thomas cum eis. Venit Iesus ianuis clausis et stetit in medio et dixit: " Pax vobis! ".
JOHN|20|27|Deinde dicit Thomae: " Infer digitum tuum huc et vide manus meas et affer manum tuam et mitte in latus meum; et noli fieri incredulus sed fidelis! ".
JOHN|20|28|Respondit Thomas et dixit ei: " Dominus meus et Deus meus! ".
JOHN|20|29|Dicit ei Iesus: " Quia vidisti me, credidisti. Beati, qui non viderunt et crediderunt! ".
JOHN|20|30|Multa quidem et alia signa fecit Iesus in conspectu discipulorum suorum, quae non sunt scripta in libro hoc;
JOHN|20|31|haec autem scripta sunt, ut credatis quia Iesus est Christus Filius Dei et ut credentes vitam habeatis in nomine eius.
JOHN|21|1|Postea manifestavit se ite rum Iesus discipulis ad mare Tiberiadis; manifestavit autem sic.
JOHN|21|2|Erant simul Simon Petrus et Thomas, qui dicitur Didymus, et Nathanael, qui erat a Cana Galilaeae, et filii Zebedaei et alii ex discipulis eius duo.
JOHN|21|3|Dicit eis Simon Petrus: " Vado piscari ". Dicunt ei: " Venimus et nos tecum ". Exierunt et ascenderunt in navem; et illa nocte nihil prendiderunt.
JOHN|21|4|Mane autem iam facto, stetit Iesus in litore; non tamen sciebant discipuli quia Iesus est.
JOHN|21|5|Dicit ergo eis Iesus: " Pueri, numquid pulmentarium habetis? ". Responderunt ei: " Non ".
JOHN|21|6|Ille autem dixit eis: " Mittite in dexteram navigii rete et invenietis. Miserunt ergo et iam non valebant illud trahere a multitudine piscium.
JOHN|21|7|Dicit ergo discipulus ille, quem diligebat Iesus, Petro: " Dominus est!. Simon ergo Petrus, cum audisset quia Dominus est, tunicam succinxit se, erat enim nudus, et misit se in mare;
JOHN|21|8|alii autem discipuli navigio venerunt, non enim longe erant a terra, sed quasi cubitis ducentis, trahentes rete piscium.
JOHN|21|9|Ut ergo descenderunt in terram, vident prunas positas et piscem superpositum et panem.
JOHN|21|10|Dicit eis Iesus: " Afferte de piscibus, quos prendidistis nunc ".
JOHN|21|11|Ascendit ergo Simon Petrus et traxit rete in terram, plenum magnis piscibus centum quinquaginta tribus; et cum tanti essent, non est scissum rete.
JOHN|21|12|Dicit eis Iesus: " Venite, prandete ". Nemo autem audebat discipulorum interrogare eum: " Tu quis es? ", scientes quia Dominus est.
JOHN|21|13|Venit Iesus et accipit panem et dat eis et piscem similiter.
JOHN|21|14|Hoc iam tertio manifestatus est Iesus discipulis, cum resurrexisset a mortuis.
JOHN|21|15|Cum ergo prandissent, dicit Simoni Petro Iesus: " Simon Ioannis, diligis me plus his? ". Dicit ei: " Etiam, Domine, tu scis quia amo te ". Dicit ei: " Pasce agnos meos ".
JOHN|21|16|Dicit ei iterum secundo: " Simon Ioannis, diligis me? ". Ait illi: " Etiam, Domine, tu scis quia amo te ". Dicit ei: " Pasce oves meas ".
JOHN|21|17|Dicit ei tertio: " Simon Ioannis, amas me? ". Contristatus est Petrus quia dixit ei tertio: " Amas me? ", et dicit ei: " Domine, tu omnia scis, tu cognoscis quia amo te ". Dicit ei: " Pasce oves meas.
JOHN|21|18|Amen, amen dico tibi: Cum esses iunior, cingebas teipsum et ambulabas, ubi volebas; cum autem senueris, extendes manus tuas, et alius te cinget et ducet, quo non vis ".
JOHN|21|19|Hoc autem dixit significans qua morte clarificaturus esset Deum. Et hoc cum dixisset, dicit ei: " Sequere me ".
JOHN|21|20|Conversus Petrus videt illum discipulum, quem diligebat Iesus, sequentem, qui et recubuit in cena super pectus eius et dixit: " Domine, quis est qui tradit te? ".
JOHN|21|21|Hunc ergo cum vidisset Petrus, dicit Iesu: " Domine, hic autem quid? ".
JOHN|21|22|Dicit ei Iesus: " Si eum volo manere donec veniam, quid ad te? Tu me sequere ".
JOHN|21|23|Exivit ergo sermo iste in fratres, quia discipulus ille non moritur. Non autem dixit ei Iesus: " Non moritur ", sed: " Si eum volo manere donec veniam, quid ad te? ".
JOHN|21|24|Hic est discipulus, qui testimonium perhibet de his et scripsit haec; et scimus quia verum est testimonium eius.
JOHN|21|25|Sunt autem et alia multa, quae fecit Iesus; quae, si scribantur per singula, nec ipsum arbitror mundum capere eos, qui scribendi sunt, libros.
