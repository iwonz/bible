LUKE|1|1|quoniam quidem multi conati sunt ordinare narrationem quae in nobis conpletae sunt rerum
LUKE|1|2|sicut tradiderunt nobis qui ab initio ipsi viderunt et ministri fuerunt sermonis
LUKE|1|3|visum est et mihi adsecuto a principio omnibus diligenter ex ordine tibi scribere optime Theophile
LUKE|1|4|ut cognoscas eorum verborum de quibus eruditus es veritatem
LUKE|1|5|fuit in diebus Herodis regis Iudaeae sacerdos quidam nomine Zaccharias de vice Abia et uxor illi de filiabus Aaron et nomen eius Elisabeth
LUKE|1|6|erant autem iusti ambo ante Deum incedentes in omnibus mandatis et iustificationibus Domini sine querella
LUKE|1|7|et non erat illis filius eo quod esset Elisabeth sterilis et ambo processissent in diebus suis
LUKE|1|8|factum est autem cum sacerdotio fungeretur in ordine vicis suae ante Deum
LUKE|1|9|secundum consuetudinem sacerdotii sorte exiit ut incensum poneret ingressus in templum Domini
LUKE|1|10|et omnis multitudo erat populi orans foris hora incensi
LUKE|1|11|apparuit autem illi angelus Domini stans a dextris altaris incensi
LUKE|1|12|et Zaccharias turbatus est videns et timor inruit super eum
LUKE|1|13|ait autem ad illum angelus ne timeas Zaccharia quoniam exaudita est deprecatio tua et uxor tua Elisabeth pariet tibi filium et vocabis nomen eius Iohannem
LUKE|1|14|et erit gaudium tibi et exultatio et multi in nativitate eius gaudebunt
LUKE|1|15|erit enim magnus coram Domino et vinum et sicera non bibet et Spiritu Sancto replebitur adhuc ex utero matris suae
LUKE|1|16|et multos filiorum Israhel convertet ad Dominum Deum ipsorum
LUKE|1|17|et ipse praecedet ante illum in spiritu et virtute Heliae ut convertat corda patrum in filios et incredibiles ad prudentiam iustorum parare Domino plebem perfectam
LUKE|1|18|et dixit Zaccharias ad angelum unde hoc sciam ego enim sum senex et uxor mea processit in diebus suis
LUKE|1|19|et respondens angelus dixit ei ego sum Gabrihel qui adsto ante Deum et missus sum loqui ad te et haec tibi evangelizare
LUKE|1|20|et ecce eris tacens et non poteris loqui usque in diem quo haec fiant pro eo quod non credidisti verbis meis quae implebuntur in tempore suo
LUKE|1|21|et erat plebs expectans Zacchariam et mirabantur quod tardaret ipse in templo
LUKE|1|22|egressus autem non poterat loqui ad illos et cognoverunt quod visionem vidisset in templo et ipse erat innuens illis et permansit mutus
LUKE|1|23|et factum est ut impleti sunt dies officii eius abiit in domum suam
LUKE|1|24|post hos autem dies concepit Elisabeth uxor eius et occultabat se mensibus quinque dicens
LUKE|1|25|quia sic mihi fecit Dominus in diebus quibus respexit auferre obprobrium meum inter homines
LUKE|1|26|in mense autem sexto missus est angelus Gabrihel a Deo in civitatem Galilaeae cui nomen Nazareth
LUKE|1|27|ad virginem desponsatam viro cui nomen erat Ioseph de domo David et nomen virginis Maria
LUKE|1|28|et ingressus angelus ad eam dixit have gratia plena Dominus tecum benedicta tu in mulieribus
LUKE|1|29|quae cum vidisset turbata est in sermone eius et cogitabat qualis esset ista salutatio
LUKE|1|30|et ait angelus ei ne timeas Maria invenisti enim gratiam apud Deum
LUKE|1|31|ecce concipies in utero et paries filium et vocabis nomen eius Iesum
LUKE|1|32|hic erit magnus et Filius Altissimi vocabitur et dabit illi Dominus Deus sedem David patris eius
LUKE|1|33|et regnabit in domo Iacob in aeternum et regni eius non erit finis
LUKE|1|34|dixit autem Maria ad angelum quomodo fiet istud quoniam virum non cognosco
LUKE|1|35|et respondens angelus dixit ei Spiritus Sanctus superveniet in te et virtus Altissimi obumbrabit tibi ideoque et quod nascetur sanctum vocabitur Filius Dei
LUKE|1|36|et ecce Elisabeth cognata tua et ipsa concepit filium in senecta sua et hic mensis est sextus illi quae vocatur sterilis
LUKE|1|37|quia non erit inpossibile apud Deum omne verbum
LUKE|1|38|dixit autem Maria ecce ancilla Domini fiat mihi secundum verbum tuum et discessit ab illa angelus
LUKE|1|39|exsurgens autem Maria in diebus illis abiit in montana cum festinatione in civitatem Iuda
LUKE|1|40|et intravit in domum Zacchariae et salutavit Elisabeth
LUKE|1|41|et factum est ut audivit salutationem Mariae Elisabeth exultavit infans in utero eius et repleta est Spiritu Sancto Elisabeth
LUKE|1|42|et exclamavit voce magna et dixit benedicta tu inter mulieres et benedictus fructus ventris tui
LUKE|1|43|et unde hoc mihi ut veniat mater Domini mei ad me
LUKE|1|44|ecce enim ut facta est vox salutationis tuae in auribus meis exultavit in gaudio infans in utero meo
LUKE|1|45|et beata quae credidit quoniam perficientur ea quae dicta sunt ei a Domino
LUKE|1|46|et ait Maria magnificat anima mea Dominum
LUKE|1|47|et exultavit spiritus meus in Deo salutari meo
LUKE|1|48|quia respexit humilitatem ancillae suae ecce enim ex hoc beatam me dicent omnes generationes
LUKE|1|49|quia fecit mihi magna qui potens est et sanctum nomen eius
LUKE|1|50|et misericordia eius in progenies et progenies timentibus eum
LUKE|1|51|fecit potentiam in brachio suo dispersit superbos mente cordis sui
LUKE|1|52|deposuit potentes de sede et exaltavit humiles
LUKE|1|53|esurientes implevit bonis et divites dimisit inanes
LUKE|1|54|suscepit Israhel puerum suum memorari misericordiae
LUKE|1|55|sicut locutus est ad patres nostros Abraham et semini eius in saecula
LUKE|1|56|mansit autem Maria cum illa quasi mensibus tribus et reversa est in domum suam
LUKE|1|57|Elisabeth autem impletum est tempus pariendi et peperit filium
LUKE|1|58|et audierunt vicini et cognati eius quia magnificavit Dominus misericordiam suam cum illa et congratulabantur ei
LUKE|1|59|et factum est in die octavo venerunt circumcidere puerum et vocabant eum nomine patris eius Zacchariam
LUKE|1|60|et respondens mater eius dixit nequaquam sed vocabitur Iohannes
LUKE|1|61|et dixerunt ad illam quia nemo est in cognatione tua qui vocetur hoc nomine
LUKE|1|62|innuebant autem patri eius quem vellet vocari eum
LUKE|1|63|et postulans pugillarem scripsit dicens Iohannes est nomen eius et mirati sunt universi
LUKE|1|64|apertum est autem ilico os eius et lingua eius et loquebatur benedicens Deum
LUKE|1|65|et factus est timor super omnes vicinos eorum et super omnia montana Iudaeae divulgabantur omnia verba haec
LUKE|1|66|et posuerunt omnes qui audierant in corde suo dicentes quid putas puer iste erit etenim manus Domini erat cum illo
LUKE|1|67|et Zaccharias pater eius impletus est Spiritu Sancto et prophetavit dicens
LUKE|1|68|benedictus Deus Israhel quia visitavit et fecit redemptionem plebi suae
LUKE|1|69|et erexit cornu salutis nobis in domo David pueri sui
LUKE|1|70|sicut locutus est per os sanctorum qui a saeculo sunt prophetarum eius
LUKE|1|71|salutem ex inimicis nostris et de manu omnium qui oderunt nos
LUKE|1|72|ad faciendam misericordiam cum patribus nostris et memorari testamenti sui sancti
LUKE|1|73|iusiurandum quod iuravit ad Abraham patrem nostrum
LUKE|1|74|daturum se nobis ut sine timore de manu inimicorum nostrorum liberati serviamus illi
LUKE|1|75|in sanctitate et iustitia coram ipso omnibus diebus nostris
LUKE|1|76|et tu puer propheta Altissimi vocaberis praeibis enim ante faciem Domini parare vias eius
LUKE|1|77|ad dandam scientiam salutis plebi eius in remissionem peccatorum eorum
LUKE|1|78|per viscera misericordiae Dei nostri in quibus visitavit nos oriens ex alto
LUKE|1|79|inluminare his qui in tenebris et in umbra mortis sedent ad dirigendos pedes nostros in viam pacis
LUKE|1|80|puer autem crescebat et confortabatur spiritu et erat in deserto usque in diem ostensionis suae ad Israhel
LUKE|2|1|factum est autem in diebus illis exiit edictum a Caesare Augusto ut describeretur universus orbis
LUKE|2|2|haec descriptio prima facta est praeside Syriae Cyrino
LUKE|2|3|et ibant omnes ut profiterentur singuli in suam civitatem
LUKE|2|4|ascendit autem et Ioseph a Galilaea de civitate Nazareth in Iudaeam civitatem David quae vocatur Bethleem eo quod esset de domo et familia David
LUKE|2|5|ut profiteretur cum Maria desponsata sibi uxore praegnate
LUKE|2|6|factum est autem cum essent ibi impleti sunt dies ut pareret
LUKE|2|7|et peperit filium suum primogenitum et pannis eum involvit et reclinavit eum in praesepio quia non erat eis locus in diversorio
LUKE|2|8|et pastores erant in regione eadem vigilantes et custodientes vigilias noctis supra gregem suum
LUKE|2|9|et ecce angelus Domini stetit iuxta illos et claritas Dei circumfulsit illos et timuerunt timore magno
LUKE|2|10|et dixit illis angelus nolite timere ecce enim evangelizo vobis gaudium magnum quod erit omni populo
LUKE|2|11|quia natus est vobis hodie salvator qui est Christus Dominus in civitate David
LUKE|2|12|et hoc vobis signum invenietis infantem pannis involutum et positum in praesepio
LUKE|2|13|et subito facta est cum angelo multitudo militiae caelestis laudantium Deum et dicentium
LUKE|2|14|gloria in altissimis Deo et in terra pax in hominibus bonae voluntatis
LUKE|2|15|et factum est ut discesserunt ab eis angeli in caelum pastores loquebantur ad invicem transeamus usque Bethleem et videamus hoc verbum quod factum est quod fecit Dominus et ostendit nobis
LUKE|2|16|et venerunt festinantes et invenerunt Mariam et Ioseph et infantem positum in praesepio
LUKE|2|17|videntes autem cognoverunt de verbo quod dictum erat illis de puero hoc
LUKE|2|18|et omnes qui audierunt mirati sunt et de his quae dicta erant a pastoribus ad ipsos
LUKE|2|19|Maria autem conservabat omnia verba haec conferens in corde suo
LUKE|2|20|et reversi sunt pastores glorificantes et laudantes Deum in omnibus quae audierant et viderant sicut dictum est ad illos
LUKE|2|21|et postquam consummati sunt dies octo ut circumcideretur vocatum est nomen eius Iesus quod vocatum est ab angelo priusquam in utero conciperetur
LUKE|2|22|et postquam impleti sunt dies purgationis eius secundum legem Mosi tulerunt illum in Hierusalem ut sisterent eum Domino
LUKE|2|23|sicut scriptum est in lege Domini quia omne masculinum adaperiens vulvam sanctum Domino vocabitur
LUKE|2|24|et ut darent hostiam secundum quod dictum est in lege Domini par turturum aut duos pullos columbarum
LUKE|2|25|et ecce homo erat in Hierusalem cui nomen Symeon et homo iste iustus et timoratus expectans consolationem Israhel et Spiritus Sanctus erat in eo
LUKE|2|26|et responsum acceperat ab Spiritu Sancto non visurum se mortem nisi prius videret Christum Domini
LUKE|2|27|et venit in Spiritu in templum et cum inducerent puerum Iesum parentes eius ut facerent secundum consuetudinem legis pro eo
LUKE|2|28|et ipse accepit eum in ulnas suas et benedixit Deum et dixit
LUKE|2|29|nunc dimittis servum tuum Domine secundum verbum tuum in pace
LUKE|2|30|quia viderunt oculi mei salutare tuum
LUKE|2|31|quod parasti ante faciem omnium populorum
LUKE|2|32|lumen ad revelationem gentium et gloriam plebis tuae Israhel
LUKE|2|33|et erat pater eius et mater mirantes super his quae dicebantur de illo
LUKE|2|34|et benedixit illis Symeon et dixit ad Mariam matrem eius ecce positus est hic in ruinam et resurrectionem multorum in Israhel et in signum cui contradicetur
LUKE|2|35|et tuam ipsius animam pertransiet gladius ut revelentur ex multis cordibus cogitationes
LUKE|2|36|et erat Anna prophetissa filia Phanuhel de tribu Aser haec processerat in diebus multis et vixerat cum viro suo annis septem a virginitate sua
LUKE|2|37|et haec vidua usque ad annos octoginta quattuor quae non discedebat de templo ieiuniis et obsecrationibus serviens nocte ac die
LUKE|2|38|et haec ipsa hora superveniens confitebatur Domino et loquebatur de illo omnibus qui expectabant redemptionem Hierusalem
LUKE|2|39|et ut perfecerunt omnia secundum legem Domini reversi sunt in Galilaeam in civitatem suam Nazareth
LUKE|2|40|puer autem crescebat et confortabatur plenus sapientia et gratia Dei erat in illo
LUKE|2|41|et ibant parentes eius per omnes annos in Hierusalem in die sollemni paschae
LUKE|2|42|et cum factus esset annorum duodecim ascendentibus illis in Hierosolymam secundum consuetudinem diei festi
LUKE|2|43|consummatisque diebus cum redirent remansit puer Iesus in Hierusalem et non cognoverunt parentes eius
LUKE|2|44|existimantes autem illum esse in comitatu venerunt iter diei et requirebant eum inter cognatos et notos
LUKE|2|45|et non invenientes regressi sunt in Hierusalem requirentes eum
LUKE|2|46|et factum est post triduum invenerunt illum in templo sedentem in medio doctorum audientem illos et interrogantem
LUKE|2|47|stupebant autem omnes qui eum audiebant super prudentia et responsis eius
LUKE|2|48|et videntes admirati sunt et dixit mater eius ad illum fili quid fecisti nobis sic ecce pater tuus et ego dolentes quaerebamus te
LUKE|2|49|et ait ad illos quid est quod me quaerebatis nesciebatis quia in his quae Patris mei sunt oportet me esse
LUKE|2|50|et ipsi non intellexerunt verbum quod locutus est ad illos
LUKE|2|51|et descendit cum eis et venit Nazareth et erat subditus illis et mater eius conservabat omnia verba haec in corde suo
LUKE|2|52|et Iesus proficiebat sapientia aetate et gratia apud Deum et homines
LUKE|3|1|anno autem quintodecimo imperii Tiberii Caesaris procurante Pontio Pilato Iudaeam tetrarcha autem Galilaeae Herode Philippo autem fratre eius tetrarcha Itureae et Trachonitidis regionis et Lysania Abilinae tetrarcha
LUKE|3|2|sub principibus sacerdotum Anna et Caiapha factum est verbum Dei super Iohannem Zacchariae filium in deserto
LUKE|3|3|et venit in omnem regionem Iordanis praedicans baptismum paenitentiae in remissionem peccatorum
LUKE|3|4|sicut scriptum est in libro sermonum Esaiae prophetae vox clamantis in deserto parate viam Domini rectas facite semitas eius
LUKE|3|5|omnis vallis implebitur et omnis mons et collis humiliabitur et erunt prava in directa et aspera in vias planas
LUKE|3|6|et videbit omnis caro salutare Dei
LUKE|3|7|dicebat ergo ad turbas quae exiebant ut baptizarentur ab ipso genimina viperarum quis ostendit vobis fugere a ventura ira
LUKE|3|8|facite ergo fructus dignos paenitentiae et ne coeperitis dicere patrem habemus Abraham dico enim vobis quia potest Deus de lapidibus istis suscitare filios Abrahae
LUKE|3|9|iam enim securis ad radicem arborum posita est omnis ergo arbor non faciens fructum exciditur et in ignem mittitur
LUKE|3|10|et interrogabant eum turbae dicentes quid ergo faciemus
LUKE|3|11|respondens autem dicebat illis qui habet duas tunicas det non habenti et qui habet escas similiter faciat
LUKE|3|12|venerunt autem et publicani ut baptizarentur et dixerunt ad illum magister quid faciemus
LUKE|3|13|at ille dixit ad eos nihil amplius quam quod constitutum est vobis faciatis
LUKE|3|14|interrogabant autem eum et milites dicentes quid faciemus et nos et ait illis neminem concutiatis neque calumniam faciatis et contenti estote stipendiis vestris
LUKE|3|15|existimante autem populo et cogitantibus omnibus in cordibus suis de Iohanne ne forte ipse esset Christus
LUKE|3|16|respondit Iohannes dicens omnibus ego quidem aqua baptizo vos venit autem fortior me cuius non sum dignus solvere corrigiam calciamentorum eius ipse vos baptizabit in Spiritu Sancto et igni
LUKE|3|17|cuius ventilabrum in manu eius et purgabit aream suam et congregabit triticum in horreum suum paleas autem conburet igni inextinguibili
LUKE|3|18|multa quidem et alia exhortans evangelizabat populum
LUKE|3|19|Herodes autem tetrarcha cum corriperetur ab illo de Herodiade uxore fratris sui et de omnibus malis quae fecit Herodes
LUKE|3|20|adiecit et hoc supra omnia et inclusit Iohannem in carcere
LUKE|3|21|factum est autem cum baptizaretur omnis populus et Iesu baptizato et orante apertum est caelum
LUKE|3|22|et descendit Spiritus Sanctus corporali specie sicut columba in ipsum et vox de caelo facta est tu es Filius meus dilectus in te conplacuit mihi
LUKE|3|23|et ipse Iesus erat incipiens quasi annorum triginta ut putabatur filius Ioseph qui fuit Heli
LUKE|3|24|qui fuit Matthat qui fuit Levi qui fuit Melchi qui fuit Iannae qui fuit Ioseph
LUKE|3|25|qui fuit Matthathiae qui fuit Amos qui fuit Naum qui fuit Esli qui fuit Naggae
LUKE|3|26|qui fuit Maath qui fuit Matthathiae qui fuit Semei qui fuit Iosech qui fuit Ioda
LUKE|3|27|qui fuit Iohanna qui fuit Resa qui fuit Zorobabel qui fuit Salathihel qui fuit Neri
LUKE|3|28|qui fuit Melchi qui fuit Addi qui fuit Cosam qui fuit Helmadam qui fuit Her
LUKE|3|29|qui fuit Iesu qui fuit Eliezer qui fuit Iorim qui fuit Matthat qui fuit Levi
LUKE|3|30|qui fuit Symeon qui fuit Iuda qui fuit Ioseph qui fuit Iona qui fuit Eliachim
LUKE|3|31|qui fuit Melea qui fuit Menna qui fuit Matthata qui fuit Nathan qui fuit David
LUKE|3|32|qui fuit Iesse qui fuit Obed qui fuit Booz qui fuit Salmon qui fuit Naasson
LUKE|3|33|qui fuit Aminadab qui fuit Aram qui fuit Esrom qui fuit Phares qui fuit Iudae
LUKE|3|34|qui fuit Iacob qui fuit Isaac qui fuit Abraham qui fuit Thare qui fuit Nachor
LUKE|3|35|qui fuit Seruch qui fuit Ragau qui fuit Phalec qui fuit Eber qui fuit Sale
LUKE|3|36|qui fuit Cainan qui fuit Arfaxat qui fuit Sem qui fuit Noe qui fuit Lamech
LUKE|3|37|qui fuit Mathusalae qui fuit Enoch qui fuit Iared qui fuit Malelehel qui fuit Cainan
LUKE|3|38|qui fuit Enos qui fuit Seth qui fuit Adam qui fuit Dei
LUKE|4|1|Iesus autem plenus Spiritu Sancto regressus est ab Iordane et agebatur in Spiritu in desertum
LUKE|4|2|diebus quadraginta et temptabatur a diabolo et nihil manducavit in diebus illis et consummatis illis esuriit
LUKE|4|3|dixit autem illi diabolus si Filius Dei es dic lapidi huic ut panis fiat
LUKE|4|4|et respondit ad illum Iesus scriptum est quia non in pane solo vivet homo sed in omni verbo Dei
LUKE|4|5|et duxit illum diabolus et ostendit illi omnia regna orbis terrae in momento temporis
LUKE|4|6|et ait ei tibi dabo potestatem hanc universam et gloriam illorum quia mihi tradita sunt et cui volo do illa
LUKE|4|7|tu ergo si adoraveris coram me erunt tua omnia
LUKE|4|8|et respondens Iesus dixit illi scriptum est Dominum Deum tuum adorabis et illi soli servies
LUKE|4|9|et duxit illum in Hierusalem et statuit eum supra pinnam templi et dixit illi si Filius Dei es mitte te hinc deorsum
LUKE|4|10|scriptum est enim quod angelis suis mandabit de te ut conservent te
LUKE|4|11|et quia in manibus tollent te ne forte offendas ad lapidem pedem tuum
LUKE|4|12|et respondens Iesus ait illi dictum est non temptabis Dominum Deum tuum
LUKE|4|13|et consummata omni temptatione diabolus recessit ab illo usque ad tempus
LUKE|4|14|et regressus est Iesus in virtute Spiritus in Galilaeam et fama exiit per universam regionem de illo
LUKE|4|15|et ipse docebat in synagogis eorum et magnificabatur ab omnibus
LUKE|4|16|et venit Nazareth ubi erat nutritus et intravit secundum consuetudinem suam die sabbati in synagogam et surrexit legere
LUKE|4|17|et traditus est illi liber prophetae Esaiae et ut revolvit librum invenit locum ubi scriptum erat
LUKE|4|18|Spiritus Domini super me propter quod unxit me evangelizare pauperibus misit me
LUKE|4|19|praedicare captivis remissionem et caecis visum dimittere confractos in remissionem praedicare annum Domini acceptum et diem retributionis
LUKE|4|20|et cum plicuisset librum reddidit ministro et sedit et omnium in synagoga oculi erant intendentes in eum
LUKE|4|21|coepit autem dicere ad illos quia hodie impleta est haec scriptura in auribus vestris
LUKE|4|22|et omnes testimonium illi dabant et mirabantur in verbis gratiae quae procedebant de ore ipsius et dicebant nonne hic filius est Ioseph
LUKE|4|23|et ait illis utique dicetis mihi hanc similitudinem medice cura te ipsum quanta audivimus facta in Capharnaum fac et hic in patria tua
LUKE|4|24|ait autem amen dico vobis quia nemo propheta acceptus est in patria sua
LUKE|4|25|in veritate dico vobis multae viduae erant in diebus Heliae in Israhel quando clusum est caelum annis tribus et mensibus sex cum facta est fames magna in omni terra
LUKE|4|26|et ad nullam illarum missus est Helias nisi in Sareptha Sidoniae ad mulierem viduam
LUKE|4|27|et multi leprosi erant in Israhel sub Heliseo propheta et nemo eorum mundatus est nisi Neman Syrus
LUKE|4|28|et repleti sunt omnes in synagoga ira haec audientes
LUKE|4|29|et surrexerunt et eiecerunt illum extra civitatem et duxerunt illum usque ad supercilium montis supra quem civitas illorum erat aedificata ut praecipitarent eum
LUKE|4|30|ipse autem transiens per medium illorum ibat
LUKE|4|31|et descendit in Capharnaum civitatem Galilaeae ibique docebat illos sabbatis
LUKE|4|32|et stupebant in doctrina eius quia in potestate erat sermo ipsius
LUKE|4|33|et in synagoga erat homo habens daemonium inmundum et exclamavit voce magna
LUKE|4|34|dicens sine quid nobis et tibi Iesu Nazarene venisti perdere nos scio te qui sis Sanctus Dei
LUKE|4|35|et increpavit illi Iesus dicens obmutesce et exi ab illo et cum proiecisset illum daemonium in medium exiit ab illo nihilque illum nocuit
LUKE|4|36|et factus est pavor in omnibus et conloquebantur ad invicem dicentes quod est hoc verbum quia in potestate et virtute imperat inmundis spiritibus et exeunt
LUKE|4|37|et divulgabatur fama de illo in omnem locum regionis
LUKE|4|38|surgens autem de synagoga introivit in domum Simonis socrus autem Simonis tenebatur magnis febribus et rogaverunt illum pro ea
LUKE|4|39|et stans super illam imperavit febri et dimisit illam et continuo surgens ministrabat illis
LUKE|4|40|cum sol autem occidisset omnes qui habebant infirmos variis languoribus ducebant illos ad eum at ille singulis manus inponens curabat eos
LUKE|4|41|exiebant autem etiam daemonia a multis clamantia et dicentia quia tu es Filius Dei et increpans non sinebat ea loqui quia sciebant ipsum esse Christum
LUKE|4|42|facta autem die egressus ibat in desertum locum et turbae requirebant eum et venerunt usque ad ipsum et detinebant illum ne discederet ab eis
LUKE|4|43|quibus ille ait quia et aliis civitatibus oportet me evangelizare regnum Dei quia ideo missus sum
LUKE|4|44|et erat praedicans in synagogis Galilaeae
LUKE|5|1|factum est autem cum turbae inruerent in eum ut audirent verbum Dei et ipse stabat secus stagnum Gennesareth
LUKE|5|2|et vidit duas naves stantes secus stagnum piscatores autem descenderant et lavabant retia
LUKE|5|3|ascendens autem in unam navem quae erat Simonis rogavit eum a terra reducere pusillum et sedens docebat de navicula turbas
LUKE|5|4|ut cessavit autem loqui dixit ad Simonem duc in altum et laxate retia vestra in capturam
LUKE|5|5|et respondens Simon dixit illi praeceptor per totam noctem laborantes nihil cepimus in verbo autem tuo laxabo rete
LUKE|5|6|et cum hoc fecissent concluserunt piscium multitudinem copiosam rumpebatur autem rete eorum
LUKE|5|7|et annuerunt sociis qui erant in alia navi ut venirent et adiuvarent eos et venerunt et impleverunt ambas naviculas ita ut mergerentur
LUKE|5|8|quod cum videret Simon Petrus procidit ad genua Iesu dicens exi a me quia homo peccator sum Domine
LUKE|5|9|stupor enim circumdederat eum et omnes qui cum illo erant in captura piscium quam ceperant
LUKE|5|10|similiter autem Iacobum et Iohannem filios Zebedaei qui erant socii Simonis et ait ad Simonem Iesus noli timere ex hoc iam homines eris capiens
LUKE|5|11|et subductis ad terram navibus relictis omnibus secuti sunt illum
LUKE|5|12|et factum est cum esset in una civitatum et ecce vir plenus lepra et videns Iesum et procidens in faciem rogavit eum dicens Domine si vis potes me mundare
LUKE|5|13|et extendens manum tetigit illum dicens volo mundare et confestim lepra discessit ab illo
LUKE|5|14|et ipse praecepit illi ut nemini diceret sed vade ostende te sacerdoti et offer pro emundatione tua sicut praecepit Moses in testimonium illis
LUKE|5|15|perambulabat autem magis sermo de illo et conveniebant turbae multae ut audirent et curarentur ab infirmitatibus suis
LUKE|5|16|ipse autem secedebat in deserto et orabat
LUKE|5|17|et factum est in una dierum et ipse sedebat docens et erant Pharisaei sedentes et legis doctores qui venerant ex omni castello Galilaeae et Iudaeae et Hierusalem et virtus erat Domini ad sanandum eos
LUKE|5|18|et ecce viri portantes in lecto hominem qui erat paralyticus et quaerebant eum inferre et ponere ante eum
LUKE|5|19|et non invenientes qua parte illum inferrent prae turba ascenderunt supra tectum per tegulas submiserunt illum cum lecto in medium ante Iesum
LUKE|5|20|quorum fidem ut vidit dixit homo remittuntur tibi peccata tua
LUKE|5|21|et coeperunt cogitare scribae et Pharisaei dicentes quis est hic qui loquitur blasphemias quis potest dimittere peccata nisi solus Deus
LUKE|5|22|ut cognovit autem Iesus cogitationes eorum respondens dixit ad illos quid cogitatis in cordibus vestris
LUKE|5|23|quid est facilius dicere dimittuntur tibi peccata an dicere surge et ambula
LUKE|5|24|ut autem sciatis quia Filius hominis potestatem habet in terra dimittere peccata ait paralytico tibi dico surge tolle lectum tuum et vade in domum tuam
LUKE|5|25|et confestim surgens coram illis tulit in quo iacebat et abiit in domum suam magnificans Deum
LUKE|5|26|et stupor adprehendit omnes et magnificabant Deum et repleti sunt timore dicentes quia vidimus mirabilia hodie
LUKE|5|27|et post haec exiit et vidit publicanum nomine Levi sedentem ad teloneum et ait illi sequere me
LUKE|5|28|et relictis omnibus surgens secutus est eum
LUKE|5|29|et fecit ei convivium magnum Levi in domo sua et erat turba multa publicanorum et aliorum qui cum illis erant discumbentes
LUKE|5|30|et murmurabant Pharisaei et scribae eorum dicentes ad discipulos eius quare cum publicanis et peccatoribus manducatis et bibitis
LUKE|5|31|et respondens Iesus dixit ad illos non egent qui sani sunt medico sed qui male habent
LUKE|5|32|non veni vocare iustos sed peccatores in paenitentiam
LUKE|5|33|at illi dixerunt ad eum quare discipuli Iohannis ieiunant frequenter et obsecrationes faciunt similiter et Pharisaeorum tui autem edunt et bibunt
LUKE|5|34|quibus ipse ait numquid potestis filios sponsi dum cum illis est sponsus facere ieiunare
LUKE|5|35|venient autem dies et cum ablatus fuerit ab illis sponsus tunc ieiunabunt in illis diebus
LUKE|5|36|dicebat autem et similitudinem ad illos quia nemo commissuram a vestimento novo inmittit in vestimentum vetus alioquin et novum rumpit et veteri non convenit commissura a novo
LUKE|5|37|et nemo mittit vinum novum in utres veteres alioquin rumpet vinum novum utres et ipsum effundetur et utres peribunt
LUKE|5|38|sed vinum novum in utres novos mittendum est et utraque conservantur
LUKE|5|39|et nemo bibens vetus statim vult novum dicit enim vetus melius est
LUKE|6|1|factum est autem in sabbato secundoprimo cum transiret per sata vellebant discipuli eius spicas et manducabant confricantes manibus
LUKE|6|2|quidam autem Pharisaeorum dicebant illis quid facitis quod non licet in sabbatis
LUKE|6|3|et respondens Iesus ad eos dixit nec hoc legistis quod fecit David cum esurisset ipse et qui cum eo erant
LUKE|6|4|quomodo intravit in domum Dei et panes propositionis sumpsit et manducavit et dedit his qui cum ipso erant quos non licet manducare nisi tantum sacerdotibus
LUKE|6|5|et dicebat illis quia dominus est Filius hominis etiam sabbati
LUKE|6|6|factum est autem et in alio sabbato ut intraret in synagogam et doceret et erat ibi homo et manus eius dextra erat arida
LUKE|6|7|observabant autem scribae et Pharisaei si in sabbato curaret ut invenirent accusare illum
LUKE|6|8|ipse vero sciebat cogitationes eorum et ait homini qui habebat manum aridam surge et sta in medium et surgens stetit
LUKE|6|9|ait autem ad illos Iesus interrogo vos si licet sabbato bene facere an male animam salvam facere an perdere
LUKE|6|10|et circumspectis omnibus dixit homini extende manum tuam et extendit et restituta est manus eius
LUKE|6|11|ipsi autem repleti sunt insipientia et conloquebantur ad invicem quidnam facerent Iesu
LUKE|6|12|factum est autem in illis diebus exiit in montem orare et erat pernoctans in oratione Dei
LUKE|6|13|et cum dies factus esset vocavit discipulos suos et elegit duodecim ex ipsis quos et apostolos nominavit
LUKE|6|14|Simonem quem cognominavit Petrum et Andream fratrem eius Iacobum et Iohannem Philippum et Bartholomeum
LUKE|6|15|Mattheum et Thomam Iacobum Alphei et Simonem qui vocatur Zelotes
LUKE|6|16|Iudam Iacobi et Iudam Scarioth qui fuit proditor
LUKE|6|17|et descendens cum illis stetit in loco campestri et turba discipulorum eius et multitudo copiosa plebis ab omni Iudaea et Hierusalem et maritimae Tyri et Sidonis
LUKE|6|18|qui venerunt ut audirent eum et sanarentur a languoribus suis et qui vexabantur ab spiritibus inmundis curabantur
LUKE|6|19|et omnis turba quaerebant eum tangere quia virtus de illo exiebat et sanabat omnes
LUKE|6|20|et ipse elevatis oculis in discipulos suos dicebat beati pauperes quia vestrum est regnum Dei
LUKE|6|21|beati qui nunc esuritis quia saturabimini beati qui nunc fletis quia ridebitis
LUKE|6|22|beati eritis cum vos oderint homines et cum separaverint vos et exprobraverint et eiecerint nomen vestrum tamquam malum propter Filium hominis
LUKE|6|23|gaudete in illa die et exultate ecce enim merces vestra multa in caelo secundum haec enim faciebant prophetis patres eorum
LUKE|6|24|verumtamen vae vobis divitibus quia habetis consolationem vestram
LUKE|6|25|vae vobis qui saturati estis quia esurietis vae vobis qui ridetis nunc quia lugebitis et flebitis
LUKE|6|26|vae cum bene vobis dixerint omnes homines secundum haec faciebant prophetis patres eorum
LUKE|6|27|sed vobis dico qui auditis diligite inimicos vestros benefacite his qui vos oderunt
LUKE|6|28|benedicite maledicentibus vobis orate pro calumniantibus vos
LUKE|6|29|ei qui te percutit in maxillam praebe et alteram et ab eo qui aufert tibi vestimentum etiam tunicam noli prohibere
LUKE|6|30|omni autem petenti te tribue et qui aufert quae tua sunt ne repetas
LUKE|6|31|et prout vultis ut faciant vobis homines et vos facite illis similiter
LUKE|6|32|et si diligitis eos qui vos diligunt quae vobis est gratia nam et peccatores diligentes se diligunt
LUKE|6|33|et si benefeceritis his qui vobis benefaciunt quae vobis est gratia siquidem et peccatores hoc faciunt
LUKE|6|34|et si mutuum dederitis his a quibus speratis recipere quae gratia est vobis nam et peccatores peccatoribus fenerantur ut recipiant aequalia
LUKE|6|35|verumtamen diligite inimicos vestros et benefacite et mutuum date nihil desperantes et erit merces vestra multa et eritis filii Altissimi quia ipse benignus est super ingratos et malos
LUKE|6|36|estote ergo misericordes sicut et Pater vester misericors est
LUKE|6|37|nolite iudicare et non iudicabimini nolite condemnare et non condemnabimini dimittite et dimittemini
LUKE|6|38|date et dabitur vobis mensuram bonam confersam et coagitatam et supereffluentem dabunt in sinum vestrum eadem quippe mensura qua mensi fueritis remetietur vobis
LUKE|6|39|dicebat autem illis et similitudinem numquid potest caecus caecum ducere nonne ambo in foveam cadent
LUKE|6|40|non est discipulus super magistrum perfectus autem omnis erit sicut magister eius
LUKE|6|41|quid autem vides festucam in oculo fratris tui trabem autem quae in oculo tuo est non consideras
LUKE|6|42|et quomodo potes dicere fratri tuo frater sine eiciam festucam de oculo tuo ipse in oculo tuo trabem non videns hypocrita eice primum trabem de oculo tuo et tunc perspicies ut educas festucam de oculo fratris tui
LUKE|6|43|non est enim arbor bona quae facit fructus malos neque arbor mala faciens fructum bonum
LUKE|6|44|unaquaeque enim arbor de fructu suo cognoscitur neque enim de spinis colligunt ficus neque de rubo vindemiant uvam
LUKE|6|45|bonus homo de bono thesauro cordis sui profert bonum et malus homo de malo profert malum ex abundantia enim cordis os loquitur
LUKE|6|46|quid autem vocatis me Domine Domine et non facitis quae dico
LUKE|6|47|omnis qui venit ad me et audit sermones meos et facit eos ostendam vobis cui similis est
LUKE|6|48|similis est homini aedificanti domum qui fodit in altum et posuit fundamenta supra petram inundatione autem facta inlisum est flumen domui illi et non potuit eam movere fundata enim erat supra petram
LUKE|6|49|qui autem audivit et non fecit similis est homini aedificanti domum suam supra terram sine fundamento in quam inlisus est fluvius et continuo concidit et facta est ruina domus illius magna
LUKE|7|1|cum autem implesset omnia verba sua in aures plebis intravit Capharnaum
LUKE|7|2|centurionis autem cuiusdam servus male habens erat moriturus qui illi erat pretiosus
LUKE|7|3|et cum audisset de Iesu misit ad eum seniores Iudaeorum rogans eum ut veniret et salvaret servum eius
LUKE|7|4|at illi cum venissent ad Iesum rogabant eum sollicite dicentes ei quia dignus est ut hoc illi praestes
LUKE|7|5|diligit enim gentem nostram et synagogam ipse aedificavit nobis
LUKE|7|6|Iesus autem ibat cum illis et cum iam non longe esset a domo misit ad eum centurio amicos dicens Domine noli vexari non enim dignus sum ut sub tectum meum intres
LUKE|7|7|propter quod et me ipsum non sum dignum arbitratus ut venirem ad te sed dic verbo et sanabitur puer meus
LUKE|7|8|nam et ego homo sum sub potestate constitutus habens sub me milites et dico huic vade et vadit et alio veni et venit et servo meo fac hoc et facit
LUKE|7|9|quo audito Iesus miratus est et conversus sequentibus se turbis dixit amen dico vobis nec in Israhel tantam fidem inveni
LUKE|7|10|et reversi qui missi fuerant domum invenerunt servum qui languerat sanum
LUKE|7|11|et factum est deinceps ibat in civitatem quae vocatur Naim et ibant cum illo discipuli eius et turba copiosa
LUKE|7|12|cum autem adpropinquaret portae civitatis et ecce defunctus efferebatur filius unicus matri suae et haec vidua erat et turba civitatis multa cum illa
LUKE|7|13|quam cum vidisset Dominus misericordia motus super ea dixit illi noli flere
LUKE|7|14|et accessit et tetigit loculum hii autem qui portabant steterunt et ait adulescens tibi dico surge
LUKE|7|15|et resedit qui erat mortuus et coepit loqui et dedit illum matri suae
LUKE|7|16|accepit autem omnes timor et magnificabant Deum dicentes quia propheta magnus surrexit in nobis et quia Deus visitavit plebem suam
LUKE|7|17|et exiit hic sermo in universam Iudaeam de eo et omnem circa regionem
LUKE|7|18|et nuntiaverunt Iohanni discipuli eius de omnibus his
LUKE|7|19|et convocavit duos de discipulis suis Iohannes et misit ad Dominum dicens tu es qui venturus es an alium expectamus
LUKE|7|20|cum autem venissent ad eum viri dixerunt Iohannes Baptista misit nos ad te dicens tu es qui venturus es an alium expectamus
LUKE|7|21|in ipsa autem hora curavit multos a languoribus et plagis et spiritibus malis et caecis multis donavit visum
LUKE|7|22|et respondens dixit illis euntes nuntiate Iohanni quae vidistis et audistis quia caeci vident claudi ambulant leprosi mundantur surdi audiunt mortui resurgunt pauperes evangelizantur
LUKE|7|23|et beatus est quicumque non fuerit scandalizatus in me
LUKE|7|24|et cum discessissent nuntii Iohannis coepit dicere de Iohanne ad turbas quid existis in desertum videre harundinem vento moveri
LUKE|7|25|sed quid existis videre hominem mollibus vestimentis indutum ecce qui in veste pretiosa sunt et deliciis in domibus regum sunt
LUKE|7|26|sed quid existis videre prophetam utique dico vobis et plus quam prophetam
LUKE|7|27|hic est de quo scriptum est ecce mitto angelum meum ante faciem tuam qui praeparabit viam tuam ante te
LUKE|7|28|dico enim vobis maior inter natos mulierum propheta Iohanne Baptista nemo est qui autem minor est in regno Dei maior est illo
LUKE|7|29|et omnis populus audiens et publicani iustificaverunt Deum baptizati baptismo Iohannis
LUKE|7|30|Pharisaei autem et legis periti consilium Dei spreverunt in semet ipsos non baptizati ab eo
LUKE|7|31|cui ergo similes dicam homines generationis huius et cui similes sunt
LUKE|7|32|similes sunt pueris sedentibus in foro et loquentibus ad invicem et dicentibus cantavimus vobis tibiis et non saltastis lamentavimus et non plorastis
LUKE|7|33|venit enim Iohannes Baptista neque manducans panem neque bibens vinum et dicitis daemonium habet
LUKE|7|34|venit Filius hominis manducans et bibens et dicitis ecce homo devorator et bibens vinum amicus publicanorum et peccatorum
LUKE|7|35|et iustificata est sapientia ab omnibus filiis suis
LUKE|7|36|rogabat autem illum quidam de Pharisaeis ut manducaret cum illo et ingressus domum Pharisaei discubuit
LUKE|7|37|et ecce mulier quae erat in civitate peccatrix ut cognovit quod accubuit in domo Pharisaei adtulit alabastrum unguenti
LUKE|7|38|et stans retro secus pedes eius lacrimis coepit rigare pedes eius et capillis capitis sui tergebat et osculabatur pedes eius et unguento unguebat
LUKE|7|39|videns autem Pharisaeus qui vocaverat eum ait intra se dicens hic si esset propheta sciret utique quae et qualis mulier quae tangit eum quia peccatrix est
LUKE|7|40|et respondens Iesus dixit ad illum Simon habeo tibi aliquid dicere at ille ait magister dic
LUKE|7|41|duo debitores erant cuidam feneratori unus debebat denarios quingentos alius quinquaginta
LUKE|7|42|non habentibus illis unde redderent donavit utrisque quis ergo eum plus diliget
LUKE|7|43|respondens Simon dixit aestimo quia is cui plus donavit at ille dixit ei recte iudicasti
LUKE|7|44|et conversus ad mulierem dixit Simoni vides hanc mulierem intravi in domum tuam aquam pedibus meis non dedisti haec autem lacrimis rigavit pedes meos et capillis suis tersit
LUKE|7|45|osculum mihi non dedisti haec autem ex quo intravit non cessavit osculari pedes meos
LUKE|7|46|oleo caput meum non unxisti haec autem unguento unxit pedes meos
LUKE|7|47|propter quod dico tibi remittentur ei peccata multa quoniam dilexit multum cui autem minus dimittitur minus diligit
LUKE|7|48|dixit autem ad illam remittuntur tibi peccata
LUKE|7|49|et coeperunt qui simul accumbebant dicere intra se quis est hic qui etiam peccata dimittit
LUKE|7|50|dixit autem ad mulierem fides tua te salvam fecit vade in pace
LUKE|8|1|et factum est deinceps et ipse iter faciebat per civitatem et castellum praedicans et evangelizans regnum Dei et duodecim cum illo
LUKE|8|2|et mulieres aliquae quae erant curatae ab spiritibus malignis et infirmitatibus Maria quae vocatur Magdalene de qua daemonia septem exierant
LUKE|8|3|et Iohanna uxor Chuza procuratoris Herodis et Susanna et aliae multae quae ministrabant eis de facultatibus suis
LUKE|8|4|cum autem turba plurima conveniret et de civitatibus properarent ad eum dixit per similitudinem
LUKE|8|5|exiit qui seminat seminare semen suum et dum seminat aliud cecidit secus viam et conculcatum est et volucres caeli comederunt illud
LUKE|8|6|et aliud cecidit supra petram et natum aruit quia non habebat humorem
LUKE|8|7|et aliud cecidit inter spinas et simul exortae spinae suffocaverunt illud
LUKE|8|8|et aliud cecidit in terram bonam et ortum fecit fructum centuplum haec dicens clamabat qui habet aures audiendi audiat
LUKE|8|9|interrogabant autem eum discipuli eius quae esset haec parabola
LUKE|8|10|quibus ipse dixit vobis datum est nosse mysterium regni Dei ceteris autem in parabolis ut videntes non videant et audientes non intellegant
LUKE|8|11|est autem haec parabola semen est verbum Dei
LUKE|8|12|qui autem secus viam sunt qui audiunt deinde venit diabolus et tollit verbum de corde eorum ne credentes salvi fiant
LUKE|8|13|nam qui supra petram qui cum audierint cum gaudio suscipiunt verbum et hii radices non habent qui ad tempus credunt et in tempore temptationis recedunt
LUKE|8|14|quod autem in spinis cecidit hii sunt qui audierunt et a sollicitudinibus et divitiis et voluptatibus vitae euntes suffocantur et non referunt fructum
LUKE|8|15|quod autem in bonam terram hii sunt qui in corde bono et optimo audientes verbum retinent et fructum adferunt in patientia
LUKE|8|16|nemo autem lucernam accendens operit eam vaso aut subtus lectum ponit sed supra candelabrum ponit ut intrantes videant lumen
LUKE|8|17|non enim est occultum quod non manifestetur nec absconditum quod non cognoscatur et in palam veniat
LUKE|8|18|videte ergo quomodo auditis qui enim habet dabitur illi et quicumque non habet etiam quod putat se habere auferetur ab illo
LUKE|8|19|venerunt autem ad illum mater et fratres eius et non poterant adire ad eum prae turba
LUKE|8|20|et nuntiatum est illi mater tua et fratres tui stant foris volentes te videre
LUKE|8|21|qui respondens dixit ad eos mater mea et fratres mei hii sunt qui verbum Dei audiunt et faciunt
LUKE|8|22|factum est autem in una dierum et ipse ascendit in naviculam et discipuli eius et ait ad illos transfretemus trans stagnum et ascenderunt
LUKE|8|23|navigantibus autem illis obdormiit et descendit procella venti in stagnum et conplebantur et periclitabantur
LUKE|8|24|accedentes autem suscitaverunt eum dicentes praeceptor perimus at ille surgens increpavit ventum et tempestatem aquae et cessavit et facta est tranquillitas
LUKE|8|25|dixit autem illis ubi est fides vestra qui timentes mirati sunt dicentes ad invicem quis putas hic est quia et ventis imperat et mari et oboediunt ei
LUKE|8|26|enavigaverunt autem ad regionem Gerasenorum quae est contra Galilaeam
LUKE|8|27|et cum egressus esset ad terram occurrit illi vir quidam qui habebat daemonium iam temporibus multis et vestimento non induebatur neque in domo manebat sed in monumentis
LUKE|8|28|is ut vidit Iesum procidit ante illum et exclamans voce magna dixit quid mihi et tibi est Iesu Fili Dei altissimi obsecro te ne me torqueas
LUKE|8|29|praecipiebat enim spiritui inmundo ut exiret ab homine multis enim temporibus arripiebat illum et vinciebatur catenis et conpedibus custoditus et ruptis vinculis agebatur a daemonio in deserta
LUKE|8|30|interrogavit autem illum Iesus dicens quod tibi nomen est at ille dixit Legio quia intraverunt daemonia multa in eum
LUKE|8|31|et rogabant illum ne imperaret illis ut in abyssum irent
LUKE|8|32|erat autem ibi grex porcorum multorum pascentium in monte et rogabant eum ut permitteret eos in illos ingredi et permisit illos
LUKE|8|33|exierunt ergo daemonia ab homine et intraverunt in porcos et impetu abiit grex per praeceps in stagnum et suffocatus est
LUKE|8|34|quod ut viderunt factum qui pascebant fugerunt et nuntiaverunt in civitatem et in villas
LUKE|8|35|exierunt autem videre quod factum est et venerunt ad Iesum et invenerunt hominem sedentem a quo daemonia exierant vestitum ac sana mente ad pedes eius et timuerunt
LUKE|8|36|nuntiaverunt autem illis et qui viderant quomodo sanus factus esset a Legione
LUKE|8|37|et rogaverunt illum omnis multitudo regionis Gerasenorum ut discederet ab ipsis quia timore magno tenebantur ipse autem ascendens navem reversus est
LUKE|8|38|et rogabat illum vir a quo daemonia exierant ut cum eo esset dimisit autem eum Iesus dicens
LUKE|8|39|redi domum tuam et narra quanta tibi fecit Deus et abiit per universam civitatem praedicans quanta illi fecisset Iesus
LUKE|8|40|factum est autem cum redisset Iesus excepit illum turba erant enim omnes expectantes eum
LUKE|8|41|et ecce venit vir cui nomen Iairus et ipse princeps synagogae erat et cecidit ad pedes Iesu rogans eum ut intraret in domum eius
LUKE|8|42|quia filia unica erat illi fere annorum duodecim et haec moriebatur et contigit dum iret a turbis conprimebatur
LUKE|8|43|et mulier quaedam erat in fluxu sanguinis ab annis duodecim quae in medicos erogaverat omnem substantiam suam nec ab ullo potuit curari
LUKE|8|44|accessit retro et tetigit fimbriam vestimenti eius et confestim stetit fluxus sanguinis eius
LUKE|8|45|et ait Iesus quis est qui me tetigit negantibus autem omnibus dixit Petrus et qui cum illo erant praeceptor turbae te conprimunt et adfligunt et dicis quis me tetigit
LUKE|8|46|et dixit Iesus tetigit me aliquis nam ego novi virtutem de me exisse
LUKE|8|47|videns autem mulier quia non latuit tremens venit et procidit ante pedes illius et ob quam causam tetigerit eum indicavit coram omni populo et quemadmodum confestim sanata sit
LUKE|8|48|at ipse dixit illi filia fides tua te salvam fecit vade in pace
LUKE|8|49|adhuc illo loquente venit a principe synagogae dicens ei quia mortua est filia tua noli vexare illum
LUKE|8|50|Iesus autem audito hoc verbo respondit patri puellae noli timere crede tantum et salva erit
LUKE|8|51|et cum venisset domum non permisit intrare secum quemquam nisi Petrum et Iohannem et Iacobum et patrem et matrem puellae
LUKE|8|52|flebant autem omnes et plangebant illam at ille dixit nolite flere non est mortua sed dormit
LUKE|8|53|et deridebant eum scientes quia mortua esset
LUKE|8|54|ipse autem tenens manum eius clamavit dicens puella surge
LUKE|8|55|et reversus est spiritus eius et surrexit continuo et iussit illi dari manducare
LUKE|8|56|et stupuerunt parentes eius quibus praecepit ne alicui dicerent quod factum erat
LUKE|9|1|convocatis autem duodecim apostolis dedit illis virtutem et potestatem super omnia daemonia et ut languores curarent
LUKE|9|2|et misit illos praedicare regnum Dei et sanare infirmos
LUKE|9|3|et ait ad illos nihil tuleritis in via neque virgam neque peram neque panem neque pecuniam neque duas tunicas habeatis
LUKE|9|4|et in quamcumque domum intraveritis ibi manete et inde ne exeatis
LUKE|9|5|et quicumque non receperint vos exeuntes de civitate illa etiam pulverem pedum vestrorum excutite in testimonium supra illos
LUKE|9|6|egressi autem circumibant per castella evangelizantes et curantes ubique
LUKE|9|7|audivit autem Herodes tetrarcha omnia quae fiebant ab eo et haesitabat eo quod diceretur
LUKE|9|8|a quibusdam quia Iohannes surrexit a mortuis a quibusdam vero quia Helias apparuit ab aliis autem quia propheta unus de antiquis surrexit
LUKE|9|9|et ait Herodes Iohannem ego decollavi quis autem est iste de quo audio ego talia et quaerebat videre eum
LUKE|9|10|et reversi apostoli narraverunt illi quaecumque fecerunt et adsumptis illis secessit seorsum in locum desertum qui est Bethsaida
LUKE|9|11|quod cum cognovissent turbae secutae sunt illum et excepit illos et loquebatur illis de regno Dei et eos qui cura indigebant sanabat
LUKE|9|12|dies autem coeperat declinare et accedentes duodecim dixerunt illi dimitte turbas ut euntes in castella villasque quae circa sunt devertant et inveniant escas quia hic in loco deserto sumus
LUKE|9|13|ait autem ad illos vos date illis manducare at illi dixerunt non sunt nobis plus quam quinque panes et duo pisces nisi forte nos eamus et emamus in omnem hanc turbam escas
LUKE|9|14|erant autem fere viri quinque milia ait autem ad discipulos suos facite illos discumbere per convivia quinquagenos
LUKE|9|15|et ita fecerunt et discumbere fecerunt omnes
LUKE|9|16|acceptis autem quinque panibus et duobus piscibus respexit in caelum et benedixit illis et fregit et distribuit discipulis suis ut ponerent ante turbas
LUKE|9|17|et manducaverunt omnes et saturati sunt et sublatum est quod superfuit illis fragmentorum cofini duodecim
LUKE|9|18|et factum est cum solus esset orans erant cum illo et discipuli et interrogavit illos dicens quem me dicunt esse turbae
LUKE|9|19|at illi responderunt et dixerunt Iohannem Baptistam alii autem Heliam alii quia propheta unus de prioribus surrexit
LUKE|9|20|dixit autem illis vos autem quem me esse dicitis respondens Simon Petrus dixit Christum Dei
LUKE|9|21|at ille increpans illos praecepit ne cui dicerent hoc
LUKE|9|22|dicens quia oportet Filium hominis multa pati et reprobari a senioribus et principibus sacerdotum et scribis et occidi et tertia die resurgere
LUKE|9|23|dicebat autem ad omnes si quis vult post me venire abneget se ipsum et tollat crucem suam cotidie et sequatur me
LUKE|9|24|qui enim voluerit animam suam salvam facere perdet illam nam qui perdiderit animam suam propter me salvam faciet illam
LUKE|9|25|quid enim proficit homo si lucretur universum mundum se autem ipsum perdat et detrimentum sui faciat
LUKE|9|26|nam qui me erubuerit et meos sermones hunc Filius hominis erubescet cum venerit in maiestate sua et Patris et sanctorum angelorum
LUKE|9|27|dico autem vobis vere sunt aliqui hic stantes qui non gustabunt mortem donec videant regnum Dei
LUKE|9|28|factum est autem post haec verba fere dies octo et adsumpsit Petrum et Iohannem et Iacobum et ascendit in montem ut oraret
LUKE|9|29|et factum est dum oraret species vultus eius altera et vestitus eius albus refulgens
LUKE|9|30|et ecce duo viri loquebantur cum illo erant autem Moses et Helias
LUKE|9|31|visi in maiestate et dicebant excessum eius quem conpleturus erat in Hierusalem
LUKE|9|32|Petrus vero et qui cum illo gravati erant somno et evigilantes viderunt maiestatem eius et duos viros qui stabant cum illo
LUKE|9|33|et factum est cum discederent ab illo ait Petrus ad Iesum praeceptor bonum est nos hic esse et faciamus tria tabernacula unum tibi et unum Mosi et unum Heliae nesciens quid diceret
LUKE|9|34|haec autem illo loquente facta est nubes et obumbravit eos et timuerunt intrantibus illis in nubem
LUKE|9|35|et vox facta est de nube dicens hic est Filius meus electus ipsum audite
LUKE|9|36|et dum fieret vox inventus est Iesus solus et ipsi tacuerunt et nemini dixerunt in illis diebus quicquam ex his quae viderant
LUKE|9|37|factum est autem in sequenti die descendentibus illis de monte occurrit illi turba multa
LUKE|9|38|et ecce vir de turba exclamavit dicens magister obsecro te respice in filium meum quia unicus est mihi
LUKE|9|39|et ecce spiritus adprehendit illum et subito clamat et elidit et dissipat eum cum spuma et vix discedit dilanians eum
LUKE|9|40|et rogavi discipulos tuos ut eicerent illum et non potuerunt
LUKE|9|41|respondens autem Iesus dixit o generatio infidelis et perversa usquequo ero apud vos et patiar vos adduc huc filium tuum
LUKE|9|42|et cum accederet elisit illum daemonium et dissipavit
LUKE|9|43|et increpavit Iesus spiritum inmundum et sanavit puerum et reddidit illum patri eius
LUKE|9|44|stupebant autem omnes in magnitudine Dei omnibusque mirantibus in omnibus quae faciebat dixit ad discipulos suos ponite vos in cordibus vestris sermones istos Filius enim hominis futurum est ut tradatur in manus hominum
LUKE|9|45|at illi ignorabant verbum istud et erat velatum ante eos ut non sentirent illud et timebant interrogare eum de hoc verbo
LUKE|9|46|intravit autem cogitatio in eos quis eorum maior esset
LUKE|9|47|at Iesus videns cogitationes cordis illorum adprehendens puerum statuit eum secus se
LUKE|9|48|et ait illis quicumque susceperit puerum istum in nomine meo me recipit et quicumque me recipit recipit eum qui me misit nam qui minor est inter omnes vos hic maior est
LUKE|9|49|respondens autem Iohannes dixit praeceptor vidimus quendam in nomine tuo eicientem daemonia et prohibuimus eum quia non sequitur nobiscum
LUKE|9|50|et ait ad illum Iesus nolite prohibere qui enim non est adversum vos pro vobis est
LUKE|9|51|factum est autem dum conplerentur dies adsumptionis eius et ipse faciem suam firmavit ut iret Hierusalem
LUKE|9|52|et misit nuntios ante conspectum suum et euntes intraverunt in civitatem Samaritanorum ut pararent illi
LUKE|9|53|et non receperunt eum quia facies eius erat euntis Hierusalem
LUKE|9|54|cum vidissent autem discipuli eius Iacobus et Iohannes dixerunt Domine vis dicimus ut ignis descendat de caelo et consumat illos
LUKE|9|55|et conversus increpavit illos
LUKE|9|56|et abierunt in aliud castellum
LUKE|9|57|factum est autem ambulantibus illis in via dixit quidam ad illum sequar te quocumque ieris
LUKE|9|58|et ait illi Iesus vulpes foveas habent et volucres caeli nidos Filius autem hominis non habet ubi caput reclinet
LUKE|9|59|ait autem ad alterum sequere me ille autem dixit Domine permitte mihi primum ire sepelire patrem meum
LUKE|9|60|dixitque ei Iesus sine ut mortui sepeliant mortuos suos tu autem vade adnuntia regnum Dei
LUKE|9|61|et ait alter sequar te Domine sed primum permitte mihi renuntiare his qui domi sunt
LUKE|9|62|ait ad illum Iesus nemo mittens manum suam in aratrum et aspiciens retro aptus est regno Dei
LUKE|10|1|post haec autem designavit Dominus et alios septuaginta duos et misit illos binos ante faciem suam in omnem civitatem et locum quo erat ipse venturus
LUKE|10|2|et dicebat illis messis quidem multa operarii autem pauci rogate ergo Dominum messis ut mittat operarios in messem
LUKE|10|3|ite ecce ego mitto vos sicut agnos inter lupos
LUKE|10|4|nolite portare sacculum neque peram neque calciamenta et neminem per viam salutaveritis
LUKE|10|5|in quamcumque domum intraveritis primum dicite pax huic domui
LUKE|10|6|et si ibi fuerit filius pacis requiescet super illam pax vestra sin autem ad vos revertetur
LUKE|10|7|in eadem autem domo manete edentes et bibentes quae apud illos sunt dignus enim est operarius mercede sua nolite transire de domo in domum
LUKE|10|8|et in quamcumque civitatem intraveritis et susceperint vos manducate quae adponuntur vobis
LUKE|10|9|et curate infirmos qui in illa sunt et dicite illis adpropinquavit in vos regnum Dei
LUKE|10|10|in quamcumque civitatem intraveritis et non receperint vos exeuntes in plateas eius dicite
LUKE|10|11|etiam pulverem qui adhesit nobis de civitate vestra extergimus in vos tamen hoc scitote quia adpropinquavit regnum Dei
LUKE|10|12|dico vobis quia Sodomis in die illa remissius erit quam illi civitati
LUKE|10|13|vae tibi Corazain vae tibi Bethsaida quia si in Tyro et Sidone factae fuissent virtutes quae in vobis factae sunt olim in cilicio et cinere sedentes paeniterent
LUKE|10|14|verumtamen Tyro et Sidoni remissius erit in iudicio quam vobis
LUKE|10|15|et tu Capharnaum usque in caelum exaltata usque ad infernum demergeris
LUKE|10|16|qui vos audit me audit et qui vos spernit me spernit qui autem me spernit spernit eum qui me misit
LUKE|10|17|reversi sunt autem septuaginta duo cum gaudio dicentes Domine etiam daemonia subiciuntur nobis in nomine tuo
LUKE|10|18|et ait illis videbam Satanan sicut fulgur de caelo cadentem
LUKE|10|19|ecce dedi vobis potestatem calcandi supra serpentes et scorpiones et supra omnem virtutem inimici et nihil vobis nocebit
LUKE|10|20|verumtamen in hoc nolite gaudere quia spiritus vobis subiciuntur gaudete autem quod nomina vestra scripta sunt in caelis
LUKE|10|21|in ipsa hora exultavit Spiritu Sancto et dixit confiteor tibi Pater Domine caeli et terrae quod abscondisti haec a sapientibus et prudentibus et revelasti ea parvulis etiam Pater quia sic placuit ante te
LUKE|10|22|omnia mihi tradita sunt a Patre meo et nemo scit qui sit Filius nisi Pater et qui sit Pater nisi Filius et cui voluerit Filius revelare
LUKE|10|23|et conversus ad discipulos suos dixit beati oculi qui vident quae videtis
LUKE|10|24|dico enim vobis quod multi prophetae et reges voluerunt videre quae vos videtis et non viderunt et audire quae auditis et non audierunt
LUKE|10|25|et ecce quidam legis peritus surrexit temptans illum et dicens magister quid faciendo vitam aeternam possidebo
LUKE|10|26|at ille dixit ad eum in lege quid scriptum est quomodo legis
LUKE|10|27|ille respondens dixit diliges Dominum Deum tuum ex toto corde tuo et ex tota anima tua et ex omnibus viribus tuis et ex omni mente tua et proximum tuum sicut te ipsum
LUKE|10|28|dixitque illi recte respondisti hoc fac et vives
LUKE|10|29|ille autem volens iustificare se ipsum dixit ad Iesum et quis est meus proximus
LUKE|10|30|suscipiens autem Iesus dixit homo quidam descendebat ab Hierusalem in Hiericho et incidit in latrones qui etiam despoliaverunt eum et plagis inpositis abierunt semivivo relicto
LUKE|10|31|accidit autem ut sacerdos quidam descenderet eadem via et viso illo praeterivit
LUKE|10|32|similiter et Levita cum esset secus locum et videret eum pertransiit
LUKE|10|33|Samaritanus autem quidam iter faciens venit secus eum et videns eum misericordia motus est
LUKE|10|34|et adpropians alligavit vulnera eius infundens oleum et vinum et inponens illum in iumentum suum duxit in stabulum et curam eius egit
LUKE|10|35|et altera die protulit duos denarios et dedit stabulario et ait curam illius habe et quodcumque supererogaveris ego cum rediero reddam tibi
LUKE|10|36|quis horum trium videtur tibi proximus fuisse illi qui incidit in latrones
LUKE|10|37|at ille dixit qui fecit misericordiam in illum et ait illi Iesus vade et tu fac similiter
LUKE|10|38|factum est autem dum irent et ipse intravit in quoddam castellum et mulier quaedam Martha nomine excepit illum in domum suam
LUKE|10|39|et huic erat soror nomine Maria quae etiam sedens secus pedes Domini audiebat verbum illius
LUKE|10|40|Martha autem satagebat circa frequens ministerium quae stetit et ait Domine non est tibi curae quod soror mea reliquit me solam ministrare dic ergo illi ut me adiuvet
LUKE|10|41|et respondens dixit illi Dominus Martha Martha sollicita es et turbaris erga plurima
LUKE|10|42|porro unum est necessarium Maria optimam partem elegit quae non auferetur ab ea
LUKE|11|1|et factum est cum esset in loco quodam orans ut cessavit dixit unus ex discipulis eius ad eum Domine doce nos orare sicut et Iohannes docuit discipulos suos
LUKE|11|2|et ait illis cum oratis dicite Pater sanctificetur nomen tuum adveniat regnum tuum
LUKE|11|3|panem nostrum cotidianum da nobis cotidie
LUKE|11|4|et dimitte nobis peccata nostra siquidem et ipsi dimittimus omni debenti nobis et ne nos inducas in temptationem
LUKE|11|5|et ait ad illos quis vestrum habebit amicum et ibit ad illum media nocte et dicit illi amice commoda mihi tres panes
LUKE|11|6|quoniam amicus meus venit de via ad me et non habeo quod ponam ante illum
LUKE|11|7|et ille de intus respondens dicat noli mihi molestus esse iam ostium clausum est et pueri mei mecum sunt in cubili non possum surgere et dare tibi
LUKE|11|8|dico vobis et si non dabit illi surgens eo quod amicus eius sit propter inprobitatem tamen eius surget et dabit illi quotquot habet necessarios
LUKE|11|9|et ego vobis dico petite et dabitur vobis quaerite et invenietis pulsate et aperietur vobis
LUKE|11|10|omnis enim qui petit accipit et qui quaerit invenit et pulsanti aperietur
LUKE|11|11|quis autem ex vobis patrem petet panem numquid lapidem dabit illi aut piscem numquid pro pisce serpentem dabit illi
LUKE|11|12|aut si petierit ovum numquid porriget illi scorpionem
LUKE|11|13|si ergo vos cum sitis mali nostis bona data dare filiis vestris quanto magis Pater vester de caelo dabit spiritum bonum petentibus se
LUKE|11|14|et erat eiciens daemonium et illud erat mutum et cum eiecisset daemonium locutus est mutus et admiratae sunt turbae
LUKE|11|15|quidam autem ex eis dixerunt in Beelzebub principe daemoniorum eicit daemonia
LUKE|11|16|et alii temptantes signum de caelo quaerebant ab eo
LUKE|11|17|ipse autem ut vidit cogitationes eorum dixit eis omne regnum in se ipsum divisum desolatur et domus supra domum cadet
LUKE|11|18|si autem et Satanas in se ipsum divisus est quomodo stabit regnum ipsius quia dicitis in Beelzebub eicere me daemonia
LUKE|11|19|si autem ego in Beelzebub eicio daemonia filii vestri in quo eiciunt ideo ipsi iudices vestri erunt
LUKE|11|20|porro si in digito Dei eicio daemonia profecto praevenit in vos regnum Dei
LUKE|11|21|cum fortis armatus custodit atrium suum in pace sunt ea quae possidet
LUKE|11|22|si autem fortior illo superveniens vicerit eum universa arma eius aufert in quibus confidebat et spolia eius distribuit
LUKE|11|23|qui non est mecum adversum me est et qui non colligit mecum dispergit
LUKE|11|24|cum inmundus spiritus exierit de homine perambulat per loca inaquosa quaerens requiem et non inveniens dicit revertar in domum meam unde exivi
LUKE|11|25|et cum venerit invenit scopis mundatam
LUKE|11|26|et tunc vadit et adsumit septem alios spiritus nequiores se et ingressi habitant ibi et sunt novissima hominis illius peiora prioribus
LUKE|11|27|factum est autem cum haec diceret extollens vocem quaedam mulier de turba dixit illi beatus venter qui te portavit et ubera quae suxisti
LUKE|11|28|at ille dixit quippini beati qui audiunt verbum Dei et custodiunt
LUKE|11|29|turbis autem concurrentibus coepit dicere generatio haec generatio nequam est signum quaerit et signum non dabitur illi nisi signum Ionae
LUKE|11|30|nam sicut Ionas fuit signum Ninevitis ita erit et Filius hominis generationi isti
LUKE|11|31|regina austri surget in iudicio cum viris generationis huius et condemnabit illos quia venit a finibus terrae audire sapientiam Salomonis et ecce plus Salomone hic
LUKE|11|32|viri ninevitae surgent in iudicio cum generatione hac et condemnabunt illam quia paenitentiam egerunt ad praedicationem Ionae et ecce plus Iona hic
LUKE|11|33|nemo lucernam accendit et in abscondito ponit neque sub modio sed supra candelabrum ut qui ingrediuntur lumen videant
LUKE|11|34|lucerna corporis tui est oculus tuus si oculus tuus fuerit simplex totum corpus tuum lucidum erit si autem nequam fuerit etiam corpus tuum tenebrosum erit
LUKE|11|35|vide ergo ne lumen quod in te est tenebrae sint
LUKE|11|36|si ergo corpus tuum totum lucidum fuerit non habens aliquam partem tenebrarum erit lucidum totum et sicut lucerna fulgoris inluminabit te
LUKE|11|37|et cum loqueretur rogavit illum quidam Pharisaeus ut pranderet apud se et ingressus recubuit
LUKE|11|38|Pharisaeus autem coepit intra se reputans dicere quare non baptizatus esset ante prandium
LUKE|11|39|et ait Dominus ad illum nunc vos Pharisaei quod de foris est calicis et catini mundatis quod autem intus est vestrum plenum est rapina et iniquitate
LUKE|11|40|stulti nonne qui fecit quod de foris est etiam id quod de intus est fecit
LUKE|11|41|verumtamen quod superest date elemosynam et ecce omnia munda sunt vobis
LUKE|11|42|sed vae vobis Pharisaeis quia decimatis mentam et rutam et omne holus et praeteritis iudicium et caritatem Dei haec autem oportuit facere et illa non omittere
LUKE|11|43|vae vobis Pharisaeis quia diligitis primas cathedras in synagogis et salutationes in foro
LUKE|11|44|vae vobis quia estis ut monumenta quae non parent et homines ambulantes supra nesciunt
LUKE|11|45|respondens autem quidam ex legis peritis ait illi magister haec dicens etiam nobis contumeliam facis
LUKE|11|46|at ille ait et vobis legis peritis vae quia oneratis homines oneribus quae portari non possunt et ipsi uno digito vestro non tangitis sarcinas
LUKE|11|47|vae vobis quia aedificatis monumenta prophetarum patres autem vestri occiderunt illos
LUKE|11|48|profecto testificamini quod consentitis operibus patrum vestrorum quoniam quidem ipsi eos occiderunt vos autem aedificatis eorum sepulchra
LUKE|11|49|propterea et sapientia Dei dixit mittam ad illos prophetas et apostolos et ex illis occident et persequentur
LUKE|11|50|ut inquiratur sanguis omnium prophetarum qui effusus est a constitutione mundi a generatione ista
LUKE|11|51|a sanguine Abel usque ad sanguinem Zacchariae qui periit inter altare et aedem ita dico vobis requiretur ab hac generatione
LUKE|11|52|vae vobis legis peritis quia tulistis clavem scientiae ipsi non introistis et eos qui introibant prohibuistis
LUKE|11|53|cum haec ad illos diceret coeperunt Pharisaei et legis periti graviter insistere et os eius opprimere de multis
LUKE|11|54|insidiantes et quaerentes capere aliquid ex ore eius ut accusarent eum
LUKE|12|1|multis autem turbis circumstantibus ita ut se invicem conculcarent coepit dicere ad discipulos suos adtendite a fermento Pharisaeorum quae est hypocrisis
LUKE|12|2|nihil autem opertum est quod non reveletur neque absconditum quod non sciatur
LUKE|12|3|quoniam quae in tenebris dixistis in lumine dicentur et quod in aurem locuti estis in cubiculis praedicabitur in tectis
LUKE|12|4|dico autem vobis amicis meis ne terreamini ab his qui occidunt corpus et post haec non habent amplius quod faciant
LUKE|12|5|ostendam autem vobis quem timeatis timete eum qui postquam occiderit habet potestatem mittere in gehennam ita dico vobis hunc timete
LUKE|12|6|nonne quinque passeres veneunt dipundio et unus ex illis non est in oblivione coram Deo
LUKE|12|7|sed et capilli capitis vestri omnes numerati sunt nolite ergo timere multis passeribus pluris estis
LUKE|12|8|dico autem vobis omnis quicumque confessus fuerit in me coram hominibus et Filius hominis confitebitur in illo coram angelis Dei
LUKE|12|9|qui autem negaverit me coram hominibus denegabitur coram angelis Dei
LUKE|12|10|et omnis qui dicit verbum in Filium hominis remittetur illi ei autem qui in Spiritum Sanctum blasphemaverit non remittetur
LUKE|12|11|cum autem inducent vos in synagogas et ad magistratus et potestates nolite solliciti esse qualiter aut quid respondeatis aut quid dicatis
LUKE|12|12|Spiritus enim Sanctus docebit vos in ipsa hora quae oporteat dicere
LUKE|12|13|ait autem quidam ei de turba magister dic fratri meo ut dividat mecum hereditatem
LUKE|12|14|at ille dixit ei homo quis me constituit iudicem aut divisorem super vos
LUKE|12|15|dixitque ad illos videte et cavete ab omni avaritia quia non in abundantia cuiusquam vita eius est ex his quae possidet
LUKE|12|16|dixit autem similitudinem ad illos dicens hominis cuiusdam divitis uberes fructus ager adtulit
LUKE|12|17|et cogitabat intra se dicens quid faciam quod non habeo quo congregem fructus meos
LUKE|12|18|et dixit hoc faciam destruam horrea mea et maiora faciam et illuc congregabo omnia quae nata sunt mihi et bona mea
LUKE|12|19|et dicam animae meae anima habes multa bona posita in annos plurimos requiesce comede bibe epulare
LUKE|12|20|dixit autem illi Deus stulte hac nocte animam tuam repetunt a te quae autem parasti cuius erunt
LUKE|12|21|sic est qui sibi thesaurizat et non est in Deum dives
LUKE|12|22|dixitque ad discipulos suos ideo dico vobis nolite solliciti esse animae quid manducetis neque corpori quid vestiamini
LUKE|12|23|anima plus est quam esca et corpus quam vestimentum
LUKE|12|24|considerate corvos quia non seminant neque metunt quibus non est cellarium neque horreum et Deus pascit illos quanto magis vos pluris estis illis
LUKE|12|25|quis autem vestrum cogitando potest adicere ad staturam suam cubitum unum
LUKE|12|26|si ergo neque quod minimum est potestis quid de ceteris solliciti estis
LUKE|12|27|considerate lilia quomodo crescunt non laborant non nent dico autem vobis nec Salomon in omni gloria sua vestiebatur sicut unum ex istis
LUKE|12|28|si autem faenum quod hodie in agro est et cras in clibanum mittitur Deus sic vestit quanto magis vos pusillae fidei
LUKE|12|29|et vos nolite quaerere quid manducetis aut quid bibatis et nolite in sublime tolli
LUKE|12|30|haec enim omnia gentes mundi quaerunt Pater autem vester scit quoniam his indigetis
LUKE|12|31|verumtamen quaerite regnum Dei et haec omnia adicientur vobis
LUKE|12|32|nolite timere pusillus grex quia conplacuit Patri vestro dare vobis regnum
LUKE|12|33|vendite quae possidetis et date elemosynam facite vobis sacculos qui non veterescunt thesaurum non deficientem in caelis quo fur non adpropiat neque tinea corrumpit
LUKE|12|34|ubi enim thesaurus vester est ibi et cor vestrum erit
LUKE|12|35|sint lumbi vestri praecincti et lucernae ardentes
LUKE|12|36|et vos similes hominibus expectantibus dominum suum quando revertatur a nuptiis ut cum venerit et pulsaverit confestim aperiant ei
LUKE|12|37|beati servi illi quos cum venerit dominus invenerit vigilantes amen dico vobis quod praecinget se et faciet illos discumbere et transiens ministrabit illis
LUKE|12|38|et si venerit in secunda vigilia et si in tertia vigilia venerit et ita invenerit beati sunt servi illi
LUKE|12|39|hoc autem scitote quia si sciret pater familias qua hora fur veniret vigilaret utique et non sineret perfodiri domum suam
LUKE|12|40|et vos estote parati quia qua hora non putatis Filius hominis venit
LUKE|12|41|ait autem ei Petrus Domine ad nos dicis hanc parabolam an et ad omnes
LUKE|12|42|dixit autem Dominus quis putas est fidelis dispensator et prudens quem constituet dominus super familiam suam ut det illis in tempore tritici mensuram
LUKE|12|43|beatus ille servus quem cum venerit dominus invenerit ita facientem
LUKE|12|44|vere dico vobis quia supra omnia quae possidet constituet illum
LUKE|12|45|quod si dixerit servus ille in corde suo moram facit dominus meus venire et coeperit percutere pueros et ancillas et edere et bibere et inebriari
LUKE|12|46|veniet dominus servi illius in die qua non sperat et hora qua nescit et dividet eum partemque eius cum infidelibus ponet
LUKE|12|47|ille autem servus qui cognovit voluntatem domini sui et non praeparavit et non fecit secundum voluntatem eius vapulabit multas
LUKE|12|48|qui autem non cognovit et fecit digna plagis vapulabit paucis omni autem cui multum datum est multum quaeretur ab eo et cui commendaverunt multum plus petent ab eo
LUKE|12|49|ignem veni mittere in terram et quid volo si accendatur
LUKE|12|50|baptisma autem habeo baptizari et quomodo coartor usque dum perficiatur
LUKE|12|51|putatis quia pacem veni dare in terram non dico vobis sed separationem
LUKE|12|52|erunt enim ex hoc quinque in domo una divisi tres in duo et duo in tres
LUKE|12|53|dividentur pater in filium et filius in patrem suum mater in filiam et filia in matrem socrus in nurum suam et nurus in socrum suam
LUKE|12|54|dicebat autem et ad turbas cum videritis nubem orientem ab occasu statim dicitis nimbus venit et ita fit
LUKE|12|55|et cum austrum flantem dicitis quia aestus erit et fit
LUKE|12|56|hypocritae faciem terrae et caeli nostis probare hoc autem tempus quomodo non probatis
LUKE|12|57|quid autem et a vobis ipsis non iudicatis quod iustum est
LUKE|12|58|cum autem vadis cum adversario tuo ad principem in via da operam liberari ab illo ne forte trahat te apud iudicem et iudex tradat te exactori et exactor mittat te in carcerem
LUKE|12|59|dico tibi non exies inde donec etiam novissimum minutum reddas
LUKE|13|1|aderant autem quidam ipso in tempore nuntiantes illi de Galilaeis quorum sanguinem Pilatus miscuit cum sacrificiis eorum
LUKE|13|2|et respondens dixit illis putatis quod hii Galilaei prae omnibus Galilaeis peccatores fuerunt quia talia passi sunt
LUKE|13|3|non dico vobis sed nisi paenitentiam habueritis omnes similiter peribitis
LUKE|13|4|sicut illi decem et octo supra quos cecidit turris in Siloam et occidit eos putatis quia et ipsi debitores fuerunt praeter omnes homines habitantes in Hierusalem
LUKE|13|5|non dico vobis sed si non paenitentiam egeritis omnes similiter peribitis
LUKE|13|6|dicebat autem hanc similitudinem arborem fici habebat quidam plantatam in vinea sua et venit quaerens fructum in illa et non invenit
LUKE|13|7|dixit autem ad cultorem vineae ecce anni tres sunt ex quo venio quaerens fructum in ficulnea hac et non invenio succide ergo illam ut quid etiam terram occupat
LUKE|13|8|at ille respondens dixit illi domine dimitte illam et hoc anno usque dum fodiam circa illam et mittam stercora
LUKE|13|9|et si quidem fecerit fructum sin autem in futurum succides eam
LUKE|13|10|erat autem docens in synagoga eorum sabbatis
LUKE|13|11|et ecce mulier quae habebat spiritum infirmitatis annis decem et octo et erat inclinata nec omnino poterat sursum respicere
LUKE|13|12|quam cum videret Iesus vocavit ad se et ait illi mulier dimissa es ab infirmitate tua
LUKE|13|13|et inposuit illi manus et confestim erecta est et glorificabat Deum
LUKE|13|14|respondens autem archisynagogus indignans quia sabbato curasset Iesus dicebat turbae sex dies sunt in quibus oportet operari in his ergo venite et curamini et non in die sabbati
LUKE|13|15|respondit autem ad illum Dominus et dixit hypocritae unusquisque vestrum sabbato non solvit bovem suum aut asinum a praesepio et ducit adaquare
LUKE|13|16|hanc autem filiam Abrahae quam alligavit Satanas ecce decem et octo annis non oportuit solvi a vinculo isto die sabbati
LUKE|13|17|et cum haec diceret erubescebant omnes adversarii eius et omnis populus gaudebat in universis quae gloriose fiebant ab eo
LUKE|13|18|dicebat ergo cui simile est regnum Dei et cui simile esse existimabo illud
LUKE|13|19|simile est grano sinapis quod acceptum homo misit in hortum suum et crevit et factum est in arborem magnam et volucres caeli requieverunt in ramis eius
LUKE|13|20|et iterum dixit cui simile aestimabo regnum Dei
LUKE|13|21|simile est fermento quod acceptum mulier abscondit in farinae sata tria donec fermentaretur totum
LUKE|13|22|et ibat per civitates et castella docens et iter faciens in Hierusalem
LUKE|13|23|ait autem illi quidam Domine si pauci sunt qui salvantur ipse autem dixit ad illos
LUKE|13|24|contendite intrare per angustam portam quia multi dico vobis quaerunt intrare et non poterunt
LUKE|13|25|cum autem intraverit pater familias et cluserit ostium et incipietis foris stare et pulsare ostium dicentes Domine aperi nobis et respondens dicet vobis nescio vos unde sitis
LUKE|13|26|tunc incipietis dicere manducavimus coram te et bibimus et in plateis nostris docuisti
LUKE|13|27|et dicet vobis nescio vos unde sitis discedite a me omnes operarii iniquitatis
LUKE|13|28|ibi erit fletus et stridor dentium cum videritis Abraham et Isaac et Iacob et omnes prophetas in regno Dei vos autem expelli foras
LUKE|13|29|et venient ab oriente et occidente et aquilone et austro et accumbent in regno Dei
LUKE|13|30|et ecce sunt novissimi qui erunt primi et sunt primi qui erunt novissimi
LUKE|13|31|in ipsa die accesserunt quidam Pharisaeorum dicentes illi exi et vade hinc quia Herodes vult te occidere
LUKE|13|32|et ait illis ite dicite vulpi illi ecce eicio daemonia et sanitates perficio hodie et cras et tertia consummor
LUKE|13|33|verumtamen oportet me hodie et cras et sequenti ambulare quia non capit prophetam perire extra Hierusalem
LUKE|13|34|Hierusalem Hierusalem quae occidis prophetas et lapidas eos qui mittuntur ad te quotiens volui congregare filios tuos quemadmodum avis nidum suum sub pinnis et noluisti
LUKE|13|35|ecce relinquitur vobis domus vestra dico autem vobis quia non videbitis me donec veniat cum dicetis benedictus qui venit in nomine Domini
LUKE|14|1|et factum est cum intraret in domum cuiusdam principis Pharisaeorum sabbato manducare panem et ipsi observabant eum
LUKE|14|2|et ecce homo quidam hydropicus erat ante illum
LUKE|14|3|et respondens Iesus dixit ad legis peritos et Pharisaeos dicens si licet sabbato curare
LUKE|14|4|at illi tacuerunt ipse vero adprehensum sanavit eum ac dimisit
LUKE|14|5|et respondens ad illos dixit cuius vestrum asinus aut bos in puteum cadet et non continuo extrahet illum die sabbati
LUKE|14|6|et non poterant ad haec respondere illi
LUKE|14|7|dicebat autem et ad invitatos parabolam intendens quomodo primos accubitus eligerent dicens ad illos
LUKE|14|8|cum invitatus fueris ad nuptias non discumbas in primo loco ne forte honoratior te sit invitatus ab eo
LUKE|14|9|et veniens is qui te et illum vocavit dicat tibi da huic locum et tunc incipias cum rubore novissimum locum tenere
LUKE|14|10|sed cum vocatus fueris vade recumbe in novissimo loco ut cum venerit qui te invitavit dicat tibi amice ascende superius tunc erit tibi gloria coram simul discumbentibus
LUKE|14|11|quia omnis qui se exaltat humiliabitur et qui se humiliat exaltabitur
LUKE|14|12|dicebat autem et ei qui se invitaverat cum facis prandium aut cenam noli vocare amicos tuos neque fratres tuos neque cognatos neque vicinos divites ne forte et ipsi te reinvitent et fiat tibi retributio
LUKE|14|13|sed cum facis convivium voca pauperes debiles claudos caecos
LUKE|14|14|et beatus eris quia non habent retribuere tibi retribuetur enim tibi in resurrectione iustorum
LUKE|14|15|haec cum audisset quidam de simul discumbentibus dixit illi beatus qui manducabit panem in regno Dei
LUKE|14|16|at ipse dixit ei homo quidam fecit cenam magnam et vocavit multos
LUKE|14|17|et misit servum suum hora cenae dicere invitatis ut venirent quia iam parata sunt omnia
LUKE|14|18|et coeperunt simul omnes excusare primus dixit ei villam emi et necesse habeo exire et videre illam rogo te habe me excusatum
LUKE|14|19|et alter dixit iuga boum emi quinque et eo probare illa rogo te habe me excusatum
LUKE|14|20|et alius dixit uxorem duxi et ideo non possum venire
LUKE|14|21|et reversus servus nuntiavit haec domino suo tunc iratus pater familias dixit servo suo exi cito in plateas et vicos civitatis et pauperes ac debiles et caecos et claudos introduc huc
LUKE|14|22|et ait servus domine factum est ut imperasti et adhuc locus est
LUKE|14|23|et ait dominus servo exi in vias et sepes et conpelle intrare ut impleatur domus mea
LUKE|14|24|dico autem vobis quod nemo virorum illorum qui vocati sunt gustabit cenam meam
LUKE|14|25|ibant autem turbae multae cum eo et conversus dixit ad illos
LUKE|14|26|si quis venit ad me et non odit patrem suum et matrem et uxorem et filios et fratres et sorores adhuc autem et animam suam non potest esse meus discipulus
LUKE|14|27|et qui non baiulat crucem suam et venit post me non potest esse meus discipulus
LUKE|14|28|quis enim ex vobis volens turrem aedificare non prius sedens conputat sumptus qui necessarii sunt si habet ad perficiendum
LUKE|14|29|ne posteaquam posuerit fundamentum et non potuerit perficere omnes qui vident incipiant inludere ei
LUKE|14|30|dicentes quia hic homo coepit aedificare et non potuit consummare
LUKE|14|31|aut qui rex iturus committere bellum adversus alium regem non sedens prius cogitat si possit cum decem milibus occurrere ei qui cum viginti milibus venit ad se
LUKE|14|32|alioquin adhuc illo longe agente legationem mittens rogat ea quae pacis sunt
LUKE|14|33|sic ergo omnis ex vobis qui non renuntiat omnibus quae possidet non potest meus esse discipulus
LUKE|14|34|bonum est sal si autem sal quoque evanuerit in quo condietur
LUKE|14|35|neque in terram neque in sterquilinium utile est sed foras mittetur qui habet aures audiendi audiat
LUKE|15|1|erant autem adpropinquantes ei publicani et peccatores ut audirent illum
LUKE|15|2|et murmurabant Pharisaei et scribae dicentes quia hic peccatores recipit et manducat cum illis
LUKE|15|3|et ait ad illos parabolam istam dicens
LUKE|15|4|quis ex vobis homo qui habet centum oves et si perdiderit unam ex illis nonne dimittit nonaginta novem in deserto et vadit ad illam quae perierat donec inveniat illam
LUKE|15|5|et cum invenerit eam inponit in umeros suos gaudens
LUKE|15|6|et veniens domum convocat amicos et vicinos dicens illis congratulamini mihi quia inveni ovem meam quae perierat
LUKE|15|7|dico vobis quod ita gaudium erit in caelo super uno peccatore paenitentiam habente quam super nonaginta novem iustis qui non indigent paenitentia
LUKE|15|8|aut quae mulier habens dragmas decem si perdiderit dragmam unam nonne accendit lucernam et everrit domum et quaerit diligenter donec inveniat
LUKE|15|9|et cum invenerit convocat amicas et vicinas dicens congratulamini mihi quia inveni dragmam quam perdideram
LUKE|15|10|ita dico vobis gaudium erit coram angelis Dei super uno peccatore paenitentiam agente
LUKE|15|11|ait autem homo quidam habuit duos filios
LUKE|15|12|et dixit adulescentior ex illis patri pater da mihi portionem substantiae quae me contingit et divisit illis substantiam
LUKE|15|13|et non post multos dies congregatis omnibus adulescentior filius peregre profectus est in regionem longinquam et ibi dissipavit substantiam suam vivendo luxuriose
LUKE|15|14|et postquam omnia consummasset facta est fames valida in regione illa et ipse coepit egere
LUKE|15|15|et abiit et adhesit uni civium regionis illius et misit illum in villam suam ut pasceret porcos
LUKE|15|16|et cupiebat implere ventrem suum de siliquis quas porci manducabant et nemo illi dabat
LUKE|15|17|in se autem reversus dixit quanti mercennarii patris mei abundant panibus ego autem hic fame pereo
LUKE|15|18|surgam et ibo ad patrem meum et dicam illi pater peccavi in caelum et coram te
LUKE|15|19|et iam non sum dignus vocari filius tuus fac me sicut unum de mercennariis tuis
LUKE|15|20|et surgens venit ad patrem suum cum autem adhuc longe esset vidit illum pater ipsius et misericordia motus est et adcurrens cecidit supra collum eius et osculatus est illum
LUKE|15|21|dixitque ei filius pater peccavi in caelum et coram te iam non sum dignus vocari filius tuus
LUKE|15|22|dixit autem pater ad servos suos cito proferte stolam primam et induite illum et date anulum in manum eius et calciamenta in pedes
LUKE|15|23|et adducite vitulum saginatum et occidite et manducemus et epulemur
LUKE|15|24|quia hic filius meus mortuus erat et revixit perierat et inventus est et coeperunt epulari
LUKE|15|25|erat autem filius eius senior in agro et cum veniret et adpropinquaret domui audivit symphoniam et chorum
LUKE|15|26|et vocavit unum de servis et interrogavit quae haec essent
LUKE|15|27|isque dixit illi frater tuus venit et occidit pater tuus vitulum saginatum quia salvum illum recepit
LUKE|15|28|indignatus est autem et nolebat introire pater ergo illius egressus coepit rogare illum
LUKE|15|29|at ille respondens dixit patri suo ecce tot annis servio tibi et numquam mandatum tuum praeterii et numquam dedisti mihi hedum ut cum amicis meis epularer
LUKE|15|30|sed postquam filius tuus hic qui devoravit substantiam suam cum meretricibus venit occidisti illi vitulum saginatum
LUKE|15|31|at ipse dixit illi fili tu semper mecum es et omnia mea tua sunt
LUKE|15|32|epulari autem et gaudere oportebat quia frater tuus hic mortuus erat et revixit perierat et inventus est
LUKE|16|1|dicebat autem et ad discipulos suos homo quidam erat dives qui habebat vilicum et hic diffamatus est apud illum quasi dissipasset bona ipsius
LUKE|16|2|et vocavit illum et ait illi quid hoc audio de te redde rationem vilicationis tuae iam enim non poteris vilicare
LUKE|16|3|ait autem vilicus intra se quid faciam quia dominus meus aufert a me vilicationem fodere non valeo mendicare erubesco
LUKE|16|4|scio quid faciam ut cum amotus fuero a vilicatione recipiant me in domos suas
LUKE|16|5|convocatis itaque singulis debitoribus domini sui dicebat primo quantum debes domino meo
LUKE|16|6|at ille dixit centum cados olei dixitque illi accipe cautionem tuam et sede cito scribe quinquaginta
LUKE|16|7|deinde alio dixit tu vero quantum debes qui ait centum choros tritici ait illi accipe litteras tuas et scribe octoginta
LUKE|16|8|et laudavit dominus vilicum iniquitatis quia prudenter fecisset quia filii huius saeculi prudentiores filiis lucis in generatione sua sunt
LUKE|16|9|et ego vobis dico facite vobis amicos de mamona iniquitatis ut cum defeceritis recipiant vos in aeterna tabernacula
LUKE|16|10|qui fidelis est in minimo et in maiori fidelis est et qui in modico iniquus est et in maiori iniquus est
LUKE|16|11|si ergo in iniquo mamona fideles non fuistis quod verum est quis credet vobis
LUKE|16|12|et si in alieno fideles non fuistis quod vestrum est quis dabit vobis
LUKE|16|13|nemo servus potest duobus dominis servire aut enim unum odiet et alterum diliget aut uni adherebit et alterum contemnet non potestis Deo servire et mamonae
LUKE|16|14|audiebant autem omnia haec Pharisaei qui erant avari et deridebant illum
LUKE|16|15|et ait illis vos estis qui iustificatis vos coram hominibus Deus autem novit corda vestra quia quod hominibus altum est abominatio est ante Deum
LUKE|16|16|lex et prophetae usque ad Iohannem ex eo regnum Dei evangelizatur et omnis in illud vim facit
LUKE|16|17|facilius est autem caelum et terram praeterire quam de lege unum apicem cadere
LUKE|16|18|omnis qui dimittit uxorem suam et ducit alteram moechatur et qui dimissam a viro ducit moechatur
LUKE|16|19|homo quidam erat dives et induebatur purpura et bysso et epulabatur cotidie splendide
LUKE|16|20|et erat quidam mendicus nomine Lazarus qui iacebat ad ianuam eius ulceribus plenus
LUKE|16|21|cupiens saturari de micis quae cadebant de mensa divitis sed et canes veniebant et lingebant ulcera eius
LUKE|16|22|factum est autem ut moreretur mendicus et portaretur ab angelis in sinum Abrahae mortuus est autem et dives et sepultus est in inferno
LUKE|16|23|elevans oculos suos cum esset in tormentis videbat Abraham a longe et Lazarum in sinu eius
LUKE|16|24|et ipse clamans dixit pater Abraham miserere mei et mitte Lazarum ut intinguat extremum digiti sui in aqua ut refrigeret linguam meam quia crucior in hac flamma
LUKE|16|25|et dixit illi Abraham fili recordare quia recepisti bona in vita tua et Lazarus similiter mala nunc autem hic consolatur tu vero cruciaris
LUKE|16|26|et in his omnibus inter nos et vos chasma magnum firmatum est ut hii qui volunt hinc transire ad vos non possint neque inde huc transmeare
LUKE|16|27|et ait rogo ergo te pater ut mittas eum in domum patris mei
LUKE|16|28|habeo enim quinque fratres ut testetur illis ne et ipsi veniant in locum hunc tormentorum
LUKE|16|29|et ait illi Abraham habent Mosen et prophetas audiant illos
LUKE|16|30|at ille dixit non pater Abraham sed si quis ex mortuis ierit ad eos paenitentiam agent
LUKE|16|31|ait autem illi si Mosen et prophetas non audiunt neque si quis ex mortuis resurrexerit credent
LUKE|17|1|et ad discipulos suos ait inpossibile est ut non veniant scandala vae autem illi per quem veniunt
LUKE|17|2|utilius est illi si lapis molaris inponatur circa collum eius et proiciatur in mare quam ut scandalizet unum de pusillis istis
LUKE|17|3|adtendite vobis si peccaverit frater tuus increpa illum et si paenitentiam egerit dimitte illi
LUKE|17|4|et si septies in die peccaverit in te et septies in die conversus fuerit ad te dicens paenitet me dimitte illi
LUKE|17|5|et dixerunt apostoli Domino adauge nobis fidem
LUKE|17|6|dixit autem Dominus si haberetis fidem sicut granum sinapis diceretis huic arbori moro eradicare et transplantare in mare et oboediret vobis
LUKE|17|7|quis autem vestrum habens servum arantem aut pascentem qui regresso de agro dicet illi statim transi recumbe
LUKE|17|8|et non dicet ei para quod cenem et praecinge te et ministra mihi donec manducem et bibam et post haec tu manducabis et bibes
LUKE|17|9|numquid gratiam habet servo illi quia fecit quae sibi imperaverat non puto
LUKE|17|10|sic et vos cum feceritis omnia quae praecepta sunt vobis dicite servi inutiles sumus quod debuimus facere fecimus
LUKE|17|11|et factum est dum iret in Hierusalem transiebat per mediam Samariam et Galilaeam
LUKE|17|12|et cum ingrederetur quoddam castellum occurrerunt ei decem viri leprosi qui steterunt a longe
LUKE|17|13|et levaverunt vocem dicentes Iesu praeceptor miserere nostri
LUKE|17|14|quos ut vidit dixit ite ostendite vos sacerdotibus et factum est dum irent mundati sunt
LUKE|17|15|unus autem ex illis ut vidit quia mundatus est regressus est cum magna voce magnificans Deum
LUKE|17|16|et cecidit in faciem ante pedes eius gratias agens et hic erat Samaritanus
LUKE|17|17|respondens autem Iesus dixit nonne decem mundati sunt et novem ubi sunt
LUKE|17|18|non est inventus qui rediret et daret gloriam Deo nisi hic alienigena
LUKE|17|19|et ait illi surge vade quia fides tua te salvum fecit
LUKE|17|20|interrogatus autem a Pharisaeis quando venit regnum Dei respondit eis et dixit non venit regnum Dei cum observatione
LUKE|17|21|neque dicent ecce hic aut ecce illic ecce enim regnum Dei intra vos est
LUKE|17|22|et ait ad discipulos venient dies quando desideretis videre unum diem Filii hominis et non videbitis
LUKE|17|23|et dicent vobis ecce hic ecce illic nolite ire neque sectemini
LUKE|17|24|nam sicut fulgur coruscans de sub caelo in ea quae sub caelo sunt fulget ita erit Filius hominis in die sua
LUKE|17|25|primum autem oportet illum multa pati et reprobari a generatione hac
LUKE|17|26|et sicut factum est in diebus Noe ita erit et in diebus Filii hominis
LUKE|17|27|edebant et bibebant uxores ducebant et dabantur ad nuptias usque in diem qua intravit Noe in arcam et venit diluvium et perdidit omnes
LUKE|17|28|similiter sicut factum est in diebus Loth edebant et bibebant emebant et vendebant plantabant aedificabant
LUKE|17|29|qua die autem exiit Loth a Sodomis pluit ignem et sulphur de caelo et omnes perdidit
LUKE|17|30|secundum haec erit qua die Filius hominis revelabitur
LUKE|17|31|in illa hora qui fuerit in tecto et vasa eius in domo ne descendat tollere illa et qui in agro similiter non redeat retro
LUKE|17|32|memores estote uxoris Loth
LUKE|17|33|quicumque quaesierit animam suam salvare perdet illam et qui perdiderit illam vivificabit eam
LUKE|17|34|dico vobis illa nocte erunt duo in lecto uno unus adsumetur et alter relinquetur
LUKE|17|35|duae erunt molentes in unum una adsumetur et altera relinquetur duo in agro unus adsumetur et alter relinquetur
LUKE|17|36|respondentes dicunt illi ubi Domine
LUKE|17|37|qui dixit eis ubicumque fuerit corpus illuc congregabuntur aquilae
LUKE|18|1|dicebat autem et parabolam ad illos quoniam oportet semper orare et non deficere
LUKE|18|2|dicens iudex quidam erat in quadam civitate qui Deum non timebat et hominem non verebatur
LUKE|18|3|vidua autem quaedam erat in civitate illa et veniebat ad eum dicens vindica me de adversario meo
LUKE|18|4|et nolebat per multum tempus post haec autem dixit intra se et si Deum non timeo nec hominem revereor
LUKE|18|5|tamen quia molesta est mihi haec vidua vindicabo illam ne in novissimo veniens suggillet me
LUKE|18|6|ait autem Dominus audite quid iudex iniquitatis dicit
LUKE|18|7|Deus autem non faciet vindictam electorum suorum clamantium ad se die ac nocte et patientiam habebit in illis
LUKE|18|8|dico vobis quia cito faciet vindictam illorum verumtamen Filius hominis veniens putas inveniet fidem in terra
LUKE|18|9|dixit autem et ad quosdam qui in se confidebant tamquam iusti et aspernabantur ceteros parabolam istam
LUKE|18|10|duo homines ascenderunt in templum ut orarent unus Pharisaeus et alter publicanus
LUKE|18|11|Pharisaeus stans haec apud se orabat Deus gratias ago tibi quia non sum sicut ceteri hominum raptores iniusti adulteri vel ut etiam hic publicanus
LUKE|18|12|ieiuno bis in sabbato decimas do omnium quae possideo
LUKE|18|13|et publicanus a longe stans nolebat nec oculos ad caelum levare sed percutiebat pectus suum dicens Deus propitius esto mihi peccatori
LUKE|18|14|dico vobis descendit hic iustificatus in domum suam ab illo quia omnis qui se exaltat humiliabitur et qui se humiliat exaltabitur
LUKE|18|15|adferebant autem ad illum et infantes ut eos tangeret quod cum viderent discipuli increpabant illos
LUKE|18|16|Iesus autem convocans illos dixit sinite pueros venire ad me et nolite eos vetare talium est enim regnum Dei
LUKE|18|17|amen dico vobis quicumque non acceperit regnum Dei sicut puer non intrabit in illud
LUKE|18|18|et interrogavit eum quidam princeps dicens magister bone quid faciens vitam aeternam possidebo
LUKE|18|19|dixit autem ei Iesus quid me dicis bonum nemo bonus nisi solus Deus
LUKE|18|20|mandata nosti non occides non moechaberis non furtum facies non falsum testimonium dices honora patrem tuum et matrem
LUKE|18|21|qui ait haec omnia custodivi a iuventute mea
LUKE|18|22|quo audito Iesus ait ei adhuc unum tibi deest omnia quaecumque habes vende et da pauperibus et habebis thesaurum in caelo et veni sequere me
LUKE|18|23|his ille auditis contristatus est quia dives erat valde
LUKE|18|24|videns autem illum Iesus tristem factum dixit quam difficile qui pecunias habent in regnum Dei intrabunt
LUKE|18|25|facilius est enim camelum per foramen acus transire quam divitem intrare in regnum Dei
LUKE|18|26|et dixerunt qui audiebant et quis potest salvus fieri
LUKE|18|27|ait illis quae inpossibilia sunt apud homines possibilia sunt apud Deum
LUKE|18|28|ait autem Petrus ecce nos dimisimus omnia et secuti sumus te
LUKE|18|29|qui dixit eis amen dico vobis nemo est qui reliquit domum aut parentes aut fratres aut uxorem aut filios propter regnum Dei
LUKE|18|30|et non recipiat multo plura in hoc tempore et in saeculo venturo vitam aeternam
LUKE|18|31|adsumpsit autem Iesus duodecim et ait illis ecce ascendimus Hierosolyma et consummabuntur omnia quae scripta sunt per prophetas de Filio hominis
LUKE|18|32|tradetur enim gentibus et inludetur et flagellabitur et conspuetur
LUKE|18|33|et postquam flagellaverint occident eum et die tertia resurget
LUKE|18|34|et ipsi nihil horum intellexerunt et erat verbum istud absconditum ab eis et non intellegebant quae dicebantur
LUKE|18|35|factum est autem cum adpropinquaret Hiericho caecus quidam sedebat secus viam mendicans
LUKE|18|36|et cum audiret turbam praetereuntem interrogabat quid hoc esset
LUKE|18|37|dixerunt autem ei quod Iesus Nazarenus transiret
LUKE|18|38|et clamavit dicens Iesu Fili David miserere mei
LUKE|18|39|et qui praeibant increpabant eum ut taceret ipse vero multo magis clamabat Fili David miserere mei
LUKE|18|40|stans autem Iesus iussit illum adduci ad se et cum adpropinquasset interrogavit illum
LUKE|18|41|dicens quid tibi vis faciam at ille dixit Domine ut videam
LUKE|18|42|et Iesus dixit illi respice fides tua te salvum fecit
LUKE|18|43|et confestim vidit et sequebatur illum magnificans Deum et omnis plebs ut vidit dedit laudem Deo
LUKE|19|1|et ingressus perambulabat Hiericho
LUKE|19|2|et ecce vir nomine Zaccheus et hic erat princeps publicanorum et ipse dives
LUKE|19|3|et quaerebat videre Iesum quis esset et non poterat prae turba quia statura pusillus erat
LUKE|19|4|et praecurrens ascendit in arborem sycomorum ut videret illum quia inde erat transiturus
LUKE|19|5|et cum venisset ad locum suspiciens Iesus vidit illum et dixit ad eum Zacchee festinans descende quia hodie in domo tua oportet me manere
LUKE|19|6|et festinans descendit et excepit illum gaudens
LUKE|19|7|et cum viderent omnes murmurabant dicentes quod ad hominem peccatorem devertisset
LUKE|19|8|stans autem Zaccheus dixit ad Dominum ecce dimidium bonorum meorum Domine do pauperibus et si quid aliquem defraudavi reddo quadruplum
LUKE|19|9|ait Iesus ad eum quia hodie salus domui huic facta est eo quod et ipse filius sit Abrahae
LUKE|19|10|venit enim Filius hominis quaerere et salvum facere quod perierat
LUKE|19|11|haec illis audientibus adiciens dixit parabolam eo quod esset prope Hierusalem et quia existimarent quod confestim regnum Dei manifestaretur
LUKE|19|12|dixit ergo homo quidam nobilis abiit in regionem longinquam accipere sibi regnum et reverti
LUKE|19|13|vocatis autem decem servis suis dedit illis decem mnas et ait ad illos negotiamini dum venio
LUKE|19|14|cives autem eius oderant illum et miserunt legationem post illum dicentes nolumus hunc regnare super nos
LUKE|19|15|et factum est ut rediret accepto regno et iussit vocari servos quibus dedit pecuniam ut sciret quantum quisque negotiatus esset
LUKE|19|16|venit autem primus dicens domine mna tua decem mnas adquisivit
LUKE|19|17|et ait illi euge bone serve quia in modico fidelis fuisti eris potestatem habens supra decem civitates
LUKE|19|18|et alter venit dicens domine mna tua fecit quinque mnas
LUKE|19|19|et huic ait et tu esto supra quinque civitates
LUKE|19|20|et alter venit dicens domine ecce mna tua quam habui repositam in sudario
LUKE|19|21|timui enim te quia homo austeris es tollis quod non posuisti et metis quod non seminasti
LUKE|19|22|dicit ei de ore tuo te iudico serve nequam sciebas quod ego austeris homo sum tollens quod non posui et metens quod non seminavi
LUKE|19|23|et quare non dedisti pecuniam meam ad mensam et ego veniens cum usuris utique exegissem illud
LUKE|19|24|et adstantibus dixit auferte ab illo mnam et date illi qui decem mnas habet
LUKE|19|25|et dixerunt ei domine habet decem mnas
LUKE|19|26|dico autem vobis quia omni habenti dabitur ab eo autem qui non habet et quod habet auferetur ab eo
LUKE|19|27|verumtamen inimicos meos illos qui noluerunt me regnare super se adducite huc et interficite ante me
LUKE|19|28|et his dictis praecedebat ascendens in Hierosolyma
LUKE|19|29|et factum est cum adpropinquasset ad Bethfage et Bethania ad montem qui vocatur Oliveti misit duos discipulos suos
LUKE|19|30|dicens ite in castellum quod contra est in quod introeuntes invenietis pullum asinae alligatum cui nemo umquam hominum sedit solvite illum et adducite
LUKE|19|31|et si quis vos interrogaverit quare solvitis sic dicetis ei quia Dominus operam eius desiderat
LUKE|19|32|abierunt autem qui missi erant et invenerunt sicut dixit illis stantem pullum
LUKE|19|33|solventibus autem illis pullum dixerunt domini eius ad illos quid solvitis pullum
LUKE|19|34|at illi dixerunt quia Dominus eum necessarium habet
LUKE|19|35|et duxerunt illum ad Iesum et iactantes vestimenta sua supra pullum inposuerunt Iesum
LUKE|19|36|eunte autem illo substernebant vestimenta sua in via
LUKE|19|37|et cum adpropinquaret iam ad descensum montis Oliveti coeperunt omnes turbae discentium gaudentes laudare Deum voce magna super omnibus quas viderant virtutibus
LUKE|19|38|dicentes benedictus qui venit rex in nomine Domini pax in caelo et gloria in excelsis
LUKE|19|39|et quidam Pharisaeorum de turbis dixerunt ad illum magister increpa discipulos tuos
LUKE|19|40|quibus ipse ait dico vobis quia si hii tacuerint lapides clamabunt
LUKE|19|41|et ut adpropinquavit videns civitatem flevit super illam dicens
LUKE|19|42|quia si cognovisses et tu et quidem in hac die tua quae ad pacem tibi nunc autem abscondita sunt ab oculis tuis
LUKE|19|43|quia venient dies in te et circumdabunt te inimici tui vallo et circumdabunt te et coangustabunt te undique
LUKE|19|44|ad terram prosternent te et filios qui in te sunt et non relinquent in te lapidem super lapidem eo quod non cognoveris tempus visitationis tuae
LUKE|19|45|et ingressus in templum coepit eicere vendentes in illo et ementes
LUKE|19|46|dicens illis scriptum est quia domus mea domus orationis est vos autem fecistis illam speluncam latronum
LUKE|19|47|et erat docens cotidie in templo principes autem sacerdotum et scribae et principes plebis quaerebant illum perdere
LUKE|19|48|et non inveniebant quid facerent illi omnis enim populus suspensus erat audiens illum
LUKE|20|1|et factum est in una dierum docente illo populum in templo et evangelizante convenerunt principes sacerdotum et scribae cum senioribus
LUKE|20|2|et aiunt dicentes ad illum dic nobis in qua potestate haec facis aut quis est qui dedit tibi hanc potestatem
LUKE|20|3|respondens autem dixit ad illos interrogabo vos et ego verbum respondete mihi
LUKE|20|4|baptismum Iohannis de caelo erat an ex hominibus
LUKE|20|5|at illi cogitabant inter se dicentes quia si dixerimus de caelo dicet quare ergo non credidistis illi
LUKE|20|6|si autem dixerimus ex hominibus plebs universa lapidabit nos certi sunt enim Iohannem prophetam esse
LUKE|20|7|et responderunt se nescire unde esset
LUKE|20|8|et Iesus ait illis neque ego dico vobis in qua potestate haec facio
LUKE|20|9|coepit autem dicere ad plebem parabolam hanc homo plantavit vineam et locavit eam colonis et ipse peregre fuit multis temporibus
LUKE|20|10|et in tempore misit ad cultores servum ut de fructu vineae darent illi qui caesum dimiserunt eum inanem
LUKE|20|11|et addidit alterum servum mittere illi autem hunc quoque caedentes et adficientes contumelia dimiserunt inanem
LUKE|20|12|et addidit tertium mittere qui et illum vulnerantes eiecerunt
LUKE|20|13|dixit autem dominus vineae quid faciam mittam filium meum dilectum forsitan cum hunc viderint verebuntur
LUKE|20|14|quem cum vidissent coloni cogitaverunt inter se dicentes hic est heres occidamus illum ut nostra fiat hereditas
LUKE|20|15|et eiectum illum extra vineam occiderunt quid ergo faciet illis dominus vineae
LUKE|20|16|veniet et perdet colonos istos et dabit vineam aliis quo audito dixerunt illi absit
LUKE|20|17|ille autem aspiciens eos ait quid est ergo hoc quod scriptum est lapidem quem reprobaverunt aedificantes hic factus est in caput anguli
LUKE|20|18|omnis qui ceciderit supra illum lapidem conquassabitur supra quem autem ceciderit comminuet illum
LUKE|20|19|et quaerebant principes sacerdotum et scribae mittere in illum manus illa hora et timuerunt populum cognoverunt enim quod ad ipsos dixerit similitudinem istam
LUKE|20|20|et observantes miserunt insidiatores qui se iustos simularent ut caperent eum in sermone et traderent illum principatui et potestati praesidis
LUKE|20|21|et interrogaverunt illum dicentes magister scimus quia recte dicis et doces et non accipis personam sed in veritate viam Dei doces
LUKE|20|22|licet nobis dare tributum Caesari an non
LUKE|20|23|considerans autem dolum illorum dixit ad eos quid me temptatis
LUKE|20|24|ostendite mihi denarium cuius habet imaginem et inscriptionem respondentes dixerunt Caesaris
LUKE|20|25|et ait illis reddite ergo quae Caesaris sunt Caesari et quae Dei sunt Deo
LUKE|20|26|et non potuerunt verbum eius reprehendere coram plebe et mirati in responso eius tacuerunt
LUKE|20|27|accesserunt autem quidam Sadducaeorum qui negant esse resurrectionem et interrogaverunt eum
LUKE|20|28|dicentes magister Moses scripsit nobis si frater alicuius mortuus fuerit habens uxorem et hic sine filiis fuerit ut accipiat eam frater eius uxorem et suscitet semen fratri suo
LUKE|20|29|septem ergo fratres erant et primus accepit uxorem et mortuus est sine filiis
LUKE|20|30|et sequens accepit illam et ipse mortuus est sine filio
LUKE|20|31|et tertius accepit illam similiter et omnes septem et non reliquerunt semen et mortui sunt
LUKE|20|32|novissima omnium mortua est et mulier
LUKE|20|33|in resurrectione ergo cuius eorum erit uxor siquidem septem habuerunt eam uxorem
LUKE|20|34|et ait illis Iesus filii saeculi huius nubunt et traduntur ad nuptias
LUKE|20|35|illi autem qui digni habebuntur saeculo illo et resurrectione ex mortuis neque nubunt neque ducunt uxores
LUKE|20|36|neque enim ultra mori poterunt aequales enim angelis sunt et filii sunt Dei cum sint filii resurrectionis
LUKE|20|37|quia vero resurgant mortui et Moses ostendit secus rubum sicut dicit Dominum Deum Abraham et Deum Isaac et Deum Iacob
LUKE|20|38|Deus autem non est mortuorum sed vivorum omnes enim vivunt ei
LUKE|20|39|respondentes autem quidam scribarum dixerunt magister bene dixisti
LUKE|20|40|et amplius non audebant eum quicquam interrogare
LUKE|20|41|dixit autem ad illos quomodo dicunt Christum Filium David esse
LUKE|20|42|et ipse David dicit in libro Psalmorum dixit Dominus Domino meo sede a dextris meis
LUKE|20|43|donec ponam inimicos tuos scabillum pedum tuorum
LUKE|20|44|David ergo Dominum illum vocat et quomodo filius eius est
LUKE|20|45|audiente autem omni populo dixit discipulis suis
LUKE|20|46|adtendite a scribis qui volunt ambulare in stolis et amant salutationes in foro et primas cathedras in synagogis et primos discubitus in conviviis
LUKE|20|47|qui devorant domos viduarum simulantes longam orationem hii accipient damnationem maiorem
LUKE|21|1|respiciens autem vidit eos qui mittebant munera sua in gazofilacium divites
LUKE|21|2|vidit autem et quandam viduam pauperculam mittentem aera minuta duo
LUKE|21|3|et dixit vere dico vobis quia vidua haec pauper plus quam omnes misit
LUKE|21|4|nam omnes hii ex abundanti sibi miserunt in munera Dei haec autem ex eo quod deest illi omnem victum suum quem habuit misit
LUKE|21|5|et quibusdam dicentibus de templo quod lapidibus bonis et donis ornatum esset dixit
LUKE|21|6|haec quae videtis venient dies in quibus non relinquetur lapis super lapidem qui non destruatur
LUKE|21|7|interrogaverunt autem illum dicentes praeceptor quando haec erunt et quod signum cum fieri incipient
LUKE|21|8|qui dixit videte ne seducamini multi enim venient in nomine meo dicentes quia ego sum et tempus adpropinquavit nolite ergo ire post illos
LUKE|21|9|cum autem audieritis proelia et seditiones nolite terreri oportet primum haec fieri sed non statim finis
LUKE|21|10|tunc dicebat illis surget gens contra gentem et regnum adversus regnum
LUKE|21|11|terraemotus magni erunt per loca et pestilentiae et fames terroresque de caelo et signa magna erunt
LUKE|21|12|sed ante haec omnia inicient vobis manus suas et persequentur tradentes in synagogas et custodias trahentes ad reges et praesides propter nomen meum
LUKE|21|13|continget autem vobis in testimonium
LUKE|21|14|ponite ergo in cordibus vestris non praemeditari quemadmodum respondeatis
LUKE|21|15|ego enim dabo vobis os et sapientiam cui non poterunt resistere et contradicere omnes adversarii vestri
LUKE|21|16|trademini autem a parentibus et fratribus et cognatis et amicis et morte adficient ex vobis
LUKE|21|17|et eritis odio omnibus propter nomen meum
LUKE|21|18|et capillus de capite vestro non peribit
LUKE|21|19|in patientia vestra possidebitis animas vestras
LUKE|21|20|cum autem videritis circumdari ab exercitu Hierusalem tunc scitote quia adpropinquavit desolatio eius
LUKE|21|21|tunc qui in Iudaea sunt fugiant in montes et qui in medio eius discedant et qui in regionibus non intrent in eam
LUKE|21|22|quia dies ultionis hii sunt ut impleantur omnia quae scripta sunt
LUKE|21|23|vae autem praegnatibus et nutrientibus in illis diebus erit enim pressura magna supra terram et ira populo huic
LUKE|21|24|et cadent in ore gladii et captivi ducentur in omnes gentes et Hierusalem calcabitur a gentibus donec impleantur tempora nationum
LUKE|21|25|et erunt signa in sole et luna et stellis et in terris pressura gentium prae confusione sonitus maris et fluctuum
LUKE|21|26|arescentibus hominibus prae timore et expectatione quae supervenient universo orbi nam virtutes caelorum movebuntur
LUKE|21|27|et tunc videbunt Filium hominis venientem in nube cum potestate magna et maiestate
LUKE|21|28|his autem fieri incipientibus respicite et levate capita vestra quoniam adpropinquat redemptio vestra
LUKE|21|29|et dixit illis similitudinem videte ficulneam et omnes arbores
LUKE|21|30|cum producunt iam ex se fructum scitis quoniam prope est aestas
LUKE|21|31|ita et vos cum videritis haec fieri scitote quoniam prope est regnum Dei
LUKE|21|32|amen dico vobis quia non praeteribit generatio haec donec omnia fiant
LUKE|21|33|caelum et terra transibunt verba autem mea non transient
LUKE|21|34|adtendite autem vobis ne forte graventur corda vestra in crapula et ebrietate et curis huius vitae et superveniat in vos repentina dies illa
LUKE|21|35|tamquam laqueus enim superveniet in omnes qui sedent super faciem omnis terrae
LUKE|21|36|vigilate itaque omni tempore orantes ut digni habeamini fugere ista omnia quae futura sunt et stare ante Filium hominis
LUKE|21|37|erat autem diebus docens in templo noctibus vero exiens morabatur in monte qui vocatur Oliveti
LUKE|21|38|et omnis populus manicabat ad eum in templo audire eum
LUKE|22|1|adpropinquabat autem dies festus azymorum qui dicitur pascha
LUKE|22|2|et quaerebant principes sacerdotum et scribae quomodo eum interficerent timebant vero plebem
LUKE|22|3|intravit autem Satanas in Iudam qui cognominatur Scarioth unum de duodecim
LUKE|22|4|et abiit et locutus est cum principibus sacerdotum et magistratibus quemadmodum illum traderet eis
LUKE|22|5|et gavisi sunt et pacti sunt pecuniam illi dare
LUKE|22|6|et spopondit et quaerebat oportunitatem ut traderet illum sine turbis
LUKE|22|7|venit autem dies azymorum in qua necesse erat occidi pascha
LUKE|22|8|et misit Petrum et Iohannem dicens euntes parate nobis pascha ut manducemus
LUKE|22|9|at illi dixerunt ubi vis paremus
LUKE|22|10|et dixit ad eos ecce introeuntibus vobis in civitatem occurret vobis homo amphoram aquae portans sequimini eum in domum in qua intrat
LUKE|22|11|et dicetis patri familias domus dicit tibi magister ubi est diversorium ubi pascha cum discipulis meis manducem
LUKE|22|12|et ipse vobis ostendet cenaculum magnum stratum et ibi parate
LUKE|22|13|euntes autem invenerunt sicut dixit illis et paraverunt pascha
LUKE|22|14|et cum facta esset hora discubuit et duodecim apostoli cum eo
LUKE|22|15|et ait illis desiderio desideravi hoc pascha manducare vobiscum antequam patiar
LUKE|22|16|dico enim vobis quia ex hoc non manducabo illud donec impleatur in regno Dei
LUKE|22|17|et accepto calice gratias egit et dixit accipite et dividite inter vos
LUKE|22|18|dico enim vobis quod non bibam de generatione vitis donec regnum Dei veniat
LUKE|22|19|et accepto pane gratias egit et fregit et dedit eis dicens hoc est corpus meum quod pro vobis datur hoc facite in meam commemorationem
LUKE|22|20|similiter et calicem postquam cenavit dicens hic est calix novum testamentum in sanguine meo quod pro vobis funditur
LUKE|22|21|verumtamen ecce manus tradentis me mecum est in mensa
LUKE|22|22|et quidem Filius hominis secundum quod definitum est vadit verumtamen vae illi homini per quem traditur
LUKE|22|23|et ipsi coeperunt quaerere inter se quis esset ex eis qui hoc facturus esset
LUKE|22|24|facta est autem et contentio inter eos quis eorum videretur esse maior
LUKE|22|25|dixit autem eis reges gentium dominantur eorum et qui potestatem habent super eos benefici vocantur
LUKE|22|26|vos autem non sic sed qui maior est in vobis fiat sicut iunior et qui praecessor est sicut ministrator
LUKE|22|27|nam quis maior est qui recumbit an qui ministrat nonne qui recumbit ego autem in medio vestrum sum sicut qui ministrat
LUKE|22|28|vos autem estis qui permansistis mecum in temptationibus meis
LUKE|22|29|et ego dispono vobis sicut disposuit mihi Pater meus regnum
LUKE|22|30|ut edatis et bibatis super mensam meam in regno et sedeatis super thronos iudicantes duodecim tribus Israhel
LUKE|22|31|ait autem Dominus Simon Simon ecce Satanas expetivit vos ut cribraret sicut triticum
LUKE|22|32|ego autem rogavi pro te ut non deficiat fides tua et tu aliquando conversus confirma fratres tuos
LUKE|22|33|qui dixit ei Domine tecum paratus sum et in carcerem et in mortem ire
LUKE|22|34|et ille dixit dico tibi Petre non cantabit hodie gallus donec ter abneges nosse me
LUKE|22|35|et dixit eis quando misi vos sine sacculo et pera et calciamentis numquid aliquid defuit vobis at illi dixerunt nihil
LUKE|22|36|dixit ergo eis sed nunc qui habet sacculum tollat similiter et peram et qui non habet vendat tunicam suam et emat gladium
LUKE|22|37|dico enim vobis quoniam adhuc hoc quod scriptum est oportet impleri in me et quod cum iniustis deputatus est etenim ea quae sunt de me finem habent
LUKE|22|38|at illi dixerunt Domine ecce gladii duo hic at ille dixit eis satis est
LUKE|22|39|et egressus ibat secundum consuetudinem in montem Olivarum secuti sunt autem illum et discipuli
LUKE|22|40|et cum pervenisset ad locum dixit illis orate ne intretis in temptationem
LUKE|22|41|et ipse avulsus est ab eis quantum iactus est lapidis et positis genibus orabat
LUKE|22|42|dicens Pater si vis transfer calicem istum a me verumtamen non mea voluntas sed tua fiat
LUKE|22|43|apparuit autem illi angelus de caelo confortans eum et factus in agonia prolixius orabat
LUKE|22|44|et factus est sudor eius sicut guttae sanguinis decurrentis in terram
LUKE|22|45|et cum surrexisset ab oratione et venisset ad discipulos suos invenit eos dormientes prae tristitia
LUKE|22|46|et ait illis quid dormitis surgite orate ne intretis in temptationem
LUKE|22|47|adhuc eo loquente ecce turba et qui vocabatur Iudas unus de duodecim antecedebat eos et adpropinquavit Iesu ut oscularetur eum
LUKE|22|48|Iesus autem dixit ei Iuda osculo Filium hominis tradis
LUKE|22|49|videntes autem hii qui circa ipsum erant quod futurum erat dixerunt ei Domine si percutimus in gladio
LUKE|22|50|et percussit unus ex illis servum principis sacerdotum et amputavit auriculam eius dextram
LUKE|22|51|respondens autem Iesus ait sinite usque huc et cum tetigisset auriculam eius sanavit eum
LUKE|22|52|dixit autem Iesus ad eos qui venerant ad se principes sacerdotum et magistratus templi et seniores quasi ad latronem existis cum gladiis et fustibus
LUKE|22|53|cum cotidie vobiscum fuerim in templo non extendistis manus in me sed haec est hora vestra et potestas tenebrarum
LUKE|22|54|conprehendentes autem eum duxerunt ad domum principis sacerdotum Petrus vero sequebatur a longe
LUKE|22|55|accenso autem igni in medio atrio et circumsedentibus illis erat Petrus in medio eorum
LUKE|22|56|quem cum vidisset ancilla quaedam sedentem ad lumen et eum fuisset intuita dixit et hic cum illo erat
LUKE|22|57|at ille negavit eum dicens mulier non novi illum
LUKE|22|58|et post pusillum alius videns eum dixit et tu de illis es Petrus vero ait o homo non sum
LUKE|22|59|et intervallo facto quasi horae unius alius quidam adfirmabat dicens vere et hic cum illo erat nam et Galilaeus est
LUKE|22|60|et ait Petrus homo nescio quod dicis et continuo adhuc illo loquente cantavit gallus
LUKE|22|61|et conversus Dominus respexit Petrum et recordatus est Petrus verbi Domini sicut dixit quia priusquam gallus cantet ter me negabis
LUKE|22|62|et egressus foras Petrus flevit amare
LUKE|22|63|et viri qui tenebant illum inludebant ei caedentes
LUKE|22|64|et velaverunt eum et percutiebant faciem eius et interrogabant eum dicentes prophetiza quis est qui te percussit
LUKE|22|65|et alia multa blasphemantes dicebant in eum
LUKE|22|66|et ut factus est dies convenerunt seniores plebis et principes sacerdotum et scribae et duxerunt illum in concilium suum dicentes si tu es Christus dic nobis
LUKE|22|67|et ait illis si vobis dixero non creditis mihi
LUKE|22|68|si autem et interrogavero non respondebitis mihi neque dimittetis
LUKE|22|69|ex hoc autem erit Filius hominis sedens a dextris virtutis Dei
LUKE|22|70|dixerunt autem omnes tu ergo es Filius Dei qui ait vos dicitis quia ego sum
LUKE|22|71|at illi dixerunt quid adhuc desideramus testimonium ipsi enim audivimus de ore eius
LUKE|23|1|et surgens omnis multitudo eorum duxerunt illum ad Pilatum
LUKE|23|2|coeperunt autem accusare illum dicentes hunc invenimus subvertentem gentem nostram et prohibentem tributa dari Caesari et dicentem se Christum regem esse
LUKE|23|3|Pilatus autem interrogavit eum dicens tu es rex Iudaeorum at ille respondens ait tu dicis
LUKE|23|4|ait autem Pilatus ad principes sacerdotum et turbas nihil invenio causae in hoc homine
LUKE|23|5|at illi invalescebant dicentes commovet populum docens per universam Iudaeam et incipiens a Galilaea usque huc
LUKE|23|6|Pilatus autem audiens Galilaeam interrogavit si homo Galilaeus esset
LUKE|23|7|et ut cognovit quod de Herodis potestate esset remisit eum ad Herodem qui et ipse Hierosolymis erat illis diebus
LUKE|23|8|Herodes autem viso Iesu gavisus est valde erat enim cupiens ex multo tempore videre eum eo quod audiret multa de illo et sperabat signum aliquod videre ab eo fieri
LUKE|23|9|interrogabat autem illum multis sermonibus at ipse nihil illi respondebat
LUKE|23|10|stabant etiam principes sacerdotum et scribae constanter accusantes eum
LUKE|23|11|sprevit autem illum Herodes cum exercitu suo et inlusit indutum veste alba et remisit ad Pilatum
LUKE|23|12|et facti sunt amici Herodes et Pilatus in ipsa die nam antea inimici erant ad invicem
LUKE|23|13|Pilatus autem convocatis principibus sacerdotum et magistratibus et plebe
LUKE|23|14|dixit ad illos obtulistis mihi hunc hominem quasi avertentem populum et ecce ego coram vobis interrogans nullam causam inveni in homine isto ex his in quibus eum accusatis
LUKE|23|15|sed neque Herodes nam remisi vos ad illum et ecce nihil dignum morte actum est ei
LUKE|23|16|emendatum ergo illum dimittam
LUKE|23|17|necesse autem habebat dimittere eis per diem festum unum
LUKE|23|18|exclamavit autem simul universa turba dicens tolle hunc et dimitte nobis Barabban
LUKE|23|19|qui erat propter seditionem quandam factam in civitate et homicidium missus in carcerem
LUKE|23|20|iterum autem Pilatus locutus est ad illos volens dimittere Iesum
LUKE|23|21|at illi succlamabant dicentes crucifige crucifige illum
LUKE|23|22|ille autem tertio dixit ad illos quid enim mali fecit iste nullam causam mortis invenio in eo corripiam ergo illum et dimittam
LUKE|23|23|at illi instabant vocibus magnis postulantes ut crucifigeretur et invalescebant voces eorum
LUKE|23|24|et Pilatus adiudicavit fieri petitionem eorum
LUKE|23|25|dimisit autem illis eum qui propter homicidium et seditionem missus fuerat in carcerem quem petebant Iesum vero tradidit voluntati eorum
LUKE|23|26|et cum ducerent eum adprehenderunt Simonem quendam Cyrenensem venientem de villa et inposuerunt illi crucem portare post Iesum
LUKE|23|27|sequebatur autem illum multa turba populi et mulierum quae plangebant et lamentabant eum
LUKE|23|28|conversus autem ad illas Iesus dixit filiae Hierusalem nolite flere super me sed super vos ipsas flete et super filios vestros
LUKE|23|29|quoniam ecce venient dies in quibus dicent beatae steriles et ventres qui non genuerunt et ubera quae non lactaverunt
LUKE|23|30|tunc incipient dicere montibus cadite super nos et collibus operite nos
LUKE|23|31|quia si in viridi ligno haec faciunt in arido quid fiet
LUKE|23|32|ducebantur autem et alii duo nequam cum eo ut interficerentur
LUKE|23|33|et postquam venerunt in locum qui vocatur Calvariae ibi crucifixerunt eum et latrones unum a dextris et alterum a sinistris
LUKE|23|34|Iesus autem dicebat Pater dimitte illis non enim sciunt quid faciunt dividentes vero vestimenta eius miserunt sortes
LUKE|23|35|et stabat populus expectans et deridebant illum principes cum eis dicentes alios salvos fecit se salvum faciat si hic est Christus Dei electus
LUKE|23|36|inludebant autem ei et milites accedentes et acetum offerentes illi
LUKE|23|37|dicentes si tu es rex Iudaeorum salvum te fac
LUKE|23|38|erat autem et superscriptio inscripta super illum litteris graecis et latinis et hebraicis hic est rex Iudaeorum
LUKE|23|39|unus autem de his qui pendebant latronibus blasphemabat eum dicens si tu es Christus salvum fac temet ipsum et nos
LUKE|23|40|respondens autem alter increpabat illum dicens neque tu times Deum quod in eadem damnatione es
LUKE|23|41|et nos quidem iuste nam digna factis recipimus hic vero nihil mali gessit
LUKE|23|42|et dicebat ad Iesum Domine memento mei cum veneris in regnum tuum
LUKE|23|43|et dixit illi Iesus amen dico tibi hodie mecum eris in paradiso
LUKE|23|44|erat autem fere hora sexta et tenebrae factae sunt in universa terra usque in nonam horam
LUKE|23|45|et obscuratus est sol et velum templi scissum est medium
LUKE|23|46|et clamans voce magna Iesus ait Pater in manus tuas commendo spiritum meum et haec dicens exspiravit
LUKE|23|47|videns autem centurio quod factum fuerat glorificavit Deum dicens vere hic homo iustus erat
LUKE|23|48|et omnis turba eorum qui simul aderant ad spectaculum istud et videbant quae fiebant percutientes pectora sua revertebantur
LUKE|23|49|stabant autem omnes noti eius a longe et mulieres quae secutae erant eum a Galilaea haec videntes
LUKE|23|50|et ecce vir nomine Ioseph qui erat decurio vir bonus et iustus
LUKE|23|51|hic non consenserat consilio et actibus eorum ab Arimathia civitate Iudaeae qui expectabat et ipse regnum Dei
LUKE|23|52|hic accessit ad Pilatum et petiit corpus Iesu
LUKE|23|53|et depositum involvit sindone et posuit eum in monumento exciso in quo nondum quisquam positus fuerat
LUKE|23|54|et dies erat parasceves et sabbatum inlucescebat
LUKE|23|55|subsecutae autem mulieres quae cum ipso venerant de Galilaea viderunt monumentum et quemadmodum positum erat corpus eius
LUKE|23|56|et revertentes paraverunt aromata et unguenta et sabbato quidem siluerunt secundum mandatum
LUKE|24|1|una autem sabbati valde diluculo venerunt ad monumentum portantes quae paraverant aromata
LUKE|24|2|et invenerunt lapidem revolutum a monumento
LUKE|24|3|et ingressae non invenerunt corpus Domini Iesu
LUKE|24|4|et factum est dum mente consternatae essent de isto ecce duo viri steterunt secus illas in veste fulgenti
LUKE|24|5|cum timerent autem et declinarent vultum in terram dixerunt ad illas quid quaeritis viventem cum mortuis
LUKE|24|6|non est hic sed surrexit recordamini qualiter locutus est vobis cum adhuc in Galilaea esset
LUKE|24|7|dicens quia oportet Filium hominis tradi in manus hominum peccatorum et crucifigi et die tertia resurgere
LUKE|24|8|et recordatae sunt verborum eius
LUKE|24|9|et regressae a monumento nuntiaverunt haec omnia illis undecim et ceteris omnibus
LUKE|24|10|erat autem Maria Magdalene et Iohanna et Maria Iacobi et ceterae quae cum eis erant quae dicebant ad apostolos haec
LUKE|24|11|et visa sunt ante illos sicut deliramentum verba ista et non credebant illis
LUKE|24|12|Petrus autem surgens cucurrit ad monumentum et procumbens videt linteamina sola posita et abiit secum mirans quod factum fuerat
LUKE|24|13|et ecce duo ex illis ibant ipsa die in castellum quod erat in spatio stadiorum sexaginta ab Hierusalem nomine Emmaus
LUKE|24|14|et ipsi loquebantur ad invicem de his omnibus quae acciderant
LUKE|24|15|et factum est dum fabularentur et secum quaererent et ipse Iesus adpropinquans ibat cum illis
LUKE|24|16|oculi autem illorum tenebantur ne eum agnoscerent
LUKE|24|17|et ait ad illos qui sunt hii sermones quos confertis ad invicem ambulantes et estis tristes
LUKE|24|18|et respondens unus cui nomen Cleopas dixit ei tu solus peregrinus es in Hierusalem et non cognovisti quae facta sunt in illa his diebus
LUKE|24|19|quibus ille dixit quae et dixerunt de Iesu Nazareno qui fuit vir propheta potens in opere et sermone coram Deo et omni populo
LUKE|24|20|et quomodo eum tradiderunt summi sacerdotum et principes nostri in damnationem mortis et crucifixerunt eum
LUKE|24|21|nos autem sperabamus quia ipse esset redempturus Israhel et nunc super haec omnia tertia dies hodie quod haec facta sunt
LUKE|24|22|sed et mulieres quaedam ex nostris terruerunt nos quae ante lucem fuerunt ad monumentum
LUKE|24|23|et non invento corpore eius venerunt dicentes se etiam visionem angelorum vidisse qui dicunt eum vivere
LUKE|24|24|et abierunt quidam ex nostris ad monumentum et ita invenerunt sicut mulieres dixerunt ipsum vero non viderunt
LUKE|24|25|et ipse dixit ad eos o stulti et tardi corde ad credendum in omnibus quae locuti sunt prophetae
LUKE|24|26|nonne haec oportuit pati Christum et ita intrare in gloriam suam
LUKE|24|27|et incipiens a Mose et omnibus prophetis interpretabatur illis in omnibus scripturis quae de ipso erant
LUKE|24|28|et adpropinquaverunt castello quo ibant et ipse se finxit longius ire
LUKE|24|29|et coegerunt illum dicentes mane nobiscum quoniam advesperascit et inclinata est iam dies et intravit cum illis
LUKE|24|30|et factum est dum recumberet cum illis accepit panem et benedixit ac fregit et porrigebat illis
LUKE|24|31|et aperti sunt oculi eorum et cognoverunt eum et ipse evanuit ex oculis eorum
LUKE|24|32|et dixerunt ad invicem nonne cor nostrum ardens erat in nobis dum loqueretur in via et aperiret nobis scripturas
LUKE|24|33|et surgentes eadem hora regressi sunt in Hierusalem et invenerunt congregatos undecim et eos qui cum ipsis erant
LUKE|24|34|dicentes quod surrexit Dominus vere et apparuit Simoni
LUKE|24|35|et ipsi narrabant quae gesta erant in via et quomodo cognoverunt eum in fractione panis
LUKE|24|36|dum haec autem loquuntur Iesus stetit in medio eorum et dicit eis pax vobis ego sum nolite timere
LUKE|24|37|conturbati vero et conterriti existimabant se spiritum videre
LUKE|24|38|et dixit eis quid turbati estis et cogitationes ascendunt in corda vestra
LUKE|24|39|videte manus meas et pedes quia ipse ego sum palpate et videte quia spiritus carnem et ossa non habet sicut me videtis habere
LUKE|24|40|et cum hoc dixisset ostendit eis manus et pedes
LUKE|24|41|adhuc autem illis non credentibus et mirantibus prae gaudio dixit habetis hic aliquid quod manducetur
LUKE|24|42|at illi obtulerunt ei partem piscis assi et favum mellis
LUKE|24|43|et cum manducasset coram eis sumens reliquias dedit eis
LUKE|24|44|et dixit ad eos haec sunt verba quae locutus sum ad vos cum adhuc essem vobiscum quoniam necesse est impleri omnia quae scripta sunt in lege Mosi et prophetis et psalmis de me
LUKE|24|45|tunc aperuit illis sensum ut intellegerent scripturas
LUKE|24|46|et dixit eis quoniam sic scriptum est et sic oportebat Christum pati et resurgere a mortuis die tertia
LUKE|24|47|et praedicari in nomine eius paenitentiam et remissionem peccatorum in omnes gentes incipientibus ab Hierosolyma
LUKE|24|48|vos autem estis testes horum
LUKE|24|49|et ego mitto promissum Patris mei in vos vos autem sedete in civitate quoadusque induamini virtutem ex alto
LUKE|24|50|eduxit autem eos foras in Bethaniam et elevatis manibus suis benedixit eis
LUKE|24|51|et factum est dum benediceret illis recessit ab eis et ferebatur in caelum
LUKE|24|52|et ipsi adorantes regressi sunt in Hierusalem cum gaudio magno
LUKE|24|53|et erant semper in templo laudantes et benedicentes Deum amen
