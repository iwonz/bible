ISA|1|1|当 乌西雅 、 约坦 、 亚哈斯 、 希西家 作 犹大 王的时候， 亚摩斯 的儿子 以赛亚 见异象，论到 犹大 和 耶路撒冷 。
ISA|1|2|天哪，要听！地啊，侧耳而听！ 因为耶和华说： “我养育儿女，将他们养大， 他们竟悖逆我。
ISA|1|3|牛认识主人， 驴认识主人的槽； 以色列 却不认识， 我的民却不明白。”
ISA|1|4|祸哉！犯罪的国民， 担着罪孽的百姓， 行恶的族类， 败坏的儿女！ 他们离弃耶和华， 藐视 以色列 的圣者， 背向他，与他疏远。
ISA|1|5|你们为什么屡次悖逆，继续受责打呢？ 你们已经满头疼痛， 全心发昏；
ISA|1|6|从脚掌到头顶， 没有一处是完好的， 尽是创伤、瘀青，与流血的伤口， 未曾挤净，未曾包扎， 也没有用膏滋润。
ISA|1|7|你们的土地荒芜， 城镇被火烧毁； 你们的田地在你们眼前被陌生人侵吞， 既被陌生人倾覆，就成为荒芜 。
ISA|1|8|仅存的 锡安 ， 好似葡萄园的草棚， 如瓜田中的茅屋， 又如被围困的城。
ISA|1|9|若不是万军之耶和华为我们留下一些幸存者， 我们早已变成 所多玛 ，像 蛾摩拉 一样了。
ISA|1|10|所多玛 的官长啊， 你们要听耶和华的言语！ 蛾摩拉 的百姓啊， 要侧耳听我们上帝的教诲！
ISA|1|11|耶和华说： “你们许多的祭物于我何益呢？ 公绵羊的燔祭和肥畜的油脂， 我已经腻烦了； 公牛、羔羊、公山羊的血， 我都不喜悦。
ISA|1|12|“你们来朝见我， 谁向你们的手要求这些， 使你们践踏我的院宇呢？
ISA|1|13|不要再献无谓的供物了， 香是我所憎恶的。 我不能容忍行恶又守严肃会： 初一、安息日和召集的大会。
ISA|1|14|你们的初一和节期，我心里恨恶， 它们成了我的重担， 担当这些，令我厌烦。
ISA|1|15|你们举手祷告，我必遮眼不看， 就算你们多多祈祷，我也不听； 你们的手沾满了血。
ISA|1|16|你们要洗涤、自洁， 从我眼前除掉恶行； 要停止作恶，
ISA|1|17|学习行善， 寻求公平， 帮助受欺压的 ， 替孤儿伸冤， 为寡妇辩护。”
ISA|1|18|耶和华说： “来吧，我们彼此辩论。 你们的罪虽像朱红，必变成雪白； 虽红如丹颜，必白如羊毛。
ISA|1|19|你们若甘心听从， 必吃地上的美物；
ISA|1|20|若不听从，反倒悖逆， 必被刀剑吞灭； 这是耶和华亲口说的。”
ISA|1|21|忠信的城竟然变为妓女！ 从前充满了公平， 公义居在其中， 现今却有凶手居住。
ISA|1|22|你的银子变为渣滓， 你的酒用水冲淡。
ISA|1|23|你的官长悖逆， 与盗贼为伍， 全都喜爱贿赂， 追求赃物； 他们不为孤儿伸冤， 寡妇的案件也呈不到他们面前。
ISA|1|24|因此，主－万军之耶和华、 以色列 的大能者说： “唉！我要向我的对头雪恨， 向我的敌人报仇。
ISA|1|25|我必反手对付你， 如碱炼净你的渣滓， 除尽你的杂质。
ISA|1|26|我必回复你的审判官，像起初一样， 回复你的谋士，如起先一般。 然后，你必称为公义之城， 忠信之邑。”
ISA|1|27|锡安 必因公平得蒙救赎， 其中归正的人必因公义得蒙救赎。
ISA|1|28|但悖逆的和犯罪的必一同败亡， 离弃耶和华的必致消灭。
ISA|1|29|那等人必因所喜爱的圣树抱愧； 你们必因所选择的园子 蒙羞，
ISA|1|30|因为你们必如叶子枯干的橡树， 如无水的园子。
ISA|1|31|有权势的必如麻线， 他的作为好像火花， 都要一同焚烧，无人扑灭。
ISA|2|1|亚摩斯 的儿子 以赛亚 所见，有关 犹大 和 耶路撒冷 的事。
ISA|2|2|末后的日子，耶和华殿的山必坚立， 超乎诸山，高举过于万岭； 万国都要流归这山。
ISA|2|3|必有许多民族前往，说： “来吧，我们登耶和华的山， 到 雅各 上帝的殿。 他必将他的道教导我们， 我们也要行他的路。” 因为教诲必出于 锡安 ， 耶和华的言语必出于 耶路撒冷 。
ISA|2|4|他必在万国中施行审判， 为许多民族断定是非。 他们要将刀打成犁头， 把枪打成镰刀； 这国不举刀攻击那国， 他们也不再学习战事。
ISA|2|5|雅各 家啊， 来吧！让我们在耶和华的光明中行走。
ISA|2|6|你离弃了你的百姓 雅各 家， 因为他们充满了东方的习俗 ， 又像 非利士 人一样观星象， 并与外邦人击掌。
ISA|2|7|他们的国满了金银， 财宝也无穷； 他们的地满了马匹， 战车也无数。
ISA|2|8|他们的地满了偶像； 他们跪拜自己手所造的， 就是自己手指所做的。
ISA|2|9|有人屈膝， 有人下跪； 所以，不要饶恕他们。
ISA|2|10|当进入磐石，藏在土中， 躲避耶和华的惊吓和他威严的荣光。
ISA|2|11|到那日，眼目高傲的必降卑， 狂妄的人必屈膝； 惟独耶和华被尊崇。
ISA|2|12|因万军之耶和华的一个日子 要临到所有骄傲狂妄的， 临到一切自高的， 使他们降为卑；
ISA|2|13|临到 黎巴嫩 高大的香柏树、 巴珊 的橡树，
ISA|2|14|临到一切高山、 一切峻岭，
ISA|2|15|临到一切碉堡、 一切坚固的城墙，
ISA|2|16|临到 他施 一切的船只、 一切华丽的船艇。
ISA|2|17|人的骄傲必屈膝， 人的狂妄必降卑； 在那日，惟独耶和华被尊崇，
ISA|2|18|偶像必全然废弃。
ISA|2|19|耶和华兴起使地大震动的时候， 人就进入石洞和土穴里， 躲避耶和华的惊吓和他威严的荣光。
ISA|2|20|到那日，人必将造来敬拜的金偶像、银偶像 抛给田鼠和蝙蝠。
ISA|2|21|耶和华兴起使地大震动的时候， 人就进入磐缝和岩隙里， 躲避耶和华的惊吓和他威严的荣光。
ISA|2|22|你们不要倚靠世人， 他只不过鼻孔里有气息， 算得了什么呢？
ISA|3|1|看哪，主－万军之耶和华要从 耶路撒冷 和 犹大 除掉众人所倚靠的，所仰赖的， 就是所倚靠的粮，所仰赖的水；
ISA|3|2|除掉勇士和战士， 审判官和先知， 占卜的和长老，
ISA|3|3|除掉五十夫长和显要、 谋士和巧匠， 以及擅长法术的人。
ISA|3|4|我必使孩童作他们的领袖， 幼儿管辖他们。
ISA|3|5|百姓要彼此欺压， 各人欺压邻舍； 青年要侮慢老人， 卑贱的要侮慢尊贵的。
ISA|3|6|人在父家拉住自己的兄弟： “你有外衣，来作我们的官长， 让这些败坏的事归于你的手下吧！”
ISA|3|7|那时，他必扬声说： “我不作医治你们的人； 我家里没有粮食，也没有衣服， 你们不可立我作百姓的官长。”
ISA|3|8|耶路撒冷 败落， 犹大 倾倒； 因为他们的舌头和行为与耶和华相悖， 无视于他荣光的眼目。
ISA|3|9|他们的脸色证明自己不正， 他们述说自己像 所多玛 一样的罪恶，毫不隐瞒。 他们有祸了！因为作恶自害。
ISA|3|10|你们要对义人说，他是有福的， 因为他必吃自己行为所结的果实。
ISA|3|11|恶人有祸了！他必遭灾难！ 因为他要按自己手所做的受报应。
ISA|3|12|至于我的百姓， 统治者剥削你们， 放高利贷的人管辖你们 。 我的百姓啊，引导你的使你走错， 并毁坏你所行的道路。
ISA|3|13|耶和华兴起诉讼， 站着审判万民。
ISA|3|14|耶和华必审问他国中的长老和领袖： “你们，你们摧毁葡萄园， 抢夺困苦人，囤积在你们家中。
ISA|3|15|你们为何压碎我的百姓， 碾磨困苦人的脸呢？” 这是万军之主耶和华说的。
ISA|3|16|耶和华说： 因为 锡安 狂傲， 行走挺项，卖弄眼目， 俏步徐行，脚下玎珰，
ISA|3|17|主必使 锡安 头顶长疮， 耶和华又暴露其下体。
ISA|3|18|到那日，主必除掉华美的足饰、额带、月牙圈、
ISA|3|19|耳环、手镯、面纱、
ISA|3|20|头巾、足链、华带、香盒、符囊、
ISA|3|21|戒指、鼻环、
ISA|3|22|礼服、外套、披肩、皮包、
ISA|3|23|手镜、细麻衣、头饰、纱巾。
ISA|3|24|必有腐烂代替馨香， 绳子代替腰带， 光秃代替美发， 麻衣系腰代替华服， 烙痕代替美貌。
ISA|3|25|你的男丁必倒在刀下， 你的勇士必死在阵上。
ISA|3|26|锡安 的城门必悲伤、哀号； 它必荒凉，坐在地上。
ISA|4|1|在那日，七个女人必拉住一个男人，说：“我们吃自己的食物，穿自己的衣服，但求你允许我们归你名下，除掉我们的羞耻。”
ISA|4|2|在那日，耶和华的苗必华美尊荣，地的出产必成为幸存的 以色列 民的骄傲和光荣。
ISA|4|3|主以公平的灵和焚烧的灵洗净 锡安 居民 的污秽，又除净在 耶路撒冷 流人血的罪。那时，剩在 锡安 、留在 耶路撒冷 的，就是一切住 耶路撒冷 、在生命册上记名的，必称为圣。
ISA|4|4|
ISA|4|5|耶和华必在整座 锡安山 ，在会众之上，白天造云，黑夜发出烟和火焰的光，因为在一切荣耀之上必有华盖；
ISA|4|6|这要作为棚子，白天可以遮荫避暑，暴风雨侵袭时，可作藏身处和避难所。
ISA|5|1|我要为我亲爱的唱歌， 我所爱的、他的葡萄园之歌。 我亲爱的有葡萄园 在肥沃的山冈上。
ISA|5|2|他刨挖园子，清除石头， 栽种上等的葡萄树， 在园中盖了一座楼， 又凿出酒池； 指望它结葡萄， 反倒结了野葡萄。
ISA|5|3|耶路撒冷 的居民和 犹大 人哪， 现在，请你们在我与我的葡萄园之间断定是非。
ISA|5|4|我为我葡萄园所做的之外， 还有什么可做的呢？ 我指望它结葡萄， 怎么倒结了野葡萄呢？
ISA|5|5|现在我告诉你们， 我要向我的葡萄园怎么做。 我必撤去篱笆，使它被烧毁； 拆毁围墙，使它被践踏。
ISA|5|6|我必使它荒废，不再修剪， 不再锄草，任荆棘蒺藜生长； 我也必吩咐密云， 不再降雨在其上。
ISA|5|7|万军之耶和华的葡萄园就是 以色列 家； 他所喜爱的树就是 犹大 人。 他指望公平， 看哪，却有流血； 指望公义， 看哪，却有冤声。
ISA|5|8|祸哉！你们以房接房， 以地连地， 以致不留余地， 只顾自己独居境内。
ISA|5|9|我耳闻万军之耶和华说： “许多房屋必然荒废； 宏伟华丽，无人居住。
ISA|5|10|十亩 的葡萄园只酿出一罢特的酒， 一贺梅珥的谷种只结一伊法粮食。”
ISA|5|11|祸哉！那些清晨早起，追寻烈酒， 因酒狂热，流连到深夜的人，
ISA|5|12|他们在宴席上 弹琴，鼓瑟，击鼓，吹笛，饮酒， 却不留意耶和华的作为， 也不留心他手所做的。
ISA|5|13|所以，我的百姓因无知就被掳去； 尊贵的人甚是饥饿， 平民也极其干渴。
ISA|5|14|因此，阴间胃口 大开， 张开无限量的口； 令 耶路撒冷 的贵族与平民、狂欢的与作乐的人 都掉落其中。
ISA|5|15|人为之屈膝， 人就降为卑； 高傲的眼目也降为卑。
ISA|5|16|惟有万军之耶和华因公平显为崇高， 神圣的上帝因公义显为圣。
ISA|5|17|羔羊必来吃草，如同在自己的草场； 在富有人的废墟，流浪的牲畜也来吃 。
ISA|5|18|祸哉！那些以虚假的绳子牵引罪孽， 以套车的绳索紧拉罪恶的人。
ISA|5|19|他们说： “任 以色列 的圣者急速前行，快快成就他的作为， 好让我们看看； 任他的筹算临近成就， 好使我们知道。”
ISA|5|20|祸哉！那些称恶为善，称善为恶， 以暗为光，以光为暗， 以苦为甜，以甜为苦的人。
ISA|5|21|祸哉！那些在自己眼中有智慧， 在自己面前有通达的人。
ISA|5|22|祸哉！那些以饮酒称雄， 以调烈酒称霸的人。
ISA|5|23|他们因受贿赂，就称恶人为义， 将义人的义夺去。
ISA|5|24|火苗怎样吞灭碎秸， 干草怎样落在火焰之中， 照样，他们的根必然腐朽， 他们的花像灰尘扬起； 因为他们厌弃万军之耶和华的教诲， 藐视 以色列 圣者的言语。
ISA|5|25|因此，耶和华的怒气向他的百姓发作。 他伸手攻击他们，山岭就震动； 他们的尸首在街市上好像粪土。 虽然如此，他的怒气并未转消， 他的手依然伸出。
ISA|5|26|他必竖立大旗，召集远方的国民， 把他们从地极叫来。 看哪，他们必急速奔来，
ISA|5|27|其中没有疲倦的，绊跌的； 没有打盹的，睡觉的； 腰带并不放松， 鞋带也不拉断。
ISA|5|28|他们的箭锐利， 弓也上了弦； 马蹄如坚石， 车轮像旋风。
ISA|5|29|他们要吼叫，像母狮， 咆哮，像少壮狮子； 他们要咆哮，抓取猎物， 稳稳叼走，无人能救回。
ISA|5|30|那日，他们要向 以色列 人咆哮， 像海浪澎湃； 人若望地，看哪，只有黑暗与祸患， 光明因密云而变黑暗。
ISA|6|1|当 乌西雅 王崩的那年，我看见主坐在高高的宝座上。他的衣裳下摆遮满圣殿。
ISA|6|2|上有撒拉弗侍立，各有六个翅膀：两个翅膀遮脸，两个翅膀遮脚，两个翅膀飞翔，
ISA|6|3|彼此呼喊说： “圣哉！圣哉！圣哉！万军之耶和华； 他的荣光遍满全地！”
ISA|6|4|因呼喊者的声音，门槛的根基震动，殿里充满了烟云。
ISA|6|5|那时我说：“祸哉！我灭亡了！因为我是嘴唇不洁的人，住在嘴唇不洁的民中，又因我亲眼看见大君王－万军之耶和华。”
ISA|6|6|有一撒拉弗向我飞来，手里拿着烧红的炭，是用火钳从坛上取下来的，
ISA|6|7|用炭沾我的口，说：“看哪，这炭沾了你的嘴唇，你的罪孽便除掉，你的罪恶就赦免了。”
ISA|6|8|我听见主的声音说：“我可以差遣谁呢？谁肯为我们去呢？”我说：“我在这里，请差遣我！”
ISA|6|9|他说：“你去告诉这百姓说： ‘你们听了又听，却不明白； 看了又看，却不晓得。’
ISA|6|10|要使这百姓心蒙油脂， 耳朵发沉， 眼睛昏花； 恐怕他们眼睛看见， 耳朵听见， 心里明白， 回转过来，就得医治。”
ISA|6|11|我就说：“主啊，这到几时为止呢？”他说： “直到城镇荒凉，无人居住， 房屋空无一人，土地极其荒芜；
ISA|6|12|耶和华将人迁到远方， 国内被撇弃的土地很多。
ISA|6|13|国内剩下的人若还有十分之一， 也必被吞灭。 然而如同大树与橡树，虽被砍伐， 残干却仍存留， 圣洁的苗裔是它的残干。”
ISA|7|1|乌西雅 的孙子， 约坦 的儿子， 犹大 王 亚哈斯 在位的时候， 亚兰 王 利汛 和 利玛利 的儿子 以色列 王 比加 上来攻打 耶路撒冷 ，却不能攻取。
ISA|7|2|有人告诉 大卫 家说：“ 亚兰 与 以法莲 已经结盟。”王的心和百姓的心就都颤动，好像林中的树被风吹动一样。
ISA|7|3|耶和华对 以赛亚 说：“你和你的儿子 施亚．雅述 要出去，到 上池 的水沟尽头，往漂布地的大路上，迎见 亚哈斯 ，
ISA|7|4|对他说：‘你要谨慎，要镇定，不要害怕，不要因 利汛 和 亚兰 ，以及 利玛利 的儿子这两个冒烟火把的头所发的烈怒而心里胆怯。
ISA|7|5|因为 亚兰 、 以法莲 ，和 利玛利 的儿子设恶谋要害你，说：
ISA|7|6|我们要上去攻击 犹大 ，扰乱它，攻破它来归我们，在其中立 他比勒 的儿子为王。
ISA|7|7|主耶和华如此说： 这事必站立不住， 也不得成就。
ISA|7|8|因为 亚兰 的首都是 大马士革 ， 大马士革 的领袖是 利汛 ； 六十五年之内， 以法莲 必然国破族亡，
ISA|7|9|以法莲 的首都是 撒玛利亚 ； 撒玛利亚 的领袖是 利玛利 的儿子。 你们若是不信， 必站立不稳。’”
ISA|7|10|耶和华又吩咐 亚哈斯 ：
ISA|7|11|“你向耶和华－你的上帝求一个预兆：在阴间的深渊，或往上的高处。”
ISA|7|12|但 亚哈斯 说：“我不求；我不试探耶和华。”
ISA|7|13|以赛亚 说：“听啊， 大卫 家！你们使人厌烦岂算小事，还要使我的上帝厌烦吗？
ISA|7|14|因此，主自己要给你们一个预兆，看哪，必有童女怀孕生子，给他起名叫 以马内利 。
ISA|7|15|到他晓得弃恶择善的时候，他必吃乳酪与蜂蜜。
ISA|7|16|因为在这孩子还不晓得弃恶择善之先，你所憎恶的那两个王的土地必被撇弃。
ISA|7|17|耶和华必使 亚述 王临到你和你的百姓，并你的父家，自从 以法莲 脱离 犹大 的时候，未曾有过这样的日子。
ISA|7|18|“那时，耶和华要呼叫，召来 埃及 江河源头的苍蝇和 亚述 地的蜂；
ISA|7|19|它们都必飞来，停在陡峭的谷中、岩石缝里、一切荆棘丛中和片片草场上。
ISA|7|20|“那时，主必用 大河 外雇来的剃刀，就是 亚述 王，剃去你的头发和脚毛，并要剃净你的胡须。
ISA|7|21|“那时，每一个人要养活一头母牛犊和两只母羊；
ISA|7|22|因为奶量充足，他就有乳酪可吃，国内剩余的人也都能吃乳酪与蜂蜜。
ISA|7|23|“那时，凡种一千棵葡萄树、价值一千银子的地方，必长出荆棘和蒺藜。
ISA|7|24|人到那里去，必带弓箭，因为遍地长满了荆棘和蒺藜。
ISA|7|25|所有锄头刨过的山地，你因惧怕荆棘和蒺藜，不敢到那里去；只能作放牛之处，羊群践踏之地。”
ISA|8|1|耶和华对我说：“你取一块大板子，拿人的笔 ，写上‘玛黑珥．沙拉勒．哈施．罢斯’ 。
ISA|8|2|我 要用可靠的证人， 乌利亚 祭司和 耶比利家 的儿子 撒迦利亚 为我作证。”
ISA|8|3|我亲近女先知 ；她就怀孕生子，耶和华对我说：“给他起名叫 玛黑珥．沙拉勒．哈施．罢斯 ；
ISA|8|4|因为在这孩子还不晓得叫爸爸妈妈以前， 大马士革 的财宝和 撒玛利亚 的掳物必被 亚述 王掠夺一空。”
ISA|8|5|耶和华又吩咐我：
ISA|8|6|“这百姓既厌弃 西罗亚 缓流的水，喜欢 利汛 以及 利玛利 的儿子，
ISA|8|7|因此，看哪，主必使 亚述 王和他的威势如 大河 翻腾汹涌的水上涨，盖过他们，必上涨超过一切水道，涨过两岸，
ISA|8|8|必冲入 犹大 ，涨溢泛滥，直到颈项。他展开翅膀，遮蔽你的全地。 以马内利 啊！”
ISA|8|9|万民哪，任凭你们行恶 ，终必毁灭； 远方的众人哪，当侧耳而听！ 任凭你们束腰，终必毁灭； 你们束起腰来，终必毁灭。
ISA|8|10|任凭你们筹算什么，终必无效； 不管你们讲定什么，总不成立； 因为上帝与我们同在。
ISA|8|11|耶和华以大能的手训诫我不可行 这百姓所行的道，对我这样说：
ISA|8|12|“这百姓说同谋背叛的，你们不要说同谋背叛。他们所怕的，你们不要怕，也不要畏惧；
ISA|8|13|但要尊万军之耶和华为圣，他才是你们所当怕的，所当畏惧的。
ISA|8|14|他必作为圣所，却向 以色列 的两家成为绊脚的石头，使人跌倒的磐石；作 耶路撒冷 居民的罗网和圈套。
ISA|8|15|许多人在其上绊倒，他们跌倒，甚至跌伤，并且落入陷阱，被抓住了。”
ISA|8|16|你要卷起律法书，在我门徒中间封住教诲。
ISA|8|17|我要等候那转脸不顾 雅各 家的耶和华，也要仰望他。
ISA|8|18|看哪，我与耶和华所赐给我的儿女成了 以色列 的预兆和奇迹，这是从住在 锡安山 万军之耶和华来的。
ISA|8|19|有人对你们说：“当求问招魂的与行巫术的，他们唧唧喳喳，念念有词。”然而，百姓不当求问自己的上帝吗？岂可为活人求问死人呢？
ISA|8|20|当以教诲和律法书为准；人所说的若不与此相符，必没有黎明。
ISA|8|21|他必经过这地，遇艰难，受饥饿；饥饿的时候，心中焦躁，咒骂自己的君王和上帝。他仰观上天，
ISA|8|22|俯察下地，看哪，尽是艰难、黑暗和骇人的昏暗。他必被赶入幽暗中去。
ISA|9|1|但那受过痛苦的必不再见幽暗。 从前上帝使 西布伦 地和 拿弗他利 地被藐视，末后却使这沿海的路， 约旦河 东，外邦人居住的 加利利 地得荣耀。
ISA|9|2|在黑暗中行走的百姓看见了大光； 住在死荫之地的人有光照耀他们。
ISA|9|3|你使这国民众多 ， 使他们喜乐大增； 他们在你面前欢喜， 好像收割时的欢喜， 又像人分战利品那样的快乐。
ISA|9|4|因为他们所负的重轭 和肩头上的杖， 并欺压者的棍， 你都已经折断， 如同在 米甸 的日子一般。
ISA|9|5|战士在战乱中所穿的靴子， 以及那滚在血中的衣服， 都必当作柴火燃烧。
ISA|9|6|因有一婴孩为我们而生； 有一子赐给我们。 政权必担在他的肩头上； 他名称为“奇妙策士、全能的上帝、永在的父、和平的君”。
ISA|9|7|他的政权与平安必加增无穷。 他必在 大卫 的宝座上治理他的国， 以公平公义使国坚定稳固， 从今直到永远。 万军之耶和华的热心必成就这事。
ISA|9|8|主向 雅各 家发出言语， 主的话临到 以色列 家。
ISA|9|9|众百姓，就是 以法莲 和 撒玛利亚 的居民， 都将知道； 他们凭骄傲自大的心说：
ISA|9|10|“砖块掉落了，我们要凿石头重建； 桑树砍了，我们要改种香柏树。”
ISA|9|11|因此，耶和华兴起 利汛 的敌人 前来攻击 以色列 ， 要激起它的仇敌，
ISA|9|12|东有 亚兰 人，西有 非利士 人； 他们张口吞吃 以色列 。 虽然如此，耶和华的怒气并未转消； 他的手依然伸出。
ISA|9|13|这百姓还没有归向击打他们的主， 也没有寻求万军之耶和华。
ISA|9|14|耶和华在一日之间 从 以色列 中剪除了头与尾－ 棕树枝与芦苇－
ISA|9|15|长老和显要就是头， 以谎言教人的先知就是尾。
ISA|9|16|因为引导这百姓的使他们走入迷途， 被引导的都必被吞灭。
ISA|9|17|所以，主不喜爱 他们的青年， 也不怜悯他们的孤儿和寡妇； 因为他们都是亵渎的，行恶的， 并且各人的口都说愚妄的话。 虽然如此，耶和华的怒气并未转消； 他的手依然伸出。
ISA|9|18|邪恶如火焚烧， 吞灭荆棘和蒺藜， 在稠密的树林中点燃， 成为烟柱，旋转上腾。
ISA|9|19|因万军之耶和华的烈怒，地都烧遍了； 百姓成为柴火， 无人怜惜弟兄。
ISA|9|20|有人右边抢夺，犹受饥饿； 左边吞吃，仍不饱足， 各人吃自己膀臂上的肉。
ISA|9|21|玛拿西 吞吃 以法莲 ， 以法莲 吞吃 玛拿西 ， 他们又一同攻击 犹大 。 虽然如此，耶和华的怒气并未转消； 他的手依然伸出。
ISA|10|1|祸哉！那些设立不义之律例的， 和记录奸诈之判词的，
ISA|10|2|为要扭曲贫寒人的案件， 夺去我民中困苦人的理， 以寡妇当作掳物， 以孤儿当作掠物。
ISA|10|3|到降罚的日子，灾祸从远方临到， 那时，你们要怎么办呢？ 你们要向谁逃奔求救呢？ 你们的财宝要存放何处呢？
ISA|10|4|他们只得屈身在被掳的人之下， 仆倒在被杀的人中间 。 虽然如此，耶和华的怒气并未转消； 他的手依然伸出。
ISA|10|5|祸哉！ 亚述 ，我怒气的棍！ 他们手中的杖是我的恼恨。
ISA|10|6|我要差遣他攻击亵渎的国， 吩咐他对付我所恼怒的民， 抢走掳物，夺取掠物， 将他们践踏，如同街上的泥土一般。
ISA|10|7|然而，这并非他的意念， 他的心不是这样打算； 他的心要摧毁， 要剪除不少的国家。
ISA|10|8|他说：“我的官长岂不都是君王吗？
ISA|10|9|迦勒挪 岂不像 迦基米施 吗？ 哈马 岂不像 亚珥拔 吗？ 撒玛利亚 岂不像 大马士革 吗？
ISA|10|10|既然我的手已伸到了这些有偶像的国， 他们所雕刻的偶像 过于 耶路撒冷 和 撒玛利亚 的偶像，
ISA|10|11|我岂不照样待 耶路撒冷 和其中的偶像， 如同我待 撒玛利亚 和其中的偶像吗？”
ISA|10|12|主在 锡安山 和 耶路撒冷 成就他一切工作的时候，说：“我必惩罚 亚述 王自大的心和他高傲尊贵的眼目。”
ISA|10|13|因为他说： “我所成就的事是靠我手的能力 和我的智慧， 因为我本有聪明。 我挪移列国的地界， 抢夺他们所积蓄的财宝， 并且像勇士，使坐宝座的降为卑。
ISA|10|14|我的手夺取列国的财宝， 好像人夺取鸟窝； 我得了全地， 好像人拾起被弃的鸟蛋； 没有振动翅膀的， 没有张嘴的，也没有鸣叫的。”
ISA|10|15|斧岂可向用斧砍伐的自夸呢？ 锯岂可向拉锯的自大呢？ 这好比棍挥动那举棍的， 好比杖举起那不是木头的人。
ISA|10|16|因此，主－万军之耶和华 必使 亚述 王的壮士变为瘦弱， 在他的荣华之下必有火点燃， 如同火在燃烧一般。
ISA|10|17|以色列 的光必变成火， 它的圣者必成为火焰； 一日之间，将 亚述 王的荆棘和蒺藜焚烧净尽，
ISA|10|18|又毁灭树林和田园的荣华， 连魂带体，好像病重的人消逝 一样。
ISA|10|19|他林中只剩下稀少的树木， 连孩童也能写其数目。
ISA|10|20|到那日， 以色列 所剩下的和 雅各 家所逃脱的，必不再倚靠那击打他们的，却要诚心仰赖耶和华－ 以色列 的圣者。
ISA|10|21|所剩下的，就是 雅各 家的余民，必归回全能的上帝。
ISA|10|22|以色列 啊，你的百姓虽多如海沙，惟有剩下的归回。灭绝之事已成定局，公义必如水涨溢。
ISA|10|23|因为万军之主耶和华在全地必成就所定的灭绝之事。
ISA|10|24|所以，万军之主耶和华如此说：“住 锡安 我的百姓啊， 亚述 王虽然用棍击打你，又如 埃及 举杖攻击你，你不要怕他。
ISA|10|25|因为还有一点点时候，我向你们发的愤怒就要结束，我的怒气要使他们灭亡。
ISA|10|26|万军之耶和华要举起鞭子来攻击他，好像在 俄立 磐石那里击打 米甸 人一样。他的杖向海伸出，他必把杖举起，如在 埃及 一般。
ISA|10|27|到那日， 亚述 王的重担必离开你的肩头，他的轭必离开你的颈项；那轭必因肥壮而撑断 。”
ISA|10|28|亚述 王来到 亚叶 ， 经过 米矶仑 ， 在 密抹 安放辎重。
ISA|10|29|他们过了隘口， 要在 迦巴 住宿。 拉玛 战兢， 扫罗 的 基比亚 逃命。
ISA|10|30|迦琳 哪，要高声呼喊！ 注意听， 莱煞 啊！ 困苦的 亚拿突 啊 ！
ISA|10|31|玛得米那 躲避， 基柄 的居民逃遁。
ISA|10|32|当那日， 亚述 王要在 挪伯 停留， 挥手攻击 锡安 的山， 就是 耶路撒冷 的山。
ISA|10|33|看哪，主－万军之耶和华 以猛撞削断树枝； 巨木必被砍下， 高大的树必降为低。
ISA|10|34|稠密的树林，他要用铁器砍下， 黎巴嫩 必被大能者伐倒 。
ISA|11|1|从 耶西 的残干必长出嫩枝， 他的根所抽的枝子必结果实。
ISA|11|2|耶和华的灵必住在他身上， 就是智慧和聪明的灵， 谋略和能力的灵， 知识和敬畏耶和华的灵。
ISA|11|3|他必以敬畏耶和华为乐； 行审判不凭眼见， 断是非也不凭耳闻；
ISA|11|4|却要以公义审判贫寒人， 以正直判断地上的困苦人， 以口中的棍击打全地， 以嘴里的气杀戮恶人。
ISA|11|5|公义必当他的腰带， 信实必作他胁下的带子。
ISA|11|6|野狼必与小绵羊同住， 豹子与小山羊同卧； 少壮狮子、牛犊和肥畜同群 ； 孩童要牵引它们。
ISA|11|7|牛必与熊同食， 牛犊与小熊同卧； 狮子与牛一样吃草。
ISA|11|8|吃奶的婴孩在虺蛇的洞口玩耍， 断奶的幼儿必按手在毒蛇的穴上。
ISA|11|9|在我圣山各处， 它们都不伤人，不害物； 因为认识耶和华的知识要遍满全地， 好像水充满海洋一般。
ISA|11|10|到那日， 耶西 的根立作万民的大旗；列国的人必寻求他，他安歇之所大有荣耀。
ISA|11|11|当那日，主必再度伸手救回自己百姓中所剩余的，就是在 亚述 、 埃及 、 巴特罗 、 古实 、 以拦 、 示拿 、 哈马 ，并众海岛所剩下的。
ISA|11|12|他要向列国竖立大旗， 召集 以色列 被赶散的人， 又从地极四方聚集分散的 犹大 人。
ISA|11|13|以法莲 的嫉妒必消散， 苦待 犹大 的也被剪除； 以法莲 必不嫉妒 犹大 ， 犹大 也不苦待 以法莲 。
ISA|11|14|他们要飞向西方， 扑在 非利士 人的肩头上， 他们要一同掳掠东方人， 他们的手伸到 以东 和 摩押 ； 亚扪 人也必顺服他们。
ISA|11|15|耶和华必使 埃及 的海湾全然毁坏 ， 他举手在 大河 之上刮起了暴热的风， 击打它，使它分成七条溪流， 人穿鞋便可渡过。
ISA|11|16|必有一条大道， 为百姓中从 亚述 逃脱生还的余民而开， 如当日为 以色列 从 埃及 上来一样。
ISA|12|1|在那日，你要说： “耶和华啊，我要称谢你！ 因为你虽然向我发怒， 你的怒气却已转消； 你又安慰了我。
ISA|12|2|“看哪！上帝是我的拯救； 我要倚靠他，并不惧怕。 因为主耶和华是我的力量， 是我的诗歌， 他也成了我的拯救。”
ISA|12|3|你们必从救恩的泉源欢然取水。
ISA|12|4|在那日，你们要说： “当称谢耶和华，求告他的名； 在万民中传扬他的作为， 宣告他的名已被尊崇。
ISA|12|5|“你们要向耶和华唱歌， 因他所做的十分宏伟； 但愿这事遍传全地。
ISA|12|6|锡安 的居民哪，当扬声欢呼， 因为在你们当中的 以色列 圣者最为伟大。”
ISA|13|1|亚摩斯 的儿子 以赛亚 所见，有关 巴比伦 的默示。
ISA|13|2|你们要在荒凉的山上竖立大旗， 向他们扬声， 挥手招呼他们进入贵族之门。
ISA|13|3|我吩咐我所分别为圣的人， 召唤我的勇士， 就是我那狂喜高傲的人， 为要执行我的怒气。
ISA|13|4|听啊，山间有喧闹的声音， 好像有许多百姓聚集， 听啊，多国之民聚集闹哄的声音； 这是万军之耶和华召集作战的军队。
ISA|13|5|他们从远方来， 从天边来， 耶和华和他恼恨的兵器 要毁灭全地。
ISA|13|6|你们要哀号， 因为耶和华的日子临近了！ 这日来到，好像毁灭从全能者来到。
ISA|13|7|因此，人的手都变软弱， 人的心都必惶惶。
ISA|13|8|他们必惊恐， 悲痛和愁苦将他们抓住。 他们阵痛，好像临产的妇人一样， 彼此惊奇对看，脸如火焰。
ISA|13|9|看哪！耶和华的日子临到， 必有残忍、愤恨、烈怒， 使这地荒芜， 除灭其中的罪人。
ISA|13|10|天上的星宿都不发光， 太阳一升起就变黑暗， 月亮也不放光。
ISA|13|11|我必因邪恶惩罚世界， 因罪孽惩罚恶人， 我要止息骄傲人的狂妄， 制伏残暴者的傲慢。
ISA|13|12|我要使人比纯金更少， 比 俄斐 的赤金还少。
ISA|13|13|我，万军之耶和华狂怒，就是发烈怒的日子， 要令天震动， 地必摇撼，离其本位。
ISA|13|14|人如被追赶的羚羊， 像无人聚集的羊群， 各自归回本族， 逃到本地。
ISA|13|15|凡被追上的必被刺死， 凡被捉拿的必倒在刀下。
ISA|13|16|他们的婴孩必在他们眼前被摔死， 他们的房屋被抢劫， 他们的妻子被污辱。
ISA|13|17|看哪，我必激起 玛代 人攻击他们， 玛代 人并不看重银子， 也不喜爱金子。
ISA|13|18|他们必用弓击溃青年， 不怜悯妇人所生的； 眼也不顾惜孩子。
ISA|13|19|巴比伦 为列国的荣耀， 为 迦勒底 人所夸耀的华美， 必像上帝所倾覆的 所多玛 、 蛾摩拉 一样；
ISA|13|20|国中必永无人烟， 世世代代无人居住； 阿拉伯 人不在那里支搭帐棚， 牧羊的人也不使羊群躺卧在那里。
ISA|13|21|旷野的走兽躺卧在那里， 咆哮的动物挤满栖身之所； 鸵鸟住在那里， 山羊鬼魔也在那里跳舞。
ISA|13|22|土狼必在它的宫殿 呼号， 野狗在华美的殿里吼叫。 巴比伦 的时辰临近了， 它的日子必不长久。
ISA|14|1|耶和华要怜悯 雅各 ，再度拣选 以色列 ，将他们安顿在本地。寄居的必与他们联合，加入 雅各 家。
ISA|14|2|外邦人要将他们带回本地。 以色列 家必在耶和华的地上得外邦人为仆婢，也要掳掠先前掳掠他们的，辖制先前欺压他们的。
ISA|14|3|当耶和华使你得享安息，脱离愁苦、烦恼，和被迫做苦工的日子，
ISA|14|4|你必唱这诗歌嘲讽 巴比伦 王说： “欺压人的竟然灭亡！ 他的凶暴 竟然止息！
ISA|14|5|耶和华折断恶人的杖， 打断统治者的权杖；
ISA|14|6|他们在愤怒中连连攻击万民， 在怒气中辖制列国， 逼迫他们，毫不留情。
ISA|14|7|现在全地得安息，享平静， 人都出声欢呼。
ISA|14|8|松树和 黎巴嫩 的香柏树 都因你欢乐： 自从你仆倒， 再也无人上来砍伐我们。
ISA|14|9|下面的阴间因你震动， 迎接你的到来； 在世曾为领袖的阴魂为你惊动， 那曾为列国君王的，都从宝座起立。
ISA|14|10|他们都要发言，对你说： ‘你也变为软弱，像我们一样吗？ 你也成了我们的样子吗？’
ISA|14|11|你的威严和琴瑟的声音都下到阴间。 你下面铺的是虫，上面盖的是蛆。
ISA|14|12|“明亮之星，早晨之子啊， 你竟然从天坠落！ 你这攻败列国的，竟然被砍倒在地上！
ISA|14|13|你心里曾说： ‘我要升到天上， 我要高举我的宝座在上帝的众星之上， 我要坐在会众聚集的山上，在极北的地方。
ISA|14|14|我要升到高云之上， 我要与至高者同等。’
ISA|14|15|然而，你必坠落阴间， 到地府极深之处。
ISA|14|16|凡看见你的都要定睛望你， 留意看你，说： ‘就是这个人吗？ 他使大地颤抖， 使列国震动，
ISA|14|17|使世界如同荒野， 使城镇倾覆； 是他，不释放被掳的人归家。’
ISA|14|18|列国的君王各自在自己的坟墓中， 在尊荣里长眠。
ISA|14|19|惟独你被抛弃在你的坟墓之外， 有如被厌恶的枝子 ， 被许多用刀刺透杀死的人覆盖着， 一同坠落地府的石头那里， 像被践踏的尸首。
ISA|14|20|你不得与君王同葬， 因为你毁坏你的国，杀戮你的民。 “恶人的后裔永不留名。
ISA|14|21|为了祖先的罪孽， 要预备他子孙的屠宰场， 免得他们兴起，夺得全地， 使城市遍满地面。”
ISA|14|22|万军之耶和华说： “我必起来攻击他们， 将 巴比伦 的名号和剩余的人， 连子带孙一并剪除； 这是耶和华说的。
ISA|14|23|“我必使 巴比伦 为豪猪占据， 成为泥沼之地； 我要用灭命的扫帚扫净它； 这是万军之耶和华说的。”
ISA|14|24|万军之耶和华起誓说： “我怎样思想，必照样成就； 我怎样定意，必照样坚立，
ISA|14|25|要在我的地上击破 亚述 ， 在我的山上将它践踏。 它的轭必离开受压制的人， 它的重担必离开他们的肩头。”
ISA|14|26|这是向全地所定的旨意， 向万国所伸出的手。
ISA|14|27|万军之耶和华既然定意，谁能阻挠呢？ 他的手已经伸出，谁能使它缩回呢？
ISA|14|28|亚哈斯 王崩的那年，有默示如下：
ISA|14|29|“全 非利士 啊， 不要因击打你的杖折断就喜乐。 因为蛇必生出毒蛇， 它所生的是会飞的火蛇。
ISA|14|30|贫寒人的长子必有得吃； 贫穷人必安然躺卧。 我必以饥荒灭绝你的根， 它 必杀尽你所剩余的人。
ISA|14|31|门哪，哀号吧！ 城啊，呼喊吧！ 全 非利士 都熔化了！ 因为有烟从北方而来， 在它的行伍中没有掉队的。”
ISA|14|32|当如何回答外邦的使者呢？ “耶和华建立了 锡安 ， 在其中他困苦的百姓必有倚靠。”
ISA|15|1|论 摩押 的默示。 一夜之间， 摩押 的 亚珥 变为荒废， 归于无有； 一夜之间， 摩押 的 基珥 变为荒废， 归于无有。
ISA|15|2|摩押 上到神庙和 底本 的丘坛去哭泣； 它因 尼波 和 米底巴 哀号， 各人头上光秃，胡须剃净。
ISA|15|3|他们在街市上腰束麻布， 都在房顶和广场上哀号， 泪流不停。
ISA|15|4|希实本 和 以利亚利 呼喊， 他们的声音达到 雅杂 ， 所以 摩押 的士兵高声喊叫， 他们的心战兢。
ISA|15|5|我的心 为 摩押 哀号； 它的难民逃到 琐珥 ， 逃到 伊基拉．施利施亚 。 他们上 鲁希坡 ，随走随哭， 在 何罗念 的路上，因毁灭发出哀声。
ISA|15|6|宁林 的水干涸， 青草枯干，嫩草死光， 青绿之物，一无所有。
ISA|15|7|因此， 摩押 人所得的财物和积蓄 都要运过 柳树河 。
ISA|15|8|哀声遍传 摩押 四境， 哀号的声音达到 以基莲 ， 哀号的声音远及 比珥．以琳 。
ISA|15|9|底们 的水充满了血， 然而我还要加添 底们 的灾难， 让狮子追上 摩押 的难民 和那地 剩余的人。
ISA|16|1|你们当将 羔羊奉送给那地的掌权者， 从 西拉 往旷野，送到 锡安 的山。
ISA|16|2|摩押 的居民 来到 亚嫩 渡口， 如逃遁的飞鸟，被赶离鸟巢 。
ISA|16|3|求你赐谋略，行公平， 使你的影子在正午如黑夜， 掩护逃亡的人，不泄露逃难者的行踪。
ISA|16|4|愿我 摩押 逃亡的人 寄居在你那里， 你作他们的避难所，躲避灭命者的面。 勒索的人消失， 毁灭的事止息， 欺压者从国中除灭，
ISA|16|5|在 大卫 帐幕中必有宝座因慈爱坚立， 必有一位君王凭信实坐在其上， 施行审判，寻求公平，迅速行公义。
ISA|16|6|我们听闻 摩押 的骄傲， 极其骄傲； 它狂妄、骄傲、自大， 它夸大的言词都是空的。
ISA|16|7|因此， 摩押 人必为 摩押 哀号， 人人都要哀号。 你们要为 吉珥．哈列设 的葡萄饼哀叹， 极其忧伤。
ISA|16|8|因为 希实本 的田地 和 西比玛 的葡萄树都衰残了， 列国的君主折断它的枝干， 这枝子曾长到 雅谢 ，延伸到旷野， 嫩枝向外伸出，直伸过海；
ISA|16|9|所以，我要为 西比玛 的葡萄树哀哭， 像 雅谢 人一样哀哭。 希实本 、 以利亚利 啊， 我要以眼泪浇灌你， 你因夏天果子和收割的庄稼， 欢呼声已经止息了。
ISA|16|10|田园中不再有欢喜快乐， 葡萄园里必无人歌唱，无人欢呼， 在压酒池中踹酒的不再踹酒了， 我使欢呼的声音止息了 。
ISA|16|11|因此，我的心肠为 摩押 哀鸣如琴， 我的内心为 吉珥．哈列设 哀哭。
ISA|16|12|当 摩押 人出现在丘坛，筋疲力尽时，虽然到自己的圣所祈祷，却仍无济于事。
ISA|16|13|这是耶和华曾论到 摩押 的话。
ISA|16|14|但现在，耶和华说：“三年之内，按照雇工年数的算法， 摩押 的荣华必变为羞辱，人口虽曾众多，剩余的又少又弱。”
ISA|17|1|论 大马士革 的默示。 看哪， 大马士革 不再为城市， 变为废墟。
ISA|17|2|亚罗珥 的城镇被撇弃 ， 将成为牧羊之处， 羊群在那里躺卧， 无人使它们惊吓。
ISA|17|3|以法莲 不再有堡垒， 大马士革 失去其王国， 亚兰 的百姓所剩无几， 如 以色列 人的荣美消失一般； 这是万军之耶和华说的。
ISA|17|4|到那日， 雅各 的荣美必失色， 它肥胖的身躯渐渐消瘦；
ISA|17|5|像人收割成熟的禾稼， 用手臂割取麦穗， 又像人在 利乏音谷 拾取穗子；
ISA|17|6|其间所剩不多，好像人打橄榄树， 在最高的树梢上只剩两、三颗橄榄， 在多结果子的旁枝上只剩四、五颗； 这是耶和华－ 以色列 的上帝说的。
ISA|17|7|当那日，人必仰望造他们的主，眼目看着 以色列 的圣者。
ISA|17|8|他们必不仰望自己手所筑的祭坛，也不理会自己指头所造的 亚舍拉 和香坛。
ISA|17|9|当那日，他们坚固的城必因 以色列 人的缘故，如同树林中和山顶上所撇弃的地方 。这样，地就荒芜了。
ISA|17|10|因你忘记拯救你的上帝， 忘记那保护你的磐石； 所以，你虽栽上佳美的树苗， 插上别样的枝子，
ISA|17|11|栽种的日子，你使它生长， 栽种的早晨，你使它开花， 但在愁苦、极其伤痛的日子， 所收割的都归无有。
ISA|17|12|唉！万民闹哄，好像海浪澎湃， 列邦喧闹，如同洪水滔滔，
ISA|17|13|列邦喧闹，如同大水滔滔； 但上帝一斥责，他们就远远躲避， 他们被追赶，如同山上风前的糠秕， 又如暴风前的碎秸；
ISA|17|14|看哪，晚上有惊吓，未到早晨它就消失无踪。 这是掳掠我们之人的厄运，是抢夺我们之人的报应。
ISA|18|1|祸哉！ 古实河 的那一边、翅膀刷刷作响之地，
ISA|18|2|差遣使者在水面上， 坐蒲草船过海。 你们这些疾行的使者， 要到高大光滑的民那里去； 那民远近都畏惧， 是强大好征服的国， 土地有河流穿过。
ISA|18|3|世上所有的居民，住在地上的人哪， 山上大旗竖起时，你们要看， 号角吹响时，你们要听。
ISA|18|4|耶和华对我如此说： “我要安静，从我的居所观看， 如同日光下闪烁的热气， 又如收割时 露水蒸发的云雾。”
ISA|18|5|收割之前，花蕾先谢， 花成了将熟的葡萄； 他必用刀削去嫩枝， 砍掉蔓延的枝条，
ISA|18|6|一起丢给山间的鸷鸟和地上的野兽； 鸷鸟要在其上避暑， 地上一切的野兽都在那里过冬。
ISA|18|7|到那时，这高大光滑的民， 远近都畏惧的民、 强大好征服之国、 土地有河流穿过； 他们必被当作 礼物献给万军之耶和华， 献到 锡安山 － 万军之耶和华立他名的地方。
ISA|19|1|论 埃及 的默示。 看哪，耶和华乘驾快云， 临到 埃及 ； 埃及 的偶像在他面前战兢， 埃及 人的心在里面消溶。
ISA|19|2|我要激起 埃及 人攻击 埃及 人， 弟兄攻击弟兄， 邻舍攻击邻舍， 这城攻击那城， 这国攻击那国。
ISA|19|3|埃及 人的心神在里面耗尽， 我要破坏他们的计谋。 他们必求问偶像和念咒的， 求问招魂的与行巫术的人。
ISA|19|4|我要将 埃及 人交在严厉的主人手中， 残暴的君王必管辖他们； 这是主－万军之耶和华说的。
ISA|19|5|海水枯竭， 河流干涸，
ISA|19|6|江河发臭， 埃及 的河水必然减少而枯干。 芦苇和芦荻枯萎，
ISA|19|7|尼罗河 旁的植物 ，在 尼罗河 的沿岸， 并 尼罗河 旁所种的一切 全都枯焦，被风吹去，归于无有。
ISA|19|8|打鱼的哀哭， 所有在 尼罗河 钓鱼的都必悲伤， 在水上撒网的也都衰残。
ISA|19|9|以细致的麻编织的必羞愧， 织布的必变苍白 ；
ISA|19|10|织布的心情沮丧 ， 所有的佣工心都愁烦。
ISA|19|11|琐安 的官长极其愚昧， 法老智慧的谋士筹划愚谋； 你们怎敢对法老说： “我是智慧人的子孙， 是古代国王的后裔？”
ISA|19|12|你的智慧人在哪里？ 万军之耶和华向 埃及 所定的旨意， 他们既然知道，就让他们告诉你吧！
ISA|19|13|琐安 的官长愚昧， 挪弗 的官长受蒙蔽； 作 埃及 支派栋梁的， 带领 埃及 走错了路。
ISA|19|14|耶和华使歪曲的灵渗入 埃及 中间， 让他们使 埃及 一切所做的都出差错， 好像醉酒之人呕吐时东倒西歪一样。
ISA|19|15|在 埃及 ，无论是头是尾， 棕树枝与芦苇，所做的事都不得成就。
ISA|19|16|到那日， 埃及 必像妇人一样，因万军之耶和华挥手攻击而战兢惧怕。
ISA|19|17|犹大 地必使 埃及 惊恐，不论向谁提起，他都惧怕。这是因万军之耶和华向 埃及 所定的旨意。
ISA|19|18|当那日， 埃及 地必有五个城市的人说 迦南 的语言，又指着万军之耶和华起誓。有一城必称为“太阳城” 。
ISA|19|19|在那日，在 埃及 地将有献给耶和华的一座坛，边界上必有为耶和华立的一根柱子。
ISA|19|20|这都要在 埃及 地为万军之耶和华作记号和证据。 埃及 人因受欺压哀求耶和华，他就差遣一位救主作护卫者，拯救他们，
ISA|19|21|耶和华就被 埃及 所认识。在那日， 埃及 人要认识耶和华，献牲祭和素祭敬拜他，并向耶和华许愿还愿。
ISA|19|22|耶和华必击打 埃及 ，又击打又医治， 埃及 人就归向耶和华。他必应允他们的祷告，医治他们。
ISA|19|23|在那日，必有从 埃及 通往 亚述 的大道。 亚述 人要进入 埃及 ， 埃及 人也要进入 亚述 ； 埃及 人要与 亚述 人一同敬拜。
ISA|19|24|在那日， 以色列 将与 埃及 、 亚述 三国一起，使地上的人得福。
ISA|19|25|万军之耶和华必赐福给他们，说：“ 埃及 －我的百姓， 亚述 －我手的工作， 以色列 －我的产业，都有福了！”
ISA|20|1|亚述 元帅 受 亚述 王 撒珥根 派遣往 亚实突 的那年，他攻打 亚实突 ，将城攻取。
ISA|20|2|那时，耶和华吩咐 亚摩斯 的儿子 以赛亚 说：“你去解掉你腰间的麻布，脱下你脚上的鞋。” 以赛亚 就这样做，赤身赤脚行走。
ISA|20|3|耶和华说：“我仆人 以赛亚 怎样赤身赤脚行走三年，作为关于 埃及 和 古实 的预兆奇迹，
ISA|20|4|照样， 亚述 王必掳去 埃及 人，掠去 古实 人，无论老少，都赤身赤脚，露出下体，使 埃及 蒙羞。
ISA|20|5|以色列 人必惊惶羞愧，因为他们仰望 古实 ，以 埃及 为荣。
ISA|20|6|“那时，沿海一带的居民必说：‘看哪，我们素来所仰望的，就是为躲避 亚述 王所逃往 求救的，不过如此！我们怎能逃脱呢？’”
ISA|21|1|论海边旷野的默示。 它像 尼革夫 的旋风扫过， 从旷野，从可怕之地而来。
ISA|21|2|有凄惨的异象向我揭示： “诡诈的在行诡诈，毁灭的在行毁灭。 以拦 哪，前进吧！ 玛代 啊，围攻吧！ 我使它一切的叹息停止了。”
ISA|21|3|为此，我腰部满是疼痛， 痛苦将我抓住， 好像临产的妇人一样的痛。 我疼痛甚至不能听， 我惊惶甚至不能看 。
ISA|21|4|我心慌乱，惊恐威吓我。 我所渴望的黄昏，反成为我的恐惧。
ISA|21|5|有人摆设筵席， 铺上地毯，又吃又喝。 “官长啊，起来， 抹亮盾牌。”
ISA|21|6|主对我如此说： “你去设立守望者， 让他报告他所看见的。
ISA|21|7|他会看见一对一对骑着马的军队， 又看见驴队，骆驼队， 他要留心听，仔细地听。”
ISA|21|8|他如狮子般吼叫 ： “主啊，我白天常站在暸望楼， 彻夜立在我的暸望台。”
ISA|21|9|看哪，有一对一对骑着马的军队前来。 他就回应说：“ 巴比伦 倾倒了！倾倒了！ 他把 巴比伦 神明的一切雕刻偶像都打碎在地上了。”
ISA|21|10|我被打的禾稼，我禾场上的谷物啊， 我从万军之耶和华－ 以色列 的上帝那里所听见的，都告诉你们了。
ISA|21|11|论 度玛 的默示。 有人声从 西珥 呼喊： “守望的啊，夜里如何？ 守望的啊，夜里如何？”
ISA|21|12|守望者说： “早晨来到，黑夜将临。 你们若要问，问吧， 也可以回头再来。”
ISA|21|13|论 阿拉伯 的默示。 底但 的旅行商队啊， 你们在 阿拉伯 的树林中住宿。
ISA|21|14|提玛 地的居民哪， 提水来迎接口渴的人， 带饼来迎接难民。
ISA|21|15|他们躲避刀剑和出了鞘的刀， 躲避上了弦的弓与战争的重灾。
ISA|21|16|主对我这样说：“一年之内，按照雇工年数的算法， 基达 一切的繁华必归无有。
ISA|21|17|基达 人中强壮弓箭手剩下的数目甚为稀少，这是耶和华－ 以色列 的上帝说的。”
ISA|22|1|论异象谷的默示。 什么事使你们上去， 全都上到屋顶呢？
ISA|22|2|你这四处呐喊、大声喧哗的城、 欢乐的邑啊， 你被杀的并非被刀所杀， 也不是因打仗阵亡。
ISA|22|3|你所有的官长一同奔逃， 不用弓箭就被捆绑 ； 你们即使逃往远方， 也要被找到，一同被捆绑。
ISA|22|4|因此我说： “不要看我， 让我痛哭吧！ 不要因我百姓 的毁灭竭力安慰我。”
ISA|22|5|因为这是万军之主耶和华使异象谷 混乱、践踏、烦扰的日子； 城墙被攻破， 哀声达到山上。
ISA|22|6|以拦 提着箭袋， 有战车、士兵、骑兵； 吉珥 亮出盾牌，
ISA|22|7|你佳美的山谷遍布战车， 骑兵排列在城门前。
ISA|22|8|他除掉 犹大 的防御。 那时，你指望森林库里的兵器。
ISA|22|9|你们看见 大卫城 缺口很多，就汇集 下池 的水；
ISA|22|10|你们数点 耶路撒冷 的房屋，拆毁房屋，用以修补城墙，
ISA|22|11|又在两道城墙中间挖水池，用以盛旧池的水，却不仰望成就这事的主，也不顾念从古时定这事的主。
ISA|22|12|当那日，万军之主耶和华使人哭泣哀号， 头上光秃，身披麻布。
ISA|22|13|看哪，人却欢喜快乐， 宰牛杀羊，吃肉喝酒： “让我们吃吃喝喝吧！因为明天要死了。”
ISA|22|14|万军之耶和华开启我的耳朵： “这罪孽直到你们死，断不得赦免！” 这是万军之主耶和华说的。
ISA|22|15|万军之主耶和华如此说：“你到 舍伯那 宫廷总管那里去，说：
ISA|22|16|‘你在这里凭什么？你在这里靠谁？竟敢在这里为自己凿坟墓，在高处为自己凿坟墓，在岩石中为自己挖安身之所！
ISA|22|17|你这伟大的人，看哪，耶和华必将你用力抛出，将你紧紧缠裹。
ISA|22|18|他必将你卷成一团，好像抛球一样抛向宽阔之地。你这主人家的羞辱啊，你必死在那里，你引以为荣的战车也毁在那里。
ISA|22|19|我要革除你的官职，你必从原位被逐 。’
ISA|22|20|“到那日，我要召 希勒家 的儿子─我的仆人 以利亚敬 来，
ISA|22|21|将你的外袍给他穿上，将你的腰带给他系紧，将你的政权交在他手中。他必作 耶路撒冷 居民和 犹大 家的父。
ISA|22|22|我要将 大卫 家的钥匙放在他肩头上。他开了，无人能关；他关了，无人能开。
ISA|22|23|我要使他立稳，像钉子钉在坚固的地方；他必成为他父家荣耀的宝座。
ISA|22|24|他父家所有的荣耀，连儿女带子孙，有如杯碗、瓶罐的小器皿，都挂在他身上。
ISA|22|25|当那日，万军之耶和华说，钉在坚固处的钉子必挪移，被砍断落地，挂在上面的各样重担都被切断。这是耶和华说的。”
ISA|23|1|论 推罗 的默示。 哀号吧， 他施 的船只！ 因为 推罗 已成废墟，没有房屋存留， 他们从 基提 地来的时候，得到这个消息 。
ISA|23|2|沿海的居民， 西顿 的商家啊， 当静默无声。 你差人航海 ，
ISA|23|3|在大水之上， 西曷河 的粮食、 尼罗河 的庄稼是 推罗 的进项， 它就成为列国的商埠。
ISA|23|4|西顿 ，你这海洋中的堡垒啊，应当羞愧， 因为大海说 ： “我未经历产痛，也没有生产， 未曾养育男孩，也没有抚养女孩。”
ISA|23|5|推罗 的风声传到 埃及 时， 他们为这风声极其疼痛。
ISA|23|6|你们当渡到 他施 去， 哀号吧，沿海的居民！
ISA|23|7|这就是你们那古老欢乐的城市吗？ 它的脚曾带人到远方居住。
ISA|23|8|谁定意 推罗 有这样的遭遇呢？ 它本是赐冠冕的， 它的商家是王子， 生意人是世上尊贵的人。
ISA|23|9|这是万军之耶和华所定的， 为要贬抑一切荣耀的狂傲， 使地上一切尊贵的人被藐视。
ISA|23|10|他施 啊， 你要像 尼罗河 一样在你的地泛滥， 不再有腰带的束缚了。
ISA|23|11|耶和华已经向海伸手， 震动列国； 他出令对付 迦南 ， 要拆毁其中的堡垒。
ISA|23|12|他说：“受欺压的少女 西顿 哪， 你必不再欢乐。 起来！渡到 基提 去， 就是在那里也不得安歇。
ISA|23|13|看哪， 迦勒底 人之地，这国民如今已不复存在。 亚述 人使它 成为住旷野者的居所。他们建筑自己的了望楼，拆毁它的宫殿，使它成为荒凉。
ISA|23|14|哀号吧， 他施 的船只！ 因你们的堡垒已成废墟。
ISA|23|15|到那时， 推罗 必被忘记七十年，就是一位君王的年数。七十年后， 推罗 的景况必如妓女之歌：
ISA|23|16|“你这被遗忘的妓女啊， 带着琴周游城内， 弹得美妙，唱许多歌， 好让人记得你。”
ISA|23|17|七十年后，耶和华必巡视 推罗 ，使它再度获利 ，与地面上的世界各国贸易 。
ISA|23|18|它的收益和获利都要归耶和华为圣，不再私自屯积存留；因为它的收益必归给住在耶和华面前的人，使他们吃饱，穿华丽的衣服。
ISA|24|1|看哪，耶和华使地空虚，变为荒芜， 地面扭曲，居民四散。
ISA|24|2|那时，百姓如何，祭司也如何； 仆人如何，主人也如何； 婢女如何，主母也如何； 买主如何，卖主也如何； 放债的如何，借贷的也如何； 债主如何，欠债的也如何。
ISA|24|3|地必全然空虚，尽都荒芜， 因为这话是耶和华说的。
ISA|24|4|大地悲哀凋零， 世界败落衰残， 地上居高位的人也没落了。
ISA|24|5|地被其上的居民所污秽， 因为他们犯了律法， 废了律例，背了永约。
ISA|24|6|所以，诅咒吞灭大地， 住在其上的都有罪； 地上的居民被火焚烧， 剩下的人稀少。
ISA|24|7|新酒悲哀，葡萄树凋残， 心中欢乐的都叹息。
ISA|24|8|击鼓之乐停止， 狂欢者的喧哗止住， 弹琴之乐也停止了。
ISA|24|9|人不再饮酒唱歌， 喝烈酒的，必以为苦。
ISA|24|10|荒凉的城拆毁了， 各家关闭，无法进入。
ISA|24|11|有人在街上嚷着要酒喝， 一切的喜乐变为昏暗， 地上的欢乐全都消失。
ISA|24|12|城里尽是荒凉， 城门全都摧毁。
ISA|24|13|地上的万民正像打过的橄榄树， 又如葡萄酿酒以后再去摘取，所剩无几。
ISA|24|14|他们要高声欢呼， 从海那边扬声赞美耶和华的威严。
ISA|24|15|因此，你们要在日出之地荣耀耶和华， 在众海岛荣耀耶和华－ 以色列 上帝的名。
ISA|24|16|我们听见从地极有人歌唱： “荣耀归于公义的那一位！” 我却说：“我灭亡了！ 我灭亡了，我有祸了！ 诡诈的还在行诡诈， 诡诈的还在大行诡诈。”
ISA|24|17|地上的居民哪， 惊吓、陷阱、罗网都临到你；
ISA|24|18|躲过惊吓之声的坠入陷阱， 逃离陷阱的又被罗网缠住， 因为天上的窗户都打开， 地的根基也震动。
ISA|24|19|地必全然破坏，尽都崩裂， 剧烈震动。
ISA|24|20|地要摇摇晃晃，好像醉酒的人， 又如小屋子摇来摇去； 罪过重压其上， 它就塌陷，不能复起。
ISA|24|21|到那日，耶和华在天上必惩罚天上的军队， 在地上必惩罚地上的列王。
ISA|24|22|他们必被聚集， 像囚犯困在牢里， 他们被关在监狱， 多日之后便受惩罚。
ISA|24|23|那时，月亮要蒙羞，太阳要惭愧， 因为万军之耶和华必在 锡安山 ， 在 耶路撒冷 作王， 在他众长老面前彰显荣耀。
ISA|25|1|耶和华啊，你是我的上帝， 我要尊崇你，称颂你的名。 因为你以信实忠信 行远古所定奇妙的事。
ISA|25|2|你使城市变为废墟， 使坚固的城荒凉， 使外邦人的城堡不再为城， 永远不再重建。
ISA|25|3|所以，强大的民必尊敬你， 残暴之国的城必敬畏你。
ISA|25|4|因为你是贫寒人的保障， 贫穷人急难中的保障， 暴风雨之避难所， 炎热地之阴凉处。 当残暴者盛气凌人的时候， 如暴风直吹墙壁，
ISA|25|5|如干旱地的热气， 你要制止外邦人的喧嚷， 残暴者的歌要停止， 好像热气因云的阴影而消失。
ISA|25|6|在这山上，万军之耶和华必为万民摆设宴席，有肥甘与美酒，就是满有骨髓的肥甘与精酿的美酒。
ISA|25|7|在这山上，他必吞灭缠裹万民的面纱和那遮盖列国的遮蔽物。
ISA|25|8|他已吞灭死亡直到永远。主耶和华必擦干各人脸上的眼泪，在全地除去他百姓的羞辱；这是耶和华说的。
ISA|25|9|到那日，人必说：“看哪，这是我们的上帝，我们向来等候他，他必拯救我们。这是耶和华，我们向来等候他，我们必因他的救恩欢喜快乐。”
ISA|25|10|耶和华的手必按住这山， 摩押 人要被践踏在他底下，好像干草被践踏在粪池 里。
ISA|25|11|他们要在其中伸展双手，好像游泳的人伸手游泳。他们的手虽灵巧，耶和华却使他们的骄傲降为卑下。
ISA|25|12|他使你城墙上坚固的碉堡倾倒，夷为平地，化为尘土。
ISA|26|1|当那日，在 犹大 地，人必唱这歌： “我们有坚固的城， 耶和华赐救恩为城墙，为城郭。
ISA|26|2|你们要敞开城门， 使守信的公义之民得以进入。
ISA|26|3|坚心倚赖你的，你必保守他十分平安， 因为他倚靠你。
ISA|26|4|你们当倚靠耶和华，直到永远， 因为耶和华，耶和华是永远的磐石。
ISA|26|5|他使居住高处的与高处的城市一同降为卑下， 将城拆毁，夷为平地，化为尘土，
ISA|26|6|使它被脚践踏， 就是被困苦人和贫寒人的脚践踏。”
ISA|26|7|义人的道是正直的， 正直的主啊，你修平义人的路。
ISA|26|8|耶和华啊，我们在你行审判的路上等候你 ， 我们心里所渴慕的，就是你的名和你的称号 。
ISA|26|9|夜间，我的心渴想你， 我里面的灵切切寻求你。 因为你在地上行审判的时候， 世上的居民就学习公义。
ISA|26|10|恶人虽然领受恩惠， 仍未学到公义。 在正直之地，他行不义， 也不看耶和华的威严。
ISA|26|11|耶和华啊，你的手高举，他们不观看； 愿他们观看你为百姓发的热心而羞愧， 愿火吞灭你的敌人。
ISA|26|12|耶和华啊，你必赏赐我们平安， 因为我们所做的一切，都是你为我们成就的。
ISA|26|13|耶和华－我们的上帝啊， 在你以外曾有别的主管辖我们， 但我们惟独称扬你的名。
ISA|26|14|死去的不能再复活， 阴魂不能再兴起； 你惩罚他们，使他们毁灭， 他们的名号 就全然消灭。
ISA|26|15|耶和华啊，你增添国民， 你增添国民，得了荣耀， 又拓展国土的疆界。
ISA|26|16|耶和华啊，他们在急难中寻求你。 你的管教临到他们身上时， 他们倾吐低声的祷告。
ISA|26|17|妇人怀孕，临产疼痛， 在痛苦之中喊叫； 耶和华啊，我们在你面前也是如此。
ISA|26|18|我们曾怀孕，曾疼痛， 所生产的竟像风一样， 并未带给地上任何拯救； 世上也未曾有居民生下来 。
ISA|26|19|你的死人要复活， 我的尸首要起来。 睡在尘土里的啊，要醒起歌唱！ 你的甘露好像晨曦 的甘露， 地要交出阴魂。
ISA|26|20|我的百姓啊，要进入内室， 关上你的门，躲避片刻， 等到愤怒过去。
ISA|26|21|因为，看哪，耶和华从他的居所出来， 要惩罚地上居民的罪孽。 地必露出其中的血， 不再掩盖被杀的人。
ISA|27|1|到那日，耶和华必用他坚硬锐利的大刀惩罚 力威亚探 ，就是那爬得快的蛇，惩罚 力威亚探 ，就是那弯弯曲曲的蛇，并杀死海里的大鱼。
ISA|27|2|当那日，你们要唱这美好 葡萄园的歌：
ISA|27|3|“我－耶和华看守葡萄园，按时灌溉， 昼夜看守，免得有人损害。
ISA|27|4|我心中不存愤怒。 惟愿在战争中我有荆棘和蒺藜， 我就起步攻击他， 把他一同焚烧；
ISA|27|5|或者让他紧靠我，以我为避难所， 与我和好， 与我和好。”
ISA|27|6|将来 雅各 要扎根， 以色列 要发芽开花， 果实遍满地面。
ISA|27|7|耶和华击打 以色列 ， 岂像击打那些击打他们的人吗？ 以色列 被杀戮， 岂像其他人所遭遇的杀戮吗？
ISA|27|8|你驱赶他们，放逐他们， 与他们相争。 在刮东风的日子， 他以暴风赶逐他们。
ISA|27|9|所以， 雅各 的罪孽藉此得赦免， 除罪的效果尽在乎此； 他使祭坛的石头变为粉碎的石灰， 使 亚舍拉 和香坛不再立起。
ISA|27|10|因为坚固的城变为荒凉， 成了被撇弃的居所，像旷野一样； 牛犊在那里吃草， 在那里躺卧，吃尽其中的树枝。
ISA|27|11|它的枝条一枯干，就被折断， 妇女用以点火燃烧。 因为这百姓蒙昧无知， 所以，造他们的必不怜悯他们， 造成他们的也不施恩给他们。
ISA|27|12|到那日， 以色列 人哪，耶和华必像人打树拾果一般，从 大河 的支流，直到 埃及 的溪谷，将你们一一收集。
ISA|27|13|当那日，号角大响；在 亚述 地将亡的，与被赶散至 埃及 地的，都要前来，在 耶路撒冷 圣山上敬拜耶和华。
ISA|28|1|祸哉！ 以法莲 酒徒高傲的冠冕， 其荣美竟如花凋残； 他们在肥沃的山谷顶上， 被酒击败。
ISA|28|2|看哪，主有一位大能大力者， 如强烈的冰雹， 如毁灭的暴风雨， 如涨溢的洪水， 他必亲手将他们摔落在地。
ISA|28|3|以法莲 酒徒高傲的冠冕， 必被脚践踏；
ISA|28|4|那如凋残之花的荣美， 在肥沃的山谷顶上， 必如夏令前初熟的无花果， 让看见的人注意， 摘到手里，随即吞吃。
ISA|28|5|到那日，万军之耶和华 必成为他余民的荣冠华冕，
ISA|28|6|成为在位审判者的公平之灵， 和城门口制敌的力量。
ISA|28|7|这些人也因酒摇晃， 因烈酒东倒西歪。 祭司和先知因烈酒摇晃， 被酒所困， 因烈酒东倒西歪。 他们错解默示， 审判时不分是非。
ISA|28|8|筵席上都满了呕吐的污秽， 没有一处干净。
ISA|28|9|“他要将知识指教谁呢？ 要向谁阐明信息呢？ 是向那些刚断奶的， 离开母亲胸怀的吗？
ISA|28|10|因为他咕哝咕哝，咕哝咕哝， 唠唠叨叨，唠唠叨叨， 这里一点，那里一点。”
ISA|28|11|耶和华要藉嘲弄的嘴唇和外邦人的舌头， 向这百姓说话。
ISA|28|12|他曾对他们说： “这是安歇之所， 你们要使疲乏的人得安歇， 这是歇息之处。” 他们却不肯听。
ISA|28|13|耶和华的话对他们而言是 “咕哝咕哝，咕哝咕哝， 唠唠叨叨， 唠唠叨叨， 这里一点，那里一点”； 以致他们往前行， 却后仰跌倒，甚至跌伤， 落入陷阱，被抓住了。
ISA|28|14|因此，你们这些傲慢的人， 就是管辖住 耶路撒冷 这百姓的， 要听耶和华的话。
ISA|28|15|你们曾说： “我们已与死亡立约， 与阴间结盟， 不可挡的鞭子挥过时， 必不临到我们； 因我们以谎言为避难所， 靠虚假来藏身”；
ISA|28|16|所以，主耶和华如此说： “看哪，我在 锡安 放一块石头作为根基， 是衡量的石头， 是宝贵的房角石，稳固的根基； 信靠他的人必不致惊恐。
ISA|28|17|我以公平为准绳， 以公义为铅垂线； 冰雹必冲去谎言的避难所， 大水必漫过藏身之处。
ISA|28|18|你们与死亡所立的约必废除， 与阴间所结的盟不得坚立； 不可挡的鞭子挥过时， 你们必被践踏。
ISA|28|19|每逢它挥来，必将你们掳去； 每早晨它必挥过， 白昼黑夜都是如此。 明白这信息的都必惊恐。”
ISA|28|20|床榻短，人不能伸展； 被子窄，人无从裹身。
ISA|28|21|耶和华必兴起，像在 毗拉心山 ， 他必发怒，如在 基遍谷 ； 为要做成他的工，就是非常的工， 成就他的事，就是奇异的事。
ISA|28|22|现在你们不可傲慢， 免得捆绑你们的绳索更结实， 因为我从万军之主耶和华那里听见， 在全地施行灭绝的事已定。
ISA|28|23|你们当侧耳听我的声音， 留心听我的言语。
ISA|28|24|那为撒种而耕地的 会不停地耕地，松土，耙地吗？
ISA|28|25|他铲平了地面， 岂不就种小茴香， 播种大茴香， 按行列种小麦， 在定处种大麦， 在田边种粗麦吗？
ISA|28|26|他的上帝教导他， 指导他合宜的方法。
ISA|28|27|原来打小茴香，不用尖利的器具， 轧大茴香，也不是用车轮； 却要用杖打小茴香， 用棍打大茴香。
ISA|28|28|谷要打， 但不能持续地捣， 用车轮和马轧， 却不轧碎它。
ISA|28|29|这也是出于万军之耶和华， 他的谋略奇妙， 他的智慧广大。
ISA|29|1|祸哉！ 亚利伊勒 ， 亚利伊勒 ， 大卫 安营的城， 任凭你年复一年， 节期照常循环，
ISA|29|2|我却要使 亚利伊勒 遭难； 它必悲伤哀号， 它对我是 亚利伊勒 。
ISA|29|3|我必四围安营攻击你， 筑台围困你， 堆垒攻击你。
ISA|29|4|你必败落，从地里说话， 你的言语细微出于尘埃。 你的声音必像那招魂者的声音出于地， 你的言语呢喃出于尘埃。
ISA|29|5|你那成群的陌生人 要像细尘， 暴民要像吹起的糠秕； 这事必顷刻之间忽然临到。
ISA|29|6|万军之耶和华必使雷轰、地震、巨响、旋风、暴风， 并吞灭的火焰临到它。
ISA|29|7|那时，攻击 亚利伊勒 列国的军队， 与一切攻击 亚利伊勒 和它城堡， 并带给它患难的， 必如梦，如夜间的异象；
ISA|29|8|又像饥饿的人在梦中吃饭， 醒了仍觉饥肠辘辘； 或像口渴的人在梦中喝水， 醒了仍觉发昏，心里想喝。 攻击 锡安山 列国的军队也必如此。
ISA|29|9|你们等候惊奇吧！ 你们沉迷宴乐吧！ 他们醉了，却非因酒； 东倒西歪，却非因烈酒。
ISA|29|10|因为耶和华将沉睡的灵浇灌你们， 遮住你们的眼， 眼就是先知， 覆盖你们的头， 头就是先见。
ISA|29|11|所有的默示，在你们看来都如封住的书卷，人将这书卷交给识字的人，说：“请念吧！”他说：“我不能念，因为它封住了。”
ISA|29|12|又将这书卷交给不识字的人，说：“请念吧！”他说：“我不识字。”
ISA|29|13|主说：“因这百姓以口亲近我， 用嘴唇尊敬我， 心却远离我； 他们敬畏我， 不过是领受前人的命令。
ISA|29|14|所以，看哪，我要在这百姓中行奇妙的事， 就是奇妙又奇妙的事。 他们智慧人的智慧必然消灭， 聪明人的聪明必然消失。”
ISA|29|15|祸哉！那些向耶和华深藏谋略的， 他们在暗中行事，说： “有谁看见我们呢？ 谁会注意我们呢？”
ISA|29|16|你们把事情颠倒了， 岂可看陶匠如陶土呢？ 受造物岂可论创造者说， “他并没有造我”？ 制成物岂可论制作者说， “他根本不懂”？
ISA|29|17|黎巴嫩 变为田园， 田园看似森林， 不是只需要一些时间吗？
ISA|29|18|那时，聋子必听见这书上的话； 盲人的眼必从迷蒙黑暗中看见。
ISA|29|19|困苦的人必因耶和华增添欢喜， 人间贫穷的必因 以色列 的圣者快乐。
ISA|29|20|因为残暴的人归于无有， 傲慢的人已经灭绝， 一切存心作恶的都被剪除。
ISA|29|21|他们凭一句话定一个人有罪， 为在城门口断是非的设下罗网， 又用虚无的事屈枉义人。
ISA|29|22|所以，救赎 亚伯拉罕 的耶和华 论到 雅各 家时如此说： “ 雅各 必不再羞愧， 面容也不再变色。
ISA|29|23|当他的儿女看见 我的手在他们当中所成就的事情 ， 他们就必尊我的名为圣， 尊 雅各 的圣者为圣， 他们必敬畏 以色列 的上帝。
ISA|29|24|心中迷糊的必明白， 发怨言的必领受训诲。”
ISA|30|1|耶和华说： “祸哉！这悖逆的儿女。 他们同谋，却不出于我， 结盟，却不出于我的灵， 以致罪上加罪。
ISA|30|2|他们没有寻求我的指示，就起身下 埃及 去， 要倚靠法老的庇护坚固自己， 并投在 埃及 的荫下。
ISA|30|3|但法老的庇护反成为你们的羞辱； 你们投在 埃及 荫下，反使你们惭愧。
ISA|30|4|他们的领袖已在 琐安 ， 他们的使臣到了 哈内斯 。
ISA|30|5|他们必因那无益于他们的民蒙羞； 那民并非帮助，也非有益， 只带来羞耻和凌辱。”
ISA|30|6|论 尼革夫 牲畜的默示。 他们将财物驮在驴背上， 将宝物驮在骆驼的背脊， 经过艰难困苦之地， 就是母狮、公狮、毒蛇、飞蛇之地， 往那无益于他们的民那里去。
ISA|30|7|埃及 的帮助是徒然的， 因此，我称它为“毫不中用的 拉哈伯 ” 。
ISA|30|8|现在你要去， 在他们面前将这话刻在版上， 写在书上， 以便流传后世，直到永永远远 。
ISA|30|9|因为他们是悖逆的百姓、说谎的儿女， 是不肯听从耶和华训诲的儿女。
ISA|30|10|他们对先见说：“不要再看了”； 对先知说：“不要向我们预言正直的事； 要对我们说好听的话， 预言虚幻的事。
ISA|30|11|要离开这道，偏离这路， 不要在我们面前再提说 以色列 的圣者。”
ISA|30|12|所以， 以色列 的圣者如此说： “因你们藐视这话， 倚赖欺压和诡诈，以此为可靠，
ISA|30|13|因此，这罪孽在你们身上， 好像高墙里有凸起的裂缝， 顷刻之间忽然坍下来了；
ISA|30|14|它被砸碎，好像把陶匠的瓦器摔碎， 毫不顾惜， 甚至在碎块中找不到一片 可用以从炉内取火，或从池中舀水。
ISA|30|15|主耶和华－ 以色列 的圣者如此说： “你们得救在乎归回安息， 得力在乎平静安稳。” 你们却是不肯，
ISA|30|16|你们说：“不然，我们要骑马奔走”， 所以你们必然奔走。 你们又说：“我们要骑快马”， 所以追赶你们的，也必飞快。
ISA|30|17|一人叱喝，令千人逃跑， 五人叱喝，你们都逃跑； 以致剩下的如山顶的旗杆， 如山冈上的大旗。
ISA|30|18|耶和华必然等候，要施恩给你们； 必然兴起，好怜悯你们。 因为耶和华是公平的上帝； 凡等候他的都是有福的！
ISA|30|19|住在 锡安 、居于 耶路撒冷 的百姓啊，你必不再哭泣。主必因你哀求的声音施恩给你，他听见的时候就必应允你。
ISA|30|20|主虽然以艰难给你当饼，以困苦给你当水，你的教师却不再隐藏，你的眼睛必看见你的教师。
ISA|30|21|你或向左或向右，必听见后边有声音说：“这是正路，要行在其间。”
ISA|30|22|你要玷污那雕刻偶像所包的银子和铸造偶像所镀的金子。你要抛弃它们，如抛弃污秽之物；对偶像说：“去吧！”
ISA|30|23|你撒种在地里，主必降雨在其上，使地所出的粮食肥美丰盛。那时，你的牲畜必在辽阔的草场吃草。
ISA|30|24|耕地的牛和驴必吃加盐的饲料，是用铲子和杈子扬净的。
ISA|30|25|在大行杀戮的日子，城楼倒塌的时候，高山峻岭必有川河涌流。
ISA|30|26|当耶和华包扎他百姓的伤口，医治他所击打伤痕的日子，月光必像日光，日光必加七倍，像七日的光一样。
ISA|30|27|看哪，耶和华的名从远方来， 他的怒气烧起，浓烟上腾。 他的嘴唇满有愤恨， 他的舌头像吞灭的火。
ISA|30|28|他的气息如涨溢的河水，直涨到颈项， 要用毁灭的筛网筛净列国， 并在众民口中安放导错方向的嚼环。
ISA|30|29|你们必唱歌，像守圣节的夜间一样；并且心中喜乐，像人吹笛，来到耶和华的山，到 以色列 的磐石那里。
ISA|30|30|耶和华必使人听见他威严的声音，又以极大的愤怒、吞灭的火焰、雷雨、暴风和像石块的冰雹，使人看见他降罚的膀臂。
ISA|30|31|亚述 必因耶和华的声音惊惶，耶和华必用杖击打它。
ISA|30|32|耶和华必将定规要打 的杖加在它身上；每打一下，都必配合击鼓弹琴的节奏。打仗时，耶和华必振臂与它交战。
ISA|30|33|原来 陀斐特 早已预备好了，是为君王预备的；又深又宽，堆满了火和木柴；耶和华的气息犹如一股硫磺使它燃起。
ISA|31|1|祸哉！那些下 埃及 求帮助的， 他们仰赖马匹，倚靠甚多的战车， 并倚靠强壮的骑兵， 却不仰望 以色列 的圣者， 也不求问耶和华。
ISA|31|2|其实，耶和华有智慧， 他降灾祸， 并不撤回自己的话， 却要兴起攻击作恶之家， 攻击那帮助人作恶的。
ISA|31|3|埃及 人不过是人，并非上帝， 他们的马不过是血肉，并不是灵。 耶和华一伸手， 那帮助人的必绊跌，受帮助的也必跌倒， 都一同灭亡。
ISA|31|4|耶和华对我如此说， 狮子和少壮狮子为猎物而咆哮， 许多牧人被召来攻击它， 它总不因他们的声音惊惶， 也不因他们的喧嚷退缩； 万军之耶和华也必如此 降临在 锡安 的大小山冈上争战。
ISA|31|5|雀鸟盘旋护卫， 万军之耶和华也必照样保护 耶路撒冷 ； 他必保护拯救， 必逾越而搭救。
ISA|31|6|以色列 人哪，要归向你们严重悖逆的那一位！
ISA|31|7|到那日，你们各人要抛弃亲手所造、陷自己于罪中的金偶像和银偶像。
ISA|31|8|亚述 必倒在刀下，并非人的刀； 有刀要将它吞灭，并非人的刀。 它要逃避这刀， 它的年轻人必做苦工。
ISA|31|9|它的磐石必因惊吓而消失， 它的领袖必因大旗惊惶； 这是那有火在 锡安 、 有炉在 耶路撒冷 的耶和华说的。
ISA|32|1|看哪，必有一位君王凭公义执政， 必有王子藉公平掌权。
ISA|32|2|必有一人如避风港， 如暴风雨的藏身处； 如干旱地的溪流， 又如干燥地巨石的阴影。
ISA|32|3|看的人眼睛不再昏花， 听的人耳朵必留心听。
ISA|32|4|性急的人懂得分辨， 口吃的人说话流畅。
ISA|32|5|愚顽人不再称为君子， 流氓不再称为绅士。
ISA|32|6|因为愚顽人必说愚妄的话， 他的心作恶 ， 行亵渎的事， 传播恶言攻击耶和华， 使饥饿的人仍然饥饿， 口渴的人无水可喝。
ISA|32|7|流氓的手段邪恶， 他图谋恶计， 用谎言毁灭困苦人； 贫穷人讲求公理时， 他也是如此行。
ISA|32|8|君子却图谋高尚的事， 他必因高尚的事站立得稳。
ISA|32|9|安逸的妇女啊，起来听我的声音！ 无虑的女子啊，侧耳听我的言语！
ISA|32|10|无虑的女子啊，再过一年，你们必颤栗， 因为无葡萄可摘， 也无果实可收。
ISA|32|11|安逸的妇女啊，要战兢； 无虑的女子啊，要颤栗， 要脱去衣服，赤着身体， 腰束麻布。
ISA|32|12|你们要为美好的田地 和多结果子的葡萄树捶胸哀哭。
ISA|32|13|刺草和荆棘要长在我百姓的田地上， 长在欢乐城中一切快乐家园上。
ISA|32|14|宫殿必被撇下， 繁华的城必被抛弃， 堡垒和了望楼永为洞穴， 成为野驴的乐土， 羊群的草场。
ISA|32|15|等到圣灵从高处浇灌我们， 旷野将变为田园， 田园看似森林。
ISA|32|16|公平要居住在旷野， 公义要安歇在田园。
ISA|32|17|公义的果实是平安， 公义的效果是平静和安稳，直到永远。
ISA|32|18|我的百姓要住在平安的居所， 安稳的住处，宁静的安歇之地。
ISA|32|19|虽有冰雹击倒树林， 城也夷为平地；
ISA|32|20|然而你们在水边撒种， 牧放牛驴的有福了！
ISA|33|1|祸哉！你这未遭毁灭而毁灭人的人， 人未以诡诈待你而你以诡诈待人的人！ 等你行完了毁灭， 自己必被毁灭； 你行完了诡诈， 人必以诡诈待你。
ISA|33|2|耶和华啊，求你施恩给我们， 我们等候你。 求你每早晨作我们的膀臂， 遭难时作我们的拯救。
ISA|33|3|轰然之声一发出，万民就奔逃； 你一兴起 ，列国就四散。
ISA|33|4|你们的掳物必被敛尽， 有如蚂蚱敛尽禾稼； 人为掳物奔走，宛如蝗虫蹦跳。
ISA|33|5|耶和华受尊崇，居高处， 使公平和公义充满 锡安 。
ISA|33|6|他是你这世代安定的力量， 丰盛的救恩、 智慧和知识； 敬畏耶和华是 锡安 的至宝。
ISA|33|7|看哪，他们的英雄在外面哀号 ， 求和的使臣在痛哭。
ISA|33|8|大路荒凉，行人止息； 盟约撕毁，见证 被弃， 人也不受尊重。
ISA|33|9|大地悲哀衰残， 黎巴嫩 羞愧且枯干， 沙仑 好像旷野， 巴珊 和 迦密 必凋残。
ISA|33|10|耶和华说： “现在我要兴起， 要高升， 要受尊崇。
ISA|33|11|你们怀的是糠秕，生的是碎秸； 你们的气息如火吞灭自己。
ISA|33|12|万民必像烧着的石灰， 又如斩断的荆棘，在火里燃烧。”
ISA|33|13|你们远方的人，当听我所做的事； 你们近处的人，当承认我的大能。
ISA|33|14|锡安 的罪人都惧怕， 战兢抓住不敬虔的人。 我们中间有谁能与吞噬的火同住？ 我们中间有谁能与不灭的火共存呢？
ISA|33|15|那行事公义、说话正直、 憎恶欺压所得之财、 摇手不受贿赂、 掩耳不听流血的计谋、 闭眼不看邪恶之事的，
ISA|33|16|这人必居高处， 他的保障是磐石的堡垒， 必有粮食赐给他， 饮水也不致断绝。
ISA|33|17|你必亲眼看见君王的荣美， 看见辽阔之地。
ISA|33|18|你的心必回想那些恐怖的事： “那数算的人在哪里？ 秤重的人在哪里？ 数点城楼的又在哪里呢？”
ISA|33|19|你必不再看见那凶暴的民， 他们嘴唇说艰涩的言语，难以理解； 舌头结巴，说无意义的话。
ISA|33|20|你要注视 锡安 ，我们守圣节的城！ 你必亲眼看见 耶路撒冷 成为安静的居所， 成为不挪移的帐幕， 橛子永不拔出， 绳索一根也不折断。
ISA|33|21|在那里，威严的耶和华对我们是宽阔的江河， 其中必没有摇桨的小船来往， 也没有巨大的船舶经过。
ISA|33|22|耶和华是审判我们的， 耶和华为我们设立律法； 耶和华是我们的君王， 他必拯救我们。
ISA|33|23|船上的绳索松开， 不能稳住桅杆， 也无法扬起船帆。 那时许多掳物被瓜分， 连瘸腿的也能夺走掠物。
ISA|33|24|城内的居民无人说：“我病了”； 城里居住的百姓，罪孽都蒙赦免。
ISA|34|1|列国啊，要近前来听！ 万民哪，要侧耳而听！ 全地和其上所充满的， 世界和其中所出的，都应当听！
ISA|34|2|因为耶和华向列国发怒， 向他们的全军发烈怒， 要将他们灭尽，任人杀戮。
ISA|34|3|被杀的人必被抛弃， 尸首臭气上腾， 诸山为他们的血所融化。
ISA|34|4|天上万象都要朽坏， 天被卷起，有如书卷， 其上的万象尽都衰残； 如葡萄树的叶子凋落， 又如无花果树枯萎一样。
ISA|34|5|因为我的刀在天上将要显现 ； 看哪，这刀临到 以东 和我所诅咒的民， 要施行审判。
ISA|34|6|耶和华的刀沾满了血， 是用油脂和羔羊、公山羊的血， 并公绵羊肾上的油脂滋润的； 因为在 波斯拉 有祭物献给耶和华， 在 以东 地有大屠杀。
ISA|34|7|野牛与他们一起倒下， 牛犊和壮牛也一同倒下。 他们的地被血染遍， 他们的尘土因油脂肥润。
ISA|34|8|这是耶和华报仇之日， 为 锡安 伸冤的报应之年。
ISA|34|9|它的河水要变为柏油， 尘埃变为硫磺， 大地成为燃烧的柏油，
ISA|34|10|昼夜总不熄灭， 它的烟永远上腾， 必世世代代成为荒废， 永永远远无人经过。
ISA|34|11|鹈鹕、豪猪要得它为业， 猫头鹰、乌鸦要住在其间。 耶和华必将空虚的准绳、 混沌的石垂线，拉在 以东 之上。
ISA|34|12|人必宣称那里没有王国， 它的贵族和所有领袖都归于无有。
ISA|34|13|以东 的宫殿要长出荆棘， 城堡要生长蒺藜和刺草； 成为野狗的住处， 鸵鸟的居所。
ISA|34|14|野兽要和土狼相遇， 山羊鬼魔要与同伴对唱， 莉莉丝 必在那里栖身， 为自己寻找安歇之处。
ISA|34|15|箭头蛇要在那里做窝， 下蛋，孵蛋，并招聚幼蛇在其保护之下； 鹞鹰也与伴侣聚集在那里。
ISA|34|16|你们要查考并诵读耶和华的书； 这些现象必然存在， 没有一样动物缺少伴侣。 因为是他，藉着我的口 吩咐， 他的灵将它们聚集。
ISA|34|17|他为它们抽签， 亲手用准绳为它们分地； 直到它们永远得地为业， 世世代代住在其间。
ISA|35|1|旷野和干旱之地必然欢喜， 沙漠也必快乐； 又如玫瑰绽放，
ISA|35|2|朵朵繁茂， 其乐融融，而且欢呼。 黎巴嫩 的荣耀， 并 迦密 与 沙仑 的华美，必赐给它。 人要看见耶和华的荣耀， 看见我们上帝的荣美。
ISA|35|3|你们要使软弱的手强壮， 使无力的膝盖稳固；
ISA|35|4|对心里焦急的人说： “要刚强，不要惧怕。 看哪，你们的上帝要来施报， 要施行极大的报应， 他必来拯救你们。”
ISA|35|5|那时，盲人的眼必睁开， 聋子的耳必开通。
ISA|35|6|那时，瘸子必跳跃如鹿， 哑巴的舌头必欢呼。 在旷野有水喷出， 在沙漠有江河涌流。
ISA|35|7|火热之地要变为水池， 干渴之地要变为泉源。 野狗躺卧休息之处 必长出青草、芦苇和蒲草。
ISA|35|8|在那里必有一条大道， 就是一条路 ，称为圣路。 污秽的人不得经过， 是专为走路的人 预备的， 愚昧的人也不会迷路。
ISA|35|9|在那里没有狮子， 猛兽也不经过； 在那里它们未现踪迹， 只有救赎的民在那里行走。
ISA|35|10|耶和华救赎的民必归回， 歌唱来到 锡安 ； 永远的快乐必归到他们头上， 他们必得着欢喜快乐， 忧伤叹息尽都逃避。
ISA|36|1|希西家 王十四年， 亚述 王 西拿基立 上来攻击 犹大 的一切坚固的城，将城攻取。
ISA|36|2|亚述 王从 拉吉 差遣将军 率领大军前往 耶路撒冷 ，到 希西家 王那里去。将军站在 上池 的水沟旁，在往漂布地的大路上。
ISA|36|3|希勒家 的儿子 以利亚敬 宫廷总管、 舍伯那 书记和 亚萨 的儿子 约亚 史官，出来见他。
ISA|36|4|将军对他们说：“你们去告诉 希西家 ，大王 亚述 王如此说：‘你倚靠什么，让你如此自信满满？
ISA|36|5|我说 ，你有打仗的计谋和能力，我看不过是空话。你到底倚靠谁，竟敢背叛我呢？
ISA|36|6|看哪，你所倚靠的 埃及 是那断裂的苇杖，人若倚靠这杖，它就刺进他的手，穿透它。 埃及 王法老向所有倚靠他的人都是这样。
ISA|36|7|你若对我说：我们倚靠耶和华－我们的上帝， 希西家 岂不是将上帝的丘坛和祭坛废去，并且吩咐 犹大 和 耶路撒冷 的人说：你们只当在这一个坛前敬拜吗？
ISA|36|8|现在你与我主 亚述 王打赌，我给你两千匹马，看你能否派得出骑士来骑它们。
ISA|36|9|若不然，怎能使我主臣仆中最小的一个军官转脸而逃呢？你难道要倚靠 埃及 的战车和骑兵吗？
ISA|36|10|现在我上来攻击毁灭这地，岂不是出于耶和华吗？耶和华吩咐我说，你上去攻击这地，毁灭它吧！’”
ISA|36|11|以利亚敬 、 舍伯那 、 约亚 对将军说：“求你用 亚兰 话对仆人说，因为我们听得懂；不要用 犹大 话对我们说，免得传到城墙上百姓的耳中。”
ISA|36|12|将军说：“我主差遣我来，岂是单对你和你的主人说这些话吗？不也是对这些坐在城墙上，要与你们一同吃自己粪、喝自己尿的人说的吗？”
ISA|36|13|于是 亚述 将军站着，用 犹大 话大声喊着说：“你们当听大王 亚述 王的话，
ISA|36|14|王如此说：‘你们不要被 希西家 欺哄了，因他不能拯救你们。
ISA|36|15|不要听凭 希西家 说服你们倚靠耶和华，他说，耶和华必要拯救我们，这城必不交在 亚述 王的手中。’
ISA|36|16|你们不要听 希西家 的话！因 亚述 王如此说：‘你们要与我讲和，出来投降，各人就可以吃自己葡萄树和无花果树的果子，喝自己井里的水，
ISA|36|17|等我来领你们到一个地方，与你们本地一样，就是有五谷和新酒之地，有粮食和葡萄园之地。
ISA|36|18|恐怕 希西家 误导你们说，耶和华必拯救我们。列国的神明有哪一个曾救它本国脱离 亚述 王的手呢？
ISA|36|19|哈马 和 亚珥拔 的神明在哪里呢？ 西法瓦音 的神明在哪里呢？它们曾救 撒玛利亚 脱离我的手吗？
ISA|36|20|这些国的神明有谁曾救自己的国家脱离我的手呢？难道耶和华能救 耶路撒冷 脱离我的手吗？’”
ISA|36|21|百姓静默不言，一句不答，因为 希西家 王曾吩咐说：“不要回答他。”
ISA|36|22|当下 希勒家 的儿子 以利亚敬 宫廷总管、 舍伯那 书记，和 亚萨 的儿子 约亚 史官都撕裂衣服，来到 希西家 那里，将 亚述 将军的话告诉他。
ISA|37|1|希西家 王听见了，就撕裂衣服，披上麻布，进了耶和华的殿。
ISA|37|2|他差遣 以利亚敬 宫廷总管和 舍伯那 书记，并祭司中年长的，都披上麻布，到 亚摩斯 的儿子 以赛亚 先知那里去。
ISA|37|3|他们对他说：“ 希西家 如此说：‘今日是急难、惩罚、凌辱的日子，就如婴孩快要出生，却没有力气生产。
ISA|37|4|或许耶和华－你的上帝听见 亚述 将军的话，就是他主人 亚述 王差他来辱骂永生上帝的话，耶和华－你的上帝就斥责所听见的这些话。求你为幸存的余民扬声祷告。’”
ISA|37|5|希西家 王的臣仆就来到 以赛亚 那里。
ISA|37|6|以赛亚 对他们说：“要对你们的主人这样说，耶和华如此说：‘你听见 亚述 王的仆人亵渎我的话，不要惧怕。
ISA|37|7|看哪，因为我必惊动他的心 ，他要听见风声就归回本地，在那里我必使他倒在刀下。’”
ISA|37|8|亚述 将军听见 亚述 王已拔营离开 拉吉 ，就启程返回，正遇见 亚述 王去攻打 立拿 。
ISA|37|9|亚述 王听见有人谈论 古实 王 特哈加 说：“他出来要与你争战。” 亚述 王一听见，就差使者去见 希西家 ，说：
ISA|37|10|“你们要对 犹大 王 希西家 如此说：‘不要听你所倚靠的上帝欺哄你说： 耶路撒冷 必不交在 亚述 王的手中。
ISA|37|11|看哪，你总听说 亚述 诸王向列国所行的是尽行灭绝，难道你能幸免吗？
ISA|37|12|我祖先所毁灭的，就是 歌散 、 哈兰 、 利色 和 提．拉撒 的 伊甸 人；这些国的神明何曾拯救他们呢？
ISA|37|13|哈马 的王， 亚珥拔 的王， 西法瓦音城 的王， 希拿 和 以瓦 的王，都在哪里呢？’”
ISA|37|14|希西家 从使者手里接过书信，看完了，就上耶和华的殿，在耶和华面前展开书信。
ISA|37|15|希西家 向耶和华祷告说：
ISA|37|16|“坐在基路伯之上万军之耶和华－ 以色列 的上帝啊，你，惟有你是地上万国的上帝，你创造了天和地。
ISA|37|17|耶和华啊，求你侧耳而听；耶和华啊，求你睁眼而看，听 西拿基立 差遣使者辱骂永生上帝的一切话。
ISA|37|18|耶和华啊， 亚述 诸王果然使列国和列国之地变为荒芜，
ISA|37|19|将列国的神明扔在火里，因为它们不是神明，是人手所造的，是木头、石头，所以被灭绝了。
ISA|37|20|耶和华－我们的上帝啊，现在求你救我们脱离 亚述 王的手，使地上万国都知道惟有你是耶和华。”
ISA|37|21|亚摩斯 的儿子 以赛亚 就差人去见 希西家 ，说：“耶和华－ 以色列 的上帝如此说，你因 亚述 王 西拿基立 的事向我祈求，
ISA|37|22|所以耶和华论他这样说： ‘少女 锡安 藐视你，嘲笑你； 耶路撒冷 向你摇头。
ISA|37|23|“‘你辱骂谁，亵渎谁， 扬起声来，高举眼目攻击谁呢？ 你攻击的是 以色列 的圣者。
ISA|37|24|你藉臣仆辱骂主说： 我率领许多战车登上高山， 到 黎巴嫩 的顶端； 我要砍伐其中高大的香柏树 和上好的松树。 我必上到极高之处， 进入茂盛的森林里。
ISA|37|25|我已经挖井喝水 我必用脚掌踏干 埃及 一切的河流。
ISA|37|26|“‘你岂没有听见 我早先所定、古时所立、现今实现的事吗？ 就是让你去毁坏坚固的城镇，使它们变为废墟；
ISA|37|27|城里居民的力量甚小， 他们惊惶羞愧； 像野草，像青菜， 如房顶上的草， 被东风刮散 。
ISA|37|28|“‘你站起，你坐下，你出去，你进来， 你向我发烈怒，我都知道。
ISA|37|29|因你向我发烈怒， 你的狂傲上达我耳中， 我要用钩子钩住你的鼻子， 将嚼环放在你口里， 使你从原路转回去。’
ISA|37|30|“我赐给你的预兆：你们今年要吃野生的，明年也要吃自长的；后年，你们就要耕种收割，栽葡萄园，吃其中的果子。
ISA|37|31|犹大 家所逃脱剩余的，仍要往下扎根，向上结果。
ISA|37|32|必有剩余的民从 耶路撒冷 而出；有逃脱的人从 锡安山 而来。万军之耶和华的热心必成就这事。
ISA|37|33|“所以耶和华论 亚述 王如此说：他必不得来到这城，也不在这里射箭，不得拿盾牌到城前，也不能建土堆攻城。
ISA|37|34|他从哪条路来，必从那条路回去，必不得来到这城。这是耶和华说的。
ISA|37|35|因我为自己的缘故，又为我仆人 大卫 的缘故，必保护拯救这城。”
ISA|37|36|耶和华的使者出去，在 亚述 营中杀了十八万五千人。清早有人起来，看哪，都是死尸。
ISA|37|37|亚述 王 西拿基立 就拔营回去，住在 尼尼微 。
ISA|37|38|一日，他在他的神明 尼斯洛 庙里叩拜，他儿子 亚得米勒 和 沙利色 用刀杀了他，然后逃到 亚拉腊 地；他儿子 以撒．哈顿 接续他作王。
ISA|38|1|那些日子， 希西家 病得要死， 亚摩斯 的儿子 以赛亚 先知来见他，对他说：“耶和华如此说：‘你当留遗嘱给你的家，因为你必死，不能活了。’”
ISA|38|2|希西家 就转脸朝墙，向耶和华祷告，
ISA|38|3|说：“耶和华啊，求你记念我在你面前怎样存完全的心，按诚实行事，又做你眼中看为善的事。” 希西家 就痛哭。
ISA|38|4|耶和华的话临到 以赛亚 说：
ISA|38|5|“你去告诉 希西家 说，耶和华－你祖先 大卫 的上帝如此说：‘我听见了你的祷告，看见了你的眼泪。看哪，我必加添你十五年的寿数；
ISA|38|6|我要救你和这城脱离 亚述 王的手，也要保护这城。’
ISA|38|7|“耶和华必成就他所说的这话。这是耶和华给你的预兆：
ISA|38|8|看哪，我要使 亚哈斯 日晷上随太阳前进的影子，往后退十度。”于是，在日晷上照下来的日影果然往后退了十度。
ISA|38|9|犹大 王 希西家 患病痊愈后的诗：
ISA|38|10|我说，在如日中天的时候我就走了， 将剩余的年岁交给阴间的门。
ISA|38|11|我说，我必不得见耶和华，不得在活人之地见耶和华， 也不再看见世人，就是短暂世界 中的居民。
ISA|38|12|我的住处好像牧人的帐棚， 遭人掀起，离我而去； 我将性命卷起， 像织布的卷布一样。 他从织布机头那里将我剪断， 你使我命丧于旦夕。
ISA|38|13|我令自己安静 直到天亮； 他像狮子折断我所有的骨头， 你使我命丧于旦夕。
ISA|38|14|我像燕子呢喃， 像白鹤鸣叫， 又如鸽子哀鸣； 我因仰望，眼睛困倦。 主啊，我受欺压， 求你为我作保。
ISA|38|15|我还有什么可说的呢？ 他应许我的 ，他已成就了。 我因心里的苦楚， 在一生的年日必谦卑而行 。
ISA|38|16|主啊，人得存活是在乎此， 我的灵存活也全在乎此 ； 求你使我痊愈，仍然存活。
ISA|38|17|看哪，我受大苦是为使我得平安； 你爱我，救我的性命脱离败坏的地府， 将我一切的罪扔在你背后。
ISA|38|18|原来，阴间不能称谢你， 死亡不能颂扬你， 下到地府的人也不能盼望你的信实。
ISA|38|19|只有活人，活人必称谢你， 像我今日称谢你一样。 为父的，必使儿女知道你的信实。
ISA|38|20|耶和华肯救我， 所以，我们要一生一世 在耶和华殿中 弹奏我弦乐的歌。
ISA|38|21|以赛亚 说：“拿一块无花果饼来，贴在疮上，王必痊愈。”
ISA|38|22|希西家 说：“我能上耶和华的殿，有什么预兆呢？”
ISA|39|1|那时， 巴拉但 的儿子， 巴比伦 王 米罗达．巴拉但 听见 希西家 病得痊愈，就送书信和礼物给他。
ISA|39|2|希西家 欢喜见使者，就将自己宝库里的金子、银子、香料、贵重的膏油和他军械库里一切的兵器，以及他所有的财宝，都给他们看；在他家中和全国之内， 希西家 没有一样不给他们看的。
ISA|39|3|于是 以赛亚 先知到 希西家 王那里去，对他说：“这些人说了些什么？他们从哪里来见你？” 希西家 说：“他们从远方的 巴比伦 来见我。”
ISA|39|4|以赛亚 说：“他们在你家里看见了什么？” 希西家 说：“凡我家中所有的，他们都看见了；我财宝中没有一样东西不给他们看的。”
ISA|39|5|以赛亚 对 希西家 说：“你要听万军之耶和华的话，
ISA|39|6|耶和华说：‘看哪，日子将到，凡你家里所有的，并你祖先积蓄到如今的一切，都要被掳到 巴比伦 去，不留下一样；
ISA|39|7|从你本身所生的孩子，其中必有被掳到 巴比伦 王宫当太监的。’”
ISA|39|8|希西家 对 以赛亚 说：“你所说耶和华的话甚好。”因为他想：“在我有生之年必有太平和安稳。”
ISA|40|1|你们的上帝说： “要安慰，安慰我的百姓。
ISA|40|2|要对 耶路撒冷 说安慰的话， 向它宣告， 它的战争已结束， 它的罪孽已赦免； 它为自己一切的罪， 已从耶和华手中加倍受罚。”
ISA|40|3|有声音呼喊着： “要在旷野为耶和华预备道路， 在沙漠为我们的上帝修直大道。
ISA|40|4|一切山洼都要填满， 大小山冈都要削平； 陡峭的要变为平坦， 崎岖的必成为平原。
ISA|40|5|耶和华的荣耀必然显现， 凡有血肉之躯的都一同看见， 因为这是耶和华亲口说的。”
ISA|40|6|有声音说：“你喊叫吧！” 我 说：“我喊叫什么呢？” 凡有血肉之躯的尽都如草， 他的一切荣美像野地的花。
ISA|40|7|耶和华吹一口气， 草就枯干，花也凋谢。 百姓诚然是草；
ISA|40|8|草必枯干，花必凋谢， 惟有我们上帝的话永远立定。
ISA|40|9|报好信息的 锡安 哪， 要登高山； 报好信息的 耶路撒冷 啊， 要极力扬声。 扬声不要惧怕， 对 犹大 的城镇说： “看哪，你们的上帝！”
ISA|40|10|看哪，主耶和华必以大能临到， 他的膀臂必为他掌权； 看哪，他的赏赐在他那里， 他的报应在他面前。
ISA|40|11|他要像牧人牧养自己的羊群， 用膀臂聚集羔羊，抱在胸怀， 慢慢引导那乳养小羊的。
ISA|40|12|谁曾用手心量诸水， 用手虎口量苍天， 用升斗盛大地的尘土， 用秤称山岭， 用天平称冈陵呢？
ISA|40|13|谁曾测度耶和华的灵， 或作他的谋士指教他呢？
ISA|40|14|他与谁商议， 谁教导他， 以公平的路指示他， 将知识传授与他， 又将通达的道指教他呢？
ISA|40|15|看哪，列国都像水桶里的一滴， 又如天平上的微尘； 看哪，他举起众海岛，好像举起极微小之物。
ISA|40|16|黎巴嫩 不够当柴烧， 其中的走兽也不够作燔祭。
ISA|40|17|列国在他面前如同不存在， 在他看来微不足道，只是虚空。
ISA|40|18|你们究竟将谁比上帝， 用什么形像与他相较呢？
ISA|40|19|至于偶像，匠人铸造它， 银匠用金子包裹它， 又为它铸造银链。
ISA|40|20|没有能力捐献的人， 就挑选不易朽坏的木头， 为自己寻找巧匠， 竖立不会倒的偶像。
ISA|40|21|你们岂不知道吗？ 岂未曾听见吗？ 难道没有人从起头就告诉你们吗？ 自从地的根基立定， 你们岂不明白吗？
ISA|40|22|上帝坐在地的穹窿之上， 地上的居民有如蚱蜢。 他铺张穹苍如幔子， 展开诸天如可住的帐棚。
ISA|40|23|他使君王归于虚无， 使地上的审判官成为虚空。
ISA|40|24|他们刚栽上， 刚种好， 根也刚扎在地里， 经他一吹，就都枯干； 旋风将他们吹去，像碎秸一样。
ISA|40|25|那圣者说：“你们将谁与我相比， 与我相等呢？”
ISA|40|26|你们要向上举目， 看是谁创造这万象， 按数目领出它们， 一一称其名， 以他的权能 和他的大能大力， 使它们一个都不缺。
ISA|40|27|雅各 啊，你为何说， 以色列 啊，你为何言， “我的道路向耶和华隐藏， 我的冤屈上帝并不查问”？
ISA|40|28|你岂不曾知道吗？ 你岂未曾听见吗？ 永在的上帝耶和华，创造地极的主， 他不疲乏，也不困倦； 他的智慧无法测度。
ISA|40|29|疲乏的，他赐能力； 软弱的，他加力量。
ISA|40|30|就是年轻人也要疲乏困倦， 强壮的也必全然跌倒。
ISA|40|31|但那等候耶和华的必重新得力。 他们必如鹰展翅上腾； 他们奔跑却不困倦， 行走却不疲乏。
ISA|41|1|众海岛啊，在我面前静默； 万民要重新得力， 让他们近前来陈述， 我们可以彼此辩论。
ISA|41|2|谁从东方兴起一人， 凭公义召他来到脚前？ 谁将列国交给他， 使他管辖列王， 把他们如灰尘交与他的刀， 如风吹的碎秸交与他的弓？
ISA|41|3|他追赶君王， 安然走过， 快速地脚不落地 。
ISA|41|4|谁做成这事， 从起初宣召历代呢？ 就是我－耶和华！ 我是首先的， 也与末后的同在。
ISA|41|5|众海岛看见就都害怕， 地极也都战兢， 他们近前来；
ISA|41|6|各人互相帮助， 对弟兄说：“壮胆吧！”
ISA|41|7|木匠鼓励银匠， 用锤子打光的鼓励打砧的， 对焊工说：“焊得好！” 又用钉子钉稳，免得它倒下。
ISA|41|8|惟你 以色列 ，我的仆人， 雅各 ，我所拣选的， 我朋友 亚伯拉罕 的后裔，
ISA|41|9|你是我从地极领来， 从地角召来的， 我对你说：“你是我的仆人； 我拣选你，并不弃绝你。”
ISA|41|10|你不要害怕，因为我与你同在； 不要惊惶，因为我是你的上帝。 我必坚固你，帮助你， 用我公义的右手扶持你。
ISA|41|11|看哪，凡向你发怒的都抱愧蒙羞， 与你相争的必如无有，并要灭亡。
ISA|41|12|与你争斗的，你要寻找他们，却遍寻不着； 与你争战的必如无有，成为虚无。
ISA|41|13|因为我耶和华－你的上帝 必搀扶你的右手， 对你说：“不要害怕！ 我必帮助你。”
ISA|41|14|虫子 雅各 ， 以色列 人哪， 不要害怕！ 我必帮助你； 救赎你的是 以色列 的圣者。 这是耶和华说的。
ISA|41|15|看哪，我使你成为 全新的打谷机，齿轮锐利； 你要把山岭打得粉碎， 使冈陵如同糠秕。
ISA|41|16|你要簸扬它们，风要将它们吹去； 旋风要刮散它们。 你却要以耶和华为喜乐， 因 以色列 的圣者夸耀。
ISA|41|17|困苦贫穷人寻找水，却寻不着； 他们因口渴，舌头干燥。 我－耶和华必应允他们， 我─ 以色列 的上帝必不离弃他们。
ISA|41|18|我要在光秃的高地开江河， 在谷中开泉源； 我要使沙漠变为水池， 使干地变为涌泉。
ISA|41|19|我要在旷野栽植香柏树、 皂荚树、番石榴树，和野橄榄树。 在沙漠一同栽上松树、杉树， 和黄杨树，
ISA|41|20|好叫人看见，知道， 思想，明白； 这是耶和华亲手做的， 是 以色列 的圣者所造的。
ISA|41|21|耶和华说： “你们要呈上你们的案件。” 雅各 的君王说： “你们要提出你们的理由。”
ISA|41|22|让它们近前来，告诉我们将来要发生什么事！ 你们要说明先前发生的事，好让我们思索； 或者告诉我们将来的事，使我们得知事情的结局。
ISA|41|23|你们要指明未来的事， 使我们知道你们是神明！ 你们或降福，或降祸， 好使我们惊奇，一同观看。
ISA|41|24|看哪，你们属乎虚无， 你们的作为也属虚空； 那选择你们的是可憎恶的。
ISA|41|25|我从北方兴起一人， 他从日出之地而来， 是求告我名的； 他必踩踏 掌权者，如踩踏泥土， 又如陶匠踹泥一般。
ISA|41|26|有谁从起初宣布这事，使我们知道呢？ 有谁从先前指明，使我们说“他是对的”呢？ 没有人宣布， 没有人指明， 也没有人听见你们的话。
ISA|41|27|我首先对 锡安 说，看哪，他们在此！ 我要将一位报好信息的赐给 耶路撒冷 。
ISA|41|28|然而我观看，并无一人； 我询问的时候， 他们中间也没有谋士可回答。
ISA|41|29|看哪，他们尽是麻烦 ， 所做的工都属虚无； 所铸的偶像是风，是虚空。
ISA|42|1|看哪，我的仆人， 我所扶持、所拣选、心所喜悦的！ 我已将我的灵赐给他， 他必将公理传给万邦。
ISA|42|2|他不喧嚷，不扬声， 也不使街上听见他的声音。
ISA|42|3|压伤的芦苇，他不折断； 将残的灯火，他不吹灭。 他凭信实将公理传开。
ISA|42|4|他不灰心，也不丧胆， 直到他在地上设立公理； 众海岛都等候他的训诲。
ISA|42|5|那创造诸天，铺张穹苍， 铺开地与地的出产， 赐气息给地上众人， 赐生命给行走其上之人的 上帝耶和华如此说：
ISA|42|6|“我－耶和华凭公义召你， 要搀扶你的手，保护你， 要藉着你与百姓立约， 使你成为万邦之光，
ISA|42|7|开盲人的眼， 领囚犯出监狱， 领坐在黑暗中的出地牢。
ISA|42|8|我是耶和华，这是我的名； 我必不将我的荣耀归给别神 ， 也不将我所得的颂赞归给雕刻的偶像。
ISA|42|9|看哪，先前的事已经成就， 现在我要指明新事， 告诉你们尚未发生的事。
ISA|42|10|航海的人和海中一切所有的， 众海岛和其中的居民， 都当向耶和华唱新歌， 从地极赞美他。
ISA|42|11|旷野和其中的城镇， 并 基达 人居住的村庄都当扬声 ； 西拉 的居民当欢呼， 在山顶上大声呼喊。
ISA|42|12|愿他们将荣耀归给耶和华， 在海岛中传扬颂赞他的话。
ISA|42|13|耶和华必如勇士出征， 如战士激起愤恨， 他要喊叫，大声呐喊， 击败他的敌人。
ISA|42|14|我许久闭口不言，沉默不语； 现在我要像临产的妇人，大声喊叫， 呼吸急促而喘气。
ISA|42|15|我要使大小山冈变为荒芜， 使其上的花草都枯干； 我要使江河变为沙洲， 使水池尽都干涸。
ISA|42|16|我要引导盲人行他们所不认识的道， 引领他们走他们未曾走过的路； 我在他们面前使黑暗变为光明， 使弯曲变为平直。 这些事我都要做， 并不离弃他们。
ISA|42|17|但那倚靠雕刻的偶像， 对铸造的偶像说： “你是我们的神明”； 这种人要退后，大大蒙羞。
ISA|42|18|你们这耳聋的，听吧！ 你们这眼瞎的，看吧， 使你们得以看见！
ISA|42|19|谁比我的仆人眼瞎呢？ 谁比我所差遣的使者耳聋呢？ 谁瞎眼像那献身给我的人？ 谁瞎眼 像耶和华的仆人呢？
ISA|42|20|看见许多事却不领会， 耳朵开通却听不见。
ISA|42|21|耶和华因自己的公义， 乐意使律法为大为尊。
ISA|42|22|但这百姓是被抢被夺的， 全都陷在洞穴中，关在监牢里； 他们成了掠物，无人拯救， 成了掳物，无人索还。
ISA|42|23|你们中间谁肯侧耳听这话， 谁肯留心听，以防将来呢？
ISA|42|24|谁将 雅各 交出作为掳物， 将 以色列 交给抢夺者呢？ 岂不是耶和华 ─我们所得罪的那位吗？ 他们不肯遵行他的道， 也不听从他的训诲。
ISA|42|25|所以，他将猛烈的怒气和战争的威力 倾倒在 以色列 身上； 在他周围如火燃起，他竟然不知， 烧着了，他也不在意。
ISA|43|1|雅各 啊，创造你的耶和华， 以色列 啊，造成你的那位， 现在如此说： “你不要害怕，因为我救赎了你； 我曾提你的名召你，你是属我的。
ISA|43|2|你从水中经过，我必与你同在， 你渡过江河，水必不漫过你； 你在火中行走，也不被烧伤， 火焰必不烧着你身。
ISA|43|3|因为我是耶和华－你的上帝， 是 以色列 的圣者－你的救主； 我使 埃及 作你的赎价， 使 古实 和 西巴 代替你。
ISA|43|4|因我看你为宝贝为尊贵； 又因我爱你， 所以使人代替你， 使万民替换你的生命。
ISA|43|5|你不要害怕，因我与你同在； 我必领你的后裔从东方来， 又从西方召集你。
ISA|43|6|我要对北方说，交出来！ 对南方说，不可扣留！ 要将我的儿子从远方带来， 将我的女儿从地极领回，
ISA|43|7|就是凡称为我名下的人， 是我为自己的荣耀创造的， 是我所塑造，所做成的。”
ISA|43|8|你要将有眼却瞎、 有耳却聋的民都带出来！
ISA|43|9|任凭万国聚集， 任凭万民会合。 他们当中谁能说明， 并将先前的事指示我们呢？ 让他们带来见证，显明他们有理， 看是否听见的人会说：“果然是真的。”
ISA|43|10|你们是我的见证， 是我所拣选的仆人， 为了要使你们知道，且信服我， 又明白我就是耶和华。 在我以前没有任何被造的真神， 在我以后也必没有。 这是耶和华说的。
ISA|43|11|我，惟有我是耶和华； 除我以外没有救主。
ISA|43|12|我曾指示，我曾拯救，我曾说明， 并没有外族的神明 在你们中间。 你们是我的见证， 我是上帝。 这是耶和华说的。
ISA|43|13|自有日子以来，我就是上帝， 谁也不能救人脱离我的手。 我要行事，谁能逆转呢？
ISA|43|14|耶和华─你们的救赎主、 以色列 的圣者如此说： “因你们的缘故， 我已派遣人到 巴比伦 去； 要使 迦勒底 人都如难民， 坐自己素来宴乐的船下来。
ISA|43|15|我是耶和华－你们的圣者， 是创造 以色列 的，是你们的君王。”
ISA|43|16|那在沧海中开道， 在大水中开路， 使战车、马匹、军兵、勇士一同出来， 使他们仆倒，不再起来， 使他们灭没，好像熄灭之灯火的耶和华如此说：
ISA|43|17|
ISA|43|18|“你们不要追念从前的事， 也不要思想古时的事。
ISA|43|19|看哪，我要行一件新事， 如今就要显明，你们岂不知道吗？ 我必在旷野开道路， 在沙漠开江河 。
ISA|43|20|野地的走兽要尊敬我， 野狗和鸵鸟也必尊敬我。 因我使旷野有水， 使沙漠有河， 好赐给我的百姓、我的选民喝。
ISA|43|21|这百姓是我为自己造的， 为要述说我的美德。”
ISA|43|22|“ 雅各 啊，你并没有求告我； 以色列 啊，你倒厌烦我。
ISA|43|23|你并没有将你的羊带来献给我做燔祭， 也没有用牲祭尊敬我； 我未曾因素祭使你操劳， 也没有因乳香使你厌烦。
ISA|43|24|你没有用银子为我买香菖蒲， 也没有用祭物的油脂使我饱足； 倒使我因你的罪恶操劳， 使我因你的罪孽厌烦。
ISA|43|25|我，惟有我为自己的缘故涂去你的过犯， 我也不再记得你的罪恶。
ISA|43|26|你尽管提醒我，让我们来辩论； 尽管陈述，自显为义。
ISA|43|27|你的始祖犯罪， 你的师傅违背我；
ISA|43|28|因此，我要凌辱圣所的领袖 ， 使 雅各 遭毁灭， 使 以色列 受辱骂。”
ISA|44|1|“我的仆人 雅各 ， 我所拣选的 以色列 啊， 现在你当听。
ISA|44|2|那位造你，使你在母腹中成形， 并要帮助你的耶和华如此说： 我的仆人 雅各 ， 我所拣选的 耶书仑 哪， 不要害怕！
ISA|44|3|因为我要把水浇灌干渴的地方， 使水涌流在干旱之地。 我要将我的灵浇灌你的后裔， 使我的福临到你的子孙。
ISA|44|4|他们要在草丛中生长 ， 如溪水旁的柳树。
ISA|44|5|这个要说：‘我是属耶和华的’， 那个要以 雅各 的名自称， 又有一个在手上写着：‘归耶和华’， 并自称为 以色列 。”
ISA|44|6|耶和华－ 以色列 的君王， 以色列 的救赎主－万军之耶和华如此说： “我是首先的，也是末后的； 除我以外再没有上帝。
ISA|44|7|自从古时我设立了人， 谁能像我宣告，指明，又为自己陈说呢？ 让他指明未来的事和必成的事吧！
ISA|44|8|你们不要恐惧，也不要害怕。 我岂不是从上古就告诉并指示你们了吗？ 你们是我的见证人！ 除我以外，岂有上帝呢？ 诚然没有磐石，就我所知，一个也没有！”
ISA|44|9|制造偶像的人尽都虚空，他们所喜悦的全无益处；偶像的见证人毫无所见，毫无所知，以致他们羞愧。
ISA|44|10|谁制造神像，铸造偶像？这些都是无益的。
ISA|44|11|看哪，他的同伙都必羞愧。工匠不过是人，任他们聚集，任他们站立吧！他们都必惧怕，一同羞愧。
ISA|44|12|铁匠用工具在火炭上工作 ，用锤打出形状，用他有力的膀臂来锤。他因饥饿而无力气；因未喝水而疲倦。
ISA|44|13|木匠拉线，用笔划出样子，用刨子刨成形状，又用圆规划了模样。他仿照人的体态，做出美妙的人形，放在庙里。
ISA|44|14|他砍伐香柏树，又取杉树和橡树，在树林中让它茁壮；或栽种松树，得雨水滋润长大。
ISA|44|15|这树，人可用以生火；他拿一些来取暖，又搧火烤饼，而且做神像供跪拜，做雕刻的偶像向它叩拜。
ISA|44|16|他将一半的木头烧在火中，用它烤肉来吃；吃饱了，就自己取暖说：“啊哈，我暖和了，我看到火了！”
ISA|44|17|然后又用剩下的一半做了一个神明，就是雕刻的偶像，向这偶像俯伏叩拜，向它祷告说：“求你拯救我，因你是我的神明。”
ISA|44|18|他们既无知，又不思想；因为耶和华蒙蔽他们的眼，使他们看不见，塞住他们的心，使他们不明白。
ISA|44|19|没有一个心里醒悟，有知识，有聪明，能说：“我曾拿一部分用火燃烧，在炭火上烤饼，也烤肉来吃。这剩下的，我岂要做可憎之像吗？我岂可向木头叩拜呢？”
ISA|44|20|他以灰尘为食，心里迷糊，以致偏邪，不能自救，也不能说：“我右手中岂不是有虚谎吗？”
ISA|44|21|雅各 啊，要思念这些事； 以色列 啊，你是我的仆人。 我造了你，你是我的仆人， 以色列 啊，我必不忘记你 。
ISA|44|22|我涂去你的过犯，像厚云消散； 涂去你的罪恶，如薄雾消失。 你当归向我，因我救赎了你。
ISA|44|23|诸天哪，应当歌唱， 因为耶和华成就这事。 地的深处啊，应当欢呼； 众山哪，要出声歌唱； 树林和其中所有的树木啊，你们都当歌唱！ 因为耶和华救赎了 雅各 ， 并要因 以色列 荣耀自己。
ISA|44|24|从你在母腹中就造了你，你的救赎主－耶和华如此说： “我－耶和华创造万物， 独自铺张诸天，亲自展开大地 ；
ISA|44|25|我使虚谎的预兆失效， 愚弄占卜的人， 使智慧人退后， 使他的知识变为愚拙；
ISA|44|26|却使我仆人的话站得住， 成就我使者的筹算。 我论 耶路撒冷 说：‘必有人居住’； 论 犹大 的城镇说：‘必被建造， 我必重建其中的废墟。’
ISA|44|27|我对深渊说：‘干了吧！ 我要使你的江河干涸’；
ISA|44|28|论 居鲁士 说：‘他是我的牧人， 他要成就我所喜悦的， 下令建造 耶路撒冷 ， 发命令立稳圣殿的根基。’”
ISA|45|1|耶和华对所膏的 居鲁士 如此说， 他的右手我曾搀扶， 使列国降服在他面前， 列王的腰带我曾松开， 使城门在他面前敞开， 不得关闭：
ISA|45|2|“我要在你前面行， 修平崎岖之地。 我必打破铜门， 砍断铁闩。
ISA|45|3|我要将暗中的宝物和隐藏的财富赐给你， 使你知道提名召你的 就是我－耶和华， 以色列 的上帝。
ISA|45|4|因我的仆人 雅各 ， 我所拣选的 以色列 ， 我提名召你； 你虽不认识我， 我也加给你名号。
ISA|45|5|我是耶和华，再没有别的了； 除了我以外再没有上帝。 你虽不认识我， 我必给你束腰。
ISA|45|6|从日出之地到日落之处使人都知道 除我以外，没有别的。 我是耶和华，再没有别的了。
ISA|45|7|我造光，又造暗； 施平安，又降灾祸； 做成这一切的是我－耶和华。
ISA|45|8|“诸天哪，要如雨倾盆而降， 云要降下公义， 地要裂开，救恩涌出 ， 使公义也一同滋长； 这都是我－耶和华造的。”
ISA|45|9|“那与造他的主争论的人有祸了！ 他不过是地上瓦块中的一片 。 泥土岂可对塑造它的说：‘你做的是什么？ 你所做的物怎么没有把手呢？ ’
ISA|45|10|有人对父亲说， ‘你生的是什么’， 对母亲 说， ‘你生产的是什么’； 这人有祸了！”
ISA|45|11|耶和华－ 以色列 的圣者， 就是造 以色列 的如此说： “难道我孩子的未来，你们能质问我， 我手的工作，你们可以吩咐我吗？
ISA|45|12|我造大地，又创造人在地上。 我亲手铺张诸天， 天上万象也是我所任命的。
ISA|45|13|我凭公义兴起 居鲁士 ， 又要修直他一切的道路。 他必建造我的城， 释放我被掳的民， 不为工价，也不为奖赏。” 这是万军之耶和华说的。
ISA|45|14|耶和华如此说： “ 埃及 的出产和 古实 的货物必归你； 身量高大的 西巴 人，他们必过来归你，为你所有。 他们必带着锁链过来跟随你， 向你下拜，祈求你说： ‘上帝真是在你中间，再没有别的， 没有别的上帝。’”
ISA|45|15|救主－ 以色列 的上帝啊， 你诚然是隐藏自己的上帝。
ISA|45|16|制造偶像的都要抱愧蒙羞， 他们要一同归于惭愧。
ISA|45|17|惟有 以色列 必蒙耶和华拯救， 得永远的救恩。 你们必不蒙羞，也不抱愧， 直到永世无尽。
ISA|45|18|耶和华如此说， 他创造诸天，他是上帝； 他造了地，形成它，坚固它， 并非创造它为荒凉， 而是要给人居住： “我是耶和华，再没有别的。
ISA|45|19|我不在隐密黑暗之地说话， 也没有对 雅各 的后裔说， ‘你们寻求我是徒然的’， 我－耶和华所讲的是公义， 所说的是正直。”
ISA|45|20|“你们从列国逃脱的人， 要一同聚集前来。 那些抬着雕刻的木偶、 祈求不能救人之神明的， 毫无知识。
ISA|45|21|你们要近前来说明， 让他们彼此商议。 谁从古时指明这事？ 谁从上古述说它？ 不是我－耶和华吗？ 除了我以外，再没有上帝； 我是公义的上帝，又是救主； 除了我以外，再没有别的了。
ISA|45|22|“地的四极都当转向我， 就必得救； 因为我是上帝，再没有别的。
ISA|45|23|我指着自己起誓， 公义从我的口发出，这话并不返回： ‘万膝必向我跪拜， 万口必凭我起誓。’
ISA|45|24|人论我说 ， “公义、能力，惟独在乎耶和华。 人必归向他， 凡向他发怒的都必蒙羞。
ISA|45|25|以色列 的后裔必因耶和华得称为义， 并要彼此夸耀。”
ISA|46|1|彼勒 叩拜， 尼波 屈身； 巴比伦 的偶像驮在走兽和牲畜背上。 你们所抬的成了重驮， 使牲畜疲乏。
ISA|46|2|这些神明一同屈身叩拜， 不能救自己 ， 反倒遭人掳去。
ISA|46|3|雅各 家， 以色列 家所有的余民哪， 你们自从生下就蒙我抱， 自出母胎便由我来背， 你们都要听从我。
ISA|46|4|直到你们年老，我不改变； 直到你们发白，我仍扶持。 我已造你，就必背你； 我必抱你，也必拯救。
ISA|46|5|你们将谁与我相比，与我相等， 将谁与我相较，使我们相似呢？
ISA|46|6|他们从钱囊中倒出金子， 用天平秤出银子， 雇银匠造成神像， 他们又俯伏，又叩拜。
ISA|46|7|他们抬起神像，扛在肩上， 安置在定处，使它站立， 不离本位； 人呼求它，它却不回答， 也无法救人脱离灾难。
ISA|46|8|你们当记得这事，立定心意 。 叛逆的人哪，要留心思想。
ISA|46|9|要追念上古的事， 因为我是上帝，并无别的； 我是上帝，没有能与我相比的。
ISA|46|10|我从起初就指明末后的事， 从古时便言明未成的事， 说：“我的筹算必立定； 凡我所喜悦的，我必成就。”
ISA|46|11|我召鸷鸟从东方来， 召那成就我筹算的人从远方来。 我已说出，就必成就； 我已谋定，也必做成。
ISA|46|12|你们这些心中顽固、 远离公义的人，要听从我。
ISA|46|13|我使我的公义临近，它已不远。 我的救恩必不迟延。 我要为 以色列 －我的荣耀 在 锡安 施行救恩。
ISA|47|1|少女 巴比伦 哪， 下来坐在尘埃； 迦勒底 啊， 没有宝座，要坐在地上； 你不再称为柔弱娇嫩。
ISA|47|2|要用磨磨面， 揭去面纱， 脱去长裙， 露腿渡河。
ISA|47|3|你的下体必被露出； 你的羞辱必被看见。 我要报复， 谁也不宽容 。
ISA|47|4|我们的救赎主是 以色列 的圣者， 他的名为万军之耶和华。
ISA|47|5|迦勒底 啊， 你要静坐，进入黑暗中， 因你不再称为万国之后。
ISA|47|6|我向我的百姓发怒， 使我的产业受凌辱， 将他们交在你手中； 然而你毫不怜悯他们， 连老年人你也加极重的轭。
ISA|47|7|你说：“我必永远为后。” 你不将这事放在心上， 也不思想事情的结局。
ISA|47|8|你这专好宴乐、以为地位稳固的， 现在当听这话。 你心中说： “惟有我，除我以外再没有别的。 我必不致寡居， 也不经历丧子之痛。”
ISA|47|9|哪知，丧子、寡居这两件事 一日之间忽然临到你； 你虽多行邪术、广施魔咒， 这两件事必全然临到你身上。
ISA|47|10|你倚靠自己的恶行，说： “无人看见我。” 你的智慧聪明使你走偏， 你心里说： “惟有我，除我以外再没有别的了。”
ISA|47|11|但灾祸临到你， 你不知如何驱除； 灾害落在你身上， 你也无法除掉， 你所不知道的毁灭必忽然临到你身上。
ISA|47|12|尽管使用从幼年就施行的魔符和众多的邪术吧！ 或许有些帮助， 或许可以致胜。
ISA|47|13|你筹划太多，以致疲倦。 让那些观天象，看星宿， 在初一说预言的都起来， 救你脱离所要临到你的事！
ISA|47|14|看哪，他们要像碎秸被火焚烧， 无法救自己脱离火焰的魔掌； 没有炭火可以取暖 ， 你也不能坐在火旁。
ISA|47|15|你所操劳的事都像这样； 从你幼年以来与你交易的都各奔己路， 没有一人来救你。
ISA|48|1|雅各 家，称为 以色列 名下， 从 犹大 的源头而出的啊， 你们指着耶和华的名起誓， 提说 以色列 的上帝， 却不凭诚信，也不凭公义； 你们自称为圣城之民， 倚靠名为万军之耶和华－ 以色列 的上帝； 现在，当听我言：
ISA|48|2|
ISA|48|3|“先前的事，我自古已说明， 已从我口而出， 是我所指示的； 我瞬间行事，事便成就。
ISA|48|4|因为我知道你是顽梗的； 你的颈项是铁的， 你的额头是铜的。
ISA|48|5|所以，我自古就给你说明， 在事未成以先指示你， 免得你说：‘这些事是我的偶像所行的， 是我雕刻的偶像和铸造的神像所命定的。’
ISA|48|6|“你既已听见，现在要察看这一切； 你们不是要说明吗？ 从今以后，我要指示你新事， 就是你所不知道的隐密事。
ISA|48|7|这事是现今造的，并非自古就有， 在今日以先，你未曾听见； 免得你说：‘看哪，这事我早已知道了。’
ISA|48|8|诚然你未曾听见，也未曾知道； 你的耳朵从来未曾开通。 我原知道你行事极其诡诈， 你自从出母胎以来， 就称为悖逆的。
ISA|48|9|“我为我的名暂且忍怒， 为了我的荣耀向你容忍， 不将你剪除。
ISA|48|10|看哪，我熬炼你，却不像熬炼银子； 你在苦难的火炉中，我试炼 你。
ISA|48|11|我为自己的缘故必做这事， 我岂能被亵渎？ 我必不将我的荣耀归给别神 。
ISA|48|12|雅各 －我所选召的 以色列 啊， 当听从我： 我是耶和华， “我是首先的，也是末后的。
ISA|48|13|我亲手立了地的根基， 以右手铺张诸天； 我一召唤，天地就都立定。
ISA|48|14|你们都当聚集而听， 偶像 之中谁曾说明这些事？ 耶和华爱他，他必向 巴比伦 成就耶和华的旨意， 耶和华的膀臂也要加在 迦勒底 人身上 。
ISA|48|15|我，惟有我曾说过， 我选召他，领他来， 他的道路必亨通。
ISA|48|16|你们要接近我来听这话， 我从起初就未曾在隐密之处说话， 万事之始，我就在那里。” 现在，主耶和华差遣了我， 带着他的灵而来 。
ISA|48|17|耶和华－你的救赎主， 以色列 的圣者如此说： “我是耶和华－你的上帝， 我教导你，使你得益处， 指引你当走的路。
ISA|48|18|甚愿你听从我的命令， 你的平安就会如河水， 你的公义如海浪，
ISA|48|19|你的后裔必多如海沙， 你腹中所生的必多如沙粒。 他的名绝不从我面前剪除， 也不灭绝。”
ISA|48|20|你们要从 巴比伦 出来， 从 迦勒底 人中逃脱， 以欢呼的声音宣告， 将这事传扬到地极，说： 耶和华救赎了他的仆人 雅各 ！
ISA|48|21|他引导他们经过沙漠， 他们却未尝干渴； 他为他们使水从磐石流出， 磐石裂开，水就涌出。
ISA|48|22|耶和华说： “恶人必不得平安！”
ISA|49|1|众海岛啊，当听从我！ 远方的众民哪，要留心听！ 自出母胎，耶和华就选召我； 自出母腹，他就称呼我的名。
ISA|49|2|他使我的口如快刀， 把我藏在他手荫之下； 又使我成为磨利的箭， 把我藏在他箭袋之中；
ISA|49|3|对我说：“你是我的仆人 以色列 ； 我必因你得荣耀。”
ISA|49|4|我却说：“我劳碌是徒然， 我尽力是虚无虚空。 耶和华诚然以公平待我， 我的赏赐在我的上帝那里。”
ISA|49|5|现在耶和华说话，他从我出母胎，就造我作他的仆人， 要使 雅各 归向他， 使 以色列 聚集在他那里。 耶和华看我为尊贵， 我的上帝是我的力量。
ISA|49|6|他说：“你作我的仆人， 使 雅各 众支派复兴， 使 以色列 中蒙保存的人归回； 然而此事尚小， 我还要使你作万邦之光， 使你施行我的救恩，直到地极。”
ISA|49|7|救赎主－ 以色列 的圣者耶和华 对那被人藐视、本国憎恶、 统治者奴役的如此说： “君王看见就站起来， 领袖也要下拜； 这都是因信实的耶和华， 因拣选你的 以色列 的圣者。”
ISA|49|8|耶和华如此说： “在悦纳的时候，我应允了你； 在拯救的日子，我帮助了你。 我要保护你， 要藉着你与百姓立约， 为了复兴遍地， 使人承受荒芜之地为业；
ISA|49|9|对那被捆绑的人说：‘出来吧！’ 对在黑暗里的人说：‘显现吧！’ 他们在路上必得饮食， 在光秃的高地必有食物。
ISA|49|10|他们不饥不渴， 炎热和烈日必不伤害他们； 因为怜悯他们的必引导他们， 领他们到水泉旁边。
ISA|49|11|我必在众山开辟路径， 大道也要填高。
ISA|49|12|看哪，他们从远方来； 有些从北方来，有些从西方来， 有些从 色弗尼 地来。”
ISA|49|13|诸天哪，应当欢呼！ 大地啊，应当快乐！ 众山哪，应当扬声歌唱！ 因为耶和华已经安慰他的百姓， 他要怜悯他的困苦之民。
ISA|49|14|锡安 说：“耶和华离弃了我， 主忘记了我。”
ISA|49|15|妇人焉能忘记她吃奶的婴孩， 不怜悯她所生的儿子？ 即或有忘记的， 我却不忘记你。
ISA|49|16|看哪，我将你铭刻在我掌上， 你的城墙常在我眼前。
ISA|49|17|建立你的胜过毁坏你的， 使你荒废的必都离你而去。
ISA|49|18|你举目向四围观看， 他们都聚集来到你这里。 我指着我的永生起誓， 你定要以他们为妆饰佩戴， 带着他们，像新娘一样。 这是耶和华说的。
ISA|49|19|至于你荒废凄凉之处， 并你被毁坏之地， 如今居民必嫌太窄， 吞灭你的必离你遥远。
ISA|49|20|你要再听见丧失子女后所生的儿女说： “这地方我居住太窄， 请你给我地方居住。”
ISA|49|21|那时你心里必说：“我既丧子不育， 被掳，飘流在外 ， 谁给我生了这些？ 谁将他们养大呢？ 看哪，我被撇下独自一人时， 他们都在哪里呢？”
ISA|49|22|主耶和华如此说： “看哪，我必向列国举手， 向万民竖立大旗； 他们必将你的儿子抱在怀中带来， 将你的女儿背在肩上扛来。
ISA|49|23|列王必作你的养父， 王后必作你的乳母。 他们必以脸伏地，向你下拜， 并舔你脚上的尘土。 你就知道我是耶和华， 等候我的必不致羞愧。”
ISA|49|24|勇士抢去的岂能夺回？ 被残暴者掳掠的岂能得解救呢？
ISA|49|25|但耶和华如此说： “就是勇士所掳掠的，也可以夺回； 残暴者所抢的，也可以得解救。 与你相争的，我必与他相争， 我也要拯救你的儿女。
ISA|49|26|我必使那欺压你的吃自己的肉， 饮自己的血，如喝甜酒喝醉一样。 凡有血肉之躯的都必知道我－耶和华是你的救主， 是你的救赎主，是 雅各 的大能者。”
ISA|50|1|耶和华如此说： “我休了你们的母亲， 她的休书在哪里呢？ 我将你们卖给了我哪一个债主呢？ 看哪，你们被卖是因你们的罪孽； 你们的母亲被休，是因你们的过犯。
ISA|50|2|我来的时候，为何没有人呢？ 我呼唤的时候，为何无人回应呢？ 我的膀臂岂是过短、不能救赎吗？ 我岂无拯救之力吗？ 看哪，我一斥责，海就干了； 我使江河变为旷野， 其中的鱼因无水腥臭，干渴而死。
ISA|50|3|我使诸天以黑暗为衣， 以麻布为遮盖。”
ISA|50|4|主耶和华赐我受教者的舌头， 使我知道怎样用言语扶助疲乏的人。 主每天早晨唤醒，唤醒我的耳朵， 使我能听，像受教者一样。
ISA|50|5|主耶和华开启我的耳朵， 我并未违背，也未退后。
ISA|50|6|人打我的背，我任他打； 人拔我两颊的胡须，我由他拔； 人侮辱我，向我吐唾沫，我并不掩面。
ISA|50|7|主耶和华必帮助我， 所以我不抱愧。 我硬着脸面好像坚石， 也知道我必不致蒙羞。
ISA|50|8|称我为义的与我相近； 谁与我争论， 让我们来对质； 谁与我作对， 让他近前来吧！
ISA|50|9|看哪，主耶和华必帮助我， 谁能定我有罪呢？ 看哪，他们都要像衣服渐渐破旧， 被蛀虫蛀光。
ISA|50|10|你们当中有谁是敬畏耶和华， 听从他仆人的话语， 却行在黑暗中，没有亮光的， 当倚靠耶和华的名， 仰赖自己的上帝。
ISA|50|11|看哪，你们当中所有点火、以火把围绕自己的人， 当行走在你们的火焰 里， 并你们所点的火把中。 这是我亲手为你们定的： 你们必躺卧在悲惨之中。
ISA|51|1|追求公义、 寻求耶和华的人哪， 当听从我！ 你们要追想自己是从哪块磐石凿出， 从哪个岩穴挖掘而来；
ISA|51|2|要追想你们的祖宗 亚伯拉罕 和生你们的 撒拉 ； 因为我选召 亚伯拉罕 时，他只有一个人， 但我赐福给他， 使他增多。
ISA|51|3|耶和华已经安慰 锡安 ， 安慰了 锡安 一切的废墟， 使旷野如 伊甸 ， 使沙漠像耶和华的园子； 其中必有欢喜、快乐、感谢， 和歌唱的声音。
ISA|51|4|我的民哪，要留心听我， 我的国啊，要向我侧耳； 因为训诲必从我而出， 我必使我的公理成为万民之光。
ISA|51|5|我的公义临近， 我的救恩发出。 我的膀臂要审判万民， 众海岛都要等候我，倚赖我的膀臂。
ISA|51|6|你们要向天举目， 观看下面的地； 天必像烟云消散， 地必如衣服渐渐破旧； 其上的居民也要如此 死亡。 惟有我的救恩永远长存， 我的公义也不废掉。
ISA|51|7|知道公义、将我的训诲存在心中的人哪， 当听从我！ 不要怕人的辱骂， 也不要因人的毁谤惊惶。
ISA|51|8|因为他们必像衣服被蛀虫蛀； 像羊毛被虫子咬。 惟有我的公义永远长存， 我的救恩直到万代。
ISA|51|9|耶和华的膀臂啊，兴起，兴起！ 以能力为衣穿上， 像古时的年日，像上古的世代一样兴起！ 从前砍碎 拉哈伯 、 刺透大鱼的，不是你吗？
ISA|51|10|使海与深渊的水干涸， 在海的深处开路， 使救赎的民走过的，不是你吗？
ISA|51|11|耶和华救赎的民必归回， 歌唱来到 锡安 ； 永恒的喜乐必归到他们头上。 他们必得着欢喜快乐， 忧伤叹息尽都逃避。
ISA|51|12|我，惟有我是安慰你们的。 你是谁，竟怕那必死的人， 怕那生命如草的世人，
ISA|51|13|却忘记铺张诸天、立定地基、 造你的耶和华？ 你因欺压者图谋毁灭所发的暴怒， 终日害怕， 其实那欺压者的暴怒在哪里呢？
ISA|51|14|被掳的即将得释放， 不至于死而下入地府， 也不致缺乏食物。
ISA|51|15|我是耶和华－你的上帝， 我搅动大海，使海中的波浪澎湃， 万军之耶和华是我的名。
ISA|51|16|我已将我的话放在你口中， 用我的手影遮蔽你， 为要安定诸天，立定地基， 并对 锡安 说：“你是我的百姓。”
ISA|51|17|耶路撒冷 啊，兴起，兴起！ 站起来！ 你从耶和华手中喝了他愤怒的杯， 那使人东倒西歪的杯，直到喝尽。
ISA|51|18|她所生育的孩子中，没有一个搀她的； 她所抚养的孩子中，没有一个扶她的。
ISA|51|19|这双重的灾难临到你， 有谁怜悯你呢？ 破坏和毁灭，饥荒和战争临到， 我如何能安慰你呢 ？
ISA|51|20|你的孩子发昏， 在各街头躺卧， 如同网罗里的羚羊， 满了耶和华的愤怒， 满了你上帝的斥责。
ISA|51|21|因此，你这困苦却非因酒而醉的， 当听这话，
ISA|51|22|你的主，耶和华， 就是为他百姓辩护的上帝如此说： “看哪，我已从你手中接过 那使人东倒西歪的杯， 就是我愤怒的杯， 你必不再喝。
ISA|51|23|我必将这杯递在苦待你的人 手中。 他们曾对你说：‘你屈身， 任我们践踏过去吧！’ 你就以背为地， 又如街道，任人走过。
ISA|52|1|锡安 哪，兴起！兴起！ 穿上你的能力！ 圣城 耶路撒冷 啊，穿上你华美的衣服！ 因为从今以后， 未受割礼、不洁净的必不再进入你中间。
ISA|52|2|耶路撒冷 啊，抖去尘埃， 起来坐在王位上！ 被掳的 锡安 哪， 解开你颈上的锁链！
ISA|52|3|耶和华如此说：“你们白白地被卖，也必不用银子赎回。”
ISA|52|4|主耶和华如此说：“先前我的百姓下到 埃及 ，在那里寄居，末后又有 亚述 人欺压他们。”
ISA|52|5|我的百姓既是白白地被掳，如今我在这里做什么呢？这是耶和华说的。辖制他们的人欢呼 ，我的名终日不断受亵渎，这是耶和华说的。
ISA|52|6|因此，我的百姓必认识我的名；在那日，他们必知道说这话的就是我。看哪，是我！”
ISA|52|7|在山上报佳音，传平安， 报好信息，传扬救恩， 那人的脚踪何等佳美啊！ 他对 锡安 说：“你的上帝作王了！”
ISA|52|8|听啊，你守望之人的声音， 他们扬声一同欢唱； 因为他们必亲眼看见耶和华返回 锡安 。
ISA|52|9|耶路撒冷 的废墟啊， 要出声一同欢唱； 因为耶和华安慰了他的百姓， 救赎了 耶路撒冷 。
ISA|52|10|耶和华在万国眼前露出圣臂， 地的四极都要看见我们上帝的救恩。
ISA|52|11|离开吧！离开吧！ 你们要从 巴比伦 出来。 你们扛抬耶和华器皿的人哪， 不要沾不洁净的东西， 离去时务要保持洁净。
ISA|52|12|你们出来必不致匆忙， 也不致奔逃； 因为耶和华要在你们前头行， 以色列 的上帝必作你们的后盾。
ISA|52|13|看哪，我的仆人行事必有智慧， 他必被高升，高举， 升到至高之处。
ISA|52|14|许多人因他 惊奇 ─他的面貌比别人憔悴， 他的外表比世人枯槁─
ISA|52|15|同样，他也必使许多国家惊奇 ， 君王要向他闭口。 未曾传给他们的，他们必看见； 未曾听见过的事，他们要明白。
ISA|53|1|我们所传的有谁信呢？ 耶和华的膀臂向谁显露呢？
ISA|53|2|他在耶和华面前生长如嫩芽， 像根出于干地。 他无佳形美容使我们注视他， 也无美貌使我们仰慕他。
ISA|53|3|他被藐视，被人厌弃； 多受痛苦，常经忧患。 他被藐视， 好像被人掩面不看的一样， 我们也不尊重他。
ISA|53|4|他诚然担当我们的忧患， 背负我们的痛苦； 我们却以为他受责罚， 是被上帝击打苦待。
ISA|53|5|他为我们的过犯受害， 为我们的罪孽被压伤。 因他受的惩罚，我们得平安； 因他受的鞭伤，我们得医治。
ISA|53|6|我们都如羊走迷， 各人偏行己路； 耶和华使我们众人的罪孽都归在他身上。
ISA|53|7|他被欺压受苦， 却不开口； 他像羔羊被牵去宰杀， 又像羊在剪毛的人手下无声， 他也是这样不开口。
ISA|53|8|因受欺压和审判，他被夺去， 谁能想到他的世代呢？ 因为他从活人之地被剪除， 为我百姓 的罪过他被带到死里 。
ISA|53|9|他虽然未行残暴， 口中也没有诡诈， 人还使他与恶人同穴， 与财主同墓 。
ISA|53|10|耶和华的旨意要压伤他， 使他受苦。 当他的生命作为赎罪祭时 ， 他必看见后裔，他的年日必然长久。 耶和华所喜悦的事，必在他手中亨通。
ISA|53|11|因自己的劳苦，他必看见光 就心满意足。 因自己的认识，我的义仆使许多人得称为义， 他要担当他们的罪孽。
ISA|53|12|因此，我要使他与位大的同份， 与强盛的均分掳物。 因为他倾倒自己的生命，以致于死， 也列在罪犯之中。 他却担当多人的罪， 为他们的过犯代求 。
ISA|54|1|你这不怀孕、不生育的，要欢呼； 你这未曾经过产难的，要欢呼，扬声呼喊； 因为被遗弃的妇人， 比有丈夫的人儿女更多； 这是耶和华说的。
ISA|54|2|要扩张你帐幕之地， 伸展你居所的幔子，不要缩回； 要放长你的绳子， 坚固你的橛子。
ISA|54|3|因为你要向左向右开展， 你的后裔必得列国为业， 又使荒废的城镇有人居住。
ISA|54|4|不要惧怕，因你必不致蒙羞； 不要抱愧，因你必不致受辱。 你必忘记年轻时的羞愧， 不再记得守寡的耻辱。
ISA|54|5|因为造你的是你的丈夫， 万军之耶和华是他的名； 救赎你的是 以色列 的圣者， 他必称为全地之上帝。
ISA|54|6|耶和华召你， 如同召回心中忧伤遭遗弃的妇人， 就是年轻时所娶被遗弃的妻子； 这是你的上帝说的。
ISA|54|7|我离弃你不过片时， 却要大施怜悯将你寻回。
ISA|54|8|我因涨溢的怒气， 一时向你转脸， 但我要以永远的慈爱怜悯你； 这是耶和华－你的救赎主说的。
ISA|54|9|这事于我有如 挪亚 的洪水； 我怎样起誓不再使 挪亚 的洪水淹没全地， 也照样起誓不再向你发怒， 且不斥责你。
ISA|54|10|大山可以挪开， 小山可以迁移， 但我的慈爱必不离开你， 我平安的约也不迁移； 这是怜悯你的耶和华说的。
ISA|54|11|你这受困苦、被暴风卷走、不得怜悯的城， 看哪，我必以灰泥来做你的石头， 以蓝宝石立你的根基，
ISA|54|12|又以红宝石造你的女墙， 以晶莹的珠玉造你的城门， 以珍贵的宝石造你四围的边界。
ISA|54|13|你的儿女都要领受耶和华的教导， 你的儿女必大享平安。
ISA|54|14|你必因公义得坚立， 必远离欺压，毫不惧怕； 你必远离惊吓，惊吓必不临近你。
ISA|54|15|若有人攻击你，这非出于我； 凡攻击你的，必因你仆倒。
ISA|54|16|看哪，我造了那吹炭火、打造合用兵器的铁匠； 我也造了那残害人、行毁灭的人。
ISA|54|17|凡为攻击你而造的兵器必无效用； 在审判时兴起用口舌攻击你的， 你必驳倒他。 这是耶和华仆人的产业， 是他们从我所得的义； 这是耶和华说的。
ISA|55|1|来！你们所有干渴的，都当来到水边； 没有银钱的也可以来。 你们都来，买了吃； 不用银钱，不付代价， 就可买酒和奶。
ISA|55|2|你们为何花钱买那不是食物的东西， 用劳碌得来的买那无法使人饱足的呢？ 你们要留意听从我的话，就能吃那美物， 得享肥甘，心中喜乐。
ISA|55|3|当侧耳而听，来到我这里； 要听，就必存活。 我要与你们立永约， 就是应许给 大卫 那可靠的慈爱。
ISA|55|4|看哪，我已立他作万民的见证， 立他作万民的君王和发令者。
ISA|55|5|看哪，你要召集素不认识的国民， 素不认识的国民要奔向你； 这都因耶和华─你的上帝， 因 以色列 的圣者已经荣耀了你。
ISA|55|6|当趁耶和华可寻找的时候寻找他， 在他接近的时候求告他。
ISA|55|7|恶人当离弃自己的道路， 不义的人应除掉自己的意念。 归向耶和华，耶和华就必怜悯他； 当归向我们的上帝，因为他必广行赦免。
ISA|55|8|我的意念非同你们的意念， 我的道路非同你们的道路。 这是耶和华说的。
ISA|55|9|天怎样高过地， 照样，我的道路高过你们的道路， 我的意念高过你们的意念。
ISA|55|10|雨雪从天而降，并不返回， 却要滋润土地，使地面发芽结实， 使撒种的有种，使要吃的有粮。
ISA|55|11|我口所出的话也必如此， 绝不徒然返回， 却要成就我的旨意， 达成我差它的目的。
ISA|55|12|你们必欢欢喜喜出来， 平平安安蒙引导。 大山小山必在你们面前欢呼， 田野的树木也都拍掌。
ISA|55|13|松树长出，代替荆棘； 番石榴长出，代替蒺藜。 这要为耶和华留名， 作为永不磨灭的证据。
ISA|56|1|耶和华如此说： “你们当守公平，行公义； 因我的救恩临近， 我的公义将要显现。
ISA|56|2|谨守安息日不予干犯， 禁止己手不作恶， 如此行、如此持守的人有福了！”
ISA|56|3|与耶和华联合的外邦人不要说： “耶和华将我和他的子民分别出来。” 太监也不要说：“看哪，我是枯树。”
ISA|56|4|因为耶和华如此说： “那些谨守我的安息日， 选择我旨意， 持守我约的太监，
ISA|56|5|我必使他们在我殿中，在我墙内， 有纪念碑，有名号， 胜过有儿有女； 我必赐他们永远的名，不能剪除。
ISA|56|6|“那些与耶和华联合， 事奉他，爱他名， 作他仆人的外邦人， 凡谨守安息日不予干犯， 又持守我约的人，
ISA|56|7|我必领他们到我的圣山， 使他们在我的祷告的殿中喜乐。 他们的燔祭和祭物， 在我坛上必蒙悦纳， 因我的殿必称为万民祷告的殿。
ISA|56|8|我还要召集更多的人 归并到这些被召集的人中。 这是召集被赶散的 以色列 人的 主耶和华说的。”
ISA|56|9|野地的走兽，你们都来吞吃吧！ 林中的野兽，你们也来吞吃！
ISA|56|10|以色列 的守望者都瞎了眼， 没有知识； 都是哑狗，不会吠叫， 只知做梦，躺卧，贪睡，
ISA|56|11|这些狗贪食，不知饱足。 这些牧人不知明辨， 他们都偏行己路， 人人追求自己的利益。
ISA|56|12|他们说：“来吧！我去拿酒， 让我们畅饮烈酒吧！ 明天必和今天一样， 甚至更好！”
ISA|57|1|义人死亡， 无人放在心上； 虔诚的人被接去， 无人理解； 义人被接去，以免祸患。
ISA|57|2|行为正直的人进入平安， 得以在床上安歇 。
ISA|57|3|到这里来吧！ 你们这些巫婆的儿子， 奸夫和妓女的后代；
ISA|57|4|你们向谁戏笑？ 向谁张口吐舌呢？ 你们岂不是叛逆所生的儿女， 虚谎所生的后代吗？
ISA|57|5|你们在橡树 中间，在各青翠的树下欲火攻心； 在山谷间，在岩隙下杀了儿女；
ISA|57|6|去拜谷中光滑的石头有你们的份， 这些就是你们的命运。 你向它们献浇酒祭，献供物， 这事我岂能容忍吗？
ISA|57|7|你在高而又高的山上安设床铺， 上那里去献祭。
ISA|57|8|你在门后，在门框后， 立起你的牌来； 你离弃了我，赤露己身， 又爬上自己所铺宽阔的床铺， 与它们立约； 你喜爱它们的床，看着它们的赤体 。
ISA|57|9|你带了油到 摩洛 那里， 加上许多香水。 你派遣使者往远方去， 甚至降到阴间，
ISA|57|10|因路途遥远，你就疲倦， 却不说，这是枉然， 以为能找到复兴之力， 所以不觉疲惫。
ISA|57|11|你怕谁，因谁恐惧， 竟说谎，不记得我， 不将这事放在心上。 是否因我许久闭口不言， 你就不怕我了呢？
ISA|57|12|我可以宣告你的公义和你的作为， 但它们与你无益。
ISA|57|13|你哀求的时候， 让你所搜集的神像 拯救你吧！ 风要把它们全都刮散， 吹一口气就都吹走。 但那投靠我的必得地产， 承受我的圣山为业。
ISA|57|14|耶和华说： “你们要修筑，修筑，要预备道路， 除掉我百姓路中的绊脚石。”
ISA|57|15|那至高无上、永远长存、 名为圣者的如此说： “我住在至高至圣的所在， 却与心灵痛悔的谦卑人同住； 要使谦卑的人心灵苏醒， 使痛悔的人内心复苏。
ISA|57|16|我必不长久控诉，也不永远怀怒， 因为我虽使灵性发昏，我也造了人的气息。
ISA|57|17|我因人贪婪的罪孽，发怒击打他； 我转脸向他发怒， 他却仍随意背道而行。
ISA|57|18|我看见他的行为， 要医治他，引导他 ， 使他和与他一同哀伤的人都得安慰。
ISA|57|19|我要医治他， 他要结出嘴唇的果实。 平安，平安，归给远处和近处的人！ 这是耶和华说的。”
ISA|57|20|但是恶人好像翻腾的海， 不得平静； 其中的水常涌出污秽和淤泥。
ISA|57|21|我的上帝说：“恶人必不得平安！”
ISA|58|1|你要大声喊叫，不要停止； 要扬声，好像吹角； 向我的百姓宣告他们的过犯， 向 雅各 家陈述他们的罪恶。
ISA|58|2|他们天天寻求我， 乐意明白我的道， 好像行义的国家， 未离弃它的上帝的典章； 他们向我求问公义的判词， 喜悦亲近上帝。
ISA|58|3|“我们禁食，你为何不看呢？ 我们刻苦己心，你为何不理会呢？” 看哪，你们禁食的时候仍追求私利， 剥削为你们做苦工的人。
ISA|58|4|看哪，你们禁食，却起纷争兴讼， 以凶恶的拳头打人。 你们今日这种禁食 无法使你们的声音听闻于高处。
ISA|58|5|这岂是我所要的禁食， 为人所用以刻苦己心的日子吗？ 我难道只是叫人如芦苇般低头， 铺上麻布和灰烬吗？ 你能称此为禁食， 为耶和华所悦纳的日子吗？
ISA|58|6|我所要的禁食，岂不是要你松开凶恶的绳， 解开轭上的索， 使被欺压的得自由， 折断一切的轭吗？
ISA|58|7|岂不是要你把食物分给饥饿的人， 将流浪的穷人接到家中， 见赤身的给他衣服遮体， 而不隐藏自己避开你的骨肉吗？
ISA|58|8|这样，必有光如晨光破晓照耀你， 你也要快快得到医治； 你的公义在你前面行， 耶和华的荣光必作你的后盾。
ISA|58|9|那时你求告，耶和华必应允； 你呼求，他必说：“我在这里。” 你若从你中间除掉重轭 和指摘人的指头，并发恶言的事，
ISA|58|10|向饥饿的人施怜悯， 使困苦的人得满足； 你在黑暗中就必得着光明， 你的幽暗必变如正午。
ISA|58|11|耶和华必时常引导你， 在干旱之地使你心满意足， 又使你骨头强壮。 你必如有水浇灌的园子， 又像水流不绝的泉源。
ISA|58|12|你们中间必有人起来修造久已荒废之处， 立起代代相承的根基。 你必称为修补裂痕的， 和重修路径给人居住的。
ISA|58|13|你若禁止自己的脚践踏安息日， 不在我的圣日做自己高兴的事， 称安息日为“可喜乐的”， 称耶和华的圣日为“可尊重的”， 尊敬这日， 不走自己的道路， 不求自己的喜悦， 也不随意说话；
ISA|58|14|那么，你就会以耶和华为乐。 耶和华要使你乘驾于地的高处， 又要以你祖先 雅各 的产业养育你； 这是耶和华亲口说的。
ISA|59|1|看哪，耶和华的膀臂并非过短，不能拯救， 耳朵并非发沉，不能听见，
ISA|59|2|但你们的罪孽使你们与上帝隔绝， 你们的罪恶使他转脸不听你们。
ISA|59|3|因你们的手掌被血沾染， 你们的指头被罪玷污， 你们的嘴唇说谎言， 你们的舌头出恶语。
ISA|59|4|无人按公义控诉， 也无人凭诚实辩白； 却倚靠虚妄，口说谎言， 怀毒害，生罪孽。
ISA|59|5|他们孵毒蛇蛋， 结蜘蛛网。 凡吃这蛋的必死， 蛋一打破，就孵出蛇来。
ISA|59|6|所结的网不能当衣服， 无法掩盖自己所作所为。 他们的行为全是邪恶， 手所做的尽都残暴。
ISA|59|7|他们的脚奔跑行恶， 急速流无辜者的血； 他们的思想全是恶念， 走过的路尽是破坏与毁灭。
ISA|59|8|平安的路，他们不知道， 所行的事无一公平。 他们为自己修筑弯曲的路， 凡走这路的都不得平安。
ISA|59|9|因此，公平离我们甚远， 公义追不上我们。 我们指望光亮，看哪，却只有黑暗， 指望光明，却行在幽暗中。
ISA|59|10|我们用手摸墙，好像盲人， 四处摸索，如同失明的人； 中午时我们绊倒，如在黄昏一样， 在强壮的人中，我们好像死人一般。
ISA|59|11|我们全都咆哮如熊， 哀鸣如鸽子； 指望公平，却得不着； 指望救恩，它却远离。
ISA|59|12|我们的过犯在你面前增加， 罪恶作证控告我们； 过犯与我们同在。 至于我们的罪孽，我们都知道：
ISA|59|13|就是悖逆，否认耶和华， 转去不跟从我们的上帝， 口说欺压和叛逆的话， 心怀谎言，随即说出；
ISA|59|14|公平转而退后， 公义站在远处， 诚实仆倒在广场上， 正直不得进入；
ISA|59|15|诚实少见， 离弃邪恶的人反成掠物。 那时，耶和华见没有公平， 就不喜悦。
ISA|59|16|他见无人， 竟无一人代求，甚为诧异， 就用自己的膀臂拯救他， 以公义扶持他。
ISA|59|17|他穿上公义为铠甲， 戴上救恩为头盔， 穿上报复为衣服， 披戴热心为外袍。
ISA|59|18|他必按人的行为报应， 恼怒他的敌人， 报复他的仇敌， 向众海岛施行报应。
ISA|59|19|在日落之处，人必敬畏耶和华的名； 在日出之地，人必敬畏他的荣耀。 他必如湍急的河流冲来， 耶和华的灵催逼他自己。
ISA|59|20|必有一位救赎主来到 锡安 ， 来到 雅各 族中离弃过犯的人那里； 这是耶和华说的。
ISA|59|21|耶和华说：“这就是我与他们所立的约：我加给你的灵，传给你的话，必不离你的口，也不离你后裔与你后裔之后裔的口，从今直到永远；这是耶和华说的。”
ISA|60|1|兴起，发光！因为你的光已来到！ 耶和华的荣光发出照耀着你。
ISA|60|2|看哪，黑暗笼罩大地， 幽暗遮盖万民， 耶和华却要升起照耀你， 他的荣光要显在你身上。
ISA|60|3|列国要来就你的光， 列王要来就你发出的光辉。
ISA|60|4|你举目向四围观看， 众人都聚集到你这里。 你的儿子从远方来， 你的女儿也被抱着带来。
ISA|60|5|那时，你看见就有光荣， 你的心兴奋欢畅 ； 因为大海那边的财富必归你， 列国的财宝也来归你。
ISA|60|6|成群的骆驼， 并 米甸 和 以法 的独峰驼遮满你； 示巴 的众人都必来到， 要奉上黄金和乳香， 又要传扬赞美耶和华的话。
ISA|60|7|基达 的羊群都聚集到你这里， 尼拜约 的公羊供你使用， 献在我坛上蒙悦纳； 我必荣耀我那荣耀的殿。
ISA|60|8|那些飞来如云、 又像鸽子飞向窗户的是谁呢？
ISA|60|9|众海岛必等候我 ， 他施 的船只领先， 将你的儿女，连同他们的金银从远方带来， 这都因 以色列 的圣者、耶和华－你上帝的名， 因为他已经荣耀了你。
ISA|60|10|外邦人要建造你的城墙， 他们的君王必服事你。 我曾发怒击打你， 如今却施恩怜悯你。
ISA|60|11|你的城门必时常开放， 昼夜不关， 使人将列国的财物带来归你， 他们的君王也被牵引而来。
ISA|60|12|不事奉你的那邦、那国要灭亡， 那些国家必全然荒废。
ISA|60|13|黎巴嫩 的荣耀， 就是松树、杉树、黄杨树， 都必一同归你， 用以装饰我圣所坐落之处； 我也要使我脚所踏之地得荣耀。
ISA|60|14|压制你的，他的子孙必来向你屈身； 藐视你的，都要在你脚前下拜。 人要称你为“耶和华的城”， 为“ 以色列 圣者的 锡安 ”。
ISA|60|15|你虽曾被抛弃，被恨恶， 甚至无人经过， 我却使你有永远的荣华， 成为世世代代的喜乐。
ISA|60|16|你要吃列国的奶， 吃列王的乳。 你就知道我－耶和华是你的救主， 是你的救赎主，是 雅各 的大能者。
ISA|60|17|我要赏赐金子代替铜， 赏赐银子代替铁， 铜代替木头， 铁代替石头。 我要以和平为你的官长， 以公义为你的监督。
ISA|60|18|你的地不再听闻残暴的事， 境内不再听见破坏与毁灭。 你必称你的墙为“拯救”， 称你的门为“赞美”。
ISA|60|19|白昼太阳不再作你的光， 月亮 也不再发光照耀你； 耶和华却要作你永远的光， 你的上帝要成为你的荣耀。
ISA|60|20|你的太阳不再落下， 月亮也不消失； 因为耶和华必作你永远的光。 你悲哀的日子定要结束。
ISA|60|21|你的居民全是义人， 永远得地为业； 他们是我栽的苗，是我手的工作， 为了彰显我的荣耀。
ISA|60|22|稀少的要成为大族， 弱小的要变为强国。 我－耶和华到了时候必速速成就这事。
ISA|61|1|主耶和华的灵在我身上， 因为耶和华用膏膏我， 叫我报好信息给贫穷的人， 差遣我医好伤心的人， 报告被掳的得释放， 被捆绑的得自由；
ISA|61|2|宣告耶和华的恩年 和我们的上帝报仇的日子； 安慰所有悲哀的人，
ISA|61|3|为 锡安 悲哀的人，赐华冠代替灰烬， 喜乐的油代替悲哀， 赞美为衣代替忧伤的灵； 称他们为“公义树”， 是耶和华所栽植的，为要彰显他的荣耀。
ISA|61|4|他们必修造久已荒凉的废墟， 建立先前凄凉之处， 重修历代荒凉之城。
ISA|61|5|那时，陌生人要伺候、牧放你们的羊群； 外邦人必为你们耕种田地， 修整你们的葡萄园。
ISA|61|6|但你们要称为“耶和华的祭司”， 称作“我们上帝的仆人”。 你们必享用列国的财物， 必承受他们的财富 。
ISA|61|7|因为他们所受双倍的羞辱， 凌辱被称为他们的命运， 因此，他们在境内必得双倍的产业， 永远之乐必归给他们。
ISA|61|8|因为我－耶和华喜爱公平， 恨恶抢夺与恶行 ； 我要凭诚实施行报偿， 与我的百姓立永约。
ISA|61|9|他们的后裔必在列国中为人所知， 他们的子孙在万民中为人所识； 凡看见他们的必承认他们是耶和华所赐福的后裔。
ISA|61|10|我因耶和华大大欢喜， 我的心因上帝喜乐； 因他以拯救为衣给我穿上， 以公义为外袍给我披上， 好像新郎戴上华冠， 又如新娘佩戴首饰。
ISA|61|11|地怎样使芽长出， 园子怎样使所栽种的生长， 主耶和华也必照样 使公义和赞美在万国中发出。
ISA|62|1|我因 锡安 必不静默， 为 耶路撒冷 必不安宁， 直到它的公义如光辉发出， 它的救恩如火把燃烧。
ISA|62|2|列国要看见你的公义， 列王要看见你的荣耀。 你必得新的名字， 是耶和华亲口起的。
ISA|62|3|你在耶和华的手中成为华冠， 在你上帝的掌上成为冠冕。
ISA|62|4|你不再称为“被撇弃的”， 你的地也不再称为“荒芜的”； 你要称为“我所喜悦的”， 你的地要称为“有归属的”。 因为耶和华喜悦你， 你的地必归属于他。
ISA|62|5|年轻人怎样娶童女， 你的百姓也要照样娶你； 新郎怎样因新娘而喜乐， 你的上帝也要如此以你为乐。
ISA|62|6|耶路撒冷 啊， 我在你城墙上设立守望者， 他们昼夜不停地呼喊。 呼求耶和华的啊，你们不要歇息，
ISA|62|7|也不要使他歇息， 直等他建立 耶路撒冷 ， 使 耶路撒冷 在地上为人所赞美。
ISA|62|8|耶和华指着自己的右手和大能的膀臂起誓说： “我必不再将你的五谷给仇敌作食物， 外邦人也必不再喝你劳碌得来的新酒。
ISA|62|9|惟有那收割的要吃，并赞美耶和华； 那储藏葡萄的要在我圣所院内喝。”
ISA|62|10|你们当从门经过，经过， 预备百姓的路。 你们要修筑，修筑大道， 清除石头， 为万民竖立大旗。
ISA|62|11|看哪，耶和华曾宣告到地极， 你们要对 锡安 说： “看哪，你的拯救者已来到。 看哪，他的赏赐在他那里， 他的报偿在他面前。”
ISA|62|12|人称他们为“圣民”，为“耶和华救赎的民”， 你也必称为“受眷顾的”，为“不被撇弃的城”。
ISA|63|1|这从 以东 的 波斯拉 来， 穿红衣服， 装扮华美， 能力广大， 大步向前迈进的是谁呢？ 就是我， 凭公义说话， 以大能施行拯救的。
ISA|63|2|你为何以红色装扮？ 你的衣服为何像踹醡酒池的人呢？
ISA|63|3|我独自踹醡酒池， 万民中并无一人与我同在。 我发怒，将他们踹下， 发烈怒将他们践踏。 他们的血溅在我的衣服上， 玷污了我一切的衣裳。
ISA|63|4|因为报仇之日在我心中， 救赎我民之年已经来到。
ISA|63|5|我仰望，见无人帮助； 我诧异，竟无人扶持。 因此，我的膀臂为我施行拯救； 我的烈怒将我扶持。
ISA|63|6|我发怒，踹下众民； 发烈怒，使他们喝醉， 又将他们的血倒在地上。
ISA|63|7|我要照耶和华一切所赐给我们的， 并他凭怜悯与丰盛的慈爱 所赐给 以色列 家的大恩， 述说他的慈爱和美德。
ISA|63|8|他说：“他们诚然是我的百姓， 未行虚假的子民。” 这样，他就作了他们的救主。
ISA|63|9|他们在一切苦难当中， 他也同受苦难， 并且他面前的使者拯救他们 。 他以慈爱和怜悯救赎他们， 在古时的日子时常抱他们，背他们。
ISA|63|10|他们竟然悖逆，使他的圣灵忧伤。 他就转变，成为他们的仇敌， 亲自攻击他们。
ISA|63|11|那时，他的百姓想起古时 摩西 的日子： “那将百姓和牧养群羊的人 从海里领上来的在哪里呢？ 那将圣灵降在他们中间，
ISA|63|12|以荣耀的膀臂在 摩西 右边行动， 在百姓面前将水分开， 为要建立自己永远的名，
ISA|63|13|又带领他们经过深处的在哪里呢？” 他们如马行走旷野，不致绊跌；
ISA|63|14|又如牲畜下到山谷， 耶和华的灵使他们得安息； 照样，你也引导你的百姓， 为要建立自己荣耀的名。
ISA|63|15|求你从天上， 从你神圣荣耀的居所垂顾观看。 你的热心和你大能的作为在哪里呢？ 你内心的关怀和你的怜悯向我们停止了。
ISA|63|16|亚伯拉罕 虽然不承认我们， 以色列 也不承认我们， 你却是我们的父。 耶和华啊，你是我们的父； 自古以来，你的名是“我们的救赎主”。
ISA|63|17|耶和华啊，你为何使我们偏离你的道， 使我们心里刚硬、不敬畏你呢？ 求你为你的仆人， 为你产业的支派而回转。
ISA|63|18|你的圣民暂时得你的圣所， 但我们的敌人践踏了它。
ISA|63|19|我们就成了你未曾治理的人， 成了未曾称为你名下的人。
ISA|64|1|愿你破天而降， 愿山在你面前震动，
ISA|64|2|好像火烧干柴， 又如火将水烧开， 使你敌人知道你的名， 列国必在你面前发颤！
ISA|64|3|你曾做我们不能逆料可畏的事； 那时你降临，山岭在你面前震动。
ISA|64|4|自古以来，人未曾听见，未曾耳闻，未曾眼见， 除你以外，还有上帝能为等候他的人行事。
ISA|64|5|你迎见那欢喜行义、记念你道的人； 看哪，你曾发怒，因我们犯了罪； 这景况已久，我们还能得救吗？
ISA|64|6|我们都如不洁净的人， 所行的义都像污秽的衣服。 我们如叶子渐渐枯干， 罪孽像风把我们吹走。
ISA|64|7|无人求告你的名， 无人奋力抓住你。 你转脸不顾我们， 你使我们因罪孽而融化 。
ISA|64|8|但耶和华啊，现在你仍是我们的父！ 我们是泥，你是陶匠； 我们都是你亲手所造的。
ISA|64|9|耶和华啊，求你不要大发震怒， 也不要永远记得罪孽； 看哪，求你垂顾我们， 因我们都是你的百姓。
ISA|64|10|你的圣城已变为旷野； 锡安 变为旷野， 耶路撒冷 成为废墟。
ISA|64|11|我们那神圣华美的殿， 就是我们祖先赞美你的地方，已被火焚烧； 我们所羡慕的美地尽都荒芜。
ISA|64|12|耶和华啊，有这些事，你还能忍受吗？ 你还静默，使我们大受苦难吗？
ISA|65|1|没有求问我的，我要让他们找到； 没有寻找我的，我要让他们寻见； 我对没有呼求我名的国 说： “我在这里！我在这里！”
ISA|65|2|我整天向那悖逆的百姓招手， 他们随自己的意念行不善之道。
ISA|65|3|这百姓时常当面惹我发怒， 在园中献祭， 在砖上烧香，
ISA|65|4|在坟墓间停留， 在隐密处过夜， 吃猪肉， 器皿中有不洁净之肉熬的汤；
ISA|65|5|且对人说：“你站开吧！ 不要挨近我，因为我对你来说太神圣了 。” 这些人惹我鼻中冒烟， 如终日燃烧的火。
ISA|65|6|看哪，这些都写在我面前。 我必不静默，却要施行报应， 将你们和你们祖先的罪孽 全都报应在后人身上； 因为他们在山上烧香， 在冈上亵渎我， 我要按他们先前所行的，报应在他们身上 ； 这是耶和华说的。
ISA|65|7|
ISA|65|8|耶和华如此说： “人在葡萄中寻得新酒时会说： ‘不要毁坏它，因为它还有用处’； 同样，我必因我仆人的缘故， 不将他们全然毁灭。
ISA|65|9|我必从 雅各 中领出后裔， 从 犹大 中领出那要继承我众山的； 我的选民要继承它， 我的仆人要在那里居住。
ISA|65|10|沙仑 必成为羊群的圈， 亚割谷 成为牛群躺卧之处， 都为寻求我的民所得。
ISA|65|11|但你们这些离弃耶和华， 就是忘记我的圣山、 为‘幸运之神’摆设筵席、 为‘命运之神’装满调和酒的，
ISA|65|12|我命定你们归于刀下， 你们都要屈身被杀； 因为我呼唤，你们不回应； 我说话，你们不听从； 反倒做我眼中看为恶的事， 选择我所不喜悦的事。”
ISA|65|13|所以，主耶和华如此说： “看哪，我的仆人必得吃，你们却饥饿； 看哪，我的仆人必得喝，你们却干渴； 看哪，我的仆人必欢喜，你们却蒙羞。
ISA|65|14|看哪，我的仆人因心中喜乐而欢呼， 你们却因心里悲痛而哀哭， 因灵里忧伤而哀号。
ISA|65|15|你们必留下自己的名 给我选民指着赌咒： 主耶和华必杀你们， 另起别名称呼他的仆人。
ISA|65|16|在地上为自己求福的， 必凭真实的上帝求福； 在地上起誓的， 必指着真实的上帝起誓。 因为从前的患难已被遗忘， 从我眼前消逝。”
ISA|65|17|“看哪，我造新天新地！ 从前的事不再被记念，也不被人放在心上；
ISA|65|18|当因我所造的欢喜快乐，直到永远； 看哪，因为我造 耶路撒冷 为人所喜， 造其中的居民为人所乐。
ISA|65|19|我必因 耶路撒冷 欢喜， 因我的百姓快乐， 那里不再听见哭泣和哀号的声音。
ISA|65|20|那里没有数日夭折的婴孩， 也没有寿数不满的老人； 因为百岁死的仍算孩童， 未达百岁而亡的 算是被诅咒的。
ISA|65|21|他们建造房屋，居住其中， 栽葡萄园，吃园中的果子；
ISA|65|22|并非造了给别人居住， 也非栽种给别人享用； 因为我百姓的日子必长久如树木， 我的选民必享受亲手劳碌得来的。
ISA|65|23|他们必不徒然劳碌， 所生产的，也不遭灾害， 因为他们和他们的子孙 都是蒙耶和华赐福的后裔。
ISA|65|24|他们尚未求告，我就应允； 正说话的时候，我就垂听。
ISA|65|25|野狼必与羔羊同食， 狮子必吃草，与牛一样， 蛇必以尘土为食物； 在我圣山的遍处， 它们都不伤人，也不害物； 这是耶和华说的。”
ISA|66|1|耶和华如此说： “天是我的座位； 地是我的脚凳。 你们能为我造怎样的殿宇呢？ 哪里是我安歇的地方呢？
ISA|66|2|这一切是我手所造的， 这一切就都存在了。 我所看顾的是困苦、灵里痛悔、 因我言语而战兢的人。 这是耶和华说的。
ISA|66|3|“至于那些宰牛，杀人， 献羔羊，打断狗颈项， 献猪血为供物， 烧乳香，称颂偶像的， 他们选择自己的道路， 心里喜爱可憎恶的事；
ISA|66|4|我也必选择苦待他们， 使他们所惧怕的临到他们； 因为我呼唤，无人回应； 我说话，他们不听从； 反倒做我眼中看为恶的事， 选择我所不喜悦的事。”
ISA|66|5|你们因耶和华言语而战兢的人哪，当听他的话： “你们的弟兄，就是恨恶你们， 因我名赶出你们的，曾说： ‘愿耶和华彰显荣耀 ， 好让我们看见你们的喜乐。’ 但蒙羞的终究是他们！
ISA|66|6|“有喧哗的声音出自城中！ 有声音来自殿里！ 是耶和华向仇敌施行报应的声音！
ISA|66|7|“ 锡安 未曾阵痛就生产， 疼痛尚未来到，就生出男孩。
ISA|66|8|国岂能一日而生？ 民岂能一时而产？ 但 锡安 一阵痛就生下儿女， 这样的事有谁听见， 有谁看见呢？
ISA|66|9|耶和华说：我使人临产， 岂不让她 生产呢？ 你的上帝说：我使人生产， 难道还让她关闭 不生吗？
ISA|66|10|“你们所有爱慕 耶路撒冷 的啊， 要与她一同欢喜，为她高兴； 你们所有为她悲哀的啊， 都要与她一同乐上加乐；
ISA|66|11|使你们在她安慰的怀中吃奶得饱， 尽情吸取她丰盛的荣耀，满心喜乐。”
ISA|66|12|耶和华如此说： “看哪，我要使平安临到她，好像江河； 使列国的荣耀及于她，如同涨溢的溪流。 你们要尽情吸吮； 你们必被抱在身旁 ，摇弄在膝上。
ISA|66|13|我要安慰你们，如同母亲安慰儿女； 你们也必在 耶路撒冷 得安慰。
ISA|66|14|你们看见，心里就喜乐， 你们的骨头必如草生长； 耶和华的手在他仆人身上彰显， 他却要向他的仇敌发怒。”
ISA|66|15|看哪，耶和华必在火中降临， 他的战车宛如暴风， 以烈怒施行报应， 以火焰施行责罚；
ISA|66|16|耶和华必以火与刀审判凡有血肉之躯的， 被耶和华所杀的很多。
ISA|66|17|那些洁净自己献给偶像，进入园内，跟随其中一个人去吃猪肉和鼠肉，并可憎之物的，他们必一同灭绝。这是耶和华说的。
ISA|66|18|我知道他们的行为和他们的意念。聚集万国万族 的时候到了 ，他们要来瞻仰我的荣耀；
ISA|66|19|我要在他们中间显神迹，差遣他们当中的幸存者到列国去，就是到 他施 、 普勒 、以善射闻名的 路德 、 土巴 、 雅完 ，和未曾听见我名声，未曾看见我荣耀的遥远海岛那里去；他们必在列国中传扬我的荣耀。
ISA|66|20|他们要将你们的弟兄从列国中带回，或骑马，或坐车，或乘蓬车，或骑骡子，或骑独峰驼，到我的圣山 耶路撒冷 ，作为供物献给耶和华。这是耶和华说的。正如 以色列 人用洁净的器皿盛供物奉到耶和华的殿中，
ISA|66|21|我也必从他们中间立人作祭司，作 利未 人。这是耶和华说的。
ISA|66|22|“我所造的新天新地在我面前长存， 你们的后裔和你们的名号也必照样长存。 这是耶和华说的。
ISA|66|23|每逢初一、安息日， 凡有血肉之躯的必前来，在我面前下拜； 这是耶和华说的。
ISA|66|24|“他们要出去观看那些违背我的人的尸首， 他们的虫是不死的， 他们的火是不灭的， 凡有血肉之躯的都必憎恶他们。”
