JER|1|1|The words of Jeremiah, the son of Hilkiah, one of the priests who were in Anathoth in the land of Benjamin,
JER|1|2|to whom the word of the LORD came in the days of Josiah the son of Amon, king of Judah, in the thirteenth year of his reign.
JER|1|3|It came also in the days of Jehoiakim the son of Josiah, king of Judah, and until the end of the eleventh year of Zedekiah, the son of Josiah, king of Judah, until the captivity of Jerusalem in the fifth month.
JER|1|4|Now the word of the LORD came to me, saying,
JER|1|5|"Before I formed you in the womb I knew you, and before you were born I consecrated you; I appointed you a prophet to the nations."
JER|1|6|Then I said, "Ah, Lord GOD! Behold, I do not know how to speak, for I am only a youth."
JER|1|7|But the LORD said to me, "Do not say, 'I am only a youth'; for to all to whom I send you, you shall go, and whatever I command you, you shall speak.
JER|1|8|Do not be afraid of them, for I am with you to deliver you, declares the LORD."
JER|1|9|Then the LORD put out his hand and touched my mouth. And the LORD said to me, "Behold, I have put my words in your mouth.
JER|1|10|See, I have set you this day over nations and over kingdoms, to pluck up and to break down, to destroy and to overthrow, to build and to plant."
JER|1|11|And the word of the LORD came to me, saying, "Jeremiah, what do you see?" And I said, "I see an almond branch."
JER|1|12|Then the LORD said to me, "You have seen well, for I am watching over my word to perform it."
JER|1|13|The word of the LORD came to me a second time, saying, "What do you see?" And I said, "I see a boiling pot, facing away from the north."
JER|1|14|Then the LORD said to me, "Out of the north disaster shall be let loose upon all the inhabitants of the land.
JER|1|15|For behold, I am calling all the tribes of the kingdoms of the north, declares the LORD, and they shall come, and every one shall set his throne at the entrance of the gates of Jerusalem, against all its walls all around and against all the cities of Judah.
JER|1|16|And I will declare my judgments against them, for all their evil in forsaking me. They have made offerings to other gods and worshiped the works of their own hands.
JER|1|17|But you, dress yourself for work; arise, and say to them everything that I command you. Do not be dismayed by them, lest I dismay you before them.
JER|1|18|And I, behold, I make you this day a fortified city, an iron pillar, and bronze walls, against the whole land, against the kings of Judah, its officials, its priests, and the people of the land.
JER|1|19|They will fight against you, but they shall not prevail against you, for I am with you, declares the LORD, to deliver you."
JER|2|1|The word of the LORD came to me, saying,
JER|2|2|"Go and proclaim in the hearing of Jerusalem, Thus says the LORD, "I remember the devotion of your youth, your love as a bride, how you followed me in the wilderness, in a land not sown.
JER|2|3|Israel was holy to the LORD, the firstfruits of his harvest. All who ate of it incurred guilt; disaster came upon them, declares the LORD."
JER|2|4|Hear the word of the LORD, O house of Jacob, and all the clans of the house of Israel.
JER|2|5|Thus says the LORD: "What wrong did your fathers find in me that they went far from me, and went after worthlessness, and became worthless?
JER|2|6|They did not say, 'Where is the LORD who brought us up from the land of Egypt, who led us in the wilderness, in a land of deserts and pits, in a land of drought and deep darkness, in a land that none passes through, where no man dwells?'
JER|2|7|And I brought you into a plentiful land to enjoy its fruits and its good things. But when you came in, you defiled my land and made my heritage an abomination.
JER|2|8|The priests did not say, 'Where is the LORD?' Those who handle the law did not know me; the shepherds transgressed against me; the prophets prophesied by Baal and went after things that do not profit.
JER|2|9|"Therefore I still contend with you, declares the LORD, and with your children's children I will contend.
JER|2|10|For cross to the coasts of Cyprus and see, or send to Kedar and examine with care; see if there has been such a thing.
JER|2|11|Has a nation changed its gods, even though they are no gods? But my people have changed their glory for that which does not profit.
JER|2|12|Be appalled, O heavens, at this; be shocked, be utterly desolate, declares the LORD,
JER|2|13|for my people have committed two evils: they have forsaken me, the fountain of living waters, and hewed out cisterns for themselves, broken cisterns that can hold no water.
JER|2|14|"Is Israel a slave? Is he a homeborn servant? Why then has he become a prey?
JER|2|15|The lions have roared against him; they have roared loudly. They have made his land a waste; his cities are in ruins, without inhabitant.
JER|2|16|Moreover, the men of Memphis and Tahpanhes have shaved the crown of your head.
JER|2|17|Have you not brought this upon yourself by forsaking the LORD your God, when he led you in the way?
JER|2|18|And now what do you gain by going to Egypt to drink the waters of the Nile? Or what do you gain by going to Assyria to drink the waters of the Euphrates?
JER|2|19|Your evil will chastise you, and your apostasy will reprove you. Know and see that it is evil and bitter for you to forsake the LORD your God; the fear of me is not in you, declares the Lord GOD of hosts.
JER|2|20|"For long ago I broke your yoke and burst your bonds; but you said, 'I will not serve.' yes, on every high hill and under every green tree you bowed down like a whore.
JER|2|21|Yet I planted you a choice vine, wholly of pure seed. How then have you turned degenerate and become a wild vine?
JER|2|22|Though you wash yourself with lye and use much soap, the stain of your guilt is still before me, declares the Lord GOD.
JER|2|23|How can you say, 'I am not unclean, I have not gone after the Baals'? Look at your way in the valley; know what you have done- a restless young camel running here and there,
JER|2|24|a wild donkey used to the wilderness, in her heat sniffing the wind! Who can restrain her lust? None who seek her need weary themselves; in her month they will find her.
JER|2|25|Keep your feet from going unshod and your throat from thirst. But you said, 'It is hopeless, for I have loved foreigners, and after them I will go.'
JER|2|26|"As a thief is shamed when caught, so the house of Israel shall be shamed: they, their kings, their officials, their priests, and their prophets,
JER|2|27|who say to a tree, 'You are my father,' and to a stone, 'You gave me birth.' For they have turned their back to me, and not their face. But in the time of their trouble they say, 'Arise and save us!'
JER|2|28|But where are your gods that you made for yourself? Let them arise, if they can save you, in your time of trouble; for as many as your cities are your gods, O Judah.
JER|2|29|"Why do you contend with me? You have all transgressed against me, declares the LORD.
JER|2|30|In vain have I struck your children; they took no correction; your own sword devoured your prophets like a ravening lion.
JER|2|31|And you, O generation, behold the word of the LORD. Have I been a wilderness to Israel, or a land of thick darkness? Why then do my people say, 'We are free, we will come no more to you'?
JER|2|32|Can a virgin forget her ornaments, or a bride her attire? Yet my people have forgotten me days without number.
JER|2|33|"How well you direct your course to seek love! So that even to wicked women you have taught your ways.
JER|2|34|Also on your skirts is found the lifeblood of the guiltless poor; you did not find them breaking in. Yet in spite of all these things
JER|2|35|you say, 'I am innocent; surely his anger has turned from me.' Behold, I will bring you to judgment for saying, 'I have not sinned.'
JER|2|36|How much you go about, changing your way! You shall be put to shame by Egypt as you were put to shame by Assyria.
JER|2|37|From it too you will come away with your hands on your head, for the LORD has rejected those in whom you trust, and you will not prosper by them.
JER|3|1|"If a man divorces his wife and she goes from him and becomes another man's wife, will he return to her? Would not that land be greatly polluted? You have played the whore with many lovers; and would you return to me? declares the LORD.
JER|3|2|Lift up your eyes to the bare heights, and see! Where have you not been ravished? By the waysides you have sat awaiting lovers like an Arab in the wilderness. You have polluted the land with your vile whoredom.
JER|3|3|Therefore the showers have been withheld, and the spring rain has not come; yet you have the forehead of a whore; you refuse to be ashamed.
JER|3|4|Have you not just now called to me, 'My father, you are the friend of my youth-
JER|3|5|will he be angry forever, will he be indignant to the end?' Behold, you have spoken, but you have done all the evil that you could."
JER|3|6|The LORD said to me in the days of King Josiah: "Have you seen what she did, that faithless one, Israel, how she went up on every high hill and under every green tree, and there played the whore?
JER|3|7|And I thought, 'After she has done all this she will return to me,' but she did not return, and her treacherous sister Judah saw it.
JER|3|8|She saw that for all the adulteries of that faithless one, Israel, I had sent her away with a decree of divorce. Yet her treacherous sister Judah did not fear, but she too went and played the whore.
JER|3|9|Because she took her whoredom lightly, she polluted the land, committing adultery with stone and tree.
JER|3|10|Yet for all this her treacherous sister Judah did not return to me with her whole heart, but in pretense, declares the LORD."
JER|3|11|And the LORD said to me, "Faithless Israel has shown herself more righteous than treacherous Judah.
JER|3|12|Go, and proclaim these words toward the north, and say, "' Return, faithless Israel, declares the LORD. I will not look on you in anger, for I am merciful, declares the LORD; I will not be angry forever.
JER|3|13|Only acknowledge your guilt, that you rebelled against the LORD your God and scattered your favors among foreigners under every green tree, and that you have not obeyed my voice, declares the LORD.
JER|3|14|Return, O faithless children, declares the LORD; for I am your master; I will take you, one from a city and two from a family, and I will bring you to Zion.
JER|3|15|"'And I will give you shepherds after my own heart, who will feed you with knowledge and understanding.
JER|3|16|And when you have multiplied and increased in the land, in those days, declares the LORD, they shall no more say, "The ark of the covenant of the LORD." It shall not come to mind or be remembered or missed; it shall not be made again.
JER|3|17|At that time Jerusalem shall be called the throne of the LORD, and all nations shall gather to it, to the presence of the LORD in Jerusalem, and they shall no more stubbornly follow their own evil heart.
JER|3|18|In those days the house of Judah shall join the house of Israel, and together they shall come from the land of the north to the land that I gave your fathers for a heritage.
JER|3|19|"'I said How I would set you among my sons, and give you a pleasant land, a heritage most beautiful of all nations. And I thought you would call me, My Father, and would not turn from following me.
JER|3|20|Surely, as a treacherous wife leaves her husband, so have you been treacherous to me, O house of Israel, declares the LORD.'"
JER|3|21|A voice on the bare heights is heard, the weeping and pleading of Israel's sons because they have perverted their way; they have forgotten the LORD their God.
JER|3|22|"Return, O faithless sons; I will heal your faithlessness." "Behold, we come to you, for you are the LORD our God.
JER|3|23|Truly the hills are a delusion, the orgies on the mountains. Truly in the LORD our God is the salvation of Israel.
JER|3|24|"But from our youth the shameful thing has devoured all for which our fathers labored, their flocks and their herds, their sons and their daughters.
JER|3|25|Let us lie down in our shame, and let our dishonor cover us. For we have sinned against the LORD our God, we and our fathers, from our youth even to this day, and we have not obeyed the voice of the LORD our God."
JER|4|1|"If you return, O Israel, declares the LORD, to me you should return. If you remove your detestable things from my presence, and do not waver,
JER|4|2|and if you swear, 'As the LORD lives,' in truth, in justice, and in righteousness, then nations shall bless themselves in him, and in him shall they glory."
JER|4|3|For thus says the LORD to the men of Judah and Jerusalem: "Break up your fallow ground, and sow not among thorns.
JER|4|4|Circumcise yourselves to the LORD; remove the foreskin of your hearts, O men of Judah and inhabitants of Jerusalem; lest my wrath go forth like fire, and burn with none to quench it, because of the evil of your deeds."
JER|4|5|Declare in Judah, and proclaim in Jerusalem, and say, "Blow the trumpet through the land; cry aloud and say, 'Assemble, and let us go into the fortified cities!'
JER|4|6|Raise a standard toward Zion, flee for safety, stay not, for I bring disaster from the north, and great destruction.
JER|4|7|A lion has gone up from his thicket, a destroyer of nations has set out; he has gone out from his place to make your land a waste; your cities will be ruins without inhabitant.
JER|4|8|For this put on sackcloth, lament, and wail, for the fierce anger of the LORD has not turned back from us."
JER|4|9|"In that day, declares the LORD, courage shall fail both king and officials. The priests shall be appalled and the prophets astounded."
JER|4|10|Then I said, "Ah, Lord GOD, surely you have utterly deceived this people and Jerusalem, saying, 'It shall be well with you,' whereas the sword has reached their very life."
JER|4|11|At that time it will be said to this people and to Jerusalem, "A hot wind from the bare heights in the desert toward the daughter of my people, not to winnow or cleanse,
JER|4|12|a wind too full for this comes for me. Now it is I who speak in judgment upon them."
JER|4|13|Behold, he comes up like clouds; his chariots like the whirlwind; his horses are swifter than eagles- woe to us, for we are ruined!
JER|4|14|O Jerusalem, wash your heart from evil, that you may be saved. How long shall your wicked thoughts lodge within you?
JER|4|15|For a voice declares from Dan and proclaims trouble from Mount Ephraim.
JER|4|16|Warn the nations that he is coming; announce to Jerusalem, "Besiegers come from a distant land; they shout against the cities of Judah.
JER|4|17|Like keepers of a field are they against her all around, because she has rebelled against me, declares the LORD.
JER|4|18|Your ways and your deeds have brought this upon you. This is your doom, and it is bitter; it has reached your very heart."
JER|4|19|My anguish, my anguish! I writhe in pain! Oh the walls of my heart! My heart is beating wildly; I cannot keep silent, for I hear the sound of the trumpet, the alarm of war.
JER|4|20|Crash follows hard on crash; the whole land is laid waste. Suddenly my tents are laid waste, my curtains in a moment.
JER|4|21|How long must I see the standard and hear the sound of the trumpet?
JER|4|22|"For my people are foolish; they know me not; they are stupid children; they have no understanding. They are 'wise'- in doing evil! But how to do good they know not."
JER|4|23|I looked on the earth, and behold, it was without form and void; and to the heavens, and they had no light.
JER|4|24|I looked on the mountains, and behold, they were quaking, and all the hills moved to and fro.
JER|4|25|I looked, and behold, there was no man, and all the birds of the air had fled.
JER|4|26|I looked, and behold, the fruitful land was a desert, and all its cities were laid in ruins before the LORD, before his fierce anger.
JER|4|27|For thus says the LORD, "The whole land shall be a desolation; yet I will not make a full end.
JER|4|28|"For this the earth shall mourn, and the heavens above be dark; for I have spoken; I have purposed; I have not relented, nor will I turn back."
JER|4|29|At the noise of horseman and archer every city takes to flight; they enter thickets; they climb among rocks; all the cities are forsaken, and no man dwells in them.
JER|4|30|And you, O desolate one, what do you mean that you dress in scarlet, that you adorn yourself with ornaments of gold, that you enlarge your eyes with paint? In vain you beautify yourself. Your lovers despise you; they seek your life.
JER|4|31|For I heard a cry as of a woman in labor, anguish as of one giving birth to her first child, the cry of the daughter of Zion gasping for breath, stretching out her hands, "Woe is me! I am fainting before murderers."
JER|5|1|Run to and fro through the streets of Jerusalem, look and take note! Search her squares to see if you can find a man, one who does justice and seeks truth, that I may pardon her.
JER|5|2|Though they say, "As the LORD lives," yet they swear falsely.
JER|5|3|O LORD, do not your eyes look for truth? You have struck them down, but they felt no anguish; you have consumed them, but they refused to take correction. They have made their faces harder than rock; they have refused to repent.
JER|5|4|Then I said, "These are only the poor; they have no sense; for they do not know the way of the LORD, the justice of their God.
JER|5|5|I will go to the great and will speak to them, for they know the way of the LORD, the justice of their God." But they all alike had broken the yoke; they had burst the bonds.
JER|5|6|Therefore a lion from the forest shall strike them down; a wolf from the desert shall devastate them. A leopard is watching their cities; everyone who goes out of them shall be torn in pieces, because their transgressions are many, their apostasies are great.
JER|5|7|"How can I pardon you? Your children have forsaken me and have sworn by those who are no gods. When I fed them to the full, they committed adultery and trooped to the houses of whores.
JER|5|8|They were well-fed, lusty stallions, each neighing for his neighbor's wife.
JER|5|9|Shall I not punish them for these things? declares the LORD; and shall I not avenge myself on a nation such as this?
JER|5|10|"Go up through her vine rows and destroy, but make not a full end; strip away her branches, for they are not the LORD's.
JER|5|11|For the house of Israel and the house of Judah have been utterly treacherous to me, declares the LORD.
JER|5|12|They have spoken falsely of the LORD and have said, 'He will do nothing; no disaster will come upon us, nor shall we see sword or famine.
JER|5|13|The prophets will become wind; the word is not in them. Thus shall it be done to them!'"
JER|5|14|Therefore thus says the LORD, the God of hosts: "Because you have spoken this word, behold, I am making my words in your mouth a fire, and this people wood, and the fire shall consume them.
JER|5|15|Behold, I am bringing against you a nation from afar, O house of Israel, declares the LORD. It is an enduring nation; it is an ancient nation, a nation whose language you do not know, nor can you understand what they say.
JER|5|16|Their quiver is like an open tomb; they are all mighty warriors.
JER|5|17|They shall eat up your harvest and your food; they shall eat up your sons and your daughters; they shall eat up your flocks and your herds; they shall eat up your vines and your fig trees; your fortified cities in which you trust they shall beat down with the sword."
JER|5|18|"But even in those days, declares the LORD, I will not make a full end of you.
JER|5|19|And when your people say, 'Why has the LORD our God done all these things to us?' you shall say to them, 'As you have forsaken me and served foreign gods in your land, so you shall serve foreigners in a land that is not yours.'"
JER|5|20|Declare this in the house of Jacob; proclaim it in Judah:
JER|5|21|"Hear this, O foolish and senseless people, who have eyes, but see not, who have ears, but hear not.
JER|5|22|Do you not fear me? declares the LORD; Do you not tremble before me? I placed the sand as the boundary for the sea, a perpetual barrier that it cannot pass; though the waves toss, they cannot prevail; though they roar, they cannot pass over it.
JER|5|23|But this people has a stubborn and rebellious heart; they have turned aside and gone away.
JER|5|24|They do not say in their hearts, 'Let us fear the LORD our God, who gives the rain in its season, the autumn rain and the spring rain, and keeps for us the weeks appointed for the harvest.'
JER|5|25|Your iniquities have turned these away, and your sins have kept good from you.
JER|5|26|For wicked men are found among my people; they lurk like fowlers lying in wait. They set a trap; they catch men.
JER|5|27|Like a cage full of birds, their houses are full of deceit; therefore they have become great and rich;
JER|5|28|they have grown fat and sleek. They know no bounds in deeds of evil; they judge not with justice the cause of the fatherless, to make it prosper, and they do not defend the rights of the needy.
JER|5|29|Shall I not punish them for these things? declares the LORD, and shall I not avenge myself on a nation such as this?"
JER|5|30|An appalling and horrible thing has happened in the land:
JER|5|31|the prophets prophesy falsely, and the priests rule at their direction; my people love to have it so, but what will you do when the end comes?
JER|6|1|Flee for safety, O people of Benjamin, from the midst of Jerusalem! Blow the trumpet in Tekoa, and raise a signal on Beth-haccherem, for disaster looms out of the north, and great destruction.
JER|6|2|The lovely and delicately bred I will destroy, the daughter of Zion.
JER|6|3|Shepherds with their flocks shall come against her; they shall pitch their tents around her; they shall pasture, each in his place.
JER|6|4|"Prepare war against her; arise, and let us attack at noon! Woe to us, for the day declines, for the shadows of evening lengthen!
JER|6|5|Arise, and let us attack by night and destroy her palaces!"
JER|6|6|For thus says the LORD of hosts: "Cut down her trees; cast up a siege mound against Jerusalem. This is the city that must be punished; there is nothing but oppression within her.
JER|6|7|As a well keeps its water fresh, so she keeps fresh her evil; violence and destruction are heard within her; sickness and wounds are ever before me.
JER|6|8|Be warned, O Jerusalem, lest I turn from you in disgust, lest I make you a desolation, an uninhabited land."
JER|6|9|Thus says the LORD of hosts: "They shall glean thoroughly as a vine the remnant of Israel; like a grape-gatherer pass your hand again over its branches."
JER|6|10|To whom shall I speak and give warning, that they may hear? Behold, their ears are uncircumcised, they cannot listen; behold, the word of the LORD is to them an object of scorn; they take no pleasure in it.
JER|6|11|Therefore I am full of the wrath of the LORD; I am weary of holding it in. "Pour it out upon the children in the street, and upon the gatherings of young men, also; both husband and wife shall be taken, the elderly and the very aged.
JER|6|12|Their houses shall be turned over to others, their fields and wives together, for I will stretch out my hand against the inhabitants of the land," declares the LORD.
JER|6|13|"For from the least to the greatest of them, everyone is greedy for unjust gain; and from prophet to priest, everyone deals falsely.
JER|6|14|They have healed the wound of my people lightly, saying, 'Peace, peace,' when there is no peace.
JER|6|15|Were they ashamed when they committed abomination? No, they were not at all ashamed; they did not know how to blush. Therefore they shall fall among those who fall; at the time that I punish them, they shall be overthrown," says the LORD.
JER|6|16|Thus says the LORD: "Stand by the roads, and look, and ask for the ancient paths, where the good way is; and walk in it, and find rest for your souls. But they said, 'We will not walk in it.'
JER|6|17|I set watchmen over you, saying, 'Pay attention to the sound of the trumpet!' But they said, 'We will not pay attention.'
JER|6|18|Therefore hear, O nations, and know, O congregation, what will happen to them.
JER|6|19|Hear, O earth; behold, I am bringing disaster upon this people, the fruit of their devices, because they have not paid attention to my words; and as for my law, they have rejected it.
JER|6|20|What use to me is frankincense that comes from Sheba, or sweet cane from a distant land? Your burnt offerings are not acceptable, nor your sacrifices pleasing to me.
JER|6|21|Therefore thus says the LORD: 'Behold, I will lay before this people stumbling blocks against which they shall stumble; fathers and sons together, neighbor and friend shall perish.'"
JER|6|22|Thus says the LORD: "Behold, a people is coming from the north country, a great nation is stirring from the farthest parts of the earth.
JER|6|23|They lay hold on bow and javelin; they are cruel and have no mercy; the sound of them is like the roaring sea; they ride on horses, set in array as a man for battle, against you, O daughter of Zion!"
JER|6|24|We have heard the report of it; our hands fall helpless; anguish has taken hold of us, pain as of a woman in labor.
JER|6|25|Go not out into the field, nor walk on the road, for the enemy has a sword; terror is on every side.
JER|6|26|O daughter of my people, put on sackcloth, and roll in ashes; make mourning as for an only son, most bitter lamentation, for suddenly the destroyer will come upon us.
JER|6|27|"I have made you a tester of metals among my people, that you may know and test their ways.
JER|6|28|They are all stubbornly rebellious, going about with slanders; they are bronze and iron; all of them act corruptly.
JER|6|29|The bellows blow fiercely; the lead is consumed by the fire; in vain the refining goes on, for the wicked are not removed.
JER|6|30|Rejected silver they are called, for the LORD has rejected them."
JER|7|1|The word that came to Jeremiah from the LORD:
JER|7|2|"Stand in the gate of the LORD's house, and proclaim there this word, and say, Hear the word of the LORD, all you men of Judah who enter these gates to worship the LORD.
JER|7|3|Thus says the LORD of hosts, the God of Israel: Amend your ways and your deeds, and I will let you dwell in this place.
JER|7|4|Do not trust in these deceptive words: 'This is the temple of the LORD, the temple of the LORD, the temple of the LORD.'
JER|7|5|"For if you truly amend your ways and your deeds, if you truly execute justice one with another,
JER|7|6|if you do not oppress the sojourner, the fatherless, or the widow, or shed innocent blood in this place, and if you do not go after other gods to your own harm,
JER|7|7|then I will let you dwell in this place, in the land that I gave of old to your fathers forever.
JER|7|8|"Behold, you trust in deceptive words to no avail.
JER|7|9|Will you steal, murder, commit adultery, swear falsely, make offerings to Baal, and go after other gods that you have not known,
JER|7|10|and then come and stand before me in this house, which is called by my name, and say, 'We are delivered!'- only to go on doing all these abominations?
JER|7|11|Has this house, which is called by my name, become a den of robbers in your eyes? Behold, I myself have seen it, declares the LORD.
JER|7|12|Go now to my place that was in Shiloh, where I made my name dwell at first, and see what I did to it because of the evil of my people Israel.
JER|7|13|And now, because you have done all these things, declares the LORD, and when I spoke to you persistently you did not listen, and when I called you, you did not answer,
JER|7|14|therefore I will do to the house that is called by my name, and in which you trust, and to the place that I gave to you and to your fathers, as I did to Shiloh.
JER|7|15|And I will cast you out of my sight, as I cast out all your kinsmen, all the offspring of Ephraim.
JER|7|16|"As for you, do not pray for this people, or lift up a cry or prayer for them, and do not intercede with me, for I will not hear you.
JER|7|17|Do you not see what they are doing in the cities of Judah and in the streets of Jerusalem?
JER|7|18|The children gather wood, the fathers kindle fire, and the women knead dough, to make cakes for the queen of heaven. And they pour out drink offerings to other gods, to provoke me to anger.
JER|7|19|Is it I whom they provoke? declares the LORD. Is it not themselves, to their own shame?
JER|7|20|Therefore thus says the Lord GOD: behold, my anger and my wrath will be poured out on this place, upon man and beast, upon the trees of the field and the fruit of the ground; it will burn and not be quenched."
JER|7|21|Thus says the LORD of hosts, the God of Israel: "Add your burnt offerings to your sacrifices, and eat the flesh.
JER|7|22|For in the day that I brought them out of the land of Egypt, I did not speak to your fathers or command them concerning burnt offerings and sacrifices.
JER|7|23|But this command I gave them: 'Obey my voice, and I will be your God, and you shall be my people. And walk in all the way that I command you, that it may be well with you.'
JER|7|24|But they did not obey or incline their ear, but walked in their own counsels and the stubbornness of their evil hearts, and went backward and not forward.
JER|7|25|From the day that your fathers came out of the land of Egypt to this day, I have persistently sent all my servants the prophets to them, day after day.
JER|7|26|Yet they did not listen to me or incline their ear, but stiffened their neck. They did worse than their fathers.
JER|7|27|"So you shall speak all these words to them, but they will not listen to you. You shall call to them, but they will not answer you.
JER|7|28|And you shall say to them, 'This is the nation that did not obey the voice of the LORD their God, and did not accept discipline; truth has perished; it is cut off from their lips.
JER|7|29|"' Cut off your hair and cast it away; raise a lamentation on the bare heights, for the LORD has rejected and forsaken the generation of his wrath.'
JER|7|30|"For the sons of Judah have done evil in my sight, declares the LORD. They have set their detestable things in the house that is called by my name, to defile it.
JER|7|31|And they have built the high places of Topheth, which is in the Valley of the Son of Hinnom, to burn their sons and their daughters in the fire, which I did not command, nor did it come into my mind.
JER|7|32|Therefore, behold, the days are coming, declares the LORD, when it will no more be called Topheth, or the Valley of the Son of Hinnom, but the Valley of Slaughter; for they will bury in Topheth, because there is no room elsewhere.
JER|7|33|And the dead bodies of this people will be food for the birds of the air, and for the beasts of the earth, and none will frighten them away.
JER|7|34|And I will silence in the cities of Judah and in the streets of Jerusalem the voice of mirth and the voice of gladness, the voice of the bridegroom and the voice of the bride, for the land shall become a waste.
JER|8|1|"At that time, declares the LORD, the bones of the kings of Judah, the bones of its officials, the bones of the priests, the bones of the prophets, and the bones of the inhabitants of Jerusalem shall be brought out of their tombs.
JER|8|2|And they shall be spread before the sun and the moon and all the host of heaven, which they have loved and served, which they have gone after, and which they have sought and worshiped. And they shall not be gathered or buried. They shall be as dung on the surface of the ground.
JER|8|3|Death shall be preferred to life by all the remnant that remains of this evil family in all the places where I have driven them, declares the LORD of hosts.
JER|8|4|"You shall say to them, Thus says the LORD: When men fall, do they not rise again? If one turns away, does he not return?
JER|8|5|Why then has this people turned away in perpetual backsliding? They hold fast to deceit; they refuse to return.
JER|8|6|I have paid attention and listened, but they have not spoken rightly; no man relents of his evil, saying, 'What have I done?' Everyone turns to his own course, like a horse plunging headlong into battle.
JER|8|7|Even the stork in the heavens knows her times, and the turtledove, swallow, and crane keep the time of their coming, but my people know not the rules of the LORD.
JER|8|8|"How can you say, 'We are wise, and the law of the LORD is with us'? But behold, the lying pen of the scribes has made it into a lie.
JER|8|9|The wise men shall be put to shame; they shall be dismayed and taken; behold, they have rejected the word of the LORD, so what wisdom is in them?
JER|8|10|Therefore I will give their wives to others and their fields to conquerors, because from the least to the greatest everyone is greedy for unjust gain; from prophet to priest, everyone deals falsely.
JER|8|11|They have healed the wound of my people lightly, saying, 'Peace, peace,' when there is no peace.
JER|8|12|Were they ashamed when they committed abomination? No, they were not at all ashamed; they did not know how to blush. Therefore they shall fall among the fallen; when I punish them, they shall be overthrown, says the LORD.
JER|8|13|When I would gather them, declares the LORD, there are no grapes on the vine, nor figs on the fig tree; even the leaves are withered, and what I gave them has passed away from them."
JER|8|14|Why do we sit still? Gather together; let us go into the fortified cities and perish there, for the LORD our God has doomed us to perish and has given us poisoned water to drink, because we have sinned against the LORD.
JER|8|15|We looked for peace, but no good came; for a time of healing, but behold, terror.
JER|8|16|"The snorting of their horses is heard from Dan; at the sound of the neighing of their stallions the whole land quakes. They come and devour the land and all that fills it, the city and those who dwell in it.
JER|8|17|For behold, I am sending among you serpents, adders that cannot be charmed, and they shall bite you," declares the LORD.
JER|8|18|My joy is gone; grief is upon me; my heart is sick within me.
JER|8|19|Behold, the cry of the daughter of my people from the length and breadth of the land: "Is the LORD not in Zion? Is her King not in her?" "Why have they provoked me to anger with their carved images and with their foreign idols?"
JER|8|20|"The harvest is past, the summer is ended, and we are not saved."
JER|8|21|For the wound of the daughter of my people is my heart wounded; I mourn, and dismay has taken hold on me.
JER|8|22|Is there no balm in Gilead? Is there no physician there? Why then has the health of the daughter of my people not been restored?
JER|9|1|Oh that my head were waters, and my eyes a fountain of tears, that I might weep day and night for the slain of the daughter of my people!
JER|9|2|Oh that I had in the desert a travelers' lodging place, that I might leave my people and go away from them! For they are all adulterers, a company of treacherous men.
JER|9|3|They bend their tongue like a bow; falsehood and not truth has grown strong in the land; for they proceed from evil to evil, and they do not know me, declares the LORD.
JER|9|4|Let everyone beware of his neighbor, and put no trust in any brother, for every brother is a deceiver, and every neighbor goes about as a slanderer.
JER|9|5|Everyone deceives his neighbor, and no one speaks the truth; they have taught their tongue to speak lies; they weary themselves committing iniquity.
JER|9|6|Heaping oppression upon oppression, and deceit upon deceit, they refuse to know me, declares the LORD.
JER|9|7|Therefore thus says the LORD of hosts: "Behold, I will refine them and test them, for what else can I do, because of my people?
JER|9|8|Their tongue is a deadly arrow; it speaks deceitfully; with his mouth each speaks peace to his neighbor, but in his heart he plans an ambush for him.
JER|9|9|Shall I not punish them for these things? declares the LORD, and shall I not avenge myself on a nation such as this?
JER|9|10|"I will take up weeping and wailing for the mountains, and a lamentation for the pastures of the wilderness, because they are laid waste so that no one passes through, and the lowing of cattle is not heard; both the birds of the air and the beasts have fled and are gone.
JER|9|11|I will make Jerusalem a heap of ruins, a lair of jackals, and I will make the cities of Judah a desolation, without inhabitant."
JER|9|12|Who is the man so wise that he can understand this? To whom has the mouth of the LORD spoken, that he may declare it? Why is the land ruined and laid waste like a wilderness, so that no one passes through?
JER|9|13|And the LORD says: "Because they have forsaken my law that I set before them, and have not obeyed my voice or walked in accord with it,
JER|9|14|but have stubbornly followed their own hearts and have gone after the Baals, as their fathers taught them.
JER|9|15|Therefore thus says the LORD of hosts, the God of Israel: Behold, I will feed this people with bitter food, and give them poisonous water to drink.
JER|9|16|I will scatter them among the nations whom neither they nor their fathers have known, and I will send the sword after them, until I have consumed them."
JER|9|17|Thus says the LORD of hosts: "Consider, and call for the mourning women to come; send for the skillful women to come;
JER|9|18|let them make haste and raise a wailing over us, that our eyes may run down with tears and our eyelids flow with water.
JER|9|19|For a sound of wailing is heard from Zion: 'How we are ruined! We are utterly shamed, because we have left the land, because they have cast down our dwellings.'"
JER|9|20|Hear, O women, the word of the LORD, and let your ear receive the word of his mouth; teach to your daughters a lament, and each to her neighbor a dirge.
JER|9|21|For death has come up into our windows; it has entered our palaces, cutting off the children from the streets and the young men from the squares.
JER|9|22|Speak, "Thus declares the LORD: 'The dead bodies of men shall fall like dung upon the open field, like sheaves after the reaper, and none shall gather them.'"
JER|9|23|Thus says the LORD: "Let not the wise man boast in his wisdom, let not the mighty man boast in his might, let not the rich man boast in his riches,
JER|9|24|but let him who boasts boast in this, that he understands and knows me, that I am the LORD who practices steadfast love, justice, and righteousness in the earth. For in these things I delight, declares the LORD."
JER|9|25|"Behold, the days are coming, declares the LORD, when I will punish all those who are circumcised merely in the flesh-
JER|9|26|Egypt, Judah, Edom, the sons of Ammon, Moab, and all who dwell in the desert who cut the corners of their hair, for all these nations are uncircumcised, and all the house of Israel is uncircumcised in heart."
JER|10|1|Hear the word that the LORD speaks to you, O house of Israel.
JER|10|2|Thus says the LORD: "Learn not the way of the nations, nor be dismayed at the signs of the heavens because the nations are dismayed at them,
JER|10|3|for the customs of the peoples are vanity. A tree from the forest is cut down and worked with an axe by the hands of a craftsman.
JER|10|4|They decorate it with silver and gold; they fasten it with hammer and nails so that it cannot move.
JER|10|5|Their idols are like scarecrows in a cucumber field, and they cannot speak; they have to be carried, for they cannot walk. Do not be afraid of them, for they cannot do evil, neither is it in them to do good."
JER|10|6|There is none like you, O LORD; you are great, and your name is great in might.
JER|10|7|Who would not fear you, O King of the nations? For this is your due; for among all the wise ones of the nations and in all their kingdoms there is none like you.
JER|10|8|They are both stupid and foolish; the instruction of idols is but wood!
JER|10|9|Beaten silver is brought from Tarshish, and gold from Uphaz. They are the work of the craftsman and of the hands of the goldsmith; their clothing is violet and purple; they are all the work of skilled men.
JER|10|10|But the LORD is the true God; he is the living God and the everlasting King. At his wrath the earth quakes, and the nations cannot endure his indignation.
JER|10|11|Thus shall you say to them: "The gods who did not make the heavens and the earth shall perish from the earth and from under the heavens."
JER|10|12|It is he who made the earth by his power, who established the world by his wisdom, and by his understanding stretched out the heavens.
JER|10|13|When he utters his voice, there is a tumult of waters in the heavens, and he makes the mist rise from the ends of the earth. He makes lightning for the rain, and he brings forth the wind from his storehouses.
JER|10|14|Every man is stupid and without knowledge; every goldsmith is put to shame by his idols, for his images are false, and there is no breath in them.
JER|10|15|They are worthless, a work of delusion; at the time of their punishment they shall perish.
JER|10|16|Not like these is he who is the portion of Jacob, for he is the one who formed all things, and Israel is the tribe of his inheritance; the LORD of hosts is his name.
JER|10|17|Gather up your bundle from the ground, O you who dwell under siege!
JER|10|18|For thus says the LORD: "Behold, I am slinging out the inhabitants of the land at this time, and I will bring distress on them, that they may feel it."
JER|10|19|Woe is me because of my hurt! My wound is grievous. But I said, "Truly this is an affliction, and I must bear it."
JER|10|20|My tent is destroyed, and all my cords are broken; my children have gone from me, and they are not; there is no one to spread my tent again and to set up my curtains.
JER|10|21|For the shepherds are stupid and do not inquire of the LORD; therefore they have not prospered, and all their flock is scattered.
JER|10|22|A voice, a rumor! Behold, it comes!- a great commotion out of the north country to make the cities of Judah a desolation, a lair of jackals.
JER|10|23|I know, O LORD, that the way of man is not in himself, that it is not in man who walks to direct his steps.
JER|10|24|Correct me, O LORD, but in justice; not in your anger, lest you bring me to nothing.
JER|10|25|Pour out your wrath on the nations that know you not, and on the peoples that call not on your name, for they have devoured Jacob; they have devoured him and consumed him, and have laid waste his habitation.
JER|11|1|The word that came to Jeremiah from the LORD:
JER|11|2|"Hear the words of this covenant, and speak to the men of Judah and the inhabitants of Jerusalem.
JER|11|3|You shall say to them, Thus says the LORD, the God of Israel: Cursed be the man who does not hear the words of this covenant
JER|11|4|that I commanded your fathers when I brought them out of the land of Egypt, from the iron furnace, saying, Listen to my voice, and do all that I command you. So shall you be my people, and I will be your God,
JER|11|5|that I may confirm the oath that I swore to your fathers, to give them a land flowing with milk and honey, as at this day." Then I answered, "So be it, LORD."
JER|11|6|And the LORD said to me, "Proclaim all these words in the cities of Judah and in the streets of Jerusalem: Hear the words of this covenant and do them.
JER|11|7|For I solemnly warned your fathers when I brought them up out of the land of Egypt, warning them persistently, even to this day, saying, Obey my voice.
JER|11|8|Yet they did not obey or incline their ear, but everyone walked in the stubbornness of his evil heart. Therefore I brought upon them all the words of this covenant, which I commanded them to do, but they did not."
JER|11|9|Again the LORD said to me, "A conspiracy exists among the men of Judah and the inhabitants of Jerusalem.
JER|11|10|They have turned back to the iniquities of their forefathers, who refused to hear my words. They have gone after other gods to serve them. The house of Israel and the house of Judah have broken my covenant that I made with their fathers.
JER|11|11|Therefore, thus says the LORD, behold, I am bringing disaster upon them that they cannot escape. Though they cry to me, I will not listen to them.
JER|11|12|Then the cities of Judah and the inhabitants of Jerusalem will go and cry to the gods to whom they make offerings, but they cannot save them in the time of their trouble.
JER|11|13|For your gods have become as many as your cities, O Judah, and as many as the streets of Jerusalem are the altars you have set up to shame, altars to make offerings to Baal.
JER|11|14|"Therefore do not pray for this people, or lift up a cry or prayer on their behalf, for I will not listen when they call to me in the time of their trouble.
JER|11|15|What right has my beloved in my house, when she has done many vile deeds? Can even sacrificial flesh avert your doom? Can you then exult?
JER|11|16|The LORD once called you 'a green olive tree, beautiful with good fruit.' But with the roar of a great tempest he will set fire to it, and its branches will be consumed.
JER|11|17|The LORD of hosts, who planted you, has decreed disaster against you, because of the evil that the house of Israel and the house of Judah have done, provoking me to anger by making offerings to Baal."
JER|11|18|The LORD made it known to me and I knew; then you showed me their deeds.
JER|11|19|But I was like a gentle lamb led to the slaughter. I did not know it was against me they devised schemes, saying, "Let us destroy the tree with its fruit, let us cut him off from the land of the living, that his name be remembered no more."
JER|11|20|But, O LORD of hosts, who judges righteously, who tests the heart and the mind, let me see your vengeance upon them, for to you have I committed my cause.
JER|11|21|Therefore thus says the LORD concerning the men of Anathoth, who seek your life, and say, "Do not prophesy in the name of the LORD, or you will die by our hand"-
JER|11|22|therefore thus says the LORD of hosts: "Behold, I will punish them. The young men shall die by the sword, their sons and their daughters shall die by famine,
JER|11|23|and none of them shall be left. For I will bring disaster upon the men of Anathoth, the year of their punishment."
JER|12|1|Righteous are you, O LORD, when I complain to you; yet I would plead my case before you. Why does the way of the wicked prosper? Why do all who are treacherous thrive?
JER|12|2|You plant them, and they take root; they grow and produce fruit; you are near in their mouth and far from their heart.
JER|12|3|But you, O LORD, know me; you see me, and test my heart toward you. Pull them out like sheep for the slaughter, and set them apart for the day of slaughter.
JER|12|4|How long will the land mourn and the grass of every field wither? For the evil of those who dwell in it the beasts and the birds are swept away, because they said, "He will not see our latter end."
JER|12|5|"If you have raced with men on foot, and they have wearied you, how will you compete with horses? And if in a safe land you are so trusting, what will you do in the thicket of the Jordan?
JER|12|6|For even your brothers and the house of your father, even they have dealt treacherously with you; they are in full cry after you; do not believe them, though they speak friendly words to you."
JER|12|7|"I have forsaken my house; I have abandoned my heritage; I have given the beloved of my soul into the hands of her enemies.
JER|12|8|My heritage has become to me like a lion in the forest; she has lifted up her voice against me; therefore I hate her.
JER|12|9|Is my heritage to me like a hyena's lair? Are the birds of prey against her all around? Go, assemble all the wild beasts; bring them to devour.
JER|12|10|Many shepherds have destroyed my vineyard; they have trampled down my portion; they have made my pleasant portion a desolate wilderness.
JER|12|11|They have made it a desolation; desolate, it mourns to me. The whole land is made desolate, but no man lays it to heart.
JER|12|12|Upon all the bare heights in the desert destroyers have come, for the sword of the LORD devours from one end of the land to the other; no flesh has peace.
JER|12|13|They have sown wheat and have reaped thorns; they have tired themselves out but profit nothing. They shall be ashamed of their harvests because of the fierce anger of the LORD."
JER|12|14|Thus says the LORD concerning all my evil neighbors who touch the heritage that I have given my people Israel to inherit: "Behold, I will pluck them up from their land, and I will pluck up the house of Judah from among them.
JER|12|15|And after I have plucked them up, I will again have compassion on them, and I will bring them again each to his heritage and each to his land.
JER|12|16|And it shall come to pass, if they will diligently learn the ways of my people, to swear by my name, 'As the LORD lives,' even as they taught my people to swear by Baal, then they shall be built up in the midst of my people.
JER|12|17|But if any nation will not listen, then I will utterly pluck it up and destroy it, declares the LORD."
JER|13|1|Thus says the LORD to me, "Go and buy a linen loincloth and put it around your waist, and do not dip it in water."
JER|13|2|So I bought a loincloth according to the word of the LORD, and put it around my waist.
JER|13|3|And the word of the LORD came to me a second time,
JER|13|4|"Take the loincloth that you have bought, which is around your waist, and arise, go to the Euphrates and hide it there in a cleft of the rock."
JER|13|5|So I went and hid it by the Euphrates, as the LORD commanded me.
JER|13|6|And after many days the LORD said to me, "Arise, go to the Euphrates, and take from there the loincloth that I commanded you to hide there."
JER|13|7|Then I went to the Euphrates, and dug, and I took the loincloth from the place where I had hidden it. And behold, the loincloth was spoiled; it was good for nothing.
JER|13|8|Then the word of the LORD came to me:
JER|13|9|"Thus says the LORD: Even so will I spoil the pride of Judah and the great pride of Jerusalem.
JER|13|10|This evil people, who refuse to hear my words, who stubbornly follow their own heart and have gone after other gods to serve them and worship them, shall be like this loincloth, which is good for nothing.
JER|13|11|For as the loincloth clings to the waist of a man, so I made the whole house of Israel and the whole house of Judah cling to me, declares the LORD, that they might be for me a people, a name, a praise, and a glory, but they would not listen.
JER|13|12|"You shall speak to them this word: 'Thus says the LORD, the God of Israel, "Every jar shall be filled with wine."' And they will say to you, 'Do we not indeed know that every jar will be filled with wine?'
JER|13|13|Then you shall say to them, 'Thus says the LORD: Behold, I will fill with drunkenness all the inhabitants of this land: the kings who sit on David's throne, the priests, the prophets, and all the inhabitants of Jerusalem.
JER|13|14|And I will dash them one against another, fathers and sons together, declares the LORD. I will not pity or spare or have compassion, that I should not destroy them.'"
JER|13|15|Hear and give ear; be not proud, for the LORD has spoken.
JER|13|16|Give glory to the LORD your God before he brings darkness, before your feet stumble on the twilight mountains, and while you look for light he turns it into gloom and makes it deep darkness.
JER|13|17|But if you will not listen, my soul will weep in secret for your pride; my eyes will weep bitterly and run down with tears, because the LORD's flock has been taken captive.
JER|13|18|Say to the king and the queen mother: "Take a lowly seat, for your beautiful crown has come down from your head."
JER|13|19|The cities of the Negeb are shut up, with none to open them; all Judah is taken into exile, wholly taken into exile.
JER|13|20|"Lift up your eyes and see those who come from the north. Where is the flock that was given you, your beautiful flock?
JER|13|21|What will you say when they set as head over you those whom you yourself have taught to be friends to you? Will not pangs take hold of you like those of a woman in labor?
JER|13|22|And if you say in your heart, 'Why have these things come upon me?' it is for the greatness of your iniquity that your skirts are lifted up and you suffer violence.
JER|13|23|Can the Ethiopian change his skin or the leopard his spots? Then also you can do good who are accustomed to do evil.
JER|13|24|I will scatter you like chaff driven by the wind from the desert.
JER|13|25|This is your lot, the portion I have measured out to you, declares the LORD, because you have forgotten me and trusted in lies.
JER|13|26|I myself will lift up your skirts over your face, and your shame will be seen.
JER|13|27|I have seen your abominations, your adulteries and neighings, your lewd whorings, on the hills in the field. Woe to you, O Jerusalem! How long will it be before you are made clean?"
JER|14|1|The word of the LORD that came to Jeremiah concerning the drought:
JER|14|2|"Judah mourns and her gates languish; her people lament on the ground, and the cry of Jerusalem goes up.
JER|14|3|Her nobles send their servants for water; they come to the cisterns; they find no water; they return with their vessels empty; they are ashamed and confounded and cover their heads.
JER|14|4|Because of the ground that is dismayed, since there is no rain on the land, the farmers are ashamed; they cover their heads.
JER|14|5|Even the doe in the field forsakes her newborn fawn because there is no grass.
JER|14|6|The wild donkeys stand on the bare heights; they pant for air like jackals; their eyes fail because there is no vegetation.
JER|14|7|"Though our iniquities testify against us, act, O LORD, for your name's sake; for our backslidings are many; we have sinned against you.
JER|14|8|O you hope of Israel, its savior in time of trouble, why should you be like a stranger in the land, like a traveler who turns aside to tarry for a night?
JER|14|9|Why should you be like a man confused, like a mighty warrior who cannot save? Yet you, O LORD, are in the midst of us, and we are called by your name; do not leave us."
JER|14|10|Thus says the LORD concerning this people: "They have loved to wander thus; they have not restrained their feet; therefore the LORD does not accept them; now he will remember their iniquity and punish their sins."
JER|14|11|The LORD said to me: "Do not pray for the welfare of this people.
JER|14|12|Though they fast, I will not hear their cry, and though they offer burnt offering and grain offering, I will not accept them. But I will consume them by the sword, by famine, and by pestilence."
JER|14|13|Then I said: "Ah, Lord GOD, behold, the prophets say to them, 'You shall not see the sword, nor shall you have famine, but I will give you assured peace in this place.'"
JER|14|14|And the LORD said to me: "The prophets are prophesying lies in my name. I did not send them, nor did I command them or speak to them. They are prophesying to you a lying vision, worthless divination, and the deceit of their own minds.
JER|14|15|Therefore thus says the LORD concerning the prophets who prophesy in my name although I did not send them, and who say, 'Sword and famine shall not come upon this land': By sword and famine those prophets shall be consumed.
JER|14|16|And the people to whom they prophesy shall be cast out in the streets of Jerusalem, victims of famine and sword, with none to bury them- them, their wives, their sons, and their daughters. For I will pour out their evil upon them.
JER|14|17|"You shall say to them this word: 'Let my eyes run down with tears night and day, and let them not cease, for the virgin daughter of my people is shattered with a great wound, with a very grievous blow.
JER|14|18|If I go out into the field, behold, those pierced by the sword! And if I enter the city, behold, the diseases of famine! For both prophet and priest ply their trade through the land and have no knowledge.'"
JER|14|19|Have you utterly rejected Judah? Does your soul loathe Zion? Why have you struck us down so that there is no healing for us? We looked for peace, but no good came; for a time of healing, but behold, terror.
JER|14|20|We acknowledge our wickedness, O LORD, and the iniquity of our fathers, for we have sinned against you.
JER|14|21|Do not spurn us, for your name's sake; do not dishonor your glorious throne; remember and do not break your covenant with us.
JER|14|22|Are there any among the false gods of the nations that can bring rain? Or can the heavens give showers? Are you not he, O LORD our God? We set our hope on you, for you do all these things.
JER|15|1|Then the LORD said to me, "Though Moses and Samuel stood before me, yet my heart would not turn toward this people. Send them out of my sight, and let them go!
JER|15|2|And when they ask you, 'Where shall we go?' you shall say to them, 'Thus says the LORD: "' Those who are for pestilence, to pestilence, and those who are for the sword, to the sword; those who are for famine, to famine, and those who are for captivity, to captivity.'
JER|15|3|I will appoint over them four kinds of destroyers, declares the LORD: the sword to kill, the dogs to tear, and the birds of the air and the beasts of the earth to devour and destroy.
JER|15|4|And I will make them a horror to all the kingdoms of the earth because of what Manasseh the son of Hezekiah, king of Judah, did in Jerusalem.
JER|15|5|"Who will have pity on you, O Jerusalem, or who will grieve for you? Who will turn aside to ask about your welfare?
JER|15|6|You have rejected me, declares the LORD; you keep going backward, so I have stretched out my hand against you and destroyed you- I am weary of relenting.
JER|15|7|I have winnowed them with a winnowing fork in the gates of the land; I have bereaved them; I have destroyed my people; they did not turn from their ways.
JER|15|8|I have made their widows more in number than the sand of the seas; I have brought against the mothers of young men a destroyer at noonday; I have made anguish and terror fall upon them suddenly.
JER|15|9|She who bore seven has grown feeble; she has fainted away; her sun went down while it was yet day; she has been shamed and disgraced. And the rest of them I will give to the sword before their enemies, declares the LORD."
JER|15|10|Woe is me, my mother, that you bore me, a man of strife and contention to the whole land! I have not lent, nor have I borrowed, yet all of them curse me.
JER|15|11|The LORD said, "Have I not set you free for their good? Have I not pleaded for you before the enemy in the time of trouble and in the time of distress?
JER|15|12|Can one break iron, iron from the north, and bronze?
JER|15|13|"Your wealth and your treasures I will give as spoil, without price, for all your sins, throughout all your territory.
JER|15|14|I will make you serve your enemies in a land that you do not know, for in my anger a fire is kindled that shall burn forever."
JER|15|15|O LORD, you know; remember me and visit me, and take vengeance for me on my persecutors. In your forbearance take me not away; know that for your sake I bear reproach.
JER|15|16|Your words were found, and I ate them, and your words became to me a joy and the delight of my heart, for I am called by your name, O LORD, God of hosts.
JER|15|17|I did not sit in the company of revelers, nor did I rejoice; I sat alone, because your hand was upon me, for you had filled me with indignation.
JER|15|18|Why is my pain unceasing, my wound incurable, refusing to be healed? Will you be to me like a deceitful brook, like waters that fail?
JER|15|19|Therefore thus says the LORD: "If you return, I will restore you, and you shall stand before me. If you utter what is precious, and not what is worthless, you shall be as my mouth. They shall turn to you, but you shall not turn to them.
JER|15|20|And I will make you to this people a fortified wall of bronze; they will fight against you, but they shall not prevail over you, for I am with you to save you and deliver you, declares the LORD.
JER|15|21|I will deliver you out of the hand of the wicked, and redeem you from the grasp of the ruthless."
JER|16|1|The word of the LORD came to me:
JER|16|2|"You shall not take a wife, nor shall you have sons or daughters in this place.
JER|16|3|For thus says the LORD concerning the sons and daughters who are born in this place, and concerning the mothers who bore them and the fathers who fathered them in this land:
JER|16|4|They shall die of deadly diseases. They shall not be lamented, nor shall they be buried. They shall be as dung on the surface of the ground. They shall perish by the sword and by famine, and their dead bodies shall be food for the birds of the air and for the beasts of the earth.
JER|16|5|"For thus says the LORD: Do not enter the house of mourning, or go to lament or grieve for them, for I have taken away my peace from this people, my steadfast love and mercy, declares the LORD.
JER|16|6|Both great and small shall die in this land. They shall not be buried, and no one shall lament for them or cut himself or make himself bald for them.
JER|16|7|No one shall break bread for the mourner, to comfort him for the dead, nor shall anyone give him the cup of consolation to drink for his father or his mother.
JER|16|8|You shall not go into the house of feasting to sit with them, to eat and drink.
JER|16|9|For thus says the LORD of hosts, the God of Israel: Behold, I will silence in this place, before your eyes and in your days, the voice of mirth and the voice of gladness, the voice of the bridegroom and the voice of the bride.
JER|16|10|"And when you tell this people all these words, and they say to you, 'Why has the LORD pronounced all this great evil against us? What is our iniquity? What is the sin that we have committed against the LORD our God?'
JER|16|11|then you shall say to them: 'Because your fathers have forsaken me, declares the LORD, and have gone after other gods and have served and worshiped them, and have forsaken me and have not kept my law,
JER|16|12|and because you have done worse than your fathers, for behold, every one of you follows his stubborn, evil will, refusing to listen to me.
JER|16|13|Therefore I will hurl you out of this land into a land that neither you nor your fathers have known, and there you shall serve other gods day and night, for I will show you no favor.'
JER|16|14|"Therefore, behold, the days are coming, declares the LORD, when it shall no longer be said, 'As the LORD lives who brought up the people of Israel out of the land of Egypt,'
JER|16|15|but 'As the LORD lives who brought up the people of Israel out of the north country and out of all the countries where he had driven them.' For I will bring them back to their own land that I gave to their fathers.
JER|16|16|"Behold, I am sending for many fishers, declares the LORD, and they shall catch them. And afterward I will send for many hunters, and they shall hunt them from every mountain and every hill, and out of the clefts of the rocks.
JER|16|17|For my eyes are on all their ways. They are not hidden from me, nor is their iniquity concealed from my eyes.
JER|16|18|But first I will doubly repay their iniquity and their sin, because they have polluted my land with the carcasses of their detestable idols, and have filled my inheritance with their abominations."
JER|16|19|O LORD, my strength and my stronghold, my refuge in the day of trouble, to you shall the nations come from the ends of the earth and say: "Our fathers have inherited nothing but lies, worthless things in which there is no profit.
JER|16|20|Can man make for himself gods? Such are not gods!"
JER|16|21|"Therefore, behold, I will make them know, this once I will make them know my power and my might, and they shall know that my name is the LORD."
JER|17|1|"The sin of Judah is written with a pen of iron; with a point of diamond it is engraved on the tablet of their heart, and on the horns of their altars,
JER|17|2|while their children remember their altars and their Asherim, beside every green tree and on the high hills,
JER|17|3|on the mountains in the open country. Your wealth and all your treasures I will give for spoil as the price of your high places for sin throughout all your territory.
JER|17|4|You shall loosen your hand from your heritage that I gave to you, and I will make you serve your enemies in a land that you do not know, for in my anger a fire is kindled that shall burn forever."
JER|17|5|Thus says the LORD: "Cursed is the man who trusts in man and makes flesh his strength, whose heart turns away from the LORD.
JER|17|6|He is like a shrub in the desert, and shall not see any good come. He shall dwell in the parched places of the wilderness, in an uninhabited salt land.
JER|17|7|"Blessed is the man who trusts in the LORD, whose trust is the LORD.
JER|17|8|He is like a tree planted by water, that sends out its roots by the stream, and does not fear when heat comes, for its leaves remain green, and is not anxious in the year of drought, for it does not cease to bear fruit."
JER|17|9|The heart is deceitful above all things, and desperately sick; who can understand it?
JER|17|10|"I the LORD search the heart and test the mind, to give every man according to his ways, according to the fruit of his deeds."
JER|17|11|Like the partridge that gathers a brood that she did not hatch, so is he who gets riches but not by justice; in the midst of his days they will leave him, and at his end he will be a fool.
JER|17|12|A glorious throne set on high from the beginning is the place of our sanctuary.
JER|17|13|O LORD, the hope of Israel, all who forsake you shall be put to shame; those who turn away from you shall be written in the earth, for they have forsaken the LORD, the fountain of living water.
JER|17|14|Heal me, O LORD, and I shall be healed; save me, and I shall be saved, for you are my praise.
JER|17|15|Behold, they say to me, "Where is the word of the LORD? Let it come!"
JER|17|16|I have not run away from being your shepherd, nor have I desired the day of sickness. You know what came out of my lips; it was before your face.
JER|17|17|Be not a terror to me; you are my refuge in the day of disaster.
JER|17|18|Let those be put to shame who persecute me, but let me not be put to shame; let them be dismayed, but let me not be dismayed; bring upon them the day of disaster; destroy them with double destruction!
JER|17|19|Thus said the LORD to me: "Go and stand in the People's Gate, by which the kings of Judah enter and by which they go out, and in all the gates of Jerusalem,
JER|17|20|and say: 'Hear the word of the LORD, you kings of Judah, and all Judah, and all the inhabitants of Jerusalem, who enter by these gates.
JER|17|21|Thus says the LORD: Take care for the sake of your lives, and do not bear a burden on the Sabbath day or bring it in by the gates of Jerusalem.
JER|17|22|And do not carry a burden out of your houses on the Sabbath or do any work, but keep the Sabbath day holy, as I commanded your fathers.
JER|17|23|Yet they did not listen or incline their ear, but stiffened their neck, that they might not hear and receive instruction.
JER|17|24|"'But if you listen to me, declares the LORD, and bring in no burden by the gates of this city on the Sabbath day, but keep the Sabbath day holy and do no work on it,
JER|17|25|then there shall enter by the gates of this city kings and princes who sit on the throne of David, riding in chariots and on horses, they and their officials, the men of Judah and the inhabitants of Jerusalem. And this city shall be inhabited forever.
JER|17|26|And people shall come from the cities of Judah and the places around Jerusalem, from the land of Benjamin, from the Shephelah, from the hill country, and from the Negeb, bringing burnt offerings and sacrifices, grain offerings and frankincense, and bringing thank offerings to the house of the LORD.
JER|17|27|But if you do not listen to me, to keep the Sabbath day holy, and not to bear a burden and enter by the gates of Jerusalem on the Sabbath day, then I will kindle a fire in its gates, and it shall devour the palaces of Jerusalem and shall not be quenched.'"
JER|18|1|The word that came to Jeremiah from the LORD:
JER|18|2|"Arise, and go down to the potter's house, and there I will let you hear my words."
JER|18|3|So I went down to the potter's house, and there he was working at his wheel.
JER|18|4|And the vessel he was making of clay was spoiled in the potter's hand, and he reworked it into another vessel, as it seemed good to the potter to do.
JER|18|5|Then the word of the LORD came to me:
JER|18|6|"O house of Israel, can I not do with you as this potter has done? declares the LORD. Behold, like the clay in the potter's hand, so are you in my hand, O house of Israel.
JER|18|7|If at any time I declare concerning a nation or a kingdom, that I will pluck up and break down and destroy it,
JER|18|8|and if that nation, concerning which I have spoken, turns from its evil, I will relent of the disaster that I intended to do to it.
JER|18|9|And if at any time I declare concerning a nation or a kingdom that I will build and plant it,
JER|18|10|and if it does evil in my sight, not listening to my voice, then I will relent of the good that I had intended to do to it.
JER|18|11|Now, therefore, say to the men of Judah and the inhabitants of Jerusalem: 'Thus says the LORD, behold, I am shaping disaster against you and devising a plan against you. Return, every one from his evil way, and amend your ways and your deeds.'
JER|18|12|"But they say, 'That is in vain! We will follow our own plans, and will every one act according to the stubbornness of his evil heart.'
JER|18|13|"Therefore thus says the LORD: Ask among the nations, Who has heard the like of this? The virgin Israel has done a very horrible thing.
JER|18|14|Does the snow of Lebanon leave the crags of Sirion? Do the mountain waters run dry, the cold flowing streams?
JER|18|15|But my people have forgotten me; they make offerings to false gods; they made them stumble in their ways, in the ancient roads, and to walk into side roads, not the highway,
JER|18|16|making their land a horror, a thing to be hissed at forever. Everyone who passes by it is horrified and shakes his head.
JER|18|17|Like the east wind I will scatter them before the enemy. I will show them my back, not my face, in the day of their calamity."
JER|18|18|Then they said, "Come, let us make plots against Jeremiah, for the law shall not perish from the priest, nor counsel from the wise, nor the word from the prophet. Come, let us strike him with the tongue, and let us not pay attention to any of his words."
JER|18|19|Hear me, O LORD, and listen to the voice of my adversaries.
JER|18|20|Should good be repaid with evil? Yet they have dug a pit for my life. Remember how I stood before you to speak good for them, to turn away your wrath from them.
JER|18|21|Therefore deliver up their children to famine; give them over to the power of the sword; let their wives become childless and widowed. May their men meet death by pestilence, their youths be struck down by the sword in battle.
JER|18|22|May a cry be heard from their houses, when you bring the plunderer suddenly upon them! For they have dug a pit to take me and laid snares for my feet.
JER|18|23|Yet you, O LORD, know all their plotting to kill me. Forgive not their iniquity, nor blot out their sin from your sight. Let them be overthrown before you; deal with them in the time of your anger.
JER|19|1|Thus says the LORD, "Go, buy a potter's earthenware flask, and take some of the elders of the people and some of the elders of the priests,
JER|19|2|and go out to the Valley of the Son of Hinnom at the entry of the Potsherd Gate, and proclaim there the words that I tell you.
JER|19|3|You shall say, 'Hear the word of the LORD, O kings of Judah and inhabitants of Jerusalem. Thus says the LORD of hosts, the God of Israel: Behold, I am bringing such disaster upon this place that the ears of everyone who hears of it will tingle.
JER|19|4|Because the people have forsaken me and have profaned this place by making offerings in it to other gods whom neither they nor their fathers nor the kings of Judah have known; and because they have filled this place with the blood of innocents,
JER|19|5|and have built the high places of Baal to burn their sons in the fire as burnt offerings to Baal, which I did not command or decree, nor did it come into my mind-
JER|19|6|therefore, behold, days are coming, declares the LORD, when this place shall no more be called Topheth, or the Valley of the Son of Hinnom, but the Valley of Slaughter.
JER|19|7|And in this place I will make void the plans of Judah and Jerusalem, and will cause their people to fall by the sword before their enemies, and by the hand of those who seek their life. I will give their dead bodies for food to the birds of the air and to the beasts of the earth.
JER|19|8|And I will make this city a horror, a thing to be hissed at. Everyone who passes by it will be horrified and will hiss because of all its wounds.
JER|19|9|And I will make them eat the flesh of their sons and their daughters, and everyone shall eat the flesh of his neighbor in the siege and in the distress, with which their enemies and those who seek their life afflict them.'
JER|19|10|"Then you shall break the flask in the sight of the men who go with you,
JER|19|11|and shall say to them, 'Thus says the LORD of hosts: So will I break this people and this city, as one breaks a potter's vessel, so that it can never be mended. Men shall bury in Topheth because there will be no place else to bury.
JER|19|12|Thus will I do to this place, declares the LORD, and to its inhabitants, making this city like Topheth.
JER|19|13|The houses of Jerusalem and the houses of the kings of Judah- all the houses on whose roofs offerings have been offered to all the host of heaven, and drink offerings have been poured out to other gods- shall be defiled like the place of Topheth.'"
JER|19|14|Then Jeremiah came from Topheth, where the LORD had sent him to prophesy, and he stood in the court of the LORD's house and said to all the people:
JER|19|15|"Thus says the LORD of hosts, the God of Israel, behold, I am bringing upon this city and upon all its towns all the disaster that I have pronounced against it, because they have stiffened their neck, refusing to hear my words."
JER|20|1|Now Pashhur the priest, the son of Immer, who was chief officer in the house of the LORD, heard Jeremiah prophesying these things.
JER|20|2|Then Pashhur beat Jeremiah the prophet, and put him in the stocks that were in the upper Benjamin Gate of the house of the LORD.
JER|20|3|The next day, when Pashhur released Jeremiah from the stocks, Jeremiah said to him, "The LORD does not call your name Pashhur, but Terror On Every Side.
JER|20|4|For thus says the LORD: Behold, I will make you a terror to yourself and to all your friends. They shall fall by the sword of their enemies while you look on. And I will give all Judah into the hand of the king of Babylon. He shall carry them captive to Babylon, and shall strike them down with the sword.
JER|20|5|Moreover, I will give all the wealth of the city, all its gains, all its prized belongings, and all the treasures of the kings of Judah into the hand of their enemies, who shall plunder them and seize them and carry them to Babylon.
JER|20|6|And you, Pashhur, and all who dwell in your house, shall go into captivity. To Babylon you shall go, and there you shall die, and there you shall be buried, you and all your friends, to whom you have prophesied falsely."
JER|20|7|O LORD, you have deceived me, and I was deceived; you are stronger than I, and you have prevailed. I have become a laughingstock all the day; everyone mocks me.
JER|20|8|For whenever I speak, I cry out, I shout, "Violence and destruction!" For the word of the LORD has become for me a reproach and derision all day long.
JER|20|9|If I say, "I will not mention him, or speak any more in his name," there is in my heart as it were a burning fire shut up in my bones, and I am weary with holding it in, and I cannot.
JER|20|10|For I hear many whispering. Terror is on every side! "Denounce him! Let us denounce him!" say all my close friends, watching for my fall. "Perhaps he will be deceived; then we can overcome him and take our revenge on him."
JER|20|11|But the LORD is with me as a dread warrior; therefore my persecutors will stumble; they will not overcome me. They will be greatly shamed, for they will not succeed. Their eternal dishonor will never be forgotten.
JER|20|12|O LORD of hosts, who tests the righteous, who sees the heart and the mind, let me see your vengeance upon them, for to you have I committed my cause.
JER|20|13|Sing to the LORD; praise the LORD! For he has delivered the life of the needy from the hand of evildoers.
JER|20|14|Cursed be the day on which I was born! The day when my mother bore me, let it not be blessed!
JER|20|15|Cursed be the man who brought the news to my father, "A son is born to you," making him very glad.
JER|20|16|Let that man be like the cities that the LORD overthrew without pity; let him hear a cry in the morning and an alarm at noon,
JER|20|17|because he did not kill me in the womb; so my mother would have been my grave, and her womb forever great.
JER|20|18|Why did I come out from the womb to see toil and sorrow, and spend my days in shame?
JER|21|1|This is the word that came to Jeremiah from the LORD, when King Zedekiah sent to him Pashhur the son of Malchiah and Zephaniah the priest, the son of Maaseiah, saying,
JER|21|2|"Inquire of the LORD for us, for Nebuchadnezzar king of Babylon is making war against us. Perhaps the LORD will deal with us according to all his wonderful deeds and will make him withdraw from us."
JER|21|3|Then Jeremiah said to them:
JER|21|4|"Thus you shall say to Zedekiah, 'Thus says the LORD, the God of Israel: Behold, I will turn back the weapons of war that are in your hands and with which you are fighting against the king of Babylon and against the Chaldeans who are besieging you outside the walls. And I will bring them together into the midst of this city.
JER|21|5|I myself will fight against you with outstretched hand and strong arm, in anger and in fury and in great wrath.
JER|21|6|And I will strike down the inhabitants of this city, both man and beast. They shall die of a great pestilence.
JER|21|7|Afterward, declares the LORD, I will give Zedekiah king of Judah and his servants and the people in this city who survive the pestilence, sword, and famine into the hand of Nebuchadnezzar king of Babylon and into the hand of their enemies, into the hand of those who seek their lives. He shall strike them down with the edge of the sword. He shall not pity them or spare them or have compassion.'
JER|21|8|"And to this people you shall say: 'Thus says the LORD: Behold, I set before you the way of life and the way of death.
JER|21|9|He who stays in this city shall die by the sword, by famine, and by pestilence, but he who goes out and surrenders to the Chaldeans who are besieging you shall live and shall have his life as a prize of war.
JER|21|10|For I have set my face against this city for harm and not for good, declares the LORD: it shall be given into the hand of the king of Babylon, and he shall burn it with fire.'
JER|21|11|"And to the house of the king of Judah say, 'Hear the word of the LORD,
JER|21|12|O house of David! Thus says the LORD: "' Execute justice in the morning, and deliver from the hand of the oppressor him who has been robbed, lest my wrath go forth like fire, and burn with none to quench it, because of your evil deeds.'"
JER|21|13|"Behold, I am against you, O inhabitant of the valley, O rock of the plain, declares the LORD; you who say, 'Who shall come down against us, or who shall enter our habitations?'
JER|21|14|I will punish you according to the fruit of your deeds, declares the LORD; I will kindle a fire in her forest, and it shall devour all that is around her."
JER|22|1|Thus says the LORD: "Go down to the house of the king of Judah and speak there this word,
JER|22|2|and say, 'Hear the word of the LORD, O King of Judah, who sits on the throne of David, you, and your servants, and your people who enter these gates.
JER|22|3|Thus says the LORD: Do justice and righteousness, and deliver from the hand of the oppressor him who has been robbed. And do no wrong or violence to the resident alien, the fatherless, and the widow, nor shed innocent blood in this place.
JER|22|4|For if you will indeed obey this word, then there shall enter the gates of this house kings who sit on the throne of David, riding in chariots and on horses, they and their servants and their people.
JER|22|5|But if you will not obey these words, I swear by myself, declares the LORD, that this house shall become a desolation.
JER|22|6|For thus says the LORD concerning the house of the king of Judah: "' You are like Gilead to me, like the summit of Lebanon, yet surely I will make you a desert, an uninhabited city.
JER|22|7|I will prepare destroyers against you, each with his weapons, and they shall cut down your choicest cedars and cast them into the fire.
JER|22|8|"'And many nations will pass by this city, and every man will say to his neighbor, "Why has the LORD dealt thus with this great city?"
JER|22|9|And they will answer, "Because they have forsaken the covenant of the LORD their God and worshiped other gods and served them."'"
JER|22|10|Weep not for him who is dead, nor grieve for him, but weep bitterly for him who goes away, for he shall return no more to see his native land.
JER|22|11|For thus says the LORD concerning Shallum the son of Josiah, king of Judah, who reigned instead of Josiah his father, and who went away from this place: "He shall return here no more,
JER|22|12|but in the place where they have carried him captive, there shall he die, and he shall never see this land again."
JER|22|13|"Woe to him who builds his house by unrighteousness, and his upper rooms by injustice, who makes his neighbor serve him for nothing and does not give him his wages,
JER|22|14|who says, 'I will build myself a great house with spacious upper rooms,' who cuts out windows for it, paneling it with cedar and painting it with vermilion.
JER|22|15|Do you think you are a king because you compete in cedar? Did not your father eat and drink and do justice and righteousness? Then it was well with him.
JER|22|16|He judged the cause of the poor and needy; then it was well. Is not this to know me? declares the LORD.
JER|22|17|But you have eyes and heart only for your dishonest gain, for shedding innocent blood, and for practicing oppression and violence."
JER|22|18|Therefore thus says the LORD concerning Jehoiakim the son of Josiah, king of Judah: "They shall not lament for him, saying, 'Ah, my brother!' or 'Ah, sister!' They shall not lament for him, saying, 'Ah, lord!' or 'Ah, his majesty!'
JER|22|19|With the burial of a donkey he shall be buried, dragged and dumped beyond the gates of Jerusalem."
JER|22|20|"Go up to Lebanon, and cry out, and lift up your voice in Bashan; cry out from Abarim, for all your lovers are destroyed.
JER|22|21|I spoke to you in your prosperity, but you said, 'I will not listen.' This has been your way from your youth, that you have not obeyed my voice.
JER|22|22|The wind shall shepherd all your shepherds, and your lovers shall go into captivity; then you will be ashamed and confounded because of all your evil.
JER|22|23|O inhabitant of Lebanon, nested among the cedars, how you will be pitied when pangs come upon you, pain as of a woman in labor!"
JER|22|24|"As I live, declares the LORD, though Coniah the son of Jehoiakim, king of Judah, were the signet ring on my right hand, yet I would tear you off
JER|22|25|and give you into the hand of those who seek your life, into the hand of those of whom you are afraid, even into the hand of Nebuchadnezzar king of Babylon and into the hand of the Chaldeans.
JER|22|26|I will hurl you and the mother who bore you into another country, where you were not born, and there you shall die.
JER|22|27|But to the land to which they will long to return, there they shall not return."
JER|22|28|Is this man Coniah a despised, broken pot, a vessel no one cares for? Why are he and his children hurled and cast into a land that they do not know?
JER|22|29|O land, land, land, hear the word of the LORD!
JER|22|30|Thus says the LORD: "Write this man down as childless, a man who shall not succeed in his days, for none of his offspring shall succeed in sitting on the throne of David and ruling again in Judah."
JER|23|1|"Woe to the shepherds who destroy and scatter the sheep of my pasture!" declares the LORD.
JER|23|2|Therefore thus says the LORD, the God of Israel, concerning the shepherds who care for my people: "You have scattered my flock and have driven them away, and you have not attended to them. Behold, I will attend to you for your evil deeds, declares the LORD.
JER|23|3|Then I will gather the remnant of my flock out of all the countries where I have driven them, and I will bring them back to their fold, and they shall be fruitful and multiply.
JER|23|4|I will set shepherds over them who will care for them, and they shall fear no more, nor be dismayed, neither shall any be missing, declares the LORD.
JER|23|5|"Behold, the days are coming, declares the LORD, when I will raise up for David a righteous Branch, and he shall reign as king and deal wisely, and shall execute justice and righteousness in the land.
JER|23|6|In his days Judah will be saved, and Israel will dwell securely. And this is the name by which he will be called: 'The LORD is our righteousness.'
JER|23|7|"Therefore, behold, the days are coming, declares the LORD, when they shall no longer say, 'As the LORD lives who brought up the people of Israel out of the land of Egypt,'
JER|23|8|but 'As the LORD lives who brought up and led the offspring of the house of Israel out of the north country and out of all the countries where he had driven them.' Then they shall dwell in their own land."
JER|23|9|Concerning the prophets: My heart is broken within me; all my bones shake; I am like a drunken man, like a man overcome by wine, because of the LORD and because of his holy words.
JER|23|10|For the land is full of adulterers; because of the curse the land mourns, and the pastures of the wilderness are dried up. Their course is evil, and their might is not right.
JER|23|11|"Both prophet and priest are ungodly; even in my house I have found their evil, declares the LORD.
JER|23|12|Therefore their way shall be to them like slippery paths in the darkness, into which they shall be driven and fall, for I will bring disaster upon them in the year of their punishment, declares the LORD.
JER|23|13|In the prophets of Samaria I saw an unsavory thing: they prophesied by Baal and led my people Israel astray.
JER|23|14|But in the prophets of Jerusalem I have seen a horrible thing: they commit adultery and walk in lies; they strengthen the hands of evildoers, so that no one turns from his evil; all of them have become like Sodom to me, and its inhabitants like Gomorrah."
JER|23|15|Therefore thus says the LORD of hosts concerning the prophets: "Behold, I will feed them with bitter food and give them poisoned water to drink, for from the prophets of Jerusalem ungodliness has gone out into all the land."
JER|23|16|Thus says the LORD of hosts: "Do not listen to the words of the prophets who prophesy to you, filling you with vain hopes. They speak visions of their own minds, not from the mouth of the LORD.
JER|23|17|They say continually to those who despise the word of the LORD, 'It shall be well with you'; and to everyone who stubbornly follows his own heart, they say, 'No disaster shall come upon you.'"
JER|23|18|For who among them has stood in the council of the LORD to see and to hear his word, or who has paid attention to his word and listened?
JER|23|19|Behold, the storm of the LORD! Wrath has gone forth, a whirling tempest; it will burst upon the head of the wicked.
JER|23|20|The anger of the LORD will not turn back until he has executed and accomplished the intents of his heart. In the latter days you will understand it clearly.
JER|23|21|"I did not send the prophets, yet they ran; I did not speak to them, yet they prophesied.
JER|23|22|But if they had stood in my council, then they would have proclaimed my words to my people, and they would have turned them from their evil way, and from the evil of their deeds.
JER|23|23|"Am I a God at hand, declares the LORD, and not a God afar off?
JER|23|24|Can a man hide himself in secret places so that I cannot see him? declares the LORD. Do I not fill heaven and earth? declares the LORD.
JER|23|25|I have heard what the prophets have said who prophesy lies in my name, saying, 'I have dreamed, I have dreamed!'
JER|23|26|How long shall there be lies in the heart of the prophets who prophesy lies, and who prophesy the deceit of their own heart,
JER|23|27|who think to make my people forget my name by their dreams that they tell one another, even as their fathers forgot my name for Baal?
JER|23|28|Let the prophet who has a dream tell the dream, but let him who has my word speak my word faithfully. What has straw in common with wheat? declares the LORD.
JER|23|29|Is not my word like fire, declares the LORD, and like a hammer that breaks the rock in pieces?
JER|23|30|Therefore, behold, I am against the prophets, declares the LORD, who steal my words from one another.
JER|23|31|Behold, I am against the prophets, declares the LORD, who use their tongues and declare, 'declares the LORD.'
JER|23|32|Behold, I am against those who prophesy lying dreams, declares the LORD, and who tell them and lead my people astray by their lies and their recklessness, when I did not send them or charge them. So they do not profit this people at all, declares the LORD.
JER|23|33|"When one of this people, or a prophet or a priest asks you, 'What is the burden of the LORD?' you shall say to them, 'You are the burden, and I will cast you off, declares the LORD.'
JER|23|34|And as for the prophet, priest, or one of the people who says, 'The burden of the LORD,' I will punish that man and his household.
JER|23|35|Thus shall you say, every one to his neighbor and every one to his brother, 'What has the LORD answered?' or 'What has the LORD spoken?'
JER|23|36|But 'the burden of the LORD' you shall mention no more, for the burden is every man's own word, and you pervert the words of the living God, the LORD of hosts, our God.
JER|23|37|Thus you shall say to the prophet, 'What has the LORD answered you?' or 'What has the LORD spoken?'
JER|23|38|But if you say, 'The burden of the LORD,' thus says the LORD, 'Because you have said these words, "The burden of the LORD," when I sent to you, saying, "You shall not say, 'The burden of the LORD,'"
JER|23|39|therefore, behold, I will surely lift you up and cast you away from my presence, you and the city that I gave to you and your fathers.
JER|23|40|And I will bring upon you everlasting reproach and perpetual shame, which shall not be forgotten.'"
JER|24|1|After Nebuchadnezzar king of Babylon had taken into exile from Jerusalem Jeconiah the son of Jehoiakim, king of Judah, together with the officials of Judah, the craftsmen, and the metal workers, and had brought them to Babylon, the LORD showed me this vision: behold, two baskets of figs placed before the temple of the LORD.
JER|24|2|One basket had very good figs, like first-ripe figs, but the other basket had very bad figs, so bad that they could not be eaten.
JER|24|3|And the LORD said to me, "What do you see, Jeremiah?" I said, "Figs, the good figs very good, and the bad figs very bad, so bad that they cannot be eaten."
JER|24|4|Then the word of the LORD came to me:
JER|24|5|"Thus says the LORD, the God of Israel: Like these good figs, so I will regard as good the exiles from Judah, whom I have sent away from this place to the land of the Chaldeans.
JER|24|6|I will set my eyes on them for good, and I will bring them back to this land. I will build them up, and not tear them down; I will plant them, and not uproot them.
JER|24|7|I will give them a heart to know that I am the LORD, and they shall be my people and I will be their God, for they shall return to me with their whole heart.
JER|24|8|"But thus says the LORD: Like the bad figs that are so bad they cannot be eaten, so will I treat Zedekiah the king of Judah, his officials, the remnant of Jerusalem who remain in this land, and those who dwell in the land of Egypt.
JER|24|9|I will make them a horror to all the kingdoms of the earth, to be a reproach, a byword, a taunt, and a curse in all the places where I shall drive them.
JER|24|10|And I will send sword, famine, and pestilence upon them, until they shall be utterly destroyed from the land that I gave to them and their fathers."
JER|25|1|The word that came to Jeremiah concerning all the people of Judah, in the fourth year of Jehoiakim the son of Josiah, king of Judah (that was the first year of Nebuchadnezzar king of Babylon),
JER|25|2|which Jeremiah the prophet spoke to all the people of Judah and all the inhabitants of Jerusalem:
JER|25|3|"For twenty-three years, from the thirteenth year of Josiah the son of Amon, king of Judah, to this day, the word of the LORD has come to me, and I have spoken persistently to you, but you have not listened.
JER|25|4|You have neither listened nor inclined your ears to hear, although the LORD persistently sent to you all his servants the prophets,
JER|25|5|saying, 'Turn now, every one of you, from his evil way and evil deeds, and dwell upon the land that the LORD has given to you and your fathers from of old and forever.
JER|25|6|Do not go after other gods to serve and worship them, or provoke me to anger with the work of your hands. Then I will do you no harm.'
JER|25|7|Yet you have not listened to me, declares the LORD, that you might provoke me to anger with the work of your hands to your own harm.
JER|25|8|"Therefore thus says the LORD of hosts: Because you have not obeyed my words,
JER|25|9|behold, I will send for all the tribes of the north, declares the LORD, and for Nebuchadnezzar the king of Babylon, my servant, and I will bring them against this land and its inhabitants, and against all these surrounding nations. I will devote them to destruction, and make them a horror, a hissing, and an everlasting desolation.
JER|25|10|Moreover, I will banish from them the voice of mirth and the voice of gladness, the voice of the bridegroom and the voice of the bride, the grinding of the millstones and the light of the lamp.
JER|25|11|This whole land shall become a ruin and a waste, and these nations shall serve the king of Babylon seventy years.
JER|25|12|Then after seventy years are completed, I will punish the king of Babylon and that nation, the land of the Chaldeans, for their iniquity, declares the LORD, making the land an everlasting waste.
JER|25|13|I will bring upon that land all the words that I have uttered against it, everything written in this book, which Jeremiah prophesied against all the nations.
JER|25|14|For many nations and great kings shall make slaves even of them, and I will recompense them according to their deeds and the work of their hands."
JER|25|15|Thus the LORD, the God of Israel, said to me: "Take from my hand this cup of the wine of wrath, and make all the nations to whom I send you drink it.
JER|25|16|They shall drink and stagger and be crazed because of the sword that I am sending among them."
JER|25|17|So I took the cup from the LORD's hand, and made all the nations to whom the LORD sent me drink it:
JER|25|18|Jerusalem and the cities of Judah, its kings and officials, to make them a desolation and a waste, a hissing and a curse, as at this day;
JER|25|19|Pharaoh king of Egypt, his servants, his officials, all his people,
JER|25|20|and all the mixed tribes among them; all the kings of the land of Uz and all the kings of the land of the Philistines (Ashkelon, Gaza, Ekron, and the remnant of Ashdod);
JER|25|21|Edom, Moab, and the sons of Ammon;
JER|25|22|all the kings of Tyre, all the kings of Sidon, and the kings of the coastland across the sea;
JER|25|23|Dedan, Tema, Buz, and all who cut the corners of their hair;
JER|25|24|all the kings of Arabia and all the kings of the mixed tribes who dwell in the desert;
JER|25|25|all the kings of Zimri, all the kings of Elam, and all the kings of Media;
JER|25|26|all the kings of the north, far and near, one after another, and all the kingdoms of the world that are on the face of the earth. And after them the king of Babylon shall drink.
JER|25|27|"Then you shall say to them, 'Thus says the LORD of hosts, the God of Israel: Drink, be drunk and vomit, fall and rise no more, because of the sword that I am sending among you.'
JER|25|28|"And if they refuse to accept the cup from your hand to drink, then you shall say to them, 'Thus says the LORD of hosts: You must drink!
JER|25|29|For behold, I begin to work disaster at the city that is called by my name, and shall you go unpunished? You shall not go unpunished, for I am summoning a sword against all the inhabitants of the earth, declares the LORD of hosts.'
JER|25|30|"You, therefore, shall prophesy against them all these words, and say to them: "' The LORD will roar from on high, and from his holy habitation utter his voice; he will roar mightily against his fold, and shout, like those who tread grapes, against all the inhabitants of the earth.
JER|25|31|The clamor will resound to the ends of the earth, for the LORD has an indictment against the nations; he is entering into judgment with all flesh, and the wicked he will put to the sword, declares the LORD.'
JER|25|32|"Thus says the LORD of hosts: Behold, disaster is going forth from nation to nation, and a great tempest is stirring from the farthest parts of the earth!
JER|25|33|"And those pierced by the LORD on that day shall extend from one end of the earth to the other. They shall not be lamented, or gathered, or buried; they shall be dung on the surface of the ground.
JER|25|34|"Wail, you shepherds, and cry out, and roll in ashes, you lords of the flock, for the days of your slaughter and dispersion have come, and you shall fall like a choice vessel.
JER|25|35|No refuge will remain for the shepherds, nor escape for the lords of the flock.
JER|25|36|A voice- the cry of the shepherds, and the wail of the lords of the flock! For the LORD is laying waste their pasture,
JER|25|37|and the peaceful folds are devastated because of the fierce anger of the LORD.
JER|25|38|Like a lion he has left his lair, for their land has become a waste because of the sword of the oppressor, and because of his fierce anger."
JER|26|1|In the beginning of the reign of Jehoiakim the son of Josiah, king of Judah, this word came from the LORD:
JER|26|2|"Thus says the LORD: Stand in the court of the LORD's house, and speak to all the cities of Judah that come to worship in the house of the LORD all the words that I command you to speak to them; do not hold back a word.
JER|26|3|It may be they will listen, and every one turn from his evil way, that I may relent of the disaster that I intend to do to them because of their evil deeds.
JER|26|4|You shall say to them, 'Thus says the LORD: If you will not listen to me, to walk in my law that I have set before you,
JER|26|5|and to listen to the words of my servants the prophets whom I send to you urgently, though you have not listened,
JER|26|6|then I will make this house like Shiloh, and I will make this city a curse for all the nations of the earth.'"
JER|26|7|The priests and the prophets and all the people heard Jeremiah speaking these words in the house of the LORD.
JER|26|8|And when Jeremiah had finished speaking all that the LORD had commanded him to speak to all the people, then the priests and the prophets and all the people laid hold of him, saying, "You shall die!
JER|26|9|Why have you prophesied in the name of the LORD, saying, 'This house shall be like Shiloh, and this city shall be desolate, without inhabitant'?" And all the people gathered around Jeremiah in the house of the LORD.
JER|26|10|When the officials of Judah heard these things, they came up from the king's house to the house of the LORD and took their seat in the entry of the New Gate of the house of the LORD.
JER|26|11|Then the priests and the prophets said to the officials and to all the people, "This man deserves the sentence of death, because he has prophesied against this city, as you have heard with your own ears."
JER|26|12|Then Jeremiah spoke to all the officials and all the people, saying, "The LORD sent me to prophesy against this house and this city all the words you have heard.
JER|26|13|Now therefore mend your ways and your deeds, and obey the voice of the LORD your God, and the LORD will relent of the disaster that he has pronounced against you.
JER|26|14|But as for me, behold, I am in your hands. Do with me as seems good and right to you.
JER|26|15|Only know for certain that if you put me to death, you will bring innocent blood upon yourselves and upon this city and its inhabitants, for in truth the LORD sent me to you to speak all these words in your ears."
JER|26|16|Then the officials and all the people said to the priests and the prophets, "This man does not deserve the sentence of death, for he has spoken to us in the name of the LORD our God."
JER|26|17|And certain of the elders of the land arose and spoke to all the assembled people, saying,
JER|26|18|"Micah of Moresheth prophesied in the days of Hezekiah king of Judah, and said to all the people of Judah: 'Thus says the LORD of hosts, "' Zion shall be plowed as a field; Jerusalem shall become a heap of ruins, and the mountain of the house a wooded height.'
JER|26|19|Did Hezekiah king of Judah and all Judah put him to death? Did he not fear the LORD and entreat the favor of the LORD, and did not the LORD relent of the disaster that he had pronounced against them? But we are about to bring great disaster upon ourselves."
JER|26|20|There was another man who prophesied in the name of the LORD, Uriah the son of Shemaiah from Kiriath-jearim. He prophesied against this city and against this land in words like those of Jeremiah.
JER|26|21|And when King Jehoiakim, with all his warriors and all the officials, heard his words, the king sought to put him to death. But when Uriah heard of it, he was afraid and fled and escaped to Egypt.
JER|26|22|Then King Jehoiakim sent to Egypt certain men, Elnathan the son of Achbor and others with him,
JER|26|23|and they took Uriah from Egypt and brought him to King Jehoiakim, who struck him down with the sword and dumped his dead body into the burial place of the common people.
JER|26|24|But the hand of Ahikam the son of Shaphan was with Jeremiah so that he was not given over to the people to be put to death.
JER|27|1|In the beginning of the reign of Zedekiah the son of Josiah, king of Judah, this word came to Jeremiah from the LORD.
JER|27|2|Thus the LORD said to me: "Make yourself straps and yoke-bars, and put them on your neck.
JER|27|3|Send word to the king of Edom, the king of Moab, the king of the sons of Ammon, the king of Tyre, and the king of Sidon by the hand of the envoys who have come to Jerusalem to Zedekiah king of Judah.
JER|27|4|Give them this charge for their masters: 'Thus says the LORD of hosts, the God of Israel: This is what you shall say to your masters:
JER|27|5|"It is I who by my great power and my outstretched arm have made the earth, with the men and animals that are on the earth, and I give it to whomever it seems right to me.
JER|27|6|Now I have given all these lands into the hand of Nebuchadnezzar, the king of Babylon, my servant, and I have given him also the beasts of the field to serve him.
JER|27|7|All the nations shall serve him and his son and his grandson, until the time of his own land comes. Then many nations and great kings shall make him their slave.
JER|27|8|"'"But if any nation or kingdom will not serve this Nebuchadnezzar king of Babylon, and put its neck under the yoke of the king of Babylon, I will punish that nation with the sword, with famine, and with pestilence, declares the LORD, until I have consumed it by his hand.
JER|27|9|So do not listen to your prophets, your diviners, your dreamers, your fortunetellers, or your sorcerers, who are saying to you, 'You shall not serve the king of Babylon.'
JER|27|10|For it is a lie that they are prophesying to you, with the result that you will be removed far from your land, and I will drive you out, and you will perish.
JER|27|11|But any nation that will bring its neck under the yoke of the king of Babylon and serve him, I will leave on its own land, to work it and dwell there, declares the LORD."'"
JER|27|12|To Zedekiah king of Judah I spoke in like manner: "Bring your necks under the yoke of the king of Babylon, and serve him and his people and live.
JER|27|13|Why will you and your people die by the sword, by famine, and by pestilence, as the LORD has spoken concerning any nation that will not serve the king of Babylon?
JER|27|14|Do not listen to the words of the prophets who are saying to you, 'You shall not serve the king of Babylon,' for it is a lie that they are prophesying to you.
JER|27|15|I have not sent them, declares the LORD, but they are prophesying falsely in my name, with the result that I will drive you out and you will perish, you and the prophets who are prophesying to you."
JER|27|16|Then I spoke to the priests and to all this people, saying, "Thus says the LORD: Do not listen to the words of your prophets who are prophesying to you, saying, 'Behold, the vessels of the LORD's house will now shortly be brought back from Babylon,' for it is a lie that they are prophesying to you.
JER|27|17|Do not listen to them; serve the king of Babylon and live. Why should this city become a desolation?
JER|27|18|If they are prophets, and if the word of the LORD is with them, then let them intercede with the LORD of hosts, that the vessels that are left in the house of the LORD, in the house of the king of Judah, and in Jerusalem may not go to Babylon.
JER|27|19|For thus says the LORD of hosts concerning the pillars, the sea, the stands, and the rest of the vessels that are left in this city,
JER|27|20|which Nebuchadnezzar king of Babylon did not take away, when he took into exile from Jerusalem to Babylon Jeconiah the son of Jehoiakim, king of Judah, and all the nobles of Judah and Jerusalem-
JER|27|21|thus says the LORD of hosts, the God of Israel, concerning the vessels that are left in the house of the LORD, in the house of the king of Judah, and in Jerusalem:
JER|27|22|They shall be carried to Babylon and remain there until the day when I visit them, declares the LORD. Then I will bring them back and restore them to this place."
JER|28|1|In that same year, at the beginning of the reign of Zedekiah king of Judah, in the fifth month of the fourth year, Hananiah the son of Azzur, the prophet from Gibeon, spoke to me in the house of the LORD, in the presence of the priests and all the people, saying,
JER|28|2|"Thus says the LORD of hosts, the God of Israel: I have broken the yoke of the king of Babylon.
JER|28|3|Within two years I will bring back to this place all the vessels of the LORD's house, which Nebuchadnezzar king of Babylon took away from this place and carried to Babylon.
JER|28|4|I will also bring back to this place Jeconiah the son of Jehoiakim, king of Judah, and all the exiles from Judah who went to Babylon, declares the LORD, for I will break the yoke of the king of Babylon."
JER|28|5|Then the prophet Jeremiah spoke to Hananiah the prophet in the presence of the priests and all the people who were standing in the house of the LORD,
JER|28|6|and the prophet Jeremiah said, "Amen! May the LORD do so; may the LORD make the words that you have prophesied come true, and bring back to this place from Babylon the vessels of the house of the LORD, and all the exiles.
JER|28|7|Yet hear now this word that I speak in your hearing and in the hearing of all the people.
JER|28|8|The prophets who preceded you and me from ancient times prophesied war, famine, and pestilence against many countries and great kingdoms.
JER|28|9|As for the prophet who prophesies peace, when the word of that prophet comes to pass, then it will be known that the LORD has truly sent the prophet."
JER|28|10|Then the prophet Hananiah took the yoke-bars from the neck of Jeremiah the prophet and broke them.
JER|28|11|And Hananiah spoke in the presence of all the people, saying, "Thus says the LORD: Even so will I break the yoke of Nebuchadnezzar king of Babylon from the neck of all the nations within two years." But Jeremiah the prophet went his way.
JER|28|12|Sometime after the prophet Hananiah had broken the yoke-bars from off the neck of Jeremiah the prophet, the word of the LORD came to Jeremiah:
JER|28|13|"Go, tell Hananiah, 'Thus says the LORD: You have broken wooden bars, but you have made in their place bars of iron.
JER|28|14|For thus says the LORD of hosts, the God of Israel: I have put upon the neck of all these nations an iron yoke to serve Nebuchadnezzar king of Babylon, and they shall serve him, for I have given to him even the beasts of the field.'"
JER|28|15|And Jeremiah the prophet said to the prophet Hananiah, "Listen, Hananiah, the LORD has not sent you, and you have made this people trust in a lie.
JER|28|16|Therefore thus says the LORD: 'Behold, I will remove you from the face of the earth. This year you shall die, because you have uttered rebellion against the LORD.'"
JER|28|17|In that same year, in the seventh month, the prophet Hananiah died.
JER|29|1|These are the words of the letter that Jeremiah the prophet sent from Jerusalem to the surviving elders of the exiles, and to the priests, the prophets, and all the people, whom Nebuchadnezzar had taken into exile from Jerusalem to Babylon.
JER|29|2|This was after King Jeconiah and the queen mother, the eunuchs, the officials of Judah and Jerusalem, the craftsmen, and the metal workers had departed from Jerusalem.
JER|29|3|The letter was sent by the hand of Elasah the son of Shaphan and Gemariah the son of Hilkiah, whom Zedekiah king of Judah sent to Babylon to Nebuchadnezzar king of Babylon. It said:
JER|29|4|"Thus says the LORD of hosts, the God of Israel, to all the exiles whom I have sent into exile from Jerusalem to Babylon:
JER|29|5|Build houses and live in them; plant gardens and eat their produce.
JER|29|6|Take wives and have sons and daughters; take wives for your sons, and give your daughters in marriage, that they may bear sons and daughters; multiply there, and do not decrease.
JER|29|7|But seek the welfare of the city where I have sent you into exile, and pray to the LORD on its behalf, for in its welfare you will find your welfare.
JER|29|8|For thus says the LORD of hosts, the God of Israel: Do not let your prophets and your diviners who are among you deceive you, and do not listen to the dreams that they dream,
JER|29|9|for it is a lie that they are prophesying to you in my name; I did not send them, declares the LORD.
JER|29|10|"For thus says the LORD: When seventy years are completed for Babylon, I will visit you, and I will fulfill to you my promise and bring you back to this place.
JER|29|11|For I know the plans I have for you, declares the LORD, plans for wholeness and not for evil, to give you a future and a hope.
JER|29|12|Then you will call upon me and come and pray to me, and I will hear you.
JER|29|13|You will seek me and find me. When you seek me with all your heart,
JER|29|14|I will be found by you, declares the LORD, and I will restore your fortunes and gather you from all the nations and all the places where I have driven you, declares the LORD, and I will bring you back to the place from which I sent you into exile.
JER|29|15|"Because you have said, 'The LORD has raised up prophets for us in Babylon,'
JER|29|16|thus says the LORD concerning the king who sits on the throne of David, and concerning all the people who dwell in this city, your kinsmen who did not go out with you into exile:
JER|29|17|'Thus says the LORD of hosts, behold, I am sending on them sword, famine, and pestilence, and I will make them like vile figs that are so rotten they cannot be eaten.
JER|29|18|I will pursue them with sword, famine, and pestilence, and will make them a horror to all the kingdoms of the earth, to be a curse, a terror, a hissing, and a reproach among all the nations where I have driven them,
JER|29|19|because they did not pay attention to my words, declares the LORD, that I persistently sent to you by my servants the prophets, but you would not listen, declares the LORD.'
JER|29|20|Hear the word of the LORD, all you exiles whom I sent away from Jerusalem to Babylon:
JER|29|21|'Thus says the LORD of hosts, the God of Israel, concerning Ahab the son of Kolaiah and Zedekiah the son of Maaseiah, who are prophesying a lie to you in my name: Behold, I will deliver them into the hand of Nebuchadnezzar king of Babylon, and he shall strike them down before your eyes.
JER|29|22|Because of them this curse shall be used by all the exiles from Judah in Babylon: "The LORD make you like Zedekiah and Ahab, whom the king of Babylon roasted in the fire,"
JER|29|23|because they have done an outrageous thing in Israel, they have committed adultery with their neighbors' wives, and they have spoken in my name lying words that I did not command them. I am the one who knows, and I am witness, declares the LORD.'"
JER|29|24|To Shemaiah of Nehelam you shall say:
JER|29|25|"Thus says the LORD of hosts, the God of Israel: You have sent letters in your name to all the people who are in Jerusalem, and to Zephaniah the son of Maaseiah the priest, and to all the priests, saying,
JER|29|26|'The LORD has made you priest instead of Jehoiada the priest, to have charge in the house of the LORD over every madman who prophesies, to put him in the stocks and neck irons.
JER|29|27|Now why have you not rebuked Jeremiah of Anathoth who is prophesying to you?
JER|29|28|For he has sent to us in Babylon, saying, "Your exile will be long; build houses and live in them, and plant gardens and eat their produce."'"
JER|29|29|Zephaniah the priest read this letter in the hearing of Jeremiah the prophet.
JER|29|30|Then the word of the LORD came to Jeremiah:
JER|29|31|"Send to all the exiles, saying, 'Thus says the LORD concerning Shemaiah of Nehelam: Because Shemaiah had prophesied to you when I did not send him, and has made you trust in a lie,
JER|29|32|therefore thus says the LORD: Behold, I will punish Shemaiah of Nehelam and his descendants. He shall not have anyone living among this people, and he shall not see the good that I will do to my people, declares the LORD, for he has spoken rebellion against the LORD.'"
JER|30|1|The word that came to Jeremiah from the LORD:
JER|30|2|"Thus says the LORD, the God of Israel: Write in a book all the words that I have spoken to you.
JER|30|3|For behold, days are coming, declares the LORD, when I will restore the fortunes of my people, Israel and Judah, says the LORD, and I will bring them back to the land that I gave to their fathers, and they shall take possession of it."
JER|30|4|These are the words that the LORD spoke concerning Israel and Judah:
JER|30|5|"Thus says the LORD: We have heard a cry of panic, of terror, and no peace.
JER|30|6|Ask now, and see, can a man bear a child? Why then do I see every man with his hands on his stomach like a woman in labor? Why has every face turned pale?
JER|30|7|Alas! That day is so great there is none like it; it is a time of distress for Jacob; yet he shall be saved out of it.
JER|30|8|"And it shall come to pass in that day, declares the LORD of hosts, that I will break his yoke from off your neck, and I will burst your bonds, and foreigners shall no more make a servant of him.
JER|30|9|But they shall serve the LORD their God and David their king, whom I will raise up for them.
JER|30|10|"Then fear not, O Jacob my servant, declares the LORD, nor be dismayed, O Israel; for behold, I will save you from far away, and your offspring from the land of their captivity. Jacob shall return and have quiet and ease, and none shall make him afraid.
JER|30|11|For I am with you to save you, declares the LORD; I will make a full end of all the nations among whom I scattered you, but of you I will not make a full end. I will discipline you in just measure, and I will by no means leave you unpunished.
JER|30|12|"For thus says the LORD: Your hurt is incurable, and your wound is grievous.
JER|30|13|There is none to uphold your cause, no medicine for your wound, no healing for you.
JER|30|14|All your lovers have forgotten you; they care nothing for you; for I have dealt you the blow of an enemy, the punishment of a merciless foe, because your guilt is great, because your sins are flagrant.
JER|30|15|Why do you cry out over your hurt? Your pain is incurable. Because your guilt is great, because your sins are flagrant, I have done these things to you.
JER|30|16|Therefore all who devour you shall be devoured, and all your foes, every one of them, shall go into captivity; those who plunder you shall be plundered, and all who prey on you I will make a prey.
JER|30|17|For I will restore health to you, and your wounds I will heal, declares the LORD, because they have called you an outcast: 'It is Zion, for whom no one cares!'
JER|30|18|"Thus says the LORD: Behold, I will restore the fortunes of the tents of Jacob and have compassion on his dwellings; the city shall be rebuilt on its mound, and the palace shall stand where it used to be.
JER|30|19|Out of them shall come songs of thanksgiving, and the voices of those who celebrate. I will multiply them, and they shall not be few; I will make them honored, and they shall not be small.
JER|30|20|Their children shall be as they were of old, and their congregation shall be established before me, and I will punish all who oppress them.
JER|30|21|Their prince shall be one of themselves; their ruler shall come out from their midst; I will make him draw near, and he shall approach me, for who would dare of himself to approach me? declares the LORD.
JER|30|22|And you shall be my people, and I will be your God."
JER|30|23|Behold the storm of the LORD! Wrath has gone forth, a whirling tempest; it will burst upon the head of the wicked.
JER|30|24|The fierce anger of the LORD will not turn back until he has executed and accomplished the intentions of his mind. In the latter days you will understand this.
JER|31|1|"At that time, declares the LORD, I will be the God of all the clans of Israel, and they shall be my people."
JER|31|2|Thus says the LORD: "The people who survived the sword found grace in the wilderness; when Israel sought for rest,
JER|31|3|the LORD appeared to him from far away. I have loved you with an everlasting love; therefore I have continued my faithfulness to you.
JER|31|4|Again I will build you, and you shall be built, O virgin Israel! Again you shall adorn yourself with tambourines and shall go forth in the dance of the merrymakers.
JER|31|5|Again you shall plant vineyards on the mountains of Samaria; the planters shall plant and shall enjoy the fruit.
JER|31|6|For there shall be a day when watchmen will call in the hill country of Ephraim: 'Arise, and let us go up to Zion, to the LORD our God.'"
JER|31|7|For thus says the LORD: "Sing aloud with gladness for Jacob, and raise shouts for the chief of the nations; proclaim, give praise, and say, 'O LORD, save your people, the remnant of Israel.'
JER|31|8|Behold, I will bring them from the north country and gather them from the farthest parts of the earth, among them the blind and the lame, the pregnant woman and her who is in labor, together; a great company, they shall return here.
JER|31|9|With weeping they shall come, and with pleas for mercy I will lead them back, I will make them walk by brooks of water, in a straight path in which they shall not stumble, for I am a father to Israel, and Ephraim is my firstborn.
JER|31|10|"Hear the word of the LORD, O nations, and declare it in the coastlands far away; say, 'He who scattered Israel will gather him, and will keep him as a shepherd keeps his flock.'
JER|31|11|For the LORD has ransomed Jacob and has redeemed him from hands too strong for him.
JER|31|12|They shall come and sing aloud on the height of Zion, and they shall be radiant over the goodness of the LORD, over the grain, the wine, and the oil, and over the young of the flock and the herd; their life shall be like a watered garden, and they shall languish no more.
JER|31|13|Then shall the young women rejoice in the dance, and the young men and the old shall be merry. I will turn their mourning into joy; I will comfort them, and give them gladness for sorrow.
JER|31|14|I will feast the soul of the priests with abundance, and my people shall be satisfied with my goodness, declares the LORD."
JER|31|15|Thus says the LORD: "A voice is heard in Ramah, lamentation and bitter weeping. Rachel is weeping for her children; she refuses to be comforted for her children, because they are no more."
JER|31|16|Thus says the LORD: "Keep your voice from weeping, and your eyes from tears, for there is a reward for your work, declares the LORD, and they shall come back from the land of the enemy.
JER|31|17|There is hope for your future, declares the LORD, and your children shall come back to their own country.
JER|31|18|I have heard Ephraim grieving, 'You have disciplined me, and I was disciplined, like an untrained calf; bring me back that I may be restored, for you are the LORD my God.
JER|31|19|For after I had turned away, I relented, and after I was instructed, I slapped my thigh; I was ashamed, and I was confounded, because I bore the disgrace of my youth.'
JER|31|20|Is Ephraim my dear son? Is he my darling child? For as often as I speak against him, I do remember him still. Therefore my heart yearns for him; I will surely have mercy on him, declares the LORD.
JER|31|21|"Set up road markers for yourself; make yourself guideposts; consider well the highway, the road by which you went. Return, O virgin Israel, return to these your cities.
JER|31|22|How long will you waver, O faithless daughter? For the LORD has created a new thing on the earth: a woman encircles a man."
JER|31|23|Thus says the LORD of hosts, the God of Israel: "Once more they shall use these words in the land of Judah and in its cities, when I restore their fortunes: "' The LORD bless you, O habitation of righteousness, O holy hill!'
JER|31|24|And Judah and all its cities shall dwell there together, and the farmers and those who wander with their flocks.
JER|31|25|For I will satisfy the weary soul, and every languishing soul I will replenish."
JER|31|26|At this I awoke and looked, and my sleep was pleasant to me.
JER|31|27|"Behold, the days are coming, declares the LORD, when I will sow the house of Israel and the house of Judah with the seed of man and the seed of beast.
JER|31|28|And it shall come to pass that as I have watched over them to pluck up and break down, to overthrow, destroy, and bring harm, so I will watch over them to build and to plant, declares the LORD.
JER|31|29|In those days they shall no longer say: "' The fathers have eaten sour grapes, and the children's teeth are set on edge.'
JER|31|30|But everyone shall die for his own sin. Each man who eats sour grapes, his teeth shall be set on edge.
JER|31|31|"Behold, the days are coming, declares the LORD, when I will make a new covenant with the house of Israel and the house of Judah,
JER|31|32|not like the covenant that I made with their fathers on the day when I took them by the hand to bring them out of the land of Egypt, my covenant that they broke, though I was their husband, declares the LORD.
JER|31|33|But this is the covenant that I will make with the house of Israel after those days, declares the LORD: I will put my law within them, and I will write it on their hearts. And I will be their God, and they shall be my people.
JER|31|34|And no longer shall each one teach his neighbor and each his brother, saying, 'Know the LORD,' for they shall all know me, from the least of them to the greatest, declares the LORD. For I will forgive their iniquity, and I will remember their sin no more."
JER|31|35|Thus says the LORD, who gives the sun for light by day and the fixed order of the moon and the stars for light by night, who stirs up the sea so that its waves roar- the LORD of hosts is his name:
JER|31|36|"If this fixed order departs from before me, declares the LORD, then shall the offspring of Israel cease from being a nation before me forever."
JER|31|37|Thus says the LORD: "If the heavens above can be measured, and the foundations of the earth below can be explored, then I will cast off all the offspring of Israel for all that they have done, declares the LORD."
JER|31|38|"Behold, the days are coming, declares the LORD, when the city shall be rebuilt for the LORD from the tower of Hananel to the Corner Gate.
JER|31|39|And the measuring line shall go out farther, straight to the hill Gareb, and shall then turn to Goah.
JER|31|40|The whole valley of the dead bodies and the ashes, and all the fields as far as the brook Kidron, to the corner of the Horse Gate toward the east, shall be sacred to the LORD. It shall not be uprooted or overthrown anymore forever."
JER|32|1|The word that came to Jeremiah from the LORD in the tenth year of Zedekiah king of Judah, which was the eighteenth year of Nebuchadnezzar.
JER|32|2|At that time the army of the king of Babylon was besieging Jerusalem, and Jeremiah the prophet was shut up in the court of the guard that was in the palace of the king of Judah.
JER|32|3|For Zedekiah king of Judah had imprisoned him, saying, "Why do you prophesy and say, 'Thus says the LORD: Behold, I am giving this city into the hand of the king of Babylon, and he shall capture it;
JER|32|4|Zedekiah king of Judah shall not escape out of the hand of the Chaldeans, but shall surely be given into the hand of the king of Babylon, and shall speak with him face to face and see him eye to eye.
JER|32|5|And he shall take Zedekiah to Babylon, and there he shall remain until I visit him, declares the LORD. Though you fight against the Chaldeans, you shall not succeed'?"
JER|32|6|Jeremiah said, "The word of the LORD came to me:
JER|32|7|Behold, Hanamel the son of Shallum your uncle will come to you and say, 'Buy my field that is at Anathoth, for the right of redemption by purchase is yours.'
JER|32|8|Then Hanamel my cousin came to me in the court of the guard, in accordance with the word of the LORD, and said to me, 'Buy my field that is at Anathoth in the land of Benjamin, for the right of possession and redemption is yours; buy it for yourself.' Then I knew that this was the word of the LORD.
JER|32|9|"And I bought the field at Anathoth from Hanamel my cousin, and weighed out the money to him, seventeen shekels of silver.
JER|32|10|I signed the deed, sealed it, got witnesses, and weighed the money on scales.
JER|32|11|Then I took the sealed deed of purchase, containing the terms and conditions and the open copy.
JER|32|12|And I gave the deed of purchase to Baruch the son of Neriah son of Mahseiah, in the presence of Hanamel my cousin, in the presence of the witnesses who signed the deed of purchase, and in the presence of all the Judeans who were sitting in the court of the guard.
JER|32|13|I charged Baruch in their presence, saying,
JER|32|14|'Thus says the LORD of hosts, the God of Israel: Take these deeds, both this sealed deed of purchase and this open deed, and put them in an earthenware vessel, that they may last for a long time.
JER|32|15|For thus says the LORD of hosts, the God of Israel: Houses and fields and vineyards shall again be bought in this land.'
JER|32|16|"After I had given the deed of purchase to Baruch the son of Neriah, I prayed to the LORD, saying:
JER|32|17|'Ah, Lord GOD! It is you who has made the heavens and the earth by your great power and by your outstretched arm! Nothing is too hard for you.
JER|32|18|You show steadfast love to thousands, but you repay the guilt of fathers to their children after them, O great and mighty God, whose name is the LORD of hosts,
JER|32|19|great in counsel and mighty in deed, whose eyes are open to all the ways of the children of man, rewarding each one according to his ways and according to the fruit of his deeds.
JER|32|20|You have shown signs and wonders in the land of Egypt, and to this day in Israel and among all mankind, and have made a name for yourself, as at this day.
JER|32|21|You brought your people Israel out of the land of Egypt with signs and wonders, with a strong hand and outstretched arm, and with great terror.
JER|32|22|And you gave them this land, which you swore to their fathers to give them, a land flowing with milk and honey.
JER|32|23|And they entered and took possession of it. But they did not obey your voice or walk in your law. They did nothing of all you commanded them to do. Therefore you have made all this disaster come upon them.
JER|32|24|Behold, the siege mounds have come up to the city to take it, and because of sword and famine and pestilence the city is given into the hands of the Chaldeans who are fighting against it. What you spoke has come to pass, and behold, you see it.
JER|32|25|Yet you, O Lord GOD, have said to me, "Buy the field for money and get witnesses"- though the city is given into the hands of the Chaldeans.'"
JER|32|26|The word of the LORD came to Jeremiah:
JER|32|27|"Behold, I am the LORD, the God of all flesh. Is anything too hard for me?
JER|32|28|Therefore, thus says the LORD: Behold, I am giving this city into the hands of the Chaldeans and into the hand of Nebuchadnezzar king of Babylon, and he shall capture it.
JER|32|29|The Chaldeans who are fighting against this city shall come and set this city on fire and burn it, with the houses on whose roofs offerings have been made to Baal and drink offerings have been poured out to other gods, to provoke me to anger.
JER|32|30|For the children of Israel and the children of Judah have done nothing but evil in my sight from their youth. The children of Israel have done nothing but provoke me to anger by the work of their hands, declares the LORD.
JER|32|31|This city has aroused my anger and wrath, from the day it was built to this day, so that I will remove it from my sight
JER|32|32|because of all the evil of the children of Israel and the children of Judah that they did to provoke me to anger- their kings and their officials, their priests and their prophets, the men of Judah and the inhabitants of Jerusalem.
JER|32|33|They have turned to me their back and not their face. And though I have taught them persistently, they have not listened to receive instruction.
JER|32|34|They set up their abominations in the house that is called by my name, to defile it.
JER|32|35|They built the high places of Baal in the Valley of the Son of Hinnom, to offer up their sons and daughters to Molech, though I did not command them, nor did it enter into my mind, that they should do this abomination, to cause Judah to sin.
JER|32|36|"Now therefore thus says the LORD, the God of Israel, concerning this city of which you say, 'It is given into the hand of the king of Babylon by sword, by famine, and by pestilence':
JER|32|37|Behold, I will gather them from all the countries to which I drove them in my anger and my wrath and in great indignation. I will bring them back to this place, and I will make them dwell in safety.
JER|32|38|And they shall be my people, and I will be their God.
JER|32|39|I will give them one heart and one way, that they may fear me forever, for their own good and the good of their children after them.
JER|32|40|I will make with them an everlasting covenant, that I will not turn away from doing good to them. And I will put the fear of me in their hearts, that they may not turn from me.
JER|32|41|I will rejoice in doing them good, and I will plant them in this land in faithfulness, with all my heart and all my soul.
JER|32|42|"For thus says the LORD: Just as I have brought all this great disaster upon this people, so I will bring upon them all the good that I promise them.
JER|32|43|Fields shall be bought in this land of which you are saying, 'It is a desolation, without man or beast; it is given into the hand of the Chaldeans.'
JER|32|44|Fields shall be bought for money, and deeds shall be signed and sealed and witnessed, in the land of Benjamin, in the places about Jerusalem, and in the cities of Judah, in the cities of the hill country, in the cities of the Shephelah, and in the cities of the Negeb; for I will restore their fortunes, declares the LORD."
JER|33|1|The word of the LORD came to Jeremiah a second time, while he was still shut up in the court of the guard:
JER|33|2|"Thus says the LORD who made the earth, the LORD who formed it to establish it- the LORD is his name:
JER|33|3|Call to me and I will answer you, and will tell you great and hidden things that you have not known.
JER|33|4|For thus says the LORD, the God of Israel, concerning the houses of this city and the houses of the kings of Judah that were torn down to make a defense against the siege mounds and against the sword:
JER|33|5|They are coming in to fight against the Chaldeans and to fill them with the dead bodies of men whom I shall strike down in my anger and my wrath, for I have hidden my face from this city because of all their evil.
JER|33|6|Behold, I will bring to it health and healing, and I will heal them and reveal to them abundance of prosperity and security.
JER|33|7|I will restore the fortunes of Judah and the fortunes of Israel, and rebuild them as they were at first.
JER|33|8|I will cleanse them from all the guilt of their sin against me, and I will forgive all the guilt of their sin and rebellion against me.
JER|33|9|And this city shall be to me a name of joy, a praise and a glory before all the nations of the earth who shall hear of all the good that I do for them. They shall fear and tremble because of all the good and all the prosperity I provide for it.
JER|33|10|"Thus says the LORD: In this place of which you say, 'It is a waste without man or beast,' in the cities of Judah and the streets of Jerusalem that are desolate, without man or inhabitant or beast, there shall be heard again
JER|33|11|the voice of mirth and the voice of gladness, the voice of the bridegroom and the voice of the bride, the voices of those who sing, as they bring thank offerings to the house of the LORD: "' Give thanks to the LORD of hosts, for the LORD is good, for his steadfast love endures forever!' For I will restore the fortunes of the land as at first, says the LORD.
JER|33|12|"Thus says the LORD of hosts: In this place that is waste, without man or beast, and in all of its cities, there shall again be habitations of shepherds resting their flocks.
JER|33|13|In the cities of the hill country, in the cities of the Shephelah, and in the cities of the Negeb, in the land of Benjamin, the places about Jerusalem, and in the cities of Judah, flocks shall again pass under the hands of the one who counts them, says the LORD.
JER|33|14|"Behold, the days are coming, declares the LORD, when I will fulfill the promise I made to the house of Israel and the house of Judah.
JER|33|15|In those days and at that time I will cause a righteous Branch to spring up for David, and he shall execute justice and righteousness in the land.
JER|33|16|In those days Judah will be saved and Jerusalem will dwell securely. And this is the name by which it will be called: 'The LORD is our righteousness.'
JER|33|17|"For thus says the LORD: David shall never lack a man to sit on the throne of the house of Israel,
JER|33|18|and the Levitical priests shall never lack a man in my presence to offer burnt offerings, to burn grain offerings, and to make sacrifices forever."
JER|33|19|The word of the LORD came to Jeremiah:
JER|33|20|"Thus says the LORD: If you can break my covenant with the day and my covenant with the night, so that day and night will not come at their appointed time,
JER|33|21|then also my covenant with David my servant may be broken, so that he shall not have a son to reign on his throne, and my covenant with the Levitical priests my ministers.
JER|33|22|As the host of heaven cannot be numbered and the sands of the sea cannot be measured, so I will multiply the offspring of David my servant, and the Levitical priests who minister to me."
JER|33|23|The word of the LORD came to Jeremiah:
JER|33|24|"Have you not observed that these people are saying, 'The LORD has rejected the two clans that he chose'? Thus they have despised my people so that they are no longer a nation in their sight.
JER|33|25|Thus says the LORD: If I have not established my covenant with day and night and the fixed order of heaven and earth,
JER|33|26|then I will reject the offspring of Jacob and David my servant and will not choose one of his offspring to rule over the offspring of Abraham, Isaac, and Jacob. For I will restore their fortunes and will have mercy on them."
JER|34|1|The word that came to Jeremiah from the LORD, when Nebuchadnezzar king of Babylon and all his army and all the kingdoms of the earth under his dominion and all the peoples were fighting against Jerusalem and all of its cities:
JER|34|2|"Thus says the LORD, the God of Israel: Go and speak to Zedekiah king of Judah and say to him, 'Thus says the LORD: Behold, I am giving this city into the hand of the king of Babylon, and he shall burn it with fire.
JER|34|3|You shall not escape from his hand but shall surely be captured and delivered into his hand. You shall see the king of Babylon eye to eye and speak with him face to face. And you shall go to Babylon.'
JER|34|4|Yet hear the word of the LORD, O Zedekiah king of Judah! Thus says the LORD concerning you: 'You shall not die by the sword.
JER|34|5|You shall die in peace. And as spices were burned for your fathers, the former kings who were before you, so people shall burn spices for you and lament for you, saying, "Alas, lord!"'For I have spoken the word, declares the LORD."
JER|34|6|Then Jeremiah the prophet spoke all these words to Zedekiah king of Judah, in Jerusalem,
JER|34|7|when the army of the king of Babylon was fighting against Jerusalem and against all the cities of Judah that were left, Lachish and Azekah, for these were the only fortified cities of Judah that remained.
JER|34|8|The word that came to Jeremiah from the LORD, after King Zedekiah had made a covenant with all the people in Jerusalem to make a proclamation of liberty to them,
JER|34|9|that everyone should set free his Hebrew slaves, male and female, so that no one should enslave a Jew, his brother.
JER|34|10|And they obeyed, all the officials and all the people who had entered into the covenant that everyone would set free his slave, male or female, so that they would not be enslaved again. They obeyed and set them free.
JER|34|11|But afterward they turned around and took back the male and female slaves they had set free, and brought them into subjection as slaves.
JER|34|12|The word of the LORD came to Jeremiah from the LORD:
JER|34|13|"Thus says the LORD, the God of Israel: I myself made a covenant with your fathers when I brought them out of the land of Egypt, out of the house of bondage, saying,
JER|34|14|'At the end of seven years each of you must set free the fellow Hebrew who has been sold to you and has served you six years; you must set him free from your service.' But your fathers did not listen to me or incline their ears to me.
JER|34|15|You recently repented and did what was right in my eyes by proclaiming liberty, each to his neighbor, and you made a covenant before me in the house that is called by my name,
JER|34|16|but then you turned around and profaned my name when each of you took back his male and female slaves, whom you had set free according to their desire, and you brought them into subjection to be your slaves.
JER|34|17|"Therefore, thus says the LORD: You have not obeyed me by proclaiming liberty, every one to his brother and to his neighbor; behold, I proclaim to you liberty to the sword, to pestilence, and to famine, declares the LORD. I will make you a horror to all the kingdoms of the earth.
JER|34|18|And the men who transgressed my covenant and did not keep the terms of the covenant that they made before me, I will make them like the calf that they cut in two and passed between its parts-
JER|34|19|the officials of Judah, the officials of Jerusalem, the eunuchs, the priests, and all the people of the land who passed between the parts of the calf.
JER|34|20|And I will give them into the hand of their enemies and into the hand of those who seek their lives. Their dead bodies shall be food for the birds of the air and the beasts of the earth.
JER|34|21|And Zedekiah king of Judah and his officials I will give into the hand of their enemies and into the hand of those who seek their lives, into the hand of the army of the king of Babylon which has withdrawn from you.
JER|34|22|Behold, I will command, declares the LORD, and will bring them back to this city. And they will fight against it and take it and burn it with fire. I will make the cities of Judah a desolation without inhabitant."
JER|35|1|The word that came to Jeremiah from the LORD in the days of Jehoiakim the son of Josiah, king of Judah:
JER|35|2|"Go to the house of the Rechabites and speak with them and bring them to the house of the LORD, into one of the chambers; then offer them wine to drink."
JER|35|3|So I took Jaazaniah the son of Jeremiah, son of Habazziniah and his brothers and all his sons and the whole house of the Rechabites.
JER|35|4|I brought them to the house of the LORD into the chamber of the sons of Hanan the son of Igdaliah, the man of God, which was near the chamber of the officials, above the chamber of Maaseiah the son of Shallum, keeper of the threshold.
JER|35|5|Then I set before the Rechabites pitchers full of wine, and cups, and I said to them, "Drink wine."
JER|35|6|But they answered, "We will drink no wine, for Jonadab the son of Rechab, our father, commanded us, 'You shall not drink wine, neither you nor your sons forever.
JER|35|7|You shall not build a house; you shall not sow seed; you shall not plant or have a vineyard; but you shall live in tents all your days, that you may live many days in the land where you sojourn.'
JER|35|8|We have obeyed the voice of Jonadab the son of Rechab, our father, in all that he commanded us, to drink no wine all our days, ourselves, our wives, our sons, or our daughters,
JER|35|9|and not to build houses to dwell in. We have no vineyard or field or seed,
JER|35|10|but we have lived in tents and have obeyed and done all that Jonadab our father commanded us.
JER|35|11|But when Nebuchadnezzar king of Babylon came up against the land, we said, 'Come, and let us go to Jerusalem for fear of the army of the Chaldeans and the army of the Syrians.' So we are living in Jerusalem."
JER|35|12|Then the word of the LORD came to Jeremiah:
JER|35|13|"Thus says the LORD of hosts, the God of Israel: Go and say to the people of Judah and the inhabitants of Jerusalem, Will you not receive instruction and listen to my words? declares the LORD.
JER|35|14|The command that Jonadab the son of Rechab gave to his sons, to drink no wine, has been kept, and they drink none to this day, for they have obeyed their father's command. I have spoken to you persistently, but you have not listened to me.
JER|35|15|I have sent to you all my servants the prophets, sending them persistently, saying, 'Turn now every one of you from his evil way, and amend your deeds, and do not go after other gods to serve them, and then you shall dwell in the land that I gave to you and your fathers.' But you did not incline your ear or listen to me.
JER|35|16|The sons of Jonadab the son of Rechab have kept the command that their father gave them, but this people has not obeyed me.
JER|35|17|Therefore, thus says the LORD, the God of hosts, the God of Israel: Behold, I am bringing upon Judah and all the inhabitants of Jerusalem all the disaster that I have pronounced against them, because I have spoken to them and they have not listened, I have called to them and they have not answered."
JER|35|18|But to the house of the Rechabites Jeremiah said, "Thus says the LORD of hosts, the God of Israel: Because you have obeyed the command of Jonadab your father and kept all his precepts and done all that he commanded you,
JER|35|19|therefore thus says the LORD of hosts, the God of Israel: Jonadab the son of Rechab shall never lack a man to stand before me."
JER|36|1|In the fourth year of Jehoiakim the son of Josiah, king of Judah, this word came to Jeremiah from the LORD:
JER|36|2|"Take a scroll and write on it all the words that I have spoken to you against Israel and Judah and all the nations, from the day I spoke to you, from the days of Josiah until today.
JER|36|3|It may be that the house of Judah will hear all the disaster that I intend to do to them, so that every one may turn from his evil way, and that I may forgive their iniquity and their sin."
JER|36|4|Then Jeremiah called Baruch the son of Neriah, and Baruch wrote on a scroll at the dictation of Jeremiah all the words of the LORD that he had spoken to him.
JER|36|5|And Jeremiah ordered Baruch, saying, "I am banned from going to the house of the LORD,
JER|36|6|so you are to go, and on a day of fasting in the hearing of all the people in the LORD's house you shall read the words of the LORD from the scroll that you have written at my dictation. You shall read them also in the hearing of all the men of Judah who come out of their cities.
JER|36|7|It may be that their plea for mercy will come before the LORD, and that every one will turn from his evil way, for great is the anger and wrath that the LORD has pronounced against this people."
JER|36|8|And Baruch the son of Neriah did all that Jeremiah the prophet ordered him about reading from the scroll the words of the LORD in the LORD's house.
JER|36|9|In the fifth year of Jehoiakim the son of Josiah, king of Judah, in the ninth month, all the people in Jerusalem and all the people who came from the cities of Judah to Jerusalem proclaimed a fast before the LORD.
JER|36|10|Then, in the hearing of all the people, Baruch read the words of Jeremiah from the scroll, in the house of the LORD, in the chamber of Gemariah the son of Shaphan the secretary, which was in the upper court, at the entry of the New Gate of the LORD's house.
JER|36|11|When Micaiah the son of Gemariah, son of Shaphan, heard all the words of the LORD from the scroll,
JER|36|12|he went down to the king's house, into the secretary's chamber, and all the officials were sitting there: Elishama the secretary, Delaiah the son of Shemaiah, Elnathan the son of Achbor, Gemariah the son of Shaphan, Zedekiah the son of Hananiah, and all the officials.
JER|36|13|And Micaiah told them all the words that he had heard, when Baruch read the scroll in the hearing of the people.
JER|36|14|Then all the officials sent Jehudi the son of Nethaniah, son of Shelemiah, son of Cushi, to say to Baruch, "Take in your hand the scroll that you read in the hearing of the people, and come." So Baruch the son of Neriah took the scroll in his hand and came to them.
JER|36|15|And they said to him, "Sit down and read it." So Baruch read it to them.
JER|36|16|When they heard all the words, they turned one to another in fear. And they said to Baruch, "We must report all these words to the king."
JER|36|17|Then they asked Baruch, "Tell us, please, how did you write all these words? Was it at his dictation?"
JER|36|18|Baruch answered them, "He dictated all these words to me, while I wrote them with ink on the scroll."
JER|36|19|Then the officials said to Baruch, "Go and hide, you and Jeremiah, and let no one know where you are."
JER|36|20|So they went into the court to the king, having put the scroll in the chamber of Elishama the secretary, and they reported all the words to the king.
JER|36|21|Then the king sent Jehudi to get the scroll, and he took it from the chamber of Elishama the secretary. And Jehudi read it to the king and all the officials who stood beside the king.
JER|36|22|It was the ninth month, and the king was sitting in the winter house, and there was a fire burning in the fire pot before him.
JER|36|23|As Jehudi read three or four columns, the king would cut them off with a knife and throw them into the fire in the fire pot, until the entire scroll was consumed in the fire that was in the fire pot.
JER|36|24|Yet neither the king nor any of his servants who heard all these words was afraid, nor did they tear their garments.
JER|36|25|Even when Elnathan and Delaiah and Gemariah urged the king not to burn the scroll, he would not listen to them.
JER|36|26|And the king commanded Jerahmeel the king's son and Seraiah the son of Azriel and Shelemiah the son of Abdeel to seize Baruch the secretary and Jeremiah the prophet, but the LORD hid them.
JER|36|27|Now after the king had burned the scroll with the words that Baruch wrote at Jeremiah's dictation, the word of the LORD came to Jeremiah:
JER|36|28|"Take another scroll and write on it all the former words that were in the first scroll, which Jehoiakim the king of Judah has burned.
JER|36|29|And concerning Jehoiakim king of Judah you shall say, 'Thus says the LORD, You have burned this scroll, saying, "Why have you written in it that the king of Babylon will certainly come and destroy this land, and will cut off from it man and beast?"
JER|36|30|Therefore thus says the LORD concerning Jehoiakim king of Judah: He shall have none to sit on the throne of David, and his dead body shall be cast out to the heat by day and the frost by night.
JER|36|31|And I will punish him and his offspring and his servants for their iniquity. I will bring upon them and upon the inhabitants of Jerusalem and upon the people of Judah all the disaster that I have pronounced against them, but they would not hear.'"
JER|36|32|Then Jeremiah took another scroll and gave it to Baruch the scribe, the son of Neriah, who wrote on it at the dictation of Jeremiah all the words of the scroll that Jehoiakim king of Judah had burned in the fire. And many similar words were added to them.
JER|37|1|Zedekiah the son of Josiah, whom Nebuchadnezzar king of Babylon made king in the land of Judah, reigned instead of Coniah the son of Jehoiakim.
JER|37|2|But neither he nor his servants nor the people of the land listened to the words of the LORD that he spoke through Jeremiah the prophet.
JER|37|3|King Zedekiah sent Jehucal the son of Shelemiah, and Zephaniah the priest, the son of Maaseiah, to Jeremiah the prophet, saying, "Please pray for us to the LORD our God."
JER|37|4|Now Jeremiah was still going in and out among the people, for he had not yet been put in prison.
JER|37|5|The army of Pharaoh had come out of Egypt. And when the Chaldeans who were besieging Jerusalem heard news about them, they withdrew from Jerusalem.
JER|37|6|Then the word of the LORD came to Jeremiah the prophet:
JER|37|7|"Thus says the LORD, God of Israel: Thus shall you say to the king of Judah who sent you to me to inquire of me, 'Behold, Pharaoh's army that came to help you is about to return to Egypt, to its own land.
JER|37|8|And the Chaldeans shall come back and fight against this city. They shall capture it and burn it with fire.
JER|37|9|Thus says the LORD, Do not deceive yourselves, saying, "The Chaldeans will surely go away from us," for they will not go away.
JER|37|10|For even if you should defeat the whole army of Chaldeans who are fighting against you, and there remained of them only wounded men, every man in his tent, they would rise up and burn this city with fire.'"
JER|37|11|Now when the Chaldean army had withdrawn from Jerusalem at the approach of Pharaoh's army,
JER|37|12|Jeremiah set out from Jerusalem to go to the land of Benjamin to receive his portion there among the people.
JER|37|13|When he was at the Benjamin Gate, a sentry there named Irijah the son of Shelemiah, son of Hananiah, seized Jeremiah the prophet, saying, "You are deserting to the Chaldeans."
JER|37|14|And Jeremiah said, "It is a lie; I am not deserting to the Chaldeans." But Irijah would not listen to him, and seized Jeremiah and brought him to the officials.
JER|37|15|And the officials were enraged at Jeremiah, and they beat him and imprisoned him in the house of Jonathan the secretary, for it had been made a prison.
JER|37|16|When Jeremiah had come to the dungeon cells and remained there many days,
JER|37|17|King Zedekiah sent for him and received him. The king questioned him secretly in his house and said, "Is there any word from the LORD?" Jeremiah said, "There is." Then he said, "You shall be delivered into the hand of the king of Babylon."
JER|37|18|Jeremiah also said to King Zedekiah, "What wrong have I done to you or your servants or this people, that you have put me in prison?
JER|37|19|Where are your prophets who prophesied to you, saying, 'The king of Babylon will not come against you and against this land'?
JER|37|20|Now hear, please, O my lord the king: let my humble plea come before you and do not send me back to the house of Jonathan the secretary, lest I die there."
JER|37|21|So King Zedekiah gave orders, and they committed Jeremiah to the court of the guard. And a loaf of bread was given him daily from the bakers' street, until all the bread of the city was gone. So Jeremiah remained in the court of the guard.
JER|38|1|Now Shephatiah the son of Mattan, Gedaliah the son of Pashhur, Jucal the son of Shelemiah, and Pashhur the son of Malchiah heard the words that Jeremiah was saying to all the people,
JER|38|2|"Thus says the LORD: He who stays in this city shall die by the sword, by famine, and by pestilence, but he who goes out to the Chaldeans shall live. He shall have his life as a prize of war, and live.
JER|38|3|Thus says the LORD: This city shall surely be given into the hand of the army of the king of Babylon and be taken."
JER|38|4|Then the officials said to the king, "Let this man be put to death, for he is weakening the hands of the soldiers who are left in this city, and the hands of all the people, by speaking such words to them. For this man is not seeking the welfare of this people, but their harm."
JER|38|5|King Zedekiah said, "Behold, he is in your hands, for the king can do nothing against you."
JER|38|6|So they took Jeremiah and cast him into the cistern of Malchiah, the king's son, which was in the court of the guard, letting Jeremiah down by ropes. And there was no water in the cistern, but only mud, and Jeremiah sank in the mud.
JER|38|7|When Ebed-melech the Ethiopian, a eunuch who was in the king's house, heard that they had put Jeremiah into the cistern- the king was sitting in the Benjamin Gate-
JER|38|8|Ebed-melech went from the king's house and said to the king,
JER|38|9|"My lord the king, these men have done evil in all that they did to Jeremiah the prophet by casting him into the cistern, and he will die there of hunger, for there is no bread left in the city."
JER|38|10|Then the king commanded Ebed-melech the Ethiopian, "Take three men with you from here, and lift Jeremiah the prophet out of the cistern before he dies."
JER|38|11|So Ebed-melech took the men with him and went to the house of the king, to a wardrobe in the storehouse, and took from there old rags and worn-out clothes, which he let down to Jeremiah in the cistern by ropes.
JER|38|12|Then Ebed-melech the Ethiopian said to Jeremiah, "Put the rags and clothes between your armpits and the ropes." Jeremiah did so.
JER|38|13|Then they drew Jeremiah up with ropes and lifted him out of the cistern. And Jeremiah remained in the court of the guard.
JER|38|14|King Zedekiah sent for Jeremiah the prophet and received him at the third entrance of the temple of the LORD. The king said to Jeremiah, "I will ask you a question; hide nothing from me."
JER|38|15|Jeremiah said to Zedekiah, "If I tell you, will you not surely put me to death? And if I give you counsel, you will not listen to me."
JER|38|16|Then King Zedekiah swore secretly to Jeremiah, "As the LORD lives, who made our souls, I will not put you to death or deliver you into the hand of these men who seek your life."
JER|38|17|Then Jeremiah said to Zedekiah, "Thus says the LORD, the God of hosts, the God of Israel: If you will surrender to the officials of the king of Babylon, then your life shall be spared, and this city shall not be burned with fire, and you and your house shall live.
JER|38|18|But if you do not surrender to the officials of the king of Babylon, then this city shall be given into the hand of the Chaldeans, and they shall burn it with fire, and you shall not escape from their hand."
JER|38|19|King Zedekiah said to Jeremiah, "I am afraid of the Judeans who have deserted to the Chaldeans, lest I be handed over to them and they deal cruelly with me."
JER|38|20|Jeremiah said, "You shall not be given to them. Obey now the voice of the LORD in what I say to you, and it shall be well with you, and your life shall be spared.
JER|38|21|But if you refuse to surrender, this is the vision which the LORD has shown to me:
JER|38|22|Behold, all the women left in the house of the king of Judah were being led out to the officials of the king of Babylon and were saying, "' Your trusted friends have deceived you and prevailed against you; now that your feet are sunk in the mud, they turn away from you.'
JER|38|23|All your wives and your sons shall be led out to the Chaldeans, and you yourself shall not escape from their hand, but shall be seized by the king of Babylon, and this city shall be burned with fire."
JER|38|24|Then Zedekiah said to Jeremiah, "Let no one know of these words, and you shall not die.
JER|38|25|If the officials hear that I have spoken with you and come to you and say to you, 'Tell us what you said to the king and what the king said to you; hide nothing from us and we will not put you to death,'
JER|38|26|then you shall say to them, 'I made a humble plea to the king that he would not send me back to the house of Jonathan to die there.'"
JER|38|27|Then all the officials came to Jeremiah and asked him, and he answered them as the king had instructed him. So they stopped speaking with him, for the conversation had not been overheard.
JER|38|28|And Jeremiah remained in the court of the guard until the day that Jerusalem was taken.
JER|39|1|In the ninth year of Zedekiah king of Judah, in the tenth month, Nebuchadnezzar king of Babylon and all his army came against Jerusalem and besieged it.
JER|39|2|In the eleventh year of Zedekiah, in the fourth month, on the ninth day of the month, a breach was made in the city.
JER|39|3|Then all the officials of the king of Babylon came and sat in the middle gate: Nergal-sar-ezer, Samgar-nebu, Sar-sekim the Rab-saris, Nergal-sar-ezer the Rab-mag, with all the rest of the officers of the king of Babylon.
JER|39|4|When Zedekiah king of Judah and all the soldiers saw them, they fled, going out of the city at night by way of the king's garden through the gate between the two walls; and they went toward the Arabah.
JER|39|5|But the army of the Chaldeans pursued them and overtook Zedekiah in the plains of Jericho. And when they had taken him, they brought him up to Nebuchadnezzar king of Babylon, at Riblah, in the land of Hamath; and he passed sentence on him.
JER|39|6|The king of Babylon slaughtered the sons of Zedekiah at Riblah before his eyes, and the king of Babylon slaughtered all the nobles of Judah.
JER|39|7|He put out the eyes of Zedekiah and bound him in chains to take him to Babylon.
JER|39|8|The Chaldeans burned the king's house and the house of the people, and broke down the walls of Jerusalem.
JER|39|9|Then Nebuzaradan, the captain of the guard, carried into exile to Babylon the rest of the people who were left in the city, those who had deserted to him, and the people who remained.
JER|39|10|Nebuzaradan, the captain of the guard, left in the land of Judah some of the poor people who owned nothing, and gave them vineyards and fields at the same time.
JER|39|11|Nebuchadnezzar king of Babylon gave command concerning Jeremiah through Nebuzaradan, the captain of the guard, saying,
JER|39|12|"Take him, look after him well, and do him no harm, but deal with him as he tells you."
JER|39|13|So Nebuzaradan the captain of the guard, Nebushazban the Rab-saris, Nergal-sar-ezer the Rab-mag, and all the chief officers of the king of Babylon
JER|39|14|sent and took Jeremiah from the court of the guard. They entrusted him to Gedaliah the son of Ahikam, son of Shaphan, that he should take him home. So he lived among the people.
JER|39|15|The word of the LORD came to Jeremiah while he was shut up in the court of the guard:
JER|39|16|"Go, and say to Ebed-melech the Ethiopian, 'Thus says the LORD of hosts, the God of Israel: Behold, I will fulfill my words against this city for harm and not for good, and they shall be accomplished before you on that day.
JER|39|17|But I will deliver you on that day, declares the LORD, and you shall not be given into the hand of the men of whom you are afraid.
JER|39|18|For I will surely save you, and you shall not fall by the sword, but you shall have your life as a prize of war, because you have put your trust in me, declares the LORD.'"
JER|40|1|The word that came to Jeremiah from the LORD after Nebuzaradan the captain of the guard had let him go from Ramah, when he took him bound in chains along with all the captives of Jerusalem and Judah who were being exiled to Babylon.
JER|40|2|The captain of the guard took Jeremiah and said to him, "The LORD your God pronounced this disaster against this place.
JER|40|3|The LORD has brought it about, and has done as he said. Because you sinned against the LORD and did not obey his voice, this thing has come upon you.
JER|40|4|Now, behold, I release you today from the chains on your hands. If it seems good to you to come with me to Babylon, come, and I will look after you well, but if it seems wrong to you to come with me to Babylon, do not come. See, the whole land is before you; go wherever you think it good and right to go.
JER|40|5|If you remain, then return to Gedaliah the son of Ahikam, son of Shaphan, whom the king of Babylon appointed governor of the cities of Judah, and dwell with him among the people. Or go wherever you think it right to go." So the captain of the guard gave him an allowance of food and a present, and let him go.
JER|40|6|Then Jeremiah went to Gedaliah the son of Ahikam, at Mizpah, and lived with him among the people who were left in the land.
JER|40|7|When all the captains of the forces in the open country and their men heard that the king of Babylon had appointed Gedaliah the son of Ahikam governor in the land and had committed to him men, women, and children, those of the poorest of the land who had not been taken into exile to Babylon,
JER|40|8|they went to Gedaliah at Mizpah- Ishmael the son of Nethaniah, Johanan the son of Kareah, Seraiah the son of Tanhumeth, the sons of Ephai the Netophathite, Jezaniah the son of the Maacathite, they and their men.
JER|40|9|Gedaliah the son of Ahikam, son of Shaphan, swore to them and their men, saying, "Do not be afraid to serve the Chaldeans. Dwell in the land and serve the king of Babylon, and it shall be well with you.
JER|40|10|As for me, I will dwell at Mizpah, to represent you before the Chaldeans who will come to us. But as for you, gather wine and summer fruits and oil, and store them in your vessels, and dwell in your cities that you have taken."
JER|40|11|Likewise, when all the Judeans who were in Moab and among the Ammonites and in Edom and in other lands heard that the king of Babylon had left a remnant in Judah and had appointed Gedaliah the son of Ahikam, son of Shaphan, as governor over them,
JER|40|12|then all the Judeans returned from all the places to which they had been driven and came to the land of Judah, to Gedaliah at Mizpah. And they gathered wine and summer fruits in great abundance.
JER|40|13|Now Johanan the son of Kareah and all the leaders of the forces in the open country came to Gedaliah at Mizpah
JER|40|14|and said to him, "Do you know that Baalis the king of the Ammonites has sent Ishmael the son of Nethaniah to take your life?" But Gedaliah the son of Ahikam would not believe them.
JER|40|15|Then Johanan the son of Kareah spoke secretly to Gedaliah at Mizpah, "Please let me go and strike down Ishmael the son of Nethaniah, and no one will know it. Why should he take your life, so that all the Judeans who are gathered about you would be scattered, and the remnant of Judah would perish?"
JER|40|16|But Gedaliah the son of Ahikam said to Johanan the son of Kareah, "You shall not do this thing, for you are speaking falsely of Ishmael."
JER|41|1|In the seventh month, Ishmael the son of Nethaniah, son of Elishama, of the royal family, one of the chief officers of the king, came with ten men to Gedaliah the son of Ahikam, at Mizpah. As they ate bread together there at Mizpah,
JER|41|2|Ishmael the son of Nethaniah and the ten men with him rose up and struck down Gedaliah the son of Ahikam, son of Shaphan, with the sword, and killed him, whom the king of Babylon had appointed governor in the land.
JER|41|3|Ishmael also struck down all the Judeans who were with Gedaliah at Mizpah, and the Chaldean soldiers who happened to be there.
JER|41|4|On the day after the murder of Gedaliah, before anyone knew of it,
JER|41|5|eighty men arrived from Shechem and Shiloh and Samaria, with their beards shaved and their clothes torn, and their bodies gashed, bringing grain offerings and incense to present at the temple of the LORD.
JER|41|6|And Ishmael the son of Nethaniah came out from Mizpah to meet them, weeping as he came. As he met them, he said to them, "Come in to Gedaliah the son of Ahikam."
JER|41|7|When they came into the city, Ishmael the son of Nethaniah and the men with him slaughtered them and cast them into a cistern.
JER|41|8|But there were ten men among them who said to Ishmael, "Do not put us to death, for we have stores of wheat, barley, oil, and honey hidden in the fields." So he refrained and did not put them to death with their companions.
JER|41|9|Now the cistern into which Ishmael had thrown all the bodies of the men whom he had struck down along with Gedaliah was the large cistern that King Asa had made for defense against Baasha king of Israel; Ishmael the son of Nethaniah filled it with the slain.
JER|41|10|Then Ishmael took captive all the rest of the people who were in Mizpah, the king's daughters and all the people who were left at Mizpah, whom Nebuzaradan, the captain of the guard, had committed to Gedaliah the son of Ahikam. Ishmael the son of Nethaniah took them captive and set out to cross over to the Ammonites.
JER|41|11|But when Johanan the son of Kareah and all the leaders of the forces with him heard of all the evil that Ishmael the son of Nethaniah had done,
JER|41|12|they took all their men and went to fight against Ishmael the son of Nethaniah. They came upon him at the great pool that is in Gibeon.
JER|41|13|And when all the people who were with Ishmael saw Johanan the son of Kareah and all the leaders of the forces with him, they rejoiced.
JER|41|14|So all the people whom Ishmael had carried away captive from Mizpah turned around and came back, and went to Johanan the son of Kareah.
JER|41|15|But Ishmael the son of Nethaniah escaped from Johanan with eight men, and went to the Ammonites.
JER|41|16|Then Johanan the son of Kareah and all the leaders of the forces with him took from Mizpah all the rest of the people whom he had recovered from Ishmael the son of Nethaniah, after he had struck down Gedaliah the son of Ahikam- soldiers, women, children, and eunuchs, whom Johanan brought back from Gibeon.
JER|41|17|And they went and stayed at Geruth Chimham near Bethlehem, intending to go to Egypt
JER|41|18|because of the Chaldeans. For they were afraid of them, because Ishmael the son of Nethaniah had struck down Gedaliah the son of Ahikam, whom the king of Babylon had made governor over the land.
JER|42|1|Then all the commanders of the forces, and Johanan the son of Kareah and Jezaniah the son of Hoshaiah, and all the people from the least to the greatest, came near
JER|42|2|and said to Jeremiah the prophet, "Let our plea for mercy come before you, and pray to the LORD your God for us, for all this remnant- because we are left with but a few, as your eyes see us-
JER|42|3|that the LORD your God may show us the way we should go, and the thing that we should do."
JER|42|4|Jeremiah the prophet said to them, "I have heard you. Behold, I will pray to the LORD your God according to your request, and whatever the LORD answers you I will tell you. I will keep nothing back from you."
JER|42|5|Then they said to Jeremiah, "May the LORD be a true and faithful witness against us if we do not act according to all the word with which the LORD your God sends you to us.
JER|42|6|Whether it is good or bad, we will obey the voice of the LORD our God to whom we are sending you, that it may be well with us when we obey the voice of the LORD our God."
JER|42|7|At the end of ten days the word of the LORD came to Jeremiah.
JER|42|8|Then he summoned Johanan the son of Kareah and all the commanders of the forces who were with him, and all the people from the least to the greatest,
JER|42|9|and said to them, "Thus says the LORD, the God of Israel, to whom you sent me to present your plea for mercy before him:
JER|42|10|If you will remain in this land, then I will build you up and not pull you down; I will plant you, and not pluck you up; for I relent of the disaster that I did to you.
JER|42|11|Do not fear the king of Babylon, of whom you are afraid. Do not fear him, declares the LORD, for I am with you, to save you and to deliver you from his hand.
JER|42|12|I will grant you mercy, that he may have mercy on you and let you remain in your own land.
JER|42|13|But if you say, 'We will not remain in this land,' disobeying the voice of the LORD your God
JER|42|14|and saying, 'No, we will go to the land of Egypt, where we shall not see war or hear the sound of the trumpet or be hungry for bread, and we will dwell there,'
JER|42|15|then hear the word of the LORD, O remnant of Judah. Thus says the LORD of hosts, the God of Israel: If you set your faces to enter Egypt and go to live there,
JER|42|16|then the sword that you fear shall overtake you there in the land of Egypt, and the famine of which you are afraid shall follow close after you to Egypt, and there you shall die.
JER|42|17|All the men who set their faces to go to Egypt to live there shall die by the sword, by famine, and by pestilence. They shall have no remnant or survivor from the disaster that I will bring upon them.
JER|42|18|"For thus says the LORD of hosts, the God of Israel: As my anger and my wrath were poured out on the inhabitants of Jerusalem, so my wrath will be poured out on you when you go to Egypt. You shall become an execration, a horror, a curse, and a taunt. You shall see this place no more.
JER|42|19|The LORD has said to you, O remnant of Judah, 'Do not go to Egypt.' Know for a certainty that I have warned you this day
JER|42|20|that you have gone astray at the cost of your lives. For you sent me to the LORD your God, saying, 'Pray for us to the LORD our God, and whatever the LORD our God says declare to us and we will do it.'
JER|42|21|And I have this day declared it to you, but you have not obeyed the voice of the LORD your God in anything that he sent me to tell you.
JER|42|22|Now therefore know for a certainty that you shall die by the sword, by famine, and by pestilence in the place where you desire to go to live."
JER|43|1|When Jeremiah finished speaking to all the people all these words of the LORD their God, with which the LORD their God had sent him to them,
JER|43|2|Azariah the son of Hoshaiah and Johanan the son of Kareah and all the insolent men said to Jeremiah, "You are telling a lie. The LORD our God did not send you to say, 'Do not go to Egypt to live there,'
JER|43|3|but Baruch the son of Neriah has set you against us, to deliver us into the hand of the Chaldeans, that they may kill us or take us into exile in Babylon."
JER|43|4|So Johanan the son of Kareah and all the commanders of the forces and all the people did not obey the voice of the LORD, to remain in the land of Judah.
JER|43|5|But Johanan the son of Kareah and all the commanders of the forces took all the remnant of Judah who had returned to live in the land of Judah from all the nations to which they had been driven-
JER|43|6|the men, the women, the children, the princesses, and every person whom Nebuzaradan the captain of the guard had left with Gedaliah the son of Ahikam, son of Shaphan; also Jeremiah the prophet and Baruch the son of Neriah.
JER|43|7|And they came into the land of Egypt, for they did not obey the voice of the LORD. And they arrived at Tahpanhes.
JER|43|8|Then the word of the LORD came to Jeremiah in Tahpanhes:
JER|43|9|"Take in your hands large stones and hide them in the mortar in the pavement that is at the entrance to Pharaoh's palace in Tahpanhes, in the sight of the men of Judah,
JER|43|10|and say to them, 'Thus says the LORD of hosts, the God of Israel: Behold, I will send and take Nebuchadnezzar the king of Babylon, my servant, and I will set his throne above these stones that I have hidden, and he will spread his royal canopy over them.
JER|43|11|He shall come and strike the land of Egypt, giving over to the pestilence those who are doomed to the pestilence, to captivity those who are doomed to captivity, and to the sword those who are doomed to the sword.
JER|43|12|I shall kindle a fire in the temples of the gods of Egypt, and he shall burn them and carry them away captive. And he shall clean the land of Egypt as a shepherd cleans his cloak of vermin, and he shall go away from there in peace.
JER|43|13|He shall break the obelisks of Heliopolis, which is in the land of Egypt, and the temples of the gods of Egypt he shall burn with fire.'"
JER|44|1|The word that came to Jeremiah concerning all the Judeans who lived in the land of Egypt, at Migdol, at Tahpanhes, at Memphis, and in the land of Pathros,
JER|44|2|"Thus says the LORD of hosts, the God of Israel: You have seen all the disaster that I brought upon Jerusalem and upon all the cities of Judah. Behold, this day they are a desolation, and no one dwells in them,
JER|44|3|because of the evil that they committed, provoking me to anger, in that they went to make offerings and serve other gods that they knew not, neither they, nor you, nor your fathers.
JER|44|4|Yet I persistently sent to you all my servants the prophets, saying, 'Oh, do not do this abomination that I hate!'
JER|44|5|But they did not listen or incline their ear, to turn from their evil and make no offerings to other gods.
JER|44|6|Therefore my wrath and my anger were poured out and kindled in the cities of Judah and in the streets of Jerusalem, and they became a waste and a desolation, as at this day.
JER|44|7|And now thus says the Lord GOD of hosts, the God of Israel: Why do you commit this great evil against yourselves, to cut off from you man and woman, infant and child, from the midst of Judah, leaving you no remnant?
JER|44|8|Why do you provoke me to anger with the works of your hands, making offerings to other gods in the land of Egypt where you have come to live, so that you may be cut off and become a curse and a taunt among all the nations of the earth?
JER|44|9|Have you forgotten the evil of your fathers, the evil of the kings of Judah, the evil of their wives, your own evil, and the evil of your wives, which they committed in the land of Judah and in the streets of Jerusalem?
JER|44|10|They have not humbled themselves even to this day, nor have they feared, nor walked in my law and my statutes that I set before you and before your fathers.
JER|44|11|"Therefore thus says the LORD of hosts, the God of Israel: Behold, I will set my face against you for harm, to cut off all Judah.
JER|44|12|I will take the remnant of Judah who have set their faces to come to the land of Egypt to live, and they shall all be consumed. In the land of Egypt they shall fall; by the sword and by famine they shall be consumed. From the least to the greatest, they shall die by the sword and by famine, and they shall become an oath, a horror, a curse, and a taunt.
JER|44|13|I will punish those who dwell in the land of Egypt, as I have punished Jerusalem, with the sword, with famine, and with pestilence,
JER|44|14|so that none of the remnant of Judah who have come to live in the land of Egypt shall escape or survive or return to the land of Judah, to which they desire to return to dwell there. For they shall not return, except some fugitives."
JER|44|15|Then all the men who knew that their wives had made offerings to other gods, and all the women who stood by, a great assembly, all the people who lived in Pathros in the land of Egypt, answered Jeremiah:
JER|44|16|"As for the word that you have spoken to us in the name of the LORD, we will not listen to you.
JER|44|17|But we will do everything that we have vowed, make offerings to the queen of heaven and pour out drink offerings to her, as we did, both we and our fathers, our kings and our officials, in the cities of Judah and in the streets of Jerusalem. For then we had plenty of food, and prospered, and saw no disaster.
JER|44|18|But since we left off making offerings to the queen of heaven and pouring out drink offerings to her, we have lacked everything and have been consumed by the sword and by famine."
JER|44|19|And the women said, "When we made offerings to the queen of heaven and poured out drink offerings to her, was it without our husbands' approval that we made cakes for her bearing her image and poured out drink offerings to her?"
JER|44|20|Then Jeremiah said to all the people, men and women, all the people who had given him this answer:
JER|44|21|"As for the offerings that you offered in the cities of Judah and in the streets of Jerusalem, you and your fathers, your kings and your officials, and the people of the land, did not the LORD remember them? Did it not come into his mind?
JER|44|22|The LORD could no longer bear your evil deeds and the abominations that you committed. Therefore your land has become a desolation and a waste and a curse, without inhabitant, as it is this day.
JER|44|23|It is because you made offerings and because you sinned against the LORD and did not obey the voice of the LORD or walk in his law and in his statutes and in his testimonies that this disaster has happened to you, as at this day."
JER|44|24|Jeremiah said to all the people and all the women, "Hear the word of the LORD, all you of Judah who are in the land of Egypt.
JER|44|25|Thus says the LORD of hosts, the God of Israel: You and your wives have declared with your mouths, and have fulfilled it with your hands, saying, 'We will surely perform our vows that we have made, to make offerings to the queen of heaven and to pour out drink offerings to her.' Then confirm your vows and perform your vows!
JER|44|26|Therefore hear the word of the LORD, all you of Judah who dwell in the land of Egypt: Behold, I have sworn by my great name, says the LORD, that my name shall no more be invoked by the mouth of any man of Judah in all the land of Egypt, saying, 'As the Lord GOD lives.'
JER|44|27|Behold, I am watching over them for disaster and not for good. All the men of Judah who are in the land of Egypt shall be consumed by the sword and by famine, until there is an end of them.
JER|44|28|And those who escape the sword shall return from the land of Egypt to the land of Judah, few in number; and all the remnant of Judah, who came to the land of Egypt to live, shall know whose word will stand, mine or theirs.
JER|44|29|This shall be the sign to you, declares the LORD, that I will punish you in this place, in order that you may know that my words will surely stand against you for harm:
JER|44|30|Thus says the LORD, behold, I will give Pharaoh Hophra king of Egypt into the hand of his enemies and into the hand of those who seek his life, as I gave Zedekiah king of Judah into the hand of Nebuchadnezzar king of Babylon, who was his enemy and sought his life."
JER|45|1|The word that Jeremiah the prophet spoke to Baruch the son of Neriah, when he wrote these words in a book at the dictation of Jeremiah, in the fourth year of Jehoiakim the son of Josiah, king of Judah:
JER|45|2|"Thus says the LORD, the God of Israel, to you, O Baruch:
JER|45|3|You said, 'Woe is me! For the LORD has added sorrow to my pain. I am weary with my groaning, and I find no rest.'
JER|45|4|Thus shall you say to him, Thus says the LORD: Behold, what I have built I am breaking down, and what I have planted I am plucking up- that is, the whole land.
JER|45|5|And do you seek great things for yourself? Seek them not, for behold, I am bringing disaster upon all flesh, declares the LORD. But I will give you your life as a prize of war in all places to which you may go."
JER|46|1|The word of the LORD that came to Jeremiah the prophet concerning the nations.
JER|46|2|About Egypt. Concerning the army of Pharaoh Neco, king of Egypt, which was by the river Euphrates at Carchemish and which Nebuchadnezzar king of Babylon defeated in the fourth year of Jehoiakim the son of Josiah, king of Judah:
JER|46|3|"Prepare buckler and shield, and advance for battle!
JER|46|4|Harness the horses; mount, O horsemen! Take your stations with your helmets, polish your spears, put on your armor!
JER|46|5|Why have I seen it? They are dismayed and have turned backward. Their warriors are beaten down and have fled in haste; they look not back- terror on every side! declares the LORD.
JER|46|6|The swift cannot flee away, nor the warrior escape; in the north by the river Euphrates they have stumbled and fallen.
JER|46|7|"Who is this, rising like the Nile, like rivers whose waters surge?
JER|46|8|Egypt rises like the Nile, like rivers whose waters surge. He said, 'I will rise, I will cover the earth, I will destroy cities and their inhabitants.'
JER|46|9|Advance, O horses, and rage, O chariots! Let the warriors go out: men of Cush and Put who handle the shield, men of Lud, skilled in handling the bow.
JER|46|10|That day is the day of the Lord GOD of hosts, a day of vengeance, to avenge himself on his foes. The sword shall devour and be sated and drink its fill of their blood. For the Lord GOD of hosts holds a sacrifice in the north country by the river Euphrates.
JER|46|11|Go up to Gilead, and take balm, O virgin daughter of Egypt! In vain you have used many medicines; there is no healing for you.
JER|46|12|The nations have heard of your shame, and the earth is full of your cry; for warrior has stumbled against warrior; they have both fallen together."
JER|46|13|The word that the LORD spoke to Jeremiah the prophet about the coming of Nebuchadnezzar king of Babylon to strike the land of Egypt:
JER|46|14|"Declare in Egypt, and proclaim in Migdol; proclaim in Memphis and Tahpanhes; Say, 'Stand ready and be prepared, for the sword shall devour around you.'
JER|46|15|Why are your mighty ones face down? They do not stand because the LORD thrust them down.
JER|46|16|He made many stumble, and they fell, and they said one to another, 'Arise, and let us go back to our own people and to the land of our birth, because of the sword of the oppressor.'
JER|46|17|Call the name of Pharaoh, king of Egypt, 'Noisy one who lets the hour go by.'
JER|46|18|"As I live, declares the King, whose name is the LORD of hosts, like Tabor among the mountains and like Carmel by the sea, shall one come.
JER|46|19|Prepare yourselves baggage for exile, O inhabitants of Egypt! For Memphis shall become a waste, a ruin, without inhabitant.
JER|46|20|"A beautiful heifer is Egypt, but a biting fly from the north has come upon her.
JER|46|21|Even her hired soldiers in her midst are like fattened calves; yes, they have turned and fled together; they did not stand, for the day of their calamity has come upon them, the time of their punishment.
JER|46|22|"She makes a sound like a serpent gliding away; for her enemies march in force and come against her with axes like those who fell trees.
JER|46|23|They shall cut down her forest, declares the LORD, though it is impenetrable, because they are more numerous than locusts; they are without number.
JER|46|24|The daughter of Egypt shall be put to shame; she shall be delivered into the hand of a people from the north."
JER|46|25|The LORD of hosts, the God of Israel, said: "Behold, I am bringing punishment upon Amon of Thebes, and Pharaoh and Egypt and her gods and her kings, upon Pharaoh and those who trust in him.
JER|46|26|I will deliver them into the hand of those who seek their life, into the hand of Nebuchadnezzar king of Babylon and his officers. Afterward Egypt shall be inhabited as in the days of old, declares the LORD.
JER|46|27|"But fear not, O Jacob my servant, nor be dismayed, O Israel, for behold, I will save you from far away, and your offspring from the land of their captivity. Jacob shall return and have quiet and ease, and none shall make him afraid.
JER|46|28|Fear not, O Jacob my servant, declares the LORD, for I am with you. I will make a full end of all the nations to which I have driven you, but of you I will not make a full end. I will discipline you in just measure, and I will by no means leave you unpunished."
JER|47|1|The word of the LORD that came to Jeremiah the prophet concerning the Philistines, before Pharaoh struck down Gaza.
JER|47|2|"Thus says the LORD: Behold, waters are rising out of the north, and shall become an overflowing torrent; they shall overflow the land and all that fills it, the city and those who dwell in it. Men shall cry out, and every inhabitant of the land shall wail.
JER|47|3|At the noise of the stamping of the hoofs of his stallions, at the rushing of his chariots, at the rumbling of their wheels, the fathers look not back to their children, so feeble are their hands,
JER|47|4|because of the day that is coming to destroy all the Philistines, to cut off from Tyre and Sidon every helper that remains. For the LORD is destroying the Philistines, the remnant of the coastland of Caphtor.
JER|47|5|Baldness has come upon Gaza; Ashkelon has perished. O remnant of their valley, how long will you gash yourselves?
JER|47|6|Ah, sword of the LORD! How long till you are quiet? Put yourself into your scabbard; rest and be still!
JER|47|7|How can it be quiet when the LORD has given it a charge? Against Ashkelon and against the seashore he has appointed it."
JER|48|1|Concerning Moab.Thus says the LORD of hosts, the God of Israel: "Woe to Nebo, for it is laid waste! Kiriathaim is put to shame, it is taken; the fortress is put to shame and broken down;
JER|48|2|the renown of Moab is no more. In Heshbon they planned disaster against her: 'Come, let us cut her off from being a nation!' You also, O Madmen, shall be brought to silence; the sword shall pursue you.
JER|48|3|"Hark! A cry from Horonaim, 'Desolation and great destruction!'
JER|48|4|Moab is destroyed; her little ones have made a cry.
JER|48|5|For at the ascent of Luhith they go up weeping; for at the descent of Horonaim they have heard the distressed cry of destruction.
JER|48|6|Flee! Save yourselves! You will be like a juniper in the desert!
JER|48|7|For, because you trusted in your works and your treasures, you also shall be taken; and Chemosh shall go into exile with his priests and his officials.
JER|48|8|The destroyer shall come upon every city, and no city shall escape; the valley shall perish, and the plain shall be destroyed, as the LORD has spoken.
JER|48|9|"Give wings to Moab, for she would fly away; her cities shall become a desolation, with no inhabitant in them.
JER|48|10|"Cursed is he who does the work of the LORD with slackness, and cursed is he who keeps back his sword from bloodshed.
JER|48|11|"Moab has been at ease from his youth and has settled on his dregs; he has not been emptied from vessel to vessel, nor has he gone into exile; so his taste remains in him, and his scent is not changed.
JER|48|12|"Therefore, behold, the days are coming, declares the LORD, when I shall send to him pourers who will pour him, and empty his vessels and break his jars in pieces.
JER|48|13|Then Moab shall be ashamed of Chemosh, as the house of Israel was ashamed of Bethel, their confidence.
JER|48|14|"How do you say, 'We are heroes and mighty men of war'?
JER|48|15|The destroyer of Moab and his cities has come up, and the choicest of his young men have gone down to slaughter, declares the King, whose name is the LORD of hosts.
JER|48|16|The calamity of Moab is near at hand, and his affliction hastens swiftly.
JER|48|17|Grieve for him, all you who are around him, and all who know his name; say, 'How the mighty scepter is broken, the glorious staff.'
JER|48|18|"Come down from your glory, and sit on the parched ground, O inhabitant of Dibon! For the destroyer of Moab has come up against you; he has destroyed your strongholds.
JER|48|19|Stand by the way and watch, O inhabitant of Aroer! Ask him who flees and her who escapes; say, 'What has happened?'
JER|48|20|Moab is put to shame, for it is broken; wail and cry! Tell it beside the Arnon, that Moab is laid waste.
JER|48|21|"Judgment has come upon the tableland, upon Holon, and Jahzah, and Mephaath,
JER|48|22|and Dibon, and Nebo, and Beth-diblathaim,
JER|48|23|and Kiriathaim, and Beth-gamul, and Beth-meon,
JER|48|24|and Kerioth, and Bozrah, and all the cities of the land of Moab, far and near.
JER|48|25|The horn of Moab is cut off, and his arm is broken, declares the LORD.
JER|48|26|"Make him drunk, because he magnified himself against the LORD, so that Moab shall wallow in his vomit, and he too shall be held in derision.
JER|48|27|Was not Israel a derision to you? Was he found among thieves, that whenever you spoke of him you wagged your head?
JER|48|28|"Leave the cities, and dwell in the rock, O inhabitants of Moab! Be like the dove that nests in the sides of the mouth of a gorge.
JER|48|29|We have heard of the pride of Moab- he is very proud- of his loftiness, his pride, and his arrogance, and the haughtiness of his heart.
JER|48|30|I know his insolence, declares the LORD; his boasts are false, his deeds are false.
JER|48|31|Therefore I wail for Moab; I cry out for all Moab; for the men of Kir-hareseth I mourn.
JER|48|32|More than for Jazer I weep for you, O vine of Sibmah! Your branches passed over the sea, reached to the Sea of Jazer; on your summer fruits and your grapes the destroyer has fallen.
JER|48|33|Gladness and joy have been taken away from the fruitful land of Moab; I have made the wine cease from the wine presses; no one treads them with shouts of joy; the shouting is not the shout of joy.
JER|48|34|"From the outcry at Heshbon even to Elealeh, as far as Jahaz they utter their voice, from Zoar to Horonaim and Eglath-shelishiyah. For the waters of Nimrim also have become desolate.
JER|48|35|And I will bring to an end in Moab, declares the LORD, him who offers sacrifice in the high place and makes offerings to his god.
JER|48|36|Therefore my heart moans for Moab like a flute, and my heart moans like a flute for the men of Kir-hareseth. Therefore the riches they gained have perished.
JER|48|37|"For every head is shaved and every beard cut off. On all the hands are gashes, and around the waist is sackcloth.
JER|48|38|On all the housetops of Moab and in the squares there is nothing but lamentation, for I have broken Moab like a vessel for which no one cares, declares the LORD.
JER|48|39|How it is broken! How they wail! How Moab has turned his back in shame! So Moab has become a derision and a horror to all that are around him."
JER|48|40|For thus says the LORD: "Behold, one shall fly swiftly like an eagle and spread his wings against Moab;
JER|48|41|the cities shall be taken and the strongholds seized. The heart of the warriors of Moab shall be in that day like the heart of a woman in her birth pains;
JER|48|42|Moab shall be destroyed and be no longer a people, because he magnified himself against the LORD.
JER|48|43|Terror, pit, and snare are before you, O inhabitant of Moab! declares the LORD.
JER|48|44|He who flees from the terror shall fall into the pit, and he who climbs out of the pit shall be caught in the snare. For I will bring these things upon Moab, the year of their punishment, declares the LORD.
JER|48|45|"In the shadow of Heshbon fugitives stop without strength, for fire came out from Heshbon, flame from the house of Sihon; it has destroyed the forehead of Moab, the crown of the sons of tumult.
JER|48|46|Woe to you, O Moab! The people of Chemosh are undone, for your sons have been taken captive, and your daughters into captivity.
JER|48|47|Yet I will restore the fortunes of Moab in the latter days, declares the LORD." Thus far is the judgment on Moab.
JER|49|1|Concerning the Ammonites.Thus says the LORD: "Has Israel no sons? Has he no heir? Why then has Milcom dispossessed Gad, and his people settled in its cities?
JER|49|2|Therefore, behold, the days are coming, declares the LORD, when I will cause the battle cry to be heard against Rabbah of the Ammonites; it shall become a desolate mound, and its villages shall be burned with fire; then Israel shall dispossess those who dispossessed him, says the LORD.
JER|49|3|"Wail, O Heshbon, for Ai is laid waste! Cry out, O daughters of Rabbah! put on sackcloth, lament, and run to and fro among the hedges! For Milcom shall go into exile, with his priests and his officials.
JER|49|4|Why do you boast of your valleys, O faithless daughter, who trusted in her treasures, saying, 'Who will come against me?'
JER|49|5|Behold, I will bring terror upon you, declares the Lord GOD of hosts, from all who are around you, and you shall be driven out, every man straight before him, with none to gather the fugitives.
JER|49|6|"But afterward I will restore the fortunes of the Ammonites, declares the LORD."
JER|49|7|Concerning Edom. Thus says the LORD of hosts: "Is wisdom no more in Teman? Has counsel perished from the prudent? Has their wisdom vanished?
JER|49|8|Flee, turn back, dwell in the depths, O inhabitants of Dedan! For I will bring the calamity of Esau upon him, the time when I punish him.
JER|49|9|If grape-gatherers came to you, would they not leave gleanings? If thieves came by night, would they not destroy only enough for themselves?
JER|49|10|But I have stripped Esau bare; I have uncovered his hiding places, and he is not able to conceal himself. His children are destroyed, and his brothers, and his neighbors; and he is no more.
JER|49|11|Leave your fatherless children; I will keep them alive; and let your widows trust in me."
JER|49|12|For thus says the LORD: "If those who did not deserve to drink the cup must drink it, will you go unpunished? You shall not go unpunished, but you must drink.
JER|49|13|For I have sworn by myself, declares the LORD, that Bozrah shall become a horror, a taunt, a waste, and a curse, and all her cities shall be perpetual wastes."
JER|49|14|I have heard a message from the LORD, and an envoy has been sent among the nations: "Gather yourselves together and come against her, and rise up for battle!
JER|49|15|For behold, I will make you small among the nations, despised among mankind.
JER|49|16|The horror you inspire has deceived you, and the pride of your heart, you who live in the clefts of the rock, who hold the height of the hill. Though you make your nest as high as the eagle's, I will bring you down from there, declares the LORD.
JER|49|17|"Edom shall become a horror. Everyone who passes by it will be horrified and will hiss because of all its disasters.
JER|49|18|As when Sodom and Gomorrah and their neighboring cities were overthrown, says the LORD, no man shall dwell there, no man shall sojourn in her.
JER|49|19|Behold, like a lion coming up from the jungle of the Jordan against a perennial pasture, I will suddenly make him run away from her. And I will appoint over her whomever I choose. For who is like me? Who will summon me? What shepherd can stand before me?
JER|49|20|Therefore hear the plan that the LORD has made against Edom and the purposes that he has formed against the inhabitants of Teman: Even the little ones of the flock shall be dragged away. Surely their fold shall be appalled at their fate.
JER|49|21|At the sound of their fall the earth shall tremble; the sound of their cry shall be heard at the Red Sea.
JER|49|22|Behold, one shall mount up and fly swiftly like an eagle and spread his wings against Bozrah, and the heart of the warriors of Edom shall be in that day like the heart of a woman in her birth pains."
JER|49|23|Concerning Damascus: "Hamath and Arpad are confounded, for they have heard bad news; they melt in fear, they are troubled like the sea that cannot be quiet.
JER|49|24|Damascus has become feeble, she turned to flee, and panic seized her; anguish and sorrows have taken hold of her, as of a woman in labor.
JER|49|25|How is the famous city not forsaken, the city of my joy?
JER|49|26|Therefore her young men shall fall in her squares, and all her soldiers shall be destroyed in that day, declares the LORD of hosts.
JER|49|27|And I will kindle a fire in the wall of Damascus, and it shall devour the strongholds of Ben-hadad."
JER|49|28|Concerning Kedar and the kingdoms of Hazor that Nebuchadnezzar king of Babylon struck down. Thus says the LORD: "Rise up, advance against Kedar! Destroy the people of the east!
JER|49|29|Their tents and their flocks shall be taken, their curtains and all their goods; their camels shall be led away from them, and men shall cry to them: 'Terror on every side!'
JER|49|30|Flee, wander far away, dwell in the depths, O inhabitants of Hazor! declares the LORD. For Nebuchadnezzar king of Babylon has made a plan against you and formed a purpose against you.
JER|49|31|"Rise up, advance against a nation at ease, that dwells securely, declares the LORD, that has no gates or bars, that dwells alone.
JER|49|32|Their camels shall become plunder, their herds of livestock a spoil. I will scatter to every wind those who cut the corners of their hair, and I will bring their calamity from every side of them, declares the LORD.
JER|49|33|Hazor shall become a haunt of jackals, an everlasting waste; no man shall dwell there; no man shall sojourn in her."
JER|49|34|The word of the LORD that came to Jeremiah the prophet concerning Elam, in the beginning of the reign of Zedekiah king of Judah.
JER|49|35|Thus says the LORD of hosts: "Behold, I will break the bow of Elam, the mainstay of their might.
JER|49|36|And I will bring upon Elam the four winds from the four quarters of heaven. And I will scatter them to all those winds, and there shall be no nation to which those driven out of Elam shall not come.
JER|49|37|I will terrify Elam before their enemies and before those who seek their life. I will bring disaster upon them, my fierce anger, declares the LORD. I will send the sword after them, until I have consumed them,
JER|49|38|and I will set my throne in Elam and destroy their king and officials, declares the LORD.
JER|49|39|"But in the latter days I will restore the fortunes of Elam, declares the LORD."
JER|50|1|The word that the LORD spoke concerning Babylon, concerning the land of the Chaldeans, by Jeremiah the prophet:
JER|50|2|"Declare among the nations and proclaim, set up a banner and proclaim, conceal it not, and say: 'Babylon is taken, Bel is put to shame, Merodach is dismayed. Her images are put to shame, her idols are dismayed.'
JER|50|3|"For out of the north a nation has come up against her, which shall make her land a desolation, and none shall dwell in it; both man and beast shall flee away.
JER|50|4|"In those days and in that time, declares the LORD, the people of Israel and the people of Judah shall come together, weeping as they come, and they shall seek the LORD their God.
JER|50|5|They shall ask the way to Zion, with faces turned toward it, saying, 'Come, let us join ourselves to the LORD in an everlasting covenant that will never be forgotten.'
JER|50|6|"My people have been lost sheep. Their shepherds have led them astray, turning them away on the mountains. From mountain to hill they have gone. They have forgotten their fold.
JER|50|7|All who found them have devoured them, and their enemies have said, 'We are not guilty, for they have sinned against the LORD, their habitation of righteousness, the LORD, the hope of their fathers.'
JER|50|8|"Flee from the midst of Babylon, and go out of the land of the Chaldeans, and be as male goats before the flock.
JER|50|9|For behold, I am stirring up and bringing against Babylon a gathering of great nations, from the north country. And they shall array themselves against her. From there she shall be taken. Their arrows are like a skilled warrior who does not return empty-handed.
JER|50|10|Chaldea shall be plundered; all who plunder her shall be sated, declares the LORD.
JER|50|11|"Though you rejoice, though you exult, O plunderers of my heritage, though you frolic like a heifer in the pasture, and neigh like stallions,
JER|50|12|your mother shall be utterly shamed, and she who bore you shall be disgraced. Behold, she shall be the last of the nations, a wilderness, a dry land, and a desert.
JER|50|13|Because of the wrath of the LORD she shall not be inhabited but shall be an utter desolation; everyone who passes by Babylon shall be appalled, and hiss because of all her wounds.
JER|50|14|Set yourselves in array against Babylon all around, all you who bend the bow; shoot at her, spare no arrows, for she has sinned against the LORD.
JER|50|15|Raise a shout against her all around; she has surrendered; her bulwarks have fallen; her walls are thrown down. For this is the vengeance of the LORD: take vengeance on her; do to her as she has done.
JER|50|16|Cut off from Babylon the sower, and the one who handles the sickle in time of harvest; because of the sword of the oppressor, every one shall turn to his own people, and every one shall flee to his own land.
JER|50|17|"Israel is a hunted sheep driven away by lions. First the king of Assyria devoured him, and now at last Nebuchadnezzar king of Babylon has gnawed his bones.
JER|50|18|Therefore, thus says the LORD of hosts, the God of Israel: Behold, I am bringing punishment on the king of Babylon and his land, as I punished the king of Assyria.
JER|50|19|I will restore Israel to his pasture, and he shall feed on Carmel and in Bashan, and his desire shall be satisfied on the hills of Ephraim and in Gilead.
JER|50|20|In those days and in that time, declares the LORD, iniquity shall be sought in Israel, and there shall be none. And sin in Judah, and none shall be found, for I will pardon those whom I leave as a remnant.
JER|50|21|"Go up against the land of Merathaim, and against the inhabitants of Pekod. Kill, and devote them to destruction, declares the LORD, and do all that I have commanded you.
JER|50|22|The noise of battle is in the land, and great destruction!
JER|50|23|How the hammer of the whole earth is cut down and broken! How Babylon has become a horror among the nations!
JER|50|24|I set a snare for you and you were taken, O Babylon, and you did not know it; you were found and caught, because you opposed the LORD.
JER|50|25|The LORD has opened his armory and brought out the weapons of his wrath, for the Lord GOD of hosts has a work to do in the land of the Chaldeans.
JER|50|26|Come against her from every quarter; open her granaries; pile her up like heaps of grain, and devote her to destruction; let nothing be left of her.
JER|50|27|Kill all her bulls; let them go down to the slaughter. Woe to them, for their day has come, the time of their punishment.
JER|50|28|"A voice! They flee and escape from the land of Babylon, to declare in Zion the vengeance of the LORD our God, vengeance for his temple.
JER|50|29|"Summon archers against Babylon, all those who bend the bow. Encamp around her; let no one escape. Repay her according to her deeds; do to her according to all that she has done. For she has proudly defied the LORD, the Holy One of Israel.
JER|50|30|Therefore her young men shall fall in her squares, and all her soldiers shall be destroyed on that day, declares the LORD.
JER|50|31|"Behold, I am against you, O proud one, declares the Lord GOD of hosts, for your day has come, the time when I will punish you.
JER|50|32|The proud one shall stumble and fall, with none to raise him up, and I will kindle a fire in his cities, and it will devour all that is around him.
JER|50|33|"Thus says the LORD of hosts: The people of Israel are oppressed, and the people of Judah with them. All who took them captive have held them fast; they refuse to let them go.
JER|50|34|Their Redeemer is strong; the LORD of hosts is his name. He will surely plead their cause, that he may give rest to the earth, but unrest to the inhabitants of Babylon.
JER|50|35|"A sword against the Chaldeans, declares the LORD, and against the inhabitants of Babylon, and against her officials and her wise men!
JER|50|36|A sword against the diviners, that they may become fools! A sword against her warriors, that they may be destroyed!
JER|50|37|A sword against her horses and against her chariots, and against all the foreign troops in her midst, that they may become women! A sword against all her treasures, that they may be plundered!
JER|50|38|A drought against her waters, that they may be dried up! For it is a land of images, and they are mad over idols.
JER|50|39|"Therefore wild beasts shall dwell with hyenas in Babylon, and ostriches shall dwell in her. She shall never again have people, nor be inhabited for all generations.
JER|50|40|As when God overthrew Sodom and Gomorrah and their neighboring cities, declares the LORD, so no man shall dwell there, and no son of man shall sojourn in her.
JER|50|41|"Behold, a people comes from the north; a mighty nation and many kings are stirring from the farthest parts of the earth.
JER|50|42|They lay hold of bow and spear; they are cruel and have no mercy. The sound of them is like the roaring of the sea; they ride on horses, arrayed as a man for battle against you, O daughter of Babylon!
JER|50|43|"The king of Babylon heard the report of them, and his hands fell helpless; anguish seized him, pain as of a woman in labor.
JER|50|44|"Behold, like a lion coming up from the thicket of the Jordan against a perennial pasture, I will suddenly make them run away from her, and I will appoint over her whomever I choose. For who is like me? Who will summon me? What shepherd can stand before me?
JER|50|45|Therefore hear the plan that the LORD has made against Babylon, and the purposes that he has formed against the land of the Chaldeans: Surely the little ones of their flock shall be dragged away; surely their fold shall be appalled at their fate.
JER|50|46|At the sound of the capture of Babylon the earth shall tremble, and her cry shall be heard among the nations."
JER|51|1|Thus says the LORD: "Behold, I will stir up the spirit of a destroyer against Babylon, against the inhabitants of Leb-kamai,
JER|51|2|and I will send to Babylon winnowers, and they shall winnow her, and they shall empty her land, when they come against her from every side on the day of trouble.
JER|51|3|Let not the archer bend his bow, and let him not stand up in his armor. Spare not her young men; devote to destruction all her army.
JER|51|4|They shall fall down slain in the land of the Chaldeans, and wounded in her streets.
JER|51|5|For Israel and Judah have not been forsaken by their God, the LORD of hosts, but the land of the Chaldeans is full of guilt against the Holy One of Israel.
JER|51|6|"Flee from the midst of Babylon; let every one save his life! Be not cut off in her punishment, for this is the time of the LORD's vengeance, the repayment he is rendering her.
JER|51|7|Babylon was a golden cup in the LORD's hand, making all the earth drunken; the nations drank of her wine; therefore the nations went mad.
JER|51|8|Suddenly Babylon has fallen and been broken; wail for her! Take balm for her pain; perhaps she may be healed.
JER|51|9|We would have healed Babylon, but she was not healed. Forsake her, and let us go each to his own country, for her judgment has reached up to heaven and has been lifted up even to the skies.
JER|51|10|The LORD has brought about our vindication; come, let us declare in Zion the work of the LORD our God.
JER|51|11|"Sharpen the arrows! Take up the shields! The LORD has stirred up the spirit of the kings of the Medes, because his purpose concerning Babylon is to destroy it, for that is the vengeance of the LORD, the vengeance for his temple.
JER|51|12|"Set up a standard against the walls of Babylon; make the watch strong; set up watchmen; prepare the ambushes; for the LORD has both planned and done what he spoke concerning the inhabitants of Babylon.
JER|51|13|O you who dwell by many waters, rich in treasures, your end has come; the thread of your life is cut.
JER|51|14|The LORD of hosts has sworn by himself: Surely I will fill you with men, as many as locusts, and they shall raise the shout of victory over you.
JER|51|15|"It is he who made the earth by his power, who established the world by his wisdom, and by his understanding stretched out the heavens.
JER|51|16|When he utters his voice there is a tumult of waters in the heavens, and he makes the mist rise from the ends of the earth. He makes lightning for the rain, and he brings forth the wind from his storehouses.
JER|51|17|Every man is stupid and without knowledge; every goldsmith is put to shame by his idols, for his images are false, and there is no breath in them.
JER|51|18|They are worthless, a work of delusion; at the time of their punishment they shall perish.
JER|51|19|Not like these is he who is the portion of Jacob, for he is the one who formed all things, and Israel is the tribe of his inheritance; the LORD of hosts is his name.
JER|51|20|"You are my hammer and weapon of war: with you I break nations in pieces; with you I destroy kingdoms;
JER|51|21|with you I break in pieces the horse and his rider; with you I break in pieces the chariot and the charioteer;
JER|51|22|with you I break in pieces man and woman; with you I break in pieces the old man and the youth; with you I break in pieces the young man and the young woman;
JER|51|23|with you I break in pieces the shepherd and his flock; with you I break in pieces the farmer and his team; with you I break in pieces governors and commanders.
JER|51|24|"I will repay Babylon and all the inhabitants of Chaldea before your very eyes for all the evil that they have done in Zion, declares the LORD.
JER|51|25|"Behold, I am against you, O destroying mountain, declares the LORD, which destroys the whole earth; I will stretch out my hand against you, and roll you down from the crags, and make you a burnt mountain.
JER|51|26|No stone shall be taken from you for a corner and no stone for a foundation, but you shall be a perpetual waste, declares the LORD.
JER|51|27|"Set up a standard on the earth; blow the trumpet among the nations; prepare the nations for war against her; summon against her the kingdoms, Ararat, Minni, and Ashkenaz; appoint a marshal against her; bring up horses like bristling locusts.
JER|51|28|Prepare the nations for war against her, the kings of the Medes, with their governors and deputies, and every land under their dominion.
JER|51|29|The land trembles and writhes in pain, for the LORD's purposes against Babylon stand, to make the land of Babylon a desolation, without inhabitant.
JER|51|30|The warriors of Babylon have ceased fighting; they remain in their strongholds; their strength has failed; they have become women; her dwellings are on fire; her bars are broken.
JER|51|31|One runner runs to meet another, and one messenger to meet another, to tell the king of Babylon that his city is taken on every side;
JER|51|32|the fords have been seized, the marshes are burned with fire, and the soldiers are in panic.
JER|51|33|For thus says the LORD of hosts, the God of Israel: The daughter of Babylon is like a threshing floor at the time when it is trodden; yet a little while and the time of her harvest will come."
JER|51|34|"Nebuchadnezzar the king of Babylon has devoured me; he has crushed me; he has made me an empty vessel; he has swallowed me like a monster; he has filled his stomach with my delicacies; he has rinsed me out.
JER|51|35|The violence done to me and to my kinsmen be upon Babylon," let the inhabitant of Zion say. "My blood be upon the inhabitants of Chaldea," let Jerusalem say.
JER|51|36|Therefore thus says the LORD: "Behold, I will plead your cause and take vengeance for you. I will dry up her sea and make her fountain dry,
JER|51|37|and Babylon shall become a heap of ruins, the haunt of jackals, a horror and a hissing, without inhabitant.
JER|51|38|"They shall roar together like lions; they shall growl like lions' cubs.
JER|51|39|While they are inflamed I will prepare them a feast and make them drunk, that they may become merry, then sleep a perpetual sleep and not wake, declares the LORD.
JER|51|40|I will bring them down like lambs to the slaughter, like rams and male goats.
JER|51|41|"How Babylon is taken, the praise of the whole earth seized! How Babylon has become a horror among the nations!
JER|51|42|The sea has come up on Babylon; she is covered with its tumultuous waves.
JER|51|43|Her cities have become a horror, a land of drought and a desert, a land in which no one dwells, and through which no son of man passes.
JER|51|44|And I will punish Bel in Babylon, and take out of his mouth what he has swallowed. The nations shall no longer flow to him; the wall of Babylon has fallen.
JER|51|45|"Go out of the midst of her, my people! Let every one save his life from the fierce anger of the LORD!
JER|51|46|Let not your heart faint, and be not fearful at the report heard in the land, when a report comes in one year and afterward a report in another year, and violence is in the land, and ruler is against ruler.
JER|51|47|"Therefore, behold, the days are coming when I will punish the images of Babylon; her whole land shall be put to shame, and all her slain shall fall in the midst of her.
JER|51|48|Then the heavens and the earth, and all that is in them, shall sing for joy over Babylon, for the destroyers shall come against them out of the north, declares the LORD.
JER|51|49|Babylon must fall for the slain of Israel, just as for Babylon have fallen the slain of all the earth.
JER|51|50|"You who have escaped from the sword, go, do not stand still! Remember the LORD from far away, and let Jerusalem come into your mind:
JER|51|51|'We are put to shame, for we have heard reproach; dishonor has covered our face, for foreigners have come into the holy places of the LORD's house.'
JER|51|52|"Therefore, behold, the days are coming, declares the LORD, when I will execute judgment upon her images, and through all her land the wounded shall groan.
JER|51|53|Though Babylon should mount up to heaven, and though she should fortify her strong height, yet destroyers would come from me against her, declares the LORD.
JER|51|54|"A voice! A cry from Babylon! The noise of great destruction from the land of the Chaldeans!
JER|51|55|For the LORD is laying Babylon waste and stilling her mighty voice. Their waves roar like many waters; the noise of their voice is raised,
JER|51|56|for a destroyer has come upon her, upon Babylon; her warriors are taken; their bows are broken in pieces, for the LORD is a God of recompense; he will surely repay.
JER|51|57|I will make drunk her officials and her wise men, her governors, her commanders, and her warriors; they shall sleep a perpetual sleep and not wake, declares the King, whose name is the LORD of hosts.
JER|51|58|"Thus says the LORD of hosts: The broad wall of Babylon shall be leveled to the ground, and her high gates shall be burned with fire. The peoples labor for nothing, and the nations weary themselves only for fire."
JER|51|59|The word that Jeremiah the prophet commanded Seraiah the son of Neriah, son of Mahseiah, when he went with Zedekiah king of Judah to Babylon, in the fourth year of his reign. Seraiah was the quartermaster.
JER|51|60|Jeremiah wrote in a book all the disaster that should come upon Babylon, all these words that are written concerning Babylon.
JER|51|61|And Jeremiah said to Seraiah: "When you come to Babylon, see that you read all these words,
JER|51|62|and say, 'O LORD, you have said concerning this place that you will cut it off, so that nothing shall dwell in it, neither man nor beast, and it shall be desolate forever.'
JER|51|63|When you finish reading this book, tie a stone to it and cast it into the midst of the Euphrates,
JER|51|64|and say, 'Thus shall Babylon sink, to rise no more, because of the disaster that I am bringing upon her, and they shall become exhausted.'"Thus far are the words of Jeremiah.
JER|52|1|Zedekiah was twenty-one years old when he became king; and he reigned eleven years in Jerusalem. His mother's name was Hamutal the daughter of Jeremiah of Libnah.
JER|52|2|And he did what was evil in the sight of the LORD, according to all that Jehoiakim had done.
JER|52|3|For because of the anger of the LORD things came to the point in Jerusalem and Judah that he cast them out from his presence. And Zedekiah rebelled against the king of Babylon.
JER|52|4|And in the ninth year of his reign, in the tenth month, on the tenth day of the month, Nebuchadnezzar king of Babylon came with all his army against Jerusalem, and laid siege to it. And they built siegeworks all around it.
JER|52|5|So the city was besieged till the eleventh year of King Zedekiah.
JER|52|6|On the ninth day of the fourth month the famine was so severe in the city that there was no food for the people of the land.
JER|52|7|Then a breach was made in the city, and all the men of war fled and went out from the city by night by the way of a gate between the two walls, by the king's garden, while the Chaldeans were around the city. And they went in the direction of the Arabah.
JER|52|8|But the army of the Chaldeans pursued the king and overtook Zedekiah in the plains of Jericho. And all his army was scattered from him.
JER|52|9|Then they captured the king and brought him up to the king of Babylon at Riblah in the land of Hamath, and he passed sentence on him.
JER|52|10|The king of Babylon slaughtered the sons of Zedekiah before his eyes, and also slaughtered all the officials of Judah at Riblah.
JER|52|11|He put out the eyes of Zedekiah, and bound him in chains, and the king of Babylon took him to Babylon, and put him in prison till the day of his death.
JER|52|12|In the fifth month, on the tenth day of the month- that was the nineteenth year of King Nebuchadnezzar, king of Babylon- Nebuzaradan the captain of the bodyguard, who served the king of Babylon, entered Jerusalem.
JER|52|13|And he burned the house of the LORD, and the king's house and all the houses of Jerusalem; every great house he burned down.
JER|52|14|And all the army of the Chaldeans, who were with the captain of the guard, broke down all the walls around Jerusalem.
JER|52|15|And Nebuzaradan the captain of the guard carried away captive some of the poorest of the people and the rest of the people who were left in the city and the deserters who had deserted to the king of Babylon, together with the rest of the artisans.
JER|52|16|But Nebuzaradan the captain of the guard left some of the poorest of the land to be vinedressers and plowmen.
JER|52|17|And the pillars of bronze that were in the house of the LORD, and the stands and the bronze sea that were in the house of the LORD, the Chaldeans broke in pieces, and carried all the bronze to Babylon.
JER|52|18|And they took away the pots and the shovels and the snuffers and the basins and the dishes for incense and all the vessels of bronze used in the temple service;
JER|52|19|also the small bowls and the fire pans and the basins and the pots and the lampstands and the dishes for incense and the bowls for drink offerings. What was of gold the captain of the guard took away as gold, and what was of silver, as silver.
JER|52|20|As for the two pillars, the one sea, the twelve bronze bulls that were under the sea, and the stands, which Solomon the king had made for the house of the LORD, the bronze of all these things was beyond weight.
JER|52|21|As for the pillars, the height of the one pillar was eighteen cubits, its circumference was twelve cubits, and its thickness was four fingers, and it was hollow.
JER|52|22|On it was a capital of bronze. The height of the one capital was five cubits. A network and pomegranates, all of bronze, were around the capital. And the second pillar had the same, with pomegranates.
JER|52|23|There were ninety-six pomegranates on the sides; all the pomegranates were a hundred upon the network all around.
JER|52|24|And the captain of the guard took Seraiah the chief priest, and Zephaniah the second priest, and the three keepers of the threshold;
JER|52|25|and from the city he took an officer who had been in command of the men of war, and seven men of the king's council, who were found in the city; and the secretary of the commander of the army who mustered the people of the land; and sixty men of the people of the land, who were found in the midst of the city.
JER|52|26|And Nebuzaradan the captain of the guard took them and brought them to the king of Babylon at Riblah.
JER|52|27|And the king of Babylon struck them down, and put them to death at Riblah in the land of Hamath. So Judah was taken into exile out of its land.
JER|52|28|This is the number of the people whom Nebuchadnezzar carried away captive: in the seventh year, 3,023 Judeans;
JER|52|29|in the eighteenth year of Nebuchadnezzar he carried away captive from Jerusalem 832 persons;
JER|52|30|in the twenty-third year of Nebuchadnezzar, Nebuzaradan the captain of the guard carried away captive of the Judeans 745 persons; all the persons were 4,600.
JER|52|31|And in the thirty-seventh year of the exile of Jehoiachin king of Judah, in the twelfth month, on the twenty-fifth day of the month, Evil-merodach king of Babylon, in the year that he became king, lifted up the head of Jehoiachin king of Judah and brought him out of prison.
JER|52|32|And he spoke kindly to him, and gave him a seat above the seats of the kings who were with him in Babylon.
JER|52|33|So Jehoiachin put off his prison garments. And every day of his life he dined regularly at the king's table,
JER|52|34|and for his allowance, a regular allowance was given him by the king according to his daily need, until the day of his death as long as he lived.
