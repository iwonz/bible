1SAM|1|1|以法莲 山区有一个 拉玛 的 琐非 人 ，名叫 以利加拿 ，他是 苏弗 的玄孙， 托户 的曾孙， 以利户 的孙子， 耶罗罕 的儿子，是 以法莲 人。
1SAM|1|2|他有两个妻子：一个名叫 哈拿 ，另一个名叫 毗尼拿 。 毗尼拿 有孩子， 哈拿 却没有孩子。
1SAM|1|3|这人每年从本城上到 示罗 ，敬拜万军之耶和华，向他献祭。在那里有 以利 的两个儿子 何弗尼 和 非尼哈 当耶和华的祭司。
1SAM|1|4|每逢献祭的日子， 以利加拿 把祭肉分给他的妻子 毗尼拿 和 毗尼拿 所生的儿女。
1SAM|1|5|他给 哈拿 的却是双分，因为他爱 哈拿 。耶和华却不使 哈拿 生育。
1SAM|1|6|她的对头 毗尼拿 因耶和华不使 哈拿 生育，就常常惹她发怒，要使她生气。
1SAM|1|7|年年都是如此。每当她上到耶和华殿的时候， 毗尼拿 就这样惹她发怒，以致她哭泣不吃饭。
1SAM|1|8|她丈夫 以利加拿 对她说：“ 哈拿 ，你为何哭泣？为何不吃饭？为何伤心难过呢？有我不比有十个儿子更好吗？”
1SAM|1|9|他们在 示罗 吃喝完了， 哈拿 就站起来。祭司 以利 坐在耶和华殿门框旁边的位子上。
1SAM|1|10|哈拿 心里愁苦，就痛痛哭泣，向耶和华祈祷。
1SAM|1|11|她许愿说：“万军之耶和华啊，你若垂顾你使女的苦情，眷念不忘你的使女，赐你的使女一个子嗣，我必使他终生归给耶和华，不用剃刀剃他的头。”
1SAM|1|12|哈拿 在耶和华面前不住地祈祷， 以利 注意她的嘴。
1SAM|1|13|哈拿 心中默祷，只动嘴唇，听不到她的声音，因此 以利 以为她喝醉了。
1SAM|1|14|以利 对她说：“你要醉到几时呢？不要再喝酒了！”
1SAM|1|15|哈拿 回答说：“我主啊，不是这样。我是心里愁苦的妇人，清酒烈酒都没有喝，只在耶和华面前倾心吐意。
1SAM|1|16|不要将你的使女看作不正经的女子。我因极其难过和生气，所以一直祷告到如今。”
1SAM|1|17|以利 回答说：“平平安安地回去吧。愿 以色列 的上帝允准你向他所求的！”
1SAM|1|18|哈拿 说：“愿你的婢女在你眼前蒙恩。”于是妇人上路，去吃饭，脸上不再带愁容了。
1SAM|1|19|他们清早起来，在耶和华面前敬拜，就回去，往 拉玛 自己的家里。 以利加拿 和妻子 哈拿 同房，耶和华顾念 哈拿 。
1SAM|1|20|时候到了， 哈拿 怀孕生了一个儿子， 哈拿 给他起名叫 撒母耳 ，说：“这是我从耶和华那里求来的。”
1SAM|1|21|以利加拿 和他全家都上去，要向耶和华献年祭和还愿祭。
1SAM|1|22|哈拿 却没有上去，因为她对丈夫说：“等孩子断了奶，我就带他上去朝见耶和华，让他永远住在那里。”
1SAM|1|23|她丈夫 以利加拿 对她说：“就照你看为好的去做吧！可以留到儿子断了奶，愿耶和华应验他的话。”于是妇人留在家里乳养儿子，直到断了奶。
1SAM|1|24|断奶之后，她就带着孩子，连同一头三岁的公牛 ，一伊法细面 ，一皮袋酒，上 示罗 耶和华的殿去。那时，孩子还小。
1SAM|1|25|他们宰了公牛，就领孩子到 以利 面前。
1SAM|1|26|妇人说：“我主啊，请容许我说，我向你，我的主起誓，从前在你这里站着祈求耶和华的那妇人就是我。
1SAM|1|27|我祈求为要得这孩子，耶和华已将我向他所求的赐给我了。
1SAM|1|28|所以，我将这孩子献给耶和华，使他终生归给耶和华。” 他就在那里敬拜耶和华。
1SAM|2|1|哈拿 祷告说： “我的心因耶和华快乐， 我的角因耶和华高举。 我的口向仇敌张开； 我因你的救恩欢欣。
1SAM|2|2|“没有一位圣者像耶和华， 除你以外没有别的了， 也没有磐石像我们的上帝。
1SAM|2|3|不要夸口说骄傲的话， 也不要口出狂妄的言语， 因耶和华是有知识的上帝， 人的行为被他衡量。
1SAM|2|4|勇士的弓折断， 跌倒的人以力量束腰。
1SAM|2|5|饱足的人作雇工求食； 饥饿的人也不再饥饿。 不生育的生了七个； 儿女多的反倒孤独。
1SAM|2|6|耶和华使人死，也使人活， 使人下阴间，也使人往上升。
1SAM|2|7|耶和华使人贫穷，也使人富足； 使人降卑，也使人升高。
1SAM|2|8|他从灰尘里抬举贫寒人， 从粪堆中提拔贫穷人， 使他们与贵族同坐， 继承荣耀的座位。 地的柱子属耶和华， 他将世界立在其上。
1SAM|2|9|“他必保护他圣民的脚步， 但恶人却在黑暗中毁灭， 因为人不是靠力量得胜。
1SAM|2|10|与耶和华相争的，必被打碎； 他必从天上打雷攻击他们。 耶和华审判地极的人， 将力量赐给所立的王， 高举受膏者的角。”
1SAM|2|11|以利加拿 往 拉玛 回自己的家去了。那孩子在 以利 祭司面前事奉耶和华。
1SAM|2|12|以利 的两个儿子是无赖，不认识耶和华。
1SAM|2|13|这二祭司对待百姓的规矩是这样：凡有人献祭，正煮肉的时候，祭司的仆人就手拿三齿的叉子来，
1SAM|2|14|将叉子往盆里，或锅里，或釜里，或壶里一插，插上来的肉，祭司都拿了去。他们对所有上到 示罗 的 以色列 人都这样做。
1SAM|2|15|甚至在未烧脂肪之前，祭司的仆人就来对献祭的人说：“把肉给祭司，让他烤吧。他不要拿你煮过的肉，要生的。”
1SAM|2|16|献祭的人若说：“他们必须先烧脂肪，然后你才可以随意拿。”仆人就说：“不，你立刻给我，不然我就要抢了。”
1SAM|2|17|这些年轻人的罪在耶和华面前非常严重，因为这些人藐视耶和华的祭物。
1SAM|2|18|那时， 撒母耳 还是孩子，穿着细麻布的以弗得，侍立在耶和华面前。
1SAM|2|19|他母亲每年为他做一件小外袍，同丈夫上来献年祭的时候带来给他。
1SAM|2|20|以利 为 以利加拿 和他妻子祝福，说：“愿耶和华由这妇人再赐你后裔，代替从耶和华求来的孩子。”他们就回自己的地方去了。
1SAM|2|21|耶和华眷顾 哈拿 ，她就怀孕生了三个儿子，两个女儿。那孩子 撒母耳 在耶和华面前渐渐长大。
1SAM|2|22|以利 年纪老迈，听见他两个儿子对 以色列 众人所做一切的事，又听见他们与会幕门前伺候的妇人同寝，
1SAM|2|23|就对他们说：“你们为何做这样的事呢？我从这众百姓听见了你们的恶行。
1SAM|2|24|我儿啊，不可这样！我听到耶和华的百姓传出你们不好的名声 。
1SAM|2|25|人若得罪人，有上帝 可以裁决；人若得罪耶和华，谁能为他代求呢？”然而他们还是不听父亲的话，因为耶和华想要他们死。
1SAM|2|26|撒母耳 这孩子渐渐长大，耶和华与人越发喜爱他。
1SAM|2|27|有神人来见 以利 ，对他说：“耶和华如此说：‘你祖宗的家在 埃及 法老家 的时候，我不是向他们显现吗？
1SAM|2|28|在 以色列 众支派中，我不是拣选他作我的祭司，上我的祭坛，烧香，在我面前穿以弗得吗？我不是将 以色列 人所献的火祭都赐给你祖宗的家吗？
1SAM|2|29|你们为何践踏我所吩咐献在我居所的祭物和供物呢 ？你为何尊重你的儿子过于尊重我，将我百姓 以色列 所献美好的祭物都拿去养肥你们自己呢？’
1SAM|2|30|因此，耶和华－ 以色列 的上帝说：‘我确实说过，你和你祖宗的家必永远行在我面前，但现在耶和华却说，我绝不会这样做。因为尊重我的，我必尊重他；藐视我的，他必被轻视。
1SAM|2|31|看哪，日子将到，我要折断你的膀臂和你祖宗家的膀臂，使你家中没有一个老年人。
1SAM|2|32|你在 以色列 人享福的时候必看见我居所的衰败 ，你家中必永远没有一个老年人。
1SAM|2|33|你家中的人，我没有从我坛前剪除的，必使你眼睛失明，心中忧伤。你家中所添的人口都必夭折。
1SAM|2|34|你的两个儿子 何弗尼 、 非尼哈 所遭遇的事是给你的预兆：他们二人必在同一日死亡。
1SAM|2|35|我要为自己立一个忠心的祭司，他行事必照我的心、如我的意。我要为他建立坚固的家，他必天天行走在我受膏者的面前。
1SAM|2|36|你家所剩下的人都必来叩拜他，求一块银子，一个饼，说：求你给我一个祭司的职分，好使我得点饼吃。’”
1SAM|3|1|那孩子 撒母耳 在 以利 面前事奉耶和华。在那些日子，耶和华的言语稀少，不常有异象。
1SAM|3|2|那时， 以利 在自己的地方睡觉；他眼目开始昏花，不能看见。
1SAM|3|3|上帝的灯还没有熄灭， 撒母耳 睡在耶和华的殿内，上帝的约柜就在那里。
1SAM|3|4|耶和华呼唤 撒母耳 ， 撒母耳 说：“我在这里！”
1SAM|3|5|他跑到 以利 那里，说：“你叫我吗？我在这里。” 以利 说：“我没有叫你，回去睡吧。”他就回去睡了。
1SAM|3|6|耶和华又呼唤 撒母耳 。 撒母耳 起来，到 以利 那里，说：“你叫我吗？我在这里。” 以利 说：“我儿，我没有叫你，回去睡吧。”
1SAM|3|7|那时 撒母耳 还未认识耶和华，耶和华的话也未曾向他启示。
1SAM|3|8|耶和华第三次再呼唤 撒母耳 。 撒母耳 起来，到 以利 那里，说：“你叫我吗？我在这里。” 以利 才明白是耶和华呼唤这小孩。
1SAM|3|9|以利 对 撒母耳 说：“你回去睡吧。他若再叫你，你就说：‘耶和华啊，请说，仆人敬听！’” 撒母耳 就回去，仍睡在原处。
1SAM|3|10|耶和华来站着，像前几次呼唤：“ 撒母耳 ！ 撒母耳 ！” 撒母耳 说：“请说，仆人敬听！”
1SAM|3|11|耶和华对 撒母耳 说：“看哪，我在 以色列 中必行一件事，凡听见的人都必双耳齐鸣。
1SAM|3|12|我指着 以利 家所说的话，到了时候，必从头到尾应验在 以利 身上。
1SAM|3|13|我曾告诉他，我必永远惩罚他的家，因为他知道自己的儿子作恶，亵渎上帝 ，却不禁止他们。
1SAM|3|14|所以我向 以利 家起誓：‘ 以利 家的罪孽，就是献祭物和供物，也永不得赎。’”
1SAM|3|15|撒母耳 睡到天亮，就开了耶和华殿的门。 撒母耳 害怕，不敢将异象告诉 以利 。
1SAM|3|16|以利 呼唤 撒母耳 说：“我儿 撒母耳 ！” 撒母耳 说：“我在这里！”
1SAM|3|17|以利 说：“他对你说了什么话，你不要向我隐瞒。你若将他对你所说的话向我隐瞒一句，愿上帝重重惩罚你。”
1SAM|3|18|撒母耳 就把一切话都告诉 以利 ，并没有隐瞒。 以利 说：“他是耶和华，愿他照他看为好的去做。”
1SAM|3|19|撒母耳 长大了，耶和华与他同在，使他所说的话一句都不落空。
1SAM|3|20|从 但 到 别是巴 ，所有的 以色列 人都知道耶和华立 撒母耳 为先知。
1SAM|3|21|耶和华又在 示罗 显现，因为耶和华在 示罗 藉他的话向 撒母耳 启示他自己。
1SAM|4|1|撒母耳 的话传遍了全 以色列 。 以色列 人出去与 非利士 人打仗，安营在 以便．以谢 ， 非利士 人安营在 亚弗 。
1SAM|4|2|非利士 人向 以色列 人摆阵。两军交战的时候， 以色列 人败在 非利士 人面前； 非利士 人在战场上杀了他们约四千人。
1SAM|4|3|百姓回到营里， 以色列 的长老说：“耶和华今日为何使我们败在 非利士 人面前呢？我们要将耶和华的约柜从 示罗 抬到我们这里来，好让他来到我们中间，救我们脱离敌人的手掌。”
1SAM|4|4|于是百姓派人到 示罗 ，从那里将坐在二基路伯上万军之耶和华的约柜抬来。 以利 的两个儿子 何弗尼 、 非尼哈 也与上帝的约柜同来。
1SAM|4|5|耶和华的约柜到了营中，全 以色列 就大声欢呼，连地都震动。
1SAM|4|6|非利士 人听见欢呼的声音，就说：“为何 希伯来 人在营里这么大声欢呼呢？”他们知道耶和华的约柜到了营中。
1SAM|4|7|非利士 人就惧怕，说：“有神明到了他们营中。”又说：“我们有祸了！从来不曾有这样的事。
1SAM|4|8|我们有祸了！谁能救我们脱离这些大能之神明的手呢？从前在旷野用各样灾祸击打 埃及 人的，就是这些神明。
1SAM|4|9|非利士 人哪，要刚强，要作大丈夫，免得作 希伯来 人的奴仆，如同他们作你们的奴仆一样。你们要作大丈夫，与他们争战。”
1SAM|4|10|非利士 人进攻， 以色列 人败了，各往自己的家逃跑。被杀的人很多， 以色列 倒下的步兵有三万。
1SAM|4|11|上帝的约柜被掳去， 以利 的两个儿子 何弗尼 、 非尼哈 也都被杀了。
1SAM|4|12|有一个 便雅悯 人从战场上逃跑，衣服撕裂，头蒙灰尘，当日来到 示罗 。
1SAM|4|13|他到了的时候，看哪， 以利 正坐在路旁的位子上观望，为上帝的约柜心里担忧。那人进城报信，全城的人就都呼喊起来。
1SAM|4|14|以利 听见呼喊的声音就说：“这喧嚷的声音是什么呢？”那人急忙来报信给 以利 。
1SAM|4|15|那时 以利 九十八岁了，两眼发直，不能看见。
1SAM|4|16|那人对 以利 说：“我是从战场上来的，今日刚从战场上逃回来。” 以利 说：“我儿，事情怎样了？”
1SAM|4|17|报信的回答说：“ 以色列 人在 非利士 人面前逃跑，百姓中被杀的很多！你的两个儿子 何弗尼 和 非尼哈 也都死了，并且上帝的约柜已经被掳去了。”
1SAM|4|18|他一提到上帝的约柜， 以利 就从城门旁自己的位子上往后跌倒，折断颈项而死，因为他年纪老迈，身体沉重。 以利 作 以色列 的士师四十年。
1SAM|4|19|以利 的媳妇， 非尼哈 的妻子怀孕将到产期，她听见上帝的约柜被掳，公公和丈夫都死了，就曲身生产，极其疼痛。
1SAM|4|20|她将要死的时候，旁边站着的妇人们对她说：“不要怕！你生了男孩了。”她不回答，也不放在心上。
1SAM|4|21|她给孩子起名叫 以迦博 ，说：“荣耀离开 以色列 了！”这是因为上帝的约柜被掳去，又因为她公公和丈夫都死了。
1SAM|4|22|她又说：“荣耀离开 以色列 ，因为上帝的约柜被掳去了。”
1SAM|5|1|非利士 人掳去上帝的约柜，从 以便．以谢 带到 亚实突 。
1SAM|5|2|非利士 人掳了上帝的约柜，带进 大衮 庙，放在 大衮 的旁边。
1SAM|5|3|次日， 亚实突 人清早起来，看哪， 大衮 仆倒在耶和华的约柜前，脸伏于地，他们就扶起 大衮 ，把它放回原处。
1SAM|5|4|又次日，他们清早起来，看哪， 大衮 仆倒在耶和华的约柜前，脸伏于地，并且 大衮 的头和两手都在门槛上折断，只剩下 大衮 的躯干。
1SAM|5|5|因此， 大衮 的祭司和所有进 大衮 庙的人，都不踏 亚实突 的 大衮 庙的门槛，直到今日。
1SAM|5|6|耶和华的手重重击打 亚实突 人，使他们恐惧，使 亚实突 和 亚实突 周围的人都生痔疮。
1SAM|5|7|亚实突 人见这情况，就说：“ 以色列 上帝的约柜不可留在我们这里，因为他的手重重击打我们和我们的神明 大衮 ”。
1SAM|5|8|他们就派人去请 非利士 的众领袖来聚集，对他们说：“我们向 以色列 上帝的约柜应当怎样做呢？”他们说：“可以把 以色列 上帝的约柜运到 迦特 去。”于是他们把 以色列 上帝的约柜运到那里。
1SAM|5|9|运到之后，耶和华的手击打那城，使那城的人非常惊慌，无论大小都生痔疮。
1SAM|5|10|他们就把上帝的约柜送到 以革伦 。上帝的约柜到了 以革伦 ， 以革伦 人就呼喊说：“他们把 以色列 上帝的约柜运到我这里，要害我和我的百姓！”
1SAM|5|11|于是他们派人去请 非利士 的众领袖来，说：“请你们把 以色列 上帝的约柜送回原处，免得害死我和我的百姓！”原来上帝的手重重攻击那城，死亡的恐惧弥漫全城，
1SAM|5|12|没有死的人都受痔疮的折磨。城里的哀声上达于天。
1SAM|6|1|耶和华的约柜在 非利士 人之地七个月。
1SAM|6|2|非利士 人召了祭司和占卜的来，说：“我们向耶和华的约柜应当怎样做呢？请指示我们要用什么方法把约柜送回原处。”
1SAM|6|3|他们说：“若要将 以色列 上帝的约柜送回去，不可空手送回，一定要给他献赔罪的礼物，然后你们才可以得痊愈，并且知道他的手为何不离开你们。”
1SAM|6|4|非利士 人说：“应当用什么献为赔罪的礼物呢？”他们说：“当按照 非利士 领袖的数目，献五个金痔疮和五个金老鼠，因为你们众人和领袖所遭遇的都是一样的灾祸。
1SAM|6|5|当制造你们痔疮的像和毁坏田地老鼠的像，并要将荣耀归给 以色列 的上帝，或者他向你们和你们的神明，以及你们的田地，把手放轻些。
1SAM|6|6|你们为何硬着心，像 埃及 人和法老硬着心一样呢？上帝岂不是严厉对付 埃及 ，使 埃及 人释放 以色列 人，他们就走了吗？
1SAM|6|7|现在你们应当造一辆新车，把两头未曾负轭，还在哺乳的母牛套在车上，赶牛犊离开母牛，回家去。
1SAM|6|8|你们要把耶和华的约柜放在车上，把所献赔罪的金器装在匣子里，放在柜旁，送走柜子，让它去。
1SAM|6|9|你们要观察：车若直行过 以色列 的边界，上到 伯．示麦 去，这大灾祸就是耶和华降在我们身上的；若不然，我们就知道，这不是他的手击打我们，而是我们偶然遭遇的。”
1SAM|6|10|非利士 人就照样做了。他们取了两头哺乳的母牛套在车上，把牛犊关在家里，
1SAM|6|11|把耶和华的约柜和装金老鼠以及金痔疮像的匣子都放在车上。
1SAM|6|12|牛直行大路，在往 伯．示麦 的一条大道上，一面走一面叫，不偏左右。 非利士 的领袖跟在后面，直到 伯．示麦 的地界。
1SAM|6|13|那时， 伯．示麦 人正在平原收割麦子，举目看见约柜，就欢欢喜喜地迎见它。
1SAM|6|14|车到了 伯．示麦 人 约书亚 的田间，就在那里停了。在那里有一块大磐石，他们把车的木头劈了，把两头母牛献给耶和华为燔祭。
1SAM|6|15|利未 人将耶和华的约柜和柜子旁边装金器的匣子拿下来，放在大磐石上。当日 伯．示麦 人献上燔祭，又献其他祭物给耶和华。
1SAM|6|16|非利士 人的五个领袖看见了，当日就回 以革伦 去。
1SAM|6|17|非利士 人献给耶和华作赔罪的金痔疮像如下：一个为 亚实突 ，一个为 迦萨 ，一个为 亚实基伦 ，一个为 迦特 ，一个为 以革伦 。
1SAM|6|18|金老鼠的数目是按照 非利士 五个领袖的城镇，就是坚固的城镇和乡村，以及大磐石。这磐石是安放耶和华约柜的，到今日还在 伯．示麦 人 约书亚 的田间。
1SAM|6|19|耶和华击杀 伯．示麦 人，因为他们观看他的约柜。他击杀了百姓七十人 。百姓因耶和华大大击杀他们，就哀哭了。
1SAM|6|20|伯．示麦 人说：“谁能在耶和华这位圣洁的上帝面前侍立呢？这约柜可以从我们这里上到谁那里去呢？”
1SAM|6|21|于是他们派使者到 基列．耶琳 的居民那里，说：“ 非利士 人将耶和华的约柜送回来了，你们下来将约柜接了，上到你们那里去吧！”
1SAM|7|1|基列．耶琳 人就来了，将耶和华的约柜接上去，抬到山上 亚比拿达 的家中，将他儿子 以利亚撒 分别为圣，看守耶和华的约柜。
1SAM|7|2|从约柜留在 基列．耶琳 的那天起，经过了许多日子，有二十年； 以色列 全家都哀哭归向耶和华。
1SAM|7|3|撒母耳 对 以色列 全家说：“你们若全心回转归向耶和华，就要从你们中间除掉外邦的神明和 亚斯她录 ，预备你们的心归向耶和华，单单事奉他，他必救你们脱离 非利士 人的手。”
1SAM|7|4|以色列 人就除掉诸 巴力 和 亚斯她录 ，单单事奉耶和华。
1SAM|7|5|撒母耳 说：“要召集 以色列 众人到 米斯巴 去，我好为你们向耶和华祷告。”
1SAM|7|6|他们就聚集在 米斯巴 ，打水浇在耶和华面前。当日他们禁食，说：“我们得罪了耶和华。” 撒母耳 在 米斯巴 作 以色列 人的士师。
1SAM|7|7|非利士 人听见 以色列 人聚集在 米斯巴 ， 非利士 的领袖就上来要攻击 以色列 。 以色列 人听见，就惧怕 非利士 人。
1SAM|7|8|以色列 人对 撒母耳 说：“愿你不住为我们呼求耶和华－我们的上帝，救我们脱离 非利士 人的手。”
1SAM|7|9|撒母耳 就把一只吃奶的羔羊献给耶和华作全牲的燔祭，为 以色列 人呼求耶和华，耶和华就应允他。
1SAM|7|10|撒母耳 正献燔祭的时候， 非利士 人前来要与 以色列 争战。当日，耶和华打雷，发出极大的声音，使 非利士 人溃乱，他们就败在 以色列 面前。
1SAM|7|11|以色列 人从 米斯巴 出来，追赶 非利士 人，击杀他们，直到 伯．甲 的下边。
1SAM|7|12|撒母耳 拿一块石头立在 米斯巴 和 善 的中间，给石头起名叫 以便．以谢 ，说：“到如今耶和华都帮助我们。”
1SAM|7|13|因此， 非利士 人被制伏了，不再入侵 以色列 境内。 撒母耳 有生之年，耶和华的手攻击 非利士 人。
1SAM|7|14|非利士 人所夺取 以色列 的城镇，从 以革伦 直到 迦特 ，都归回 以色列 了。 以色列 也从 非利士 人手中收回这些城所属的地界。那时 以色列 与 亚摩利 人和平相处。
1SAM|7|15|撒母耳 一生作 以色列 的士师。
1SAM|7|16|他每年巡行到 伯特利 、 吉甲 、 米斯巴 ，在这些地方审判 以色列 人。
1SAM|7|17|随后他回到 拉玛 ，因为他的家在那里；他在那里审判 以色列 人，并且在那里为耶和华筑了一座坛。
1SAM|8|1|撒母耳 年纪老迈，就立他的儿子作 以色列 的士师。
1SAM|8|2|他的长子名叫 约珥 ，次子名叫 亚比亚 ；他们在 别是巴 作士师。
1SAM|8|3|他的儿子不行他的道，贪图财利，收取贿赂，屈枉正直。
1SAM|8|4|以色列 的长老都聚集在 拉玛 ，来到 撒母耳 那里，
1SAM|8|5|对他说：“看哪，你年纪老了，你的儿子又不行你的道。现在请你为我们立一个王治理我们，像列国一样。”
1SAM|8|6|撒母耳 不喜悦他们说“立一个王治理我们”，他就向耶和华祷告。
1SAM|8|7|耶和华对 撒母耳 说：“你只管听从百姓向你说的一切话，因为他们不是厌弃你，而是厌弃我，不要我作他们的王。
1SAM|8|8|自从我领他们出 埃及 的日子到如今，他们离弃我，事奉别神；正像他们从前所做的一切事，现在他们也照样向你做了。
1SAM|8|9|现在你只管听从他们的话，不过要严厉警告他们，告诉他们将来王会用什么方式管辖他们。”
1SAM|8|10|撒母耳 将耶和华一切的话转告求他立王的百姓。
1SAM|8|11|他说：“管辖你们的王必用这样的方式：他必派你们的儿子为他驾车，赶马，在他的战车前奔跑。
1SAM|8|12|他要为自己立千夫长、五十夫长；耕种他的田地，收割他的庄稼；打造他的兵器和车上的器械。
1SAM|8|13|他必叫你们的女儿为他制造香膏，作厨师与烤饼的，
1SAM|8|14|也必取你们最好的田地、葡萄园、橄榄园，赐给他的臣仆。
1SAM|8|15|你们的粮食和葡萄园所出产的，他必征收十分之一给他的官员和臣仆，
1SAM|8|16|又必叫你们的仆人婢女，健壮的青年和你们的驴为他做工。
1SAM|8|17|你们的羊群，他必征收十分之一，你们自己也必作他的仆人。
1SAM|8|18|那日，你们必因自己所选的王哀求耶和华，但那日耶和华却不应允你们。”
1SAM|8|19|百姓却不肯听 撒母耳 的话，说：“不！我们一定要一个王治理我们，
1SAM|8|20|使我们像列国一样，有王治理我们，率领我们，为我们争战。”
1SAM|8|21|撒母耳 听见百姓这一切话，就禀告给耶和华听。
1SAM|8|22|耶和华对 撒母耳 说：“你只管听从他们的话，为他们立一个王。” 撒母耳 对 以色列 人说：“去，你们各归各城吧！”
1SAM|9|1|有一个 便雅悯 人名叫 基士 ，是 便雅悯 人 亚斐亚 的玄孙， 比歌拉 的曾孙， 洗罗 的孙子， 亚别 的儿子，是个大能的勇士 。
1SAM|9|2|他有一个儿子名叫 扫罗 ，又健壮、又英俊，在 以色列 人中没有一个可以与他相比；他比众百姓高出一个头 。
1SAM|9|3|扫罗 的父亲 基士 丢失了几匹母驴，他就吩咐儿子 扫罗 说：“起来，带一个仆人去寻找驴子。”
1SAM|9|4|扫罗 走过 以法莲 山区，又过 沙利沙 地，都没有找着。他们走过 沙琳 地，驴不在那里，又走过 便雅悯 地，也没有找到。
1SAM|9|5|到了 苏弗 地， 扫罗 对跟随他的仆人说：“我们不如回去，免得我父亲不为驴挂虑，反为我们担忧。”
1SAM|9|6|仆人对他说：“看哪，这城里有一位神人，受人敬重，凡他所说的全都应验。现在让我们到他那里去，或者他能指示我们当走的路。”
1SAM|9|7|扫罗 对仆人说：“看哪，我们若去，送什么给那人呢？我们袋子里的食物都吃完了，也没有礼物可以送给神人，我们还有些什么呢？”
1SAM|9|8|仆人又回答 扫罗 说：“看哪，我手里还有四分之一舍客勒的银子，可以送给神人，请他指示我们当走的路。”
1SAM|9|9|从前 以色列 中，若有人去求问上帝，就这么说：“来，我们到先见那里去吧！”因现在的先知，从前称为先见。
1SAM|9|10|扫罗 对仆人说：“好主意！来，我们去吧。”于是他们往神人所住的城里去了。
1SAM|9|11|他们上坡要进城，遇见几个少女出来打水，就问她们说：“先见有没有在这里呢？”
1SAM|9|12|她们回答说：“有的，看哪，他就在你们前面。快！他今日正来到城里，因为今日百姓要在丘坛献祭。
1SAM|9|13|你们一进城，他还没有上丘坛吃祭物之前，就会遇见他。因为他没有到，百姓不能吃，必须等他先为祭物祝谢，然后受邀的人才可以吃。现在就上去吧，因为这时候你们会遇见他。”
1SAM|9|14|他们就上到那城，进入城中的时候，看哪， 撒母耳 正迎着他们来，要上丘坛去。
1SAM|9|15|扫罗 还没有到的前一日，耶和华已经对 撒母耳 启示说：
1SAM|9|16|“明日这时候，我必使一个人从 便雅悯 地到你这里来，你要膏他作我百姓 以色列 的君王。他必救我的百姓脱离 非利士 人的手，因为我眷顾我的百姓 ，他们的哀声已上达于我。”
1SAM|9|17|撒母耳 看见 扫罗 的时候，耶和华对他说：“看哪，这就是我对你所说的人，他必治理我的百姓。”
1SAM|9|18|扫罗 在城门中走到 撒母耳 跟前，说：“请告诉我，先见的家在哪里？”
1SAM|9|19|撒母耳 回答扫罗说：“我就是先见。你在我前面先上丘坛去，因为你们今日必跟我同席。明日早晨我送你走，会把你心里一切的事都告诉你。
1SAM|9|20|至于你前三日所丢失的几匹母驴，你心里不必挂虑，都已经找到了。 以色列 众人所仰慕的是谁呢？不是仰慕你和你父的全家吗？”
1SAM|9|21|扫罗 回答说：“我不是 以色列 支派中最小的 便雅悯 人吗？我的家族不是 便雅悯 支派中最小的家族吗？你为何对我说这样的话呢？”
1SAM|9|22|撒母耳 领 扫罗 和他的仆人进了大厅，使他们在受邀的人中坐首位；受邀者约有三十个。
1SAM|9|23|撒母耳 对厨师说：“我交给你的那一份祭肉，吩咐你收存的，现在可以拿来。”
1SAM|9|24|厨师就举起祭肉的腿和腿上的部分 ，摆在 扫罗 面前。 撒母耳 说：“看哪，所存留的摆在你面前了。吃吧！因为这是为你保留到这特定的时候的，好让你说，是我请了这百姓来，” 当日， 扫罗 就与 撒母耳 同席。
1SAM|9|25|他们从丘坛下来进城， 撒母耳 和 扫罗 在房顶上说话。
1SAM|9|26|次日他们清早起来。黎明的时候， 撒母耳 呼叫在房顶上的 扫罗 ，说：“起来，我好送你回去。” 扫罗 就起来，和 撒母耳 二人一同到外面去。
1SAM|9|27|二人下到城边， 撒母耳 对 扫罗 说：“你要吩咐仆人先走，仆人走了以后， 你要留在这里，这时候我要将上帝的话传给你听。”
1SAM|10|1|撒母耳 拿一瓶膏油倒在 扫罗 的头上，亲吻他，说：“耶和华岂不是膏你作他产业的君王吗？
1SAM|10|2|你今日离开我之后，会在 便雅悯 境内的 谢撒 ，靠近 拉结 的坟墓，遇见两个人。他们会对你说：‘你要找的几匹母驴已经找到了。看哪，你父亲不为驴子的事挂虑，反为你担忧，说：我为儿子该做些什么呢？’
1SAM|10|3|你从那里往前走，到了 他泊 的橡树那里，会遇见三个往 伯特利 去敬拜上帝的人：一个带着三只小山羊，一个带着三个饼，一个带着一皮袋酒。
1SAM|10|4|他们会向你问安，给你两个饼，你就从他们手中接过来。
1SAM|10|5|然后你要到上帝的山去，在那里有 非利士 的驻军。你到了城里的时候，会遇见一队先知从丘坛下来，前面有鼓瑟的、击鼓的、吹笛的、弹琴的，他们都受感说话。
1SAM|10|6|耶和华的灵必大大感动你，你就与他们一同受感说话，转变成另一个人。
1SAM|10|7|这征兆临到你，你就要趁机做该做的事，因为上帝与你同在。
1SAM|10|8|你要在我以先下到 吉甲 。看哪，我必下到你那里献燔祭和平安祭。你要等候七日，等我到你那里指示你当做的事。”
1SAM|10|9|扫罗 转身离开 撒母耳 ，上帝就改变他，赐给他另一颗心。当日这一切征兆都应验了。
1SAM|10|10|他们来到那座山，看哪，有一队先知遇见 扫罗 。上帝的灵大大感动他，他就在先知中受感说话。
1SAM|10|11|所有先前认识 扫罗 的人看见了，看哪，他和先知一同受感说话，百姓就彼此说：“ 基士 的儿子遇见了什么呢？ 扫罗 也在先知中吗？”
1SAM|10|12|那地方有一个人说：“这些人的父亲是谁呢？”因此就有一句俗语说：“ 扫罗 也在先知中吗？”
1SAM|10|13|扫罗 受感说完了话，就上丘坛去了。
1SAM|10|14|扫罗 的叔叔问 扫罗 和他的仆人说：“你们到哪里去了？”他说：“我们找驴子去了。但我们找不到，就去了 撒母耳 那里。”
1SAM|10|15|扫罗 的叔叔说：“告诉我 撒母耳 对你们说了些什么。”
1SAM|10|16|扫罗 对他的叔叔说：“他明明告诉我们，驴子已经找到了。”至于 撒母耳 所说君王的事， 扫罗 没有告诉叔叔。
1SAM|10|17|撒母耳 召集百姓到 米斯巴 耶和华那里。
1SAM|10|18|他对 以色列 众人说：“耶和华－ 以色列 的上帝如此说：‘我领 以色列 出 埃及 ，救你们脱离 埃及 人的手，以及脱离欺压你们各国之人的手。’
1SAM|10|19|你们今日却厌弃救你们脱离一切灾祸和患难的上帝，对他说：‘求你立一个王治理我们。’现在你们应当按支派和宗族站在耶和华面前。”
1SAM|10|20|于是， 撒母耳 叫 以色列 众支派近前来抽签，抽到了 便雅悯 支派。
1SAM|10|21|然后，他叫 便雅悯 支派按宗族近前来，抽到了 玛特利 族，接着又抽到了 基士 的儿子 扫罗 。众人寻找他却找不到，
1SAM|10|22|就再问耶和华说：“那人来到这里了没有？”耶和华说：“看哪，他藏在物品堆中。”
1SAM|10|23|众人就跑去从那里领他出来。他站在百姓中间，比众百姓高出一个头。
1SAM|10|24|撒母耳 对众百姓说：“你们看到了耶和华所拣选的人吗？众百姓中没有人可以与他相比。”众百姓就欢呼说：“愿王万岁！”
1SAM|10|25|撒母耳 将君王的典章对百姓说明，又记在书上，放在耶和华面前，然后 撒母耳 遣散众百姓，各回自己的家去了。
1SAM|10|26|扫罗 也往 基比亚 自己的家去，有一群心中被上帝感动的勇士跟随他。
1SAM|10|27|但有些无赖之辈说：“这人怎么能救我们呢？”他们就藐视他，不送礼物给他。 扫罗 却保持沉默。
1SAM|11|1|亚扪 人 拿辖 上来，对着 基列 的 雅比 安营。 雅比 众人对 拿辖 说：“你与我们立约，我们就服事你。”
1SAM|11|2|亚扪 人 拿辖 对他们说：“你们若由我挖出你们各人的右眼，以此凌辱 以色列 众人，我就与你们立约。”
1SAM|11|3|雅比 的长老对他说：“求你宽容我们七日，等我们派人到 以色列 的全境去。若没有人来救我们，我们就出来归顺你。”
1SAM|11|4|使者到了 扫罗 住的 基比亚 ，把这事说给百姓听，众百姓就都放声大哭。
1SAM|11|5|看哪， 扫罗 正从田间赶牛回来，说：“百姓为什么哭呢？”众人把 雅比 人的话告诉他。
1SAM|11|6|扫罗 听见这些话，就被上帝的灵催逼，大发怒气。
1SAM|11|7|他把一对牛切成小块，吩咐使者传送到 以色列 全境，说：“凡不出来跟随 扫罗 和 撒母耳 的，就必这样待他的牛。”耶和华使百姓惧怕，他们就都出来如同一人。
1SAM|11|8|扫罗 在 比色 数点他们： 以色列 人有三十万， 犹大 人有三万。
1SAM|11|9|他们对那些来的使者说：“你们要对 基列 的 雅比 人这样说，明天太阳快到中午的时候，你们必得解救。”使者回去告诉 雅比 人，他们就欢喜了。
1SAM|11|10|于是 雅比 人对 亚扪 人说：“明日我们出来归顺你们，可以照你们看为好的待我们。”
1SAM|11|11|第二日， 扫罗 把百姓分为三队，在清晨换岗哨的时候入侵 亚扪 人的军营，击杀他们直到中午的时候。逃脱的人都分散了，甚至没有两个人同在一起。
1SAM|11|12|百姓对 撒母耳 说：“那说‘ 扫罗 岂能作我们的王’的是谁呢？把他们交出来，我们好处死他们。”
1SAM|11|13|扫罗 说：“今日耶和华在 以色列 中施行拯救，所以今日不可处死人。”
1SAM|11|14|撒母耳 对百姓说：“来，我们到 吉甲 去，在那里开始新的王国。”
1SAM|11|15|众百姓到了 吉甲 那里，在耶和华面前拥立 扫罗 为王，又在耶和华面前献平安祭。 扫罗 和 以色列 众人在那里都非常欢喜。
1SAM|12|1|撒母耳 对 以色列 众人说：“看哪，我已听了你们对我所说一切的话，为你们立了一个王。
1SAM|12|2|现在，看哪，有这王行走在你们前面。我已年老发白，看哪，我的儿子都在你们这里。我从幼年直到今日都行走在你们前面。
1SAM|12|3|我在这里，你们要在耶和华和他的受膏者面前为我作证，我夺过谁的牛，抢过谁的驴，欺负过谁，虐待过谁，从谁手里收过贿赂而蒙蔽自己的眼目呢？若有，我必偿还。”
1SAM|12|4|众人说：“你未曾欺负我们，虐待我们，也未曾从任何人手里收过任何东西。”
1SAM|12|5|撒母耳 对他们说：“你们在我手里没有找着什么，有耶和华在你们中间作证，也有他的受膏者今日作证。”他们说 ：“愿耶和华作证。”
1SAM|12|6|撒母耳 对百姓说：“从前立 摩西 和 亚伦 ，又领你们祖先出 埃及 地的是耶和华。
1SAM|12|7|现在你们要站住，让我在耶和华面前，以耶和华向你们和你们祖先所行一切公义的事来和你们争辩。
1SAM|12|8|从前 雅各 到了 埃及 ，后来你们的祖先呼求耶和华，耶和华就差遣 摩西 和 亚伦 领你们的祖先出 埃及 ，来到这地方居住。
1SAM|12|9|他们却忘记耶和华－他们的上帝，他就把他们交给 夏琐 将军 西西拉 的手中，以及 非利士 人和 摩押 王的手中 。于是这些人常来攻击他们。
1SAM|12|10|他们呼求耶和华说：‘我们离弃了耶和华去事奉诸 巴力 和 亚斯她录 ，我们有罪了。现在求你救我们脱离仇敌的手，我们必事奉你。’
1SAM|12|11|耶和华就差遣 耶路巴力 、 比但 、 耶弗他 、 撒母耳 救你们脱离四围仇敌的手，你们才安然居住。
1SAM|12|12|你们见 亚扪 人的王 拿辖 来攻击你们，就对我说：‘不，要有一个王治理我们。’其实耶和华－你们的上帝是你们的王。
1SAM|12|13|现在，看哪，这就是你们所选的、你们所求的王。看哪，耶和华已经为你们立王了。
1SAM|12|14|你们若敬畏耶和华，事奉他，听从他的话，不违背耶和华的命令，你们和治理你们的王也都跟从耶和华－你们的上帝就好了。
1SAM|12|15|倘若不听从耶和华的话，违背他的命令，耶和华的手必攻击你们，像从前攻击你们祖先一样。
1SAM|12|16|现在你们要站住，看耶和华在你们眼前要行的一件大事。
1SAM|12|17|这不是割麦子的时候吗？我求告耶和华，他必打雷降雨，让你们知道并且看出，你们为自己求立王的事在耶和华眼前是犯大罪了。”
1SAM|12|18|于是 撒母耳 求告耶和华，耶和华就在这日打雷降雨，众百姓就非常惧怕耶和华和 撒母耳 。
1SAM|12|19|众百姓对 撒母耳 说：“请你为仆人向耶和华－你的上帝祷告，免得我们死亡，因为我们求立王的事，正是罪上加罪了。”
1SAM|12|20|撒母耳 对百姓说：“不要惧怕！你们虽然行了这恶，却不要偏离耶和华，只要尽心事奉他。
1SAM|12|21|不可偏离去随从那没有益处、不能救人的虚无的神明 ，因为它们是虚无的。
1SAM|12|22|耶和华必因他大名的缘故不撇弃他的子民，因为耶和华喜悦你们作他的子民。
1SAM|12|23|至于我，我如果停止为你们祷告，就得罪耶和华了，我绝不会这样做。我必以善道正路指教你们。
1SAM|12|24|但你们要敬畏耶和华，诚诚实实地尽心事奉他，因你们要留意，他向你们所行的事何等大。
1SAM|12|25|你们若不断作恶，你们和你们的王必一同灭亡。”
1SAM|13|1|扫罗 登基的时候年三十 岁，作 以色列 王二年 。
1SAM|13|2|扫罗 从 以色列 中选出三千人：二千跟随 扫罗 在 密抹 和 伯特利 山区，一千跟随 约拿单 在 便雅悯 的 基比亚 。其余的百姓， 扫罗 打发他们各自回自己的帐棚去了。
1SAM|13|3|约拿单 攻击 非利士 人在 迦巴 的驻军， 非利士 人听见了这事。 扫罗 就在遍地吹角，说：“让 希伯来 人都听见。”
1SAM|13|4|以色列 众人听见 扫罗 攻击 非利士 的驻军，又听见 以色列 为 非利士 人所憎恶，百姓就跟随 扫罗 ，在 吉甲 集合。
1SAM|13|5|非利士 人集合，要与 以色列 人作战。他们有战车三万辆，骑兵六千，士兵像海边的沙那样多。他们上来，在 伯．亚文 东边的 密抹 安营。
1SAM|13|6|以色列 人见自己危急，军队被围攻，百姓就藏在山洞、丛林、岩隙、地窖和深坑中。
1SAM|13|7|有些 希伯来 人过了 约旦河 ，逃到 迦得 和 基列 地。 扫罗 还在 吉甲 ，所有的人都战战兢兢地跟随他。
1SAM|13|8|扫罗 照着 撒母耳 所定的日期等了七日。但是， 撒母耳 还没有来到 吉甲 ，百姓就离开 扫罗 散去了。
1SAM|13|9|于是 扫罗 说：“把燔祭和平安祭带到我这里来。” 扫罗 就献上燔祭。
1SAM|13|10|他刚献完燔祭，看哪， 撒母耳 就到了。 扫罗 出去迎接他，向他问安。
1SAM|13|11|撒母耳 说：“你做了什么事啊？” 扫罗 说：“因为我见百姓离开我散去，你又不照所定的日期来到，而且 非利士 人已在 密抹 集合；
1SAM|13|12|我说：‘现在 非利士 人已经下到 吉甲 来攻击我，可是我还没有向耶和华祷告。’所以我就勉强献上燔祭。”
1SAM|13|13|撒母耳 对 扫罗 说：“你做了糊涂事了，没有遵守耶和华－你上帝吩咐你的命令。不然，耶和华会在 以色列 中坚立你的国度，直到永远。
1SAM|13|14|现在你的国度必不长久。耶和华已经寻着一个合他心意的人，立他作百姓的君王，因为你没有遵守耶和华所吩咐你的。”
1SAM|13|15|撒母耳 就起来，从 吉甲 上到 便雅悯 的 基比亚 。 扫罗 数点跟随他的百姓，约有六百人。
1SAM|13|16|扫罗 和他儿子 约拿单 ，以及跟随他们的百姓，都住在 便雅悯 的 迦巴 ， 非利士 人却在 密抹 安营。
1SAM|13|17|有突击队从 非利士 营中出来，分成三队：一队往 俄弗拉 到 书亚 地去，
1SAM|13|18|一队往 伯．和仑 去，一队往边界，下望朝着旷野的 洗波音谷 。
1SAM|13|19|那时， 以色列 全地找不到一个铁匠，因为 非利士 人说：“恐怕 希伯来 人制造刀枪。”
1SAM|13|20|以色列 众人要磨锄、犁、斧、铲，就各自下到 非利士 人那里去磨。
1SAM|13|21|磨锄或犁的价钱是三分之二舍客勒，磨斧或修整刺棒的价钱是三分之一舍客勒。
1SAM|13|22|所以到了战争的日子，所有跟随 扫罗 和 约拿单 的百姓找不到一个手里有刀有枪的，惟 扫罗 和他儿子 约拿单 有。
1SAM|13|23|非利士 人的一队驻军出来，到 密抹 的隘口。
1SAM|14|1|有一日， 扫罗 的儿子 约拿单 对拿他兵器的青年说：“来，我们过去到 非利士 的驻军那里。”但他没有告诉父亲。
1SAM|14|2|扫罗 在 基比亚 的郊外，坐在 米矶仑 的石榴树下，跟随他的百姓约有六百人。
1SAM|14|3|在那里有 亚希突 的儿子 亚希亚 ，穿着以弗得。 亚希突 是 以迦博 的哥哥， 非尼哈 的儿子， 以利 的孙子。 以利 从前在 示罗 作耶和华的祭司。 约拿单 去了，百姓却不知道。
1SAM|14|4|约拿单 要从隘口过到 非利士 驻军那里去。这隘口两边各有一座齿状峭壁：一座名叫 播薛 ，另一座名叫 西尼 ；
1SAM|14|5|一座向北，对着 密抹 ，一座向南，对着 迦巴 。
1SAM|14|6|约拿单 对拿兵器的青年说：“来，我们过去到那些未受割礼之人的驻军那里，或者耶和华为我们施展能力，因为耶和华使人得胜，不在乎人多人少 。”
1SAM|14|7|拿兵器的对他说：“随你的心意做吧。你上去，看哪，我一定跟随你，与你同心。”
1SAM|14|8|约拿单 说：“看哪，我们要过去到那些人那里，在他们那里展现我们自己。
1SAM|14|9|他们若对我们这么说：‘站住，等我们到你们那里去’，我们就站在原地，不上他们那里去；
1SAM|14|10|但他们若这么说：‘上到我们这里来吧’，我们就上去，因为耶和华把他们交在我们手里了。这就是我们的凭据。”
1SAM|14|11|二人就让 非利士 的驻军看见。 非利士 人说：“看哪， 希伯来 人从躲藏的洞穴里出来了！”
1SAM|14|12|站岗的士兵对 约拿单 和拿兵器的人说：“上到这里来，我们有一件事要告诉你们。” 约拿单 就对拿兵器的人说：“跟我上去，因为耶和华把他们交在 以色列 人手里了。”
1SAM|14|13|约拿单 手脚并用爬上去，拿兵器的人跟随他。 非利士 人仆倒在 约拿单 面前，拿兵器的人跟着他，杀死他们。
1SAM|14|14|约拿单 和拿兵器的人第一次击杀的约有二十人，都在一亩 地的半犁沟之内。
1SAM|14|15|于是在军营、在田野、在众百姓中，人心惶惶，驻军和突击队都战兢；地也震动，这是从上帝那里来的惊恐 。
1SAM|14|16|在 便雅悯 的 基比亚 ， 扫罗 的哨兵观看，看哪， 非利士 全军溃乱，四处乱窜。
1SAM|14|17|扫罗 就对跟随他的百姓说：“你们去数点人数，看是谁从我们这里出去。”他们一数点，看哪， 约拿单 和拿兵器的人不在其中。
1SAM|14|18|那时上帝的约柜 在 以色列 人那里。 扫罗 对 亚希亚 说：“你把上帝的约柜请到这里来。”
1SAM|14|19|扫罗 正与祭司说话的时候， 非利士 营中的骚乱越来越剧烈； 扫罗 就对祭司说：“停手吧！”
1SAM|14|20|扫罗 和所有跟随他的百姓都集合，来到战场，看哪， 非利士 人用刀互相击杀，大大混乱。
1SAM|14|21|那先前由四方来跟随 非利士 人、在他们营中的 希伯来 人，现在也转过来帮助跟随 扫罗 和 约拿单 的 以色列 人了。
1SAM|14|22|那藏在 以法莲 山区的 以色列 众人听说 非利士 人逃跑，就出来紧紧地追击他们。
1SAM|14|23|那日，耶和华使 以色列 人得胜，战争一直打到 伯．亚文 。
1SAM|14|24|那日， 以色列 人非常困惫，因为 扫罗 叫百姓起誓说：“凡不等到晚上我向敌人报完了仇就吃东西的，必受诅咒。”因此所有的百姓都没有尝食物。
1SAM|14|25|所有的百姓 进入树林，见地面上有蜜。
1SAM|14|26|百姓进了树林，看哪，有蜜流出来，却没有人敢用手取蜜入口，因为百姓怕那誓言。
1SAM|14|27|约拿单 没有听见他父亲叫百姓起誓，所以他伸出手中的杖，以杖头蘸在蜂房里，用手取回送入口内，他的眼睛就明亮了。
1SAM|14|28|百姓中有一人对他说：“你父亲曾叫百姓严严地起誓说，今日吃东西的人必受诅咒；因此百姓就疲乏了。”
1SAM|14|29|约拿单 说：“我父亲给这地添麻烦了。你们看，我尝了这一点蜜，眼睛就明亮了。
1SAM|14|30|今日百姓若随意吃了从仇敌夺来的东西，现在击杀的 非利士 人岂不更多吗？”
1SAM|14|31|这日， 以色列 人击杀 非利士 人，从 密抹 直到 亚雅仑 。但百姓非常疲乏，
1SAM|14|32|就急着扑向掠物，夺取牛羊和牛犊，宰于地上，连肉带血吃了。
1SAM|14|33|有人告诉 扫罗 说：“看哪，百姓吃带血的肉，得罪耶和华了。” 扫罗 说：“你们行了诡诈，今日把一块大石头滚到我这里来吧。”
1SAM|14|34|扫罗 又说：“你们分散到百姓中，对他们说，你们各人把牛羊牵到我这里来宰了吃，不可吃带血的肉得罪耶和华。”那夜，所有的百姓把自己手中的牛 牵到那里宰了。
1SAM|14|35|扫罗 为耶和华筑了一座坛，这是他开始为耶和华筑的坛。
1SAM|14|36|扫罗 说：“我们要在夜里下去追赶 非利士 人，抢掠他们，直到天亮，不给他们留下一人。”众百姓说：“你看怎样好就做吧！”祭司说：“我们要先在这里亲近上帝。”
1SAM|14|37|扫罗 求问上帝说：“我可以下去追赶 非利士 人吗？你把他们交在 以色列 人手里吗？”这日上帝没有回答他。
1SAM|14|38|扫罗 说：“百姓中的众领袖，你们都要近前来到这里，查明今日这罪是怎样发生的。
1SAM|14|39|我指着拯救 以色列 的永生的耶和华起誓，就是我儿子 约拿单 犯了罪，他也必被处死。”但众百姓中无人回答他。
1SAM|14|40|扫罗 对 以色列 众人说：“你们站在一边，我与我儿子 约拿单 也站在一边。”百姓对 扫罗 说：“你看怎样好就做吧！”
1SAM|14|41|扫罗 向耶和华－ 以色列 的上帝祷告说：“求你指示正确的答案。”抽中的是 扫罗 和 约拿单 ，百姓尽都无事。
1SAM|14|42|扫罗 说：“你们再抽签，看是我，还是我儿子 约拿单 。”抽中的是 约拿单 。
1SAM|14|43|扫罗 对 约拿单 说：“你告诉我，你做了什么事？” 约拿单 说：“我只是用手中的杖，以杖头蘸了一点蜜尝尝，看哪，我就要死吗？”
1SAM|14|44|扫罗 说：“ 约拿单 哪，你一定要死！若不然，愿上帝重重惩罚我。”
1SAM|14|45|百姓对 扫罗 说：“ 约拿单 在 以色列 中大行拯救，岂可死呢？绝对不可！我们指着永生的耶和华起誓，连他的一根头发也不可落地，因为他今日与上帝一同做事。”于是百姓救 约拿单 免了死亡。
1SAM|14|46|扫罗 上去，不追赶 非利士 人， 非利士 人也回本地去了。
1SAM|14|47|扫罗 执掌 以色列 的国权，攻打他四围所有的仇敌，就是 摩押 人、 亚扪 人、 以东 人和 琐巴 诸王，以及 非利士 人。他无论往何处去，都打败他们。
1SAM|14|48|扫罗 奋勇作战，击败 亚玛力 人，救了 以色列 脱离抢掠他们之人的手。
1SAM|14|49|扫罗 的儿子是 约拿单 、 亦施韦 、 麦基．舒亚 。他的两个女儿：长女名叫 米拉 ，次女名叫 米甲 。
1SAM|14|50|扫罗 的妻子名叫 亚希暖 ，是 亚希玛斯 的女儿。 扫罗 军队的元帅名叫 押尼珥 ，是 扫罗 的叔叔 尼珥 的儿子。
1SAM|14|51|扫罗 的父亲 基士 ， 押尼珥 的父亲 尼珥 ，都是 亚别 的儿子。
1SAM|14|52|扫罗 有生之年常与 非利士 人激烈争战，他看到任何有能力的人或勇士，都招募来跟随他。
1SAM|15|1|撒母耳 对 扫罗 说：“耶和华差遣我膏你为王，治理他的百姓 以色列 ，现在你要听从耶和华的话。
1SAM|15|2|万军之耶和华如此说：‘ 以色列 人从 埃及 上来的时候，在路上 亚玛力 人怎样待他们，怎样抵挡他们，我都要惩罚。
1SAM|15|3|现在你要去攻打 亚玛力 人，灭尽他们所有的，不可怜惜他们，将男女、孩童、吃奶的，以及牛、羊、骆驼和驴全都杀死。’”
1SAM|15|4|于是 扫罗 在 提拉因 召集百姓，数点他们，共有二十万步兵和一万 犹大 人。
1SAM|15|5|扫罗 到了 亚玛力 的京城，在谷中设下埋伏。
1SAM|15|6|扫罗 对 基尼 人说：“你们离开 亚玛力 人下去吧，免得我把你们和 亚玛力 人一同杀灭，因为 以色列 众人从 埃及 上来的时候，你们曾恩待他们。”于是 基尼 人离开了 亚玛力 人。
1SAM|15|7|扫罗 攻打 亚玛力 人，从 哈腓拉 直到 埃及 东边的 书珥 ，
1SAM|15|8|生擒了 亚玛力 王 亚甲 ，用刀杀尽 亚玛力 的众百姓。
1SAM|15|9|扫罗 和百姓却怜惜 亚甲 ，爱惜上好的牛、羊、牛犊、羔羊，以及一切美物，不肯灭绝。但是凡看不上眼和没有价值的，他们尽都杀了。
1SAM|15|10|耶和华的话临到 撒母耳 说：
1SAM|15|11|“我立 扫罗 为王，我感到遗憾，因为他转去不跟从我，不遵守我的命令。” 撒母耳 就很生气，终夜哀求耶和华。
1SAM|15|12|撒母耳 清早起来，去见 扫罗 。有人告诉 撒母耳 说：“ 扫罗 到了 迦密 ，看哪，他在那里为自己立了纪念碑，又转身下到 吉甲 。”
1SAM|15|13|撒母耳 到了 扫罗 那里， 扫罗 对他说：“愿耶和华赐福给你，耶和华的命令我已遵守了。”
1SAM|15|14|撒母耳 说：“我耳中听见有羊叫、牛鸣的声音，又是什么呢？”
1SAM|15|15|扫罗 说：“这是百姓从 亚玛力 人那里带来的，因为他们爱惜上好的牛羊，要献给耶和华－你的上帝。其余的，我们都灭尽了。”
1SAM|15|16|撒母耳 对 扫罗 说：“住口吧！等我把耶和华昨夜向我所说的话告诉你。” 扫罗 说：“请说。”
1SAM|15|17|撒母耳 说：“你虽然看自己为小，你岂不是作了 以色列 诸支派的元首吗？耶和华膏你作了 以色列 的王。
1SAM|15|18|耶和华差遣你，吩咐你说：‘你去除灭那些犯罪的 亚玛力 人，攻打他们，直到把他们完全灭尽。’
1SAM|15|19|你为何没有听从耶和华的话呢？你为何急着扑向掠物，行耶和华眼中看为恶的事呢？”
1SAM|15|20|扫罗 对 撒母耳 说：“我听从了耶和华的话，行了耶和华派我行的路，擒了 亚玛力 王 亚甲 来，灭尽了 亚玛力 人。
1SAM|15|21|百姓却从掠物中取了牛羊，是当灭之物中最好的，要在 吉甲 献给耶和华－你的上帝。”
1SAM|15|22|撒母耳 说： “耶和华喜爱燔祭和祭物， 岂如喜爱人听从他的话呢？ 看哪，听命胜于献祭， 顺从胜于公羊的脂肪。
1SAM|15|23|悖逆与占卜的罪相等， 顽梗与拜偶像的罪孽相同。 因为你厌弃耶和华的命令， 耶和华也厌弃你作王。”
1SAM|15|24|扫罗 对 撒母耳 说：“我有罪了！我违背了耶和华的指示和你的命令；因为我惧怕百姓，听从了他们的话。
1SAM|15|25|现在求你赦免我的罪，同我回去，我好敬拜耶和华。”
1SAM|15|26|撒母耳 对 扫罗 说：“我不同你回去，因为你厌弃耶和华的命令，耶和华也厌弃你作 以色列 的王。”
1SAM|15|27|撒母耳 转身要走， 扫罗 抓住他外袍的衣角，外袍就断裂了。
1SAM|15|28|撒母耳 对他说：“今日耶和华使 以色列 国与你断绝，把这国赐给另一个比你更好的人。
1SAM|15|29|以色列 的大能者必不说谎，也不后悔，因为他不是世人，绝不后悔。”
1SAM|15|30|扫罗 说：“我有罪了。现在求你在我百姓的长老和 以色列 人面前尊重我，同我回去，我好敬拜耶和华－你的上帝。”
1SAM|15|31|于是 撒母耳 转身跟随 扫罗 回去， 扫罗 就敬拜耶和华。
1SAM|15|32|撒母耳 说：“把 亚玛力 王 亚甲 带到我这里来。” 亚甲 就欢欢喜喜地来到他面前，说：“死亡的苦难必定过去了。”
1SAM|15|33|撒母耳 说：“你既用刀使妇人丧子，你母亲在妇人中也必照样丧子。”于是， 撒母耳 在 吉甲 耶和华面前把 亚甲 砍碎了。
1SAM|15|34|撒母耳 回了 拉玛 。 扫罗 上他所住的 基比亚 ，回自己的家去了。
1SAM|15|35|撒母耳 直到死的日子，再没有见 扫罗 。但 撒母耳 为 扫罗 悲伤，因为耶和华遗憾立 扫罗 为 以色列 的王。
1SAM|16|1|耶和华对 撒母耳 说：“我既厌弃 扫罗 作 以色列 的王，你为他悲伤要到几时呢？你将膏油盛满了角；来，我差遣你到 伯利恒 人 耶西 那里去，因为我在他儿子中已看中了一个为我作王的。”
1SAM|16|2|撒母耳 说：“我怎么能去呢？ 扫罗 一听见，就会杀我。”耶和华说：“你可以手里牵一头小母牛去，说：‘我来是要向耶和华献祭。’
1SAM|16|3|你要请 耶西 来一同献祭，我会指示你当做的事。我对你说的那个人，你要为我膏他。”
1SAM|16|4|撒母耳 遵照耶和华的话去做，来到 伯利恒 ，城里的长老都战战兢兢出来迎接他，有人问他说：“你是为平安来的吗？”
1SAM|16|5|他说：“为平安来的，我来是要向耶和华献祭。你们要使自己分别为圣，来跟我一同献祭。” 撒母耳 把 耶西 和他众儿子分别为圣，请他们来一同献祭。
1SAM|16|6|他们来的时候， 撒母耳 看见 以利押 ，就心里说，耶和华的受膏者一定在耶和华面前了。
1SAM|16|7|耶和华却对 撒母耳 说：“不要只看他的外貌和他身材高大，我不拣选他。因为耶和华不像人看人，人是看外貌 ，耶和华是看内心。”
1SAM|16|8|耶西 叫 亚比拿达 从 撒母耳 面前经过， 撒母耳 说：“耶和华也不拣选他。”
1SAM|16|9|耶西 又叫 沙玛 经过， 撒母耳 说：“耶和华也不拣选他。”
1SAM|16|10|耶西 叫他七个儿子都从 撒母耳 面前经过， 撒母耳 对 耶西 说：“这些都不是耶和华所拣选的。”
1SAM|16|11|撒母耳 对 耶西 说：“你的儿子都在这里了吗？”他说：“还有一个最小的，看哪，他正在放羊。” 撒母耳 对 耶西 说：“你派人去叫他来；他若不来这里，我们必不坐席。”
1SAM|16|12|耶西 就派人去叫他来。他面色红润，双目清秀，容貌俊美。耶和华说：“起来，膏他，因为这就是他了。”
1SAM|16|13|撒母耳 就用角里的膏油，在他的兄长中膏了他。从这日起，耶和华的灵就大大感动 大卫 。 撒母耳 起身回 拉玛 去了。
1SAM|16|14|耶和华的灵离开 扫罗 ，有邪灵从耶和华那里来扰乱他。
1SAM|16|15|扫罗 的臣仆对他说：“看哪，有邪灵从上帝那里来扰乱你。
1SAM|16|16|我们的主可以吩咐你面前的臣仆，去找一个善于弹琴的来。上帝那里来的邪灵临到你身上的时候，他用手弹琴，你就会感觉爽快。”
1SAM|16|17|扫罗 对臣仆说：“你们给我找一个善于弹琴的，带到我这里来。”
1SAM|16|18|仆人中有一个回答说：“看哪，我曾见 伯利恒 人 耶西 的一个儿子善于弹琴，是大能的勇士，说话合宜，容貌俊美，耶和华也与他同在。”
1SAM|16|19|于是 扫罗 差遣使者到 耶西 那里，说：“叫你放羊的儿子 大卫 到我这里来。”
1SAM|16|20|耶西 把几个饼和一皮袋酒，以及一只小山羊，驮在驴上，由儿子 大卫 的手送给 扫罗 。
1SAM|16|21|大卫 到了 扫罗 那里，就侍立在 扫罗 面前。 扫罗 很喜欢他，他就作了 扫罗 拿兵器的人。
1SAM|16|22|扫罗 派人到 耶西 那里，说：“让 大卫 侍立在我面前，因为他在我眼前蒙了恩宠。”
1SAM|16|23|从上帝那里来的邪灵临到 扫罗 身上的时候， 大卫 就拿琴，用手弹奏，使 扫罗 舒畅，感觉爽快，那邪灵就离开他了。
1SAM|17|1|非利士 人召集他们的军队来争战。他们聚集在 犹大 的 梭哥 ，在 梭哥 和 亚西加 中间的 以弗．大悯 安营。
1SAM|17|2|扫罗 和 以色列 人也聚集，在 以拉谷 安营，摆阵迎战，要与 非利士 人打仗。
1SAM|17|3|非利士 人站在这边的山上， 以色列 人站在那边的山上，当中有谷。
1SAM|17|4|从 非利士 营中出来一个挑战的人，名叫 歌利亚 ，是 迦特 人，身高六肘一虎口。
1SAM|17|5|他头戴铜盔，身穿铠甲，甲重五千舍客勒铜。
1SAM|17|6|他腿上有铜护膝，两肩之中背负铜矛。
1SAM|17|7|他的枪杆粗如织布机的轴，枪头的铁重六百舍客勒。有一个拿盾牌的人走在他前面。
1SAM|17|8|歌利亚 站着，对 以色列 的军队喊叫，对他们说：“你们出来摆阵作战是为了什么呢？我不是 非利士 人吗？你们不是 扫罗 的仆人吗？你们选一个人出来，叫他下来到我这里吧。
1SAM|17|9|他若能与我决斗，把我杀死，我们就作你们的奴隶；我若胜了他，把他杀死，你们就作我们的奴隶，服事我们。”
1SAM|17|10|那 非利士 人又说：“我今日向 以色列 的军队骂阵。你们叫一个人出来，跟我决斗吧。”
1SAM|17|11|扫罗 和 以色列 众人听见 非利士 人这些话就惊惶，非常害怕。
1SAM|17|12|大卫 是 犹大 伯利恒 的 以法他 人 耶西 的儿子， 耶西 有八个儿子。在 扫罗 的时候，这人年老，在众人中受敬重 。
1SAM|17|13|耶西 最大的三个儿子跟随 扫罗 出征。出征的三个儿子名字是：长子 以利押 ，次子 亚比拿达 ，三子 沙玛 。
1SAM|17|14|大卫 是最小的，最大的三个儿子跟随 扫罗 。
1SAM|17|15|大卫 有时离开 扫罗 ，回 伯利恒 为他父亲放羊。
1SAM|17|16|那 非利士 人早晚都出来站着，共四十日。
1SAM|17|17|耶西 对他儿子 大卫 说：“你拿一伊法烘了的穗子和十个饼，跑到营里去，交给你的哥哥，
1SAM|17|18|再拿这十块奶饼，送给他们的千夫长，并要问你哥哥好，向他们要个凭据回来。”
1SAM|17|19|扫罗 和 大卫 的三个哥哥，以及 以色列 众人，都在 以拉谷 与 非利士 人打仗。
1SAM|17|20|大卫 早晨起来，把羊交托一个看守的人，照 耶西 所吩咐的带着食物去了。到了军营，军队刚出到战场，呐喊叫阵。
1SAM|17|21|以色列 人和 非利士 人都摆列阵势，彼此相对。
1SAM|17|22|大卫 把东西留在看守物件的人手中，跑到战场，问他哥哥好。
1SAM|17|23|他与他们说话的时候，看哪，那挑战的人，就是 迦特 的 非利士 人 歌利亚 ，从 非利士 队伍中上来，说了同样的话， 大卫 听见了。
1SAM|17|24|以色列 众人看见那人就非常害怕，从他面前逃跑。
1SAM|17|25|以色列 人说：“这上来的人你看见了吗？他上来是要向 以色列 人骂阵。若有人能杀他，王必赏赐他大财，将自己的女儿嫁给他，并在 以色列 人中免除他父家纳粮服役。”
1SAM|17|26|大卫 对站在旁边的人说：“若有人杀这 非利士 人，除掉 以色列 人的羞辱，他会怎样呢？这未受割礼的 非利士 人是谁，竟敢向永生上帝的军队骂阵！”
1SAM|17|27|百姓照同样的话对他说：“若有人杀了那人，必这样待他。”
1SAM|17|28|大卫 的长兄 以利押 听见 大卫 与他们所说的话，就向他发怒，说：“你下来做什么呢？在旷野的那几只羊，你交托谁了呢？我知道你的骄傲和你心里的恶意，你下来只是为了看战争！”
1SAM|17|29|大卫 说：“我现在做了什么呢？只是问一句话也不可以吗？”
1SAM|17|30|大卫 离开他转向别人，问了同样的事，百姓也照先前的话回答他。
1SAM|17|31|有人听见 大卫 所说的话，就在 扫罗 面前报告； 扫罗 就派人叫他来。
1SAM|17|32|大卫 对 扫罗 说：“人不必因那 非利士 人灰心。你的仆人要去与他决斗。”
1SAM|17|33|扫罗 对 大卫 说：“你不能去与那 非利士 人决斗，因为你年纪太轻，他从小就是战士。”
1SAM|17|34|大卫 对 扫罗 说：“你仆人为父亲放羊，有时狮子来了，有时熊来了，从群中抓走一只羔羊。
1SAM|17|35|我就追赶它，击打它，把羔羊从它口中救出来。它起来攻击我，我就揪它的胡子，打死它。
1SAM|17|36|你仆人曾打死狮子和熊，这未受割礼的 非利士 人必像狮子和熊一样，因为他向永生上帝的军队骂阵。”
1SAM|17|37|大卫 又说：“耶和华救我脱离狮子和熊的爪，他必救我脱离这 非利士 人的手。” 扫罗 对 大卫 说：“你去吧！耶和华必与你同在。”
1SAM|17|38|扫罗 把自己的战衣给 大卫 穿上，将铜盔戴在他头上，又给他穿上铠甲。
1SAM|17|39|大卫 佩刀在战衣上，试着走走看。因 大卫 没有试过，就对 扫罗 说：“我穿戴这些不能走路，因为我没有试过。”于是他脱下身上的这些军装。
1SAM|17|40|他手中拿杖，又在溪中挑选了五块光滑的石子，放在袋里，就是牧人带的囊里，手里拿着甩石的机弦，迎向那 非利士 人。
1SAM|17|41|那 非利士 人渐渐走近 大卫 ，拿盾牌的人在他前面。
1SAM|17|42|非利士 人观看，见了 大卫 ，就藐视他，因为他年轻，面色红润，容貌俊美。
1SAM|17|43|非利士 人对 大卫 说：“你拿着杖到我这里来，我岂是狗吗？” 非利士 人就指着自己的神明诅咒 大卫 。
1SAM|17|44|非利士 人又对 大卫 说：“来吧！我要把你的肉给空中的飞鸟和田野的走兽。”
1SAM|17|45|大卫 对 非利士 人说：“你来攻击我，是靠着刀枪和铜矛，但我来攻击你，是靠着万军之耶和华的名，就是你所辱骂、带领 以色列 军队的上帝。
1SAM|17|46|今日耶和华必将你交在我手里。我必杀你，砍下你的头，今日我要把 非利士 军兵的尸体给空中的飞鸟和地上的野兽，使全地的人都知道以色列中有上帝，
1SAM|17|47|又使这里的全会众知道，耶和华使人得胜，不是用刀用枪，因为战争全在乎耶和华。他必将你们交在我们手里。”
1SAM|17|48|那 非利士 人起来，迎向 大卫 ，走近前来。 大卫 急忙往战场，迎向 非利士 人跑去。
1SAM|17|49|大卫 伸手入囊中，从里面掏出一块石子来，用机弦甩去，击中 非利士 人的前额，石子进入额内，他就仆倒，面伏于地。
1SAM|17|50|这样， 大卫 用机弦和石子胜了那 非利士 人，击中了他，把他杀死； 大卫 手中没有刀。
1SAM|17|51|大卫 跑去，站在那 非利士 人身旁，把他的刀从鞘中拔出来，杀死他，用刀割下他的头。 非利士 众人看见他们的勇士死了，就都逃跑。
1SAM|17|52|以色列 人和 犹大 人就起来呐喊，追赶 非利士 人，直到 该 和 以革伦 的城门。被杀的 非利士 人倒在路上，从 沙拉音 直到 迦特 和 以革伦 。
1SAM|17|53|以色列 人追赶 非利士 人回来，抢夺了他们的军营。
1SAM|17|54|大卫 拿着那 非利士 人的头带到 耶路撒冷 ，却把那 非利士 人的军装放在自己的帐棚里。
1SAM|17|55|扫罗 看见 大卫 去迎战 非利士 人，就问 押尼珥 元帅说：“ 押尼珥 ，那年轻人是谁的儿子？” 押尼珥 说：“王啊，我在你面前起誓，我不知道。”
1SAM|17|56|王说：“你可以问问那孩子是谁的儿子。”
1SAM|17|57|大卫 打死那 非利士 人回来， 押尼珥 领他到 扫罗 面前， 大卫 手中拿着 非利士 人的头。
1SAM|17|58|扫罗 问他说：“年轻人，你是谁的儿子？” 大卫 说：“我是你仆人 伯利恒 人 耶西 的儿子。”
1SAM|18|1|大卫 对 扫罗 说完了话， 约拿单 的心与 大卫 的心深相契合。 约拿单 爱 大卫 ，如同爱自己的性命。
1SAM|18|2|那日 扫罗 留住 大卫 ，不让他回父家。
1SAM|18|3|约拿单 爱 大卫 如同爱自己的性命，就与他立约。
1SAM|18|4|约拿单 从身上脱下外袍，给了 大卫 ，又把战衣、刀、弓、腰带都给了他。
1SAM|18|5|扫罗 无论差遣 大卫 往何处去，他都做事精明。 扫罗 立他作军队的指挥官，众百姓和 扫罗 的臣仆都看为美。
1SAM|18|6|大卫 打死了那 非利士 人，同众人回来的时候，妇女们从 以色列 各城里出来，欢欢喜喜，打鼓奏乐，唱歌跳舞，迎接 扫罗 王。
1SAM|18|7|众妇女欢乐唱和，说： “ 扫罗 杀死千千， 大卫 杀死万万。”
1SAM|18|8|扫罗 非常愤怒，不喜欢这话。他说：“将万万归给 大卫 ，千千归给我，只剩下王国没有给他！”
1SAM|18|9|从这日起， 扫罗 就敌视 大卫 。
1SAM|18|10|次日，从上帝来的邪灵紧抓住 扫罗 ，他就在家中胡言乱语。 大卫 照常弹琴， 扫罗 手里拿着枪。
1SAM|18|11|扫罗 把枪一掷，心里说：“我要将 大卫 刺透，钉在墙上。” 大卫 闪避了他两次。
1SAM|18|12|扫罗 惧怕 大卫 ，因为耶和华离开自己，与 大卫 同在。
1SAM|18|13|所以 扫罗 叫 大卫 离开自己，立他为千夫长，他就领兵出入。
1SAM|18|14|大卫 所做的每一件事都精明，耶和华也与他同在。
1SAM|18|15|扫罗 见 大卫 做事精明，就更怕他。
1SAM|18|16|但 以色列 和 犹大 众人都爱 大卫 ，因为他领他们出入。
1SAM|18|17|扫罗 对 大卫 说：“看哪，我将大女儿 米拉 嫁给你，只要你作我的勇士，为耶和华争战。” 扫罗 心里说：“我不好亲手害他，要藉 非利士 人的手害他。”
1SAM|18|18|大卫 对 扫罗 说：“我是谁，我是什么出身，我父家在 以色列 中算什么，岂敢作王的女婿呢？”
1SAM|18|19|扫罗 的女儿 米拉 到了当嫁给 大卫 的时候， 扫罗 却将她嫁给了 米何拉 人 亚得列 。
1SAM|18|20|扫罗 的女儿 米甲 爱 大卫 。有人告诉 扫罗 ，这件事在 扫罗 眼中看为合宜。
1SAM|18|21|扫罗 心里说：“我把这女儿嫁给 大卫 ，作他的圈套，好藉 非利士 人的手害他。”所以 扫罗 第二次对 大卫 说：“你今日可以作我的女婿。”
1SAM|18|22|扫罗 吩咐臣仆：“你们暗中对 大卫 说：‘看哪，王喜欢你，王的臣仆也都爱戴你，现在你就作王的女婿吧。’”
1SAM|18|23|扫罗 的臣仆照这话说给 大卫 听。 大卫 说：“你们把作王的女婿看为小事吗？我是贫穷卑微的人。”
1SAM|18|24|扫罗 的臣仆回奏说， 大卫 说了这样的话。
1SAM|18|25|扫罗 说：“你们要对 大卫 这样说：‘王不要什么聘礼，只要一百 非利士 人的包皮，好在王的仇敌身上报仇。’” 扫罗 的意图是要 大卫 落在 非利士 人的手中。
1SAM|18|26|扫罗 的臣仆把这话告诉 大卫 ， 大卫 就欢喜作王的女婿。日期还没有到，
1SAM|18|27|大卫 和跟随他的人起来前往，杀了二百 非利士 人，将包皮足数交给王，为要作王的女婿。于是 扫罗 将女儿 米甲 嫁给 大卫 。
1SAM|18|28|扫罗 见耶和华与 大卫 同在，女儿 米甲 又爱 大卫 ，
1SAM|18|29|就更怕 大卫 ，常常与 大卫 为敌。
1SAM|18|30|每逢 非利士 的军官出来打仗， 大卫 做事比 扫罗 任何臣仆更精明，因此他的名极受尊重。
1SAM|19|1|扫罗 吩咐他儿子 约拿单 和众臣仆要杀 大卫 ，但 扫罗 的儿子 约拿单 却很喜爱 大卫 。
1SAM|19|2|约拿单 告诉 大卫 说：“我父 扫罗 想要杀你，现在你要小心，明日早晨留在一个僻静的地方藏起来。
1SAM|19|3|我会出去，到你所藏的田里，站在我父亲旁边，与父亲谈论到你。我看情形怎样，会告诉你。”
1SAM|19|4|约拿单 向他父亲 扫罗 说 大卫 的好话，对他说：“王不可得罪王的仆人 大卫 ，因为他未曾得罪你，他所行的对你都很有益处。
1SAM|19|5|他拚了命杀那 非利士 人，并且耶和华为全 以色列 大施拯救。那时你看见，也很欢喜，现在为何要犯罪，流无辜人的血，无缘无故杀 大卫 呢？”
1SAM|19|6|扫罗 听了 约拿单 的话，就指着永生的耶和华起誓：“我绝不杀他。”
1SAM|19|7|约拿单 叫 大卫 来，把这一切事告诉他。 约拿单 带他去见 扫罗 ，他就像以前一样侍立在 扫罗 面前。
1SAM|19|8|此后又有战争， 大卫 出去与 非利士 人打仗。他大大击败他们，他们就在他面前逃跑。
1SAM|19|9|从耶和华来的邪灵又降在 扫罗 身上， 扫罗 手里拿枪坐在屋里， 大卫 正用手弹琴。
1SAM|19|10|扫罗 想要用枪刺透 大卫 ，把他钉在墙上，他却躲开 扫罗 ， 扫罗 的枪刺入墙内。当夜 大卫 逃走，躲起来了。
1SAM|19|11|扫罗 派一些使者到 大卫 的房屋那里守着他，等到天亮要杀他。 大卫 的妻子 米甲 对 大卫 说：“你今夜若不逃命，明日就要被杀。”
1SAM|19|12|于是 米甲 将 大卫 从窗户缒下去，让他走； 大卫 就逃走，躲起来了。
1SAM|19|13|米甲 把家中的神像放在床上，头枕在山羊毛的枕头上，用衣服盖起来。
1SAM|19|14|扫罗 派一些使者去捉拿 大卫 ， 米甲 说：“他病了。”
1SAM|19|15|扫罗 又派一些使者去看 大卫 ，说：“把他连床一起抬到我这里，我好杀他。”
1SAM|19|16|使者进去，看哪，神像在床上，头枕在山羊毛的枕头上。
1SAM|19|17|扫罗 对 米甲 说：“你为什么这样欺骗我，放我仇敌逃走呢？” 米甲 对 扫罗 说：“他对我说：‘你放我走吧，我何必要杀你呢？’”
1SAM|19|18|大卫 逃跑躲避，来到 拉玛 的 撒母耳 那里，把 扫罗 向他所行的事全告诉他。他和 撒母耳 就去，住在 拿约 。
1SAM|19|19|有人告诉 扫罗 说：“看哪， 大卫 在 拉玛 的 拿约 ”。
1SAM|19|20|扫罗 派一些使者去捉拿 大卫 。去的人见一队先知受感说话， 撒母耳 站在当中领导他们， 扫罗 派去的使者也受上帝的灵感动说话。
1SAM|19|21|有人把这事告诉 扫罗 ，他又派另一些使者去，他们也受感说话。 扫罗 第三次派使者去，他们也受感说话。
1SAM|19|22|然后 扫罗 亲自往 拉玛 去，到了 西沽 的大井，问人说：“ 撒母耳 和 大卫 在哪里？”有人说：“看哪，在 拉玛 的 拿约 。”
1SAM|19|23|他就往那里去，到了 拉玛 的 拿约 。上帝的灵也临到他，他一面走一面受感说话，直到 拉玛 的 拿约 。
1SAM|19|24|他也脱了衣服，也在 撒母耳 面前受感说话，一日一夜赤身躺卧。因此有人说：“ 扫罗 也在先知中吗？”
1SAM|20|1|大卫 从 拉玛 的 拿约 逃跑，来到 约拿单 面前，对他说：“我做了什么，有什么罪孽，在你父亲面前犯了什么罪，他竟要寻索我的性命呢？”
1SAM|20|2|约拿单 对他说：“绝无此事！你必不至于死。看哪，我父做事，无论大小，没有不告诉我的。我父亲为什么要隐瞒我这件事呢？不会这样的！”
1SAM|20|3|大卫 又起誓说：“你父亲确实知道我在你眼前蒙恩。所以他说，‘这事不要让 约拿单 知道，免得他愁烦。’我指着永生的耶和华起誓，又指着你的性命起誓，我离死只差一步而已。”
1SAM|20|4|约拿单 对 大卫 说：“你心里所求的，我必为你成就。”
1SAM|20|5|大卫 对 约拿单 说：“看哪，明日是初一，我必须与王同席用餐，求你让我去藏在田野，直到第三日傍晚。
1SAM|20|6|你父亲若见我不在席上，你就说：‘ 大卫 恳求我允许他赶回本城 伯利恒 去，因为他全家在那里献年祭。’
1SAM|20|7|你父亲若说好，你的仆人就平安了；他若大怒，你就知道他决意行恶。
1SAM|20|8|求你施恩于仆人，因你在耶和华面前曾与仆人立约。我若有罪孽，你就亲自杀死我，何必把我交给你父亲呢？”
1SAM|20|9|约拿单 说：“绝无此事！我若确实知道我父亲决意害你，怎么会不告诉你呢？”
1SAM|20|10|大卫 对 约拿单 说：“你父亲若严厉回答你，谁来告诉我呢？”
1SAM|20|11|约拿单 对 大卫 说：“来，让我们到田野去。”二人就往田野去了。
1SAM|20|12|约拿单 对 大卫 说：“愿耶和华－ 以色列 的上帝作证。明日约在这时候，或第三日，我一探出我父亲的心意，看哪，若对 大卫 是好意，我怎么会不派人来告诉你呢？
1SAM|20|13|我父亲若有意害你，而我不告诉你，送你平安地离开，愿耶和华重重惩罚 约拿单 。愿耶和华与你同在，如同从前与我父亲同在一样。
1SAM|20|14|你要照耶和华的慈爱恩待我，不但我活着的时候免我死亡，
1SAM|20|15|就是耶和华从地面逐一剪除 大卫 仇敌的时候，你也永不可向我家断绝恩惠。”
1SAM|20|16|于是 约拿单 与 大卫 家立约：“愿耶和华从 大卫 仇敌 的手来追讨。”
1SAM|20|17|约拿单 因爱 大卫 如同爱自己的性命，就叫他再起誓。
1SAM|20|18|约拿单 对他说：“明日是初一，你的座位空着，人必察觉你不在。
1SAM|20|19|到第三日，就要走一段长路下去 ，去到你遇事那天所藏的地方，在 以色 磐石 的旁边等候。
1SAM|20|20|我会向磐石旁边射三箭，如同射箭靶一样。
1SAM|20|21|看哪，我会派僮仆，说：‘去把箭找来。’我若对僮仆喊说：‘看哪，箭在你的这边，把箭拿来’，你就可以平安回来；我指着永生的耶和华起誓，你一定没有事。
1SAM|20|22|我若对孩子说：‘看哪，箭在你的前方’，你就要离开，因为是耶和华差你去的。
1SAM|20|23|至于你和我，我们所说的话，看哪，耶和华在你我中间作证，直到永远。”
1SAM|20|24|大卫 就去藏在田野。到了初一，王要坐席用餐。
1SAM|20|25|王照常坐在靠墙的位子上， 约拿单 在对面 ， 押尼珥 坐在 扫罗 旁边， 大卫 的座位却是空的。
1SAM|20|26|这日 扫罗 没有说什么，因为他说：“ 大卫 或许有事，偶染不洁，还未得洁净。”
1SAM|20|27|初二， 大卫 的座位还空着。 扫罗 对他儿子 约拿单 说：“ 耶西 的儿子为何昨日、今日都没有来用餐呢？”
1SAM|20|28|约拿单 回答 扫罗 说：“ 大卫 恳求我允许他回 伯利恒 去，
1SAM|20|29|说：‘求你让我去，因为我家在城里有献祭的事，我哥哥吩咐我去。如今我若在你眼前蒙恩，求你让我去见我的兄弟。’所以 大卫 没有来赴王的筵席。”
1SAM|20|30|扫罗 向 约拿单 怒气大发，对他说：“你这顽梗悖逆之妇人所生的，我怎么会不知道你选择 耶西 的儿子 ，自取羞辱，也使你母亲露体蒙羞呢？
1SAM|20|31|只要 耶西 的儿子还活在世上一天，你和你的国必保不住。现在你要派人去，把他带到我这里来，因为他是该死的。”
1SAM|20|32|约拿单 回答父亲 扫罗 说：“他为什么该死呢？他做了什么呢？”
1SAM|20|33|扫罗 向 约拿单 掷枪要刺他， 约拿单 就知道他父亲决意要杀死 大卫 。
1SAM|20|34|于是 约拿单 气愤愤地从席上起来。他在初二这天没有吃饭，因为他为 大卫 愁烦，又因为他父亲羞辱了他。
1SAM|20|35|次日早晨， 约拿单 按着与 大卫 约定的时候到田野去，有一个小僮仆跟随他。
1SAM|20|36|约拿单 对僮仆说：“你跑去把我所射的箭找来。”僮仆跑去， 约拿单 就把箭射在僮仆的前方。
1SAM|20|37|僮仆到了 约拿单 落箭之地， 约拿单 呼叫僮仆说：“箭不是在你的前方吗？”
1SAM|20|38|约拿单 又呼叫僮仆说：“快去，不要站在那里！”僮仆就捡起箭来，回到主人那里。
1SAM|20|39|僮仆不知道这是什么意思，只有 约拿单 和 大卫 知道这事。
1SAM|20|40|约拿单 把他的弓箭交给僮仆，吩咐他说：“你拿到城里去。”
1SAM|20|41|僮仆一去， 大卫 就从南边 出来，俯伏在地，拜了三拜。他们彼此亲吻，一起哭泣， 大卫 哭得更悲哀。
1SAM|20|42|约拿单 对 大卫 说：“你平平安安地去吧！因为我们二人曾指着耶和华的名起誓说：‘愿耶和华在你我中间，以及你我后裔中间作证，直到永远。’” 大卫 就起身走了， 约拿单 也回城里去了。
1SAM|21|1|大卫 到了 挪伯 的 亚希米勒 祭司那里， 亚希米勒 战战兢兢地出来迎接他，对他说：“你为什么独自一人，没有人跟随你呢？”
1SAM|21|2|大卫 对 亚希米勒 祭司说：“王吩咐我一件事，对我说：‘我差遣你，吩咐你的这件事，不可让任何人知道。’因此我已告诉一些仆人到某处去 。
1SAM|21|3|现在你手中有什么？请你给我五个饼或是可以找到的食物。”
1SAM|21|4|祭司对 大卫 说：“我手中没有普通的饼，只有圣饼，只能给没有亲近妇人的年轻人。”
1SAM|21|5|大卫 回答祭司说：“我们确实没有亲近妇人，如同往常我出征的时候一样。平常行路，仆人的身体 都还分别为圣，何况今日岂不更使自己分别为圣吗？”
1SAM|21|6|祭司拿圣饼给他，因为在那里没有别的饼，只有那从耶和华面前撤下的供饼，就是换上热饼的日子取下来的。
1SAM|21|7|当日，有 扫罗 的一个臣仆在那里，他留在耶和华的面前，名叫 多益 ，是 以东 人，作 扫罗 的畜牧长。
1SAM|21|8|大卫 对 亚希米勒 说：“你手中有没有枪或刀？因为王的事紧急，连刀剑兵器我都没有带。”
1SAM|21|9|祭司说：“你在 以拉谷 所杀的 非利士 人 歌利亚 的那刀，看哪，裹在布中，放在以弗得后边。你若要可以拿去，除此以外，再没有别的了。” 大卫 说：“没有什么可以跟它比的了！请你给我。”
1SAM|21|10|那日 大卫 起来，躲避 扫罗 ，逃到 迦特 王 亚吉 那里。
1SAM|21|11|亚吉 的臣仆对他说：“这不是那地的国王 大卫 吗？那里的人跳舞唱和： ‘ 扫罗 杀死千千， 大卫 杀死万万’， 不是指着他说的吗？”
1SAM|21|12|大卫 把这些话放在心里，就很惧怕 迦特 王 亚吉 。
1SAM|21|13|于是他在众人眼前一反常态，在他们中间 装疯作癫，在城门的门扇上胡写乱画，任由唾沫流在胡子上。
1SAM|21|14|亚吉 对臣仆说：“看哪，你们看这人疯了，为什么带他到我这里来呢？
1SAM|21|15|我岂缺少疯子，你们竟然带这人到我面前疯癫吗？这个人可以进我的家吗？”
1SAM|22|1|大卫 离开那里，逃到 亚杜兰 洞。他的兄弟和他父亲全家听见了，都下到他那里去。
1SAM|22|2|凡生活窘迫的、欠债的、心里苦恼的都聚集到 大卫 那里，他就作他们的领袖，跟随他的约有四百人。
1SAM|22|3|大卫 从那里往 摩押 的 米斯巴 去，对 摩押 王说：“请你让我父母搬来，跟你们在一起，等我知道上帝要为我怎样做。”
1SAM|22|4|大卫 领他父母到 摩押 王面前。 大卫 住山寨一切的日子，他父母也都住在 摩押 王那里。
1SAM|22|5|先知 迦得 对 大卫 说：“你不要住在山寨，要到 犹大 地去。” 大卫 就去，来到 哈列 的树林。
1SAM|22|6|扫罗 听见 大卫 和跟随他之人的下落， 扫罗 正在 基比亚 ，坐在山顶 的柳树下，手里拿着枪，众臣仆侍立在左右。
1SAM|22|7|扫罗 对左右侍立的臣仆说：“ 便雅悯 人哪，听着！ 耶西 的儿子也能把田地和葡萄园赐给你们各人吗？他能立你们各人作千夫长和百夫长吗？
1SAM|22|8|你们竟都结党害我！我儿子与 耶西 的儿子立约的时候，无人告诉我；我儿子挑唆我的臣仆谋害我，像今日这样，也无人告诉我，为我忧虑。”
1SAM|22|9|那时 以东 人 多益 站在 扫罗 的臣仆中，回答说：“我曾看见 耶西 的儿子往 挪伯 去，到了 亚希突 的儿子 亚希米勒 那里。
1SAM|22|10|亚希米勒 为他求问耶和华，给他食物，又把 非利士 人 歌利亚 的刀给了他。”
1SAM|22|11|王就派人把 亚希突 的儿子 亚希米勒 祭司和他父亲的全家，就是在 挪伯 的祭司都召了来，他们都来到王那里。
1SAM|22|12|扫罗 说：“ 亚希突 的儿子，听着！”他说：“我主，我在这里。”
1SAM|22|13|扫罗 对他说：“你为什么与 耶西 的儿子结党害我，把食物和刀给他，又为他求问上帝，使他起来谋害我，像今日这样？”
1SAM|22|14|亚希米勒 回答王说：“王的众臣仆中有谁比 大卫 忠心呢？他是王的女婿，又是你的侍卫长 ，并且是你宫中受敬重的人。
1SAM|22|15|我今日才开始为他求问上帝吗？绝非如此！王不要归罪于我和我父全家，因为这事，无论大小，仆人都不知情。”
1SAM|22|16|王说：“ 亚希米勒 ，你和你父全家都是该死的！”
1SAM|22|17|王吩咐左右的侍卫说：“你们转身去杀耶和华的祭司吧！因为他们帮助 大卫 ，知道 大卫 逃跑却不告诉我。”但王的臣仆都不愿动手杀耶和华的祭司。
1SAM|22|18|王吩咐 多益 说：“你转身去杀祭司吧！” 以东 人 多益 就转身去杀祭司，那日杀了穿细麻布以弗得的，共八十五人，
1SAM|22|19|又用刀把祭司城 挪伯 中的男女、孩童和吃奶的都杀了，又用刀杀了牛、羊和驴子。
1SAM|22|20|亚希突 的儿子 亚希米勒 有一个儿子逃脱了；他名叫 亚比亚他 ，逃到 大卫 那里。
1SAM|22|21|亚比亚他 把 扫罗 杀耶和华祭司的事告诉 大卫 。
1SAM|22|22|大卫 对 亚比亚他 说：“那日我见 以东 人 多益 在那里，就知道他一定会告诉 扫罗 。你父的全家丧命，都是因我的缘故。
1SAM|22|23|你可以住在我这里，不要惧怕。因为寻索你命的也要寻索我的命，你在我这里可得保护。”
1SAM|23|1|有人告诉 大卫 说：“看哪， 非利士 人攻击 基伊拉 ，抢夺禾场。”
1SAM|23|2|大卫 求问耶和华说：“我可以去吗？我可以去攻打那些 非利士 人吗？”耶和华对 大卫 说：“你可以去攻打 非利士 人，拯救 基伊拉 。”
1SAM|23|3|大卫 的人对他说：“看哪，我们在 犹大 这里尚且惧怕，何况到 基伊拉 去攻打 非利士 人的军队呢？”
1SAM|23|4|大卫 又再求问耶和华，耶和华回答说：“你起身下 基伊拉 去，我必将 非利士 人交在你手里。”
1SAM|23|5|于是 大卫 和他的人往 基伊拉 去，与 非利士 人打仗，大大击败他们，夺取他们的牲畜。这样， 大卫 救了 基伊拉 的居民。
1SAM|23|6|亚希米勒 的儿子 亚比亚他 逃往 基伊拉 到 大卫 那里的时候，手里拿着以弗得。
1SAM|23|7|有人告诉 扫罗 ， 大卫 到了 基伊拉 。 扫罗 说：“上帝将他交在我手里了，因为他进了有门有闩的城，把自己关起来了。”
1SAM|23|8|于是 扫罗 召集众百姓，要下去攻打 基伊拉 ，围困 大卫 和他的人。
1SAM|23|9|大卫 知道 扫罗 设计陷害他，就对 亚比亚他 祭司说：“把以弗得拿过来。”
1SAM|23|10|大卫 说：“耶和华－ 以色列 的上帝啊，你仆人确实听见 扫罗 设法要到 基伊拉 来，为我的缘故毁灭这城。
1SAM|23|11|基伊拉 人会把我交在 扫罗 手里吗？ 扫罗 会下来，正如你仆人所听见的吗？耶和华－ 以色列 的上帝啊，求你指示仆人！”耶和华说：“他会下来。”
1SAM|23|12|大卫 又说：“ 基伊拉 人会把我和我的人交在 扫罗 手里吗？”耶和华说：“他们会交出来。”
1SAM|23|13|于是 大卫 和他的人约有六百名起身离开 基伊拉 ，往他们所能去的地方去。有人告诉 扫罗 ， 大卫 离开 基伊拉 逃走了， 扫罗 就停止出发了。
1SAM|23|14|大卫 住在旷野的山寨里，在 西弗 旷野的山区。 扫罗 天天寻索 大卫 ，上帝却不将 大卫 交在他手里。
1SAM|23|15|大卫 看到 扫罗 出来寻索他的命。那时，他住在 西弗 旷野的树林里 ；
1SAM|23|16|扫罗 的儿子 约拿单 起身，到树林里去见 大卫 ，使他的手倚靠上帝得以坚固，
1SAM|23|17|对他说：“不要惧怕！我父 扫罗 的手无法害你 ，你必作 以色列 的王，我必作你的宰相。我父 扫罗 也知道这事。”
1SAM|23|18|于是二人在耶和华面前立约。 大卫 仍住在树林里， 约拿单 就回家去了。
1SAM|23|19|西弗 人上 基比亚 到 扫罗 那里，说：“ 大卫 不是在我们那里，在树林里的山寨中，在荒野 南边的 哈基拉山 藏着吗？
1SAM|23|20|现在，王啊，请随你的心愿要下来，就请下来；至于我们，一定会把他交在王的手里。”
1SAM|23|21|扫罗 说：“愿耶和华赐福给你们，因为你们体恤我。
1SAM|23|22|请你们回去，再确定一下，调查并看清楚他落脚的地方，是谁看见他在那里 ，因为有人告诉我他很狡猾。
1SAM|23|23|你们要看清楚，调查他藏匿的每一个地方，回来给我确实的报告，我就与你们同去。他若在境内，我必从 犹大 的千门万户中搜出他来。”
1SAM|23|24|西弗 人动身，在 扫罗 以先往 西弗 去。 大卫 和他的人却在 玛云 旷野，在荒野南边的 亚拉巴 。
1SAM|23|25|扫罗 和他的人去寻索 大卫 。有人告诉 大卫 ，他就下到岩石那里，留在 玛云 的旷野。 扫罗 听见了，就在 玛云 的旷野追赶 大卫 。
1SAM|23|26|扫罗 在山的这一边走， 大卫 和他的人在山的那一边。 大卫 急忙躲避 扫罗 ， 扫罗 和他的人正四面围住 大卫 和他的人，要捉拿他们。
1SAM|23|27|有使者来对 扫罗 说：“ 非利士 人入境抢掠，请快快回去！”
1SAM|23|28|于是 扫罗 不再追赶 大卫 ，回去迎击 非利士 人。因此那地方名叫 西拉．哈玛希罗结 。
1SAM|23|29|大卫 从那里上去，住在 隐．基底 的山寨里。
1SAM|24|1|扫罗 追赶 非利士 人回来，有人告诉他说：“看哪， 大卫 在 隐．基底 的旷野。”
1SAM|24|2|扫罗 就从全 以色列 中挑选三千精兵，往 野山羊磐石 的东边 去，寻索 大卫 和他的人。
1SAM|24|3|到了路旁的羊圈，在那里有个洞， 扫罗 进去大解。 大卫 和他的人正藏在洞里的深处。
1SAM|24|4|大卫 的人对 大卫 说：“看哪，这日子到了！耶和华曾对你说：‘看哪，我要将你的仇敌交在你手里，你可以照你看为好的对待他。’” 大卫 就起来，悄悄地割下 扫罗 外袍的衣角。
1SAM|24|5|随后 大卫 心中自责，因为他割下了 扫罗 的衣角。
1SAM|24|6|他对他的人说：“耶和华绝不允许我对我的主，耶和华的受膏者做这事，伸手害他，因为他是耶和华的受膏者。”
1SAM|24|7|大卫 用这话劝阻他的人，不许他们起来害 扫罗 。 扫罗 起来，从洞里出去，预备上路。
1SAM|24|8|然后 大卫 也起来，从洞里出去，呼唤 扫罗 说：“我主，我王！” 扫罗 回头观看， 大卫 就屈身，脸伏于地下拜。
1SAM|24|9|大卫 对 扫罗 说：“你为何听信人的谗言，说‘看哪， 大卫 想要害你’呢？
1SAM|24|10|看哪，今日你亲眼看见，在洞中耶和华将你交在我手里。有人要我杀你，我却爱惜你，说：‘我不敢伸手害我的主，因为他是耶和华的受膏者。’
1SAM|24|11|我父啊，请看，看你外袍的衣角在我手中。我割下你外袍的衣角，却没有杀你。你知道，并且看见我没有恶意要悖逆你。你虽然要猎取我的命，我却没有得罪你。
1SAM|24|12|愿耶和华在你我中间判断，愿耶和华在你身上为我伸冤，我却不亲手加害于你。
1SAM|24|13|古人有句俗语说：‘恶事出于恶人。’我却不亲手加害于你。
1SAM|24|14|以色列 王出来要寻找谁呢？你要追赶谁呢？不过是一条死狗，一只跳蚤而已。
1SAM|24|15|愿耶和华作仲裁者，在你我中间判断。愿他鉴察，为我伸冤，救我脱离你的手。”
1SAM|24|16|大卫 向 扫罗 说完了这些话， 扫罗 说：“我儿 大卫 ，这是你的声音吗？”于是 扫罗 放声大哭，
1SAM|24|17|对 大卫 说：“你比我公义，因为你以善待我，我却以恶待你。
1SAM|24|18|今日你已显明是以善待我，因为耶和华将我交在你手里，你却没有杀我。
1SAM|24|19|人若遇见仇敌，岂肯放他平安上路呢？愿耶和华因你今日向我所做的，以善回报你。
1SAM|24|20|现在，看哪，我知道你一定会作王， 以色列 的国必要坚立在你手里。
1SAM|24|21|现在你要指着耶和华向我起誓，你必不剪除我的后裔，必不从我父家除去我的名。”
1SAM|24|22|于是 大卫 向 扫罗 起誓， 扫罗 就回家去， 大卫 和他的人也上山寨去了。
1SAM|25|1|撒母耳 死了， 以色列 众人聚集，为他哀哭，把他葬在 拉玛 他的家里。 大卫 动身，下到 巴兰 的旷野。
1SAM|25|2|在 玛云 有一个人，他的产业在 迦密 。这人是一个大富翁，有三千只绵羊，一千只山羊；他正在 迦密 剪羊毛。
1SAM|25|3|这人名叫 拿八 ，他的妻子名叫 亚比该 。 拿八 的妻子有美好的见识，又有美丽的容貌，但 拿八 为人刚愎凶恶，是 迦勒 族的人。
1SAM|25|4|大卫 在旷野听见 拿八 正在剪羊毛，
1SAM|25|5|就派十个仆人，对他们说：“你们上 迦密 到 拿八 那里，提我的名向他问安。
1SAM|25|6|你们要如此说：‘愿你来年平安 ，愿你家平安，愿你一切所有的都平安。
1SAM|25|7|现在我听说你有剪羊毛的人，你的牧人和我们在一起，他们在 迦密 一切的日子，我们没有欺负过他们，他们也未曾失去什么。
1SAM|25|8|你问你的仆人，他们会告诉你。愿我的仆人在你眼前得欢心，因为我们是在好日子来的。请你随手分点食物给仆人和你儿子 大卫 。’”
1SAM|25|9|大卫 的仆人到了，就提 大卫 的名，把这一切话告诉 拿八 ，他们就停顿下来。
1SAM|25|10|拿八 回答 大卫 的仆人说：“ 大卫 是谁？ 耶西 的儿子是谁？今日悖逆主人奔逃的仆人很多。
1SAM|25|11|我岂可把饮食，以及我为剪羊毛的人所宰的肉给那些我不知道从哪里来的人呢？”
1SAM|25|12|大卫 的仆人转身从原路回去，照这一切的话告诉 大卫 。
1SAM|25|13|大卫 对他的人说：“你们各人都要佩上刀！”各人就都佩上刀， 大卫 也佩上刀。跟随 大卫 上去的约有四百人，留下二百人看守物件。
1SAM|25|14|拿八 的一个仆人告诉 拿八 的妻子 亚比该 说：“看哪， 大卫 从旷野派使者来向我主人问安，主人却辱骂他们。
1SAM|25|15|但是那些人待我们真好；我们在田野与他们一切来往的日子，没有受他们欺负，也未曾失去什么。
1SAM|25|16|我们在他们那里牧羊，一切的日子他们昼夜保护我们 。
1SAM|25|17|现在，你当知道，看怎样做才好。不然，祸患必定临到我主人和他全家。他性情凶暴，无人敢与他说话。”
1SAM|25|18|亚比该 急忙将二百个饼，两皮袋酒，五只宰好的羊，五细亚烘熟的穗子，一百个葡萄干饼，二百个无花果饼，都驮在驴上，
1SAM|25|19|对仆人说：“你们在我前面走，看哪，我跟着你们去。”她却没有告诉丈夫 拿八 。
1SAM|25|20|亚比该 骑着驴，正下山坡，看哪， 大卫 和他的人正迎着 亚比该 下来，她就去迎接他们。
1SAM|25|21|大卫 曾说：“我在旷野为那人看守他一切所有的，以致他未失去任何一样东西，实在是徒然了！他竟然向我以恶报善。
1SAM|25|22|凡属 拿八 的男丁，我若留一个到明日早晨，愿上帝重重惩罚 大卫 ！”
1SAM|25|23|亚比该 看见 大卫 ，就急忙下驴，在 大卫 面前脸伏于地叩拜。
1SAM|25|24|她俯伏在 大卫 的脚前，说：“我主啊，愿这罪归于我！求你容许使女向你进言，更求你听使女的话。
1SAM|25|25|我主不必理会 拿八 这性情凶暴的人，他就像他的名字一样；他名叫 拿八 ，为人也真是愚顽。至于我，你的使女并没有看见我主所派来的仆人。
1SAM|25|26|现在，我主啊，耶和华既然阻止你亲手报仇，避免流人的血，我指着永生的耶和华起誓，又指着你的性命起誓：‘现在，愿你的仇敌和谋害我主的人都像 拿八 一样。’
1SAM|25|27|现在求我主把婢女送来的礼物给跟随我主的仆人。
1SAM|25|28|求你原谅使女的冒犯。耶和华必为我主建立坚固的家，因为我主为耶和华争战，并且你一生的日子查不出有什么恶来。
1SAM|25|29|虽有人起来追逼你，要寻索你的性命，我主的性命在耶和华－你的上帝那里，如同藏在生命的宝藏中。至于你仇敌的性命，耶和华必甩去，如用机弦甩石一样。
1SAM|25|30|耶和华照所应许你的福气赐给我主，立你作 以色列 王的时候，
1SAM|25|31|我主就不至于因为亲手报仇，流了无辜人的血，而心里不安，良心有亏了。耶和华赐福给我主的时候，求你记得你的使女。”
1SAM|25|32|大卫 对 亚比该 说：“耶和华－ 以色列 的上帝是应当称颂的，因为他今日派你来迎接我。
1SAM|25|33|你和你的见识也配得称赞，因为你今日拦阻我亲手报仇、流人的血。
1SAM|25|34|我指着阻止我加害于你的耶和华－ 以色列 永生的上帝起誓，若不是你很快地来迎接我，到早晨天亮的时候，凡属 拿八 的男丁，必定一个也不留。”
1SAM|25|35|大卫 从 亚比该 手中收了她带来的礼物，对她说：“平平安安上你的家去吧！你看，我看了你的情面，听了你的话。”
1SAM|25|36|亚比该 到 拿八 那里，看哪，他在家里摆设宴席，如同王的宴席。 拿八 心情舒畅，酩酊大醉。所以 亚比该 大小事都没有告诉他，直等到早晨天亮的时候。
1SAM|25|37|到了早晨， 拿八 酒醒了，他的妻子把这些事都告诉他，他就发心脏病快死了，僵如石头。
1SAM|25|38|过了十天，耶和华击打 拿八 ，他就死了。
1SAM|25|39|大卫 听见 拿八 死了，就说：“耶和华是应当称颂的，因为我从 拿八 手中受了羞辱，他为我伸冤，又阻止他的仆人行恶；耶和华使 拿八 的恶归到他自己头上。”于是 大卫 派人去向 亚比该 说，要娶她为妻。
1SAM|25|40|大卫 的仆人来到 迦密 ，到 亚比该 那里，对她说：“ 大卫 派我们到你这里，要娶你作他的妻子。”
1SAM|25|41|亚比该 起来叩拜，俯伏在地，说：“看哪，你的使女情愿作婢女，为我主的仆人洗脚。”
1SAM|25|42|亚比该 立刻起身，骑上驴，五个女仆跟着她走。她跟从 大卫 的使者去，就作了 大卫 的妻子。
1SAM|25|43|大卫 先前娶了 耶斯列 人 亚希暖 ，她们二人都作了他的妻子。
1SAM|25|44|扫罗 已把他的女儿 米甲 ，就是 大卫 的妻子，给了 迦琳 人 拉亿 的儿子 帕提 为妻。
1SAM|26|1|西弗 人来到 基比亚 ，到 扫罗 那里，说：“ 大卫 不是在荒野 东边 的 哈基拉山 藏着吗？”
1SAM|26|2|扫罗 动身，带领 以色列 人中挑选的三千精兵下到 西弗 的旷野，要在那里寻索 大卫 。
1SAM|26|3|扫罗 在荒野东边的 哈基拉山 ，在路旁安营。那时 大卫 住在旷野，看见 扫罗 到旷野来追赶他，
1SAM|26|4|大卫 就派人去探听，知道 扫罗 果然来了。
1SAM|26|5|大卫 起来，到 扫罗 安营的地方，看见 扫罗 和 尼珥 的儿子 押尼珥 元帅躺卧之处； 扫罗 睡在军营里，士兵安营在他周围。
1SAM|26|6|大卫 对 赫 人 亚希米勒 和 洗鲁雅 的儿子 约押 的兄弟 亚比筛 说：“谁同我下到 扫罗 营里去？” 亚比筛 说：“我同你下去。”
1SAM|26|7|于是 大卫 和 亚比筛 夜间到了士兵那里；看哪， 扫罗 睡在军营里，他的枪在头旁，插在地上。 押尼珥 和士兵睡在他周围。
1SAM|26|8|亚比筛 对 大卫 说：“上帝将你的仇敌交在你手里，现在让我拿枪把他刺透在地上，一刺就成，不用再刺他了。”
1SAM|26|9|大卫 对 亚比筛 说：“不可杀害他！有谁伸手害耶和华的受膏者而无罪呢？”
1SAM|26|10|大卫 又说：“我指着永生的耶和华起誓，他或被耶和华击杀，或死期到了，或出战阵亡，
1SAM|26|11|耶和华绝不允许我伸手害耶和华的受膏者。现在你可以把他头旁的枪和水壶拿来，我们就走。”
1SAM|26|12|大卫 从 扫罗 的头旁拿了枪和水壶，他们就走了。没有人看见，没有人知道，也没有人醒过来。他们都睡着了，因为耶和华使他们沉睡了。
1SAM|26|13|大卫 过到另一边去，远远地站在山顶上，与他们相离很远。
1SAM|26|14|大卫 呼叫百姓和 尼珥 的儿子 押尼珥 说：“ 押尼珥 ，你为何不回答呢？” 押尼珥 回答说：“你是谁？竟敢呼唤王呢？”
1SAM|26|15|大卫 对 押尼珥 说：“你不是个大丈夫吗？ 以色列 中谁能比你呢？百姓中有一个人进来要害死你主你王，你为何没有保护你主你王呢？
1SAM|26|16|你做的这件事不好！我指着永生的耶和华起誓，你们都是该死的，因为你们没有保护你们的主，就是耶和华的受膏者。现在你看，王头旁的枪和水壶在哪里？”
1SAM|26|17|扫罗 认出 大卫 的声音，就说：“我儿 大卫 ，这是你的声音吗？” 大卫 说：“我主我王啊，是我的声音。”
1SAM|26|18|又说：“我主为何要追赶仆人呢？我做了什么？我手做了什么恶事呢？
1SAM|26|19|现在求我主我王听仆人的话：若是耶和华激发你来攻击我，愿耶和华悦纳供物；若是出于人，愿他们在耶和华面前受诅咒，因为他们今日赶逐我，不让我在耶和华的产业中有分，说：‘你去事奉别神吧！’
1SAM|26|20|现在不要使我的血流在远离耶和华面的地上。因为 以色列 王出来，只不过是寻找一只跳蚤，如同人在山上猎取一只鹧鸪。”
1SAM|26|21|扫罗 说：“我有罪了！我儿 大卫 ，回来吧！我必不再加害于你，因为你今日看我的性命为宝贵。看哪，我是个糊涂人，大大错了。”
1SAM|26|22|大卫 回答说：“看哪，这是王的枪，可以吩咐一个仆人过来拿去。
1SAM|26|23|今日耶和华将王交在我手里，我却不肯伸手害耶和华的受膏者。耶和华必照各人的公义诚实报应他。
1SAM|26|24|看哪，我今日看重你的性命，愿耶和华也照样看重我的性命，并且拯救我脱离一切患难。”
1SAM|26|25|扫罗 对 大卫 说：“我儿 大卫 ，愿你得福！你必做大事，也必得胜。”于是 大卫 上路， 扫罗 也回自己的地方去了。
1SAM|27|1|大卫 心里说：“总有一天我会死在 扫罗 手里，现在我最好逃到 非利士 人的地去， 扫罗 就会绝望，不会继续在 以色列 全境内寻索我了。这样，我才可以脱离他的手。”
1SAM|27|2|于是 大卫 动身，和跟随他的六百人投奔 玛俄 的儿子 迦特 王 亚吉 去了。
1SAM|27|3|大卫 和他的两个妻子，就是 耶斯列 人 亚希暖 和作过 拿八 妻子的 迦密 人 亚比该 ，以及他的人，连同各人的眷属，都住在 迦特 的 亚吉 那里。
1SAM|27|4|有人告诉 扫罗 ：“ 大卫 逃到 迦特 。” 扫罗 就不再寻索他了。
1SAM|27|5|大卫 对 亚吉 说：“我若蒙你看得起，求你在郊外的城镇中赐我一个地方，让我住在那里。仆人何必与王同住京城呢？”
1SAM|27|6|当日 亚吉 把 洗革拉 赐给他，因此 洗革拉 属于 犹大 王，直到今日。
1SAM|27|7|大卫 在 非利士 人的地，住的期间有一年四个月。
1SAM|27|8|大卫 和他的人上去，侵夺 基述 人、 基色 人、 亚玛力 人，这些是从 帖兰 经过 书珥 直到 埃及 地的居民 。
1SAM|27|9|大卫 攻击那地，无论男女没有留下一个活口，又夺获牛、羊、驴、骆驼和衣服，回来到 亚吉 那里。
1SAM|27|10|亚吉 说：“今日你们没有去抢夺什么地方吧 ？” 大卫 说：“侵夺了 犹大 、 耶拉篾 、 基尼 等地的南方。”
1SAM|27|11|无论男女， 大卫 没有留下一个活口带到 迦特 来。他说：“恐怕他们把我们的事告诉人，说：‘ 大卫 如此做了。’”这是他住在 非利士 人之地一切日子的惯例。
1SAM|27|12|亚吉 信了 大卫 ，说：“ 大卫 已经使本族 以色列 人憎恶他，所以他必永远作我的仆人了。”
1SAM|28|1|那时， 非利士 人召集军队，要与 以色列 打仗。 亚吉 对 大卫 说：“你当知道，你和你的人都要随我出征。”
1SAM|28|2|大卫 对 亚吉 说：“好，仆人所能做的事，王都知道。” 亚吉 对 大卫 说：“好，我立你终生作我 的侍卫。”
1SAM|28|3|那时 撒母耳 已经死了， 以色列 众人为他哀哭，把他葬在他的本城 拉玛 。 扫罗 曾在国内驱除招魂的和行巫术的人。
1SAM|28|4|非利士 人集合，来到 书念 安营； 扫罗 集合 以色列 众人在 基利波 安营。
1SAM|28|5|扫罗 看见 非利士 的军队，就惧怕，心中大大战兢。
1SAM|28|6|扫罗 求问耶和华，耶和华却不藉梦，或乌陵，或先知回答他。
1SAM|28|7|扫罗 吩咐臣仆说：“为我找一个招魂的妇人，我好去问她。”臣仆对他说：“看哪，在 隐．多珥 有一个招魂的妇人。”
1SAM|28|8|于是 扫罗 改了装，穿上别的衣服，带着两个人，夜里去见那妇人。 扫罗 说：“请你用招魂的法术，把我所告诉你的死人，为我招上来。”
1SAM|28|9|妇人对他说：“看哪，你知道 扫罗 所做的，他从国中剪除招魂的和行巫术的。你为何为我的性命设下罗网，要害死我呢？”
1SAM|28|10|扫罗 向妇人指着耶和华起誓说：“我指着永生的耶和华起誓，你必不因这事受罚。”
1SAM|28|11|妇人说：“我为你招谁上来呢？”他说：“为我招 撒母耳 上来。”
1SAM|28|12|妇人看见 撒母耳 ，就大声喊叫。妇人对 扫罗 说：“你是 扫罗 ，为什么欺骗我呢？”
1SAM|28|13|王对妇人说：“不要惧怕，你看见什么呢？”妇人对 扫罗 说：“我看见有神明从地里上来。”
1SAM|28|14|扫罗 说：“他是怎样的形状？”妇人说：“有一个老人上来，身穿长袍。” 扫罗 知道是 撒母耳 ，就屈身，脸伏于地下拜。
1SAM|28|15|撒母耳 对 扫罗 说：“你为什么搅扰我，招我上来呢？” 扫罗 说：“我十分为难，因为 非利士 人攻击我，上帝离开我，不再藉先知或梦回答我。因此请你上来，好指示我应当怎样做。”
1SAM|28|16|撒母耳 说：“耶和华已经离开你，与你为敌，你何必问我呢？
1SAM|28|17|耶和华照他藉我所说的话为他自己 实现了。耶和华已经从你手里夺去国权，赐给别人，就是 大卫 。
1SAM|28|18|因为你没有听从耶和华的话，没有执行他对 亚玛力 人的恼怒，所以今日耶和华向你做这事。
1SAM|28|19|耶和华也必将你和 以色列 交在 非利士 人手里。明日你和你儿子们必与我在一处了；耶和华也必将 以色列 的军兵交在 非利士 人手里。”
1SAM|28|20|扫罗 突然全身仆倒在地，因为 撒母耳 的话令他十分惧怕。他毫无气力，因为他一日一夜都没有吃什么。
1SAM|28|21|妇人到 扫罗 面前，见他极其惊恐，对他说：“看哪，婢女听从了你，不顾惜自己的性命，遵从你吩咐我的话。
1SAM|28|22|现在求你也听婢女的话，让我在你面前摆上一点食物，你吃了才有气力上路。”
1SAM|28|23|扫罗 不肯，说：“我不吃。”但他的仆人和那妇人再三劝他，他才听他们的话，从地上起来，坐在床上。
1SAM|28|24|妇人急忙把家里的一只肥牛犊宰了，又拿面来揉，烤成无酵饼，
1SAM|28|25|摆在 扫罗 和他仆人面前。他们吃了，当夜就起身走了。
1SAM|29|1|非利士 人聚集他们所有的军队到 亚弗 ； 以色列 人在 耶斯列 的泉旁安营。
1SAM|29|2|非利士 人的领袖各率队伍，或百或千的前进； 大卫 和他的人同 亚吉 跟在后边前进。
1SAM|29|3|非利士 人的领袖说：“这些 希伯来 人在这里做什么呢？” 亚吉 对 非利士 人的领袖说：“这不是 以色列 王 扫罗 的臣仆 大卫 吗？他在我这里有些年日了。自从他投降直到今日，我未曾见他有什么过错。”
1SAM|29|4|非利士 人的领袖向 亚吉 发怒，对他说：“叫这人回去！叫他回到你指派他的地方去，不可让他同我们出征，免得他在阵上反成为我们的敌人。他用什么与他主人复和呢？岂不是用我们这些人的首级吗？
1SAM|29|5|有人跳舞唱和说： ‘ 扫罗 杀死千千， 大卫 杀死万万’， 不就是这个 大卫 吗？”
1SAM|29|6|亚吉 叫 大卫 来，对他说：“我指着永生的耶和华起誓，你是个正直人。你随我在军中出入，我也很满意。自从你投奔我到如今，我未曾看见你有什么过失，但是众领袖看你不顺眼。
1SAM|29|7|现在你平平安安地回去，不要做 非利士 人领袖眼中看为恶的事。”
1SAM|29|8|大卫 对 亚吉 说：“但我做了什么呢？自从仆人到你面前，直到今日，你查出我有什么过错，使我不去攻击我主我王的仇敌呢？”
1SAM|29|9|亚吉 回答 大卫 说：“我知道你在我眼中是好人，如同上帝的使者一样，只是 非利士 人的领袖说：‘这人不可同我们上战场。’
1SAM|29|10|现在，你和跟随你来的，就是你主人的仆人，清晨要早早起来，回到我所指派你的地方去，不要把中伤的话放在心上，因为你在我面前很好 。你们清晨早早起来，天一亮就回去吧！”
1SAM|29|11|于是 大卫 和他的人清晨早早起来，回到 非利士 人的地去。 非利士 人也上 耶斯列 去了。
1SAM|30|1|第三日， 大卫 和他的人到了 洗革拉 。 亚玛力 人已经侵夺 尼革夫 和 洗革拉 。他们攻破 洗革拉 ，用火焚烧。
1SAM|30|2|他们掳去城内的妇女和城中的大小人口，一个都没有杀，全都带走，他们就上路去了。
1SAM|30|3|大卫 和他的人到了那城，看哪，城已被火烧毁，他们的妻子儿女都被掳去了。
1SAM|30|4|大卫 和跟随他的百姓就放声大哭，直到没有气力再哭。
1SAM|30|5|大卫 的两个妻子， 耶斯列 人 亚希暖 和作过 拿八 妻子的 迦密 人 亚比该 ，也被掳去了。
1SAM|30|6|大卫 非常焦急，因为众百姓为自己的儿女痛心，说要用石头打死他。 大卫 却倚靠耶和华－他的上帝，坚定自己。
1SAM|30|7|大卫 对 亚希米勒 的儿子 亚比亚他 祭司说：“请你把以弗得拿来给我。” 亚比亚他 就把以弗得拿给 大卫 。
1SAM|30|8|大卫 求问耶和华说：“我追赶这群人，是否追得上呢？”耶和华对他说：“你可以追，一定追得上，也一定救得回来。”
1SAM|30|9|于是， 大卫 出发，他和跟随他的六百人来到 比梭溪 ，那些不能前去的就留在那里。
1SAM|30|10|大卫 带着四百人往前追赶；有二百人疲乏，不能过 比梭溪 ，留在那里。
1SAM|30|11|这四百人在田野遇见一个 埃及 人，就带他到 大卫 面前，给他饼吃，给他水喝，
1SAM|30|12|又给他一块无花果饼，两个葡萄干饼。他吃了，精神就恢复了，因为他三日三夜没有吃饼，没有喝水。
1SAM|30|13|大卫 对他说：“你是谁的人？你从哪里来？”他说：“我是 埃及 的青年，是 亚玛力 人的奴仆。因为我三天前生病，我主人就把我撇弃了。
1SAM|30|14|我们侵夺了 基利提 的南方和属 犹大 的地，以及 迦勒 地的南方，又用火烧了 洗革拉 。”
1SAM|30|15|大卫 对他说：“你肯领我们下到那群人那里吗？”他说：“你要向我指着上帝起誓，你不杀我，也不把我交在我主人手里，我就领你下到那群人那里。”
1SAM|30|16|那人领 大卫 下去，看哪，他们分散在全地面，吃喝跳舞，因为他们从 非利士 人的地和 犹大 地掳来的财物非常多。
1SAM|30|17|大卫 击杀他们，从黎明直到次日晚上，除了四百个骑骆驼逃走的青年之外，一个也没有逃脱。
1SAM|30|18|亚玛力 人所掳去的财物， 大卫 全都夺回，并救回他的两个妻子。
1SAM|30|19|凡 亚玛力 人所掳去的，无论大小、儿女、掠物和一切被掳去的， 大卫 全都夺回来。
1SAM|30|20|大卫 所夺来的牛群羊群，有人赶在群畜前面，说：“这是 大卫 的掠物。”
1SAM|30|21|大卫 到了那疲乏不能跟随、留在 比梭溪 的二百人那里。他们出来迎接 大卫 和跟随他的百姓。 大卫 上前向他们问安。
1SAM|30|22|跟随 大卫 去的人中，每一个恶人和无赖都说：“这些人既然没有和我同去，我们所夺的财物就不分给他们，只把他们各人的妻子儿女给他们，让他们带回去就好了。”
1SAM|30|23|大卫 说：“我的弟兄，耶和华所赐给我们的，你们不可这么做，因为他保佑了我们，把那群来攻击我们的人交在我们手里。
1SAM|30|24|谁肯在这事上听你们呢？上阵的分得多少，留下看守物件的也分得多少，大家应当平分。”
1SAM|30|25|从那日起， 大卫 定此为 以色列 的律例典章，直到今日。
1SAM|30|26|大卫 到了 洗革拉 ，从掠物中取些送给他的朋友，就是 犹大 的长老，说：“看哪，这是从耶和华仇敌那里夺来的，送给你们作礼物。”
1SAM|30|27|有在 伯特利 的， 尼革夫 之 拉末 的， 雅提珥 的，
1SAM|30|28|有在 亚罗珥 的， 息末 的， 以实提莫 的，
1SAM|30|29|有在 拉哈勒 的， 耶拉篾 各城的， 基尼 各城的，
1SAM|30|30|有在 何珥玛 的， 坡拉珊 的， 亚挞 的，
1SAM|30|31|有在 希伯仑 的，以及 大卫 和跟随他的人经常进出之处的。
1SAM|31|1|非利士 人攻打 以色列 。 以色列 人在 非利士 人面前逃跑，很多人 在 基利波山 被杀仆倒。
1SAM|31|2|非利士 人紧追 扫罗 和他的儿子，杀了 扫罗 的儿子 约拿单 、 亚比拿达 、 麦基．舒亚 。
1SAM|31|3|攻击 扫罗 的战事激烈，弓箭手追上他，他被弓箭手射中，伤势很重 。
1SAM|31|4|扫罗 吩咐拿他兵器的人说：“你拔出刀来，把我刺死，免得那些未受割礼的人来刺我，凌辱我。”但拿兵器的人不肯，因为他非常惧怕。于是 扫罗 拿起刀来，伏在刀上。
1SAM|31|5|拿兵器的人见 扫罗 已死，也伏在刀上跟他一起死。
1SAM|31|6|这样， 扫罗 和他三个儿子，与拿他兵器的人，以及他所有的人 ，都在那日一起死了。
1SAM|31|7|住平原那边和 约旦河 那边的 以色列 人，见 以色列 军兵逃跑， 扫罗 和他儿子都死了，就弃城逃跑。 非利士 人前来住在其中。
1SAM|31|8|次日， 非利士 人来剥那些被杀之人的衣服，看见 扫罗 和他三个儿子仆倒在 基利波山 。
1SAM|31|9|他们割下他的首级，剥了他的盔甲，派人到 非利士 人之地的四境，报信给他们庙里的偶像和百姓。
1SAM|31|10|他们将 扫罗 的盔甲放在 亚斯她录 庙里，把他的尸身钉在 伯．珊 的城墙上。
1SAM|31|11|基列 的 雅比 居民听见 非利士 人向 扫罗 所行的事，
1SAM|31|12|他们所有的勇士就起身，走了一夜，把 扫罗 和他儿子的尸身从 伯．珊 城墙上取下来，送到 雅比 ，在那里用火烧了，
1SAM|31|13|把骸骨葬在 雅比 的柳树下，并且禁食七日。
