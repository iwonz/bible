DAN|1|1|anno tertio regni Ioachim regis Iuda venit Nabuchodonosor rex Babylonis Hierusalem et obsedit eam
DAN|1|2|et tradidit Dominus in manu eius Ioachim regem Iudae et partem vasorum domus Dei et asportavit ea in terram Sennaar in domum dei sui et vasa intulit in domum thesauri dei sui
DAN|1|3|et ait rex Asfanaz praeposito eunuchorum suorum ut introduceret de filiis Israhel et de semine regio et tyrannorum
DAN|1|4|pueros in quibus nulla esset macula decoros forma et eruditos omni sapientia cautos scientia et doctos disciplina et qui possent stare in palatio regis ut doceret eos litteras et linguam Chaldeorum
DAN|1|5|et constituit eis rex annonam per singulos dies de cibis suis et de vino unde bibebat ipse ut enutriti tribus annis postea starent in conspectu regis
DAN|1|6|fuerunt ergo inter eos de filiis Iuda Danihel Ananias Misahel et Azarias
DAN|1|7|et inposuit eis praepositus eunuchorum nomina Daniheli Balthasar et Ananiae Sedrac Misaheli Misac et Azariae Abdenago
DAN|1|8|proposuit autem Danihel in corde suo ne pollueretur de mensa regis neque de vino potus eius et rogavit eunuchorum praepositum ne contaminaretur
DAN|1|9|dedit autem Deus Daniheli gratiam et misericordiam in conspectu principis eunuchorum
DAN|1|10|et ait princeps eunuchorum ad Danihel timeo ego dominum meum regem qui constituit vobis cibum et potum qui si viderit vultus vestros macilentiores prae ceteris adulescentibus coaevis vestris condemnabitis caput meum regi
DAN|1|11|et dixit Danihel ad Malassar quem constituerat princeps eunuchorum super Danihel Ananiam Misahel et Azariam
DAN|1|12|tempta nos obsecro servos tuos diebus decem et dentur nobis legumina ad vescendum et aqua ad bibendum
DAN|1|13|et contemplare vultus nostros et vultus puerorum qui vescuntur cibo regio et sicut videris facies cum servis tuis
DAN|1|14|qui audito sermone huiuscemodi temptavit eos diebus decem
DAN|1|15|post dies autem decem apparuerunt vultus eorum meliores et corpulentiores prae omnibus pueris qui vescebantur cibo regio
DAN|1|16|porro Malassar tollebat cibaria et vinum potus eorum dabatque eis legumina
DAN|1|17|pueris autem his dedit Deus scientiam et disciplinam in omni libro et sapientia Daniheli autem intellegentiam omnium visionum et somniorum
DAN|1|18|conpletis itaque diebus post quos dixerat rex ut introducerentur introduxit eos praepositus eunuchorum in conspectu Nabuchodonosor
DAN|1|19|cumque locutus eis fuisset rex non sunt inventi de universis tales ut Danihel Ananias Misahel et Azarias et steterunt in conspectu regis
DAN|1|20|et omne verbum sapientiae et intellectus quod sciscitatus est ab eis rex invenit in eis decuplum super cunctos ariolos et magos qui erant in universo regno eius
DAN|1|21|fuit autem Danihel usque ad annum primum Cyri regis
DAN|2|1|in anno secundo regni Nabuchodonosor vidit Nabuchodonosor somnium et conterritus est spiritus eius et somnium eius fugit ab eo
DAN|2|2|praecepit ergo rex ut convocarentur arioli et magi et malefici et Chaldei et indicarent regi somnia sua qui cum venissent steterunt coram rege
DAN|2|3|et dixit ad eos rex vidi somnium et mente confusus ignoro quid viderim
DAN|2|4|responderuntque Chaldei regi syriace rex in sempiternum vive dic somnium servis tuis et interpretationem eius indicabimus
DAN|2|5|et respondens rex ait Chaldeis sermo recessit a me nisi indicaveritis mihi somnium et coniecturam eius peribitis vos et domus vestrae publicabuntur
DAN|2|6|si autem somnium et coniecturam eius narraveritis praemia et dona et honorem multum accipietis a me somnium igitur et interpretationem eius indicate mihi
DAN|2|7|responderunt secundo atque dixerunt rex somnium dicat servis suis et interpretationem illius indicabimus
DAN|2|8|respondit rex et ait certo novi quia tempus redimitis scientes quod recesserit a me sermo
DAN|2|9|si ergo somnium non indicaveritis mihi una est de vobis sententia quod interpretationem quoque fallacem et deceptione plenam conposueritis ut loquamini mihi donec tempus pertranseat somnium itaque dicite mihi ut sciam quod interpretationem quoque eius veram loquamini
DAN|2|10|respondentes ergo Chaldei coram rege dixerunt non est homo super terram qui sermonem tuum rex possit implere sed neque regum quisquam magnus et potens verbum huiuscemodi sciscitatur ab omni ariolo et mago et Chaldeo
DAN|2|11|sermo enim quem tu rex quaeris gravis est nec repperietur quisquam qui indicet illum in conspectu regis exceptis diis quorum non est cum hominibus conversatio
DAN|2|12|quo audito rex in furore et in ira magna praecepit ut perirent omnes sapientes Babylonis
DAN|2|13|et egressa sententia sapientes interficiebantur quaerebaturque Danihel et socii eius ut perirent
DAN|2|14|tunc Danihel requisivit de lege atque sententia ab Arioch principe militiae regis qui egressus fuerat ad interficiendos sapientes Babylonis
DAN|2|15|et interrogavit eum qui a rege acceperat potestatem quam ob causam tam crudelis sententia a facie esset regis egressa cum ergo rem indicasset Arioch Daniheli
DAN|2|16|Danihel ingressus rogavit regem ut tempus daret sibi ad solutionem indicandam regi
DAN|2|17|et ingressus est domum suam Ananiaeque Misaheli et Azariae sociis suis indicavit negotium
DAN|2|18|ut quaererent misericordiam a facie Dei caeli super sacramento isto et non perirent Danihel et socii eius cum ceteris sapientibus Babylonis
DAN|2|19|tunc Daniheli per visionem nocte mysterium revelatum est et Danihel benedixit Deo caeli
DAN|2|20|et locutus ait sit nomen Domini benedictum a saeculo et usque in saeculum quia sapientia et fortitudo eius sunt
DAN|2|21|et ipse mutat tempora et aetates transfert regna atque constituit dat sapientiam sapientibus et scientiam intellegentibus disciplinam
DAN|2|22|ipse revelat profunda et abscondita et novit in tenebris constituta et lux cum eo est
DAN|2|23|tibi Deus patrum meorum confiteor teque laudo quia sapientiam et fortitudinem dedisti mihi et nunc ostendisti mihi quae rogavimus te quia sermonem regis aperuisti nobis
DAN|2|24|post haec Danihel ingressus ad Arioch quem constituerat rex ut perderet sapientes Babylonis sic ei locutus est sapientes Babylonis ne perdas introduc me in conspectu regis et solutionem regi enarrabo
DAN|2|25|tunc Arioch festinus introduxit Danihelem ad regem et dixit ei inveni hominem de filiis transmigrationis Iudae qui solutionem regi adnuntiet
DAN|2|26|respondit rex et dixit Daniheli cuius nomen erat Balthasar putasne vere potes indicare mihi somnium quod vidi et interpretationem eius
DAN|2|27|et respondens Danihel coram rege ait mysterium quod rex interrogat sapientes magi et arioli et aruspices non queunt indicare regi
DAN|2|28|sed est Deus in caelo revelans mysteria qui indicavit tibi rex Nabuchodonosor quae ventura sunt novissimis temporibus somnium tuum et visiones capitis tui in cubili tuo huiuscemodi sunt
DAN|2|29|tu rex cogitare coepisti in stratu tuo quid esset futurum post haec et qui revelat mysteria ostendit tibi quae ventura sunt
DAN|2|30|mihi quoque non in sapientia quae est in me plus quam in cunctis viventibus sacramentum hoc revelatum est sed ut interpretatio regi manifesta fieret et cogitationes mentis tuae scires
DAN|2|31|tu rex videbas et ecce quasi statua una grandis statua illa magna et statura sublimis stabat contra te et intuitus eius erat terribilis
DAN|2|32|huius statuae caput ex auro optimo erat pectus autem et brachia de argento porro venter et femora ex aere
DAN|2|33|tibiae autem ferreae pedum quaedam pars erat ferrea quaedam fictilis
DAN|2|34|videbas ita donec abscisus est lapis sine manibus et percussit statuam in pedibus eius ferreis et fictilibus et comminuit eos
DAN|2|35|tunc contrita sunt pariter ferrum testa aes argentum et aurum et redacta quasi in favillam aestivae areae rapta sunt vento nullusque locus inventus est eis lapis autem qui percusserat statuam factus est mons magnus et implevit universam terram
DAN|2|36|hoc est somnium interpretationem quoque eius dicemus coram te rex
DAN|2|37|tu rex regum es et Deus caeli regnum fortitudinem et imperium et gloriam dedit tibi
DAN|2|38|et omnia in quibus habitant filii hominum et bestiae agri volucresque caeli dedit in manu tua et sub dicione tua universa constituit tu es ergo caput aureum
DAN|2|39|et post te consurget regnum aliud minus te et regnum tertium aliud aereum quod imperabit universae terrae
DAN|2|40|et regnum quartum erit velut ferrum quomodo ferrum comminuit et domat omnia sic comminuet omnia haec et conteret
DAN|2|41|porro quia vidisti pedum et digitorum partem testae figuli et partem ferream regnum divisum erit quod tamen de plantario ferri orietur secundum quod vidisti ferrum mixtum testae ex luto
DAN|2|42|et digitos pedum ex parte ferreos et ex parte fictiles ex parte regnum erit solidum et ex parte contritum
DAN|2|43|quia autem vidisti ferrum mixtum testae ex luto commiscebuntur quidem humano semine sed non adherebunt sibi sicuti ferrum misceri non potest testae
DAN|2|44|in diebus autem regnorum illorum suscitabit Deus caeli regnum quod in aeternum non dissipabitur et regnum eius populo alteri non tradetur comminuet et consumet universa regna haec et ipsum stabit in aeternum
DAN|2|45|secundum quod vidisti quod de monte abscisus est lapis sine manibus et comminuit testam et ferrum et aes et argentum et aurum Deus magnus ostendit regi quae futura sunt postea et verum est somnium et fidelis interpretatio eius
DAN|2|46|tunc rex Nabuchodonosor cecidit in faciem suam et Danihelum adoravit et hostias et incensum praecepit ut sacrificarent ei
DAN|2|47|loquens ergo rex ait Daniheli vere Deus vester Deus deorum est et Dominus regum et revelans mysteria quoniam potuisti aperire sacramentum hoc
DAN|2|48|tunc rex Danihelum in sublime extulit et munera multa et magna dedit ei et constituit eum principem super omnes provincias Babylonis et praefectum magistratuum super cunctos sapientes Babylonis
DAN|2|49|Danihel autem postulavit a rege et constituit super opera provinciae Babylonis Sedrac Misac et Abdenago ipse autem Danihel erat in foribus regis
DAN|3|1|Nabuchodonosor rex fecit statuam auream altitudine cubitorum sexaginta latitudine cubitorum sex et statuit eam in campo Duram provinciae Babylonis
DAN|3|2|itaque Nabuchodonosor rex misit ad congregandos satrapas magistratus et iudices duces et tyrannos et praefectos omnesque principes regionum ut convenirent ad dedicationem statuae quam erexerat Nabuchodonosor rex
DAN|3|3|tunc congregati sunt satrapae magistratus et iudices duces et tyranni et optimates qui erant in potestatibus constituti et universi principes regionum ut convenirent ad dedicationem statuae quam erexerat Nabuchodonosor rex stabant autem in conspectu statuae quam posuerat Nabuchodonosor
DAN|3|4|et praeco clamabat valenter vobis dicitur populis tribubus et linguis
DAN|3|5|in hora qua audieritis sonitum tubae et fistulae et citharae sambucae et psalterii et symphoniae et universi generis musicorum cadentes adorate statuam auream quam constituit Nabuchodonosor rex
DAN|3|6|si quis autem non prostratus adoraverit eadem hora mittetur in fornacem ignis ardentis
DAN|3|7|post haec igitur statim ut audierunt omnes populi sonitum tubae fistulae et citharae sambucae et psalterii et symphoniae et omnis generis musicorum cadentes omnes populi et tribus et linguae adoraverunt statuam auream quam constituerat Nabuchodonosor rex
DAN|3|8|statimque et in ipso tempore accedentes viri chaldei accusaverunt Iudaeos
DAN|3|9|dixeruntque Nabuchodonosor regi rex in aeternum vive
DAN|3|10|tu rex posuisti decretum ut omnis homo qui audierit sonitum tubae fistulae et citharae sambucae et psalterii et symphoniae et universi generis musicorum prosternat se et adoret statuam auream
DAN|3|11|si quis autem non procidens adoraverit mittatur in fornacem ignis ardentem
DAN|3|12|sunt ergo viri iudaei quos constituisti super opera regionis Babyloniae Sedrac Misac et Abdenago viri isti contempserunt rex decretum tuum deos tuos non colunt et statuam auream quam erexisti non adorant
DAN|3|13|tunc Nabuchodonosor in furore et in ira praecepit ut adducerentur Sedrac Misac et Abdenago qui confestim adducti sunt in conspectu regis
DAN|3|14|pronuntiansque Nabuchodonosor rex ait eis verene Sedrac Misac et Abdenago deos meos non colitis et statuam auream quam constitui non adoratis
DAN|3|15|nunc ergo si estis parati quacumque hora audieritis sonitum tubae fistulae et citharae sambucae psalterii et symphoniae omnisque generis musicorum prosternite vos et adorate statuam quam feci quod si non adoraveritis eadem hora mittemini in fornacem ignis ardentem et quis est Deus qui eripiat vos de manu mea
DAN|3|16|respondentes Sedrac Misac et Abdenago dixerunt regi Nabuchodonosor non oportet nos de hac re respondere tibi
DAN|3|17|ecce enim Deus noster quem colimus potest eripere nos de camino ignis ardentis et de manibus tuis rex liberare
DAN|3|18|quod si noluerit notum tibi sit rex quia deos tuos non colimus et statuam auream quam erexisti non adoramus
DAN|3|19|tunc Nabuchodonosor repletus est furore et aspectus faciei illius inmutatus est super Sedrac Misac et Abdenago et praecepit ut succenderetur fornax septuplum quam succendi consuerat
DAN|3|20|et viris fortissimis de exercitu suo iussit ut ligatis pedibus Sedrac Misac et Abdenago mitterent eos in fornacem ignis ardentem
DAN|3|21|et confestim viri illi vincti cum bracis suis et tiaris et calciamentis et vestibus missi sunt in medium fornacis ignis ardentis
DAN|3|22|nam iussio regis urguebat fornax autem succensa erat nimis porro viros illos qui miserant Sedrac Misac et Abdenago interfecit flamma ignis
DAN|3|23|viri autem hii id est tres Sedrac Misac et Abdenago ceciderunt in medio camini ignis ardentis conligati
DAN|3|24|et ambulabant in medio flammae laudantes Deum et benedicentes Domino
DAN|3|25|stans autem Azarias oravit sic aperiensque os suum in medio ignis ait
DAN|3|26|benedictus es Domine Deus patrum nostrorum et laudabilis et gloriosum nomen tuum in saecula
DAN|3|27|quia iustus es in omnibus quae fecisti nobis et universa opera tua vera et viae tuae rectae et omnia iudicia tua vera
DAN|3|28|iudicia enim vera fecisti iuxta omnia quae induxisti super nos et super civitatem sanctam patrum nostrorum Hierusalem quia in veritate et in iudicio induxisti omnia haec propter peccata nostra
DAN|3|29|peccavimus enim et inique egimus recedentes a te et deliquimus in omnibus
DAN|3|30|et praecepta tua non audivimus nec observavimus nec fecimus sicut praeceperas nobis ut bene nobis esset
DAN|3|31|omnia ergo quae induxisti super nos et universa quae fecisti nobis vero iudicio fecisti
DAN|3|32|et tradidisti nos in manibus inimicorum iniquorum et pessimorum praevaricatorumque et regi iniusto et pessimo ultra omnem terram
DAN|3|33|et nunc non possumus aperire os confusio et obprobrium facti sumus servis tuis et his qui colunt te
DAN|3|34|ne quaesumus tradas nos in perpetuum propter nomen tuum et ne dissipes testamentum tuum
DAN|3|35|neque auferas misericordiam tuam a nobis propter Abraham dilectum tuum et Isaac servum tuum et Israhel sanctum tuum
DAN|3|36|quibus locutus es pollicens quod multiplicares semen eorum sicut stellas caeli et sicut harenam quae est in litore maris
DAN|3|37|quia Domine inminuti sumus plus quam omnes gentes sumusque humiles in universa terra hodie propter peccata nostra
DAN|3|38|et non est in tempore hoc princeps et propheta et dux neque holocaustum neque sacrificium neque oblatio neque incensum neque locus primitiarum coram te
DAN|3|39|ut possimus invenire misericordiam sed in anima contrita et spiritu humilitatis suscipiamur
DAN|3|40|sicut in holocaustum arietum et taurorum et sicut in milibus agnorum pinguium sic fiat sacrificium nostrum in conspectu tuo hodie ut placeat tibi quoniam non est confusio confidentibus in te
DAN|3|41|et nunc sequimur in toto corde et timemus te et quaerimus faciem tuam
DAN|3|42|ne confundas nos sed fac nobiscum iuxta mansuetudinem tuam et secundum multitudinem misericordiae tuae
DAN|3|43|et erue nos in mirabilibus tuis et da gloriam nomini tuo Domine
DAN|3|44|et confundantur omnes qui ostendunt servis tuis mala confundantur in omni potentia et robur eorum conteratur
DAN|3|45|sciant quia tu Domine Deus solus et gloriosus super orbem terrarum
DAN|3|46|et non cessabant qui inmiserant eos ministri regis succendere fornacem naptha et stuppa et pice et malleolis
DAN|3|47|et effundebatur flamma super fornacem cubitis quadraginta novem
DAN|3|48|et erupit et incendit quos repperit iuxta fornacem de Chaldeis
DAN|3|49|angelus autem descendit cum Azaria et sociis eius in fornacem et excussit flammam ignis de fornace
DAN|3|50|et fecit medium fornacis quasi ventum roris flantem et non tetigit eos omnino ignis neque contristavit nec quicquam molestiae intulit
DAN|3|51|tunc hii tres quasi ex uno ore laudabant et glorificabant et benedicebant Deo in fornace dicentes
DAN|3|52|benedictus es Domine Deus patrum nostrorum et laudabilis et superexaltatus in saecula et benedictum nomen gloriae tuae sanctum et laudabile et superexaltatum in omnibus saeculis
DAN|3|53|benedictus es in templo sancto gloriae tuae et superlaudabilis et supergloriosus in saecula
DAN|3|54|benedictus es in throno regni tui et superlaudabilis et superexaltatus in saecula
DAN|3|55|benedictus es qui intueris abyssos et sedes super cherubin et laudabilis et superexaltatus in saecula
DAN|3|56|benedictus es in firmamento caeli et laudabilis et gloriosus in saecula
DAN|3|57|benedicite omnia opera Domini Domino laudate et superexaltate eum in saecula
DAN|3|58|benedicite angeli Domino laudate et superexaltate eum in saecula
DAN|3|59|benedicite caeli Domino laudate et superexaltate eum in saecula
DAN|3|60|benedicite aquae omnes quae super caelos sunt Domino laudate et superexaltate eum in saecula
DAN|3|61|benedicite omnes virtutes Domini Domino laudate et superexaltate eum in saecula
DAN|3|62|benedicite sol et luna Domino laudate et superexaltate eum in saecula
DAN|3|63|benedicite stellae caeli Domino laudate et superexaltate eum in saecula
DAN|3|64|benedicite omnis imber et ros Domino laudate et superexaltate eum in saecula
DAN|3|65|benedicite omnis spiritus Domino laudate et superexaltate eum in saecula
DAN|3|66|benedicite ignis et aestus Domino laudate et superexaltate eum in saecula
DAN|3|67|benedicite frigus et aestus Domino laudate et superexaltate eum in saecula
DAN|3|68|benedicite rores et pruina Domino laudate et superexaltate eum in saecula
DAN|3|69|benedicite gelu et frigus Domino laudate et superexaltate eum in saecula
DAN|3|70|benedicite glacies et nives Domino laudate et superexaltate eum in saecula
DAN|3|71|benedicite noctes et dies Domino laudate et superexaltate eum in saecula
DAN|3|72|benedicite lux et tenebrae Domino laudate et superexaltate eum in saecula
DAN|3|73|benedicite fulgura et nubes Domino laudate et superexaltate eum in saecula
DAN|3|74|benedicat terra Dominum laudet et superexaltet eum in saecula
DAN|3|75|benedicite montes et colles Domino laudate et superexaltate eum in saecula
DAN|3|76|benedicite universa germinantia in terra Domino laudate et superexaltate eum in saecula
DAN|3|77|benedicite fontes Domino laudate et superexaltate eum in saecula
DAN|3|78|benedicite maria et flumina Domino laudate et superexaltate eum in saecula
DAN|3|79|benedicite cete et omnia quae moventur in aquis Domino laudate et superexaltate eum in saecula
DAN|3|80|benedicite omnes volucres caeli Domino laudate et superexaltate eum in saecula
DAN|3|81|benedicite omnes bestiae et pecora Domino laudate et superexaltate eum in saecula
DAN|3|82|benedicite filii hominum Domino laudate et superexaltate eum in saecula
DAN|3|83|benedic Israhel Domino laudate et superexaltate eum in saecula
DAN|3|84|benedicite sacerdotes Domini Domino laudate et superexaltate eum in saecula
DAN|3|85|benedicite servi Domini Domino laudate et superexaltate eum in saecula
DAN|3|86|benedicite spiritus et animae iustorum Domino laudate et superexaltate eum in saecula
DAN|3|87|benedicite sancti et humiles corde Domino laudate et superexaltate eum in saecula
DAN|3|88|benedicite Anania Azaria et Misahel Domino laudate et superexaltate eum in saecula quia eruit nos de inferno et salvos fecit de manu mortis et liberavit de medio ardentis flammae et de medio ignis eruit nos
DAN|3|89|confitemini Domino quoniam bonus quoniam in saeculum misericordia eius
DAN|3|90|benedicite omnes religiosi Domino Deo deorum laudate et confitemini quia in omnia saecula misericordia eius
DAN|3|91|tunc Nabuchodonosor rex obstipuit et surrexit propere et ait optimatibus suis nonne tres viros misimus in medio ignis conpeditos qui respondentes dixerunt regi vere rex
DAN|3|92|respondit et ait ecce ego video viros quattuor solutos et ambulantes in medio ignis et nihil corruptionis in eis est et species quarti similis filio Dei
DAN|3|93|tunc accessit Nabuchodonosor ad ostium fornacis ignis ardentis et ait Sedrac Misac et Abdenago servi Dei excelsi egredimini et venite statimque egressi sunt Sedrac Misac et Abdenago de medio ignis
DAN|3|94|et congregati satrapae magistratus et iudices et potentes regis contemplabantur viros illos quoniam nihil potestatis habuisset ignis in corporibus eorum et capillus capitis eorum non esset adustus et sarabara eorum non fuissent inmutata et odor ignis non transisset per eos
DAN|3|95|et erumpens Nabuchodonosor ait benedictus Deus eorum Sedrac videlicet Misac et Abdenago qui misit angelum suum et eruit servos suos quia crediderunt in eo et verbum regis inmutaverunt et tradiderunt corpora sua ne servirent et ne adorarent omnem deum excepto Deo suo
DAN|3|96|a me ergo positum est hoc decretum ut omnis populus et tribus et lingua quaecumque locuta fuerit blasphemiam contra Deum Sedrac Misac et Abdenago dispereat et domus eius vastetur neque enim est Deus alius qui possit ita salvare
DAN|3|97|tunc rex promovit Sedrac Misac et Abdenago in provincia Babylonis
DAN|3|98|Nabuchodonosor rex omnibus populis gentibus et linguis quae habitant in universa terra pax vobis multiplicetur
DAN|3|99|signa et mirabilia fecit apud me Deus excelsus placuit ergo mihi praedicare
DAN|3|100|signa eius quia magna sunt et mirabilia eius quia fortia et regnum eius regnum sempiternum et potestas eius in generationem et generationem
DAN|4|1|ego Nabuchodonosor quietus eram in domo mea et florens in palatio meo
DAN|4|2|somnium vidi quod perterruit me et cogitationes meae in stratu meo et visiones capitis mei conturbaverunt me
DAN|4|3|et per me propositum est decretum ut introducerentur in conspectu meo cuncti sapientes Babylonis et ut solutionem somnii indicarent mihi
DAN|4|4|tunc ingrediebantur arioli magi Chaldei et aruspices et somnium narravi in conspectu eorum et solutionem eius non indicaverunt mihi
DAN|4|5|donec collega ingressus est in conspectu meo Danihel cuius nomen Balthasar secundum nomen dei mei qui habet spiritum deorum sanctorum in semet ipso et somnium coram eo locutus sum
DAN|4|6|Balthasar princeps ariolorum quem ego scio quod spiritum deorum sanctorum habeas in te et omne sacramentum non est inpossibile tibi visiones somniorum meorum quas vidi et solutionem eorum narra
DAN|4|7|visio capitis mei in cubili meo videbam et ecce arbor in medio terrae et altitudo eius nimia
DAN|4|8|magna arbor et fortis et proceritas eius contingens caelum aspectus illius erat usque ad terminos universae terrae
DAN|4|9|folia eius pulcherrima et fructus eius nimius et esca universorum in ea subter eam habitabant animalia et bestiae et in ramis eius conversabantur volucres caeli et ex ea vescebatur omnis caro
DAN|4|10|videbam in visione capitis mei super stratum meum et ecce vigil et sanctus de caelo descendit
DAN|4|11|clamavit fortiter et sic ait succidite arborem et praecidite ramos eius excutite folia eius et dispergite fructum eius fugiant bestiae quae subter eam sunt et volucres de ramis eius
DAN|4|12|verumtamen germen radicum eius in terra sinite et alligetur vinculo ferreo et aereo in herbis quae foris sunt et rore caeli tinguatur et cum feris pars eius in herba terrae
DAN|4|13|cor eius ab humano commutetur et cor ferae detur ei et septem tempora mutentur super eum
DAN|4|14|in sententia vigilum decretum est et sermo sanctorum et petitio donec cognoscant viventes quoniam dominatur Excelsus in regno hominum et cuicumque voluerit dabit illud et humillimum hominem constituet super eo
DAN|4|15|hoc somnium vidi ego rex Nabuchodonosor tu ergo Balthasar interpretationem narra festinus quia omnes sapientes regni mei non queunt solutionem edicere mihi tu autem potes quia spiritus deorum sanctorum in te est
DAN|4|16|tunc Danihel cuius nomen Balthasar coepit intra semet ipsum tacitus cogitare quasi hora una et cogitationes eius conturbabant eum respondens autem rex ait Balthasar somnium et interpretatio eius non conturbent te respondit Balthasar et dixit domine mi somnium his qui te oderunt et interpretatio eius hostibus tuis sit
DAN|4|17|arborem quam vidisti sublimem atque robustam cuius altitudo pertingit ad caelum et aspectus illius in omnem terram
DAN|4|18|et rami eius pulcherrimi et fructus eius nimius et esca omnium in ea subter eam habitantes bestiae agri et in ramis eius commorantes aves caeli
DAN|4|19|tu es rex qui magnificatus es et invaluisti et magnitudo tua crevit et pervenit usque ad caelum et potestas tua in terminos universae terrae
DAN|4|20|quod autem vidit rex vigilem et sanctum descendere de caelo et dicere succidite arborem et dissipate illam attamen germen radicum eius in terra dimittite et vinciatur ferro et aere in herbis foris et rore caeli conspergatur et cum feris sit pabulum eius donec septem tempora commutentur super eum
DAN|4|21|haec est interpretatio sententiae Altissimi quae pervenit super dominum meum regem
DAN|4|22|eicient te ab hominibus et cum bestiis feris erit habitatio tua et faenum ut bos comedes et rore caeli infunderis septem quoque tempora mutabuntur super te donec scias quod dominetur Excelsus super regnum hominum et cuicumque voluerit det illud
DAN|4|23|quod autem praecepit ut relinqueretur germen radicum eius id est arboris regnum tuum tibi manebit postquam cognoveris potestatem esse caelestem
DAN|4|24|quam ob rem rex consilium meum placeat tibi et peccata tua elemosynis redime et iniquitates tuas misericordiis pauperum forsitan ignoscat delictis tuis
DAN|4|25|omnia venerunt super Nabuchodonosor regem
DAN|4|26|post finem mensuum duodecim in aula Babylonis deambulabat
DAN|4|27|responditque rex et ait nonne haec est Babylon magna quam ego aedificavi in domum regni in robore fortitudinis meae et in gloria decoris mei
DAN|4|28|cum adhuc sermo esset in ore regis vox de caelo ruit tibi dicitur Nabuchodonosor rex regnum transiit a te
DAN|4|29|et ab hominibus te eicient et cum bestiis feris erit habitatio tua faenum quasi bos comedes et septem tempora mutabuntur super te donec scias quod dominetur Excelsus in regno hominum et cuicumque voluerit det illud
DAN|4|30|eadem hora sermo conpletus est super Nabuchodonosor ex hominibus abiectus est et faenum ut bos comedit et rore caeli corpus eius infectum est donec capilli eius in similitudinem aquilarum crescerent et ungues eius quasi avium
DAN|4|31|igitur post finem dierum ego Nabuchodonosor oculos meos ad caelum levavi et sensus meus redditus est mihi et Altissimo benedixi et viventem in sempiternum laudavi et glorificavi quia potestas eius potestas sempiterna et regnum eius in generationem et generationem
DAN|4|32|et omnes habitatores terrae apud eum in nihilum reputati sunt iuxta voluntatem enim suam facit tam in virtutibus caeli quam in habitatoribus terrae et non est qui resistat manui eius et dicat ei quare fecisti
DAN|4|33|in ipso tempore sensus meus reversus est ad me et ad honorem regni mei decoremque perveni et figura mea reversa est ad me et optimates mei et magistratus mei requisierunt me et in regno meo constitutus sum et magnificentia amplior addita est mihi
DAN|4|34|nunc igitur ego Nabuchodonosor laudo et magnifico et glorifico Regem caeli quia omnia opera eius vera et viae eius iudicia et gradientes in superbia potest humiliare
DAN|5|1|Balthasar rex fecit grande convivium optimatibus suis mille et unusquisque secundum suam bibebat aetatem
DAN|5|2|praecepit ergo iam temulentus ut adferrentur vasa aurea et argentea quae asportaverat Nabuchodonosor pater eius de templo quod fuit in Hierusalem ut biberent in eis rex et optimates eius uxoresque eius et concubinae
DAN|5|3|tunc adlata sunt vasa aurea quae asportaverat de templo quod fuerat in Hierusalem et biberunt in eis rex et optimates eius uxores et concubinae illius
DAN|5|4|bibebant vinum et laudabant deos suos aureos et argenteos et aereos ferreos ligneosque et lapideos
DAN|5|5|in eadem hora apparuerunt digiti quasi manus hominis scribentis contra candelabrum in superficie parietis aulae regiae et rex aspiciebat articulos manus scribentis
DAN|5|6|tunc regis facies commutata est et cogitationes eius conturbabant eum et conpages renum eius solvebantur et genua eius ad se invicem conlidebantur
DAN|5|7|exclamavit itaque rex fortiter ut introducerent magos Chaldeos et aruspices et proloquens rex ait sapientibus Babylonis quicumque legerit scripturam hanc et interpretationem eius manifestam mihi fecerit purpura vestietur et torquem auream habebit in collo et tertius in regno meo erit
DAN|5|8|tunc ingressi omnes sapientes regis non potuerunt nec scripturam legere nec interpretationem indicare regi
DAN|5|9|unde rex Balthasar satis conturbatus est et vultus illius inmutatus est sed et optimates eius turbabantur
DAN|5|10|regina autem pro re quae acciderat regi et optimatibus eius domum convivii ingressa est et proloquens ait rex in aeternum vive non te conturbent cogitationes tuae neque facies tua inmutetur
DAN|5|11|est vir in regno tuo qui spiritum deorum sanctorum habet in se et in diebus patris tui scientia et sapientia inventae sunt in eo nam et rex Nabuchodonosor pater tuus principem magorum incantatorum Chaldeorum et aruspicum constituit eum pater inquam tuus o rex
DAN|5|12|quia spiritus amplior et prudentia intellegentiaque interpretatio somniorum et ostensio secretorum ac solutio ligatorum inventae sunt in eo hoc est in Danihelo cui rex posuit nomen Balthasar nunc itaque Danihel vocetur et interpretationem narrabit
DAN|5|13|igitur introductus est Danihel coram rege ad quem praefatus rex ait tu es Danihel de filiis captivitatis Iudae quam adduxit rex pater meus de Iudaea
DAN|5|14|audivi de te quoniam spiritum deorum habeas et scientia intellegentiaque ac sapientia ampliores inventae sint in te
DAN|5|15|et nunc introgressi sunt in conspectu meo sapientes magi ut scripturam hanc legerent et interpretationem eius indicarent mihi et nequiverunt sensum sermonis huius edicere
DAN|5|16|porro ego audivi de te quod possis obscura interpretari et ligata dissolvere si ergo vales scripturam legere et interpretationem indicare mihi purpura vestieris et torquem auream circa collum tuum habebis et tertius in regno meo princeps eris
DAN|5|17|ad quae respondens Danihel ait coram rege munera tua sint tibi et dona domus tuae alteri da scripturam autem legam tibi rex et interpretationem eius ostendam tibi
DAN|5|18|o rex Deus altissimus regnum et magnificentiam gloriam et honorem dedit Nabuchodonosor patri tuo
DAN|5|19|et propter magnificentiam quam dederat ei universi populi tribus et linguae tremebant et metuebant eum quos volebat interficiebat et quos volebat percutiebat quos volebat exaltabat et quos volebat humiliabat
DAN|5|20|quando autem elevatum est cor eius et spiritus illius obfirmatus est ad superbiam depositus est de solio regni sui et gloria eius ablata est
DAN|5|21|et a filiis hominum eiectus est sed et cor eius cum bestiis positum est et cum onagris erat habitatio eius faenum quoque ut bos comedebat et rore caeli corpus eius infectum est donec cognosceret quod potestatem habeat Altissimus in regno hominum et quemcumque voluerit suscitabit super illud
DAN|5|22|tu quoque filius eius Balthasar non humiliasti cor tuum cum scires haec omnia
DAN|5|23|sed adversum Dominatorem caeli elevatus es et vasa domus eius adlata sunt coram te et tu et optimates tui et uxores tuae et concubinae vinum bibistis in eis deos quoque argenteos et aureos et aereos ferreos ligneosque et lapideos qui non vident neque audiunt neque sentiunt laudasti porro Deum qui habet flatum tuum in manu sua et omnes vias tuas non glorificasti
DAN|5|24|idcirco ab eo missus est articulus manus quae scripsit hoc quod exaratum est
DAN|5|25|haec est autem scriptura quae digesta est mane thecel fares
DAN|5|26|et haec interpretatio sermonis mane numeravit Deus regnum tuum et conplevit illud
DAN|5|27|thecel adpensum est in statera et inventus es minus habens
DAN|5|28|fares divisum est regnum tuum et datum est Medis et Persis
DAN|5|29|tunc iubente rege indutus est Danihel purpura et circumdata est torques aurea collo eius et praedicatum est de eo quod haberet potestatem tertius in regno
DAN|5|30|eadem nocte interfectus est Balthasar rex Chaldeus
DAN|5|31|et Darius Medus successit in regnum annos natus sexaginta duo
DAN|6|1|placuit Dario et constituit supra regnum satrapas centum viginti ut essent in toto regno suo
DAN|6|2|et super eos principes tres ex quibus Danihel unus erat ut satrapae illis redderent rationem et rex non sustineret molestiam
DAN|6|3|igitur Danihel superabat omnes principes et satrapas quia spiritus Dei amplior erat in eo
DAN|6|4|porro rex cogitabat constituere eum super omne regnum unde principes et satrapae quaerebant occasionem ut invenirent Daniheli ex latere regni nullamque causam et suspicionem repperire potuerunt eo quod fidelis esset et omnis culpa et suspicio non inveniretur in eo
DAN|6|5|dixerunt ergo viri illi non inveniemus Daniheli huic aliquam occasionem nisi forte in lege Dei sui
DAN|6|6|tunc principes et satrapae subripuerunt regi et sic locuti sunt ei Darie rex in aeternum vive
DAN|6|7|consilium inierunt cuncti principes regni magistratus et satrapae senatores et iudices ut decretum imperatorium exeat et edictum ut omnis qui petierit aliquam petitionem a quocumque deo et homine usque ad dies triginta nisi a te rex mittatur in lacum leonum
DAN|6|8|nunc itaque rex confirma sententiam et scribe decretum ut non inmutetur quod statutum est a Medis atque Persis nec praevaricari cuiquam liceat
DAN|6|9|porro rex Darius proposuit edictum et statuit
DAN|6|10|quod cum Danihel conperisset id est constitutam legem ingressus est domum suam et fenestris apertis in cenaculo suo contra Hierusalem tribus temporibus in die flectebat genua sua et adorabat confitebaturque coram Deo suo sicut et ante facere consueverat
DAN|6|11|viri igitur illi curiosius inquirentes invenerunt Danihel orantem et obsecrantem Deum suum
DAN|6|12|et accedentes locuti sunt regi super edicto rex numquid non constituisti ut omnis homo qui rogaret quemquam de diis et hominibus usque ad dies triginta nisi a te rex mitteretur in lacum leonum ad quod respondens rex ait verus sermo iuxta decretum Medorum atque Persarum quod praevaricari non licet
DAN|6|13|tunc respondentes dixerunt coram rege Danihel de filiis captivitatis Iudae non curavit de lege tua et de edicto quod constituisti sed tribus temporibus per diem orat obsecratione sua
DAN|6|14|quod verbum cum audisset rex satis contristatus est et pro Danihel posuit cor ut liberaret eum et usque ad occasum solis laborabat ut erueret illum
DAN|6|15|viri autem illi intellegentes regem dixerunt ei scito rex quia lex Medorum est atque Persarum ut omne decretum quod constituit rex non liceat inmutari
DAN|6|16|tunc rex praecepit et adduxerunt Danihelem et miserunt eum in lacum leonum dixitque rex Daniheli Deus tuus quem colis semper ipse liberabit te
DAN|6|17|adlatusque est lapis unus et positus est super os laci quem obsignavit rex anulo suo et anulo optimatum suorum ne quid fieret contra Danihel
DAN|6|18|et abiit rex in domum suam et dormivit incenatus cibique non sunt inlati coram eo insuper et somnus recessit ab eo
DAN|6|19|tunc rex primo diluculo consurgens festinus ad lacum leonum perrexit
DAN|6|20|adpropinquansque lacui Danihelem voce lacrimabili inclamavit et affatus est eum Danihel serve Dei viventis Deus tuus cui tu servis semper putasne valuit liberare te a leonibus
DAN|6|21|et Danihel regi respondens ait rex in aeternum vive
DAN|6|22|Deus meus misit angelum suum et conclusit ora leonum et non nocuerunt mihi quia coram eo iustitia inventa est in me sed et coram te rex delictum non feci
DAN|6|23|tunc rex vehementer gavisus est super eo et Danihelem praecepit educi de lacu eductusque est Danihel de lacu et nulla laesio inventa est in eo quia credidit Deo suo
DAN|6|24|iubente autem rege adducti sunt viri illi qui accusaverant Danihelem et in lacum leonum missi sunt ipsi et filii et uxores eorum et non pervenerunt usque ad pavimentum laci donec arriperent eos leones et omnia ossa eorum comminuerunt
DAN|6|25|tunc Darius rex scripsit universis populis tribubus et linguis habitantibus in universa terra pax vobis multiplicetur
DAN|6|26|a me constitutum est decretum ut in universo imperio et regno meo tremescant et paveant Deum Danihelis ipse est enim Deus vivens et aeternus in saecula et regnum eius non dissipabitur et potestas eius usque in aeternum
DAN|6|27|ipse liberator atque salvator faciens signa et mirabilia in caelo et in terra qui liberavit Danihelem de manu leonum
DAN|6|28|porro Danihel perseveravit usque ad regnum Darii regnumque Cyri Persae
DAN|7|1|anno primo Balthasar regis Babylonis Danihel somnium vidit visio autem capitis eius in cubili suo et somnium scribens brevi sermone conprehendit summatimque perstringens ait
DAN|7|2|videbam in visione mea nocte et ecce quattuor venti caeli pugnabant in mari magno
DAN|7|3|et quattuor bestiae grandes ascendebant de mari diversae inter se
DAN|7|4|prima quasi leaena et alas habebat aquilae aspiciebam donec evulsae sunt alae eius et sublata est de terra et super pedes quasi homo stetit et cor eius datum est ei
DAN|7|5|et ecce bestia alia similis urso in parte stetit et tres ordines erant in ore eius et in dentibus eius et sic dicebant ei surge comede carnes plurimas
DAN|7|6|post hoc aspiciebam et ecce alia quasi pardus et alas habebat avis quattuor super se et quattuor capita erant in bestia et potestas data est ei
DAN|7|7|post hoc aspiciebam in visione noctis et ecce bestia quarta terribilis atque mirabilis et fortis nimis dentes ferreos habebat magnos comedens atque comminuens et reliqua pedibus suis conculcans dissimilis autem erat ceteris bestiis quas videram ante eam et habebat cornua decem
DAN|7|8|considerabam cornua et ecce cornu aliud parvulum ortum est de medio eorum et tria de cornibus primis evulsa sunt a facie eius et ecce oculi quasi oculi hominis erant in cornu isto et os loquens ingentia
DAN|7|9|aspiciebam donec throni positi sunt et antiquus dierum sedit vestimentum eius quasi nix candidum et capilli capitis eius quasi lana munda thronus eius flammae ignis rotae eius ignis accensus
DAN|7|10|fluvius igneus rapidusque egrediebatur a facie eius milia milium ministrabant ei et decies milies centena milia adsistebant ei iudicium sedit et libri aperti sunt
DAN|7|11|aspiciebam propter vocem sermonum grandium quos cornu illud loquebatur et vidi quoniam interfecta esset bestia et perisset corpus eius et traditum esset ad conburendum igni
DAN|7|12|aliarum quoque bestiarum ablata esset potestas et tempora vitae constituta essent eis usque ad tempus et tempus
DAN|7|13|aspiciebam ergo in visione noctis et ecce cum nubibus caeli quasi filius hominis veniebat et usque ad antiquum dierum pervenit et in conspectu eius obtulerunt eum
DAN|7|14|et dedit ei potestatem et honorem et regnum et omnes populi tribus ac linguae ipsi servient potestas eius potestas aeterna quae non auferetur et regnum eius quod non corrumpetur
DAN|7|15|horruit spiritus meus ego Danihel territus sum in his et visiones capitis mei conturbaverunt me
DAN|7|16|accessi ad unum de adsistentibus et veritatem quaerebam ab eo de omnibus his qui dixit mihi interpretationem sermonum et edocuit me
DAN|7|17|hae bestiae magnae quattuor quattuor regna consurgent de terra
DAN|7|18|suscipient autem regnum sancti Dei altissimi et obtinebunt regnum usque in saeculum et saeculum saeculorum
DAN|7|19|post hoc volui diligenter discere de bestia quarta quia erat dissimilis valde ab omnibus et terribilis nimis dentes et ungues eius ferrei comedebat et comminuebat et reliquias pedibus suis conculcabat
DAN|7|20|et de cornibus decem quae habebat in capite et de alio quod ortum fuerat ante quod ceciderant tria cornua de cornu illo quod habebat oculos et os loquens grandia et maius erat ceteris
DAN|7|21|aspiciebam et ecce cornu illud faciebat bellum adversus sanctos et praevalebat eis
DAN|7|22|donec venit antiquus dierum et iudicium dedit sanctis Excelsi et tempus advenit et regnum obtinuerunt sancti
DAN|7|23|et sic ait bestia quarta regnum quartum erit in terra quod maius erit omnibus regnis et devorabit universam terram et conculcabit et comminuet eam
DAN|7|24|porro cornua decem ipsius regni decem reges erunt et alius consurget post eos et ipse potentior erit prioribus et tres reges humiliabit
DAN|7|25|et sermones contra Excelsum loquetur et sanctos Altissimi conteret et putabit quod possit mutare tempora et leges et tradentur in manu eius usque ad tempus et tempora et dimidium temporis
DAN|7|26|et iudicium sedebit ut auferatur potentia et conteratur et dispereat usque in finem
DAN|7|27|regnum autem et potestas et magnitudo regni quae est subter omne caelum detur populo sanctorum Altissimi cuius regnum regnum sempiternum est et omnes reges servient ei et oboedient
DAN|7|28|hucusque finis verbi ego Danihel multum cogitationibus meis conturbabar et facies mea mutata est in me verbum autem in corde meo conservavi
DAN|8|1|anno tertio regni Balthasar regis visio apparuit mihi ego Danihel post id quod videram in principio
DAN|8|2|vidi in visione mea cum essem in Susis castro quod est in Aelam civitate vidi autem in visione esse me super portam Ulai
DAN|8|3|et levavi oculos meos et vidi et ecce aries unus stabat ante paludem habens cornua excelsa et unum excelsius altero atque succrescens postea
DAN|8|4|vidi arietem cornibus ventilantem contra occidentem et contra aquilonem et contra meridiem et omnes bestiae non poterant resistere ei neque liberari de manu eius fecitque secundum voluntatem suam et magnificatus est
DAN|8|5|et ego intellegebam ecce autem hircus caprarum veniebat ab occidente super faciem totius terrae et non tangebat terram porro hircus habebat cornu insigne inter oculos suos
DAN|8|6|et venit usque ad arietem illum cornutum quem videram stantem ante portam et cucurrit ad eum in impetu fortitudinis suae
DAN|8|7|cumque adpropinquasset prope arietem efferatus est in eum et percussit arietem et comminuit duo cornua eius et non poterat aries resistere ei cumque eum misisset in terram conculcavit et nemo quibat liberare arietem de manu eius
DAN|8|8|hircus autem caprarum magnus factus est nimis cumque crevisset fractum est cornu magnum et orta sunt cornua quattuor subter illud per quattuor ventos caeli
DAN|8|9|de uno autem ex eis egressum est cornu unum modicum et factum est grande contra meridiem et contra orientem et contra fortitudinem
DAN|8|10|et magnificatum est usque ad fortitudinem caeli et deiecit de fortitudine et de stellis et conculcavit eas
DAN|8|11|et usque ad principem fortitudinis magnificatus est et ab eo tulit iuge sacrificium et deiecit locum sanctificationis eius
DAN|8|12|robur autem datum est contra iuge sacrificium propter peccata et prosternetur veritas in terra et faciet et prosperabitur
DAN|8|13|et audivi unum de sanctis loquentem et dixit unus sanctus alteri nescio cui loquenti usquequo visio et iuge sacrificium et peccatum desolationis quae facta est et sanctuarium et fortitudo conculcabitur
DAN|8|14|et dixit ei usque ad vesperam et mane duo milia trecenti et mundabitur sanctuarium
DAN|8|15|factum est autem cum viderem ego Danihel visionem et quaererem intellegentiam ecce stetit in conspectu meo quasi species viri
DAN|8|16|et audivi vocem viri inter Ulai et clamavit et ait Gabrihel fac intellegere istum visionem
DAN|8|17|et venit et stetit iuxta ubi ego stabam cumque venisset pavens corrui in faciem meam et ait ad me intellege fili hominis quoniam in tempore finis conplebitur visio
DAN|8|18|cumque loqueretur ad me conlapsus sum pronus in terram et tetigit me et statuit me in gradu meo
DAN|8|19|dixitque mihi ego ostendam tibi quae futura sint in novissimo maledictionis quoniam habet tempus finem suum
DAN|8|20|aries quem vidisti habere cornua rex Medorum est atque Persarum
DAN|8|21|porro hircus caprarum rex Graecorum est et cornu grande quod erat inter oculos eius ipse est rex primus
DAN|8|22|quod autem fracto illo surrexerunt quattuor pro eo quattuor reges de gente eius consurgent sed non in fortitudine eius
DAN|8|23|et post regnum eorum cum creverint iniquitates consurget rex inpudens facie et intellegens propositiones
DAN|8|24|et roborabitur fortitudo eius sed non in viribus suis et supra quam credi potest universa vastabit et prosperabitur et faciet et interficiet robustos et populum sanctorum
DAN|8|25|secundum voluntatem suam et dirigetur dolus in manu eius et cor suum magnificabit et in copia rerum omnium occidet plurimos et contra principem principum consurget et sine manu conteretur
DAN|8|26|et visio vespere et mane quae dicta est vera est tu ergo signa visionem quia post dies multos erit
DAN|8|27|et ego Danihel langui et aegrotavi per dies cumque surrexissem faciebam opera regis et stupebam ad visionem et non erat qui interpretaretur
DAN|9|1|in anno primo Darii filii Asueri de semine Medorum qui imperavit super regnum Chaldeorum
DAN|9|2|anno uno regni eius ego Danihel intellexi in libris numerum annorum de quo factus est sermo Domini ad Hieremiam prophetam ut conplerentur desolationes Hierusalem septuaginta anni
DAN|9|3|et posui faciem meam ad Dominum Deum rogare et deprecari in ieiuniis sacco et cinere
DAN|9|4|et oravi Dominum Deum meum et confessus sum et dixi obsecro Domine Deus magne et terribilis custodiens pactum et misericordiam diligentibus te et custodientibus mandata tua
DAN|9|5|peccavimus inique fecimus impie egimus et recessimus et declinavimus a mandatis tuis ac iudiciis
DAN|9|6|non oboedivimus servis tuis prophetis qui locuti sunt in nomine tuo regibus nostris principibus nostris patribus nostris omnique populo terrae
DAN|9|7|tibi Domine iustitia nobis autem confusio faciei sicut est hodie viro Iuda et habitatoribus Hierusalem et omni Israhel his qui prope sunt et his qui procul in universis terris ad quas eiecisti eos propter iniquitates eorum in quibus peccaverunt in te
DAN|9|8|Domine nobis confusio faciei regibus nostris principibus nostris et patribus nostris qui peccaverunt
DAN|9|9|tibi autem Domino Deo nostro misericordia et propitiatio quia recessimus a te
DAN|9|10|et non audivimus vocem Domini Dei nostri ut ambularemus in lege eius quam posuit nobis per servos suos prophetas
DAN|9|11|et omnis Israhel praevaricati sunt legem tuam et declinaverunt ne audirent vocem tuam et stillavit super nos maledictio et detestatio quae scripta est in libro Mosi servi Dei quia peccavimus ei
DAN|9|12|et statuit sermones suos quos locutus est super nos et super principes nostros qui iudicaverunt nos ut superducerent in nos malum magnum quale numquam fuit sub omni caelo secundum quod factum est in Hierusalem
DAN|9|13|sicut scriptum est in lege Mosi omne malum hoc venit super nos et non rogavimus faciem tuam Domine Deus noster ut reverteremur ab iniquitatibus nostris et cogitaremus veritatem tuam
DAN|9|14|et vigilavit Dominus et adduxit eam super nos iustus Dominus Deus noster in omnibus operibus suis quae fecit non enim audivimus vocem eius
DAN|9|15|et nunc Domine Deus noster qui eduxisti populum tuum de terra Aegypti in manu forti et fecisti tibi nomen secundum diem hanc peccavimus iniquitatem fecimus
DAN|9|16|Domine in omnem iustitiam tuam avertatur obsecro ira tua et furor tuus a civitate tua Hierusalem et monte sancto tuo propter peccata enim nostra et iniquitates patrum nostrorum Hierusalem et populus tuus in obprobrium sunt omnibus per circuitum nostrum
DAN|9|17|nunc ergo exaudi Deus noster orationem servi tui et preces eius et ostende faciem tuam super sanctuarium tuum quod desertum est propter temet ipsum
DAN|9|18|inclina Deus meus aurem tuam et audi aperi oculos tuos et vide desolationem nostram et civitatem super quam invocatum est nomen tuum neque enim in iustificationibus nostris prosternimus preces ante faciem tuam sed in miserationibus tuis multis
DAN|9|19|exaudi Domine placare Domine adtende et fac ne moreris propter temet ipsum Deus meus quia nomen tuum invocatum est super civitatem et super populum tuum
DAN|9|20|cumque adhuc loquerer et orarem et confiterer peccata mea et peccata populi mei Israhel ut prosternerem preces meas in conspectu Dei mei pro monte sancto Dei mei
DAN|9|21|adhuc me loquente in oratione ecce vir Gabrihel quem videram in visione principio cito volans tetigit me in tempore sacrificii vespertini
DAN|9|22|et docuit me et locutus est mihi dixitque Danihel nunc egressus sum ut docerem te et intellegeres
DAN|9|23|ab exordio precum tuarum egressus est sermo ego autem veni ut indicarem tibi quia vir desideriorum es tu ergo animadverte sermonem et intellege visionem
DAN|9|24|septuaginta ebdomades adbreviatae sunt super populum tuum et super urbem sanctam tuam ut consummetur praevaricatio et finem accipiat peccatum et deleatur iniquitas et adducatur iustitia sempiterna et impleatur visio et prophetes et unguatur sanctus sanctorum
DAN|9|25|scito ergo et animadverte ab exitu sermonis ut iterum aedificetur Hierusalem usque ad christum ducem ebdomades septem et ebdomades sexaginta duae erunt et rursum aedificabitur platea et muri in angustia temporum
DAN|9|26|et post ebdomades sexaginta duas occidetur christus et non erit eius et civitatem et sanctuarium dissipabit populus cum duce venturo et finis eius vastitas et post finem belli statuta desolatio
DAN|9|27|confirmabit autem pactum multis ebdomas una et in dimidio ebdomadis deficiet hostia et sacrificium et in templo erit abominatio desolationis et usque ad consummationem et finem perseverabit desolatio
DAN|10|1|anno tertio Cyri regis Persarum verbum revelatum est Daniheli cognomento Balthasar et verum verbum et fortitudo magna intellexitque sermonem intellegentia est enim opus in visione
DAN|10|2|in diebus illis ego Danihel lugebam trium ebdomadarum diebus
DAN|10|3|panem desiderabilem non comedi et caro et vinum non introierunt in os meum sed neque unguento unctus sum donec conplerentur trium ebdomadarum dies
DAN|10|4|die autem vicesima et quarta mensis primi eram iuxta fluvium magnum qui est Tigris
DAN|10|5|et levavi oculos meos et vidi et ecce vir unus vestitus lineis et renes eius accincti auro obrizo
DAN|10|6|et corpus eius quasi chrysolitus et facies eius velut species fulgoris et oculi eius ut lampas ardens et brachia eius et quae deorsum usque ad pedes quasi species aeris candentis et vox sermonum eius ut vox multitudinis
DAN|10|7|vidi autem ego Danihel solus visionem porro viri qui erant mecum non viderunt sed terror nimius inruit super eos et fugerunt in absconditum
DAN|10|8|ego autem relictus solus vidi visionem grandem hanc et non remansit in me fortitudo sed et species mea inmutata est in me et emarcui nec habui quicquam virium
DAN|10|9|et audivi vocem sermonum eius et audiens iacebam consternatus super faciem meam vultusque meus herebat terrae
DAN|10|10|et ecce manus tetigit me et erexit me super genua mea et super articulos manuum mearum
DAN|10|11|et dixit ad me Danihel vir desideriorum intellege verba quae ego loquor ad te et sta in gradu tuo nunc enim sum missus ad te cumque dixisset mihi sermonem istum steti tremens
DAN|10|12|et ait ad me noli metuere Danihel quia ex die primo quo posuisti cor tuum ad intellegendum ut te adfligeres in conspectu Dei tui exaudita sunt verba tua et ego veni propter sermones tuos
DAN|10|13|princeps autem regni Persarum restitit mihi viginti et uno diebus et ecce Michahel unus de principibus primis venit in adiutorium meum et ego remansi ibi iuxta regem Persarum
DAN|10|14|veni autem ut docerem te quae ventura sunt populo tuo in novissimis diebus quoniam adhuc visio in dies
DAN|10|15|cumque loqueretur mihi huiuscemodi verbis deieci vultum meum ad terram et tacui
DAN|10|16|et ecce quasi similitudo filii hominis tetigit labia mea et aperiens os meum locutus sum et dixi ad eum qui stabat contra me domine mi in visione tua dissolutae sunt conpages meae et nihil in me remansit virium
DAN|10|17|et quomodo poterit servus domini mei loqui cum domino meo nihil enim in me remansit virium sed et halitus meus intercluditur
DAN|10|18|rursum ergo tetigit me quasi visio hominis et confortavit me
DAN|10|19|et dixit noli timere vir desideriorum pax tibi confortare et esto robustus cumque loqueretur mecum convalui et dixi loquere domine mi quia confortasti me
DAN|10|20|et ait numquid scis quare venerim ad te et nunc revertar ut proelier adversum principem Persarum cum enim egrederer apparuit princeps Graecorum veniens
DAN|10|21|verumtamen adnuntiabo tibi quod expressum est in scriptura veritatis et nemo est adiutor meus in omnibus his nisi Michahel princeps vester
DAN|11|1|ego autem ab anno primo Darii Medi stabam ut confortaretur et roboraretur
DAN|11|2|et nunc veritatem adnuntiabo tibi ecce adhuc tres reges stabunt in Perside et quartus ditabitur opibus nimiis super omnes et cum invaluerit divitiis suis concitabit omnes adversum regnum Graeciae
DAN|11|3|surget vero rex fortis et dominabitur potestate multa et faciet quod placuerit ei
DAN|11|4|et cum steterit conteretur regnum eius et dividetur in quattuor ventos caeli sed non in posteros eius neque secundum potentiam illius qua dominatus est lacerabitur enim regnum eius etiam in externos exceptis his
DAN|11|5|et confortabitur rex austri et de principibus eius praevalebit super eum et dominabitur dicione multa enim dominatio eius
DAN|11|6|et post finem annorum foederabuntur filiaque regis austri veniet ad regem aquilonis facere amicitiam et non obtinebit fortitudinem brachii nec stabit semen eius et tradetur ipsa et qui adduxerunt eam adulescentes eius et qui confortabant eam in temporibus
DAN|11|7|et stabit de germine radicum eius plantatio et veniet cum exercitu et ingredietur provinciam regis aquilonis et abutetur eis et obtinebit
DAN|11|8|insuper et deos eorum et sculptilia vasa quoque pretiosa argenti et auri captiva ducet in Aegyptum ipse praevalebit adversum regem aquilonis
DAN|11|9|et intrabit in regnum rex austri et revertetur ad terram suam
DAN|11|10|filii autem eius provocabuntur et congregabunt multitudinem exercituum plurimorum et veniet properans et inundans et revertetur et concitabitur et congredietur cum robore eius
DAN|11|11|et provocatus rex austri egredietur et pugnabit adversum regem aquilonis et praeparabit multitudinem nimiam et dabitur multitudo in manu eius
DAN|11|12|et capiet multitudinem et exaltabitur cor eius et deiciet multa milia sed non praevalebit
DAN|11|13|convertetur enim rex aquilonis et praeparabit multitudinem multo maiorem quam prius et in fine temporum annorumque veniet properans cum exercitu magno et opibus nimiis
DAN|11|14|et in temporibus illis multi consurgent adversum regem austri filii quoque praevaricatorum populi tui extollentur ut impleant visionem et corruent
DAN|11|15|et veniet rex aquilonis et conportabit aggerem et capiet urbes munitissimas et brachia austri non sustinebunt et consurgent electi eius ad resistendum et non erit fortitudo
DAN|11|16|et faciet veniens super eum iuxta placitum suum et non erit qui stet contra faciem eius et stabit in terra inclita et consumetur in manu eius
DAN|11|17|et ponet faciem suam ut veniat ad tenendum universum regnum eius et recta faciet cum eo et filiam feminarum dabit ei ut evertat illud et non stabit nec illius erit
DAN|11|18|et convertet faciem suam ad insulas et capiet multas et cessare faciet principem obprobrii sui et obprobrium eius convertetur in eum
DAN|11|19|et convertet faciem suam ad imperium terrae suae et inpinget et corruet et non invenietur
DAN|11|20|et stabit in loco eius vilissimus et indignus decore regio et in paucis diebus conteretur non in furore nec in proelio
DAN|11|21|et stabit in loco eius despectus et non tribuetur ei honor regius et veniet clam et obtinebit regnum in fraudulentia
DAN|11|22|et brachia pugnantis expugnabuntur a facie eius et conterentur insuper et dux foederis
DAN|11|23|et post amicitias cum eo faciet dolum et ascendet et superabit in modico populo
DAN|11|24|abundantes et uberes urbes ingredietur et faciet quae non fecerunt patres eius et patres patrum eius rapinas et praedam et divitias eorum dissipabit et contra firmissimas cogitationes iniet et hoc usque ad tempus
DAN|11|25|et concitabitur fortitudo eius et cor eius adversum regem austri in exercitu magno et rex austri provocabitur ad bellum multis auxiliis et fortibus nimis et non stabunt quia inibunt adversum eum consilia
DAN|11|26|et comedentes panem cum eo conterent illum exercitusque eius opprimetur et cadent interfecti plurimi
DAN|11|27|duorum quoque regum cor erit ut malefaciant et ad mensam unam mendacium loquentur et non proficient quia adhuc finis in aliud tempus
DAN|11|28|et revertetur in terram suam cum opibus multis et cor eius adversus testamentum sanctum et faciet et revertetur in terram suam
DAN|11|29|statuto tempore revertetur et veniet ad austrum et non erit priori simile novissimum
DAN|11|30|et venient super eum trieres et Romani et percutietur et revertetur et indignabitur contra testamentum sanctuarii et faciet reverteturque et cogitabit adversum eos qui dereliquerunt testamentum sanctuarii
DAN|11|31|et brachia ex eo stabunt et polluent sanctuarium fortitudinis et auferent iuge sacrificium et dabunt abominationem in desolationem
DAN|11|32|et impii in testamentum simulabunt fraudulenter populus autem sciens Deum suum obtinebit et faciet
DAN|11|33|et docti in populo docebunt plurimos et ruent in gladio et in flamma in captivitate et rapina dierum
DAN|11|34|cumque corruerint sublevabuntur auxilio parvulo et adplicabuntur eis plurimi fraudulenter
DAN|11|35|et de eruditis ruent ut conflentur et eligantur et dealbentur usque ad tempus praefinitum quia adhuc aliud tempus erit
DAN|11|36|et faciet iuxta voluntatem suam rex et elevabitur et magnificabitur adversum omnem deum et adversum Deum deorum loquetur magnifica et diriget donec conpleatur iracundia perpetrata est quippe definitio
DAN|11|37|et Deum patrum suorum non reputabit et erit in concupiscentiis feminarum nec quemquam deorum curabit quia adversum universa consurget
DAN|11|38|deum autem Maozim in loco suo venerabitur et deum quem ignoraverunt patres eius colet auro et argento et lapide pretioso rebusque pretiosis
DAN|11|39|et faciet ut muniat Maozim cum deo alieno quem cognovit et multiplicabit gloriam et dabit eis potestatem in multis et terram dividet gratuito
DAN|11|40|et in tempore praefinito proeliabitur adversum eum rex austri et quasi tempestas veniet contra illum rex aquilonis in curribus et in equitibus et in classe magna et ingredietur terras et conteret et pertransiet
DAN|11|41|et introibit in terram gloriosam et multae corruent hae autem solae salvabuntur de manu eius Edom et Moab et principium filiorum Ammon
DAN|11|42|et mittet manum suam in terras et terra Aegypti non effugiet
DAN|11|43|et dominabitur thesaurorum auri et argenti et in omnibus pretiosis Aegypti per Lybias quoque et Aethiopias transibit
DAN|11|44|et fama turbabit eum ab oriente et ab aquilone et veniet in multitudine magna ut conterat et interficiat plurimos
DAN|11|45|et figet tabernaculum suum Apedno inter maria super montem inclitum et sanctum et veniet usque ad summitatem eius et nemo auxiliabitur ei
DAN|12|1|in tempore autem illo consurget Michahel princeps magnus qui stat pro filiis populi tui et veniet tempus quale non fuit ab eo quo gentes esse coeperunt usque ad tempus illud et in tempore illo salvabitur populus tuus omnis qui inventus fuerit scriptus in libro
DAN|12|2|et multi de his qui dormiunt in terrae pulvere evigilabunt alii in vitam aeternam et alii in obprobrium ut videant semper
DAN|12|3|qui autem docti fuerint fulgebunt quasi splendor firmamenti et qui ad iustitiam erudiunt multos quasi stellae in perpetuas aeternitates
DAN|12|4|tu autem Danihel clude sermones et signa librum usque ad tempus statutum pertransibunt plurimi et multiplex erit scientia
DAN|12|5|et vidi ego Danihel et ecce quasi duo alii stabant unus hinc super ripam fluminis et alius inde ex altera ripa fluminis
DAN|12|6|et dixi viro qui indutus erat lineis qui stabat super aquas fluminis usquequo finis horum mirabilium
DAN|12|7|et audivi virum qui indutus erat lineis qui stabat super aquas fluminis cum levasset dexteram et sinistram suam in caelum et iurasset per viventem in aeternum quia in tempus temporum et dimidium temporis et cum conpleta fuerit dispersio manus populi sancti conplebuntur universa haec
DAN|12|8|et ego audivi et non intellexi et dixi domine mi quid erit post haec
DAN|12|9|et ait vade Danihel quia clausi sunt signatique sermones usque ad tempus praefinitum
DAN|12|10|eligentur et dealbabuntur et quasi ignis probabuntur multi et impie agent impii neque intellegent omnes impii porro docti intellegent
DAN|12|11|et a tempore cum ablatum fuerit iuge sacrificium et posita fuerit abominatio in desolatione dies mille ducenti nonaginta
DAN|12|12|beatus qui expectat et pervenit ad dies mille trecentos triginta quinque
DAN|12|13|tu autem vade ad praefinitum et requiesce et stabis in sorte tua in fine dierum
