PROV|1|1|The proverbs of Solomon, son of David, king of Israel:
PROV|1|2|To know wisdom and instruction, to understand words of insight,
PROV|1|3|to receive instruction in wise dealing, in righteousness, justice, and equity;
PROV|1|4|to give prudence to the simple, knowledge and discretion to the youth-
PROV|1|5|Let the wise hear and increase in learning, and the one who understands obtain guidance,
PROV|1|6|to understand a proverb and a saying, the words of the wise and their riddles.
PROV|1|7|The fear of the LORD is the beginning of knowledge; fools despise wisdom and instruction.
PROV|1|8|Hear, my son, your father's instruction, and forsake not your mother's teaching,
PROV|1|9|for they are a graceful garland for your head and pendants for your neck.
PROV|1|10|My son, if sinners entice you, do not consent.
PROV|1|11|If they say, "Come with us, let us lie in wait for blood; let us ambush the innocent without reason;
PROV|1|12|like Sheol let us swallow them alive, and whole, like those who go down to the pit;
PROV|1|13|we shall find all precious goods, we shall fill our houses with plunder;
PROV|1|14|throw in your lot among us; we will all have one purse"-
PROV|1|15|my son, do not walk in the way with them; hold back your foot from their paths,
PROV|1|16|for their feet run to evil, and they make haste to shed blood.
PROV|1|17|For in vain is a net spread in the sight of any bird,
PROV|1|18|but these men lie in wait for their own blood; they set an ambush for their own lives.
PROV|1|19|Such are the ways of everyone who is greedy for unjust gain; it takes away the life of its possessors.
PROV|1|20|Wisdom cries aloud in the street, in the markets she raises her voice;
PROV|1|21|at the head of the noisy streets she cries out; at the entrance of the city gates she speaks:
PROV|1|22|"How long, O simple ones, will you love being simple? How long will scoffers delight in their scoffing and fools hate knowledge?
PROV|1|23|If you turn at my reproof, behold, I will pour out my spirit to you; I will make my words known to you.
PROV|1|24|Because I have called and you refused to listen, have stretched out my hand and no one has heeded,
PROV|1|25|because you have ignored all my counsel and would have none of my reproof,
PROV|1|26|I also will laugh at your calamity; I will mock when terror strikes you,
PROV|1|27|when terror strikes you like a storm and your calamity comes like a whirlwind, when distress and anguish come upon you.
PROV|1|28|Then they will call upon me, but I will not answer; they will seek me diligently but will not find me.
PROV|1|29|Because they hated knowledge and did not choose the fear of the LORD,
PROV|1|30|would have none of my counsel and despised all my reproof,
PROV|1|31|therefore they shall eat the fruit of their way, and have their fill of their own devices.
PROV|1|32|For the simple are killed by their turning away, and the complacency of fools destroys them;
PROV|1|33|but whoever listens to me will dwell secure and will be at ease, without dread of disaster."
PROV|2|1|My son, if you receive my words and treasure up my commandments with you,
PROV|2|2|making your ear attentive to wisdom and inclining your heart to understanding;
PROV|2|3|yes, if you call out for insight and raise your voice for understanding,
PROV|2|4|if you seek it like silver and search for it as for hidden treasures,
PROV|2|5|then you will understand the fear of the LORD and find the knowledge of God.
PROV|2|6|For the LORD gives wisdom; from his mouth come knowledge and understanding;
PROV|2|7|he stores up sound wisdom for the upright; he is a shield to those who walk in integrity,
PROV|2|8|guarding the paths of justice and watching over the way of his saints.
PROV|2|9|Then you will understand righteousness and justice and equity, every good path;
PROV|2|10|for wisdom will come into your heart, and knowledge will be pleasant to your soul;
PROV|2|11|discretion will watch over you, understanding will guard you,
PROV|2|12|delivering you from the way of evil, from men of perverted speech,
PROV|2|13|who forsake the paths of uprightness to walk in the ways of darkness,
PROV|2|14|who rejoice in doing evil and delight in the perverseness of evil,
PROV|2|15|men whose paths are crooked, and who are devious in their ways.
PROV|2|16|So you will be delivered from the forbidden woman, from the adulteress with her smooth words,
PROV|2|17|who forsakes the companion of her youth and forgets the covenant of her God;
PROV|2|18|for her house sinks down to death, and her paths to the departed;
PROV|2|19|none who go to her come back, nor do they regain the paths of life.
PROV|2|20|So you will walk in the way of the good and keep to the paths of the righteous.
PROV|2|21|For the upright will inhabit the land, and those with integrity will remain in it,
PROV|2|22|but the wicked will be cut off from the land, and the treacherous will be rooted out of it.
PROV|3|1|My son, do not forget my teaching, but let your heart keep my commandments,
PROV|3|2|for length of days and years of life and peace they will add to you.
PROV|3|3|Let not steadfast love and faithfulness forsake you; bind them around your neck; write them on the tablet of your heart.
PROV|3|4|So you will find favor and good success in the sight of God and man.
PROV|3|5|Trust in the LORD with all your heart, and do not lean on your own understanding.
PROV|3|6|In all your ways acknowledge him, and he will make straight your paths.
PROV|3|7|Be not wise in your own eyes; fear the LORD, and turn away from evil.
PROV|3|8|It will be healing to your flesh and refreshment to your bones.
PROV|3|9|Honor the LORD with your wealth and with the firstfruits of all your produce;
PROV|3|10|then your barns will be filled with plenty, and your vats will be bursting with wine.
PROV|3|11|My son, do not despise the LORD's discipline or be weary of his reproof,
PROV|3|12|for the LORD reproves him whom he loves, as a father the son in whom he delights.
PROV|3|13|Blessed is the one who finds wisdom, and the one who gets understanding,
PROV|3|14|for the gain from her is better than gain from silver and her profit better than gold.
PROV|3|15|She is more precious than jewels, and nothing you desire can compare with her.
PROV|3|16|Long life is in her right hand; in her left hand are riches and honor.
PROV|3|17|Her ways are ways of pleasantness, and all her paths are peace.
PROV|3|18|She is a tree of life to those who lay hold of her; those who hold her fast are called blessed.
PROV|3|19|The LORD by wisdom founded the earth; by understanding he established the heavens;
PROV|3|20|by his knowledge the deeps broke open, and the clouds drop down the dew.
PROV|3|21|My son, do not lose sight of these- keep sound wisdom and discretion,
PROV|3|22|and they will be life for your soul and adornment for your neck.
PROV|3|23|Then you will walk on your way securely, and your foot will not stumble.
PROV|3|24|If you lie down, you will not be afraid; when you lie down, your sleep will be sweet.
PROV|3|25|Do not be afraid of sudden terror or of the ruin of the wicked, when it comes,
PROV|3|26|for the LORD will be your confidence and will keep your foot from being caught.
PROV|3|27|Do not withhold good from those to whom it is due, when it is in your power to do it.
PROV|3|28|Do not say to your neighbor, "Go, and come again, tomorrow I will give it"- when you have it with you.
PROV|3|29|Do not plan evil against your neighbor, who dwells trustingly beside you.
PROV|3|30|Do not contend with a man for no reason, when he has done you no harm.
PROV|3|31|Do not envy a man of violence and do not choose any of his ways,
PROV|3|32|for the devious person is an abomination to the LORD, but the upright are in his confidence.
PROV|3|33|The LORD's curse is on the house of the wicked, but he blesses the dwelling of the righteous.
PROV|3|34|Toward the scorners he is scornful, but to the humble he gives favor.
PROV|3|35|The wise will inherit honor, but fools get disgrace.
PROV|4|1|Hear, O sons, a father's instruction, and be attentive, that you may gain insight,
PROV|4|2|for I give you good precepts; do not forsake my teaching.
PROV|4|3|When I was a son with my father, tender, the only one in the sight of my mother,
PROV|4|4|he taught me and said to me, "Let your heart hold fast my words; keep my commandments, and live.
PROV|4|5|Get wisdom; get insight; do not forget, and do not turn away from the words of my mouth.
PROV|4|6|Do not forsake her, and she will keep you; love her, and she will guard you.
PROV|4|7|The beginning of wisdom is this: Get wisdom, and whatever you get, get insight.
PROV|4|8|Prize her highly, and she will exalt you; she will honor you if you embrace her.
PROV|4|9|She will place on your head a graceful garland; she will bestow on you a beautiful crown."
PROV|4|10|Hear, my son, and accept my words, that the years of your life may be many.
PROV|4|11|I have taught you the way of wisdom; I have led you in the paths of uprightness.
PROV|4|12|When you walk, your step will not be hampered, and if you run, you will not stumble.
PROV|4|13|Keep hold of instruction; do not let go; guard her, for she is your life.
PROV|4|14|Do not enter the path of the wicked, and do not walk in the way of the evil.
PROV|4|15|Avoid it; do not go on it; turn away from it and pass on.
PROV|4|16|For they cannot sleep unless they have done wrong; they are robbed of sleep unless they have made someone stumble.
PROV|4|17|For they eat the bread of wickedness and drink the wine of violence.
PROV|4|18|But the path of the righteous is like the light of dawn, which shines brighter and brighter until full day.
PROV|4|19|The way of the wicked is like deep darkness; they do not know over what they stumble.
PROV|4|20|My son, be attentive to my words; incline your ear to my sayings.
PROV|4|21|Let them not escape from your sight; keep them within your heart.
PROV|4|22|For they are life to those who find them, and healing to all their flesh.
PROV|4|23|Keep your heart with all vigilance, for from it flow the springs of life.
PROV|4|24|Put away from you crooked speech, and put devious talk far from you.
PROV|4|25|Let your eyes look directly forward, and your gaze be straight before you.
PROV|4|26|Ponder the path of your feet; then all your ways will be sure.
PROV|4|27|Do not swerve to the right or to the left; turn your foot away from evil.
PROV|5|1|My son, be attentive to my wisdom; incline your ear to my understanding,
PROV|5|2|that you may keep discretion, and your lips may guard knowledge.
PROV|5|3|For the lips of a forbidden woman drip honey, and her speech is smoother than oil,
PROV|5|4|but in the end she is bitter as wormwood, sharp as a two-edged sword.
PROV|5|5|Her feet go down to death; her steps follow the path to Sheol;
PROV|5|6|she does not ponder the path of life; her ways wander, and she does not know it.
PROV|5|7|And now, O sons, listen to me, and do not depart from the words of my mouth.
PROV|5|8|Keep your way far from her, and do not go near the door of her house,
PROV|5|9|lest you give your honor to others and your years to the merciless,
PROV|5|10|lest strangers take their fill of your strength, and your labors go to the house of a foreigner,
PROV|5|11|and at the end of your life you groan, when your flesh and body are consumed,
PROV|5|12|and you say, "How I hated discipline, and my heart despised reproof!
PROV|5|13|I did not listen to the voice of my teachers or incline my ear to my instructors.
PROV|5|14|I am at the brink of utter ruin in the assembled congregation."
PROV|5|15|Drink water from your own cistern, flowing water from your own well.
PROV|5|16|Should your springs be scattered abroad, streams of water in the streets?
PROV|5|17|Let them be for yourself alone, and not for strangers with you.
PROV|5|18|Let your fountain be blessed, and rejoice in the wife of your youth,
PROV|5|19|a lovely deer, a graceful doe. Let her breasts fill you at all times with delight; be intoxicated always in her love.
PROV|5|20|Why should you be intoxicated, my son, with a forbidden woman and embrace the bosom of an adulteress?
PROV|5|21|For a man's ways are before the eyes of the LORD, and he ponders all his paths.
PROV|5|22|The iniquities of the wicked ensnare him, and he is held fast in the cords of his sin.
PROV|5|23|He dies for lack of discipline, and because of his great folly he is led astray.
PROV|6|1|My son, if you have put up security for your neighbor, have given your pledge for a stranger,
PROV|6|2|if you are snared in the words of your mouth, caught in the words of your mouth,
PROV|6|3|then do this, my son, and save yourself, for you have come into the hand of your neighbor: go, hasten, and plead urgently with your neighbor.
PROV|6|4|Give your eyes no sleep and your eyelids no slumber;
PROV|6|5|save yourself like a gazelle from the hand of the hunter, like a bird from the hand of the fowler.
PROV|6|6|Go to the ant, O sluggard; consider her ways, and be wise.
PROV|6|7|Without having any chief, officer, or ruler,
PROV|6|8|she prepares her bread in summer and gathers her food in harvest.
PROV|6|9|How long will you lie there, O sluggard? When will you arise from your sleep?
PROV|6|10|A little sleep, a little slumber, a little folding of the hands to rest,
PROV|6|11|and poverty will come upon you like a robber, and want like an armed man.
PROV|6|12|A worthless person, a wicked man, goes about with crooked speech,
PROV|6|13|winks with his eyes, signals with his feet, points with his finger,
PROV|6|14|with perverted heart devises evil, continually sowing discord;
PROV|6|15|therefore calamity will come upon him suddenly; in a moment he will be broken beyond healing.
PROV|6|16|There are six things that the LORD hates, seven that are an abomination to him:
PROV|6|17|haughty eyes, a lying tongue, and hands that shed innocent blood,
PROV|6|18|a heart that devises wicked plans, feet that make haste to run to evil,
PROV|6|19|a false witness who breathes out lies, and one who sows discord among brothers.
PROV|6|20|My son, keep your father's commandment, and forsake not your mother's teaching.
PROV|6|21|Bind them on your heart always; tie them around your neck.
PROV|6|22|When you walk, they will lead you; when you lie down, they will watch over you; and when you awake, they will talk with you.
PROV|6|23|For the commandment is a lamp and the teaching a light, and the reproofs of discipline are the way of life,
PROV|6|24|to preserve you from the evil woman, from the smooth tongue of the adulteress.
PROV|6|25|Do not desire her beauty in your heart, and do not let her capture you with her eyelashes;
PROV|6|26|for the price of a prostitute is only a loaf of bread, but a married woman hunts down a precious life.
PROV|6|27|Can a man carry fire next to his chest and his clothes not be burned?
PROV|6|28|Or can one walk on hot coals and his feet not be scorched?
PROV|6|29|So is he who goes in to his neighbor's wife; none who touches her will go unpunished.
PROV|6|30|People do not despise a thief if he steals to satisfy his appetite when he is hungry,
PROV|6|31|but if he is caught, he will pay sevenfold; he will give all the goods of his house.
PROV|6|32|He who commits adultery lacks sense; he who does it destroys himself.
PROV|6|33|Wounds and dishonor will he get, and his disgrace will not be wiped away.
PROV|6|34|For jealousy makes a man furious, and he will not spare when he takes revenge.
PROV|6|35|He will accept no compensation; he will refuse though you multiply gifts.
PROV|7|1|My son, keep my wordsand treasure up my commandments with you;
PROV|7|2|keep my commandments and live; keep my teaching as the apple of your eye;
PROV|7|3|bind them on your fingers; write them on the tablet of your heart.
PROV|7|4|Say to wisdom, "You are my sister," and call insight your intimate friend,
PROV|7|5|to keep you from the forbidden woman, from the adulteress with her smooth words.
PROV|7|6|For at the window of my house I have looked out through my lattice,
PROV|7|7|and I have seen among the simple, I have perceived among the youths, a young man lacking sense,
PROV|7|8|passing along the street near her corner, taking the road to her house
PROV|7|9|in the twilight, in the evening, at the time of night and darkness.
PROV|7|10|And behold, the woman meets him, dressed as a prostitute, wily of heart.
PROV|7|11|She is loud and wayward; her feet do not stay at home;
PROV|7|12|now in the street, now in the market, and at every corner she lies in wait.
PROV|7|13|She seizes him and kisses him, and with bold face she says to him,
PROV|7|14|"I had to offer sacrifices, and today I have paid my vows;
PROV|7|15|so now I have come out to meet you, to seek you eagerly, and I have found you.
PROV|7|16|I have spread my couch with coverings, colored linens from Egyptian linen;
PROV|7|17|I have perfumed my bed with myrrh, aloes, and cinnamon.
PROV|7|18|Come, let us take our fill of love till morning; let us delight ourselves with love.
PROV|7|19|For my husband is not at home; he has gone on a long journey;
PROV|7|20|he took a bag of money with him; at full moon he will come home."
PROV|7|21|With much seductive speech she persuades him; with her smooth talk she compels him.
PROV|7|22|All at once he follows her, as an ox goes to the slaughter, or as a stag is caught fast
PROV|7|23|till an arrow pierces its liver; as a bird rushes into a snare; he does not know that it will cost him his life.
PROV|7|24|And now, O sons, listen to me, and be attentive to the words of my mouth.
PROV|7|25|Let not your heart turn aside to her ways; do not stray into her paths,
PROV|7|26|for many a victim has she laid low, and all her slain are a mighty throng.
PROV|7|27|Her house is the way to Sheol, going down to the chambers of death.
PROV|8|1|Does not wisdom call?Does not understanding raise her voice?
PROV|8|2|On the heights beside the way, at the crossroads she takes her stand;
PROV|8|3|beside the gates in front of the town, at the entrance of the portals she cries aloud:
PROV|8|4|"To you, O men, I call, and my cry is to the children of man.
PROV|8|5|O simple ones, learn prudence; O fools, learn sense.
PROV|8|6|Hear, for I will speak noble things, and from my lips will come what is right,
PROV|8|7|for my mouth will utter truth; wickedness is an abomination to my lips.
PROV|8|8|All the words of my mouth are righteous; there is nothing twisted or crooked in them.
PROV|8|9|They are all straight to him who understands, and right to those who find knowledge.
PROV|8|10|Take my instruction instead of silver, and knowledge rather than choice gold,
PROV|8|11|for wisdom is better than jewels, and all that you may desire cannot compare with her.
PROV|8|12|"I, wisdom, dwell with prudence, and I find knowledge and discretion.
PROV|8|13|The fear of the LORD is hatred of evil. Pride and arrogance and the way of evil and perverted speech I hate.
PROV|8|14|I have counsel and sound wisdom; I have insight; I have strength.
PROV|8|15|By me kings reign, and rulers decree what is just;
PROV|8|16|by me princes rule, and nobles, all who govern justly.
PROV|8|17|I love those who love me, and those who seek me diligently find me.
PROV|8|18|Riches and honor are with me, enduring wealth and righteousness.
PROV|8|19|My fruit is better than gold, even fine gold, and my yield than choice silver.
PROV|8|20|I walk in the way of righteousness, in the paths of justice,
PROV|8|21|granting an inheritance to those who love me, and filling their treasuries.
PROV|8|22|"The LORD possessed me at the beginning of his work, the first of his acts of old.
PROV|8|23|Ages ago I was set up, at the first, before the beginning of the earth.
PROV|8|24|When there were no depths I was brought forth, when there were no springs abounding with water.
PROV|8|25|Before the mountains had been shaped, before the hills, I was brought forth,
PROV|8|26|before he had made the earth with its fields, or the first of the dust of the world.
PROV|8|27|When he established the heavens, I was there; when he drew a circle on the face of the deep,
PROV|8|28|when he made firm the skies above, when he established the fountains of the deep,
PROV|8|29|when he assigned to the sea its limit, so that the waters might not transgress his command, when he marked out the foundations of the earth,
PROV|8|30|then I was beside him, like a master workman, and I was daily his delight, rejoicing before him always,
PROV|8|31|rejoicing in his inhabited world and delighting in the children of man.
PROV|8|32|"And now, O sons, listen to me: blessed are those who keep my ways.
PROV|8|33|Hear instruction and be wise, and do not neglect it.
PROV|8|34|Blessed is the one who listens to me, watching daily at my gates, waiting beside my doors.
PROV|8|35|For whoever finds me finds life and obtains favor from the LORD,
PROV|8|36|but he who fails to find me injures himself; all who hate me love death."
PROV|9|1|Wisdom has built her house;she has hewn her seven pillars.
PROV|9|2|She has slaughtered her beasts; she has mixed her wine; she has also set her table.
PROV|9|3|She has sent out her young women to call from the highest places in the town,
PROV|9|4|"Whoever is simple, let him turn in here!" To him who lacks sense she says,
PROV|9|5|"Come, eat of my bread and drink of the wine I have mixed.
PROV|9|6|Leave your simple ways, and live, and walk in the way of insight."
PROV|9|7|Whoever corrects a scoffer gets himself abuse, and he who reproves a wicked man incurs injury.
PROV|9|8|Do not reprove a scoffer, or he will hate you; reprove a wise man, and he will love you.
PROV|9|9|Give instruction to a wise man, and he will be still wiser; teach a righteous man, and he will increase in learning.
PROV|9|10|The fear of the LORD is the beginning of wisdom, and the knowledge of the Holy One is insight.
PROV|9|11|For by me your days will be multiplied, and years will be added to your life.
PROV|9|12|If you are wise, you are wise for yourself; if you scoff, you alone will bear it.
PROV|9|13|The woman Folly is loud; she is seductive and knows nothing.
PROV|9|14|She sits at the door of her house; she takes a seat on the highest places of the town,
PROV|9|15|calling to those who pass by, who are going straight on their way,
PROV|9|16|"Whoever is simple, let him turn in here!" And to him who lacks sense she says,
PROV|9|17|"Stolen water is sweet, and bread eaten in secret is pleasant."
PROV|9|18|But he does not know that the dead are there, that her guests are in the depths of Sheol.
PROV|10|1|The proverbs of Solomon. A wise son makes a glad father, but a foolish son is a sorrow to his mother.
PROV|10|2|Treasures gained by wickedness do not profit, but righteousness delivers from death.
PROV|10|3|The LORD does not let the righteous go hungry, but he thwarts the craving of the wicked.
PROV|10|4|A slack hand causes poverty, but the hand of the diligent makes rich.
PROV|10|5|He who gathers in summer is a prudent son, but he who sleeps in harvest is a son who brings shame.
PROV|10|6|Blessings are on the head of the righteous, but the mouth of the wicked conceals violence.
PROV|10|7|The memory of the righteous is a blessing, but the name of the wicked will rot.
PROV|10|8|The wise of heart will receive commandments, but a babbling fool will come to ruin.
PROV|10|9|Whoever walks in integrity walks securely, but he who makes his ways crooked will be found out.
PROV|10|10|Whoever winks the eye causes trouble, but a babbling fool will come to ruin.
PROV|10|11|The mouth of the righteous is a fountain of life, but the mouth of the wicked conceals violence.
PROV|10|12|Hatred stirs up strife, but love covers all offenses.
PROV|10|13|On the lips of him who has understanding, wisdom is found, but a rod is for the back of him who lacks sense.
PROV|10|14|The wise lay up knowledge, but the mouth of a fool brings ruin near.
PROV|10|15|A rich man's wealth is his strong city; the poverty of the poor is their ruin.
PROV|10|16|The wage of the righteous leads to life, the gain of the wicked to sin.
PROV|10|17|Whoever heeds instruction is on the path to life, but he who rejects reproof leads others astray.
PROV|10|18|The one who conceals hatred has lying lips, and whoever utters slander is a fool.
PROV|10|19|When words are many, transgression is not lacking, but whoever restrains his lips is prudent.
PROV|10|20|The tongue of the righteous is choice silver; the heart of the wicked is of little worth.
PROV|10|21|The lips of the righteous feed many, but fools die for lack of sense.
PROV|10|22|The blessing of the LORD makes rich, and he adds no sorrow with it.
PROV|10|23|Doing wrong is like a joke to a fool, but wisdom is pleasure to a man of understanding.
PROV|10|24|What the wicked dreads will come upon him, but the desire of the righteous will be granted.
PROV|10|25|When the tempest passes, the wicked is no more, but the righteous is established forever.
PROV|10|26|Like vinegar to the teeth and smoke to the eyes, so is the sluggard to those who send him.
PROV|10|27|The fear of the LORD prolongs life, but the years of the wicked will be short.
PROV|10|28|The hope of the righteous brings joy, but the expectation of the wicked will perish.
PROV|10|29|The way of the LORD is a stronghold to the blameless, but destruction to evildoers.
PROV|10|30|The righteous will never be removed, but the wicked will not dwell in the land.
PROV|10|31|The mouth of the righteous brings forth wisdom, but the perverse tongue will be cut off.
PROV|10|32|The lips of the righteous know what is acceptable, but the mouth of the wicked, what is perverse.
PROV|11|1|A false balance is an abomination to the LORD, but a just weight is his delight.
PROV|11|2|When pride comes, then comes disgrace, but with the humble is wisdom.
PROV|11|3|The integrity of the upright guides them, but the crookedness of the treacherous destroys them.
PROV|11|4|Riches do not profit in the day of wrath, but righteousness delivers from death.
PROV|11|5|The righteousness of the blameless keeps his way straight, but the wicked falls by his own wickedness.
PROV|11|6|The righteousness of the upright delivers them, but the treacherous are taken captive by their lust.
PROV|11|7|When the wicked dies, his hope will perish, and the expectation of wealth perishes too.
PROV|11|8|The righteous is delivered from trouble, and the wicked walks into it instead.
PROV|11|9|With his mouth the godless man would destroy his neighbor, but by knowledge the righteous are delivered.
PROV|11|10|When it goes well with the righteous, the city rejoices, and when the wicked perish there are shouts of gladness.
PROV|11|11|By the blessing of the upright a city is exalted, but by the mouth of the wicked it is overthrown.
PROV|11|12|Whoever belittles his neighbor lacks sense, but a man of understanding remains silent.
PROV|11|13|Whoever goes about slandering reveals secrets, but he who is trustworthy in spirit keeps a thing covered.
PROV|11|14|Where there is no guidance, a people falls, but in an abundance of counselors there is safety.
PROV|11|15|Whoever puts up security for a stranger will surely suffer harm, but he who hates striking hands in pledge is secure.
PROV|11|16|A gracious woman gets honor, and violent men get riches.
PROV|11|17|A man who is kind benefits himself, but a cruel man hurts himself.
PROV|11|18|The wicked earns deceptive wages, but one who sows righteousness gets a sure reward.
PROV|11|19|Whoever is steadfast in righteousness will live, but he who pursues evil will die.
PROV|11|20|Those of crooked heart are an abomination to the LORD, but those of blameless ways are his delight.
PROV|11|21|Be assured, an evil person will not go unpunished, but the offspring of the righteous will be delivered.
PROV|11|22|Like a gold ring in a pig's snout is a beautiful woman without discretion.
PROV|11|23|The desire of the righteous ends only in good; the expectation of the wicked in wrath.
PROV|11|24|One gives freely, yet grows all the richer; another withholds what he should give, and only suffers want.
PROV|11|25|Whoever brings blessing will be enriched, and one who waters will himself be watered.
PROV|11|26|The people curse him who holds back grain, but a blessing is on the head of him who sells it.
PROV|11|27|Whoever diligently seeks good seeks favor, but evil comes to him who searches for it.
PROV|11|28|Whoever trusts in his riches will fall, but the righteous will flourish like a green leaf.
PROV|11|29|Whoever troubles his own household will inherit the wind, and the fool will be servant to the wise of heart.
PROV|11|30|The fruit of the righteous is a tree of life, and whoever captures souls is wise.
PROV|11|31|If the righteous is repaid on earth, how much more the wicked and the sinner!
PROV|12|1|Whoever loves discipline loves knowledge, but he who hates reproof is stupid.
PROV|12|2|A good man obtains favor from the LORD, but a man of evil devices he condemns.
PROV|12|3|No one is established by wickedness, but the root of the righteous will never be moved.
PROV|12|4|An excellent wife is the crown of her husband, but she who brings shame is like rottenness in his bones.
PROV|12|5|The thoughts of the righteous are just; the counsels of the wicked are deceitful.
PROV|12|6|The words of the wicked lie in wait for blood, but the mouth of the upright delivers them.
PROV|12|7|The wicked are overthrown and are no more, but the house of the righteous will stand.
PROV|12|8|A man is commended according to his good sense, but one of twisted mind is despised.
PROV|12|9|Better to be lowly and have a servant than to play the great man and lack bread.
PROV|12|10|Whoever is righteous has regard for the life of his beast, but the mercy of the wicked is cruel.
PROV|12|11|Whoever works his land will have plenty of bread, but he who follows worthless pursuits lacks sense.
PROV|12|12|Whoever is wicked covets the spoil of evildoers, but the root of the righteous bears fruit.
PROV|12|13|An evil man is ensnared by the transgression of his lips, but the righteous escapes from trouble.
PROV|12|14|From the fruit of his mouth a man is satisfied with good, and the work of a man's hand comes back to him.
PROV|12|15|The way of a fool is right in his own eyes, but a wise man listens to advice.
PROV|12|16|The vexation of a fool is known at once, but the prudent ignores an insult.
PROV|12|17|Whoever speaks the truth gives honest evidence, but a false witness utters deceit.
PROV|12|18|There is one whose rash words are like sword thrusts, but the tongue of the wise brings healing.
PROV|12|19|Truthful lips endure forever, but a lying tongue is but for a moment.
PROV|12|20|Deceit is in the heart of those who devise evil, but those who plan peace have joy.
PROV|12|21|No ill befalls the righteous, but the wicked are filled with trouble.
PROV|12|22|Lying lips are an abomination to the LORD, but those who act faithfully are his delight.
PROV|12|23|A prudent man conceals knowledge, but the heart of fools proclaims folly.
PROV|12|24|The hand of the diligent will rule, while the slothful will be put to forced labor.
PROV|12|25|Anxiety in a man's heart weighs him down, but a good word makes him glad.
PROV|12|26|One who is righteous is a guide to his neighbor, but the way of the wicked leads them astray.
PROV|12|27|Whoever is slothful will not roast his game, but the diligent man will get precious wealth.
PROV|12|28|In the path of righteousness is life, and in its pathway there is no death.
PROV|13|1|A wise son hears his father's instruction, but a scoffer does not listen to rebuke.
PROV|13|2|From the fruit of his mouth a man eats what is good, but the desire of the treacherous is for violence.
PROV|13|3|Whoever guards his mouth preserves his life; he who opens wide his lips comes to ruin.
PROV|13|4|The soul of the sluggard craves and gets nothing, while the soul of the diligent is richly supplied.
PROV|13|5|The righteous hates falsehood, but the wicked brings shame and disgrace.
PROV|13|6|Righteousness guards him whose way is blameless, but sin overthrows the wicked.
PROV|13|7|One pretends to be rich, yet has nothing; another pretends to be poor, yet has great wealth.
PROV|13|8|The ransom of a man's life is his wealth, but a poor man hears no threat.
PROV|13|9|The light of the righteous rejoices, but the lamp of the wicked will be put out.
PROV|13|10|By insolence comes nothing but strife, but with those who take advice is wisdom.
PROV|13|11|Wealth gained hastily will dwindle, but whoever gathers little by little will increase it.
PROV|13|12|Hope deferred makes the heart sick, but a desire fulfilled is a tree of life.
PROV|13|13|Whoever despises the word brings destruction on himself, but he who reveres the commandment will be rewarded.
PROV|13|14|The teaching of the wise is a fountain of life, that one may turn away from the snares of death.
PROV|13|15|Good sense wins favor, but the way of the treacherous is their ruin.
PROV|13|16|In everything the prudent acts with knowledge, but a fool flaunts his folly.
PROV|13|17|A wicked messenger falls into trouble, but a faithful envoy brings healing.
PROV|13|18|Poverty and disgrace come to him who ignores instruction, but whoever heeds reproof is honored.
PROV|13|19|A desire fulfilled is sweet to the soul, but to turn away from evil is an abomination to fools.
PROV|13|20|Whoever walks with the wise becomes wise, but the companion of fools will suffer harm.
PROV|13|21|Disaster pursues sinners, but the righteous are rewarded with good.
PROV|13|22|A good man leaves an inheritance to his children's children, but the sinner's wealth is laid up for the righteous.
PROV|13|23|The fallow ground of the poor would yield much food, but it is swept away through injustice.
PROV|13|24|Whoever spares the rod hates his son, but he who loves him is diligent to discipline him.
PROV|13|25|The righteous has enough to satisfy his appetite, but the belly of the wicked suffers want.
PROV|14|1|The wisest of women builds her house, but folly with her own hands tears it down.
PROV|14|2|Whoever walks in uprightness fears the LORD, but he who is devious in his ways despises him.
PROV|14|3|By the mouth of a fool comes a rod for his back, but the lips of the wise will preserve them.
PROV|14|4|Where there are no oxen, the manger is clean, but abundant crops come by the strength of the ox.
PROV|14|5|A faithful witness does not lie, but a false witness breathes out lies.
PROV|14|6|A scoffer seeks wisdom in vain, but knowledge is easy for a man of understanding.
PROV|14|7|Leave the presence of a fool, for there you do not meet words of knowledge.
PROV|14|8|The wisdom of the prudent is to discern his way, but the folly of fools is deceiving.
PROV|14|9|Fools mock at the guilt offering, but the upright enjoy acceptance.
PROV|14|10|The heart knows its own bitterness, and no stranger shares its joy.
PROV|14|11|The house of the wicked will be destroyed, but the tent of the upright will flourish.
PROV|14|12|There is a way that seems right to a man, but its end is the way to death.
PROV|14|13|Even in laughter the heart may ache, and the end of joy may be grief.
PROV|14|14|The backslider in heart will be filled with the fruit of his ways, and a good man will be filled with the fruit of his ways.
PROV|14|15|The simple believes everything, but the prudent gives thought to his steps.
PROV|14|16|One who is wise is cautious and turns away from evil, but a fool is reckless and careless.
PROV|14|17|A man of quick temper acts foolishly, and a man of evil devices is hated.
PROV|14|18|The simple inherit folly, but the prudent are crowned with knowledge.
PROV|14|19|The evil bow down before the good, the wicked at the gates of the righteous.
PROV|14|20|The poor is disliked even by his neighbor, but the rich has many friends.
PROV|14|21|Whoever despises his neighbor is a sinner, but blessed is he who is generous to the poor.
PROV|14|22|Do they not go astray who devise evil? Those who devise good meet steadfast love and faithfulness.
PROV|14|23|In all toil there is profit, but mere talk tends only to poverty.
PROV|14|24|The crown of the wise is their wealth, but the folly of fools brings folly.
PROV|14|25|A truthful witness saves lives, but one who breathes out lies is deceitful.
PROV|14|26|In the fear of the LORD one has strong confidence, and his children will have a refuge.
PROV|14|27|The fear of the LORD is a fountain of life, that one may turn away from the snares of death.
PROV|14|28|In a multitude of people is the glory of a king, but without people a prince is ruined.
PROV|14|29|Whoever is slow to anger has great understanding, but he who has a hasty temper exalts folly.
PROV|14|30|A tranquil heart gives life to the flesh, but envy makes the bones rot.
PROV|14|31|Whoever oppresses a poor man insults his Maker, but he who is generous to the needy honors him.
PROV|14|32|The wicked is overthrown through his evildoing, but the righteous finds refuge in his death.
PROV|14|33|Wisdom rests in the heart of a man of understanding, but it makes itself known even in the midst of fools.
PROV|14|34|Righteousness exalts a nation, but sin is a reproach to any people.
PROV|14|35|A servant who deals wisely has the king's favor, but his wrath falls on one who acts shamefully.
PROV|15|1|A soft answer turns away wrath, but a harsh word stirs up anger.
PROV|15|2|The tongue of the wise commends knowledge, but the mouths of fools pour out folly.
PROV|15|3|The eyes of the LORD are in every place, keeping watch on the evil and the good.
PROV|15|4|A gentle tongue is a tree of life, but perverseness in it breaks the spirit.
PROV|15|5|A fool despises his father's instruction, but whoever heeds reproof is prudent.
PROV|15|6|In the house of the righteous there is much treasure, but trouble befalls the income of the wicked.
PROV|15|7|The lips of the wise spread knowledge; not so the hearts of fools.
PROV|15|8|The sacrifice of the wicked is an abomination to the LORD, but the prayer of the upright is acceptable to him.
PROV|15|9|The way of the wicked is an abomination to the LORD, but he loves him who pursues righteousness.
PROV|15|10|There is severe discipline for him who forsakes the way; whoever hates reproof will die.
PROV|15|11|Sheol and Abaddon lie open before the LORD; how much more the hearts of the children of man!
PROV|15|12|A scoffer does not like to be reproved; he will not go to the wise.
PROV|15|13|A glad heart makes a cheerful face, but by sorrow of heart the spirit is crushed.
PROV|15|14|The heart of him who has understanding seeks knowledge, but the mouths of fools feed on folly.
PROV|15|15|All the days of the afflicted are evil, but the cheerful of heart has a continual feast.
PROV|15|16|Better is a little with the fear of the LORD than great treasure and trouble with it.
PROV|15|17|Better is a dinner of herbs where love is than a fattened ox and hatred with it.
PROV|15|18|A hot-tempered man stirs up strife, but he who is slow to anger quiets contention.
PROV|15|19|The way of a sluggard is like a hedge of thorns, but the path of the upright is a level highway.
PROV|15|20|A wise son makes a glad father, but a foolish man despises his mother.
PROV|15|21|Folly is a joy to him who lacks sense, but a man of understanding walks straight ahead.
PROV|15|22|Without counsel plans fail, but with many advisers they succeed.
PROV|15|23|To make an apt answer is a joy to a man, and a word in season, how good it is!
PROV|15|24|The path of life leads upward for the prudent, that he may turn away from Sheol beneath.
PROV|15|25|The LORD tears down the house of the proud but maintains the widow's boundaries.
PROV|15|26|The thoughts of the wicked are an abomination to the LORD, but gracious words are pure.
PROV|15|27|Whoever is greedy for unjust gain troubles his own household, but he who hates bribes will live.
PROV|15|28|The heart of the righteous ponders how to answer, but the mouth of the wicked pours out evil things.
PROV|15|29|The LORD is far from the wicked, but he hears the prayer of the righteous.
PROV|15|30|The light of the eyes rejoices the heart, and good news refreshes the bones.
PROV|15|31|The ear that listens to life-giving reproof will dwell among the wise.
PROV|15|32|Whoever ignores instruction despises himself, but he who listens to reproof gains intelligence.
PROV|15|33|The fear of the LORD is instruction in wisdom, and humility comes before honor.
PROV|16|1|The plans of the heart belong to man, but the answer of the tongue is from the LORD.
PROV|16|2|All the ways of a man are pure in his own eyes, but the LORD weighs the spirit.
PROV|16|3|Commit your work to the LORD, and your plans will be established.
PROV|16|4|The LORD has made everything for its purpose, even the wicked for the day of trouble.
PROV|16|5|Everyone who is arrogant in heart is an abomination to the LORD; be assured, he will not go unpunished.
PROV|16|6|By steadfast love and faithfulness iniquity is atoned for, and by the fear of the LORD one turns away from evil.
PROV|16|7|When a man's ways please the LORD, he makes even his enemies to be at peace with him.
PROV|16|8|Better is a little with righteousness than great revenues with injustice.
PROV|16|9|The heart of man plans his way, but the LORD establishes his steps.
PROV|16|10|An oracle is on the lips of a king; his mouth does not sin in judgment.
PROV|16|11|A just balance and scales are the LORD's; all the weights in the bag are his work.
PROV|16|12|It is an abomination to kings to do evil, for the throne is established by righteousness.
PROV|16|13|Righteous lips are the delight of a king, and he loves him who speaks what is right.
PROV|16|14|A king's wrath is a messenger of death, and a wise man will appease it.
PROV|16|15|In the light of a king's face there is life, and his favor is like the clouds that bring the spring rain.
PROV|16|16|How much better to get wisdom than gold! To get understanding is to be chosen rather than silver.
PROV|16|17|The highway of the upright turns aside from evil; whoever guards his way preserves his life.
PROV|16|18|Pride goes before destruction, and a haughty spirit before a fall.
PROV|16|19|It is better to be of a lowly spirit with the poor than to divide the spoil with the proud.
PROV|16|20|Whoever gives thought to the word will discover good, and blessed is he who trusts in the LORD.
PROV|16|21|The wise of heart is called discerning, and sweetness of speech increases persuasiveness.
PROV|16|22|Good sense is a fountain of life to him who has it, but the instruction of fools is folly.
PROV|16|23|The heart of the wise makes his speech judicious and adds persuasiveness to his lips.
PROV|16|24|Gracious words are like a honeycomb, sweetness to the soul and health to the body.
PROV|16|25|There is a way that seems right to a man, but its end is the way to death.
PROV|16|26|A worker's appetite works for him; his mouth urges him on.
PROV|16|27|A worthless man plots evil, and his speech is like a scorching fire.
PROV|16|28|A dishonest man spreads strife, and a whisperer separates close friends.
PROV|16|29|A man of violence entices his neighbor and leads him in a way that is not good.
PROV|16|30|Whoever winks his eyes plans dishonest things; he who purses his lips brings evil to pass.
PROV|16|31|Gray hair is a crown of glory; it is gained in a righteous life.
PROV|16|32|Whoever is slow to anger is better than the mighty, and he who rules his spirit than he who takes a city.
PROV|16|33|The lot is cast into the lap, but its every decision is from the LORD.
PROV|17|1|Better is a dry morsel with quiet than a house full of feasting with strife.
PROV|17|2|A servant who deals wisely will rule over a son who acts shamefully and will share the inheritance as one of the brothers.
PROV|17|3|The crucible is for silver, and the furnace is for gold, and the LORD tests hearts.
PROV|17|4|An evildoer listens to wicked lips, and a liar gives ear to a mischievous tongue.
PROV|17|5|Whoever mocks the poor insults his Maker; he who is glad at calamity will not go unpunished.
PROV|17|6|Grandchildren are the crown of the aged, and the glory of children is their fathers.
PROV|17|7|Fine speech is not becoming to a fool; still less is false speech to a prince.
PROV|17|8|A bribe is like a magic stone in the eyes of the one who gives it; wherever he turns he prospers.
PROV|17|9|Whoever covers an offense seeks love, but he who repeats a matter separates close friends.
PROV|17|10|A rebuke goes deeper into a man of understanding than a hundred blows into a fool.
PROV|17|11|An evil man seeks only rebellion, and a cruel messenger will be sent against him.
PROV|17|12|Let a man meet a she-bear robbed of her cubs rather than a fool in his folly.
PROV|17|13|If anyone returns evil for good, evil will not depart from his house.
PROV|17|14|The beginning of strife is like letting out water, so quit before the quarrel breaks out.
PROV|17|15|He who justifies the wicked and he who condemns the righteous are both alike an abomination to the LORD.
PROV|17|16|Why should a fool have money in his hand to buy wisdom when he has no sense?
PROV|17|17|A friend loves at all times, and a brother is born for adversity.
PROV|17|18|One who lacks sense gives a pledge and puts up security in the presence of his neighbor.
PROV|17|19|Whoever loves transgression loves strife; he who makes his door high seeks destruction.
PROV|17|20|A man of crooked heart does not discover good, and one with a dishonest tongue falls into calamity.
PROV|17|21|He who sires a fool gets himself sorrow, and the father of a fool has no joy.
PROV|17|22|A joyful heart is good medicine, but a crushed spirit dries up the bones.
PROV|17|23|The wicked accepts a bribe in secret to pervert the ways of justice.
PROV|17|24|The discerning sets his face toward wisdom, but the eyes of a fool are on the ends of the earth.
PROV|17|25|A foolish son is a grief to his father and bitterness to her who bore him.
PROV|17|26|To impose a fine on a righteous man is not good, nor to strike the noble for their uprightness.
PROV|17|27|Whoever restrains his words has knowledge, and he who has a cool spirit is a man of understanding.
PROV|17|28|Even a fool who keeps silent is considered wise; when he closes his lips, he is deemed intelligent.
PROV|18|1|Whoever isolates himself seeks his own desire; he breaks out against all sound judgment.
PROV|18|2|A fool takes no pleasure in understanding, but only in expressing his opinion.
PROV|18|3|When wickedness comes, contempt comes also, and with dishonor comes disgrace.
PROV|18|4|The words of a man's mouth are deep waters; the fountain of wisdom is a bubbling brook.
PROV|18|5|It is not good to be partial to the wicked or to deprive the righteous of justice.
PROV|18|6|A fool's lips walk into a fight, and his mouth invites a beating.
PROV|18|7|A fool's mouth is his ruin, and his lips are a snare to his soul.
PROV|18|8|The words of a whisperer are like delicious morsels; they go down into the inner parts of the body.
PROV|18|9|Whoever is slack in his work is a brother to him who destroys.
PROV|18|10|The name of the LORD is a strong tower; the righteous man runs into it and is safe.
PROV|18|11|A rich man's wealth is his strong city, and like a high wall in his imagination.
PROV|18|12|Before destruction a man's heart is haughty, but humility comes before honor.
PROV|18|13|If one gives an answer before he hears, it is his folly and shame.
PROV|18|14|A man's spirit will endure sickness, but a crushed spirit who can bear?
PROV|18|15|An intelligent heart acquires knowledge, and the ear of the wise seeks knowledge.
PROV|18|16|A man's gift makes room for him and brings him before the great.
PROV|18|17|The one who states his case first seems right, until the other comes and examines him.
PROV|18|18|The lot puts an end to quarrels and decides between powerful contenders.
PROV|18|19|A brother offended is more unyielding than a strong city, and quarreling is like the bars of a castle.
PROV|18|20|From the fruit of a man's mouth his stomach is satisfied; he is satisfied by the yield of his lips.
PROV|18|21|Death and life are in the power of the tongue, and those who love it will eat its fruits.
PROV|18|22|He who finds a wife finds a good thing and obtains favor from the LORD.
PROV|18|23|The poor use entreaties, but the rich answer roughly.
PROV|18|24|A man of many companions may come to ruin, but there is a friend who sticks closer than a brother.
PROV|19|1|Better is a poor person who walks in his integrity than one who is crooked in speech and is a fool.
PROV|19|2|Desire without knowledge is not good, and whoever makes haste with his feet misses his way.
PROV|19|3|When a man's folly brings his way to ruin, his heart rages against the LORD.
PROV|19|4|Wealth brings many new friends, but a poor man is deserted by his friend.
PROV|19|5|A false witness will not go unpunished, and he who breathes out lies will not escape.
PROV|19|6|Many seek the favor of a generous man, and everyone is a friend to a man who gives gifts.
PROV|19|7|All a poor man's brothers hate him; how much more do his friends go far from him! He pursues them with words, but does not have them.
PROV|19|8|Whoever gets sense loves his own soul; he who keeps understanding will discover good.
PROV|19|9|A false witness will not go unpunished, and he who breathes out lies will perish.
PROV|19|10|It is not fitting for a fool to live in luxury, much less for a slave to rule over princes.
PROV|19|11|Good sense makes one slow to anger, and it is his glory to overlook an offense.
PROV|19|12|A king's wrath is like the growling of a lion, but his favor is like dew on the grass.
PROV|19|13|A foolish son is ruin to his father, and a wife's quarreling is a continual dripping of rain.
PROV|19|14|House and wealth are inherited from fathers, but a prudent wife is from the LORD.
PROV|19|15|Slothfulness casts into a deep sleep, and an idle person will suffer hunger.
PROV|19|16|Whoever keeps the commandment keeps his life; he who despises his ways will die.
PROV|19|17|Whoever is generous to the poor lends to the LORD, and he will repay him for his deed.
PROV|19|18|Discipline your son, for there is hope; do not set your heart on putting him to death.
PROV|19|19|A man of great wrath will pay the penalty, for if you deliver him, you will only have to do it again.
PROV|19|20|Listen to advice and accept instruction, that you may gain wisdom in the future.
PROV|19|21|Many are the plans in the mind of a man, but it is the purpose of the LORD that will stand.
PROV|19|22|What is desired in a man is steadfast love, and a poor man is better than a liar.
PROV|19|23|The fear of the LORD leads to life, and whoever has it rests satisfied; he will not be visited by harm.
PROV|19|24|The sluggard buries his hand in the dish and will not even bring it back to his mouth.
PROV|19|25|Strike a scoffer, and the simple will learn prudence; reprove a man of understanding, and he will gain knowledge.
PROV|19|26|He who does violence to his father and chases away his mother is a son who brings shame and reproach.
PROV|19|27|Cease to hear instruction, my son, and you will stray from the words of knowledge.
PROV|19|28|A worthless witness mocks at justice, and the mouth of the wicked devours iniquity.
PROV|19|29|Condemnation is ready for scoffers, and beating for the backs of fools.
PROV|20|1|Wine is a mocker, strong drink a brawler, and whoever is led astray by it is not wise.
PROV|20|2|The terror of a king is like the growling of a lion; whoever provokes him to anger forfeits his life.
PROV|20|3|It is an honor for a man to keep aloof from strife, but every fool will be quarreling.
PROV|20|4|The sluggard does not plow in the autumn; he will seek at harvest and have nothing.
PROV|20|5|The purpose in a man's heart is like deep water, but a man of understanding will draw it out.
PROV|20|6|Many a man proclaims his own steadfast love, but a faithful man who can find?
PROV|20|7|The righteous who walks in his integrity- blessed are his children after him!
PROV|20|8|A king who sits on the throne of judgment winnows all evil with his eyes.
PROV|20|9|Who can say, "I have made my heart pure; I am clean from my sin"?
PROV|20|10|Unequal weights and unequal measures are both alike an abomination to the LORD.
PROV|20|11|Even a child makes himself known by his acts, by whether his conduct is pure and upright.
PROV|20|12|The hearing ear and the seeing eye, the LORD has made them both.
PROV|20|13|Love not sleep, lest you come to poverty; open your eyes, and you will have plenty of bread.
PROV|20|14|"Bad, Bad," says the buyer, but when he goes away, then he boasts.
PROV|20|15|There is gold and abundance of costly stones, but the lips of knowledge are a precious jewel.
PROV|20|16|Take a man's garment when he has put up security for a stranger, and hold it in pledge when he puts up security for foreigners.
PROV|20|17|Bread gained by deceit is sweet to a man, but afterward his mouth will be full of gravel.
PROV|20|18|Plans are established by counsel; by wise guidance wage war.
PROV|20|19|Whoever goes about slandering reveals secrets; therefore do not associate with a simple babbler.
PROV|20|20|If one curses his father or his mother, his lamp will be put out in utter darkness.
PROV|20|21|An inheritance gained hastily in the beginning will not be blessed in the end.
PROV|20|22|Do not say, "I will repay evil"; wait for the LORD, and he will deliver you.
PROV|20|23|Unequal weights are an abomination to the LORD, and false scales are not good.
PROV|20|24|A man's steps are from the LORD; how then can man understand his way?
PROV|20|25|It is a snare to say rashly, "It is holy," and to reflect only after making vows.
PROV|20|26|A wise king winnows the wicked and drives the wheel over them.
PROV|20|27|The spirit of man is the lamp of the LORD, searching all his innermost parts.
PROV|20|28|Steadfast love and faithfulness preserve the king, and by steadfast love his throne is upheld.
PROV|20|29|The glory of young men is their strength, but the splendor of old men is their gray hair.
PROV|20|30|Blows that wound cleanse away evil; strokes make clean the innermost parts.
PROV|21|1|The king's heart is a stream of water in the hand of the LORD; he turns it wherever he will.
PROV|21|2|Every way of a man is right in his own eyes, but the LORD weighs the heart.
PROV|21|3|To do righteousness and justice is more acceptable to the LORD than sacrifice.
PROV|21|4|Haughty eyes and a proud heart, the lamp of the wicked, are sin.
PROV|21|5|The plans of the diligent lead surely to abundance, but everyone who is hasty comes only to poverty.
PROV|21|6|The getting of treasures by a lying tongue is a fleeting vapor and a snare of death.
PROV|21|7|The violence of the wicked will sweep them away, because they refuse to do what is just.
PROV|21|8|The way of the guilty is crooked, but the conduct of the pure is upright.
PROV|21|9|It is better to live in a corner of the housetop than in a house shared with a quarrelsome wife.
PROV|21|10|The soul of the wicked desires evil; his neighbor finds no mercy in his eyes.
PROV|21|11|When a scoffer is punished, the simple becomes wise; when a wise man is instructed, he gains knowledge.
PROV|21|12|The Righteous One observes the house of the wicked; he throws the wicked down to ruin.
PROV|21|13|Whoever closes his ear to the cry of the poor will himself call out and not be answered.
PROV|21|14|A gift in secret averts anger, and a concealed bribe, strong wrath.
PROV|21|15|When justice is done, it is a joy to the righteous but terror to evildoers.
PROV|21|16|One who wanders from the way of good sense will rest in the assembly of the dead.
PROV|21|17|Whoever loves pleasure will be a poor man; he who loves wine and oil will not be rich.
PROV|21|18|The wicked is a ransom for the righteous, and the traitor for the upright.
PROV|21|19|It is better to live in a desert land than with a quarrelsome and fretful woman.
PROV|21|20|Precious treasure and oil are in a wise man's dwelling, but a foolish man devours it.
PROV|21|21|Whoever pursues righteousness and kindness will find life, righteousness, and honor.
PROV|21|22|A wise man scales the city of the mighty and brings down the stronghold in which they trust.
PROV|21|23|Whoever keeps his mouth and his tongue keeps himself out of trouble.
PROV|21|24|"Scoffer" is the name of the arrogant, haughty man who acts with arrogant pride.
PROV|21|25|The desire of the sluggard kills him, for his hands refuse to labor.
PROV|21|26|All day long he craves and craves, but the righteous gives and does not hold back.
PROV|21|27|The sacrifice of the wicked is an abomination; how much more when he brings it with evil intent.
PROV|21|28|A false witness will perish, but the word of a man who hears will endure.
PROV|21|29|A wicked man puts on a bold face, but the upright gives thought to his ways.
PROV|21|30|No wisdom, no understanding, no counsel can avail against the LORD.
PROV|21|31|The horse is made ready for the day of battle, but the victory belongs to the LORD.
PROV|22|1|A good name is to be chosen rather than great riches, and favor is better than silver or gold.
PROV|22|2|The rich and the poor meet together; the LORD is the maker of them all.
PROV|22|3|The prudent sees danger and hides himself, but the simple go on and suffer for it.
PROV|22|4|The reward for humility and fear of the LORD is riches and honor and life.
PROV|22|5|Thorns and snares are in the way of the crooked; whoever guards his soul will keep far from them.
PROV|22|6|Train up a child in the way he should go; even when he is old he will not depart from it.
PROV|22|7|The rich rules over the poor, and the borrower is the slave of the lender.
PROV|22|8|Whoever sows injustice will reap calamity, and the rod of his fury will fail.
PROV|22|9|Whoever has a bountiful eye will be blessed, for he shares his bread with the poor.
PROV|22|10|Drive out a scoffer, and strife will go out, and quarreling and abuse will cease.
PROV|22|11|He who loves purity of heart, and whose speech is gracious, will have the king as his friend.
PROV|22|12|The eyes of the LORD keep watch over knowledge, but he overthrows the words of the traitor.
PROV|22|13|The sluggard says, "There is a lion outside! I shall be killed in the streets!"
PROV|22|14|The mouth of forbidden women is a deep pit; he with whom the LORD is angry will fall into it.
PROV|22|15|Folly is bound up in the heart of a child, but the rod of discipline drives it far from him.
PROV|22|16|Whoever oppresses the poor to increase his own wealth, or gives to the rich, will only come to poverty.
PROV|22|17|Incline your ear, and hear the words of the wise, and apply your heart to my knowledge,
PROV|22|18|for it will be pleasant if you keep them within you, if all of them are ready on your lips.
PROV|22|19|That your trust may be in the LORD, I have made them known to you today, even to you.
PROV|22|20|Have I not written for you thirty sayings of counsel and knowledge,
PROV|22|21|to make you know what is right and true, that you may give a true answer to those who sent you?
PROV|22|22|Do not rob the poor, because he is poor, or crush the afflicted at the gate,
PROV|22|23|for the LORD will plead their cause and rob of life those who rob them.
PROV|22|24|Make no friendship with a man given to anger, nor go with a wrathful man,
PROV|22|25|lest you learn his ways and entangle yourself in a snare.
PROV|22|26|Be not one of those who give pledges, who put up security for debts.
PROV|22|27|If you have nothing with which to pay, why should your bed be taken from under you?
PROV|22|28|Do not move the ancient landmark that your fathers have set.
PROV|22|29|Do you see a man skillful in his work? He will stand before kings; he will not stand before obscure men.
PROV|23|1|When you sit down to eat with a ruler, observe carefully what is before you,
PROV|23|2|and put a knife to your throat if you are given to appetite.
PROV|23|3|Do not desire his delicacies, for they are deceptive food.
PROV|23|4|Do not toil to acquire wealth; be discerning enough to desist.
PROV|23|5|When your eyes light on it, it is gone, for suddenly it sprouts wings, flying like an eagle toward heaven.
PROV|23|6|Do not eat the bread of a man who is stingy; do not desire his delicacies,
PROV|23|7|for he is like one who is inwardly calculating. "Eat and drink!" he says to you, but his heart is not with you.
PROV|23|8|You will vomit up the morsels that you have eaten, and waste your pleasant words.
PROV|23|9|Do not speak in the hearing of a fool, for he will despise the good sense of your words.
PROV|23|10|Do not move an ancient landmark or enter the fields of the fatherless,
PROV|23|11|for their Redeemer is strong; he will plead their cause against you.
PROV|23|12|Apply your heart to instruction and your ear to words of knowledge.
PROV|23|13|Do not withhold discipline from a child; if you strike him with a rod, he will not die.
PROV|23|14|If you strike him with the rod, you will save his soul from Sheol.
PROV|23|15|My son, if your heart is wise, my heart too will be glad.
PROV|23|16|My inmost being will exult when your lips speak what is right.
PROV|23|17|Let not your heart envy sinners, but continue in the fear of the LORD all the day.
PROV|23|18|Surely there is a future, and your hope will not be cut off.
PROV|23|19|Hear, my son, and be wise, and direct your heart in the way.
PROV|23|20|Be not among drunkards or among gluttonous eaters of meat,
PROV|23|21|for the drunkard and the glutton will come to poverty, and slumber will clothe them with rags.
PROV|23|22|Listen to your father who gave you life, and do not despise your mother when she is old.
PROV|23|23|Buy truth, and do not sell it; buy wisdom, instruction, and understanding.
PROV|23|24|The father of the righteous will greatly rejoice; he who fathers a wise son will be glad in him.
PROV|23|25|Let your father and mother be glad; let her who bore you rejoice.
PROV|23|26|My son, give me your heart, and let your eyes observe my ways.
PROV|23|27|For a prostitute is a deep pit; an adulteress is a narrow well.
PROV|23|28|She lies in wait like a robber and increases the traitors among mankind.
PROV|23|29|Who has woe? Who has sorrow? Who has strife? Who has complaining? Who has wounds without cause? Who has redness of eyes?
PROV|23|30|Those who tarry long over wine; those who go to try mixed wine.
PROV|23|31|Do not look at wine when it is red, when it sparkles in the cup and goes down smoothly.
PROV|23|32|In the end it bites like a serpent and stings like an adder.
PROV|23|33|Your eyes will see strange things, and your heart utter perverse things.
PROV|23|34|You will be like one who lies down in the midst of the sea, like one who lies on the top of a mast.
PROV|23|35|"They struck me," you will say, "but I was not hurt; they beat me, but I did not feel it. When shall I awake? I must have another drink."
PROV|24|1|Be not envious of evil men, nor desire to be with them,
PROV|24|2|for their hearts devise violence, and their lips talk of trouble.
PROV|24|3|By wisdom a house is built, and by understanding it is established;
PROV|24|4|by knowledge the rooms are filled with all precious and pleasant riches.
PROV|24|5|A wise man is full of strength, and a man of knowledge enhances his might,
PROV|24|6|for by wise guidance you can wage your war, and in abundance of counselors there is victory.
PROV|24|7|Wisdom is too high for a fool; in the gate he does not open his mouth.
PROV|24|8|Whoever plans to do evil will be called a schemer.
PROV|24|9|The devising of folly is sin, and the scoffer is an abomination to mankind.
PROV|24|10|If you faint in the day of adversity, your strength is small.
PROV|24|11|Rescue those who are being taken away to death; hold back those who are stumbling to the slaughter.
PROV|24|12|If you say, "Behold, we did not know this," does not he who weighs the heart perceive it? Does not he who keeps watch over your soul know it, and will he not repay man according to his work?
PROV|24|13|My son, eat honey, for it is good, and the drippings of the honeycomb are sweet to your taste.
PROV|24|14|Know that wisdom is such to your soul; if you find it, there will be a future, and your hope will not be cut off.
PROV|24|15|Lie not in wait as a wicked man against the dwelling of the righteous; do no violence to his home;
PROV|24|16|for the righteous falls seven times and rises again, but the wicked stumble in times of calamity.
PROV|24|17|Do not rejoice when your enemy falls, and let not your heart be glad when he stumbles,
PROV|24|18|lest the LORD see it and be displeased, and turn away his anger from him.
PROV|24|19|Fret not yourself because of evildoers, and be not envious of the wicked,
PROV|24|20|for the evil man has no future; the lamp of the wicked will be put out.
PROV|24|21|My son, fear the LORD and the king, and do not join with those who do otherwise,
PROV|24|22|for disaster from them will rise suddenly, and who knows the ruin that will come from them both?
PROV|24|23|These also are sayings of the wise. Partiality in judging is not good.
PROV|24|24|Whoever says to the wicked, "You are in the right," will be cursed by peoples, abhorred by nations,
PROV|24|25|but those who rebuke the wicked will have delight, and a good blessing will come upon them.
PROV|24|26|Whoever gives an honest answer kisses the lips.
PROV|24|27|Prepare your work outside; get everything ready for yourself in the field, and after that build your house.
PROV|24|28|Be not a witness against your neighbor without cause, and do not deceive with your lips.
PROV|24|29|Do not say, "I will do to him as he has done to me; I will pay the man back for what he has done."
PROV|24|30|I passed by the field of a sluggard, by the vineyard of a man lacking sense,
PROV|24|31|and behold, it was all overgrown with thorns; the ground was covered with nettles, and its stone wall was broken down.
PROV|24|32|Then I saw and considered it; I looked and received instruction.
PROV|24|33|A little sleep, a little slumber, a little folding of the hands to rest,
PROV|24|34|and poverty will come upon you like a robber, and want like an armed man.
PROV|25|1|These also are proverbs of Solomon which the men of Hezekiah king of Judah copied.
PROV|25|2|It is the glory of God to conceal things, but the glory of kings is to search things out.
PROV|25|3|As the heavens for height, and the earth for depth, so the heart of kings is unsearchable.
PROV|25|4|Take away the dross from the silver, and the smith has material for a vessel;
PROV|25|5|take away the wicked from the presence of the king, and his throne will be established in righteousness.
PROV|25|6|Do not put yourself forward in the king's presence or stand in the place of the great,
PROV|25|7|for it is better to be told, "Come up here," than to be put lower in the presence of a noble. What your eyes have seen
PROV|25|8|do not hastily bring into court, for what will you do in the end, when your neighbor puts you to shame?
PROV|25|9|Argue your case with your neighbor himself, and do not reveal another's secret,
PROV|25|10|lest he who hears you bring shame upon you, and your ill repute have no end.
PROV|25|11|A word fitly spoken is like apples of gold in a setting of silver.
PROV|25|12|Like a gold ring or an ornament of gold is a wise reprover to a listening ear.
PROV|25|13|Like the cold of snow in the time of harvest is a faithful messenger to those who send him; he refreshes the soul of his masters.
PROV|25|14|Like clouds and wind without rain is a man who boasts of a gift he does not give.
PROV|25|15|With patience a ruler may be persuaded, and a soft tongue will break a bone.
PROV|25|16|If you have found honey, eat only enough for you, lest you have your fill of it and vomit it.
PROV|25|17|Let your foot be seldom in your neighbor's house, lest he have his fill of you and hate you.
PROV|25|18|A man who bears false witness against his neighbor is like a war club, or a sword, or a sharp arrow.
PROV|25|19|Trusting in a treacherous man in time of trouble is like a bad tooth or a foot that slips.
PROV|25|20|Whoever sings songs to a heavy heart is like one who takes off a garment on a cold day, and like vinegar on soda.
PROV|25|21|If your enemy is hungry, give him bread to eat, and if he is thirsty, give him water to drink,
PROV|25|22|for you will heap burning coals on his head, and the LORD will reward you.
PROV|25|23|The north wind brings forth rain, and a backbiting tongue, angry looks.
PROV|25|24|It is better to live in a corner of the housetop than in a house shared with a quarrelsome wife.
PROV|25|25|Like cold water to a thirsty soul, so is good news from a far country.
PROV|25|26|Like a muddied spring or a polluted fountain is a righteous man who gives way before the wicked.
PROV|25|27|It is not good to eat much honey, nor is it glorious to seek one's own glory.
PROV|25|28|A man without self-control is like a city broken into and left without walls.
PROV|26|1|Like snow in summer or rain in harvest, so honor is not fitting for a fool.
PROV|26|2|Like a sparrow in its flitting, like a swallow in its flying, a curse that is causeless does not alight.
PROV|26|3|A whip for the horse, a bridle for the donkey, and a rod for the back of fools.
PROV|26|4|Answer not a fool according to his folly, lest you be like him yourself.
PROV|26|5|Answer a fool according to his folly, lest he be wise in his own eyes.
PROV|26|6|Whoever sends a message by the hand of a fool cuts off his own feet and drinks violence.
PROV|26|7|Like a lame man's legs, which hang useless, is a proverb in the mouth of fools.
PROV|26|8|Like one who binds the stone in the sling is one who gives honor to a fool.
PROV|26|9|Like a thorn that goes up into the hand of a drunkard is a proverb in the mouth of fools.
PROV|26|10|Like an archer who wounds everybody is one who hires a passing fool or drunkard.
PROV|26|11|Like a dog that returns to his vomit is a fool who repeats his folly.
PROV|26|12|Do you see a man who is wise in his own eyes? There is more hope for a fool than for him.
PROV|26|13|The sluggard says, "There is a lion in the road! There is a lion in the streets!"
PROV|26|14|As a door turns on its hinges, so does a sluggard on his bed.
PROV|26|15|The sluggard buries his hand in the dish; it wears him out to bring it back to his mouth.
PROV|26|16|The sluggard is wiser in his own eyes than seven men who can answer sensibly.
PROV|26|17|Whoever meddles in a quarrel not his own is like one who takes a passing dog by the ears.
PROV|26|18|Like a madman who throws firebrands, arrows, and death
PROV|26|19|is the man who deceives his neighbor and says, "I am only joking!"
PROV|26|20|For lack of wood the fire goes out, and where there is no whisperer, quarreling ceases.
PROV|26|21|As charcoal to hot embers and wood to fire, so is a quarrelsome man for kindling strife.
PROV|26|22|The words of a whisperer are like delicious morsels; they go down into the inner parts of the body.
PROV|26|23|Like the glaze covering an earthen vessel are fervent lips with an evil heart.
PROV|26|24|Whoever hates disguises himself with his lips and harbors deceit in his heart;
PROV|26|25|when he speaks graciously, believe him not, for there are seven abominations in his heart;
PROV|26|26|though his hatred be covered with deception, his wickedness will be exposed in the assembly.
PROV|26|27|Whoever digs a pit will fall into it, and a stone will come back on him who starts it rolling.
PROV|26|28|A lying tongue hates its victims, and a flattering mouth works ruin.
PROV|27|1|Do not boast about tomorrow, for you do not know what a day may bring.
PROV|27|2|Let another praise you, and not your own mouth; a stranger, and not your own lips.
PROV|27|3|A stone is heavy, and sand is weighty, but a fool's provocation is heavier than both.
PROV|27|4|Wrath is cruel, anger is overwhelming, but who can stand before jealousy?
PROV|27|5|Better is open rebuke than hidden love.
PROV|27|6|Faithful are the wounds of a friend; profuse are the kisses of an enemy.
PROV|27|7|One who is full loathes honey, but to one who is hungry everything bitter is sweet.
PROV|27|8|Like a bird that strays from its nest is a man who strays from his home.
PROV|27|9|Oil and perfume make the heart glad, and the sweetness of a friend comes from his earnest counsel.
PROV|27|10|Do not forsake your friend and your father's friend, and do not go to your brother's house in the day of your calamity. Better is a neighbor who is near than a brother who is far away.
PROV|27|11|Be wise, my son, and make my heart glad, that I may answer him who reproaches me.
PROV|27|12|The prudent sees danger and hides himself, but the simple go on and suffer for it.
PROV|27|13|Take a man's garment when he has put up security for a stranger, and hold it in pledge when he puts up security for an adulteress.
PROV|27|14|Whoever blesses his neighbor with a loud voice, rising early in the morning, will be counted as cursing.
PROV|27|15|A continual dripping on a rainy day and a quarrelsome wife are alike;
PROV|27|16|to restrain her is to restrain the wind or to grasp oil in one's right hand.
PROV|27|17|Iron sharpens iron, and one man sharpens another.
PROV|27|18|Whoever tends a fig tree will eat its fruit, and he who guards his master will be honored.
PROV|27|19|As in water face reflects face, so the heart of man reflects the man.
PROV|27|20|Sheol and Abaddon are never satisfied, and never satisfied are the eyes of man.
PROV|27|21|The crucible is for silver, and the furnace is for gold, and a man is tested by his praise.
PROV|27|22|Crush a fool in a mortar with a pestle along with crushed grain, yet his folly will not depart from him.
PROV|27|23|Know well the condition of your flocks, and give attention to your herds,
PROV|27|24|for riches do not last forever; and does a crown endure to all generations?
PROV|27|25|When the grass is gone and the new growth appears and the vegetation of the mountains is gathered,
PROV|27|26|the lambs will provide your clothing, and the goats the price of a field.
PROV|27|27|There will be enough goats' milk for your food, for the food of your household and maintenance for your girls.
PROV|28|1|The wicked flee when no one pursues, but the righteous are bold as a lion.
PROV|28|2|When a land transgresses, it has many rulers, but with a man of understanding and knowledge, its stability will long continue.
PROV|28|3|A poor man who oppresses the poor is a beating rain that leaves no food.
PROV|28|4|Those who forsake the law praise the wicked, but those who keep the law strive against them.
PROV|28|5|Evil men do not understand justice, but those who seek the LORD understand it completely.
PROV|28|6|Better is a poor man who walks in his integrity than a rich man who is crooked in his ways.
PROV|28|7|The one who keeps the law is a son with understanding, but a companion of gluttons shames his father.
PROV|28|8|Whoever multiplies his wealth by interest and profit gathers it for him who is generous to the poor.
PROV|28|9|If one turns away his ear from hearing the law, even his prayer is an abomination.
PROV|28|10|Whoever misleads the upright into an evil way will fall into his own pit, but the blameless will have a goodly inheritance.
PROV|28|11|A rich man is wise in his own eyes, but a poor man who has understanding will find him out.
PROV|28|12|When the righteous triumph, there is great glory, but when the wicked rise, people hide themselves.
PROV|28|13|Whoever conceals his transgressions will not prosper, but he who confesses and forsakes them will obtain mercy.
PROV|28|14|Blessed is the one who fears the LORD always, but whoever hardens his heart will fall into calamity.
PROV|28|15|Like a roaring lion or a charging bear is a wicked ruler over a poor people.
PROV|28|16|A ruler who lacks understanding is a cruel oppressor, but he who hates unjust gain will prolong his days.
PROV|28|17|If one is burdened with the blood of another, he will be a fugitive until death; let no one help him.
PROV|28|18|Whoever walks in integrity will be delivered, but he who is crooked in his ways will suddenly fall.
PROV|28|19|Whoever works his land will have plenty of bread, but he who follows worthless pursuits will have plenty of poverty.
PROV|28|20|A faithful man will abound with blessings, but whoever hastens to be rich will not go unpunished.
PROV|28|21|To show partiality is not good, but for a piece of bread a man will do wrong.
PROV|28|22|A stingy man hastens after wealth and does not know that poverty will come upon him.
PROV|28|23|Whoever rebukes a man will afterward find more favor than he who flatters with his tongue.
PROV|28|24|Whoever robs his father or his mother and says, "That is no transgression," is a companion to a man who destroys.
PROV|28|25|A greedy man stirs up strife, but the one who trusts in the LORD will be enriched.
PROV|28|26|Whoever trusts in his own mind is a fool, but he who walks in wisdom will be delivered.
PROV|28|27|Whoever gives to the poor will not want, but he who hides his eyes will get many a curse.
PROV|28|28|When the wicked rise, people hide themselves, but when they perish, the righteous increase.
PROV|29|1|He who is often reproved, yet stiffens his neck, will suddenly be broken beyond healing.
PROV|29|2|When the righteous increase, the people rejoice, but when the wicked rule, the people groan.
PROV|29|3|He who loves wisdom makes his father glad, but a companion of prostitutes squanders his wealth.
PROV|29|4|By justice a king builds up the land, but he who exacts gifts tears it down.
PROV|29|5|A man who flatters his neighbor spreads a net for his feet.
PROV|29|6|An evil man is ensnared in his transgression, but a righteous man sings and rejoices.
PROV|29|7|A righteous man knows the rights of the poor; a wicked man does not understand such knowledge.
PROV|29|8|Scoffers set a city aflame, but the wise turn away wrath.
PROV|29|9|If a wise man has an argument with a fool, the fool only rages and laughs, and there is no quiet.
PROV|29|10|Bloodthirsty men hate one who is blameless and seek the life of the upright.
PROV|29|11|A fool gives full vent to his spirit, but a wise man quietly holds it back.
PROV|29|12|If a ruler listens to falsehood, all his officials will be wicked.
PROV|29|13|The poor man and the oppressor meet together; the LORD gives light to the eyes of both.
PROV|29|14|If a king faithfully judges the poor, his throne will be established forever.
PROV|29|15|The rod and reproof give wisdom, but a child left to himself brings shame to his mother.
PROV|29|16|When the wicked increase, transgression increases, but the righteous will look upon their downfall.
PROV|29|17|Discipline your son, and he will give you rest; he will give delight to your heart.
PROV|29|18|Where there is no prophetic vision the people cast off restraint, but blessed is he who keeps the law.
PROV|29|19|By mere words a servant is not disciplined, for though he understands, he will not respond.
PROV|29|20|Do you see a man who is hasty in his words? There is more hope for a fool than for him.
PROV|29|21|Whoever pampers his servant from childhood will in the end find him his heir.
PROV|29|22|A man of wrath stirs up strife, and one given to anger causes much transgression.
PROV|29|23|One's pride will bring him low, but he who is lowly in spirit will obtain honor.
PROV|29|24|The partner of a thief hates his own life; he hears the curse, but discloses nothing.
PROV|29|25|The fear of man lays a snare, but whoever trusts in the LORD is safe.
PROV|29|26|Many seek the face of a ruler, but it is from the LORD that a man gets justice.
PROV|29|27|An unjust man is an abomination to the righteous, but one whose way is straight is an abomination to the wicked.
PROV|30|1|The words of Agur son of Jakeh. The oracle. The man declares, I am weary, O God; I am weary, O God, and worn out.
PROV|30|2|Surely I am too stupid to be a man. I have not the understanding of a man.
PROV|30|3|I have not learned wisdom, nor have I knowledge of the Holy One.
PROV|30|4|Who has ascended to heaven and come down? Who has gathered the wind in his fists? Who has wrapped up the waters in a garment? Who has established all the ends of the earth? What is his name, and what is his son's name? Surely you know!
PROV|30|5|Every word of God proves true; he is a shield to those who take refuge in him.
PROV|30|6|Do not add to his words, lest he rebuke you and you be found a liar.
PROV|30|7|Two things I ask of you; deny them not to me before I die:
PROV|30|8|Remove far from me falsehood and lying; give me neither poverty nor riches; feed me with the food that is needful for me,
PROV|30|9|lest I be full and deny you and say, "Who is the LORD?" or lest I be poor and steal and profane the name of my God.
PROV|30|10|Do not slander a servant to his master, lest he curse you and you be held guilty.
PROV|30|11|There are those who curse their fathers and do not bless their mothers.
PROV|30|12|There are those who are clean in their own eyes but are not washed of their filth.
PROV|30|13|There are those- how lofty are their eyes, how high their eyelids lift!
PROV|30|14|There are those whose teeth are swords, whose fangs are knives, to devour the poor from off the earth, the needy from among mankind.
PROV|30|15|The leech has two daughters; "Give" and "Give," they cry. Three things are never satisfied; four never say, "Enough":
PROV|30|16|Sheol, the barren womb, the land never satisfied with water, and the fire that never says, "Enough."
PROV|30|17|The eye that mocks a father and scorns to obey a mother will be picked out by the ravens of the valley and eaten by the vultures.
PROV|30|18|Three things are too wonderful for me; four I do not understand:
PROV|30|19|the way of an eagle in the sky, the way of a serpent on a rock, the way of a ship on the high seas, and the way of a man with a virgin.
PROV|30|20|This is the way of an adulteress: she eats and wipes her mouth and says, "I have done no wrong."
PROV|30|21|Under three things the earth trembles; under four it cannot bear up:
PROV|30|22|a slave when he becomes king, and a fool when he is filled with food;
PROV|30|23|an unloved woman when she gets a husband, and a maidservant when she displaces her mistress.
PROV|30|24|Four things on earth are small, but they are exceedingly wise:
PROV|30|25|the ants are a people not strong, yet they provide their food in the summer;
PROV|30|26|the rock badgers are a people not mighty, yet they make their homes in the cliffs;
PROV|30|27|the locusts have no king, yet all of them march in rank;
PROV|30|28|the lizard you can take in your hands, yet it is in kings' palaces.
PROV|30|29|Three things are stately in their tread; four are stately in their stride:
PROV|30|30|the lion, which is mightiest among beasts and does not turn back before any;
PROV|30|31|the strutting rooster, the he-goat, and a king whose army is with him.
PROV|30|32|If you have been foolish, exalting yourself, or if you have been devising evil, put your hand on your mouth.
PROV|30|33|For pressing milk produces curds, pressing the nose produces blood, and pressing anger produces strife.
PROV|31|1|The words of King Lemuel. An oracle that his mother taught him:
PROV|31|2|What are you doing, my son? What are you doing, son of my womb? What are you doing, son of my vows?
PROV|31|3|Do not give your strength to women, your ways to those who destroy kings.
PROV|31|4|It is not for kings, O Lemuel, it is not for kings to drink wine, or for rulers to take strong drink,
PROV|31|5|lest they drink and forget what has been decreed and pervert the rights of all the afflicted.
PROV|31|6|Give strong drink to the one who is perishing, and wine to those in bitter distress;
PROV|31|7|let them drink and forget their poverty and remember their misery no more.
PROV|31|8|Open your mouth for the mute, for the rights of all who are destitute.
PROV|31|9|Open your mouth, judge righteously, defend the rights of the poor and needy.
PROV|31|10|An excellent wife who can find? She is far more precious than jewels.
PROV|31|11|The heart of her husband trusts in her, and he will have no lack of gain.
PROV|31|12|She does him good, and not harm, all the days of her life.
PROV|31|13|She seeks wool and flax, and works with willing hands.
PROV|31|14|She is like the ships of the merchant; she brings her food from afar.
PROV|31|15|She rises while it is yet night and provides food for her household and portions for her maidens.
PROV|31|16|She considers a field and buys it; with the fruit of her hands she plants a vineyard.
PROV|31|17|She dresses herself with strength and makes her arms strong.
PROV|31|18|She perceives that her merchandise is profitable. Her lamp does not go out at night.
PROV|31|19|She puts her hands to the distaff, and her hands hold the spindle.
PROV|31|20|She opens her hand to the poor and reaches out her hands to the needy.
PROV|31|21|She is not afraid of snow for her household, for all her household are clothed in scarlet.
PROV|31|22|She makes bed coverings for herself; her clothing is fine linen and purple.
PROV|31|23|Her husband is known in the gates when he sits among the elders of the land.
PROV|31|24|She makes linen garments and sells them; she delivers sashes to the merchant.
PROV|31|25|Strength and dignity are her clothing, and she laughs at the time to come.
PROV|31|26|She opens her mouth with wisdom, and the teaching of kindness is on her tongue.
PROV|31|27|She looks well to the ways of her household and does not eat the bread of idleness.
PROV|31|28|Her children rise up and call her blessed; her husband also, and he praises her:
PROV|31|29|"Many women have done excellently, but you surpass them all."
PROV|31|30|Charm is deceitful, and beauty is vain, but a woman who fears the LORD is to be praised.
PROV|31|31|Give her of the fruit of her hands, and let her works praise her in the gates.
