1JOHN|1|1|論到從起初原有的生命之道，就是我們所聽見、所看見、親眼看過、親手摸過的－
1JOHN|1|2|這生命已經顯現出來，我們看見了，現在又作見證，把原與父同在，並且向我們顯現過的那永遠的生命傳揚給你們－
1JOHN|1|3|我們把所看見、所聽見的傳揚給你們，為要使你們也與我們有團契，而我們的團契是與父和他兒子耶穌基督所共有的。
1JOHN|1|4|我們把這些事寫給你們，使我們 的喜樂得以滿足。
1JOHN|1|5|上帝就是光，在他毫無黑暗；這是我們從主所聽見，又報給你們的信息。
1JOHN|1|6|我們若說，我們與上帝有團契，卻仍在黑暗裏行走，就是說謊話，不實行真理了。
1JOHN|1|7|我們若在光明中行走，如同上帝在光明中，就彼此有團契，他兒子耶穌的血就洗淨我們一切的罪。
1JOHN|1|8|我們若說自己沒有罪，就是欺騙自己，真理就不在我們裏面了。
1JOHN|1|9|我們若認自己的罪，上帝是信實的，是公義的，必要赦免我們的罪，洗淨我們一切的不義。
1JOHN|1|10|我們若說自己沒有犯過罪，就是把上帝當作說謊的，他的道就不在我們裏面了。
1JOHN|2|1|我的孩子們哪，我把這些話寫給你們，是要你們不犯罪。若有人犯罪，在父那裏我們有一位中保，就是那義者耶穌基督。
1JOHN|2|2|他為我們的罪作了贖罪祭，不單是為我們的罪，也是為普天下人的罪。
1JOHN|2|3|我們若遵守上帝的命令，就知道我們確實認識他。
1JOHN|2|4|人若說「我認識他」，卻不遵守他的命令，就是說謊話的，真理就不在他裏面了。
1JOHN|2|5|凡遵守他的道的，愛上帝的心確實地在他裏面達到完全了。由此我們知道我們是在他裏面。
1JOHN|2|6|凡說自己住在他裏面的，就該照著他所行的去行。
1JOHN|2|7|親愛的，我寫給你們的不是一條新命令，而是你們從起初所受的舊命令；這舊命令就是你們所聽過的道。
1JOHN|2|8|然而，我寫給你們的是一條新命令，在基督裏是真實的，在你們也是真實的，因為黑暗漸漸消逝，真光已經在照耀。
1JOHN|2|9|人若說自己在光明中，卻恨他的弟兄，他到如今還是在黑暗裏。
1JOHN|2|10|那愛弟兄的，就是住在光明中，他不會使人失足犯罪 。
1JOHN|2|11|惟獨那恨弟兄的，是在黑暗裏，也在黑暗裏行走，不知道往哪裏去，因為黑暗使他的眼睛瞎了。
1JOHN|2|12|孩子們哪，我寫信給你們， 因為你們的罪藉著基督的名得了赦免。
1JOHN|2|13|父老們啊，我寫信給你們， 因為你們認識從起初就有的那一位。 青年們哪，我寫信給你們， 因為你們勝過了那惡者。
1JOHN|2|14|孩子們哪，我曾寫信給你們， 因為你們認識父。 父老們啊，我曾寫信給你們， 因為你們認識從起初就有的那一位。 青年們哪，我曾寫信給你們， 因為你們剛強， 上帝的道常存在你們心裏， 你們也勝過了那惡者。
1JOHN|2|15|不要愛世界和世界上的東西，若有人愛世界，愛父的心就不在他裏面了。
1JOHN|2|16|因為凡世界上的東西，好比肉體的情慾、眼目的情慾和今生的驕傲，都不是從父來的，而是從世界來的。
1JOHN|2|17|這世界和世上的情慾都要消逝，惟獨那遵行上帝旨意的人永遠常存。
1JOHN|2|18|孩子們哪，如今是末世的時光了。你們曾聽過那敵基督者要來，現在有好些敵基督者已經出來了；由此我們就知道，如今是末世的時光了。
1JOHN|2|19|他們從我們中間出去，卻不是屬我們的，若是屬我們的，就必仍舊與我們同在。他們出去，這就顯明他們都不是屬我們的。
1JOHN|2|20|你們從那聖者受了恩膏，並且你們大家都知道 。
1JOHN|2|21|我寫信給你們，不是因你們不認識真理，而是因你們認識，並且知道一切虛謊都不是從真理出來的。
1JOHN|2|22|誰是說謊話的呢？不就是那不認耶穌為基督的嗎？那不認父與子的，這個人就是敵基督的。
1JOHN|2|23|凡不認子的，就沒有父；宣認子的，連父也有了。
1JOHN|2|24|論到你們，務要將那從起初所聽見的常存在心裏；若將從起初所聽見的存在心裏，你們就會住在子裏面，也會住在父裏面。
1JOHN|2|25|基督所應許我們的就是永生。
1JOHN|2|26|我將這些話寫給你們，是論到那些迷惑你們的人說的。
1JOHN|2|27|至於你們，你們從基督所受的恩膏常存在你們心裏，並不用人教導你們，自有他的恩膏在凡事上教導你們。這恩膏是真的，不是假的，你們要按這恩膏的教導住在他裏面。
1JOHN|2|28|孩子們哪，你們要住在基督裏面。這樣，他若顯現，我們就可以坦然無懼；當他來臨的時候，在他面前不至於慚愧。
1JOHN|2|29|你們若知道他是公義的，就知道凡行公義的人都是他所生的。
1JOHN|3|1|你們看父賜給我們的是何等的慈愛，讓我們得以稱為上帝的兒女；我們也真是他的兒女。世人不認識我們 的理由，是因他們未曾認識父。
1JOHN|3|2|親愛的，我們現在是上帝的兒女，將來如何還未顯明。我們所知道的是：基督顯現的時候，我們會像他，因為我們將見到他的本相。
1JOHN|3|3|凡對他有這指望的，就潔淨自己，像他是潔淨的一樣。
1JOHN|3|4|凡犯罪的，就是做違背律法的事；違背律法就是罪。
1JOHN|3|5|你們知道，基督曾顯現是要除掉罪 ；在他並沒有罪。
1JOHN|3|6|凡住在他裏面的，不犯罪；凡犯罪的，未曾看見他，也未曾認識他。
1JOHN|3|7|孩子們哪，不要讓人迷惑了你們；行義的才是義人，正如基督是義的。
1JOHN|3|8|犯罪的是出於魔鬼，因為魔鬼從起初就犯罪。上帝的兒子顯現出來，是為了要毀滅魔鬼的作為。
1JOHN|3|9|凡從上帝生的，不犯罪，因上帝的道 存在他裏面，他也不能犯罪，因為他是由上帝所生的。
1JOHN|3|10|這就顯明誰是上帝的兒女，誰是魔鬼的兒女了。凡不行義的，不是出於上帝，不愛他弟兄的，也是如此。
1JOHN|3|11|我們要彼此相愛。這就是你們從起初所聽到的信息。
1JOHN|3|12|不要像 該隱 ；他是屬那邪惡者，殺了自己的弟弟。為甚麼殺了他呢？因為自己的行為是邪惡的，而弟弟的行為是正直的。
1JOHN|3|13|弟兄們，世人若恨你們，不要驚訝。
1JOHN|3|14|我們知道，我們已經出死入生了，因為我們愛弟兄。沒有愛心的，仍住在死中。
1JOHN|3|15|凡恨自己弟兄的，就是殺人的；你們知道，凡殺人的，沒有永生住在他裏面。
1JOHN|3|16|基督為我們捨命，我們從此就知道何為愛；我們也當為弟兄捨命。
1JOHN|3|17|凡有世上財物的，看見弟兄缺乏，卻關閉了惻隱的心，上帝的愛怎能住在他裏面呢？
1JOHN|3|18|孩子們哪，我們相愛，不要只在言語或舌頭上，總要以行為和真誠表現出來。
1JOHN|3|19|從這一點，我們會知道，我們是出於真理的，並且我們在上帝面前可以安心，
1JOHN|3|20|即使我們的心責備自己，上帝比我們的心大，他知道一切。
1JOHN|3|21|親愛的，我們的心若不責備我們，在上帝面前就可以坦然無懼了。
1JOHN|3|22|我們一切所求的，就從他得著，因為我們遵守他的命令，行他所喜悅的事。
1JOHN|3|23|上帝的命令就是：我們要信他兒子耶穌基督的名，並且照他所賜給我們的命令彼此相愛。
1JOHN|3|24|遵守上帝命令的，住在上帝裏面，而上帝也住在他裏面。從這一點，我們知道上帝住在我們裏面，這是由於他所賜給我們的聖靈。
1JOHN|4|1|親愛的，一切的靈不可都信，總要察驗那些靈是否出於上帝，因為有許多假先知已經來到世上。
1JOHN|4|2|凡宣認耶穌基督是成了肉身而來的靈就是出於上帝的，由此你們可以認出上帝的靈來；
1JOHN|4|3|凡不宣認耶穌的靈，不是出於上帝。這是那敵基督者的靈；你們從前聽見他要來，現在他已經在世上了。
1JOHN|4|4|孩子們哪，你們是屬上帝的，並且勝過了假先知，因為那在你們裏面的比那在世界上的更大。
1JOHN|4|5|他們是屬世界的，所以講論世界的事，而世人也聽從他們。
1JOHN|4|6|我們是屬上帝的，認識上帝的就聽從我們；不屬上帝的就不聽從我們。從此我們可以認出真理的靈和錯謬的靈來。
1JOHN|4|7|親愛的，我們要彼此相愛，因為愛是從上帝來的。凡有愛的都是由上帝而生，並且認識上帝。
1JOHN|4|8|沒有愛的就不認識上帝，因為上帝就是愛。
1JOHN|4|9|上帝差他獨一的兒子到世上來，使我們藉著他得生命；由此，上帝對我們的愛就顯明了。
1JOHN|4|10|不是我們愛上帝，而是上帝愛我們，差他的兒子為我們的罪作了贖罪祭；這就是愛。
1JOHN|4|11|親愛的，既然上帝這樣愛我們，我們也要彼此相愛。
1JOHN|4|12|從來沒有人見過上帝，我們若彼此相愛，上帝就住在我們裏面，他的愛在我們裏面得以完滿了。
1JOHN|4|13|因為上帝將他的靈賜給我們，由此我們知道我們是住在他裏面，而他也住在我們裏面。
1JOHN|4|14|父差子作世人的救主，這是我們所看見並且作見證的。
1JOHN|4|15|凡宣認耶穌為上帝兒子的，上帝就住在他裏面，而他也住在上帝裏面。
1JOHN|4|16|我們知道並且深信上帝是愛我們的。 上帝就是愛，住在愛裏面的就是住在上帝裏面；上帝也住在他裏面。
1JOHN|4|17|由此，愛在我們裏面得以完滿：我們可以在審判的日子坦然無懼，因為基督如何，我們在這世上也如何。
1JOHN|4|18|在愛裏沒有懼怕；完滿的愛把懼怕驅逐出去，因為懼怕裏含著懲罰，懼怕的人在愛裏尚未得到完滿。
1JOHN|4|19|我們愛，因為上帝先愛我們。
1JOHN|4|20|人若說「我愛上帝」，卻恨他的弟兄，就是說謊了；不愛他看得見的弟兄，就不能愛看不見的上帝 。
1JOHN|4|21|愛上帝的，也要愛弟兄；這是我們從上帝所受的命令。
1JOHN|5|1|凡信耶穌是基督的，都是從上帝生的；凡愛生他之上帝的，也必愛從上帝生的 。
1JOHN|5|2|我們愛上帝，又實行 他的命令，由此就知道我們愛上帝的兒女了。
1JOHN|5|3|我們遵守上帝的命令，這就是愛他了，而且他的命令並不是難守的。
1JOHN|5|4|因為凡從上帝生的就勝過世界；使我們勝過世界的就是我們的信心。
1JOHN|5|5|勝過世界的是誰呢？不就是那信耶穌是上帝兒子的嗎？
1JOHN|5|6|這藉著水和血而來的，就是耶穌基督，不是單用水，而是用水又用血，並且有聖靈作見證，因為聖靈就是真理。
1JOHN|5|7|作見證的有三：
1JOHN|5|8|就是聖靈、水與血，這三樣也都是一致的。
1JOHN|5|9|既然我們領受人的見證，上帝的見證更該領受 了，因為上帝的見證是為他兒子作的。
1JOHN|5|10|信上帝兒子的，就有這見證在他心裏；不信上帝的，就是把上帝當作說謊的，因為不信上帝為他兒子作的見證。
1JOHN|5|11|這見證就是：上帝賜給我們永生，而這永生是在他兒子裏面的。
1JOHN|5|12|那有上帝兒子的，就有生命；沒有上帝兒子的，就沒有生命。
1JOHN|5|13|我把這些話寫給你們信奉上帝兒子之名的人，要讓你們知道自己有永生。
1JOHN|5|14|我們若照著上帝的旨意祈求，他就垂聽我們；這就是我們對他所存坦然無懼的心。
1JOHN|5|15|既然我們知道他聽我們一切所求的，就知道我們所求於他的，無不得著。
1JOHN|5|16|人若看見弟兄犯了不至於死的罪，就要為他祈求，上帝必將生命賜給他—有些人犯的罪是不至於死的；有的是至於死的罪，我不是說要為這罪祈求。
1JOHN|5|17|一切不義的事都是罪，但也有不至於死的罪。
1JOHN|5|18|我們知道，凡從上帝生的，必不犯罪；從上帝生的那一位，必保守他，那邪惡者無法加害於他。
1JOHN|5|19|我們知道，我們是屬上帝的，而全世界都伏在那邪惡者的權勢之下。
1JOHN|5|20|我們知道，上帝的兒子已經來到，並且將悟性賜給我們，使我們認識那位真實者，我們也在那位真實者裏面，就是在他兒子耶穌基督裏面。這是真神，也是永生。
1JOHN|5|21|孩子們哪，你們要遠避偶像。
