EXOD|1|1|These are the names of the sons of Israel who went to Egypt with Jacob, each with his family:
EXOD|1|2|Reuben, Simeon, Levi and Judah;
EXOD|1|3|Issachar, Zebulun and Benjamin;
EXOD|1|4|Dan and Naphtali; Gad and Asher.
EXOD|1|5|The descendants of Jacob numbered seventy in all; Joseph was already in Egypt.
EXOD|1|6|Now Joseph and all his brothers and all that generation died,
EXOD|1|7|but the Israelites were fruitful and multiplied greatly and became exceedingly numerous, so that the land was filled with them.
EXOD|1|8|Then a new king, who did not know about Joseph, came to power in Egypt.
EXOD|1|9|"Look," he said to his people, "the Israelites have become much too numerous for us.
EXOD|1|10|Come, we must deal shrewdly with them or they will become even more numerous and, if war breaks out, will join our enemies, fight against us and leave the country."
EXOD|1|11|So they put slave masters over them to oppress them with forced labor, and they built Pithom and Rameses as store cities for Pharaoh.
EXOD|1|12|But the more they were oppressed, the more they multiplied and spread; so the Egyptians came to dread the Israelites
EXOD|1|13|and worked them ruthlessly.
EXOD|1|14|They made their lives bitter with hard labor in brick and mortar and with all kinds of work in the fields; in all their hard labor the Egyptians used them ruthlessly.
EXOD|1|15|The king of Egypt said to the Hebrew midwives, whose names were Shiphrah and Puah,
EXOD|1|16|"When you help the Hebrew women in childbirth and observe them on the delivery stool, if it is a boy, kill him; but if it is a girl, let her live."
EXOD|1|17|The midwives, however, feared God and did not do what the king of Egypt had told them to do; they let the boys live.
EXOD|1|18|Then the king of Egypt summoned the midwives and asked them, "Why have you done this? Why have you let the boys live?"
EXOD|1|19|The midwives answered Pharaoh, "Hebrew women are not like Egyptian women; they are vigorous and give birth before the midwives arrive."
EXOD|1|20|So God was kind to the midwives and the people increased and became even more numerous.
EXOD|1|21|And because the midwives feared God, he gave them families of their own.
EXOD|1|22|Then Pharaoh gave this order to all his people: "Every boy that is born you must throw into the Nile, but let every girl live."
EXOD|2|1|Now a man of the house of Levi married a Levite woman,
EXOD|2|2|and she became pregnant and gave birth to a son. When she saw that he was a fine child, she hid him for three months.
EXOD|2|3|But when she could hide him no longer, she got a papyrus basket for him and coated it with tar and pitch. Then she placed the child in it and put it among the reeds along the bank of the Nile.
EXOD|2|4|His sister stood at a distance to see what would happen to him.
EXOD|2|5|Then Pharaoh's daughter went down to the Nile to bathe, and her attendants were walking along the river bank. She saw the basket among the reeds and sent her slave girl to get it.
EXOD|2|6|She opened it and saw the baby. He was crying, and she felt sorry for him. "This is one of the Hebrew babies," she said.
EXOD|2|7|Then his sister asked Pharaoh's daughter, "Shall I go and get one of the Hebrew women to nurse the baby for you?"
EXOD|2|8|"Yes, go," she answered. And the girl went and got the baby's mother.
EXOD|2|9|Pharaoh's daughter said to her, "Take this baby and nurse him for me, and I will pay you." So the woman took the baby and nursed him.
EXOD|2|10|When the child grew older, she took him to Pharaoh's daughter and he became her son. She named him Moses, saying, "I drew him out of the water."
EXOD|2|11|One day, after Moses had grown up, he went out to where his own people were and watched them at their hard labor. He saw an Egyptian beating a Hebrew, one of his own people.
EXOD|2|12|Glancing this way and that and seeing no one, he killed the Egyptian and hid him in the sand.
EXOD|2|13|The next day he went out and saw two Hebrews fighting. He asked the one in the wrong, "Why are you hitting your fellow Hebrew?"
EXOD|2|14|The man said, "Who made you ruler and judge over us? Are you thinking of killing me as you killed the Egyptian?" Then Moses was afraid and thought, "What I did must have become known."
EXOD|2|15|When Pharaoh heard of this, he tried to kill Moses, but Moses fled from Pharaoh and went to live in Midian, where he sat down by a well.
EXOD|2|16|Now a priest of Midian had seven daughters, and they came to draw water and fill the troughs to water their father's flock.
EXOD|2|17|Some shepherds came along and drove them away, but Moses got up and came to their rescue and watered their flock.
EXOD|2|18|When the girls returned to Reuel their father, he asked them, "Why have you returned so early today?"
EXOD|2|19|They answered, "An Egyptian rescued us from the shepherds. He even drew water for us and watered the flock."
EXOD|2|20|"And where is he?" he asked his daughters. "Why did you leave him? Invite him to have something to eat."
EXOD|2|21|Moses agreed to stay with the man, who gave his daughter Zipporah to Moses in marriage.
EXOD|2|22|Zipporah gave birth to a son, and Moses named him Gershom, saying, "I have become an alien in a foreign land."
EXOD|2|23|During that long period, the king of Egypt died. The Israelites groaned in their slavery and cried out, and their cry for help because of their slavery went up to God.
EXOD|2|24|God heard their groaning and he remembered his covenant with Abraham, with Isaac and with Jacob.
EXOD|2|25|So God looked on the Israelites and was concerned about them.
EXOD|3|1|Now Moses was tending the flock of Jethro his father-in-law, the priest of Midian, and he led the flock to the far side of the desert and came to Horeb, the mountain of God.
EXOD|3|2|There the angel of the LORD appeared to him in flames of fire from within a bush. Moses saw that though the bush was on fire it did not burn up.
EXOD|3|3|So Moses thought, "I will go over and see this strange sight-why the bush does not burn up."
EXOD|3|4|When the LORD saw that he had gone over to look, God called to him from within the bush, "Moses! Moses!" And Moses said, "Here I am."
EXOD|3|5|"Do not come any closer," God said. "Take off your sandals, for the place where you are standing is holy ground."
EXOD|3|6|Then he said, "I am the God of your father, the God of Abraham, the God of Isaac and the God of Jacob." At this, Moses hid his face, because he was afraid to look at God.
EXOD|3|7|The LORD said, "I have indeed seen the misery of my people in Egypt. I have heard them crying out because of their slave drivers, and I am concerned about their suffering.
EXOD|3|8|So I have come down to rescue them from the hand of the Egyptians and to bring them up out of that land into a good and spacious land, a land flowing with milk and honey-the home of the Canaanites, Hittites, Amorites, Perizzites, Hivites and Jebusites.
EXOD|3|9|And now the cry of the Israelites has reached me, and I have seen the way the Egyptians are oppressing them.
EXOD|3|10|So now, go. I am sending you to Pharaoh to bring my people the Israelites out of Egypt."
EXOD|3|11|But Moses said to God, "Who am I, that I should go to Pharaoh and bring the Israelites out of Egypt?"
EXOD|3|12|And God said, "I will be with you. And this will be the sign to you that it is I who have sent you: When you have brought the people out of Egypt, you will worship God on this mountain."
EXOD|3|13|Moses said to God, "Suppose I go to the Israelites and say to them, 'The God of your fathers has sent me to you,' and they ask me, 'What is his name?' Then what shall I tell them?"
EXOD|3|14|God said to Moses, "I am who I am. This is what you are to say to the Israelites: 'I AM has sent me to you.'"
EXOD|3|15|God also said to Moses, "Say to the Israelites, 'The LORD, the God of your fathers-the God of Abraham, the God of Isaac and the God of Jacob-has sent me to you.' This is my name forever, the name by which I am to be remembered from generation to generation.
EXOD|3|16|"Go, assemble the elders of Israel and say to them, 'The LORD, the God of your fathers-the God of Abraham, Isaac and Jacob-appeared to me and said: I have watched over you and have seen what has been done to you in Egypt.
EXOD|3|17|And I have promised to bring you up out of your misery in Egypt into the land of the Canaanites, Hittites, Amorites, Perizzites, Hivites and Jebusites-a land flowing with milk and honey.'
EXOD|3|18|"The elders of Israel will listen to you. Then you and the elders are to go to the king of Egypt and say to him, 'The LORD, the God of the Hebrews, has met with us. Let us take a three-day journey into the desert to offer sacrifices to the LORD our God.'
EXOD|3|19|But I know that the king of Egypt will not let you go unless a mighty hand compels him.
EXOD|3|20|So I will stretch out my hand and strike the Egyptians with all the wonders that I will perform among them. After that, he will let you go.
EXOD|3|21|"And I will make the Egyptians favorably disposed toward this people, so that when you leave you will not go empty-handed.
EXOD|3|22|Every woman is to ask her neighbor and any woman living in her house for articles of silver and gold and for clothing, which you will put on your sons and daughters. And so you will plunder the Egyptians."
EXOD|4|1|Moses answered, "What if they do not believe me or listen to me and say, 'The LORD did not appear to you'?"
EXOD|4|2|Then the LORD said to him, "What is that in your hand?A staff," he replied.
EXOD|4|3|The LORD said, "Throw it on the ground." Moses threw it on the ground and it became a snake, and he ran from it.
EXOD|4|4|Then the LORD said to him, "Reach out your hand and take it by the tail." So Moses reached out and took hold of the snake and it turned back into a staff in his hand.
EXOD|4|5|"This," said the LORD, "is so that they may believe that the LORD, the God of their fathers-the God of Abraham, the God of Isaac and the God of Jacob-has appeared to you."
EXOD|4|6|Then the LORD said, "Put your hand inside your cloak." So Moses put his hand into his cloak, and when he took it out, it was leprous, like snow.
EXOD|4|7|"Now put it back into your cloak," he said. So Moses put his hand back into his cloak, and when he took it out, it was restored, like the rest of his flesh.
EXOD|4|8|Then the LORD said, "If they do not believe you or pay attention to the first miraculous sign, they may believe the second.
EXOD|4|9|But if they do not believe these two signs or listen to you, take some water from the Nile and pour it on the dry ground. The water you take from the river will become blood on the ground."
EXOD|4|10|Moses said to the LORD, "O Lord, I have never been eloquent, neither in the past nor since you have spoken to your servant. I am slow of speech and tongue."
EXOD|4|11|The LORD said to him, "Who gave man his mouth? Who makes him deaf or mute? Who gives him sight or makes him blind? Is it not I, the LORD?
EXOD|4|12|Now go; I will help you speak and will teach you what to say."
EXOD|4|13|But Moses said, "O Lord, please send someone else to do it."
EXOD|4|14|Then the LORD's anger burned against Moses and he said, "What about your brother, Aaron the Levite? I know he can speak well. He is already on his way to meet you, and his heart will be glad when he sees you.
EXOD|4|15|You shall speak to him and put words in his mouth; I will help both of you speak and will teach you what to do.
EXOD|4|16|He will speak to the people for you, and it will be as if he were your mouth and as if you were God to him.
EXOD|4|17|But take this staff in your hand so you can perform miraculous signs with it."
EXOD|4|18|Then Moses went back to Jethro his father-in-law and said to him, "Let me go back to my own people in Egypt to see if any of them are still alive." Jethro said, "Go, and I wish you well."
EXOD|4|19|Now the LORD had said to Moses in Midian, "Go back to Egypt, for all the men who wanted to kill you are dead."
EXOD|4|20|So Moses took his wife and sons, put them on a donkey and started back to Egypt. And he took the staff of God in his hand.
EXOD|4|21|The LORD said to Moses, "When you return to Egypt, see that you perform before Pharaoh all the wonders I have given you the power to do. But I will harden his heart so that he will not let the people go.
EXOD|4|22|Then say to Pharaoh, 'This is what the LORD says: Israel is my firstborn son,
EXOD|4|23|and I told you, "Let my son go, so he may worship me." But you refused to let him go; so I will kill your firstborn son.'"
EXOD|4|24|At a lodging place on the way, the LORD met {Moses} and was about to kill him.
EXOD|4|25|But Zipporah took a flint knife, cut off her son's foreskin and touched {Moses'} feet with it. "Surely you are a bridegroom of blood to me," she said.
EXOD|4|26|So the LORD let him alone. (At that time she said "bridegroom of blood," referring to circumcision.)
EXOD|4|27|The LORD said to Aaron, "Go into the desert to meet Moses." So he met Moses at the mountain of God and kissed him.
EXOD|4|28|Then Moses told Aaron everything the LORD had sent him to say, and also about all the miraculous signs he had commanded him to perform.
EXOD|4|29|Moses and Aaron brought together all the elders of the Israelites,
EXOD|4|30|and Aaron told them everything the LORD had said to Moses. He also performed the signs before the people,
EXOD|4|31|and they believed. And when they heard that the LORD was concerned about them and had seen their misery, they bowed down and worshiped.
EXOD|5|1|Afterward Moses and Aaron went to Pharaoh and said, "This is what the LORD, the God of Israel, says: 'Let my people go, so that they may hold a festival to me in the desert.'"
EXOD|5|2|Pharaoh said, "Who is the LORD, that I should obey him and let Israel go? I do not know the LORD and I will not let Israel go."
EXOD|5|3|Then they said, "The God of the Hebrews has met with us. Now let us take a three-day journey into the desert to offer sacrifices to the LORD our God, or he may strike us with plagues or with the sword."
EXOD|5|4|But the king of Egypt said, "Moses and Aaron, why are you taking the people away from their labor? Get back to your work!"
EXOD|5|5|Then Pharaoh said, "Look, the people of the land are now numerous, and you are stopping them from working."
EXOD|5|6|That same day Pharaoh gave this order to the slave drivers and foremen in charge of the people:
EXOD|5|7|"You are no longer to supply the people with straw for making bricks; let them go and gather their own straw.
EXOD|5|8|But require them to make the same number of bricks as before; don't reduce the quota. They are lazy; that is why they are crying out, 'Let us go and sacrifice to our God.'
EXOD|5|9|Make the work harder for the men so that they keep working and pay no attention to lies."
EXOD|5|10|Then the slave drivers and the foremen went out and said to the people, "This is what Pharaoh says: 'I will not give you any more straw.
EXOD|5|11|Go and get your own straw wherever you can find it, but your work will not be reduced at all.'"
EXOD|5|12|So the people scattered all over Egypt to gather stubble to use for straw.
EXOD|5|13|The slave drivers kept pressing them, saying, "Complete the work required of you for each day, just as when you had straw."
EXOD|5|14|The Israelite foremen appointed by Pharaoh's slave drivers were beaten and were asked, "Why didn't you meet your quota of bricks yesterday or today, as before?"
EXOD|5|15|Then the Israelite foremen went and appealed to Pharaoh: "Why have you treated your servants this way?
EXOD|5|16|Your servants are given no straw, yet we are told, 'Make bricks!' Your servants are being beaten, but the fault is with your own people."
EXOD|5|17|Pharaoh said, "Lazy, that's what you are-lazy! That is why you keep saying, 'Let us go and sacrifice to the LORD.'
EXOD|5|18|Now get to work. You will not be given any straw, yet you must produce your full quota of bricks."
EXOD|5|19|The Israelite foremen realized they were in trouble when they were told, "You are not to reduce the number of bricks required of you for each day."
EXOD|5|20|When they left Pharaoh, they found Moses and Aaron waiting to meet them,
EXOD|5|21|and they said, "May the LORD look upon you and judge you! You have made us a stench to Pharaoh and his officials and have put a sword in their hand to kill us."
EXOD|5|22|Moses returned to the LORD and said, "O Lord, why have you brought trouble upon this people? Is this why you sent me?
EXOD|5|23|Ever since I went to Pharaoh to speak in your name, he has brought trouble upon this people, and you have not rescued your people at all."
EXOD|6|1|Then the LORD said to Moses, "Now you will see what I will do to Pharaoh: Because of my mighty hand he will let them go; because of my mighty hand he will drive them out of his country."
EXOD|6|2|God also said to Moses, "I am the LORD.
EXOD|6|3|I appeared to Abraham, to Isaac and to Jacob as God Almighty, but by my name the LORD I did not make myself known to them.
EXOD|6|4|I also established my covenant with them to give them the land of Canaan, where they lived as aliens.
EXOD|6|5|Moreover, I have heard the groaning of the Israelites, whom the Egyptians are enslaving, and I have remembered my covenant.
EXOD|6|6|"Therefore, say to the Israelites: 'I am the LORD, and I will bring you out from under the yoke of the Egyptians. I will free you from being slaves to them, and I will redeem you with an outstretched arm and with mighty acts of judgment.
EXOD|6|7|I will take you as my own people, and I will be your God. Then you will know that I am the LORD your God, who brought you out from under the yoke of the Egyptians.
EXOD|6|8|And I will bring you to the land I swore with uplifted hand to give to Abraham, to Isaac and to Jacob. I will give it to you as a possession. I am the LORD.'"
EXOD|6|9|Moses reported this to the Israelites, but they did not listen to him because of their discouragement and cruel bondage.
EXOD|6|10|Then the LORD said to Moses,
EXOD|6|11|"Go, tell Pharaoh king of Egypt to let the Israelites go out of his country."
EXOD|6|12|But Moses said to the LORD, "If the Israelites will not listen to me, why would Pharaoh listen to me, since I speak with faltering lips?"
EXOD|6|13|Now the LORD spoke to Moses and Aaron about the Israelites and Pharaoh king of Egypt, and he commanded them to bring the Israelites out of Egypt.
EXOD|6|14|These were the heads of their families: The sons of Reuben the firstborn son of Israel were Hanoch and Pallu, Hezron and Carmi. These were the clans of Reuben.
EXOD|6|15|The sons of Simeon were Jemuel, Jamin, Ohad, Jakin, Zohar and Shaul the son of a Canaanite woman. These were the clans of Simeon.
EXOD|6|16|These were the names of the sons of Levi according to their records: Gershon, Kohath and Merari. Levi lived 137 years.
EXOD|6|17|The sons of Gershon, by clans, were Libni and Shimei.
EXOD|6|18|The sons of Kohath were Amram, Izhar, Hebron and Uzziel. Kohath lived 133 years.
EXOD|6|19|The sons of Merari were Mahli and Mushi. These were the clans of Levi according to their records.
EXOD|6|20|Amram married his father's sister Jochebed, who bore him Aaron and Moses. Amram lived 137 years.
EXOD|6|21|The sons of Izhar were Korah, Nepheg and Zicri.
EXOD|6|22|The sons of Uzziel were Mishael, Elzaphan and Sithri.
EXOD|6|23|Aaron married Elisheba, daughter of Amminadab and sister of Nahshon, and she bore him Nadab and Abihu, Eleazar and Ithamar.
EXOD|6|24|The sons of Korah were Assir, Elkanah and Abiasaph. These were the Korahite clans.
EXOD|6|25|Eleazar son of Aaron married one of the daughters of Putiel, and she bore him Phinehas. These were the heads of the Levite families, clan by clan.
EXOD|6|26|It was this same Aaron and Moses to whom the LORD said, "Bring the Israelites out of Egypt by their divisions."
EXOD|6|27|They were the ones who spoke to Pharaoh king of Egypt about bringing the Israelites out of Egypt. It was the same Moses and Aaron.
EXOD|6|28|Now when the LORD spoke to Moses in Egypt,
EXOD|6|29|he said to him, "I am the LORD. Tell Pharaoh king of Egypt everything I tell you."
EXOD|6|30|But Moses said to the LORD, "Since I speak with faltering lips, why would Pharaoh listen to me?"
EXOD|7|1|Then the LORD said to Moses, "See, I have made you like God to Pharaoh, and your brother Aaron will be your prophet.
EXOD|7|2|You are to say everything I command you, and your brother Aaron is to tell Pharaoh to let the Israelites go out of his country.
EXOD|7|3|But I will harden Pharaoh's heart, and though I multiply my miraculous signs and wonders in Egypt,
EXOD|7|4|he will not listen to you. Then I will lay my hand on Egypt and with mighty acts of judgment I will bring out my divisions, my people the Israelites.
EXOD|7|5|And the Egyptians will know that I am the LORD when I stretch out my hand against Egypt and bring the Israelites out of it."
EXOD|7|6|Moses and Aaron did just as the LORD commanded them.
EXOD|7|7|Moses was eighty years old and Aaron eighty-three when they spoke to Pharaoh.
EXOD|7|8|The LORD said to Moses and Aaron,
EXOD|7|9|"When Pharaoh says to you, 'Perform a miracle,' then say to Aaron, 'Take your staff and throw it down before Pharaoh,' and it will become a snake."
EXOD|7|10|So Moses and Aaron went to Pharaoh and did just as the LORD commanded. Aaron threw his staff down in front of Pharaoh and his officials, and it became a snake.
EXOD|7|11|Pharaoh then summoned wise men and sorcerers, and the Egyptian magicians also did the same things by their secret arts:
EXOD|7|12|Each one threw down his staff and it became a snake. But Aaron's staff swallowed up their staffs.
EXOD|7|13|Yet Pharaoh's heart became hard and he would not listen to them, just as the LORD had said.
EXOD|7|14|Then the LORD said to Moses, "Pharaoh's heart is unyielding; he refuses to let the people go.
EXOD|7|15|Go to Pharaoh in the morning as he goes out to the water. Wait on the bank of the Nile to meet him, and take in your hand the staff that was changed into a snake.
EXOD|7|16|Then say to him, 'The LORD, the God of the Hebrews, has sent me to say to you: Let my people go, so that they may worship me in the desert. But until now you have not listened.
EXOD|7|17|This is what the LORD says: By this you will know that I am the LORD: With the staff that is in my hand I will strike the water of the Nile, and it will be changed into blood.
EXOD|7|18|The fish in the Nile will die, and the river will stink; the Egyptians will not be able to drink its water.'"
EXOD|7|19|The LORD said to Moses, "Tell Aaron, 'Take your staff and stretch out your hand over the waters of Egypt-over the streams and canals, over the ponds and all the reservoirs'-and they will turn to blood. Blood will be everywhere in Egypt, even in the wooden buckets and stone jars."
EXOD|7|20|Moses and Aaron did just as the LORD had commanded. He raised his staff in the presence of Pharaoh and his officials and struck the water of the Nile, and all the water was changed into blood.
EXOD|7|21|The fish in the Nile died, and the river smelled so bad that the Egyptians could not drink its water. Blood was everywhere in Egypt.
EXOD|7|22|But the Egyptian magicians did the same things by their secret arts, and Pharaoh's heart became hard; he would not listen to Moses and Aaron, just as the LORD had said.
EXOD|7|23|Instead, he turned and went into his palace, and did not take even this to heart.
EXOD|7|24|And all the Egyptians dug along the Nile to get drinking water, because they could not drink the water of the river.
EXOD|7|25|Seven days passed after the LORD struck the Nile.
EXOD|8|1|Then the LORD said to Moses, "Go to Pharaoh and say to him, 'This is what the LORD says: Let my people go, so that they may worship me.
EXOD|8|2|If you refuse to let them go, I will plague your whole country with frogs.
EXOD|8|3|The Nile will teem with frogs. They will come up into your palace and your bedroom and onto your bed, into the houses of your officials and on your people, and into your ovens and kneading troughs.
EXOD|8|4|The frogs will go up on you and your people and all your officials.'"
EXOD|8|5|Then the LORD said to Moses, "Tell Aaron, 'Stretch out your hand with your staff over the streams and canals and ponds, and make frogs come up on the land of Egypt.'"
EXOD|8|6|So Aaron stretched out his hand over the waters of Egypt, and the frogs came up and covered the land.
EXOD|8|7|But the magicians did the same things by their secret arts; they also made frogs come up on the land of Egypt.
EXOD|8|8|Pharaoh summoned Moses and Aaron and said, "Pray to the LORD to take the frogs away from me and my people, and I will let your people go to offer sacrifices to the LORD."
EXOD|8|9|Moses said to Pharaoh, "I leave to you the honor of setting the time for me to pray for you and your officials and your people that you and your houses may be rid of the frogs, except for those that remain in the Nile."
EXOD|8|10|"Tomorrow," Pharaoh said. Moses replied, "It will be as you say, so that you may know there is no one like the LORD our God.
EXOD|8|11|The frogs will leave you and your houses, your officials and your people; they will remain only in the Nile."
EXOD|8|12|After Moses and Aaron left Pharaoh, Moses cried out to the LORD about the frogs he had brought on Pharaoh.
EXOD|8|13|And the LORD did what Moses asked. The frogs died in the houses, in the courtyards and in the fields.
EXOD|8|14|They were piled into heaps, and the land reeked of them.
EXOD|8|15|But when Pharaoh saw that there was relief, he hardened his heart and would not listen to Moses and Aaron, just as the LORD had said.
EXOD|8|16|Then the LORD said to Moses, "Tell Aaron, 'Stretch out your staff and strike the dust of the ground,' and throughout the land of Egypt the dust will become gnats."
EXOD|8|17|They did this, and when Aaron stretched out his hand with the staff and struck the dust of the ground, gnats came upon men and animals. All the dust throughout the land of Egypt became gnats.
EXOD|8|18|But when the magicians tried to produce gnats by their secret arts, they could not. And the gnats were on men and animals.
EXOD|8|19|The magicians said to Pharaoh, "This is the finger of God." But Pharaoh's heart was hard and he would not listen, just as the LORD had said.
EXOD|8|20|Then the LORD said to Moses, "Get up early in the morning and confront Pharaoh as he goes to the water and say to him, 'This is what the LORD says: Let my people go, so that they may worship me.
EXOD|8|21|If you do not let my people go, I will send swarms of flies on you and your officials, on your people and into your houses. The houses of the Egyptians will be full of flies, and even the ground where they are.
EXOD|8|22|"'But on that day I will deal differently with the land of Goshen, where my people live; no swarms of flies will be there, so that you will know that I, the LORD, am in this land.
EXOD|8|23|I will make a distinction between my people and your people. This miraculous sign will occur tomorrow.'"
EXOD|8|24|And the LORD did this. Dense swarms of flies poured into Pharaoh's palace and into the houses of his officials, and throughout Egypt the land was ruined by the flies.
EXOD|8|25|Then Pharaoh summoned Moses and Aaron and said, "Go, sacrifice to your God here in the land."
EXOD|8|26|But Moses said, "That would not be right. The sacrifices we offer the LORD our God would be detestable to the Egyptians. And if we offer sacrifices that are detestable in their eyes, will they not stone us?
EXOD|8|27|We must take a three-day journey into the desert to offer sacrifices to the LORD our God, as he commands us."
EXOD|8|28|Pharaoh said, "I will let you go to offer sacrifices to the LORD your God in the desert, but you must not go very far. Now pray for me."
EXOD|8|29|Moses answered, "As soon as I leave you, I will pray to the LORD, and tomorrow the flies will leave Pharaoh and his officials and his people. Only be sure that Pharaoh does not act deceitfully again by not letting the people go to offer sacrifices to the LORD."
EXOD|8|30|Then Moses left Pharaoh and prayed to the LORD,
EXOD|8|31|and the LORD did what Moses asked: The flies left Pharaoh and his officials and his people; not a fly remained.
EXOD|8|32|But this time also Pharaoh hardened his heart and would not let the people go.
EXOD|9|1|Then the LORD said to Moses, "Go to Pharaoh and say to him, 'This is what the LORD, the God of the Hebrews, says: "Let my people go, so that they may worship me."
EXOD|9|2|If you refuse to let them go and continue to hold them back,
EXOD|9|3|the hand of the LORD will bring a terrible plague on your livestock in the field-on your horses and donkeys and camels and on your cattle and sheep and goats.
EXOD|9|4|But the LORD will make a distinction between the livestock of Israel and that of Egypt, so that no animal belonging to the Israelites will die.'"
EXOD|9|5|The LORD set a time and said, "Tomorrow the LORD will do this in the land."
EXOD|9|6|And the next day the LORD did it: All the livestock of the Egyptians died, but not one animal belonging to the Israelites died.
EXOD|9|7|Pharaoh sent men to investigate and found that not even one of the animals of the Israelites had died. Yet his heart was unyielding and he would not let the people go.
EXOD|9|8|Then the LORD said to Moses and Aaron, "Take handfuls of soot from a furnace and have Moses toss it into the air in the presence of Pharaoh.
EXOD|9|9|It will become fine dust over the whole land of Egypt, and festering boils will break out on men and animals throughout the land."
EXOD|9|10|So they took soot from a furnace and stood before Pharaoh. Moses tossed it into the air, and festering boils broke out on men and animals.
EXOD|9|11|The magicians could not stand before Moses because of the boils that were on them and on all the Egyptians.
EXOD|9|12|But the LORD hardened Pharaoh's heart and he would not listen to Moses and Aaron, just as the LORD had said to Moses.
EXOD|9|13|Then the LORD said to Moses, "Get up early in the morning, confront Pharaoh and say to him, 'This is what the LORD, the God of the Hebrews, says: Let my people go, so that they may worship me,
EXOD|9|14|or this time I will send the full force of my plagues against you and against your officials and your people, so you may know that there is no one like me in all the earth.
EXOD|9|15|For by now I could have stretched out my hand and struck you and your people with a plague that would have wiped you off the earth.
EXOD|9|16|But I have raised you up for this very purpose, that I might show you my power and that my name might be proclaimed in all the earth.
EXOD|9|17|You still set yourself against my people and will not let them go.
EXOD|9|18|Therefore, at this time tomorrow I will send the worst hailstorm that has ever fallen on Egypt, from the day it was founded till now.
EXOD|9|19|Give an order now to bring your livestock and everything you have in the field to a place of shelter, because the hail will fall on every man and animal that has not been brought in and is still out in the field, and they will die.'"
EXOD|9|20|Those officials of Pharaoh who feared the word of the LORD hurried to bring their slaves and their livestock inside.
EXOD|9|21|But those who ignored the word of the LORD left their slaves and livestock in the field.
EXOD|9|22|Then the LORD said to Moses, "Stretch out your hand toward the sky so that hail will fall all over Egypt-on men and animals and on everything growing in the fields of Egypt."
EXOD|9|23|When Moses stretched out his staff toward the sky, the LORD sent thunder and hail, and lightning flashed down to the ground. So the LORD rained hail on the land of Egypt;
EXOD|9|24|hail fell and lightning flashed back and forth. It was the worst storm in all the land of Egypt since it had become a nation.
EXOD|9|25|Throughout Egypt hail struck everything in the fields-both men and animals; it beat down everything growing in the fields and stripped every tree.
EXOD|9|26|The only place it did not hail was the land of Goshen, where the Israelites were.
EXOD|9|27|Then Pharaoh summoned Moses and Aaron. "This time I have sinned," he said to them. "The LORD is in the right, and I and my people are in the wrong.
EXOD|9|28|Pray to the LORD, for we have had enough thunder and hail. I will let you go; you don't have to stay any longer."
EXOD|9|29|Moses replied, "When I have gone out of the city, I will spread out my hands in prayer to the LORD. The thunder will stop and there will be no more hail, so you may know that the earth is the LORD's.
EXOD|9|30|But I know that you and your officials still do not fear the LORD God."
EXOD|9|31|(The flax and barley were destroyed, since the barley had headed and the flax was in bloom.
EXOD|9|32|The wheat and spelt, however, were not destroyed, because they ripen later.)
EXOD|9|33|Then Moses left Pharaoh and went out of the city. He spread out his hands toward the LORD; the thunder and hail stopped, and the rain no longer poured down on the land.
EXOD|9|34|When Pharaoh saw that the rain and hail and thunder had stopped, he sinned again: He and his officials hardened their hearts.
EXOD|9|35|So Pharaoh's heart was hard and he would not let the Israelites go, just as the LORD had said through Moses.
EXOD|10|1|Then the LORD said to Moses, "Go to Pharaoh, for I have hardened his heart and the hearts of his officials so that I may perform these miraculous signs of mine among them
EXOD|10|2|that you may tell your children and grandchildren how I dealt harshly with the Egyptians and how I performed my signs among them, and that you may know that I am the LORD."
EXOD|10|3|So Moses and Aaron went to Pharaoh and said to him, "This is what the LORD, the God of the Hebrews, says: 'How long will you refuse to humble yourself before me? Let my people go, so that they may worship me.
EXOD|10|4|If you refuse to let them go, I will bring locusts into your country tomorrow.
EXOD|10|5|They will cover the face of the ground so that it cannot be seen. They will devour what little you have left after the hail, including every tree that is growing in your fields.
EXOD|10|6|They will fill your houses and those of all your officials and all the Egyptians-something neither your fathers nor your forefathers have ever seen from the day they settled in this land till now.'" Then Moses turned and left Pharaoh.
EXOD|10|7|Pharaoh's officials said to him, "How long will this man be a snare to us? Let the people go, so that they may worship the LORD their God. Do you not yet realize that Egypt is ruined?"
EXOD|10|8|Then Moses and Aaron were brought back to Pharaoh. "Go, worship the LORD your God," he said. "But just who will be going?"
EXOD|10|9|Moses answered, "We will go with our young and old, with our sons and daughters, and with our flocks and herds, because we are to celebrate a festival to the LORD."
EXOD|10|10|Pharaoh said, "The LORD be with you-if I let you go, along with your women and children! Clearly you are bent on evil.
EXOD|10|11|No! Have only the men go; and worship the LORD, since that's what you have been asking for." Then Moses and Aaron were driven out of Pharaoh's presence.
EXOD|10|12|And the LORD said to Moses, "Stretch out your hand over Egypt so that locusts will swarm over the land and devour everything growing in the fields, everything left by the hail."
EXOD|10|13|So Moses stretched out his staff over Egypt, and the LORD made an east wind blow across the land all that day and all that night. By morning the wind had brought the locusts;
EXOD|10|14|they invaded all Egypt and settled down in every area of the country in great numbers. Never before had there been such a plague of locusts, nor will there ever be again.
EXOD|10|15|They covered all the ground until it was black. They devoured all that was left after the hail-everything growing in the fields and the fruit on the trees. Nothing green remained on tree or plant in all the land of Egypt.
EXOD|10|16|Pharaoh quickly summoned Moses and Aaron and said, "I have sinned against the LORD your God and against you.
EXOD|10|17|Now forgive my sin once more and pray to the LORD your God to take this deadly plague away from me."
EXOD|10|18|Moses then left Pharaoh and prayed to the LORD.
EXOD|10|19|And the LORD changed the wind to a very strong west wind, which caught up the locusts and carried them into the Red Sea. Not a locust was left anywhere in Egypt.
EXOD|10|20|But the LORD hardened Pharaoh's heart, and he would not let the Israelites go.
EXOD|10|21|Then the LORD said to Moses, "Stretch out your hand toward the sky so that darkness will spread over Egypt-darkness that can be felt."
EXOD|10|22|So Moses stretched out his hand toward the sky, and total darkness covered all Egypt for three days.
EXOD|10|23|No one could see anyone else or leave his place for three days. Yet all the Israelites had light in the places where they lived.
EXOD|10|24|Then Pharaoh summoned Moses and said, "Go, worship the LORD. Even your women and children may go with you; only leave your flocks and herds behind."
EXOD|10|25|But Moses said, "You must allow us to have sacrifices and burnt offerings to present to the LORD our God.
EXOD|10|26|Our livestock too must go with us; not a hoof is to be left behind. We have to use some of them in worshiping the LORD our God, and until we get there we will not know what we are to use to worship the LORD."
EXOD|10|27|But the LORD hardened Pharaoh's heart, and he was not willing to let them go.
EXOD|10|28|Pharaoh said to Moses, "Get out of my sight! Make sure you do not appear before me again! The day you see my face you will die."
EXOD|10|29|"Just as you say," Moses replied, "I will never appear before you again."
EXOD|11|1|Now the LORD had said to Moses, "I will bring one more plague on Pharaoh and on Egypt. After that, he will let you go from here, and when he does, he will drive you out completely.
EXOD|11|2|Tell the people that men and women alike are to ask their neighbors for articles of silver and gold."
EXOD|11|3|(The LORD made the Egyptians favorably disposed toward the people, and Moses himself was highly regarded in Egypt by Pharaoh's officials and by the people.)
EXOD|11|4|So Moses said, "This is what the LORD says: 'About midnight I will go throughout Egypt.
EXOD|11|5|Every firstborn son in Egypt will die, from the firstborn son of Pharaoh, who sits on the throne, to the firstborn son of the slave girl, who is at her hand mill, and all the firstborn of the cattle as well.
EXOD|11|6|There will be loud wailing throughout Egypt-worse than there has ever been or ever will be again.
EXOD|11|7|But among the Israelites not a dog will bark at any man or animal.' Then you will know that the LORD makes a distinction between Egypt and Israel.
EXOD|11|8|All these officials of yours will come to me, bowing down before me and saying, 'Go, you and all the people who follow you!' After that I will leave." Then Moses, hot with anger, left Pharaoh.
EXOD|11|9|The LORD had said to Moses, "Pharaoh will refuse to listen to you-so that my wonders may be multiplied in Egypt."
EXOD|11|10|Moses and Aaron performed all these wonders before Pharaoh, but the LORD hardened Pharaoh's heart, and he would not let the Israelites go out of his country.
EXOD|12|1|The LORD said to Moses and Aaron in Egypt,
EXOD|12|2|"This month is to be for you the first month, the first month of your year.
EXOD|12|3|Tell the whole community of Israel that on the tenth day of this month each man is to take a lamb for his family, one for each household.
EXOD|12|4|If any household is too small for a whole lamb, they must share one with their nearest neighbor, having taken into account the number of people there are. You are to determine the amount of lamb needed in accordance with what each person will eat.
EXOD|12|5|The animals you choose must be year-old males without defect, and you may take them from the sheep or the goats.
EXOD|12|6|Take care of them until the fourteenth day of the month, when all the people of the community of Israel must slaughter them at twilight.
EXOD|12|7|Then they are to take some of the blood and put it on the sides and tops of the doorframes of the houses where they eat the lambs.
EXOD|12|8|That same night they are to eat the meat roasted over the fire, along with bitter herbs, and bread made without yeast.
EXOD|12|9|Do not eat the meat raw or cooked in water, but roast it over the fire-head, legs and inner parts.
EXOD|12|10|Do not leave any of it till morning; if some is left till morning, you must burn it.
EXOD|12|11|This is how you are to eat it: with your cloak tucked into your belt, your sandals on your feet and your staff in your hand. Eat it in haste; it is the LORD's Passover.
EXOD|12|12|"On that same night I will pass through Egypt and strike down every firstborn-both men and animals-and I will bring judgment on all the gods of Egypt. I am the LORD.
EXOD|12|13|The blood will be a sign for you on the houses where you are; and when I see the blood, I will pass over you. No destructive plague will touch you when I strike Egypt.
EXOD|12|14|"This is a day you are to commemorate; for the generations to come you shall celebrate it as a festival to the LORD -a lasting ordinance.
EXOD|12|15|For seven days you are to eat bread made without yeast. On the first day remove the yeast from your houses, for whoever eats anything with yeast in it from the first day through the seventh must be cut off from Israel.
EXOD|12|16|On the first day hold a sacred assembly, and another one on the seventh day. Do no work at all on these days, except to prepare food for everyone to eat-that is all you may do.
EXOD|12|17|"Celebrate the Feast of Unleavened Bread, because it was on this very day that I brought your divisions out of Egypt. Celebrate this day as a lasting ordinance for the generations to come.
EXOD|12|18|In the first month you are to eat bread made without yeast, from the evening of the fourteenth day until the evening of the twenty-first day.
EXOD|12|19|For seven days no yeast is to be found in your houses. And whoever eats anything with yeast in it must be cut off from the community of Israel, whether he is an alien or native-born.
EXOD|12|20|Eat nothing made with yeast. Wherever you live, you must eat unleavened bread."
EXOD|12|21|Then Moses summoned all the elders of Israel and said to them, "Go at once and select the animals for your families and slaughter the Passover lamb.
EXOD|12|22|Take a bunch of hyssop, dip it into the blood in the basin and put some of the blood on the top and on both sides of the doorframe. Not one of you shall go out the door of his house until morning.
EXOD|12|23|When the LORD goes through the land to strike down the Egyptians, he will see the blood on the top and sides of the doorframe and will pass over that doorway, and he will not permit the destroyer to enter your houses and strike you down.
EXOD|12|24|"Obey these instructions as a lasting ordinance for you and your descendants.
EXOD|12|25|When you enter the land that the LORD will give you as he promised, observe this ceremony.
EXOD|12|26|And when your children ask you, 'What does this ceremony mean to you?'
EXOD|12|27|then tell them, 'It is the Passover sacrifice to the LORD, who passed over the houses of the Israelites in Egypt and spared our homes when he struck down the Egyptians.'" Then the people bowed down and worshiped.
EXOD|12|28|The Israelites did just what the LORD commanded Moses and Aaron.
EXOD|12|29|At midnight the LORD struck down all the firstborn in Egypt, from the firstborn of Pharaoh, who sat on the throne, to the firstborn of the prisoner, who was in the dungeon, and the firstborn of all the livestock as well.
EXOD|12|30|Pharaoh and all his officials and all the Egyptians got up during the night, and there was loud wailing in Egypt, for there was not a house without someone dead.
EXOD|12|31|During the night Pharaoh summoned Moses and Aaron and said, "Up! Leave my people, you and the Israelites! Go, worship the LORD as you have requested.
EXOD|12|32|Take your flocks and herds, as you have said, and go. And also bless me."
EXOD|12|33|The Egyptians urged the people to hurry and leave the country. "For otherwise," they said, "we will all die!"
EXOD|12|34|So the people took their dough before the yeast was added, and carried it on their shoulders in kneading troughs wrapped in clothing.
EXOD|12|35|The Israelites did as Moses instructed and asked the Egyptians for articles of silver and gold and for clothing.
EXOD|12|36|The LORD had made the Egyptians favorably disposed toward the people, and they gave them what they asked for; so they plundered the Egyptians.
EXOD|12|37|The Israelites journeyed from Rameses to Succoth. There were about six hundred thousand men on foot, besides women and children.
EXOD|12|38|Many other people went up with them, as well as large droves of livestock, both flocks and herds.
EXOD|12|39|With the dough they had brought from Egypt, they baked cakes of unleavened bread. The dough was without yeast because they had been driven out of Egypt and did not have time to prepare food for themselves.
EXOD|12|40|Now the length of time the Israelite people lived in Egypt was 430 years.
EXOD|12|41|At the end of the 430 years, to the very day, all the LORD's divisions left Egypt.
EXOD|12|42|Because the LORD kept vigil that night to bring them out of Egypt, on this night all the Israelites are to keep vigil to honor the LORD for the generations to come.
EXOD|12|43|The LORD said to Moses and Aaron, "These are the regulations for the Passover: "No foreigner is to eat of it.
EXOD|12|44|Any slave you have bought may eat of it after you have circumcised him,
EXOD|12|45|but a temporary resident and a hired worker may not eat of it.
EXOD|12|46|"It must be eaten inside one house; take none of the meat outside the house. Do not break any of the bones.
EXOD|12|47|The whole community of Israel must celebrate it.
EXOD|12|48|"An alien living among you who wants to celebrate the LORD's Passover must have all the males in his household circumcised; then he may take part like one born in the land. No uncircumcised male may eat of it.
EXOD|12|49|The same law applies to the native-born and to the alien living among you."
EXOD|12|50|All the Israelites did just what the LORD had commanded Moses and Aaron.
EXOD|12|51|And on that very day the LORD brought the Israelites out of Egypt by their divisions.
EXOD|13|1|The LORD said to Moses,
EXOD|13|2|"Consecrate to me every firstborn male. The first offspring of every womb among the Israelites belongs to me, whether man or animal."
EXOD|13|3|Then Moses said to the people, "Commemorate this day, the day you came out of Egypt, out of the land of slavery, because the LORD brought you out of it with a mighty hand. Eat nothing containing yeast.
EXOD|13|4|Today, in the month of Abib, you are leaving.
EXOD|13|5|When the LORD brings you into the land of the Canaanites, Hittites, Amorites, Hivites and Jebusites-the land he swore to your forefathers to give you, a land flowing with milk and honey-you are to observe this ceremony in this month:
EXOD|13|6|For seven days eat bread made without yeast and on the seventh day hold a festival to the LORD.
EXOD|13|7|Eat unleavened bread during those seven days; nothing with yeast in it is to be seen among you, nor shall any yeast be seen anywhere within your borders.
EXOD|13|8|On that day tell your son, 'I do this because of what the LORD did for me when I came out of Egypt.'
EXOD|13|9|This observance will be for you like a sign on your hand and a reminder on your forehead that the law of the LORD is to be on your lips. For the LORD brought you out of Egypt with his mighty hand.
EXOD|13|10|You must keep this ordinance at the appointed time year after year.
EXOD|13|11|"After the LORD brings you into the land of the Canaanites and gives it to you, as he promised on oath to you and your forefathers,
EXOD|13|12|you are to give over to the LORD the first offspring of every womb. All the firstborn males of your livestock belong to the LORD.
EXOD|13|13|Redeem with a lamb every firstborn donkey, but if you do not redeem it, break its neck. Redeem every firstborn among your sons.
EXOD|13|14|"In days to come, when your son asks you, 'What does this mean?' say to him, 'With a mighty hand the LORD brought us out of Egypt, out of the land of slavery.
EXOD|13|15|When Pharaoh stubbornly refused to let us go, the LORD killed every firstborn in Egypt, both man and animal. This is why I sacrifice to the LORD the first male offspring of every womb and redeem each of my firstborn sons.'
EXOD|13|16|And it will be like a sign on your hand and a symbol on your forehead that the LORD brought us out of Egypt with his mighty hand."
EXOD|13|17|When Pharaoh let the people go, God did not lead them on the road through the Philistine country, though that was shorter. For God said, "If they face war, they might change their minds and return to Egypt."
EXOD|13|18|So God led the people around by the desert road toward the Red Sea. The Israelites went up out of Egypt armed for battle.
EXOD|13|19|Moses took the bones of Joseph with him because Joseph had made the sons of Israel swear an oath. He had said, "God will surely come to your aid, and then you must carry my bones up with you from this place."
EXOD|13|20|After leaving Succoth they camped at Etham on the edge of the desert.
EXOD|13|21|By day the LORD went ahead of them in a pillar of cloud to guide them on their way and by night in a pillar of fire to give them light, so that they could travel by day or night.
EXOD|13|22|Neither the pillar of cloud by day nor the pillar of fire by night left its place in front of the people.
EXOD|14|1|Then the LORD said to Moses,
EXOD|14|2|"Tell the Israelites to turn back and encamp near Pi Hahiroth, between Migdol and the sea. They are to encamp by the sea, directly opposite Baal Zephon.
EXOD|14|3|Pharaoh will think, 'The Israelites are wandering around the land in confusion, hemmed in by the desert.'
EXOD|14|4|And I will harden Pharaoh's heart, and he will pursue them. But I will gain glory for myself through Pharaoh and all his army, and the Egyptians will know that I am the LORD." So the Israelites did this.
EXOD|14|5|When the king of Egypt was told that the people had fled, Pharaoh and his officials changed their minds about them and said, "What have we done? We have let the Israelites go and have lost their services!"
EXOD|14|6|So he had his chariot made ready and took his army with him.
EXOD|14|7|He took six hundred of the best chariots, along with all the other chariots of Egypt, with officers over all of them.
EXOD|14|8|The LORD hardened the heart of Pharaoh king of Egypt, so that he pursued the Israelites, who were marching out boldly.
EXOD|14|9|The Egyptians-all Pharaoh's horses and chariots, horsemen and troops-pursued the Israelites and overtook them as they camped by the sea near Pi Hahiroth, opposite Baal Zephon.
EXOD|14|10|As Pharaoh approached, the Israelites looked up, and there were the Egyptians, marching after them. They were terrified and cried out to the LORD.
EXOD|14|11|They said to Moses, "Was it because there were no graves in Egypt that you brought us to the desert to die? What have you done to us by bringing us out of Egypt?
EXOD|14|12|Didn't we say to you in Egypt, 'Leave us alone; let us serve the Egyptians'? It would have been better for us to serve the Egyptians than to die in the desert!"
EXOD|14|13|Moses answered the people, "Do not be afraid. Stand firm and you will see the deliverance the LORD will bring you today. The Egyptians you see today you will never see again.
EXOD|14|14|The LORD will fight for you; you need only to be still."
EXOD|14|15|Then the LORD said to Moses, "Why are you crying out to me? Tell the Israelites to move on.
EXOD|14|16|Raise your staff and stretch out your hand over the sea to divide the water so that the Israelites can go through the sea on dry ground.
EXOD|14|17|I will harden the hearts of the Egyptians so that they will go in after them. And I will gain glory through Pharaoh and all his army, through his chariots and his horsemen.
EXOD|14|18|The Egyptians will know that I am the LORD when I gain glory through Pharaoh, his chariots and his horsemen."
EXOD|14|19|Then the angel of God, who had been traveling in front of Israel's army, withdrew and went behind them. The pillar of cloud also moved from in front and stood behind them,
EXOD|14|20|coming between the armies of Egypt and Israel. Throughout the night the cloud brought darkness to the one side and light to the other side; so neither went near the other all night long.
EXOD|14|21|Then Moses stretched out his hand over the sea, and all that night the LORD drove the sea back with a strong east wind and turned it into dry land. The waters were divided,
EXOD|14|22|and the Israelites went through the sea on dry ground, with a wall of water on their right and on their left.
EXOD|14|23|The Egyptians pursued them, and all Pharaoh's horses and chariots and horsemen followed them into the sea.
EXOD|14|24|During the last watch of the night the LORD looked down from the pillar of fire and cloud at the Egyptian army and threw it into confusion.
EXOD|14|25|He made the wheels of their chariots come off so that they had difficulty driving. And the Egyptians said, "Let's get away from the Israelites! The LORD is fighting for them against Egypt."
EXOD|14|26|Then the LORD said to Moses, "Stretch out your hand over the sea so that the waters may flow back over the Egyptians and their chariots and horsemen."
EXOD|14|27|Moses stretched out his hand over the sea, and at daybreak the sea went back to its place. The Egyptians were fleeing toward it, and the LORD swept them into the sea.
EXOD|14|28|The water flowed back and covered the chariots and horsemen-the entire army of Pharaoh that had followed the Israelites into the sea. Not one of them survived.
EXOD|14|29|But the Israelites went through the sea on dry ground, with a wall of water on their right and on their left.
EXOD|14|30|That day the LORD saved Israel from the hands of the Egyptians, and Israel saw the Egyptians lying dead on the shore.
EXOD|14|31|And when the Israelites saw the great power the LORD displayed against the Egyptians, the people feared the LORD and put their trust in him and in Moses his servant.
EXOD|15|1|Then Moses and the Israelites sang this song to the LORD: "I will sing to the LORD, for he is highly exalted. The horse and its rider he has hurled into the sea.
EXOD|15|2|The LORD is my strength and my song; he has become my salvation. He is my God, and I will praise him, my father's God, and I will exalt him.
EXOD|15|3|The LORD is a warrior; the LORD is his name.
EXOD|15|4|Pharaoh's chariots and his army he has hurled into the sea. The best of Pharaoh's officers are drowned in the Red Sea.
EXOD|15|5|The deep waters have covered them; they sank to the depths like a stone.
EXOD|15|6|"Your right hand, O LORD, was majestic in power. Your right hand, O LORD, shattered the enemy.
EXOD|15|7|In the greatness of your majesty you threw down those who opposed you. You unleashed your burning anger; it consumed them like stubble.
EXOD|15|8|By the blast of your nostrils the waters piled up. The surging waters stood firm like a wall; the deep waters congealed in the heart of the sea.
EXOD|15|9|"The enemy boasted, 'I will pursue, I will overtake them. I will divide the spoils; I will gorge myself on them. I will draw my sword and my hand will destroy them.'
EXOD|15|10|But you blew with your breath, and the sea covered them. They sank like lead in the mighty waters.
EXOD|15|11|"Who among the gods is like you, O LORD? Who is like you- majestic in holiness, awesome in glory, working wonders?
EXOD|15|12|You stretched out your right hand and the earth swallowed them.
EXOD|15|13|"In your unfailing love you will lead the people you have redeemed. In your strength you will guide them to your holy dwelling.
EXOD|15|14|The nations will hear and tremble; anguish will grip the people of Philistia.
EXOD|15|15|The chiefs of Edom will be terrified, the leaders of Moab will be seized with trembling, the people of Canaan will melt away;
EXOD|15|16|terror and dread will fall upon them. By the power of your arm they will be as still as a stone- until your people pass by, O LORD, until the people you bought pass by.
EXOD|15|17|You will bring them in and plant them on the mountain of your inheritance- the place, O LORD, you made for your dwelling, the sanctuary, O Lord, your hands established.
EXOD|15|18|The LORD will reign for ever and ever."
EXOD|15|19|When Pharaoh's horses, chariots and horsemen went into the sea, the LORD brought the waters of the sea back over them, but the Israelites walked through the sea on dry ground.
EXOD|15|20|Then Miriam the prophetess, Aaron's sister, took a tambourine in her hand, and all the women followed her, with tambourines and dancing.
EXOD|15|21|Miriam sang to them: "Sing to the LORD, for he is highly exalted. The horse and its rider he has hurled into the sea."
EXOD|15|22|Then Moses led Israel from the Red Sea and they went into the Desert of Shur. For three days they traveled in the desert without finding water.
EXOD|15|23|When they came to Marah, they could not drink its water because it was bitter. (That is why the place is called Marah. )
EXOD|15|24|So the people grumbled against Moses, saying, "What are we to drink?"
EXOD|15|25|Then Moses cried out to the LORD, and the LORD showed him a piece of wood. He threw it into the water, and the water became sweet. There the LORD made a decree and a law for them, and there he tested them.
EXOD|15|26|He said, "If you listen carefully to the voice of the LORD your God and do what is right in his eyes, if you pay attention to his commands and keep all his decrees, I will not bring on you any of the diseases I brought on the Egyptians, for I am the LORD, who heals you."
EXOD|15|27|Then they came to Elim, where there were twelve springs and seventy palm trees, and they camped there near the water.
EXOD|16|1|The whole Israelite community set out from Elim and came to the Desert of Sin, which is between Elim and Sinai, on the fifteenth day of the second month after they had come out of Egypt.
EXOD|16|2|In the desert the whole community grumbled against Moses and Aaron.
EXOD|16|3|The Israelites said to them, "If only we had died by the LORD's hand in Egypt! There we sat around pots of meat and ate all the food we wanted, but you have brought us out into this desert to starve this entire assembly to death."
EXOD|16|4|Then the LORD said to Moses, "I will rain down bread from heaven for you. The people are to go out each day and gather enough for that day. In this way I will test them and see whether they will follow my instructions.
EXOD|16|5|On the sixth day they are to prepare what they bring in, and that is to be twice as much as they gather on the other days."
EXOD|16|6|So Moses and Aaron said to all the Israelites, "In the evening you will know that it was the LORD who brought you out of Egypt,
EXOD|16|7|and in the morning you will see the glory of the LORD, because he has heard your grumbling against him. Who are we, that you should grumble against us?"
EXOD|16|8|Moses also said, "You will know that it was the LORD when he gives you meat to eat in the evening and all the bread you want in the morning, because he has heard your grumbling against him. Who are we? You are not grumbling against us, but against the LORD."
EXOD|16|9|Then Moses told Aaron, "Say to the entire Israelite community, 'Come before the LORD, for he has heard your grumbling.'"
EXOD|16|10|While Aaron was speaking to the whole Israelite community, they looked toward the desert, and there was the glory of the LORD appearing in the cloud.
EXOD|16|11|The LORD said to Moses,
EXOD|16|12|"I have heard the grumbling of the Israelites. Tell them, 'At twilight you will eat meat, and in the morning you will be filled with bread. Then you will know that I am the LORD your God.'"
EXOD|16|13|That evening quail came and covered the camp, and in the morning there was a layer of dew around the camp.
EXOD|16|14|When the dew was gone, thin flakes like frost on the ground appeared on the desert floor.
EXOD|16|15|When the Israelites saw it, they said to each other, "What is it?" For they did not know what it was. Moses said to them, "It is the bread the LORD has given you to eat.
EXOD|16|16|This is what the LORD has commanded: 'Each one is to gather as much as he needs. Take an omer for each person you have in your tent.'"
EXOD|16|17|The Israelites did as they were told; some gathered much, some little.
EXOD|16|18|And when they measured it by the omer, he who gathered much did not have too much, and he who gathered little did not have too little. Each one gathered as much as he needed.
EXOD|16|19|Then Moses said to them, "No one is to keep any of it until morning."
EXOD|16|20|However, some of them paid no attention to Moses; they kept part of it until morning, but it was full of maggots and began to smell. So Moses was angry with them.
EXOD|16|21|Each morning everyone gathered as much as he needed, and when the sun grew hot, it melted away.
EXOD|16|22|On the sixth day, they gathered twice as much-two omers for each person-and the leaders of the community came and reported this to Moses.
EXOD|16|23|He said to them, "This is what the LORD commanded: 'Tomorrow is to be a day of rest, a holy Sabbath to the LORD. So bake what you want to bake and boil what you want to boil. Save whatever is left and keep it until morning.'"
EXOD|16|24|So they saved it until morning, as Moses commanded, and it did not stink or get maggots in it.
EXOD|16|25|"Eat it today," Moses said, "because today is a Sabbath to the LORD. You will not find any of it on the ground today.
EXOD|16|26|Six days you are to gather it, but on the seventh day, the Sabbath, there will not be any."
EXOD|16|27|Nevertheless, some of the people went out on the seventh day to gather it, but they found none.
EXOD|16|28|Then the LORD said to Moses, "How long will you refuse to keep my commands and my instructions?
EXOD|16|29|Bear in mind that the LORD has given you the Sabbath; that is why on the sixth day he gives you bread for two days. Everyone is to stay where he is on the seventh day; no one is to go out."
EXOD|16|30|So the people rested on the seventh day.
EXOD|16|31|The people of Israel called the bread manna. It was white like coriander seed and tasted like wafers made with honey.
EXOD|16|32|Moses said, "This is what the LORD has commanded: 'Take an omer of manna and keep it for the generations to come, so they can see the bread I gave you to eat in the desert when I brought you out of Egypt.'"
EXOD|16|33|So Moses said to Aaron, "Take a jar and put an omer of manna in it. Then place it before the LORD to be kept for the generations to come."
EXOD|16|34|As the LORD commanded Moses, Aaron put the manna in front of the Testimony, that it might be kept.
EXOD|16|35|The Israelites ate manna forty years, until they came to a land that was settled; they ate manna until they reached the border of Canaan.
EXOD|16|36|(An omer is one tenth of an ephah.)
EXOD|17|1|The whole Israelite community set out from the Desert of Sin, traveling from place to place as the LORD commanded. They camped at Rephidim, but there was no water for the people to drink.
EXOD|17|2|So they quarreled with Moses and said, "Give us water to drink." Moses replied, "Why do you quarrel with me? Why do you put the LORD to the test?"
EXOD|17|3|But the people were thirsty for water there, and they grumbled against Moses. They said, "Why did you bring us up out of Egypt to make us and our children and livestock die of thirst?"
EXOD|17|4|Then Moses cried out to the LORD, "What am I to do with these people? They are almost ready to stone me."
EXOD|17|5|The LORD answered Moses, "Walk on ahead of the people. Take with you some of the elders of Israel and take in your hand the staff with which you struck the Nile, and go.
EXOD|17|6|I will stand there before you by the rock at Horeb. Strike the rock, and water will come out of it for the people to drink." So Moses did this in the sight of the elders of Israel.
EXOD|17|7|And he called the place Massah and Meribah because the Israelites quarreled and because they tested the LORD saying, "Is the LORD among us or not?"
EXOD|17|8|The Amalekites came and attacked the Israelites at Rephidim.
EXOD|17|9|Moses said to Joshua, "Choose some of our men and go out to fight the Amalekites. Tomorrow I will stand on top of the hill with the staff of God in my hands."
EXOD|17|10|So Joshua fought the Amalekites as Moses had ordered, and Moses, Aaron and Hur went to the top of the hill.
EXOD|17|11|As long as Moses held up his hands, the Israelites were winning, but whenever he lowered his hands, the Amalekites were winning.
EXOD|17|12|When Moses' hands grew tired, they took a stone and put it under him and he sat on it. Aaron and Hur held his hands up-one on one side, one on the other-so that his hands remained steady till sunset.
EXOD|17|13|So Joshua overcame the Amalekite army with the sword.
EXOD|17|14|Then the LORD said to Moses, "Write this on a scroll as something to be remembered and make sure that Joshua hears it, because I will completely blot out the memory of Amalek from under heaven."
EXOD|17|15|Moses built an altar and called it The LORD is my Banner.
EXOD|17|16|He said, "For hands were lifted up to the throne of the LORD. The LORD will be at war against the Amalekites from generation to generation."
EXOD|18|1|Now Jethro, the priest of Midian and father-in-law of Moses, heard of everything God had done for Moses and for his people Israel, and how the LORD had brought Israel out of Egypt.
EXOD|18|2|After Moses had sent away his wife Zipporah, his father-in-law Jethro received her
EXOD|18|3|and her two sons. One son was named Gershom, for Moses said, "I have become an alien in a foreign land";
EXOD|18|4|and the other was named Eliezer, for he said, "My father's God was my helper; he saved me from the sword of Pharaoh."
EXOD|18|5|Jethro, Moses' father-in-law, together with Moses' sons and wife, came to him in the desert, where he was camped near the mountain of God.
EXOD|18|6|Jethro had sent word to him, "I, your father-in-law Jethro, am coming to you with your wife and her two sons."
EXOD|18|7|So Moses went out to meet his father-in-law and bowed down and kissed him. They greeted each other and then went into the tent.
EXOD|18|8|Moses told his father-in-law about everything the LORD had done to Pharaoh and the Egyptians for Israel's sake and about all the hardships they had met along the way and how the LORD had saved them.
EXOD|18|9|Jethro was delighted to hear about all the good things the LORD had done for Israel in rescuing them from the hand of the Egyptians.
EXOD|18|10|He said, "Praise be to the LORD, who rescued you from the hand of the Egyptians and of Pharaoh, and who rescued the people from the hand of the Egyptians.
EXOD|18|11|Now I know that the LORD is greater than all other gods, for he did this to those who had treated Israel arrogantly."
EXOD|18|12|Then Jethro, Moses' father-in-law, brought a burnt offering and other sacrifices to God, and Aaron came with all the elders of Israel to eat bread with Moses' father-in-law in the presence of God.
EXOD|18|13|The next day Moses took his seat to serve as judge for the people, and they stood around him from morning till evening.
EXOD|18|14|When his father-in-law saw all that Moses was doing for the people, he said, "What is this you are doing for the people? Why do you alone sit as judge, while all these people stand around you from morning till evening?"
EXOD|18|15|Moses answered him, "Because the people come to me to seek God's will.
EXOD|18|16|Whenever they have a dispute, it is brought to me, and I decide between the parties and inform them of God's decrees and laws."
EXOD|18|17|Moses' father-in-law replied, "What you are doing is not good.
EXOD|18|18|You and these people who come to you will only wear yourselves out. The work is too heavy for you; you cannot handle it alone.
EXOD|18|19|Listen now to me and I will give you some advice, and may God be with you. You must be the people's representative before God and bring their disputes to him.
EXOD|18|20|Teach them the decrees and laws, and show them the way to live and the duties they are to perform.
EXOD|18|21|But select capable men from all the people-men who fear God, trustworthy men who hate dishonest gain-and appoint them as officials over thousands, hundreds, fifties and tens.
EXOD|18|22|Have them serve as judges for the people at all times, but have them bring every difficult case to you; the simple cases they can decide themselves. That will make your load lighter, because they will share it with you.
EXOD|18|23|If you do this and God so commands, you will be able to stand the strain, and all these people will go home satisfied."
EXOD|18|24|Moses listened to his father-in-law and did everything he said.
EXOD|18|25|He chose capable men from all Israel and made them leaders of the people, officials over thousands, hundreds, fifties and tens.
EXOD|18|26|They served as judges for the people at all times. The difficult cases they brought to Moses, but the simple ones they decided themselves.
EXOD|18|27|Then Moses sent his father-in-law on his way, and Jethro returned to his own country.
EXOD|19|1|In the third month after the Israelites left Egypt-on the very day-they came to the Desert of Sinai.
EXOD|19|2|After they set out from Rephidim, they entered the Desert of Sinai, and Israel camped there in the desert in front of the mountain.
EXOD|19|3|Then Moses went up to God, and the LORD called to him from the mountain and said, "This is what you are to say to the house of Jacob and what you are to tell the people of Israel:
EXOD|19|4|'You yourselves have seen what I did to Egypt, and how I carried you on eagles' wings and brought you to myself.
EXOD|19|5|Now if you obey me fully and keep my covenant, then out of all nations you will be my treasured possession. Although the whole earth is mine,
EXOD|19|6|you will be for me a kingdom of priests and a holy nation.' These are the words you are to speak to the Israelites."
EXOD|19|7|So Moses went back and summoned the elders of the people and set before them all the words the LORD had commanded him to speak.
EXOD|19|8|The people all responded together, "We will do everything the LORD has said." So Moses brought their answer back to the LORD.
EXOD|19|9|The LORD said to Moses, "I am going to come to you in a dense cloud, so that the people will hear me speaking with you and will always put their trust in you." Then Moses told the LORD what the people had said.
EXOD|19|10|And the LORD said to Moses, "Go to the people and consecrate them today and tomorrow. Have them wash their clothes
EXOD|19|11|and be ready by the third day, because on that day the LORD will come down on Mount Sinai in the sight of all the people.
EXOD|19|12|Put limits for the people around the mountain and tell them, 'Be careful that you do not go up the mountain or touch the foot of it. Whoever touches the mountain shall surely be put to death.
EXOD|19|13|He shall surely be stoned or shot with arrows; not a hand is to be laid on him. Whether man or animal, he shall not be permitted to live.' Only when the ram's horn sounds a long blast may they go up to the mountain."
EXOD|19|14|After Moses had gone down the mountain to the people, he consecrated them, and they washed their clothes.
EXOD|19|15|Then he said to the people, "Prepare yourselves for the third day. Abstain from sexual relations."
EXOD|19|16|On the morning of the third day there was thunder and lightning, with a thick cloud over the mountain, and a very loud trumpet blast. Everyone in the camp trembled.
EXOD|19|17|Then Moses led the people out of the camp to meet with God, and they stood at the foot of the mountain.
EXOD|19|18|Mount Sinai was covered with smoke, because the LORD descended on it in fire. The smoke billowed up from it like smoke from a furnace, the whole mountain trembled violently,
EXOD|19|19|and the sound of the trumpet grew louder and louder. Then Moses spoke and the voice of God answered him.
EXOD|19|20|The LORD descended to the top of Mount Sinai and called Moses to the top of the mountain. So Moses went up
EXOD|19|21|and the LORD said to him, "Go down and warn the people so they do not force their way through to see the LORD and many of them perish.
EXOD|19|22|Even the priests, who approach the LORD, must consecrate themselves, or the LORD will break out against them."
EXOD|19|23|Moses said to the LORD, "The people cannot come up Mount Sinai, because you yourself warned us, 'Put limits around the mountain and set it apart as holy.'"
EXOD|19|24|The LORD replied, "Go down and bring Aaron up with you. But the priests and the people must not force their way through to come up to the LORD, or he will break out against them."
EXOD|19|25|So Moses went down to the people and told them.
EXOD|20|1|And God spoke all these words:
EXOD|20|2|"I am the LORD your God, who brought you out of Egypt, out of the land of slavery.
EXOD|20|3|"You shall have no other gods before me.
EXOD|20|4|"You shall not make for yourself an idol in the form of anything in heaven above or on the earth beneath or in the waters below.
EXOD|20|5|You shall not bow down to them or worship them; for I, the LORD your God, am a jealous God, punishing the children for the sin of the fathers to the third and fourth generation of those who hate me,
EXOD|20|6|but showing love to a thousand {generations} of those who love me and keep my commandments.
EXOD|20|7|"You shall not misuse the name of the LORD your God, for the LORD will not hold anyone guiltless who misuses his name.
EXOD|20|8|"Remember the Sabbath day by keeping it holy.
EXOD|20|9|Six days you shall labor and do all your work,
EXOD|20|10|but the seventh day is a Sabbath to the LORD your God. On it you shall not do any work, neither you, nor your son or daughter, nor your manservant or maidservant, nor your animals, nor the alien within your gates.
EXOD|20|11|For in six days the LORD made the heavens and the earth, the sea, and all that is in them, but he rested on the seventh day. Therefore the LORD blessed the Sabbath day and made it holy.
EXOD|20|12|"Honor your father and your mother, so that you may live long in the land the LORD your God is giving you.
EXOD|20|13|"You shall not murder.
EXOD|20|14|"You shall not commit adultery.
EXOD|20|15|"You shall not steal.
EXOD|20|16|"You shall not give false testimony against your neighbor.
EXOD|20|17|"You shall not covet your neighbor's house. You shall not covet your neighbor's wife, or his manservant or maidservant, his ox or donkey, or anything that belongs to your neighbor."
EXOD|20|18|When the people saw the thunder and lightning and heard the trumpet and saw the mountain in smoke, they trembled with fear. They stayed at a distance
EXOD|20|19|and said to Moses, "Speak to us yourself and we will listen. But do not have God speak to us or we will die."
EXOD|20|20|Moses said to the people, "Do not be afraid. God has come to test you, so that the fear of God will be with you to keep you from sinning."
EXOD|20|21|The people remained at a distance, while Moses approached the thick darkness where God was.
EXOD|20|22|Then the LORD said to Moses, "Tell the Israelites this: 'You have seen for yourselves that I have spoken to you from heaven:
EXOD|20|23|Do not make any gods to be alongside me; do not make for yourselves gods of silver or gods of gold.
EXOD|20|24|"'Make an altar of earth for me and sacrifice on it your burnt offerings and fellowship offerings, your sheep and goats and your cattle. Wherever I cause my name to be honored, I will come to you and bless you.
EXOD|20|25|If you make an altar of stones for me, do not build it with dressed stones, for you will defile it if you use a tool on it.
EXOD|20|26|And do not go up to my altar on steps, lest your nakedness be exposed on it.'
EXOD|21|1|"These are the laws you are to set before them:
EXOD|21|2|"If you buy a Hebrew servant, he is to serve you for six years. But in the seventh year, he shall go free, without paying anything.
EXOD|21|3|If he comes alone, he is to go free alone; but if he has a wife when he comes, she is to go with him.
EXOD|21|4|If his master gives him a wife and she bears him sons or daughters, the woman and her children shall belong to her master, and only the man shall go free.
EXOD|21|5|"But if the servant declares, 'I love my master and my wife and children and do not want to go free,'
EXOD|21|6|then his master must take him before the judges. He shall take him to the door or the doorpost and pierce his ear with an awl. Then he will be his servant for life.
EXOD|21|7|"If a man sells his daughter as a servant, she is not to go free as menservants do.
EXOD|21|8|If she does not please the master who has selected her for himself, he must let her be redeemed. He has no right to sell her to foreigners, because he has broken faith with her.
EXOD|21|9|If he selects her for his son, he must grant her the rights of a daughter.
EXOD|21|10|If he marries another woman, he must not deprive the first one of her food, clothing and marital rights.
EXOD|21|11|If he does not provide her with these three things, she is to go free, without any payment of money.
EXOD|21|12|"Anyone who strikes a man and kills him shall surely be put to death.
EXOD|21|13|However, if he does not do it intentionally, but God lets it happen, he is to flee to a place I will designate.
EXOD|21|14|But if a man schemes and kills another man deliberately, take him away from my altar and put him to death.
EXOD|21|15|"Anyone who attacks his father or his mother must be put to death.
EXOD|21|16|"Anyone who kidnaps another and either sells him or still has him when he is caught must be put to death.
EXOD|21|17|"Anyone who curses his father or mother must be put to death.
EXOD|21|18|"If men quarrel and one hits the other with a stone or with his fist and he does not die but is confined to bed,
EXOD|21|19|the one who struck the blow will not be held responsible if the other gets up and walks around outside with his staff; however, he must pay the injured man for the loss of his time and see that he is completely healed.
EXOD|21|20|"If a man beats his male or female slave with a rod and the slave dies as a direct result, he must be punished,
EXOD|21|21|but he is not to be punished if the slave gets up after a day or two, since the slave is his property.
EXOD|21|22|"If men who are fighting hit a pregnant woman and she gives birth prematurely but there is no serious injury, the offender must be fined whatever the woman's husband demands and the court allows.
EXOD|21|23|But if there is serious injury, you are to take life for life,
EXOD|21|24|eye for eye, tooth for tooth, hand for hand, foot for foot,
EXOD|21|25|burn for burn, wound for wound, bruise for bruise.
EXOD|21|26|"If a man hits a manservant or maidservant in the eye and destroys it, he must let the servant go free to compensate for the eye.
EXOD|21|27|And if he knocks out the tooth of a manservant or maidservant, he must let the servant go free to compensate for the tooth.
EXOD|21|28|"If a bull gores a man or a woman to death, the bull must be stoned to death, and its meat must not be eaten. But the owner of the bull will not be held responsible.
EXOD|21|29|If, however, the bull has had the habit of goring and the owner has been warned but has not kept it penned up and it kills a man or woman, the bull must be stoned and the owner also must be put to death.
EXOD|21|30|However, if payment is demanded of him, he may redeem his life by paying whatever is demanded.
EXOD|21|31|This law also applies if the bull gores a son or daughter.
EXOD|21|32|If the bull gores a male or female slave, the owner must pay thirty shekels of silver to the master of the slave, and the bull must be stoned.
EXOD|21|33|"If a man uncovers a pit or digs one and fails to cover it and an ox or a donkey falls into it,
EXOD|21|34|the owner of the pit must pay for the loss; he must pay its owner, and the dead animal will be his.
EXOD|21|35|"If a man's bull injures the bull of another and it dies, they are to sell the live one and divide both the money and the dead animal equally.
EXOD|21|36|However, if it was known that the bull had the habit of goring, yet the owner did not keep it penned up, the owner must pay, animal for animal, and the dead animal will be his.
EXOD|22|1|"If a man steals an ox or a sheep and slaughters it or sells it, he must pay back five head of cattle for the ox and four sheep for the sheep.
EXOD|22|2|"If a thief is caught breaking in and is struck so that he dies, the defender is not guilty of bloodshed;
EXOD|22|3|but if it happens after sunrise, he is guilty of bloodshed. "A thief must certainly make restitution, but if he has nothing, he must be sold to pay for his theft.
EXOD|22|4|"If the stolen animal is found alive in his possession-whether ox or donkey or sheep-he must pay back double.
EXOD|22|5|"If a man grazes his livestock in a field or vineyard and lets them stray and they graze in another man's field, he must make restitution from the best of his own field or vineyard.
EXOD|22|6|"If a fire breaks out and spreads into thornbushes so that it burns shocks of grain or standing grain or the whole field, the one who started the fire must make restitution.
EXOD|22|7|"If a man gives his neighbor silver or goods for safekeeping and they are stolen from the neighbor's house, the thief, if he is caught, must pay back double.
EXOD|22|8|But if the thief is not found, the owner of the house must appear before the judges to determine whether he has laid his hands on the other man's property.
EXOD|22|9|In all cases of illegal possession of an ox, a donkey, a sheep, a garment, or any other lost property about which somebody says, 'This is mine,' both parties are to bring their cases before the judges. The one whom the judges declare guilty must pay back double to his neighbor.
EXOD|22|10|"If a man gives a donkey, an ox, a sheep or any other animal to his neighbor for safekeeping and it dies or is injured or is taken away while no one is looking,
EXOD|22|11|the issue between them will be settled by the taking of an oath before the LORD that the neighbor did not lay hands on the other person's property. The owner is to accept this, and no restitution is required.
EXOD|22|12|But if the animal was stolen from the neighbor, he must make restitution to the owner.
EXOD|22|13|If it was torn to pieces by a wild animal, he shall bring in the remains as evidence and he will not be required to pay for the torn animal.
EXOD|22|14|"If a man borrows an animal from his neighbor and it is injured or dies while the owner is not present, he must make restitution.
EXOD|22|15|But if the owner is with the animal, the borrower will not have to pay. If the animal was hired, the money paid for the hire covers the loss.
EXOD|22|16|"If a man seduces a virgin who is not pledged to be married and sleeps with her, he must pay the bride-price, and she shall be his wife.
EXOD|22|17|If her father absolutely refuses to give her to him, he must still pay the bride-price for virgins.
EXOD|22|18|"Do not allow a sorceress to live.
EXOD|22|19|"Anyone who has sexual relations with an animal must be put to death.
EXOD|22|20|"Whoever sacrifices to any god other than the LORD must be destroyed.
EXOD|22|21|"Do not mistreat an alien or oppress him, for you were aliens in Egypt.
EXOD|22|22|"Do not take advantage of a widow or an orphan.
EXOD|22|23|If you do and they cry out to me, I will certainly hear their cry.
EXOD|22|24|My anger will be aroused, and I will kill you with the sword; your wives will become widows and your children fatherless.
EXOD|22|25|"If you lend money to one of my people among you who is needy, do not be like a moneylender; charge him no interest.
EXOD|22|26|If you take your neighbor's cloak as a pledge, return it to him by sunset,
EXOD|22|27|because his cloak is the only covering he has for his body. What else will he sleep in? When he cries out to me, I will hear, for I am compassionate.
EXOD|22|28|"Do not blaspheme God or curse the ruler of your people.
EXOD|22|29|"Do not hold back offerings from your granaries or your vats. "You must give me the firstborn of your sons.
EXOD|22|30|Do the same with your cattle and your sheep. Let them stay with their mothers for seven days, but give them to me on the eighth day.
EXOD|22|31|"You are to be my holy people. So do not eat the meat of an animal torn by wild beasts; throw it to the dogs.
EXOD|23|1|"Do not spread false reports. Do not help a wicked man by being a malicious witness.
EXOD|23|2|"Do not follow the crowd in doing wrong. When you give testimony in a lawsuit, do not pervert justice by siding with the crowd,
EXOD|23|3|and do not show favoritism to a poor man in his lawsuit.
EXOD|23|4|"If you come across your enemy's ox or donkey wandering off, be sure to take it back to him.
EXOD|23|5|If you see the donkey of someone who hates you fallen down under its load, do not leave it there; be sure you help him with it.
EXOD|23|6|"Do not deny justice to your poor people in their lawsuits.
EXOD|23|7|Have nothing to do with a false charge and do not put an innocent or honest person to death, for I will not acquit the guilty.
EXOD|23|8|"Do not accept a bribe, for a bribe blinds those who see and twists the words of the righteous.
EXOD|23|9|"Do not oppress an alien; you yourselves know how it feels to be aliens, because you were aliens in Egypt.
EXOD|23|10|"For six years you are to sow your fields and harvest the crops,
EXOD|23|11|but during the seventh year let the land lie unplowed and unused. Then the poor among your people may get food from it, and the wild animals may eat what they leave. Do the same with your vineyard and your olive grove.
EXOD|23|12|"Six days do your work, but on the seventh day do not work, so that your ox and your donkey may rest and the slave born in your household, and the alien as well, may be refreshed.
EXOD|23|13|"Be careful to do everything I have said to you. Do not invoke the names of other gods; do not let them be heard on your lips.
EXOD|23|14|"Three times a year you are to celebrate a festival to me.
EXOD|23|15|"Celebrate the Feast of Unleavened Bread; for seven days eat bread made without yeast, as I commanded you. Do this at the appointed time in the month of Abib, for in that month you came out of Egypt. "No one is to appear before me empty-handed.
EXOD|23|16|"Celebrate the Feast of Harvest with the firstfruits of the crops you sow in your field. "Celebrate the Feast of Ingathering at the end of the year, when you gather in your crops from the field.
EXOD|23|17|"Three times a year all the men are to appear before the Sovereign LORD.
EXOD|23|18|"Do not offer the blood of a sacrifice to me along with anything containing yeast. "The fat of my festival offerings must not be kept until morning.
EXOD|23|19|"Bring the best of the firstfruits of your soil to the house of the LORD your God. "Do not cook a young goat in its mother's milk.
EXOD|23|20|"See, I am sending an angel ahead of you to guard you along the way and to bring you to the place I have prepared.
EXOD|23|21|Pay attention to him and listen to what he says. Do not rebel against him; he will not forgive your rebellion, since my Name is in him.
EXOD|23|22|If you listen carefully to what he says and do all that I say, I will be an enemy to your enemies and will oppose those who oppose you.
EXOD|23|23|My angel will go ahead of you and bring you into the land of the Amorites, Hittites, Perizzites, Canaanites, Hivites and Jebusites, and I will wipe them out.
EXOD|23|24|Do not bow down before their gods or worship them or follow their practices. You must demolish them and break their sacred stones to pieces.
EXOD|23|25|Worship the LORD your God, and his blessing will be on your food and water. I will take away sickness from among you,
EXOD|23|26|and none will miscarry or be barren in your land. I will give you a full life span.
EXOD|23|27|"I will send my terror ahead of you and throw into confusion every nation you encounter. I will make all your enemies turn their backs and run.
EXOD|23|28|I will send the hornet ahead of you to drive the Hivites, Canaanites and Hittites out of your way.
EXOD|23|29|But I will not drive them out in a single year, because the land would become desolate and the wild animals too numerous for you.
EXOD|23|30|Little by little I will drive them out before you, until you have increased enough to take possession of the land.
EXOD|23|31|"I will establish your borders from the Red Sea to the Sea of the Philistines, and from the desert to the River. I will hand over to you the people who live in the land and you will drive them out before you.
EXOD|23|32|Do not make a covenant with them or with their gods.
EXOD|23|33|Do not let them live in your land, or they will cause you to sin against me, because the worship of their gods will certainly be a snare to you."
EXOD|24|1|Then he said to Moses, "Come up to the LORD, you and Aaron, Nadab and Abihu, and seventy of the elders of Israel. You are to worship at a distance,
EXOD|24|2|but Moses alone is to approach the LORD; the others must not come near. And the people may not come up with him."
EXOD|24|3|When Moses went and told the people all the LORD's words and laws, they responded with one voice, "Everything the LORD has said we will do."
EXOD|24|4|Moses then wrote down everything the LORD had said. He got up early the next morning and built an altar at the foot of the mountain and set up twelve stone pillars representing the twelve tribes of Israel.
EXOD|24|5|Then he sent young Israelite men, and they offered burnt offerings and sacrificed young bulls as fellowship offerings to the LORD.
EXOD|24|6|Moses took half of the blood and put it in bowls, and the other half he sprinkled on the altar.
EXOD|24|7|Then he took the Book of the Covenant and read it to the people. They responded, "We will do everything the LORD has said; we will obey."
EXOD|24|8|Moses then took the blood, sprinkled it on the people and said, "This is the blood of the covenant that the LORD has made with you in accordance with all these words."
EXOD|24|9|Moses and Aaron, Nadab and Abihu, and the seventy elders of Israel went up
EXOD|24|10|and saw the God of Israel. Under his feet was something like a pavement made of sapphire, clear as the sky itself.
EXOD|24|11|But God did not raise his hand against these leaders of the Israelites; they saw God, and they ate and drank.
EXOD|24|12|The LORD said to Moses, "Come up to me on the mountain and stay here, and I will give you the tablets of stone, with the law and commands I have written for their instruction."
EXOD|24|13|Then Moses set out with Joshua his aide, and Moses went up on the mountain of God.
EXOD|24|14|He said to the elders, "Wait here for us until we come back to you. Aaron and Hur are with you, and anyone involved in a dispute can go to them."
EXOD|24|15|When Moses went up on the mountain, the cloud covered it,
EXOD|24|16|and the glory of the LORD settled on Mount Sinai. For six days the cloud covered the mountain, and on the seventh day the LORD called to Moses from within the cloud.
EXOD|24|17|To the Israelites the glory of the LORD looked like a consuming fire on top of the mountain.
EXOD|24|18|Then Moses entered the cloud as he went on up the mountain. And he stayed on the mountain forty days and forty nights.
EXOD|25|1|The LORD said to Moses,
EXOD|25|2|"Tell the Israelites to bring me an offering. You are to receive the offering for me from each man whose heart prompts him to give.
EXOD|25|3|These are the offerings you are to receive from them: gold, silver and bronze;
EXOD|25|4|blue, purple and scarlet yarn and fine linen; goat hair;
EXOD|25|5|ram skins dyed red and hides of sea cows; acacia wood;
EXOD|25|6|olive oil for the light; spices for the anointing oil and for the fragrant incense;
EXOD|25|7|and onyx stones and other gems to be mounted on the ephod and breastpiece.
EXOD|25|8|"Then have them make a sanctuary for me, and I will dwell among them.
EXOD|25|9|Make this tabernacle and all its furnishings exactly like the pattern I will show you.
EXOD|25|10|"Have them make a chest of acacia wood-two and a half cubits long, a cubit and a half wide, and a cubit and a half high.
EXOD|25|11|Overlay it with pure gold, both inside and out, and make a gold molding around it.
EXOD|25|12|Cast four gold rings for it and fasten them to its four feet, with two rings on one side and two rings on the other.
EXOD|25|13|Then make poles of acacia wood and overlay them with gold.
EXOD|25|14|Insert the poles into the rings on the sides of the chest to carry it.
EXOD|25|15|The poles are to remain in the rings of this ark; they are not to be removed.
EXOD|25|16|Then put in the ark the Testimony, which I will give you.
EXOD|25|17|"Make an atonement cover of pure gold-two and a half cubits long and a cubit and a half wide.
EXOD|25|18|And make two cherubim out of hammered gold at the ends of the cover.
EXOD|25|19|Make one cherub on one end and the second cherub on the other; make the cherubim of one piece with the cover, at the two ends.
EXOD|25|20|The cherubim are to have their wings spread upward, overshadowing the cover with them. The cherubim are to face each other, looking toward the cover.
EXOD|25|21|Place the cover on top of the ark and put in the ark the Testimony, which I will give you.
EXOD|25|22|There, above the cover between the two cherubim that are over the ark of the Testimony, I will meet with you and give you all my commands for the Israelites.
EXOD|25|23|"Make a table of acacia wood-two cubits long, a cubit wide and a cubit and a half high.
EXOD|25|24|Overlay it with pure gold and make a gold molding around it.
EXOD|25|25|Also make around it a rim a handbreadth wide and put a gold molding on the rim.
EXOD|25|26|Make four gold rings for the table and fasten them to the four corners, where the four legs are.
EXOD|25|27|The rings are to be close to the rim to hold the poles used in carrying the table.
EXOD|25|28|Make the poles of acacia wood, overlay them with gold and carry the table with them.
EXOD|25|29|And make its plates and dishes of pure gold, as well as its pitchers and bowls for the pouring out of offerings.
EXOD|25|30|Put the bread of the Presence on this table to be before me at all times.
EXOD|25|31|"Make a lampstand of pure gold and hammer it out, base and shaft; its flowerlike cups, buds and blossoms shall be of one piece with it.
EXOD|25|32|Six branches are to extend from the sides of the lampstand-three on one side and three on the other.
EXOD|25|33|Three cups shaped like almond flowers with buds and blossoms are to be on one branch, three on the next branch, and the same for all six branches extending from the lampstand.
EXOD|25|34|And on the lampstand there are to be four cups shaped like almond flowers with buds and blossoms.
EXOD|25|35|One bud shall be under the first pair of branches extending from the lampstand, a second bud under the second pair, and a third bud under the third pair-six branches in all.
EXOD|25|36|The buds and branches shall all be of one piece with the lampstand, hammered out of pure gold.
EXOD|25|37|"Then make its seven lamps and set them up on it so that they light the space in front of it.
EXOD|25|38|Its wick trimmers and trays are to be of pure gold.
EXOD|25|39|A talent of pure gold is to be used for the lampstand and all these accessories.
EXOD|25|40|See that you make them according to the pattern shown you on the mountain.
EXOD|26|1|"Make the tabernacle with ten curtains of finely twisted linen and blue, purple and scarlet yarn, with cherubim worked into them by a skilled craftsman.
EXOD|26|2|All the curtains are to be the same size-twenty-eight cubits long and four cubits wide.
EXOD|26|3|Join five of the curtains together, and do the same with the other five.
EXOD|26|4|Make loops of blue material along the edge of the end curtain in one set, and do the same with the end curtain in the other set.
EXOD|26|5|Make fifty loops on one curtain and fifty loops on the end curtain of the other set, with the loops opposite each other.
EXOD|26|6|Then make fifty gold clasps and use them to fasten the curtains together so that the tabernacle is a unit.
EXOD|26|7|"Make curtains of goat hair for the tent over the tabernacle-eleven altogether.
EXOD|26|8|All eleven curtains are to be the same size-thirty cubits long and four cubits wide.
EXOD|26|9|Join five of the curtains together into one set and the other six into another set. Fold the sixth curtain double at the front of the tent.
EXOD|26|10|Make fifty loops along the edge of the end curtain in one set and also along the edge of the end curtain in the other set.
EXOD|26|11|Then make fifty bronze clasps and put them in the loops to fasten the tent together as a unit.
EXOD|26|12|As for the additional length of the tent curtains, the half curtain that is left over is to hang down at the rear of the tabernacle.
EXOD|26|13|The tent curtains will be a cubit longer on both sides; what is left will hang over the sides of the tabernacle so as to cover it.
EXOD|26|14|Make for the tent a covering of ram skins dyed red, and over that a covering of hides of sea cows.
EXOD|26|15|"Make upright frames of acacia wood for the tabernacle.
EXOD|26|16|Each frame is to be ten cubits long and a cubit and a half wide,
EXOD|26|17|with two projections set parallel to each other. Make all the frames of the tabernacle in this way.
EXOD|26|18|Make twenty frames for the south side of the tabernacle
EXOD|26|19|and make forty silver bases to go under them-two bases for each frame, one under each projection.
EXOD|26|20|For the other side, the north side of the tabernacle, make twenty frames
EXOD|26|21|and forty silver bases-two under each frame.
EXOD|26|22|Make six frames for the far end, that is, the west end of the tabernacle,
EXOD|26|23|and make two frames for the corners at the far end.
EXOD|26|24|At these two corners they must be double from the bottom all the way to the top, and fitted into a single ring; both shall be like that.
EXOD|26|25|So there will be eight frames and sixteen silver bases-two under each frame.
EXOD|26|26|"Also make crossbars of acacia wood: five for the frames on one side of the tabernacle,
EXOD|26|27|five for those on the other side, and five for the frames on the west, at the far end of the tabernacle.
EXOD|26|28|The center crossbar is to extend from end to end at the middle of the frames.
EXOD|26|29|Overlay the frames with gold and make gold rings to hold the crossbars. Also overlay the crossbars with gold.
EXOD|26|30|"Set up the tabernacle according to the plan shown you on the mountain.
EXOD|26|31|"Make a curtain of blue, purple and scarlet yarn and finely twisted linen, with cherubim worked into it by a skilled craftsman.
EXOD|26|32|Hang it with gold hooks on four posts of acacia wood overlaid with gold and standing on four silver bases.
EXOD|26|33|Hang the curtain from the clasps and place the ark of the Testimony behind the curtain. The curtain will separate the Holy Place from the Most Holy Place.
EXOD|26|34|Put the atonement cover on the ark of the Testimony in the Most Holy Place.
EXOD|26|35|Place the table outside the curtain on the north side of the tabernacle and put the lampstand opposite it on the south side.
EXOD|26|36|"For the entrance to the tent make a curtain of blue, purple and scarlet yarn and finely twisted linen-the work of an embroiderer.
EXOD|26|37|Make gold hooks for this curtain and five posts of acacia wood overlaid with gold. And cast five bronze bases for them.
EXOD|27|1|"Build an altar of acacia wood, three cubits high; it is to be square, five cubits long and five cubits wide.
EXOD|27|2|Make a horn at each of the four corners, so that the horns and the altar are of one piece, and overlay the altar with bronze.
EXOD|27|3|Make all its utensils of bronze-its pots to remove the ashes, and its shovels, sprinkling bowls, meat forks and firepans.
EXOD|27|4|Make a grating for it, a bronze network, and make a bronze ring at each of the four corners of the network.
EXOD|27|5|Put it under the ledge of the altar so that it is halfway up the altar.
EXOD|27|6|Make poles of acacia wood for the altar and overlay them with bronze.
EXOD|27|7|The poles are to be inserted into the rings so they will be on two sides of the altar when it is carried.
EXOD|27|8|Make the altar hollow, out of boards. It is to be made just as you were shown on the mountain.
EXOD|27|9|"Make a courtyard for the tabernacle. The south side shall be a hundred cubits long and is to have curtains of finely twisted linen,
EXOD|27|10|with twenty posts and twenty bronze bases and with silver hooks and bands on the posts.
EXOD|27|11|The north side shall also be a hundred cubits long and is to have curtains, with twenty posts and twenty bronze bases and with silver hooks and bands on the posts.
EXOD|27|12|"The west end of the courtyard shall be fifty cubits wide and have curtains, with ten posts and ten bases.
EXOD|27|13|On the east end, toward the sunrise, the courtyard shall also be fifty cubits wide.
EXOD|27|14|Curtains fifteen cubits long are to be on one side of the entrance, with three posts and three bases,
EXOD|27|15|and curtains fifteen cubits long are to be on the other side, with three posts and three bases.
EXOD|27|16|"For the entrance to the courtyard, provide a curtain twenty cubits long, of blue, purple and scarlet yarn and finely twisted linen-the work of an embroiderer-with four posts and four bases.
EXOD|27|17|All the posts around the courtyard are to have silver bands and hooks, and bronze bases.
EXOD|27|18|The courtyard shall be a hundred cubits long and fifty cubits wide, with curtains of finely twisted linen five cubits high, and with bronze bases.
EXOD|27|19|All the other articles used in the service of the tabernacle, whatever their function, including all the tent pegs for it and those for the courtyard, are to be of bronze.
EXOD|27|20|"Command the Israelites to bring you clear oil of pressed olives for the light so that the lamps may be kept burning.
EXOD|27|21|In the Tent of Meeting, outside the curtain that is in front of the Testimony, Aaron and his sons are to keep the lamps burning before the LORD from evening till morning. This is to be a lasting ordinance among the Israelites for the generations to come.
EXOD|28|1|"Have Aaron your brother brought to you from among the Israelites, along with his sons Nadab and Abihu, Eleazar and Ithamar, so they may serve me as priests.
EXOD|28|2|Make sacred garments for your brother Aaron, to give him dignity and honor.
EXOD|28|3|Tell all the skilled men to whom I have given wisdom in such matters that they are to make garments for Aaron, for his consecration, so he may serve me as priest.
EXOD|28|4|These are the garments they are to make: a breastpiece, an ephod, a robe, a woven tunic, a turban and a sash. They are to make these sacred garments for your brother Aaron and his sons, so they may serve me as priests.
EXOD|28|5|Have them use gold, and blue, purple and scarlet yarn, and fine linen.
EXOD|28|6|"Make the ephod of gold, and of blue, purple and scarlet yarn, and of finely twisted linen-the work of a skilled craftsman.
EXOD|28|7|It is to have two shoulder pieces attached to two of its corners, so it can be fastened.
EXOD|28|8|Its skillfully woven waistband is to be like it-of one piece with the ephod and made with gold, and with blue, purple and scarlet yarn, and with finely twisted linen.
EXOD|28|9|"Take two onyx stones and engrave on them the names of the sons of Israel
EXOD|28|10|in the order of their birth-six names on one stone and the remaining six on the other.
EXOD|28|11|Engrave the names of the sons of Israel on the two stones the way a gem cutter engraves a seal. Then mount the stones in gold filigree settings
EXOD|28|12|and fasten them on the shoulder pieces of the ephod as memorial stones for the sons of Israel. Aaron is to bear the names on his shoulders as a memorial before the LORD.
EXOD|28|13|Make gold filigree settings
EXOD|28|14|and two braided chains of pure gold, like a rope, and attach the chains to the settings.
EXOD|28|15|"Fashion a breastpiece for making decisions-the work of a skilled craftsman. Make it like the ephod: of gold, and of blue, purple and scarlet yarn, and of finely twisted linen.
EXOD|28|16|It is to be square-a span long and a span wide-and folded double.
EXOD|28|17|Then mount four rows of precious stones on it. In the first row there shall be a ruby, a topaz and a beryl;
EXOD|28|18|in the second row a turquoise, a sapphire and an emerald;
EXOD|28|19|in the third row a jacinth, an agate and an amethyst;
EXOD|28|20|in the fourth row a chrysolite, an onyx and a jasper. Mount them in gold filigree settings.
EXOD|28|21|There are to be twelve stones, one for each of the names of the sons of Israel, each engraved like a seal with the name of one of the twelve tribes.
EXOD|28|22|"For the breastpiece make braided chains of pure gold, like a rope.
EXOD|28|23|Make two gold rings for it and fasten them to two corners of the breastpiece.
EXOD|28|24|Fasten the two gold chains to the rings at the corners of the breastpiece,
EXOD|28|25|and the other ends of the chains to the two settings, attaching them to the shoulder pieces of the ephod at the front.
EXOD|28|26|Make two gold rings and attach them to the other two corners of the breastpiece on the inside edge next to the ephod.
EXOD|28|27|Make two more gold rings and attach them to the bottom of the shoulder pieces on the front of the ephod, close to the seam just above the waistband of the ephod.
EXOD|28|28|The rings of the breastpiece are to be tied to the rings of the ephod with blue cord, connecting it to the waistband, so that the breastpiece will not swing out from the ephod.
EXOD|28|29|"Whenever Aaron enters the Holy Place, he will bear the names of the sons of Israel over his heart on the breastpiece of decision as a continuing memorial before the LORD.
EXOD|28|30|Also put the Urim and the Thummim in the breastpiece, so they may be over Aaron's heart whenever he enters the presence of the LORD. Thus Aaron will always bear the means of making decisions for the Israelites over his heart before the LORD.
EXOD|28|31|"Make the robe of the ephod entirely of blue cloth,
EXOD|28|32|with an opening for the head in its center. There shall be a woven edge like a collar around this opening, so that it will not tear.
EXOD|28|33|Make pomegranates of blue, purple and scarlet yarn around the hem of the robe, with gold bells between them.
EXOD|28|34|The gold bells and the pomegranates are to alternate around the hem of the robe.
EXOD|28|35|Aaron must wear it when he ministers. The sound of the bells will be heard when he enters the Holy Place before the LORD and when he comes out, so that he will not die.
EXOD|28|36|"Make a plate of pure gold and engrave on it as on a seal:HOLY TO THE LORD.
EXOD|28|37|Fasten a blue cord to it to attach it to the turban; it is to be on the front of the turban.
EXOD|28|38|It will be on Aaron's forehead, and he will bear the guilt involved in the sacred gifts the Israelites consecrate, whatever their gifts may be. It will be on Aaron's forehead continually so that they will be acceptable to the LORD.
EXOD|28|39|"Weave the tunic of fine linen and make the turban of fine linen. The sash is to be the work of an embroiderer.
EXOD|28|40|Make tunics, sashes and headbands for Aaron's sons, to give them dignity and honor.
EXOD|28|41|After you put these clothes on your brother Aaron and his sons, anoint and ordain them. Consecrate them so they may serve me as priests.
EXOD|28|42|"Make linen undergarments as a covering for the body, reaching from the waist to the thigh.
EXOD|28|43|Aaron and his sons must wear them whenever they enter the Tent of Meeting or approach the altar to minister in the Holy Place, so that they will not incur guilt and die. "This is to be a lasting ordinance for Aaron and his descendants.
EXOD|29|1|"This is what you are to do to consecrate them, so they may serve me as priests: Take a young bull and two rams without defect.
EXOD|29|2|And from fine wheat flour, without yeast, make bread, and cakes mixed with oil, and wafers spread with oil.
EXOD|29|3|Put them in a basket and present them in it-along with the bull and the two rams.
EXOD|29|4|Then bring Aaron and his sons to the entrance to the Tent of Meeting and wash them with water.
EXOD|29|5|Take the garments and dress Aaron with the tunic, the robe of the ephod, the ephod itself and the breastpiece. Fasten the ephod on him by its skillfully woven waistband.
EXOD|29|6|Put the turban on his head and attach the sacred diadem to the turban.
EXOD|29|7|Take the anointing oil and anoint him by pouring it on his head.
EXOD|29|8|Bring his sons and dress them in tunics
EXOD|29|9|and put headbands on them. Then tie sashes on Aaron and his sons. The priesthood is theirs by a lasting ordinance. In this way you shall ordain Aaron and his sons.
EXOD|29|10|"Bring the bull to the front of the Tent of Meeting, and Aaron and his sons shall lay their hands on its head.
EXOD|29|11|Slaughter it in the LORD's presence at the entrance to the Tent of Meeting.
EXOD|29|12|Take some of the bull's blood and put it on the horns of the altar with your finger, and pour out the rest of it at the base of the altar.
EXOD|29|13|Then take all the fat around the inner parts, the covering of the liver, and both kidneys with the fat on them, and burn them on the altar.
EXOD|29|14|But burn the bull's flesh and its hide and its offal outside the camp. It is a sin offering.
EXOD|29|15|"Take one of the rams, and Aaron and his sons shall lay their hands on its head.
EXOD|29|16|Slaughter it and take the blood and sprinkle it against the altar on all sides.
EXOD|29|17|Cut the ram into pieces and wash the inner parts and the legs, putting them with the head and the other pieces.
EXOD|29|18|Then burn the entire ram on the altar. It is a burnt offering to the LORD, a pleasing aroma, an offering made to the LORD by fire.
EXOD|29|19|"Take the other ram, and Aaron and his sons shall lay their hands on its head.
EXOD|29|20|Slaughter it, take some of its blood and put it on the lobes of the right ears of Aaron and his sons, on the thumbs of their right hands, and on the big toes of their right feet. Then sprinkle blood against the altar on all sides.
EXOD|29|21|And take some of the blood on the altar and some of the anointing oil and sprinkle it on Aaron and his garments and on his sons and their garments. Then he and his sons and their garments will be consecrated.
EXOD|29|22|"Take from this ram the fat, the fat tail, the fat around the inner parts, the covering of the liver, both kidneys with the fat on them, and the right thigh. (This is the ram for the ordination.)
EXOD|29|23|From the basket of bread made without yeast, which is before the LORD, take a loaf, and a cake made with oil, and a wafer.
EXOD|29|24|Put all these in the hands of Aaron and his sons and wave them before the LORD as a wave offering.
EXOD|29|25|Then take them from their hands and burn them on the altar along with the burnt offering for a pleasing aroma to the LORD, an offering made to the LORD by fire.
EXOD|29|26|After you take the breast of the ram for Aaron's ordination, wave it before the LORD as a wave offering, and it will be your share.
EXOD|29|27|"Consecrate those parts of the ordination ram that belong to Aaron and his sons: the breast that was waved and the thigh that was presented.
EXOD|29|28|This is always to be the regular share from the Israelites for Aaron and his sons. It is the contribution the Israelites are to make to the LORD from their fellowship offerings.
EXOD|29|29|"Aaron's sacred garments will belong to his descendants so that they can be anointed and ordained in them.
EXOD|29|30|The son who succeeds him as priest and comes to the Tent of Meeting to minister in the Holy Place is to wear them seven days.
EXOD|29|31|"Take the ram for the ordination and cook the meat in a sacred place.
EXOD|29|32|At the entrance to the Tent of Meeting, Aaron and his sons are to eat the meat of the ram and the bread that is in the basket.
EXOD|29|33|They are to eat these offerings by which atonement was made for their ordination and consecration. But no one else may eat them, because they are sacred.
EXOD|29|34|And if any of the meat of the ordination ram or any bread is left over till morning, burn it up. It must not be eaten, because it is sacred.
EXOD|29|35|"Do for Aaron and his sons everything I have commanded you, taking seven days to ordain them.
EXOD|29|36|Sacrifice a bull each day as a sin offering to make atonement. Purify the altar by making atonement for it, and anoint it to consecrate it.
EXOD|29|37|For seven days make atonement for the altar and consecrate it. Then the altar will be most holy, and whatever touches it will be holy.
EXOD|29|38|"This is what you are to offer on the altar regularly each day: two lambs a year old.
EXOD|29|39|Offer one in the morning and the other at twilight.
EXOD|29|40|With the first lamb offer a tenth of an ephah of fine flour mixed with a quarter of a hin of oil from pressed olives, and a quarter of a hin of wine as a drink offering.
EXOD|29|41|Sacrifice the other lamb at twilight with the same grain offering and its drink offering as in the morning-a pleasing aroma, an offering made to the LORD by fire.
EXOD|29|42|"For the generations to come this burnt offering is to be made regularly at the entrance to the Tent of Meeting before the LORD. There I will meet you and speak to you;
EXOD|29|43|there also I will meet with the Israelites, and the place will be consecrated by my glory.
EXOD|29|44|"So I will consecrate the Tent of Meeting and the altar and will consecrate Aaron and his sons to serve me as priests.
EXOD|29|45|Then I will dwell among the Israelites and be their God.
EXOD|29|46|They will know that I am the LORD their God, who brought them out of Egypt so that I might dwell among them. I am the LORD their God.
EXOD|30|1|"Make an altar of acacia wood for burning incense.
EXOD|30|2|It is to be square, a cubit long and a cubit wide, and two cubits high -its horns of one piece with it.
EXOD|30|3|Overlay the top and all the sides and the horns with pure gold, and make a gold molding around it.
EXOD|30|4|Make two gold rings for the altar below the molding-two on opposite sides-to hold the poles used to carry it.
EXOD|30|5|Make the poles of acacia wood and overlay them with gold.
EXOD|30|6|Put the altar in front of the curtain that is before the ark of the Testimony-before the atonement cover that is over the Testimony-where I will meet with you.
EXOD|30|7|"Aaron must burn fragrant incense on the altar every morning when he tends the lamps.
EXOD|30|8|He must burn incense again when he lights the lamps at twilight so incense will burn regularly before the LORD for the generations to come.
EXOD|30|9|Do not offer on this altar any other incense or any burnt offering or grain offering, and do not pour a drink offering on it.
EXOD|30|10|Once a year Aaron shall make atonement on its horns. This annual atonement must be made with the blood of the atoning sin offering for the generations to come. It is most holy to the LORD."
EXOD|30|11|Then the LORD said to Moses,
EXOD|30|12|"When you take a census of the Israelites to count them, each one must pay the LORD a ransom for his life at the time he is counted. Then no plague will come on them when you number them.
EXOD|30|13|Each one who crosses over to those already counted is to give a half shekel, according to the sanctuary shekel, which weighs twenty gerahs. This half shekel is an offering to the LORD.
EXOD|30|14|All who cross over, those twenty years old or more, are to give an offering to the LORD.
EXOD|30|15|The rich are not to give more than a half shekel and the poor are not to give less when you make the offering to the LORD to atone for your lives.
EXOD|30|16|Receive the atonement money from the Israelites and use it for the service of the Tent of Meeting. It will be a memorial for the Israelites before the LORD, making atonement for your lives."
EXOD|30|17|Then the LORD said to Moses,
EXOD|30|18|"Make a bronze basin, with its bronze stand, for washing. Place it between the Tent of Meeting and the altar, and put water in it.
EXOD|30|19|Aaron and his sons are to wash their hands and feet with water from it.
EXOD|30|20|Whenever they enter the Tent of Meeting, they shall wash with water so that they will not die. Also, when they approach the altar to minister by presenting an offering made to the LORD by fire,
EXOD|30|21|they shall wash their hands and feet so that they will not die. This is to be a lasting ordinance for Aaron and his descendants for the generations to come."
EXOD|30|22|Then the LORD said to Moses,
EXOD|30|23|"Take the following fine spices: 500 shekels of liquid myrrh, half as much (that is, 250 shekels) of fragrant cinnamon, 250 shekels of fragrant cane,
EXOD|30|24|500 shekels of cassia-all according to the sanctuary shekel-and a hin of olive oil.
EXOD|30|25|Make these into a sacred anointing oil, a fragrant blend, the work of a perfumer. It will be the sacred anointing oil.
EXOD|30|26|Then use it to anoint the Tent of Meeting, the ark of the Testimony,
EXOD|30|27|the table and all its articles, the lampstand and its accessories, the altar of incense,
EXOD|30|28|the altar of burnt offering and all its utensils, and the basin with its stand.
EXOD|30|29|You shall consecrate them so they will be most holy, and whatever touches them will be holy.
EXOD|30|30|"Anoint Aaron and his sons and consecrate them so they may serve me as priests.
EXOD|30|31|Say to the Israelites, 'This is to be my sacred anointing oil for the generations to come.
EXOD|30|32|Do not pour it on men's bodies and do not make any oil with the same formula. It is sacred, and you are to consider it sacred.
EXOD|30|33|Whoever makes perfume like it and whoever puts it on anyone other than a priest must be cut off from his people.'"
EXOD|30|34|Then the LORD said to Moses, "Take fragrant spices-gum resin, onycha and galbanum-and pure frankincense, all in equal amounts,
EXOD|30|35|and make a fragrant blend of incense, the work of a perfumer. It is to be salted and pure and sacred.
EXOD|30|36|Grind some of it to powder and place it in front of the Testimony in the Tent of Meeting, where I will meet with you. It shall be most holy to you.
EXOD|30|37|Do not make any incense with this formula for yourselves; consider it holy to the LORD.
EXOD|30|38|Whoever makes any like it to enjoy its fragrance must be cut off from his people."
EXOD|31|1|Then the LORD said to Moses,
EXOD|31|2|"See, I have chosen Bezalel son of Uri, the son of Hur, of the tribe of Judah,
EXOD|31|3|and I have filled him with the Spirit of God, with skill, ability and knowledge in all kinds of crafts-
EXOD|31|4|to make artistic designs for work in gold, silver and bronze,
EXOD|31|5|to cut and set stones, to work in wood, and to engage in all kinds of craftsmanship.
EXOD|31|6|Moreover, I have appointed Oholiab son of Ahisamach, of the tribe of Dan, to help him. Also I have given skill to all the craftsmen to make everything I have commanded you:
EXOD|31|7|the Tent of Meeting, the ark of the Testimony with the atonement cover on it, and all the other furnishings of the tent-
EXOD|31|8|the table and its articles, the pure gold lampstand and all its accessories, the altar of incense,
EXOD|31|9|the altar of burnt offering and all its utensils, the basin with its stand-
EXOD|31|10|and also the woven garments, both the sacred garments for Aaron the priest and the garments for his sons when they serve as priests,
EXOD|31|11|and the anointing oil and fragrant incense for the Holy Place. They are to make them just as I commanded you."
EXOD|31|12|Then the LORD said to Moses,
EXOD|31|13|"Say to the Israelites, 'You must observe my Sabbaths. This will be a sign between me and you for the generations to come, so you may know that I am the LORD, who makes you holy.
EXOD|31|14|"'Observe the Sabbath, because it is holy to you. Anyone who desecrates it must be put to death; whoever does any work on that day must be cut off from his people.
EXOD|31|15|For six days, work is to be done, but the seventh day is a Sabbath of rest, holy to the LORD. Whoever does any work on the Sabbath day must be put to death.
EXOD|31|16|The Israelites are to observe the Sabbath, celebrating it for the generations to come as a lasting covenant.
EXOD|31|17|It will be a sign between me and the Israelites forever, for in six days the LORD made the heavens and the earth, and on the seventh day he abstained from work and rested.'"
EXOD|31|18|When the LORD finished speaking to Moses on Mount Sinai, he gave him the two tablets of the Testimony, the tablets of stone inscribed by the finger of God.
EXOD|32|1|When the people saw that Moses was so long in coming down from the mountain, they gathered around Aaron and said, "Come, make us gods who will go before us. As for this fellow Moses who brought us up out of Egypt, we don't know what has happened to him."
EXOD|32|2|Aaron answered them, "Take off the gold earrings that your wives, your sons and your daughters are wearing, and bring them to me."
EXOD|32|3|So all the people took off their earrings and brought them to Aaron.
EXOD|32|4|He took what they handed him and made it into an idol cast in the shape of a calf, fashioning it with a tool. Then they said, "These are your gods, O Israel, who brought you up out of Egypt."
EXOD|32|5|When Aaron saw this, he built an altar in front of the calf and announced, "Tomorrow there will be a festival to the LORD."
EXOD|32|6|So the next day the people rose early and sacrificed burnt offerings and presented fellowship offerings. Afterward they sat down to eat and drink and got up to indulge in revelry.
EXOD|32|7|Then the LORD said to Moses, "Go down, because your people, whom you brought up out of Egypt, have become corrupt.
EXOD|32|8|They have been quick to turn away from what I commanded them and have made themselves an idol cast in the shape of a calf. They have bowed down to it and sacrificed to it and have said, 'These are your gods, O Israel, who brought you up out of Egypt.'
EXOD|32|9|"I have seen these people," the LORD said to Moses, "and they are a stiff-necked people.
EXOD|32|10|Now leave me alone so that my anger may burn against them and that I may destroy them. Then I will make you into a great nation."
EXOD|32|11|But Moses sought the favor of the LORD his God. "O LORD," he said, "why should your anger burn against your people, whom you brought out of Egypt with great power and a mighty hand?
EXOD|32|12|Why should the Egyptians say, 'It was with evil intent that he brought them out, to kill them in the mountains and to wipe them off the face of the earth'? Turn from your fierce anger; relent and do not bring disaster on your people.
EXOD|32|13|Remember your servants Abraham, Isaac and Israel, to whom you swore by your own self: 'I will make your descendants as numerous as the stars in the sky and I will give your descendants all this land I promised them, and it will be their inheritance forever.'"
EXOD|32|14|Then the LORD relented and did not bring on his people the disaster he had threatened.
EXOD|32|15|Moses turned and went down the mountain with the two tablets of the Testimony in his hands. They were inscribed on both sides, front and back.
EXOD|32|16|The tablets were the work of God; the writing was the writing of God, engraved on the tablets.
EXOD|32|17|When Joshua heard the noise of the people shouting, he said to Moses, "There is the sound of war in the camp."
EXOD|32|18|Moses replied: "It is not the sound of victory, it is not the sound of defeat; it is the sound of singing that I hear."
EXOD|32|19|When Moses approached the camp and saw the calf and the dancing, his anger burned and he threw the tablets out of his hands, breaking them to pieces at the foot of the mountain.
EXOD|32|20|And he took the calf they had made and burned it in the fire; then he ground it to powder, scattered it on the water and made the Israelites drink it.
EXOD|32|21|He said to Aaron, "What did these people do to you, that you led them into such great sin?"
EXOD|32|22|"Do not be angry, my lord," Aaron answered. "You know how prone these people are to evil.
EXOD|32|23|They said to me, 'Make us gods who will go before us. As for this fellow Moses who brought us up out of Egypt, we don't know what has happened to him.'
EXOD|32|24|So I told them, 'Whoever has any gold jewelry, take it off.' Then they gave me the gold, and I threw it into the fire, and out came this calf!"
EXOD|32|25|Moses saw that the people were running wild and that Aaron had let them get out of control and so become a laughingstock to their enemies.
EXOD|32|26|So he stood at the entrance to the camp and said, "Whoever is for the LORD, come to me." And all the Levites rallied to him.
EXOD|32|27|Then he said to them, "This is what the LORD, the God of Israel, says: 'Each man strap a sword to his side. Go back and forth through the camp from one end to the other, each killing his brother and friend and neighbor.'"
EXOD|32|28|The Levites did as Moses commanded, and that day about three thousand of the people died.
EXOD|32|29|Then Moses said, "You have been set apart to the LORD today, for you were against your own sons and brothers, and he has blessed you this day."
EXOD|32|30|The next day Moses said to the people, "You have committed a great sin. But now I will go up to the LORD; perhaps I can make atonement for your sin."
EXOD|32|31|So Moses went back to the LORD and said, "Oh, what a great sin these people have committed! They have made themselves gods of gold.
EXOD|32|32|But now, please forgive their sin-but if not, then blot me out of the book you have written."
EXOD|32|33|The LORD replied to Moses, "Whoever has sinned against me I will blot out of my book.
EXOD|32|34|Now go, lead the people to the place I spoke of, and my angel will go before you. However, when the time comes for me to punish, I will punish them for their sin."
EXOD|32|35|And the LORD struck the people with a plague because of what they did with the calf Aaron had made.
EXOD|33|1|Then the LORD said to Moses, "Leave this place, you and the people you brought up out of Egypt, and go up to the land I promised on oath to Abraham, Isaac and Jacob, saying, 'I will give it to your descendants.'
EXOD|33|2|I will send an angel before you and drive out the Canaanites, Amorites, Hittites, Perizzites, Hivites and Jebusites.
EXOD|33|3|Go up to the land flowing with milk and honey. But I will not go with you, because you are a stiff-necked people and I might destroy you on the way."
EXOD|33|4|When the people heard these distressing words, they began to mourn and no one put on any ornaments.
EXOD|33|5|For the LORD had said to Moses, "Tell the Israelites, 'You are a stiff-necked people. If I were to go with you even for a moment, I might destroy you. Now take off your ornaments and I will decide what to do with you.'"
EXOD|33|6|So the Israelites stripped off their ornaments at Mount Horeb.
EXOD|33|7|Now Moses used to take a tent and pitch it outside the camp some distance away, calling it the "tent of meeting." Anyone inquiring of the LORD would go to the tent of meeting outside the camp.
EXOD|33|8|And whenever Moses went out to the tent, all the people rose and stood at the entrances to their tents, watching Moses until he entered the tent.
EXOD|33|9|As Moses went into the tent, the pillar of cloud would come down and stay at the entrance, while the LORD spoke with Moses.
EXOD|33|10|Whenever the people saw the pillar of cloud standing at the entrance to the tent, they all stood and worshiped, each at the entrance to his tent.
EXOD|33|11|The LORD would speak to Moses face to face, as a man speaks with his friend. Then Moses would return to the camp, but his young aide Joshua son of Nun did not leave the tent.
EXOD|33|12|Moses said to the LORD, "You have been telling me, 'Lead these people,' but you have not let me know whom you will send with me. You have said, 'I know you by name and you have found favor with me.'
EXOD|33|13|If you are pleased with me, teach me your ways so I may know you and continue to find favor with you. Remember that this nation is your people."
EXOD|33|14|The LORD replied, "My Presence will go with you, and I will give you rest."
EXOD|33|15|Then Moses said to him, "If your Presence does not go with us, do not send us up from here.
EXOD|33|16|How will anyone know that you are pleased with me and with your people unless you go with us? What else will distinguish me and your people from all the other people on the face of the earth?"
EXOD|33|17|And the LORD said to Moses, "I will do the very thing you have asked, because I am pleased with you and I know you by name."
EXOD|33|18|Then Moses said, "Now show me your glory."
EXOD|33|19|And the LORD said, "I will cause all my goodness to pass in front of you, and I will proclaim my name, the LORD, in your presence. I will have mercy on whom I will have mercy, and I will have compassion on whom I will have compassion.
EXOD|33|20|But," he said, "you cannot see my face, for no one may see me and live."
EXOD|33|21|Then the LORD said, "There is a place near me where you may stand on a rock.
EXOD|33|22|When my glory passes by, I will put you in a cleft in the rock and cover you with my hand until I have passed by.
EXOD|33|23|Then I will remove my hand and you will see my back; but my face must not be seen."
EXOD|34|1|The LORD said to Moses, "Chisel out two stone tablets like the first ones, and I will write on them the words that were on the first tablets, which you broke.
EXOD|34|2|Be ready in the morning, and then come up on Mount Sinai. Present yourself to me there on top of the mountain.
EXOD|34|3|No one is to come with you or be seen anywhere on the mountain; not even the flocks and herds may graze in front of the mountain."
EXOD|34|4|So Moses chiseled out two stone tablets like the first ones and went up Mount Sinai early in the morning, as the LORD had commanded him; and he carried the two stone tablets in his hands.
EXOD|34|5|Then the LORD came down in the cloud and stood there with him and proclaimed his name, the LORD.
EXOD|34|6|And he passed in front of Moses, proclaiming, "The LORD, the LORD, the compassionate and gracious God, slow to anger, abounding in love and faithfulness,
EXOD|34|7|maintaining love to thousands, and forgiving wickedness, rebellion and sin. Yet he does not leave the guilty unpunished; he punishes the children and their children for the sin of the fathers to the third and fourth generation."
EXOD|34|8|Moses bowed to the ground at once and worshiped.
EXOD|34|9|"O Lord, if I have found favor in your eyes," he said, "then let the Lord go with us. Although this is a stiff-necked people, forgive our wickedness and our sin, and take us as your inheritance."
EXOD|34|10|Then the LORD said: "I am making a covenant with you. Before all your people I will do wonders never before done in any nation in all the world. The people you live among will see how awesome is the work that I, the LORD, will do for you.
EXOD|34|11|Obey what I command you today. I will drive out before you the Amorites, Canaanites, Hittites, Perizzites, Hivites and Jebusites.
EXOD|34|12|Be careful not to make a treaty with those who live in the land where you are going, or they will be a snare among you.
EXOD|34|13|Break down their altars, smash their sacred stones and cut down their Asherah poles.
EXOD|34|14|Do not worship any other god, for the LORD, whose name is Jealous, is a jealous God.
EXOD|34|15|"Be careful not to make a treaty with those who live in the land; for when they prostitute themselves to their gods and sacrifice to them, they will invite you and you will eat their sacrifices.
EXOD|34|16|And when you choose some of their daughters as wives for your sons and those daughters prostitute themselves to their gods, they will lead your sons to do the same.
EXOD|34|17|"Do not make cast idols.
EXOD|34|18|"Celebrate the Feast of Unleavened Bread. For seven days eat bread made without yeast, as I commanded you. Do this at the appointed time in the month of Abib, for in that month you came out of Egypt.
EXOD|34|19|"The first offspring of every womb belongs to me, including all the firstborn males of your livestock, whether from herd or flock.
EXOD|34|20|Redeem the firstborn donkey with a lamb, but if you do not redeem it, break its neck. Redeem all your firstborn sons. "No one is to appear before me empty-handed.
EXOD|34|21|"Six days you shall labor, but on the seventh day you shall rest; even during the plowing season and harvest you must rest.
EXOD|34|22|"Celebrate the Feast of Weeks with the firstfruits of the wheat harvest, and the Feast of Ingathering at the turn of the year.
EXOD|34|23|Three times a year all your men are to appear before the Sovereign LORD, the God of Israel.
EXOD|34|24|I will drive out nations before you and enlarge your territory, and no one will covet your land when you go up three times each year to appear before the LORD your God.
EXOD|34|25|"Do not offer the blood of a sacrifice to me along with anything containing yeast, and do not let any of the sacrifice from the Passover Feast remain until morning.
EXOD|34|26|"Bring the best of the firstfruits of your soil to the house of the LORD your God. "Do not cook a young goat in its mother's milk."
EXOD|34|27|Then the LORD said to Moses, "Write down these words, for in accordance with these words I have made a covenant with you and with Israel."
EXOD|34|28|Moses was there with the LORD forty days and forty nights without eating bread or drinking water. And he wrote on the tablets the words of the covenant-the Ten Commandments.
EXOD|34|29|When Moses came down from Mount Sinai with the two tablets of the Testimony in his hands, he was not aware that his face was radiant because he had spoken with the LORD.
EXOD|34|30|When Aaron and all the Israelites saw Moses, his face was radiant, and they were afraid to come near him.
EXOD|34|31|But Moses called to them; so Aaron and all the leaders of the community came back to him, and he spoke to them.
EXOD|34|32|Afterward all the Israelites came near him, and he gave them all the commands the LORD had given him on Mount Sinai.
EXOD|34|33|When Moses finished speaking to them, he put a veil over his face.
EXOD|34|34|But whenever he entered the LORD's presence to speak with him, he removed the veil until he came out. And when he came out and told the Israelites what he had been commanded,
EXOD|34|35|they saw that his face was radiant. Then Moses would put the veil back over his face until he went in to speak with the LORD.
EXOD|35|1|Moses assembled the whole Israelite community and said to them, "These are the things the LORD has commanded you to do:
EXOD|35|2|For six days, work is to be done, but the seventh day shall be your holy day, a Sabbath of rest to the LORD. Whoever does any work on it must be put to death.
EXOD|35|3|Do not light a fire in any of your dwellings on the Sabbath day."
EXOD|35|4|Moses said to the whole Israelite community, "This is what the LORD has commanded:
EXOD|35|5|From what you have, take an offering for the LORD. Everyone who is willing is to bring to the LORD an offering of gold, silver and bronze;
EXOD|35|6|blue, purple and scarlet yarn and fine linen; goat hair;
EXOD|35|7|ram skins dyed red and hides of sea cows; acacia wood;
EXOD|35|8|olive oil for the light; spices for the anointing oil and for the fragrant incense;
EXOD|35|9|and onyx stones and other gems to be mounted on the ephod and breastpiece.
EXOD|35|10|"All who are skilled among you are to come and make everything the LORD has commanded:
EXOD|35|11|the tabernacle with its tent and its covering, clasps, frames, crossbars, posts and bases;
EXOD|35|12|the ark with its poles and the atonement cover and the curtain that shields it;
EXOD|35|13|the table with its poles and all its articles and the bread of the Presence;
EXOD|35|14|the lampstand that is for light with its accessories, lamps and oil for the light;
EXOD|35|15|the altar of incense with its poles, the anointing oil and the fragrant incense; the curtain for the doorway at the entrance to the tabernacle;
EXOD|35|16|the altar of burnt offering with its bronze grating, its poles and all its utensils; the bronze basin with its stand;
EXOD|35|17|the curtains of the courtyard with its posts and bases, and the curtain for the entrance to the courtyard;
EXOD|35|18|the tent pegs for the tabernacle and for the courtyard, and their ropes;
EXOD|35|19|the woven garments worn for ministering in the sanctuary-both the sacred garments for Aaron the priest and the garments for his sons when they serve as priests."
EXOD|35|20|Then the whole Israelite community withdrew from Moses' presence,
EXOD|35|21|and everyone who was willing and whose heart moved him came and brought an offering to the LORD for the work on the Tent of Meeting, for all its service, and for the sacred garments.
EXOD|35|22|All who were willing, men and women alike, came and brought gold jewelry of all kinds: brooches, earrings, rings and ornaments. They all presented their gold as a wave offering to the LORD.
EXOD|35|23|Everyone who had blue, purple or scarlet yarn or fine linen, or goat hair, ram skins dyed red or hides of sea cows brought them.
EXOD|35|24|Those presenting an offering of silver or bronze brought it as an offering to the LORD, and everyone who had acacia wood for any part of the work brought it.
EXOD|35|25|Every skilled woman spun with her hands and brought what she had spun-blue, purple or scarlet yarn or fine linen.
EXOD|35|26|And all the women who were willing and had the skill spun the goat hair.
EXOD|35|27|The leaders brought onyx stones and other gems to be mounted on the ephod and breastpiece.
EXOD|35|28|They also brought spices and olive oil for the light and for the anointing oil and for the fragrant incense.
EXOD|35|29|All the Israelite men and women who were willing brought to the LORD freewill offerings for all the work the LORD through Moses had commanded them to do.
EXOD|35|30|Then Moses said to the Israelites, "See, the LORD has chosen Bezalel son of Uri, the son of Hur, of the tribe of Judah,
EXOD|35|31|and he has filled him with the Spirit of God, with skill, ability and knowledge in all kinds of crafts-
EXOD|35|32|to make artistic designs for work in gold, silver and bronze,
EXOD|35|33|to cut and set stones, to work in wood and to engage in all kinds of artistic craftsmanship.
EXOD|35|34|And he has given both him and Oholiab son of Ahisamach, of the tribe of Dan, the ability to teach others.
EXOD|35|35|He has filled them with skill to do all kinds of work as craftsmen, designers, embroiderers in blue, purple and scarlet yarn and fine linen, and weavers-all of them master craftsmen and designers.
EXOD|36|1|So Bezalel, Oholiab and every skilled person to whom the LORD has given skill and ability to know how to carry out all the work of constructing the sanctuary are to do the work just as the LORD has commanded."
EXOD|36|2|Then Moses summoned Bezalel and Oholiab and every skilled person to whom the LORD had given ability and who was willing to come and do the work.
EXOD|36|3|They received from Moses all the offerings the Israelites had brought to carry out the work of constructing the sanctuary. And the people continued to bring freewill offerings morning after morning.
EXOD|36|4|So all the skilled craftsmen who were doing all the work on the sanctuary left their work
EXOD|36|5|and said to Moses, "The people are bringing more than enough for doing the work the LORD commanded to be done."
EXOD|36|6|Then Moses gave an order and they sent this word throughout the camp: "No man or woman is to make anything else as an offering for the sanctuary." And so the people were restrained from bringing more,
EXOD|36|7|because what they already had was more than enough to do all the work.
EXOD|36|8|All the skilled men among the workmen made the tabernacle with ten curtains of finely twisted linen and blue, purple and scarlet yarn, with cherubim worked into them by a skilled craftsman.
EXOD|36|9|All the curtains were the same size-twenty-eight cubits long and four cubits wide.
EXOD|36|10|They joined five of the curtains together and did the same with the other five.
EXOD|36|11|Then they made loops of blue material along the edge of the end curtain in one set, and the same was done with the end curtain in the other set.
EXOD|36|12|They also made fifty loops on one curtain and fifty loops on the end curtain of the other set, with the loops opposite each other.
EXOD|36|13|Then they made fifty gold clasps and used them to fasten the two sets of curtains together so that the tabernacle was a unit.
EXOD|36|14|They made curtains of goat hair for the tent over the tabernacle-eleven altogether.
EXOD|36|15|All eleven curtains were the same size-thirty cubits long and four cubits wide.
EXOD|36|16|They joined five of the curtains into one set and the other six into another set.
EXOD|36|17|Then they made fifty loops along the edge of the end curtain in one set and also along the edge of the end curtain in the other set.
EXOD|36|18|They made fifty bronze clasps to fasten the tent together as a unit.
EXOD|36|19|Then they made for the tent a covering of ram skins dyed red, and over that a covering of hides of sea cows.
EXOD|36|20|They made upright frames of acacia wood for the tabernacle.
EXOD|36|21|Each frame was ten cubits long and a cubit and a half wide,
EXOD|36|22|with two projections set parallel to each other. They made all the frames of the tabernacle in this way.
EXOD|36|23|They made twenty frames for the south side of the tabernacle
EXOD|36|24|and made forty silver bases to go under them-two bases for each frame, one under each projection.
EXOD|36|25|For the other side, the north side of the tabernacle, they made twenty frames
EXOD|36|26|and forty silver bases-two under each frame.
EXOD|36|27|They made six frames for the far end, that is, the west end of the tabernacle,
EXOD|36|28|and two frames were made for the corners of the tabernacle at the far end.
EXOD|36|29|At these two corners the frames were double from the bottom all the way to the top and fitted into a single ring; both were made alike.
EXOD|36|30|So there were eight frames and sixteen silver bases-two under each frame.
EXOD|36|31|They also made crossbars of acacia wood: five for the frames on one side of the tabernacle,
EXOD|36|32|five for those on the other side, and five for the frames on the west, at the far end of the tabernacle.
EXOD|36|33|They made the center crossbar so that it extended from end to end at the middle of the frames.
EXOD|36|34|They overlaid the frames with gold and made gold rings to hold the crossbars. They also overlaid the crossbars with gold.
EXOD|36|35|They made the curtain of blue, purple and scarlet yarn and finely twisted linen, with cherubim worked into it by a skilled craftsman.
EXOD|36|36|They made four posts of acacia wood for it and overlaid them with gold. They made gold hooks for them and cast their four silver bases.
EXOD|36|37|For the entrance to the tent they made a curtain of blue, purple and scarlet yarn and finely twisted linen-the work of an embroiderer;
EXOD|36|38|and they made five posts with hooks for them. They overlaid the tops of the posts and their bands with gold and made their five bases of bronze.
EXOD|37|1|Bezalel made the ark of acacia wood-two and a half cubits long, a cubit and a half wide, and a cubit and a half high.
EXOD|37|2|He overlaid it with pure gold, both inside and out, and made a gold molding around it.
EXOD|37|3|He cast four gold rings for it and fastened them to its four feet, with two rings on one side and two rings on the other.
EXOD|37|4|Then he made poles of acacia wood and overlaid them with gold.
EXOD|37|5|And he inserted the poles into the rings on the sides of the ark to carry it.
EXOD|37|6|He made the atonement cover of pure gold-two and a half cubits long and a cubit and a half wide.
EXOD|37|7|Then he made two cherubim out of hammered gold at the ends of the cover.
EXOD|37|8|He made one cherub on one end and the second cherub on the other; at the two ends he made them of one piece with the cover.
EXOD|37|9|The cherubim had their wings spread upward, overshadowing the cover with them. The cherubim faced each other, looking toward the cover.
EXOD|37|10|They made the table of acacia wood-two cubits long, a cubit wide, and a cubit and a half high.
EXOD|37|11|Then they overlaid it with pure gold and made a gold molding around it.
EXOD|37|12|They also made around it a rim a handbreadth wide and put a gold molding on the rim.
EXOD|37|13|They cast four gold rings for the table and fastened them to the four corners, where the four legs were.
EXOD|37|14|The rings were put close to the rim to hold the poles used in carrying the table.
EXOD|37|15|The poles for carrying the table were made of acacia wood and were overlaid with gold.
EXOD|37|16|And they made from pure gold the articles for the table-its plates and dishes and bowls and its pitchers for the pouring out of drink offerings.
EXOD|37|17|They made the lampstand of pure gold and hammered it out, base and shaft; its flowerlike cups, buds and blossoms were of one piece with it.
EXOD|37|18|Six branches extended from the sides of the lampstand-three on one side and three on the other.
EXOD|37|19|Three cups shaped like almond flowers with buds and blossoms were on one branch, three on the next branch and the same for all six branches extending from the lampstand.
EXOD|37|20|And on the lampstand were four cups shaped like almond flowers with buds and blossoms.
EXOD|37|21|One bud was under the first pair of branches extending from the lampstand, a second bud under the second pair, and a third bud under the third pair-six branches in all.
EXOD|37|22|The buds and the branches were all of one piece with the lampstand, hammered out of pure gold.
EXOD|37|23|They made its seven lamps, as well as its wick trimmers and trays, of pure gold.
EXOD|37|24|They made the lampstand and all its accessories from one talent of pure gold.
EXOD|37|25|They made the altar of incense out of acacia wood. It was square, a cubit long and a cubit wide, and two cubits high -its horns of one piece with it.
EXOD|37|26|They overlaid the top and all the sides and the horns with pure gold, and made a gold molding around it.
EXOD|37|27|They made two gold rings below the molding-two on opposite sides-to hold the poles used to carry it.
EXOD|37|28|They made the poles of acacia wood and overlaid them with gold.
EXOD|37|29|They also made the sacred anointing oil and the pure, fragrant incense-the work of a perfumer.
EXOD|38|1|They built the altar of burnt offering of acacia wood, three cubits high; it was square, five cubits long and five cubits wide.
EXOD|38|2|They made a horn at each of the four corners, so that the horns and the altar were of one piece, and they overlaid the altar with bronze.
EXOD|38|3|They made all its utensils of bronze-its pots, shovels, sprinkling bowls, meat forks and firepans.
EXOD|38|4|They made a grating for the altar, a bronze network, to be under its ledge, halfway up the altar.
EXOD|38|5|They cast bronze rings to hold the poles for the four corners of the bronze grating.
EXOD|38|6|They made the poles of acacia wood and overlaid them with bronze.
EXOD|38|7|They inserted the poles into the rings so they would be on the sides of the altar for carrying it. They made it hollow, out of boards.
EXOD|38|8|They made the bronze basin and its bronze stand from the mirrors of the women who served at the entrance to the Tent of Meeting.
EXOD|38|9|Next they made the courtyard. The south side was a hundred cubits long and had curtains of finely twisted linen,
EXOD|38|10|with twenty posts and twenty bronze bases, and with silver hooks and bands on the posts.
EXOD|38|11|The north side was also a hundred cubits long and had twenty posts and twenty bronze bases, with silver hooks and bands on the posts.
EXOD|38|12|The west end was fifty cubits wide and had curtains, with ten posts and ten bases, with silver hooks and bands on the posts.
EXOD|38|13|The east end, toward the sunrise, was also fifty cubits wide.
EXOD|38|14|Curtains fifteen cubits long were on one side of the entrance, with three posts and three bases,
EXOD|38|15|and curtains fifteen cubits long were on the other side of the entrance to the courtyard, with three posts and three bases.
EXOD|38|16|All the curtains around the courtyard were of finely twisted linen.
EXOD|38|17|The bases for the posts were bronze. The hooks and bands on the posts were silver, and their tops were overlaid with silver; so all the posts of the courtyard had silver bands.
EXOD|38|18|The curtain for the entrance to the courtyard was of blue, purple and scarlet yarn and finely twisted linen-the work of an embroiderer. It was twenty cubits long and, like the curtains of the courtyard, five cubits high,
EXOD|38|19|with four posts and four bronze bases. Their hooks and bands were silver, and their tops were overlaid with silver.
EXOD|38|20|All the tent pegs of the tabernacle and of the surrounding courtyard were bronze.
EXOD|38|21|These are the amounts of the materials used for the tabernacle, the tabernacle of the Testimony, which were recorded at Moses' command by the Levites under the direction of Ithamar son of Aaron, the priest.
EXOD|38|22|(Bezalel son of Uri, the son of Hur, of the tribe of Judah, made everything the LORD commanded Moses;
EXOD|38|23|with him was Oholiab son of Ahisamach, of the tribe of Dan-a craftsman and designer, and an embroiderer in blue, purple and scarlet yarn and fine linen.)
EXOD|38|24|The total amount of the gold from the wave offering used for all the work on the sanctuary was 29 talents and 730 shekels, according to the sanctuary shekel.
EXOD|38|25|The silver obtained from those of the community who were counted in the census was 100 talents and 1,775 shekels, according to the sanctuary shekel-
EXOD|38|26|one beka per person, that is, half a shekel, according to the sanctuary shekel, from everyone who had crossed over to those counted, twenty years old or more, a total of 603,550 men.
EXOD|38|27|The 100 talents of silver were used to cast the bases for the sanctuary and for the curtain-100 bases from the 100 talents, one talent for each base.
EXOD|38|28|They used the 1,775 shekels to make the hooks for the posts, to overlay the tops of the posts, and to make their bands.
EXOD|38|29|The bronze from the wave offering was 70 talents and 2,400 shekels.
EXOD|38|30|They used it to make the bases for the entrance to the Tent of Meeting, the bronze altar with its bronze grating and all its utensils,
EXOD|38|31|the bases for the surrounding courtyard and those for its entrance and all the tent pegs for the tabernacle and those for the surrounding courtyard.
EXOD|39|1|From the blue, purple and scarlet yarn they made woven garments for ministering in the sanctuary. They also made sacred garments for Aaron, as the LORD commanded Moses.
EXOD|39|2|They made the ephod of gold, and of blue, purple and scarlet yarn, and of finely twisted linen.
EXOD|39|3|They hammered out thin sheets of gold and cut strands to be worked into the blue, purple and scarlet yarn and fine linen-the work of a skilled craftsman.
EXOD|39|4|They made shoulder pieces for the ephod, which were attached to two of its corners, so it could be fastened.
EXOD|39|5|Its skillfully woven waistband was like it-of one piece with the ephod and made with gold, and with blue, purple and scarlet yarn, and with finely twisted linen, as the LORD commanded Moses.
EXOD|39|6|They mounted the onyx stones in gold filigree settings and engraved them like a seal with the names of the sons of Israel.
EXOD|39|7|Then they fastened them on the shoulder pieces of the ephod as memorial stones for the sons of Israel, as the LORD commanded Moses.
EXOD|39|8|They fashioned the breastpiece-the work of a skilled craftsman. They made it like the ephod: of gold, and of blue, purple and scarlet yarn, and of finely twisted linen.
EXOD|39|9|It was square-a span long and a span wide-and folded double.
EXOD|39|10|Then they mounted four rows of precious stones on it. In the first row there was a ruby, a topaz and a beryl;
EXOD|39|11|in the second row a turquoise, a sapphire and an emerald;
EXOD|39|12|in the third row a jacinth, an agate and an amethyst;
EXOD|39|13|in the fourth row a chrysolite, an onyx and a jasper. They were mounted in gold filigree settings.
EXOD|39|14|There were twelve stones, one for each of the names of the sons of Israel, each engraved like a seal with the name of one of the twelve tribes.
EXOD|39|15|For the breastpiece they made braided chains of pure gold, like a rope.
EXOD|39|16|They made two gold filigree settings and two gold rings, and fastened the rings to two of the corners of the breastpiece.
EXOD|39|17|They fastened the two gold chains to the rings at the corners of the breastpiece,
EXOD|39|18|and the other ends of the chains to the two settings, attaching them to the shoulder pieces of the ephod at the front.
EXOD|39|19|They made two gold rings and attached them to the other two corners of the breastpiece on the inside edge next to the ephod.
EXOD|39|20|Then they made two more gold rings and attached them to the bottom of the shoulder pieces on the front of the ephod, close to the seam just above the waistband of the ephod.
EXOD|39|21|They tied the rings of the breastpiece to the rings of the ephod with blue cord, connecting it to the waistband so that the breastpiece would not swing out from the ephod-as the LORD commanded Moses.
EXOD|39|22|They made the robe of the ephod entirely of blue cloth-the work of a weaver-
EXOD|39|23|with an opening in the center of the robe like the opening of a collar, and a band around this opening, so that it would not tear.
EXOD|39|24|They made pomegranates of blue, purple and scarlet yarn and finely twisted linen around the hem of the robe.
EXOD|39|25|And they made bells of pure gold and attached them around the hem between the pomegranates.
EXOD|39|26|The bells and pomegranates alternated around the hem of the robe to be worn for ministering, as the LORD commanded Moses.
EXOD|39|27|For Aaron and his sons, they made tunics of fine linen-the work of a weaver-
EXOD|39|28|and the turban of fine linen, the linen headbands and the undergarments of finely twisted linen.
EXOD|39|29|The sash was of finely twisted linen and blue, purple and scarlet yarn-the work of an embroiderer-as the LORD commanded Moses.
EXOD|39|30|They made the plate, the sacred diadem, out of pure gold and engraved on it, like an inscription on a seal: HOLY TO THE LORD.
EXOD|39|31|Then they fastened a blue cord to it to attach it to the turban, as the LORD commanded Moses.
EXOD|39|32|So all the work on the tabernacle, the Tent of Meeting, was completed. The Israelites did everything just as the LORD commanded Moses.
EXOD|39|33|Then they brought the tabernacle to Moses: the tent and all its furnishings, its clasps, frames, crossbars, posts and bases;
EXOD|39|34|the covering of ram skins dyed red, the covering of hides of sea cows and the shielding curtain;
EXOD|39|35|the ark of the Testimony with its poles and the atonement cover;
EXOD|39|36|the table with all its articles and the bread of the Presence;
EXOD|39|37|the pure gold lampstand with its row of lamps and all its accessories, and the oil for the light;
EXOD|39|38|the gold altar, the anointing oil, the fragrant incense, and the curtain for the entrance to the tent;
EXOD|39|39|the bronze altar with its bronze grating, its poles and all its utensils; the basin with its stand;
EXOD|39|40|the curtains of the courtyard with its posts and bases, and the curtain for the entrance to the courtyard; the ropes and tent pegs for the courtyard; all the furnishings for the tabernacle, the Tent of Meeting;
EXOD|39|41|and the woven garments worn for ministering in the sanctuary, both the sacred garments for Aaron the priest and the garments for his sons when serving as priests.
EXOD|39|42|The Israelites had done all the work just as the LORD had commanded Moses.
EXOD|39|43|Moses inspected the work and saw that they had done it just as the LORD had commanded. So Moses blessed them.
EXOD|40|1|Then the LORD said to Moses:
EXOD|40|2|"Set up the tabernacle, the Tent of Meeting, on the first day of the first month.
EXOD|40|3|Place the ark of the Testimony in it and shield the ark with the curtain.
EXOD|40|4|Bring in the table and set out what belongs on it. Then bring in the lampstand and set up its lamps.
EXOD|40|5|Place the gold altar of incense in front of the ark of the Testimony and put the curtain at the entrance to the tabernacle.
EXOD|40|6|"Place the altar of burnt offering in front of the entrance to the tabernacle, the Tent of Meeting;
EXOD|40|7|place the basin between the Tent of Meeting and the altar and put water in it.
EXOD|40|8|Set up the courtyard around it and put the curtain at the entrance to the courtyard.
EXOD|40|9|"Take the anointing oil and anoint the tabernacle and everything in it; consecrate it and all its furnishings, and it will be holy.
EXOD|40|10|Then anoint the altar of burnt offering and all its utensils; consecrate the altar, and it will be most holy.
EXOD|40|11|Anoint the basin and its stand and consecrate them.
EXOD|40|12|"Bring Aaron and his sons to the entrance to the Tent of Meeting and wash them with water.
EXOD|40|13|Then dress Aaron in the sacred garments, anoint him and consecrate him so he may serve me as priest.
EXOD|40|14|Bring his sons and dress them in tunics.
EXOD|40|15|Anoint them just as you anointed their father, so they may serve me as priests. Their anointing will be to a priesthood that will continue for all generations to come."
EXOD|40|16|Moses did everything just as the LORD commanded him.
EXOD|40|17|So the tabernacle was set up on the first day of the first month in the second year.
EXOD|40|18|When Moses set up the tabernacle, he put the bases in place, erected the frames, inserted the crossbars and set up the posts.
EXOD|40|19|Then he spread the tent over the tabernacle and put the covering over the tent, as the LORD commanded him.
EXOD|40|20|He took the Testimony and placed it in the ark, attached the poles to the ark and put the atonement cover over it.
EXOD|40|21|Then he brought the ark into the tabernacle and hung the shielding curtain and shielded the ark of the Testimony, as the LORD commanded him.
EXOD|40|22|Moses placed the table in the Tent of Meeting on the north side of the tabernacle outside the curtain
EXOD|40|23|and set out the bread on it before the LORD, as the LORD commanded him.
EXOD|40|24|He placed the lampstand in the Tent of Meeting opposite the table on the south side of the tabernacle
EXOD|40|25|and set up the lamps before the LORD, as the LORD commanded him.
EXOD|40|26|Moses placed the gold altar in the Tent of Meeting in front of the curtain
EXOD|40|27|and burned fragrant incense on it, as the LORD commanded him.
EXOD|40|28|Then he put up the curtain at the entrance to the tabernacle.
EXOD|40|29|He set the altar of burnt offering near the entrance to the tabernacle, the Tent of Meeting, and offered on it burnt offerings and grain offerings, as the LORD commanded him.
EXOD|40|30|He placed the basin between the Tent of Meeting and the altar and put water in it for washing,
EXOD|40|31|and Moses and Aaron and his sons used it to wash their hands and feet.
EXOD|40|32|They washed whenever they entered the Tent of Meeting or approached the altar, as the LORD commanded Moses.
EXOD|40|33|Then Moses set up the courtyard around the tabernacle and altar and put up the curtain at the entrance to the courtyard. And so Moses finished the work.
EXOD|40|34|Then the cloud covered the Tent of Meeting, and the glory of the Lord filled the tabernacle.
EXOD|40|35|Moses could not enter the Tent of Meeting because the cloud had settled upon it, and the glory of the LORD filled the tabernacle.
EXOD|40|36|In all the travels of the Israelites, whenever the cloud lifted from above the tabernacle, they would set out;
EXOD|40|37|but if the cloud did not lift, they did not set out-until the day it lifted.
EXOD|40|38|So the cloud of the LORD was over the tabernacle by day, and fire was in the cloud by night, in the sight of all the house of Israel during all their travels.
