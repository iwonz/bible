1TIM|1|1|Paulus, apostolus Christi Iesu secundum praeceptum Dei sal vatoris nostri et Christi Iesu spei nostrae,
1TIM|1|2|Timotheo germano filio in fide: gratia, misericordia, pax a Deo Patre et Christo Iesu Domino nostro.
1TIM|1|3|Sicut rogavi te, ut remaneres Ephesi, cum irem in Macedoniam, ut praeciperes quibusdam, ne aliter docerent
1TIM|1|4|neque intenderent fabulis et genealogiis interminatis, quae quaestiones praestant magis quam dispensationem Dei, quae est in fide;
1TIM|1|5|finis autem praecepti est caritas de corde puro et conscientia bona et fide non ficta,
1TIM|1|6|a quibus quidam aberrantes conversi sunt in vaniloquium,
1TIM|1|7|volentes esse legis doctores, non intellegentes neque quae loquuntur neque de quibus affirmant.
1TIM|1|8|Scimus autem quia bona est lex, si quis ea legitime utatur,
1TIM|1|9|sciens hoc quia iusto lex non est posita sed iniustis et non subiectis, impiis et peccatoribus, sceleratis et contaminatis, patricidis et matricidis, homicidis,
1TIM|1|10|fornicariis, masculorum concubitoribus, plagiariis, mendacibus, periuris et si quid aliud sanae doctrinae adversatur,
1TIM|1|11|secundum evangelium gloriae beati Dei, quod creditum est mihi.
1TIM|1|12|Gratiam habeo ei, qui me confortavit, Christo Iesu Domino nostro, quia fidelem me existimavit ponens in ministerio,
1TIM|1|13|qui prius fui blasphemus et persecutor et contumeliosus; sed misericordiam consecutus sum, quia ignorans feci in incredulitate;
1TIM|1|14|superabundavit autem gratia Domini nostri cum fide et dilectione, quae sunt in Christo Iesu.
1TIM|1|15|Fidelis sermo et omni acceptione dignus: Christus Iesus venit in mundum peccatores salvos facere; quorum primus ego sum,
1TIM|1|16|sed ideo misericordiam consecutus sum, ut in me primo ostenderet Christus Iesus omnem longanimitatem, ad informationem eorum, qui credituri sunt illi in vitam aeternam.
1TIM|1|17|Regi autem saeculorum, incorruptibili, invisibili, soli Deo honor et gloria in saecula saeculorum. Amen.
1TIM|1|18|Hoc praeceptum commendo tibi, fili Timothee, secundum praecedentes super te prophetias, ut milites in illis bonam militiam
1TIM|1|19|habens fidem et bonam conscientiam, quam quidam repellentes circa fidem naufragaverunt;
1TIM|1|20|ex quibus est Hymenaeus et Alexander, quos tradidi Satanae, ut discant non blasphemare.
1TIM|2|1|Obsecro igitur primo omnium fieri obsecrationes, orationes, postulationes, gratiarum actiones pro omnibus hominibus,
1TIM|2|2|pro regibus et omnibus, qui in sublimitate sunt, ut quietam et tranquillam vitam agamus in omni pietate et castitate.
1TIM|2|3|Hoc bonum est et acceptum coram salvatore nostro Deo,
1TIM|2|4|qui omnes homines vult salvos fieri et ad agnitionem veritatis venire.
1TIM|2|5|Unus enim Deus, unus et mediator Dei et hominum, homo Christus Iesus,
1TIM|2|6|qui dedit redemptionem semetipsum pro omnibus, testimonium temporibus suis;
1TIM|2|7|in quod positus sum ego praedicator et apostolus - veritatem dico, non mentior - doctor gentium in fide et veritate.
1TIM|2|8|Volo ergo viros orare in omni loco levantes puras manus sine ira et disceptatione;
1TIM|2|9|similiter et mulieres in habitu ornato cum verecundia et sobrietate ornantes se, non in tortis crinibus et auro aut margaritis vel veste pretiosa,
1TIM|2|10|sed, quod decet mulieres, profitentes pietatem per opera bona.
1TIM|2|11|Mulier in tranquillitate discat cum omni subiectione;
1TIM|2|12|docere autem mulieri non permitto neque dominari in virum, sed esse in tranquillitate.
1TIM|2|13|Adam enim primus formatus est, deinde Eva;
1TIM|2|14|et Adam non est seductus, mulier autem seducta in praevaricatione fuit.
1TIM|2|15|Salvabitur autem per filiorum generationem, si permanserint in fide et dilectione et sanctificatione cum sobrietate.
1TIM|3|1|Fidelis sermo: si quis episco patum appetit, bonum opus de siderat.
1TIM|3|2|Oportet ergo episcopum irreprehensibilem esse, unius uxoris virum, sobrium, prudentem, ornatum, hospitalem, doctorem,
1TIM|3|3|non vinolentum, non percussorem sed modestum, non litigiosum, non cupidum,
1TIM|3|4|suae domui bene praepositum, filios habentem in subiectione cum omni castitate
1TIM|3|5|- si quis autem domui suae praeesse nescit, quomodo ecclesiae Dei curam habebit? C,
1TIM|3|6|non neophytum, ne in superbia elatus in iudicium incidat Diaboli.
1TIM|3|7|Oportet autem illum et testimonium habere bonum ab his, qui foris sunt, ut non in opprobrium incidat et laqueum Diaboli.
1TIM|3|8|Diaconos similiter pudicos, non bilingues, non multo vino deditos, non turpe lucrum sectantes,
1TIM|3|9|habentes mysterium fidei in conscientia pura.
1TIM|3|10|Et hi autem probentur primum, deinde ministrent nullum crimen habentes.
1TIM|3|11|Mulieres similiter pudicas, non detrahentes, sobrias, fideles in omnibus.
1TIM|3|12|Diaconi sint unius uxoris viri, qui filiis suis bene praesint et suis domibus;
1TIM|3|13|qui enim bene ministraverint, gradum sibi bonum acquirent et multam fiduciam in fide, quae est in Christo Iesu.
1TIM|3|14|Haec tibi scribo sperans venire ad te cito;
1TIM|3|15|si autem tardavero, ut scias quomodo oporteat in domo Dei conversari, quae est ecclesia Dei vivi, columna et firmamentum veritatis.
1TIM|3|16|Et omnium confessione magnum est pietatis mysterium:Qui manifestatus est in carne,iustificatus est in Spiritu,apparuit angelis,praedicatus est in gentibus,creditus est in mumdo,assumptus est in gloria.
1TIM|4|1|Spiritus autem manifeste dicit, quia in novissimis temporibus discedent quidam a fide, attendentes spiritibus seductoribus et doctrinis daemoniorum,
1TIM|4|2|in hypocrisi loquentium mendacium et cauteriatam habentium suam conscientiam,
1TIM|4|3|prohibentium nubere, abstinere a cibis, quos Deus creavit ad percipiendum cum gratiarum actione fidelibus et his, qui cognoverunt veritatem.
1TIM|4|4|Quia omnis creatura Dei bona, et nihil reiciendum, quod cum gratiarum actione percipitur;
1TIM|4|5|sanctificatur enim per verbum Dei et orationem.
1TIM|4|6|Haec proponens fratribus bonus eris minister Christi Iesu, enutritus verbis fidei et bonae doctrinae, quam assecutus es;
1TIM|4|7|profanas autem et aniles fabulas devita.Exerce teipsum ad pietatem;
1TIM|4|8|nam corporalis exercitatio ad modicum utilis est, pietas autem ad omnia utilis est promissionem habens vitae, quae nunc est, et futurae.
1TIM|4|9|Fidelis sermo et omni acceptione dignus:
1TIM|4|10|in hoc enim laboramus et certamus, quia sperantes sumus in Deum vivum, qui est salvator omnium hominum, maxime fidelium.
1TIM|4|11|Praecipe haec et doce.
1TIM|4|12|Nemo adulescentiam tuam contemnat; sed exemplum esto fidelium in verbo, in conversatione, in caritate, in fide, in castitate.
1TIM|4|13|Dum venio, attende lectioni, exhortationi, doctrinae.
1TIM|4|14|Noli neglegere donationem, quae in te est, quae data est tibi per prophetiam cum impositione manuum presbyterii.
1TIM|4|15|Haec meditare, in his esto, ut profectus tuus manifestus sit omnibus.
1TIM|4|16|Attende tibi et doctrinae; insta in illis; hoc enim faciens et teipsum salvum facies et eos, qui te audiunt.
1TIM|5|1|Seniorem ne increpaveris, sed obsecra ut patrem, iuvenes ut fratres,
1TIM|5|2|anus ut matres, iuvenculas ut sorores in omni castitate.
1TIM|5|3|Viduas honora, quae vere viduae sunt.
1TIM|5|4|Si qua autem vidua filios aut nepotes habet, discant primum domum suam pie regere et mutuam vicem reddere parentibus; hoc enim acceptum est coram Deo.
1TIM|5|5|Quae autem vere vidua est et desolata, sperat in Deum et instat obsecrationibus et orationibus nocte ac die;
1TIM|5|6|nam quae in deliciis est vivens, mortua est.
1TIM|5|7|Et haec praecipe, ut irreprehensibiles sint.
1TIM|5|8|Si quis autem suorum et maxime domesticorum curam non habet, fidem negavit et est infideli deterior.
1TIM|5|9|Vidua adscribatur non minus sexaginta annorum, quae fuerit unius viri uxor,
1TIM|5|10|in operibus bonis testimonium habens: si filios educavit, si hospitio recepit, si sanctorum pedes lavit, si tribulationem patientibus subministravit, si omne opus bonum subsecuta est.
1TIM|5|11|Adulescentiores autem viduas devita; cum enim luxuriatae fuerint adversus Christum, nubere volunt,
1TIM|5|12|habentes damnationem, quia primam fidem irritam fecerunt;
1TIM|5|13|simul autem et otiosae discunt circumire domos, non solum otiosae sed et verbosae et curiosae, loquentes quae non oportet.
1TIM|5|14|Volo ergo iuniores nubere, filios procreare, dominas domus esse, nullam occasionem dare adversario maledicti gratia;
1TIM|5|15|iam enim quaedam conversae sunt retro Satanam.
1TIM|5|16|Si qua fidelis habet viduas, subministret illis, et non gravetur ecclesia, ut his, quae vere viduae sunt, sufficiat.
1TIM|5|17|Qui bene praesunt presbyteri, duplici honore digni habeantur, maxime qui laborant in verbo et doctrina;
1TIM|5|18|dicit enim Scriptura: " Non infrenabis os bovi trituranti " et: " Dignus operarius mercede sua ".
1TIM|5|19|Adversus presbyterum accusationem noli recipere, nisi sub duobus vel tribus testibus.
1TIM|5|20|Peccantes coram omnibus argue, ut et ceteri timorem habeant.
1TIM|5|21|Testificor coram Deo et Christo Iesu et electis angelis, ut haec custodias sine praeiudicio nihil faciens in aliquam partem declinando.
1TIM|5|22|Manus cito nemini imposueris neque communicaveris peccatis alienis; teipsum castum custodi.
1TIM|5|23|Noli adhuc aquam bibere, sed vino modico utere propter stomachum et frequentes tuas infirmitates.
1TIM|5|24|Quorundam hominum peccata manifesta sunt praecedentia ad iudicium, quosdam autem et subsequuntur;
1TIM|5|25|similiter et facta bona manifesta sunt, et, quae aliter se habent, abscondi non possunt.
1TIM|6|1|Quicumque sunt sub iugo, servi dominos suos omni honore di gnos arbitrentur, ne nomen Dei et doctrina blasphemetur.
1TIM|6|2|Qui autem fideles habent dominos, non contemnant, quia fratres sunt, sed magis serviant, quia fideles sunt et dilecti, qui beneficii participes sunt. Haec doce et exhortare.
1TIM|6|3|Si quis aliter docet et non accedit sanis sermonibus Domini nostri Iesu Christi et ei, quae secundum pietatem est, doctrinae,
1TIM|6|4|superbus est, nihil sciens, sed languens circa quaestiones et pugnas verborum, ex quibus oriuntur invidiae, contentiones, blasphemiae, suspiciones malae,
1TIM|6|5|conflictationes hominum mente corruptorum et qui veritate privati sunt, existimantium quaestum esse pietatem.
1TIM|6|6|Est autem quaestus magnus pietas cum sufficientia.
1TIM|6|7|Nihil enim intulimus in mundum, quia nec auferre quid possumus;
1TIM|6|8|habentes autem alimenta et quibus tegamur, his contenti erimus.
1TIM|6|9|Nam qui volunt divites fieri, incidunt in tentationem et laqueum et desideria multa stulta et nociva, quae mergunt homines in interitum et perditionem;
1TIM|6|10|radix enim omnium malorum est cupiditas, quam quidam appetentes erraverunt a fide et inseruerunt se doloribus multis.
1TIM|6|11|Tu autem, o homo Dei, haec fuge; sectare vero iustitiam, pietatem, fidem, caritatem, patientiam, mansuetudinem.
1TIM|6|12|Certa bonum certamen fidei, apprehende vitam aeternam, ad quam vocatus es, et confessus es bonam confessionem coram multis testibus.
1TIM|6|13|Praecipio tibi coram Deo, qui vivificat omnia, et Christo Iesu, qui testimonium reddidit sub Pontio Pilato bonam confessionem,
1TIM|6|14|ut serves mandatum sine macula irreprehensibile usque in adventum Domini nostri Iesu Christi,
1TIM|6|15|quem suis temporibus ostendet beatus et solus potens, Rex regnantium et Dominus dominantium,
1TIM|6|16|qui solus habet immortalitatem, lucem habitans inaccessibilem, quem vidit nullus hominum nec videre potest; cui honor et imperium sempiternum. Amen.
1TIM|6|17|Divitibus huius saeculi praecipe non superbe sapere neque sperare in incerto divitiarum sed in Deo, qui praestat nobis omnia abunde ad fruendum,
1TIM|6|18|bene agere, divites fieri in operibus bonis, facile tribuere, communicare,
1TIM|6|19|thesaurizare sibi fundamentum bonum in futurum, ut apprehendant veram vitam.
1TIM|6|20|O Timothee, depositum custodi, devitans profanas vocum novitates et oppositiones falsi nominis scientiae,
1TIM|6|21|quam quidam profitentes circa fidem aberraverunt.Gratia vobiscum.
