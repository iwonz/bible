EXOD|1|1|Haec sunt nomina filiorum Is rael, qui ingressi sunt Aegyp tum cum Iacob; singuli cum domibus suis introierunt:
EXOD|1|2|Ruben, Simeon, Levi, Iuda,
EXOD|1|3|Issachar, Zabulon et Beniamin,
EXOD|1|4|Dan et Nephthali, Gad et Aser.
EXOD|1|5|Erant igitur omnes animae eorum, qui egressi sunt de femore Iacob, septuaginta; Ioseph autem in Aegypto erat.
EXOD|1|6|Quo mortuo et universis fratribus eius omnique cognatione illa,
EXOD|1|7|filii Israel creverunt et pullulantes multiplicati sunt ac roborati nimis impleverunt terram.
EXOD|1|8|Surrexit interea rex novus super Aegyptum, qui ignorabat Ioseph;
EXOD|1|9|et ait ad populum suum: " Ecce, populus filiorum Israel multus et fortior nobis est;
EXOD|1|10|venite, prudenter agamus cum eo, ne forte multiplicetur et, si ingruerit contra nos bellum, addatur inimicis nostris, expugnatisque nobis, egrediatur de terra ".
EXOD|1|11|Praeposuit itaque eis magistros operum, ut affligerent eos oneribus; aedificaveruntque urbes promptuarias pharaoni, Phithom et Ramesses.
EXOD|1|12|Quantoque opprimebant eos, tanto magis multiplicabantur et crescebant.
EXOD|1|13|Formidaveruntque filios Israel Aegyptii et in servitutem redegerunt eos
EXOD|1|14|atque ad amaritudinem perducebant vitam eorum operibus duris luti et lateris omnique famulatu, quo in terrae operibus premebantur.
EXOD|1|15|Dixit autem rex Aegypti obstetricibus Hebraeorum, quarum una vocabatur Sephra, altera Phua,
EXOD|1|16|praecipiens eis: " Quando obstetricabitis Hebraeas, et partus tempus advenerit, si masculus fuerit, interficite eum; si femina, reservate ".
EXOD|1|17|Timuerunt autem obstetrices Deum et non fecerunt iuxta praeceptum regis Aegypti, sed conservabant mares.
EXOD|1|18|Quibus ad se accersitis rex ait: " Quidnam est hoc, quod facere voluistis, ut pueros servaretis? ".
EXOD|1|19|Quae responderunt: " Non sunt Hebraeae sicut Aegyptiae mulieres; ipsae enim robustae sunt et, priusquam veniamus ad eas, pariunt ".
EXOD|1|20|Bene ergo fecit Deus obstetricibus, et crevit populus confortatusque est nimis;
EXOD|1|21|et, quia timuerunt obstetrices Deum, aedificavit illis domos.
EXOD|1|22|Praecepit ergo pharao omni populo suo dicens: " Quidquid masculini sexus natum fuerit, in flumen proicite; quidquid feminei, reservate ".
EXOD|2|1|Egressus est vir de domo Levi et accepit uxorem stirpis suae;
EXOD|2|2|quae concepit et peperit filium et videns eum elegantem abscondit tribus mensibus.
EXOD|2|3|Cumque iam celare non posset, sumpsit fiscellam scirpeam et linivit eam bitumine ac pice; posuitque intus infantulum et exposuit eum in carecto ripae fluminis,
EXOD|2|4|stante procul sorore eius et considerante eventum rei.
EXOD|2|5|Ecce autem descendebat filia pharaonis, ut lavaretur in flumine, et puellae eius gradiebantur per crepidinem alvei. Quae cum vidisset fiscellam in papyrione, misit unam e famulabus suis; et allatam
EXOD|2|6|aperiens cernensque in ea parvulum vagientem, miserta eius ait: " De infantibus Hebraeorum est hic ".
EXOD|2|7|Cui soror pueri: " Vis, inquit, ut vadam et vocem tibi mulierem Hebraeam, quae nutrire possit tibi infantulum? ".
EXOD|2|8|Respondit: " Vade ". Perrexit puella et vocavit matrem infantis.
EXOD|2|9|Ad quam locuta filia pharaonis: " Accipe, ait, puerum istum et nutri mihi; ego dabo tibi mercedem tuam ". Suscepit mulier et nutrivit puerum adultumque tradidit filiae pharaonis.
EXOD|2|10|Quem illa adoptavit in locum filii vocavitque nomen eius Moysen dicens: " Quia de aqua tuli eum ".
EXOD|2|11|In diebus illis, postquam creverat, Moyses egressus est ad fratres suos; viditque afflictionem eorum et virum Aegyptium percutientem quendam de Hebraeis fratribus suis.
EXOD|2|12|Cumque circumspexisset huc atque illuc et nullum adesse vidisset, percussum Aegyptium abscondit sabulo.
EXOD|2|13|Et egressus die altero conspexit duos Hebraeos rixantes dixitque ei, qui faciebat iniuriam: " Quare percutis proximum tuum? ".
EXOD|2|14|Qui respondit: " Quis te constituit principem et iudicem super nos? Num occidere me tu vis, sicut occidisti Aegyptium? ". Timuit Moyses et ait: " Quomodo palam factum est verbum istud? ".
EXOD|2|15|Audivitque pharao sermonem hunc et quaerebat occidere Moysen. Qui fugiens de conspectu eius moratus est in terra Madian; venit ergo in terram Madian et sedit iuxta puteum.
EXOD|2|16|Erant autem sacerdoti Madian septem filiae, quae venerunt ad hauriendam aquam; et impletis canalibus adaquare cupiebant greges patris sui.
EXOD|2|17|Supervenere pastores et eiecerunt eas: surrexitque Moyses et, defensis puellis, adaquavit oves earum.
EXOD|2|18|Quae cum revertissent ad Raguel patrem suum, dixit ad eas: " Cur velocius venistis solito? ".
EXOD|2|19|Responderunt: " Vir Aegyptius liberavit nos de manu pastorum; insuper et hausit aquam nobis potumque dedit ovibus ".
EXOD|2|20|At ille: " Ubi est? ", inquit. " Quare dimisistis hominem? Vocate eum, ut comedat panem ".
EXOD|2|21|Consensit ergo Moyses habitare cum eo accepitque Sephoram filiam eius uxorem.
EXOD|2|22|Quae peperit ei filium, quem vocavit Gersam dicens: " Advena sum in terra aliena ".
EXOD|2|23|Post multum vero temporis mortuus est rex Aegypti; et ingemiscentes filii Israel propter opera vociferati sunt, ascenditque clamor eorum ad Deum ab operibus.
EXOD|2|24|Et audivit gemitum eorum ac recordatus est foederis, quod pepigit cum Abraham, Isaac et Iacob;
EXOD|2|25|et respexit Dominus filios Israel et apparuit eis.
EXOD|3|1|Moyses autem pascebat oves Iethro soceri sui sacerdotis Ma dian; cumque minasset gregem ultra desertum, venit ad montem Dei Horeb.
EXOD|3|2|Apparuitque ei angelus Domini in flamma ignis de medio rubi; et videbat quod rubus arderet et non combureretur.
EXOD|3|3|Dixit ergo Moyses: " Vadam et videbo visionem hanc magnam, quare non comburatur rubus ".
EXOD|3|4|Cernens autem Dominus quod pergeret ad videndum, vocavit eum Deus de medio rubi et ait: " Moyses, Moyses ". Qui respondit: " Adsum ".
EXOD|3|5|At ille: " Ne appropies, inquit, huc; solve calceamentum de pedibus tuis; locus enim, in quo stas, terra sancta est ".
EXOD|3|6|Et ait: " Ego sum Deus patris tui, Deus Abraham, Deus Isaac et Deus Iacob ". Abscondit Moyses faciem suam; non enim audebat aspicere contra Deum.
EXOD|3|7|Cui ait Dominus: " Vidi afflictionem populi mei in Aegypto et clamorem eius audivi propter duritiam exactorum eorum.
EXOD|3|8|Et sciens dolorem eius descendi, ut liberem eum de manibus Aegyptiorum et educam de terra illa in terram bonam et spatiosam, in terram, quae fluit lacte et melle, ad loca Chananaei et Hetthaei et Amorraei et Pherezaei et Hevaei et Iebusaei.
EXOD|3|9|Clamor ergo filiorum Israel venit ad me, vidique afflictionem eorum, qua ab Aegyptiis opprimuntur;
EXOD|3|10|sed veni, mittam te ad pharaonem, ut educas populum meum, filios Israel, de Aegypto ".
EXOD|3|11|Dixitque Moyses ad Deum: " Quis sum ego, ut vadam ad pharaonem et educam filios Israel de Aegypto? ".
EXOD|3|12|Qui dixit ei: " Ego ero tecum; et hoc habebis signum quod miserim te: cum eduxeris populum de Aegypto, servietis Deo super montem istum ".
EXOD|3|13|Ait Moyses ad Deum: " Ecce, ego vadam ad filios Israel et dicam eis: Deus patrum vestrorum misit me ad vos. Si dixerint mihi: "Quod est nomen eius?" quid dicam eis? ".
EXOD|3|14|Dixit Deus ad Moysen: " Ego sum qui sum ". Ait: " Sic dices filiis Israel: Qui sum misit me ad vos ".
EXOD|3|15|Dixitque iterum Deus ad Moysen: " Haec dices filiis Israel: Dominus, Deus patrum vestrorum, Deus Abraham, Deus Isaac et Deus lacob, misit me ad vos; hoc nomen mihi est in aeternum, et hoc memoriale meum in generationem et generationem.
EXOD|3|16|Vade et congrega seniores Israel et dices ad eos: Dominus, Deus patrum vestrorum, apparuit mihi, Deus Abraham, Deus Isaac et Deus Iacob, dicens: Visitans visitavi vos et vidi omnia, quae acciderunt vobis in Aegypto;
EXOD|3|17|et dixi: Educam vos de afflictione Aegypti in terram Chananaei et Hetthaei et Amorraei et Pherezaei et Hevaei et Iebusaei, ad terram fluentem lacte et melle.
EXOD|3|18|Et audient vocem tuam; ingredierisque tu et seniores Israel ad regem Aegypti, et dicetis ad eum: Dominus, Deus Hebraeorum, occurrit nobis; et nunc eamus viam trium dierum in solitudinem, ut immolemus Domino Deo nostro.
EXOD|3|19|Sed ego scio quod non dimittet vos rex Aegypti, ut eatis, nisi per manum validam.
EXOD|3|20|Extendam enim manum meam et percutiam Aegyptum in cunctis mirabilibus meis, quae facturus sum in medio eius; post haec dimittet vos.
EXOD|3|21|Daboque gratiam populo huic coram Aegyptiis, et, cum egrediemini, non exibitis vacui.
EXOD|3|22|Sed postulabit mulier a vicina sua et ab hospita sua vasa argentea et aurea ac vestes; ponetisque eas super filios et filias vestras et spoliabitis Aegyptum ".
EXOD|4|1|Respondens Moyses ait: " Quid autem, si non credent mihi ne que audient vocem meam, sed dicent: "Non apparuit tibi Dominus?" ".
EXOD|4|2|Dixit ergo ad eum: " Quid est quod tenes in manu tua? ". Respondit: " Virga ".
EXOD|4|3|Dixitque Dominus: " Proice eam in terram! ". Proiecit, et versa est in serpentem, ita ut fugeret Moyses.
EXOD|4|4|Dixitque Dominus: " Extende manum tuam et apprehende caudam eius! ". Extendit et tenuit, versaque est in virgam.
EXOD|4|5|" Ut credant, inquit, quod apparuerit tibi Dominus, Deus patrum suorum, Deus Abraham, Deus Isaac et Deus Iacob ".
EXOD|4|6|Dixitque Dominus rursum: " Mitte manum tuam in sinum tuum! ". Quam cum misisset in sinum, protulit leprosam instar nivis.
EXOD|4|7|" Retrahe, ait, manum tuam in sinum tuum! ". Retraxit et protulit iterum, et erat similis carni reliquae.
EXOD|4|8|" Si non crediderint, inquit, tibi, neque audierint sermonem signi prioris, credent verbo signi sequentis.
EXOD|4|9|Quod si nec duobus quidem his signis crediderint neque audierint vocem tuam, sume aquam fluminis et effunde eam super aridam, et, quidquid hauseris de fluvio, vertetur in sanguinem ".
EXOD|4|10|Ait Moyses: " Obsecro, Domine, non sum eloquens ab heri et nudiustertius et ex quo locutus es ad servum tuum, nam impeditioris et tardioris linguae sum ".
EXOD|4|11|Dixit Dominus ad eum: " Quis fecit os hominis? Aut quis fabricatus est mutum vel surdum vel videntem vel caecum? Nonne ego?
EXOD|4|12|Perge igitur, et ego ero in ore tuo; doceboque te quid loquaris ".
EXOD|4|13|At ille: " Obsecro, inquit, Domine, mitte quem missurus es ".
EXOD|4|14|Iratus Dominus in Moysen ait: " Aaron, frater tuus Levites, scio quod eloquens sit; ecce ipse egreditur in occursum tuum vidensque te laetabitur corde.
EXOD|4|15|Loquere ad eum et pone verba mea in ore eius; et ego ero in ore tuo et in ore illius et ostendam vobis quid agere debeatis.
EXOD|4|16|Ipse loquetur pro te ad populum et erit os tuum; tu autem eris ei ut Deus.
EXOD|4|17|Virgam quoque hanc sume in manu tua, in qua facturus es signa ".
EXOD|4|18|Abiit Moyses et reversus est ad Iethro socerum suum dixitque ei: " Vadam, quaeso, et revertar ad fratres meos in Aegyptum, ut videam, si adhuc vivant ". Cui ait Iethro: " Vade in pace ".
EXOD|4|19|Dixit ergo Dominus ad Moysen in Madian: " Vade, revertere in Aegyptum; mortui sunt enim omnes, qui quaerebant animam tuam ".
EXOD|4|20|Tulit Moyses uxorem suam et filios suos et imposuit eos super asinum; reversusque est in Aegyptum portans virgam Dei in manu sua.
EXOD|4|21|Dixitque ei Dominus revertenti in Aegyptum: " Vide, ut omnia ostenta, quae posui in manu tua, facias coram pharaone; ego indurabo cor eius, et non dimittet populum.
EXOD|4|22|Dicesque ad eum: Haec dicit Dominus: Filius meus primogenitus Israel.
EXOD|4|23|Dico tibi: Dimitte filium meum, ut serviat mihi; si autem non vis dimittere eum, ecce ego interficiam filium tuum primogenitum ".
EXOD|4|24|Cumque esset in itinere, in deversorio, occurrit ei Dominus et volebat occidere eum.
EXOD|4|25|Tulit ilico Sephora acutissimam petram et circumcidit praeputium filii sui; tetigitque pedes eius et ait: " Sponsus sanguinum tu mihi es ".
EXOD|4|26|Et dimisit eum, postquam dixerat: " Sponsus sanguinum ", ob circumcisionem.
EXOD|4|27|Dixit autem Dominus ad Aaron: " Vade in occursum Moysi in desertum ". Qui perrexit obviam ei in montem Dei et osculatus est eum.
EXOD|4|28|Narravitque Moyses Aaron omnia verba Domini, quibus miserat eum, et signa, quae mandaverat.
EXOD|4|29|Veneruntque simul et congregaverunt cunctos seniores filiorum Israel.
EXOD|4|30|Locutusque est Aaron omnia verba, quae dixerat Dominus ad Moysen, et fecit signa coram populo.
EXOD|4|31|Et credidit populus, audieruntque quod visitasset Dominus filios Israel et quod respexisset afflictionem eorum; et proni adoraverunt.
EXOD|5|1|Post haec ingressi sunt Moyses et Aaron et dixerunt pharaoni: " Haec dicit Dominus, Deus Israel: Dimitte populum meum, ut sacrificet mihi in deserto ".
EXOD|5|2|At ille responclit: " Quis est Dominus, ut audiam vocem eius et dimittam Israel? Nescio Dominum et Israel non dimittam ".
EXOD|5|3|Dixeruntque: " Deus Hebraeorum occurrit nobis; eamus, quaeso, viam trium dierum in solitudinem et sacrificemus Domino Deo nostro, ne forte accidat nobis pestis aut gladius ".
EXOD|5|4|Ait ad eos rex Aegypti: " Quare, Moyses et Aaron, sollicitatis populum ab operibus suis? Ite ad onera vestra ".
EXOD|5|5|Dixitque pharao: " Multus nimis iam est populus terrae; videtis quod turba succreverit; quanto magis si dederitis eis requiem ab operibus? ".
EXOD|5|6|Praecepit ergo in die illo exactoribus populi et praefectis eius dicens:
EXOD|5|7|" Nequaquam ultra dabitis paleas populo ad conficiendos lateres sicut prius, sed ipsi vadant et colligant stipulas.
EXOD|5|8|Et mensuram laterum, quam prius faciebant, imponetis super eos; nec minuetis quidquam. Vacant enim et idcirco vociferantur dicentes: "Eamus et sacrificemus Deo nostro".
EXOD|5|9|Opprimantur operibus et expleant ea, ut non acquiescant verbis mendacibus ".
EXOD|5|10|Igitur egressi exactores populi et praefecti eius dixerunt ad populum: " Sic dicit pharao: "Non do vobis paleas.
EXOD|5|11|Ite et colligite, sicubi invenire poteritis, nec minuetur quid quam de opere vestro" ".
EXOD|5|12|Dispersusque est populus per omnem terram Aegypti ad colligendas paleas.
EXOD|5|13|Exactores quoque instabant dicentes: " Complete opus vestrum cotidie, ut prius facere solebatis, quando dabantur vobis paleae ".
EXOD|5|14|Flagellatique sunt praefecti filiorum Israel, quos constituerant super eos exactores pharaonis dicentes: " Quare non implestis mensuram laterum sicut prius, nec heri nec hodie? ".
EXOD|5|15|Veneruntque praefecti filiorum Israel et vociferati sunt ad pharaonem dicentes: " Cur ita agis contra servos tuos?
EXOD|5|16|Paleae non dantur nobis, et lateres similiter imperantur; en famuli tui flagellis caedimur, et populus tuus est in culpa ".
EXOD|5|17|Qui ait: " Vacatis otio et idcirco dicitis: "Eamus et sacrificemus Domino".
EXOD|5|18|Ite ergo et operamini; paleae non dabuntur vobis, et reddetis consuetum numerum laterum ".
EXOD|5|19|Videbantque se praefecti filiorum Israel in malo, eo quod diceretur eis: " Non minuetur quidquam de lateribus per singulos dies ";
EXOD|5|20|occurreruntque Moysi et Aaron, qui stabant ex adverso egredientibus a pharaone,
EXOD|5|21|et dixerunt ad eos: " Videat Dominus et iudicet, quoniam foetere fecistis odorem nostrum coram pharaone et servis eius; et praebuistis ei gladium, ut occideret nos ".
EXOD|5|22|Reversusque est Moyses ad Dominum et ait: " Domine, cur afflixisti populum istum? Quare misisti me?
EXOD|5|23|Ex eo enim quo ingressus sum ad pharaonem, ut loquerer in nomine tuo, afflixit populum tuum; et non liberasti eos ".
EXOD|6|1|Dixitque Dominus ad Moysen: " Nunc videbis quae facturus sim pharaoni; per manum enim fortem dimittet eos et in manu robusta eiciet illos de terra sua ".
EXOD|6|2|Locutusque est Dominus ad Moysen dicens: " Ego Dominus,
EXOD|6|3|qui apparui Abraham, Isaac et Iacob ut Deus omnipotens; et nomen meum Dominum non indicavi eis.
EXOD|6|4|Pepigique cum eis foedus, ut darem illis terram Chanaan, terram peregrinationis eorum, in qua fuerunt advenae.
EXOD|6|5|Ego audivi gemitum filiorum Israel, quia Aegyptii oppresserunt eos, et recordatus sum pacti mei.
EXOD|6|6|Ideo dic filiis Israel: Ego Dominus, qui educam vos de ergastulo Aegyptiorum; et eruam de servitute ac redimam in brachio excelso et iudiciis magnis.
EXOD|6|7|Et assumam vos mihi in populum et ero vester Deus; et scietis quod ego sum Dominus Deus vester, qui eduxerim vos de ergastulo Aegyptiorum
EXOD|6|8|et induxerim in terram, super quam levavi manum meam, ut darem eam Abraham, Isaac et Iacob; daboque illam vobis possidendam, ego Dominus ".
EXOD|6|9|Narravit ergo Moyses omnia filiis Israel; qui non acquieverunt ei propter angustiam spiritus et opus durissimum.
EXOD|6|10|Locutusque est Dominus ad Moysen dicens:
EXOD|6|11|" Ingredere et loquere ad pharaonem regem Aegypti, ut dimittat filios Israel de terra sua ".
EXOD|6|12|Respondit Moyses coram Domino: " Ecce, filii Israel non audiunt me, et quomodo audiet me pharao, praesertim cum incircumcisus sim labiis? ".
EXOD|6|13|Locutusque est Dominus ad Moysen et Aaron et dedit mandatum ad filios Israel et ad pharaonem regem Aegypti, ut educerent filios Israel de terra Aegypti.
EXOD|6|14|Isti sunt principes domorum per familias suas.Filii Ruben primogeniti Israelis: Henoch et Phallu, Hesron et Charmi; hae cognationes Ruben.
EXOD|6|15|Filii Simeon: Iamuel et Iamin et Ahod et Iachin et Sohar er Saul filius Chananitidis; hae progenies Simeon.
EXOD|6|16|Et haec nomina filiorum Levi per cognationes suas: Gerson et Caath et Merari; anni autem vitae Levi fuerunt centum triginta septem.
EXOD|6|17|Filii Gerson: Lobni et Semei per cognationes suas.
EXOD|6|18|Filii Caath: Amram et Isaar et Hebron et Oziel; anni quoque vitae Caath centum triginta tres.
EXOD|6|19|Filii Merari: Moholi et Musi; hae cognationes Levi per familias suas.
EXOD|6|20|Accepit autem Amram uxorem Iochabed amitam suam, quae peperit ei Aaron et Moysen; fueruntque anni vitae Amram centum triginta septem.
EXOD|6|21|Filii quoque Isaar: Core et Napheg et Zechri.
EXOD|6|22|Filii quoque Oziel: Misael et Elisaphan et Sethri.
EXOD|6|23|Accepit autem Aaron uxorem Elisabeth filiam Aminadab sororem Naasson, quae peperit ei Nadab et Abiu et Eleazar et Ithamar.
EXOD|6|24|Filii quoque Core: Asir et Elcana et Abiasaph; hae sunt cognationes Coritarum.
EXOD|6|25|At vero Eleazar filius Aaron accepit uxorem de filiabus Phutiel, quae peperit ei Phinees; hi sunt principes familiarum Leviticarum per cognationes suas.
EXOD|6|26|Iste est Aaron et Moyses, quibus praecepit Dominus, ut educerent filios Israel de terra Aegypti per turmas suas.
EXOD|6|27|Hi sunt qui loquuntur ad pharaonem regem Aegypti, ut educant filios Israel de Aegypto; iste est Moyses et Aaron
EXOD|6|28|in die, qua locutus est Dominus ad Moysen in terra Aegypti.
EXOD|6|29|Et locutus est Dominus ad Moysen dicens: " Ego Dominus; loquere ad pharaonem regem Aegypti omnia, quae ego loquor tibi ".
EXOD|6|30|Et ait Moyses coram Domino: " En incircumcisus labiis sum. Quomodo audiet me pharao? ".
EXOD|7|1|Dixitque Dominus ad Moysen: " Ecce constitui te deum pha raonis, et Aaron frater tuus erit propheta tuus.
EXOD|7|2|Tu loqueris omnia, quae mando tibi; et ille loquetur ad pharaonem, ut dimittat filios Israel de terra sua.
EXOD|7|3|Sed ego indurabo cor eius et multiplicabo signa et ostenta mea in terra Aegypti.
EXOD|7|4|Et non audiet vos; immittamque manum meam super Aegyptum et educam exercitum et populum meum, filios Israel, de terra Aegypti per iudicia maxima.
EXOD|7|5|Et scient Aegyptii quia ego sum Dominus, qui extenderim manum meam super Aegyptum et eduxerim filios Israel de medio eorum ".
EXOD|7|6|Fecit itaque Moyses et Aaron, sicut praeceperat Dominus; ita egerunt.
EXOD|7|7|Erat autem Moyses octoginta annorum, et Aaron octoginta trium, quando locuti sunt ad pharaonem.
EXOD|7|8|Dixitque Dominus ad Moysen et Aaron:
EXOD|7|9|" Cum dixerit vobis pharao: "Ostendite signum", dices ad Aaron: Tolle virgam tuam et proice eam coram pharaone, ac vertetur in colubrum ".
EXOD|7|10|Ingressi itaque Moyses et Aaron ad pharaonem fecerunt, sicut praeceperat Dominus; proiecitque Aaron virgam coram pharaone et servis eius, quae versa est in colubrum.
EXOD|7|11|Vocavit autem pharao sapientes et maleficos, et fecerunt etiam ipsi magi Aegypti per incantationes suas similiter.
EXOD|7|12|Proieceruntque singuli virgas suas, quae versae sunt in colubros; sed devoravit virga Aaron virgas eorum.
EXOD|7|13|Induratumque est cor pharaonis, et non audivit eos, sicut dixerat Dominus.
EXOD|7|14|Dixit autem Dominus ad Moysen: " Ingravatum est cor pharaonis: non vult dimittere populum.
EXOD|7|15|Vade ad eum mane. Ecce egredietur ad aquas; et stabis in occursum eius super ripam fluminis. Et virgam, quae conversa est in serpentem, tolles in manu tua
EXOD|7|16|dicesque ad eum: Dominus, Deus Hebraeorum, misit me ad te dicens: Dimitte populum meum, ut sacrificet mihi in deserto; et usque ad praesens audire noluisti.
EXOD|7|17|Haec igitur dicit Dominus: In hoc scies quod sim Dominus: ecce percutiam virga, quae in manu mea est, aquam fluminis; et vertetur in sanguinem.
EXOD|7|18|Pisces quoque, qui sunt in fluvio, morientur, et computrescent aquae, et taedebit Aegyptios bibere aquam fluminis ".
EXOD|7|19|Dixit quoque Dominus ad Moysen: " Dic ad Aaron: Tolle virgam tuam et extende manum tuam super aquas Aegypti, super fluvios eorum et rivos ac paludes et omnes lacus aquarum, ut vertantur in sanguinem; et sit cruor in omni terra Aegypti, tam in ligneis vasis quam in saxeis ".
EXOD|7|20|Feceruntque ita Moyses et Aaron, sicut praeceperat Dominus. Et elevans virgam percussit aquam fluminis coram pharaone et servis eius; quae versa est in sanguinem.
EXOD|7|21|Et pisces, qui erant in flumine, mortui sunt, computruitque fluvius, et non poterant Aegyptii bibere aquam fluminis; et fuit sanguis in tota terra Aegypti.
EXOD|7|22|Feceruntque similiter malefici Aegyptiorum incantationibus suis; et induratum est cor pharaonis, nec audivit eos, sicut dixerat Dominus.
EXOD|7|23|Avertitque se et ingressus est domum suam nec ad hoc apposuit cor suum.
EXOD|7|24|Foderunt autem omnes Aegyptii per circuitum fluminis aquam, ut biberent; non enim poterant bibere de aqua fluminis.
EXOD|7|25|Impletique sunt septem dies, postquam percussit Dominus fluvium.
EXOD|7|26|Dixit quoque Dominus ad Moysen: " Ingredere ad pharaonem et dices ad eum: Haec dicit Dominus: Dimitte populum meum, ut sacrificet mihi.
EXOD|7|27|Sin autem nolueris dimittere, ecce ego percutiam omnes terminos tuos ranis.
EXOD|7|28|Et ebulliet fluvius ranas, quae ascendent et ingredientur domum tuam et cubiculum lectuli tui et super stratum tuum et in domos servorum tuorum et in populum tuum et in furnos tuos et in pistrina tua;
EXOD|7|29|et ad te et ad populum tuum et ad omnes servos tuos intrabunt ranae ".
EXOD|8|1|Dixitque Dominus ad Moysen: " Dic ad Aaron: Extende ma num tuam cum baculo tuo super fluvios, super rivos ac paludes et educ ranas super terram Aegypti ".
EXOD|8|2|Et extendit Aaron manum super aquas Aegypti, et ascenderunt ranae operueruntque terram Aegypti.
EXOD|8|3|Fecerunt autem et malefici per incantationes suas similiter eduxeruntque ranas super terram Aegypti.
EXOD|8|4|Vocavit autem pharao Moysen et Aaron et dixit: " Orate Dominum, ut auferat ranas a me et a populo meo, et dimittam populum, ut sacrificet Domino ".
EXOD|8|5|Dixitque Moyses ad pharaonem: " Constitue mihi, quando deprecer pro te et pro servis et pro populo tuo, ut abigantur ranae a te et a domo tua et tantum in flumine remaneant ".
EXOD|8|6|Qui respondit: " Cras ". At ille: " Iuxta verbum, inquit, tuum faciam, ut scias quoniam non est sicut Dominus Deus noster.
EXOD|8|7|Et recedent ranae a te et a domo tua et a servis tuis et a populo tuo; tantum in flumine remanebunt ".
EXOD|8|8|Egressique sunt Moyses et Aaron a pharaone; et clamavit Moyses ad Dominum pro sponsione ranarum, quam condixerat pharaoni.
EXOD|8|9|Fecitque Dominus iuxta verbum Moysi, et mortuae sunt ranae de domibus et de villis et de agris;
EXOD|8|10|congregaveruntque eas in immensos aggeres, et computruit terra.
EXOD|8|11|Videns autem pharao quod data esset requies, ingravavit cor suum et non audivit eos, sicut dixerat Dominus.
EXOD|8|12|Dixitque Dominus ad Moysen: " Loquere ad Aaron: Extende virgam tuam et percute pulverem terrae, et sint scinifes in universa terra Aegypti ".
EXOD|8|13|Feceruntque ita; et extendit Aaron manum virgam tenens percussitque pulverem terrae. Et facti sunt scinifes in hominibus et in iumentis; omnis pulvis terrae versus est in scinifes per totam terram Aegypti.
EXOD|8|14|Feceruntque similiter malefici incantationibus suis, ut educerent scinifes; et non potuerunt. Erantque scinifes tam in hominibus quam in iumentis;
EXOD|8|15|et dixerunt malefici ad pharaonem: " Digitus Dei est hic ". Induratumque est cor pharaonis et non audivit eos, sicut praeceperat Dominus.
EXOD|8|16|Dixit quoque Dominus ad Moysen: " Consurge diluculo et sta coram pharaone. Egredietur enim ad aquas, et dices ad eum: Haec dicit Dominus: Dimitte populum meum, ut sacrificet mihi.
EXOD|8|17|Quod si non dimiseris eum, ecce ego immittam in te et in servos tuos et in populum tuum et in domos tuas omne genus muscarum; et implebuntur domus Aegyptiorum muscis et etiam humus, in qua fuerint.
EXOD|8|18|Et segregabo in die illa terram Gessen, in qua populus meus est, ut non sint ibi muscae, et scias quoniam ego Dominus in medio terrae;
EXOD|8|19|ponamque divi sionem inter populum meum et populum tuum; cras erit signum istud ".
EXOD|8|20|Fecitque Dominus ita; et venit musca gravissima in domos pharaonis et servorum eius et in omnem terram Aegypti, corruptaque est terra ab huiuscemodi muscis.
EXOD|8|21|Vocavitque pharao Moysen et Aaron et ait eis: " Ite, sacrificate Deo vestro in terra ".
EXOD|8|22|Et ait Moyses: " Non potest ita fieri: abominationes enim Aegyptiorum immolabimus Domino Deo nostro; quod si mactaverimus ea, quae colunt Aegyptii, coram eis, lapidibus nos obruent.
EXOD|8|23|Viam trium dierum pergemus in solitudinem et sacrificabimus Domino Deo nostro, sicut praecepit nobis ".
EXOD|8|24|Dixitque pharao: " Ego dimittam vos, ut sacrificetis Domino Deo vestro in deserto, verumtamen longius ne abeatis; rogate pro me ".
EXOD|8|25|Et ait Moyses: " Egressus a te, orabo Dominum, et recedet musca a pharaone et a servis suis et a populo eius cras; verumtamen noli ultra fallere, ut non dimittas populum sacrificare Domino ".
EXOD|8|26|Egressusque Moyses a pharaone oravit Dominum;
EXOD|8|27|qui fecit iuxta verbum illius et abstulit muscas a pharaone et a servis suis et a populo eius; non superfuit ne una quidem.
EXOD|8|28|Et ingravatum est cor pharaonis, ita ut ne hac quidem vice dimitteret populum.
EXOD|9|1|Dixit autem Dominus ad Moysen: " Ingredere ad pharaonem et loquere ad eum: Haec dicit Dominus, Deus Hebraeorum: Dimitte populum meum, ut sacrificet mihi.
EXOD|9|2|Quod si adhuc renuis et retines eos,
EXOD|9|3|ecce manus Domini erit super possessionem tuam in agris, super equos et asinos et camelos et boves et oves, pestis valde gravis;
EXOD|9|4|et distinguet Dominus inter possessiones Israel et possessiones Aegyptiorum, ut nihil omnino pereat ex his, quae pertinent ad filios Israel.
EXOD|9|5|Constituitque Dominus tempus dicens: Cras faciet Dominus verbum istud in terra ".
EXOD|9|6|Fecit ergo Dominus verbum hoc altera die, mortuaque sunt omnia animantia Aegyptiorum; de animalibus vero filiorum Israel nihil omnino periit.
EXOD|9|7|Et misit pharao ad videndum; nec erat quidquam mortuum de his, quae possidebat Israel. Ingravatumque est cor pharaonis, et non dimisit populum.
EXOD|9|8|Et dixit Dominus ad Moysen et Aaron: " Tollite plenas manus cineris de camino, et spargat illum Moyses in caelum coram pharaone;
EXOD|9|9|sitque pulvis super omnem terram Aegypti; erunt enim in hominibus et iumentis ulcera et vesicae turgentes in universa terra Aegypti ".
EXOD|9|10|Tuleruntque cinerem de camino et steterunt coram pharaone, et sparsit illum Moyses in caelum; factaque sunt ulcera vesicarum turgentium in hominibus et iumentis.
EXOD|9|11|Nec poterant malefici stare coram Moyse propter ulcera, quae in illis erant et in omni terra Aegypti.
EXOD|9|12|Induravitque Dominus cor pharaonis, et non audivit eos, sicut locutus est Dominus ad Moysen.
EXOD|9|13|Dixitque Dominus ad Moysen: " Mane consurge et sta coram pharaone et dices ad eum: Haec dicit Dominus, Deus Hebraeorum: Dimitte populum meum, ut sacrificet mihi;
EXOD|9|14|quia in hac vice mittam omnes plagas meas super cor tuum et super servos tuos et super populum tuum, ut scias quod non sit similis mei in omni terra.
EXOD|9|15|Nunc enim extendens manum si percussissem te et populum tuum peste, perisses de terra.
EXOD|9|16|Idcirco autem servavi te, ut ostendam in te fortitudinem meam, et narretur nomen meum in omni terra.
EXOD|9|17|Adhuc retines populum meum et non vis dimittere eum?
EXOD|9|18|En pluam cras, hac ipsa hora, grandinem multam nimis, qualis non fuit in Aegypto a die, qua fundata est, usque in praesens tempus.
EXOD|9|19|Mitte ergo iam nunc et congrega iumenta tua et omnia, quae habes in agro; homines enim et iumenta universa, quae inventa fuerint foris nec congregata de agris, cadet super ea grando, et morientur ".
EXOD|9|20|Qui timuit verbum Domini de servis pharaonis, fecit confugere servos suos et iumenta in domos;
EXOD|9|21|qui autem neglexit sermonem Domini, dimisit servos suos et iumenta in agris.
EXOD|9|22|Et dixit Dominus ad Moysen: " Extende manum tuam in caelum, ut fiat grando in universa terra Aegypti super homines et super iumenta et super omnem herbam agri in terra Aegypti ".
EXOD|9|23|Extenditque Moyses virgam in caelum, et Dominus dedit tonitrua et grandinem ac discurrentia fulgura super terram; pluitque Dominus grandinem super terram Aegypti.
EXOD|9|24|Et grando et ignis immixta pariter ferebantur; tantaeque fuit magnitudinis, quanta ante numquam apparuit in universa terra Aegypti, ex quo gens illa condita est.
EXOD|9|25|Et percussit grando in omni terra Aegypti cuncta, quae fuerunt in agris, ab homine usque ad iumentum; cunctamque herbam agri percussit grando et omne lignum regionis confregit.
EXOD|9|26|Tantum in terra Gessen, ubi erant filii Israel, grando non cecidit.
EXOD|9|27|Misitque pharao et vocavit Moysen et Aaron dicens ad eos: " Nunc peccavi; Dominus iustus, ego et populus meus rei.
EXOD|9|28|Orate Dominum, ut desinant tonitrua Dei et grando, et dimittam vos, et nequaquam hic ultra manebitis ".
EXOD|9|29|Ait Moyses: " Cum egressus fuero de urbe, extendam palmas meas ad Dominum; et cessabunt tonitrua, et grando non erit, ut scias quia Domini est terra.
EXOD|9|30|Novi autem quod et tu et servi tui necdum timeatis Dominum Deum ".
EXOD|9|31|Linum ergo et hordeum laesum est, eo quod hordeum iam spicas et linum iam folliculos germinaret;
EXOD|9|32|triticum autem et far non sunt laesa, quia serotina erant.
EXOD|9|33|Egressusque Moyses a pharaone ex urbe tetendit manus ad Dominum; et cessaverunt tonitrua et grando, nec ultra effundebatur pluvia super terram. 34 Videns autem pharao quod cessasset pluvia et grando et tonitrua, auxit peccatum; 35 et ingravatum est cor eius et servorum illius et induratum nimis; nec dimisit filios Israel, sicut dixerat Dominus per manum Moysi.
EXOD|10|1|Et dixit Dominus ad Moy sen: " Ingredere ad pharao nem: ego enim induravi cor eius et servorum illius, ut faciam signa mea haec in medio eorum,
EXOD|10|2|et narres in auribus filii tui et nepotum tuorum, quotiens contriverim Aegyptios et signa mea fecerim in eis; et sciatis quia ego Dominus ".
EXOD|10|3|Introierunt ergo Moyses et Aaron ad pharaonem et dixerunt ei: " Haec dicit Dominus, Deus Hebraeorum: Usquequo non vis subici mihi? Dimitte populum meum, ut sacrificet mihi.
EXOD|10|4|Sin autem resistis et non vis dimittere eum, ecce ego inducam cras locustam in fines tuos,
EXOD|10|5|quae operiat superficiem terrae, ne quidquam eius appareat, sed comedatur, quod residuum fuerit grandini; corrodet enim omnia ligna, quae germinant in agris.
EXOD|10|6|Et implebunt domos tuas et servorum tuorum et omnium Aegyptiorum, quantam non viderunt patres tui et avi, ex quo orti sunt super terram usque in praesentem diem ". Avertitque se et egressus est a pharaone.
EXOD|10|7|Dixerunt autem servi pharaonis ad eum: " Usquequo patiemur hoc scandalum? Dimitte homines, ut sacrificent Domino Deo suo; nonne vides quod perierit Aegyptus? ".
EXOD|10|8|Revocaveruntque Moysen et Aaron ad pharaonem, qui dixit eis: " Ite, sacrificate Domino Deo vestro. Quinam sunt qui ituri sunt? ".
EXOD|10|9|Ait Moyses: " Cum parvulis nostris et senioribus pergemus, cum filiis et filiabus, cum ovibus et armentis; est enim sollemnitas Domini nobis ".
EXOD|10|10|Et respondit eis: " Sic Dominus sit vobiscum, quomodo ego dimittam vos et parvulos vestros. Cui dubium est quod pessime cogitetis?
EXOD|10|11|Non fiet ita, sed ite tantum viri et sacrificate Domino; hoc enim et ipsi petistis ". Statimque eiecti sunt de conspectu pharaonis.
EXOD|10|12|Dixit autem Dominus ad Moysen: " Extende manum tuam super terram Aegypti, ut veniat locusta et ascendat super eam et devoret omnem herbam, quidquid residuum fuerit grandini ".
EXOD|10|13|Et extendit Moyses virgam super terram Aegypti, et Dominus induxit ventum urentem tota die illa et nocte. Et mane facto, ventus urens levavit locustas;
EXOD|10|14|quae ascenderunt super universam terram Aegypti et sederunt in cunctis finibus Aegyptiorum innumerabiles, quales ante illud tempus non fuerant nec postea futurae sunt.
EXOD|10|15|Operueruntque universam superficiem terrae, et obscurata est terra. Devoraverunt igitur omnem herbam terrae et, quidquid pomorum in arboribus fuit, quae grando dimiserat; nihilque omnino virens relictum est in lignis et in herbis terrae in cuncta Aegypto.
EXOD|10|16|Quam ob rem festinus pharao vocavit Moysen et Aaron et dixit eis: " Peccavi in Dominum Deum vestrum et in vos.
EXOD|10|17|Sed nunc dimittite peccatum mihi tantum hac vice et rogate Dominum Deum vestrum, ut auferat a me saltem mortem istam ".
EXOD|10|18|Egressusque Moyses de conspectu pharaonis oravit Dominum,
EXOD|10|19|qui flare fecit ventum ab occidente vehementissimum et arreptam locustam proiecit in mare Rubrum; non remansit ne una quidem in cunctis finibus Aegypti.
EXOD|10|20|Et induravit Dominus cor pharaonis, nec dimisit filios Israel.
EXOD|10|21|Dixit autem Dominus ad Moysen: " Extende manum tuam in caelum, et sint tenebrae super terram Aegypti tam densae ut palpari queant ".
EXOD|10|22|Extenditque Moyses manum in caelum, et factae sunt tenebrae horribiles in universa terra Aegypti tribus diebus.
EXOD|10|23|Nemo vidit fratrem suum nec movit se de loco, in quo erat. Ubicumque autem habitabant filii Israel, lux erat.
EXOD|10|24|Vocavitque pharao Moysen et Aaron et dixit eis: " Ite, sacrificate Domino; oves tantum vestrae et armenta remaneant, parvuli vestri eant vobiscum ".
EXOD|10|25|Ait Moyses: " Etiamsi tu hostias et holocausta dares nobis, quae offeramus Domino Deo nostro,
EXOD|10|26|tamen et greges nostri pergent nobiscum; non remanebit ex eis ungula, quoniam ex ipsis sumemus, quae necessaria sunt in cultum Domini Dei nostri; praesertim cum ignoremus quid debeat immolari, donec ad ipsum locum perveniamus ".
EXOD|10|27|Induravit autem Dominus cor pharaonis, et noluit dimittere eos.
EXOD|10|28|Dixitque pharao ad eum: " Recede a me. Cave, ne ultra videas faciem meam; quocumque die apparueris mihi, morieris ".
EXOD|10|29|Respondit Moyses: " Ita fiet, ut locutus es; non videbo ultra faciem tuam ".
EXOD|11|1|Et dixit Dominus ad Moy sen: " Adhuc una plaga tan gam pharaonem et Aegyptum, et post haec dimittet vos utique, immo et exire compellet.
EXOD|11|2|Dices ergo omni plebi, ut postulet vir ab amico suo et mulier a vicina sua vasa argentea et aurea;
EXOD|11|3|dabit autem Dominus gratiam populo coram Aegyptiis ". Fuitque Moyses vir magnus valde in terra Aegypti coram servis pharaonis et omni populo.
EXOD|11|4|Et ait Moyses: " Haec dicit Dominus: Media nocte egrediar in Aegyptum;
EXOD|11|5|et morietur omne primogenitum in terra Aegyptiorum, a primogenito pharaonis, qui sedet in solio eius, usque ad primogenitum ancillae, quae est ad molam, et omnia primogenita iumentorum.
EXOD|11|6|Eritque clamor magnus in universa terra Aegypti, qualis nec ante fuit nec postea futurus est.
EXOD|11|7|Apud omnes autem filios Israel non mutiet canis contra hominem et pecus, ut sciatis quanto miraculo dividat Dominus Aegyptios et Israel.
EXOD|11|8|Descendentque omnes servi tui isti ad me et adorabunt me dicentes: "Egredere tu et omnis populus, qui sequitur te". Post haec egrediar ". Et exivit a pharaone iratus nimis.
EXOD|11|9|Dixit autem Dominus ad Moysen: " Non audiet vos pharao, ut multa signa fiant in terra Aegypti ".
EXOD|11|10|Moyses autem et Aaron fecerunt omnia ostenta haec coram pharaone; et induravit Dominus cor pharaonis, nec dimisit filios Israel de terra sua.
EXOD|12|1|Dixit Dominus ad Moysen et Aaron in terra Aegypti:
EXOD|12|2|" Mensis iste vobis principium mensium, primus erit in mensibus anni.
EXOD|12|3|Loquimini ad universum coetum filiorum Israel et dicite eis: Decima die mensis huius tollat unusquisque agnum per familias et domos suas.
EXOD|12|4|Sin autem minor est numerus, ut sufficere possit ad vescendum agnum, assumet vicinum suum, qui iunctus est domui suae, iuxta numerum animarum, quae sufficere possunt ad esum agni.
EXOD|12|5|Erit autem vobis agnus absque macula, masculus, anniculus; quem de agnis vel haedis tolletis
EXOD|12|6|et servabitis eum usque ad quartam decimam diem mensis huius; immolabitque eum universa congregatio filiorum Israel ad vesperam.
EXOD|12|7|Et sument de sanguine eius ac ponent super utrumque postem et in superliminaribus domorum, in quibus comedent illum;
EXOD|12|8|et edent carnes nocte illa assas igni et azymos panes cum lactucis amaris.
EXOD|12|9|Non comedetis ex eo crudum quid nec coctum aqua, sed tantum assum igni; caput cum pedibus eius et intestinis vorabitis.
EXOD|12|10|Nec remanebit quidquam ex eo usque mane; si quid residuum fuerit, igne comburetis.
EXOD|12|11|Sic autem comedetis illum: renes vestros accingetis, calceamenta habebitis in pedibus, tenentes baculos in manibus, et comedetis festinanter; est enim Pascha (id est Transitus) Domini!
EXOD|12|12|Et transibo per terram Aegypti nocte illa percutiamque omne primogenitum in terra Aegypti ab homine usque ad pecus; et in cunctis diis Aegypti faciam iudicia, ego Dominus.
EXOD|12|13|Erit autem sanguis vobis in signum in aedibus, in quibus eritis; et videbo sanguinem et transibo vos, nec erit in vobis plaga disperdens, quando percussero terram Aegypti.
EXOD|12|14|Habebitis autem hanc diem in monumentum et celebrabitis eam sollemnem Domino in generationibus vestris cultu sempiterno.
EXOD|12|15|Septem diebus azyma comedetis. Iam in die primo non erit fermentum in domibus vestris; quicumque comederit fermentatum, a primo die usque ad diem septimum, peribit anima illa de Israel.
EXOD|12|16|Dies prima erit sancta atque sollemnis, et dies septima eadem festivitate venerabilis. Nihil operis facietis in eis, exceptis his, quae ad vescendum pertinent.
EXOD|12|17|Et observabitis azyma, in eadem enim ipsa die eduxi exercitum vestrum de terra Aegypti; et custodietis diem istum in generationes vestras ritu perpetuo.
EXOD|12|18|Primo mense, quarta decima die mensis ad vesperam comedetis azyma; usque ad diem vicesimam primam eiusdem mensis ad vesperam.
EXOD|12|19|Septem diebus fermentum non invenietur in domibus vestris. Qui comederit fermentatum, peribit anima eius de coetu Israel, tam de advenis quam de indigenis terrae.
EXOD|12|20|Omne fermentatum non comedetis; in cunctis habitaculis vestris edetis azyma ".
EXOD|12|21|Vocavit autem Moyses omnes seniores filiorum Israel et dixit ad eos: " Ite tollentes animal per familias vestras et immolate Pascha.
EXOD|12|22|Fasciculumque hyssopi tingite in sanguine, qui est in pelvi, et aspergite ex eo superliminare et utrumque postem. Nullus vestrum egrediatur ostium domus suae usque mane.
EXOD|12|23|Transibit enim Dominus percutiens Aegyptios; cumque viderit sanguinem in superliminari et in utroque poste, transcendet ostium et non sinet percussorem ingredi domos vestras et laedere.
EXOD|12|24|Custodite verbum istud legitimum tibi et filiis tuis usque in aeternum.
EXOD|12|25|Cumque introieritis terram, quam Dominus daturus est vobis, ut pollicitus est, observabitis caeremonias istas;
EXOD|12|26|et, cum dixerint vobis filii vestri: "Quae est ista religio?",
EXOD|12|27|dicetis eis: "Victima Paschae Domino est, quando transivit super domos filiorum Israel in Aegypto percutiens Aegyptios et domos nostras liberans" ". Incurvatusque populus adoravit;
EXOD|12|28|et egressi filii Israel fecerunt, sicut praeceperat Dominus Moysi et Aaron.
EXOD|12|29|Factum est autem in noctis medio, percussit Dominus omne primogenitum in terra Aegypti, a primogenito pharaonis, qui in solio eius sedebat, usque ad primogenitum captivi, qui erat in carcere, et omne primogenitum iumentorum.
EXOD|12|30|Surrexitque pharao nocte et omnes servi eius cunctaque Aegyptus, et ortus est clamor magnus in Aegypto, neque enim erat domus, in qua non iaceret mortuus.
EXOD|12|31|Vocatisque pharao Moyse et Aaron nocte, ait: " Surgite, egredimini a populo meo, vos et filii Israel; ite, immolate Domino, sicut dicitis.
EXOD|12|32|Oves vestras et armenta assumite, ut petieratis, et abeuntes benedicite mihi ".
EXOD|12|33|Urgebantque Aegyptii populum de terra exire velociter dicentes: " Omnes moriemur ".
EXOD|12|34|Tulit igitur populus conspersam farinam, antequam fermentaretur; et ligans pistrina in palliis suis posuit super umeros suos.
EXOD|12|35|Feceruntque filii Israel, sicut praeceperat Moyses, et petierunt ab Aegyptiis vasa argentea et aurea vestemque plurimam.
EXOD|12|36|Dominus autem dedit gratiam populo coram Aegyptiis, ut commodarent eis; et spoliaverunt Aegyptios.
EXOD|12|37|Profectique sunt filii Israel de Ramesse in Succoth, sescenta fere milia peditum virorum absque parvulis.
EXOD|12|38|Sed et vulgus promiscuum innumerabile ascendit cum eis, oves et armenta, animantia multa nimis.
EXOD|12|39|Coxeruntque farinam, quam dudum de Aegypto conspersam tulerant, et fecerunt subcinericios panes azymos; neque enim poterant fermentari, cogentibus exire Aegyptiis et nullam facere sinentibus moram; nec pulmenti quidquam occurrerant praeparare.
EXOD|12|40|Habitatio autem filiorum Israel, qua manserant in Aegypto, fuit quadringentorum triginta annorum.
EXOD|12|41|Quibus expletis, eadem die egressus est omnis exercitus Domini de terra Aegypti.
EXOD|12|42|Nox ista vigiliarum Domino, quando eduxit eos de terra Aegypti: hanc observare debent Domino omnes filii Israel in generationibus suis.
EXOD|12|43|Dixitque Dominus ad Moysen et Aaron: " Haec est religio Paschae: Omnis alienigena non comedet ex eo;
EXOD|12|44|omnis autem servus empticius circumcidetur et sic comedet;
EXOD|12|45|advena et mercennarius non edent ex eo.
EXOD|12|46|In una domo comedetur, nec efferetis de carnibus eius foras nec os illius confringetis.
EXOD|12|47|Omnis coetus filiorum Israel faciet illud.
EXOD|12|48|Quod si quis peregrinorum in vestram voluerit transire coloniam et facere Pascha Domini, circumcidetur prius omne masculinum eius, et tunc rite celebrabit eritque sicut indigena terrae; si quis autem circumcisus non fuerit, non vescetur ex eo.
EXOD|12|49|Eadem lex erit indigenae et colono, qui peregrinatur apud vos ".
EXOD|12|50|Feceruntque omnes filii Israel, sicut praeceperat Dominus Moysi et Aaron;
EXOD|12|51|et in eadem die eduxit Dominus filios Israel de terra Aegypti per turmas suas.
EXOD|13|1|Locutusque est Dominus ad Moysen dicens:
EXOD|13|2|" Sanctifica mihi omne primogenitum, quod aperit vulvam in filiis Israel, tam de hominibus quam de iumentis: mea sunt enim omnia ".
EXOD|13|3|Et ait Moyses ad populum: " Mementote diei huius, in qua egressi estis de Aegypto et de domo servitutis, quoniam in manu forti eduxit vos Dominus de loco isto, ut non comedatis fermentatum panem.
EXOD|13|4|Hodie egredimini, mense Abib (id est novarum Frugum).
EXOD|13|5|Cumque introduxerit te Dominus in terram Chananaei et Hetthaei et Amorraei et Hevaei et Iebusaei, quam iuravit patribus tuis, ut daret tibi, terram fluentem lacte et melle; celebrabis hunc morem sacrorum mense isto.
EXOD|13|6|Septem diebus vesceris azymis, et in die septimo erit sollemnitas Domini.
EXOD|13|7|Azyma comedetis septem diebus: non apparebit apud te aliquid fermentatum nec in cunctis finibus tuis.
EXOD|13|8|Narrabisque filio tuo in die illo dicens: "Propter hoc, quod fecit mihi Dominus, quando egressus sum de Aegypto".
EXOD|13|9|Et erit quasi signum in manu tua et quasi monumentum inter oculos tuos, ut lex Domini semper sit in ore tuo; in manu enim forti eduxit te Dominus de Aegypto.
EXOD|13|10|Custodies huiuscemodi cultum statuto tempore a diebus in dies.
EXOD|13|11|Cumque introduxerit te Dominus in terram Chananaei, sicut iuravit tibi et patribus tuis, et dederit tibi eam,
EXOD|13|12|separabis omne, quod aperit vulvam, Domino et quod primitivum est in pecoribus tuis; quidquid habueris masculini sexus, consecrabis Domino.
EXOD|13|13|Primogenitum asini mutabis ove; quod, si non redemeris, interficies. Omne autem primogenitum hominis de filiis tuis pretio redimes.
EXOD|13|14|Cumque interrogaverit te filius tuus cras dicens: "Quid est hoc?", respondebis ei: "In manu forti eduxit nos Dominus de Aegypto, de domo servitutis.
EXOD|13|15|Nam, cum induratus esset pharao et nollet nos dimittere, occidit Dominus omne primogenitum in terra Aegypti, a primogenito hominis usque ad primogenitum iumentorum; idcirco immolo Domino omne, quod aperit vulvam, masculini sexus, et omnia primogenita filiorum meorum redimo".
EXOD|13|16|Erit igitur quasi signum in manu tua et quasi appensum quid ob recordationem inter oculos tuos, eo quod in manu forti eduxit nos Dominus de Aegypto ".
EXOD|13|17|Igitur cum emisisset pharao populum, non eos duxit Deus per viam terrae Philisthim, quae vicina est, reputans ne forte paeniteret populum, si vidisset adversum se bella consurgere, et reverteretur in Aegyptum,
EXOD|13|18|sed circumduxit per viam deserti, quae est iuxta mare Rubrum. Et armati ascenderunt filii Israel de terra Aegypti.
EXOD|13|19|Tulit quoque Moyses ossa Ioseph secum, eo quod adiurasset filios Israel dicens: " Visitabit vos Deus; efferte ossa mea hinc vobiscum ".
EXOD|13|20|Profectique de Succoth castrametati sunt in Etham, in extremis finibus solitudinis.
EXOD|13|21|Dominus autem praecedebat eos ad ostendendam viam per diem in columna nubis et per noctem in columna ignis, ut dux esset itineris utroque tempore.
EXOD|13|22|Nunquam defuit columna nubis per diem, nec columna ignis per noctem, coram populo.
EXOD|14|1|Locutus est autem Dominus ad Moysen dicens:
EXOD|14|2|" Lo quere filiis Israel: Reversi castrametentur e regione Phihahiroth, quae est inter Magdolum et mare contra Beelsephon; in conspectu eius castra ponetis super mare.
EXOD|14|3|Dicturusque est pharao super filiis Israel: "Errant in terra, conclusit eos desertum".
EXOD|14|4|Et indurabo cor eius, ac persequetur eos, et glorificabor in pharaone et in omni exercitu eius; scientque Aegyptii quia ego sum Dominus ". Feceruntque ita.
EXOD|14|5|Et nuntiatum est regi Aegyptiorum quod fugisset populus; immutatumque est cor pharaonis et servorum eius super populo, et dixerunt: " Quid hoc fecimus, ut dimitteremus Israel, ne servirent nobis? ".
EXOD|14|6|Iunxit ergo currum et omnem populum suum assumpsit secum;
EXOD|14|7|tulitque sescentos currus electos et quidquid in Aegypto curruum fuit et bellatores in singulis curribus.
EXOD|14|8|Induravitque Dominus cor pharaonis regis Aegypti, et persecutus est filios Israel; at illi egressi erant in manu excelsa.
EXOD|14|9|Cumque persequerentur Aegyptii vestigia praecedentium, reppererunt eos in castris super mare; omnes equi et currus pharaonis, equites et exercitus eius erant in Phihahiroth contra Beelsephon.
EXOD|14|10|Cumque appropinquasset pharao, levantes filii Israel oculos viderunt Aegyptios post se et timuerunt valde clamaveruntque ad Dominum
EXOD|14|11|et dixerunt ad Moysen: " Forsitan non erant sepulcra in Aegypto? Ideo tulisti nos, ut moreremur in solitudine. Quid hoc fecisti, ut educeres nos ex Aegypto?
EXOD|14|12|Nonne iste est sermo, quem loquebamur ad te in Aegypto dicentes: Recede a nobis, ut serviamus Aegyptiis? Multo enim melius erat servire eis quam mori in solitudine ".
EXOD|14|13|Et ait Moyses ad populum: " Nolite timere; state et videte salutem Domini, quam facturus est vobis hodie; Aegyptios enim, quos nunc videtis, nequaquam ultra videbitis usque in sempiternum.
EXOD|14|14|Dominus pugnabit pro vobis, et vos silebitis ".
EXOD|14|15|Dixitque Dominus ad Moysen: " Quid clamas ad me? Loquere filiis Israel, ut proficiscantur.
EXOD|14|16|Tu autem eleva virgam tuam et extende manum tuam super mare et divide illud, ut gradiantur filii Israel in medio mari per siccum.
EXOD|14|17|Ego autem indurabo cor Aegyptiorum, ut persequantur eos; et glorificabor in pharaone et in omni exercitu eius, in curribus et in equitibus illius.
EXOD|14|18|Et scient Aegyptii quia ego sum Dominus, cum glorificatus fuero in pharaone, in curribus atque in equitibus eius ".
EXOD|14|19|Tollensque se angelus Dei, qui praecedebat castra Israel, abiit post eos; et cum eo pariter columna nubis, priora dimittens, post tergum.
EXOD|14|20|Stetit inter castra Aegyptiorum et castra Israel; et erat nubes tenebrosa et illuminans noctem, ita ut ad se invicem toto noctis tempore accedere non valerent.
EXOD|14|21|Cumque extendisset Moyses manum super mare, reppulit illud Dominus, flante vento vehementi et urente tota nocte, et vertit in siccum; divisaque est aqua.
EXOD|14|22|Et ingressi sunt filii Israel per medium maris sicci; erat enim aqua quasi murus a dextra eorum et laeva.
EXOD|14|23|Persequentesque Aegyptii ingressi sunt post eos, omnis equitatus pharaonis, currus eius et equites per medium maris.
EXOD|14|24|Iamque advenerat vigilia matutina, et ecce respiciens Dominus super castra Aegyptiorum per columnam ignis et nubis perturbavit exercitum eorum;
EXOD|14|25|et impedivit rotas curruum, ita ut difficile moverentur. Dixerunt ergo Aegyptii: " Fugiamus Israelem! Dominus enim pugnat pro eis contra nos ".
EXOD|14|26|Et ait Dominus ad Moysen: " Extende manum tuam super mare, ut revertantur aquae ad Aegyptios super currus et equites eorum ".
EXOD|14|27|Cumque extendisset Moyses manum contra mare, reversum est primo diluculo ad priorem locum; fugientibusque Aegyptiis occurrerunt aquae, et involvit eos Dominus in mediis fluctibus.
EXOD|14|28|Reversaeque sunt aquae et operuerunt currus et equites cuncti exercitus pharaonis, qui sequentes ingressi fuerant mare; ne unus quidem superfuit ex eis.
EXOD|14|29|Filii autem Israel perrexerunt per medium sicci maris, et aquae eis erant quasi pro muro a dextris et a sinistris.
EXOD|14|30|Liberavitque Dominus in die illo Israel de manu Aegyptiorum. Et viderunt Aegyptios mortuos super litus maris
EXOD|14|31|et manum magnam, quam exercuerat Dominus contra eos; timuitque populus Dominum et crediderunt Domino et Moysi servo eius.
EXOD|15|1|Tunc cecinit Moyses et filii Israel carmen hoc Domino, et dixerunt:" Cantemus Domino,gloriose enim magnificatus est:equum et ascensorem eiusdeiecit in mare!
EXOD|15|2|Fortitudo mea et robur meum Dominus,et factus est mihi in salutem.Iste Deus meus,et glorificabo eum;Deus patris mei,et exaltabo eum!
EXOD|15|3|Dominus quasi vir pugnator;Dominus nomen eius!
EXOD|15|4|Currus pharaonis et exercitum eiusproiecit in mare;electi bellatores eiussubmersi sunt in mari Rubro.
EXOD|15|5|Abyssi operuerunt eos,descenderunt in profundum quasi lapis.
EXOD|15|6|Dextera tua, Domine,magnifice in fortitudine,dextera tua, Domine,percussit inimicum.
EXOD|15|7|Et in multitudine gloriae tuaedeposuisti adversarios tuos;misisti iram tuam,quae devoravit eos sicut stipulam.
EXOD|15|8|Et in spiritu furoris tuicongregatae sunt aquae;stetit ut aggerunda fluens,coagulatae sunt abyssiin medio mari.
EXOD|15|9|Dixit inimicus:"Persequar, comprehendam,dividam spolia,implebitur anima mea;evaginabo gladium meum,interficiet eos manus mea!".
EXOD|15|10|Flavit spiritus tuus,et operuit eos mare;submersi sunt quasi plumbumin aquis vehementibus.
EXOD|15|11|Quis similis tuiin diis, Domine?Quis similis tui,magnificus in sanctitate,terribilis atque laudabilis,faciens mirabilia?
EXOD|15|12|Extendisti manum tuam,devoravit eos terra.
EXOD|15|13|Dux fuisti in misericordia tuapopulo, quem redemisti,et portasti eum in fortitudine tuaad habitaculum sanctum tuum.
EXOD|15|14|Attenderunt populi et commoti sunt,dolores obtinuerunt habitatores Philisthaeae.
EXOD|15|15|Tunc conturbati sunt principes Edom,potentes Moab obtinuit tremor,obriguerunt omnes habitatores Chanaan.
EXOD|15|16|Irruit super eosformido et pavor;in magnitudine brachii tuifiunt immobiles quasi lapis,donec pertranseat populus tuus, Domine,donec pertranseat populus tuus iste,quem possedisti.
EXOD|15|17|Introduces eos et plantabisin monte hereditatis tuae,firmissimo habitaculo tuo,quod operatus es, Domine,sanctuario, Domine,quod firmaverunt manus tuae.
EXOD|15|18|Dominus regnabitin aeternum et ultra! ".
EXOD|15|19|Ingressi sunt enim equi pharaonis cum curribus et equitibus eius in mare, et reduxit super eos Dominus aquas maris; filii autem Israel ambu laverunt per siccum in medio eius.
EXOD|15|20|Sumpsit ergo Maria prophetissa soror Aaron tympanum in manu sua; egressaeque sunt omnes mulieres post eam cum tympanis et choris,
EXOD|15|21|quibus praecinebat dicens:" Cantemus Domino,gloriose enim magnificatus est:equum et ascensorem eiusdeiecit in mare! ".
EXOD|15|22|Tulit autem Moyses Israel de mari Rubro, et egressi sunt in desertum Sur; ambulaveruntque tribus diebus per solitudinem et non inveniebant aquam.
EXOD|15|23|Et venerunt in Mara nec poterant bibere aquas de Mara, eo quod essent amarae; unde vocatum est nomen eius Mara (id est Amaritudo).
EXOD|15|24|Et murmuravit populus contra Moysen dicens: " Quid bibemus? ".
EXOD|15|25|At ille clamavit ad Dominum, qui ostendit ei lignum; quod cum misisset in aquas, in dulcedinem versae sunt. Ibi constituit ei praecepta atque iudicia et ibi tentavit eum
EXOD|15|26|dicens: " Si audieris vocem Domini Dei tui et, quod rectum est coram eo, feceris et oboedieris mandatis eius custodierisque omnia praecepta illius, cunctum languorem, quem posui in Aegypto, non inducam super te: Ego enim Dominus sanator tuus ".
EXOD|15|27|Venerunt autem in Elim, ubi erant duodecim fontes aquarum et septuaginta palmae; et castrametati sunt iuxta aquas.
EXOD|16|1|Profectique sunt de Elim, et venit omnis congregatio filio rum Israel in desertum Sin, quod est inter Elim et Sinai, quinto decimo die mensis secundi postquam egressi sunt de terra Aegypti.
EXOD|16|2|Et murmuravit omnis congregatio filiorum Israel contra Moysen et Aaron in solitudine,
EXOD|16|3|dixeruntque filii Israel ad eos: " Utinam mortui essemus per manum Domini in terra Aegypti, quando sedebamus super ollas carnium et comedebamus panem in saturitate. Cur eduxistis nos in desertum istud, ut occideretis omnem coetum fame? ".
EXOD|16|4|Dixit autem Dominus ad Moysen: " Ecce ego pluam vobis panes de caelo; egrediatur populus et colligat, quae sufficiunt per singulos dies, ut tentem eum, utrum ambulet in lege mea an non.
EXOD|16|5|Die autem sexta parabunt quod intulerint, et duplum erit quam colligere solebant per singulos dies ".
EXOD|16|6|Dixeruntque Moyses et Aaron ad omnes filios Israel:" Vespere scietisquod Dominus eduxerit vosde terra Aegypti;
EXOD|16|7|et mane videbitisgloriam Domini.Audivit enim murmur vestrum contra Dominum. Nos vero quid sumus, quia mussitatis contra nos? ".
EXOD|16|8|Et ait Moyses:" Dabit Dominus vobisvespere carnes edereet mane panes in saturitate,eo quod audierit murmurationes vestras, quibus murmurati estis contra eum. Nos enim quid sumus? Nec contra nos est murmur vestrum, sed contra Dominum ".
EXOD|16|9|Dixitque Moyses ad Aaron: " Dic universae congregationi filiorum Israel: Accedite coram Domino; audivit enim murmur ve strum ".
EXOD|16|10|Cumque loqueretur Aaron ad omnem coetum filiorum Israel, respexerunt ad solitudinem, et ecce gloria Domini apparuit in nube.
EXOD|16|11|Locutus est autem Dominus ad Moysen dicens:
EXOD|16|12|" Audivi murmurationes filiorum Israel. Loquere ad eos: Vespere comedetis carnes et mane saturabimini panibus scietisque quod ego sum Dominus Deus vester ".
EXOD|16|13|Factum est ergo vespere, et ascendens coturnix operuit castra; mane quoque ros iacuit per circuitum castrorum.
EXOD|16|14|Cumque operuisset superficiem deserti, apparuit minutum et squamatum in similitudinem pruinae super terram.
EXOD|16|15|Quod cum vidissent filii Israel, dixerunt ad invicem: " Manhu? " (quod significat: " Quid est hoc? "). Ignorabant enim quid esset. Quibus ait Moyses: " Iste est panis, quem dedit Dominus vobis ad vescendum.
EXOD|16|16|Hic est sermo, quem praecepit Dominus: "Colligat ex eo unusquisque quantum sufficiat ad vescendum; gomor per singula capita iuxta numerum animarum vestrarum, quae habitant in tabernaculo, sic tolletis" ".
EXOD|16|17|Feceruntque ita filii Israel; et collegerunt alius plus, alius minus.
EXOD|16|18|Et mensi sunt ad mensuram gomor; nec qui plus collegerat, habuit amplius, nec qui minus paraverat, repperit minus, sed singuli, iuxta id quod edere poterant, congregaverunt.
EXOD|16|19|Dixitque Moyses ad eos: " Nullus relinquat ex eo in mane ".
EXOD|16|20|Qui non audierunt eum, sed dimiserunt quidam ex eis usque mane, et scatere coepit vermibus atque computruit; et iratus est contra eos Moyses.
EXOD|16|21|Colligebant autem mane singuli, quantum sufficere poterat ad vescendum; cumque incaluisset sol, liquefiebat.
EXOD|16|22|In die autem sexta collegerunt cibos duplices, id est duo gomor per singulos homines. Venerunt autem omnes principes congregationis et narraverunt Moysi.
EXOD|16|23|Qui ait eis: " Hoc est quod locutus est Dominus: Requies, sabbatum sanctum Domino cras; quodcumque torrendum est, torrete et, quae coquenda sunt, coquite; quidquid autem reliquum fuerit, reponite usque in mane ".
EXOD|16|24|Feceruntque ita, ut praeceperat Moyses, et non computruit, neque vermis inventus est in eo.
EXOD|16|25|Dixitque Moyses: " Comedite illud hodie, quia sabbatum est Domino; non invenietur hodie in agro.
EXOD|16|26|Sex diebus colligite; in die autem septimo sabbatum est Domino, idcirco non invenietur in eo ".
EXOD|16|27|Venitque septima dies; et egressi de populo, ut colligerent, non invenerunt.
EXOD|16|28|Dixit autem Dominus ad Moysen: " Usquequo non vultis custodire mandata mea et legem meam?
EXOD|16|29|Videte quod Dominus dederit vobis sabbatum et propter hoc die sexta tribuit vobis cibos duplices; maneat unusquisque apud semetipsum, nullus egrediatur de loco suo die septimo ".
EXOD|16|30|Et sabbatizavit populus die septimo.
EXOD|16|31|Appellavitque domus Israel nomen eius Man: quod erat quasi semen coriandri album, gustusque eius quasi similae cum melle.
EXOD|16|32|Dixit autem Moyses: " Iste est sermo, quem praecepit Dominus: "Imple gomor ex eo, et custodiatur in generationes vestras, ut noverint panem, quo alui vos in solitudine, quando educti estis de terra Aegypti" ".
EXOD|16|33|Dixitque Moyses ad Aaron: " Sume vas unum et mitte ibi man, quantum potest capere gomor; et repone coram Domino ad servandum in generationes vestras ".
EXOD|16|34|Sicut praecepit Dominus Moysi, posuit illud Aaron coram testimonio reservandum.
EXOD|16|35|Filii autem Israel comederunt man quadraginta annis, donec venirent in terram habitabilem; hoc cibo aliti sunt, usquequo tangerent fines terrae Chanaan.
EXOD|16|36|Gomor autem decima pars est ephi.
EXOD|17|1|Igitur profecta omnis congregatio filiorum Israel de deserto Sin per mansiones suas iuxta sermonem Domini, castrametati sunt in Raphidim, ubi non erat aqua ad bibendum populo.
EXOD|17|2|Qui iurgatus contra Moysen ait: " Da nobis aquam, ut bibamus ". Quibus respondit Moyses: " Quid iurgamini contra me? Cur tentatis Dominum? ".
EXOD|17|3|Sitivit ergo ibi populus prae aquae penuria et murmuravit contra Moysen dicens: " Cur fecisti nos exire de Aegypto, ut occideres nos et liberos nostros ac iumenta siti? ".
EXOD|17|4|Clamavit autem Moyses ad Dominum dicens: " Quid faciam populo huic? Adhuc paululum et lapidabunt me ".
EXOD|17|5|Et ait Dominus ad Moysen: " Antecede populum et sume tecum de senioribus Israel, et virgam, qua percussisti fluvium, tolle in manu tua et vade.
EXOD|17|6|En ego stabo coram te ibi super petram Horeb; percutiesque petram, et exibit ex ea aqua, ut bibat populus ". Fecit Moyses ita coram senioribus Israel.
EXOD|17|7|Et vocavit nomen loci illius Massa et Meriba, propter iurgium filiorum Israel et quia tentaverunt Dominum dicentes: " Estne Dominus in nobis an non? ".
EXOD|17|8|Venit autem Amalec et pugnabat contra Israel in Raphidim.
EXOD|17|9|Dixitque Moyses ad Iosue: " Elige nobis viros et egressus pugna contra Amalec; cras ego stabo in vertice collis habens virgam Dei in manu mea ".
EXOD|17|10|Fecit Iosue, ut locutus erat ei Moyses, et pugnavit contra Amalec; Moyses autem et Aaron et Hur ascenderunt super verticem collis.
EXOD|17|11|Cumque levaret Moyses manus, vincebat Israel; sin autem remisisset, superabat Amalec.
EXOD|17|12|Manus autem Moysi erant graves; sumentes igitur lapidem posuerunt subter eum, in quo sedit; Aaron autem et Hur sustentabant manus eius ex utraque parte. Et factum est ut manus eius non lassarentur usque ad occasum solis.
EXOD|17|13|Vicitque Iosue Amalec et populum eius in ore gladii.
EXOD|17|14|Dixit autem Dominus ad Moysen: " Scribe hoc ob monumentum in libro et trade auribus Iosue; delebo enim memoriam Amalec sub caelo ".
EXOD|17|15|Aedificavitque Moyses altare et vocavit nomen eius Dominus Nissi "Dominus vexillum meum)
EXOD|17|16|dicens:" Quia manus contra solium Domini:bellum Domino erit contra Amalec a generatione in generationem ".
EXOD|18|1|Cumque audisset Iethro sacerdos Madian socer Moysi omnia, quae fecerat Deus Moysi et Israel populo suo, eo quod eduxisset Dominus Israel de Aegypto,
EXOD|18|2|tulit Sephoram uxorem Moysi, quam remiserat,
EXOD|18|3|et duos filios eius, quorum unus vocabatur Gersam, dicente patre: " Advena fui in terra aliena ",
EXOD|18|4|alter vero Eliezer: " Deus enim, ait, patris mei adiutor meus, et eruit me de gladio pharaonis ".
EXOD|18|5|Venit ergo Iethro socer Moysi et filii eius et uxor eius ad Moysen in desertum, ubi erat castrametatus iuxta montem Dei;
EXOD|18|6|et mandavit Moysi dicens: " Ego socer tuus Iethro venio ad te et uxor tua et duo filii tui cum ea ".
EXOD|18|7|Qui egressus in occursum soceri sui adoravit et osculatus est eum, salutaveruntque se mutuo verbis pacificis. Cumque intrasset tabernaculum,
EXOD|18|8|narravit Moyses socero suo cuncta, quae fecerat Dominus pharaoni et Aegyptiis propter Israel, universumque laborem, qui accidisset eis in itinere, et quod liberaverat eos Dominus.
EXOD|18|9|Laetatusque est Iethro super omnibus bonis, quae fecerat Dominus Israel, eo quod eruisset eum de manu Aegyptiorum,
EXOD|18|10|et ait: " Benedictus Dominus, qui liberavit vos de manu Aegyptiorum et de manu pharaonis.
EXOD|18|11|Nunc cognovi quia magnus Dominus super omnes deos, eo quod eruerit populum de manu Aegyptiorum, qui superbe egerunt contra illos ".
EXOD|18|12|Obtulit ergo Iethro socer Moysi holocausta et hostias Deo; veneruntque Aaron et omnes seniores Israel, ut comederent panem cum eo coram Deo.
EXOD|18|13|Altero autem die sedit Moyses, ut iudicaret populum, qui assistebat Moysi de mane usque ad vesperam.
EXOD|18|14|Quod cum vidisset socer eius, omnia scilicet, quae agebat in populo, ait: " Quid est hoc, quod facis in plebe? Cur solus sedes, et omnis populus praestolatur de mane usque ad vesperam? ".
EXOD|18|15|Cui respondit Moyses: " Venit ad me populus quaerens sententiam Dei.
EXOD|18|16|Cumque acciderit eis aliqua disceptatio, veniunt ad me, ut iudicem inter eos et ostendam praecepta Dei et leges eius ".
EXOD|18|17|At ille: " Non bonam, inquit, rem facis.
EXOD|18|18|Consumeris et tu et populus iste, qui tecum est. Ultra vires tuas est negotium; solus illud non poteris sustinere.
EXOD|18|19|Sed audi verba mea atque consilia, et erit Deus tecum: Esto tu populo in his, quae ad Deum pertinent, ut referas causas ad Deum
EXOD|18|20|ostendasque populo praecepta et leges viamque, per quam ingredi debeant, et opus, quod facere debeant.
EXOD|18|21|Provide autem de omni plebe viros strenuos et timentes Deum, in quibus sit veritas, et qui oderint avaritiam, et constitue ex eis tribunos et centuriones et quinquagenarios et decanos,
EXOD|18|22|qui iudicent populum omni tempore. Quidquid autem maius fuerit, referant ad te, et ipsi minora tantummodo iudicent; leviusque sit tibi, partito cum aliis onere.
EXOD|18|23|Si hoc feceris, implebis imperium Dei et praecepta eius poteris sustentare, et omnis hic populus revertetur ad loca sua cum pace ".
EXOD|18|24|Quibus auditis, Moyses fecit omnia, quae ille suggesserat;
EXOD|18|25|et, electis viris strenuis de cuncto Israel, constituit eos principes populi, tribunos et centuriones et quinquagenarios et decanos,
EXOD|18|26|qui iudicabant plebem omni tempore. Quidquid autem gravius erat, referebant ad eum, faciliora tantummodo iudicantes.
EXOD|18|27|Dimisitque socerum suum, qui reversus abiit in terram suam.
EXOD|19|1|Mense tertio egressionis Israel de terra Aegypti, in die hac venerunt in solitudinem Sinai.
EXOD|19|2|Nam profecti de Raphidim et pervenientes usque in desertum Sinai, castrametati sunt in eodem loco,ibique Israel fixit tentoria e regione montis.
EXOD|19|3|Moyses autem ascendit ad Deum, vocavitque eum Dominus de monte et ait:" Haec dices domui Iacobet annuntiabis filiis Israel:
EXOD|19|4|Vos ipsi vidistis, quae fecerim Aegyptiis,quomodo portaverim vos super alas aquilarumet adduxerim ad me.
EXOD|19|5|Si ergo audieritis vocem meamet custodieritis pactum meum,eritis mihi in peculium de cunctis populis;mea est enim omnis terra.
EXOD|19|6|Et vos eritis mihi regnum sacerdotumet gens sancta.Haec sunt verba, quae loqueris ad filios Israel ".
EXOD|19|7|Venit Moyses et, convocatis maioribus natu populi, exposuit omnes sermones, quos mandaverat Dominus.
EXOD|19|8|Responditque universus populus simul: " Cuncta, quae locutus est Dominus, faciemus ". Cumque rettulisset Moyses verba populi ad Dominum,
EXOD|19|9|ait ei Dominus: " Ecce ego veniam ad te in caligine nubis, ut audiat me populus loquentem ad te et tibi quoque credat in perpetuum ".Nuntiavit ergo Moyses verba populi ad Dominum,
EXOD|19|10|qui dixit ei: " Vade ad populum et sanctifica illos hodie et cras; laventque vestimenta sua
EXOD|19|11|et sint parati in diem tertium. In die enim tertio descendet Dominus coram omni plebe super montem Sinai.
EXOD|19|12|Constituesque terminos populo per circuitum et dices: Cavete, ne ascendatis in montem nec tangatis fines illius; omnis, qui tetigerit montem, morte morietur.
EXOD|19|13|Manus non tanget eum, sed lapidibus opprimetur aut confodietur iaculis; sive iumentum fuerit, sive homo, non vivet. Cum coeperit clangere bucina, tunc ascendant in montem ".
EXOD|19|14|Descenditque Moyses de monte ad populum et sanctificavit eum; cumque lavissent vestimenta sua,
EXOD|19|15|ait ad eos: " Estote parati in diem tertium; ne appropinquetis uxoribus vestris ".
EXOD|19|16|Iamque advenerat tertius dies, et mane inclaruerat; et ecce coeperunt audiri tonitrua ac micare fulgura et nubes densissima operire montem, clangorque bucinae vehementius perstrepebat; et timuit populus, qui erat in castris.
EXOD|19|17|Cumque eduxisset eos Moyses in occursum Dei de loco castrorum, steterunt ad radices montis.
EXOD|19|18|Totus autem mons Sinai fumabat, eo quod descendisset Dominus super eum in igne, et ascenderet fumus ex eo quasi de fornace. Et tremuit omnis mons vehementer.
EXOD|19|19|Et sonitus bucinae paulatim crescebat in maius; Moyses loquebatur, et Deus respondebat ei cum voce.
EXOD|19|20|Descenditque Dominus super montem Sinai in ipso montis vertice et vocavit Moysen in cacumen eius. Quo cum ascendisset,
EXOD|19|21|dixit ad eum: " Descende et contestare populum, ne velit transcendere terminos ad videndum Dominum, et pereat ex eis plurima multitudo.
EXOD|19|22|Sacerdotes quoque, qui accedunt ad Dominum, sanctificentur, ne percutiat eos ".
EXOD|19|23|Dixitque Moyses ad Dominum: " Non poterit vulgus ascendere in montem Sinai, tu enim testificatus es et iussisti dicens: "Pone terminos circa montem et sanctifica illum" ".
EXOD|19|24|Cui ait Dominus: " Vade, descende; ascendesque tu et Aaron tecum, sacerdotes autem et populus ne transeant terminos nec ascendant ad Dominum, ne interficiat illos ".
EXOD|19|25|Descenditque Moyses ad populum et omnia narravit eis.
EXOD|20|1|Locutusque est Deus cunctos sermones hos:
EXOD|20|2|" Ego sum Dominus Deus tuus, qui eduxi te de terra Aegypti, de domo servitutis.
EXOD|20|3|Non habebis deos alienos coram me.
EXOD|20|4|Non facies tibi sculptile neque omnem similitudinem eorum, quae sunt in caelo desuper et quae in terra deorsum et quae in aquis sub terra.
EXOD|20|5|Non adorabis ea neque coles, quia ego sum Dominus Deus tuus, Deus zelotes, visitans iniquitatem patrum in filiis in tertiam et quartam generationem eorum, qui oderunt me,
EXOD|20|6|et faciens misericordiam in milia his, qui diligunt me et custodiunt praecepta mea.
EXOD|20|7|Non assumes nomen Domini Dei tui in vanum, nec enim habebit insontem Dominus eum, qui assumpserit nomen Domini Dei sui frustra.
EXOD|20|8|Memento, ut diem sabbati sanctifices.
EXOD|20|9|Sex diebus operaberis et facies omnia opera tua;
EXOD|20|10|septimus autem dies sabbatum Domino Deo tuo est; non facies omne opus tu et filius tuus et filia tua, servus tuus et ancilla tua, iumentum tuum et advena, qui est intra portas tuas.
EXOD|20|11|Sex enim diebus fecit Dominus caelum et terram et mare et omnia, quae in eis sunt, et requievit in die septimo; idcirco benedixit Dominus diei sabbati et sanctificavit eum.
EXOD|20|12|Honora patrem tuum et matrem tuam, ut sis longaevus super terram, quam Dominus Deus tuus dabit tibi.
EXOD|20|13|Non occides.
EXOD|20|14|Non moechaberis.
EXOD|20|15|Non furtum facies.
EXOD|20|16|Non loqueris contra proximum tuum falsum testimonium.
EXOD|20|17|Non concupisces domum proximi tui: non desiderabis uxorem eius, non servum, non ancillam, non bovem, non asinum nec omnia, quae illius sunt ".
EXOD|20|18|Cunctus autem populus videbat voces et lampades et sonitum bucinae montemque fumantem; et perterriti ac pavore concussi steterunt procul
EXOD|20|19|dicentes Moysi: " Loquere tu nobis, et audiemus; non loquatur nobis Deus, ne moriamur ".
EXOD|20|20|Et ait Moyses ad populum: " Nolite timere; ut enim probaret vos, venit Deus, et ut timor illius esset in vobis, ne peccaretis ".
EXOD|20|21|Stetitque populus de longe; Moyses autem accessit ad caliginem, in qua erat Deus.
EXOD|20|22|Dixit praeterea Dominus ad Moysen: " Haec dices filiis Israel: Vos vidistis quod de caelo locutus sim vobis.
EXOD|20|23|Non facietis praeter me deos argenteos nec deos aureos facietis vobis.
EXOD|20|24|Altare de terra facietis mihi et offeretis super eo holocausta et pacifica vestra, oves vestras et boves; in omni loco, in quo memoriam fecero nominis mei, veniam ad te et benedicam tibi.
EXOD|20|25|Quod si altare lapideum feceris mihi, non aedificabis illud de sectis lapidibus; si enim levaveris cultrum super eo, polluetur.
EXOD|20|26|Non ascendes per gradus ad altare meum, ne reveletur turpitudo tua.
EXOD|21|1|Haec sunt iudicia, quae propones eis:
EXOD|21|2|Si emeris servum Hebraeum, sex annis serviet tibi; in septimo egredietur liber gratis.
EXOD|21|3|Si solus intraverit, solus exeat; si habens uxorem, et uxor egredietur simul.
EXOD|21|4|Sin autem dominus dederit illi uxorem, et pepererit filios et filias, mulier et liberi eius erunt domini sui; ipse vero exibit solus.
EXOD|21|5|Quod si dixerit servus: "Diligo dominum meum et uxorem ac liberos, non egrediar liber",
EXOD|21|6|afferet eum dominus ad Deum et applicabit eum ad ostium vel postes perforabitque aurem eius subula; et erit ei servus in saeculum.
EXOD|21|7|Si quis vendiderit filiam suam in famulam, non egredietur sicut servi exire consueverunt.
EXOD|21|8|Si displicuerit oculis domini sui, cui tradita fuerat, faciat eam redimi; populo autem alieno vendendi non habebit potestatem, quia fraudavit eam.
EXOD|21|9|Sin autem filio suo desponderit eam, iuxta morem filiarum faciet illi.
EXOD|21|10|Quod si alteram sibi acceperit, cibum et vestimentum et concubitum non negabit.
EXOD|21|11|Si tria ista non fecerit ei, egredietur gratis absque pretio.
EXOD|21|12|Qui percusserit hominem, et ille mortuus fuerit, morte moriatur.
EXOD|21|13|Qui autem non est insidiatus, sed Deus illum tradidit in manus eius, constituam tibi locum, in quem fugere debeat.
EXOD|21|14|Si quis de industria occiderit proximum suum et per insidias, ab altari meo evelles eum, ut moriatur.
EXOD|21|15|Qui percusserit patrem suum aut matrem, morte moriatur.
EXOD|21|16|Qui furatus fuerit hominem sive vendiderit eum sive inventus fuerit in manu eius, morte moriatur.
EXOD|21|17|Qui maledixerit patri suo vel matri, morte moriatur.
EXOD|21|18|Si rixati fuerint viri, et percusserit alter proximum suum lapide vel pugno, et ille mortuus non fuerit, sed iacuerit in lectulo,
EXOD|21|19|si surrexerit et ambulaverit foris super baculum suum, impunitus erit, qui percusserit, ita tamen, ut operas eius deperditas et impensas pro medela restituat.
EXOD|21|20|Qui percusserit servum suum vel ancillam virga, et mortui fuerint in manibus eius, ultioni subiacetur.
EXOD|21|21|Sin autem uno die vel duobus supervixerit, non subiacebit poenae, quia pecunia illius est.
EXOD|21|22|Si rixati fuerint viri, et percusserit quis mulierem praegnantem et abortivum quidem fecerit, sed aliud quid adversi non acciderit, subiacebit damno, quantum maritus mulieris expetierit, et arbitri iudicaverint.
EXOD|21|23|Sin autem quid adversi acciderit, reddet animam pro anima,
EXOD|21|24|oculum pro oculo, dentem pro dente, manum pro manu, pedem pro pede,
EXOD|21|25|adustionem pro adustione, vulnus pro vulnere, livorem pro livore.
EXOD|21|26|Si percusserit quispiam oculum servi sui aut ancillae et luscos eos fecerit, dimittet eos liberos pro oculo.
EXOD|21|27|Dentem quoque si excusserit servo vel ancillae suae, dimittet eos liberos pro dente.
EXOD|21|28|Si bos cornu percusserit virum aut mulierem, et mortui fuerint, lapidibus obruetur, et non comedentur carnes eius; dominus autem bovis innocens erit.
EXOD|21|29|Quod si bos cornupeta fuerit ab heri et nudiustertius, et contestati sunt dominum eius, nec recluserit eum, occideritque virum aut mulierem: et bos lapidibus obruetur, et dominum illius occident.
EXOD|21|30|Quod si pretium ei fuerit impositum, dabit pro anima sua, quidquid fuerit postulatus.
EXOD|21|31|Filium quoque vel filiam si cornu percusserit, simili sententiae subiacebit.
EXOD|21|32|Si servum vel ancillam invaserit, triginta siclos argenti dabit domino; bos vero lapidibus opprimetur.
EXOD|21|33|Si quis aperuerit cisternam vel foderit et non operuerit eam, cedideritque bos vel asinus in eam,
EXOD|21|34|dominus cisternae reddet pretium iumentorum; quod autem mortuum est, ipsius erit.
EXOD|21|35|Si bos alienus bovem alterius vulneraverit, et ille mortuus fuerit, vendent bovem vivum et divident pretium; cadaver autem mortui inter se dispertient.
EXOD|21|36|Sin autem notum erat quod bos cornupeta esset ab heri et nudiustertius, et non custodivit eum dominus suus, reddet bovem pro bove et cadaver integrum accipiet.
EXOD|21|37|Si quis furatus fuerit bovem aut ovem et occiderit vel vendiderit, quinque boves pro uno bove restituet et quattuor oves pro una ove.
EXOD|22|1|Si effringens fur domum sive suffodiens fuerit inventus et, accepto vulnere, mortuus fuerit, percussor non erit reus sanguinis.
EXOD|22|2|Quod si orto sole hoc fecerit, erit reus sanguinis. Fur plene restituet. Si non habuerit, quod reddat, venumdabitur pro furto.
EXOD|22|3|Si inventum fuerit apud eum, quod furatus est, vivens sive bos sive asinus sive ovis, duplum restituet.
EXOD|22|4|Si quispiam depasci permiserit agrum vel vineam et dimiserit iumentum suum, ut depascatur agrum alienum, restituet plene ex agro suo secundum fruges eius; si autem totum agrum depastum fuerit, quidquid optimum habuerit in agro suo vel in vinea, restituet.
EXOD|22|5|Si egressus ignis invenerit spinas et comprehenderit acervos frugum sive stantes segetes sive agrum, reddet damnum, qui ignem succenderit.
EXOD|22|6|Si quis commendaverit amico pecuniam aut vasa in custodiam, et ab eo, qui susceperat, furto ablata fuerint, si invenitur fur, duplum reddet.
EXOD|22|7|Si latet fur, dominus domus applicabitur ad Deum et iurabit quod non extenderit manum in rem proximi sui.
EXOD|22|8|In omni causa fraudis tam de bove quam de asino et ove ac vestimento et, quidquid damnum inferre potest, si quis dixerit: " Hoc est! ", ad Deum utriusque causa perveniet, et, quem Deus condemnaverit, duplum restituet proximo suo.
EXOD|22|9|Si quis commendaverit proximo suo asinum, bovem, ovem vel omne iumentum ad custodiam, et mortuum fuerit aut fractum vel captum ab hostibus, nullusque hoc viderit,
EXOD|22|10|iusiurandum per Dominum erit in medio quod non extenderit manum ad rem proximi sui; suscipietque dominus iuramentum, et ille reddere non cogetur.
EXOD|22|11|Quod si furto ablatum fuerit, restituet damnum domino;
EXOD|22|12|si dilaceratum a bestia, deferat, quod occisum est, in testimonium et non restituet.
EXOD|22|13|Qui a proximo suo quidquam horum mutuo postulaverit, et fractum aut mortuum fuerit, domino non praesente, reddere compelletur.
EXOD|22|14|Quod si impraesentiarum dominus fuerit, non restituet. Si mercennarius est, venit in mercedem operis sui.
EXOD|22|15|Si seduxerit quis virginem necdum desponsatam dormieritque cum ea, pretio acquiret eam sibi uxorem.
EXOD|22|16|Si pater virginis eam dare noluerit, appendet ei pecuniam iuxta pretium pro virginibus dandum.
EXOD|22|17|Maleficam non patieris vivere.
EXOD|22|18|Qui coierit cum iumento, morte moriatur.
EXOD|22|19|Qui immolat diis, occidetur, praeter Domino soli.
EXOD|22|20|Advenam non opprimes neque affliges eum; advenae enim et ipsi fuistis in terra Aegypti.
EXOD|22|21|Viduae et pupillo non nocebitis.
EXOD|22|22|Si laeseritis eos, vociferabuntur ad me, et ego audiam clamorem eorum;
EXOD|22|23|et indignabitur furor meus, percutiamque vos gladio, et erunt uxores vestrae viduae et filii vestri pupilli.
EXOD|22|24|Si pecuniam mutuam dederis in populo meo pauperi, qui habitat tecum, non eris ei quasi creditor; non imponetis ei usuram.
EXOD|22|25|Si pignus a proximo tuo acceperis pallium, ante solis occasum reddes ei;
EXOD|22|26|ipsum enim est solum, quo operitur, indumentum carnis eius, nec habet aliud, in quo dormiat; si clamaverit ad me, exaudiam eum, quia misericors sum.
EXOD|22|27|Deo non detrahes et principi populi tui non maledices.
EXOD|22|28|Abundantiam areae tuae et torcularis tui non tardabis reddere.Primogenitum filiorum tuorum dabis mihi.
EXOD|22|29|De bobus quoque et ovibus similiter facies: septem diebus sit cum matre sua, die octavo reddes illum mihi.
EXOD|22|30|Viri sancti eritis mihi; carnem animalis in agro dilacerati non comedetis, sed proicietis canibus.
EXOD|23|1|Non suscipies famam falsam nec iunges manum tuam cum impio, ut dicas falsum testimonium.
EXOD|23|2|Non sequeris turbam ad faciendum malum; nec in iudicio plurimorum acquiesces sententiae, ut a vero devies.
EXOD|23|3|Pauperis quoque non misereberis in iudicio.
EXOD|23|4|Si occurreris bovi inimici tui aut asino erranti, reduc ad eum.
EXOD|23|5|Si videris asinum odientis te iacere sub onere suo, non pertransibis, sed sublevabis cum eo.
EXOD|23|6|Non pervertes iudicium pauperis in lite eius.
EXOD|23|7|Mendacium fugies. Insontem et iustum non occides, quia aversor impium.
EXOD|23|8|Nec accipies munera, quae excaecant etiam prudentes et subvertunt verba iustorum.
EXOD|23|9|Peregrinum non opprimes; scitis enim advenarum animas, quia et ipsi peregrini fuistis in terra Aegypti.
EXOD|23|10|Sex annis seminabis terram tuam et congregabis fruges eius.
EXOD|23|11|Anno autem septimo dimittes eam et requiescere facies, ut comedant pauperes populi tui; et quidquid reliquum fuerit, edant bestiae agri. Ita facies in vinea et in oliveto tuo.
EXOD|23|12|Sex diebus operaberis; septima die cessabis, ut requiescat bos et asinus tuus, et refrigeretur filius ancillae tuae et advena.
EXOD|23|13|Omnia, quae dixi vobis, custodite, et nomen externorum deorum non invocabitis, neque audietur ex ore tuo.
EXOD|23|14|Tribus vicibus per singulos annos mihi festa celebrabitis.
EXOD|23|15|Sollemnitatem Azymorum custodies: septem diebus comedes azyma, sicut praecepi tibi, tempore statuto mensis Abib, quando egressus es de Aegypto.Non apparebis in conspectu meo vacuus.
EXOD|23|16|Et sollemnitatem Messis primitivorum operis tui, quaecumque seminaveris in agro; sollemnitatem quoque Collectae in exitu anni, quando congregaveris omnes fruges tuas de agro.
EXOD|23|17|Ter in anno apparebit omne masculinum tuum coram Domino Deo.
EXOD|23|18|Non immolabis super fermento sanguinem victimae meae, nec remanebit adeps sollemnitatis meae usque mane.
EXOD|23|19|Primitias primarum frugum terrae tuae deferes in domum Domini Dei tui.Non coques haedum in lacte matris suae.
EXOD|23|20|Ecce ego mittam angelum, qui praecedat te et custodiat in via et introducat ad locum, quem paravi.
EXOD|23|21|Observa eum et audi vocem eius nec contemnendum putes; quia non dimittet, cum peccaveritis, quia est nomen meum in illo.
EXOD|23|22|Quod si audieris vocem eius et feceris omnia, quae loquor, inimicus ero inimicis tuis et affligam affligentes te.
EXOD|23|23|Praecedet enim te angelus meus et introducet te ad Amorraeum et Hetthaeum et Pherezaeum Chananaeumque et Hevaeum et Iebusaeum, quos ego conteram.
EXOD|23|24|Non adorabis deos eorum nec coles eos; non facies secundum opera eorum, sed destrues eos et confringes lapides eorum.
EXOD|23|25|Servietisque Domino Deo vestro, ut benedicam panibus tuis et aquis et auferam infirmitatem de medio tui.
EXOD|23|26|Non erit abortiens nec sterilis in terra tua; numerum dierum tuorum implebo.
EXOD|23|27|Terrorem meum mittam in praecursum tuum et perturbabo omnem populum, ad quem ingre dieris; cunctorumque inimicorum tuorum coram te terga vertam
EXOD|23|28|emittens crabrones prius, qui fugabunt Hevaeum et Chananaeum et Hetthaeum, antequam introeas.
EXOD|23|29|Non eiciam eos a facie tua anno uno, ne terra in solitudinem redigatur, et multiplicentur contra te bestiae agri.
EXOD|23|30|Paulatim expellam eos de conspectu tuo, donec augearis et possideas terram.
EXOD|23|31|Ponam autem terminos tuos a mari Rubro usque ad mare Palaestinorum et a deserto usque ad Fluvium. Tradam manibus vestris habitatores terrae et eiciam eos de conspectu vestro.
EXOD|23|32|Non inibis cum eis foedus nec cum diis eorum.
EXOD|23|33|Non habitent in terra tua, ne peccare te faciant in me, si servieris diis eorum; quod tibi certo erit in scandalum ".
EXOD|24|1|Moysi quoque dixit: " Ascende ad Dominum, tu et Aa ron, Nadab et Abiu et septuaginta senes ex Israel, et adorabitis procul.
EXOD|24|2|Solusque Moyses ascendet ad Dominum, et illi non appropinquabunt, nec populus ascendet cum eo ".
EXOD|24|3|Venit ergo Moyses et narravit plebi omnia verba Domini atque iudicia; responditque omnis populus una voce: " Omnia verba Domini, quae locutus est, faciemus ".
EXOD|24|4|Scripsit autem Moyses universos sermones Domini; et mane consurgens aedificavit altare ad radices montis et duodecim lapides per duodecim tribus Israel.
EXOD|24|5|Misitque iuvenes de filiis Israel, et obtulerunt holocausta; immolaveruntque victimas pacificas Domino vitulos.
EXOD|24|6|Tulit itaque Moyses dimidiam partem sanguinis et misit in crateras; partem autem residuam respersit super altare.
EXOD|24|7|Assumensque volumen foederis legit, audiente populo, qui dixerunt: " Omnia, quae locutus est Dominus, faciemus et erimus oboedientes ".
EXOD|24|8|Ille vero sumptum sanguinem respersit in populum et ait: " Hic est sanguis foederis, quod pepigit Dominus vobiscum super cunctis sermonibus his ".
EXOD|24|9|Ascenderuntque Moyses et Aaron, Nadab et Abiu et septuaginta de senioribus Israel.
EXOD|24|10|Et viderunt Deum Israel, et sub pedibus eius quasi opus lapidis sapphirini et quasi ipsum caelum, cum serenum est.
EXOD|24|11|Nec in electos filiorum Israel misit manum suam; videruntque Deum et comederunt ac biberunt.
EXOD|24|12|Dixit autem Dominus ad Moysen: " Ascende ad me in montem et esto ibi; daboque tibi tabulas lapideas et legem ac mandata, quae scripsi, ut doceas eos ".
EXOD|24|13|Surrexerunt Moyses et Iosue minister eius; ascendensque Moyses in montem Dei
EXOD|24|14|senioribus ait: " Exspectate hic, donec revertamur ad vos. Habetis Aaron et Hur vobiscum; si quid natum fuerit quaestionis, referetis ad eos ".
EXOD|24|15|Cumque ascendisset Moyses in montem, operuit nubes montem;
EXOD|24|16|et habitavit gloria Domini super Sinai tegens illum nube sex diebus; septimo autem die vocavit eum de medio caliginis.
EXOD|24|17|Erat autem species gloriae Domini quasi ignis ardens super verticem montis in conspectu filiorum Israel.
EXOD|24|18|Ingressusque Moyses medium nebulae ascendit in montem; et fuit ibi quadraginta diebus et quadraginta noctibus.
EXOD|25|1|Locutusque est Dominus ad Moysen dicens:
EXOD|25|2|" Loquere filiis Israel, ut tollant mihi donaria; ab omni homine, qui offert ultroneus, accipietis ea.
EXOD|25|3|Haec sunt autem, quae accipere debetis: aurum et argentum et aes,
EXOD|25|4|hyacinthum et purpuram coccumque et byssum, pilos caprarum
EXOD|25|5|et pelles arietum rubricatas pellesque delphini et ligna acaciae,
EXOD|25|6|oleum ad luminaria concinnanda, aromata in unguentum et in thymiama boni odoris,
EXOD|25|7|lapides onychinos et gemmas ad ornandum ephod ac pectorale.
EXOD|25|8|Facientque mihi sanctuarium, et habitabo in medio eorum.
EXOD|25|9|Iuxta omnem similitudinem habitaculi, quam ostendam tibi, et omnium vasorum in cultum eius: sicque facietis illud.
EXOD|25|10|Arcam de lignis acaciae compingent; cuius longitudo habeat duos semis cubitos, latitudo cubitum et dimidium, altitudo cubitum similiter ac semissem.
EXOD|25|11|Et deaurabis eam auro mundissimo intus et foris; faciesque supra coronam auream per circuitum
EXOD|25|12|et conflabis ei quattuor circulos aureos, quos pones in quattuor arcae pedibus: duo circuli sint in latere uno et duo in altero.
EXOD|25|13|Facies quoque vectes de lignis acaciae et operies eos auro;
EXOD|25|14|inducesque per circulos, qui sunt in arcae lateribus, ut portetur in eis;
EXOD|25|15|qui semper erunt in circulis nec umquam extrahentur ab eis.
EXOD|25|16|Ponesque in arcam testimonium, quod dabo tibi.
EXOD|25|17|Facies et propitiatorium de auro mundissimo; duos cubitos et dimidium tenebit longitudo eius, et cubitum ac semissem latitudo.
EXOD|25|18|Duos quoque cherubim aureos et productiles facies ex utraque parte propitiatorii,
EXOD|25|19|cherub unus sit in latere uno et alter in altero; ex propitiatorio facies cherubim in utraque parte eius.
EXOD|25|20|Expandent alas sursum et operient alis suis propitiatorium; respicientque se mutuo, versis vultibus in propitiatorium,
EXOD|25|21|quo operienda est arca, in qua pones testimonium, quod dabo tibi.
EXOD|25|22|Et conveniam te ibi et loquar ad te supra propitiatorium de medio duorum cherubim, qui erunt super arcam testimonii, cuncta, quae mandabo per te filiis Israel.
EXOD|25|23|Facies et mensam de lignis acaciae habentem duos cubitos longitudinis et in latitudine cubitum et in altitudine cubitum ac semissem.
EXOD|25|24|Et inaurabis eam auro purissimo; faciesque illi coronam auream per circuitum.
EXOD|25|25|Facies quoque ei limbum altum quattuor digitis per circuitum et super illum coronam auream.
EXOD|25|26|Quattuor quoque circulos aureos praeparabis et pones eos in quattuor angulis eiusdem mensae per singulos pedes.
EXOD|25|27|Iuxta limbum erunt circuli aurei, ut mittantur vectes per eos, et possit mensa portari.
EXOD|25|28|Ipsosque vectes facies de lignis acaciae et circumdabis auro, et per ipsos subvehitur mensa.
EXOD|25|29|Parabis et acetabula ac phialas, vasa et cyathos, in quibus offerenda sunt libamina, ex auro purissimo.
EXOD|25|30|Et pones super mensam panes propositionis in conspectu meo semper.
EXOD|25|31|Facies et candelabrum ductile de auro mundissimo: basis et hastile eius, scyphi et sphaerulae ac flores in unum efformentur.
EXOD|25|32|Sex calami egredientur de lateribus, tres ex uno latere et tres ex altero.
EXOD|25|33|Tres scyphi quasi in nucis modum in calamo uno sphaerulaeque simul et flores; et tres similiter scyphi instar nucis in calamo altero sphaerulaeque simul et flores: hoc erit opus sex calamorum, qui producendi sunt de hastili.
EXOD|25|34|In ipso autem hastili candelabri erunt quattuor scyphi in nucis modum sphaerulaeque et flores.
EXOD|25|35|Singulae sphaerulae sub binis calamis per tria loca, qui simul sex fiunt, procedentes de hastili uno.
EXOD|25|36|Sphaerulae igitur et calami unum cum ipso erunt, totum ductile de auro purissimo.
EXOD|25|37|Facies et lucernas septem et pones eas super candelabrum, ut luceant in locum ex adverso.
EXOD|25|38|Emunctoria quoque et vasa, in quibus emuncta condantur, fient de auro purissimo.
EXOD|25|39|Omne pondus candelabri cum universis vasis suis habebit talentum auri purissimi.
EXOD|25|40|Inspice et fac secundum exemplar, quod tibi in monte monstratum est.
EXOD|26|1|Habitaculum vero ita facies: decem cortinas de bysso re torta et hyacintho ac purpura coccoque cum cherubim opere polymito facies.
EXOD|26|2|Longitudo cortinae unius habebit viginti octo cubitos, latitudo quattuor cubitorum erit. Unius mensurae fient universae cortinae.
EXOD|26|3|Quinque cortinae sibi iungentur mutuo, et aliae quinque nexu simili cohaerebunt.
EXOD|26|4|Ansulas hyacinthinas in latere facies cortinae unius in extremitate iuncturae et similiter facies in latere cortinae extremae in iunctura altera.
EXOD|26|5|Quinquaginta ansulas facies in cortina una et quinquaginta ansulas facies in summitate cortinae, quae est in iunctura altera, ita insertas, ut ansa contra ansam veniat.
EXOD|26|6|Facies et quinquaginta fibulas aureas, quibus cortinarum vela iungenda sunt, ut unum habitaculum fiat.
EXOD|26|7|Facies et saga cilicina undecim pro tabernaculo super habitaculum.
EXOD|26|8|Longitudo sagi unius habebit triginta cubitos et latitudo quattuor; aequa erit mensura sagorum omnium.
EXOD|26|9|E quibus quinque iunges seorsum et sex sibi mutuo copulabis, ita ut sextum sagum in fronte tecti duplices.
EXOD|26|10|Facies et quinquaginta ansas in ora sagi ultimi iuncturae unius et quinquaginta ansas in ora sagi iuncturae alterius.
EXOD|26|11|Facies et quinquaginta fibulas aeneas, quibus iungantur ansae, ut unum ex omnibus tabernaculum fiat.
EXOD|26|12|Quod autem superfuerit in sagis, quae parantur tecto, id est unum sagum, quod amplius est, ex medietate eius operies posteriora habitaculi;
EXOD|26|13|et cubitus ex una parte pendebit, et alter ex altera, qui plus est in longitudine sagorum tabernaculi utrumque latus habitaculi protegens.
EXOD|26|14|Facies et operimentum aliud pro tabernaculo de pellibus arietum rubricatis et super hoc rursum aliud operimentum de pellibus delphini.
EXOD|26|15|Facies et tabulas stantes habitaculi de lignis acaciae,
EXOD|26|16|quae singulae denos cubitos in longitudine habeant et in latitudine singulos ac semissem.
EXOD|26|17|In tabula una duo pedes fient, quibus tabula alteri tabulae conectatur; atque in hunc modum cunctae tabulae habitaculi parabuntur.
EXOD|26|18|Quarum viginti erunt in latere meridiano, quod vergit ad austrum;
EXOD|26|19|quibus quadraginta bases argenteas fundes, ut binae bases singulis pedibus singularum tabularum subiciantur.
EXOD|26|20|In latere quoque secundo habitaculi, quod vergit ad aquilonem, viginti tabulae erunt,
EXOD|26|21|quadraginta habentes bases argenteas; binae bases singulis tabulis supponentur.
EXOD|26|22|Ad occidentalem vero plagam in tergo habitaculi facies sex tabulas;
EXOD|26|23|et rursum alias duas, quae in angulis erigantur, post tergum habitaculi.
EXOD|26|24|Eruntque geminae a deorsum usque sursum in compaginem unam; ita erit duabus istis, pro duabus angulis erunt.
EXOD|26|25|Et erunt simul tabulae octo, bases earum argenteae sedecim, duabus basibus per unam tabulam supputatis.
EXOD|26|26|Facies et vectes de lignis acaciae, quinque ad continendas tabulas in uno latere habitaculi
EXOD|26|27|et quinque alios in altero et eiusdem numeri in tergo ad occidentalem plagam;
EXOD|26|28|vectis autem medius transibit per medias tabulas a summo usque ad summum.
EXOD|26|29|Ipsasque tabulas deaurabis et fundes eis anulos aureos, per quos vectes tabulata contineant, quos operies laminis aureis.
EXOD|26|30|Et eriges habitaculum iuxta exemplar, quod tibi in monte monstratum est.
EXOD|26|31|Facies et velum de hyacintho et purpura coccoque et bysso retorta, opere polymito, cum cherubim intextis.
EXOD|26|32|Quod appendes in quattuor columnis de lignis acaciae, quae ipsae quidem deauratae erunt et habebunt uncos aureos, sed bases argenteas.
EXOD|26|33|Inseres autem velum subter fibulas, intra quod pones arcam testimonii et quo sanctum et sanctum sanctorum dividentur.
EXOD|26|34|Pones et propitiatorium super arcam testimonii in sancto sanctorum
EXOD|26|35|mensamque extra velum et contra mensam candelabrum in latere habitaculi meridiano; mensa enim stabit in parte aquilonis.
EXOD|26|36|Facies et velum in introitu tabernaculi de hyacintho et purpura coccoque et bysso retorta opere plumarii.
EXOD|26|37|Et quinque columnas deaurabis lignorum acaciae, ante quas ducetur velum, quarum erunt unci aurei et bases aeneae.
EXOD|27|1|Facies et altare de lignis acaciae, quod habebit quinque cubitos in longitudine et totidem in latitudine, id est quadrum, et tres cubitos in altitudine.
EXOD|27|2|Cornua autem per quattuor angulos ex ipso erunt, et operies illud aere.
EXOD|27|3|Faciesque in usus eius lebetes ad suscipiendos cineres et vatilla et pateras atque fuscinulas et ignium receptacula; omnia vasa ex aere fabricabis.
EXOD|27|4|Craticulamque facies ei in modum retis aeneam, per cuius quattuor angulos erunt quattuor anuli aenei,
EXOD|27|5|et pones eam subter marginem altaris; eritque craticula usque ad altaris medium.
EXOD|27|6|Facies et vectes altaris de lignis acaciae duos, quos operies laminis aeneis,
EXOD|27|7|et induces per anulos; eruntque ex utroque latere altaris ad portandum.
EXOD|27|8|Cavum ex tabulis facies illud; sicut tibi in monte monstratum est, sic facient.
EXOD|27|9|Facies et atrium habitaculi, in cuius plaga australi contra meridiem erunt tentoria de bysso retorta: centum cubitos unum latus tenebit in longitudine
EXOD|27|10|et columnas viginti et bases totidem aeneas et uncos columnarum anulosque earum argenteos.
EXOD|27|11|Similiter in latere aquilonis: per longum erunt tentoria centum cubitorum, columnae viginti et bases aeneae eiusdem numeri et unci columnarum anulique earum argentei.
EXOD|27|12|In latitudine vero atrii, quae respicit ad occidentem, erunt tentoria per quinquaginta cubitos et columnae decem basesque totidem.
EXOD|27|13|In ea quoque atrii latitudine, quae respicit ad orientem, quinquaginta cubiti erunt,
EXOD|27|14|in quibus quindecim cubitorum tentoria lateri uno deputabuntur columnaeque tres et bases totidem;
EXOD|27|15|et in latere altero erunt tentoria, cubitos obtinentia quindecim, columnae tres et bases totidem.
EXOD|27|16|In introitu vero atrii fiet velum cubitorum viginti, ex hyacintho et purpura coccoque et bysso retorta opere plumarii; columnas habebit quattuor cum basibus totidem.
EXOD|27|17|Omnes columnae atrii per circuitum cinctae erunt anulis argenteis, et unci earum erunt argentei et bases aeneae.
EXOD|27|18|In longitudine occupabit atrium cubitos centum, in latitudine quinquaginta, altitudo quinque cubitorum erit; fietque de bysso retorta, et habebit bases aeneas.
EXOD|27|19|Cuncta vasa habitaculi in omnes usus eius et omnes paxillos eius et omnes paxillos atrii ex aere facies.
EXOD|27|20|Praecipe filiis Israel, ut afferant tibi oleum de arboribus olivarum purissimum piloque contusum, ut ardeat lucerna semper
EXOD|27|21|in tabernaculo conventus, extra velum, quod oppansum est testimonio. Et parabunt eam Aaron et filii eius, ut a vespere usque mane luceat coram Domino. Perpetuus erit cultus per successiones eorum a filiis Israel.
EXOD|28|1|Applica quoque ad te Aaron fratrem tuum cum filiis suis de medio filiorum Israel, ut sacerdotio fungantur mihi: Aaron, Nadab et Abiu, Eleazar et Ithamar.
EXOD|28|2|Faciesque vestes sanctas Aaron fratri tuo in gloriam et decorem;
EXOD|28|3|et loqueris cunctis sapientibus corde, quos replevi spiritu prudentiae, ut faciant vestes Aaron, in quibus sanctificatus ministret mihi.
EXOD|28|4|Haec autem erunt vestimenta, quae facient: pectorale et ephod, tunicam et subuculam textam, tiaram et balteum. Facient vestimenta sancta Aaron fratri tuo et filiis eius, ut sacerdotio fungantur mihi;
EXOD|28|5|accipientque aurum et hyacinthum et purpuram coccumque et byssum.
EXOD|28|6|Facient autem ephod de auro et hyacintho ac purpura coccoque bysso retorta opere polymito.
EXOD|28|7|Duas fascias umerales habebit et in utroque latere summitatum suarum copulabitur cum eis.
EXOD|28|8|Et balteus super ephod ad constringendum, eiusdem operis et unum cum eo, erit ex auro et hyacintho et purpura coccoque et bysso retorta.
EXOD|28|9|Sumesque duos lapides onychinos et sculpes in eis nomina filiorum Israel:
EXOD|28|10|sex nomina in lapide uno et sex reliqua in altero, iuxta ordinem nativitatis eorum.
EXOD|28|11|Opere sculptoris et caelatura gemmarii sculpes eos nominibus filiorum Israel, inclusos textura aurea;
EXOD|28|12|et pones duos lapides super fascias umerales ephod, lapides memorialis filiorum Israel. Portabitque Aaron nomina eorum coram Domino super utrumque umerum ob recordationem.
EXOD|28|13|Facies ergo margines textas ex auro
EXOD|28|14|et duas catenulas ex auro purissimo quasi funiculos opus tortile et inseres catenulas tortas marginibus.
EXOD|28|15|Pectorale quoque iudicii facies opere polymito, iuxta texturam ephod, ex auro, hyacintho et purpura coccoque et bysso retorta.
EXOD|28|16|Quadrangulum erit et duplex; mensuram palmi habebit tam in longitudine quam in latitudine.
EXOD|28|17|Ponesque in eo quattuor ordines lapidum: in primo versu erit lapis sardius et topazius et smaragdus;
EXOD|28|18|in secundo carbunculus, sapphirus et iaspis;
EXOD|28|19|in tertio hyacinthus, achates et amethystus;
EXOD|28|20|in quarto chrysolithus, onychinus et beryllus. Inclusi auro erunt per ordines suos.
EXOD|28|21|Habebuntque nomina filiorum Israel: duodecim nominibus caelabuntur, singuli lapides nominibus singulorum per duodecim tribus.
EXOD|28|22|Facies in pectorali catenas quasi funiculos, opus tortile, ex auro purissimo;
EXOD|28|23|et duos anulos aureos, quos pones in utraque pectoralis summitate;
EXOD|28|24|catenasque aureas iunges anulis, qui sunt in marginalibus eius;
EXOD|28|25|et ipsarum catenarum extrema duobus copulabis marginibus in fasciis umeralibus ephod in parte eius anteriore.
EXOD|28|26|Facies et duos anulos aureos, quos pones in summitatibus pectoralis in ora interiore, quae respicit ephod.
EXOD|28|27|Necnon et alios duos anulos aureos, qui ponendi sunt in utraque fascia umerali ephod deorsum, versus partem anteriorem eius iuxta iuncturam eius supra balteum ephod,
EXOD|28|28|et stringatur pectorale anulis suis cum anulis ephod vitta hyacinthina, ut maneat supra balteum ephod, et a se invicem pectorale et ephod nequeant separari.
EXOD|28|29|Portabitque Aaron nomina filiorum Israel in pectorali iudicii super cor suum, quando ingredietur sanctuarium: memoriale coram Domino in aeternum.
EXOD|28|30|Pones autem in pectorali iudicii Urim et Tummim, quae erunt super cor Aaron, quando ingredietur coram Domino; et gestabit iudicium filiorum Israel super cor suum in conspectu Domini semper.
EXOD|28|31|Facies et pallium ephod totum hyacinthinum,
EXOD|28|32|in cuius medio supra erit capitium et ora per gyrum eius textilis, sicut in capitio loricae, ne rumpatur.
EXOD|28|33|Deorsum vero, ad pedes eiusdem pallii per circuitum, quasi mala punica facies ex hyacintho et purpura et cocco, mixtis in medio tintinnabulis aureis;
EXOD|28|34|ita ut sit tintinnabulum aureum inter singula mala punica.
EXOD|28|35|Et vestietur eo Aaron in officio ministerii, ut audiatur sonitus, quando ingreditur et egreditur sanctuarium in conspectu Domini, et non moriatur.
EXOD|28|36|Facies et laminam de auro purissimo, in qua sculpes opere caelatoris: "Sanctum Domino".
EXOD|28|37|Ligabisque eam vitta hyacinthina, et erit super tiaram
EXOD|28|38|super frontem Aaron. Portabitque Aaron iniquitatem contra sancta, quae sanctificabunt filii Israel in cunctis muneribus et donariis suis. Eritque lamina semper in fronte eius, ut placatus eis sit Dominus.
EXOD|28|39|Texesque tunicam bysso et tiaram byssinam facies et balteum opere plumarii.
EXOD|28|40|Porro filiis Aaron tunicas lineas parabis et balteos ac mitras in gloriam et decorem;
EXOD|28|41|vestiesque his omnibus Aaron fratrem tuum et filios eius cum eo. Et unges eos et implebis manus eorum sanctificabisque illos, ut sacerdotio fungantur mihi.
EXOD|28|42|Facies eis et feminalia linea, ut operiant carnem turpitudinis suae a renibus usque ad femora;
EXOD|28|43|et utentur eis Aaron et filii eius, quando ingredientur tabernaculum conventus, vel quando appropinquant ad altare, ut ministrent in sanctuario, ne iniquitatis rei moriantur: legitimum sempiternum erit Aaron et semini eius post eum.
EXOD|29|1|Sed et hoc facies eis, ut mihi in sacerdotio consecrentur: tolle vitulum unum de armento et arietes duos immaculatos
EXOD|29|2|panesque azymos et crustulas absque fermento, quae conspersa sint oleo, lagana quoque azyma oleo lita; de simila triticea cuncta facies
EXOD|29|3|et posita in canistro offeres, vitulum quoque et duos arietes.
EXOD|29|4|Aaron ac filios eius applicabis ad ostium tabernaculi conventus. Cumque laveris patrem cum filiis suis aqua,
EXOD|29|5|indues Aaron vestimentis suis, id est subucula et tunica ephod et ephod et pectorali, quod constringes ei cingulo ephod;
EXOD|29|6|et pones tiaram in capite eius et diadema sanctum super tiaram
EXOD|29|7|et oleum unctionis fundes super caput eius; atque hoc ritu consecrabitur.
EXOD|29|8|Filios quoque illius applicabis et indues tunicis lineis cingesque balteo
EXOD|29|9|et impones eis mitras; eruntque sacerdotes mihi iure perpetuo.Postquam impleveris manus Aaron et filiorum eius,
EXOD|29|10|applicabis et vitulum coram tabernaculo conventus; imponentque Aaron et filii eius manus super caput illius,
EXOD|29|11|et mactabis eum in conspectu Domini, iuxta ostium tabernaculi conventus.
EXOD|29|12|Sumptumque de sanguine vituli, pones super cornua altaris digito tuo, reliquum autem sanguinem fundes iuxta basim eius.
EXOD|29|13|Sumes et adipem totum, qui operit intestina, et reticulum iecoris ac duos renes et adipem, qui super eos est, et offeres comburens super altare;
EXOD|29|14|carnes vero vituli et corium et fimum combures foris extra castra, eo quod pro peccato sit.
EXOD|29|15|Unum quoque arietem sumes, super cuius caput ponent Aaron et filii eius manus;
EXOD|29|16|quem cum mactaveris, tolles sanguinem eius et fundes super altare per circuitum.
EXOD|29|17|Ipsum autem arietem secabis in frusta lotaque intestina eius ac pedes pones super concisas carnes et super caput illius.
EXOD|29|18|Et adolebis totum arietem super altare: holocaustum est Domino, odor suavissimus, incensum est Domino.
EXOD|29|19|Tolles quoque arietem alterum, super cuius caput Aaron et filii eius ponent manus;
EXOD|29|20|quem cum immolaveris, sumes de sanguine ipsius et pones super extremum auriculae dextrae Aaron et filiorum eius et super pollices manus eorum ac pedis dextri; fundesque sanguinem super altare per circuitum.
EXOD|29|21|Cumque tuleris de sanguine, qui est super altare, et de oleo unctionis, asperges Aaron et vestes eius, filios et vestimenta eorum cum ipso. Et sanctus erit ipse et vestimenta eius et filii eius et vestimenta eorum cum ipso.
EXOD|29|22|Tollesque adipem de ariete et caudam et arvinam, quae operit intestina, ac reticulum iecoris et duos renes atque adipem, qui super eos est, armumque dextrum, eo quod sit aries consecrationis,
EXOD|29|23|tortamque panis unam, crustulam unam conspersam oleo, laganum unum de canistro azymorum, quod positum est in conspectu Domini;
EXOD|29|24|ponesque omnia super manus Aaron et filiorum eius, ut agitent ea coram Domino.
EXOD|29|25|Suscipiesque universa de manibus eorum et incendes in altari super holocausto in odorem suavissimum in conspectu Domini; quia incensum est Domino.
EXOD|29|26|Sumes quoque pectusculum de ariete, quo initiatus est Aaron, elevabisque illud coram Domino; et cedet in partem tuam.
EXOD|29|27|Sanctificabisque pectusculum elevatum et armum oblatum, quem de ariete separasti,
EXOD|29|28|quo initiatus est Aaron et filii eius; cedentque in partem Aaron et filiorum eius iure perpetuo a filiis Israel; quia oblatio est et oblatio erit a filiis Israel de victimis eorum pacificis, oblatio eorum Domino.
EXOD|29|29|Vestem autem sanctam, qua utetur Aaron, habebunt filii eius post eum, ut ungantur in ea, et impleantur in ea manus eorum.
EXOD|29|30|Septem diebus utetur illa, qui pontifex pro eo fuerit constitutus de filiis eius, qui ingredietur tabernaculum conventus, ut ministret in sanctuario.
EXOD|29|31|Arietem autem consecrationis tolles et coques carnes eius in loco sancto.
EXOD|29|32|Et vescetur Aaron et filii eius carnibus arietis et panibus, qui sunt in canistro, in vestibulo tabernaculi conventus.
EXOD|29|33|Et comedent ea, quibus expiatio facta fuerit ad implendum manus eorum, ad sanctificandum eos. Alienigena non vescetur ex eis, quia sancta sunt.
EXOD|29|34|Quod si remanserit de carnibus consecrationis sive de panibus usque mane, combures reliquias igni; non comedentur, quia sancta sunt.
EXOD|29|35|Omnia, quae praecepi tibi, facies super Aaron et filiis eius. Septem diebus consecrabis manus eorum
EXOD|29|36|et vitulum pro peccato offeres per singulos dies ad expiandum. Mundabisque altare expians illud et unges illud in sanctificationem.
EXOD|29|37|Septem diebus expiabis altare et sanctificabis; et erit sanctum sanctorum: omnis, qui tetigerit illud, sanctificabitur.
EXOD|29|38|Hoc est quod facies in altari: agnos anniculos duos per singulos dies iugiter,
EXOD|29|39|unum agnum mane et alterum vespere;
EXOD|29|40|decimam partem similae conspersae oleo tunso, quod habeat mensuram quartam partem hin, et vinum ad libandum eiusdem mensurae in agno uno.
EXOD|29|41|Alterum vero agnum offeres ad vesperam iuxta ritum matutinae oblationis et libationis in odorem suavitatis, incensum Domino,
EXOD|29|42|holocaustum perpetuum in generationes vestras, ad ostium tabernaculi conventus coram Domino, ubi conveniam vos, ut loquar ad te.
EXOD|29|43|Ibi conveniam filios Israel, et sanctificabitur locus in gloria mea.
EXOD|29|44|Sanctificabo et tabernaculum conventus cum altari et Aaron cum filiis eius, ut sacerdotio fungantur mihi.
EXOD|29|45|Et habitabo in medio filiorum Israel eroque eis Deus;
EXOD|29|46|et scient quia ego Dominus Deus eorum, qui eduxi eos de terra Aegypti, ut manerem inter illos: ego Dominus Deus ipsorum.
EXOD|30|1|Facies quoque altare ad adolendum thymiama de lignis acaciae
EXOD|30|2|habens cubitum longitudinis et alterum latitudinis, id est quadrangulum, et duos cubitos in altitudine; cornua ex ipso procedent.
EXOD|30|3|Vestiesque illud auro purissimo, tam craticulam eius quam parietes per circuitum et cornua. Faciesque ei coronam aureolam per gyrum
EXOD|30|4|et duos anulos aureos sub corona in duobus lateribus, ut mittantur in eos vectes, et altare portetur.
EXOD|30|5|Ipsos quoque vectes facies de lignis acaciae et inaurabis.
EXOD|30|6|Ponesque altare contra velum, quod ante arcam pendet testimonii, coram propitiatorio, quo tegitur testimonium, ubi conveniam ad te.
EXOD|30|7|Et adolebit incensum super eo Aaron suave fragrans mane. Quando componet lucernas, incendet illud;
EXOD|30|8|et quando collocabit eas ad vesperum, uret thymiama sempiternum coram Domino in generationes vestras.
EXOD|30|9|Non offeretis super eo thymiama compositionis alterius nec holocaustum nec oblationem, nec libabitis libamina.
EXOD|30|10|Et expiabit Aaron super cornua eius semel per annum in sanguine sacrificii pro peccato; et placabit super eo in generationibus vestris: sanctum sanctorum erit Domino ".
EXOD|30|11|Locutusque est Dominus ad Moysen dicens:
EXOD|30|12|" Quando tuleris summam filiorum Israel iuxta numerum, dabunt singuli pretium expiationis pro animabus suis Domino; et non erit plaga in eis, cum fuerint recensiti.
EXOD|30|13|Hoc autem dabit omnis, qui transit ad censum, dimidium sicli iuxta mensuram sanctuarii ­ siclus viginti obolos habet ­; media pars sicli offeretur Domino.
EXOD|30|14|Qui habetur in numero a viginti annis et supra, dabit pretium;
EXOD|30|15|dives non addet ad medium sicli, et pauper nihil minuet, quando dabitis oblationem Domino in expiationem animarum vestrarum.
EXOD|30|16|Susceptamque expiationis pecuniam, quae collata est a filiis Israel, trades in usus tabernaculi conventus, ut sit monumentum eorum coram Domino et propitietur animabus illorum ".
EXOD|30|17|Locutusque est Dominus ad Moysen dicens:
EXOD|30|18|" Facies et labrum aeneum cum basi aenea ad lavandum; ponesque illud inter tabernaculum conventus et altare. Et, missa aqua,
EXOD|30|19|lavabunt in eo Aaron et filii eius manus suas ac pedes.
EXOD|30|20|Quando ingressuri sunt tabernaculum conventus, lavabunt se aqua, ne moriantur; vel quando accessuri sunt ad altare, ut ministrent, ut adoleant victimam Domino.
EXOD|30|21|Et lavabunt manus et pedes, ne moriantur: legitimum sempiternum erit, ipsi et semini eius per successiones ".
EXOD|30|22|Locutusque est Dominus ad Moysen
EXOD|30|23|dicens: " Sume tibi aromata prima myrrhae electae quingentos siclos et cinnamomi boni odoris medium, id est ducentos quinquaginta siclos, calami suave olentis similiter ducentos quinquaginta,
EXOD|30|24|casiae autem quingentos siclos, in pondere sanctuarii, olei de olivetis mensuram hin.
EXOD|30|25|Faciesque unctionis oleum sanctum, unguentum compositum opere unguentarii; unctionis oleum sanctum erit.
EXOD|30|26|Et unges ex eo tabernaculum conventus et arcam testamenti
EXOD|30|27|mensamque cum vasis suis, candelabrum et utensilia eius, altaria thymiamatis
EXOD|30|28|et holocausti et universam supellectilem, quae ad cultum eorum pertinet, et labrum cum basi sua.
EXOD|30|29|Sanctificabisque omnia, et erunt sancta sanctorum: qui tetigerit ea, sanctificabitur.
EXOD|30|30|Aaron et filios eius unges sanctificabisque eos, ut sacerdotio fungantur mihi.
EXOD|30|31|Filiis quoque Israel dices: Hoc oleum unctionis sanctum erit mihi in generationes vestras.
EXOD|30|32|Caro hominis non ungetur ex eo, et iuxta compositionem eius non facietis aliud, quia sanctum est et sanctum erit vobis.
EXOD|30|33|Homo quicumque tale composuerit et dederit ex eo super alienum, exterminabitur de populo suo ".
EXOD|30|34|Dixitque Dominus ad Moysen: " Sume tibi aromata, stacten et onycha, galbanum boni odoris et tus lucidissimum; aequalis ponderis erunt omnia.
EXOD|30|35|Faciesque thymiama compositum opere unguentarii, sale conditum et purum et sanctum.
EXOD|30|36|Cumque in tenuissimum pulverem ex parte contuderis, pones ex eo coram testimonio in tabernaculo conventus, in quo conveniam ad te: sanctum sanctorum erit vobis thymiama.
EXOD|30|37|Talem compositionem non facietis in usus vestros, quia tibi sanctum erit pro Domino;
EXOD|30|38|homo quicumque fecerit simile, ut odore illius perfruatur, peribit de populis suis ".
EXOD|31|1|Locutusque est Dominus ad Moysen dicens:
EXOD|31|2|" Ecce voca vi ex nomine Beseleel filium Uri filii Hur de tribu Iudae
EXOD|31|3|et implevi eum spiritu Dei, sapientia et intellegentia et scientia in omni opere
EXOD|31|4|ad excogitandum, quidquid fabrefieri potest ex auro et argento et aere,
EXOD|31|5|ad scindendum et includendum gemmas et ad sculpendum ligna, ad faciendum omne opus;
EXOD|31|6|dedique ei socium Ooliab filium Achisamech de tribu Dan et in corde omnis eruditi posui sapientiam, ut faciant cuncta, quae praecepi tibi:
EXOD|31|7|tabernaculum conventus et arcam testimonii et propitiatorium, quod super eam est, et cuncta vasa tabernaculi
EXOD|31|8|mensamque et vasa eius, candelabrum purissimum cum vasis suis et altaria thymiamatis
EXOD|31|9|et holocausti et omnia vasa eorum, labrum cum basi sua
EXOD|31|10|et vestes textas et vestes sanctas Aaron sacerdoti et vestes filiorum eius, ut fungantur officio suo in sacris,
EXOD|31|11|oleum unctionis et thymiama aromatum in sanctuario: omnia, quae praecepi tibi, facient ".
EXOD|31|12|Et locutus est Dominus ad Moysen dicens:
EXOD|31|13|" Loquere filiis Israel et dices ad eos: Videte ut sabbatum meum custodiatis, quia signum est inter me et vos in generationibus vestris, ut sciatis quia ego Dominus, qui sanctifico vos.
EXOD|31|14|Custodite sabbatum, sanctum est enim vobis. Qui polluerit illud, morte morietur; qui fecerit in eo opus, peribit anima illius de medio populi sui.
EXOD|31|15|Sex diebus facietis opus; in die septimo sabbatum est, requies sancta Domino: omnis, qui fecerit opus in hac die, morietur.
EXOD|31|16|Custodiant filii Israel sabbatum et celebrent illud in generationibus suis: pactum est sempiternum
EXOD|31|17|inter me et filios Israel signumque perpetuum; sex enim diebus fecit Dominus caelum et terram et in septimo ab opere cessavit et respiravit ".
EXOD|31|18|Deditque Dominus Moysi, completis huiuscemodi sermonibus in monte Sinai, duas tabulas testimonii lapideas scriptas digito Dei.
EXOD|32|1|Videns autem populus quod moram faceret descendendi de monte Moyses, congregatus ad Aaron dixit: " Surge, fac nobis deos, qui nos praecedant; Moysi enim, huic viro, qui nos eduxit de terra Aegypti, ignoramus quid acciderit ".
EXOD|32|2|Dixitque ad eos Aaron: " Tollite inaures aureas de uxorum filiorumque et filiarum vestrarum auribus et afferte ad me ".
EXOD|32|3|Fecitque omnis populus, quae iusserat, deferens inaures ad Aaron.
EXOD|32|4|Quas cum ille accepisset, formavit stilo imaginem et fecit ex eis vitulum conflatilem. Dixeruntque: " Hi sunt dii tui, Israel, qui te eduxerunt de terra Aegypti! ".
EXOD|32|5|Quod cum vidisset Aaron, aedificavit altare coram eo et praeconis voce clamavit dicens: " Cras sollemnitas Domini est ".
EXOD|32|6|Surgen tesque mane altero die obtulerunt holocausta et hostias pacificas; et sedit populus manducare et bibere et surrexerunt ludere.
EXOD|32|7|Locutus est autem Dominus ad Moysen: " Vade, descende; peccavit populus tuus, quem eduxisti de terra Aegypti.
EXOD|32|8|Recesserunt cito de via, quam praecepi eis, feceruntque sibi vitulum conflatilem et adoraverunt atque immolantes ei hostias dixerunt: "Isti sunt dii tui, Israel, qui te eduxerunt de terra Aegypti!" ".
EXOD|32|9|Rursumque ait Dominus ad Moysen: " Cerno quod populus iste durae cervicis sit;
EXOD|32|10|dimitte me, ut irascatur furor meus contra eos et deleam eos faciamque te in gentem magnam ".
EXOD|32|11|Moyses autem orabat Dominum Deum suum dicens: " Cur, Domine, irascitur furor tuus contra populum tuum, quem eduxisti de terra Aegypti in fortitudine magna et in manu robusta?
EXOD|32|12|Ne, quaeso, dicant Aegyptii: "Callide eduxit eos, ut interficeret in montibus et deleret e terra". Quiescat ira tua, et esto placabilis super nequitia populi tui.
EXOD|32|13|Recordare Abraham, Isaac et Israel servorum tuorum, quibus iurasti per temetipsum dicens: "Multiplicabo semen vestrum sicut stellas caeli; et universam terram hanc, de qua locutus sum, dabo semini vestro, et possidebitis eam semper" ".
EXOD|32|14|Placatusque est Dominus, ne faceret malum, quod locutus fuerat adversus populum suum.
EXOD|32|15|Et reversus est Moyses de monte portans duas tabulas testimonii in manu sua scriptas ex utraque parte
EXOD|32|16|et factas opere Dei; scriptura quoque Dei erat sculpta in tabulis.
EXOD|32|17|Audiens autem Iosue tumultum populi vociferantis dixit ad Moysen: " Ululatus pugnae auditur in castris ".
EXOD|32|18|Qui respondit:" Non est clamor vincentiumneque clamor fugientium,sed clamorem cantantiumego audio ".
EXOD|32|19|Cumque appropinquasset ad castra, vidit vitulum et choros; iratusque valde proiecit de manu tabulas et confregit eas ad radices montis.
EXOD|32|20|Arripiensque vitulum, quem fecerant, combussit et contrivit usque ad pulverem, quem sparsit in aquam et dedit ex eo potum filiis Israel.
EXOD|32|21|Dixitque ad Aaron: " Quid tibi fecit hic populus, ut induceres super eum peccatum maximum? ".
EXOD|32|22|Cui ille respondit: " Ne indignetur dominus meus; tu enim nosti populum istum, quod pronus sit ad malum.
EXOD|32|23|Dixerunt mihi: "Fac nobis deos, qui nos praecedant; huic enim Moysi, qui nos eduxit de terra Aegypti, nescimus quid acciderit".
EXOD|32|24|Quibus ego dixi: Quis vestrum habet aurum? Abstulerunt et dederunt mihi, et proieci illud in ignem; egressusque est hic vitulus ".
EXOD|32|25|Vidit ergo Moyses populum quod esset effrenatus; relaxaverat enim ei Aaron frenum in ludibrium hostium eorum.
EXOD|32|26|Et stans in porta castrorum ait: " Si quis est Domini, iungatur mihi! ". Congregatique sunt ad eum omnes filii Levi.
EXOD|32|27|Quibus ait: " Haec dicit Dominus, Deus Israel: Ponat unusquisque gladium super femur suum. Ite et redite de porta usque ad portam per medium castrorum, et occidat unusquisque fratrem et amicum et proximum suum ".
EXOD|32|28|Fecerunt filii Levi iuxta sermonem Moysi; cecideruntque de populo in die illa quasi tria milia hominum.
EXOD|32|29|Et ait Moyses: " Implestis manus vestras hodie Domino unusquisque in filio et in fratre suo, ut detur vobis benedictio ".
EXOD|32|30|Facto autem altero die, locutus est Moyses ad populum: " Peccastis peccatum maximum; ascendam ad Dominum, si quo modo quivero eum deprecari pro scelere vestro ".
EXOD|32|31|Reversusque ad Dominum ait: " Obsecro, peccavit populus iste peccatum maximum, feceruntque sibi deos aureos; aut dimitte eis hanc noxam
EXOD|32|32|aut, si non facis, dele me de libro tuo, quem scripsisti ".
EXOD|32|33|Cui respondit Dominus: " Qui peccaverit mihi, delebo eum de libro meo.
EXOD|32|34|Tu autem vade et duc populum istum, quo locutus sum tibi: angelus meus praecedet te; ego autem in die ultionis visitabo et hoc peccatum eorum ".
EXOD|32|35|Percussit ergo Dominus populum pro reatu vituli, quem fecerat Aaron.
EXOD|33|1|Locutusque est Dominus ad Moysen: " Vade, ascende de loco isto, tu et populus tuus, quem eduxisti de terra Aegypti, in terram, quam iuravi Abraham, Isaac et Iacob dicens: Semini tuo dabo eam.
EXOD|33|2|Et mittam praecursorem tui angelum et eiciam Chananaeum et Amorraeum et Hetthaeum et Pherezaeum et Hevaeum et Iebusaeum,
EXOD|33|3|et intres in terram fluentem lacte et melle. Non enim ascendam tecum, quia populus durae cervicis es, ne forte disperdam te in via ".
EXOD|33|4|Audiens populus sermonem hunc pessimum luxit, et nullus ex more indutus est cultu suo.
EXOD|33|5|Dixitque Dominus ad Moysen: " Loquere filiis Israel: Populus durae cervicis es; uno momento, si ascendam in medio tui, delebo te. Nunc autem depone ornatum tuum, ut sciam quid faciam tibi ".
EXOD|33|6|Deposuerunt ergo filii Israel ornatum suum a monte Horeb.
EXOD|33|7|Moyses autem tollens tabernaculum tetendit ei extra castra procul; vocavitque nomen eius Tabernaculum conventus. Et omnis, qui quaerebat Dominum, egrediebatur ad tabernaculum conventus extra castra.
EXOD|33|8|Cumque egrederetur Moyses ad tabernaculum, surgebat universa plebs, et stabat unusquisque in ostio papilionis sui; aspiciebantque tergum Moysi, donec ingrederetur tabernaculum.
EXOD|33|9|Ingresso autem illo tabernaculum, descendebat columna nubis et stabat ad ostium; loquebaturque cum Moyse,
EXOD|33|10|cernentibus universis quod columna nubis staret ad ostium tabernaculi. Stabantque ipsi et adorabant per fores tabernaculorum suorum.
EXOD|33|11|Loquebatur autem Dominus ad Moysen facie ad faciem, sicut solet loqui homo ad amicum suum. Cumque ille reverteretur in castra, minister eius Iosue filius Nun puer non recedebat de medio tabernaculi.
EXOD|33|12|Dixit autem Moyses ad Dominum: " Praecipis, ut educam populum istum, et non indicas mihi, quem missurus es mecum; cum dixeris: "Novi te ex nomine, et invenisti gratiam coram me".
EXOD|33|13|Si ergo inveni gratiam in conspectu tuo, ostende mihi viam tuam, ut sciam te et inveniam gratiam ante oculos tuos; respice quia populus tuus est natio haec ".
EXOD|33|14|Dixitque Dominus: " Facies mea ibit, et requiem dabo tibi ".
EXOD|33|15|Et ait Moyses: " Si non tu ipse eas, ne educas nos de loco isto;
EXOD|33|16|in quo enim scietur me et populum tuum invenisse gratiam in conspectu tuo, nisi ambulaveris nobiscum, ut glorificemur ego et populus tuus prae omnibus populis, qui habitant super terram? ".
EXOD|33|17|Dixitque Dominus ad Moysen: " Et verbum istud, quod locutus es, faciam; invenisti enim gratiam coram me, et teipsum novi ex nomine ".
EXOD|33|18|Qui ait: " Ostende mihi gloriam tuam ".
EXOD|33|19|Respondit: " Ego ostendam omne bonum tibi et vocabo in nomine Domini coram te; et miserebor, cui voluero, et clemens ero, in quem mihi placuerit ".
EXOD|33|20|Rursumque ait: " Non poteris videre faciem meam; non enim videbit me homo et vivet ".
EXOD|33|21|Et iterum: " Ecce, inquit, est locus apud me, stabis super petram;
EXOD|33|22|cumque transibit gloria mea, ponam te in foramine petrae et protegam dextera mea, donec transeam;
EXOD|33|23|tollamque manum meam, et videbis posteriora mea; faciem autem meam videre non poteris ".
EXOD|34|1|Dixitque Dominus ad Moy sen: " Praecide tibi duas ta bulas lapideas instar priorum, et scribam super eas verba, quae habuerunt tabulae, quas fregisti.
EXOD|34|2|Esto paratus mane, ut ascendas statim in montem Sinai; stabisque mihi super verticem montis.
EXOD|34|3|Nullus ascendat tecum, nec videatur quispiam per totum montem; oves quoque et boves non pascantur e contra ".
EXOD|34|4|Excidit ergo duas tabulas lapideas, quales antea fuerant; et de nocte consurgens ascendit in montem Sinai, sicut praeceperat ei Dominus, portans secum tabulas.
EXOD|34|5|Cumque descendisset Dominus per nubem, stetit cum eo vocans in nomine Domini.
EXOD|34|6|Et transiens coram eo clamavit: " Dominus, Dominus Deus, misericors et clemens, patiens et multae miserationis ac verax,
EXOD|34|7|qui custodit misericordiam in milia, qui aufert iniquitatem et scelera atque peccata, nihil autem impunitum sinit, qui reddit iniquitatem patrum in filiis ac nepotibus in tertiam et quartam progeniem ".
EXOD|34|8|Festinusque Moyses curvatus est pronus in terram et adorans
EXOD|34|9|ait: " Si inveni gratiam in conspectu tuo, Domine, obsecro, ut gradiaris nobiscum; populus quidem durae cervicis est, sed tu auferes iniquitates nostras atque peccata nosque possidebis ".
EXOD|34|10|Respondit Dominus: " Ego inibo pactum coram universo populo tuo; mirabilia faciam, quae numquam visa sunt super totam terram nec in ullis gentibus, ut cernat cunctus populus, in cuius es medio, opus Domini terribile, quod facturus sum tecum.
EXOD|34|11|Observa cuncta, quae hodie mando tibi: ego ipse eiciam ante faciem tuam Amorraeum et Chananaeum et Hetthaeum, Pherezaeum quoque et Hevaeum et Iebusaeum.
EXOD|34|12|Cave, ne umquam cum habitatoribus terrae, quam intraveris, iungas amicitias, quae tibi sint in ruinam;
EXOD|34|13|sed aras eorum destrue, confringe lapides palosque succide.
EXOD|34|14|Noli adorare deum alienum: Dominus Zelotes nomen eius, Deus est aemulator.
EXOD|34|15|Ne ineas pactum cum hominibus illarum regionum, ne, cum fornicati fuerint cum diis suis et sacrificaverint eis, vocet te quispiam, et comedas de immolatis.
EXOD|34|16|Nec uxorem de filiabus eorum accipies filiis tuis, ne, postquam ipsae fuerint fornicatae cum diis suis, fornicari faciant et filios tuos in deos suos.
EXOD|34|17|Deos conflatiles non facies tibi.
EXOD|34|18|Sollemnitatem Azymorum custodies: septem diebus vesceris azymis, sicut praecepi tibi, in tempore constituto mensis Abib; mense enim verni temporis egressus es de Aegypto.
EXOD|34|19|Omne, quod aperit vulvam generis masculini, meum erit; de cuncto grege tuo tam de bobus quam de ovibus meum erit.
EXOD|34|20|Primogenitum asini redimes ove, sin autem nec pretium pro eo dederis, franges cervicem eius. Primogenitum filiorum tuorum redimes; nec apparebis in conspectu meo vacuus.
EXOD|34|21|Sex diebus operaberis, die septimo cessabis etiam arare et metere.
EXOD|34|22|Sollemnitatem Hebdomadarum facies tibi in primitiis frugum messis tuae triticeae et sollemnitatem Collectae, quando, redeunte anni tempore, cuncta conduntur.
EXOD|34|23|Tribus temporibus anni apparebit omne masculinum tuum in conspectu omnipotentis Domini, Dei Israel.
EXOD|34|24|Cum enim tulero gentes a facie tua et dilatavero terminos tuos, nullus insidiabitur terrae tuae, ascendente te et apparente in conspectu Domini Dei tui ter in anno.
EXOD|34|25|Non immolabis super fermento sanguinem hostiae meae; neque residebit mane de victima sollemnitatis Paschae.
EXOD|34|26|Primitias frugum terrae tuae afferes in domum Domini Dei tui.Non coques haedum in lacte matris suae ".
EXOD|34|27|Dixitque Dominus ad Moysen: " Scribe tibi verba haec, quibus et tecum et cum Israel pepigi foedus ".
EXOD|34|28|Fuit ergo ibi cum Domino quadraginta dies et quadraginta noctes; panem non comedit et aquam non bibit et scripsit in tabulis verba foederis, decem verba.
EXOD|34|29|Cumque descenderet Moyses de monte Sinai, tenebat duas tabulas testimonii et ignorabat quod resplenderet cutis faciei suae ex consortio sermonis Domini.
EXOD|34|30|Videntes autem Aaron et filii Israel resplendere cutem faciei Moysi, timuerunt prope accedere;
EXOD|34|31|vocatique ab eo reversi sunt tam Aaron quam principes synagogae. Et postquam locutus est ad eos,
EXOD|34|32|venerunt ad eum etiam omnes filii Israel; quibus praecepit cuncta, quae audierat a Domino in monte Sinai.
EXOD|34|33|Impletisque sermonibus, posuit velamen super faciem suam,
EXOD|34|34|quod ingressus ad Dominum et loquens cum eo auferebat, donec exiret; et tunc loquebatur ad filios Israel omnia, quae sibi fuerant imperata.
EXOD|34|35|Qui videbant cutem faciei Moysi resplendere, sed operiebat ille rursus faciem suam, donec ingressus loqueretur cum eo.
EXOD|35|1|Igitur, congregato omni coetu filiorum Israel, dixit ad eos: " Haec sunt, quae iussit Dominus fieri:
EXOD|35|2|sex diebus facietis opus, septimus dies erit vobis sanctus, sabbatum et requies Domino; qui fecerit opus in eo, occidetur.
EXOD|35|3|Non succendetis ignem in omnibus habitaculis vestris per diem sabbati ".
EXOD|35|4|Et ait Moyses ad omnem coetum filiorum Israel: " Iste est sermo, quem praecepit Dominus dicens:
EXOD|35|5|"Separate apud vos donaria Domino". Omnis voluntarius et proni animi offerat ea Domino: aurum et argentum et aes,
EXOD|35|6|hyacinthum et purpuram coccumque et byssum, pilos caprarum
EXOD|35|7|et pelles arietum rubricatas et pelles delphini, ligna acaciae
EXOD|35|8|et oleum ad luminaria concinnanda et aromata, ut conficiatur unguentum et thymiama suavissimum,
EXOD|35|9|lapides onychinos et gemmas ad ornatum ephod et pectoralis.
EXOD|35|10|Quisquis vestrum sapiens est, veniat et faciat, quod Dominus imperavit,
EXOD|35|11|habitaculum scilicet et tentorium eius atque operimentum, fibulas et tabulata cum vectibus, columnas et bases;
EXOD|35|12|arcam et vectes, propitiatorium et velum, quod ante illud oppanditur;
EXOD|35|13|mensam cum vectibus et vasis et propositionis panibus;
EXOD|35|14|candelabrum ad luminaria sustentanda, vasa illius et lucernas et oleum ad nutrimenta luminarium;
EXOD|35|15|altare thymiamatis et vectes et oleum unctionis et thymiama ex aromatibus; velum ad ostium habitaculi;
EXOD|35|16|altare holocausti et craticulam eius aeneam cum vectibus et vasis suis, labrum et basim eius;
EXOD|35|17|cortinas atrii cum columnis et basibus, velum in foribus atrii;
EXOD|35|18|paxillos habitaculi et atrii cum funiculis suis;
EXOD|35|19|vestimenta texta, quorum usus est in ministerio sanctuarii, vestes sanctas Aaron pontificis ac vestes filiorum eius, ut sacerdotio fungantur mihi ".
EXOD|35|20|Egressus est omnis coetus filiorum Israel de conspectu Moysi,
EXOD|35|21|et venit, quisquis erat mentis promptissimae, et attulit sponte sua donaria Domino ad faciendum opus tabernaculi conventus et quidquid ad cultum et ad vestes sanctas necessarium erat.
EXOD|35|22|Viri cum mulieribus, omnes voluntarii praebuerunt fibulas et inaures, anulos et dextralia; omne vas aureum in donaria Domini separatum est.
EXOD|35|23|Si quis habebat hyacinthum et purpuram coccumque, byssum et pilos caprarum, pelles arietum rubricatas et pelles delphini,
EXOD|35|24|argenti aerisque metalla, obtulerunt Domino lignaque acaciae in varios usus.
EXOD|35|25|Sed et mulieres eruditae dederunt, quae neverant, hyacinthum, purpuram et coccum ac byssum
EXOD|35|26|et pilos caprarum, sponte propria cuncta tribuentes.
EXOD|35|27|Principes vero obtulerunt lapides onychinos et gemmas ad ephod et pectorale
EXOD|35|28|aromataque et oleum ad luminaria concinnanda et ad praeparandum unguentum ac thymiama odoris suavissimi componendum.
EXOD|35|29|Omnes viri et mulieres mente prompta obtulerunt donaria, ut fierent opera, quae iusserat Dominus per manum Moysi. Cuncti filii Israel voluntaria Domino dedicaverunt.
EXOD|35|30|Dixitque Moyses ad filios Israel: " Ecce vocavit Dominus ex nomine Beseleel filium Uri filii Hur de tribu Iudae;
EXOD|35|31|implevitque eum spiritu Dei, sapientia et intellegentia et scientia ad omne opus,
EXOD|35|32|ad excogitandum et faciendum opus in auro et argento et aere,
EXOD|35|33|ad scindendum et includendum gemmas et ad sculpendum ligna, quidquid fabre adinveniri potest.
EXOD|35|34|Dedit quoque in corde eius, ut alios doceret, ipsi et Ooliab filio Achisamech de tribu Dan.
EXOD|35|35|Ambos implevit sapientia, ut faciant opera fabri polymitarii ac plumarii de hyacintho ac purpura coccoque et bysso et textoris, facientes omne opus ac nova quaeque reperientes ".
EXOD|36|1|Fecit ergo Beseleel et Ooliab et omnis vir sapiens, quibus dedit Dominus sapientiam et intellectum, ut scirent fabre operari, quae in usus sanctuarii necessaria sunt et quae praecepit Dominus.
EXOD|36|2|Cumque vocasset Moyses Beseleel et Ooliab et omnem eruditum virum, cui dederat Dominus sapientiam, omnes, qui sponte sua obtulerant se ad faciendum opus,
EXOD|36|3|acceperunt ab ipso universa donaria, quae attulerant filii Israel ad faciendum opus in cultum sanctuarii. Ipsi autem cotidie mane donaria ei offerebant.
EXOD|36|4|Unde omnes sapientes artifices venerunt singuli de opere suo pro sanctuario
EXOD|36|5|et dixerunt Moysi: " Plus offert populus quam necessarium est operi, quod Dominus iussit facere ".
EXOD|36|6|Iussit ergo Moyses praeconis voce per castra clamari: " Nec vir nec mulier quidquam offerat ultra pro omni opere sanctuario ". Sicque cessatum est a muneribus offerendis,
EXOD|36|7|eo quod oblata sufficerent et superabundarent.
EXOD|36|8|Feceruntque omnes corde sapientes inter artifices habitaculi cortinas decem de bysso retorta et hyacintho et purpura coccoque, cum cherubim intextis arte polymita;
EXOD|36|9|quarum una habebat in longitudine viginti octo cubitos et in latitudine quattuor: una mensura erat omnium cortinarum.
EXOD|36|10|Coniunxitque cortinas quinque alteram alteri et alias quinque sibi invicem copulavit.
EXOD|36|11|Fecit et ansas hyacinthinas in ora cortinae unius in extremitate iuncturae et in ora cortinae extremae in iunctura altera similiter.
EXOD|36|12|Quinquagenas ansas fecit pro utraque cortina, ut contra se invicem venirent ansae et mutuo iungerentur.
EXOD|36|13|Unde et quinquaginta fudit fibulas aureas, quae morderent cortinarum ansas, et fieret unum habitaculum.
EXOD|36|14|Fecit et saga undecim de pilis caprarum pro tentorio super habitaculum;
EXOD|36|15|unum sagum in longitudine habebat cubitos triginta et in latitudine cubitos quattuor: unius mensurae erant omnia saga.
EXOD|36|16|Quorum quinque iunxit seorsum et sex alia separatim.
EXOD|36|17|Fecitque ansas quinquaginta in ora sagi ultimi iuncturae unius et quinquaginta in ora sagi iuncturae alterius, ut sibi invicem iungerentur;
EXOD|36|18|et fecit fibulas aeneas quinquaginta, quibus necteretur tentorium, ut esset unum.
EXOD|36|19|Fecit et opertorium tentorio de pellibus arietum rubricatis aliudque desuper velamentum de pellibus delphini.
EXOD|36|20|Fecit et tabulas habitaculi de lignis acaciae stantes.
EXOD|36|21|Decem cubitorum erat longitudo tabulae unius, et unum ac semis cubitum latitudo retinebat.
EXOD|36|22|Bini pedes erant per singulas tabulas, ut altera alteri iungeretur: sic fecit in omnibus tabulis habitaculi.
EXOD|36|23|E quibus viginti ad plagam meridianam erant contra austrum
EXOD|36|24|cum quadraginta basibus argenteis. Duae bases sub singulis tabulis ponebantur pro duabus pedibus.
EXOD|36|25|Ad plagam quoque habitaculi, quae respicit ad aquilonem, fecit viginti tabulas
EXOD|36|26|cum quadraginta basibus argenteis: duas bases per singulas tabulas.
EXOD|36|27|Contra occidentem vero, id est ad eam partem habitaculi quae mare respicit, fecit sex tabulas
EXOD|36|28|et duas alias per singulos angulos habitaculi retro;
EXOD|36|29|quae gemellae erant a deorsum usque sursum in unam compaginem. Ita fecit duas tabulas in duobus angulis,
EXOD|36|30|ut octo essent simul tabulae et haberent bases argenteas sedecim: binas scilicet bases sub singulis tabulis.
EXOD|36|31|Fecit et vectes de lignis acaciae quinque ad continendas tabulas unius lateris habitaculi
EXOD|36|32|et quinque alios ad alterius lateris coaptandas tabulas; et extra hos quinque alios vectes ad occidentalem plagam habitaculi contra mare.
EXOD|36|33|Fecit autem vectem medium, qui per medias tabulas ab una extremitate usque ad alteram perveniret.
EXOD|36|34|Ipsa autem tabulata deauravit. Et anulos eorum fecit aureos, per quos vectes induci possent; quos et ipsos laminis aureis operuit.
EXOD|36|35|Fecit et velum de hyacintho et purpura coccoque ac bysso retorta, opere polymitario, cum cherubim intextis;
EXOD|36|36|et quattuor columnas de lignis acaciae, quas cum uncis suis deauravit, fusis basibus earum argenteis.
EXOD|36|37|Fecit et velum in introitu tabernaculi ex hyacintho, purpura, cocco byssoque retorta opere plumarii;
EXOD|36|38|et columnas quinque cum uncis suis. Et operuit auro capita et anulos earum basesque earum fudit aeneas.
EXOD|37|1|Fecit autem Beseleel et ar cam de lignis acaciae haben tem duos semis cubitos in longitudine et cubitum ac semissem in latitudine, altitudo quoque unius cubiti fuit et dimidii; vestivitque eam auro purissimo intus ac foris.
EXOD|37|2|Et fecit illi coronam auream per gyrum,
EXOD|37|3|conflans quattuor anulos aureos in quattuor pedibus eius; duos anulos in latere uno et duos in altero.
EXOD|37|4|Vectes quoque fecit de lignis acaciae, quos vestivit auro
EXOD|37|5|et quos misit in anulos, qui erant in lateribus arcae, ad portandum eam.
EXOD|37|6|Fecit et propitiatorium de auro mundissimo: duorum cubitorum et dimidii in longitudine et cubiti ac semis in latitudine.
EXOD|37|7|Duos etiam cherubim ex auro ductili fecit ex utraque parte propitiatorii:
EXOD|37|8|cherub unum ex summitate unius partis et cherub alterum ex summitate partis alterius; duos cherubim ex singulis summitatibus propitiatorii
EXOD|37|9|extendentes alas sursum et tegentes alis suis propitiatorium seque mutuo et illud respicientes.
EXOD|37|10|Fecit et mensam de lignis acaciae in longitudine duorum cubitorum et in latitudine unius cubiti, quae habebat in altitudine cubitum ac semissem;
EXOD|37|11|circumdeditque eam auro mundissimo et fecit illi coronam auream per gyrum.
EXOD|37|12|Fecit ei quoque limbum aureum quattuor digitorum per circuitum et super illum coronam auream.
EXOD|37|13|Fudit et quattuor circulos aureos, quos posuit in quattuor angulis per singulos pedes mensae
EXOD|37|14|iuxta limbum; misitque in eos vectes, ut possit mensa portari.
EXOD|37|15|Ipsos quoque vectes fecit de lignis acaciae et circumdedit eos auro;
EXOD|37|16|et vasa ad diversos usus mensae, acetabula, phialas et cyathos et crateras ex auro puro, in quibus offerenda sunt libamina.
EXOD|37|17|Fecit et candelabrum ductile de auro mundissimo, basim et hastile eius; scyphi sphaerulaeque ac flores unum cum ipso erant:
EXOD|37|18|sex in utroque latere, tres calami ex parte una et tres ex altera;
EXOD|37|19|tres scyphi in nucis modum in calamo uno sphaerulaeque simul et flores et tres scyphi instar nucis in calamo altero sphaerulaeque simul et flores. Aequum erat opus sex calamorum, qui procedebant de hastili candelabri.
EXOD|37|20|In ipso autem hastili erant quattuor scyphi in nucis modum sphaerulaeque et flores;
EXOD|37|21|singulae sphaerulae sub binis calamis per loca tria, qui simul sex fiunt calami procedentes de hastili uno.
EXOD|37|22|Sphaerulae igitur et calami unum cum ipso erant, totum ductile ex auro purissimo.
EXOD|37|23|Fecit et lucernas septem cum emunctoriis suis et vasa, ubi emuncta condantur, de auro mundissimo.
EXOD|37|24|Talentum auri purissimi appendebat candelabrum cum omnibus vasis suis.
EXOD|37|25|Fecit et altare thymiamatis de lignis acaciae habens per quadrum singulos cubitos et in altitudine duos; e cuius angulis procedebant cornua.
EXOD|37|26|Vestivitque illud auro purissimo cum craticula ac parietibus et cornibus.
EXOD|37|27|Fecitque ei coronam aureolam per gyrum et binos anulos aureos sub corona in duobus lateribus, ut mittantur in eos vectes, et possit altare portari.
EXOD|37|28|Ipsos autem vectes fecit de lignis acaciae et operuit laminis aureis.
EXOD|37|29|Composuit et oleum ad sanctificationis unguentum et thymiama de aromatibus mundissimis opere pigmentarii.
EXOD|38|1|Fecit et altare holocausti de lignis acaciae quinque cubi torum per quadrum et trium in altitudine,
EXOD|38|2|cuius cornua de angulis procedebant; operuitque illud laminis aeneis.
EXOD|38|3|Et in usus eius paravit ex aere vasa diversa: lebetes, vatilla et pateras, fuscinulas et ignium receptacula.
EXOD|38|4|Craticulamque eius in modum retis fecit aeneam subter marginem altaris ab imo usque ad medium eius,
EXOD|38|5|fusis quattuor anulis per totidem craticulae summitates, ad immittendos vectes ad portandum.
EXOD|38|6|Quos et ipsos fecit de lignis acaciae et operuit laminis aeneis;
EXOD|38|7|induxitque in circulos, qui in lateribus altaris eminebant. Ipsum autem altare non erat solidum, sed cavum ex tabulis et intus vacuum.
EXOD|38|8|Fecit et labrum aeneum cum basi sua de speculis mulierum, quae excubabant in ostio tabernaculi conventus.
EXOD|38|9|Fecit et atrium, in cuius australi plaga erant tentoria de bysso retorta cubitorum centum;
EXOD|38|10|columnae aeneae viginti cum basibus suis; unci columnarum et anuli earum argentei.
EXOD|38|11|Aeque ad septentrionalem plagam tentoria, columnae basesque et unci anulique columnarum eiusdem mensurae et operis ac metalli erant.
EXOD|38|12|In ea vero plaga, quae ad occidentem respicit, fuerunt tentoria cubitorum quinquaginta, columnae decem cum basibus suis; et unci columnarum anulique earum argentei.
EXOD|38|13|Porro contra orientem quinquaginta cubitorum paravit tentoria,
EXOD|38|14|e quibus quindecim cubitos columnarum trium cum basibus suis unum tenebat latus;
EXOD|38|15|et in parte altera ­ quia inter utraque introitum tabernaculi fecit ­ quindecim aeque cubitorum erant tentoria columnaeque tres et bases totidem.
EXOD|38|16|Cuncta atrii tentoria in circuitu ex bysso retorta texuerat.
EXOD|38|17|Bases columnarum fuere aeneae, unci autem earum et anuli earum argentei et capita earum vestivit argento et omnes columnas atrii cinxit anulis argenteis.
EXOD|38|18|Et in introitu eius opere plumario fecit velum ex hyacintho, purpura, cocco ac bysso retorta; quod habebat viginti cubitos in longitudine, altitudo vero quinque cubitorum erat iuxta mensuram, quam cuncta atrii tentoria habebant.
EXOD|38|19|Columnae autem in ingressu fuere quattuor cum basibus aeneis, uncis argenteis; capitaque et anulos earum vestivit argento.
EXOD|38|20|Paxillos quoque habitaculi et atrii per gyrum fecit aeneos.
EXOD|38|21|Hic est census habitaculi, habitaculi testimonii, qui recensitus est iuxta praeceptum Moysi ministerio Levitarum per manum Ithamar filii Aaron sacerdotis.
EXOD|38|22|Beseleel filius Uri filii Hur de tribu Iudae fecit cuncta, quae praeceperat Dominus Moysi,
EXOD|38|23|iuncto sibi socio Ooliab filio Achisamech de tribu Dan fabro et polymitario atque plumario ex hyacintho, purpura, cocco et bysso.
EXOD|38|24|Omne aurum, quod expensum est in opere sanctuarii et quod oblatum est in donariis, viginti novem talentorum fuit et septingentorum triginta siclorum ad mensuram sicli sanctuarii.
EXOD|38|25|Argentum autem eorum, qui in congregatione recensiti sunt, centum talentorum fuit et mille septingentorum et septuaginta quinque siclorum ad mensuram sicli sanctuarii.
EXOD|38|26|Beca, id est dimidium sicli iuxta mensuram sicli sanctuarii, dedit quisquis transit ad censum a viginti annis et supra, de sescentis tribus milibus et quingentis quinquaginta armatorum.
EXOD|38|27|De talentis centum argenti conflatae sunt bases sanctuarii et veli, singulis talentis per bases singulas supputatis.
EXOD|38|28|De mille autem septingentis et septuaginta quinque siclis fecit uncos columnarum et vestivit capita earum et cinxit eas argento.
EXOD|38|29|Aeris quoque oblata sunt septuaginta talenta et duo milia et quadringenti sicli,
EXOD|38|30|ex quibus fecit bases in introitu tabernaculi conventus et altare aeneum cum craticula sua omniaque vasa, quae ad usum eius pertinent,
EXOD|38|31|et bases atrii tam in circuitu quam in ingressu eius et omnes paxillos habitaculi atque atrii per gyrum.
EXOD|39|1|De hyacintho vero et purpura, cocco ac bysso fecerunt vestes textas pro ministerio sanctuarii. Et fecerunt vestes sacras Aaron, sicut praecepit Dominus Moysi.
EXOD|39|2|Fecerunt igitur ephod de auro, hyacintho et purpura coccoque et bysso retorta
EXOD|39|3|opere polymitario tundentes bratteas aureas et extenuantes in fila, ut possent torqueri cum priorum colorum subtegmine.
EXOD|39|4|Fasciasque umerales fecerunt ei, cum quibus in utroque latere summitatum suarum copulabatur,
EXOD|39|5|et balteum, quo constringebatur ephod, eiusdem operis et unum cum eo ex auro, et hyacintho et purpura coccoque et bysso retorta, sicut praeceperat Dominus Moysi.
EXOD|39|6|Paraverunt et duos lapides onychinos, inclusos texturis aureis et sculptos arte gemmaria nominibus filiorum Israel;
EXOD|39|7|posueruntque eos in fasciis umeralibus ephod, lapides memorialis filiorum Israel, sicut praeceperat Dominus Moysi.
EXOD|39|8|Fecerunt et pectorale opere polymito iuxta opus ephod ex auro, hyacintho, purpura coccoque et bysso retorta,
EXOD|39|9|quadrangulum duplex mensurae palmi.
EXOD|39|10|Et posuerunt in eo gemmarum ordines quattuor: in primo versu erat sardius, topazius, smaragdus;
EXOD|39|11|in secundo carbunculus, sapphirus et iaspis;
EXOD|39|12|in tertio hyacinthus, achates et amethystus;
EXOD|39|13|in quarto chrysolithus, onychinus et beryllus: inclusi textura aurea per ordines suos.
EXOD|39|14|Ipsique lapides duodecim sculpti erant nominibus duodecim tribuum Israel, singuli per nomina singulorum.
EXOD|39|15|Fecerunt in pectorali catenulas quasi funiculos opus tortile de auro purissimo
EXOD|39|16|et duos margines aureos totidemque anulos aureos. Porro duos anulos posuerunt in utraque summitate pectoralis;
EXOD|39|17|duos funiculos aureos inseruerunt anulis, qui in pectoralis angulis eminebant.
EXOD|39|18|Duas summitates amborum funiculorum colligaverunt duobus marginibus in fasciis umeralibus ephod in parte eius anteriore.
EXOD|39|19|Et fecerunt duos anulos aureos et posuerunt super duas summitates pectoralis in eius margine interiore contra ephod, sicut praecepit Dominus Moysi.
EXOD|39|20|Feceruntque duos anulos aureos, quos posuerunt in duabus fasciis umeralibus ephod deorsum in latere eius anteriore secus iuncturam eius super balteum ephod.
EXOD|39|21|Et strinxerunt pectorale anulis eius ad anulos ephod vitta hyacinthina, ut esset super balteum ephod, ne amoveretur ab ephod, sicut praecepit Dominus Moysi.
EXOD|39|22|Fecerunt quoque pallium ephod opere textili totum hyacinthinum
EXOD|39|23|et capitium in medio eius supra oramque per gyrum sicut in capitio loricae;
EXOD|39|24|deorsum autem ad pedes mala punica ex hyacintho, purpura, cocco ac bysso retorta
EXOD|39|25|et tintinnabula de auro purissimo, quae posuerunt inter malogranata in inferiore parte pallii per gyrum,
EXOD|39|26|ut sit tintinnabulum inter singula mala punica, quibus ornatus incedebat pontifex, quando ministerio fungebatur, sicut praeceperat Dominus Moysi.
EXOD|39|27|Fecerunt et tunicas byssinas opere textili Aaron et filiis eius
EXOD|39|28|et tiaram et ornatum mitrarum ex bysso, feminalia quoque linea ex bysso retorta,
EXOD|39|29|cingulum vero de bysso retorta, hyacintho, purpura ac cocco, arte plumaria, sicut praeceperat Dominus Moysi.
EXOD|39|30|Fecerunt et laminam diadema sanctitatis de auro purissimo; scripseruntque in ea opere caelatoris: " Sanctum Domino ";
EXOD|39|31|et strinxerunt eam desuper cum tiara vitta hyacinthina, sicut praeceperat Dominus Moysi.
EXOD|39|32|Perfectum est igitur omne opus habitaculi et tabernaculi conventus; feceruntque filii Israel cuncta, quae praeceperat Dominus Moysi: sic fecerunt.
EXOD|39|33|Et obtulerunt habitaculum et tabernaculum et universam supellectilem, fibulas, tabulas, vectes, columnas ac bases,
EXOD|39|34|opertorium de pellibus arietum rubricatis et operimentum de pellibus delphini, velum,
EXOD|39|35|arcam testimonii, vectes, propitiatorium,
EXOD|39|36|mensam cum vasis suis et propositionis panibus,
EXOD|39|37|candelabrum ex auro puro, lucernas in ordine earum et utensilia earum cum oleo candelabri,
EXOD|39|38|altare aureum et unguentum et thymiama ex aromatibus et velum in introitu tabernaculi,
EXOD|39|39|altare aeneum, craticulam aeneam, vectes et vasa eius omnia, labrum cum basi sua,
EXOD|39|40|tentoria atrii et columnas cum basibus suis, velum in introitu atrii funiculosque illius et paxillos. Nihil ex vasis defuit, quae in ministerium habitaculi in tabernaculo conventus iussa sunt fieri.
EXOD|39|41|Vestes quoque textas, quibus sacerdotes utuntur in sanctuario, et vestes sacras Aaron sacerdotis et vestes filiorum eius
EXOD|39|42|obtulerunt filii Israel, sicut praeceperat Dominus Moysi.
EXOD|39|43|Quae postquam Moyses cuncta vidit completa, benedixit eis.
EXOD|40|1|Locutusque est Dominus ad Moysen dicens:
EXOD|40|2|" Mense pri mo, die prima mensis eriges habitaculum, tabernaculum conventus,
EXOD|40|3|et pones in eo arcam testimonii, abscondes illam velo;
EXOD|40|4|et, illata mensa, pones super eam, quae rite praecepta sunt. Candelabrum stabit cum lucernis suis
EXOD|40|5|et altare aureum, in quo adoletur incensum, coram arca testimonii. Velum in introitu habitaculi pones,
EXOD|40|6|et ante tabernaculum conventus altare holocausti,
EXOD|40|7|et labrum inter altare et tabernaculum conventus et implebis illud aqua.
EXOD|40|8|Circumdabisque atrium tentoriis et pones velum in porta eius.
EXOD|40|9|Et, assumpto unctionis oleo, unges habitaculum et omnia, quae in eo sunt, et consecrabis illud cum vasis suis, et erit sanctum.
EXOD|40|10|Unges quoque altare holocausti et omnia vasa eius et consecrabis altare, et erit sanctum sanctorum.
EXOD|40|11|Et unges labrum cum basi sua et consecrabis illud.
EXOD|40|12|Applicabisque Aaron et filios eius ad fores tabernaculi conventus; et lotos aqua
EXOD|40|13|indues Aaron sanctis vestibus, unges et consecrabis eum, ut mihi sacerdotio fungatur;
EXOD|40|14|filios eius applicabis et vesties eos tunicis
EXOD|40|15|et unges eos, sicut unxisti patrem eorum, ut mihi sacerdotio fungantur, et unctio eorum erit eis in sacerdotium sempiternum in generationibus eorum ".
EXOD|40|16|Fecitque Moyses omnia, quae praeceperat ei Dominus: sic fecit.
EXOD|40|17|Igitur mense primo anni secundi, prima die mensis collocatum est habitaculum.
EXOD|40|18|Erexitque Moyses illud et posuit bases ac tabulas et vectes statuitque columnas
EXOD|40|19|et expandit tentorium super habitaculum, imposito desuper operimento, sicut Dominus imperaverat Moysi.
EXOD|40|20|Sumpsit et posuit testimonium in arca et, subditis infra vectibus, posuit propitiatorium desuper.
EXOD|40|21|Cumque intulisset arcam in habitaculum, appendit ante eam velum, sicut iusserat Dominus Moysi.
EXOD|40|22|Posuit et mensam in tabernaculo conventus ad plagam septentrionalem extra velum,
EXOD|40|23|ordinatis coram propositionis panibus, sicut praeceperat Dominus Moysi.
EXOD|40|24|Posuit et candelabrum in tabernaculo conventus e regione mensae in parte australi,
EXOD|40|25|locatis per ordinem lucernis, sicut praeceperat Dominus Moysi.
EXOD|40|26|Posuit et altare aureum in tabernaculo conventus coram propitiatorio
EXOD|40|27|et adolevit super eo incensum aromatum, sicut iusserat Dominus Moysi.
EXOD|40|28|Posuit et velum in introitu habitaculi
EXOD|40|29|et altare holocausti in vestibulo habitaculi, tabernaculi conventus, offerens in eo holocaustum et sacrificium, sicut Dominus imperaverat Moysi.
EXOD|40|30|Labrum quoque statuit inter tabernaculum conventus et altare implens illud aqua;
EXOD|40|31|laveruntque Moyses et Aaron ac filii eius manus suas et pedes,
EXOD|40|32|cum ingrederentur tabernaculum conventus et accederent ad altare, sicut praeceperat Dominus Moysi.
EXOD|40|33|Erexit et atrium per gyrum habitaculi et altaris, ducto in introitu eius velo. Sic complevit opus.
EXOD|40|34|Et operuit nubes tabernaculum conventus, et gloria Domini implevit habitaculum.
EXOD|40|35|Nec poterat Moyses ingredi tabernaculum conventus, quia habitavit nubes super illud, et gloria Domini replevit habitaculum.
EXOD|40|36|Si quando nubes de tabernaculo ascendebat, proficiscebantur filii Israel in omnibus stationibus suis;
EXOD|40|37|si autem non ascendebat nubes, non proficiscebantur usque in diem, quo levabatur.
EXOD|40|38|Nubes quippe Domini incubabat per diem habitaculo, et ignis in nocte, ante oculos universae domus Israel per cunctas mansiones suas." "
