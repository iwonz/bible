2CHR|1|1|大衛 的兒子 所羅門 鞏固他的國度；耶和華－他的上帝與他同在，使他極其尊大。
2CHR|1|2|所羅門 吩咐全 以色列 ，就是千夫長、百夫長、審判官、全 以色列 的眾領袖和族長前來。
2CHR|1|3|所羅門 率領全會眾往 基遍 的丘壇去，因那裏有上帝的會幕，就是耶和華的僕人 摩西 在曠野所造的。
2CHR|1|4|只是上帝的約櫃， 大衛 已經從 基列‧耶琳 接到他所預備的地方，因他曾在 耶路撒冷 為約櫃支搭了帳幕，
2CHR|1|5|把 戶珥 的孫子， 烏利 的兒子 比撒列 所造的銅壇擺在 基遍 耶和華的會幕前。 所羅門 和會眾求告耶和華。
2CHR|1|6|所羅門 上到耶和華面前會幕的銅壇那裏，在壇上獻一千祭牲為燔祭。
2CHR|1|7|當夜，上帝向 所羅門 顯現，對他說：「你願我賜你甚麼，你可以求。」
2CHR|1|8|所羅門 對上帝說：「你曾向我父親 大衛 大施慈愛，使我接續他作王。
2CHR|1|9|耶和華上帝啊，現在求你實現向我父親 大衛 所應許的話；因你立我作這百姓的王，他們如同地上的塵沙那樣多。
2CHR|1|10|現在，求你賜我智慧聰明，好在這百姓面前出入；不然，誰能判斷你這麼多的百姓呢？」
2CHR|1|11|上帝對 所羅門 說：「你有這心意，不求資財、豐富、尊榮，也不求滅絕恨你之人的性命，又不求長壽；我既立你作我百姓的王，你只求智慧聰明，好審判我的百姓，
2CHR|1|12|我必賜你智慧聰明，也必賜你資財、豐富、尊榮，在你以前的列王未曾有過，在你以後也不會再有。」
2CHR|1|13|於是， 所羅門 從 基遍 丘壇會幕前回到 耶路撒冷 ，治理 以色列 。
2CHR|1|14|所羅門 聚集戰車騎兵；他有一千四百輛戰車，一萬二千名騎兵，安置在屯車城，在 耶路撒冷 的王那裏。
2CHR|1|15|王在 耶路撒冷 使金銀多如石頭，香柏木多如 謝非拉 的桑樹。
2CHR|1|16|所羅門 的馬是從 埃及 和 科威 運來的，是王的商人按著定價從 科威 買來的。
2CHR|1|17|他們從 埃及 進口戰車，每輛六百舍客勒銀子，馬每匹一百五十舍客勒； 赫 人眾王和 亞蘭 諸王的戰車和馬，也是經由他們的手出口的。
2CHR|2|1|所羅門 吩咐要為耶和華的名建造殿宇，又為自己的王國建造宮殿。
2CHR|2|2|所羅門 徵召七萬名扛抬的，八萬個在山上鑿石頭的人，三千六百個監工。
2CHR|2|3|所羅門 派人去見 推羅 王 希蘭 ，說：「你曾運香柏木給我父親 大衛 建造宮殿居住，請你也這樣待我。
2CHR|2|4|看哪，我要為耶和華－我上帝的名建造殿宇，分別為聖獻給他，在他面前燒芬芳的香，經常獻供餅，每早晚、安息日、初一，以及耶和華－我們上帝所定的節期獻燔祭。這是 以色列 人永遠的定例。
2CHR|2|5|我所要建造的殿宇宏大，因為我們的上帝至大，超乎眾神。
2CHR|2|6|天和天上的天，尚且不足他居住，誰能為他建造殿宇呢？我是誰，能為他建造殿宇嗎？不過在他面前燒香而已！
2CHR|2|7|現在請你派一個巧匠來，就是善用金、銀、銅、鐵，和紫色、朱紅色、藍色線做工，並精於雕刻之工的巧匠，與跟我一起在 猶大 和 耶路撒冷 、我父親 大衛 所預備的巧匠一同做工；
2CHR|2|8|又請你從 黎巴嫩 運香柏木、松木、檀香木到我這裏來，因我知道你的僕人擅長砍伐 黎巴嫩 的樹木。看哪，我的僕人必幫助你的僕人，
2CHR|2|9|好為我預備許多的木料，因我要建造的殿宇高大出奇。
2CHR|2|10|看哪，我必給你僕人，就是砍伐樹木的伐木工，二萬歌珥壓碎的小麥 ，二萬歌珥大麥，二萬罷特酒，二萬罷特油。」
2CHR|2|11|推羅 王 希蘭 寫信回答 所羅門 說：「耶和華因為愛他的百姓，所以立你作他們的王。」
2CHR|2|12|又說：「創造天和地的耶和華－ 以色列 的上帝是應當稱頌的！他賜給 大衛 王一個有智慧的兒子，使他有見識，有聰明，可以為耶和華建造殿宇，又為自己的王國建造宮殿。
2CHR|2|13|「現在我派一個精巧聰明的人去，他是我的師父 戶蘭 ，
2CHR|2|14|是 但 支派一個婦人的兒子，父親是 推羅 人。他善用金、銀、銅、鐵、石、木，和紫色、藍色、細麻和朱紅色線製造各物，並精於雕刻，又能設計各樣交給他做的圖案。我派這人與你的巧匠和你父親－我主 大衛 的巧匠一同做工。
2CHR|2|15|我主所說的小麥、大麥、酒、油，請運來給眾僕人。
2CHR|2|16|我們必照你所需用的，從 黎巴嫩 砍伐樹木，紮成筏子，浮海運到 約帕 ；你可以從那裏運到 耶路撒冷 。」
2CHR|2|17|所羅門 仿照他父親 大衛 數點所有在 以色列 地寄居的外邦人，共有十五萬三千六百名。
2CHR|2|18|他叫其中的七萬人作扛抬，八萬人在山上鑿石頭，三千六百人監督百姓工作。
2CHR|3|1|所羅門 在 耶路撒冷 開工建造耶和華的殿，就在耶和華向他父親 大衛 顯現的 摩利亞山 上， 耶布斯 人 阿珥楠 的禾場， 大衛 指定的地方。
2CHR|3|2|所羅門 作王第四年二月初二 開工建造。
2CHR|3|3|所羅門 所建築的上帝殿的根基是這樣：長六十肘，寬二十肘，都按著古時的尺寸。
2CHR|3|4|前面的 走廊長二十肘，與殿的寬度一樣，高一百二十肘；裏面貼上純金。
2CHR|3|5|大殿的牆都用松木板遮蔽，又貼上純金，上面刻著棕樹和鏈子。
2CHR|3|6|他用寶石裝飾這殿，使殿華美；金子都是 巴瓦音 的金子。
2CHR|3|7|他用金子貼殿和殿的棟梁、門檻、牆壁、門扇；牆上刻著基路伯。
2CHR|3|8|他建造至聖所，長二十肘，與殿的寬度一樣，寬二十肘，都貼上純金，共用了六百他連得金子。
2CHR|3|9|金的釘子重五十舍客勒。樓房都貼上金子。
2CHR|3|10|他又在至聖所用雕刻的手藝造兩個基路伯，包上金子。
2CHR|3|11|兩個基路伯的翅膀共長二十肘。這基路伯的一個翅膀長五肘，挨著殿這邊的牆；另一個翅膀也長五肘，與那基路伯翅膀相接。
2CHR|3|12|那基路伯的一個翅膀長五肘，挨著殿那邊的牆；另一個翅膀也長五肘，與這基路伯的翅膀相接。
2CHR|3|13|這兩個基路伯張開翅膀，共長二十肘，用腳站立，臉面向殿。
2CHR|3|14|他又用藍色、紫色、朱紅色線和細麻織幔子，在其上繡基路伯。
2CHR|3|15|他在殿前造了兩根柱子，高三十五肘；柱子上面的柱頂高五肘。
2CHR|3|16|他造鏈子在內殿裏，安在柱頂上，又做一百個石榴，安在鏈子上。
2CHR|3|17|他把兩根柱子立在殿前，一根在右邊，一根在左邊；右邊的起名叫 雅斤 ，左邊的起名叫 波阿斯 。
2CHR|4|1|他造一座銅壇，長二十肘，寬二十肘，高十肘。
2CHR|4|2|他又鑄一個銅海，周圍是圓的，直徑十肘，高五肘，用繩子量周圍是三十肘。
2CHR|4|3|銅海下面的周圍有牛的樣式，有十肘，繞著銅海；牛有兩行，是造銅海的時候鑄上去的。
2CHR|4|4|銅海安在十二頭銅牛上：三頭向北，三頭向西，三頭向南，三頭向東。銅海安在牛上，牛尾都向內。
2CHR|4|5|銅海厚一掌，邊如杯邊，像百合花，容量是三千罷特。
2CHR|4|6|他又造十個盆：五個放在右邊，五個放在左邊，作洗滌之用。獻燔祭所用之物都洗在盆內；但銅海是為祭司洗滌用的。
2CHR|4|7|他照所定的樣式造十個金燈臺，放在殿裏：五個在右邊，五個在左邊。
2CHR|4|8|他造十張桌子，放在殿裏：五張在右邊，五張在左邊。他又造一百個金碗。
2CHR|4|9|他建造祭司院和大院，以及院門，門扇包上銅。
2CHR|4|10|他把銅海安在殿的右邊，就是東南邊。
2CHR|4|11|戶蘭 又造了盆、鏟子和盤子。這樣， 戶蘭 為 所羅門 王做完了上帝殿的工：
2CHR|4|12|兩根柱子和柱子頂上兩個如碗的柱頂，以及蓋著如碗柱頂的兩個網子；
2CHR|4|13|四百個石榴，安在兩個網子上，每網兩行石榴，蓋著柱子上面兩個如碗的柱頂。
2CHR|4|14|他造盆座，又造其上的盆；
2CHR|4|15|銅海和其下的十二頭牛；
2CHR|4|16|盆、鏟子、肉叉。巧匠 戶蘭 給 所羅門 王為耶和華殿造的這一切器皿都是用磨亮的銅，
2CHR|4|17|是王在 約旦 平原、 疏割 和 撒利但 中間的泥巴地鑄成的。
2CHR|4|18|所羅門 造這一切器皿，數量很多，銅的重量無法計算。
2CHR|4|19|所羅門 又為上帝的殿造了各樣的器皿：金壇和獻供餅的供桌；
2CHR|4|20|純金的燈臺和燈盞，可以照定例點在內殿前；
2CHR|4|21|燈臺上的花和燈盞，以及燈剪，都是金的，而且是純金的；
2CHR|4|22|純金的鉗子、盤子、勺子、火盆。至於殿門和至聖所的門扇，以及殿的門扇，都是金的。
2CHR|5|1|所羅門 王做完了耶和華殿一切的工，就把他父親 大衛 分別為聖的金銀和一切器皿都帶來，放在上帝殿的庫房裏。
2CHR|5|2|於是， 所羅門 召集 以色列 的長老、各支派的領袖和 以色列 人的族長到 耶路撒冷 ，要把耶和華的約櫃從 大衛城 ，就是 錫安 ，接上來。
2CHR|5|3|在七月節期的時候，所有的 以色列 人都聚集到王那裏。
2CHR|5|4|以色列 眾長老一來到， 利未 人就抬起約櫃。
2CHR|5|5|祭司和 利未 人將約櫃請上來，又把會幕和會幕一切的聖器皿都帶上來。
2CHR|5|6|所羅門 王和聚集到他那裏的 以色列 全會眾都在約櫃前獻牛羊為祭，多得不可勝數，無法計算。
2CHR|5|7|祭司將耶和華的約櫃請進內殿，就是至聖所，安置在兩個基路伯的翅膀底下約櫃自己的地方。
2CHR|5|8|基路伯張開翅膀在約櫃上面的地方，從上面遮住約櫃和抬櫃的槓。
2CHR|5|9|這槓很長，從內殿前的約櫃可以看見槓頭，從外面卻看不見。這槓直到今日還在那裏。
2CHR|5|10|約櫃裏沒有別的，只有兩塊石版，就是 以色列 人出 埃及 ，耶和華與他們立約的時候， 摩西 在 何烈山 所放的。
2CHR|5|11|當時，所有在那裏的祭司，不論哪個班次供職的，都使自己分別為聖。祭司從聖所出來的時候，
2CHR|5|12|所有歌唱的 利未 人， 亞薩 、 希幔 、 耶杜頓 ，和他們的眾兒子、眾弟兄都穿細麻布衣服，站在祭壇的東邊敲鈸，鼓瑟，彈琴，和他們一起的還有一百二十個吹號的祭司。
2CHR|5|13|吹號的、歌唱的都合一齊聲，讚美稱謝耶和華。他們配合號筒、鐃鈸和其他樂器，揚聲讚美耶和華： 「耶和華本為善， 他的慈愛永遠長存！」 那時，耶和華的殿充滿了雲彩。
2CHR|5|14|祭司因雲彩的緣故不能站立供職，因為耶和華的榮光充滿了上帝的殿。
2CHR|6|1|那時， 所羅門 說： 「耶和華曾說要住在幽暗之處。
2CHR|6|2|我為你建了一座雄偉的殿宇， 作為你永遠居住的地方。」
2CHR|6|3|王轉過臉來為 以色列 全會眾祝福， 以色列 全會眾都站立。
2CHR|6|4|所羅門 說：「耶和華－ 以色列 的上帝是應當稱頌的！因他親口向我父 大衛 應許的，也親手成就了；他曾說：
2CHR|6|5|『自從那日我領我百姓出 埃及 地以來，我未曾在 以色列 各支派中選擇一城，在那裏為我的名建造殿宇，也未曾揀選一人作我百姓 以色列 的君王。
2CHR|6|6|但我選擇 耶路撒冷 ，使我的名留在那裏，又揀選 大衛 治理我的百姓 以色列 。』
2CHR|6|7|我父 大衛 的心意是要為耶和華－ 以色列 上帝的名建殿。
2CHR|6|8|耶和華卻對我父 大衛 說：『你有心為我的名建殿，這心意是好的；
2CHR|6|9|但你不可建殿，惟有你親生的兒子才可為我的名建殿。』
2CHR|6|10|現在耶和華實現了他所應許的話，使我接續我父 大衛 坐 以色列 的王位，正如耶和華所說的，我也為耶和華－ 以色列 上帝的名建造了這殿。
2CHR|6|11|我將約櫃安置在那裏，櫃內有耶和華的約，就是他與 以色列 人所立的約。」
2CHR|6|12|所羅門 當著 以色列 全會眾，站在耶和華的壇前，舉起手來。
2CHR|6|13|所羅門 曾造一個銅臺，長五肘，寬五肘，高三肘，放在院中。他站在臺上，當著 以色列 全會眾雙膝跪下，向天舉手，
2CHR|6|14|說：「耶和華－ 以色列 的上帝啊，天上地下沒有神明可與你相比！你向那些盡心行在你面前的僕人守約施慈愛，
2CHR|6|15|這約是你向你僕人 大衛 守的，是你應許他的。你親口應許，親手成就，正如今日一樣。
2CHR|6|16|耶和華－ 以色列 的上帝啊，你向你僕人我父 大衛 應許說：『你的子孫若謹慎自己的行為，遵行我的律法，像你在我面前所行的，就不斷有人在我面前坐 以色列 的王位。』現在求你信守這話。
2CHR|6|17|耶和華－ 以色列 的上帝啊，現在求你成就向你僕人 大衛 所應許的話。
2CHR|6|18|「上帝果真與世人同住在地上嗎？看哪，天和天上的天尚且不足容納你，何況我所建的這殿呢？
2CHR|6|19|惟求耶和華－我的上帝垂顧僕人的禱告祈求，俯聽僕人在你面前的祈禱呼求。
2CHR|6|20|願你的眼目晝夜看顧這殿，就是你應許立為你名的居所；求你垂聽禱告，你僕人向此處的禱告。
2CHR|6|21|你僕人和你百姓 以色列 向此處祈禱的時候，求你從天上你的居所垂聽，垂聽而赦免。
2CHR|6|22|「人若得罪鄰舍，有人強迫他，要他起誓，他來到這殿，在你的壇前起誓，
2CHR|6|23|求你從天上垂聽、處理，向你的僕人施行審判，定惡人有罪，照他所行的報應在他頭上；定義人為義，照他的義賞賜他。
2CHR|6|24|「你的百姓 以色列 若得罪你，敗在仇敵面前，卻又歸向你，宣認你的名，在這殿裏向你祈求禱告，
2CHR|6|25|求你從天上垂聽，赦免你百姓 以色列 的罪，使他們歸回你賜給他們和他們列祖之地。
2CHR|6|26|「你的百姓若得罪了你，你使天閉塞不下雨；他們若向此處禱告，宣認你的名，因你的懲罰而離開他們的罪，
2CHR|6|27|求你在天上垂聽，赦免你僕人你百姓 以色列 的罪，將當行的善道教導他們，並降雨在你的地，就是你賜給你百姓為業之地。
2CHR|6|28|「這地若有饑荒、瘟疫、焚風 、霉爛、蝗蟲、螞蚱，或有仇敵圍困這地的城門，無論遭遇甚麼災禍疾病，
2CHR|6|29|你的百姓 以色列 ，或眾人或一人，自覺災禍困苦，向這殿舉手，無論祈求甚麼，禱告甚麼，
2CHR|6|30|求你從天上你的居所垂聽赦免。因為你知道人心，惟有你知道世人的心，求你照各人所行的一切待他們，
2CHR|6|31|使他們在你賜給我們列祖的土地上一生一世敬畏你，遵行你的道。
2CHR|6|32|「論到不屬你百姓 以色列 的外邦人，若為你的大名和大能的手，以及伸出來的膀臂，從遠方而來，來向這殿禱告，
2CHR|6|33|求你從天上你的居所垂聽，照著外邦人向你所求的一切而行，使地上萬民都認識你的名，敬畏你，像你的百姓 以色列 一樣，又使他們知道我所建造的是稱為你名下的殿。
2CHR|6|34|「你的百姓若奉你的派遣出去，無論往何處與仇敵爭戰，他們若向你所選擇的這城和我為你名所建造的殿禱告，
2CHR|6|35|求你從天上垂聽他們的禱告祈求，為他們伸張正義。
2CHR|6|36|「你的百姓若得罪你，因為沒有人不犯罪，你向他們發怒，把他們交在仇敵面前，擄他們的人把他們帶到或遠或近之地；
2CHR|6|37|他們若在被擄之地那裏回心轉意，在被擄之地悔改，向你懇求說：『我們有罪了，我們悖逆了，我們作惡了』；
2CHR|6|38|他們若在被擄之地盡心盡性歸向你，又向自己的地，就是你賜給他們列祖的地和你所選擇的城，以及我為你名所建造的這殿禱告，
2CHR|6|39|求你從天上你的居所垂聽他們的禱告祈求，為他們伸張正義，赦免你的百姓向你犯的罪。
2CHR|6|40|我的上帝啊，現在求你睜眼看，側耳聽在此處所獻的禱告。
2CHR|6|41|「耶和華上帝啊，現在求你興起， 與你有能力的約櫃同入安歇之所。 耶和華上帝啊，願你的祭司披上救恩， 願你的聖民蒙福歡樂。
2CHR|6|42|耶和華上帝啊，求你不要厭棄你的受膏者， 要記得向你僕人 大衛 所施的慈愛。」
2CHR|7|1|所羅門 祈禱完畢，就有火從天降下來，燒盡燔祭和祭物。耶和華的榮光充滿了殿；
2CHR|7|2|因耶和華的榮光充滿了耶和華的殿，所以祭司不能進耶和華的殿。
2CHR|7|3|那火降下、耶和華的榮光在殿上的時候， 以色列 眾人看見，就在石板地俯伏敬拜，稱謝耶和華： 「耶和華本為善， 他的慈愛永遠長存！」
2CHR|7|4|王和眾百姓在耶和華面前獻祭。
2CHR|7|5|所羅門 王獻二萬二千頭牛，十二萬隻羊為祭。這樣，王和眾百姓為上帝的殿行了奉獻之禮。
2CHR|7|6|祭司各供其職侍立， 利未 人拿著耶和華的樂器，就是 大衛 王所造、為要頌讚耶和華的樂器，因他的慈愛永遠長存；他們為 大衛 的讚美詩奏樂；祭司在眾人面前吹號， 以色列 眾人都站立。
2CHR|7|7|所羅門 因他所造的銅壇容不下燔祭、素祭和脂肪，就將耶和華殿前院子的中間分別為聖，在那裏獻燔祭和平安祭牲的脂肪。
2CHR|7|8|那時 所羅門 守節七日，從 哈馬口 直到 埃及 溪谷的 以色列 眾人都與他同在一起，成了一個極其盛大的會。
2CHR|7|9|第八日他們舉行嚴肅會，行奉獻壇的禮七日，守節七日。
2CHR|7|10|七月二十三日，王差遣百姓回自己的帳棚去；他們為耶和華向 大衛 和 所羅門 ，以及他百姓 以色列 所施的恩惠，心裏都歡喜快樂。
2CHR|7|11|所羅門 建完了耶和華的殿和王宮；在耶和華的殿和王宮的工程上，凡他心中所要做的，都順利做成了。
2CHR|7|12|夜間耶和華向 所羅門 顯現，對他說：「我已聽了你的禱告，也選擇這地方歸我作獻祭的殿宇。
2CHR|7|13|我若使天閉塞不下雨，或使蝗蟲吃這地的出產，或降瘟疫在我子民中，
2CHR|7|14|這稱為我名下的子民，若是謙卑自己，禱告，尋求我的面，轉離他們的惡行，我必從天上垂聽，赦免他們的罪，醫治他們的地。
2CHR|7|15|我必睜眼看，側耳聽在此處所獻的禱告。
2CHR|7|16|現在我已選擇這殿，分別為聖，使我的名永在其中；我的眼、我的心也必時常在那裏。
2CHR|7|17|你若行在我面前，效法你父 大衛 所行的，遵行我一切所吩咐你的，謹守我的律例典章，
2CHR|7|18|我就必堅固你國度的王位，正如我與你父 大衛 所立的約，說：『你的子孫必不斷有人治理 以色列 。』
2CHR|7|19|「倘若你們轉去，離棄我擺在你們面前的律例誡命，去事奉別神，敬拜它們，
2CHR|7|20|我就必把 以色列 人從我賜給他們的地上連根拔起，也必從我面前捨棄那為我名所分別為聖的殿，使它在萬民中成為笑柄，被人譏誚。
2CHR|7|21|這殿雖然崇高，將來凡經過的人必驚訝說：『耶和華為何向這地和這殿如此行呢？』
2CHR|7|22|人必說：『因為此地的人離棄領他們祖先出 埃及 地的耶和華－他們的上帝，去親近別神，敬拜事奉它們，所以耶和華使這一切災禍臨到他們。』」
2CHR|8|1|所羅門 建造耶和華的殿和王宮，用了二十年才完成。
2CHR|8|2|所羅門 修築 希蘭 送給他的城鎮，使 以色列 人住在那裏。
2CHR|8|3|所羅門 往 哈馬‧瑣巴 去，攻取了那地方。
2CHR|8|4|所羅門 建造曠野的 達莫 ，建造 哈馬 一切的儲貨城，
2CHR|8|5|又建造 上伯‧和崙 、 下伯‧和崙 ，成為有牆、門、閂的堡壘城。
2CHR|8|6|所羅門 建造 巴拉 和一切的儲貨城、戰車城、戰馬城，以及他所想要建造的，在 耶路撒冷 、 黎巴嫩 ，和自己所治理全國中的一切建設。
2CHR|8|7|至於所有剩下的百姓，不屬 以色列 的 赫 人、 亞摩利 人、 比利洗 人、 希未 人、 耶布斯 人，
2CHR|8|8|那些 以色列 人在當地不能滅盡的人， 所羅門 徵召他們剩下的後代服勞役，直到今日。
2CHR|8|9|惟有 以色列 人， 所羅門 不使他們當奴僕做工，而是作他的戰士、軍官、戰車長、騎兵長。
2CHR|8|10|這些是 所羅門 王的監工，共有二百五十名百姓的監工。
2CHR|8|11|所羅門 把法老的女兒遷出 大衛城 ，上到他為她建造的宮裏，因 所羅門 說：「耶和華約櫃所到之處都是聖地，所以我的妻子不可住在 以色列 王 大衛 的宮裏。」
2CHR|8|12|那時， 所羅門 在走廊前他所築的耶和華的壇上，向耶和華獻燔祭，
2CHR|8|13|又遵照 摩西 的吩咐，在安息日、初一，以及每年在除酵節、七七節、住棚節三個節期，獻每日所當獻上的祭。
2CHR|8|14|所羅門 照著他父親 大衛 所定的條例，分派祭司的班次，擔任他們的職務，又分派 利未 人的任務，負責頌讚，並在祭司面前做每日當做的事，又派門口的守衛按著班次看守各門，因為神人 大衛 是這樣吩咐的。
2CHR|8|15|王對眾祭司和 利未 人的吩咐，無論是管理庫房或任何事務，他們都不違背。
2CHR|8|16|所羅門 所有的工作都準備就緒，從立耶和華殿的根基直到完工的日子。耶和華的殿就完成了。
2CHR|8|17|那時， 所羅門 往 以東 地海岸的 以旬‧迦別 和 以祿 去。
2CHR|8|18|希蘭 派他的臣僕，把船隻和熟悉航海的僕人送到 所羅門 那裏。他們同 所羅門 的僕人到了 俄斐 ，從那裏得了四百五十他連得金子，運到 所羅門 王那裏。
2CHR|9|1|示巴 女王聽見 所羅門 的名聲，就來到 耶路撒冷 ，要用難題考問 所羅門 。她帶著很多的隨從，有駱駝馱著香料、許多金子和寶石。她來到 所羅門 那裏，向他提出心中所有的問題。
2CHR|9|2|所羅門 回答了她所有的問題，沒有一個問題太難，是 所羅門 不能向她解答的。
2CHR|9|3|示巴 女王看見 所羅門 的智慧和他所建造的宮殿，
2CHR|9|4|席上的食物，坐著的群臣，侍立的僕人和他們的服裝，司酒長和他們的服裝，以及他上耶和華殿的臺階 ，就詫異得神不守舍。
2CHR|9|5|她對王說：「我在本國所聽到的話，論到你的事和你的智慧是真的！
2CHR|9|6|我本來不信那些話，及至我來親眼看見了，看哪，人所告訴我的，還不及你豐富智慧的一半，超過我所聽見的傳聞。
2CHR|9|7|你的人是有福的！你這些常侍立在你面前、聽你智慧話的僕人是有福的！
2CHR|9|8|耶和華－你的上帝是應當稱頌的！他喜愛你，使你坐他的王位，為耶和華－你的上帝作王；因為你的上帝愛 以色列 ，要永遠堅立它，所以立你作他們的王，使你秉公行義。」
2CHR|9|9|於是 示巴 女王把一百二十他連得金子、極多的香料和寶石送給 所羅門 王；從來沒有像 示巴 女王送給 所羅門 王那麼多的香料。
2CHR|9|10|希蘭 的僕人和 所羅門 的僕人也從 俄斐 運了金子來，又運了檀香木和寶石來。
2CHR|9|11|王用檀香木為耶和華的殿和王宮做階梯，又為歌唱的人做琴瑟； 猶大 地從來沒有見過這樣的。
2CHR|9|12|所羅門 王除了回贈 示巴 女王所帶來的，凡她所提出的一切要求， 所羅門 王都送給她。於是女王和她臣僕轉回，到本國去了。
2CHR|9|13|所羅門 每年所得的金子，重六百六十六他連得，
2CHR|9|14|另外還有從商人和貿易所收到的，以及 阿拉伯 諸王和各地的省長進貢給 所羅門 的金銀。
2CHR|9|15|所羅門 王用錘出來的金子打成二百面盾牌，每面盾牌用六百舍客勒錘出來的金子；
2CHR|9|16|又用錘出來的金子打成三百面小盾牌，每面小盾牌用三百舍客勒金子。王把它們放在 黎巴嫩林宮 裏。
2CHR|9|17|王又製造一個大的象牙寶座，包上純金。
2CHR|9|18|寶座有六層臺階，又有金腳凳，與寶座相連。座位之處兩旁有扶手，靠近扶手有兩隻獅子站立。
2CHR|9|19|六層臺階上有十二隻獅子站立，分站左邊和右邊；任何國度都沒有這樣做的。
2CHR|9|20|所羅門 王一切的飲器都是金的， 黎巴嫩林宮 裏所有的器皿都是純金的。在 所羅門 的日子，銀子算不了甚麼。
2CHR|9|21|因王的船隻與 希蘭 的僕人一同往 他施 去， 他施 船隻每三年一次把金、銀、象牙、猿猴、孔雀 運回來。
2CHR|9|22|所羅門 王的財寶與智慧勝過地上的眾王。
2CHR|9|23|地上的眾王都求見 所羅門 的面，要聽上帝放在他心裏的智慧。
2CHR|9|24|他們各帶貢物，就是銀器、金器、衣服、兵器、香料、馬、騾子，每年都有一定的數量。
2CHR|9|25|所羅門 擁有給戰車和馬用的四千個棚子，還有一萬二千名騎兵，安置在屯車城，在 耶路撒冷 的王那裏。
2CHR|9|26|所羅門 統管諸王，從 大河 到 非利士 人的地，直到 埃及 的邊界。
2CHR|9|27|王在 耶路撒冷 使銀子多如石頭，香柏木多如 謝非拉 的桑樹。
2CHR|9|28|有人從 埃及 和各國為 所羅門 把馬匹運來。
2CHR|9|29|所羅門 其餘的事，自始至終，不都寫在 拿單 先知的書上和 示羅 人 亞希雅 的《預言書》上，以及 易多 先見論 尼八 兒子 耶羅波安 的《默示書》上嗎？
2CHR|9|30|所羅門 在 耶路撒冷 作全 以色列 的王四十年。
2CHR|9|31|所羅門 與他祖先同睡，葬在他父親 大衛 的城裏，他兒子 羅波安 接續他作王。
2CHR|10|1|羅波安 往 示劍 去，因 以色列 眾人都到了 示劍 ，要立他作王。
2CHR|10|2|尼八 的兒子 耶羅波安 先前躲避 所羅門 王，逃往 埃及 ，住在那裏；他聽見這事，就從 埃及 回來。
2CHR|10|3|以色列 人派人去請他來。 耶羅波安 就和 以色列 眾人來，與 羅波安 談話，說：
2CHR|10|4|「你父親使我們負重軛，現在求你減輕你父親所加給我們的苦工和重軛，我們就服事你。」
2CHR|10|5|羅波安 對他們說：「過三天再來見我吧！」百姓就走了。
2CHR|10|6|羅波安 的父親 所羅門 在世的時候，有侍立在他面前的長者， 羅波安 王和他們商議，說：「你們出個主意，好把話帶回給這百姓。」
2CHR|10|7|他們對他說：「王若恩待這百姓，使他們喜悅，跟他們說好話，他們就永遠作王的僕人了。」
2CHR|10|8|王不採納長者給他出的主意，卻和那些與他一同長大、在他面前侍立的年輕人商議。
2CHR|10|9|他對他們說：「這百姓對我說：『你父親使我們負重軛，求你減輕一些。』你們出個甚麼主意，我們好把話帶回給他們。」
2CHR|10|10|那些與他一同長大的年輕人對他說：「這些百姓對王說：『你父親使我們負重軛，求你給我們減輕一些。』王要對他們如此說：『我的小指頭比我父親的腰還粗呢！
2CHR|10|11|我父親使你們負重軛，現在我必使你們負更重的軛！我父親用鞭子懲罰你們，我卻要用蠍子！』」
2CHR|10|12|耶羅波安 和眾百姓遵照王所說「你們第三天再來見我」的話，第三天來到 羅波安 那裏。
2CHR|10|13|王嚴厲地回答他們。 羅波安 王不採納長者所出的主意，
2CHR|10|14|卻照著年輕人所出的主意對他們說：「我 使你們負重軛，我必使你們負更重的軛！我父親用鞭子懲罰你們，我卻要用蠍子！」
2CHR|10|15|王不依從百姓，因這事件是出於上帝，為要應驗耶和華藉 示羅 人 亞希雅 對 尼八 的兒子 耶羅波安 所說的話。
2CHR|10|16|以色列 眾人見王不依從他們，百姓就回覆王說： 「我們在 大衛 中有甚麼分呢？ 我們在 耶西 的兒子中沒有產業！ 以色列 啊，各回自己的帳棚去吧！ 大衛 啊，現在你顧自己的家吧！」 於是， 以色列 眾人都回自己的帳棚去了；
2CHR|10|17|至於住 猶大 城鎮的 以色列 人， 羅波安 仍作他們的王。
2CHR|10|18|羅波安 王派監管勞役的 哈多蘭 去， 以色列 人用石頭打他，他就死了。 羅波安 王急忙上車，逃回 耶路撒冷 去了。
2CHR|10|19|這樣， 以色列 背叛 大衛 家，直到今日。
2CHR|11|1|羅波安 來到 耶路撒冷 ，召集 猶大 家和 便雅憫 家，共十八萬人，都是精選的戰士，要與 以色列 爭戰，好將國奪回再歸自己。
2CHR|11|2|但耶和華的話臨到神人 示瑪雅 ，說：
2CHR|11|3|「你去告訴 所羅門 的兒子 猶大 王 羅波安 和住 猶大 、 便雅憫 的 以色列 眾人，說：
2CHR|11|4|『耶和華如此說：你們不可上去與你們的弟兄爭戰。各自回家去吧！因為這事是出於我。』」眾人就聽從耶和華的話回去，不去與 耶羅波安 爭戰。
2CHR|11|5|羅波安 住在 耶路撒冷 ，在 猶大 為防禦修築城鎮，
2CHR|11|6|他修築 伯利恆 、 以坦 、 提哥亞 、
2CHR|11|7|伯‧夙 、 梭哥 、 亞杜蘭 、
2CHR|11|8|迦特 、 瑪利沙 、 西弗 、
2CHR|11|9|亞多萊音 、 拉吉 、 亞西加 、
2CHR|11|10|瑣拉 、 亞雅崙 、 希伯崙 。這都是 猶大 和 便雅憫 的堅固城。
2CHR|11|11|羅波安 又鞏固這些堡壘，在其中安置軍官，儲備糧食、油和酒。
2CHR|11|12|他在各城裏預備盾牌和槍，使城極其堅固。 猶大 和 便雅憫 都歸了他。
2CHR|11|13|全 以色列 的祭司和 利未 人都從四方來歸 羅波安 。
2CHR|11|14|利未 人放棄他們的郊野和產業，來到 猶大 與 耶路撒冷 ，因為 耶羅波安 和他的兒子拒絕他們，不許他們擔任祭司事奉耶和華。
2CHR|11|15|耶羅波安 為丘壇，為山羊鬼魔，為自己所造的牛犢設立祭司。
2CHR|11|16|以色列 各支派中，凡立定心意尋求耶和華－ 以色列 上帝的，都隨從 利未 人來到 耶路撒冷 獻祭給耶和華－他們列祖的上帝。
2CHR|11|17|這就鞏固了 猶大 王國，使 所羅門 的兒子 羅波安 強盛三年，因為這三年他們遵行 大衛 和 所羅門 的道。
2CHR|11|18|羅波安 娶 大衛 兒子 耶利末 的女兒 瑪哈拉 為妻，又娶 耶西 兒子 以利押 的女兒 亞比孩 為妻，
2CHR|11|19|從她生了幾個兒子，就是 耶烏施 、 示瑪利雅 和 撒罕 。
2CHR|11|20|後來他又娶 押沙龍 的女兒 瑪迦 ，從她生了 亞比雅 、 亞太 、 細撒 和 示羅密 。
2CHR|11|21|羅波安 有十八個妻和六十個妾，生了二十八個兒子，六十個女兒；他卻愛 押沙龍 的女兒 瑪迦 ，過於愛其他的妻妾。
2CHR|11|22|羅波安 立 瑪迦 的兒子 亞比雅 作太子，在他兄弟中為首，因為要立他作王。
2CHR|11|23|羅波安 辦事精明，把他眾兒子分散在 猶大 和 便雅憫 全地各堅固城裏，賜他們大量的糧食，又給他們娶許多妻子。
2CHR|12|1|羅波安 的王國穩固，他強盛的時候就離棄耶和華的律法，全 以色列 都跟從他。
2CHR|12|2|羅波安 王第五年， 埃及 王 示撒 上來攻打 耶路撒冷 ，因為他們背叛了耶和華。
2CHR|12|3|示撒 帶著一千二百輛戰車，六萬名騎兵，以及跟隨他從 埃及 出來的 路比 人、 蘇基 人和 古實 人的軍隊，多得不可勝數。
2CHR|12|4|他攻取了 猶大 的堅固城，來到 耶路撒冷 。
2CHR|12|5|那時， 猶大 的領袖因為 示撒 的緣故聚集在 耶路撒冷 ，有先知 示瑪雅 去見 羅波安 和眾領袖，對他們說：「耶和華如此說：『你們離棄了我，所以我也離棄你們，把你們交在 示撒 手裏。』」
2CHR|12|6|於是 以色列 的領袖和王都謙卑說：「耶和華是公義的。」
2CHR|12|7|耶和華見他們謙卑，耶和華的話就臨到 示瑪雅 ，說：「他們既謙卑，我必不滅絕他們；我要使他們暫時得拯救，不藉著 示撒 的手將我的怒氣倒在 耶路撒冷 。
2CHR|12|8|然而他們必作 示撒 的僕人，好叫他們知道，服事我與服事地上邦國有何分別。」
2CHR|12|9|於是， 埃及 王 示撒 上來攻取 耶路撒冷 ，奪了耶和華殿和王宮裏的寶物，盡都帶走，又奪走 所羅門 製造的金盾牌。
2CHR|12|10|羅波安 王製造銅盾牌代替那些金盾牌，交給看守王宮宮門的護衛長看管。
2CHR|12|11|每逢王進耶和華的殿，護衛兵就來，舉起這些盾牌；隨後仍將盾牌送回護衛室。
2CHR|12|12|王謙卑的時候，耶和華的怒氣就轉消了，不全然滅盡，並且在 猶大 中，情況也有好轉。
2CHR|12|13|羅波安 王自強，在 耶路撒冷 作王。他登基的時候年四十一歲，在 耶路撒冷 ，就是耶和華從 以色列 眾支派中所選擇立他名的城，作王十七年。 羅波安 的母親名叫 拿瑪 ，是 亞捫 人。
2CHR|12|14|羅波安 行惡，因他沒有立定心意尋求耶和華。
2CHR|12|15|羅波安 的事蹟，自始至終不都寫在 示瑪雅 先知和 易多 先見的《史記》上嗎？ 羅波安 與 耶羅波安 時常交戰。
2CHR|12|16|羅波安 與他祖先同睡，葬在 大衛城 ，他的兒子 亞比雅 接續他作王。
2CHR|13|1|耶羅波安 王十八年， 亞比雅 登基作 猶大 王，
2CHR|13|2|在 耶路撒冷 作王三年。他母親名叫 米該亞 ，是 基比亞 人 烏列 的女兒 。 亞比雅 常與 耶羅波安 交戰。
2CHR|13|3|有一次 亞比雅 率領四十萬精選的士兵出戰，他們都是勇敢的戰士； 耶羅波安 也率領八十萬精選的大能勇士，迎著 亞比雅 擺陣。
2CHR|13|4|亞比雅 站在 以法蓮 山區中的 洗瑪臉山 上，說：「 耶羅波安 和 以色列 眾人哪，要聽我說！
2CHR|13|5|耶和華－ 以色列 的上帝曾立鹽約，將 以色列 國永遠賜給 大衛 和他的子孫，你們不知道嗎？
2CHR|13|6|但 大衛 兒子 所羅門 的臣僕、 尼八 的兒子 耶羅波安 起來背叛他的主人。
2CHR|13|7|有些無賴的歹徒聚集跟從他，逞強攻擊 所羅門 的兒子 羅波安 ；那時 羅波安 還年輕，心志軟弱，不能抵擋他們。
2CHR|13|8|「現在你們說要抗拒 大衛 子孫手下所治理的耶和華的國，你們的人數眾多，你們那裏又有 耶羅波安 為你們所造當作神明的金牛犢。
2CHR|13|9|你們不是驅逐耶和華的祭司 亞倫 的後裔和 利未 人嗎？不是照著外邦人的惡俗為自己立祭司嗎？無論何人牽一頭公牛犢、七隻公綿羊將自己分別出來，就可作虛無神明的祭司。
2CHR|13|10|至於我們，耶和華是我們的上帝，我們並沒有離棄他。我們有事奉耶和華的祭司，都是 亞倫 的後裔，並有 利未 人各盡其職。
2CHR|13|11|他們每日早晚向耶和華獻燔祭，燒芬芳的香，又在純金的 供桌上擺供餅，每晚點燃金燈臺上的燈盞，因為我們遵守耶和華－我們上帝的命令，但你們卻離棄了他。
2CHR|13|12|看哪，率領我們的是上帝，又有他的祭司拿號向你們吹出響聲。 以色列 人哪，不要與耶和華－你們列祖的上帝爭戰，因你們必不能得勝。」
2CHR|13|13|耶羅波安 卻在 猶大 人的後頭設伏兵。這樣， 以色列 人在 猶大 人的前頭，伏兵在 猶大 人的後頭。
2CHR|13|14|猶大 人轉過來，看哪，前後都有戰事，就呼求耶和華，祭司也吹號。
2CHR|13|15|於是 猶大 人吶喊。 猶大 人吶喊的時候，上帝就擊打 耶羅波安 和 以色列 眾人，使他們敗在 亞比雅 與 猶大 人面前。
2CHR|13|16|以色列 人在 猶大 人面前逃跑，上帝將他們交在 猶大 人手裏。
2CHR|13|17|亞比雅 和他的軍兵大大擊殺 以色列 人， 以色列 人被殺仆倒的精兵有五十萬。
2CHR|13|18|那時， 以色列 人被制伏了。 猶大 人得勝，因為他們倚靠耶和華－他們列祖的上帝。
2CHR|13|19|亞比雅 追趕 耶羅波安 ，攻取了他的幾座城，就是 伯特利 和所屬的鄉鎮 ， 耶沙拿 和所屬的鄉鎮， 以法拉音 和所屬的鄉鎮。
2CHR|13|20|亞比雅 在世的時候， 耶羅波安 不再強盛；耶和華擊打他，他就死了。
2CHR|13|21|亞比雅 卻漸漸強盛。他娶了十四個妻妾，生了二十二個兒子，十六個女兒。
2CHR|13|22|亞比雅 其餘的事和他的言行都寫在 易多 先知的評傳上。
2CHR|14|1|亞比雅 與他祖先同睡，葬在 大衛城 ，他的兒子 亞撒 接續他作王。 亞撒 在位期間，國中太平十年。
2CHR|14|2|亞撒 行耶和華－他上帝眼中看為善為正的事，
2CHR|14|3|除掉外邦的祭壇和丘壇，打碎柱像，砍下 亞舍拉 ，
2CHR|14|4|吩咐 猶大 人尋求耶和華－他們列祖的上帝，遵行他的律法和誡命，
2CHR|14|5|又在 猶大 各城鎮除掉丘壇和香壇。在他治理下，國中太平。
2CHR|14|6|他在 猶大 建造了幾座堅固城。那些年間，國中太平，沒有戰爭，因為耶和華賜他平安。
2CHR|14|7|他對 猶大 人說：「我們要建造這些城鎮，四圍築牆，蓋城樓，安門，做閂；地仍屬於我們，因為我們尋求耶和華－我們的上帝；我們尋求他，他就賜我們四境平安。」於是他們建造城鎮，諸事亨通。
2CHR|14|8|亞撒 的軍兵，出自 猶大 拿盾牌拿槍的三十萬人，出自 便雅憫 拿小盾牌拉弓的二十八萬人；這些全都是大能的勇士。
2CHR|14|9|古實 人 謝拉 率領一百萬軍兵，三百輛戰車，出來攻擊 猶大 人，到了 瑪利沙 。
2CHR|14|10|亞撒 出去迎戰，在 瑪利沙 的 洗法谷 彼此擺陣。
2CHR|14|11|亞撒 呼求耶和華－他的上帝說：「耶和華啊，在強弱之間，惟有你能幫助。耶和華－我們的上帝啊，求你幫助我們，因為我們仰賴你，奉你的名來抵擋這大軍。耶和華啊，你是我們的上帝，不要讓人勝過你。」
2CHR|14|12|於是耶和華擊打 古實 人，使他們敗在 亞撒 和 猶大 人面前， 古實 人就逃跑了。
2CHR|14|13|亞撒 和跟隨他的軍兵追趕他們，直到 基拉耳 。 古實 人被殺的很多，無法復原，因為他們在耶和華與他軍兵面前被擊潰。 猶大 人奪了許多財物，
2CHR|14|14|又攻打 基拉耳 四圍一切的城鎮；城中的人都懼怕耶和華。 猶大 人擄掠了一切的城鎮，因其中的財物很多，
2CHR|14|15|又毀壞了群畜的圈，奪取許多的羊和駱駝，就回 耶路撒冷 去了。
2CHR|15|1|上帝的靈臨到 俄德 的兒子 亞撒利雅 。
2CHR|15|2|他出來迎接 亞撒 ，對他說：「 亞撒 ， 猶大 和 便雅憫 眾人哪，要聽我說：你們若順從耶和華，耶和華必與你們同在；你們若尋求他，就必尋見；你們若離棄他，他必離棄你們。
2CHR|15|3|以色列 人不信真神，沒有訓誨的祭司，也沒有律法，已經許多日子了。
2CHR|15|4|但他們在急難的時候歸向耶和華－ 以色列 的上帝，尋求他，他就被他們尋見。
2CHR|15|5|那時，出入的人不得平安，各地的居民都遭大亂；
2CHR|15|6|他們被破壞殆盡，這國攻擊那國，這城攻擊那城，因為上帝用各樣災難擾亂他們。
2CHR|15|7|現在你們要剛強，不要手軟，因你們所行的必得賞賜。」
2CHR|15|8|亞撒 聽見這些話和 俄德 先知的預言，就壯起膽來，在 猶大 和 便雅憫 全地，以及 以法蓮 山區所奪的各城，把其中的可憎之物盡都除掉，又在耶和華殿的走廊前重新修築耶和華的壇。
2CHR|15|9|他又召集 猶大 和 便雅憫 眾人，以及他們中間寄居的 以法蓮 人、 瑪拿西 人、 西緬 人。有許多 以色列 人歸順 亞撒 ，因為他們看見耶和華－他的上帝與他同在。
2CHR|15|10|亞撒 作王第十五年三月，他們都聚集在 耶路撒冷 。
2CHR|15|11|那日他們從所取的擄物中，將七百頭牛和七千隻羊獻給耶和華。
2CHR|15|12|他們立約，要盡心盡性尋求耶和華－他們列祖的上帝。
2CHR|15|13|凡不尋求耶和華－ 以色列 上帝的，無論大小、男女，必被處死。
2CHR|15|14|他們就大聲歡呼，吹號吹角，向耶和華起誓。
2CHR|15|15|猶大 眾人為所起的誓歡喜，因他們盡心起誓，盡意尋求耶和華，耶和華就被他們尋見，且賜他們四境平安。
2CHR|15|16|亞撒 王甚至廢了他祖母 瑪迦 太后的位，因 瑪迦 造了可憎的 亞舍拉 。 亞撒 砍下她的偶像，搗得粉碎，在 汲淪溪 邊燒了，
2CHR|15|17|只是丘壇還沒有從 以色列 中廢去，然而 亞撒 一生有純正的心。
2CHR|15|18|亞撒 將他父親所分別為聖與自己所分別為聖的金銀和器皿都奉到上帝的殿裏。
2CHR|15|19|亞撒 作王直到第三十五年，都沒有戰事。
2CHR|16|1|亞撒 作王第三十六年， 以色列 王 巴沙 上來攻擊 猶大 ，修築 拉瑪 ，不許人從 猶大 王 亞撒 那裏出入。
2CHR|16|2|於是 亞撒 從耶和華殿和王宮的府庫裏拿出金銀來，送給住在 大馬士革 的 亞蘭 王 便‧哈達 ，說：
2CHR|16|3|「你父曾與我父立約，我與你也要這樣立約。看哪，我把金銀送給你，請你廢掉你與 以色列 王 巴沙 所立的約，使他從我這裏撤退。」
2CHR|16|4|便‧哈達 聽從了 亞撒 王，就派遣他的軍官去攻打 以色列 的城鎮。他們攻下了 以雲 、 但 、 亞伯‧瑪音 和 拿弗他利 一切的儲貨城。
2CHR|16|5|巴沙 聽見了，就停工不修築 拉瑪 ，任由他的工程停止。
2CHR|16|6|於是 亞撒 王率領 猶大 眾人，運走 巴沙 修築 拉瑪 所用的石頭和木料，用以修築 迦巴 和 米斯巴 。
2CHR|16|7|那時， 哈拿尼 先見來見 猶大 王 亞撒 ，對他說：「因你仰賴 亞蘭 王，沒有仰賴耶和華－你的上帝，所以 亞蘭 王的軍兵逃脫了你的手。
2CHR|16|8|古實 人和 路比 人的軍隊不是非常強大嗎？他們的戰車騎兵不是極多嗎？只因你仰賴耶和華，他就將他們交在你手裏。
2CHR|16|9|因為耶和華的眼目遍察全地，要堅固向他存純正之心的人。你在這事上行得愚昧；因此，以後你必有戰爭。」
2CHR|16|10|亞撒 惱恨先見，為了這事向他發怒，將他囚在監裏。那時 亞撒 也虐待一些百姓。
2CHR|16|11|亞撒 自始至終的事蹟，看哪，都寫在《猶大和以色列諸王記》上。
2CHR|16|12|亞撒 作王三十九年的時候患了腳疾，非常嚴重。他生病的時候沒有求耶和華，只求醫生。
2CHR|16|13|他作王四十一年死了，與他祖先同睡，
2CHR|16|14|葬在 大衛城 自己所鑿的墳墓裏。人把他放在床上，床上堆滿各樣馨香的香料，就是按做香的作法調和的香料，又為他生一堆大火誌哀。
2CHR|17|1|亞撒 的兒子 約沙法 接續他作王，奮勇自強，防備 以色列 。
2CHR|17|2|他安置軍兵在 猶大 一切堅固城裏，又安置駐軍在 猶大 地和他父親 亞撒 所得 以法蓮 的城鎮中。
2CHR|17|3|耶和華與 約沙法 同在，因為他行他祖先 大衛 從前所行的道，不去尋求諸 巴力 ，
2CHR|17|4|只尋求他父親的上帝，遵行他的誡命，不效法 以色列 人的行為。
2CHR|17|5|所以耶和華堅定 約沙法 手中的國， 猶大 眾人給他進貢； 約沙法 大有財富和尊榮。
2CHR|17|6|他樂意遵行耶和華的道，並且從 猶大 再次除掉一切丘壇和 亞舍拉 。
2CHR|17|7|他作王第三年，差遣官員 便‧亥伊勒 、 俄巴底 、 撒迦利雅 、 拿坦業 、 米該亞 往 猶大 各城去教導百姓。
2CHR|17|8|跟他們一同去的有 利未 人 示瑪雅 、 尼探雅 、 西巴第雅 、 亞撒黑 、 示米拉末 、 約拿單 、 亞多尼雅 、 多比雅 、 駝‧巴多尼雅 ；跟他們一同的又有 以利沙瑪 和 約蘭 二位祭司。
2CHR|17|9|他們在 猶大 教導，帶著耶和華的律法書，走遍 猶大 各城教導百姓。
2CHR|17|10|猶大 四圍地上的邦國都懼怕耶和華，不敢與 約沙法 爭戰。
2CHR|17|11|有些 非利士 人送禮物，進貢銀子給 約沙法 。 阿拉伯 人也送他七千七百隻公綿羊，七千七百隻公山羊。
2CHR|17|12|約沙法 日漸強大，他在 猶大 建造堡壘和儲貨城。
2CHR|17|13|他在 猶大 城鎮中有許多工程，在 耶路撒冷 又有戰士，就是大能的勇士。
2CHR|17|14|他們按著父家的數目如下： 猶大 族的千夫長以 押拿 為首，率領三十萬大能的勇士；
2CHR|17|15|其次是 約哈難 千夫長，率領二十八萬；
2CHR|17|16|其次是 細基利 的兒子 亞瑪斯雅 ，他是一個自願奉獻給耶和華的人，率領二十萬大能的勇士。
2CHR|17|17|便雅憫 族有大能的勇士 以利雅大 ，率領二十萬拿弓箭和盾牌的人；
2CHR|17|18|其次是 約薩拔 ，率領十八萬預備打仗的人。
2CHR|17|19|這些都是伺候王的，還有王在全 猶大 的堅固城所安置的不在其內。
2CHR|18|1|約沙法 大有財富和尊榮，他與 亞哈 結親。
2CHR|18|2|過了幾年，他下到 撒瑪利亞 去見 亞哈 ； 亞哈 為他和跟從他的人宰了許多牛羊，勸他一同上去攻打 基列 的 拉末 。
2CHR|18|3|以色列 王 亞哈 問 猶大 王 約沙法 說：「你肯同我去攻打 基列 的 拉末 嗎？」他回答說：「你我不分彼此，我的軍隊就是你的軍隊，我們必與你一同去爭戰。」
2CHR|18|4|約沙法 對 以色列 王說：「請你先求問耶和華的話。」
2CHR|18|5|於是 以色列 王召集先知四百人，問他們說：「我可以上去攻打 基列 的 拉末 嗎？還是不要上去呢？」他們說：「可以上去，因為上帝必將那城交在王的手裏。」
2CHR|18|6|約沙法 說：「這裏還有沒有耶和華的先知，我們好求問他呢？」
2CHR|18|7|以色列 王對 約沙法 說：「還有一個人，是 音拉 的兒子 米該雅 ，我們可以託他求問耶和華。只是我真的很恨他，因為他對我說預言，從不說吉言，總是說凶信。」 約沙法 說：「請王不要這麼說。」
2CHR|18|8|以色列 王就召了一個官員來，說：「你快去，把 音拉 的兒子 米該雅 召來。」
2CHR|18|9|以色列 王和 猶大 王 約沙法 在 撒瑪利亞 城門前的禾場，各穿朝服，坐在寶座上，所有的先知都在他們面前說預言。
2CHR|18|10|基拿拿 的兒子 西底家 為自己造了鐵角，說：「耶和華如此說：『你要用這些角牴觸 亞蘭 人，直到將他們滅盡。』」
2CHR|18|11|所有的先知也都這樣預言說：「可以上 基列 的 拉末 去，必然得勝，因為耶和華必將那城交在王的手中。」
2CHR|18|12|那去召 米該雅 的使者對他說：「看哪，眾先知都異口同聲向王說吉言，你也跟他們說一樣的話，說吉言吧！」
2CHR|18|13|米該雅 說：「我指著永生的耶和華起誓，我的上帝說甚麼，我就說甚麼。」
2CHR|18|14|米該雅 來到王那裏，王問他：「 米該雅 啊，我們可以上去攻打 基列 的 拉末 嗎？還是不要上去呢？」他說：「可以上去，必然得勝，敵人必交在你們手裏。」
2CHR|18|15|王對他說：「我要你發誓多少次，你才會奉耶和華的名向我說實話呢？」
2CHR|18|16|米該雅 說：「我看見 以色列 眾人散佈在山上，如同沒有牧人的羊群一般。耶和華說：『這些人沒有主人，他們可以平安地各自回家去。』」
2CHR|18|17|以色列 王對 約沙法 說：「我豈沒有告訴你，這人對我說預言，從不說吉言，只說凶信嗎？」
2CHR|18|18|米該雅 說：「因此你們要聽耶和華的話！我看見耶和華坐在寶座上，天上的萬軍侍立在他左右。
2CHR|18|19|耶和華 說：『誰去引誘 以色列 王 亞哈 上 基列 的 拉末 去陣亡呢？』這個這樣說，那個那樣說。
2CHR|18|20|隨後有一個靈出來，站在耶和華面前，說：『我去引誘他。』耶和華問他：『用甚麼方法呢？』
2CHR|18|21|他說：『我要出去，在他眾先知的口中成為謊言的靈。』耶和華說：『這樣，你去引誘他，必能成功。你出去，照樣做吧！』
2CHR|18|22|現在，看哪，耶和華使謊言的靈入了你的這些先知的口，並且耶和華已經宣告要降禍於你。」
2CHR|18|23|基拿拿 的兒子 西底家 前來打 米該雅 一巴掌，說：「耶和華的靈從哪裏離開我向你說話呢？」
2CHR|18|24|米該雅 說：「看哪，你進入嚴密的內室躲藏的那日，就必看見。」
2CHR|18|25|以色列 王說：「把 米該雅 帶走，交回給 亞們 市長和 約阿施 王子。
2CHR|18|26|你們要說：『王如此說：把這個人關在監獄裏，使他受苦，吃不飽喝不足，直等到我平安回來。』」
2CHR|18|27|米該雅 說：「你若真的能平安回來，那就是耶和華沒有藉我說話了。」他又說：「眾百姓啊，你們都要聽！」
2CHR|18|28|以色列 王和 猶大 王 約沙法 上 基列 的 拉末 去。
2CHR|18|29|以色列 王對 約沙法 說：「我要改裝上陣，你可以仍穿王服。」於是 以色列 王改裝，他們上陣去了。
2CHR|18|30|亞蘭 王吩咐他的戰車長說：「你們不要與他們的大將或小兵交戰，只要單單攻擊 以色列 王。」
2CHR|18|31|那些戰車長看見 約沙法 就說：「這一定是 以色列 王！」他們轉過去與他交戰。 約沙法 一呼喊，耶和華就幫助他，上帝使他們轉離他。
2CHR|18|32|戰車長見他不是 以色列 王，就轉身不追他了。
2CHR|18|33|有一人開弓，並不知情，箭恰巧射入 以色列 王鎧甲的縫裏。王對駕車的說：「我受重傷了，你掉過車來，載我離開戰場！」
2CHR|18|34|那日，戰況越來越猛， 以色列 王勉強站在戰車上，面對 亞蘭 人，直到傍晚。日落的時候，王就死了。
2CHR|19|1|猶大 王 約沙法 平安回 耶路撒冷 ，到自己的宮裏。
2CHR|19|2|哈拿尼 的兒子 耶戶 先見出來迎接 約沙法 王，對他說：「你怎麼可以幫助惡人，愛那恨耶和華的人呢？因此耶和華的憤怒臨到你了。
2CHR|19|3|然而你還有善行，因你從國中除掉 亞舍拉 ，立定心意尋求上帝。」
2CHR|19|4|約沙法 住在 耶路撒冷 ，以後又出巡民間，從 別是巴 直到 以法蓮 山區，引導百姓歸向耶和華－他們列祖的上帝。
2CHR|19|5|他在國中，在 猶大 一切堅固城設立審判官，各城都是如此。
2CHR|19|6|他對審判官說：「你們應當謹慎所做的事，因為你們審判不是為人，而是為耶和華。在審判的事上，他必與你們同在。
2CHR|19|7|現在，你們應當敬畏耶和華，謹慎辦事，因為耶和華－我們的上帝沒有不義，不看人的情面，也不受賄賂。」
2CHR|19|8|約沙法 從 利未 人和祭司，以及 以色列 族長中，也委派人在 耶路撒冷 為耶和華施行審判，為 耶路撒冷 的居民聽訟斷案 。
2CHR|19|9|約沙法 吩咐他們說：「你們當這樣，以敬畏耶和華、誠實和純正的心辦事。
2CHR|19|10|你們住在各城的弟兄，若有爭訟的案件呈到你們這裏，或為流血，或犯律法、誡命、律例、典章，你們要警戒他們，免得他們得罪耶和華，以致憤怒臨到你們和你們的弟兄；你們當這樣行，就沒有罪了。
2CHR|19|11|看哪，凡屬耶和華的事，有 亞瑪利雅 祭司長管理你們；凡屬王的事，有 猶大 家的領袖 以實瑪利 的兒子 西巴第雅 管理你們；在你們面前有 利未 人作官長。你們應當壯膽辦事，願耶和華與善人同在。」
2CHR|20|1|此後， 摩押 人和 亞捫 人，連同一些 米烏尼 人 來攻擊 約沙法 。
2CHR|20|2|有人來報告 約沙法 說：「從海的那邊， 以東 有大軍來攻擊你，看哪，他們在 哈洗遜‧他瑪 ，就是 隱‧基底 。」
2CHR|20|3|約沙法 懼怕，就定意尋求耶和華，在全 猶大 宣告禁食。
2CHR|20|4|於是 猶大 人聚集，求耶和華幫助，甚至他們從 猶大 各城前來尋求耶和華。
2CHR|20|5|約沙法 站在 猶大 和 耶路撒冷 的會眾中，在耶和華殿新的院子前，
2CHR|20|6|說：「耶和華－我們列祖的上帝啊，你不是天上的上帝嗎？你不是萬邦萬國的主宰嗎？在你手中有大能大力，無人能抵擋你。
2CHR|20|7|我們的上帝啊，你不是曾在你百姓 以色列 面前驅逐這地的居民，將這地賜給你朋友 亞伯拉罕 的後裔永遠為業嗎？
2CHR|20|8|他們住在這地，又為你的名建造聖所，說：
2CHR|20|9|『若有禍患臨到我們，或刀兵的懲罰，或瘟疫饑荒，我們在急難的時候，站在這殿前向你呼求，你必垂聽並且拯救，因為你的名在這殿裏。』
2CHR|20|10|現在，看哪， 以色列 人出 埃及 地的時候，你不容許 以色列 人侵犯 亞捫 人、 摩押 人和 西珥山 人， 以色列 人就離開他們，不滅絕他們。
2CHR|20|11|看哪，他們這樣回報我們，要來驅逐我們離開你賜給我們為業之地。
2CHR|20|12|我們的上帝啊，你不懲罰他們嗎？因為我們無力抵擋這來攻擊我們的大軍。我們不知道該怎麼做，我們的眼目單仰望你。」
2CHR|20|13|猶大 眾人和他們的孩童、妻子、兒女都站在耶和華面前。
2CHR|20|14|那時，耶和華的靈在會眾中臨到 利未 人 亞薩 的後裔 雅哈悉 ，他是 瑪探雅 的玄孫， 耶利 的曾孫， 比拿雅 的孫子， 撒迦利雅 的兒子。
2CHR|20|15|他說：「 猶大 眾人、 耶路撒冷 的居民和 約沙法 王啊，你們要留心聽，耶和華對你們如此說：『不要因這大軍恐懼驚惶，因為勝敗不在乎你們，而是在乎上帝。
2CHR|20|16|明日你們要下去迎敵；看哪，他們從 洗斯坡 上來，你們必在 耶魯伊勒 曠野前的谷口遇見他們。
2CHR|20|17|猶大 和 耶路撒冷 人哪，這次你們不要爭戰，要擺陣站著，看耶和華為你們施行拯救。不要恐懼，也不要驚惶。明日當出去迎敵，因為耶和華與你們同在。』」
2CHR|20|18|約沙法 屈身，臉伏於地， 猶大 眾人和 耶路撒冷 的居民也俯伏在耶和華面前，敬拜耶和華。
2CHR|20|19|哥轄 子孫和 可拉 子孫的 利未 人都起來，用極大的聲音讚美耶和華－ 以色列 的上帝。
2CHR|20|20|清晨，眾人早起往 提哥亞 的曠野去。出去的時候， 約沙法 站著說：「 猶大 人和 耶路撒冷 的居民哪，要聽我說：信靠耶和華－你們的上帝就必站立得穩；信賴他的先知就必亨通。」
2CHR|20|21|約沙法 與百姓商議，就設立歌唱的人，頌讚耶和華，使他們穿上聖潔的禮服，走在軍隊前讚美耶和華： 「當稱謝耶和華， 因他的慈愛永遠長存！」
2CHR|20|22|他們開始唱歌讚美的時候，耶和華派伏兵擊殺那來攻擊 猶大 的 亞捫 人、 摩押 人和 西珥山 人，他們就被打敗了。
2CHR|20|23|亞捫 人和 摩押 人起來，擊殺住 西珥山 的人，把他們滅盡；滅盡住 西珥山 的人之後，他們又彼此自相擊殺。
2CHR|20|24|猶大 人來到曠野的瞭望樓，向那大軍觀看，看哪，遍地都是屍體，沒有一個逃脫的。
2CHR|20|25|約沙法 和他的百姓就來收取掠物，找到許多牲畜 、財物、衣服 和珍寶。他們取掠物歸為己有，直到無法攜帶；因為掠物太多，他們足足收取了三日。
2CHR|20|26|第四日，眾人聚集在 比拉迦谷 ，在那裏稱頌耶和華；因此那地方名叫 比拉迦谷 ，直到今日。
2CHR|20|27|在 約沙法 率領下， 猶大 人和 耶路撒冷 人都歡歡喜喜地回 耶路撒冷 ，耶和華使他們因戰勝仇敵而喜樂。
2CHR|20|28|他們彈琴、鼓瑟、吹號來到 耶路撒冷 ，進了耶和華的殿。
2CHR|20|29|地上所有的邦國聽見耶和華打敗 以色列 的仇敵，就都懼怕上帝。
2CHR|20|30|這樣， 約沙法 的國得享太平，因為上帝賜他四境平安。
2CHR|20|31|約沙法 作 猶大 王，登基的時候年三十五歲，在 耶路撒冷 作王二十五年。他母親名叫 阿蘇巴 ，是 示利希 的女兒。
2CHR|20|32|約沙法 效法他父親 亞撒 所行的道，不偏離左右，行耶和華眼中看為正的事。
2CHR|20|33|只是丘壇還沒有廢去，百姓也沒有立定心意歸向他們列祖的上帝。
2CHR|20|34|約沙法 其餘的事，看哪，自始至終都寫在 哈拿尼 的兒子 耶戶 的書上，這些事也記載在《以色列諸王記》上。
2CHR|20|35|此後， 猶大 王 約沙法 與 以色列 王 亞哈謝 結盟； 亞哈謝 多行惡事。
2CHR|20|36|他們合夥造船要往 他施 去，就在 以旬‧迦別 造船。
2CHR|20|37|瑪利沙 人 多大瓦 的兒子 以利以謝 向 約沙法 預言說：「因你與 亞哈謝 結盟，耶和華必破壞你所造的。」後來那些船果然毀壞，不能往 他施 去了。
2CHR|21|1|約沙法 與他祖先同睡，與他祖先同葬在 大衛城 ，他的兒子 約蘭 接續他作王。
2CHR|21|2|約蘭 有幾個兄弟，就是 約沙法 的兒子 亞撒利雅 、 耶歇 、 撒迦利雅 、 亞撒列夫 、 米迦勒 、 示法提雅 ；這些都是 以色列 王 約沙法 的兒子。
2CHR|21|3|他們的父親把許多禮物，金銀財寶和 猶大 的堅固城賜給他們，卻把國賜給 約蘭 ，因為他是長子。
2CHR|21|4|約蘭 起來治理他父親的國，奮勇自強，用刀殺了他所有的兄弟和 以色列 的幾個領袖。
2CHR|21|5|約蘭 登基的時候年三十二歲，在 耶路撒冷 作王八年。
2CHR|21|6|他行 以色列 諸王的道，正如 亞哈 家所行的，因他娶了 亞哈 的女兒為妻，行耶和華眼中看為惡的事。
2CHR|21|7|耶和華卻因自己與 大衛 所立的約，不肯滅絕 大衛 的家，要照他所應許的，永遠賜燈光給 大衛 和他的子孫。
2CHR|21|8|約蘭 在位期間， 以東 背叛，自己立王治理他們，脫離 猶大 的權勢。
2CHR|21|9|約蘭 就率領他的軍官和所有的戰車過去。他夜間起來，攻打圍困他的 以東 人和戰車長。
2CHR|21|10|這樣， 以東 背叛，脫離 猶大 的權勢，直到今日。那時， 立拿 也背叛了，脫離它的權勢，因為 約蘭 離棄耶和華－他列祖的上帝。
2CHR|21|11|他又在 猶大 山嶺 建造丘壇，使 耶路撒冷 的居民行淫，誘惑 猶大 。
2CHR|21|12|以利亞 先知寫信給 約蘭 說：「耶和華－你祖先 大衛 的上帝如此說：『因為你不行你父 約沙法 和 猶大 王 亞撒 的道，
2CHR|21|13|反而行 以色列 諸王的道，使 猶大 和 耶路撒冷 居民行淫，像 亞哈 家行淫一樣，又殺了你父家比你好的那些兄弟。
2CHR|21|14|看哪，耶和華必降大災於你的百姓和你的妻妾、兒女，以及你一切所有的。
2CHR|21|15|至於你，你必患許多的病 ，你的腸子也必生許多的病，日漸沉重，直到腸子墜落下來。』」
2CHR|21|16|耶和華激發 非利士 人和靠近 古實 人的 阿拉伯 人的心來攻擊 約蘭 。
2CHR|21|17|他們上來攻擊 猶大 ，侵入境內，擄掠了王宮裏所有的財物和他的妻妾、兒女，除了他的小兒子 約哈斯 之外，沒有留下一個兒子。
2CHR|21|18|這一切事以後，耶和華擊打 約蘭 ，使他的腸子患不能醫治的病。
2CHR|21|19|這病纏綿日久，過了二年，腸子墜落下來，他就病重而死。他的百姓沒有為他生火誌哀，像從前為他祖先生火一樣。
2CHR|21|20|約蘭 登基的時候年三十二歲，在 耶路撒冷 作王八年。他逝世無人思慕，眾人把他葬在 大衛城 ，只是不在列王的墳墓裏。
2CHR|22|1|耶路撒冷 的居民立 約蘭 的小兒子 亞哈謝 接續他作王，因為跟隨 阿拉伯 人來攻營的軍兵把 亞哈謝 所有的兄長都殺了； 猶大 王 約蘭 的兒子 亞哈謝 就作了王。
2CHR|22|2|亞哈謝 登基的時候年四十二歲 ，在 耶路撒冷 作王一年。他母親名叫 亞她利雅 ，是 暗利 的孫女。
2CHR|22|3|亞哈謝 也行 亞哈 家的道，因為他母親給他主謀，使他行惡。
2CHR|22|4|他行耶和華眼中看為惡的事，像 亞哈 家一樣；因他父親死後，他們給他主謀，使他敗壞。
2CHR|22|5|他也聽從他們的計謀，與 以色列 王 亞哈 的兒子 約蘭 同往 基列 的 拉末 去，與 亞蘭 王 哈薛 交戰。 亞蘭 人打傷了 約蘭 ，
2CHR|22|6|他回到 耶斯列 ，醫治在 拉末 與 亞蘭 王 哈薛 打仗時被擊打所受的傷。 約蘭 的兒子 猶大 王 亞哈謝 因為 亞哈 的兒子 約蘭 病了，就下到 耶斯列 看望他。
2CHR|22|7|亞哈謝 去見 約蘭 而遇害，這是出乎上帝；因為他一到就同 約蘭 出去攻擊 寧示 的孫子 耶戶 ；這 耶戶 是耶和華所膏，使他剪除 亞哈 家的。
2CHR|22|8|耶戶 向 亞哈 家施行懲罰的時候，遇見 猶大 的眾領袖和 亞哈謝 的姪子們正服事 亞哈謝 ，就把他們都殺了。
2CHR|22|9|亞哈謝 躲在 撒瑪利亞 ， 耶戶 尋找他，眾人把他拿住，送到 耶戶 那裏，就殺了他。他們把他埋葬，因他們說，他是那盡心尋求耶和華之 約沙法 的兒子。這樣， 亞哈謝 的家無力保住國權。
2CHR|22|10|亞哈謝 的母親 亞她利雅 見她兒子死了，就起來剿滅 猶大 王室所有的後裔。
2CHR|22|11|但王的女兒 約示巴 將 亞哈謝 的兒子 約阿施 從那被殺的王子中偷出來，把他和他的奶媽藏在臥房裏。 約示巴 是 約蘭 王的女兒， 亞哈謝 的妹妹，祭司 耶何耶大 的妻子。她藏了 約阿施 ，躲避 亞她利雅 ，免受殺害。
2CHR|22|12|亞她利雅 治理這地的時候， 約阿施 和他們一同在上帝殿裏藏了六年。
2CHR|23|1|第七年， 耶何耶大 奮勇自強，叫了 耶羅罕 的兒子 亞撒利雅 、 約哈難 的兒子 以實瑪利 、 俄備得 的兒子 亞撒利雅 、 亞大雅 的兒子 瑪西雅 ，和 細基利 的兒子 以利沙法 等眾百夫長，與他們立約。
2CHR|23|2|他們走遍 猶大 ，從 猶大 各城召集 利未 人和 以色列 的眾族長到 耶路撒冷 來。
2CHR|23|3|全會眾在上帝殿裏與王立約。 耶何耶大 對他們說：「看哪，王的兒子必作王，正如耶和華指著 大衛 子孫所應許的。
2CHR|23|4|你們要這樣做：在安息日值班的祭司和 利未 人，三分之一要把守各門，
2CHR|23|5|三分之一要在王宮，三分之一要在 根基門 ；眾百姓都要在耶和華殿的院內。
2CHR|23|6|除了祭司和供職的 利未 人之外，不准別人進耶和華的殿；只有他們可以進去，因為他們是神聖的。眾百姓都要遵守耶和華所吩咐的。
2CHR|23|7|利未 人要手中各拿兵器，四圍保護王；凡擅自進殿的，要被處死。王出入的時候，你們當跟隨他。」
2CHR|23|8|利未 人和 猶大 眾人都照著 耶何耶大 祭司一切所吩咐的去做，各帶自己的人，無論安息日值班或不值班的都來，因為 耶何耶大 祭司不許他們下班。
2CHR|23|9|耶何耶大 祭司就把上帝殿裏所藏 大衛 王的槍和大小盾牌交給百夫長，
2CHR|23|10|又分派眾百姓手中各拿兵器，在祭壇和殿那裏，從殿南到殿北，站在王的四圍；
2CHR|23|11|他們領 約阿施 出來，給他戴上冠冕，把律法書交給他，立他作王。 耶何耶大 和他的兒子們膏他，他們說：「願王萬歲！」
2CHR|23|12|亞她利雅 聽見百姓奔走讚美王的聲音，就進耶和華的殿，到百姓那裏。
2CHR|23|13|她觀看，看哪，王站在殿門的柱旁，百夫長和號手在王旁邊，國中的眾百姓都歡樂吹號，又有歌唱的人用樂器領人歌唱讚美。 亞她利雅 就撕裂衣服，喊著說：「反了！反了！」
2CHR|23|14|耶何耶大 祭司帶領管軍兵的百夫長出來，對他們說：「把她從行列之間趕出去，凡跟隨她的必用刀殺死！」因為祭司說：「不可在耶和華殿裏殺她。」
2CHR|23|15|他們就下手拿住她；她進入通往王宮的 馬門 ，他們就在那裏把她殺了。
2CHR|23|16|耶何耶大 與眾百姓，又與王立約，要作耶和華的子民。
2CHR|23|17|於是眾百姓到 巴力 廟去，拆毀了廟，打碎祭壇和偶像，又在壇前把 巴力 的祭司 瑪坦 殺了。
2CHR|23|18|耶何耶大 派官員在 利未 家的祭司手下看守耶和華的殿，他們是 大衛 所分派的，在耶和華殿中照 摩西 律法上所寫，獻燔祭給耶和華，又按 大衛 所定的，歡樂歌唱。
2CHR|23|19|耶何耶大 又設立守衛把守耶和華殿的各門，無論因何事而不潔淨的人，都不准進去。
2CHR|23|20|他又率領百夫長和貴族，與民間的官長，以及國中的眾百姓，請王從耶和華的殿下來，由 上門 正中進入王宮，使王坐在國度的王位上。
2CHR|23|21|國中的眾百姓都歡樂，合城也都平靜。他們已將 亞她利雅 用刀殺了。
2CHR|24|1|約阿施 登基的時候年方七歲，在 耶路撒冷 作王四十年。他母親名叫 西比亞 ，是 別是巴 人。
2CHR|24|2|耶何耶大 祭司在世的日子， 約阿施 行耶和華眼中看為正的事。
2CHR|24|3|耶何耶大 為他娶了兩個妻子，他生兒育女。
2CHR|24|4|此後， 約阿施 有心重修耶和華的殿，
2CHR|24|5|就召集祭司和 利未 人，吩咐他們說：「你們要往 猶大 各城去，向 以色列 眾人徵收銀子，按每年的需要整修你們上帝的殿；你們要急速辦理這事。」但 利未 人沒有急速辦理。
2CHR|24|6|王召了 耶何耶大 祭司長來，對他說：「從前耶和華的僕人 摩西 ，為法櫃的帳幕與 以色列 會眾所定的捐獻，你為何不叫 利未 人照這例向 猶大 和 耶路撒冷 徵收呢？」
2CHR|24|7|因為那惡婦 亞她利雅 的兒子們曾拆毀上帝的殿，又用耶和華殿中分別為聖的物供奉諸 巴力 。
2CHR|24|8|於是王下令造一個櫃子，放在耶和華殿的門外，
2CHR|24|9|又通告 猶大 和 耶路撒冷 ，要將上帝僕人 摩西 在曠野所吩咐 以色列 的捐獻送來給耶和華。
2CHR|24|10|眾領袖和百姓都歡歡喜喜帶捐獻來，投入櫃中，直到投滿。
2CHR|24|11|利未 人見銀子多了，把櫃子抬到王所派的官長面前；這時王的書記和祭司長的助手就會來把櫃子倒空，然後放回原處。日日都是這樣做，積蓄的銀子很多。
2CHR|24|12|王與 耶何耶大 把銀子交給耶和華殿裏辦事的人，他們就雇了石匠、木匠重修耶和華的殿，又雇了鐵匠、銅匠整修耶和華的殿。
2CHR|24|13|工人做工，修理工程在他們手中漸漸完成，他們將上帝的殿修理得如同從前一樣，非常堅固。
2CHR|24|14|他們做完了，就把多餘的銀子拿到王與 耶何耶大 面前，用以製造耶和華殿供奉所用的器皿和調羹，以及金銀的器皿。 耶何耶大 在世的日子，眾人經常在耶和華殿裏獻燔祭。
2CHR|24|15|耶何耶大 年紀老邁，日子滿足而死，死的時候年一百三十歲。
2CHR|24|16|眾人把他與列王同葬在 大衛城 ，因為他在 以色列 中為上帝和他的殿做了美善的事。
2CHR|24|17|耶何耶大 死後， 猶大 的眾領袖來叩拜王，那時王就聽了他們。
2CHR|24|18|他們離棄耶和華－他們列祖上帝的殿，去事奉 亞舍拉 和偶像；因他們這罪，就有憤怒臨到 猶大 和 耶路撒冷 。
2CHR|24|19|但上帝仍差遣先知到他們那裏，引導他們歸向耶和華。先知警戒他們，他們卻不肯聽。
2CHR|24|20|那時，上帝的靈感動 耶何耶大 的兒子 撒迦利亞 祭司，他就站在上面，對百姓說：「上帝如此說：『你們為何干犯耶和華的誡命，以致不得亨通呢？因為你們離棄耶和華，所以他也離棄你們。』」
2CHR|24|21|眾人謀害 撒迦利亞 ，照著王的吩咐，在耶和華殿的院內用石頭打死他。
2CHR|24|22|這樣， 約阿施 王不記念 撒迦利亞 的父親 耶何耶大 向自己所施的恩，殺了他的兒子。 撒迦利亞 臨死的時候說：「願耶和華鑒察伸冤！」
2CHR|24|23|年底的時候， 亞蘭 的軍兵上來攻擊 約阿施 ，來到 猶大 和 耶路撒冷 ，殺了百姓中的眾領袖，把所掠取的財物全送到 大馬士革 王那裏。
2CHR|24|24|亞蘭 的軍兵雖只來了一小隊人，耶和華卻將極大的軍隊交在他們手裏；因為 猶大 人離棄耶和華－他們列祖的上帝，所以 亞蘭 人懲罰 約阿施 。
2CHR|24|25|亞蘭 人離開 約阿施 的時候，他患重病 ；他的臣僕背叛他，要報 耶何耶大 祭司兒子 的流血之仇，在床上殺了他。他就死了，葬在 大衛城 ，只是不葬在列王的墳墓裏。
2CHR|24|26|背叛他的是 亞捫 婦人 示米押 的兒子 撒拔 和 摩押 婦人 示米利 的兒子 約薩拔 。
2CHR|24|27|至於他的兒子們和他所受的眾多警戒，以及他重修上帝殿的事，看哪，都寫在《列王評傳》上。他的兒子 亞瑪謝 接續他作王。
2CHR|25|1|亞瑪謝 登基的時候年二十五歲，在 耶路撒冷 作王二十九年。他母親名叫 約耶但 ，是 耶路撒冷 人。
2CHR|25|2|亞瑪謝 行耶和華眼中看為正的事，只是沒有純正的心。
2CHR|25|3|他的王國一鞏固，就把殺他父王的臣僕殺了，
2CHR|25|4|卻沒有處死他們的兒子，這是照 摩西 律法書上耶和華所吩咐的說：「不可因子殺父，也不可因父殺子，各人要為自己的罪而死。」
2CHR|25|5|亞瑪謝 召集 猶大 人，按著父家為全 猶大 和 便雅憫 設立千夫長、百夫長，又數點人數，從二十歲以上，能拿槍拿盾牌出去打仗的精兵共有三十萬；
2CHR|25|6|又用一百他連得銀子，從 以色列 招募了十萬大能的勇士。
2CHR|25|7|有一個神人來見 亞瑪謝 ，對他說：「王啊，不要帶領 以色列 的軍兵與你同去，因為耶和華不和 以色列 ，和任何 以法蓮 的子孫同在。
2CHR|25|8|你若一定要去，就奮勇作戰吧！但上帝必使你敗在敵人面前，因為上帝能助人得勝，也能使人落敗。」
2CHR|25|9|亞瑪謝 問神人：「我給了 以色列 軍隊的那一百他連得銀子怎麼樣呢？」神人回答：「耶和華會把比這些更多的賜給你。」
2CHR|25|10|於是 亞瑪謝 把那從 以法蓮 來的軍兵分別出來，叫他們到自己的地方去。他們非常惱怒 猶大 ，氣憤地回自己的地方去了。
2CHR|25|11|亞瑪謝 壯起膽來，率領他的軍隊到 鹽谷 ，殺了一萬 西珥 人。
2CHR|25|12|猶大 人又生擒了一萬人，把他們帶到 西拉 山頂上，從 西拉 山頂扔下去，把他們全都摔碎了。
2CHR|25|13|但 亞瑪謝 所打發回去、不許一同出征的那些軍兵劫掠 猶大 各城，從 撒瑪利亞 直到 伯‧和崙 ，殺了三千人，搶了許多財物。
2CHR|25|14|亞瑪謝 擊殺 以東 人回來以後，他把 西珥 人的神像帶回，立為自己的神明，在它們面前叩拜燒香。
2CHR|25|15|耶和華的怒氣向 亞瑪謝 發作，差派一個先知去見他，對他說：「這些神明不能救自己的百姓脫離你的手，你為何尋求它們呢？」
2CHR|25|16|先知與王說話的時候，王對他說：「難道我們立你作王的謀士嗎？你住口吧！為何要挨打呢？」先知就止住了，卻說：「我知道上帝已定意要消滅你，因為你行這事，不聽從我的勸戒。」
2CHR|25|17|猶大 王 亞瑪謝 經商議後，就派人去見 耶戶 的孫子， 約哈斯 的兒子 以色列 王 約阿施 ，說：「來，讓我們面對面較量吧！」
2CHR|25|18|以色列 王 約阿施 派人去見 猶大 王 亞瑪謝 ，說：「 黎巴嫩 的蒺藜派人去見 黎巴嫩 的香柏樹，說：『將你的女兒嫁給我的兒子。』但有一隻野獸經過 黎巴嫩 ，把蒺藜踐踏了。
2CHR|25|19|你說，看哪，你打敗了 以東 ，就心高氣傲，以此為榮。現在，你待在家裏算了吧，為何要惹禍使自己和 猶大 一同敗亡呢？」
2CHR|25|20|亞瑪謝 卻不肯聽從。這是出乎上帝，好將他們交在敵人手裏，因為他們尋求 以東 的神明。
2CHR|25|21|於是 以色列 王 約阿施 上來，在 猶大 的 伯‧示麥 與 猶大 王 亞瑪謝 面對面較量。
2CHR|25|22|猶大 敗在 以色列 面前，他們逃跑，各人逃回自己的帳棚去了。
2CHR|25|23|以色列 王 約阿施 在 伯‧示麥 擒住 約哈斯 的孫子， 約阿施 的兒子 猶大 王 亞瑪謝 ，把他帶到 耶路撒冷 ，又拆毀 耶路撒冷 的城牆，從 以法蓮門 直到 角門 共四百肘。
2CHR|25|24|他帶著 俄別‧以東 所看守上帝殿裏的一切金銀和器皿，與王宮裏的財寶，又帶著人質，回 撒瑪利亞 去了。
2CHR|25|25|約哈斯 的兒子 以色列 王 約阿施 死後， 猶大 王 約阿施 的兒子 亞瑪謝 又活了十五年。
2CHR|25|26|亞瑪謝 其餘的事，自始至終，看哪，不都寫在《猶大和以色列諸王記》上嗎？
2CHR|25|27|自從 亞瑪謝 離棄耶和華之後，在 耶路撒冷 有人背叛他，他就逃往 拉吉 ；他們卻派人追到 拉吉 ，在那裏殺了他。
2CHR|25|28|有人用馬將他馱回，把他與祖先一同葬在 猶大 的城 。
2CHR|26|1|猶大 眾百姓立 烏西雅 接續他父親 亞瑪謝 作王，那時他年十六歲。
2CHR|26|2|亞瑪謝 王與他祖先同睡之後， 烏西雅 收復 以祿 回歸 猶大 ，又重新修建。
2CHR|26|3|烏西雅 登基的時候年十六歲，在 耶路撒冷 作王五十二年。他母親名叫 耶可利雅 ，是 耶路撒冷 人。
2CHR|26|4|烏西雅 行耶和華眼中看為正的事，效法他父親 亞瑪謝 一切所行的。
2CHR|26|5|撒迦利亞 是一個通曉上帝默示的人 ，他在世的日子， 烏西雅 定意尋求上帝； 烏西雅 尋求耶和華的日子，上帝使他亨通。
2CHR|26|6|他出去攻擊 非利士 人，拆毀了 迦特 、 雅比尼 和 亞實突 的城牆，又在 非利士 人中，在 亞實突 境內建築城鎮。
2CHR|26|7|上帝幫助他攻擊 非利士 人和住在 姑珥‧巴力 的 阿拉伯 人，以及 米烏尼 人。
2CHR|26|8|米烏尼 人 向 烏西雅 進貢。他的名聲傳到 埃及 ，因他非常強盛。
2CHR|26|9|烏西雅 在 耶路撒冷 的 角門 和 谷門 ，以及城牆轉角之處建築城樓，非常堅固。
2CHR|26|10|他在曠野建築瞭望樓，又挖了許多井，因為他在 謝非拉 和平原有很多牲畜。他在山區和肥沃的土地雇用耕種田地和修整葡萄園的人，因為他喜愛土地。
2CHR|26|11|烏西雅 又有軍兵，照書記 耶利 和官長 瑪西雅 所數點的，在王的一個將軍 哈拿尼雅 手下，分隊出戰。
2CHR|26|12|族長和大能勇士的總數共二千六百人，
2CHR|26|13|他們手下的軍兵共三十萬七千五百人，都大有能力，善於作戰，幫助王攻擊仇敵。
2CHR|26|14|烏西雅 為全軍預備盾牌、頭盔、鎧甲、槍、弓和甩石的機弦，
2CHR|26|15|又在 耶路撒冷 叫巧匠設計機器，安在城樓和角樓上，用以射箭，投擲大石。 烏西雅 的名聲傳到遠方，因為他得了非凡的幫助，極其強盛。
2CHR|26|16|烏西雅 既強盛，就心高氣傲，以致敗壞。他干犯耶和華－他的上帝，進耶和華的殿，要在香壇上燒香。
2CHR|26|17|亞撒利雅 祭司率領八十名勇敢的耶和華的祭司，跟隨他進去。
2CHR|26|18|他們阻止 烏西雅 王，對他說：「 烏西雅 啊，給耶和華燒香不是你的事，而是 亞倫 子孫的事，他們是分別為聖來燒香的祭司。你出聖殿吧！因為你犯了罪，耶和華上帝必不使你得尊榮。」
2CHR|26|19|烏西雅 發怒，手拿香爐要燒香。他在耶和華殿中香壇旁向眾祭司發怒的時候，他的額頭在眾祭司面前忽然長出痲瘋 。
2CHR|26|20|亞撒利雅 祭司長和眾祭司轉向他，看哪，他的額頭長出痲瘋，就催他離開那裏；他自己也急速出去，因為耶和華降災於他。
2CHR|26|21|烏西雅 王患痲瘋直到死的那日；他因為染上痲瘋，就住在隔離的行宮裏，與耶和華的殿隔絕。他兒子 約坦 管理王的家，治理這地的百姓。
2CHR|26|22|烏西雅 其餘的事，自始至終， 亞摩斯 的兒子 以賽亞 先知都記錄下來。
2CHR|26|23|烏西雅 與他祖先同睡，與他祖先同葬在田間的王陵；因為人說，他是長痲瘋的。他的兒子 約坦 接續他作王。
2CHR|27|1|約坦 登基的時候年二十五歲，在 耶路撒冷 作王十六年。他母親名叫 耶路沙 ，是 撒督 的女兒。
2CHR|27|2|約坦 行耶和華眼中看為正的事，效法他父親 烏西雅 一切所行的，只是他不入耶和華的殿。百姓仍舊行敗壞的事。
2CHR|27|3|約坦 建造耶和華殿的 上門 ，在 俄斐勒 城牆上有很多建設，
2CHR|27|4|又在 猶大 山區建造城鎮，在樹林中建築營寨和瞭望樓。
2CHR|27|5|約坦 與 亞捫 人的王打仗，勝了他們。那年 亞捫 人向他進貢一百他連得銀子，一萬歌珥小麥，一萬歌珥大麥；第二年、第三年 亞捫 人也這樣做。
2CHR|27|6|約坦 日漸強盛，因為他在耶和華－他上帝面前行正道。
2CHR|27|7|約坦 其餘的事和一切戰役，以及他的行為，看哪，都寫在《以色列和猶大列王記》上。
2CHR|27|8|他登基的時候年二十五歲，在 耶路撒冷 作王十六年。
2CHR|27|9|約坦 與他祖先同睡，葬在 大衛城 ，他兒子 亞哈斯 接續他作王。
2CHR|28|1|亞哈斯 登基的時候年二十歲，在 耶路撒冷 作王十六年。他不像他祖先 大衛 行耶和華眼中看為正的事，
2CHR|28|2|卻行 以色列 諸王的道，又鑄造諸 巴力 的像，
2CHR|28|3|照著耶和華從 以色列 人面前趕出的外邦人所行可憎的事，在 欣嫩子谷 燒香，用火焚燒他的兒女，
2CHR|28|4|又在丘壇上、山岡上、各青翠樹下獻祭燒香。
2CHR|28|5|耶和華－他的上帝將他交在 亞蘭 王手裏。 亞蘭 王打敗他，從他擄走了許多人，帶到 大馬士革 去。上帝又將他交在 以色列 王手裏， 以色列 王向他大行殺戮。
2CHR|28|6|利瑪利 的兒子 比加 一日之內在 猶大 殺了十二萬人，都是勇士，因為他們離棄了耶和華－他們列祖的上帝。
2CHR|28|7|有一個叫 細基利 的 以法蓮 勇士，殺了 瑪西雅 王子、 押斯利甘 宮廷總管和 以利加拿 宰相。
2CHR|28|8|以色列 人擄了他們的弟兄，連婦人帶兒女共二十萬，又掠取了許多財物，把這些掠物帶到 撒瑪利亞 去。
2CHR|28|9|但那裏有耶和華的一個先知，名叫 俄德 ，出來迎接往 撒瑪利亞 去的軍兵，對他們說：「看哪，耶和華－你們列祖的上帝惱怒 猶大 人，將他們交在你們手裏，你們竟怒氣沖天，向他們大行殺戮。
2CHR|28|10|如今你們又有意強逼 猶大 人和 耶路撒冷 人作你們的奴婢，你們豈不是也得罪了耶和華－你們的上帝嗎？
2CHR|28|11|現在你們當聽我說，要將從你們弟兄中擄來的釋放回去，因耶和華的烈怒已臨到你們了。」
2CHR|28|12|於是， 以法蓮 人的幾個領袖，就是 約哈難 的兒子 亞撒利雅 、 米實利末 的兒子 比利家 、 沙龍 的兒子 耶希西家 、 哈得萊 的兒子 亞瑪撒 ，起來攔阻從戰場上回來的人，
2CHR|28|13|對他們說：「你們不可把這些被擄的人帶到這裏，因我們已經得罪耶和華了。你們還想加增我們的罪惡過犯嗎？因為我們的罪過深重，已經有烈怒臨到 以色列 了。」
2CHR|28|14|於是帶兵器的人將擄來的人口和掠取的財物都留在眾領袖和全會眾面前。
2CHR|28|15|以上提名的那些人就起來，照顧被擄的人；其中凡赤身的，就從所掠取的財物中拿出衣服和鞋來，給他們穿，又給他們吃喝，用膏抹他們；其中凡軟弱的，就使他們騎驢，送到棕樹城 耶利哥 他們弟兄那裏。然後，他們就回 撒瑪利亞 去了。
2CHR|28|16|那時， 亞哈斯 王派人去求 亞述 諸王 來幫助他，
2CHR|28|17|因為 以東 人又來攻擊 猶大 ，擄掠俘虜。
2CHR|28|18|非利士 人也來侵佔 謝非拉 和 猶大 的 尼革夫 的城鎮，攻取了 伯‧示麥 、 亞雅崙 、 基低羅 、 梭哥 和所屬的鄉鎮、 亭拿 和所屬的鄉鎮、 瑾鎖 和所屬的鄉鎮，就住在那裏。
2CHR|28|19|因為 以色列 王 亞哈斯 在 猶大 放肆，大大干犯耶和華，所以耶和華使 猶大 卑微。
2CHR|28|20|亞述 王 提革拉‧毗列色 來攻擊他，不幫助他，反倒欺負他。
2CHR|28|21|亞哈斯 從耶和華殿裏和王宮中，以及眾領袖家中取財寶送給 亞述 王，也無濟於事。
2CHR|28|22|這 亞哈斯 王在急難的時候，越發得罪耶和華。
2CHR|28|23|他向那攻擊他的 大馬士革 的神明獻祭，說：「因為 亞蘭 王的神明幫助他們，我也要向這些神明獻祭，好讓它們幫助我。」但那些神明卻使他和全 以色列 敗亡。
2CHR|28|24|亞哈斯 聚集上帝殿裏的器皿，把上帝殿裏的器皿都打碎了，並且封鎖耶和華殿的門，又在 耶路撒冷 各處的轉角為自己建築祭壇。
2CHR|28|25|他在 猶大 各城建立丘壇，向別神燒香，惹耶和華－他列祖的上帝發怒。
2CHR|28|26|亞哈斯 其餘的事和他一切的行為，自始至終，看哪，都寫在《猶大和以色列諸王記》上。
2CHR|28|27|亞哈斯 與他祖先同睡，葬在 耶路撒冷 城裏，卻沒有送入 以色列 諸王的墳墓。他的兒子 希西家 接續他作王。
2CHR|29|1|希西家 登基的時候年二十五歲，在 耶路撒冷 作王二十九年。他母親名叫 亞比雅 ，是 撒迦利雅 的女兒。
2CHR|29|2|希西家 行耶和華眼中看為正的事，效法他祖先 大衛 一切所行的。
2CHR|29|3|元年正月，他開了耶和華殿的門，重新整修。
2CHR|29|4|他召祭司和 利未 人來，聚集在東邊的廣場，
2CHR|29|5|對他們說：「 利未 人哪，當聽我說：現在你們要將自己分別為聖，又將耶和華－你們列祖上帝的殿分別為聖，從聖所中除去污穢之物。
2CHR|29|6|因我們的祖先犯了罪，行耶和華－我們上帝眼中看為惡的事，離棄他，轉臉背向耶和華的居所。
2CHR|29|7|他們又封鎖走廊的門，吹滅燈火，不在聖所中向 以色列 的上帝燒香，或獻燔祭。
2CHR|29|8|耶和華的憤怒臨到 猶大 和 耶路撒冷 ，使他們恐懼，令人驚駭，使人嗤笑，正如你們親眼所見的。
2CHR|29|9|看哪，我們的祖宗倒在刀下，我們的妻子兒女也為此被擄掠。
2CHR|29|10|現在我心中有意與耶和華－ 以色列 的上帝立約，好使他的烈怒轉離我們。
2CHR|29|11|我的眾子啊，現在不要懈怠；因為耶和華揀選你們站在他面前事奉他，作他的僕人，向他燒香。」
2CHR|29|12|於是， 利未 人起來，當中有 哥轄 的子孫， 亞瑪賽 的兒子 瑪哈 、 亞撒利雅 的兒子 約珥 ； 米拉利 的子孫， 亞伯底 的兒子 基士 、 耶哈利勒 的兒子 亞撒利雅 ； 革順 人， 薪瑪 的兒子 約亞 、 約亞 的兒子 伊甸 ；
2CHR|29|13|以利撒反 的子孫 申利 和 耶利 ； 亞薩 的子孫， 撒迦利雅 和 瑪探雅 ；
2CHR|29|14|希幔 的子孫 耶歇 和 示每 ； 耶杜頓 的子孫 示瑪雅 和 烏薛 。
2CHR|29|15|他們聚集他們的弟兄，將自己分別為聖，照著耶和華的話和王的吩咐，進去潔淨耶和華的殿。
2CHR|29|16|祭司進入耶和華的內殿要潔淨殿，把耶和華殿中所發現一切污穢之物都搬出去，搬到耶和華殿的院子，由 利未 人接走，搬出去到外頭的 汲淪溪 。
2CHR|29|17|從正月初一開始分別為聖，初八就來到耶和華殿的走廊。他們又用了八日使耶和華的殿分別為聖，到正月十六日才完成。
2CHR|29|18|於是，他們到裏面去見 希西家 王，說：「我們已將耶和華的全殿和燔祭壇，以及壇的一切器皿、供餅的供桌，與供桌的一切器皿都潔淨了；
2CHR|29|19|並且連 亞哈斯 王在位犯罪的時候所廢棄的器皿，我們也都預備齊全，分別為聖，看哪，它們都在耶和華的祭壇前。」
2CHR|29|20|希西家 王清早起來，召集城裏的領袖都上耶和華的殿。
2CHR|29|21|他們牽了七頭公牛，七隻公羊，七隻羔羊，七隻公山羊，要為國、為殿、為 猶大 作贖罪祭。王吩咐 亞倫 的子孫眾祭司在耶和華的壇上獻祭。
2CHR|29|22|他們宰了公牛，祭司將血接來，灑在壇上；他們宰了公羊，把血灑在壇上，又宰了羔羊，也把血灑在壇上。
2CHR|29|23|他們把那些作贖罪祭的公山羊牽到王和會眾面前，按手在公山羊上。
2CHR|29|24|祭司宰了羊，將血獻在壇上作贖罪祭，為全 以色列 贖罪，因為王吩咐要為全 以色列 獻上燔祭和贖罪祭。
2CHR|29|25|王又派 利未 人在耶和華殿中敲鈸，鼓瑟，彈琴，正如 大衛 和王的先見 迦得 ，以及 拿單 先知所吩咐的，就是耶和華藉先知所吩咐的。
2CHR|29|26|利未 人拿 大衛 的樂器，祭司拿號，一同站立。
2CHR|29|27|希西家 吩咐在壇上獻燔祭，開始獻燔祭的時候，他們就唱讚美耶和華的歌，吹號，並用 以色列 王 大衛 的樂器伴奏。
2CHR|29|28|全會眾都敬拜，歌唱的歌唱，吹號的吹號，如此直到燔祭獻完了。
2CHR|29|29|獻完了祭，王和所有在場跟隨他的人都俯伏敬拜。
2CHR|29|30|希西家 王與眾領袖吩咐 利未 人用 大衛 和 亞薩 先見的詩詞頌讚耶和華，他們歡歡喜喜地頌讚，低頭敬拜。
2CHR|29|31|希西家 回應說：「如今你們既承接聖職歸耶和華，就要前來把祭物和感謝祭奉到耶和華的殿裏。」會眾就奉上祭物和感謝祭，凡甘心樂意的也奉上燔祭。
2CHR|29|32|會眾所奉的燔祭數目如下：七十頭公牛，一百隻公羊，二百隻羔羊，這些全都是要作燔祭獻給耶和華的；
2CHR|29|33|又有分別為聖之物，就是六百頭公牛，三千隻綿羊。
2CHR|29|34|但祭司太少，不能剝盡所有燔祭牲的皮，所以他們的弟兄 利未 人幫助他們，直等獻祭的事完畢，直到其他的祭司也分別為聖了；因 利未 人以正直的心分別為聖，勝過祭司。
2CHR|29|35|燔祭和平安祭牲的脂肪，以及與燔祭同獻的澆酒祭很多。這樣，耶和華殿中的事務俱都齊備了。
2CHR|29|36|希西家 和眾百姓都因上帝為百姓所預備的而喜樂，因為這事辦得很迅速。
2CHR|30|1|希西家 派人去見 以色列 和 猶大 眾人，又寫信給 以法蓮 和 瑪拿西 人，要他們到 耶路撒冷 耶和華的殿，向耶和華－ 以色列 的上帝守逾越節，
2CHR|30|2|因為王和眾領袖，以及 耶路撒冷 全會眾已經商議，要在二月份守逾越節。
2CHR|30|3|那時他們不能守，因為分別為聖的祭司不夠，百姓也還沒有聚集在 耶路撒冷 。
2CHR|30|4|這事在王與全會眾眼中都看為合宜。
2CHR|30|5|於是他們下令，通告全 以色列 ，從 別是巴 直到 但 ，吩咐百姓都來，在 耶路撒冷 向耶和華－ 以色列 的上帝守逾越節，因為他們已經許久沒有照所寫的守這節了 。
2CHR|30|6|信差遵著王命，拿著王和眾領袖所發的信，送達全 以色列 和 猶大 ，說：「 以色列 人哪，當轉向耶和華－ 亞伯拉罕 、 以撒 、 以色列 的上帝，好叫他轉向你們這些脫離 亞述 諸王之手的餘民。
2CHR|30|7|不要效法你們的祖先和你們的弟兄；他們干犯耶和華－他們列祖的上帝，以致耶和華使他們令人驚駭，正如你們所見的。
2CHR|30|8|現在，不要像你們祖先硬著頸項，只要歸順耶和華，進入他的聖所，就是永遠成聖的居所，又要事奉耶和華－你們的上帝，好使他的烈怒轉離你們。
2CHR|30|9|你們若轉向耶和華，你們的弟兄和兒女必在擄掠他們的人面前蒙憐憫，得以歸回這地，因為耶和華－你們的上帝有恩惠，有憐憫。你們若轉向他，他必不會轉臉不顧你們。」
2CHR|30|10|信差從這城跑到那城，傳遍了 以法蓮 和 瑪拿西 之地，直到 西布倫 ；那裏的人卻戲笑他們，譏誚他們。
2CHR|30|11|然而 亞設 、 瑪拿西 、 西布倫 中也有人謙卑自己，來到 耶路撒冷 。
2CHR|30|12|上帝也按手在 猶大 人身上，使他們一心遵行王與眾領袖照著耶和華的話所發的命令。
2CHR|30|13|二月時，許多百姓聚集在 耶路撒冷 ，成為一個盛大的會，要守除酵節。
2CHR|30|14|他們起來，把 耶路撒冷 的祭壇和燒香的壇盡都除去，扔在 汲淪溪 中。
2CHR|30|15|二月十四日，他們宰了逾越節的羔羊。祭司與 利未 人覺得慚愧，就使自己分別為聖，把燔祭奉到耶和華的殿中。
2CHR|30|16|他們遵照神人 摩西 的律法，按定例站在自己的地方；祭司從 利未 人手裏接過血來，灑出去。
2CHR|30|17|會眾中有許多人尚未分別為聖，所以 利未 人為所有不潔的人宰逾越節的羔羊，使他們歸耶和華為聖。
2CHR|30|18|從 以法蓮 、 瑪拿西 、 以薩迦 、 西布倫 來的許多百姓尚未自潔，他們卻吃逾越節的羔羊，不合所寫的條例。 希西家 為他們禱告說：「求至善的耶和華饒恕
2CHR|30|19|那凡專心尋求上帝耶和華－他列祖的上帝，卻未照聖所潔淨禮自潔的人。」
2CHR|30|20|耶和華應允 希西家 ，醫治了百姓。
2CHR|30|21|在 耶路撒冷 的 以色列 人守除酵節七日，大大喜樂。 利未 人和祭司為耶和華演奏響亮的樂器，天天頌讚耶和華。
2CHR|30|22|希西家 慰勞所有精通禮儀，事奉耶和華的 利未 人。於是眾人吃節期的筵席七日，又獻平安祭，並且稱謝耶和華－他們列祖的上帝。
2CHR|30|23|全會眾商議，要再守節七日；於是他們歡歡喜喜地又守節七日。
2CHR|30|24|猶大 王 希西家 賜給會眾一千頭公牛，七千隻羊；眾領袖也賜給會眾一千頭公牛，一萬隻羊，並有許多祭司將自己分別為聖。
2CHR|30|25|猶大 全會眾、祭司、 利未 人和從 以色列 來的全會眾，以及那些從 以色列 地來的和住在 猶大 的寄居的人，盡都喜樂。
2CHR|30|26|這樣，在 耶路撒冷 大有喜樂，因自從 以色列 王 大衛 的兒子 所羅門 以來，在 耶路撒冷 從未有過這樣的喜樂。
2CHR|30|27|那時，祭司和 利未 人起來，為百姓祝福。他們的聲音蒙上帝垂聽，他們的禱告達到他天上的聖所。
2CHR|31|1|這一切事都完畢以後，在那裏的 以色列 眾人就到 猶大 的城鎮，打碎柱像，砍斷 亞舍拉 ，又在 猶大 、 便雅憫 、 以法蓮 、 瑪拿西 遍地把丘壇和祭壇完全拆毀。於是 以色列 眾人各回各城，各歸自己產業的地去了。
2CHR|31|2|希西家 分派祭司和 利未 人的班次，使祭司和 利未 人照各自的班次，按各自的職分獻燔祭和平安祭，又在耶和華殿 的門內事奉，稱謝頌讚耶和華。
2CHR|31|3|王又從自己的產業中分出一份來作燔祭，就是早晚的燔祭，和安息日、初一，以及節期的燔祭，都是按耶和華律法上所記載的。
2CHR|31|4|他又吩咐住 耶路撒冷 的百姓將祭司和 利未 人所應得的份給他們，使他們堅守耶和華的律法。
2CHR|31|5|命令一出， 以色列 人就把初熟的五穀、新酒、新油、蜜和田地的出產多多送來；他們把各樣出產的十分之一大量送來。
2CHR|31|6|住 猶大 各城的 以色列 人和 猶大 人也將牛羊的十分之一，以及分別為聖歸耶和華－他們上帝之物，就是十分取一之物，盡都送來，積成一堆一堆；
2CHR|31|7|他們從三月開始堆積，到七月才完成。
2CHR|31|8|希西家 和眾領袖來，看見這些堆積物，就稱頌耶和華，又為耶和華的百姓 以色列 祝福。
2CHR|31|9|希西家 向祭司和 利未 人查問這些堆積物。
2CHR|31|10|撒督 家的 亞撒利雅 祭司長告訴他說：「自從禮物開始送到耶和華的殿以來，我們不但吃飽，而且剩下的很多；因為耶和華賜福給他的百姓，所剩下的才這樣豐盛。」
2CHR|31|11|希西家 吩咐要在耶和華殿裏預備倉房，他們就預備了。
2CHR|31|12|他們誠心將禮物，十分取一之物，就是分別為聖之物，都搬入倉內。 利未 人 歌楠雅 主管這事，他的兄弟 示每 是副主管。
2CHR|31|13|耶歇 、 亞撒細雅 、 拿哈 、 亞撒黑 、 耶利摩 、 約撒拔 、 以列 、 伊斯瑪基雅 、 瑪哈 、 比拿雅 都是督辦，在 歌楠雅 和他兄弟 示每 的手下，是 希西家 王和管理上帝殿的 亞撒利雅 所委派的。
2CHR|31|14|守東門的 利未 人 音拿 的兒子 可利 ，掌管獻給上帝的甘心祭，發放獻給耶和華的禮物和至聖的物。
2CHR|31|15|在祭司的各城裏，在他手下忠心協助他的有 伊甸 、 (王民)雅(王民) 、 耶書亞 、 示瑪雅 、 亞瑪利雅 、 示迦尼雅 ，都按著班次分給他們的弟兄，無論大小，
2CHR|31|16|不論是否登錄在家譜，凡三歲以上的男丁，每日進耶和華殿、按班次供職事奉的，都分給他，
2CHR|31|17|也發放給按父家登錄在家譜的祭司；又按班次職任分給二十歲以上的 利未 人，
2CHR|31|18|又按家譜的登記，分給他們的小孩、妻子、兒女，給全體會眾；因為他們忠誠，將自己分別為聖。
2CHR|31|19|住在各城郊野 亞倫 的子孫、按名受委任的人，要把應得的份給祭司中所有的男丁和載入家譜的 利未 人。
2CHR|31|20|希西家 在全 猶大 都這樣辦理，在耶和華－他上帝面前行良善、正直、忠誠的事。
2CHR|31|21|凡他所行的，無論是開始辦上帝殿的事，是遵律法守誡命，是尋求他的上帝，他都盡心去做，無不亨通。
2CHR|32|1|在這些虔誠的事以後， 亞述 王 西拿基立 來侵犯 猶大 ，圍困堅固城，想要攻破它們。
2CHR|32|2|希西家 見 西拿基立 來，定意要攻打 耶路撒冷 ，
2CHR|32|3|就與領袖和勇士商議，塞住城外的泉源；他們都幫助他。
2CHR|32|4|於是許多百姓聚集，塞住一切泉源，以及國中流通的小河，說：「 亞述 諸王來，為何讓他們得著許多水呢？」
2CHR|32|5|希西家 奮勇自強，修築所有毀壞的城牆，升高城樓，又在城外築另一片城牆，堅固 大衛城 的 米羅 ，製造許多兵器和盾牌。
2CHR|32|6|他設立軍事將領管理百姓，召集他們在城門的廣場，勉勵他們，說：
2CHR|32|7|「你們當剛強壯膽，不要因 亞述 王和跟隨他的大軍恐懼驚慌，因為與我們同在的，比與他們同在的更大。
2CHR|32|8|與他們同在的是血肉之臂，但與我們同在的是耶和華－我們的上帝，他必幫助我們，為我們爭戰。」百姓因 猶大 王 希西家 的話就得到鼓勵。
2CHR|32|9|此後， 亞述 王 西拿基立 和跟隨他的全軍攻打 拉吉 ，派臣僕到 耶路撒冷 見 猶大 王 希西家 和所有在 耶路撒冷 的 猶大 人，說：
2CHR|32|10|「 亞述 王 西拿基立 如此說：『你們倚靠甚麼，還留在 耶路撒冷 受困嗎？
2CHR|32|11|希西家 說：耶和華－我們的上帝必救我們脫離 亞述 王的手，這不是誘惑你們，使你們受飢渴而死嗎？
2CHR|32|12|希西家 豈不是將耶和華的丘壇和祭壇廢去，並且吩咐 猶大 與 耶路撒冷 的人說：你們當在一個壇前敬拜，在其上燒香嗎？
2CHR|32|13|我與我祖先向列邦民族所行的，你們豈不知道嗎？列邦的神明何嘗能救自己的國脫離我的手呢？
2CHR|32|14|我祖先所滅的那些國的神明，有誰能救自己的百姓脫離我的手呢？難道你們的上帝能救你們脫離我的手嗎？
2CHR|32|15|現在，不要讓 希西家 這樣欺騙你們，誘惑你們，也不要相信他，因為沒有一國一邦的神明能救自己的百姓脫離我的手和我祖先的手，你們的上帝也絕不能救你們脫離我的手。』」
2CHR|32|16|西拿基立 的臣僕還說了一些話來毀謗耶和華上帝和他的僕人 希西家 。
2CHR|32|17|西拿基立 也寫信毀謗耶和華－ 以色列 的上帝，說：「列邦的神明既不能救自己的百姓脫離我的手， 希西家 的上帝也不能救他的百姓脫離我的手。」
2CHR|32|18|亞述 王的臣僕用 猶大 話向 耶路撒冷 城牆上的百姓大聲呼喊，要恐嚇他們，擾亂他們，以便取城。
2CHR|32|19|他們談論 耶路撒冷 的上帝，如同談論世上人手所造的神明一樣。
2CHR|32|20|希西家 王和 亞摩斯 的兒子 以賽亞 先知為此禱告，向天呼求。
2CHR|32|21|耶和華就差遣一個使者進入 亞述 王的營中，把所有大能的勇士、官長和將領盡都滅了。 亞述 王滿面羞愧地回到本國，進了他神明的廟中，他幾個親生的兒子在那裏用刀殺了他。
2CHR|32|22|這樣，耶和華救 希西家 和 耶路撒冷 的居民脫離 亞述 王 西拿基立 的手，也脫離一切仇敵的手，又賜他們四境平安 。
2CHR|32|23|有許多人到 耶路撒冷 將供物獻與耶和華，又將寶物送給 猶大 王 希西家 。自此之後， 希西家 在列國人的眼中受人尊崇。
2CHR|32|24|那些日子， 希西家 病得要死，就向耶和華禱告，耶和華應允他，賜他一個預兆。
2CHR|32|25|希西家 卻沒有照他所蒙的恩回報，因他心裏驕傲，所以憤怒要臨到他，臨到 猶大 和 耶路撒冷 。
2CHR|32|26|但 希西家 和 耶路撒冷 的居民為了心裏驕傲，就一同謙卑，以致耶和華的憤怒在 希西家 的日子沒有臨到他們。
2CHR|32|27|希西家 大有財富和尊榮，他為自己建造府庫，收藏金銀、寶石、香料、盾牌和各樣的寶器，
2CHR|32|28|又建造倉房，收藏五穀、新酒和新的油，又為各類牲畜蓋棚立圈，
2CHR|32|29|並且為自己建立城鎮，也擁有許多的羊群牛群，因為上帝賜他極多的財產。
2CHR|32|30|這 希西家 也塞住 基訓 的上源，引水直下，流在 大衛城 的西邊。 希西家 所行的事盡都亨通。
2CHR|32|31|但當 巴比倫 諸侯差遣使者來見 希西家 ，詢問國中所發生的奇事時，上帝離開他，要考驗他，好知道他心裏的一切。
2CHR|32|32|希西家 其餘的事和他的善行，看哪，都寫在 亞摩斯 的兒子 以賽亞 先知的《默示書》上和《猶大和以色列諸王記》上。
2CHR|32|33|希西家 與他祖先同睡，葬在 大衛 子孫陵墓的斜坡上。他死的時候， 猶大 眾人和 耶路撒冷 的居民都向他致敬。他的兒子 瑪拿西 接續他作王。
2CHR|33|1|瑪拿西 登基的時候年十二歲，在 耶路撒冷 作王五十五年。
2CHR|33|2|他行耶和華眼中看為惡的事，效法耶和華在 以色列 人面前趕出的列國那些可憎的事。
2CHR|33|3|他重新建築他父親 希西家 所拆毀的丘壇，為諸 巴力 築壇，造 亞舍拉 ，又敬拜天上的萬象，事奉它們。
2CHR|33|4|他在耶和華殿中築壇，耶和華曾指著這殿說：「我的名必永遠在 耶路撒冷 。」
2CHR|33|5|他在耶和華殿的兩個院子為天上的萬象築壇，
2CHR|33|6|並在 欣嫩子谷 使他的兒子經火，又觀星象，行法術，行邪術，求問招魂的和行巫術的，多行耶和華眼中看為惡的事，惹他發怒。
2CHR|33|7|他在上帝殿內立雕刻的偶像；上帝曾對 大衛 和他兒子 所羅門 說：「我在 以色列 眾支派中所選擇的 耶路撒冷 和這殿，必立我的名，直到永遠。
2CHR|33|8|只要 以色列 人謹守遵行我藉 摩西 吩咐他們的一切律法、律例、典章，我就不再使他們的腳挪移，離開我所賜給他們列祖之土地。」
2CHR|33|9|瑪拿西 引誘 猶大 和 耶路撒冷 的居民行惡，比耶和華在 以色列 人面前所滅的列國更嚴重。
2CHR|33|10|耶和華警戒 瑪拿西 和他的百姓，他們卻不聽。
2CHR|33|11|所以耶和華使 亞述 王的將領來攻擊他們，用手銬銬住 瑪拿西 ，用銅鏈鎖住他，把他帶到 巴比倫 去。
2CHR|33|12|他在急難的時候懇求耶和華－他的上帝，並在他列祖的上帝面前極其謙卑。
2CHR|33|13|他祈禱耶和華，耶和華就應允他，垂聽他的禱告，使他歸回 耶路撒冷 ，仍坐王位。 瑪拿西 這才知道惟獨耶和華是上帝。
2CHR|33|14|此後， 瑪拿西 在 大衛城 外，從谷內 基訓 西邊直到 魚門 口，建築城牆，環繞 俄斐勒 ；這牆建得很高。他又在 猶大 各堅固城內設立將領。
2CHR|33|15|他除掉外邦人的神像與耶和華殿中的偶像，又將他在耶和華殿的山上和 耶路撒冷 所築的各壇都拆毀，拋在城外。
2CHR|33|16|他重修耶和華的祭壇，在壇上獻平安祭和感謝祭，並吩咐 猶大 人事奉耶和華－ 以色列 的上帝。
2CHR|33|17|百姓卻仍在丘壇上獻祭，不過，他們只獻給耶和華－他們的上帝。
2CHR|33|18|瑪拿西 其餘的事和他向上帝的禱告，以及先見奉耶和華－ 以色列 上帝的名警戒他的話，看哪，都在《以色列諸王記》上。
2CHR|33|19|他的禱告，上帝怎樣應允他，他未謙卑以前的一切罪愆過犯，以及在何處建築丘壇，設立 亞舍拉 和雕刻的偶像，看哪，都寫在 何賽 的書上。
2CHR|33|20|瑪拿西 與他祖先同睡，葬在自己的宮中，他兒子 亞們 接續他作王。
2CHR|33|21|亞們 登基的時候年二十二歲，在 耶路撒冷 作王二年。
2CHR|33|22|他行耶和華眼中看為惡的事，效法他父親 瑪拿西 所行的，祭祀他父親 瑪拿西 所雕刻的一切偶像，事奉它們，
2CHR|33|23|但他不像他父親 瑪拿西 在耶和華面前那樣謙卑下來。這 亞們 的罪越犯越大。
2CHR|33|24|他的臣僕背叛他，在宮裏殺了他。
2CHR|33|25|但這地的百姓殺了所有背叛 亞們 王的人；這地的百姓立他兒子 約西亞 接續他作王。
2CHR|34|1|約西亞 登基的時候年八歲，在 耶路撒冷 作王三十一年。
2CHR|34|2|他行耶和華眼中看為正的事，行他祖先 大衛 所行的道，不偏左右。
2CHR|34|3|他作王第八年，尚且年輕，就尋求他祖先 大衛 的上帝。到了十二年，他開始潔淨 猶大 和 耶路撒冷 ，除掉丘壇、 亞舍拉 、雕刻的像和鑄造的像。
2CHR|34|4|眾人在他面前拆毀諸 巴力 的壇，砍斷壇上高高的香壇，又把 亞舍拉 和雕刻的像，以及鑄造的像打碎成灰，撒在向偶像獻祭之人的墳上，
2CHR|34|5|把祭司的骸骨燒在他們的壇上，潔淨了 猶大 和 耶路撒冷 。
2CHR|34|6|他又在 瑪拿西 、 以法蓮 、 西緬 、 拿弗他利 各城和四圍的廢墟 ，
2CHR|34|7|拆毀祭壇，把 亞舍拉 和雕刻的像打碎成灰，砍斷 以色列 全地所有的香壇。於是他回 耶路撒冷 去了。
2CHR|34|8|約西亞 王十八年，這地和殿潔淨了之後，他派 亞薩利雅 的兒子 沙番 、 瑪西雅 市長、 約哈斯 的兒子 約亞 史官去整修耶和華－他上帝的殿。
2CHR|34|9|他們去見 希勒家 大祭司，把奉到上帝殿的銀子交給他；這銀子是看守殿門的 利未 人從 瑪拿西 、 以法蓮 ，和 以色列 所有倖存的人，以及 猶大 、 便雅憫 眾人和 耶路撒冷 的居民收來的。
2CHR|34|10|他們把這銀子交給耶和華殿裏督工的，由他們轉交整修耶和華殿的工匠，
2CHR|34|11|就是交給木匠和石匠，好為 猶大 王所毀壞的殿，買鑿成的石頭和作鉤子與棟梁的木料。
2CHR|34|12|這些人辦事誠實，管理他們的是 利未 人 米拉利 的子孫 雅哈 和 俄巴底 ，又有 哥轄 人 撒迦利亞 和 米書蘭 ；還有所有善於奏樂的 利未 人。
2CHR|34|13|他們監督扛抬的人，督導一切做各樣工的人。 利未 人中也有作書記、官員、守衛的。
2CHR|34|14|他們把奉到耶和華殿的銀子運出來的時候， 希勒家 祭司發現了耶和華藉 摩西 所傳的律法書。
2CHR|34|15|希勒家 對 沙番 書記說：「我在耶和華殿裏發現了律法書。」 希勒家 把書遞給 沙番 。
2CHR|34|16|沙番 把書拿到王那裏，又把這事回覆王說：「凡交給僕人的手所辦的事，他們都辦好了。
2CHR|34|17|耶和華殿裏所發現的銀子已經倒出來，交在督工和工匠的手裏了。」
2CHR|34|18|沙番 書記又向王報告說：「 希勒家 祭司遞給我一卷書。」 沙番 就在王面前朗讀那書。
2CHR|34|19|王聽見律法的話，就撕裂衣服。
2CHR|34|20|王吩咐 希勒家 與 沙番 的兒子 亞希甘 、 米迦 的兒子 亞比頓 、 沙番 書記和王的臣僕 亞撒雅 ，說：
2CHR|34|21|「你們去，以所發現這書上的話，為我、為 以色列 和 猶大 倖存的人求問耶和華；因為我們的祖先沒有遵守耶和華的話，沒有照這書上所記的一切去做，耶和華的烈怒就倒在我們身上。」
2CHR|34|22|於是， 希勒家 和王的人 都去見 戶勒大 女先知，她是掌管禮服的 沙龍 的妻子， 沙龍 是 哈斯拉 的孫子， 特瓦 的兒子。 戶勒大 住在 耶路撒冷 第二區。他們向她說明來意。
2CHR|34|23|她對他們說：「耶和華－ 以色列 的上帝如此說：『你們可以回覆那派你們來見我的人說，
2CHR|34|24|耶和華如此說：看哪，我必照著在 猶大 王面前所讀那書上記載的一切詛咒，降禍於這地方和其上的居民。
2CHR|34|25|因為他們離棄我，向別神燒香，用他們手所做的一切惹我發怒，所以我的憤怒必倒在這地方，總不止息。』
2CHR|34|26|然而，派你們來求問耶和華的 猶大 王，你們要這樣回覆他：『耶和華－ 以色列 的上帝如此說：至於你所聽見的話，
2CHR|34|27|就是聽見我指著這地方和其上居民所說的話，你的心就軟化，在我面前謙卑下來，撕裂衣服，向我哭泣，因此我應允你。這是耶和華說的。
2CHR|34|28|看哪，我必使你歸到你祖先那裏，平安地進入墳墓，我要降於這地方和其上居民的一切災禍，你不會親眼看見。』」他們就去把這話回覆王。
2CHR|34|29|王派人召集 猶大 和 耶路撒冷 的眾長老來。
2CHR|34|30|王和 猶大 眾人、 耶路撒冷 的居民、祭司、 利未 人，以及所有的百姓，無論大小，都一同上到耶和華的殿去；王把殿裏所發現的約書上面一切的話讀給他們聽。
2CHR|34|31|王站在自己的位上，在耶和華面前立約，要盡心盡性跟從耶和華，遵守他的誡命、法度、律例，實行這書上所記這約的話；
2CHR|34|32|又使所有住 耶路撒冷 和 便雅憫 的人都服從這約。於是 耶路撒冷 的居民都遵行上帝，就是他們列祖之上帝的約。
2CHR|34|33|約西亞 從 以色列 各處把一切可憎之物盡都除掉，使 以色列 境內的人都事奉耶和華－他們的上帝。 約西亞 在世的日子，眾人都跟從耶和華－他們列祖的上帝，總不離開。
2CHR|35|1|約西亞 在 耶路撒冷 向耶和華守逾越節。正月十四日，他們宰了逾越節的羔羊。
2CHR|35|2|王分派祭司各盡其職，又勉勵他們辦耶和華殿中的事。
2CHR|35|3|他對那歸耶和華為聖、教導 以色列 眾人的 利未 人說：「你們將聖約櫃安放在 以色列 王 大衛 兒子 所羅門 建造的殿裏，不必再用肩扛抬。現在你們要服事耶和華－你們的上帝和他的百姓 以色列 。
2CHR|35|4|你們應當按著父家，照著班次，遵照 以色列 王 大衛 和他兒子 所羅門 所寫的，預備自己。
2CHR|35|5|要按著你們百姓的弟兄、父家的班次，侍立在聖所；每父家的班次中要有幾個 利未 人。
2CHR|35|6|要宰逾越節的羔羊，將自己分別為聖，為你們的弟兄預備，好遵守耶和華藉 摩西 所吩咐的話。」
2CHR|35|7|約西亞 從群畜中賜給所有在場的百姓，三萬隻小綿羊和小山羊，三千頭牛，作逾越節的祭物；這些都是出自王的產業。
2CHR|35|8|約西亞 的眾領袖也樂意把祭牲給百姓、祭司和 利未 人；管理上帝殿的 希勒家 、 撒迦利亞 、 耶歇 ，把二千六百隻羔羊和三百頭牛給祭司作逾越節的祭物。
2CHR|35|9|利未 人的族長 歌楠雅 和他兩個兄弟 示瑪雅 、 拿坦業 ，與 哈沙比雅 、 耶利 、 約撒拔 ，把五千隻羔羊和五百頭牛給 利未 人作逾越節的祭物。
2CHR|35|10|這樣，事奉的工作都安排好了，照王所吩咐的，祭司站在自己的位上， 利未 人按著班次侍立。
2CHR|35|11|他們宰了逾越節的羔羊，祭司從他們手裏接過血來 灑出去； 利未 人剝皮，
2CHR|35|12|把燔祭拿走，再按著父家的班次分給眾百姓，照 摩西 書上所寫的獻給耶和華；獻牛也是這樣。
2CHR|35|13|他們按著常例，用火烤逾越節的羔羊。至於其他的聖物，他們用盆，用鍋，用釜煮了，速速地送給眾百姓。
2CHR|35|14|然後他們為自己和祭司預備祭物，因為作祭司的 亞倫 子孫獻燔祭和脂肪，直到晚上。所以 利未 人為自己和作祭司的 亞倫 子孫預備。
2CHR|35|15|歌唱的 亞薩 子孫，照著 大衛 、 亞薩 、 希幔 和王的先見 耶杜頓 所吩咐的，站在自己的位上。守門的看守各門，不用離開他們的職守，因為他們的弟兄 利未 人給他們預備。
2CHR|35|16|當日，一切供奉耶和華、守逾越節，以及在耶和華壇上獻燔祭的事，都照 約西亞 王的吩咐預備好了。
2CHR|35|17|那時，在場的 以色列 人都守逾越節，又守除酵節七日。
2CHR|35|18|自從 撒母耳 先知的日子以來，在 以色列 中沒有守過這樣的逾越節， 以色列 諸王也沒有守過像 約西亞 、祭司、 利未 人、所有住 猶大 和 以色列 的人，以及 耶路撒冷 居民所守的逾越節。
2CHR|35|19|這逾越節是 約西亞 作王十八年時守的。
2CHR|35|20|約西亞 為殿做完這一切事以後， 埃及 王 尼哥 上來，要攻打靠近 幼發拉底河 的 迦基米施 ； 約西亞 出去迎擊他。
2CHR|35|21|他派使者來見 約西亞 ，說：「 猶大 王啊，我跟你有甚麼相干呢？我今日來不是要攻打你，而是要攻打與我爭戰之家，並且上帝吩咐我從速行事。你不要干預與我同在的上帝，免得他毀滅你。」
2CHR|35|22|約西亞 卻不轉臉離開他，反而改裝要與他打仗。他不聽從上帝藉 尼哥 的口所說的話，就來到 米吉多 平原爭戰。
2CHR|35|23|弓箭手射中 約西亞 王。王對他的臣僕說：「我受了重傷，你們載我離開戰場吧！」
2CHR|35|24|他的臣僕扶他下了戰車，上了他的副座車，送他到 耶路撒冷 。他就死了，葬在他祖先的墳墓裏。全 猶大 和 耶路撒冷 都哀悼 約西亞 。
2CHR|35|25|耶利米 為 約西亞 作哀歌，所有歌唱的男女也唱哀歌，追悼 約西亞 ，直到今日。他們在 以色列 中以此為定例；看哪，這些哀歌寫在《哀歌書》上。
2CHR|35|26|約西亞 其餘的事和他遵照耶和華律法上所記而行的善事，
2CHR|35|27|以及他自始至終所行的，看哪，都寫在《以色列和猶大列王記》上。
2CHR|36|1|這地的百姓立 約西亞 的兒子 約哈斯 在 耶路撒冷 接續他父親作王。
2CHR|36|2|約哈斯 登基的時候年二十三歲，在 耶路撒冷 作王三個月。
2CHR|36|3|埃及 王在 耶路撒冷 廢了他，又罰這地一百他連得銀子，一他連得金子。
2CHR|36|4|埃及 王 尼哥 立 約哈斯 的哥哥 以利雅敬 作 猶大 和 耶路撒冷 的王，給他改名叫 約雅敬 。 尼哥 卻將他的弟弟 約哈斯 帶到 埃及 去。
2CHR|36|5|約雅敬 登基的時候年二十五歲，在 耶路撒冷 作王十一年。他行耶和華－他上帝眼中看為惡的事。
2CHR|36|6|巴比倫 王 尼布甲尼撒 上來攻擊他，用銅鏈鎖著他，要把他帶到 巴比倫 去。
2CHR|36|7|尼布甲尼撒 又將耶和華殿裏的一些器皿帶到 巴比倫 ，放在 巴比倫 自己的宮裏 。
2CHR|36|8|約雅敬 其餘的事和他所行可憎的事，以及發生在他身上的事，看哪，都寫在《以色列和猶大列王記》上，他兒子 約雅斤 接續他作王。
2CHR|36|9|約雅斤 登基的時候年八歲 ，在 耶路撒冷 作王三個月十天，他行耶和華眼中看為惡的事。
2CHR|36|10|過了一年， 尼布甲尼撒 王差遣人將 約雅斤 和耶和華殿裏寶貴的器皿帶到 巴比倫 ，然後立 約雅斤 的叔父 西底家 作 猶大 和 耶路撒冷 的王。
2CHR|36|11|西底家 登基的時候年二十一歲，在 耶路撒冷 作王十一年。
2CHR|36|12|他行耶和華－他上帝眼中看為惡的事，沒有謙卑聽從 耶利米 先知所傳達耶和華的話。
2CHR|36|13|尼布甲尼撒 王曾叫他指著上帝起誓，他卻背叛，硬著頸項，內心頑固，不歸向耶和華－ 以色列 的上帝。
2CHR|36|14|眾祭司長和百姓也多多犯罪，效法列國一切可憎的事，玷污耶和華在 耶路撒冷 分別為聖的殿。
2CHR|36|15|耶和華－他們列祖的上帝因為愛惜自己的百姓和居所，一再差遣使者去警戒他們。
2CHR|36|16|他們卻嘲笑上帝的使者，藐視他的話，譏誚他的先知，以致耶和華向他的百姓大發烈怒，甚至無法可救。
2CHR|36|17|所以，耶和華使 迦勒底 人的王來攻擊他們，在他們聖殿裏用刀殺了他們的壯丁，不憐憫他們的少男少女、老人長者。耶和華把所有的人都交在他手裏。
2CHR|36|18|他把上帝殿裏一切的大小器皿與耶和華殿裏的財寶，以及王和眾領袖的財寶，全都帶到 巴比倫 去。
2CHR|36|19|迦勒底 人焚燒了上帝的殿，拆毀 耶路撒冷 的城牆，用火燒了城裏所有的宮殿，毀壞了城裏一切寶貴的器皿。
2CHR|36|20|凡脫離刀劍的倖存者， 迦勒底 王都擄到 巴比倫 去，作他和他子孫的僕婢，直到 波斯 國興起。
2CHR|36|21|這就應驗耶和華藉 耶利米 的口所說的話：地得享安息；在荒涼的日子，地就守安息，直到滿了七十年。
2CHR|36|22|波斯 王 居魯士 元年，耶和華為要應驗藉 耶利米 的口所說的話，就激發 波斯 王 居魯士 的心，使他下詔書通告全國，說：
2CHR|36|23|「 波斯 王 居魯士 如此說：耶和華－天上的上帝已將地上萬國賜給我，又委派我在 猶大 的 耶路撒冷 為他建造殿宇。你們中間凡作他子民的可以上去，願耶和華－他的上帝與他同在。」
