ECCL|1|1|在 耶路撒冷 作王、 大衛 的兒子、傳道者的言語。
ECCL|1|2|傳道者說：虛空的虛空， 虛空的虛空，全是虛空。
ECCL|1|3|人一切的勞碌， 就是他在日光之下的勞碌，有甚麼益處呢？
ECCL|1|4|一代過去，一代又來， 地卻永遠長存。
ECCL|1|5|太陽上升，太陽下落， 急歸所出之地。
ECCL|1|6|風往南颳，又向北轉， 不停旋轉，繞回原路。
ECCL|1|7|江河都往海裏流，海卻不滿； 江河從何處流，仍歸回原處。
ECCL|1|8|萬事令人厭倦， 人不能說盡。 眼看，看不飽； 耳聽，聽不足。
ECCL|1|9|已有的事，後必再有； 已行的事，後必再行。 日光之下並無新事。
ECCL|1|10|有一件事人指著說：「看，這是新的！」 它在我們以前的世代早已有了。
ECCL|1|11|已過的事，無人記念； 將來的事，後來的人也不記念。
ECCL|1|12|我傳道者在 耶路撒冷 作過 以色列 的王。
ECCL|1|13|我用智慧專心探尋、考察天下所發生的一切事：上帝給世人何等沉重的擔子，使他們在其中勞苦！
ECCL|1|14|我見日光之下所發生的一切事，看哪，全是虛空，全是捕風。
ECCL|1|15|彎曲的，不能變直； 缺乏的，不計其數。
ECCL|1|16|我心裏說：「看哪，我大有智慧，勝過在我以前所有統治 耶路撒冷 的人；我的心也多經歷智慧和知識的事。」
ECCL|1|17|我專心想要明白智慧，想要明白狂妄與愚昧，方知這也是捕風。
ECCL|1|18|因為多有智慧，就多有愁煩； 增加知識，就增加憂傷。
ECCL|2|1|我心裏說：「來吧，讓我用喜樂試試你，使你享福！」看哪，這也是虛空。
ECCL|2|2|論嬉笑，我說：「這是狂妄。」論享樂，「這有甚麼用呢？」
ECCL|2|3|我心以智慧引導我，我心裏探究，如何用酒使身體舒暢，如何抓住愚昧，直等我看明世人在天下短暫一生中，當行何事為美。
ECCL|2|4|我大興土木，為自己建造房屋，栽葡萄園，
ECCL|2|5|修造庭園和公園，在其中栽種各樣果樹，
ECCL|2|6|挖造水池，用以灌溉林中的幼樹。
ECCL|2|7|我買了僕婢，也有生在家中的僕婢；又有許多牛群羊群，勝過我以前所有在 耶路撒冷 的人。
ECCL|2|8|我為自己積蓄金銀，搜集各君王、各省份的財寶；又為自己得男女歌手和世人所喜愛的物，以及一個又一個的妃嬪。
ECCL|2|9|這樣，我就日漸昌盛，勝過我以前所有在 耶路撒冷 的人。我的智慧仍然存留。
ECCL|2|10|凡我眼所求的，我沒有克制它；我心所樂的，我沒有不享受。因我的心要為一切的勞碌快樂，這是我從一切勞碌中所得的報償 。
ECCL|2|11|後來，我回顧我手所經營的一切和我勞碌所做的工。看哪，全是虛空，全是捕風；在日光之下毫無益處。
ECCL|2|12|我轉而回顧智慧、狂妄和愚昧。在王以後來的人又如何呢？不過做先前所做的就是了。
ECCL|2|13|於是我看出智慧勝過愚昧，如同光明勝過黑暗。
ECCL|2|14|智慧人的眼目光明 ，愚昧人卻在黑暗裏行。但我知道他們都有相同的遭遇。
ECCL|2|15|我心裏就說：「愚昧人所遇見的，我也一樣遇見，那麼我何必更有智慧呢？」我心裏說：「這也是虛空。」
ECCL|2|16|智慧人和愚昧人一樣，不會長久被人記念，因為日後都被遺忘。可嘆！智慧人和愚昧人都一樣會死亡。
ECCL|2|17|於是我恨惡生命，因為在日光之下所發生的事我都以為煩惱，全是虛空，全是捕風。
ECCL|2|18|我恨惡一切的勞碌，就是我在日光之下所勞碌的，因為我所得的必須留給我以後的人。
ECCL|2|19|那人是智慧是愚昧，誰能知道呢？他竟要掌管我在日光之下用智慧勞碌所得的。這也是虛空。
ECCL|2|20|我轉想我在日光之下所勞碌的一切工作，心就絕望。
ECCL|2|21|因為有人用智慧、知識、靈巧勞碌工作，所得來的卻要遺留給未曾勞碌的人作產業。這也是虛空，大大不幸。
ECCL|2|22|人一切的勞碌操心，就是他在日光之下所勞碌的，又得著了甚麼呢？
ECCL|2|23|他日日憂慮，他的勞苦成為愁煩，連夜間心也不得休息。這也是虛空。
ECCL|2|24|難道一個人有吃有喝，且在勞碌中享福，不是福氣嗎？我看這也是出於上帝的手。
ECCL|2|25|論到吃用、享福，誰能勝過我呢？
ECCL|2|26|上帝喜愛誰，就給誰智慧、知識和喜樂；惟有罪人，上帝使他勞苦，將他所儲藏、所堆積的歸給上帝所喜愛的人。這也是虛空，也是捕風。
ECCL|3|1|凡事都有定期， 天下每一事務都有定時。
ECCL|3|2|生有時，死有時； 栽種有時，拔出 有時；
ECCL|3|3|殺戮有時，醫治有時； 拆毀有時，建造有時；
ECCL|3|4|哭有時，笑有時； 哀慟有時，跳舞有時；
ECCL|3|5|丟石頭有時，撿石頭有時； 懷抱有時，不抱有時；
ECCL|3|6|尋找有時，失落有時； 保存有時，拋棄有時；
ECCL|3|7|撕裂有時，縫補有時； 沉默有時，說話有時；
ECCL|3|8|喜愛有時，恨惡有時； 戰爭有時，和平有時。
ECCL|3|9|這樣，做事的人在他所勞碌的事上得到甚麼益處呢？
ECCL|3|10|我觀看上帝給世人的擔子，使他們在其中勞苦：
ECCL|3|11|上帝造萬物，各按其時成為美好，又將永恆安放在世人心裏；然而上帝從始至終的作為，人不能測透。
ECCL|3|12|我知道，人除了終身喜樂納福，沒有一件幸福的事。
ECCL|3|13|並且人人吃喝，在他的一切勞碌中享福，這也是上帝的賞賜。
ECCL|3|14|我知道上帝所做的都必存到永遠；無所增添，無所減少。上帝這樣做，是要人在他面前存敬畏的心。
ECCL|3|15|現今的事以前就有了，將來的事也早已有了，並且上帝使已過的事重新再來 。
ECCL|3|16|我又見日光之下，應有公平之處有奸惡，應有公義之處也有奸惡。
ECCL|3|17|我心裏說：「上帝必審判義人和惡人，因為在那裏，各樣事務，一切工作，都有定時。」
ECCL|3|18|我心裏說：「為世人的緣故，上帝考驗他們，讓他們看見自己不過像走獸一樣。」
ECCL|3|19|因為世人遭遇的，走獸也遭遇，所遭遇的都一樣：這個怎樣死，那個也怎樣死，他們都有一樣的氣息。人不能強於走獸，全是虛空；
ECCL|3|20|都歸一處，都是出於塵土，也都歸於塵土。
ECCL|3|21|誰知道人的氣息是往上升，走獸的氣息是下入地呢？
ECCL|3|22|總而言之，人能夠在他經營的事上喜樂，是最好不過了，因為這是他應得的報償。他身後的事誰能領他回來看呢？
ECCL|4|1|我轉而觀看日光之下所發生的一切欺壓之事。看哪，受欺壓的流淚，無人安慰；欺壓他們的有權勢，也無人安慰。
ECCL|4|2|因此，我讚歎那已死的死人，勝過那還活著的活人。
ECCL|4|3|但那尚未出生，就是未曾見過日光之下所發生之惡事的，比這兩種人更幸福。
ECCL|4|4|我見人因彼此嫉妒而有一切的勞碌和各樣工作的成就，這也是虛空，也是捕風。
ECCL|4|5|愚昧人抱著雙臂， 自食其肉。
ECCL|4|6|一掌滿滿而得享安靜， 勝過兩掌滿滿而勞碌捕風。
ECCL|4|7|我轉而觀看日光之下有一件虛空的事：
ECCL|4|8|有人孤單無雙，無子無兄弟，竟勞碌不息，眼目也不以財富為滿足。他說：「我勞碌，自己卻不享福，到底是為了誰呢？」這也是虛空，是極沉重的擔子。
ECCL|4|9|兩個人總比一個人好，他們勞碌同得美好的報償。
ECCL|4|10|若是跌倒，這人可以扶起他的同伴；倘若孤身跌倒，沒有別人扶起他來，這人就有禍了。
ECCL|4|11|再者，二人同睡就都暖和，一人獨睡怎能暖和呢？
ECCL|4|12|若遇敵攻擊，孤身難擋，二人就能抵擋他；三股合成的繩子不易折斷。
ECCL|4|13|貧窮而有智慧的年輕人，勝過年老不再納諫的愚昧王，
ECCL|4|14|那人從監牢裏出來作王，在國中原是出身貧寒。
ECCL|4|15|我見日光之下所有行走的活人，都跟隨那年輕人，就是接續作王的那位。
ECCL|4|16|他的百姓，就是他所治理的眾人，多得無數；但後來的人還是不喜歡他。這也是虛空，也是捕風。
ECCL|5|1|你到上帝的殿要謹慎你的腳步；近前聽，勝過愚昧人獻祭，他們不知道自己在作惡。
ECCL|5|2|在上帝面前你不可冒失開口，也不可心急發言；因為上帝在天上，你在地上，所以你的話語要少。
ECCL|5|3|事務多，令人做夢；話語多，顯出愚昧。
ECCL|5|4|你向上帝許願，還願不可遲延，因他不喜歡愚昧人，你許的願應當償還。
ECCL|5|5|你許願不還，不如不許。
ECCL|5|6|不可放任你的口使肉體犯罪，也不可在使者 面前說是錯許了。為何使上帝因你的聲音發怒，敗壞你手所做的呢？
ECCL|5|7|多夢多言，其中多有虛空，你只要敬畏上帝。
ECCL|5|8|你若在一個地區看見窮人受欺壓，公義公平被掠奪，不要因此驚奇；有一位高過居高位的在鑒察，在他們之上還有更高的。
ECCL|5|9|況且地的益處歸眾人，就是君王也受田地的供應。
ECCL|5|10|喜愛銀子的，不因得銀子滿足；喜愛財富的，也不因得利益知足。這也是虛空。
ECCL|5|11|貨物增添，吃的人也增添，物主得甚麼益處呢？不過眼看而已！
ECCL|5|12|勞碌的人不拘吃多吃少，睡得香甜；富人的豐足卻不容他睡覺。
ECCL|5|13|我見日光之下有一件令人憂傷的禍患，就是財主積存財富，反害自己。
ECCL|5|14|他因遭遇不幸 ，財產盡失；他生了兒子，手裏卻一無所有。
ECCL|5|15|他怎樣從母胎赤身而來，也必照樣赤身而去；他所勞碌得來的，手中分毫不能帶去。
ECCL|5|16|這是一件令人憂傷的禍患。他來的時候怎樣，去的時候也必怎樣。他為風勞碌有甚麼益處呢？
ECCL|5|17|並且他終身在黑暗中吃喝 ，多有煩惱、病痛和怒氣。
ECCL|5|18|看哪，我所見為善為美的，就是人在上帝賜他一生的日子吃喝，享受日光之下勞碌得來的好處，因為這是他應得的報償。
ECCL|5|19|而且，一個人蒙上帝賞賜財富與資產，又使他能享用，能獲取自己當有的報償 ，在他的勞碌中喜樂，這是上帝的賞賜。
ECCL|5|20|他不多思念自己一生的日子，因為上帝使他的心充滿喜樂。
ECCL|6|1|我見日光之下有一件禍患重壓在人身上，
ECCL|6|2|就是人蒙上帝賜他財富、資產和尊榮，以致他心裏所願的一樣都不缺，只是上帝使他不能享用，反被外人享用。這是虛空，也是禍患。
ECCL|6|3|人若生一百個兒子，活許多歲數；他即使壽命很長，心裏卻不因福樂而滿足，又不得埋葬；我說，那流掉的胎比他倒好。
ECCL|6|4|因為這胎虛虛而來，暗暗而去，名字被黑暗遮蔽，
ECCL|6|5|而且沒有見過天日，甚麼都不知道，這胎比那人倒享安息。
ECCL|6|6|那人雖然活千年，再活千年，卻不能享福；眾人豈不都歸同一個地方去嗎？
ECCL|6|7|人的勞碌都為口腹，心裏卻不知足。
ECCL|6|8|智慧人比愚昧人有甚麼益處呢？困苦人在眾人面前知道如何行，有甚麼益處呢？
ECCL|6|9|眼睛所看的比心裏妄想的倒好。這也是虛空，也是捕風。
ECCL|6|10|先前所有的，早已起了名，人早知道人是如何的，不能與比自己強壯的相爭。
ECCL|6|11|話語多，虛空也增多，這對人有甚麼益處呢？
ECCL|6|12|人一生虛度的日子，如影兒經過，誰知道甚麼才是對他有益呢？誰能告訴他身後在日光之下會發生甚麼事呢？
ECCL|7|1|名譽強如美好的膏油， 人死去的日子勝過他出生的日子。
ECCL|7|2|往喪家去， 強如往宴樂的家， 因為死是眾人的結局， 活人必將這事放在心上。
ECCL|7|3|憂愁強如喜笑， 因為面帶愁容，終必使心喜樂。
ECCL|7|4|智慧人的心在遭喪之家； 愚昧人的心在快樂之家。
ECCL|7|5|聽智慧人的責備， 強如聽愚昧人歌唱；
ECCL|7|6|因為愚昧人的笑聲， 好像鍋子下面燒荊棘的爆聲， 這也是虛空。
ECCL|7|7|勒索使智慧人變為愚妄， 賄賂能敗壞人的心。
ECCL|7|8|事情的終局強如它的起頭； 存心忍耐的，勝過居心驕傲的。
ECCL|7|9|你的心不要急躁惱怒， 因為惱怒存在愚昧人的懷中。
ECCL|7|10|不要說： 為甚麼先前的日子強過現今的日子呢？ 你這樣問不是出於智慧。
ECCL|7|11|智慧加上產業是美好的， 對見天日的人都有益處。
ECCL|7|12|因為智慧庇護人， 好像金錢庇護人一樣； 智慧能保全智慧者的生命， 這就是知識的益處。
ECCL|7|13|你要觀看上帝的作為， 誰能使他所彎曲的變直呢？
ECCL|7|14|順利時要喜樂；患難時當思考。上帝使這兩樣都發生，因此，人不知將會發生甚麼事。
ECCL|7|15|在虛度的日子裏，我見過各樣的事情，義人在他的義中滅亡，惡人在他的惡中倒享長壽。
ECCL|7|16|不要行義過分，也不要過於自逞智慧，何必自取敗亡呢？
ECCL|7|17|不要行惡過分，也不要為人愚昧，何必未到期而死呢？
ECCL|7|18|你持守這個，那個也不要鬆手才好。敬畏上帝的人，這一切都能兼得。
ECCL|7|19|智慧使擁有智慧的人比城中十個官長更有能力。
ECCL|7|20|其實世上沒有行善而不犯罪的義人。
ECCL|7|21|人所說的話，你不要都放在心上，免得聽見你的僕人詛咒你。
ECCL|7|22|因為你心裏知道，自己也曾屢次詛咒別人。
ECCL|7|23|我曾用智慧試驗這一切事，我說：「要得智慧。」智慧卻離我遠。
ECCL|7|24|萬事之理遙不可及，太深奧，誰能測透呢？
ECCL|7|25|我轉念，一心要知道，要考察，要尋求智慧和萬事的來由，要知道邪惡為愚昧，愚昧為狂妄。
ECCL|7|26|我發現有一種婦人比死還苦毒：她本身是陷阱，她的心是羅網，手是鎖鏈。凡蒙上帝喜愛的人必能躲開她；有罪的人卻被她纏住了。
ECCL|7|27|傳道者說：「你看，我考察一件又一件，為要尋求萬事的來由，這是我所尋得的：
ECCL|7|28|我繼續尋找，卻未找到；一千當中，我找到一個男的，但在這一切當中，卻找不到一個女的。
ECCL|7|29|你看，我所找到的只有一件，就是上帝造的人是正直的，但他們卻尋出許多詭計。」
ECCL|8|1|誰如 智慧人呢？ 誰知道事情的解釋呢？ 人的智慧使他的臉發光， 改變他臉上的暴戾之氣 。
ECCL|8|2|我勸你 因上帝誓言的緣故，當遵守王的命令。
ECCL|8|3|不要急躁離開王的面前，不要固執行惡，因為他凡事都隨自己心意而行。
ECCL|8|4|王的話本有權力，誰能對他說：「你在做甚麼？」
ECCL|8|5|凡遵守命令的，必不經歷禍患；智慧人的心知道適當的時機和必經的過程。
ECCL|8|6|各樣事務都有時機和過程，但人有苦難重壓在身。
ECCL|8|7|他不知道將來的事，其實將來如何，誰能告訴他呢？
ECCL|8|8|沒有人能掌握生命，將生命留住；也沒有人有權力掌管死期。這場爭戰無人能免；邪惡也不能救那行邪惡的人。
ECCL|8|9|這一切我都見過，我專心考察日光之下所發生的一切事，有時這人管轄那人，令他受害。
ECCL|8|10|我見惡人埋葬；從前他們進出聖地，他們在城中的作為被人忘記。這也是虛空。
ECCL|8|11|判罪之後不立刻執行，所以世人滿懷作惡的心思。
ECCL|8|12|罪人雖然作惡百次，倒享長壽；然而我也知道，福樂必臨到敬畏上帝的人，就是在他面前心存敬畏的人。
ECCL|8|13|惡人卻不得福樂，他的日子好像影兒不得長久，因為他不敬畏上帝。
ECCL|8|14|世上有一件虛空的事，就是義人所遭遇的，反而照惡人所做的；惡人所遭遇的，反而照義人所做的。我說，這也是虛空。
ECCL|8|15|我就稱讚快樂，原來人在日光之下，最大的福氣莫過於吃喝快樂；他在日光之下，上帝賜他一生的日子，要從勞碌中享受所得。
ECCL|8|16|我專心想要明白智慧，要觀看世上所發生的事。有人晝夜不得闔眼睡覺。
ECCL|8|17|我觀看上帝一切的作為，知道人不能探求日光之下所發生的事；任憑他費多少力探索，都找不出來，智慧人雖說他明白，仍不能找出來。
ECCL|9|1|我將這一切事放在心上，詳細研究這些，就知道義人和智慧人，並他們的作為都在上帝手中；或是愛，或是恨，都在他們面前，但人不能知道。
ECCL|9|2|凡臨到眾人的際遇都一樣：義人和惡人，好人 ，潔淨的人和不潔淨的人，獻祭的和不獻祭的，都一樣。好人如何，罪人也如何；起誓的如何，怕起誓的也如何。
ECCL|9|3|在日光之下發生的一切事中有一件禍患，就是眾人的際遇都一樣，並且世人的心充滿了惡；活著的時候心裏狂妄，後來就歸死人那裏去了。
ECCL|9|4|與一切活人相連的，那人還有指望，因為活著的狗勝過死了的獅子。
ECCL|9|5|活著的人知道必死；死了的人毫無所知，也不再得賞賜，因為他們的名 已被遺忘。
ECCL|9|6|他們的愛，他們的恨，他們的嫉妒，早就消滅了。在日光之下所發生的一切事，他們永不再有份了。
ECCL|9|7|你只管歡歡喜喜吃你的飯，心中快樂喝你的酒，因為上帝已經悅納你的作為。
ECCL|9|8|你的衣服要時時潔白，你頭上也不要缺少膏油。
ECCL|9|9|在你一生虛空的日子，就是上帝賜你在日光之下虛空 的日子，當與你所愛的妻快活度日，因為那是你一生中在日光之下勞碌所得的報償。
ECCL|9|10|凡你手所當做的事，要盡力去做；因為在你所必須去的陰間沒有工作，沒有謀算，沒有知識，也沒有智慧。
ECCL|9|11|我轉而回顧日光之下，快跑的未必能贏，強壯的未必戰勝，智慧的未必得糧食，聰明的未必得財富，有學問的未必得人喜悅，全在乎各人遇上的時候和機會。
ECCL|9|12|人不知道自己的定期。魚被險惡的網圈住，鳥被羅網捉住，禍患的時刻忽然臨到，世人陷在其中也是如此。
ECCL|9|13|我見日光之下有一樣智慧，在我看來是偉大的，
ECCL|9|14|就是有一人口稀少的小城，遇大君王前來攻擊，修築營壘，將城圍困。
ECCL|9|15|城中有一個貧窮的智慧人，他用智慧救了那城，卻沒有人記念那窮人。
ECCL|9|16|我就說，智慧勝過勇力；然而那貧窮人的智慧被人藐視，他的話也無人聽從。
ECCL|9|17|寧可聽智慧人安靜的話語，不聽掌權者在愚昧人中的喊聲。
ECCL|9|18|智慧勝過打仗的兵器；但一個罪人能敗壞許多善事。
ECCL|10|1|死蒼蠅使做香的膏油散發臭氣； 同樣，一點愚昧也能壓倒智慧和尊榮。
ECCL|10|2|智慧人的心居右； 愚昧人的心居左。
ECCL|10|3|愚昧人的行徑顯出無知， 對眾人說，他是愚昧人。
ECCL|10|4|掌權者的怒氣若向你發作， 不要離開你的本位， 因為鎮定能平息大過。
ECCL|10|5|我見日光之下有一件禍患， 似乎出於統治者的錯誤，
ECCL|10|6|就是愚昧人立在高位； 有錢人卻坐在低位。
ECCL|10|7|我見僕人騎馬， 王子像僕人在地上步行。
ECCL|10|8|挖陷坑的，自己必陷在其中； 拆城牆的，自己必被蛇咬。
ECCL|10|9|開鑿石頭的，會受損傷； 劈開木頭的，必遭危險。
ECCL|10|10|鐵器鈍了，若不將刃磨快，就必多費力氣； 但智慧的益處在於使人成功。
ECCL|10|11|尚未行法術，蛇若咬人， 行法術的人就得不到甚麼好處了。
ECCL|10|12|智慧人的口說出恩言； 愚昧人的嘴吞滅自己，
ECCL|10|13|他口中的話語起頭是愚昧， 終局是邪惡的狂妄。
ECCL|10|14|愚昧人多有話語。 人不知將來會發生甚麼事， 他身後的事誰能告訴他呢？
ECCL|10|15|愚昧人的勞碌使自己困乏， 連進城的路他也不知道。
ECCL|10|16|邦國啊，你的君王若年少， 你的群臣早晨宴樂， 你就有禍了！
ECCL|10|17|邦國啊，你的君王若是貴族之子， 你的群臣按時吃喝， 是為強身，不為酒醉， 你就有福了！
ECCL|10|18|因人懶惰，房頂塌下； 因人手懶，房屋滴漏。
ECCL|10|19|擺設宴席是為歡樂。 酒能使人快活， 錢能叫萬事應心。
ECCL|10|20|不可詛咒君王， 連起意也不可， 在臥室裏也不可詛咒富人； 因為空中的飛鳥必傳揚這聲音， 有翅膀的必述說這事。
ECCL|11|1|當將你的糧食撒在水面上， 因為日子久了，你必能得著它。
ECCL|11|2|將你所擁有的分給七人，或八人， 因為你不知道會有甚麼災禍臨到地上。
ECCL|11|3|雲若滿了雨，就必傾倒在地上。 樹向南倒，或向北倒， 樹倒在何處，就留在何處。
ECCL|11|4|看風的，必不撒種； 望雲的，必不收割。
ECCL|11|5|你不知道氣息如何進入孕婦的骨頭裏 ；照樣，造萬物之上帝的作為，你也無從得知。
ECCL|11|6|早晨要撒種，晚上也不要歇手，因為你不知道哪一樣發旺；前者或後者，或兩者都一樣好。
ECCL|11|7|光是甜美的，眼見日光是多麼好啊！
ECCL|11|8|人活多少年，就當快樂多少年，然而也當想到黑暗的日子；因為這樣的日子必多，所要來臨的全是虛空。
ECCL|11|9|年輕人哪，你在年少時當快樂；在年輕時使你的心歡暢，做你心所願做的，看你眼所愛看的；卻要知道，為這一切，上帝必審問你。
ECCL|11|10|所以，當從心中除掉愁煩，從肉體除去痛苦；因為年少和年輕之時，全是虛空。
ECCL|12|1|你趁著年輕、衰老的日子尚未來到，就是你所說，我毫無喜悅的那些歲月來臨之前，當記念造你的主。
ECCL|12|2|不要等到太陽、光明、月亮、星宿變為黑暗，雨後雲又返回；
ECCL|12|3|看守房屋的發顫，強壯的屈身，推磨的婦女因人少而停工，從窗戶往外看的眼光變為昏暗；
ECCL|12|4|街門關閉，推磨的聲音微小，鳥一叫，就驚醒，唱歌女子的聲音也都微弱；
ECCL|12|5|人怕高處，路上有驚慌；杏樹開花，蚱蜢成為重擔，慾望不再挑起；因為人歸他永遠的家，弔喪的在街上往來。
ECCL|12|6|不要等到銀鏈折斷 ，金罐破裂，瓶子在泉旁損壞，水輪在井口斷裂，
ECCL|12|7|塵土仍歸於地，像原來一樣，氣息仍歸於賜氣息的上帝。
ECCL|12|8|傳道者說：「虛空的虛空，全是虛空。」
ECCL|12|9|再者，傳道者因有智慧，將知識教導眾人；他思量，考察，並列舉出許多箴言。
ECCL|12|10|傳道者專心尋求可喜悅的言語，是憑正直寫的誠實話。
ECCL|12|11|智慧人的話語如同刺棒；這些嘉言好像釘穩的釘子，都是一個牧者所賜的。
ECCL|12|12|我兒，還有一點，你當受勸戒：著書多，沒有窮盡；讀書多，身體疲倦。
ECCL|12|13|這些事都已聽見了，結論就是：敬畏上帝，謹守他的誡命，這是人當盡的本分。
ECCL|12|14|因為人所做的事，連一切隱藏的事，無論是善是惡，上帝都必審問。
