1KGS|1|1|Et rex David senuerat habebat que aetatis plurimos dies; cum que operiretur vestibus, non calefiebat.
1KGS|1|2|Dixerunt ergo ei servi sui: " Quaeratur domino nostro regi adulescentula virgo et stet coram rege et curam eius agat dormiatque in sinu tuo et calefaciat dominum nostrum regem ".
1KGS|1|3|Quaesierunt igitur adulescentulam speciosam in omnibus finibus Israel et invenerunt Abisag Sunamitin et adduxerunt eam ad regem.
1KGS|1|4|Erat autem puella pulchra nimis et curam agebat regis et ministrabat ei; rex vero non cognovit eam.
1KGS|1|5|Adonias autem filius Haggith elevabatur dicens: " Ego regnabo! ". Fecitque sibi currum et equites et quinquaginta viros, qui ante eum currerent.
1KGS|1|6|Nec corripuit eum pater suus aliquando dicens: " Quare hoc fecisti? ". Erat autem et ipse pulcher valde, secundus natu post Absalom.
1KGS|1|7|Et sermo ei cum Ioab filio Sarviae et cum Abiathar sacerdote, qui adiuvabant partes Adoniae.
1KGS|1|8|Sadoc vero sacerdos et Banaias filius Ioiadae et Nathan propheta et Semei et Rei et robur exercitus David non erat cum Adonia.
1KGS|1|9|Immolatis ergo Adonias ovibus et vitulis et pinguibus iuxta lapidem Zoheleth, qui erat vicinus fonti Rogel, vocavit universos fratres suos filios regis et omnes viros Iudae servos regis;
1KGS|1|10|Nathan autem prophetam et Banaiam et robustos quosque et Salomonem fratrem suum non vocavit.
1KGS|1|11|Dixit itaque Nathan ad Bethsabee matrem Salomonis: " Num audisti quod regnaverit Adonias filius Haggith, et dominus noster David hoc ignorat?
1KGS|1|12|Nunc ergo veni, accipe a me consilium et salva animam tuam filiique tui Salomonis.
1KGS|1|13|Vade et ingredere ad regem David et dic ei: Nonne tu, domine mi rex, iurasti mihi ancillae tuae dicens: "Salomon filius tuus regnabit post me et ipse sedebit in solio meo"? Quare ergo regnat Adonias?
1KGS|1|14|Et, adhuc ibi te loquente cum rege, ego veniam post te et complebo sermones tuos ".
1KGS|1|15|Ingressa est itaque Bethsabee ad regem in cubiculo; rex autem senuerat nimis, et Abisag Sunamitis ministrabat ei.
1KGS|1|16|Inclinavit se Bethsabee et adoravit regem; ad quam rex: " Quid tibi, inquit, vis? ".
1KGS|1|17|Quae respondens ait: " Domine mi, tu iurasti per Dominum Deum tuum ancillae tuae: "Salomon filius tuus regnabit post me, et ipse sedebit in solio meo";
1KGS|1|18|et ecce nunc Adonias regnat, te, domine mi rex, ignorante.
1KGS|1|19|Mactavit boves et pinguia quaeque et oves plurimas et vocavit omnes filios regis, Abiathar quoque sacerdotem et Ioab principem militiae; Salomonem autem servum tuum non vocavit.
1KGS|1|20|Verumtamen, domine mi rex, in te oculi respiciunt totius Israel, ut indices eis quis sedere debeat in solio tuo, domine mi rex, post te.
1KGS|1|21|Eritque, cum dormierit dominus meus rex cum patribus suis, erimus ego et filius meus Salomon peccatores ".
1KGS|1|22|Adhuc illa loquente cum rege, Nathan propheta venit;
1KGS|1|23|et nuntiaverunt regi dicentes: " Adest Nathan propheta ". Cumque introisset ante conspectum regis et adorasset eum pronus in terram,
1KGS|1|24|dixit Nathan: " Domine mi rex, tu ergo dixisti: "Adonias regnet post me, et ipse sedeat super thronum meum"?
1KGS|1|25|Quia descendit hodie et immolavit boves et pinguia et arietes plurimos et vocavit universos filios regis et principes exercitus, Abiathar quoque sacerdotem; illique vescentes et bibentes coram eo dixerunt: "Vivat rex Adonias!".
1KGS|1|26|Me autem servum tuum et Sadoc sacerdotem et Banaiam filium Ioiadae et Salomonem famulum tuum non vocavit.
1KGS|1|27|Numquid a domino meo rege exivit hoc verbum, et mihi non indicasti servo tuo quis sessurus esset super thronum domini mei regis post eum? ".
1KGS|1|28|Et respondit rex David dicens: " Vocate ad me Bethsabee ". Quae cum fuisset ingressa coram rege et stetisset ante eum,
1KGS|1|29|iuravit rex et ait: " Vivit Dominus, qui eruit animam meam de omni angustia,
1KGS|1|30|quia, sicut iuravi tibi per Dominum, Deum Israel, dicens: Salomon filius tuus regnabit post me et ipse sedebit super solium meum pro me, sic faciam hodie ".
1KGS|1|31|Summissoque Bethsabee in terram vultu, adoravit regem dicens: " Vivat dominus meus rex David in aeternum! ".
1KGS|1|32|Dixit quoque rex David: " Vocate mihi Sadoc sacerdotem et Nathan prophetam et Banaiam filium Ioiadae ". Qui cum ingressi fuissent coram rege,
1KGS|1|33|dixit ad eos: " Tollite vobiscum servos domini vestri et imponite Salomonem filium meum, super mulam meam et ducite eum in Gihon,
1KGS|1|34|et ungat eum ibi Sadoc sacerdos et Nathan propheta in regem super Israel, et canetis bucina atque dicetis: "Vivat rex Salomon!".
1KGS|1|35|Et ascendetis post eum, et veniet et sedebit super solium meum, et ipse regnabit pro me; illique praecipiam, ut sit dux super Israel et super Iudam ".
1KGS|1|36|Et respondit Banaias filius Ioiadae regi dicens: " Amen, sic loquatur Dominus Deus domini mei regis.
1KGS|1|37|Quomodo fuit Dominus cum domino meo rege, sic sit cum Salomone et sublimius faciat solium eius a solio domini mei regis David ".
1KGS|1|38|Descendit ergo Sadoc sacerdos et Nathan propheta et Banaias filius Ioiadae et Cherethi et Phelethi, et imposuerunt Salomonem super mulam regis David et adduxerunt eum in Gihon.
1KGS|1|39|Sumpsitque Sadoc sacerdos cornu olei de tabernaculo et unxit Salomonem; et cecinerunt bucina, et dixit omnis populus: " Vivat rex Salomon! ".
1KGS|1|40|Et ascendit universa multitudo post eum, et populus canebat tibiis et laetabatur gaudio magno, et insonuit terra ad clamorem eorum.
1KGS|1|41|Audivit autem Adonias et omnes, qui invitati fuerant ab eo; iamque convivium finitum erat. Sed et Ioab, audita voce tubae, ait: " Quid sibi vult clamor civitatis tumultuantis? ".
1KGS|1|42|Adhuc illo loquente, Ionathan filius Abiathar sacerdotis venit; cui dixit Adonias: " Ingredere, quia vir strenuus es et bona nuntians ".
1KGS|1|43|Responditque Ionathan Adoniae: " Nequaquam! Dominus enim noster, rex David, regem constituit Salomonem
1KGS|1|44|misitque cum eo Sadoc sacerdotem et Nathan prophetam et Banaiam filium Ioiadae et Cherethi et Phelethi, et imposuerunt eum super mulam regis;
1KGS|1|45|unxeruntque eum Sadoc sacerdos et Nathan propheta regem in Gihon. Et ascenderunt inde laetantes, et insonuit civitas; haec est vox, quam audistis.
1KGS|1|46|Sed et Salomon sedit super solio regni,
1KGS|1|47|et ingressi servi regis benedixerunt domino nostro regi David dicentes: Amplificet Deus nomen Salomonis super nomen tuum et magnificet thronum eius super thronum tuum". Et adoravit rex in lectulo suo.
1KGS|1|48|Insuper et haec locutus est: "Benedictus Dominus, Deus Israel, qui dedit hodie sedentem in solio meo, videntibus oculis meis" ".
1KGS|1|49|Territi sunt ergo et surrexerunt omnes, qui invitati fuerant ab Adonia, et ivit unusquisque in viam suam.
1KGS|1|50|Adonias autem timens Salomonem surrexit et abiit tenuitque cornua altaris.
1KGS|1|51|Et nuntiaverunt Salomoni dicentes: " Ecce Adonias timens regem Salomonem tenuit cornua altaris dicens: "Iuret mihi hodie rex Salomon quod non interficiat servum suum gladio"".
1KGS|1|52|Dixitque Salomon: " Si fuerit vir bonus, non cadet ne unus quidem capillus eius in terram; sin autem malum inventum fuerit in eo, morietur.
1KGS|1|53|Misit ergo rex Salomon et eduxit eum ab altari, et ingressus adoravit regem Salomonem; dixitque ei Salomon: " Vade in domum tuam ".
1KGS|2|1|Appropinquaverant autem dies David ut moreretur, praecepit que Salomoni filio suo dicens:
1KGS|2|2|" Ego ingredior viam universae terrae; confortare et esto vir
1KGS|2|3|et observa decreta Domini Dei tui, ut ambules in viis eius et custodias statuta eius et praecepta eius et iudicia et testimonia, sicut scriptum est in lege Moysi, ut prospere agas in universis, quae facis et quocumque te verteris;
1KGS|2|4|ut confirmet Dominus sermonem suum, quem locutus est de me dicens: "Si custodierint filii tui viam suam et ambulaverint coram me in veritate, in omni corde suo et in omni anima sua, non auferetur tibi vir de solio Israel".
1KGS|2|5|Tu quoque nosti, quae fecerit mihi Ioab filius Sarviae, quae fecerit duobus principibus exercitus Israel, Abner filio Ner et Amasae filio Iether, quos occidit; et effudit sanguinem belli in pace et posuit cruorem proelii in balteo suo, qui erat circa lumbos eius, et in calceamento suo, quod erat in pedibus eius.
1KGS|2|6|Facies ergo iuxta sapientiam tuam et non deduces canitiem eius pacifice ad inferos.
1KGS|2|7|Sed filiis Berzellai Galaaditis reddes gratiam, eruntque comedentes in mensa tua; occurrerunt enim mihi, quando fugiebam a facie Absalom fratris tui.
1KGS|2|8|Habes quoque apud te Semei filium Gera de Beniamin de Bahurim, qui maledixit mihi maledictione pessima, quando ibam ad Mahanaim; sed quia descendit mihi in occursum ad Iordanem, et iuravi ei per Dominum dicens: Non te interficiam gladio.
1KGS|2|9|Tu noli pati esse eum innoxium; vir autem sapiens es et scies, quae facias ei deducesque canos eius cum sanguine ad infernum ".
1KGS|2|10|Dormivit igitur David cum patribus suis et sepultus est in civitate David.
1KGS|2|11|Dies autem, quibus regnavit David super Israel, quadraginta anni sunt: in Hebron regnavit septem annis, in Ierusalem triginta tribus.
1KGS|2|12|Salomon autem sedit super thronum David patris sui, et firmatum est regnum eius nimis.
1KGS|2|13|Et ingressus est Adonias filius Haggith ad Bethsabee matrem Salomonis, quae dixit ei: " Pacificusne ingressus tuus? ". Qui respondit: " Pacificus.
1KGS|2|14|Addiditque: " Sermo mihi est ad te ". Cui ait: " Loquere ". Et ille:
1KGS|2|15|" Tu, inquit, nosti quia meum erat regnum, et me proposuerat omnis Israel sibi in regem, sed translatum est regnum et factum est fratris mei; a Domino enim constitutum est ei.
1KGS|2|16|Nunc ergo petitionem unam deprecor a te; ne confundas faciem meam ". Quae dixit ad eum: " Loquere ".
1KGS|2|17|Et ille ait: " Precor, ut dicas Salomoni regi - neque enim negare tibi quidquam potest - ut det mihi Abisag Sunamitin uxorem ".
1KGS|2|18|Et ait Bethsabee: " Bene, ego loquar pro te regi ".
1KGS|2|19|Venit ergo Bethsabee ad regem Salomonem, ut loqueretur ei pro Adonia. Et surrexit rex in occursum eius adoravitque eam et sedit super thronum suum; positus quoque est thronus matri regis, quae sedit ad dexteram eius.
1KGS|2|20|Dixitque ei: " Petitionem unam parvulam ego deprecor a te; ne confundas faciem meam". Dixit ei rex: " Pete, mater mi, neque enim fas est, ut avertam faciem tuam ".
1KGS|2|21|Quae ait: " Detur Abisag Sunamitis Adoniae fratri tuo uxor ".
1KGS|2|22|Responditque rex Salomon et dixit matri suae: " Quare postulas Abisag Sunamitin Adoniae? Postula ei et regnum! Ipse est enim frater meus maior me et habet Abiathar sacerdotem et Ioab filium Sarviae ".
1KGS|2|23|Iuravit itaque rex Salomon per Dominum dicens: " Haec faciat mihi Deus et haec addat, certe contra animam suam locutus est Adonias verbum hoc.
1KGS|2|24|Et nunc, vivit Dominus, qui firmavit me et collocavit me super solium David patris mei et qui fecit mihi domum, sicut locutus est, certe hodie occidetur Adonias ".
1KGS|2|25|Misitque rex Salomon per manum Banaiae filii Ioiadae, qui interfecit eum, et mortuus est.
1KGS|2|26|Abiathar quoque sacerdoti dixit rex: " Vade in Anathoth ad agrum tuum; es quidem vir mortis, sed hodie te non interficiam, quia portasti arcam Domini Dei coram David patre meo et sustinuisti laborem in omnibus, in quibus laboravit pater meus ".
1KGS|2|27|Eiecit ergo Salomon Abiathar, ut non esset sacerdos Domini, ut impleretur sermo Domini, quem locutus est super domum Heli in Silo.
1KGS|2|28|Venit autem nuntius ad Ioab. Ioab autem declinaverat post Adoniam, cum post Absalom non declinasset; fugit ergo Ioab in tabernaculum Domini et apprehendit cornua altaris.
1KGS|2|29|Nuntiatumque est regi Salomoni, quod fugisset Ioab in tabernaculum Domini et esset iuxta altare; misitque Salomon Banaiam filium Ioiadae dicens: " Vade, interfice eum! ".
1KGS|2|30|Venit Banaias ad tabernaculum Domini et dixit ei: " Haec dicit rex: Egredere!". Qui ait: " Non egrediar, sed hic moriar ". Renuntiavit Banaias regi sermonem dicens: " Haec locutus est Ioab et haec respondit mihi ".
1KGS|2|31|Dixitque ei rex: " Fac, sicut locutus est, et interfice eum et sepeli; et amovebis sanguinem innocentem, qui effusus est a Ioab, a me et a domo patris mei.
1KGS|2|32|Et reddet Dominus sanguinem eius super caput eius, quia interfecit duos viros iustos melioresque se et occidit eos gladio, patre meo David ignorante: Abner filium Ner principem militiae Israel et Amasam filium Iether principem exercitus Iudae.
1KGS|2|33|Et revertetur sanguis illorum in caput Ioab et in caput seminis eius in sempiternum; David autem et semini eius et domui et throno illius sit pax usque in aeternum a Domino ".
1KGS|2|34|Ascendit itaque Banaias filius Ioiadae et aggressus eum interfecit; sepultusque est in domo sua in deserto.
1KGS|2|35|Et constituit rex Banaiam filium Ioiadae pro eo super exercitum et Sadoc sacerdotem posuit pro Abiathar.
1KGS|2|36|Misit quoque rex et vocavit Semei dixitque ei: " Aedifica tibi domum in Ierusalem et habita ibi et non egredieris inde huc atque illuc;
1KGS|2|37|quacumque autem die egressus fueris et transieris torrentem Cedron, scito te interficiendum; sanguis tuus erit super caput tuum ".
1KGS|2|38|Dixitque Semei regi: " Bonus sermo; sicut locutus est dominus meus rex, sic faciet servus tuus ". Habitavit itaque Semei in Ierusalem diebus multis.
1KGS|2|39|Factum est autem post annos tres, ut fugerent duo servi Semei ad Achis filium Maacha regem Geth; nuntiatumque est Semei quod servi eius essent in Geth.
1KGS|2|40|Et surrexit Semei et stravit asinum suum ivitque in Geth ad Achis ad requirendos servos suos et adduxit eos de Geth.
1KGS|2|41|Nuntiatum est autem Salomoni quod isset Semei in Geth de Ierusalem et redisset.
1KGS|2|42|Et mittens vocavit eum dixitque illi: " Nonne testificatus sum tibi per Dominum et praedixi tibi: Quacumque die egressus ieris huc et illuc, scito te esse moriturum? Et respondisti mihi "Bonus sermo; audivi".
1KGS|2|43|Quare ergo non custodisti iusiurandum Domini et praeceptum, quod praeceperam tibi? ".
1KGS|2|44|Dixitque rex ad Semei: " Tu nosti omne malum, cuius tibi conscium est cor tuum, quod fecisti David patri meo; reddit Dominus malitiam tuam in caput tuum.
1KGS|2|45|Et rex Salomon benedictus, et thronus David erit stabilis coram Domino usque in sempiternum ".
1KGS|2|46|Iussit itaque rex Banaiae filio Ioiadae, qui egressus percussit eum, et mortuus est. Confirmatum est igitur regnum in manu Salomonis.
1KGS|3|1|Et affinitate coniunctus est pharaoni regi Aegypti. Accepit namque filiam eius et adduxit in civitatem David, donec compleret aedificans domum suam et domum Domini et murum Ierusalem per circuitum.
1KGS|3|2|Attamen populus immolabat in excelsis; non enim aedificatum erat templum nomini Domini usque in diem illum.
1KGS|3|3|Dilexit autem Salomon Dominum ambulans in praeceptis David patris sui, excepto quod in excelsis immolabat et accendebat thymiama.
1KGS|3|4|Abiit itaque in Gabaon, ut immolaret ibi; illud quippe erat excelsum maximum. Mille hostias in holocaustum obtulit Salomon super altare illud.
1KGS|3|5|In Gabaon apparuit Dominus Salomoni per somnium nocte dicens: " Postula quod vis, ut dem tibi ".
1KGS|3|6|Et ait Salomon: " Tu fecisti cum servo tuo David patre meo misericordiam magnam, sicut ambulavit in conspectu tuo in veritate et iustitia et recto corde tecum; custodisti ei misericordiam tuam grandem et dedisti ei filium sedentem super thronum eius, sicut est hodie.
1KGS|3|7|Et nunc, Domine Deus meus, tu regnare fecisti servum tuum pro David patre meo. Ego autem sum puer parvus et ignorans egressum et introitum meum;
1KGS|3|8|et servus tuus in medio est populi, quem elegisti, populi infiniti, qui numerari et supputari non potest prae multitudine.
1KGS|3|9|Da ergo servo tuo cor docile, ut iudicare possit populum tuum et discernere inter bonum et malum. Quis enim potest iudicare populum tuum hunc multum? ".
1KGS|3|10|Placuit ergo sermo coram Domino quod Salomon rem huiuscemodi postulasset,
1KGS|3|11|et dixit Deus Salomoni: " Quia postulasti verbum hoc et non petisti tibi dies multos nec divitias aut animam inimicorum tuorum, sed postulasti tibi sapientiam ad discernendum iudicium,
1KGS|3|12|ecce feci tibi secundum sermones tuos et dedi tibi cor sapiens et intellegens, in tantum ut nullus ante te similis tui fuerit nec post te surrecturus sit;
1KGS|3|13|sed et haec, quae non postulasti, dedi tibi, divitias scilicet et gloriam, ut nemo fuerit similis tui in regibus cunctis diebus tuis.
1KGS|3|14|Si autem ambulaveris in viis meis et custodieris praecepta mea et mandata mea, sicut ambulavit David pater tuus, longos faciam dies tuos ".
1KGS|3|15|Igitur evigilavit Salomon et intellexit quod esset somnium. Cumque venisset Ierusalem, stetit coram arca foederis Domini et obtulit holocausta et fecit victimas pacificas et convivium universis famulis suis.
1KGS|3|16|Tunc venerunt duae mulieres meretrices ad regem steteruntque coram eo.
1KGS|3|17|Quarum una ait: " Obsecro, mi domine; ego et mulier haec habitabamus in domo una, et peperi apud eam in domo;
1KGS|3|18|tertia vero die, postquam ego peperi, peperit et haec; et eramus simul, nullusque alius nobiscum in domo, exceptis nobis duabus.
1KGS|3|19|Mortuus est autem filius mulieris huius nocte; dormiens quippe oppressit eum.
1KGS|3|20|Et consurgens intempesta nocte, silentio tulit filium meum de latere meo ancillae tuae dormientis et collocavit in sinu suo; suum autem filium, qui erat mortuus, posuit in sinu meo.
1KGS|3|21|Cumque surrexissem mane, ut darem lac filio meo, apparuit mortuus; quem diligentius intuens clara luce, deprehendi non esse meum, quem genueram ".
1KGS|3|22|Responditque altera mulier: " Non est ita, sed filius meus vivit, tuus autem mortuus est ". E contrario illa dicebat: " Mentiris. Filius quippe tuus mortuus est, meus autem vivit ". Atque in hunc modum contendebant coram rege.
1KGS|3|23|Tunc rex ait: " Haec dicit: "Filius meus vivit, et filius tuus mortuus est"; et ista respondit: "Non, sed filius tuus mortuus est, et filius meus vivit" ".
1KGS|3|24|Dixit ergo rex: " Afferte mihi gladium! ". Cumque attulissent gladium coram rege:
1KGS|3|25|" Dividite, inquit, infantem vivum in duas partes, et date dimidiam partem uni et dimidiam partem alteri ".
1KGS|3|26|Dixit autem mulier, cuius filius erat vivus, ad regem - commota sunt quippe viscera eius super filio suo -: " Obsecro, domine, date illi infantem vivum et nolite interficere eum ". E contrario illa dicebat: " Nec mihi nec tibi sit; dividatur ".
1KGS|3|27|Respondens rex ait: " Date huic infantem vivum, et non occidatur; haec est mater eius ".
1KGS|3|28|Audivit itaque omnis Israel iudicium, quod iudicasset rex; et timuerunt regem videntes sapientiam Dei esse in eo ad faciendum iudicium.
1KGS|4|1|Erat autem rex Salomon regnans super omnem Israel.
1KGS|4|2|Et hi principes quos habebat: Azarias filius Sadoc sacerdos;
1KGS|4|3|Elihoreph et Ahia filii Sisa scribae; Iosaphat filius Ahilud cancellarius;
1KGS|4|4|Banaias filius Ioiadae super exercitum; Sadoc autem et Abiathar sacerdotes;
1KGS|4|5|Azarias filius Nathan super praefectos; Zabud filius Nathan sacerdos amicus regis;
1KGS|4|6|et Ahisar praepositus domus et Adoniram filius Abda super tributa.
1KGS|4|7|Habebat autem Salomon duodecim praefectos super omnem Israel, qui praebebant annonam regi et domui eius; per singulos enim menses in anno singuli necessaria ministrabant.
1KGS|4|8|Et haec nomina eorum: Benhur in monte Ephraim;
1KGS|4|9|Bendecar in Maces et in Salebim et in Bethsames et in Elon et in Bethanan;
1KGS|4|10|Benhesed in Aruboth, ipsius erat Socho et omnis terra Epher;
1KGS|4|11|Benabinadab, cuius omnis regio Dor, Tapheth filiam Salomonis habebat uxorem;
1KGS|4|12|Baana filius Ahilud regebat Thanach et Mageddo et universam Bethsan, quae est iuxta Sarthan subter Iezrahel, a Bethsan usque Abelmehula et usque ultra Iecmaam;
1KGS|4|13|Bengaber in Ramoth Galaad habebat villas Iair filii Manasse in Galaad: ipse praeerat in omni regione Argob, quae est in Basan, sexaginta civitatibus magnis atque muratis, quae habebant seras aereas;
1KGS|4|14|Ahinadab filius Addo praeerat in Mahanaim;
1KGS|4|15|Achimaas in Nephthali, sed et ipse habebat Basemath filiam Salomonis in coniugio;
1KGS|4|16|Baana filius Chusai in Aser et in Baloth;
1KGS|4|17|Iosaphat filius Pharue in Issachar;
1KGS|4|18|Semei filius Ela in Beniamin;
1KGS|4|19|Gaber filius Uri in terra Galaad, in terra Sehon regis Amorraei et Og regis Basan, ut praefectus unus, qui erat in terra.
1KGS|4|20|Iuda et Israel innumerabiles, sicut arena maris in multitudine, comedentes et bibentes atque laetantes.
1KGS|5|1|Salomon autem erat in dicione sua habens omnia regna a Flu mine usque ad terram Philisthim et ad terminum Aegypti offerentium sibi munera et servientium ei cunctis diebus vitae eius.
1KGS|5|2|Erat autem cibus Salomonis per dies singulos triginta chori similae et sexaginta chori farinae,
1KGS|5|3|decem boves pingues et viginti boves pascuales et centum oves, excepta venatione cervorum, caprearum atque bubalorum et avium altilium.
1KGS|5|4|Ipse enim obtinebat omnem regionem, quae erat trans Flumen, a Thaphsa usque Gazam, et cunctos reges illarum regionum; et habebat pacem ex omni parte in circuitu.
1KGS|5|5|Habitabatque Iuda et Israel absque timore ullo, unusquisque sub vite sua et sub ficu sua a Dan usque Bersabee cunctis diebus Salomonis.
1KGS|5|6|Et habebat Salomon quattuor milia praesepia equorum currulium et duodecim milia equestres.
1KGS|5|7|Et praebebant supradicti praefecti necessaria mensae regis Salomonis et convivarum eius cum ingenti cura, unusquisque in suo mense.
1KGS|5|8|Hordeum quoque et paleas equorum et iumentorum deferebant in locum, ubi erat unicuique constitutum.
1KGS|5|9|Dedit quoque Deus sapientiam Salomoni et prudentiam multam nimis et latitudinem cordis quasi arenam, quae est in litore maris.
1KGS|5|10|Et praecedebat sapientia Salomonis sapientiam omnium Orientalium et Aegyptiorum;
1KGS|5|11|et erat sapientior cunctis hominibus, sapientior Ethan Ezrahita et Heman et Chalchol et Darda filiis Mahol et erat nominatus in universis gentibus per circuitum.
1KGS|5|12|Locutus est quoque Salomon tria milia parabolas, et fuerunt carmina eius quinque et mille.
1KGS|5|13|Et disputavit super lignis, a cedro, quae est in Libano, usque ad hyssopum, quae egreditur de pariete; et disseruit de iumentis et volucribus et reptilibus et piscibus.
1KGS|5|14|Et veniebant de cunctis populis ad audiendam sapientiam Salomonis, ab universis regibus terrae, qui audiebant sapientiam eius.
1KGS|5|15|Misit quoque Hiram rex Tyri servos suos ad Salomonem; audivit enim quod ipsum unxissent regem pro patre eius, quia amicus fuerat Hiram David omni tempore.
1KGS|5|16|Misit autem et Salomon ad Hiram dicens:
1KGS|5|17|" Tu scis voluntatem David patris mei et quia non potuerit aedificare domum nomini Domini Dei sui propter bella imminentia per circuitum, donec daret Dominus eos sub vestigio pedum eius.
1KGS|5|18|Nunc autem requiem dedit Dominus Deus meus mihi per circuitum; non est adversarius neque occursus malus.
1KGS|5|19|Quam ob rem cogito aedificare templum nomini Domini Dei mei, sicut locutus est Dominus David patri meo dicens: "Filius tuus, quem dabo pro te super solium tuum, ipse aedificabit domum nomini meo".
1KGS|5|20|Praecipe igitur, ut praecidant mihi cedros de Libano, et servi mei sint cum servis tuis; mercedem autem servorum tuorum dabo tibi quamcumque praeceperis; scis enim quoniam non est in populo meo vir, qui noverit ligna caedere sicut Sidonii ".
1KGS|5|21|Cum ergo audisset Hiram verba Salomonis, laetatus est valde et ait: " Benedictus Dominus hodie, qui dedit David filium sapientissimum super populum hunc plurimum ".
1KGS|5|22|Et misit Hiram ad Salomonem dicens: " Audivi, quaecumque mandasti mihi; ego faciam omnem voluntatem tuam in lignis cedrinis et abiegnis.
1KGS|5|23|Servi mei deponent ea de Libano ad mare, et ego componam ea in ratibus in mari usque ad locum, quem significaveris mihi, et applicabo ea ibi, et tu tolles ea; praebebisque necessaria mihi, ut detur cibus domui meae ".
1KGS|5|24|Itaque Hiram dabat Salomoni ligna cedrina et ligna abiegna iuxta omnem voluntatem eius.
1KGS|5|25|Salomon autem praebebat Hiram viginti milia chororum tritici in cibum domui eius et viginti choros purissimi olei; haec tribuebat Salomon Hiram per annos singulos.
1KGS|5|26|Dedit quoque Dominus sapientiam Salomoni, sicut locutus est ei; et erat pax inter Hiram et Salomonem, et percusserunt foedus ambo.
1KGS|5|27|Elegitque rex Salomon operas de omni Israel, et erat indictio triginta milia virorum.
1KGS|5|28|Mittebatque eos in Libanum decem milia per menses singulos vicissim, ita ut duobus mensibus essent in domibus suis; et Adoniram erat super huiuscemodi indictione.
1KGS|5|29|Fueruntque Salomoni septuaginta milia eorum, qui onera portabant, et octoginta milia latomorum in monte,
1KGS|5|30|absque praepositis, qui praeerant singulis operibus numero trium milium et trecentorum praecipientium populo, his, qui faciebant opus.
1KGS|5|31|Praecepitque rex, ut tollerent lapides grandes, lapides pretiosos in fundamentum templi, lapides quadratos;
1KGS|5|32|dolaverunt ergo caementarii Salomonis, caementarii Hiram et Giblii ligna et lapides et praeparaverunt ad aedificandam domum.
1KGS|6|1|Factum est igitur quadringente simo et octogesimo anno egres sionis filiorum Israel de terra Aegypti, in anno quarto, mense Ziv - ipse est mensis secundus - regni Salomonis super Israel, aedificare coepit domum Domino.
1KGS|6|2|Domus autem, quam aedificabat rex Salomon Domino, habebat sexaginta cubitos in longitudine et viginti cubitos in latitudine et triginta cubitos in altitudine.
1KGS|6|3|Et porticus erat ante templum viginti cubitorum longitudinis iuxta mensuram latitudinis templi et habebat decem cubitos latitudinis ante faciem templi.
1KGS|6|4|Fecitque in templo fenestras cum marginibus et cancellis.
1KGS|6|5|Et aedificavit contra parietem templi tabulata per gyrum in parietibus domus per circuitum templi et Dabir et fecit latera in circuitu.
1KGS|6|6|Tabulatum, quod subter erat, quinque cubitos habebat latitudinis et medium tabulatum sex cubitorum latitudinis et tertium tabulatum septem habens cubitos latitudinis; gradus enim posuit in domo per circuitum forinsecus, ut non ingrederentur trabes in muros templi.
1KGS|6|7|Domus autem cum aedificaretur, lapidibus dedolatis atque perfectis aedificata est; et malleus et securis et omne ferramentum non sunt audita in domo, cum aedificaretur.
1KGS|6|8|Ostium lateris inferioris in parte erat domus dextrae, et per cochleam ascendebant in medium latus et a medio in tertium.
1KGS|6|9|Et aedificavit domum et consummavit eam; texit quoque domum laquearibus cedrinis.
1KGS|6|10|Aedificavit ergo stratum contra omnem domum quinque cubitis altitudinis et iunxit domui lignis cedrinis.
1KGS|6|11|Et factus est sermo Domini ad Salomonem dicens:
1KGS|6|12|" Domus haec, quam aedificas, si ambulaveris in praeceptis meis et iudicia mea feceris et custodieris omnia mandata mea gradiens per ea, firmabo sermonem meum tibi, quem locutus sum ad David patrem tuum;
1KGS|6|13|et habitabo in medio filiorum Israel et non derelinquam populum meum Israel ".
1KGS|6|14|Igitur aedificavit Salomon domum et consummavit eam.
1KGS|6|15|Et aedificavit parietes domus intrinsecus tabulis cedrinis; a pavimento domus usque ad summitatem parietum et usque ad laquearia operuit lignis intrinsecus et texit pavimentum domus tabulis abiegnis.
1KGS|6|16|Aedificavitque viginti cubitorum a posteriore parte templi tabulis cedrinis a pavimento usque ad superiora; et fecit ei intrinsecus Dabir, id est sancta sanctorum.
1KGS|6|17|Porro quadraginta cubitorum erat ipsum templum ante illud.
1KGS|6|18|Et cedrus in domo intrinsecus sculptas habebat colocynthidas et calices apertos florum. Omnia cedrinis tabulis vestiebantur, nec omnino lapis apparere poterat in pariete.
1KGS|6|19|Dabir autem in medio domus in interiori parte fecerat, ut poneret ibi arcam foederis Domini.
1KGS|6|20|Habebat viginti cubitos longitudinis et viginti cubitos latitudinis et viginti cubitos altitudinis; et vestivit illud auro purissimo et fecit altare cedrinum ante Dabir.
1KGS|6|21|Domum quoque operuit Salomon intrinsecus auro purissimo et posuit catenas aureas ante Dabir.
1KGS|6|22|Nihilque erat in templo, quod non auro tegeretur; sed et totum altare Dabir texit auro.
1KGS|6|23|Et fecit in Dabir duos cherubim de lignis oleastri decem cubitorum altitudinis.
1KGS|6|24|Quinque cubitorum ala cherub una et quinque cubitorum ala cherub altera, id est decem cubitos habentes a summitate alae unius usque ad alae alterius summitatem.
1KGS|6|25|Decem quoque cubitorum erat cherub secundus, mensura par et effigies una erat duobus cherubim;
1KGS|6|26|altitudinem habebat unus cherub decem cubitorum et similiter cherub secundus.
1KGS|6|27|Posuitque cherubim in medio templi interioris; extendebant autem alas suas cherubim, et tangebat ala una parietem et ala cherub secundi tangebat parietem alterum; alae autem alterae in media parte templi se invicem contingebant.
1KGS|6|28|Texit quoque cherubim auro.
1KGS|6|29|Et omnes parietes templi per circuitum scalpsit variis caelaturis; et fecit in eis cherubim et palmas et calices apertos florum intrinsecus et foras.
1KGS|6|30|Sed et pavimentum domus texit auro intrinsecus et extrinsecus.
1KGS|6|31|Et pro ingressu Dabir fecit valvas de lignis oleastri postesque cum marginibus quinque.
1KGS|6|32|Et in duabus valvis de lignis oleastri scalpsit cherubim et palmas et calices apertos florum et vestivit ea auro operiens tam cherubim quam palmas et cetera auro.
1KGS|6|33|Fecitque eodem modo pro introitu templi postes cum quattuor marginibus de lignis oleastri
1KGS|6|34|et duas valvas de lignis abiegnis; et utraque valva duplex erat et versatilis.
1KGS|6|35|Et scalpsit cherubim et palmas et calices apertos florum operuitque omnia laminis aureis.
1KGS|6|36|Et aedificavit atrium interius tribus ordinibus lapidum politorum et uno ordine lignorum cedri.
1KGS|6|37|Anno quarto fundata est domus Domini in mense Ziv;
1KGS|6|38|et in anno undecimo, mense Bul - ipse est mensis octavus - perfecta est domus in omni opere suo et in universis utensilibus; aedificavitque eam annis septem.
1KGS|7|1|Domum autem suam aedificavit Salomon tredecim annis et ad perfectum usque perduxit.
1KGS|7|2|Aedificavit quoque domum Saltus Libani centum cubitorum longitudinis et quinquaginta cubitorum latitudinis et triginta cubitorum altitudinis super quattuor ordines columnarum cedrinarum, et ligna cedrina super columnas.
1KGS|7|3|Et erat tectum cedrinum in alto super tabulas quadraginta quinque, quae erant super columnas, quindecim in uno ordine,
1KGS|7|4|et marginum tres ordines, fenestra iuxta fenestram tribus vicibus.
1KGS|7|5|Ostia, id est postes, habebant quadruplicem marginem.
1KGS|7|6|Et porticum columnarum fecit quinquaginta cubitorum longitudinis et triginta cubitorum latitudinis, et alteram porticum in facie maioris porticus et columnas et cancellos ante eas.
1KGS|7|7|Porticum quoque solii, in qua tribunal erat, fecit et texit lignis cedrinis a pavimento usque ad pavimentum.
1KGS|7|8|Et domus, in qua habitabat, erat in altero atrio intro a porticu et simili opere. Domum quoque fecit filiae pharaonis, quam uxorem duxerat Salomon, tali opere quali et hanc porticum.
1KGS|7|9|Omnia lapidibus pretiosis, qui ad normam quandam atque mensuram tam intrinsecus quam extrinsecus serrati erant, a fundamento usque ad summitatem parietum, et extrinsecus usque ad atrium maius.
1KGS|7|10|Fundamenta autem de lapidibus pretiosis, lapidibus magnis decem sive octo cubitorum.
1KGS|7|11|Et desuper lapides pretiosi secundum mensuram secti et ligna cedrina.
1KGS|7|12|Et atrium maius in circuitu habebat tres ordines de lapidibus sectis et unum ordinem de dolata cedro; necnon et atrium domus Domini interius et porticus domus.
1KGS|7|13|Misit quoque rex Salomon et tulit Hiram de Tyro,
1KGS|7|14|filium mulieris viduae de tribu Nephthali, patre Tyrio, artificem aerarium et plenum sapientia et intellegentia et doctrina ad faciendum omne opus ex aere. Qui, cum venisset ad regem Salomonem, fecit omne opus eius.
1KGS|7|15|Et finxit duas columnas aereas, decem et octo cubitorum altitudinis columnam unam, et linea duodecim cubitorum ambiebat columnam, et grossitudo eius quattuor digitorum, et intrinsecus cava erat; sic et columna altera.
1KGS|7|16|Duo quoque capitella fecit, quae ponerentur super capita columnarum, fusili aere; quinque cubitorum altitudinis capitellum unum et quinque cubitorum altitudinis capitellum alterum,
1KGS|7|17|et serta quasi in modum texturae, fimbriae in modum catenarum sibi invicem miro opere contextarum in capitellis, quae erant super caput columnarum, septem in capitello uno et septem in capitello altero.
1KGS|7|18|Et fecit malogranatorum duos ordines per circuitum super sertum unum, ut tegerent capitella, quae erant super summitatem columnarum; eodem modo fecit et capitello secundo.
1KGS|7|19|Capitella autem, quae erant super capita columnarum, quasi opere lilii fabricata erant in porticu, quattuor cubitorum.
1KGS|7|20|Et rursum alia capitella in summitate duarum columnarum etiam desuper, iuxta alvum, quae erat super sertum. Malogranatorum autem ducentorum duo ordines erant in circuitu capitelli primi et eodem modo in circuitu capitelli secundi.
1KGS|7|21|Et statuit duas columnas in porticum templi; cumque statuisset columnam dexteram, vocavit eam nomine Iachin, similiter erexit columnam sinistram et vocavit nomen eius Booz.
1KGS|7|22|Et super capita columnarum opus in modum lilii posuit; per fectumque est opus columnarum.
1KGS|7|23|Fecit quoque mare fusile decem cubitorum a labio usque ad labium, rotundum in circuitu, quinque cubitorum altitudo eius; et resticula triginta cubitorum cingebat illud per circuitum.
1KGS|7|24|Et scalptura colocynthidum subter labium circuibat illud, duo ordines scalpturarum fusilium in una fusione cum mari.
1KGS|7|25|Et stabat super duodecim boves, e quibus tres respiciebant ad aquilonem et tres ad occidentem et tres ad meridiem et tres ad orientem, et mare super eos desuper erat; quorum posteriora universa intrinsecus latitabant.
1KGS|7|26|Grossitudo autem luteris habebat mensuram palmi, labiumque eius erat quasi labium calicis et folium repandi lilii; duo milia batos capiebat.
1KGS|7|27|Et fecit bases decem aereas, quattuor cubitorum longitudinis bases singulas et quattuor cubitorum latitudinis et trium cubitorum altitudinis.
1KGS|7|28|Hoc autem erat opus basium: limbos habebant, insuper et limbos inter columellas.
1KGS|7|29|Super limbos inter columellas erant leones et boves et cherubim, et super columellas similiter; supra et infra leones et boves erant coronae, opus malleatum.
1KGS|7|30|Et quattuor rotae per bases singulas et axes aerei, et quattuor pedes et quasi umeruli subter luterem fusiles, contra singulos coronae.
1KGS|7|31|Et os eius erat rotundum, opus basis, unius cubiti et dimidii; etiam in ore eius variae caelaturae erant, limbi autem eius erant quadrati, non rotundi.
1KGS|7|32|Quattuor quoque rotae subter limbis erant, et fulcra rotarum cohaerebant basi; una rota habebat altitudinis cubitum et semis.
1KGS|7|33|Tales autem rotae erant, quales solent in curru fieri, et fulcra earum et canthi et radii et modioli, omnia fusilia.
1KGS|7|34|Nam et umeruli illi quattuor per singulos angulos basis unius ex ipsa basi fusiles et coniuncti erant.
1KGS|7|35|In summitate autem basis erat quaedam rotunditas dimidii cubiti, et in summitate basis fulcra eius et limbi eius ex semetipsa.
1KGS|7|36|Scalpsit quoque in tabulatis illis, fulcris eius et super limbos eius cherubim et leones et palmas secundum vacuum singulorum, et coronas per circuitum.
1KGS|7|37|In hunc modum fecit decem bases, fusura una, et mensura scalpturaque consimili.
1KGS|7|38|Fecit quoque decem luteres aereos; quadraginta batos capiebat luter unus, eratque quattuor cubitorum; singulosque luteres per singulas, id est decem bases posuit.
1KGS|7|39|Et constituit decem bases, quinque ad dexteram partem templi et quinque ad sinistram; mare autem posuit ad dexteram partem templi contra orientem ad meridiem.
1KGS|7|40|Fecit quoque Hiram lebetes et vatilla et phialas et perfecit omne opus regi Salomoni in templo Domini;
1KGS|7|41|columnas duas et globos capitellorum super capita columnarum duos et serta duo, ut operirent duos globos, qui erant super capita columnarum;
1KGS|7|42|et malogranata quadringenta in duobus sertis, duos versus malogranatorum in sertis singulis, ad operiendos globos capitellorum, qui erant super faciem columnarum;
1KGS|7|43|et bases decem et luteres decem super bases
1KGS|7|44|et mare unum et boves duodecim subter mare;
1KGS|7|45|et lebetes et vatilla et phialas. Omnia vasa, quae fecit Hiram regi Salomoni in domo Domini, de aere polito erant.
1KGS|7|46|In campestri regione Iordanis fudit ea rex in argillosa terra inter Succoth et Sarthan.
1KGS|7|47|Et posuit Salomon omnia vasa; propter multitudinem autem nimiam ignorabatur pondus aeris.
1KGS|7|48|Fecitque Salomon omnia vasa in domo Domini: altare aureum et mensam, super quam ponerentur panes propositionis, auream;
1KGS|7|49|et candelabra, quinque ad dexteram et quinque ad sinistram contra Dabir, ex auro puro, et florem et lucernas desuper aureas; et forcipes aureos
1KGS|7|50|et pateras et cultros et phialas et sartagines et turibula de auro purissimo; et cardines ostiorum domus interioris Sancti sanctorum et ostiorum domus templi ex auro.
1KGS|7|51|Et perfecit omne opus, quod faciebat Salomon in domo Domini, et intulit Salomon, quae sanctificaverat David pater suus, argentum et aurum et vasa, reposuitque in thesauris domus Domini.
1KGS|8|1|Tunc congregavit Salomon om nes maiores natu Israel - om nes principes tribuum, duces familiarum filiorum Israel ad regem Salomonem - in Ierusalem, ut deferrent arcam foederis Domini de civitate David, id est de Sion.
1KGS|8|2|Convenitque ad regem Salomonem universus Israel in mense Ethanim in sollemnitate, ipse est mensis septimus.
1KGS|8|3|Veneruntque cuncti senes Israel, et tulerunt sacerdotes arcam
1KGS|8|4|et portaverunt arcam Domini et tabernaculum conventus et omnia vasa sanctuarii, quae erant in tabernaculo; et ferebant ea sacerdotes et Levitae.
1KGS|8|5|Rex autem Salomon et universus coetus Israel, qui convenerat ad eum, cum illo ante arcam immolabant oves et boves absque aestimatione et numero.
1KGS|8|6|Et intulerunt sacerdotes arcam foederis Domini in locum suum in Dabir templi, in sanctum sanctorum, subter alas cherubim;
1KGS|8|7|siquidem cherubim expandebant alas super locum arcae et protegebant arcam et vectes eius desuper.
1KGS|8|8|Cumque eminerent vectes et apparerent summitates eorum foris in sanctuario ante Dabir, non apparebant ultra extrinsecus; qui et fuerunt ibi usque in praesentem diem.
1KGS|8|9|In arca autem non erat aliud nisi duae tabulae lapideae, quas posuerat in ea Moyses in Horeb, quando pepigit Dominus foedus cum filiis Israel, cum egrederentur de terra Aegypti.
1KGS|8|10|Factum est autem cum exissent sacerdotes de sanctuario, nebula implevit domum Domini,
1KGS|8|11|et non poterant sacerdotes stare et ministrare propter nebulam; impleverat enim gloria Domini domum Domini.
1KGS|8|12|Tunc ait Salomon: Dominus dixit ut habitaret in nebula.
1KGS|8|13|Aedificans aedificavi domum in habitaculum tuum,firmissimum solium tuum in sempiternum ".
1KGS|8|14|Convertitque rex faciem suam et benedixit omni ecclesiae Israel; omnis enim ecclesia Israel stabat.
1KGS|8|15|Et ait: " Benedictus Dominus, Deus Israel, qui locutus est ore suo ad David patrem meum et in manibus suis perfecit dicens:
1KGS|8|16|"A die qua eduxi populum meum Israel de Aegypto, non elegi civitatem de universis tribubus Israel, ut aedificaretur domus, et esset nomen meum ibi; sed elegi David, ut esset super populum meum Israel".
1KGS|8|17|Voluitque David pater meus aedificare domum nomini Domini, Dei Israel,
1KGS|8|18|et ait Dominus ad David patrem meum: "Quod cogitasti in corde tuo aedificare domum nomini meo, bene fecisti hoc ipsum mente tractans;
1KGS|8|19|verumtamen tu non aedificabis domum sed filius tuus, qui egredietur de lumbis tuis, ipse aedificabit domum nomini meo".
1KGS|8|20|Confirmavit Dominus sermonem suum, quem locutus est; stetique pro David patre meo et sedi super thronum Israel, sicut locutus est Dominus, et aedificavi domum nomini Domini, Dei Israel.
1KGS|8|21|Et constitui ibi locum arcae, in qua foedus est Domini, quod percussit cum patribus nostris, quando eduxit eos de terra Aegypti ".
1KGS|8|22|Stetit autem Salomon ante altare Domini in conspectu omnis ecclesiae Israel et expandit manus suas in caelum
1KGS|8|23|et ait: " Domine, Deus Israel, non est similis tui Deus in caelo desuper et super terra deorsum, qui custodis pactum et misericordiam servis tuis, qui ambulant coram te in toto corde suo;
1KGS|8|24|qui custodisti servo tuo David patri meo, quae locutus es ei; ore locutus es et manibus perfecisti, ut et haec dies probat.
1KGS|8|25|Nunc igitur, Domine, Deus Israel, conserva famulo tuo David patri meo, quae locutus es ei dicens: "Non auferetur de te vir coram me, qui sedeat super thronum Israel, ita tamen, si custodierint filii tui viam suam, ut ambulent coram me, sicut tu ambulasti in conspectu meo".
1KGS|8|26|Et nunc, Domine, Deus Israel, firmentur verba tua, quae locutus es servo tuo David patri meo.
1KGS|8|27|Ergone putandum est quod vere Deus habitet super terram? Si enim caelum et caeli caelorum te capere non possunt, quanto magis domus haec, quam aedificavi!
1KGS|8|28|Sed respice ad orationem servi tui et ad preces eius, Domine Deus meus; audi clamorem et orationem, quam servus tuus orat coram te hodie,
1KGS|8|29|ut sint oculi tui aperti super domum hanc nocte ac die, super locum, de quo dixisti: "Erit nomen meum ibi", ut exaudias orationem, qua orat te servus tuus in loco isto,
1KGS|8|30|ut exaudias deprecationem servi tui et populi tui Israel, quodcumque oraverint in loco isto, et exaudies in loco habitaculi tui in caelo et, cum exaudieris, propitius eris.
1KGS|8|31|Si peccaverit homo in proximum suum et habuerit aliquod iuramentum, quo teneatur astrictus, et venerit propter iuramentum coram altari tuo in domum istam,
1KGS|8|32|tu exaudies in caelo et facies et iudicabis servos tuos condemnans impium et reddens viam suam super caput eius iustificansque iustum et retribuens ei secundum iustitiam suam.
1KGS|8|33|Si superatus fuerit populus tuus Israel ab inimicis suis, quia peccaturus est tibi, et agentes paenitentiam et confitentes nomini tuo venerint et oraverint et deprecati te fuerint in domo hac,
1KGS|8|34|exaudi in caelo et dimitte peccatum populi tui Israel et reduces eos in terram, quam dedisti patribus eorum.
1KGS|8|35|Si clausum fuerit caelum et non pluerit propter peccata eorum, et oraverint in loco isto confessi nomini tuo et a peccatis suis conversi propter afflictionem suam,
1KGS|8|36|exaudi eos in caelo et dimitte peccata servorum tuorum et populi tui Israel et ostende eis viam bonam, per quam ambulent, et da pluviam super terram tuam, quam dedisti populo tuo in possessionem.
1KGS|8|37|Fames si oborta fuerit in terra aut pestilentia aut uredo aut aurugo aut locusta vel bruchus, et afflixerit eum inimicus eius portas obsidens, omnis plaga, universa infirmitas,
1KGS|8|38|cuncta oratio et deprecatio, quae acciderit omni homini de populo tuo Israel; si quis cognoverit plagam cordis sui et expanderit manus suas in domo hac,
1KGS|8|39|tu audies in caelo in loco habitationis tuae et repropitiaberis et facies, ut des unicuique secundum omnes vias suas, sicut videris cor eius, quia tu nosti solus cor omnium filiorum hominum,
1KGS|8|40|ut timeant te cunctis diebus, quibus vivunt super faciem terrae, quam dedisti patribus nostris.
1KGS|8|41|Insuper et alienigena, qui non est de populo tuo Israel, cum venerit de terra longinqua propter nomen tuum
1KGS|8|42|- audietur enim nomen tuum magnum et manus tua fortis et brachium tuum extentum ubique - cum venerit ergo et oraverit in hoc loco,
1KGS|8|43|tu exaudies in caelo in loco habitationis tuae et facies omnia, pro quibus invocaverit te alienigena, ut sciant universi populi terrarum nomen tuum et timeant te, sicut populus tuus Israel, et probent quia nomen tuum invocatum est super domum hanc, quam aedificavi.
1KGS|8|44|Si egressus fuerit populus tuus ad bellum contra inimicos suos per viam, quocumque miseris eos, et oraverint te contra viam civitatis, quam elegisti, et contra domum, quam aedificavi nomini tuo,
1KGS|8|45|exaudies in caelo orationes eorum et preces eorum et facies iudicium eorum.
1KGS|8|46|Quod si peccaverint tibi - non est enim homo qui non peccet - et iratus tradideris eos inimicis suis, et captivi ducti fuerint in terram inimicorum longe vel prope
1KGS|8|47|et egerint paenitentiam in corde suo in loco captivitatis et conversi deprecati te fuerint in captivitate sua dicentes: "Peccavimus, inique egimus, impie gessimus";
1KGS|8|48|et reversi fuerint ad te in universo corde suo et tota anima sua in terra inimicorum suorum, ad quam captivi ducti sunt, et oraverint te contra viam terrae suae, quam dedisti patribus eorum, et civitatis, quam elegisti, et templi, quod aedificavi nomini tuo,
1KGS|8|49|exaudies in caelo in firmamento solii tui orationes eorum et preces eorum et facies iudicium eorum;
1KGS|8|50|et propitiaberis populo tuo, qui peccavit tibi, et omnibus iniquitatibus eorum, quibus praevaricati sunt in te, et dabis misericordiam coram eis, qui eos captivos habuerint, ut misereantur eis
1KGS|8|51|- populus enim tuus est et hereditas tua, quos eduxisti de terra Aegypti de medio fornacis ferreae -
1KGS|8|52|ut sint oculi tui aperti ad deprecationem servi tui et populi tui Israel, et exaudias eos in universis, pro quibus invocaverint te.
1KGS|8|53|Tu enim separasti eos tibi in hereditatem de universis populis terrae, sicut locutus es per Moysen servum tuum, quando eduxisti patres nostros de Aegypto, Domine Deus ".
1KGS|8|54|Factum est autem cum complesset Salomon orans Dominum omnem orationem et deprecationem hanc, surrexit de conspectu altaris Domini; utrumque enim genu in terram fixerat et manus expanderat in caelum.
1KGS|8|55|Stetit ergo et benedixit omni ecclesiae Israel voce magna dicens:
1KGS|8|56|" Benedictus Dominus, qui dedit requiem populo suo Israel iuxta omnia, quae locutus est; non cecidit ne unus quidem sermo ex omnibus bonis, quae locutus est per Moysen servum suum.
1KGS|8|57|Sit Dominus Deus noster nobiscum, sicut fuit cum patribus nostris, non derelinquens nos neque proiciens,
1KGS|8|58|sed inclinet corda nostra ad se, ut ambulemus in universis viis eius et custodiamus mandata eius et decreta et iudicia, quaecumque mandavit patribus nostris.
1KGS|8|59|Et sint sermones mei isti, quibus deprecatus sum coram Domino, appropinquantes Domino Deo nostro die ac nocte, ut faciat iudicium servo suo et populo suo Israel per singulos dies,
1KGS|8|60|ut sciant omnes populi terrae quia Dominus ipse est Deus, et non est ultra absque eo.
1KGS|8|61|Sit quoque cor vestrum perfectum cum Domino Deo nostro, ut ambuletis in decretis eius et custodiatis mandata eius sicut et hodie ".
1KGS|8|62|Igitur rex et omnis Israel cum eo immolabant victimas coram Domino.
1KGS|8|63|Mactavitque Salomon hostias pacificas, quas immolavit Domino, boum viginti duo milia et ovium centum viginti milia. Et dedicaverunt templum Domini rex et omnes filii Israel.
1KGS|8|64|In die illa sanctificavit rex medium atrii, quod erat ante domum Domini; fecit quippe holocaustum ibi et oblationem et adipem pacificorum, quoniam altare aereum, quod erat coram Domino, minus erat et capere non poterat holocaustum et oblationem et adipem pacificorum.
1KGS|8|65|Fecit ergo Salomon in tempore illo festivitatem celebrem, et omnis Israel cum eo, ecclesia magna ab introitu Emath usque ad rivum Aegypti, coram Domino Deo nostro septem diebus.
1KGS|8|66|Et in die octava dimisit populos; qui benedicentes regi profecti sunt in tabernacula sua laetantes et alacri corde super omnibus bonis, quae fecerat Dominus David servo suo et Israel populo suo.
1KGS|9|1|Factum est autem cum perfecisset Salomon aedificium domus Domini et aedificium regis et omne, quod optaverat et voluerat facere,
1KGS|9|2|apparuit ei Dominus secundo, sicut apparuerat ei in Gabaon.
1KGS|9|3|Dixitque Dominus ad eum: " Exaudivi orationem tuam et deprecationem tuam, quam deprecatus es coram me; sanctificavi domum hanc, quam aedificasti, ut ponerem nomen meum ibi in sempiternum; et erunt oculi mei et cor meum ibi cunctis diebus.
1KGS|9|4|Tu quoque, si ambulaveris coram me, sicut ambulavit David pater tuus in simplicitate cordis et in aequitate, et feceris omnia, quae praecepi tibi, et legitima mea et iudicia mea servaveris,
1KGS|9|5|ponam thronum regni tui super Israel in sempiternum, sicut locutus sum David patri tuo dicens: Non auferetur de genere tuo vir de solio Israel.
1KGS|9|6|Si autem aversione aversi fueritis vos et filii vestri non sequentes me nec custodientes mandata mea et decreta mea, quae proposui vobis, sed abieritis et colueritis deos alienos et adoraveritis eos,
1KGS|9|7|auferam Israel de superficie terrae, quam dedi eis, et templum, quod sanctificavi nomini meo, proiciam a conspectu meo; eritque Israel in proverbium et in fabulam cunctis populis,
1KGS|9|8|et domus haec erit in ruinas. Omnis, qui transierit per eam, stupebit et sibilabit et dicet: "Quare fecit Dominus sic terrae huic et domui huic?".
1KGS|9|9|Et respondebunt: "Quia dereliquerunt Dominum Deum suum, qui eduxit patres eorum de terra Aegypti, et secuti sunt deos alienos et adoraverunt eos et coluerunt eos; idcirco induxit Dominus super eos omne malum hoc" ".
1KGS|9|10|Expletis autem annis viginti, postquam aedificaverat Salomon duas domos, id est domum Domini et domum regis
1KGS|9|11|- Hiram rege Tyri praebente Salomoni ligna cedrina et abiegna et aurum iuxta omne quod opus habuerat - tunc dedit Salomon Hiram viginti oppida in terra Galilaeae.
1KGS|9|12|Et egressus est Hiram de Tyro, ut videret oppida, quae dederat ei Salomon, et non placuerunt ei;
1KGS|9|13|et ait: " Haeccine sunt civitates, quas dedisti mihi, frater? ". Et appellavit eas terram Chabul usque in diem hanc.
1KGS|9|14|Misit quoque Hiram ad regem centum viginti talenta auri.
1KGS|9|15|Haec est summa indictionis, quam constituit rex Salomon ad aedificandam domum Domini et domum suam et Mello et murum Ierusalem et Asor et Mageddo et Gazer.
1KGS|9|16|Pharao rex Aegypti ascendit et cepit Gazer succenditque eam igni et Chananaeum, qui habitabat in civitate, interfecit; et dedit eam in dotem filiae suae uxori Salomonis.
1KGS|9|17|Aedificavit ergo Salomon Gazer et Bethoron inferiorem
1KGS|9|18|et Baalath et Thamar in terra solitudinis
1KGS|9|19|et omnes civitates horreorum, quae ad se pertinebant, et civitates curruum et civitates equorum et quodcumque ei placuit, ut aedificaret in Ierusalem et in Libano et in omni terra potestatis suae.
1KGS|9|20|Universum populum, qui remanserat de Amorraeis et Hetthaeis et Pherezaeis et Hevaeis et Iebusaeis, qui non erant de filiis Israel,
1KGS|9|21|horum filios, qui remanserant post eos in terra, quos scilicet non potuerant filii Israel exterminare, fecit Salomon tributarios usque in diem hanc.
1KGS|9|22|De filiis autem Israel non constituit Salomon servire quemquam, sed erant viri bellatores et ministri eius et principes et pugnatores eius et praefecti curruum et equitum.
1KGS|9|23|Erant autem principes eorum, qui super omnia opera Salomonis praepositi erant, quingenti quinquaginta; qui habebant subiectum populum et statutis operibus imperabant.
1KGS|9|24|Filia autem pharaonis ascendit de civitate David in domum suam, quam aedificaverat ei; tunc aedificavit Mello.
1KGS|9|25|Offerebat quoque Salomon tribus vicibus per annos singulos holocausta et pacificas victimas super altare, quod aedificaverat Domino, et adolebat coram Domino; perfectumque est templum.
1KGS|9|26|Classem quoque fecit rex Salomon in Asiongaber, quae est iuxta Ailath in litore maris Rubri in terra Idumaea.
1KGS|9|27|Misitque Hiram in classe illa servos suos viros nauticos gnaros maris cum servis Salomonis.
1KGS|9|28|Qui, cum venissent in Ophir, sumptum inde aurum quadringentorum viginti talentorum detulerunt ad regem Salomonem.
1KGS|10|1|Sed et regina Saba, audita fama Salomonis - in hono rem nominis Domini - venit tentare eum in aenigmatibus.
1KGS|10|2|Et ingressa Ierusalem multo cum comitatu et divitiis, camelis portantibus aromata et aurum infinitum nimis et gemmas pretiosas, venit ad Salomonem et locuta est ei universa, quae habebat in corde suo.
1KGS|10|3|Et docuit eam Salomon omnia verba, quae proposuerat: non fuit sermo, qui regem posset latere, et non responderet ei.
1KGS|10|4|Videns autem regina Saba omnem sapientiam Salomonis et domum, quam aedificaverat,
1KGS|10|5|et cibos mensae eius et sessionem servorum et ordinem ministrantium vestesque eorum et pincernas et holocausta, quae offerebat in domo Domini, non habebat ultra spiritum
1KGS|10|6|dixitque ad regem: " Verus est sermo, quem audivi in terra mea super rebus tuis et super sapientia tua!
1KGS|10|7|Et non credebam narrantibus mihi, donec ipsa veni et vidi oculis meis et probavi quod media pars mihi nuntiata non fuerit; maior est sapientia et bona tua quam rumor, quem audivi.
1KGS|10|8|Beati viri tui et beati servi tui hi, qui stant coram te semper et audiunt sapientiam tuam!
1KGS|10|9|Sit Dominus Deus tuus benedictus, cui placuisti, et posuit te super thronum Israel, eo quod dilexerit Dominus Israel in sempiternum et constituit te regem, ut faceres iudicium et iustitiam ".
1KGS|10|10|Dedit ergo regi centum viginti talenta auri et aromata multa nimis et gemmas pretiosas; non sunt allata ultra aromata tam multa quam ea, quae dedit regina Saba regi Salomoni.
1KGS|10|11|Sed et classis Hiram, quae portabat aurum de Ophir, attulit ex Ophir ligna thyina multa nimis et gemmas pretiosas.
1KGS|10|12|Fecitque rex de lignis thyinis fulcra domus Domini et domus regiae et citharas lyrasque cantoribus. Non sunt allata huiuscemodi ligna thyina neque visa usque in praesentem diem.
1KGS|10|13|Rex autem Salomon dedit reginae Saba omnia, quae voluit et petivit ab eo, praeter ea, quae ultro obtulerat ei munere regio. Quae reversa est et abiit in terram suam cum servis suis.
1KGS|10|14|Erat autem pondus auri, quod afferebatur Salomoni per annos singulos, sescentorum sexaginta sex talentorum auri,
1KGS|10|15|praeter id, quod proveniebat ex tributis subiectorum et commercio negotiatorum et omnium regum Arabiae et ducum terrae.
1KGS|10|16|Fecit quoque rex Salomon ducenta scuta de auro puro, sescentos auri siclos dedit in laminas scuti unius;
1KGS|10|17|et trecentas peltas ex auro probato, tres minae auri unam peltam vestiebant; posuitque ea rex in domo Saltus Libani.
1KGS|10|18|Fecit etiam rex Salomon thronum de ebore grandem et vestivit eum auro fulvo nimis.
1KGS|10|19|Qui habebat sex gradus, et summitas throni rotunda erat in parte posteriori, et duae manus hinc atque inde tenentes sedile, et duo leones stabant iuxta manus;
1KGS|10|20|et duodecim leunculi stantes super sex gradus hinc atque inde. Non est factum tale opus in universis regnis.
1KGS|10|21|Sed et omnia vasa, quibus potabat rex Salomon, erant aurea, et universa supellex domus Saltus Libani de auro purissimo; non erat argentum nec alicuius pretii putabatur in diebus Salomonis,
1KGS|10|22|quia classis Tharsis, quae regi erat, per mare cum classe Hiram semel per tres annos redibat deferens aurum et argentum et ebur et simias et pavos.
1KGS|10|23|Magnificatus est ergo rex Salomon super omnes reges terrae divitiis et sapientia.
1KGS|10|24|Et universa terra desiderabat vultum Salomonis, ut audiret sapientiam eius, quam dederat Deus in corde eius.
1KGS|10|25|Et singuli deferebant ei munera, vasa argentea et aurea, vestes et arma bellica, aromata quoque et equos et mulos per annos singulos.
1KGS|10|26|Congregavitque Salomon currus et equites, et facti sunt ei mille quadringenti currus et duodecim milia equitum; et disposuit eos per civitates quadrigarum et cum rege in Ierusalem.
1KGS|10|27|Fecitque ut tanta esset abundantia argenti in Ierusalem quanta et lapidum; et cedrorum praebuit multitudinem quasi sycomoros, quae nascuntur in Sephela.
1KGS|10|28|Et educebantur equi Salomoni de Aegypto et de Coa; negotiatores enim regis emebant de Coa statuto pretio.
1KGS|10|29|Constabat autem et egrediebatur quadriga ex Aegypto sescentis siclis argenti, et equus centum quinquaginta; atque in hunc modum cunctis regibus Hetthaeorum et Syriae per manus suas venundabant.
1KGS|11|1|Rex autem Salomon amavit mulieres alienigenas multas, filiam quoque pharaonis et Moabitidas et Ammonitidas, Idumaeas et Sidonias et Hetthaeas,
1KGS|11|2|de gentibus, super quibus dixit Dominus filiis Israel: " Non ingrediemini ad eas, neque de illis ingredientur ad vestras; certissime enim avertent corda vestra, ut sequamini deos earum ". His itaque copulatus est Salomon amore;
1KGS|11|3|fueruntque ei uxores quasi reginae septingentae et concubinae trecentae, et averterunt mulieres cor eius.
1KGS|11|4|Cumque iam esset senex, depravatum est cor eius per mulieres, ut sequeretur deos alienos; nec erat cor eius perfectum cum Domino Deo suo sicut cor David patris eius,
1KGS|11|5|sed colebat Salomon Astharthen, deam Sidoniorum, et Melchom idolum Ammonitarum.
1KGS|11|6|Fecitque Salomon quod non placuerat coram Domino et non adimplevit ut sequeretur Dominum sicut David pater eius.
1KGS|11|7|Tunc aedificavit Salomon fanum Chamos idolo Moab in monte, qui est contra Ierusalem, et Melchom idolo filiorum Ammon;
1KGS|11|8|atque in hunc modum fecit universis uxoribus suis alienigenis, quae adolebant et immolabant diis suis.
1KGS|11|9|Igitur iratus est Dominus Salomoni, quod aversa esset mens eius a Domino, Deo Israel, qui apparuerat ei bis
1KGS|11|10|et praeceperat de verbo hoc, ne sequeretur deos alienos; et non custodivit, quae mandavit ei Dominus.
1KGS|11|11|Dixit itaque Dominus Salomoni: " Quia habuisti hoc apud te et non custodisti pactum meum et praecepta mea, quae mandavi tibi, disrumpens scindam regnum tuum a te et dabo illud servo tuo.
1KGS|11|12|Verumtamen in diebus tuis non faciam propter David patrem tuum; de manu filii tui scindam illud.
1KGS|11|13|Nec totum regnum auferam, sed tribum unam dabo filio tuo propter David servum meum et Ierusalem, quam elegi ".
1KGS|11|14|Suscitavit autem Dominus adversarium Salomoni Adad Idumaeum, qui erat de semine regio, in Edom.
1KGS|11|15|Cum enim vicisset David Idumaeam, et ascendisset Ioab princeps militiae ad sepeliendum eos, qui fuerant interfecti, et occidisset omne masculinum in Idumaea
1KGS|11|16|- sex enim mensibus ibi moratus est Ioab et omnis Israel, donec interimerent omne masculinum in Idumaea -
1KGS|11|17|fugit Adad ipse et viri Idumaei de servis patris eius cum eo, ut ingrederetur Aegyptum; erat autem Adad puer parvulus.
1KGS|11|18|Cumque surrexissent de Madian, venerunt in Pharan tuleruntque secum viros de Pharan et introierunt Aegyptum ad pharaonem regem Aegypti, qui dedit ei domum et cibos constituit et terram delegavit.
1KGS|11|19|Et invenit Adad gratiam coram pharao valde, in tantum ut daret ei uxorem sororem uxoris suae germanam Taphnes reginae.
1KGS|11|20|Genuitque ei soror Taphnes Genubath filium et ablactavit eum Taphnes in domo pharaonis, eratque Genubath habitans apud pharaonem cum filiis eius.
1KGS|11|21|Cumque audisset Adad in Aegypto dormisse David cum patribus suis et mortuum esse Ioab principem militiae, dixit pharaoni: " Dimitte me, ut vadam in terram meam ".
1KGS|11|22|Dixitque ei pharao: " Qua enim re apud me indiges, ut quaeras ire ad terram tuam? ". At ille respondit: " Nulla; sed obsecro, ut dimittas me ".
1KGS|11|23|Suscitavit quoque Deus Salomoni adversarium Razon filium Eliada, qui fugerat ab Adadezer rege Soba domino suo.
1KGS|11|24|Et congregavit ad se viros et factus est princeps turmae, cum interficeret eos David; abieruntque Damascum et habitaverunt ibi et regnaverunt in Damasco.
1KGS|11|25|Eratque adversarius Israeli cunctis diebus Salomonis; et hoc cum malo, quod erat Adad. Et detestatus est Israel regnavitque in Syria.
1KGS|11|26|Ieroboam quoque filius Nabat, Ephrathaeus de Sareda, servus Salomonis, cuius mater erat nomine Sarva mulier vidua, levavit manum contra regem.
1KGS|11|27|Et haec causa rebellionis adversus eum: Salomon aedificavit Mello et coaequavit voraginem civitatis David patris sui.
1KGS|11|28|Erat autem Ieroboam vir fortis et strenuus; vidensque Salomon adulescentem industrium constituerat eum praefectum super labores universae domus Ioseph.
1KGS|11|29|Factum est igitur in tempore illo, ut Ieroboam egrederetur de Ierusalem, et inveniret eum Ahias Silonites propheta in via opertus pallio novo; erant autem duo tantum in agro.
1KGS|11|30|Apprehendensque Ahias pallium suum novum, quo coopertus erat, scidit in duodecim partes
1KGS|11|31|et ait ad Ieroboam: " Tolle tibi decem scissuras; haec enim dicit Dominus, Deus Israel: Ecce ego scindam regnum de manu Salomonis et dabo tibi decem tribus.
1KGS|11|32|Porro una tribus remanebit ei propter servum meum David et Ierusalem civitatem, quam elegi ex omnibus tribubus Israel;
1KGS|11|33|eo quod dereliquerint me et adoraverint Astharthen deam Sidoniorum et Chamos deum Moab et Melchom deum filiorum Ammon et non ambulaverint in viis meis, ut facerent iustitiam coram me et praecepta mea et iudicia sicut David pater eius.
1KGS|11|34|Nec auferam omne regnum de manu eius, sed ducem ponam eum cunctis diebus vitae suae propter David servum meum, quem elegi, qui custodivit mandata mea et praecepta mea.
1KGS|11|35|Auferam autem regnum de manu filii eius et dabo tibi decem tribus;
1KGS|11|36|filio autem eius dabo tribum unam, ut remaneat lucerna David servo meo cunctis diebus coram me in Ierusalem civitate, quam elegi, ut esset nomen meum ibi.
1KGS|11|37|Te autem assumam, et regnabis super omnia, quae desiderat anima tua, erisque rex super Israel.
1KGS|11|38|Si igitur audieris omnia, quae praecepero tibi, et ambulaveris in viis meis et feceris, quod rectum est coram me custodiens mandata mea et praecepta mea, sicut fecit David servus meus, ero tecum et aedificabo tibi domum stabilem, quomodo aedificavi David, et tradam tibi Israel
1KGS|11|39|et affligam semen David super hoc, verumtamen non cunctis diebus ".
1KGS|11|40|Voluit ergo Salomon interficere Ieroboam, qui surrexit et aufugit in Aegyptum ad Sesac regem Aegypti et fuit in Aegypto usque ad mortem Salomonis.
1KGS|11|41|Reliqua autem gestorum Salomonis, omnia, quae fecit, et sapientia eius, ecce universa scripta sunt in libro gestorum Salomonis;
1KGS|11|42|dies autem, quos regnavit Salomon in Ierusalem super omnem Israel, quadraginta anni sunt.
1KGS|11|43|Dormivitque Salomon cum patribus suis et sepultus est in civitate David patris sui; regnavitque Roboam filius eius pro eo.
1KGS|12|1|Venit autem Roboam in Sichem; illuc enim congregatus erat omnis Israel ad constituendum eum regem.
1KGS|12|2|At Ieroboam filius Nabat, cum adhuc esset in Aegypto profugus a facie regis Salomonis, audito hoc nuntio, reversus est de Aegypto.
1KGS|12|3|Miseruntque et vocaverunt eum. Venit ergo Ieroboam et omnis multitudo Israel, et locuti sunt ad Roboam dicentes:
1KGS|12|4|" Pater tuus durissimum iugum imposuit nobis; tu itaque nunc imminue paululum de imperio patris tui durissimo et de iugo gravissimo, quod imposuit nobis, et serviemus tibi ".
1KGS|12|5|Qui ait eis: " Ite usque ad tertium diem et revertimini ad me ".Cumque abisset populus,
1KGS|12|6|iniit consilium rex Roboam cum senioribus, qui assistebant coram Salomone patre eius, cum adhuc viveret, et ait: " Quod mihi datis consilium, ut respondeam populo huic? ".
1KGS|12|7|Qui dixerunt ei: " Si hodie oboedieris populo huic et servieris et petitioni eorum cesseris locutusque fueris ad eos verba lenia, erunt tibi servi cunctis diebus ".
1KGS|12|8|Qui dereliquit consilium senum, quod dederant ei, et adhibuit adulescentes, qui nutriti fuerant cum eo et assistebant illi,
1KGS|12|9|dixitque ad eos: " Quod mihi datis consilium, ut respondeam populo huic, qui dixerunt mihi: "Levius fac iugum, quod imposuit pater tuus super nos"?.
1KGS|12|10|Et dixerunt ei iuvenes, qui nutriti fuerant cum eo: " Sic loquere populo huic, qui locuti sunt ad te dicentes: "Pater tuus aggravavit iugum nostrum, tu releva nos"; sic loqueris ad eos: Minimus digitus meus grossior est lumbis patris mei.
1KGS|12|11|Et nunc, pater meus posuit super vos iugum grave, ego autem addam super iugum vestrum; pater meus cecidit vos flagellis, ego autem caedam scorpionibus ".
1KGS|12|12|Venit ergo Ieroboam et omnis populus ad Roboam die tertia, sicut locutus fuerat rex dicens: " Revertimini ad me die tertia ".
1KGS|12|13|Responditque rex populo dura, derelicto consilio seniorum, quod ei dederant,
1KGS|12|14|et locutus est eis secundum consilium iuvenum dicens: Pater meus aggravavit iugum vestrum,ego autem addam iugo vestro;pater meus cecidit vos flagellis,ego autem caedam vos scorpionibus ".
1KGS|12|15|Ergo non acquievit rex populo, quoniam dispositum erat a Domino, ut suscitaret verbum suum, quod locutus fuerat in manu Ahiae Silonitae ad Ieroboam filium Nabat.
1KGS|12|16|Videns itaque omnis Israel quod noluisset eos audire rex, respondit ei dicens: Quae nobis pars in David,vel quae hereditas in filio Isai?Vade in tabernacula tua, Israel!Nunc vide domum tuam, David! ". Et abiit Israel in tabernacula sua.
1KGS|12|17|Super filios autem Israel, quicumque habitabant in civitatibus Iudae, regnavit Roboam.
1KGS|12|18|Misit rex Roboam Adoniram, qui erat super servitutem; et lapidavit eum omnis Israel, et mortuus est. Porro rex Roboam festinus ascendit currum et fugit in Ierusalem.
1KGS|12|19|Recessitque Israel a domo David usque in praesentem diem.
1KGS|12|20|Factum est autem cum audisset omnis Israel quod reversus esset Ieroboam, miserunt et vocaverunt eum, congregato coetu, et constituerunt eum regem super omnem Israel; nec secutus est quisquam domum David praeter tribum Iudae solam.
1KGS|12|21|Venit autem Roboam Ierusalem et congrcgavit universam domum Iudae et tribum Beniamin, centum octoginta milia electorum virorum bellatorum, ut pugnaret contra domum Israel et reduceret regnum Roboam filio Salomonis.
1KGS|12|22|Factus est vero sermo Domini ad Semeiam virum Dei dicens:
1KGS|12|23|" Loquere ad Roboam filium Salomonis regem Iudae et ad omnem domum Iudae et Beniamin et reliquos de populo dicens:
1KGS|12|24|Haec dicit Dominus: Non ascendetis neque bellabitis contra fratres vestros, filios Israel; revertatur vir in domum suam; a me enim factum est hoc ". Audierunt sermonem Domini et reversi sunt de itinere, sicut eis praeceperat Dominus.
1KGS|12|25|Aedificavit autem Ieroboam Sichem in monte Ephraim et habitavit ibi; et egressus inde aedificavit Phanuel.
1KGS|12|26|Dixitque Ieroboam in corde suo: " Nunc revertetur regnum ad domum David,
1KGS|12|27|si ascenderit populus iste, ut faciat sacrificia in domo Domini in Ierusalem, et convertetur cor populi huius ad dominum suum Roboam regem Iudae, interficientque me et revertentur ad Roboam regem Iudae ".
1KGS|12|28|Et excogitato consilio, fecit rex duos vitulos aureos et dixit ad populum: " Nolite ultra ascendere in Ierusalem! Ecce dii tui, Israel, qui te eduxerunt de terra Aegypti ".
1KGS|12|29|Posuitque unum in Bethel et alterum donavit in Dan;
1KGS|12|30|et factum est hoc in peccatum: ibat enim populus coram uno usque in Dan.
1KGS|12|31|Et fecit fana in excelsis et sacerdotes de extremis populi, qui non erant de filiis Levi.
1KGS|12|32|Constituitque diem sollemnem in mense octavo, quinta decima die mensis, in similitudinem sollemnitatis, quae celebratur in Iuda. Et ascendit altare; sic fecit in Bethel, ut immolaret vitulis, quos fabricatus erat; constituitque in Bethel sacerdotes excelsorum, quae fecerat.
1KGS|12|33|Et ascendit super altare, quod exstruxerat in Bethel, quinta decima die mensis octavi, quem finxerat de corde suo; et fecit sollemnitatem filiis Israel et ascendit super altare, ut adoleret.
1KGS|13|1|Et ecce vir Dei venit de Iuda in sermone Domini in Bethel, Ieroboam stante super altare ad adolendum;
1KGS|13|2|et exclamavit contra altare in sermone Domini et ait: " Altare, altare, haec dicit Dominus: Ecce filius nascetur domui David, Iosias nomine, et immolabit super te sacerdotes excelsorum, qui nunc in te immolant, et ossa hominum super te incendent ".
1KGS|13|3|Deditque in illa die signum dicens: " Hoc erit signum, quod locutus est Dominus: ecce altare scindetur, et effundetur cinis, qui in eo est ".
1KGS|13|4|Cumque audisset rex sermonem hominis Dei, quem inclamaverat contra altare in Bethel, extendit manum suam de altari dicens: " Apprehendite eum! ". Et exaruit manus eius, quam extenderat contra eum, nec valuit retrahere eam ad se.
1KGS|13|5|Altare quoque scissum est, et effusus est cinis de altari iuxta signum, quod praedixerat vir Dei in sermone Domini.
1KGS|13|6|Et ait rex ad virum Dei: " Deprecare faciem Domini Dei tui et ora pro me, ut restituatur manus mea mihi ". Oravit vir Dei faciem Domini, et reversa est manus regis ad eum et facta est sicut prius fuerat.
1KGS|13|7|Locutus est autem rex ad virum Dei: " Veni mecum domum, ut prandeas, et dabo tibi munera ".
1KGS|13|8|Responditque vir Dei ad regem: " Si dederis mihi mediam partem domus tuae, non veniam tecum nec comedam panem neque bibam aquam in loco isto;
1KGS|13|9|sic enim mandatum est mihi in sermone Domini praecipientis: "Non comedes panem neque bibes aquam nec reverteris per viam, qua venisti" ".
1KGS|13|10|Abiit ergo per aliam viam et non est reversus per iter, quo venerat in Bethel.
1KGS|13|11|Prophetes autem quidam senex habitabat in Bethel; ad quem venerunt filii sui et narraverunt ei omnia opera, quae fecerat vir Dei illa die in Bethel, et verba, quae locutus fuerat ad regem, narraverunt quoque patri suo.
1KGS|13|12|Et dixit eis pater eorum: " Per quam viam abiit? ". Ostenderunt ei filii sui viam, per quam abierat vir Dei, qui venerat de Iuda.
1KGS|13|13|Et ait filiis suis: " Sternite mihi asinum ". Qui cum stravissent, ascendit
1KGS|13|14|et abiit post virum Dei et invenit eum sedentem subtus terebinthum et ait illi: " Tune es vir Dei, qui venisti de Iuda?". Respondit ille: " Ego sum ".
1KGS|13|15|Dixit ad eum: " Veni mecum domum, ut comedas panem ".
1KGS|13|16|Qui ait: " Non possum reverti neque venire tecum nec comedam panem neque bibam aquam in loco isto;
1KGS|13|17|sic enim dictum est mihi in sermone Domini: "Non comedes panem et non bibes ibi aquam nec reverteris per viam, qua ieris" ".
1KGS|13|18|Qui ait illi: " Et ego propheta sum similis tui; et angelus locutus est mihi in sermone Domini dicens: "Reduc eum tecum in domum tuam, et comedat panem et bibat aquam" ". Fefellit eum
1KGS|13|19|et reduxit secum; comedit ergo panem in domo eius et bibit aquam.
1KGS|13|20|Cumque sederent ad mensam, factus est sermo Domini ad prophetam, qui reduxerat eum,
1KGS|13|21|et exclamavit ad virum Dei, qui venerat de Iuda, dicens: " Haec dicit Dominus: Quia non oboediens fuisti ori Domini et non custodisti mandatum, quod praecepit tibi Dominus Deus tuus,
1KGS|13|22|et reversus es et comedisti panem et bibisti aquam in loco, in quo praecepit tibi, ne comederes panem neque biberes aquam, non inferetur cadaver tuum in sepulcrum patrum tuorum ".
1KGS|13|23|Cumque comedisset panem et bibisset, stravit sibi asinum prophetae, qui reduxerat eum;
1KGS|13|24|et, cum abisset, invenit eum leo in via et occidit, et erat cadaver eius proiectum in itinere; asinus autem stabat iuxta illum, et leo stabat iuxta cadaver.
1KGS|13|25|Et ecce viri transeuntes viderunt cadaver proiectum in via et leonem stantem iuxta cadaver; et venerunt et divulgaverunt in civitate, in qua prophetes ille senex habitabat.
1KGS|13|26|Quod cum audisset propheta ille, qui reduxerat eum de via, ait: " Vir Dei est, qui inoboediens fuit ori Domini, et tradidit eum Dominus leoni; et confregit eum et occidit iuxta verbum Domini, quod locutus est ei ".
1KGS|13|27|Dixitque ad filios suos: " Sternite mihi asinum! ". Qui cum stravissent,
1KGS|13|28|et ille abisset, invenit cadaver eius proiectum in via et asinum et leonem stantes iuxta cadaver; non comedit leo de cadavere nec laesit asinum.
1KGS|13|29|Tulit ergo prophetes cadaver viri Dei et posuit illud super asinum et reversus intulit in civitatem prophetae senis, ut plangerent eum et sepelirent.
1KGS|13|30|Et posuit cadaver eius in sepulcro suo, et planxerunt eum: " Heu, heu, mi frater! ".
1KGS|13|31|Cumque sepelissent eum, dixit ad filios suos: " Cum mortuus fuero, sepelite me in sepulcro, in quo vir Dei sepultus est; iuxta ossa eius ponite ossa mea.
1KGS|13|32|Profecto enim veniet sermo, quem praedixit in sermone Domini contra altare, quod est in Bethel, et contra omnia fana excelsorum, quae sunt in urbibus Samariae ".
1KGS|13|33|Post haec non est reversus Ieroboam de via sua pessima, sed iterum faciebat de novissimis populi sacerdotes excelsorum; quicumque volebat, implebat eius manum, ut fieret sacerdos excelsorum.
1KGS|13|34|Et propter hanc causam peccavit domus Ieroboam, et eversa est et deleta de superficie terrae.
1KGS|14|1|In tempore illo aegrotavit Abia filius Ieroboam,
1KGS|14|2|dixitque Ieroboam uxori suae: " Surge et commuta habitum, ne cognoscaris quod sis uxor Ieroboam, et vade in Silo, ubi est Ahias propheta, qui locutus est mihi quod regnaturus essem super populum hunc.
1KGS|14|3|Tolle quoque in manu tua decem panes et crustula et vas mellis et vade ad illum: ipse indicabit tibi quid eventurum sit puero ".
1KGS|14|4|Fecit, ut dixerat, uxor Ieroboam et consurgens abiit in Silo et venit in domum Ahiae; at ille non poterat videre, quia caligaverant oculi eius prae senectute.
1KGS|14|5|Dixerat autem Dominus ad Ahiam: " Ecce uxor Ieroboam ingredietur, ut consulat te super filio suo, qui aegrotat; haec et haec loqueris ei. Cum intret, simulabit se peregrinam esse ".
1KGS|14|6|Cum ergo audiret Ahias sonitum pedum eius introeuntis per ostium, ait: " Ingredere, uxor Ieroboam. Quare aliam te esse simulas? Ego autem missus sum ad te durus nuntius.
1KGS|14|7|Vade et dic Ieroboam: "Haec dicit Dominus, Deus Israel: Quia exaltavi te de medio populi et dedi te ducem super populum meum Israel
1KGS|14|8|et scidi regnum a domo David et dedi illud tibi, et non fuisti sicut servus meus David, qui custodivit mandata mea et secutus est me in toto corde suo faciens quod placitum esset in conspectu meo,
1KGS|14|9|sed operatus es mala super omnes, qui fuerunt ante te, et fecisti tibi deos alienos et conflatiles, ut me ad iracundiam provocares, me autem proiecisti post tergum tuum:
1KGS|14|10|idcirco ecce ego inducam mala super domum Ieroboam et percutiam de Ieroboam quidquid masculini sexus, impuberem et puberem in Israel; et mundabo reliquias domus Ieroboam, sicut mundari solet fimus usque ad purum.
1KGS|14|11|Qui mortui fuerint de Ieroboam in civitate, comedent eos canes; qui autem mortui fuerint in agro, vorabunt eos aves caeli, quia Dominus locutus est.
1KGS|14|12|Tu igitur surge et vade in domum tuam, et in ipso introitu pedum tuorum in urbem morietur puer,
1KGS|14|13|et planget eum omnis Israel et sepeliet; iste enim solus inferetur de Ieroboam in sepulcrum, quia inventum est in eo, quod bonum erat Domino, Deo Israel, in domo Ieroboam.
1KGS|14|14|Constituet autem sibi Dominus regem super Israel, qui percutiat domum Ieroboam.
1KGS|14|15|Et percutiet Dominus Israel, ut moveatur sicut arundo in aqua, et evellet Israel de terra bona hac, quam dedit patribus eorum; et ventilabit eos trans Flumen, quia fecerunt sibi palos, ut irritarent Dominum.
1KGS|14|16|Et tradet Dominus Israel propter peccata Ieroboam, qui peccavit et peccare fecit Israel" ".
1KGS|14|17|Surrexit itaque uxor Ieroboam et abiit et venit in Thersa; cumque illa ingrederetur limen domus, puer mortuus est.
1KGS|14|18|Et sepelierunt eum, et planxit illum omnis Israel iuxta sermonem Domini, quem locutus est in manu servi sui Ahiae prophetae.
1KGS|14|19|Reliqua autem gestorum Ieroboam, quomodo pugnaverit et quomodo regnaverit, ecce scripta sunt in libro annalium regum Israel.
1KGS|14|20|Dies autem, quibus regnavit Ieroboam, viginti duo anni sunt; et dormivit cum patribus suis. Regnavitque Nadab filius eius pro eo.
1KGS|14|21|Porro Roboam filius Salomonis regnavit in Iuda. Quadraginta et unius anni erat Roboam, cum regnare coepisset, et decem et septem annos regnavit in Ierusalem civitate, quam elegit Dominus, ut poneret nomen suum ibi ex omnibus tribubus Israel. Nomen autem matris eius Naama Ammanites.
1KGS|14|22|Et fecit Iuda malum coram Domino, et irritaverunt eum super omnibus, quae fecerant patres eorum in peccatis suis, quae peccaverant;
1KGS|14|23|aedificaverunt enim et ipsi sibi excelsa et lapides et palos super omnem collem excelsum et subter omnem arborem frondosam.
1KGS|14|24|Sed et prostibula fuerunt in terra; feceruntque omnes abominationes gentium, quas attrivit Dominus ante faciem filiorum Israel.
1KGS|14|25|In quinto autem anno regni Roboam ascendit Sesac rex Aegypti in Ierusalem
1KGS|14|26|et tulit thesauros domus Domini et thesauros regios et universa diripuit, scuta quoque aurea omnia, quae fecerat Salomon.
1KGS|14|27|Pro quibus fecit rex Roboam scuta aerea et tradidit ea in manu ducum cursorum, qui excubabant ante ostium domus regis.
1KGS|14|28|Cumque ingrederetur rex in domum Domini, portabant ea cursores et postea reportabant ad armamentarium cursorum.
1KGS|14|29|Reliqua autem gestorum Roboam et omnia, quae fecit, ecce scripta sunt in libro annalium regum Iudae.
1KGS|14|30|Fuitque bellum inter Roboam et Ieroboam cunctis diebus.
1KGS|14|31|Dormivit itaque Roboam cum patribus suis et sepultus est cum eis in civitate David; nomen autem matris eius Naama Ammanites. Et regnavit Abiam filius eius pro eo.
1KGS|15|1|Igitur in octavo decimo anno regni Ieroboam filii Nabat regnavit Abiam super Iudam.
1KGS|15|2|Tribus annis regnavit in Ierusalem; nomen matris eius Maacha filia Abessalom.
1KGS|15|3|Ambulavitque in omnibus peccatis patris sui, quae fecerat ante eum; nec erat cor eius perfectum cum Domino Deo suo sicut cor David patris eius.
1KGS|15|4|Sed propter David dedit ei Dominus Deus suus lucernam in Ierusalem, ut suscitaret filium eius post eum et statueret Ierusalem;
1KGS|15|5|eo quod fecisset David rectum in oculis Domini et non declinasset ab omnibus, quae praeceperat ei, cunctis diebus vitae suae, excepta re Uriae Hetthaei. (6)
1KGS|15|6|attamen bellum fuit inter Roboam et inter Hieroboam omni tempore vitae eius
1KGS|15|7|Reliqua autem gestorum Abiam et omnia, quae fecit, nonne haec scripta sunt in libro annalium regum Iudae? Fuitque bellum inter Abiam et inter Ieroboam.
1KGS|15|8|Et dormivit Abiam cum patribus suis, et sepelierunt eum in civitate David; regnavitque Asa filius eius pro eo.
1KGS|15|9|In anno ergo vicesimo Ieroboam regis Israel regnavit Asa rex Iudae
1KGS|15|10|et quadraginta et uno anno regnavit in Ierusalem. Nomen matris eius Maacha filia Abessalom.
1KGS|15|11|Et fecit Asa rectum ante conspectum Domini sicut David pater eius.
1KGS|15|12|Et abstulit prostibula de terra purgavitque universas sordes idolorum, quae fecerant patres eius.
1KGS|15|13|Insuper et Maacham matrem suam amovit, ne esset domina, eo quod fecisset abominationem Aserae; confregitque Asa simulacrum turpissimum et combussit in torrente Cedron.
1KGS|15|14|Excelsa autem non abstulit; verumtamen cor Asa perfectum erat coram Domino cunctis diebus suis.
1KGS|15|15|Et intulit ea, quae sanctificaverat pater suus et quae ipse voverat, in domum Domini, argentum et aurum et vasa.
1KGS|15|16|Bellum autem erat inter Asa et Baasa regem lsrael cunctis diebus eorum.
1KGS|15|17|Ascendit quoque Baasa rex Israel in Iudam et aedificavit Rama, ut non posset quispiam egredi vel ingredi de parte Asa regis Iudae.
1KGS|15|18|Tollens itaque Asa omne argentum et aurum, quod remanserat in thesauris domus Domini et in thesauris domus regiae, dedit illud in manu servorum suorum et misit ad Benadad filium Tabremmon filii Hezion regem Syriae, qui habitabat in Damasco, dicens:
1KGS|15|19|" Foedus est inter me et te et inter patrem meum et patrem tuum; ideo misi tibi munera, argentum et aurum, et peto, ut irritum facias foedus, quod habes cum Baasa rege Israel, et recedat a me ".
1KGS|15|20|Acquiescens Benadad regi Asa misit principes exercituum suorum in civitates Israel, et percusserunt Ahion et Dan et Abelbethmaacha et universam Chenereth cum omni terra Nephthali.
1KGS|15|21|Quod cum audisset Baasa, cessavit aedificare Rama et reversus est in Thersa.
1KGS|15|22|Rex autem Asa convocavit omnem Iudam, nullo excusato; et tulerunt lapides Rama et ligna eius, quibus aedificaverat Baasa, et exstruxit de eis rex Asa Gabaa Beniamin et Maspha.
1KGS|15|23|Reliqua autem omnium gestorum Asa et universa fortitudo eius et cuncta, quae fecit, et civitates, quas exstruxit, nonne haec scripta sunt in libro annalium regum Iudae? Verumtamen in tempore senectutis suae doluit pedes;
1KGS|15|24|et dormivit cum patribus suis et sepultus est cum eis in civitate David patris sui. Regnavitque Iosaphat filius eius pro eo.
1KGS|15|25|Nadab vero filius Ieroboam regnavit super Israel anno secundo Asa regis Iudae; regnavitque super Israel duobus annis.
1KGS|15|26|Et fecit, quod malum est in conspectu Domini, et ambulavit in viis patris sui et in peccato eius, quo peccare fecit Israel.
1KGS|15|27|Insidiatus est autem ei Baasa filius Ahiae de domo Issachar et percussit eum in Gebbethon, quae est urbs Philisthinorum; siquidem Nadab et omnis Israel obsidebant Gebbethon.
1KGS|15|28|Interfecit igitur illum Baasa in anno tertio Asa regis Iudae et regnavit pro eo.
1KGS|15|29|Cumque regnasset, percussit omnem domum Ieroboam; non dimisit ne unam quidem animam de semine eius, donec deleret eam iuxta verbum Domini, quod locutus fuerat in manu servi sui Ahiae Silonitis
1KGS|15|30|propter peccata Ieroboam, quae peccaverat et quibus peccare fecerat Israel, et propter delictum, quo irritaverat Dominum, Deum Israel.
1KGS|15|31|Reliqua autem gestorum Nadab et omnia, quae fortiter operatus est, nonne haec scripta sunt in libro annalium regum Israel?
1KGS|15|32|Fuitque bellum inter Asa et Baasa regem Israel cunctis diebus eorum.
1KGS|15|33|Anno tertio Asa regis Iudae regnavit Baasa filius Ahiae super omnem Israel in Thersa viginti quattuor annis;
1KGS|15|34|et fecit malum coram Domino ambulavitque in via Ieroboam et in peccato eius, quo peccare fecit Israel.
1KGS|16|1|Factus est autem sermo Domini ad Iehu filium Hanani contra Baasa dicens:
1KGS|16|2|" Pro eo quod exaltavi te de pulvere et posui te ducem super populum meum Israel, tu autem ambulasti in via Ieroboam et peccare fecisti populum meum Israel, ut me irritares in peccatis eorum,
1KGS|16|3|ecce ego demetam posteriora Baasa et posteriora domus eius et faciam domum tuam sicut domum Ieroboam filii Nabat.
1KGS|16|4|Qui mortuus fuerit de Baasa in civitate, comedent eum canes; et, qui mortuus fuerit ex eo in agro, comedent eum volucres caeli".
1KGS|16|5|Reliqua autem gestorum Baasa et quaecumque fecit et fortitudo eius, nonne haec scripta sunt in libro annalium regum Israel?
1KGS|16|6|Dormivit ergo Baasa cum patribus suis sepultusque est in Thersa; et regnavit Ela filius eius pro eo.
1KGS|16|7|Sed et in manu Iehu filii Hanani prophetae verbum Domini factum est ad Baasa et ad domum eius propter omne malum, quod fecerat coram Domino ad irritandum eum in operibus manuum suarum, ut fieret sicut domus Ieroboam, eo quod percussisset eam.
1KGS|16|8|Anno vicesimo sexto Asa regis Iudae regnavit Ela filius Baasa super Israel in Thersa duobus annis.
1KGS|16|9|Et rebellavit contra eum servus suus Zamri dux mediae partis curruum. Erat autem Ela in Thersa bibens et temulentus in domo Arsa praefecti domus in Thersa;
1KGS|16|10|irruens ergo Zamri percussit et occidit eum anno vicesimo septimo Asa regis Iudae et regnavit pro eo.
1KGS|16|11|Cumque regnasset et sedisset super solium eius, percussit omnem domum Baasa et non dereliquit ex eo quidquid masculini sexus et propinquos et amicos eius.
1KGS|16|12|Delevitque Zamri omnem domum Baasa iuxta verbum Domini, quod locutus fuerat ad Baasa in manu Iehu prophetae,
1KGS|16|13|propter universa peccata Baasa et peccata Ela filii eius, qui peccaverunt et peccare fecerunt Israel provocantes Dominum, Deum Israel, in vanitatibus suis.
1KGS|16|14|Reliqua autem gestorum Ela et omnia, quae fecit, nonne haec scripta sunt in libro annalium regum Israel?
1KGS|16|15|Anno vicesimo septimo Asa regis Iudae regnavit Zamri septem diebus in Thersa. Porro exercitus obsidebat Gebbethon urbem Philisthinorum.
1KGS|16|16|Cumque audisset rebellasse Zamri et occidisse regem, fecit sibi regem omnis Israel Amri, qui erat princeps militiae super Israel in die illa in castris.
1KGS|16|17|Ascendit ergo Amri et omnis Israel cum eo de Gebbethon, et obsidebant Thersa;
1KGS|16|18|videns autem Zamri quod expugnanda esset civitas, ingressus est palatium et succendit super se domum regiam et mortuus est igne
1KGS|16|19|in peccatis suis, quae peccaverat faciens malum coram Domino et ambulans in via Ieroboam et in peccato eius, quo fecit peccare Israel.
1KGS|16|20|Reliqua autem gestorum Zamri et rebellio, quam fecit, nonne haec scripta sunt in libro annalium regum Israel?
1KGS|16|21|Tunc divisus est populus Israel in duas partes: media pars populi sequebatur Thebni filium Gineth, ut constitueret eum regem, et media pars Amri.
1KGS|16|22|Praevaluit autem populus, qui erat cum Amri, populo, qui sequebatur Thebni filium Gineth; mortuusque est Thebni, et regnavit Amri.
1KGS|16|23|Anno tricesimo primo Asa regis Iudae regnavit Amri super Israel duodecim annis; in Thersa regnavit sex annis.
1KGS|16|24|Emitque montem Samariae a Somer duobus talentis argenti et aedificavit eum et vocavit nomen civitatis, quam exstruxerat, nomine Somer domini montis Samariae.
1KGS|16|25|Fecit autem Amri malum in conspectu Domini et operatus est nequiter super omnes, qui fuerunt ante eum;
1KGS|16|26|ambulavitque in omni via Ieroboam filii Nabat et in peccato eius, quo peccare fecerat Israel, ut irritaret Dominum, Deum Israel, in vanitatibus suis.
1KGS|16|27|Reliqua autem gestorum Amri et proelia eius, quae fortiter gessit, nonne haec scripta sunt in libro annalium regum Israel?
1KGS|16|28|Et dormivit Amri cum patribus suis et sepultus est in Samaria; regnavitque Achab filius eius pro eo.
1KGS|16|29|Achab vero filius Amri regnavit super Israel anno tricesimo octavo Asa regis Iudae; et regnavit Achab filius Amri super Israel in Samaria viginti et duobus annis.
1KGS|16|30|Et fecit Achab filius Amri malum in conspectu Domini super omnes, qui fuerunt ante eum.
1KGS|16|31|Nec suffecit ei, ut ambularet in peccatis Ieroboam filii Nabat; insuper duxit uxorem Iezabel filiam Ethbaal regis Sidoniorum et abiit et servivit Baal et adoravit eum.
1KGS|16|32|Et posuit aram Baal in templo Baal, quod aedificaverat in Samaria,
1KGS|16|33|et fecit Achab palum. Et addidit Achab in opere suo irritans Dominum, Deum Israel, super omnes reges Israel, qui fuerant ante eum.
1KGS|16|34|In diebus eius aedificavit Hiel de Bethel Iericho; in Abiram primitivo suo fundavit eam et in Segub novissimo suo posuit portas eius, iuxta verbum Domini, quod locutus fuerat in manu Iosue filii Nun.
1KGS|17|1|Et dixit Elias Thesbites de Thesbi in Galaad ad Achab: " Vivit Dominus, Deus Israel, in cuius conspectu sto. Non erit annis his ros et pluvia, nisi iuxta oris mei verba! ".
1KGS|17|2|Et factum est verbum Domini ad eum dicens:
1KGS|17|3|" Recede hinc et vade contra orientem et abscondere in torrente Charith, qui est contra Iordanem,
1KGS|17|4|et ibi de torrente bibes; corvisque praecepi, ut pascant te ibi ".
1KGS|17|5|Abiit ergo et fecit iuxta verbum Domini; cumque abisset, sedit in torrente Charith, qui est contra Iordanem.
1KGS|17|6|Corvi quoque deferebant ei panem et carnes mane, similiter panem et carnes vesperi; et bibebat de torrente.
1KGS|17|7|Post dies autem siccatus est torrens; non enim pluerat super terram.
1KGS|17|8|Factus est igitur sermo Domini ad eum dicens:
1KGS|17|9|" Surge et vade in Sarepta Sidoniorum et manebis ibi; praecepi enim ibi mulieri viduae, ut pascat te ".
1KGS|17|10|Surrexit et abiit Sareptam. Cumque venisset ad portam civitatis, apparuit ei mulier vidua colligens ligna; et vocavit eam dixitque: " Da mihi paululum aquae in vase, ut bibam ".
1KGS|17|11|Cumque illa pergeret, ut afferret, clamavit post tergum eius dicens: " Affer mihi, obsecro, et buccellam panis in manu tua ".
1KGS|17|12|Quae respondit: " Vivit Dominus Deus tuus, non habeo panem, nisi quantum pugillus capere potest farinae in hydria et paululum olei in lecytho. En colligo duo ligna, ut ingrediar et faciam illud mihi et filio meo, ut comedamus et moriamur ".
1KGS|17|13|Ad quam Elias ait: " Noli timere, sed vade et fac, sicut dixisti; verumtamen mihi primum fac de ipsa farinula subcinericium panem parvulum et affer ad me; tibi autem et filio tuo facies postea.
1KGS|17|14|Haec autem dicit Dominus, Deus Israel: "Hydria farinae non deficiet, nec lecythus olei minuetur usque ad diem, in qua daturus est Dominus pluviam super faciem terrae" ".
1KGS|17|15|Quae abiit et fecit iuxta verbum Eliae et comedit illa et ipse et domus eius per dies.
1KGS|17|16|Hydria farinae non defecit, et lecythus olei non est imminutus iuxta verbum Domini, quod locutus fuerat in manu Eliae.
1KGS|17|17|Factum est autem post haec, aegrotavit filius mulieris matris familiae; et erat languor fortis nimis, ita ut non remaneret in eo halitus.
1KGS|17|18|Dixit ergo ad Eliam: " Quid mihi et tibi, vir Dei? Ingressus es ad me, ut rememorarentur iniquitates meae, et interficeres filium meum? ".
1KGS|17|19|Et ait ad eam: " Da mihi filium tuum ". Tulitque eum de sinu illius et portavit in cenaculum, ubi ipse manebat, et posuit super lectulum suum;
1KGS|17|20|clamavitque ad Dominum et dixit: " Domine Deus meus, etiamne viduam, apud quam ego ut hospes habito, afflixisti, ut interficeres filium eius?.
1KGS|17|21|Et expandit se atque mensus est super puerum tribus vicibus et clamavit ad Dominum et ait: " Domine Deus meus, revertatur, oro, anima pueri huius in viscera eius ".
1KGS|17|22|Et exaudivit Dominus vocem Eliae, et reversa est anima pueri intra eum, et revixit.
1KGS|17|23|Tulitque Elias puerum et deposuit eum de cenaculo in inferiorem domum et tradidit matri suae et ait illi: " En vivit filius tuus ".
1KGS|17|24|Dixitque mulier ad Eliam: " Nunc in isto cognovi quoniam vir Dei es tu, et verbum Domini in ore tuo verum est ".
1KGS|18|1|Post dies multos factum est verbum Domini ad Eliam in anno tertio dicens: " Vade et ostende te Achab, ut dem pluviam super faciem terrae ".
1KGS|18|2|Ivit ergo Elias, ut ostenderet se Achab.Erat autem fames vehemens in Samaria.
1KGS|18|3|Vocavitque Achab Abdiam dispensatorem domus suae. Abdias autem timebat Dominum valde;
1KGS|18|4|nam, cum interficeret Iezabel prophetas Domini, tulit ille centum prophetas et abscondit eos quinquagenos et quinquagenos in speluncis et pavit eos pane et aqua.
1KGS|18|5|Dixit ergo Achab ad Abdiam: " Vade in terra ad universos fontes aquarum et in cunctas valles, si forte invenire possimus herbam, ut salvemus equos et mulos et nullum de iumentis interficere debeamus ".
1KGS|18|6|Diviseruntque sibi regiones, ut circuirent eas: Achab ibat per viam unam, et Abdias per viam alteram seorsum.
1KGS|18|7|Cumque esset Abdias in via, Elias occurrit ei; qui cum cognovisset eum, cecidit super faciem suam et ait: " Num tu es, domine mi, Elias? ".
1KGS|18|8|Cui ille respondit: " Ego. Vade, dic domino tuo: "Adest Elias" ".
1KGS|18|9|Et ille: " Quid peccavi, inquit, quoniam trades me servum tuum in manu Achab, ut interficiat me?
1KGS|18|10|Vivit Dominus Deus tuus, non est gens aut regnum, quo non miserit dominus meus te requirens et, respondentibus cunctis: "Non est hic", adiuravit regna singula et gentes, eo quod minime reperireris.
1KGS|18|11|Et nunc dicis mihi: "Vade et dic domino tuo: Adest Elias".
1KGS|18|12|Cumque recessero a te, spiritus Domini asportabit te in locum, quem ego ignoro; et ingressus nuntiabo Achab, et non inveniet te et interficiet me. Servus autem tuus timet Dominum ab infantia sua.
1KGS|18|13|Numquid non indicatum est domino meo quid fecerim, cum interficeret Iezabel prophetas Domini: quod absconderim de prophetis Domini centum viros, quinquagenos et quinquagenos in speluncis et paverim eos pane et aqua?
1KGS|18|14|Et nunc tu dicis: "Vade et dic domino tuo: Adest Elias", ut interficiat me ".
1KGS|18|15|Dixit Elias: " Vivit Dominus exercituum ante cuius vultum sto: hodie apparebo ei ".
1KGS|18|16|Abiit ergo Abdias in occursum Achab et indicavit ei.Venitque Achab in occursum Eliae
1KGS|18|17|et, cum vidisset eum, ait: " Tune es, qui conturbas Israel? ".
1KGS|18|18|Et ille ait: " Non turbavi Israel, sed tu et domus patris tui, qui dereliquistis mandata Domini, et secutus es Baalim.
1KGS|18|19|Verumtamen nunc mitte et congrega ad me universum Israel in monte Carmeli et prophetas Baal quadringentos quinquaginta prophetasque Aserae quadringentos, qui comedunt de mensa Iezabel ".
1KGS|18|20|Misit Achab ad omnes filios Israel et congregavit prophetas in monte Carmeli.
1KGS|18|21|Accedens autem Elias ad omnem populum ait: " Usquequo claudicatis in duas partes? Si Dominus est Deus, sequimini eum; si autem Baal, sequimini illum ". Et non respondit ei populus verbum.
1KGS|18|22|Et ait rursus Elias ad populum: " Ego remansi propheta Domini solus; prophetae autem Baal quadringenti et quinquaginta viri sunt.
1KGS|18|23|Dentur nobis duo boves, et illi eligant sibi bovem unum et in frusta caedentes ponant super ligna; ignem autem non supponant. Et ego faciam bovem alterum et imponam super ligna; ignemque non supponam.
1KGS|18|24|Invocate nomen dei vestri, et ego invocabo nomen Domini; et Deus, qui exaudierit per ignem, ipse est Deus! ". Respondens omnis populus ait: " Optima propositio ".
1KGS|18|25|Dixit ergo Elias prophetis Baal: " Eligite vobis bovem unum et facite primi, quia vos plures estis; et invocate nomen dei vestri ignemque non supponatis ".
1KGS|18|26|Qui cum tulissent bovem, quem dederat eis, fecerunt et invocabant nomen Baal de mane usque ad meridiem dicentes: " Baal, exaudi nos! ". Et non erat vox, nec qui responderet. Saliebantque in circuitu altaris, quod fecerant.
1KGS|18|27|Cumque esset iam meridies, illudebat eis Elias dicens: " Clamate voce maiore; deus enim est et forsitan occupatus est aut secessit aut in itinere aut certe dormit, ut excitetur ".
1KGS|18|28|Clamabant ergo voce magna et incidebant se iuxta ritum suum cultris et lanceolis, donec perfunderentur sanguine.
1KGS|18|29|Postquam autem transiit meridies, et, illis prophetantibus, venerat tempus, quo sacrificium offerri solet, nec audiebatur vox, neque aliquis respondebat nec attendebat orantes,
1KGS|18|30|dixit Elias omni populo: " Venite ad me ". Et, accedente ad se populo, curavit altare Domini, quod destructum fuerat;
1KGS|18|31|et tulit duodecim lapides iuxta numerum tribuum filiorum Iacob, ad quem factus est sermo Domini dicens: " Israel erit nomen tuum ".
1KGS|18|32|Et aedificavit lapidibus altare in nomine Domini fecitque aquaeductum quasi pro duobus satis in circuitu altaris
1KGS|18|33|et composuit ligna divisitque per membra bovem et posuit super ligna
1KGS|18|34|et ait: " Implete quattuor hydrias aqua et fundite super holocaustum et super ligna ". Rursumque dixit: " Etiam secundo hoc facite ". Qui cum fecissent et secundo, ait: " Etiam tertio idipsum facite ". Feceruntque et tertio,
1KGS|18|35|et currebant aquae circum altare, et fossa aquaeductus repleta est.
1KGS|18|36|Cumque iam tempus esset, ut offerretur sacrificium, accedens Elias propheta ait: " Domine, Deus Abraham, Isaac et Israel, hodie ostende quia tu es Deus in Israel, et ego servus tuus et iuxta praeceptum tuum feci omnia haec.
1KGS|18|37|Exaudi me, Domine, exaudi me, ut discat populus iste quia tu, Domine, es Deus et tu convertisti cor eorum iterum! ".
1KGS|18|38|Cecidit autem ignis Domini et voravit holocaustum et ligna et lapides, pulverem quoque et aquam, quae erat in aquaeductu lambens.
1KGS|18|39|Quod cum vidisset omnis populus, cecidit in faciem suam et ait: " Dominus ipse est Deus, Dominus ipse est Deus! ".
1KGS|18|40|Dixitque Elias ad eos: " Apprehendite prophetas Baal, et ne unus quidem effugiat ex eis! ". Quos cum comprehendissent, duxit eos Elias ad torrentem Cison et interfecit eos ibi.
1KGS|18|41|Et ait Elias ad Achab: " Ascende, comede et bibe, quia sonus multae pluviae est ".
1KGS|18|42|Ascendit Achab, ut comederet et biberet. Elias autem ascendit in verticem Carmeli et pronus in terram posuit faciem inter genua sua
1KGS|18|43|et dixit ad puerum suum: " Ascende et prospice contra mare ". Qui, cum ascen disset et contemplatus esset, ait: " Non est quidquam ". Et rursum ait illi: " Revertere septem vicibus ".
1KGS|18|44|In septima autem vice dixit: " Ecce nubecula parva quasi manus hominis ascendit de mari ". Et ait: " Ascende et dic Achab: Iunge et descende, ne occupet te pluvia! ".
1KGS|18|45|Et factum est interea: ecce caeli contenebrati sunt, et nubes et ventus, et facta est pluvia grandis. Ascendens itaque Achab abiit in Iezrahel.
1KGS|18|46|Et manus Domini facta est super Eliam; accinctisque lumbis, currebat ante Achab, donec veniret in Iezrahel.
1KGS|19|1|Nuntiavit autem Achab Iezabel omnia, quae fecerat Elias, et quomodo occidisset universos prophetas gladio.
1KGS|19|2|Misitque Iezabel nuntium ad Eliam dicens: " Haec mihi faciant dii et haec addant, nisi hac hora cras posuero animam tuam sicut animam unius ex illis ".
1KGS|19|3|Timuit ergo Elias et surgens abiit, ut animam suam salvaret, venitque in Bersabee Iudae et dimisit ibi puerum suum.
1KGS|19|4|Et perrexit in desertum via unius diei; cumque venisset et sederet subter unam iuniperum, petivit animae suae, ut moreretur, et ait: " Sufficit mihi, Domine! Tolle animam meam; neque enim melior sum quam patres mei ".
1KGS|19|5|Proiecitque se et obdormivit in umbra iuniperi; et ecce angelus tetigit eum et dixit illi: " Surge, comede! ".
1KGS|19|6|Respexit, et ecce ad caput suum subcinericius panis et vas aquae; comedit ergo et bibit et rursum obdormivit.
1KGS|19|7|Reversusque est angelus Domini secundo et tetigit eum dixitque illi: " Surge, comede! Grandis enim tibi restat via ".
1KGS|19|8|Qui, cum surrexisset, comedit et bibit et ambulavit in fortitudine cibi illius quadraginta diebus et quadraginta noctibus usque ad montem Dei Horeb.
1KGS|19|9|Cumque venisset illuc, mansit in spelunca. Et ecce sermo Domini ad eum dixitque illi: " Quid hic agis, Elia? ".
1KGS|19|10|At ille respondit: " Zelo zelatus sum pro Domino, Deo exercituum, quia dereliquerunt pactum tuum filii Israel, altaria tua destruxerunt et prophetas tuos occiderunt gladio; et derelictus sum ego solus, et quaerunt animam meam, ut auferant eam ".
1KGS|19|11|Et ait ei: " Egredere et sta in monte coram Domino ". Et ecce Dominus transit, et ventus grandis et fortis subvertens montes et conterens petras ante Dominum; non in vento Dominus. Et post ventum, commotio; non in commotione Dominus.
1KGS|19|12|Et post commotionem, ignis; non in igne Dominus. Et post ignem, sibilus aurae tenuis.
1KGS|19|13|Quod cum audisset Elias, operuit vultum suum pallio et egressus stetit in ostio speluncae; et ecce vox ad eum dicens: " Quid agis hic, Elia? ".
1KGS|19|14|Et ille respondit: " Zelo zelatus sum pro Domino, Deo exercituum, quia dereliquerunt pactum tuum filii Israel, altaria tua destruxerunt et prophetas tuos occiderunt gladio; et derelictus sum ego solus, et quaerunt animam meam, ut auferant eam ".
1KGS|19|15|Et ait Dominus ad eum: " Vade et revertere in viam tuam per desertum in Damascum. Cumque perveneris, unges Hazael regem super Syriam;
1KGS|19|16|et Iehu filium Namsi unges regem super Israel; Eliseum autem filium Saphat, qui est de Abelmehula, unges prophetam pro te.
1KGS|19|17|Et erit: quicumque fugerit gladium Hazael, occidet eum Iehu; et, qui fugerit gladium Iehu, interficiet eum Eliseus.
1KGS|19|18|Et relinquam mihi in Israel septem milia: universorum genua, quae non sunt incurvata ante Baal, et omne os, quod non osculatum est eum ".
1KGS|19|19|Profectus ergo inde repperit Eliseum filium Saphat arantem duodecim iugis boum; et ipse cum duodecimo erat. Cumque venisset Elias ad eum, misit pallium suum super illum,
1KGS|19|20|qui statim, relictis bobus, cucurrit post Eliam et ait: " Osculer, oro, patrem meum et matrem meam, et sic sequar te ". Dixitque ei: " Vade et revertere; quid enim feci tibi? ".
1KGS|19|21|Reversus autem ab eo tulit par boum et mactavit illud et in iugo boum coxit carnes et dedit populo, et comederunt. Consurgensque abiit et secutus est Eliam et ministrabat ei.
1KGS|20|1|Porro Benadad rex Syriae congregavit omnem exerci tum suum et triginta duos reges secum et equos et currus et ascendens pugnabat contra Samariam et obsidebat eam.
1KGS|20|2|Mittensque nuntios ad Achab regem Israel in civitatem
1KGS|20|3|ait: " Haec dicit Benadad: Argentum tuum et aurum tuum meum est, et uxores tuae et filii tui optimi mei sunt ".
1KGS|20|4|Responditque rex Israel: " Iuxta verbum tuum, domine mi rex; tuus sum ego et omnia mea ".
1KGS|20|5|Revertentesque nuntii dixerunt: " Haec dicit Benadad: Quia misi ad te dicens: "Argentum tuum et aurum tuum et uxores tuas et filios tuos dabis mihi",
1KGS|20|6|profecto cras hac eadem hora mittam servos meos ad te, et scrutabuntur domum tuam et domum servorum tuorum; et omne, quod oculis tuis pretiosum est, ponent in manibus suis et auferent ".
1KGS|20|7|Vocavit autem rex Israel omnes seniores terrae et ait: " Animadvertite et videte quoniam insidietur nobis; misit enim ad me pro uxoribus meis et filiis et pro argento et auro, et non abnui ".
1KGS|20|8|Dixeruntque omnes maiores natu et universus populus ad eum: " Non audias neque acquiescas illi ".
1KGS|20|9|Respondit itaque nuntiis Benadad: " Dicite domino meo regi: Omnia, propter quae misisti ad me servum tuum initio, faciam; hanc autem rem facere non possum ". Reversique nuntii rettulerunt ei.
1KGS|20|10|Qui remisit et ait: " Haec faciant mihi dii et haec addant, si suffecerit pulvis Samariae pugillis omnis populi, qui sequitur me ".
1KGS|20|11|Et respondens rex Israel ait: " Dicite ei: Ne glorietur accinctus aeque ut discinctus ".
1KGS|20|12|Factum est autem, cum audisset verbum istud, bibebat ipse et reges in umbraculis et ait servis suis: " Circumdate civitatem! ". Et circumdederunt eam.
1KGS|20|13|Et ecce propheta unus accedens ad Achab regem Israel ait: " Haec dicit Dominus: Certe vidisti omnem multitudinem hanc nimiam. Ecce ego tradam eam in manu tua hodie, ut scias quia ego sum Dominus ".
1KGS|20|14|Et ait Achab: " Per quem? ". Dixitque ei: " Haec dicit Dominus: Per pedisequos principum provinciarum ". Et ait: " Quis incipiet proeliari? ". Et ille dixit: " Tu ".
1KGS|20|15|Recensuit ergo pueros principum provinciarum et repperit numerum ducentorum triginta duorum; et post eos recensuit populum, omnes filios Israel, septem milia.
1KGS|20|16|Et egressi sunt meridie. Benadad autem bibebat temulentus in umbraculis ipse et reges triginta duo cum eo, qui ad auxilium eius venerant.
1KGS|20|17|Egressi sunt autem pueri principum provinciarum in prima fronte. Misit itaque Benadad, qui nuntiaverunt ei dicentes: " Viri egressi sunt de Samaria ".
1KGS|20|18|At ille ait: " Sive pro pace veniunt, apprehendite eos vivos; sive ut proelientur, vivos eos capite ".
1KGS|20|19|Egressi erant ergo ex urbe pueri principum provinciarum, ac reliquus exercitus sequebatur,
1KGS|20|20|et percussit unusquisque virum, qui contra se venerat; fugeruntque Syri, et persecutus est eos Israel. Fugit quoque Benadad rex Syriae in equo cum equitibus.
1KGS|20|21|Necnon egressus rex Israel percussit equos et currus et percussit Syriam plaga magna.
1KGS|20|22|Accedens autem propheta ad regem Israel dixit ei: " Vade et confortare et scito et vide quid facias; vertente enim anno rex Syriae ascendet contra te ".
1KGS|20|23|Servi vero regis Syriae dixerunt ei: " Deus montium est Deus eorum, ideo superaverunt nos; sed pugnemus contra eos in campestribus et obtinebimus eos.
1KGS|20|24|Fac ergo hoc: Amove reges singulos a loco suo et pone principes pro eis;
1KGS|20|25|et instaura numerum militum, qui ceciderunt de tuis, et equos secundum equos pristinos et currus secundum currus, quos ante habuisti, et pugnabimus contra eos in campestribus: et videbis quod obtinebimus eos ". Credidit consilio eorum et fecit ita.
1KGS|20|26|Igitur vertente anno recensuit Benadad Syros et ascendit in Aphec, ut pugnaret contra Israel.
1KGS|20|27|Porro filii Israel recensiti sunt et, acceptis cibariis, profecti ex adverso castraque metati sunt contra eos, quasi duo parvi greges caprarum; Syri autem repleverunt terram.
1KGS|20|28|Et accedens vir Dei dixit ad regem Israel: " Haec dicit Dominus: Quia dixerunt Syri: "Deus montium est Dominus et non est Deus vallium", dabo omnem multitudinem hanc grandem in manu tua, et scietis quia ego Dominus.
1KGS|20|29|Dirigebant septem diebus ex adverso hi atque illi acies, septima autem die commissum est bellum; percusseruntque filii Israel de Syris centum milia peditum in die una.
1KGS|20|30|Fugerunt autem, qui remanserant in Aphec, in civitatem, et cecidit murus super viginti septem milia hominum, qui remanserant.Porro Benadad fugiens ingressus est civitatem in cubiculum, quod erat intra cubiculum.
1KGS|20|31|Dixeruntque ei servi sui: " Ecce audivimus quod reges domus Israel clementes sint; ponamus itaque saccos in lumbis nostris et funiculos in capitibus nostris et egrediamur ad regem Israel; forsitan salvabit animam tuam ".
1KGS|20|32|Accinxerunt saccis lumbos suos et posuerunt funes in capitibus suis veneruntque ad regem Israel et dixerunt: " Servus tuus Benadad dicit: Vivat, oro te, anima mea" ". Et ille ait: " Si adhuc vivit, frater meus est ".
1KGS|20|33|Quod acceperunt viri pro omine et festinantes rapuerunt verbum ex ore eius atque dixerunt: " Frater tuus Benadad ". Et dixit eis: " Ite et adducite eum ". Egressus est ergo ad eum Benadad, et levavit eum in currum suum.
1KGS|20|34|Qui dixit ei: " Civitates, quas tulit pater meus a patre tuo, reddam; et plateas fac tibi in Damasco, sicut fecit pater meus in Samaria ". Achab: " Ego autem, inquit, foederatum te dimittam ". Et pepigit ei foedus et dimisit eum.
1KGS|20|35|Tunc vir quidam de filiis prophetarum dixit ad socium suum in sermone Domini: " Percute me! ". At ille noluit percutere.
1KGS|20|36|Cui ait: " Quia noluisti audire vocem Domini, ecce recedes a me, et percutiet te leo ". Cumque paululum recessisset ab eo, invenit eum leo atque percussit.
1KGS|20|37|Sed et alterum inveniens virum dixit ad eum: " Percute me! ". Qui percussit eum et vulneravit.
1KGS|20|38|Abiit ergo propheta et occurrit regi in via et mutavit aspectum ponens fasciam super oculos suos.
1KGS|20|39|Cumque rex transiret, clamavit ad regem et ait: " Servus tuus egressus est ad proeliandum comminus; cumque fugisset vir unus, adduxit eum quidam ad me et ait: "Custodi virum istum! Qui si lapsus fuerit, erit anima tua pro anima eius, aut talentum argenti appendes".
1KGS|20|40|Dum autem ego turbatus huc illucque me verterem, subito non comparuit. Et ait rex Israel ad eum: " Hoc est iudicium tuum, quod ipse decrevisti.
1KGS|20|41|At ille statim abstulit fasciam de oculis suis, et cognovit eum rex Israel quod esset de prophetis.
1KGS|20|42|Qui ait ad eum: " Haec dicit Dominus: Quia dimisisti de manu tua virum, quem morti devoveram, erit anima tua pro anima eius, et populus tuus pro populo eius ".
1KGS|20|43|Reversus est igitur rex Israel in domum suam tristis et indignans venitque in Samariam.
1KGS|21|1|Postea autem factum est hoc. Vinea erat Naboth Iez rahelitae, quae erat in Iezrahel iuxta palatium Achab regis Samariae.
1KGS|21|2|Locutus est ergo Achab ad Naboth dicens: " Da mihi vineam tuam, ut faciam mihi hortum holerum, quia vicina est et prope domum meam. Daboque tibi pro ea vineam meliorem aut, si tibi commodius putas, argenti pretium quanto digna est ".
1KGS|21|3|Cui respondit Naboth: " Propitius mihi sit Dominus, ne dem hereditatem patrum meorum tibi ".
1KGS|21|4|Venit ergo Achab in domum suam tristis et indignans super verbo, quod locutus fuerat ad eum Naboth Iezrahelites dicens: " Non dabo tibi hereditatem patrum meorum ". Et proiciens se in lectulum suum avertit faciem ad parietem et non comedit panem.
1KGS|21|5|Ingressa est autem ad eum Iezabel uxor sua dixitque ei: " Quid est hoc, unde anima tua contristata est? Et quare non comedis panem? ".
1KGS|21|6|Qui respondit ei: " Quia locutus sum Naboth Iezrahelitae et dixi ei: Da mihi vineam tuam, accepta pecunia; aut, si tibi placet, dabo tibi vineam pro ea. Et ille ait: "Non dabo tibi vineam meam" ".
1KGS|21|7|Dixit ergo ad eum Iezabel uxor eius: " Grandis auctoritatis es et bene regis regnum Israel! Surge et comede panem et aequo esto animo; ego dabo tibi vineam Naboth Iezrahelitae ".
1KGS|21|8|Scripsit itaque litteras ex nomine Achab et signavit eas anulo eius et misit ad maiores natu et ad optimates, qui erant in civitate eius et habitabant cum Naboth.
1KGS|21|9|Litterarum autem haec erat sententia: " Praedicate ieiunium et sedere facite Naboth in capite populi
1KGS|21|10|et submittite duos viros filios Belial contra eum, et testimonium dicant: "Maledixisti Deum et regem"; et educite eum et lapidate, sicque moriatur ".
1KGS|21|11|Fecerunt ergo cives eius maiores natu et optimates, qui habitabant cum eo in urbe, sicut praeceperat eis Iezabel et sicut scriptum erat in litteris, quas miserat ad eos.
1KGS|21|12|Praedicaverunt ieiunium et sedere fecerunt Naboth in capite populi;
1KGS|21|13|et ingressi duo viri filii Belial sederunt contra eum et illi, ut viri diabolici, dixerunt contra eum testimonium coram multitudine: " Maledixit Naboth Deum et regem ". Quam ob rem eduxerunt eum extra civitatem et lapidibus interfecerunt;
1KGS|21|14|miseruntque ad Iezabel dicentes: " Lapidatus est Naboth et mortuus est.
1KGS|21|15|Factum est autem cum audisset Iezabel lapidatum Naboth et mortuum, locuta est ad Achab: " Surge, posside vineam Naboth Iezrahelitae, qui noluit tibi acquiescere et dare eam, accepta pecunia; non enim vivit Naboth, sed mortuus est ".
1KGS|21|16|Quod cum audisset Achab, mortuum videlicet Naboth, surrexit et descendebat in vineam Naboth Iezrahelitae, ut possideret eam.
1KGS|21|17|Factus est igitur sermo Domini ad Eliam Thesbiten dicens:
1KGS|21|18|" Surge et descende in occursum Achab regis Israel, qui est in Samaria; ecce est in vinea Naboth, ad quam descendit, ut possideat eam.
1KGS|21|19|Et loqueris ad eum dicens: Haec dicit Dominus: Occidisti, insuper et possedisti! Et post haec addes: Haec dicit Dominus: In loco, in quo linxerunt canes sanguinem Naboth, lambent tuum quoque sanguinem ".
1KGS|21|20|Et ait Achab ad Eliam: " Num invenisti me, inimice mi? ". Qui dixit: " Inveni, eo quod venumdatus sis, ut faceres malum in conspectu Domini.
1KGS|21|21|Ecce ego inducam super te malum et demetam posteriora tua et interficiam de Achab quidquid masculini sexus sive impuberem sive puberem in Israel.
1KGS|21|22|Et dabo domum tuam sicut domum Ieroboam filii Nabat et sicut domum Baasa filii Ahia, quia egisti, ut me ad iracundiam provocares, et peccare fecisti Israel.
1KGS|21|23|Sed et de Iezabel locutus est Dominus dicens: Canes comedent Iezabel in agro Iezrahel.
1KGS|21|24|Qui de Achab mortuus fuerit in civitate, comedent eum canes; qui autem mortuus fuerit in agro, comedent eum volucres caeli ".
1KGS|21|25|Igitur non fuit alter talis sicut Achab, qui venumdatus est, ut faceret malum in conspectu Domini; concitavit enim eum Iezabel uxor sua,
1KGS|21|26|et abominabilis effectus est, in tantum ut sequeretur idola secundum omnia, quae fecerant Amorraei, quos consumpsit Dominus a facie filiorum Israel.
1KGS|21|27|Itaque cum audisset Achab sermones istos, scidit vestem suam et operuit cilicio carnem suam ieiunavitque et dormivit in sacco et ambulabat demisso capite.
1KGS|21|28|Factus est autem sermo Domini ad Eliam Thesbiten dicens:
1KGS|21|29|Nonne vidisti humiliatum Achab coram me? Quia igitur humiliatus est mei causa, non inducam malum in diebus eius, sed in diebus filii sui inferam malum domui eius ".
1KGS|22|1|Transierunt igitur tres anni absque bello inter Syriam et Israel.
1KGS|22|2|In anno autem tertio descendit Iosaphat rex ludae ad regem Israel,
1KGS|22|3|dixitque rex Israel ad servos suos: " Ignoratis quod nostra sit Ramoth Galaad et neglegimus tollere eam de manu regis Syriae? ".
1KGS|22|4|Et ait ad Iosaphat: " Veniesne mecum ad proeliandum in Ramoth Galaad? ".
1KGS|22|5|Dixitque Iosaphat ad regem Israel: " Sicut ego sum, ita et tu; populus meus et populus tuus unum sunt, et equites mei et equites tui ". Dixitque Iosaphat ad regem Israel: " Quaere, oro te, hodie sermonem Domini ".
1KGS|22|6|Congregavit ergo rex Israel prophetas quadringentos circiter viros et ait ad eos: " Ire debeo in Ramoth Galaad ad bellandum, an quiescere? ". Qui responderunt: " Ascende, et dabit Dominus in manu regis ".
1KGS|22|7|Dixit autem Iosaphat: " Non est hic et alius propheta Domini, ut interrogemus per eum? ".
1KGS|22|8|Et ait rex Israel ad Iosaphat: " Remansit vir unus, per quem possimus interrogare Dominum; sed ego odi eum, quia non prophetat mihi bonum sed malum: Michaeas filius Iemla ". Cui Iosaphat ait: " Ne loquaris ita, rex.
1KGS|22|9|Vocavit ergo rex Israel eunuchum quendam et dixit ei: " Festina adducere Michaeam filium Iemla ".
1KGS|22|10|Rex autem Israel et Iosaphat rex Iudae sedebat unusquisque in solio suo vestiti cultu regio in area iuxta ostium portae Samariae; et universi prophetae prophetabant in conspectu eorum.
1KGS|22|11|Fecit quoque sibi Sedecias filius Chanaana cornua ferrea et ait: " Haec dicit Dominus: His ventilabis Syriam, donec deleas eam ".
1KGS|22|12|Omnesque prophetae similiter prophetabant dicentes: " Ascende in Ramoth Galaad et vade prospere, et tradet Dominus in manu regis ".
1KGS|22|13|Nuntius vero, qui ierat ut vocaret Michaeam, locutus est ad eum dicens: Ecce sermones prophetarum ore uno regi bona praedicant; sit ergo sermo tuus similis eorum, et loquere bona ".
1KGS|22|14|Cui Michaeas ait: " Vivit Dominus quia, quodcumque dixerit mihi Dominus, hoc loquar! ".
1KGS|22|15|Venit itaque ad regem, et ait illi rex: " Michaea, ire debemus in Ramoth Galaad ad proeliandum, an cessare? ". Cui ille respondit: " Ascende et vade prospere, et tradet Dominus in manu regis ".
1KGS|22|16|Dixit autem rex ad eum: " Iterum atque iterum adiuro te, ut non loquaris mihi, nisi quod verum est in nomine Domini ".
1KGS|22|17|Et ille ait: Vidi cunctum Israeldispersum in montibusquasi oves non habentes pastorem. Et ait Dominus: "Non habent isti dominum; revertatur unusquisque in domum suam in pace" ".
1KGS|22|18|Dixit ergo rex Israel ad Iosaphat: " Numquid non dixi tibi quia non prophetat mihi bonum sed semper malum? ".
1KGS|22|19|Ille vero addens ait: " Propterea audi sermonem Domini: Vidi Dominum sedentem super solium suum et omnem exercitum caeli assistentem ei a dextris et a sinistris.
1KGS|22|20|Et ait Dominus: "Quis decipiet Achab, ut ascendat et cadat in Ramoth Galaad?". Et dixit unus verba huiuscemodi et alius aliter.
1KGS|22|21|Egressus est autem spiritus et stetit coram Domino et ait: "Ego decipiam illum". Cui locutus est Dominus: "In quo?".
1KGS|22|22|Et ille ait: "Egrediar et ero spiritus mendax in ore omnium prophetarum eius". Et dixit Dominus: "Decipies et praevalebis; egredere et fac ita".
1KGS|22|23|Nunc igitur ecce dedit Dominus spiritum mendacii in ore omnium prophetarum tuorum, qui hic sunt, et Dominus locutus est contra te malum.
1KGS|22|24|Accessit autem Sedecias filius Chanaana et percussit Michaeam in maxillam et dixit: " Quomodo transivit spiritus Domini a me, ut loqueretur tibi? ".
1KGS|22|25|Et ait Michaeas: " Visurus es in die illa, quando ingredieris cubiculum intra cubiculum, ut abscondaris ".
1KGS|22|26|Et ait rex Israel: " Tolle Michaeam, et maneat apud Amon principem civitatis et apud Ioas filium regis,
1KGS|22|27|et dic eis: "Haec dicit rex: Mittite virum istum in carcerem et sustentate eum pane tribulationis et aqua angustiae, donec revertar in pace" ".
1KGS|22|28|Dixitque Michaeas: " Si reversus fueris in pace, non est locutus Dominus in me ". Et ait: " Audite, populi omnes! ".
1KGS|22|29|Ascendit itaque rex Israel et Iosaphat rex Iudae in Ramoth Galaad.
1KGS|22|30|Dixitque rex Israel ad Iosaphat: " Mutato aspectu ineundum est proelium; tu autem induere vestibus tuis ". Porro rex Israel mutavit aspectum et ingressus est bellum.
1KGS|22|31|Rex autem Syriae praeceperat principibus curruum triginta duobus dicens: " Non pugnabitis contra minorem et maiorem quempiam, nisi contra regem Israel solum ".
1KGS|22|32|Cum ergo vidissent principes curruum Iosaphat, suspicati sunt quod ipse esset rex Israel et impetu facto pugnabant contra eum. Et exclamavit Iosaphat;
1KGS|22|33|intellexeruntque principes curruum quod non esset rex Israel et cessaverunt ab eo.
1KGS|22|34|Vir autem quidam tetendit arcum in incertum sagittam dirigens et percussit regem Israel inter iuncturas et loricam. At ille dixit aurigae suo: " Verte manum tuam et eice me de exercitu, quia graviter vulneratus sum ".
1KGS|22|35|Aggravatum est ergo proelium in die illa; et rex Israel stabat in curru suo contra Syros et mortuus est vespere: fluebat autem sanguis plagae in sinum currus.
1KGS|22|36|Et clamor insonuit in universo exercitu ad solis occasum: " Unusquisque revertatur in civitatem et in terram suam! ".
1KGS|22|37|Mortuus est igitur rex et perlatus est Samariam; sepelieruntque regem in Samaria.
1KGS|22|38|Et laverunt currum eius in piscina Samariae; et linxerunt canes sanguinem eius, et scorta laverunt se iuxta verbum Domini, quod locutus fuerat.
1KGS|22|39|Reliqua vero gestorum Achab et universa, quae fecit, et domus eburnea, quam aedificavit, cunctaeque urbes, quas exstruxit, nonne haec scripta sunt in libro annalium regum Israel?
1KGS|22|40|Dormivit ergo Achab cum patribus suis; et regnavit Ochozias filius eius pro eo.
1KGS|22|41|Iosaphat vero filius Asa regnare coeperat super Iudam anno quarto Achab regis Israel;
1KGS|22|42|triginta quinque annorum erat, cum regnare coepisset, et viginti quinque annos regnavit in Ierusalem. Nomen matris eius Azuba filia Selachi.
1KGS|22|43|Et ambulavit in omni via Asa patris sui et non declinavit ex ea; fecitque, quod rectum erat in conspectu Domini.
1KGS|22|44|Verumtamen excelsa non abstulit; adhuc enim populus sacrificabat et adolebat in excelsis.
1KGS|22|45|Pacemque fecit Iosaphat cum rege Israel.
1KGS|22|46|Reliqua autem gestorum Iosaphat et opera eius, quae fortiter gessit, et proelia, nonne haec scripta sunt in libro annalium regum Iudae?
1KGS|22|47|Sed et reliquias prostibulorum, qui remanserant in diebus Asa patris eius, abstulit de terra.
1KGS|22|48|Nec erat tunc rex in Edom sed praefectus regius.
1KGS|22|49|Rex vero Iosaphat fecerat naves Tharsis, quae navigarent in Ophir propter aurum; et ire non potuerunt, quia confractae sunt in Asiongaber.
1KGS|22|50|Tunc ait Ochozias filius Achab ad Iosaphat: " Vadant servi mei cum servis tuis in navibus ". Et noluit Iosaphat.
1KGS|22|51|Dormivitque Iosaphat cum patribus suis et sepultus est cum eis in civitate David patris sui; regnavitque Ioram filius eius pro eo.
1KGS|22|52|Ochozias autem filius Achab regnare coeperat super Israel in Samaria anno septimo decimo Iosaphat regis Iudae regnavitque super Israel duobus annis.
1KGS|22|53|Et fecit malum in conspectu Domini et ambulavit in via patris sui et matris suae et in via Ieroboam filii Nabat, qui peccare fecit Israel;
1KGS|22|54|servivit quoque Baal et adoravit eum et irritavit Dominum, Deum Israel, iuxta omnia, quae fecerat pater eius.
