MIC|1|1|The word of the LORD that came to Micah of Moresheth in the days of Jotham, Ahaz, and Hezekiah, kings of Judah, which he saw concerning Samaria and Jerusalem.
MIC|1|2|Hear, you peoples, all of you; pay attention, O earth, and all that is in it, and let the Lord GOD be a witness against you, the Lord from his holy temple.
MIC|1|3|For behold, the LORD is coming out of his place, and will come down and tread upon the high places of the earth.
MIC|1|4|And the mountains will melt under him, and the valleys will split open, like wax before the fire, like waters poured down a steep place.
MIC|1|5|All this is for the transgression of Jacob and for the sins of the house of Israel. What is the transgression of Jacob? Is it not Samaria? And what is the high place of Judah? Is it not Jerusalem?
MIC|1|6|Therefore I will make Samaria a heap in the open country, a place for planting vineyards, and I will pour down her stones into the valley and uncover her foundations.
MIC|1|7|All her carved images shall be beaten to pieces, all her wages shall be burned with fire, and all her idols I will lay waste, for from the fee of a prostitute she gathered them, and to the fee of a prostitute they shall return.
MIC|1|8|For this I will lament and wail; I will go stripped and naked; I will make lamentation like the jackals, and mourning like the ostriches.
MIC|1|9|For her wound is incurable, and it has come to Judah; it has reached to the gate of my people, to Jerusalem.
MIC|1|10|Tell it not in Gath; weep not at all; in Beth-le-aphrah roll yourselves in the dust.
MIC|1|11|Pass on your way, inhabitants of Shaphir, in nakedness and shame; the inhabitants of Zaanan do not come out; the lamentation of Beth-ezel shall take away from you its standing place.
MIC|1|12|For the inhabitants of Maroth wait anxiously for good, because disaster has come down from the LORD to the gate of Jerusalem.
MIC|1|13|Harness the steeds to the chariots, inhabitants of Lachish; it was the beginning of sin to the daughter of Zion, for in you were found the transgressions of Israel.
MIC|1|14|Therefore you shall give parting gifts to Moresheth-gath; the houses of Achzib shall be a deceitful thing to the kings of Israel.
MIC|1|15|I will again bring a conqueror to you, inhabitants of Mareshah; the glory of Israel shall come to Adullam.
MIC|1|16|Make yourselves bald and cut off your hair, for the children of your delight; make yourselves as bald as the eagle, for they shall go from you into exile.
MIC|2|1|Woe to those who devise wickedness and work evil on their beds! When the morning dawns, they perform it, because it is in the power of their hand.
MIC|2|2|They covet fields and seize them, and houses, and take them away; they oppress a man and his house, a man and his inheritance.
MIC|2|3|Therefore thus says the LORD: behold, against this family I am devising disaster, from which you cannot remove your necks, and you shall not walk haughtily, for it will be a time of disaster.
MIC|2|4|In that day they shall take up a taunt song against you and moan bitterly, and say, "We are utterly ruined; he changes the portion of my people; how he removes it from me! To an apostate he allots our fields."
MIC|2|5|Therefore you will have none to cast the line by lot in the assembly of the LORD.
MIC|2|6|"Do not preach"- thus they preach- "one should not preach of such things; disgrace will not overtake us."
MIC|2|7|Should this be said, O house of Jacob? Has the LORD grown impatient? Are these his deeds? Do not my words do good to him who walks uprightly?
MIC|2|8|But lately my people have risen up as an enemy; you strip the rich robe from those who pass by trustingly with no thought of war.
MIC|2|9|The women of my people you drive out from their delightful houses; from their young children you take away my splendor forever.
MIC|2|10|Arise and go, for this is no place to rest, because of uncleanness that destroys with a grievous destruction.
MIC|2|11|If a man should go about and utter wind and lies, saying, "I will preach to you of wine and strong drink," he would be the preacher for this people!
MIC|2|12|I will surely assemble all of you, O Jacob; I will gather the remnant of Israel; I will set them together like sheep in a fold, like a flock in its pasture, a noisy multitude of men.
MIC|2|13|He who opens the breach goes up before them; they break through and pass the gate, going out by it. Their king passes on before them, the LORD at their head.
MIC|3|1|And I said:Hear, you heads of Jacob and rulers of the house of Israel! Is it not for you to know justice?-
MIC|3|2|you who hate the good and love the evil, who tear the skin from off my people and their flesh from off their bones,
MIC|3|3|who eat the flesh of my people, and flay their skin from off them, and break their bones in pieces and chop them up like meat in a pot, like flesh in a cauldron.
MIC|3|4|Then they will cry to the LORD, but he will not answer them; he will hide his face from them at that time, because they have made their deeds evil.
MIC|3|5|Thus says the LORD concerning the prophets who lead my people astray, who cry "Peace" when they have something to eat, but declare war against him who puts nothing into their mouths.
MIC|3|6|Therefore it shall be night to you, without vision, and darkness to you, without divination. The sun shall go down on the prophets, and the day shall be black over them;
MIC|3|7|the seers shall be disgraced, and the diviners put to shame; they shall all cover their lips, for there is no answer from God.
MIC|3|8|But as for me, I am filled with power, with the Spirit of the LORD, and with justice and might, to declare to Jacob his transgression and to Israel his sin.
MIC|3|9|Hear this, you heads of the house of Jacob and rulers of the house of Israel, who detest justice and make crooked all that is straight,
MIC|3|10|who build Zion with blood and Jerusalem with iniquity.
MIC|3|11|Its heads give judgment for a bribe; its priests teach for a price; its prophets practice divination for money; yet they lean on the LORD and say, "Is not the LORD in the midst of us? No disaster shall come upon us."
MIC|3|12|Therefore because of you Zion shall be plowed as a field; Jerusalem shall become a heap of ruins, and the mountain of the house a wooded height.
MIC|4|1|It shall come to pass in the latter days that the mountain of the house of the LORD shall be established as the highest of the mountains, and it shall be lifted up above the hills; and peoples shall flow to it,
MIC|4|2|and many nations shall come, and say: "Come, let us go up to the mountain of the LORD, to the house of the God of Jacob, that he may teach us his ways and that we may walk in his paths." For out of Zion shall go forth the law, and the word of the LORD from Jerusalem.
MIC|4|3|He shall judge between many peoples, and shall decide for strong nations afar off; and they shall beat their swords into plowshares, and their spears into pruning hooks; nation shall not lift up sword against nation, neither shall they learn war anymore;
MIC|4|4|but they shall sit every man under his vine and under his fig tree, and no one shall make them afraid, for the mouth of the LORD of hosts has spoken.
MIC|4|5|For all the peoples walk each in the name of its god, but we will walk in the name of the LORD our God forever and ever.
MIC|4|6|In that day, declares the LORD, I will assemble the lame and gather those who have been driven away and those whom I have afflicted;
MIC|4|7|and the lame I will make the remnant, and those who were cast off, a strong nation; and the LORD will reign over them in Mount Zion from this time forth and forevermore.
MIC|4|8|And you, O tower of the flock, hill of the daughter of Zion, to you shall it come, the former dominion shall come, kingship for the daughter of Jerusalem.
MIC|4|9|Now why do you cry aloud? Is there no king in you? Has your counselor perished, that pain seized you like a woman in labor?
MIC|4|10|Writhe and groan, O daughter of Zion, like a woman in labor, for now you shall go out from the city and dwell in the open country; you shall go to Babylon. There you shall be rescued; there the LORD will redeem you from the hand of your enemies.
MIC|4|11|Now many nations are assembled against you, saying, "Let her be defiled, and let our eyes gaze upon Zion."
MIC|4|12|But they do not know the thoughts of the LORD; they do not understand his plan, that he has gathered them as sheaves to the threshing floor.
MIC|4|13|Arise and thresh, O daughter of Zion, for I will make your horn iron, and I will make your hoofs bronze; you shall beat in pieces many peoples; and shall devote their gain to the LORD, their wealth to the Lord of the whole earth.
MIC|5|1|Now muster your troops, O daughter of troops; siege is laid against us; with a rod they strike the judge of Israel on the cheek.
MIC|5|2|But you, O Bethlehem Ephrathah, who are too little to be among the clans of Judah, from you shall come forth for me one who is to be ruler in Israel, whose origin is from of old, from ancient days.
MIC|5|3|Therefore he shall give them up until the time when she who is in labor has given birth; then the rest of his brothers shall return to the people of Israel.
MIC|5|4|And he shall stand and shepherd his flock in the strength of the LORD, in the majesty of the name of the LORD his God. And they shall dwell secure, for now he shall be great to the ends of the earth.
MIC|5|5|And he shall be their peace. When the Assyrian comes into our land and treads in our palaces, then we will raise against him seven shepherds and eight princes of men;
MIC|5|6|they shall shepherd the land of Assyria with the sword, and the land of Nimrod at its entrances; and he shall deliver us from the Assyrian when he comes into our land and treads within our border.
MIC|5|7|Then the remnant of Jacob shall be in the midst of many peoples like dew from the LORD, like showers on the grass, which delay not for a man nor wait for the children of man.
MIC|5|8|And the remnant of Jacob shall be among the nations, in the midst of many peoples, like a lion among the beasts of the forest, like a young lion among the flocks of sheep, which, when it goes through, treads down and tears in pieces, and there is none to deliver.
MIC|5|9|Your hand shall be lifted up over your adversaries, and all your enemies shall be cut off.
MIC|5|10|And in that day, declares the LORD, I will cut off your horses from among you and will destroy your chariots;
MIC|5|11|and I will cut off the cities of your land and throw down all your strongholds;
MIC|5|12|and I will cut off sorceries from your hand, and you shall have no more tellers of fortunes;
MIC|5|13|and I will cut off your carved images and your pillars from among you, and you shall bow down no more to the work of your hands;
MIC|5|14|and I will root out your Asherah images from among you and destroy your cities.
MIC|5|15|And in anger and wrath I will execute vengeance on the nations that did not obey.
MIC|6|1|Hear what the LORD says:Arise, plead your case before the mountains, and let the hills hear your voice.
MIC|6|2|Hear, you mountains, the indictment of the LORD, and you enduring foundations of the earth, for the LORD has an indictment against his people, and he will contend with Israel.
MIC|6|3|"O my people, what have I done to you? How have I wearied you? Answer me!
MIC|6|4|For I brought you up from the land of Egypt and redeemed you from the house of slavery, and I sent before you Moses, Aaron, and Miriam.
MIC|6|5|O my people, remember what Balak king of Moab devised, and what Balaam the son of Beor answered him, and what happened from Shittim to Gilgal, that you may know the saving acts of the LORD."
MIC|6|6|"With what shall I come before the LORD, and bow myself before God on high? Shall I come before him with burnt offerings, with calves a year old?
MIC|6|7|Will the LORD be pleased with thousands of rams, with ten thousands of rivers of oil? Shall I give my firstborn for my transgression, the fruit of my body for the sin of my soul?"
MIC|6|8|He has told you, O man, what is good; and what does the LORD require of you but to do justice, and to love kindness, and to walk humbly with your God?
MIC|6|9|The voice of the LORD cries to the city- and it is sound wisdom to fear your name: "Hear of the rod and of him who appointed it!
MIC|6|10|Can I forget any longer the treasures of wickedness in the house of the wicked, and the scant measure that is accursed?
MIC|6|11|Shall I acquit the man with wicked scales and with a bag of deceitful weights?
MIC|6|12|Your rich men are full of violence; your inhabitants speak lies, and their tongue is deceitful in their mouth.
MIC|6|13|Therefore I strike you with a grievous blow, making you desolate because of your sins.
MIC|6|14|You shall eat, but not be satisfied, and there shall be hunger within you; you shall put away, but not preserve, and what you preserve I will give to the sword.
MIC|6|15|You shall sow, but not reap; you shall tread olives, but not anoint yourselves with oil; you shall tread grapes, but not drink wine.
MIC|6|16|For you have kept the statutes of Omri, and all the works of the house of Ahab; and you have walked in their counsels, that I may make you a desolation, and your inhabitants a hissing; so you shall bear the scorn of my people."
MIC|7|1|Woe is me! For I have become as when the summer fruit has been gathered, as when the grapes have been gleaned: there is no cluster to eat, no first-ripe fig that my soul desires.
MIC|7|2|The godly has perished from the earth, and there is no one upright among mankind; they all lie in wait for blood, and each hunts the other with a net.
MIC|7|3|Their hands are on what is evil, to do it well; the prince and the judge ask for a bribe, and the great man utters the evil desire of his soul; thus they weave it together.
MIC|7|4|The best of them is like a brier, the most upright of them a thorn hedge. The day of your watchmen, of your punishment, has come; now their confusion is at hand.
MIC|7|5|Put no trust in a neighbor; have no confidence in a friend; guard the doors of your mouth from her who lies in your arms;
MIC|7|6|for the son treats the father with contempt, the daughter rises up against her mother, the daughter-in-law against her mother-in-law; a man's enemies are the men of his own house.
MIC|7|7|But as for me, I will look to the LORD; I will wait for the God of my salvation; my God will hear me.
MIC|7|8|Rejoice not over me, O my enemy; when I fall, I shall rise; when I sit in darkness, the LORD will be a light to me.
MIC|7|9|I will bear the indignation of the LORD because I have sinned against him, until he pleads my cause and executes judgment for me. He will bring me out to the light; I shall look upon his vindication.
MIC|7|10|Then my enemy will see, and shame will cover her who said to me, "Where is the LORD your God?" My eyes will look upon her; now she will be trampled down like the mire of the streets.
MIC|7|11|A day for the building of your walls! In that day the boundary shall be far extended.
MIC|7|12|In that day they will come to you, from Assyria and the cities of Egypt, and from Egypt to the River, from sea to sea and from mountain to mountain.
MIC|7|13|But the earth will be desolate because of its inhabitants, for the fruit of their deeds.
MIC|7|14|Shepherd your people with your staff, the flock of your inheritance, who dwell alone in a forest in the midst of a garden land; let them graze in Bashan and Gilead as in the days of old.
MIC|7|15|As in the days when you came out of the land of Egypt, I will show them marvelous things.
MIC|7|16|The nations shall see and be ashamed of all their might; they shall lay their hands on their mouths; their ears shall be deaf;
MIC|7|17|they shall lick the dust like a serpent, like the crawling things of the earth; they shall come trembling out of their strongholds; they shall turn in dread to the LORD our God, and they shall be in fear of you.
MIC|7|18|Who is a God like you, pardoning iniquity and passing over transgression for the remnant of his inheritance? He does not retain his anger forever, because he delights in steadfast love.
MIC|7|19|He will again have compassion on us; he will tread our iniquities under foot. You will cast all our sins into the depths of the sea.
MIC|7|20|You will show faithfulness to Jacob and steadfast love to Abraham, as you have sworn to our fathers from the days of old.
