2CHR|1|1|І зміцнився Соломон, син Давидів, над царством своїм, а Господь, Бог його, був із ним та високо звеличив його.
2CHR|1|2|І сказав Соломон до всього Ізраїля, до тисячників та сотників, і до суддів, і до всіх начальників, до всього Ізраїля, до голів батьківських родів.
2CHR|1|3|І пішли Соломон та ввесь збір із ним до пагірка, що в Ґів'оні, бо там була скинія Божого заповіту, яку зробив Мойсей, раб Господній, у пустині.
2CHR|1|4|Але Божого ковчега Давид переніс із Кір'ят-Єаріму туди, де приготовив йому місце Давид, бо він поставив йому скинію в Єрусалимі.
2CHR|1|5|А мідяного жертівника, що зробив був Веселіїл, син Урії, сина Хурового, він поставив перед скинією Господньою. І звертався до нього Соломон та збір.
2CHR|1|6|І зійшов Соломон туди перед Господнє лице на мідяний жертівник, що належав до скинії заповіту, і приніс на ньому тисячу цілопалень.
2CHR|1|7|Тієї ночі явився Бог Соломонові та й сказав йому: Зажадай, чого дати тобі!
2CHR|1|8|І сказав Соломон до Бога: Ти зробив був велику милість з батьком моїм Давидом, і настановив царем мене замість нього.
2CHR|1|9|Тепер, Господи, Боже, нехай буде виповнене слово Твоє до батька мого Давида, бо Ти настановив мене царем над народом численним, як порох землі.
2CHR|1|10|Дай тепер мені мудрість та знання, щоб умів я виходити й входити перед цим народом, бо хто зможе судити цей великий Твій народ?
2CHR|1|11|І сказав Бог до Соломона: За те, що оце було на серці твоїм, і ти не жадав багатства, маєтків та слави, ані душі ворогів своїх, а також довгих днів не жадав ти, а жадав для себе мудрости та знання, щоб судити народ Мій, над яким Я настановив тебе царем,
2CHR|1|12|то дасться тобі мудрість та знання, а багатство, і маєтки та славу Я дам тобі такі, яких не було між царями перед тобою, і по тобі не буде таких!
2CHR|1|13|І прийшов Соломон із пагірка, що в Ґів'оні, до Єрусалиму, від скинії заповіту, і зацарював над Ізраїлем.
2CHR|1|14|І зібрав Соломон колесниць та верхівців, і було в нього тисяча й чотири сотні колесниць та дванадцять тисяч верхівців, і він порозміщував їх по колесничних містах та при царі в Єрусалимі.
2CHR|1|15|І цар зібрав в Єрусалимі срібла та золота, мов каміння, а кедрів зібрав, щодо численности, як сикомор, що в Шефелі.
2CHR|1|16|А коней, що були в Соломона, приводили з Єгипту та з Кеве; царські купці купували їх з Кеве.
2CHR|1|17|І ходили вони, і вивозили з Єгипту колесницю за шість сотень срібла, а коня за сотню й п'ятдесят. І так вони вивозили все це своєю рукою для всіх царів хіттійських та царів сирійських.
2CHR|2|1|(1-18) І Соломон наказав будувати дім для Господнього Ймення та дім царський для себе.
2CHR|2|2|(2-1) І відлічив Соломон сімдесят тисяч чоловіка носіїв та вісімдесят тисяч чоловіка каменотесів у горах, а керівників над ними три тисячі й шість сотень.
2CHR|2|3|(2-2) І послав Соломон до Хірама, царя тирського, говорячи: Як зробив ти з батьком моїм Давидом, і послав був йому кедри на будову дому його, щоб сидіти в ньому, так зроби й мені.
2CHR|2|4|(2-3) Ось я будую храм для Ймення Господа, Бога мого, щоб присвятити Йому, щоб кадити перед Його лицем запашне кадило, і для постійного покладення хліба та для цілопалення на ранок і на вечір, на суботи й на молодики та на свята Господа, Бога нашого. Навіки це над Ізраїлем!
2CHR|2|5|(2-4) А храм, якого я будую, великий, бо Бог наш більший від усіх богів!
2CHR|2|6|(2-5) А хто має силу збудувати Йому храма, коли небо й небеса небес не обіймають Його? І хто я, що збудую Йому храма? Хіба тільки на кадіння перед лицем Його!
2CHR|2|7|(2-6) А тепер пошли мені чоловіка, здібного до роботи в золоті, і в сріблі, і в міді, і в залізі, і в пурпурі, і в червені, і в блакиті, і що вміє вирізувати різьби, разом із тими мистцями, що зо мною в Юді та в Єрусалимі, яких приготовив батько мій Давид.
2CHR|2|8|(2-7) І пошли мені з Ливану дерева кедрового, кипарисового та сандалового, бо я знаю, що твої раби вміють рубати дерева ливанські. І оце мої раби будуть рабами твоїми,
2CHR|2|9|(2-8) щоб наготовити мені безліч дерева, бо цей храм, що я будую, буде великий та пишний!
2CHR|2|10|(2-9) А ось дереворубам, що стинають дерева, рабам твоїм, дав я пшениці, як поживи, двадцять тисяч корів, та ячменю двадцять тисяч корів, і вина двадцять тисяч батів, і оливи двадцять тисяч батів.
2CHR|2|11|(2-10) І сказав Хірам, цар тирський, листом і послав до Соломона: Через любов Господа до народу Свого поставив Він тебе над ними за царя.
2CHR|2|12|(2-11) І сказав Хірам: Благословенний Господь, Бог Ізраїлів, що вчинив небеса та землю, що дав цареві Давидові сина мудрого, який має розум та багатий на знання, що збудує дім Господній та дім царський для себе!
2CHR|2|13|(2-12) А тепер я посилаю мудрого чоловіка, що має знання, Хурам-Аві,
2CHR|2|14|(2-13) сина жінки з Данових дочок, а батько його тирянин, що вміє робити в золоті та в сріблі, в міді, в залізі, в каміннях та в деревах, у пурпурі й у блакиті, і в віссоні, і в червені, і різати всяку різьбу, і виконувати всяку думку, що буде дана йому з мистцями твоїми та з мистцями пана мого Давида, батька твого.
2CHR|2|15|(2-14) А тепер пшеницю й ячмінь, оливу та вино, про які казав мій пан, нехай посилає своїм рабам.
2CHR|2|16|(2-15) А ми нарубаємо дерев із Ливану за всякою твоєю потребою, і спровадимо їх тобі плотами морем до Яфи, а ти спровадиш їх до Єрусалиму.
2CHR|2|17|(2-16) І перелічив Соломон усіх людей приходьків, що в Ізраїлевому Краї, за переліком, що перелічив був їх його батько Давид, і було знайдено їх сто й п'ятдесят тисяч і три тисячі й шість сотень.
2CHR|2|18|(2-17) І він зробив із них сімдесят тисяч носіїв та вісімдесят тисяч каменотесів у горах, та тридцять тисяч і шість сотень керівників, що спонукували той народ до праці.
2CHR|3|1|І зачав Соломон будувати Господній дім в Єрусалимі на горі Морійя, що вказана була батькові його Давидові, на місці, яке приготовив Давид на тоці євусеянина Орнана.
2CHR|3|2|І зачав він будувати другого місяця, другого дня, четвертого року свого царювання.
2CHR|3|3|А це основа будови Божого дому: довжина шістдесят ліктів старою мірою, а ширина двадцять ліктів.
2CHR|3|4|А притвор, щодо довжини, був за шириною храму, двадцять ліктів, а вишина сто й двадцять. І покрив він його зсередини чистим золотом.
2CHR|3|5|А великий храм він покрив кипарисовим деревом, і покрив його добрим золотом, і наробив на ньому пальм та ланцюгів.
2CHR|3|6|І покрив він той храм дорогим каменем на оздобу, а золото золото було з Парваїму.
2CHR|3|7|І покрив він золотом храм, балки, пороги, і стіни його та його двері, а на стінах повирізував херувимів.
2CHR|3|8|І зробив дім Святого Святих: довжина його за шириною храму двадцять ліктів, і ширина його двадцять ліктів. І покрив він його добрим золотом, на таланти шість сотень.
2CHR|3|9|А вага цвяхів на шеклі золота п'ятдесят; і горниці покрив золотом.
2CHR|3|10|І зробив він у домі Святого Святих двох херувимів різьб'яною роботою, і покрив їх золотом.
2CHR|3|11|А крила херувимів: довжина їх двадцять ліктів, крило одного на п'ять ліктів, дотикалося стіни храму, а крило інше п'ять ліктів, дотикалося крила другого херувима.
2CHR|3|12|А крило другого херувима п'ять ліктів, дотикалося стіни храму, а крило інше п'ять ліктів, прилягало до крила іншого херувима.
2CHR|3|13|Розтягнені крила цих херувимів двадцять ліктів; і вони стояли на ногах своїх, а їхні обличчя до храму.
2CHR|3|14|І зробив він завісу, блакить, і пурпур, і червень, і віссон, і наробив на ній херувимів.
2CHR|3|15|І зробив він перед храмом два стовпи, тридцять і п'ять ліктів завдовжки, а маковиці, що на верху його, п'ять ліктів.
2CHR|3|16|І поробив ланцюги, як у девірі, і дав їх на верхи тих стовпів. І зробив сотню гранатових яблук, і дав на ланцюги.
2CHR|3|17|І поставив стовпи перед храмом, один з правиці, а один з лівиці. І назвав ім'я правому: Яхін, а ім'я лівому Боаз.
2CHR|4|1|І зробив мідяного жертівника, двадцять ліктів довжина йому і двадцять ліктів ширина йому, і десять ліктів височина йому.
2CHR|4|2|І зробив він лите море, десять на міру ліктем від краю його до краю його, навколо круглясте, і п'ять на міру ліктем височина йому. А шнур тридцять на міру ліктем оточував його навколо.
2CHR|4|3|А під ним постать волів, що зо всіх сторін оточують його, на десять ліктів на міру ліктем оточують море навколо; два ряди волів відлиті при відливанні його.
2CHR|4|4|Воно стояло на дванадцятьох волах, три обернені на північ, і три обернені на захід, і три обернені на південь, і три обернені на схід. А море на них зверху, а всі зади їх до нутра.
2CHR|4|5|А грубина його долоня, а край його як робота краю келіха, квітки лілеї. Містило воно три тисячі батів.
2CHR|4|6|І зробив десять умивальниць, і поставив п'ять з правиці, а п'ять з лівиці, щоб мити в них, приготовлене на цілопалення полощуть у них, а море для священиків, щоб митися в ньому.
2CHR|4|7|І зробив десять золотих свічників, як належалося, і поставив їх у храмі п'ять з правиці, а п'ять з лівиці.
2CHR|4|8|І зробив десять столів, і поставив у храмі, п'ять з правиці, а п'ять з лівиці. І зробив сто золотих кропильниць.
2CHR|4|9|І зробив священиче подвір'я та подвір'я велике, і двері до подвір'я, і їхні двері покрив міддю.
2CHR|4|10|А море поставив з правого боку на південний схід.
2CHR|4|11|І поробив Хурам горнята, і лопатки, і кропильниці. І покінчив Хурам робити працю, яку зробив для царя Соломона в Божому домі:
2CHR|4|12|два стовпи, і кулі, і дві маковиці на верху тих стовпів, і дві мережки на покриття обидвох куль маковиць, що на верхах стовпів,
2CHR|4|13|і чотири сотні гранатових яблук для обох мережок, два ряди гранатових яблук для однієї мережки, щоб покрити обидві кулі маковиць, що на переді тих стовпів.
2CHR|4|14|І поробив підстави, і поробив умивальниці на тих підставах,
2CHR|4|15|одне море, і дванадцять волів під ним,
2CHR|4|16|і горнята, і лопатки, і видельця, і всі їхні речі поробив Хурам-Авів цареві Соломонові для Господнього дому з виполіруваної міді.
2CHR|4|17|На Йорданській рівнині повідливав їх цар у глинистій землі між Суккотом та між Цередою.
2CHR|4|18|І наробив Соломон усіх цих речей дуже багато, бо не досліджена була вага міді.
2CHR|4|19|І поробив Соломон усі речі, що в Божому домі, та золотого жертівника й столи, а на них хліб показний,
2CHR|4|20|і свічники, і їхні лямпадки, щоб запалювати їх за постановою перед девіром, зо щирого золота.
2CHR|4|21|А квітки, і лямпадки, і щипчики із золота, з досконалого золота.
2CHR|4|22|А ножиці, і кропильниці, і ложки, і кадильниці зо щирого золота; а вхід до дому, його внутрішні двері до Святого Святих та двері дому до храму із золота.
2CHR|5|1|І була закінчена вся праця, яку зробив Соломон для Господнього дому. І Соломон повносив освячені речі свого батька Давида, і срібло, і золото, і всі ці речі дав до скарбниці Божого дому.
2CHR|5|2|Тоді Соломон зібрав до Єрусалиму Ізраїлевих старших, і всіх голів племен, начальників батьківських родів Ізраїлевих синів, щоб перенести ковчега Господнього заповіту з Давидового Міста, воно Сіон.
2CHR|5|3|І були зібрані до царя всі ізраїльтяни в свято, воно сьомого місяця.
2CHR|5|4|І поприходили всі Ізраїлеві старші, і Левити понесли ковчега.
2CHR|5|5|І понесли ковчега та скинію заповіту, і всі святі речі, що в скинії, несли їх священики та Левити.
2CHR|5|6|А цар Соломон та вся Ізраїлева громада, що зібралася при ньому перед ковчегом, приносили в жертву худобу дрібну та худобу велику, що через многоту не була ані записувана, ані лічена!
2CHR|5|7|І священики внесли ковчега Господнього заповіту до його місця, до девіру дому, до Святого Святих, під крила херувимів.
2CHR|5|8|А херувими простягали крила над місцем ковчега, і затінювали херувими над ковчегом та над його держаками зверху.
2CHR|5|9|А ті держаки були довгі, і головки тих держаків були видні з ковчегу, що перед девіром, а назовні не були видні. І були вони там аж до цього дня.
2CHR|5|10|У ковчезі не було нічого, тільки дві таблиці, що поклав Мойсей на Хориві, коли Господь склав був заповіта з Ізраїлевими синами при виході їх із Єгипту.
2CHR|5|11|І сталося, як священики виходили із святині, а всі священики, що були там, освятилися, без додержання черг,
2CHR|5|12|а Левити співаки, усі вони, аж до Асафа, Гемана, Єдутуна, і синів їхніх та братів їхніх, убрані в віссон, з цимбалами, із арфами та з цитрами, стояли на схід від жертівника, а з ними сто й двадцять священиків, що сурмили на сурмах,
2CHR|5|13|і було воно для сурмачів та співаків як одне, щоб подати один голос на хвалу та дяку Господеві, і як загримів голос на сурмах, і на цимбалах, і на музичних знаряддях, і як хвалили Господа: Добрий бо Він, бо навіки Його милосердя! то дім, дім Господній наповнився хмарою!...
2CHR|5|14|І не могли священики стояти й служити через ту хмару, бо слава Господня наповнила дім Божий!...
2CHR|6|1|Тоді Соломон проказав: Промовив Господь, що Він пробуватиме в мряці.
2CHR|6|2|А я збудував храм оселі Твоєї, і місце Твого пробування навіки!
2CHR|6|3|І повернув цар обличчя своє, та й поблагословив увесь Ізраїлів збір, увесь же Ізраїлів збір стояв.
2CHR|6|4|А він сказав: Благословенний Господь, Бог Ізраїлів, що Своїми устами говорив був із моїм батьком Давидом, і руками Своїми виконав, кажучи:
2CHR|6|5|Від того дня, коли Я вивів Свій народ з єгипетського краю, Я не вибрав Собі міста зо всіх Ізраїлевих племен, щоб збудувати храм на пробування Мого Імени там. І не вибрав Я нікого, щоб був володарем над народом Моїм, Ізраїлем.
2CHR|6|6|Та вибрав Я Єрусалим на пробування Мого Імени там, і вибрав Я Давида, щоб був над народом Моїм, Ізраїлем.
2CHR|6|7|І було на серці мого батька Давида збудувати храм для Ймення Господа, Бога Ізраїлевого.
2CHR|6|8|Та сказав Господь до мого батька Давида: За те, що на твоєму серці було збудувати храм для Ймення Мого, ти зробив добре, що було тобі на серці.
2CHR|6|9|Тільки ти не збудуєш цього храму, але син твій, що вийде із стегон твоїх, він збудує цей храм для Ймення Мого!
2CHR|6|10|І сповнив Господь Своє слово, що Він говорив. І став я замість батька свого Давида та й сів на Ізраїлевому троні, як говорив був Господь, і я збудував оцей храм для Ймення Господа, Бога Ізраїлевого.
2CHR|6|11|І поставив я там ковчега, що в ньому Господній заповіт, якого Він склав з Ізраїлевими синами.
2CHR|6|12|І став він перед Господнім жертівником навпроти всього Ізраїлевого збору, і простяг свої руки.
2CHR|6|13|А Соломон зробив був мідяне стояло, і поставив його на середину подвір'я, п'ять ліктів довжина йому, і п'ять ліктів ширина йому, а три лікті вишина йому. І став він на ньому, і став на коліна свої навпроти всього Ізраїлевого збору, і простяг свої руки до неба,
2CHR|6|14|та й сказав: Господи, Боже Ізраїлів! Нема подібного Тобі Бога на небі та на землі! Ти стережеш заповіта та милість для Своїх рабів, що ходять перед Твоїм лицем усім своїм серцем.
2CHR|6|15|Ти сповнив Своєму рабові Давидові, батькові моєму, те, що говорив йому. І говорив Ти йому Своїми устами, а рукою Своєю виповнив, як цього дня.
2CHR|6|16|А тепер, Господи, Боже Ізраїлів, сповни для Свого раба Давида, мого батька, те, що говорив Ти йому, кажучи: Не переведеться з-перед лиця Мого ніхто з тих, що мають сидіти на Ізраїлевому троні, якщо тільки сини твої будуть додержувати своїх доріг, щоб ходити в Законі Моїм, як ти ходив перед лицем Моїм.
2CHR|6|17|А тепер, Господи, Боже Ізраїлів, нехай буде запевнене слово Твоє, яке Ти говорив рабові Своєму Давидові.
2CHR|6|18|Бо чи ж справді Бог сидить з людиною на землі? Ось небо та небо небес не обіймають Тебе, що ж тоді храм цей, що я збудував?
2CHR|6|19|І Ти звернешся до молитви Свого раба та до його благання, Господи, Боже мій, щоб почути поклик та молитву, якою раб Твій молиться перед лицем Твоїм,
2CHR|6|20|щоб очі Твої були відкриті на цей храм удень та вночі, на те місце, про яке Ти сказав, що покладеш Ім'я Своє там, щоб почути молитву, якою буде молитися Твій раб на цьому місці.
2CHR|6|21|І Ти будеш прислухатися до благань Свого раба та Свого народу, Ізраїля, що будуть молитися на цьому місці. І Ти почуєш із місця Свого пробування, із небес і почуєш, і пробачиш.
2CHR|6|22|Якщо згрішить людина про ти свого ближнього, і буде примушена принести клятву, щоб присягнути, і клятва прийде перед Твоїм жертівником у цьому храмі,
2CHR|6|23|то Ти почуєш із небес, і зробиш, і розсудиш Своїх рабів, обвинуватиш несправедливого, щоб дати його дорогу на його голову, й усправедливиш справедливого, щоб дати йому за його справедливістю.
2CHR|6|24|А якщо Твій народ, Ізраїль, буде вдарений ворогом, бо прогрішив Тобі, і коли вони звернуться, і будуть хвалити Ім'я Твоє, і будуть молитися, і будуть благати Тебе в цьому храмі,
2CHR|6|25|то Ти почуєш із небес, і простиш гріх народу Свого, Ізраїля, і вернеш їх до землі, яку дав Ти їм та їхнім батькам!
2CHR|6|26|Коли затримається небо, і не буде дощу, бо прогрішаться Тобі, то вони помоляться на цьому місці, і будуть славити Ім'я Твоє, і з гріха свого навернуться, бо Ти будеш їх впокоряти,
2CHR|6|27|то Ти почуєш на небесах, і пробачиш гріх Своїх рабів та народу Свого, Ізраїля, бо покажеш їм ту добру дорогу, якою вони підуть, і Ти даси дощ на Край Свій, якого Ти дав Своєму народові на спадщину!
2CHR|6|28|Голод коли буде в Краю, моровиця коли буде, посуха, жовтачка, сарана, черва коли буде, коли його вороги гнобитимуть його в Краї міст його, коли буде яка пораза, яка хвороба,
2CHR|6|29|усяка молитва, усяке благання, що буде від якої людини чи від усього народу Твого, Ізраїля, коли кожен буде знати поразу свою та горе своє, і простягне руки свої до цього храму,
2CHR|6|30|то Ти почуєш із небес, із місця постійного пробування Свого, і пробачиш, і даси тому чоловікові за всіма його дорогами, бо Ти знаєш серце його, бо Ти один знаєш серце людських синів,
2CHR|6|31|щоб вони боялися Тебе, і ходили Твоїми дорогами по всі дні, які вони житимуть на поверхні землі, яку Ти дав батькам нашим!
2CHR|6|32|Також і чужинця, який не з народу Твого, Ізраїля, і він прийде з далекого краю ради Ймення Твого великого, і руки Твоєї Сильної та рамена Твого витягненого, і прийде, і помолиться в цьому храмі,
2CHR|6|33|то Ти почуєш це з небес, місця постійного пробування Свого, і зробиш усе, про що буде кликати до Тебе той чужинець, щоб усі народи землі пізнали Ім'я Твоє, та щоб боялися Тебе, як народ Твій, Ізраїль, і щоб пізнали вони, що Ім'я Твоє покликане над оцім храмом, що я збудував!
2CHR|6|34|Коли народ Твій вийде на війну на своїх ворогів, дорогою, якою Ти пошлеш їх, і помоляться вони до Тебе в напрямі до цього міста, що Ти вибрав його, та храму, що я збудував для Ймення Твого,
2CHR|6|35|то почуєш Ти з небес їхню молитву та їхнє благання, і вчиниш їм суд!
2CHR|6|36|Коли вони згрішать Тобі, бо немає людини, щоб вона не згрішила, і Ти розгніваєшся на них, і даси їх ворогові, а їхні поневільники візьмуть їх до неволі до краю далекого чи близького,
2CHR|6|37|і коли вони прийдуть до розуму в краю, куди взяті до неволі, і навернуться, і будуть благати Тебе в краю своєї неволі, говорячи: Ми згрішили, скривили дорогу свою, і були ми несправедливі,
2CHR|6|38|і коли вони навернуться до Тебе всім своїм серцем і всією душею своєю в краю своєї неволі, куди їх поневолили, і помоляться в напрямі до свого Краю, що Ти дав їхнім батькам, і в напрямі міста, яке Ти вибрав, та храму, що я збудував для Ймення Твого,
2CHR|6|39|то Ти почуєш із небес, із постійного місця пробування Свого, їхню молитву та їхні благання, і вчиниш їм суд, і простиш Своєму народові, що вони згрішили Тобі!
2CHR|6|40|Тепер, Боже мій, благаю, нехай будуть очі Твої відкриті, а уші Твої наставлені на слухання молитви цього місця!
2CHR|6|41|А тепер, Устань же, о Господи, Боже, на Свій відпочинок, Ти й ковчег сили Твоєї! Священики Твої, о Господи Боже, нехай у спасіння зодягнуться, а побожні Твої хай добром веселяться!
2CHR|6|42|Господи Боже, не відвертай лиця від Свого помазанця, згадай же про милість Своєму рабові Давиду!
2CHR|7|1|А коли Соломон закінчив молитися, то зійшов огонь із небес, поїв цілопалення та жертви, а слава Господня наповнила храм той!
2CHR|7|2|І священики не могли ввійти до Господнього дому, бо слава Господня наповнила дім Господній!
2CHR|7|3|А всі Ізраїлеві сини бачили, як сходив огонь та Господня слава на храм той, і вони попадали обличчям до землі на підлогу з камінних плит, і вклонилися до землі, і дякували Господеві: Добрий бо Він, бо навіки Його милосердя!
2CHR|7|4|А цар та ввесь народ приносили жертву перед Господнім лицем.
2CHR|7|5|І приніс цар Соломон на жертву худоби великої двадцять і дві тисячі, а худоби дрібної сто й двадцять тисяч. І виконали обряд освячення Божого дому цар та ввесь народ.
2CHR|7|6|А священики стояли на вартах своїх, а Левити зо знаряддями Господньої пісні, що поробив цар Давид на подяку Господеві, Бо навіки Його милосердя, коли Давид хвалив ними; і священики сурмили навпроти них, а ввесь Ізраїль стояв...
2CHR|7|7|І посвятив Соломон середину подвір'я, що перед Господнім домом, бо приніс там цілопалення та лій мирних жертв, бо мідяний жертівник, якого зробив Соломон, не міг умістити цілопалення й хлібної жертви та лою.
2CHR|7|8|І справив Соломон того часу те свято на сім день, а ввесь Ізраїль був з ним, дуже великий збір, що зійшовся звідти, де йдеться до Хамату, аж до єгипетського потоку.
2CHR|7|9|А восьмого дня справили віддання свята, бо обряд освячення жертівника справляли сім день, і свято сім день.
2CHR|7|10|А дня двадцятого й третього сьомого місяця відпустив він народ до їхніх наметів, радісних та веселосердих через усе те добро, що Господь учинив Давидові й Соломонові, та народові Своєму Ізраїлеві.
2CHR|7|11|І закінчив Соломон дім Господній та дім царський, та все, що приходило Соломонові на серце, щоб зробити в Господньому домі та в домі своєму, пощастило йому.
2CHR|7|12|І явився Господь Соломонові вночі та й сказав йому: Вислухав Я молитви твої, та вибрав оце місце для Себе на храм жертви.
2CHR|7|13|Якщо Я замкну небеса, і не буде дощу, і якщо накажу сарані поїсти землю, і якщо нашлю моровицю на народ Мій,
2CHR|7|14|і впокоряться люди Мої, що над ними кличеться Ім'я Моє, і помоляться, і будуть шукати Ім'я Мого, і повернуть зо злих своїх доріг, то Я вислухаю з небес, і прощу їхній гріх, та й вилікую їхній Край!
2CHR|7|15|Тепер очі Мої будуть відкриті, а уші Мої наставлені на слухання молитви цього місця.
2CHR|7|16|І тепер Я вибрав, і освятив цей храм, щоб Ім'я Моє було там аж навіки, Мої ж очі та серце Моє будуть там по всі дні.
2CHR|7|17|А тепер, якщо будеш ходити перед лицем Моїм, як ходив був батько твій Давид, щоб зробити все, що наказав Я тобі, і якщо будеш дотримуватися уставів Моїх та прав Моїх,
2CHR|7|18|то поставлю певно трона царства твого, як склав Я заповіта з батьком твоїм Давидом, говорячи: Не буде в тебе переводу нікому з пануючих в Ізраїлі!
2CHR|7|19|А якщо ви відвернетеся та покинете устави Мої й заповіді Мої, що Я дав вам, і підете, і будете служити іншим богам, і будете вклонятися їм,
2CHR|7|20|то Я повириваю їх з Моєї землі, яку дав їм, а цей храм, що Я освятив для Ймення Свого, відкину від лиця Свого, і дам його за приповістку та за посміховище серед усіх народів!
2CHR|7|21|А храм цей, що був найвищий, кожен, хто проходитиме біля нього, скам'яніє та й скаже: За що Господь зробив так цьому Краєві та храмові цьому?...
2CHR|7|22|І відкажуть: За те, що вони покинули Господа, Бога батьків своїх, Який вивів їх з єгипетського краю, і держалися міцно інших богів, і вклонялися їм, і служили їм, тому Він навів на них усе оце лихо!...
2CHR|8|1|І сталося по двадцятьох роках, коли Соломон будував дім Господній та свій дім,
2CHR|8|2|то міста, які дав Хурам Соломонові, Соломон розбудував їх, і осадив там Ізраїлевих синів.
2CHR|8|3|І пішов Соломон до Хават-Цови, і переміг її.
2CHR|8|4|І збудував він Тадмора в пустині, та всі міста для запасів, що побудував у Хаматі.
2CHR|8|5|І побудував він Бет-Хорон горішній та Бет-Хорон долішній, твердинні міста, мури, двері та засуви,
2CHR|8|6|і Баалат, і всі міста для запасів, що були в Соломона, і всі міста для колесниць, і міста для верхівців, і всяке пожадання Соломона, що жадав він збудувати в Єрусалимі й на Ливані, та в усьому Краї його панування.
2CHR|8|7|Увесь народ, позосталий з хіттеян, і з амореян, і з періззеян, і з хіввеян, і з євусеян, що вони не з Ізраїля,
2CHR|8|8|з їхніх синів, що зосталися по них у Краї, що їх не повигублювали Ізраїлеві сини, то їх Соломон узяв на данину, і це позосталося аж до цього дня.
2CHR|8|9|А Ізраїлевих синів Соломон не робив рабами для своєї праці, але вони були військові, і зверхники сторожі його, і зверхники колесниць його та його верхівців.
2CHR|8|10|І оце вони були зверхники-намісники царя Соломона, двісті і п'ятдесят, що панували над народом.
2CHR|8|11|А фараонову дочку перевів Соломон із Давидового Міста до дому, що збудував для неї, як сказав: Не буде сидіти мені жінка в домі Давида, Ізраїлевого царя, бо святий він, бо Господній ковчег увійшов у нього.
2CHR|8|12|Тоді Соломон приніс цілопалення для Господа на Господньому жертівнику, якого він збудував перед притвором,
2CHR|8|13|щоб за потребою кожного дня приносити жертву за Мойсеєвим наказом, на суботи, і на молодики, і на свята три рази в році: в свято Опрісноків, і в свято Тижнів, і в свято Кучок.
2CHR|8|14|І поставив він, за розпорядком Давида, батька свого, черги священиків на їхню службу, і Левитів на їхніх вартах на хвалу та на службу відповідно до священиків за потребою кожного дня, і придверних в їхніх чергах для кожної брами, бо такий був наказ Давида, Божого чоловіка.
2CHR|8|15|І не відступали вони від наказів царя про священиків та Левитів, щодо всякої речі й щодо скарбів.
2CHR|8|16|І була зроблена вся Соломонова праця аж до цього дня, від заложення Господнього дому й аж до закінчення його, коли був закінчений дім Господній.
2CHR|8|17|Тоді пішов Соломон до Ецйон-Ґеверу та до Елоту над морським берегом в едомському краї.
2CHR|8|18|І прислав йому Хурам через своїх рабів кораблі та рабів, що знали море. І прийшли вони з Соломоновими рабами до Офіру, і взяли звідти чотири сотні й п'ятдесят талантів золота, і привезли до царя Соломона.
2CHR|9|1|А цариця Шеви почула була про славу Соломонову, і прийшла випробувати Соломона загадками в Єрусалимі. Прийшла вона з дуже великим багатством, із верблюдами, що несли пахощі та безліч золота й дорогого каміння. І прийшла вона до Соломона, і говорила з ним про все, що було на серці її.
2CHR|9|2|І Соломон вияснив їй усі її запити, і не було запиту, незнаного Соломонові, якого не порішив би він їй.
2CHR|9|3|І побачила цариця Шеви всю Соломонову мудрість та дім, що він збудував,
2CHR|9|4|і їжу столу його, і мешкання рабів його, і поставу слуг його та їхні одежі, і чашників його, та їхні одежі, і вхід його, яким він уходить до Господнього дому, і не могла вона з дива вийти!
2CHR|9|5|І сказала вона до царя: Правдою було те, що я чула в своїм краї про твої діла та про твою мудрість.
2CHR|9|6|І не повірила я їхнім словам, аж поки сама не прийшла та не побачили мої очі, і ось не була представлена мені й половина великости твоєї мудрости: ти перевищив славу, про яку я чула!
2CHR|9|7|Щасливі люди твої, і щасливі оці твої слуги, що завжди стоять перед обличчям твоїм та слухають твою мудрість!
2CHR|9|8|Нехай буде благословенний Господь, Бог твій, що вподобав тебе, щоб посадити тебе на Свого трона за царя у Господа, Бога твого, через любов Бога твого до Ізраїля, щоб утвердити його навіки. І Він настановив тебе над ними царем, щоб чинити право та справедливість!
2CHR|9|9|І дала вона цареві сто й двадцять талантів золота, і дуже багато пахощів та дороге каміння. І більш уже не було таких пахощів, як ті, що цариця Шеви дала цареві Соломонові!
2CHR|9|10|І також Хурамові раби та раби Соломонові, що довозили золото з Офіру, спроваджували алмуґове дерево та дороге каміння.
2CHR|9|11|І поробив цар з алмуґового дерева сходи для Господнього дому та для дому царського, і гусла, і арфи для співаків. І такі речі, як вони, не бачені перед тим в юдейському Краї!
2CHR|9|12|А цар Соломон дав цариці Шеви все бажання її, чого вона бажала, окрім такого, що вона привезла до царя. І пішла вона назад до свого краю, вона та слуги її.
2CHR|9|13|І була вага того золота, що приходило для Соломона в одному році, шість сотень і шістдесят і шість талантів золота,
2CHR|9|14|окрім того, що приходило від купців та з торговлі ходячих. І всі царі арабські та намісники Краю довозили золото й срібло Соломонові.
2CHR|9|15|І зробив цар Соломон дві сотні великих щитів із кутого золота, шість сотень шеклів кутого золота йшло на одного щита,
2CHR|9|16|та три сотні щитів менших із кутого золота, три сотні шеклів золота йшло на одного щита. І цар віддав їх до дому Ливанського Лісу.
2CHR|9|17|І зробив цар великого трона зо слонової кости, і покрив його чистим золотом.
2CHR|9|18|У трона було шість східців та підніжжя з золота позад трону, та поруччя з цього й з того боку при місці сидіння, та два леви, що стояли при поруччях.
2CHR|9|19|І дванадцять левів стояли там на шости ступенях з того й з того боку. По всіх царствах не було так зробленого!
2CHR|9|20|І ввесь посуд на пиття царя Соломона золото, і всі речі дому Ливанського Лісу щире золото, нічого з срібла, воно за Соломонових днів не рахувалося за щось.
2CHR|9|21|Бо цареві кораблі ходили до Таршішу з Хурамовими рабами. Раз на три роки приходили таршіські кораблі, що довозили золото та срібло, слонову кість, і мавп та пав.
2CHR|9|22|І став цар Соломон найбільшим від усіх земних царів, щодо багатства та щодо мудрости.
2CHR|9|23|І всі земні царі хотіли бачити Соломона, щоб послухати його мудрости, що Бог дав у його серце.
2CHR|9|24|І вони приносили кожен свого дара, речі срібні та речі золоті, й одежу, зброю та пахощі, коні та мули, що на рік припадало.
2CHR|9|25|І було в Соломона чотири тисячі кінських жолобів та колесниць, і дванадцять тисяч верхівців, і він порозміщував їх по колесничних містах та при царі в Єрусалимі.
2CHR|9|26|І він панував над усіма царями від Річки й аж до краю филистимлян, і аж до єгипетської границі.
2CHR|9|27|І Соломон наскладав в Єрусалимі срібла, мов того каміння, а кедрів наскладав, щодо численности, як сикомори, що в Шефелі!
2CHR|9|28|А коней приводили Соломонові з Єгипту та з усіх країв.
2CHR|9|29|А решта Соломонових діл, перших та останніх, ото вони описані в історії пророка Натана, і в пророцтві шілонянина Ахійї, і в видіннях прозорливця Єді на Єровоама, Неватового сина.
2CHR|9|30|І царював Соломон в Єрусалимі над усім Ізраїлем сорок літ.
2CHR|9|31|І спочив Соломон за своїми батьками, і поховали його в Місті Давида, батька його, а замість нього зацарював син його Рехав'ам.
2CHR|10|1|І пішов Рехав'ам до Сихему, бо до Сихему зійшовся ввесь Ізраїль, щоб настановити його царем.
2CHR|10|2|І сталося, як почув це Єровоам, Неватів син, він був в Єгипті, куди втік від царя Соломона, то вернувся Єровоам з Єгипту.
2CHR|10|3|І послали й покликали його. І прийшов Єровоам та ввесь Ізраїль, і вони говорили до Рехав'ама, кажучи:
2CHR|10|4|Твій батько вчинив був тяжким наше ярмо, а ти полегши жорстоку роботу батька свого та тяжке його ярмо, що наклав він був на нас, і ми будемо служити тобі.
2CHR|10|5|А він відказав їм: Ідіть ще на три дні, і верніться до мене. І пішов той народ.
2CHR|10|6|І радився цар Рехав'ам зо старшими, що стояли перед обличчям його батька Соломона, коли він був живий, говорячи: Як ви радите відповісти цьому народові?
2CHR|10|7|І вони говорили йому, кажучи: Якщо ти будеш добрим для цього народу, і зробиш за волею їх, і говоритимеш їм добрі слова, то вони будуть тобі рабами по всі дні.
2CHR|10|8|Та він відкинув пораду старших, що радили йому, і радився з молодиками, що виросли разом із ним, що стояли перед ним.
2CHR|10|9|І сказав він до них: Що ви радите, і що відповімо цьому народові, який говорив мені, кажучи: Полегши ярмо, яке твій батько наклав був на нас.
2CHR|10|10|І говорили з ним ті молодики, що виросли з ним, кажучи: Так скажеш тому народові, що промовляв до тебе, говорячи: Твій батько вчинив був тяжким наше ярмо, а ти дай полегшу нам. Отак скажеш до них: Мій мізинець грубший за стегна мого батька!
2CHR|10|11|А тепер: мій батько наклав був на вас тяжке ярмо, а я добавлю до вашого ярма! Батько мій карав вас бичами, а я битиму скорпіонами...
2CHR|10|12|І прийшов Єровоам та ввесь народ до Рехав'ама третього дня, як цар говорив, кажучи: Верніться до мене третього дня.
2CHR|10|13|І цар жорстоко відповів їм. І відкинув цар Рехав'ам пораду старших,
2CHR|10|14|і говорив до них за порадою тих молодиків, кажучи: Мій батько вчинив був тяжким ваше ярмо, а я добавлю до нього! Батько мій карав вас бичами, а я скорпіонами!...
2CHR|10|15|І не послухався цар народу, бо це спричинене було від Бога, щоб справдити Господеві слово Своє, яке Він говорив був через шілонянина Ахійю, Неватового сина.
2CHR|10|16|І побачив увесь Ізраїль, що цар не послухався їх, і народ відповів цареві, кажучи: Яка нам частина в Давиді? І спадщини нема нам у сині Єссея! Усі до наметів своїх, о Ізраїлю! Познай тепер дім свій, Давиде! І пішов увесь Ізраїль до наметів своїх...
2CHR|10|17|А Ізраїлеві сини, що сиділи в Юдиних містах, то над ними зацарював Рехав'ам.
2CHR|10|18|І послав цар Рехав'ам Гадорама, що був над даниною, та Ізраїлеві сини закидали його камінням, і він помер. А цар Рехав'ам поспішив сісти на колесницю та втекти до Єрусалиму...
2CHR|10|19|І відпав Ізраїль від Давидового дому, і так є аж до цього дня.
2CHR|11|1|І прийшов Рехав'ам до Єрусалиму, і зібрав дім Юдин та Веніяминів, сто й вісімдесят тисяч вибраних військових, щоб воювати з Ізраїлем, щоб вернути царство Рехав'амові.
2CHR|11|2|І було Господнє слово до Шемаї, чоловіка Божого, говорячи:
2CHR|11|3|Скажи Рехав'амові, Соломонову синові, цареві Юдиному, та всьому Ізраїлеві в Юді та в Веніямині, говорячи:
2CHR|11|4|Так сказав Господь: Не йдіть і не воюйте з своїми братами! Верніться кожен до дому свого, бо ця річ сталася від Мене! І вони послухалися Господніх слів, і вернулися з походу на Єровоама.
2CHR|11|5|І осівся Рехав'ам в Єрусалимі, і побудував твердинні міста в Юді.
2CHR|11|6|І збудував він Віфлеєма, і Етама, і Текою,
2CHR|11|7|і Бет-Цура, і Сохо, і Адуллама,
2CHR|11|8|і Ґата, і Марешу, і Зіфа,
2CHR|11|9|і Адораїма, і Лахіша, і Азеку,
2CHR|11|10|і Цор'у, і Айялона, і Хеврона, що в Юді та в Веніямині, міста твердинні.
2CHR|11|11|І зміцнив він ті твердині, і дав у них начальників, і запаси, і оливи, і вина,
2CHR|11|12|а до кожного окремого міста великі щити та ратища, і дуже сильно їх позміцнював. І був його Юда та Веніямин.
2CHR|11|13|А священики та Левити, що були в усьому Ізраїлі, зібралися до нього з усієї їхньої границі.
2CHR|11|14|Бо Левити кидали пасовиська свої та власність свою, і приходили до Юди та до Єрусалиму, бо Єровоам та сини його усунули їх від священичого служіння Господеві,
2CHR|11|15|і понаставляли собі священиків для пагірків та демонів, та для тельців, що він понароблював.
2CHR|11|16|А за ними, зо всіх Ізраїлевих племен ті, що віддавали своє серце шукати Господа, Бога Ізраїля, приходили до Єрусалиму приносити жертви Господеві, Богові батьків своїх.
2CHR|11|17|І зміцнили вони Юдине царство, і підсилили Рехав'ама, Соломонового сина, на три роки, бо вони ходили три роки дорогою Давида та Соломона.
2CHR|11|18|І взяв собі Рехав'ам жінку Махалат, дочку Єрімота, Давидового сина, та Авіхаїл, дочку Еліава, Ісаєвого сина.
2CHR|11|19|І вона породила йому синів: Єуша, і Шемарію, Загама.
2CHR|11|20|А по ній він узяв Мааху, дочку Авесаломову, і вона породила йому Авійю, і Аттая, і Зізу, і Шеломіта.
2CHR|11|21|І покохав Рехав'ам Мааху, Авесаломову дочку, над усіх жінок своїх та наложниць своїх, бо він узяв вісімнадцять жінок та шістдесят наложниць, і породив двадцять і вісім синів та шістдесят дочок.
2CHR|11|22|А за голову Рехав'ам поставив Авійю, Маахиного сина, за володаря серед братів його, бо він хотів настановити його царем.
2CHR|11|23|І мудро він чинив, і порозсилав усіх синів своїх до всіх країв Юди й Веніямина, до всіх твердинних міст, і дав їм багате утримання, і підшукав їм багато жінок.
2CHR|12|1|І сталося, як зміцніло Рехав'амове царство й став він сильний, то покинув він, і ввесь Ізраїль із ним, Господнього Закона.
2CHR|12|2|І сталося п'ятого року царя Рехав'ама, пішов Шішак, єгипетський цар, на Єрусалим, бо вони спроневірилися Господеві,
2CHR|12|3|з тисячею й двомастами колесниць та з шістдесятьма тисячами верхівців: і не було числа для народу, що прийшов із ним з Єгипту, ливіянам, суккійянам та кушанам.
2CHR|12|4|І здобув він твердинні міста, що в Юді, і прийшов аж до Єрусалиму.
2CHR|12|5|А пророк Шемая прийшов до Рехав'ама та Юдиних зверхників, що зібралися до Єрусалиму, утікаючи перед Шішаком, та й сказав до них: Так сказав Господь: Ви залишили Мене, а тому Я залишив вас і видав у Шішакову руку!
2CHR|12|6|І впокорилися Ізраїлеві зверхники та цар і сказали: Справедливий Господь!
2CHR|12|7|А коли Господь побачив, що вони впокорилися, то було Господнє слово до Шемаї, говорячи: Упокорилися вони, не нищитиму їх, але дам їм трохи людей на порятунок, і не виллється гнів Мій на Єрусалим через Шішака.
2CHR|12|8|Бо вони стануть йому за рабів, та й пізнають тоді службу Мені та службу царствам земним.
2CHR|12|9|І вийшов Шішак, єгипетський цар, на Єрусалим, і забрав скарби Господнього дому та скарби дому царевого, і все позабирав. І забрав він золоті щити, що Соломон поробив був.
2CHR|12|10|А цар Рехав'ам поробив замість них мідяні щити, і склав їх на руки зверхника сторожів, що стерегли вхід до царського дому.
2CHR|12|11|І бувало, як тільки цар ішов до Господнього дому, приходили бігуни, та й носили їх, а потім вертали їх до комори бігунів.
2CHR|12|12|А коли він впокорився, то відвернувся від нього Господній гнів, і не знищив його аж до вигублення. Та й у Юдеї були ще справи добрі.
2CHR|12|13|І зміцнився цар Рехав'ам в Єрусалимі й царював. А Рехав'ам був віку сорока й одного року, коли зацарював, і царював він сімнадцять літ в Єрусалимі, у тому місті, яке вибрав Господь зо всіх Ізраїлевих племен, щоб покласти там Своє Ймення. А ім'я його матері аммонітка Наама.
2CHR|12|14|І робив він лихе, бо не схиляв свого серця, щоб звертатися до Господа.
2CHR|12|15|А Рехав'амові діла, перші й останні, ото вони описані в історії пророка Шемаї та прозорливця Іддо: Родословні книги. І точилися війни поміж Рехав'амом та Єровоамом по всі дні.
2CHR|12|16|І спочив Рехав'ам зо своїми батьками, і був він похований у Давидовому Місті, а замість нього зацарював його син Авійя.
2CHR|13|1|Вісімнадцятого року царя Єровоама та зацарював Авійя над Юдою.
2CHR|13|2|Три роки царював він в Єрусалимі. А ім'я його матері Міхая, дочка Уріїла з Ґів'ї. І війна точилася між Авійєю та між Єровоамом.
2CHR|13|3|І зачав Авійя війну з військом хоробрих вояків, чотири сотні тисяч вибраних мужів, а Єровоам приготовився до війни з ним з вісьмома сотнями тисяч вибраних мужів, хоробрих вояків.
2CHR|13|4|І встав Авійя з-над гори Цемараїм, що в Єфремових горах, та й сказав: Послухайте мене, Єровоаме, та ввесь Ізраїлю!
2CHR|13|5|Чи ж не вам знати, що Господь, Бог Ізраїлів, дав Давидові царство над Ізраїлем навіки, йому та синам його, соляною умовою?
2CHR|13|6|Та встав Єровоам, Неватів син, раб Соломона, Давидового сина, і збунтувався на пана свого.
2CHR|13|7|І зібралися до нього люди пусті, нікчемні, і стали міцніші від Рехав'ама, Соломонового сина. А Рехав'ам був юнак та м'якосердий, і не був сильним проти них.
2CHR|13|8|А тепер ви говорите, щоб бути сильними проти Господнього царства в руці Давидових синів, а вас велика кількість, і з вами золоті тельці, яких Єровоам понароблював вам за богів.
2CHR|13|9|Чи ж ви не повиганяли Господніх священиків, Ааронових синів, та Левитів? І понаставляли ви собі священиків, як ставлять народи цих країв, кожен, хто прийде, щоб посвятитися молодим бичком та сімома баранами, то стає священиком для того, що не є Богом.
2CHR|13|10|А ми, Бог наш Господь, і ми не полишили Його, а наші священики, що служать Господеві, це Ааронові сини, а Левити при службі.
2CHR|13|11|І ми приносимо Господеві цілопалення кожного ранку та кожного вечора, і запашне кадило, і укладання хліба на чистому столі, і золотий свічник та лямпади його, щоб запалювати кожного вечора, бо ми стережемо службу Господа, нашого Бога, а ви полишили Його!
2CHR|13|12|І ось з нами на чолі Бог, і священики Його, і голосні сурми, щоб сурмити на вас. Ізраїлеві сини, не воюйте з Господом, Богом вашим, бо вам не поведеться!
2CHR|13|13|А Єровоам вирядив засідку, щоб пішла позад них, і були вони перед Юдою, а засідка позад них.
2CHR|13|14|І обернулися юдеї, аж ось у них бій спереду та ззаду! І кликали вони до Господа, а священики сурмили в сурми...
2CHR|13|15|І закричали юдеї. І сталося, як юдеї закричали, то Бог ударив Єровоама та всього Ізраїля перед Авійєю та перед Юдою.
2CHR|13|16|І повтікали ізраїльтяни перед Юдою, і Бог дав їх в їхню руку.
2CHR|13|17|І вдарили в них Авійя та народ його великою поразою, і попадали трупи з Ізраїля, п'ять сотень тисяч вибраних мужів!
2CHR|13|18|І впокорилися Ізраїлеві сини того часу, а Юдині сини зміцніли, бо опиралися на Господа, Бога їхніх батьків.
2CHR|13|19|І гнався Авійя за Єровоамом, і здобув від нього міста: Бет-Ел та залежні його міста, і Єшану та залежні її міста, і Ефрон та залежні його міста.
2CHR|13|20|І Єровоам не затримав сили вже за днів Авійї. І вдарив його Господь, і він помер.
2CHR|13|21|І зміцнився Авійя, і взяв собі чотирнадцять жінок, і породив двадцять і двоє синів та шістнадцятеро дочок.
2CHR|13|22|А решта Авійєвих діл, і дороги його та слова його описані в історії пророка Іддо.
2CHR|14|1|(13-23) І спочив Авійя зо своїми батьками, і поховали його в Давидовому Місті, а замість нього зацарював син його Аса. За його днів заспокоївся Край на десять літ.
2CHR|14|2|(14-1) І робив Аса добре та вгодне в очах Господа, Бога свого.
2CHR|14|3|(14-2) І повсував він жертівники чужих богів та пагірки, і порозбивав камінні стовпи для божків, і постинав святі дерева.
2CHR|14|4|(14-3) І наказав він Юді звертатися до Господа, Бога батьків своїх, і виконувати Його Закона та заповідь.
2CHR|14|5|(14-4) І повсував він зо всіх Юдиних міст пагірки та подоби сонця. І заспокоїлося царство при ньому.
2CHR|14|6|(14-5) І побудував він твердинні міста в Юді, бо заспокоївся Край, і не було на нього війни за тих років, бо Господь дав йому мир.
2CHR|14|7|(14-6) І сказав він до Юди: Побудуймо ці міста, й оточімо муром та баштами, ворітьми та засувами. Іще він, цей Край, наш, бо зверталися ми до Господа, нашого Бога. Зверталися ми, і Він дав нам мир навколо. І побудували, і їм щастило.
2CHR|14|8|(14-7) І було в Аси війська: носіїв великих щитів та ратищ з Юди три сотні тисяч, а з Веніямина таких, що носять малого щита, та лучників двісті й вісімдесят тисяч. Усі вони хоробрі вояки.
2CHR|14|9|(14-8) І вийшов на них кушеянин Зерах із військом у тисячу тисяч та з трьома сотнями колесниць, і прибув аж до Мареші.
2CHR|14|10|(14-9) І вийшов Аса проти нього, і вони вставилися до бою в долині Цефат при Мареші.
2CHR|14|11|(14-10) І кликнув Аса до Господа. Бога свого, та й сказав: Господи, нема кому, крім Тебе, допомогти численному або безсилому. Допоможи нам, Господи, Боже наш, бо ми на Тебе опираємося, і в Ім'я Твоє ми прийшли на цю безліч. Господи, Ти Бог наш, нехай людина не має сили проти Тебе!
2CHR|14|12|(14-11) І побив Господь кушеян перед Асою та перед Юдою, і кушеяни повтікали.
2CHR|14|13|(14-12) І гнав їх Аса та народ, що був з ним, аж до Ґерару. І попадало з кушеян багато, так що ніхто з них не залишився живий, бо вони були поторощені перед Господнім лицем та перед табором Його. І понесли вони дуже багато здобичі.
2CHR|14|14|(14-13) І побили вони всі міста навколо Ґерару, бо Господній страх був на них. І пограбували вони всі ті міста, бо в них було багато здобичі.
2CHR|14|15|(14-14) Порозбивали вони також намети чередників, і зайняли дуже багато дрібної худоби та верблюдів, та й вернулися до Єрусалиму.
2CHR|15|1|А Азарія, син Оведів, злинув на нього Дух Божий.
2CHR|15|2|І вийшов він перед Асу та й сказав йому: Послухайте мене, Асо та ввесь Юдо й Веніямине! Господь з вами, якщо будете з Ним, і якщо будете Його шукати, дасть вам знайти Себе. А якщо ви полишите Його, полишить Він вас!
2CHR|15|3|У Ізраїля було багато днів, коли був він без правдивого Бога, і без священика-вчителя та без Закону.
2CHR|15|4|І вернувся він в утиску своєму до Господа, Бога Ізраїлевого, і вони шукали Його, і Він дав їм знайти Себе.
2CHR|15|5|А тими часами не було спокою ані тому, хто виходить, ані тому, хто входить, бо були великі неспокої в усіх мешканців Краю.
2CHR|15|6|І воював народ проти народу та місто проти міста, бо Бог побентежив їх усяким лихом.
2CHR|15|7|А ви будьте міцні, і нехай не слабнуть ваші руки, бо є нагорода для вашої чинности!
2CHR|15|8|А коли Аса почув оці слова та пророцтво, яке говорив пророк Азарія, син Оведів, то зміцнився, і повикидав поганські гидоти зо всього краю Юдиного та Веніяминового, та з міст, які він здобув з Єфремових гір, і відновив Господнього жертівника, що перед Господнім притвором.
2CHR|15|9|І зібрав він усього Юду й Веніямина та тих, що мешкали часово з ними з Єфрему, і з Манасії, і з Симеона, бо дуже багато поперебігали до нього з Ізраїля, коли побачили, що з ним Господь, його Бог.
2CHR|15|10|І вони зібралися до Єрусалиму третього місяця, п'ятнадцятого року царювання Аси.
2CHR|15|11|І принесли вони того дня в жертву для Господа зо здобичі, яку поприводили: худоби великої сім сотень, а худоби дрібної сім тисяч.
2CHR|15|12|І ввійшли вони в умову, щоб звертатися до Господа, Бога їхніх батьків, усім своїм серцем та всією своєю душею.
2CHR|15|13|А кожен, хто не буде звертатися до Господа, Бога Ізраїля, буде забитий від малого й аж до великого, від чоловіка й аж до жінки.
2CHR|15|14|І заприсяглися вони Господеві голосом сильним, і окликом, і сурмами, і рогами.
2CHR|15|15|І тішився ввесь Юда тією присягою, бо вони заприсяглися всім серцем своїм, і всією своєю волею шукали Його, і Він дав їм знайти Себе. І Господь дав їм мир навколо.
2CHR|15|16|І навіть Мааху, матір царя Аси, й її він позбавив права бути царицею, бо вона зробила була ідола Астарти. І Аса порубав боввана її, і розтер, і спалив у долині Кедрон.
2CHR|15|17|Та пагірки не минулися в Ізраїля, але Асине серце було все з Господом по всі його дні.
2CHR|15|18|І вніс він до Божого дому святі речі свого батька та святі речі свої, срібло, і золото, і посуд.
2CHR|15|19|А війни не було аж до тридцять й п'ятого року царювання Аси.
2CHR|16|1|Тридцятого й шостого року царювання Аси пішов Баша, Ізраїлів цар, проти Юди, і будував Раму, щоб не дати нікому від Аси, царя Юдиного, виходити та входити.
2CHR|16|2|І виніс Аса срібло та золото із скарбниць Господнього дому та дому царевого, і послав до Бен-Гадада, царя сирійського, що сидів у Дамаску, говорячи:
2CHR|16|3|Є умова між мною та між тобою, і між батьком моїм та батьком твоїм. Ось послав я тобі срібла та золота, іди, зламай умову свою з Башею, царем Ізраїлевим, і нехай він відійде від мене.
2CHR|16|4|І послухався Бен-Гадад царя Аси, і послав зверхників свого війська на Ізраїлеві міста, і вони поруйнували Іййона, і Дана, і Авел-Маїма та всі запаси міст Нефталимових.
2CHR|16|5|І сталося, як Баша це почув, то перестав будувати Раму, і спинив свою працю.
2CHR|16|6|А цар Аса взяв усього Юду, і вони повиносили каміння Рами та її дерево, що з них будував був Баша, і побудував з того Ґеву та Міцпу.
2CHR|16|7|А того часу прийшов прозорливець Ханані до Аси, Юдиного царя, та й сказав до нього: Через те, що ти спирався на сирійського царя, а не сперся на Господа, Бога свого, тому втекло з твоєї руки військо сирійського царя.
2CHR|16|8|Чи ж не були кушеяни та ливіяни військом дуже великим, колесницями й верхівцями дуже численними? Та коли ти сперся на Господа, Він дав їх у твою руку.
2CHR|16|9|Бо очі Господні дивляться по всій землі, щоб зміцнити тих, у кого все їхнє серце до Нього. Тому зробив ти нерозумно, бо відтепер будуть у тебе війни!
2CHR|16|10|І розгнівався Аса на прозорливця, і дав його до в'язниці, бо був у гніві на нього за це. І Аса тиснув декого з народу того часу.
2CHR|16|11|І оце Асині діла, перші та останні, ось вони описані в книзі Юдиних та Ізраїлевих царів.
2CHR|16|12|І занедужав Аса тридцятого й дев'ятого року свого царювання на свої ноги, і хвороба його була тяжка. Та й у хворобі своїй не звертався він до Господа, але до лікарів.
2CHR|16|13|І спочив Аса з своїми батьками, і помер сорокового й першого року свого царювання.
2CHR|16|14|І поховали його в його гробницях, які він викопав собі в Давидовому Місті. І поклали його на ложі, що він наповнив пахощами та різними, по-містецькому зробленими, мастями. І спалили йому дуже велике паління.
2CHR|17|1|А замість нього зацарював син його Йосафат, та зміцнився над Ізраїлем.
2CHR|17|2|І поставив він військо по всіх укріплених Юдиних містах, і дав залоги в Юдиному краї та в Єфремових містах, які був здобув його батько Аса.
2CHR|17|3|І був Господь з Йосафатом, бо він ходив першими дорогами батька свого Давида, і не шукав Ваалів.
2CHR|17|4|Бо він звертався до Бога свого батька, і ходив за Його заповідями, а не за чином Ізраїля.
2CHR|17|5|І Господь зміцнив його царство в руці його, і вся Юдея давала дарунка Йосафатові, і було в нього багато багатства та слави.
2CHR|17|6|І повищилось серце його на Господніх дорогах, і він іще повсовував пагірки та Астарти з Юди.
2CHR|17|7|А третього року свого царювання послав він до своїх зверхників, до Бен-Хаїла, і до Овадії, і до Захарія, і до Натанаїла, і до Міхаї, щоб вони навчали в Юдиних містах.
2CHR|17|8|А з ними були Левити: Шемая, і Натанія, і Зевадія, і Асаїл, і Шемірамот, і Єгонатан, і Адонійя, і Товійя, і Тов-Адонійя, Левити, а з ними Елішама та Єгорам, священики.
2CHR|17|9|І навчали вони в Юдеї, а з ними була книга Закону Господнього. І ходили вони довкола по всіх Юдиних містах, і навчали серед народу.
2CHR|17|10|І був страх Господній на всіх царствах краю, що навколо Юди, і вони не воювали з Йосафатом.
2CHR|17|11|А від филистимлян приносили Йосафатові дари та срібло данини; також араби приводили йому дрібну худобу: сім тисяч і сім сотень баранів та сім тисяч і сім сотень козлів.
2CHR|17|12|І Йосафат усе зростав угору. І побудував він в Юді твердині та міста на запаси.
2CHR|17|13|І мав він багато добра по Юдиних містах, і мужів військових, хоробрих вояків в Єрусалимі.
2CHR|17|14|А оце їхній перегляд, за домами їхніх батьків. Від Юди тисячники: зверхник Адна, а з ним три сотні тисяч хоробрих вояків.
2CHR|17|15|А при ньому зверхник Єгоханан, а з ним двісті й вісімдесят тисяч.
2CHR|17|16|А при ньому Амасія, син Зіхрі, що присвятив себе Господеві, а з ним двісті тисяч хоробрих вояків.
2CHR|17|17|А від Веніямина: хоробрий вояк Ел'яда, а з ним двісті тисяч узброєних луком та щитом.
2CHR|17|18|А при ньому Єгозавад, а з ним сто й вісімдесят тисяч узброєного війська.
2CHR|17|19|Оці служили цареві, опріч тих, яких цар умістив по твердинних містах по всьому Юді.
2CHR|18|1|І було в Йосафата багато багатства та слави, і він посвоячився з Ахавом.
2CHR|18|2|А по кількох роках пішов він до Ахава до Самарії. І Ахав нарізав багато худоби дрібної та худоби великої йому та народові, що з ним, і намовив його піти на ґілеадський Рамот.
2CHR|18|3|І сказав Ахав, цар Ізраїлів, до Йосафата, царя Юдиного: Чи підеш зо мною до ґілеадського Рамоту? А той відказав йому: Я як ти, народ мій як твій народ, і буду з тобою на війні.
2CHR|18|4|І сказав Йосафат до Ізраїлевого царя: Вивідай зараз слово Господнє!
2CHR|18|5|І зібрав Ізраїлів цар пророків, чотири сотні чоловіка, та й сказав до них: Чи йти нам на війну на ґілеадський Рамот, чи занехати? А ті сказали: Іди, і Бог дасть його в цареву руку!
2CHR|18|6|І сказав Йосафат: Чи нема тут іще Господнього пророка, і звернімось до нього.
2CHR|18|7|І сказав Ізраїлів цар до Йосафата: Є ще один муж, щоб через нього звернутися до Господа. Та я ненавиджу його, бо він не пророкує на мене добре, а по всі дні свої тільки лихе. Це Міхей, син Їмлин. А Йосафат відказав: Нехай цар не говорить таке!
2CHR|18|8|І покликав Ізраїлів цар одного евнуха й сказав: Приведи скоріше Міхея, Їмлиного сина!
2CHR|18|9|А цар Ізраїлів та Йосафат, цар Юдин, сиділи кожен на троні своїм, повбирані в шати; а сиділи вони при вході брами Самарії, а всі пророки пророкували перед ними.
2CHR|18|10|А Цідкійя, Кенаанин син, зробив собі залізні роги й сказав: Так сказав Господь: Оцим будеш бодати сиріян аж до вигублення їх!
2CHR|18|11|І всі пророки пророкували так, говорячи: Виходь до ґілеадського Рамоту, і май успіх, і Господь дасть його в цареву руку!
2CHR|18|12|А той посланець, що пішов покликати Міхея, говорив до нього, кажучи: Ось слова тих пророків, одноусно звіщають цареві добро. Нехай же буде слово твоє таке, як кожного з них, і ти говоритимеш добре.
2CHR|18|13|І сказав Міхей: Як живий Господь, те, що скаже Господь, тільки те говоритиму!
2CHR|18|14|І прийшов він до царя, а цар сказав до нього: Міхею, чи йти на війну до ґілеадського Рамоту, чи занехати? А той відказав: Вийдіть, і будете мати успіх, і вони будуть дані в вашу руку.
2CHR|18|15|І сказав йому цар: Аж скільки разів я заприсягав тебе, що ти не говоритимеш мені нічого, тільки правду в Ім'я Господа?
2CHR|18|16|А той відказав: Я бачив усього Ізраїля, розпорошеного по горах, немов вівці, що не мають пастуха. І сказав Господь: Немає в них пана, нехай вернуться з миром кожен до дому свого!
2CHR|18|17|І сказав Ізраїлів цар до Йосафата: Чи ж не казав я тобі, він не буде пророкувати мені доброго, а тільки лихе?
2CHR|18|18|А Міхей відказав: Тому послухайте Господнього слова: Бачив я Господа, що сидів на престолі Своїм, а все небесне військо стояло по правиці Його та по лівиці Його.
2CHR|18|19|І сказав Господь: Хто намовить Ахава, Ізраїлевого царя, і він вийде й упаде в ґілеадському Рамоті? І говорили: той говорив так, а той говорив так.
2CHR|18|20|І вийшов дух, і став перед Господнім лицем та й сказав: Я намовлю його! І сказав йому Господь: Чим?
2CHR|18|21|А той відказав: Я вийду й стану духом неправди в устах усіх його пророків. А Господь сказав: Ти намовиш, а також переможеш; вийди та й зроби так!
2CHR|18|22|А тепер оце Господь дав духа неправди в уста оцих твоїх пророків, і Господь говорив на тебе недобре...
2CHR|18|23|І підійшов Цідкійя, Кенаанин син, і вдарив Міхея по щоці та й сказав: Кудою це перейшов Дух Господній від мене, щоб говорити з тобою?
2CHR|18|24|А Міхей відказав: Ось ти побачиш це того дня, коли ввійдеш до внутрішньої кімнати, щоб сховатися...
2CHR|18|25|І сказав Ізраїлів цар: Візьміть Міхея, і відведіть його до Амона, зверхника міста, та до Йоаша, царевого сина,
2CHR|18|26|та й скажете: Отак сказав цар: Посадіть оцього до в'язничного дому, і давайте йому їсти скупо хліба й скупо води, аж поки я не вернуся з миром.
2CHR|18|27|А Міхей відказав: Якщо справді вернешся ти з миром, то не говорив Господь через мене. І до того сказав: Слухайте це, усі люди!
2CHR|18|28|І вийшов Ізраїлів цар та Йосафат, цар Юдин, до ґілеадського Рамоту.
2CHR|18|29|І сказав Ізраїлів цар до Йосафата: Я переберуся й піду на бій, а ти вбери свої шати! І перебрався Ізраїлів цар, і пішли на бій.
2CHR|18|30|А сирійський цар наказав зверхникам своїх колесниць, говорячи: Не воюйте ні з малим, ні з великим, а тільки з самим Ізраїлевим царем!
2CHR|18|31|І сталося, як зверхники колесниць побачили Йонатана, то вони сказали: Це Ізраїлів цар! І вони оточили його, щоб воювати. І закричав Йосафат, і Господь допоміг йому, і Бог звабив їх від нього.
2CHR|18|32|І сталося, як зверхники колесниць побачили, що це не Ізраїлів цар, то повернули від нього.
2CHR|18|33|А один чоловік знехотя натягнув лука, та й ударив Ізраїлевого царя між підв'язанням пояса та між панцерем. А той сказав візникові: Заверни назад, і випровадь мене від війська, бо я ранений...
2CHR|18|34|І збільшився бій того дня, а Ізраїлів цар був поставлений на колесниці проти сиріян аж до вечора. І помер він під час заходу сонця...
2CHR|19|1|І вернувся Йосафат, цар Юдин, із миром до дому свого до Єрусалиму.
2CHR|19|2|І вийшов перед нього прозорливець Єгу, син Ханані, та й сказав до царя Йосафата: Чи будеш допомагати несправедливому, а тих, хто ненавидить Господа, будеш любити? І за це на тобі гнів від Господнього лиця.
2CHR|19|3|Але й добрі речі знайшлися при тобі, бо ти повигублював Астарти з Краю, і нахилив своє серце, щоб шукати Господа.
2CHR|19|4|І осівся Йосафат в Єрусалимі, і він знову виходив між народ від Беер-Шеви аж до Єфремових гір, і навертав їх до Господа, Бога їхніх батьків.
2CHR|19|5|І понаставляв він суддів у Краю, по всіх укріплених Юдиних містах, для кожного міста.
2CHR|19|6|І сказав він до суддів: Дивіться, що ви робите, бо не для людини ви судите, але для Господа, і Він з вами в справі суду.
2CHR|19|7|А тепер нехай буде Господній страх на вас. Стережіться й робіть, бо нема в Господа, Бога нашого, кривди, ані огляду на особу, ані брання дарунка.
2CHR|19|8|А також в Єрусалимі понаставляв Йосафат з Левитів і з священиків та з голів батьківських домів Ізраїля для Господнього суду та для суперечок. І вернулися вони до Єрусалиму.
2CHR|19|9|І він наказав їм, говорячи: Отак чиніть у страху Господньому, вірністю та цілим серцем.
2CHR|19|10|А щодо всякої суперечки, що прийде до вас від ваших братів, що сидять по містах своїх, де треба розсудити чи то за кров, чи то за Закон, чи то за заповідь, устави, чи за права, то остережете їх, і вони не згрішать Господеві, і не буде гніву на вас та на ваших братів. Так робіть, і не згрішите!
2CHR|19|11|А ось священик Амарія голова над вами до всяких Господніх речей, а Завадія, син Ізмаїлів, володар Юдиного дому, до всякої царевої речі, і писарі Левити перед вами. Будьте міцні й зробіть, і нехай буде Господь з добрим!
2CHR|20|1|І сталося по тому, пішли моавітяни та аммонітяни, а з ними деякі з меунян, проти Йосафата на війну.
2CHR|20|2|І прийшли, і донесли Йосафатові, говорячи: Прийшла на тебе сила силенна з того боку моря, з Сирії, і ось вони в Хаццон-Тамарі, воно Ен-Ґеді.
2CHR|20|3|І злякався Йосафат, і постановив звернутися до Господа. І він проголосив піст на всю Юдею.
2CHR|20|4|І зібралися юдеяни просити допомоги від Господа, також поприходили зо всіх Юдиних міст просити Господа.
2CHR|20|5|І став Йосафат у зборі Юдиному та єрусалимському в Господньому домі, перед новим подвір'ям,
2CHR|20|6|та й сказав: Господи, Боже батьків наших! Чи ж не Ти Бог на небесах? І Ти пануєш над усіма царствами народів, і в руці Твоїй сила та міць, і немає такого, хто б став проти Тебе!
2CHR|20|7|Чи ж не Ти, Боже наш, повиганяв мешканців цього Краю перед народом Твоїм, Ізраїлем, і дав його Авраамовому насінню, Твоєму приятелеві навіки?
2CHR|20|8|І вони осілися в ньому, і збудували Тобі в ньому святиню для Ймення Твого, говорячи:
2CHR|20|9|Якщо прийде на нас зло, меч укарання, чи моровиця, чи голод, то ми станемо перед цим храмом та перед лицем Твоїм, бо Ім'я Твоє в цьому храмі, і будемо кликати до Тебе з нашого утиску, і Ти почуєш, і спасеш.
2CHR|20|10|А тепер ось сини Аммонові й Моавові та мешканці гори Сеїр, що через них Ти не дав ізраїльтянам іти, коли вони виходили були з єгипетського краю, і вони минули їх, і не вигубили їх,
2CHR|20|11|і оце вони відплачують нам навалою, щоб вигнати нас із спадку Твого, який Ти віддав нам.
2CHR|20|12|Боже наш, чи ж Ти не осудиш їх? Нема бо в нас сили перед цією силою силенною, що приходить на нас, і ми не знаємо, що зробимо, бо наші очі на Тебе!
2CHR|20|13|А всі юдеяни стояли перед Господнім лицем, також діти їхні, жінки їхні та їхні сини.
2CHR|20|14|А Яхазіїл, син Захарія, сина Бенаї, Єіїла, сина Маттанії, Левит із Асафових синів, був на ньому Дух Господній серед збору,
2CHR|20|15|і він сказав: Послухайте, ввесь Юдо й мешканці Єрусалиму та царю Йосафате! Так говорить до вас Господь: Не бійтеся та не жахайтеся перед цією силенною силою, бо не ваша ця війна, але Божа!
2CHR|20|16|Узавтра зійдіть на них, ось вони входять збіччям Ціцу, і ви їх знайдете на кінці долини, навпроти пустині Єруїл.
2CHR|20|17|Не вам воювати в цьому, поставтеся й станьте, і побачите, що Господнє спасіння з вами, Юдо й Єрусалиме! Не бійтеся й не жахайтеся, узавтра виходьте перед них, а Господь буде з вами!
2CHR|20|18|І вклонився Йосафат обличчям до землі, а ввесь Юда та мешканці Єрусалиму попадали перед Господнім лицем, щоб уклонитися Господеві.
2CHR|20|19|І встали Левити з синів Кегатівців та з синів Корахівців, щоб хвалити Господа, Бога Ізраїлевого сильним голосом, високим.
2CHR|20|20|І повставали вони рано вранці, і вийшли до пустині Текоя. А як вони виходили, став Йосафат та й сказав: Послухайте мене, Юда та мешканці Єрусалиму! Віруйте в Господа, вашого Бога, і будете запевнені, вірте пророкам Його, і пощаститься вам!
2CHR|20|21|І радився він з народом, і поставив співаків для Господа, і вони хвалили величність святости, коли йшли перед озброєними, і говорили: Дякуйте Господу, бо навіки Його милосердя!
2CHR|20|22|А того часу, коли зачали вони співати та хвалити, дав Господь засідку на синів Аммонових і Моавових та на мешканців гори Сеїр, що прийшли були проти Юди, і були вони побиті,
2CHR|20|23|бо повстали аммонітяни та моавітяни на мешканців гори Сеїр, щоб учинити їх закляттям, і щоб вигубити. А коли вони покінчили це з мешканцями Сеїру, стали помагати один проти одного, щоб вигубити себе.
2CHR|20|24|І коли Юда прийшов на вартівню до пустині, і поглянули вони на натовп, аж ось трупи, що попадали на землю, і не було урятованого!
2CHR|20|25|І прийшов Йосафат та народ його, щоб пограбувати їхню здобич, і знайшли серед них дуже багато і маєтку, і одежі, і коштовностей, і понабирали собі стільки, що не могли нести. І вони три дні все грабували ту здобич, бо численна була вона!
2CHR|20|26|А четвертого дня зібралися вони до долини Бераха, бо там благословляли Господа; тому назвали ім'я тому місцю: долина Бераха, і так воно зветься аж до сьогодні.
2CHR|20|27|І вернулися всі юдеяни та єрусалимляни, а Йосафат на чолі їх, щоб вернутися до Єрусалиму з радістю, бо звеселив їх Господь спасінням від їхніх ворогів.
2CHR|20|28|І прибули вони до Єрусалиму з арфами й з цитрами та сурмами до Господнього дому.
2CHR|20|29|І був Божий страх на всі царства країв, коли вони почули, що Господь воював з Ізраїлевими ворогами...
2CHR|20|30|І заспокоїлося Йосафатове царство, і дав йому його Бог мир навколо.
2CHR|20|31|І царював Йосафат над Юдою. Він був віку тридцяти й п'яти років, коли зацарював, а двадцять і п'ять літ царював в Єрусалимі. А ім'я його матері Азува, дочка Шілхи.
2CHR|20|32|І ходив він дорогою свого батька Аси, і не уступався з неї, щоб робити вгодне в Господніх очах.
2CHR|20|33|Тільки пагірки не минулися, і народ іще не вчинив свого серця міцним для Бога своїх батьків.
2CHR|20|34|А решта Йосафатових діл, перші й останні, ото вони описані в записах Єгу, сина Ханані, що внесене до книги Ізраїлевих царів.
2CHR|20|35|А по тому поєднався Йосафат, цар Юдин, з Ахазією, Ізраїлевим царем, що робив несправедливо.
2CHR|20|36|І поєднався він із ним, щоб поробити кораблі, щоб ходити до Таршішу. І поробили вони кораблі в Ецйон-Ґевері.
2CHR|20|37|Та Елієзер, син Додави, з Мареші, пророкував на Йосафата, говорячи: За те, що ти поєднався з Ахазією, поруйнував Господь чини твої! І порозбивалися ті кораблі, і не могли йти до Таршішу...
2CHR|21|1|І спочив Йосафат із своїми батьками. І був він похований із своїми батьками в Давидовому Місті, а замість нього зацарював син його Єгорам.
2CHR|21|2|І були в нього брати, Йосафатові сини: Азарія, і Єхіїл, і Захарій, і Азарія, і Михаїл, і Шефатія, усі вони сини Йосафата, Ізраїлевого царя.
2CHR|21|3|І дав їм їхній батько великі подарунки срібла, і золота, і коштовності з твердинними містами в Юді, а царство дав Єгорамові, бо він первороджений.
2CHR|21|4|І став Єгорам на царстві батька. І зміцнився він, і позабивав усіх братів своїх мечем, а також декого з Ізраїлевих зверхників.
2CHR|21|5|Єгорам був віку тридцяти й двох літ, коли зацарював, і царював вісім літ в Єрусалимі.
2CHR|21|6|І ходив він дорогою Ізраїлевих царів, як робив Ахавів дім, бо Ахавова дочка була йому за жінку. І робив він зло в Господніх очах.
2CHR|21|7|Та не хотів Господь погубити Давидів дім ради заповіту, що склав був із Давидом, і як говорив дати світильника йому та синам його по всі дні.
2CHR|21|8|За його днів відпав був Едом з-під Юдиної руки, і настановили над собою царя.
2CHR|21|9|І пішов Єгорам зо своїми зверхниками, і всі колесниці з ним. І сталося, що він устав уночі та й побив Едома, що оточив був його, та зверхників колесниць.
2CHR|21|10|І відпав Едом з-під Юдиної руки, і так є аж до цього дня. Тоді того часу відпала й Лівна з-під руки його, бо він покинув Господа, Бога своїх батьків.
2CHR|21|11|Також він наробив пагірків по Юдиних містах, і вчинив перелюбами єрусалимських мешканців, а Юду звів.
2CHR|21|12|І прийшов до нього лист від пророка Іллі такого змісту: Так говорить Господь, Бог Давида, твого батька: За те, що не ходив ти дорогами Йосафата, свого батька, і дорогами Аси, Юдиного царя,
2CHR|21|13|а ходив дорогою Ізраїлевого царя, і вчинив перелюбниками Юду та мешканців Єрусалиму, як чинив перелюбниками дім Ахавів, а також братів своїх, дім свого батька, ліпших від тебе, ти позабивав,
2CHR|21|14|то ось ударить Господь великою поразою в народі твоїм, і в синах твоїх, і в жінках твоїх, і в усьому маєтку твоєму.
2CHR|21|15|А ти будеш у великих хворобах, у хворобі нутра свого, аж вийдуть нутрощі твої через довгочасну хворобу.
2CHR|21|16|І збудив Господь на Єгорама духа филистимлян та арабів, що при етіопах.
2CHR|21|17|І вийшли вони на Юду, і ввірвалися до нього, і позабирали ввесь маєток, що знаходився в царському домі, а також синів його та жінок його. І не позосталося в нього сина, окрім Єгоахаза, наймолодшого з синів його.
2CHR|21|18|А по всьому тому вдарив його Господь у нутрощах його невидужною хворобою.
2CHR|21|19|І сталося по певному часі, коли надійшов кінець двох років, вийшли його нутрощі від хвороби його, і він помер у тяжких болях. А народ його не зробив для нього спалення пахощів, як робили спалення батькам його.
2CHR|21|20|Він був віку тридцяти й двох літ, коли зацарював, а царював вісім літ в Єрусалимі. І відійшов він, і ніхто за ним не жалував; і поховали його в Давидовому Місті, та не в царських гробах.
2CHR|22|1|А мешканці Єрусалиму настановили царем замість нього Ахазію, його найменшого сина, бо всіх перших позабивала та ватага, що приходила з арабами на табір. І зацарював Ахазія, син Єгорама, Юдиного царя.
2CHR|22|2|Ахазія був віку сорока й двох літ, коли зацарював, і царював він в Єрусалимі один рік. А ім'я його матері Аталія, дочка Омрієва.
2CHR|22|3|Також він ходив дорогою Ахавого дому, бо його мати була йому дорадниця, щоб чинити беззаконня.
2CHR|22|4|І чинив він зло в Господніх очах, як Ахавів дім, бо вони були йому дорадниками по смерті його батька, на погибіль йому.
2CHR|22|5|Також за їхньою порадою він ходив. І пішов він з Єгорамом, сином Ахава, Ізраїлевого царя, на війну на Хазаїла, сирійського царя, в ґілеадський Рамот. І побили сиріяни Йорама.
2CHR|22|6|І вернувся він лікуватися в Їзреелі від тих ран, що завдали йому в Рамі, як він воював із Хазаїлом, сирійським царем. А Азарія, Єгорамів син, цар Юдин, зійшов побачити Єгорама, Ахавого сина, в Їзреелі, бо він був слабий.
2CHR|22|7|І від Бога було на погибіль Ахазії, щоб прийти до Єгорама, бо як прийшов, вийшов з Єгорамом на Єгу, сина Німші, що Господь помазав його вигубити Ахавів дім.
2CHR|22|8|І сталося, коли Єгу чинив суд над Ахавовим домом, то знайшов він Юдиних зверхників та синів Ахазієвих братів, що служили Ахазієві, і позабивав їх.
2CHR|22|9|І відшукав він Ахазію, і схопили його, а він ховався в Самарії. І привели його до Єгу та й забили його; і поховали його, бо сказали: Він син Йосафата, що всім серцем своїм звертався до Господа. І не було в домі Ахазії нікого, хто мав би силу царювати.
2CHR|22|10|А коли Аталія, мати Ахазії, побачила, що помер її син, то встала й вигубила все цареве насіння Юдиного дому...
2CHR|22|11|А Єгосав'ат, дочка царя, взяла Йоаша, сина Ахазії, та й викрала його з-поміж вбиваних царських синів, і дала його та няньку його до спальної кімнати. І сховала його Єгосав'ат, дочка царя Єгорама, жінка священика Єгояди, бо вона була сестра Ахазії, перед Аталією, і та не забила його.
2CHR|22|12|І він був з ними в Божому домі, ховаючися шість років, а Аталія царювала над Краєм.
2CHR|23|1|А сьомого року зміцнився Єгояда й прийняв сотників: Азарію, Єрохамового сина, і Ізмаїла, сина Єгохананового, і Азарію, сина Оведового, і Маасею, сина Адаї, і Елісафата, сина Зіхрієвого, в умову з собою.
2CHR|23|2|І обійшли вони Юду, і зібрали зо всіх Юдиних міст Левитів та голів Ізраїлевих домів, і прийшли до Єрусалиму.
2CHR|23|3|І ввесь збір склав у Божому домі умову з царем. І сказав їм Єгояда: Оце царський син буде царювати, як говорив Господь про Давидових синів.
2CHR|23|4|Оце та річ, яку зробите: третина з вас, що приходите в суботу, із священиків та з Левитів, будете за придверних біля порогів.
2CHR|23|5|А третина при царському домі, а третина при брамі Єсод, а ввесь народ у подвір'ях Господнього дому.
2CHR|23|6|І нехай не входить до Господнього йому ніхто, окрім священиків та тих, хто прислуговує із Левитів, вони ввійдуть, бо освячені вони, а ввесь народ буде пильнувати Господньої сторожі.
2CHR|23|7|І оточать Левити царя навколо, кожен із своєю зброєю в руці своїй; а хто чужий увійшов би до дому, нехай буде забитий! І будете ви з царем при вході його та при виході його.
2CHR|23|8|І зробили Левити та ввесь Юда все, що наказав священик Єгояда. І взяли кожен людей своїх, що приходять у суботу та відходять у суботу, бо священик Єгояда не звільнив черг.
2CHR|23|9|І дав священик Єгояда сотникам ратища, і малі щити, і інші щити, що належали цареві Давидові, що були в Божому домі.
2CHR|23|10|І поставив він увесь народ, а кожен мав свою зброю в руці своїй, від правого боку дому аж до лівого боку дому, при жертівнику та при домі, навколо біля царя.
2CHR|23|11|І вивели вони царського сина, і поклали на нього корону та звої Закону. І зробили вони його царем, і помазали його Єгояда та сини його, та й крикнули: Нехай живе цар!
2CHR|23|12|І почула Аталія голос народу, що бігав та славив царя, і прийшла до народу до Господнього дому.
2CHR|23|13|І побачила вона, аж ось цар стоїть на помості своїм при вході, а при царі зверхники та сурми, а ввесь народ Краю радіє та сурмить у сурми, а співаки з музичними знаряддями, що подавали до відома знаки на хвалу. І роздерла Аталія шати свої та й крикнула: Змова, змова!
2CHR|23|14|А священик Єгояда наказав сотникам, поставленим над військом, і сказав до них: Виведіть її поміж шереги, а хто інший піде за нею, нехай буде забитий мечем! Бо священик сказав: Не заб'єте її в Господньому домі!
2CHR|23|15|І зробили їй прохід, і вона вийшла входом Кінської брами до царського дому, і там забили її.
2CHR|23|16|І склав Єгояда умову між собою й між усім народом та між царем, щоб бути народом Господнім.
2CHR|23|17|І ввійшов увесь народ до Ваалового дому, та й порозбивали його та жертівники його, і бовванів його зовсім поламали, а Маттана, Ваалового священика, убили перед жертівниками.
2CHR|23|18|А в Господньому домі Єгояда віддав уряди на руку священиків та Левитів, яких поділив Давид над Господнім домом, щоб приносити Господні цілопалення, як написано в Мойсеєвім Законі, з радістю та зо співом, за уставом Давидовим.
2CHR|23|19|А при брамах Господнього дому поставив він придверних, щоб не ввійшов хто будь-чим нечистий.
2CHR|23|20|І взяв він сотників, і вельмож, і тих, що старшинують над народом, та ввесь народ Краю, і відвели царя з Господнього дому. І ввійшли вони через горішню браму до царського дому, і посадили царя на троні царства.
2CHR|23|21|І радів увесь народ Краю, а місто заспокоїлося. А Аталію вбили мечем.
2CHR|24|1|Йоаш був віку семи років, коли зацарював, і сорок років царював він в Єрусалимі. А ім'я його матері Цівія, з Беер-Шеви.
2CHR|24|2|І робив Йоаш вгодне в Господніх очах по всі дні священика Єгояди.
2CHR|24|3|І взяв йому Єгояда дві жінки, а той породив синів та дочок.
2CHR|24|4|І сталося по тому, було в Йоашевому серці відновити Господній дім.
2CHR|24|5|І зібрав він священиків та Левитів, і сказав до них: Підіть по Юдиних містах, і збирайте з усього Ізраїля срібло на направу храму вашого Бога рік-річно, і ви будете спішити в цій справі! Та не спішилися Левити.
2CHR|24|6|І покликав цар Єгояду, голову священиків, і сказав до нього: Чому ти не жадаєш від Левитів, щоб приносили з Юди та з Єрусалиму дарунки, за постановою Мойсея, раба Господнього, та Ізраїлевого збору на скинію свідоцтва?
2CHR|24|7|Бо сини нечестивої Аталії вломилися були до Божого дому, і всі святощі Господнього дому вжили для Ваалів.
2CHR|24|8|І сказав цар, і зробили одну скриньку, і поставили її в брамі Господнього дому назовні.
2CHR|24|9|І проголосили в Юді та в Єрусалимі приносити для Господа даток, що його встановив на Ізраїля в пустині Мойсей, Божий раб.
2CHR|24|10|І раділи всі зверхники та ввесь народ, і приносили й кидали до скриньки, аж поки вона наповнилася.
2CHR|24|11|І бувало того часу, коли Левити приносили скриньку на царський перегляд, і як вони бачили, що численне те срібло, то приходив царський писар та призначений від священика-голови, і вони випорожнювали скриньку. Потім відносили її, і повертали її на її місце. Так робили вони день-у-день, і зібрали дуже багато срібла.
2CHR|24|12|А цар та Єгояда давали його тим, що робили працю роботи Господнього дому, і все наймали каменярів та теслів, щоб відновлювати дім Господній, а також тим, що обробляли залізо та мідь на зміцнення Господнього дому.
2CHR|24|13|І працювали робітники, і чинилася направа працею їхньої руки. І поставили вони Божий дім на міру його, і зміцнили його.
2CHR|24|14|А коли покінчили, вони принесли перед царя та Єгояду решту срібла. І поробили вони з нього речі для Господнього дому, речі для служби та для жертвоприношення, і ложки, і посуд золотий та срібний. І приносили цілопалення в Господньому домі завжди, по всі дні Єгояди.
2CHR|24|15|І постарів Єгояда, і наситився днями й помер. Він був віку ста й тридцяти літ, коли помер.
2CHR|24|16|І поховали його в Давидовому Місті з царями, бо робив він добро в Ізраїлі і для Бога, і для Його храму.
2CHR|24|17|А по Єгоядиній смерті прийшли князі Юдині, і поклонилися цареві. Тоді цар їх послухав.
2CHR|24|18|І покинули вони дім Господа, Бога своїх батьків, та й служили Астартам та божкам. І був Божий гнів на Юду та Єрусалим за цю їхню провину.
2CHR|24|19|І послав Він між них пророків, щоб привернути їх до Господа, і вони свідчили проти них, та ті не слухались.
2CHR|24|20|А Дух Господній огорнув Захарія, сина священика Єгояди, і він став перед народом та й сказав до них: Так сказав Бог: Чому ви переступаєте Господні заповіти? Ви не матимете успіху, бо ви покинули Господа, то й Він покинув вас!...
2CHR|24|21|І змовилися вони на нього, і закидали його камінням з царського наказу в подвір'ї Господнього дому...
2CHR|24|22|І не пам'ятав цар Йоаш тієї милости, яку зробив був із ним батько того Єгояда, але вбив сина його. А як той умирав, то сказав: Нехай побачить Господь, і нехай покарає!...
2CHR|24|23|І сталося наприкінці року, прийшло на нього сирійське військо, і прибули до Юди та до Єрусалиму, і позабивали всіх зверхників народу, а всю здобич із них послали цареві в Дамаск.
2CHR|24|24|Хоч з малою кількістю людей прийшло сирійське військо, проте Господь дав в їхню руку дуже велику силу, бо ті покинули Господа, Бога батьків своїх. А над Йоашем вони виконали присуд.
2CHR|24|25|А коли вони відійшли від нього, позоставивши його в тяжких хворобах, змовилися на нього його раби за кров синів священика Єгояди, і забили його на ліжку його, і він помер... І поховали його в Давидовому Місті, та не поховали його в гробах царських.
2CHR|24|26|А оце змовники на нього: Завад, син аммонітянки Шім'ат, і Єгозавад, син моавітянки Шімріт.
2CHR|24|27|А сини його, і великість тягару, покладеного на нього, і відбудова Божого дому, ото вони описані в викладі Книги Царів. А замість нього зацарював син його Амація.
2CHR|25|1|У віці двадцяти й п'яти літ зацарював Амація, і двадцять і п'ять літ царював він в Єрусалимі. А ім'я його матері Єгоаддан, з Єрусалиму.
2CHR|25|2|І робив він угодне в Господніх очах, тільки не з цілим серцем.
2CHR|25|3|І сталося, як зміцнилося царство за ним, то він повбивав своїх рабів, що забили царя свого, його батька.
2CHR|25|4|А синів їх він не позабивав, як написано в книзі Мойсеєвого Закону, що наказав був Господь, говорячи: Не помруть батьки за синів, а сини не помруть за батьків, бо кожен за гріх свій помре.
2CHR|25|5|І зібрав Амація Юду, і поставив їх за домом їхніх батьків, за тисячниками та за сотниками для всього Юди та Веніямина; і він перелічив їх від віку двадцяти років і вище, і знайшов їх три сотні тисяч вибраного, здатного до війська, хто тримає ратище та великого щита.
2CHR|25|6|І найняв він із Ізраїля сотню тисяч хоробрих вояків за сотню талантів срібла.
2CHR|25|7|І прийшов до нього Божий чоловік, говорячи: О царю, нехай не виходить з тобою Ізраїлеве військо, бо Господь не з Ізраїлем, ні з жодним із синів Єфрема.
2CHR|25|8|Але йди тільки ти, роби, будь відважний на війні! Інакше вчинить Бог, що ти спіткнешся перед ворогом, бо в Бога є сила допомагати, або робити, щоб спіткнутися.
2CHR|25|9|І сказав Амація до Божого чоловіка: А що робити з тією сотнею талантів, що я дав Ізраїлевому війську? А Божий чоловік відказав: Господь може дати тобі більше від цього!
2CHR|25|10|І відділив Амація їх, те військо, що прийшло з краю Єфремового, щоб ішло на своє місце. І дуже запалився їхній гнів на Юду, і вони вернулися на своє місце в запаленому гніві.
2CHR|25|11|А Амація зміцнився, і попровадив свій народ, і пішов до Соляної долини, і побив десять тисяч Сеїрових синів,
2CHR|25|12|а десять тисяч живих узяли Юдині сини до неволі. І привели їх на верхів'я скелі, і поскидали їх з верхів'я тієї скелі, і всі вони позабивалися...
2CHR|25|13|А люди того війська, що Амація вернув, щоб не йшли з ним на війну, розсипалися по Юдиних містах від Самарії й аж до Бет-Хорону, і повбивали з них три тисячі, і пограбували велику здобич.
2CHR|25|14|І сталося по тому, як прийшов Амація, побивши едомлян, то він приніс богів Сеїрових синів, і поставив їх собі за богів, і перед ними вклонявся, і їм кадив.
2CHR|25|15|І запалився Господній гнів на Амацію, і Він послав до нього пророка, а той сказав йому: Нащо ти звертався до богів цього народу, богів, що не врятували народу свого від твоєї руки?
2CHR|25|16|І сталося, як він говорив це до нього, сказав йому цар: Чи я поставив тебе за царевого дорадника? Перестань собі, нащо вбивати тебе? І перестав той пророк, але сказав: Я знаю, що Бог постановив погубити тебе, бо зробив ти це, і не слухав моєї поради...
2CHR|25|17|І радився Амація, цар Юдин, і послав до Йоаша, сина Єгоахаза, сина Єгу, Ізраїлевого царя, говорячи: Іди но, поміряємось!
2CHR|25|18|І послав Йоаш, Ізраїлів цар, до Амації, Юдиного царя, говорячи: Тернина, що на Ливані, послала до кедрини, що на Ливані, кажучи: Дай но дочку свою моєму синові за жінку! Та перейшла польова звірина, що на Ливані, і витоптала ту тернину...
2CHR|25|19|Ти сказав: Ось побив ти Едома, і піднесло тебе серце твоє, щоб пишатися. Тепер сиди ж у своєму домі. Нащо будеш дрочитися зо злом, і впадеш ти та Юда з тобою?
2CHR|25|20|Та не послухався Амація, бо від Бога було це, щоб віддати їх у руку ворога, бо зверталися вони до едомських богів.
2CHR|25|21|І вийшов Йоаш, Ізраїлів цар, і зустрілися він та Амація, цар Юдин, у Юдиному Бет-Шемеші.
2CHR|25|22|І був побитий Юда перед Ізраїлем, і повтікали кожен до намету свого.
2CHR|25|23|А Йоаш, цар Ізраїлів, схопив Амацію, Юдиного царя, сина Йоаша, сина Єгоахаза, у Бет-Шемеші, і привів його до Єрусалиму, і зробив пролім в єрусалимському мурі, від Єфремової брами аж до брами Наріжної, чотири сотні ліктів.
2CHR|25|24|І забрав він усе золото й срібло, та ввесь посуд, що знаходився в Божому домі в Овед-Едома, та скарби царевого дому, та закладників, і вернувся в Самарію.
2CHR|25|25|І жив Амація, Йоашів син, цар Юдин, по смерті Йоаша, Єгоахазового сина, Ізраїлевого царя, п'ятнадцять літ.
2CHR|25|26|А решта діл Амації, перші та останні, ото вони написані в Книзі Царів Юдиних та Ізраїлевих.
2CHR|25|27|А від часу, коли Амація відступив від Господа, то склали на нього змову в Єрусалимі, та він утік до Лахішу. І послали за ним до Лахішу, і вбили його там.
2CHR|25|28|І повезли його на конях, і поховали його з батьками його в Давидовому Місті.
2CHR|26|1|І взяв увесь Юдин народ Уззійю, а він був шістнадцяти літ, і настановили його царем замість батька його Амації.
2CHR|26|2|Він збудував Елота, і вернув його Юді, як цар спочив зо своїми батьками.
2CHR|26|3|Уззійя був віку шістнадцяти літ, коли він зацарював, а п'ятдесят і два роки царював в Єрусалимі. А ім'я його матері Єхолія, з Єрусалиму.
2CHR|26|4|І робив він угодне в Господніх очах, усе, що робив батько його Амація.
2CHR|26|5|І став він звертатися до Бога за днів Захарія, що розумів Божі видіння. А за днів, коли він звертався до Господа, Бог давав йому успіх.
2CHR|26|6|І він вийшов, і воював із филистимлянами, і поруйнував мур міста Ґату, і мур Явне, і мур Асдоду, і побудував міста в Асдоді та в филистимлян.
2CHR|26|7|І допоміг йому Бог над филистимлянами, і над арабами, що живуть у Ґур-Баалі, та над мецнітами.
2CHR|26|8|І давали аммонітяни данину для Уззійї, а ім'я його пронеслося аж туди, де йдеться до Єгипту, бо він сильно зміцнився.
2CHR|26|9|І збудував Уззійя башту в Єрусалимі над брамою Пінна, і над брамою Ґай, і над Мікцоа, і позміцнював їх.
2CHR|26|10|І побудував він башти в пустині, і повисікував багато ям для води, бо мав великі череди і на долині, і на рівнині, рільників, і виноградарів у горах, і садки, бо він любив хліборобство.
2CHR|26|11|І було в Уззійї військо, що провадило війну, яке виходило на війну відділом за числом їхнього переліку через писаря Єіїла та урядника Маасею, під рукою Хананії з царевих зверхників.
2CHR|26|12|Усе число голів батьківських родів, хоробрих вояків, дві тисячі й шість сотень.
2CHR|26|13|А при них війська, три сотні тисяч і сім тисяч і п'ять сотень тих, що провадять війну великою силою, щоб допомагати цареві на ворога.
2CHR|26|14|І наготовив для них Уззійя для всього війська щити малі й ратища, і шоломи, і панцери, і луки, і пращного каміння.
2CHR|26|15|І наробив він в Єрусалимі військових машин, майстерно придуманих, щоб були вони на баштах і на рогах на стріляння стрілами та великим камінням. І пронеслося ім'я його аж надто далеко, бо він дивно зробив, щоб допомогти собі, так що став сильним.
2CHR|26|16|А як він зміцнів, запишалося його серце аж до зіпсуття, і він спроневірився Господеві, Богові своєму. І ввійшов він до храму Господнього, щоб кадити на кадильному жертівнику.
2CHR|26|17|А за ним пішов священик Азарія, а з ним Господні священики, вісімдесят хоробрих мужів.
2CHR|26|18|І стали вони проти царя Узійї та й сказали йому: Не тобі, Уззійє, кадити для Господа, а священикам, синам Аароновим, посвяченим на кадіння... Вийди зо святині, бо ти спроневірився, і не за честь це буде тобі від Господа Бога!
2CHR|26|19|І розгнівався Уззійя, а в руці його була кадильниця на кадіння. А коли він розгнівався на священиків, то на чолі його показалася проказа, перед священиками в Господньому домі, при кадильному жертівнику...
2CHR|26|20|І глянув на нього первосвященик Азарія та всі священики, аж ось він прокажений на чолі своїм! І вони поспішно вигнали його звідти, та й сам він поспішив вийти, бо вразив його Господь!
2CHR|26|21|І був цар Уззійя прокажений аж до дня своєї смерти, і сидів в осібному домі прокажений, бо був вилучений від Господнього дому. А над царським домом був син його Йотам, він судив народ Краю.
2CHR|26|22|А решту діл Уззійї, перші й останні, описав пророк Ісая, син Амосів.
2CHR|26|23|І спочив Уззійя з своїми батьками, і поховали його з батьками його на погребовому царському полі, бо сказали: Він прокажений. А замість нього зацарював син його Йотам.
2CHR|27|1|Йотам був віку двадцяти й п'яти років, коли зацарював, і шістнадцять літ царював в Єрусалимі. А ім'я його матері Єруша, Садокова дочка.
2CHR|27|2|І робив він угодне в Господніх очах, усе, що робив був його батько Уззійя. Тільки він не входив до Господнього храму, та народ іще грішив.
2CHR|27|3|Він збудував горішню браму Господнього дому, і багато побудував на мурі Офел.
2CHR|27|4|І побудував він міста в Юдиних горах, а в лісах побудував твердині та башти.
2CHR|27|5|І він воював з царем аммонітян, і був сильніший від них. І дали йому аммонітяни того року сотню талантів срібла, і десять тисяч корів пшениці та десять тисяч ячменю. Це давали йому аммонітяни й року другого та третього.
2CHR|27|6|І став сильний Йотам, бо поправив дороги свої перед лицем Господа, Бога свого.
2CHR|27|7|А решта Йотамових діл, і всі війни його та дороги його, ось вони описані в Книзі Царів Ізраїлевих та Юдиних.
2CHR|27|8|Він був віку двадцяти й п'яти літ, коли зацарював, і шістнадцять літ царював в Єрусалимі.
2CHR|27|9|І спочив Йотам із своїми батьками, і поховали його в Давидовому Місті, а замість нього зацарював син його Ахаз.
2CHR|28|1|Ахаз був віку двадцяти літ, коли він зацарював, і шістнадцять літ царював в Єрусалимі.
2CHR|28|2|І ходив він дорогами Ізраїлевих царів, а також робив литих бовванів Ваалів.
2CHR|28|3|І він кадив у долині Бен-Гіннома, і палив своїх синів огнем за гидотами тих народів, що Господь повиганяв їх перед Ізраїлевими синами.
2CHR|28|4|І він приносив жертви та кадив на пагірках і на висотах, та під кожним зеленим деревом.
2CHR|28|5|І дав його Господь, Бог його, в руку сирійського царя, і вони повбивали з його війська та взяли до неволі від нього багатьох полонених, і спровадили до Дамаску. Крім того, він був виданий і в руку Ізраїлевого царя, і той уразив його великою поразою.
2CHR|28|6|І побив Пеках, син Ремалії, в Юді сто й двадцять тисяч одного дня, все мужів хоробрих, за те, що залишили вони Господа, Бога їхніх батьків.
2CHR|28|7|А Зіхрі, лицар Єфремів, забив Маасею, царського сина, й Азрікама, володаря дому, й Елкану, другого по царі.
2CHR|28|8|І Ізраїлеві сини взяли до неволі зо своїх братів двісті тисяч жінок, синів та дочок, а також пограбували від них велику здобич, і спровадили ту здобич до Самарії.
2CHR|28|9|А там був Господній пророк, Одед ім'я йому. І він вийшов перед військо, що входило до Самарії, та й сказав їм: Ось Господь, Бог ваших батьків, у гніві на Юду, віддав їх у вашу руку, а ви повибивали між ними з лютістю, яка досягла аж до небес.
2CHR|28|10|А тепер ви задумуєте здобути собі за рабів та за невільниць дітей Юди та Єрусалиму. Чи ж за вами самими нема провин проти Господа, Бога вашого?
2CHR|28|11|Отож, послухайте мене тепер, і верніть тих полонених, яких взяли ви до неволі з ваших братів, бо на вас ревність Господнього гніву!
2CHR|28|12|І встали дехто з голів Єфремових синів: Азарія, син Єгоханана, Берехія, син Мешіллемотів, і Єхізкійя, син Шаллумів, і Амаса, син Хадлаїв, проти тих, що приходили з війська,
2CHR|28|13|та й сказали до них: Не приводьте цих полонених сюди, бо на провину нам проти Господа ви задумуєте додати це до наших гріхів та до нашої провини. Бо велика наша провина та жар гніву Господнього на Ізраїля!
2CHR|28|14|І озброєні покинули тих полонених та ту здобич перед зверхниками та всім збором.
2CHR|28|15|І встали ті мужі, що були означені іменами, і взяли полонених, і всіх їхніх нагих позодягали зо здобичі, і зодягнули їх, і обули їх, і нагодували їх, і напоїли їх, і намастили їх, і кожного слабого з них повезли на ослах. І припровадили їх до Єрихону, міста пальм, до їхніх братів, а самі вернулися до Самарії.
2CHR|28|16|Того часу послав цар Ахаз до асирійських царів, щоб допомогли йому.
2CHR|28|17|Прийшли ще й едомляни, і побили багатьох між Юдою, і взяли до неволі полонених.
2CHR|28|18|А филистимляни розсипалися по містах Шефелі та Юдиного Неґеву, і здобули Бет-Шемеш, і Айялон, і Ґедерот, і Сохо та залежні міста його, і Тімну та залежні міста її, і Ґімзо та залежні міста його, й осілися там.
2CHR|28|19|Бо Господь принизив Юду через Ахаза, Ізраїлевого царя, бо завільно поступав він щодо Юди, і спроневірився великим гріхом проти Господа.
2CHR|28|20|І прийшов на нього Тіґлат Пілнеесер, цар асирійський, й утискав його, і не допоміг йому.
2CHR|28|21|Бо Ахаз пограбував був Господній дім, і дім царів, і зверхників, і дав це асирійському цареві, та не було це на поміч йому.
2CHR|28|22|А в часі утиску його, то продовжував спроневірюватися Господеві він, той цар Ахаз.
2CHR|28|23|І приносив він жертви дамаським богам, що його побили, і говорив: Через те, що боги сирійських царів допомагають їм, то буду приносити їм жертви, вони будуть допомагати мені! А вони були йому на те, щоб спотикався він та ввесь Ізраїль!
2CHR|28|24|І Ахаз зібрав посуд Божого дому, і порубав посуд Божого дому. І позамикав він двері Господнього дому, і поробив собі жертівники в кожному куті в Єрусалимі...
2CHR|28|25|І в кожному місті Юдиному поробив він пагірки, щоб кадити іншим богам, і розгнівав Господа, Бога батьків своїх.
2CHR|28|26|А решта його діл та всі дороги його, перші й останні, ото вони описані в Книзі Царів Юдиних та Ізраїлевих.
2CHR|28|27|І спочив Ахаз зо своїми батьками, і поховали його в місті, в Єрусалимі, бо не внесли його до гробів Ізраїлевих царів, а замість нього зацарював син його Єзекія.
2CHR|29|1|Єзекія зацарював у віці двадцяти й п'яти літ, а двадцять і дев'ять літ царював він в Єрусалимі. А ім'я його матері Авійя, дочка Захарії.
2CHR|29|2|І робив він угодне в Господніх очах, як усе, що робив був його батько Давид.
2CHR|29|3|Він першого року свого царювання, місяця першого відчинив двері Господнього дому, і поправив їх.
2CHR|29|4|І привів він священиків та Левитів, і зібрав їх на східню площу,
2CHR|29|5|та й сказав їм: Послухайте мене, Левити! Освятіться тепер, і освятіть дім Господа, Бога ваших батьків, і винесіть нечисть із святині.
2CHR|29|6|Бо наші батьки спроневірилися, і робили лихе в очах Господа, Бога нашого, і залишили Його, і відвернули своє обличчя від Господньої скинії, й обернулися спиною до неї.
2CHR|29|7|Також замкнули вони двері притвору, і погасили лямпадки, а кадила не кадили, і цілопалення не приносили в святині для Ізраїлевого Бога.
2CHR|29|8|І був Господній гнів на Юду та на Єрусалим, і Він дав їх на ганьбу, і на спустошення, і на посміховище, як ви бачите своїми очима.
2CHR|29|9|І ось попадали наші батьки від меча, а наші сини, і наші дочки, і жінки наші в неволі за це!
2CHR|29|10|Тепер на моєму серці лежить скласти заповіта з Господом, Ізраїлевим Богом, і нехай Він відверне від нас жар гніву Свого.
2CHR|29|11|Сини мої, не будьте недбалі тепер, бо вас Господь вибрав ставати перед лицем Його на службу Йому, та щоб служити Йому й кадити Йому!
2CHR|29|12|І встали Левити: Махат, син Амасаїв, і Йоїл, син Азарії, від синів Кегатових; а від синів Мерарієвих: Кіш, син Авдіїв, і Азарія, син Єгаллел'їлів; а від Ґершонівців: Йоах, син Зіммин, і Еден, син Йоахів;
2CHR|29|13|а від синів Еліцафанових: Шімрі, і Єіїл; а від синів Асафових: Захарій та Маттанія.
2CHR|29|14|А від Геманових синів: Єхіїл, і Шім'ї; а від синів Єдутунових: Шемая та Уззіїл.
2CHR|29|15|І зібрали вони братів своїх, і освятилися, і пішли за наказом царським у справах Господніх, щоб очистити Господній дім.
2CHR|29|16|І повходили священики до середини Господнього дому на очищення. І повиносили вони всю нечистість, яку знайшли в Господньому храмі, до подвір'я Господнього дому, а Левити взяли це, щоб винести назовні до долини Кедрон.
2CHR|29|17|І зачали вони першого дня першого місяця освящати, а восьмого дня того місяця ввійшли до Господнього притвору. І освятили вони Господній дім за вісім день, а шістнадцятого дня першого місяця закінчили.
2CHR|29|18|І ввійшли вони в середину дому до царя Єзекії та й сказали: Очистили ми ввесь Господній дім, і жертівника цілопалення, та всі його речі, і стіл укладання хлібів та всі його речі.
2CHR|29|19|А всі ті речі, які цар Ахаз занехав був за свого царювання, коли спроневірився, ми приготовили та освятили, і ось вони перед Господнім жертівником.
2CHR|29|20|І встав рано цар Єзекія, і зібрав зверхників міста та й увійшов до Господнього дому.
2CHR|29|21|І привели вони сім биків, і сім баранів, і сім овечок, і сім козлів на жертву за гріх: за царство, і за святиню, і за Юду, а він звелів Аароновим синам, священикам, принести це в жертву на Господньому жертівнику.
2CHR|29|22|І порізали ту велику худобу, а священики прийняли кров і покропили на жертівника; і порізали баранів, і покропили ту кров на жертівника; і порізали овечок, і покропили ту кров на жертівника.
2CHR|29|23|І привели козлів жертви за гріх перед царя та збори, і вони поклали свої руки на них.
2CHR|29|24|І зарізали їх священики, а їхньою кров'ю очистили жертівника, щоб очистити всього Ізраїля, бо за всього Ізраїля звелів цар принести це цілопалення та цю жертву за гріх.
2CHR|29|25|І поставив він Левитів Господнього дому з цимбалами, з арфами та з цитрами, за наказом Давида та Ґада, царевого прозорливця, та пророка Натана, бо в руці Господа наказ, що йде через пророків Його.
2CHR|29|26|І поставали Левити з Давидовим знаряддям, а священики із сурмами.
2CHR|29|27|І сказав Єзекія принести цілопалення на жертівника. А коли розпочали цілопалення, зачався спів Господеві та звуки сурем і музичного знаряддя Давида, Ізраїлевого царя.
2CHR|29|28|І ввесь збір вклонився, і співаки співали, а сурми сурмили, це все аж до кінця цілопалення!
2CHR|29|29|А як скінчили приносити жертву, попадали навколішки цар та всі, що були з ним, і вклонилися.
2CHR|29|30|І сказав цар Єзекія та зверхники до Левитів, щоб вони хвалили Господа словами Давида та прозорливця Асафа, і вони хвалили з великою радістю, і схилялися, і вклонялися до землі.
2CHR|29|31|І відповів Єзекія й сказав: Тепер ви освячені для Господа. Підійдіть, і приведіть жертви та приноси вдячні для Господнього дому. І привів збір жертви та приноси вдячні, і кожен, хто мав жертвенне серце, приносив цілопалення.
2CHR|29|32|І було число цілопалення, що спровадив збір: худоби великої сімдесят, баранів сотня, овечок двісті, для цілопалення Господеві все це.
2CHR|29|33|А для святости: худоби великої шість сотень, а худоби дрібної три тисячі.
2CHR|29|34|Тільки священиків було мало, і не могли вони обдирати шкур зо всіх цілопалень; і допомагали їм їхні брати Левити аж до скінчення праці, і поки освятилися священики, бо Левити були простосердіші на освячення, аніж священики.
2CHR|29|35|І також було багато палень серед мирних жертов і серед жертов литих до цілопалення. І так була відновлена служба Господнього дому.
2CHR|29|36|І радів Єзекія та ввесь народ тим, що Бог приготовив для народу, бо та річ сталася несподівано!
2CHR|30|1|І послав Єзекія по всьому Ізраїлю та по Юдеї, а також написав листи до країв Єфрема та Манасії, щоб прийшли до Господнього дому в Єрусалимі, щоб справити Пасху для Господа, Ізраїлевого Бога.
2CHR|30|2|І радився цар і зверхники його та ввесь збір в Єрусалимі, щоб справити Пасху другого місяця.
2CHR|30|3|Бо не могли справити її того часу, бо священики не освятилися в потрібному числі, а народ не зібрався до Єрусалиму.
2CHR|30|4|І була вгодна та річ в очах царевих та в очах усього збору.
2CHR|30|5|І вони постановили оголосити по всьому Ізраїлю від Беер-Шеви й аж до Дана, щоб приходили справити Пасху для Господа, Ізраїлевого Бога, в Єрусалим, бо не часто робили її так, як написано.
2CHR|30|6|І пішли бігуни з листами від царя та його зверхників по всьому Ізраїлі та Юдеї, та за наказом царя говорили: Ізраїлеві сини, верніться до Господа, Бога Авраамового, Ісакового та Ізраїлевого, і Він повернеться до останку, позосталого вам із руки асирійських царів.
2CHR|30|7|І не будьте такі, як ваші батьки та як ваші брати, що спроневірилися Господеві, Богові їхніх батьків, і Він дав їх на спустошення, як ви бачите.
2CHR|30|8|Тепер не будьте твердошиї, як ваші батьки. Покоріться Господеві, і ввійдіть до святині Його, яку Він освятив навіки, і служіть Господеві, Богові вашому, і Він відверне від вас жар гніву Свого.
2CHR|30|9|Бо як ви навернетесь до Господа, то брати ваші та ваші сини знайдуть милосердя в своїх поневільників, і зможуть вернутися до цього Краю, бо милостивий і милосердний Господь, Бог ваш, і Він не відверне лиця від вас, якщо ви навернетеся до Нього.
2CHR|30|10|І сторожі все переходили з міста до міста по краю Єфремовому та Манасіїному й аж до Завулона. Та люди глузували з них, і висміювали їх.
2CHR|30|11|Тільки люди з Асира, і Манасії та з Завулона впокорилися, і поприходили до Єрусалиму.
2CHR|30|12|Також в Юдеї була Божа рука, щоб дати їм одне серце для виконання наказу царя та зверхників за Господнім словом.
2CHR|30|13|І зібрався до Єрусалиму численний народ, щоб справити свято Опрісноків другого місяця, збір дуже численний.
2CHR|30|14|І встали вони, і повикидали ідольські жертівники, що були в Єрусалимі, і повикидали всі кадильниці, та й повкидали до долини Кедрон.
2CHR|30|15|І зарізали пасхальне ягня чотирнадцятого дня другого місяця, а священики та Левити засоромилися й освятилися, і принесли цілопалення до Господнього дому.
2CHR|30|16|І поставали вони на своєму місці за їхнім правом, за Законом Мойсея, чоловіка Божого. Священики кропили кров, беручи з руки Левитів.
2CHR|30|17|Багато бо було в зборі, що не освятилися, тому Левити були для різання пасхальних ягнят за кожного нечистого, щоб посвятити для Господа.
2CHR|30|18|Бо безліч народу, багато з Єфрема та Манасії, Іссахара та Завулона не очистилися, але їли Пасху, не так, як написано. Та Єзекія молився за них, говорячи: Добрий Господь простить кожному,
2CHR|30|19|хто все своє серце міцно встановив, щоб звертатися до Бога, Господа, Бога батьків своїх, хоч не зробив він за правилами чистости святині.
2CHR|30|20|І послухав Господь Єзекію, і простив народ.
2CHR|30|21|І справляли Ізраїлеві сини, що знаходилися в Єрусалимі, свято Опрісноків сім день з великою радістю, а Левити та священики день-у-день славили Господа всією силою.
2CHR|30|22|І промовляв Єзекія до серця всіх Левитів, що мали добре розуміння для Господа. І їли святкову жертву сім день, і приносили мирні жертви, і сповідалися Господеві, Богові батьків своїх.
2CHR|30|23|І ввесь збір нарадився справити свято ще другі сім день, і справляли сім день в радості.
2CHR|30|24|Бо Єзекія, цар Юдин, дав для збору тисячу биків і сім тисяч худоби дрібної, а зверхники дали для збору тисячу биків і десять тисяч худоби дрібної. І освятилося багато священиків.
2CHR|30|25|І радів увесь Юдин збір, і священики та Левити, і ввесь збір, що прийшов з Ізраїля, і приходьки, що поприходили з Ізраїлевого Краю, та ті, що сиділи в Юдеї.
2CHR|30|26|І була велика радість в Єрусалимі, бо від днів Соломона, Давидового сина, Ізраїлевого царя, не було такого, як оце в Єрусалимі!
2CHR|30|27|І встали священики та Левити, і поблагословили народ. І почутий був їхній голос, а їхня молитва дійшла до оселі святости Його, до небес!
2CHR|31|1|А коли це все скінчилося, вийшов увесь Ізраїль, що знаходився там, до Юдиних міст, і поламали стовпи для божків, і постинали посвячені дерева, і порозбивали пагірки та жертівники в усьому Юді й Веніямині, і в Єфремі та Манасії аж до кінця. Потому вернулися всі Ізраїлеві сини, кожен до своєї посілости, до своїх міст.
2CHR|31|2|І Єзекія поставив черги священиків та Левитів за їхніми відділами, кожного за його служенням, зо священиків та з Левитів, на цілопалення, і на мирні жертви, на служення й на подяку, і на хвалу в брамах Господніх таборів.
2CHR|31|3|А царева частка зо здобутку його приділена була на цілопалення: на цілопалення ранішні та вечірні, і на цілопалення на суботи й на молодики та на свята, як написано в Законі Господньому.
2CHR|31|4|І наказав він народові, мешканцям Єрусалиму, давати частку священичу та левитську, щоб вони були ревними з Законі Господньому.
2CHR|31|5|А як поширився той наказ, поназносили Ізраїлеві сини багато первоплодів збіжжя, виноградного соку, і нової оливи, і меду, і всякого полевого врожаю; і як десятину того всього багато поназносили.
2CHR|31|6|А Ізраїлеві та Юдині сини, що сиділи по Юдиних містах, також вони поприносили десятину худоби великої та худоби дрібної, і десятину святих речей, посвячених Господеві, їхньому Богові, і понадавали того багато куп.
2CHR|31|7|Третього місяця зачали складати ті купи, а місяця сьомого закінчили.
2CHR|31|8|І прийшли Єзекія та зверхники, і побачили ті купи, і поблагословили Господа та народ Його, Ізраїля.
2CHR|31|9|І вивідував Єзекія священиків та Левитів про ті купи.
2CHR|31|10|І говорив до нього священик Азарія, голова Садокового дому, і сказав: Відколи зачали приносити приношення до Господнього дому, ми їли й були ситі, і багато позосталося, бо Господь поблагословив народ Свій. А з останків складено оцю многоту.
2CHR|31|11|Тоді Єзекія наказав приготовити комори в Господньому домі, і приготовили.
2CHR|31|12|І вірно перенесли туди приношення, і десятину, і святощі, а над ними володарем був Левит Конанія, а брат його Шім'ї другим.
2CHR|31|13|А Єхіїл, і Азазія, і Нахат, і Асагел, і Єрімот, і Йозавад, і Еліїл, і Їсмахія, і Махат, і Беная були урядовцями під рукою Конанії та брата його Шім'ї, призначені царем та Азарієм, володарем при Божому домі.
2CHR|31|14|А Коре, син Їмни, Левит, придверний зо східнього боку, був над добровільними жертвами Богові, щоб видавати Господні приношення та речі найсвятіші.
2CHR|31|15|А при ньому були: Еден, і Мін'ямін, і Єшуа, і Шемая, Амарія, і Шеханія по священичих містах, щоб вірно роздавати їхнім братам за чергами, як великому, так і малому,
2CHR|31|16|окрім їхніх позаписуваних: для мужчин від віку трьох літ і вище, для кожного, хто приходив до Господнього дому на щоденне діло, на їхнє служення, за їхніми сторожами та за їхніми чергами,
2CHR|31|17|і приписаним священикам до дому їхніх батьків, та Левитам від віку двадцяти літ і вище, у сторожах їхніх та в чергах їхніх,
2CHR|31|18|і їхнім приписаним з усіма їхніми дітьми, їхніми жінками, і їхніми синами, і їхніми дочками, для всього збору, бо вони в вірності своїй посвящаються на святість.
2CHR|31|19|А синам священика Аарона, на полях пасовиська їхніх міст, у кожному місті поставлені були мужі, що зазначені поіменно, щоб давати частки кожному мужчині серед священиків та всякому приписаному серед Левитів.
2CHR|31|20|І зробив Єзекія так, як це, по всій Юдеї. І робив він добре й угодне та справедливе перед лицем Господа, Бога свого.
2CHR|31|21|І в усякому ділі, яке він зачинав, у роботі Божого дому, і в Законі, і в заповіді, щоб звертатися до Бога свого, робив він усім своїм серцем, і мав успіх.
2CHR|32|1|По цих справах та по цій вірності прийшов Санхерів, цар асирійський, і ввійшов в Юдею, і розклався табором проти укріплених міст, і думав здобути їх собі.
2CHR|32|2|І побачив Єзекія, що прийшов Санхерів, і що він задумує війну на Єрусалим,
2CHR|32|3|то він нарадився зо своїми зверхниками та своїми лицарями позатикати джерельні води, що назовні міста. І вони допомогли йому.
2CHR|32|4|І було зібрано багато народу, і вони позатикали всі джерела й потік, що плив у Краю, говорячи: Нащо б мали так багато води асирійські царі, коли прийдуть?
2CHR|32|5|І він підбадьорився, і забудував увесь виломаний мур, і поставив на нього башту, а поза тим муром інший мур, і зміцнив Мілло в Давидовому Місті, і наробив багато ратищ та щитів.
2CHR|32|6|І понаставляв він над народом військових зверхників, і зібрав їх до себе, на майдан біля міської брами, і промовляв до їхнього серця, говорячи:
2CHR|32|7|Будьте міцні та будьте мужні, не бійтеся й не жахайтеся перед асирійським царем та перед усім тим натовпом, що з ним, бо з нами більше, ніж із ним.
2CHR|32|8|З ним рамено тілесне, а з нами Господь, Бог наш, щоб допомагати нам та воювати наші війни! І оперся народ на слова Єзекії, Юдиного царя.
2CHR|32|9|По цьому послав Санхерів, асирійський цар, своїх рабів до Єрусалиму, а він сам таборував проти Лахішу, і вся сила його була з ним, до Єзекії, Юдиного царя, і до всього Юди, що в Єрусалимі, сказати:
2CHR|32|10|Так говорить Санхерів, цар асирійський: На що ви сподіваєтесь і сидите в облозі в Єрусалимі?
2CHR|32|11|Оце Єзекія намовляє вас, щоб дати вас на смерть від голоду та від спраги, кажучи: Господь, Бог наш, урятує нас від руки асирійського царя.
2CHR|32|12|Чи ж не він, Єзекія, поруйнував пагірки його та жертівники його, і сказав до Юди та до Єрусалиму, говорячи: Перед одним жертівником будете вклонятися й на ньому будете кадити?
2CHR|32|13|Чи ж ви не знаєте, що зробив я та батьки мої всім народом земель? Чи справді могли боги народів тих країв урятувати свій край від моєї руки?
2CHR|32|14|Хто з-поміж усіх богів цих народів, яких мої батьки вчинили закляттям, міг урятувати свій народ від моєї руки? Як зможе Бог ваш урятувати вас від моєї руки?
2CHR|32|15|А тепер нехай не обманює вас Єзекія, і нехай не зводить вас, як оце. І не вірте йому, бо не зміг жоден бог жодного народу та царства врятувати свого народу від моєї руки та від руки батьків моїх, то тим більше ваші боги не врятують вас від моєї руки!
2CHR|32|16|І ще говорили його раби на Господа, Бога, та на Його раба Єзекію.
2CHR|32|17|І писав він листи з лайкою на Господа, Ізраїлевого Бога, і говорив на Нього таке: Як боги народів тих країв не спасли свого народу від моєї руки, так не спасе Єзекіїн Бог народу Свого від моєї руки!
2CHR|32|18|І кликали вони сильним голосом по-юдейському до єрусалимського народу, що був на мурі, щоб настрашити їх та налякати їх, щоб здобути місто.
2CHR|32|19|І говорили вони на Бога єрусалимського, як на богів землі, чин людських рук.
2CHR|32|20|І молився цар Єзекія та пророк Ісая, син Амосів, про це, і кликали до неба.
2CHR|32|21|І послав Господь Ангола, і він вигубив кожного хороброго вояка, і володаря, і зверхника в таборі царя асирійського, і той вернувся з соромом обличчя до краю свого. А коли він прийшов до дому бога свого, то дехто з тих, що вийшли з нутра його, вбили його там мечем...
2CHR|32|22|І спас Господь Єзекію та єрусалимських мешканців від руки Санхеріва, царя асирійського, та від руки всякого, і дав їм мир навколо.
2CHR|32|23|І багато-хто приносили дара для Господа до Єрусалиму та дорогоцінні речі для Єзекії, Юдиного царя. І він по цьому піднісся в очах усіх народів!
2CHR|32|24|Тими днями занедужав Єзекія смертельно. І він молився до Господа, і Він відповів йому, і дав йому знака.
2CHR|32|25|Та Єзекія не віддав так, як було зроблено йому, бо запишнилося серце його. І був гнів Божий на нього, і на Юдею, та на Єрусалим.
2CHR|32|26|Але впокорився Єзекія в пишноті серця свого, він та мешканці Єрусалиму, і не прийшов на них Господній гнів за днів Єзекії.
2CHR|32|27|І було в Єзекії дуже багато багатства та слави, і він поробив собі скарбниці на срібло й на золото, та на камінь дорогий, і на пахощі, і на щити, і на всякі дорогі речі,
2CHR|32|28|і клуні на врожай збіжжя, і виноградного соку, і свіжої оливи, і жолоби для всякої худоби, і жолоби для черід.
2CHR|32|29|І побудував він собі міста, і мав великий набуток худоби дрібної та худоби великої, бо Бог дав йому дуже великий маєток.
2CHR|32|30|І він, Єзекія, заткнув вихід води горішнього Ґіхону, і вивів її вдолину на захід від Давидового Міста. І мав Єзекія успіх в усіх своїх ділах.
2CHR|32|31|Тільки при послах вавилонських зверхників, посланих до нього, щоб вивідати про чудо, що було в Краю, залишив був його Бог, щоб випробувати його, щоб пізнати все в його серці.
2CHR|32|32|А решта діл Єзекії та його чесноти, ото вони описані в видіннях пророка Ісаї, Амосового сина, у Книзі Царів Юдиних та Ізраїлевих.
2CHR|32|33|І спочив Єзекія з батьками своїми, і поховали його на узбіччях гробів Давидових синів, і віддали йому честь по смерті його, уся Юдея та мешканці Єрусалиму. А замість нього зацарював син його Манасія.
2CHR|33|1|Манасія був віку дванадцяти літ, коли він зацарював, і царював в Єрусалимі п'ятдесят і п'ять літ.
2CHR|33|2|І робив він лихе в Господніх очах, за поганською гидотою тих народів, яких вигнав Господь з-перед Ізраїлевих синів.
2CHR|33|3|І він знову побудував пагірки, які порозбивав був його батько Єзекія, і понаставляв жертівники для Ваалів, і поробив Астарти, і вклонявся всім небесним силам, і служив їм.
2CHR|33|4|І побудував він жертівники в Господньому домі, про якого сказав був Господь: В Єрусалимі буде Ім'я Моє навіки!
2CHR|33|5|І побудував він жертівники для всіх небесних сил на обох подвір'ях Господнього дому.
2CHR|33|6|І він перепроваджував своїх синів через огонь у долині Гінномового сина, і гадав, і ворожив, і чарував, і настановляв викликувачів духів померлих і духів віщих, і багато робив зла в очах Господа, щоб гнівити Його.
2CHR|33|7|І поставив він різаного боввана, якого зробив, у Божому домі, про якого Бог сказав був до Давида та до сина його Соломона: У цьому домі та в Єрусалимі, що його Я вибрав зо всіх міст Ізраїлевих племен, покладу Я Ім'я Своє навіки!
2CHR|33|8|І більше не виступить Ізраїлева нога з тієї землі, яку Я дав вашим батькам, якщо тільки вони будуть пильнувати робити все так, як наказав Я їм, увесь Закон, і устави, і постанови, дані через Мойсея.
2CHR|33|9|Та Манасія робив блудливими Юдею та мешканців Єрусалиму, щоб робити гірше від тих народів, яких Господь вигубив з-перед Ізраїлевих синів.
2CHR|33|10|І говорив Господь до Манасії та до народу його, та не слухались вони.
2CHR|33|11|І Господь навів на них зверхників війська асирійського царя, а вони схопили Манасію на повід, і скували його мідяними кайданами та й повели його до Вавилону.
2CHR|33|12|А як був він утискуваний, благав він лице Господа, Бога свого, і дуже впокорився перед лицем Бога своїх батьків.
2CHR|33|13|І молився він до Нього, і Він був ублаганий, і вислухав благання його, і вернув його до Єрусалиму, до царства його. І пізнав Манасія, що Господь Він Бог!
2CHR|33|14|По цьому збудував він зовнішній мур для Давидового Міста на захід від Ґіхону, в долині, до входу в Рибну браму, й оточив Офела й дуже високо підняв його. І понаставляв він військових зверхників по всіх укріплених містах Юдеї.
2CHR|33|15|І повикидав він чужих богів та подобу боввана з Господнього дому, і всі жертівники, що він побудував був на горі Господнього дому та в Єрусалимі, і викинув те поза місто.
2CHR|33|16|І збудував він Господнього жертівника, і приніс на ньому жертви приносів мирних та вдячних, і звелів юдеям служити Господеві, Богові Ізраїлевому.
2CHR|33|17|Але народ приносив жертви ще на пагірках, тільки вже Господеві, Богові своєму.
2CHR|33|18|А решта діл Манасії, і його молитва до Бога його, і слова прозорливців, що говорили до нього Ім'ям Господа, Бога Ізраїлевого, ото вони описані в історії Ізраїлевих царів.
2CHR|33|19|А молитва його, і як Він був ублаганий, і ввесь його гріх та його спроневірення, і місця, що побудував на них пагірки й поставив Астарти та боввани перед своїм упокоренням, ось вони описані в словах його прозорливців.
2CHR|33|20|І спочив Манасія з батьками своїми, і поховали його в домі його, а замість нього зацарював син його Амон.
2CHR|33|21|Амон був віку двадцяти й двох років, коли він зацарював, і царював він в Єрусалимі два роки.
2CHR|33|22|І робив він зло Господніх очах, як робив його батько Манасія. А всім бовванам, яких наробив його батько Манасія, Амон приносив жертви та служив їм.
2CHR|33|23|І не впокорився він перед Господнім лицем, як упокорився був його батько Манасія, і він, Амон, побільшив провину.
2CHR|33|24|І змовилися раби його на нього, і забили його в його домі.
2CHR|33|25|Та народ Краю перебив усіх змовників на царя Амона. І настановив народ Краю царем замість нього сина його Йосію.
2CHR|34|1|Йосія був віку восьми літ, коли він зацарював, і царював в Єрусалимі тридцять і один рік.
2CHR|34|2|І робив він угодне в Господніх очах, і ходив дорогами свого батька Давида, і не вступався ані праворуч, ані ліворуч.
2CHR|34|3|І восьмого року царювання свого, бувши ще юнаком, розпочав він звертатися до Бога батька свого Давида, а дванадцятого року розпочав очищати Юду та Єрусалим від пагірків, і Астарт, і бовванів різаних та литих.
2CHR|34|4|І порозбивали перед ним Ваалові жертівники, а стовпи сонця, що були на них, він повирубував, а Астарти, і боввани різані та литі поламав і розтер, і розкидав на гроби тих, хто приносив їм жертви.
2CHR|34|5|А кості жерців попалив на їхніх жертівниках, і очистив Юдею та Єрусалим.
2CHR|34|6|А по містах Манасії, і Єфрема, і Симеона, і аж до Нефталима по їхніх руїнах навколо
2CHR|34|7|порозбивав жертівники та Астарти, і потовк боввани на порох, а всі ідоли сонця повирубував в усьому Ізраїлевому краї, і вернувся до Єрусалиму.
2CHR|34|8|А вісімнадцятого року царювання його, по очищенні Краю та Божого дому, послав він Шафана, сина Ацалії, і Маасею, зверхника міста, та Йоаха, та канцлера Йоаха, сина Йохазового, щоб направити дім Господа, Бога його.
2CHR|34|9|І прийшли вони до первосвященика Хілкійї, і дали срібло, що було знесене до Господнього дому, яке зібрали Левити, що стерегли порога, з руки Манасії й Єфрема, та з усієї решти Ізраїля, і з усього Юди й Веніямина та мешканців Єрусалиму.
2CHR|34|10|І дали на руку робітників праці, приставлених до Господнього дому, а робітники тієї праці, що робили в Господньому домі, віддали на відбудову та на направу Божого дому.
2CHR|34|11|І дали вони теслям, і будівничим, щоб купувати тесане каміння та дерева на зв'язування та на покриття домів, що їх понищили Юдині царі.
2CHR|34|12|А ті люди чесно виконували працю, а над ними були поставлені Яхат та Овадія, Левити з синів Мерарієвих, і Захарій та Мешуллам із синів Кегатівців для керування. А всі ті Левіти, що розумілися на музичних знаряддях,
2CHR|34|13|були над носіями, і керували всіма робітниками на кожну роботу; а з Левитів були писарі й урядники та придверні.
2CHR|34|14|А коли вони виймали срібло, принесене до Господнього дому, священик Хілкійя знайшов книгу Господнього Закону, даного через Мойсея.
2CHR|34|15|І відповів Хілкійя й сказав до писаря Шафана: Я знайшов у Господньому домі книгу Закону! І дав Хілкійя ту книгу Шафанові.
2CHR|34|16|І приніс Шафан ту книгу до царя, і приніс цареві ще відповідь, говорячи: Усе, що дано через твоїх рабів, вони роблять.
2CHR|34|17|І вони висипали те срібло, що знайдене в Господньому домі, і дали його на руку приставлених та на руку робітників праці.
2CHR|34|18|І доніс писар Шафан цареві, говорячи: Священик Хілкійя дав мені книгу. І Шафан перечитав з неї перед царем.
2CHR|34|19|І сталося, як цар почув слова книги Закону, то роздер свої шати...
2CHR|34|20|І наказав цар Хілкійї, і Ахікамові, Шафановому синові, і Авдонові, Міхиному синові, і писареві Шафанові, і Асаї, царевому рабові, говорячи:
2CHR|34|21|Ідіть, зверніться до Господа про мене та про позосталих в Ізраїлі та в Юдеї, про слова цієї книги, що знайдена. Великий бо гнів Господній, що вилився на нас за те, що батьки наші це дотримували Господнього слова, щоб робити все, як написано в цій книзі.
2CHR|34|22|І пішов Хілкійя та ті, кому звелів цар, до пророчиці Хулди, жінки Шаллума, сина Токегата, сина Хасриного, сторожа шат, а вона сиділа в Єрусалимі на Новому Місті, і говорили до неї про це.
2CHR|34|23|А вона сказала до них: Так говорить Господь, Бог Ізраїлів: Скажіть чоловікові, що послав вас до мене:
2CHR|34|24|Так говорить Господь: Ось Я наведу лихо на оце місце та на мешканців його, усі ті прокляття, що написані в книзі, яку читали перед Юдиним царем,
2CHR|34|25|за те, що вони покинули Мене й кадили іншим богам, щоб гнівити Мене всіма ділами своїх рук. І вилився гнів Мій на це місце, і він не погасне...
2CHR|34|26|А Юдиному цареві, що послав вас звернутися до Господа, скажете йому так: Так говорить Господь, Бог Ізраїлів, про ті слова, які ти чув:
2CHR|34|27|За те, що зм'якло твоє серце, і ти впокорився перед лицем Бога свого, коли ти почув слова Його на це місце та на мешканців його, і ти впокорився перед лицем Моїм, і роздер свої шати та плакав перед Моїм лицем, то Я також почув, говорить Господь.
2CHR|34|28|Ось Я прилучу тебе до батьків твоїх, і ти будеш прилучений до гробів своїх у спокої, і очі твої не побачать усього того лиха, що Я наведу на оце місце та на мешканців його! І вони принесли відповідь цареві.
2CHR|34|29|А цар послав, і зібрав усіх старших Юдеї та Єрусалиму.
2CHR|34|30|І ввійшов до Господнього дому цар, і кожен муж Юдеї, і мешканці Єрусалиму, і священики, і Левити, і ввесь народ від великого й аж до малого, і він прочитав уголос слова книги Заповіту, знайденої в Господньому домі.
2CHR|34|31|І став цар на своєму місці, і склав заповіта перед Господнім лицем, щоб ходити за Господом та додержувати заповіді Його, і свідчення Його, і устави Його всім серцем своїм та всім життям своїм, щоб виконувати слова того заповіту, що написані в тій книзі.
2CHR|34|32|І наставив він кожного, хто знаходився в Єрусалимі та в Веніямині, до того. І мешканці Єрусалиму робили за заповітом Бога, Бога своїх батьків.
2CHR|34|33|І Йосія повикидав усі поганські гидоти з усіх країв, що в Ізраїлевих синів, і змусив кожного, хто знаходився в Ізраїлі, служити Господеві, їхньому Богові. За всіх днів його вони не відступали від Господа, Бога своїх батьків.
2CHR|35|1|І справив Йосія в Єрусалимі Пасху для Господа, і зарізали пасхальне ягня чотирнадцятого дня першого місяця.
2CHR|35|2|І поставив він священиків на їхні становища, і підбадьорував їх на службу Господнього дому.
2CHR|35|3|І сказав він Левитам, наставникам усього Ізраїля, посвяченим для Господа: Дайте святого ковчега до храму, що його збудував Соломон, син Давидів, цар Ізраїлів. Нема пощо вам носити його на раменах, служіть тепер Господеві, вашому Богові, та Його народові, Ізраїлеві.
2CHR|35|4|І приготуйтеся за родом ваших батьків, за вашими чергами, за писанням Давида, Ізраїлевого царя, та за писанням його сина Соломона.
2CHR|35|5|І станьте в святині за відділами батьківських родів ваших братів, синів народу, а поділ за батьківськими домами в Левитів.
2CHR|35|6|І заріжте пасхальне ягня, й освятіться, і приготуйте для ваших братів, щоб робити за Господнім словом, даним через Мойсея.
2CHR|35|7|І дав Йосія для людських синів худоби дрібної, овечок та молодих кіз, це все на пасхальне ягня для кожного, хто знаходився в Єрусалимі, числом тридцять тисяч, а худоби великої три тисячі. Це з набутку царевого.
2CHR|35|8|А його зверхники дали на жертву для народу, для священиків та для Левитів: Хілкійя, і Захарій, і Єхіїл, старші в Божому домі, дали священикам на пасхальні жертви дві тисячі й шість сотень худоби дрібної, а худоби великої три тисячі.
2CHR|35|9|А Конанія, і Шемая, і брат його Натанаїл, і Хашавія, і Єіїл, і Йозавад, зверхники Левитів, дали для Левитів на пасхальні жертви п'ять тисяч худоби дрібної, а худоби великої п'ять сотень.
2CHR|35|10|І була міцно встановлена служба, і стали священики на своїм становищі, а Левити при своїх чергах, за наказом царя.
2CHR|35|11|І різали пасхальне ягня, а священики кропили кров'ю, беручи з їхньої руки, а Левити здирали шкуру.
2CHR|35|12|І відділили, що було на цілопалення, щоб дати їх за відділами, по батьківських домах синам народу на приношення Господеві, як написано в Мойсеєвій книзі. І так зробили й з худобою великою.
2CHR|35|13|І пекли пасхальне ягня на огні, за постановою, а святі жертви варили в горшках, і в котлах, і в горнятах, і швидко несли всім синам народу.
2CHR|35|14|А потім наварили собі та священикам, бо священики, Ааронові сини, були зайняті приношенням цілопалення та лою аж до ночі, то Левити наготовили їжі собі та священикам, Аароновим синам.
2CHR|35|15|А співаки, Асафові сини, були на своїх місцях за наказом Давида, і Асафа, і Гемана, і Єдутуна, царевого прозорливця, а придверні були при кожній брамі, їм не треба було відходити від своїх робіт, бо їхні брати Левити наготовили їм.
2CHR|35|16|І була міцно встановлена вся Господня служба того дня, щоб справити Пасху й принести цілопалення на Господньому жертівнику, за наказом царя Йосії.
2CHR|35|17|І Ізраїлеві сини, що знаходилися там, справляли того часу Пасху та свято Опрісноків сім день.
2CHR|35|18|І не справлялася Пасха, як ця, в Ізраїлі від днів пророка Самуїла, а всі Ізраїлеві царі не справляли такої, як ця Пасха, що справив Йосія, і священики, і Левити, і ввесь Юда та Ізраїль, що знаходився там, та мешканці Єрусалиму.
2CHR|35|19|Вісімнадцятого року царювання Йосії справлялася ця Пасха.
2CHR|35|20|По всьому цьому, коли Йосія приготовив дім Божий, прийшов Нехо, цар єгипетський, щоб воювати в Каркеміші над Ефратом, а Йосія вийшов навпроти нього.
2CHR|35|21|І послав той до нього послів, говорячи: Що мені до тебе, царю Юдин? Не проти тебе приходжу я сьогодні, але проти дому, що воює зо мною. А Бог наказав мені спішити. Не протився Богові, що зо мною, і нехай Він не знищить тебе!
2CHR|35|22|Та Йосія не відвернувся від нього, але перебрався, щоб воювати з ним, і не послухався слів Нехо, що були з Божого наказу, і прийшов воювати в долині Меґіддо.
2CHR|35|23|І вистрілили стрільці на царя Йосію. І сказав цар до своїх рабів: Відведіть мене, бо я сильно ранений...
2CHR|35|24|І перевели його його раби з військової колесниці на його другий повіз, і відвезли його до Єрусалиму. І помер він, і був похований у гробах своїх батьків, а вся Юдея та Єрусалим були в жалобі по Йосії.
2CHR|35|25|І Єремія співав жалобну пісню по Йосії. А всі співаки та співачки оповідали в жалобних своїх піснях про Йосію, і так є аж до сьогодні, і дали їх за уставу для Ізраїля, і ось вони написані в Жалобних Піснях.
2CHR|35|26|А решта діл Йосії та його чесноти, за написаним у Господнім Законі,
2CHR|35|27|і дії його перші та останні, ото вони описані в Книзі Царів Ізраїлевих та Юдиних.
2CHR|36|1|А народ Краю взяв Йоахаза, сина Йосії, і настановив його царем в Єрусалимі замість батька його.
2CHR|36|2|Йоахаз був віку двадцяти й трьох літ, коли він зацарював, і царював в Єрусалимі три місяці.
2CHR|36|3|І скинув його єгипетський цар в Єрусалимі, і наклав кару на цей Край, сто талантів срібла та талант золота.
2CHR|36|4|І єгипетський цар настановив царем над Юдеєю та Єрусалимом брата його Ел'якима, і змінив ім'я йому на Єгояким. А брата його Йоахаза узяв Нехо й відвів його до Єгипту.
2CHR|36|5|Єгояким був віку двадцяти й п'яти літ, коли він зацарював, і одинадцять років царював в Єрусалимі. І робив він зло в очах Господа, Бога свого.
2CHR|36|6|На нього пішов Навуходоносор, цар вавилонський, і він закував його в мідяні кайдани, щоб відвести його до Вавилону.
2CHR|36|7|А дещо з посуду Господнього дому Навуходоносор відправив до Вавилону, і дав його до храму свого в Вавилоні.
2CHR|36|8|А решта Єгоякимових діл та гидоти його, які він робив, і що знайдено проти нього, ото вони описані в Книзі Царів Ізраїлевих та Юдиних. А замість нього зацарював син його Єгояхін.
2CHR|36|9|Єгояхін був віку восьми літ, коли він зацарював, і царював в Єрусалимі три місяці й десять день. І робив він лихе в Господніх очах.
2CHR|36|10|А по році послав цар Навуходоносор, і привів його до Вавилону з дорогим посудом Господнього дому, а царем над Юдеєю та Єрусалимом настановив брата його Седекію.
2CHR|36|11|Седекія був віку двадцяти й одного року, коли він зацарював, і він царював в Єрусалимі одинадцять років.
2CHR|36|12|І робив він зло в очах Господа, Бога свого, не впокорився перед пророком Єремією, що говорив із наказу Господнього.
2CHR|36|13|І він також відкинувся від царя Навуходоносора, що був заприсягнув його Господом, і вчинив твердою свою шию, і став запеклим, щоб не навертатися до Господа, Бога Ізраїлевого.
2CHR|36|14|Також усі зверхники священиків та народу ще більше грішили, шануючи гидоти поган, і вони занечистили Господній дім, якого Він освятив в Єрусалимі.
2CHR|36|15|А Господь, Бог їхніх батьків, усе посилав до них через Своїх послів слова остороги, бо Він змилосердився над народом Своїм та над оселею Своєю.
2CHR|36|16|Та вони соромили Божих послів, і погорджували їхніми словами, і насміхалися з Його пророків, аж поки не піднісся гнів Господа на народ Його так, що не було вже ліку.
2CHR|36|17|І Він навів на них халдейського царя, і той позабивав мечем їхніх вибраних у домі їхньої святині, і не змилосердився ані над юнаком, ані над дівчиною, ані над старим, ані над старезним, усе дав в його руку...
2CHR|36|18|І всі речі Божого дому, великі та малі, і скарби дому Господнього та дому царя й його зверхників, усе переніс до Вавилону.
2CHR|36|19|І спалили вони Божий дім, і порозбивали мур Єрусалиму, і всі палати його попалили огнем, а всі дорогі речі його понищили...
2CHR|36|20|І пішло на вигнання до Вавилону позостале від меча, і стали йому та синам його за рабів аж до зацарювання перського царства,
2CHR|36|21|щоб виповнилося Господнє слово, проречене Єреміїними устами, аж поки вподобає собі земля свої суботи, по всі дні її спустошення святкувала вона суботи, щоб сповнилися сімдесят літ.
2CHR|36|22|А першого року Кіра, царя перського, коли сповнилось слово Господнє, проречене устами Єреміїними, збудив Господь духа Кіра, царя перського, і він оголосив по всьому царству своєму, а також на письмі, говорячи:
2CHR|36|23|Так говорить Кір, цар перський: Усі земні царства дав мені Господь, Бог Небесний, і Він наклав на мене збудувати Йому храма в Єрусалимі, що в Юдеї. Хто між вами з усього Його народу, нехай буде Господь, Бог його, з ним, і нехай він іде до Єрусалиму!
