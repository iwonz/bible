REV|1|1|耶稣基督的启示，就是上帝赐给他，要他将必须快要发生的事指示他的众仆人。他差遣使者指明给他的仆人 约翰 ，
REV|1|2|约翰 就将上帝的道和耶稣基督的见证，凡自己所看见的，都见证出来。
REV|1|3|诵读这书上预言的，和那些听见又遵守其中所记载的，都是有福的，因为时候近了。
REV|1|4|约翰 写信给 亚细亚 的七个教会。愿那位今在、昔在、以后永在的上帝，与他宝座前的七灵，和那忠信的见证者、从死人中复活的首生者 、世上君王的元首耶稣基督，赐恩惠和平安 给你们。 他爱我们，用自己的血使我们从罪中得释放 ，
REV|1|5|
REV|1|6|又使我们成为国度，作他父上帝的祭司。愿荣耀、权能归给他，直到永永远远 。阿们！
REV|1|7|“看哪，他驾云降临； 众目都要看见他， 连刺他的人也要看见他； 地上的万族要因他哀哭。” 这是真实的。阿们！
REV|1|8|主上帝说：“我是阿拉法，我是俄梅戛 ，是今在、昔在、以后永在的全能者。”
REV|1|9|我— 约翰 就是你们的弟兄，在耶稣里和你们一同在患难、国度、忍耐里有份的，为上帝的道，并为给耶稣作的见证，曾在那名叫 拔摩 的海岛上。
REV|1|10|有一主日我被圣灵感动，听见在我后面有大声音如吹号，
REV|1|11|说：“把你所看见的写在书上，寄给 以弗所 、 士每拿 、 别迦摩 、 推雅推喇 、 撒狄 、 非拉铁非 、 老底嘉 那七个教会。”
REV|1|12|我转过身来要看看是谁的声音在跟我说话。我一转过来，看见了七个金灯台；
REV|1|13|在灯台中间有一位好像人子的，身穿垂到脚的长袍，胸间束着金带。
REV|1|14|他的头与发皆白，如白羊毛，如雪；他的眼睛好像火焰，
REV|1|15|双脚好像在炉中锻鍊得发亮的铜，声音好像众水的声音。
REV|1|16|他右手拿着七颗星，从他口中吐出一把两刃的利剑，面貌好像烈日放光。
REV|1|17|我看见了他，就仆倒在他脚前，像死人一样。他用右手按着我说：“不要怕。我是首先的，是末后的，
REV|1|18|又是永活的。我曾死过，看哪，我是活着的，直到永永远远；并且我拿着死亡和阴间的钥匙。
REV|1|19|所以，你要把所看见的事、现在的事和以后将发生的事，都写下来。
REV|1|20|至于你所看见、在我右手中的七颗星和那七个金灯台的奥秘就是：七颗星是七个教会的使者，七个灯台是七个教会。”
REV|2|1|“你要写信给 以弗所 教会的使者，说：‘那右手拿着七颗星，在七个金灯台中间行走的这样说：
REV|2|2|我知道你的行为、劳碌、忍耐，也知道你不容忍恶人。你也曾察验那自称为使徒却不是使徒的，看出他们是假的。
REV|2|3|你能忍耐，曾为我的名劳苦而不困倦。
REV|2|4|然而，有一件事我要责备你，就是你把起初的爱心抛弃了。
REV|2|5|所以你要回想你是从哪里坠落的，并且要悔改，做起初所做的工作。你若不悔改，我要到你那里去，把你的灯台从原处挪去。
REV|2|6|然而你还有一件可取的事，就是你恨恶 尼哥拉 派的行为，这种行为也是我所恨恶的。
REV|2|7|凡有耳朵的都应当听圣灵向众教会所说的话。得胜的，我必将上帝乐园中生命树的果子赐给他吃。’”
REV|2|8|“你要写信给 士每拿 教会的使者，说：‘那首先的、末后的，死过又活了的这样说：
REV|2|9|我知道你的患难和贫穷—其实你却是富足的，也知道那自称是 犹太 人的所说毁谤的话，其实他们不是 犹太 人，而是撒但会堂的人。
REV|2|10|你将要受的苦，你不用怕。看哪！魔鬼要把你们中间几个人下在监里，使你们受考验，你们要遭受苦难十日。你务要至死忠心，我就赐给你那生命的冠冕。
REV|2|11|凡有耳朵的都应当听圣灵向众教会所说的话。得胜的必不受第二次死的害。’”
REV|2|12|“你要写信给 别迦摩 教会的使者，说：‘那有两刃利剑的这样说：
REV|2|13|我知道你的居所，就是有撒但座位之处；当我忠心的见证人 安提帕 在你们中间，在撒但所住的地方被杀之时，你还坚守我的名，没有否认对我的信仰。
REV|2|14|然而，有几件事我要责备你，就是在你那里有人服从了 巴兰 的教训；这 巴兰 曾教唆 巴勒 将绊脚石放在 以色列 人面前，使他们吃祭过偶像之物，并且犯淫乱。
REV|2|15|同样，你那里也有人服从了 尼哥拉 派的教训。
REV|2|16|所以，你当悔改；若不悔改，我很快就到你那里来，用我口中的剑攻击他们。
REV|2|17|凡有耳朵的都应当听圣灵向众教会所说的话。得胜的，我必将那隐藏的吗哪赐给他，并赐他一块白石，石上写着新的名字，除了那领受的以外，没有人认识。’”
REV|2|18|“你要写信给 推雅推喇 教会的使者，说：‘上帝的儿子，那位眼睛如火焰、双脚像发亮的铜的这样说：
REV|2|19|我知道你的行为：爱心、信心、勤劳、忍耐；又知道你末后所行的善事比起初所行的更多。
REV|2|20|然而，有一件事我要责备你，就是你容忍那自称是先知的妇人 耶洗别 教唆我的仆人，引诱他们犯淫乱，吃祭过偶像之物。
REV|2|21|我曾给她悔改的机会，她却不肯悔改她的淫行。
REV|2|22|看吧，我要使她病倒在床上。那些与她犯奸淫的人若不悔改他们的行为，我也要使他们同受大患难。
REV|2|23|我又要杀死她的儿女，众教会就知道，我是那察看人肺腑心肠的，我要照你们的行为报应各人。
REV|2|24|至于你们其余的 推雅推喇 人，就是一切不随从这教训，不明白他们所谓撒但深奥之理的人，我告诉你们，我不会再把别的担子放在你们身上。
REV|2|25|你们只要持守那已经有的，直到我来。
REV|2|26|那得胜又遵守我命令到底的， 我要赐给他权柄制伏列国；
REV|2|27|他必用铁杖管辖他们， 如同打碎陶器，
REV|2|28|像我也从我父领受了权柄一样。我又要把晨星赐给他。
REV|2|29|凡有耳朵的都应当听圣灵向众教会所说的话。’”
REV|3|1|“你要写信给 撒狄 教会的使者，说：‘那有上帝的七灵和七颗星的这样说：我知道你的行为，就是名义上你是活的，实际上你是死的。
REV|3|2|你要警醒，坚固那些剩下、快要死的，因为我发现你的行为，在我上帝面前没有一样是完全的。
REV|3|3|所以，要记得你所领受和听见的；要遵守，并要悔改。你若不警醒，我必如贼一样来到；我几时来到你那里，你绝不会知道。
REV|3|4|然而，在 撒狄 你还有几位是未曾污秽自己衣服的，他们会穿白衣与我同行，因为他们是配穿的。
REV|3|5|得胜的必这样穿白衣，我也不从生命册上涂去他的名；我要在我父面前，和我父的众使者面前，宣认他的名。
REV|3|6|凡有耳朵的都应当听圣灵向众教会所说的话。’”
REV|3|7|“你要写信给 非拉铁非 教会的使者，说： ‘那神圣、真实的， 拿着 大卫 的钥匙， 开了就没有人能关， 关了就没有人能开的这样说：
REV|3|8|我知道你的行为。看哪，我在你面前给你一个敞开的门，是没有人能关的。我知道你有一点力量，也遵守我的道，没有否认我的名。
REV|3|9|那属撒但会堂的，自称是 犹太 人，其实不是 犹太 人，而是说谎话的，我要使他们来到你脚前下拜，使他们知道我已经爱你了。
REV|3|10|因为你遵守了我坚忍的道，我也必在普天下人受试炼的时候保守你免受试炼。
REV|3|11|我必快来，你要持守你所有的，免得人夺去你的冠冕。
REV|3|12|得胜的，我要使他在我上帝的殿中作柱子，他必不再从那里出去。我又要把我上帝的名和我上帝城的名—从天上我上帝那里降下来的新 耶路撒冷 ，和我的新名，都写在他上面。
REV|3|13|凡有耳朵的都应当听圣灵向众教会所说的话。’”
REV|3|14|“你要写信给 老底嘉 教会的使者，说：‘那位阿们、诚信真实的见证者、上帝创造的根源这样说：
REV|3|15|我知道你的行为，你也不冷也不热；我巴不得你或冷或热。
REV|3|16|既然你如温水，也不冷也不热，我要从我口中把你吐出去。
REV|3|17|你说：我是富足的，已经发了财，一样都不缺，却不知道你是困苦、可怜、贫穷、瞎眼、赤身的。
REV|3|18|我劝你向我买从火中锻鍊出来的金子，使你富足；又买白衣穿上，使你赤身的羞耻不露出来；又买眼药抹你的眼睛，使你能看见。
REV|3|19|凡我所疼爱的，我就责备管教。所以，你要发热心，也要悔改。
REV|3|20|看哪，我站在门外叩门，若有听见我声音而开门的，我要进到他那里去，我与他，他与我一起吃饭。
REV|3|21|得胜的，我要赐他在我宝座上与我同坐，就如我得了胜，在我父的宝座上与他同坐一般。
REV|3|22|凡有耳朵的都应当听圣灵向众教会所说的话。’”
REV|4|1|这些事以后，我观看，看见天上有一道门开着。我头一次听见的那好像吹号的声音对我说：“你上这里来，我要把此后必须发生的事指示你。”
REV|4|2|我立刻被圣灵感动，见有一个宝座安置在天上，有一位坐在宝座上。
REV|4|3|那坐着的，看来好像碧玉和红宝石；又有彩虹围着宝座，光彩好像绿宝石。
REV|4|4|宝座的周围又有二十四个座位，上面坐着二十四位长老，身穿白衣，头上戴着金冠冕。
REV|4|5|有闪电、声音、雷轰从宝座中发出。在宝座前点着七支火炬，就是上帝的七灵。
REV|4|6|宝座前有一个如同水晶的玻璃海。 宝座的周围，四边有四个活物，遍体前后都长满了眼睛。
REV|4|7|第一个活物像狮子，第二个像牛犊，第三个的脸像人脸，第四个像飞鹰。
REV|4|8|四个活物各有六个翅膀，遍体内外都长满了眼睛。他们昼夜不住地说： “圣哉！圣哉！圣哉！ 主—全能的上帝； 昔在、今在、以后永在！”
REV|4|9|每逢四活物将荣耀、尊贵、感谢归给那坐在宝座上、活到永永远远者的时候，
REV|4|10|二十四位长老就俯伏敬拜坐在宝座上活到永永远远的那一位，又把他们的冠冕放在宝座前，说：
REV|4|11|“我们的主，我们的上帝， 你配得荣耀、尊贵、权柄， 因为你创造了万物， 万物因你的旨意被创造而存在。”
REV|5|1|我看见坐在宝座那位的右手中有书卷，正反面都写着字，用七个印密封着。
REV|5|2|我又看见一位大力的天使大声宣告说：“有谁配展开那书卷，揭开那七个印呢？”
REV|5|3|在天上、地上、地底下，没有人能展开、能阅览那书卷。
REV|5|4|因为没有人配展开、阅览那书卷，我就大哭。
REV|5|5|长老中有一位对我说：“不要哭。看哪， 犹大 支派中的狮子， 大卫 的根，他已得胜，能展开那书卷，揭开那七个印。”
REV|5|6|我又看见宝座和四个活物，以及长老之中有羔羊站着，像是被杀的，有七个角七只眼睛，就是上帝的七 灵，奉差遣往普天下去的。
REV|5|7|这羔羊前来，从坐在宝座上那位的右手中拿了书卷。
REV|5|8|他一拿了书卷，四活物和二十四位长老就俯伏在羔羊面前，各拿着琴和盛满了香的金炉；这香就是众圣徒的祈祷。
REV|5|9|他们唱新歌，说： “你配拿书卷， 配揭开它的七印； 因为你曾被杀，用自己的血 从各支派、各语言、各民族、各邦国中买了人来，使他们归于上帝，
REV|5|10|又使他们成为国民和祭司，归于我们的上帝； 他们将在地上执掌王权。”
REV|5|11|我又观看，我听见宝座和活物及长老的周围有许多天使的声音；他们的数目有千千万万，
REV|5|12|大声说： “被杀的羔羊配得 权能、丰富、智慧、力量、 尊贵、荣耀、颂赞。
REV|5|13|我又听见在天上、地上、地底下、沧海里和天地间一切所有被造之物，都说： “愿颂赞、尊贵、荣耀、权势， 都归给坐在宝座上的那位和羔羊， 直到永永远远！”
REV|5|14|四活物就说：“阿们！”众长老也俯伏敬拜。
REV|6|1|我看见羔羊揭开七个印中第一个印的时候，听见四活物中的一个活物，声音如雷，说：“你来！”
REV|6|2|我就观看，看见一匹白马，骑在马上的拿着弓，并有冠冕赐给他。他出来征服，胜而又胜。
REV|6|3|羔羊揭开第二个印的时候，我听见第二个活物说：“你来！”
REV|6|4|就另有一匹马出来，是红色的；有权柄赐给了那骑马的，要从地上夺去太平，使人彼此相杀；他又接受了一把大刀。
REV|6|5|羔羊揭开第三个印的时候，我听见第三个活物说：“你来！”我就观看，看见一匹黑马；骑在马上的，手里拿着天平。
REV|6|6|我听见在四个活物中似乎有声音说：“一个银币买一升麦子，一个银币买三升大麦；油和酒不可糟蹋。”
REV|6|7|羔羊揭开第四个印的时候，我听见第四个活物说：“你来！”
REV|6|8|我就观看，看见一匹灰色马；骑在马上的，名字叫作“死”，阴间也随着他；有权柄赐给他们，可以用刀剑、饥荒、瘟疫、野兽，杀害地上四分之一的人。
REV|6|9|羔羊揭开第五个印的时候，我看见在祭坛底下有曾为上帝的道，并为作见证而被杀的人的灵魂，
REV|6|10|大声喊着说：“神圣真实的主宰啊，你不审判住在地上的人，为我们所流的血伸冤，要到几时呢？”
REV|6|11|于是有白袍赐给他们各人；又有话吩咐他们还要歇息片刻，等到与他们同作仆人的，和他们的弟兄，像他们一样被杀的人的数目凑足的时候。
REV|6|12|羔羊揭开第六个印的时候，我看见地大震动，太阳变黑像粗麻布，整个月亮变红像血，
REV|6|13|天上的星辰坠落在地上，如同无花果树被大风摇动，落下未熟的果子一样。
REV|6|14|天就裂开，好像书卷被卷起来；山岭海岛都被移动离开原位。
REV|6|15|地上的君王、臣宰、将军、富户、壮士，和一切为奴的、自主的，都藏在山洞和岩石穴里，
REV|6|16|向山和岩石说：“倒在我们身上吧！把我们藏起来，躲避坐宝座者的脸面和羔羊的愤怒；
REV|6|17|因为他们遭愤怒的大日子到了，谁能站得住呢？”
REV|7|1|此后，我看见四位天使站在地的四角，执掌地上四方的风，使风不吹在地上、海上和各种树上。
REV|7|2|我又看见另有一位天使从日出之地上来，拿着永生上帝的印。他向那得到权柄能伤害地和海的四位天使大声喊着，
REV|7|3|说：“你们不可伤害地、海和树林，等我们在我们上帝众仆人的额上盖了印。”
REV|7|4|我听见 以色列 人各支派中受印的数目有十四万四千；
REV|7|5|犹大 支派中受印的有一万二千； 吕便 支派中有一万二千； 迦得 支派中有一万二千；
REV|7|6|亚设 支派中有一万二千； 拿弗他利 支派中有一万二千； 玛拿西 支派中有一万二千；
REV|7|7|西缅 支派中有一万二千； 利未 支派中有一万二千； 以萨迦 支派中有一万二千；
REV|7|8|西布伦 支派中有一万二千； 约瑟 支派中有一万二千； 便雅悯 支派中受印的有一万二千。
REV|7|9|此后，我观看，看见有许多人，没有人能计算，是从各邦国、各支派、各民族、各语言来的，站在宝座和羔羊面前，身穿白衣，手拿棕树枝，
REV|7|10|大声喊着说： “愿救恩归于坐在宝座上我们的上帝， 也归于羔羊！”
REV|7|11|众天使都站在宝座和众长老，以及四个活物的周围，俯伏在宝座前，敬拜上帝，
REV|7|12|说： “阿们！颂赞、荣耀、智慧、 感谢、尊贵、权能、 力量都归于我们的上帝， 直到永永远远。阿们！”
REV|7|13|长老中有一位回应我说：“这些穿白衣的是谁？是从哪里来的？”
REV|7|14|我对他说：“我主啊，你是知道的。”他向我说：“这些人是从大患难中出来的，他们曾用羔羊的血把衣裳洗得洁白。
REV|7|15|所以，他们在上帝宝座前， 昼夜在他殿中事奉他； 那坐在宝座上的要用帐幕覆庇他们。
REV|7|16|他们不再饥，不再渴； 太阳必不伤害他们， 任何炎热也不伤害他们，
REV|7|17|因为宝座中的羔羊必牧养他们， 领他们到生命水的泉源； 上帝必擦去他们一切的眼泪。”
REV|8|1|羔羊揭开第七个印的时候，天上寂静约有半小时。
REV|8|2|我看见那站在上帝面前的七位天使，有七枝号赐给他们。
REV|8|3|另有一位天使拿着金香炉来，站在祭坛旁边；有许多香赐给他，要和众圣徒的祈祷一同献在宝座前的金坛上。
REV|8|4|那香的烟和众圣徒的祈祷从天使的手中一同升到上帝面前。
REV|8|5|天使拿着香炉，盛满了坛上的火，倒在地上；就有雷轰、响声、闪电、地震。
REV|8|6|拿着七枝号筒的七位天使预备好要吹号。
REV|8|7|第一位天使吹号，就有冰雹和火搀着血扔在地上；地的三分之一和树的三分之一被烧掉了，一切的青草也被烧掉了。
REV|8|8|第二位天使吹号，就有像火烧着的大山扔在海中；海的三分之一变成血，
REV|8|9|海中有生命的被造之物死了三分之一，船只也毁坏了三分之一。
REV|8|10|第三位天使吹号，就有烧着的大星好像火把从天上坠下来，落在江河的三分之一和众水的泉源上。
REV|8|11|这星名叫“苦艾”；众水的三分之一变为苦艾，许多人因水变苦而死了。
REV|8|12|第四位天使吹号，太阳的三分之一、月亮的三分之一、星辰的三分之一都被击打，以致日月星的三分之一变黑了，白昼的三分之一没有光，黑夜也是这样。
REV|8|13|我观看，听见一只在空中飞的鹰大声说：“祸哉！祸哉！祸哉！地上的居民哪，其余的三位天使快要吹号了！”
REV|9|1|第五位天使吹号，我就看见一颗星从天上坠落到地上；有无底坑的钥匙赐给它。
REV|9|2|它开了无底坑，就有烟从坑里往上冒，好像大火炉的烟；太阳和天空都因这烟昏暗了。
REV|9|3|有蝗虫从烟中出来，飞到地上，有权柄赐给它们，好像地上的蝎子有权柄一样。
REV|9|4|它们奉命不可伤害地上的草、各样绿色植物和各种树木，惟独可伤害额上没有上帝印记的人；
REV|9|5|但是不许蝗虫害死他们，只可使他们受痛苦五个月；这痛苦就像人被蝎子螫了的痛苦一样。
REV|9|6|在那些日子，人求死，却死不了；想死，死却避开他们。
REV|9|7|蝗虫的形状好像预备上阵的战马一样，头上戴的好像金冠冕，脸面好像男人的脸面，
REV|9|8|头发像女人的头发，牙齿像狮子的牙齿；
REV|9|9|它们胸前有甲，好像铁甲；又有翅膀的响声，好像许多车马奔跑上阵的声音。
REV|9|10|它们有尾巴像蝎子，长着毒刺，尾巴上的毒刺有能力伤害人五个月。
REV|9|11|它们有无底坑的使者作它们的王，按着 希伯来 话名叫 亚巴顿 ， 希腊 话名话叫 亚玻伦 。
REV|9|12|第一样灾祸过去了；看哪，还有两样灾祸要来。
REV|9|13|第六位天使吹号，我听见有声音从上帝面前金坛的四 角发出来，
REV|9|14|吩咐那吹号的第六位天使，说：“把那捆绑在 幼发拉底 大河的四个使者释放了。”
REV|9|15|那四个使者就被释放；他们原是预备好，在特定的年、月、日、时，要杀人类的三分之一。
REV|9|16|骑兵有二亿；他们的数目我听见了。
REV|9|17|我在异象中看见那些马和骑马的：骑马的穿着火红、紫玛瑙及硫磺色的胸甲；马的头好像狮子的头，有火、有烟、有硫磺从马的口中喷出来。
REV|9|18|从马的口中所喷出来的火、烟和硫磺这三样灾害杀了人类的三分之一。
REV|9|19|马的能力在于它们的口和尾巴；它们的尾巴像蛇，有头，用头来伤害人。
REV|9|20|其余未曾被这些灾难所杀的人仍旧不为自己手所做的悔改，还是去拜鬼魔和那些不能看、不能听、不能走，用金、银、铜、木、石所造的偶像。
REV|9|21|他们也不为自己所犯的那些凶杀、邪术、淫乱、偷窃的事悔改。
REV|10|1|我又看见另一位大力的天使从天降下，披着云彩，头上有彩虹，脸面像太阳，两脚像火柱。
REV|10|2|他手里拿着展开的小书卷。他右脚踏海，左脚踏地，
REV|10|3|大声呼喊，好像狮子吼叫。呼喊完了，就有七个雷发出声音。
REV|10|4|七个雷发声后，我正要写出来，就听见从天上有声音说：“七个雷所说的，你要封上，不可写出来。”
REV|10|5|我所看见的那踏海踏地的天使向天举起右手，
REV|10|6|指着创造天和天上之物、地和地上之物、海和海中之物、直活到永永远远的那位起誓，说：“不再有时日了 。”
REV|10|7|但在第七位天使要吹号的日子，上帝的奥秘就要成全了，正如上帝向他仆人众先知所宣告的。
REV|10|8|我先前从天上所听见的那声音又吩咐我说：“你去，把那踏海踏地之天使手中展开的小书卷拿过来。”
REV|10|9|我就走到天使那里，对他说，请他把小书卷给我。他对我说：“你拿去，把它吃光。它会使你肚子发苦，然而在你口中会甘甜如蜜。”
REV|10|10|于是我从天使手中把小书卷接过来，把它吃光了，在我口中果然甘甜如蜜，吃了以后，我肚子觉得发苦。
REV|10|11|天使们对我说：“你必须指着许多民族、邦国、语言、君王再说预言。”
REV|11|1|有一根芦苇，像丈量的杖，赐给我；且有话说：“起来！将上帝的殿和祭坛，以及在殿中礼拜的人，都量一量。
REV|11|2|只是殿外的院子不用量，因为这是要给外邦人的；他们将践踏圣城四十二个月。
REV|11|3|“我要赐权柄给我那两个见证人，穿着粗麻衣说预言一千二百六十天。”
REV|11|4|他们就是那站在世界之主面前的两棵橄榄树和两个灯台。
REV|11|5|若有人想要害他们，就有火从他们口中喷出来，烧灭仇敌；凡想要害他们的都必须这样被杀。
REV|11|6|这二人有权柄关闭天空，使他们说预言的日子不下雨；又有权柄使水变为血，并且能随时随意用各样的灾害击打大地世界。
REV|11|7|他们作完见证的时候，那从无底坑里上来的兽要跟他们交战，并且得胜，把他们杀了。
REV|11|8|他们的尸首将倒在大城的街道上；这城按着灵意叫 所多玛 ，又叫 埃及 ，就是他们的主钉十字架的地方。
REV|11|9|从各民族、支派、语言、邦国中有人观看他们的尸首三天半，又不许人把尸首安放在坟墓里。
REV|11|10|住在地上的人会因他们而欢喜快乐，互相馈送礼物，因为这两位先知曾使住在地上的人受痛苦。
REV|11|11|过了这三天半，有生命的气息从上帝那里进入他们里面，他们就站起来；看见他们的人都大大惧怕。
REV|11|12|两位先知听见有大声音从天上对他们说：“上这里来。”他们就驾着云上了天，他们的仇敌也看见了。
REV|11|13|正在那时候，地大震动，城倒塌了十分之一；因地震而死的有七千人，其余的都恐惧，归荣耀给天上的上帝。
REV|11|14|第二样灾祸过去了；看哪，第三样灾祸快到了。
REV|11|15|第七位天使吹号，天上就有大声音说： “世上的国已成了我们的主和他所立的基督的国了。 他要作王直到永永远远！”
REV|11|16|在上帝面前，坐在自己座位上的二十四位长老都俯伏在地上敬拜上帝，
REV|11|17|说： “今在昔在的主—全能的上帝啊， 我们感谢你！ 因你执掌大权作王了。
REV|11|18|外邦发怒， 你的愤怒临到了。 审判死人的时候也到了； 你的仆人众先知、众圣徒及敬畏你名的人， 连大带小得赏赐的时候到了； 你毁灭那些毁灭大地者的时候也到了。”
REV|11|19|于是，上帝天上的圣所开了，在他圣所中，他的约柜出现了；随后有闪电、响声、雷轰、地震、大冰雹。
REV|12|1|天上出现了一个大兆头：有一个妇人身披太阳，脚踏月亮，头戴十二颗星的冠冕；
REV|12|2|她怀了孕，在生产的阵痛中疼痛地喊叫。
REV|12|3|天上又出现了另一个兆头：有一条大红龙 ，有七个头十个角；七个头上戴着七个冠冕。
REV|12|4|它的尾巴拖拉着天上星辰的三分之一，把它们摔在地上。然后龙站在那将要生产的妇人面前，等她生产后要吞吃她的孩子。
REV|12|5|妇人生了一个男孩子，就是将来要用铁杖管辖 万国的；她的孩子被提到上帝和他宝座那里去。
REV|12|6|妇人就逃到旷野，在那里有上帝给她预备的地方，使她在那里被供养一千二百六十天。
REV|12|7|天上发生了争战。 米迦勒 同他的使者与龙作战，龙同它的使者也起来应战，
REV|12|8|它们都打败了，天上再也没有它们的地方。
REV|12|9|大龙就是那古蛇，名叫魔鬼，又叫撒但，是迷惑普天下的；它被摔在地上，它的使者也一同被摔下去。
REV|12|10|我听见在天上有大声音说： “我上帝的救恩、能力、国度， 和他所立的基督的权柄现在都来到了。 因为那个在我们上帝面前、 昼夜控告我们弟兄的， 已经被摔下去了。
REV|12|11|弟兄胜过那条龙是因羔羊的血， 和因自己所见证的道。 虽然至于死，他们也不惜自己的性命。
REV|12|12|所以，诸天和住在其中的， 你们都快乐吧！ 只是地和海有祸了！ 因为魔鬼知道自己的时候不多， 就气愤愤地下到你们那里去了。”
REV|12|13|龙见自己被摔在地上，就迫害那生男孩子的妇人。
REV|12|14|于是有大鹰的两个翅膀赐给妇人，让她能飞到旷野，到自己的地方，躲避那蛇。她在那里受供养一载二载半载。
REV|12|15|蛇在妇人背后，从口中喷出水来，像河一样，要将妇人冲走。
REV|12|16|地却帮助了妇人，开口吞了从龙口喷出来的水。
REV|12|17|于是龙向妇人发怒，去与她其余的儿女作战，就是与那些遵守上帝命令 、为耶稣作见证的 。
REV|12|18|那时龙站在海边沙滩上。
REV|13|1|我又看见一只兽从海里上来，有十个角七个头；在十个角上戴着十个冠冕，七个头上有亵渎的名号。
REV|13|2|我所看见的兽，形状像豹，脚像熊的脚，口像狮子的口。那条龙将自己的能力、座位和大权柄都给了它。
REV|13|3|我看见兽的七个头中，有一个似乎受了致命伤，那伤却医好了。全地的人都很惊讶，跟从了那只兽。
REV|13|4|他们都拜那条龙，因为它把自己的权柄给了兽；又拜那只兽，说：“谁能比这只兽，谁能与它交战呢？”
REV|13|5|龙又赐给那只兽说夸大亵渎话的口，又赐给它权柄可以任意行事四十二个月。
REV|13|6|那兽就开口向上帝说亵渎的话，亵渎上帝的名和他的帐幕，就是那些住在天上的。
REV|13|7|它又被准许与圣徒作战，并且得胜，也赐给它权柄，可以制伏各支派、各民族、各语言、各邦国。
REV|13|8|凡住在地上、名字从创世以来没有记在被杀羔羊的生命册上的人都要拜它。
REV|13|9|凡有耳朵的都听吧！
REV|13|10|该被掳掠的，必被掳掠； 该被刀杀的，必被刀杀。 在此，圣徒要有耐心和信心。
REV|13|11|我又看见另一只兽从地里上来。它有两个角如同羔羊，说话好像龙。
REV|13|12|它在第一只兽面前施行第一只兽所有的权柄，并且使地和住在地上的人拜那致命伤被医好了的第一只兽。
REV|13|13|这只兽又行大奇事，甚至在人面前使火从天降在地上。
REV|13|14|它得了权柄在第一只兽面前能行奇事，迷惑住在地上的人，告诉他们要为那受过刀伤还活着的兽造个像。
REV|13|15|又有权柄赐给它，让那只兽的像有生气，并且能说话，又使所有不拜兽像的人都被杀害。
REV|13|16|它又使众人，无论大小、贫富，自主的、为奴的，都在右手上，或是在额上，打一个印记；
REV|13|17|这样，除了那有印记，有兽的名或有兽名数字的，都不得买或卖。
REV|13|18|在此，要有智慧：让有悟性的人解开兽的数目吧，因为这是一个人的数字，那数字是六百六十六。
REV|14|1|我又观看，看见羔羊站在 锡安山 ，和他在一起的有十四万四千人，都有他的名和他父亲的名写在额上。
REV|14|2|我听见从天上有声音，像众水的声音和大雷的声音，我所听见的声音好像琴师所弹的琴声。
REV|14|3|他们在宝座前，和在四活物及众长老前唱新歌，除了从地上买来的那十四万四千人以外，没有人能学这歌。
REV|14|4|这些人未曾沾染妇女，他们原是童身。羔羊无论往哪里去，他们都跟随他。他们是从人间买来的，作为初熟的果子归给上帝和羔羊。
REV|14|5|在他们口中找不出谎言，他们是没有瑕疵的。
REV|14|6|我又看见另一位天使在空中飞翔，有永远的福音要传给住在地上的人，就是各邦国、各支派、各语言、各民族。
REV|14|7|他大声说：“要敬畏上帝，把荣耀归给他，因为他施行审判的时候已经到了。要敬拜那创造天、地、海和水源的主。”
REV|14|8|另有第二位天使接着说：“倾覆了！那曾叫列国喝淫乱、烈怒之酒的大 巴比伦 倾覆了！”
REV|14|9|另有第三位天使接着他们，大声说：“若有人拜那只兽和兽像，在额上或在手上受了印记，
REV|14|10|他也必喝上帝烈怒的酒；这酒是斟在上帝愤怒的杯中的纯酒。他要在圣天使和羔羊面前，在火与硫磺之中受痛苦。
REV|14|11|使他们受痛苦的烟往上冒，直到永永远远。那些拜兽和兽像，受了它名字的印记的人，昼夜不得安宁。”
REV|14|12|在此，遵守上帝命令 和坚信耶稣真道的圣徒要有耐心。
REV|14|13|我听见从天上有声音说：“你要写下：从今以后，在主里死去的人有福了。”圣灵说：“是的，他们要从自己的劳苦中得安息，因为工作的成果永随着他们。”
REV|14|14|我又观看，看见有一片白云，云上坐着一位好像是人子的，头上戴着金冠冕，手里拿着锋利的镰刀。
REV|14|15|另有一位天使从圣所出来，向那坐在云上的大声喊着：“伸出你的镰刀来收割吧，因为收割的时候已经到了，地上的庄稼已经熟透了。”
REV|14|16|于是那坐在云上的把镰刀向地上挥去，地上的庄稼就收割了。
REV|14|17|另有一位天使从天上的圣所出来，他也拿着锋利的镰刀。
REV|14|18|另有一位天使从祭坛出来，是有权柄管火的，向那拿着锋利镰刀的大声喊着说：“伸出锋利的镰刀来，收取地上葡萄树的果子，因为葡萄熟透了。”
REV|14|19|那天使就把镰刀向地上挥去，收取了地上的葡萄，扔进上帝愤怒的大醡酒池里。
REV|14|20|那醡酒池在城外被踹踏，有血从醡酒池里流出来，涨到马的嚼环那么高，约有一千六百斯他迪 那么远。
REV|15|1|我看见在天上有另一兆头，大而且奇，就是七位天使掌管末了的七种灾难，因为上帝的烈怒在这七种灾难中发尽了。
REV|15|2|我看见仿佛有搀杂火的玻璃海；又看见那些胜了那兽和兽像，以及它名字的数字的人，都站在玻璃海上，拿着上帝的竖琴。
REV|15|3|他们唱上帝仆人 摩西 的歌和羔羊的歌，说： “主—全能的上帝啊， 你的作为又伟大又奇妙！ 万国之王啊， 你的道路又公义又真实！
REV|15|4|主啊，谁敢不敬畏你， 不把荣耀归于你的名？ 因为只有你是神圣的。 万民都要来， 在你面前敬拜， 因你公义的作为已经彰显了。”
REV|15|5|此后，我看见在天上那存放法柜的圣所开了。
REV|15|6|那掌管七种灾难的七位天使从圣所出来，穿着洁白明亮的细麻衣 ，胸间束着金带。
REV|15|7|四个活物中，有一个把盛满了活到永永远远之上帝烈怒的七个金碗给了那七位天使。
REV|15|8|圣所中充满了上帝的荣耀和权能而来的烟。没有人能进入圣所，直等到那七位天使降完了七种灾难。
REV|16|1|我听见有大声音从圣所里出来，向那七位天使说：“你们去，把盛着上帝烈怒的七碗倾倒在地上。”
REV|16|2|第一位天使去，把碗倾倒在地上，就有又臭又毒的疮生在那些有兽的印记和拜兽像的人身上。
REV|16|3|第二位天使把碗倾倒在海里，海就变成像死人的血一样，海里所有的活物都死了。
REV|16|4|第三位天使把碗倾倒在河流和水源里，水就变成血了。
REV|16|5|我听见掌管众水的天使说： “昔在、今在的圣者啊， 你做的判断公义；
REV|16|6|因他们曾流过圣徒与先知的血， 现在你给他们血喝， 这是他们该受的。”
REV|16|7|我又听见祭坛中有声音说： “是的，主—全能的上帝啊， 你的判断又真实又公义！”
REV|16|8|第四位天使把碗倾倒在太阳上，使太阳可用火烤人。
REV|16|9|人被炎热所烤，就亵渎那有权掌管这些灾难的上帝的名，他们没有悔改，也没有把荣耀归给上帝。
REV|16|10|第五位天使把碗倾倒在兽的座位上，兽的国就变成黑暗。人因疼痛而咬自己的舌头；
REV|16|11|又因所受的疼痛和生的疮，就亵渎天上的上帝，也没有为他们的行为悔改。
REV|16|12|第六位天使把碗倾倒在大 幼发拉底河 上，河水就干了，为要给从日出之地所来的众王预备道路。
REV|16|13|我又看见三个污秽的灵，好像青蛙，从龙的口、兽的口和假先知的口中出来。
REV|16|14|他们本是鬼魔的灵，施行奇事，到普天下众王那里去，召集他们在全能者上帝的大日子作战。
REV|16|15|看哪，我来像贼一样。那警醒、穿着衣服的人有福了；他不至于赤身而行，给人看见他的羞耻。
REV|16|16|于是，那三个鬼魔把众王聚集在 希伯来 话叫作 哈米吉多顿 的地方。
REV|16|17|第七位天使把碗倾倒在空中，就有大声音从圣所的宝座上出来，说：“成了！”
REV|16|18|又有闪电、响声、雷轰、大地震，自从地上有人以来没有这样大、这样厉害的地震。
REV|16|19|那大城裂为三段，列国的城也都倒塌了。上帝记起了大 巴比伦城 ，把那盛自己烈怒的酒杯递给她。
REV|16|20|各海岛都逃避了，众山也不见了。
REV|16|21|又有大冰雹从天掉落在人身上，每一个约重一他连得，以致人因冰雹的灾难而亵渎上帝，因为那灾难太大了。
REV|17|1|拿着七个碗的七位天使中，有一位前来对我说：“来，我要让你看那坐在众水之上的大淫妇所要受的惩罚；
REV|17|2|地上的君王都曾与她行淫，住在地上的人也喝醉了她淫乱的酒。”
REV|17|3|我在圣灵感动下，被天使带到旷野去，我看见一个女人骑在朱红色的兽上；那只兽有七个头十个角，遍体有亵渎的名号。
REV|17|4|那女人穿着紫色和朱红色的衣服，用金子、宝石、珍珠作妆饰，手拿着金杯，杯中盛满了可憎之物和她淫乱的污秽。
REV|17|5|在她额上写着奥秘的名字，说：“大 巴比伦 ，世上的淫妇和一切可憎之物的母。”
REV|17|6|我又看见那女人喝醉了圣徒的血和为耶稣作见证的人的血。 我看见她，非常诧异。
REV|17|7|天使对我说：“你为什么诧异呢？我要把这女人和驮着她那七头十角的兽的奥秘告诉你。
REV|17|8|你曾看见的兽，以前有，现在没有，将来要从无底坑里上来，又归于沉沦。凡住在地上、名字从创世以来没有记在生命册上的人看见那只兽都要诧异，因为它以前有，现在没有，以后再有。
REV|17|9|在此要有智慧的心思：那七个头就是女人所坐的七座山；他们又是七个王，
REV|17|10|五个已经倒了，一个还在，一个还没有来到；他来的时候必须只暂时停留。
REV|17|11|那以前有、现在没有的兽就是第八个，他也和那七个同列，正归于沉沦。
REV|17|12|你曾看见的那十个角就是十个王；他们还没有得到国度，但他们要和那只兽同得权柄作王一个时辰。
REV|17|13|他们同心把自己的能力权柄交给那只兽。
REV|17|14|他们将与羔羊作战，羔羊必胜过他们，因为羔羊是万主之主、万王之王，而同羔羊在一起的是蒙召、被选、忠心的人。”
REV|17|15|天使又对我说：“你所看见那淫妇坐的众水，就是许多民族、人民、邦国、语言。
REV|17|16|你所看见的那十个角与兽必恨这淫妇，他们要使她孤独赤身，又要吃她的肉，用火将她烧尽。
REV|17|17|因为上帝使诸王同心执行他的旨意，把他们自己的国交给那只兽，直等到上帝的话都应验了。
REV|17|18|你所看见的那女人就是管辖地上众王的大城。”
REV|18|1|此后，我看见另一位有大权柄的天使从天降下，地由于他的荣耀而发光。
REV|18|2|他以强而有力的声音喊着说： “倾覆了！大 巴比伦 倾覆了！ 她成了鬼魔的住处， 各样污秽之灵的巢穴， 各样污秽之鸟的窝， 各样污秽可憎之兽的出没处 。
REV|18|3|因为列国都喝了她淫乱大怒的酒 ； 地上的君王和她行淫； 地上的商人因她极度奢华而发了财。”
REV|18|4|我又听见另一个声音从天上说： “我的民哪，从那城出来吧！ 免得和她在罪上有份， 受她所受的灾殃；
REV|18|5|因她的罪恶滔天， 上帝已经记得她的不义。
REV|18|6|她怎样待人，也要怎样待她， 按她所行的加倍地报应她； 用她调酒的杯加倍调给她喝。
REV|18|7|她怎样荣耀自己，怎样奢华， 也要使她照样痛苦悲哀。 因她心里说： ‘我坐了皇后的位， 并不是寡妇， 绝不至于悲哀。’
REV|18|8|所以在一天之内，她的灾殃要一齐来到， 就是死亡、悲哀、饥荒。 她将被火烧尽， 因为审判她的主上帝大有能力。”
REV|18|9|地上的君王，与她行淫、一同奢华的，看见烧她的烟，就必为她哭泣哀号；
REV|18|10|因怕她的痛苦，就远远地站着，说： “祸哉，祸哉，这大城！ 坚固的 巴比伦城 啊！ 一时之间，你的审判要来到了。”
REV|18|11|地上的商人也都为她哭泣悲哀，因为没有人再买他们的货物了；
REV|18|12|这货物就是金、银、宝石、珍珠、细麻布、丝绸、紫色和朱红色衣料、各样香木、各样象牙的器皿、各样极宝贵的木头和铜、铁、大理石的器皿，
REV|18|13|和肉桂、豆蔻、香料、香膏、乳香、酒、油、细面、麦子、牛、羊、马、马车，以及奴隶、人口。
REV|18|14|“你所贪爱的果子离开了你； 你一切的珍馐美味和华美的物件 都从你那里毁灭， 绝对见不到了。”
REV|18|15|贩卖这些货物、藉着她发财的商人，因怕她的痛苦，就远远地站着哭泣悲哀，
REV|18|16|说： “祸哉，祸哉，这大城！ 她穿着细麻、 紫色、朱红色的衣服， 用金子、宝石、珍珠为妆饰。
REV|18|17|一时之间，这么多的财富就归于无有了。” 所有的船长和到处航海的，水手以及所有靠海为业的，都远远地站着，
REV|18|18|看见烧她的烟，就喊着说：“有哪一个城能跟这大城比呢？”
REV|18|19|于是他们把灰尘撒在头上，哭泣悲哀地喊着说： “祸哉，祸哉，这大城！ 凡有船在海中的， 都因她的珍宝成了富足。 她在一时之间就成为荒芜。
REV|18|20|天哪，众圣徒、众使徒、众先知啊！ 你们都要因她欢喜， 因为上帝已经在她身上为你们伸了冤。”
REV|18|21|有一位大力的天使举起一块石头，好像大磨石，扔在海里，说： “ 巴比伦 大城 也必这样猛力地被扔下去， 绝对见不到了。
REV|18|22|弹琴、歌唱、 吹笛、吹号的声音， 在你中间绝对听不见了； 各行手艺的技工 在你中间绝对见不到了； 推磨的声音 在你中间绝对听不见了；
REV|18|23|灯台的光 在你中间绝对不再照耀了； 新郎和新娘的声音 在你中间绝对听不见了。 你的商人原来是地上的显要； 万国也被你的邪术迷惑了。
REV|18|24|先知、圣徒和地上一切被杀的人的血都在这城里找到了。”
REV|19|1|此后，我听见好像有一大群人在天上大声说： “哈利路亚 ！ 救恩、荣耀、权能都属于我们的上帝。
REV|19|2|他的判断又真实又公义； 因他判断了那大淫妇， 她用淫行败坏了世界。 上帝为他的仆人伸冤， 向淫妇讨流仆人血的罪。”
REV|19|3|他们又一次说： “哈利路亚！ 烧淫妇的烟往上冒，直到永永远远。”
REV|19|4|那二十四位长老和四活物就俯伏敬拜坐在宝座上的上帝，说： “阿们。哈利路亚！”
REV|19|5|接着，有声音从宝座出来说： “上帝的众仆人哪， 凡敬畏他的， 无论大小， 都要赞美我们的上帝！”
REV|19|6|我听见好像一大群人的声音，像众水的声音，像大雷的声音，说： “哈利路亚！ 因为主─我们的上帝 、 全能者，作王了。
REV|19|7|我们要欢喜快乐， 将荣耀归给他； 因为羔羊的婚期到了， 他的新娘也自己预备好了，
REV|19|8|她蒙恩得穿明亮洁白的细麻衣： 这细麻衣就是圣徒们的义行。”
REV|19|9|天使对我说：“你要写下来：凡被请赴羔羊婚宴的人有福了！”他又对我说：“这些都是上帝真实的话。”
REV|19|10|我就俯伏在他脚前要拜他。他对我说：“千万不可！我和你，以及那些为耶稣作见证的弟兄同是仆人。你要敬拜上帝。”因为那些为耶稣作见证的人有预言的灵。
REV|19|11|后来我看见天开了。有一匹白马，骑在马上的称为 “诚信”、“真实”，他审判和争战都凭着公义。
REV|19|12|他的眼睛如 火焰，头上戴着许多冠冕；他身上写着一个名字，除了他自己没有人知道。
REV|19|13|他穿着浸过血的衣服；他的名称为“上帝之道”。
REV|19|14|众天军都骑着白马，穿着又白又洁净的细麻衣跟随他。
REV|19|15|有利剑从他口中出来，用来击打列国。他要用铁杖管辖 他们，并且要踹全能上帝烈怒的醡酒池。
REV|19|16|在他衣服和大腿上写着“万王之王，万主之主”的名号。
REV|19|17|我又看见一位天使站在太阳中，向天空一切的飞鸟大声喊着说：“你们聚集来赴上帝的大宴席，
REV|19|18|为要吃君王的肉、将军的肉、壮士的肉、马和骑士的肉、一切自主的和为奴的，以及尊贵的和卑贱的肉。”
REV|19|19|我又看见那兽和地上的君王，和他们的军队都聚集，要与白马骑士和他的军队作战。
REV|19|20|那兽被擒拿了；那在兽面前曾行奇事、迷惑了接受兽的印记和拜兽像的人的假先知，也与兽同被擒拿。他们两个就活生生地被扔进烧着硫磺的火湖里，
REV|19|21|其余的人被白马骑士口中吐出来的剑杀了；所有的飞鸟都吃饱了他们的肉。
REV|20|1|我又看见一位天使从天降下，手里拿着无底坑的钥匙和一条大铁链。
REV|20|2|他抓住那龙，那古蛇，就是魔鬼、撒但，把它捆绑了一千年，
REV|20|3|扔在无底坑里，把无底坑关闭，用印封上，使它不再迷惑列国，等到那一千年满了。这些事以后，它必须暂时被释放。
REV|20|4|我又看见一些宝座，坐在上面的有审判的权柄赐给他们。我又看见那些因为给耶稣作见证，并为上帝之道被斩首的人的灵魂，和没有拜过那兽与兽像、也没有在额上和手上打过它印记的人的灵魂。他们都复活了，与基督一同作王一千年。
REV|20|5|这是头一次的复活。其余的死人还没有复活，直等那一千年满了。
REV|20|6|在头一次复活有份的有福了，圣洁了！第二次的死在他们身上没有权柄，但他们要作上帝和基督的祭司，也要与基督一同作王一千年。
REV|20|7|那一千年满了，撒但会从监牢里被释放，
REV|20|8|出来要迷惑地上四方的列国，就是 歌革 和 玛各 ，使他们聚集争战。他们的人数多如海沙。
REV|20|9|他们上来布满了全地，围住圣徒的营与蒙爱的城，就有火从天降下，烧灭了他们。
REV|20|10|那迷惑他们的魔鬼被扔进硫磺的火湖里，就是那兽和假先知所在的地方，他们会昼夜受折磨，直到永永远远。
REV|20|11|我又看见一个白色的大宝座和那坐在上面的；天和地都从他面前逃避，再也找不到它们的位置了。
REV|20|12|我又看见死了的人，无论大小，都站在宝座前。案卷都展开了，并另有一卷展开，就是生命册。死了的人都凭着这些案卷所记载的，照他们所行的受审判。
REV|20|13|于是海交出其中的死人，死亡和阴间也交出其中的死人；他们都照各人所行的受审判。
REV|20|14|死亡和阴间也被扔进火湖里，这火湖就是第二次的死。
REV|20|15|凡名字没有记在生命册上的人，就被扔进火湖里。
REV|21|1|我又看见一个新天新地，因为先前的天和先前的地已经过去了，海也不再有了。
REV|21|2|我又看见圣城，新 耶路撒冷 由上帝那里，从天而降，预备好了，就如新娘打扮整齐，等候丈夫。
REV|21|3|我听见有大声音从宝座出来，说： “看哪，上帝的帐幕在人间！ 他要和他们同住， 他们要作他的子民。 上帝要亲自与他们同在。
REV|21|4|上帝要擦去他们一切的眼泪； 不再有死亡， 也不再有悲哀、哭号、痛苦， 因为先前的事都过去了。”
REV|21|5|那位坐在宝座上的说：“看哪，我把一切都更新了！”他又说：“你要写下来，因为这些话是可信靠的，是真实的。”
REV|21|6|他又对我说：“成了！我是阿拉法，我是俄梅戛；我是开始，我是终结。我要把生命的泉水白白赐给那口渴的人喝。
REV|21|7|得胜的要承受这些为业；我要作他的上帝，他要作我的儿子。
REV|21|8|至于胆怯的、不信的、可憎的、杀人的、淫乱的、行邪术的、拜偶像的和一切说谎话的人，他们将在烧着硫磺的火湖里有份；这是第二次的死。”
REV|21|9|拿着七个金碗、盛满末后七种灾祸的七位天使中，有一位来对我说：“你来，我要给你看新娘，就是羔羊的妻子。”
REV|21|10|我在圣灵感动下，天使带我到一座高大的山，给我看由上帝那里、从天而降的圣城 耶路撒冷 ，
REV|21|11|这城有上帝的荣耀，它光辉如同极贵的宝石，好像碧玉，明如水晶。
REV|21|12|它有高大的墙，有十二个门，门上有十二位天使，门上又写着 以色列 人十二个支派的名字 。
REV|21|13|东边有三个门，北边有三个门，南边有三个门，西边有三个门。
REV|21|14|城墙有十二个根基，根基上有羔羊十二使徒的名字。
REV|21|15|那对我说话的天使拿着金的芦苇当尺，要量那城、城门和城墙。
REV|21|16|城是四方的，长宽一样。天使用芦苇量那城，共有一万二千斯他迪，长、宽、高都是一样。
REV|21|17|他又量了城墙，按着人的尺寸，就是天使的尺寸，共有一百四十四肘。
REV|21|18|墙是碧玉造的；城是纯金的，如同明净的玻璃。
REV|21|19|城墙的根基是用各样宝石修饰的：第一个根基是碧玉，第二是蓝宝石，第三是绿玛瑙，第四是绿宝石，
REV|21|20|第五是红玛瑙，第六是红宝石，第七是黄璧玺，第八是水苍玉，第九是红璧玺，第十是翡翠，第十一是紫玛瑙，第十二是紫晶。
REV|21|21|十二个门是十二颗珍珠；每一个门是一颗珍珠造的。城内的街道是纯金的，好像透明的玻璃。
REV|21|22|我没有看见城内有殿，因主—全能者上帝和羔羊就是城的殿。
REV|21|23|那城内不用日月光照，因为有上帝的荣耀光照，又有羔羊为城的灯。
REV|21|24|列国要藉着城的光行走；地上的君王要把自己的荣耀带给那城。
REV|21|25|城门白昼总不关闭，在那里没有黑夜。
REV|21|26|人要将列国的荣耀尊贵带给那城。
REV|21|27|凡不洁净的，和那行可憎与虚谎之事的人，都不得进那城，只有名字写在羔羊生命册上的才得进去。
REV|22|1|天使又让我看一道生命水的河，明亮如水晶，从上帝和羔羊的宝座流出来，
REV|22|2|经过城内街道的中央；在河的两边有生命树，结十二样 的果子，每月都结果子；树上的叶子可作医治万民之用。
REV|22|3|以后不再有任何诅咒。在城里将有上帝和羔羊的宝座。他的仆人都要事奉他，
REV|22|4|也要见他的面。他的名字将写在他们的额上。
REV|22|5|不再有黑夜；他们也不需要灯光或日光，因为主上帝要光照他们。他们要作王，直到永永远远。
REV|22|6|天使又对我说：“这些话是可信靠的，是真实的。主，就是赐灵感给众先知的上帝，差遣他的使者，要将必须快要发生的事指示他的众仆人。”
REV|22|7|“看哪，我必快来！凡遵守这书上预言的有福了。”
REV|22|8|这些事是我－ 约翰 所听见所看见的。当我听见看见时，就俯伏在指示我的天使脚前要拜他。
REV|22|9|他对我说：“千万不可！我与你和你的弟兄众先知，以及那些守这书上的话的人，同是作仆人。你要敬拜上帝。”
REV|22|10|他又对我说：“不可封了这书上的预言，因为时候近了。
REV|22|11|不义的，让他仍旧不义；污秽的，让他仍旧污秽；为义的，让他仍旧为义；圣洁的，让他仍旧圣洁。”
REV|22|12|“看哪，我必快来！赏罚在我，要照每个人所行的报应他。
REV|22|13|我是阿拉法，我是俄梅戛；我是首先的，我是末后的；我是开始，我是终结。”
REV|22|14|那些洗净自己衣服的有福了！他们可得权柄到生命树那里，也能从门进城。
REV|22|15|城外有犬类、行邪术的、淫乱的、杀人的、拜偶像的，以及所有喜爱和行虚谎的人。
REV|22|16|“我－耶稣差遣我的使者，为了众教会向你们证明这些事。我是 大卫 的根，是他的后裔；我是明亮的晨星。”
REV|22|17|圣灵和新娘都说：“来！”听见的人也要说：“来！”口渴的人也要来，愿意的人都可以白白取生命的水喝。
REV|22|18|我警告一切听见这书上预言的人：若有人在这预言上加添什么，上帝必将记在这书上的灾祸加在他身上。
REV|22|19|这书上的预言，若有人删去什么，上帝必从这书上所记的生命树和圣城删去他的份。
REV|22|20|证明这些事的说：“是的，我必快来！”阿们！主耶稣啊，我愿你来！
REV|22|21|愿主耶稣的恩惠与众圣徒同在。阿们！
