NUM|1|1|locutusque est Dominus ad Mosen in deserto Sinai in tabernaculo foederis prima die mensis secundi anno altero egressionis eorum ex Aegypto dicens
NUM|1|2|tollite summam universae congregationis filiorum Israhel per cognationes et domos suas et nomina singulorum quicquid sexus est masculini
NUM|1|3|a vicesimo anno et supra omnium virorum fortium ex Israhel et numerabitis eos per turmas suas tu et Aaron
NUM|1|4|eruntque vobiscum principes tribuum ac domorum in cognationibus suis
NUM|1|5|quorum ista sunt nomina de Ruben Elisur filius Sedeur
NUM|1|6|de Symeon Salamihel filius Surisaddai
NUM|1|7|de Iuda Naasson filius Aminadab
NUM|1|8|de Isachar Nathanahel filius Suar
NUM|1|9|de Zabulon Heliab filius Helon
NUM|1|10|filiorum autem Ioseph de Ephraim Helisama filius Ammiud de Manasse Gamalihel filius Phadassur
NUM|1|11|de Beniamin Abidan filius Gedeonis
NUM|1|12|de Dan Ahiezer filius Amisaddai
NUM|1|13|de Aser Phegihel filius Ochran
NUM|1|14|de Gad Heliasaph filius Duhel
NUM|1|15|de Nepthali Ahira filius Henan
NUM|1|16|hii nobilissimi principes multitudinis per tribus et cognationes suas et capita exercitus Israhel
NUM|1|17|quos tulerunt Moses et Aaron cum omni vulgi multitudine
NUM|1|18|et congregaverunt primo die mensis secundi recensentes eos per cognationes et domos ac familias et capita et nomina singulorum a vicesimo anno et supra
NUM|1|19|sicut praeceperat Dominus Mosi numeratique sunt in deserto Sinai
NUM|1|20|de Ruben primogenito Israhelis per generationes et familias ac domos suas et nomina capitum singulorum omne quod sexus est masculini a vicesimo anno et supra procedentium ad bellum
NUM|1|21|quadraginta sex milia quingenti
NUM|1|22|de filiis Symeon per generationes et familias ac domos cognationum suarum recensiti sunt per nomina et capita singulorum omne quod sexus est masculini a vicesimo anno et supra procedentium ad bellum
NUM|1|23|quinquaginta novem milia trecenti
NUM|1|24|de filiis Gad per generationes et familias ac domos cognationum suarum recensiti sunt per nomina singulorum a viginti annis et supra omnes qui ad bella procederent
NUM|1|25|quadraginta quinque milia sescenti quinquaginta
NUM|1|26|de filiis Iuda per generationes et familias ac domos cognationum suarum per nomina singulorum a vicesimo anno et supra omnes qui poterant ad bella procedere
NUM|1|27|recensiti sunt septuaginta quattuor milia sescenti
NUM|1|28|de filiis Isachar per generationes et familias ac domos cognationum suarum per nomina singulorum a vicesimo anno et supra omnes qui ad bella procederent
NUM|1|29|recensiti sunt quinquaginta quattuor milia quadringenti
NUM|1|30|de filiis Zabulon per generationes et familias ac domos cognationum suarum recensiti sunt per nomina singulorum a vicesimo anno et supra omnes qui poterant ad bella procedere
NUM|1|31|quinquaginta septem milia quadringenti
NUM|1|32|de filiis Ioseph filiorum Ephraim per generationes et familias ac domos cognationum suarum recensiti sunt per nomina singulorum a vicesimo anno et supra omnes qui poterant ad bella procedere
NUM|1|33|quadraginta milia quingenti
NUM|1|34|porro filiorum Manasse per generationes et familias ac domos cognationum suarum recensiti sunt per nomina singulorum a viginti annis et supra omnes qui poterant ad bella procedere
NUM|1|35|triginta duo milia ducenti
NUM|1|36|de filiis Beniamin per generationes et familias ac domos cognationum suarum recensiti sunt nominibus singulorum a vicesimo anno et supra omnes qui poterant ad bella procedere
NUM|1|37|triginta quinque milia quadringenti
NUM|1|38|de filiis Dan per generationes et familias ac domos cognationum suarum recensiti sunt nominibus singulorum a vicesimo anno et supra omnes qui poterant ad bella procedere
NUM|1|39|sexaginta duo milia septingenti
NUM|1|40|de filiis Aser per generationes et familias ac domos cognationum suarum recensiti sunt per nomina singulorum a vicesimo anno et supra omnes qui poterant ad bella procedere
NUM|1|41|quadraginta milia et mille quingenti
NUM|1|42|de filiis Nepthali per generationes et familias ac domos cognationum suarum recensiti sunt nominibus singulorum a vicesimo anno et supra omnes qui poterant ad bella procedere
NUM|1|43|quinquaginta tria milia quadringenti
NUM|1|44|hii sunt quos numeraverunt Moses et Aaron et duodecim principes Israhel singulos per domos cognationum suarum
NUM|1|45|fueruntque omnes filiorum Israhel per domos et familias suas a vicesimo anno et supra qui poterant ad bella procedere
NUM|1|46|sescenta tria milia virorum quingenti quinquaginta
NUM|1|47|Levitae autem in tribu familiarum suarum non sunt numerati cum eis
NUM|1|48|locutusque est Dominus ad Mosen dicens
NUM|1|49|tribum Levi noli numerare neque ponas summam eorum cum filiis Israhel
NUM|1|50|sed constitue eos super tabernaculum testimonii cuncta vasa eius et quicquid ad caerimonias pertinet ipsi portabunt tabernaculum et omnia utensilia eius et erunt in ministerio ac per gyrum tabernaculi metabuntur
NUM|1|51|cum proficiscendum fuerit deponent Levitae tabernaculum cum castra metanda erigent quisquis externorum accesserit occidetur
NUM|1|52|metabuntur autem castra filii Israhel unusquisque per turmas et cuneos atque exercitum suum
NUM|1|53|porro Levitae per gyrum tabernaculi figent tentoria ne fiat indignatio super multitudinem filiorum Israhel et excubabunt in custodiis tabernaculi testimonii
NUM|1|54|fecerunt ergo filii Israhel iuxta omnia quae praeceperat Dominus Mosi
NUM|2|1|locutusque est Dominus ad Mosen et Aaron dicens
NUM|2|2|singuli per turmas signa atque vexilla et domos cognationum suarum castrametabuntur filiorum Israhel per gyrum tabernaculi foederis
NUM|2|3|ad orientem Iudas figet tentoria per turmas exercitus sui eritque princeps filiorum eius Naasson filius Aminadab
NUM|2|4|et omnis de stirpe eius summa pugnantium septuaginta quattuor milia sescentorum
NUM|2|5|iuxta eum castrametati sunt de tribu Isachar quorum princeps fuit Nathanahel filius Suar
NUM|2|6|et omnis numerus pugnatorum eius quinquaginta quattuor milia quadringenti
NUM|2|7|in tribu Zabulon princeps fuit Heliab filius Helon
NUM|2|8|omnis de stirpe eius exercitus pugnatorum quinquaginta septem milia quadringenti
NUM|2|9|universi qui in castris Iudae adnumerati sunt fuerunt centum octoginta sex milia quadringenti et per turmas suas primi egredientur
NUM|2|10|in castris filiorum Ruben ad meridianam plagam erit princeps Elisur filius Sedeur
NUM|2|11|et cunctus exercitus pugnatorum eius qui numerati sunt quadraginta sex milia quingenti
NUM|2|12|iuxta eum castrametati sunt de tribu Symeon quorum princeps fuit Salamihel filius Surisaddai
NUM|2|13|et cunctus exercitus pugnatorum eius qui numerati sunt quinquaginta novem milia trecenti
NUM|2|14|in tribu Gad princeps fuit Heliasaph filius Duhel
NUM|2|15|et cunctus exercitus pugnatorum eius qui numerati sunt quadraginta quinque milia sescenti quinquaginta
NUM|2|16|omnes qui recensiti sunt in castris Ruben centum quinquaginta milia et mille quadringenti quinquaginta per turmas suas in secundo loco proficiscentur
NUM|2|17|levabitur autem tabernaculum testimonii per officia Levitarum et turmas eorum quomodo erigetur ita et deponetur singuli per loca et ordines suos proficiscentur
NUM|2|18|ad occidentalem plagam erunt castra filiorum Ephraim quorum princeps fuit Helisama filius Ammiud
NUM|2|19|cunctus exercitus pugnatorum eius qui numerati sunt quadraginta milia quingenti
NUM|2|20|et cum eis tribus filiorum Manasse quorum princeps fuit Gamalihel filius Phadassur
NUM|2|21|cunctus exercitus pugnatorum eius qui numerati sunt triginta duo milia ducenti
NUM|2|22|in tribu filiorum Beniamin princeps fuit Abidan filius Gedeonis
NUM|2|23|et cunctus exercitus pugnatorum eius qui recensiti sunt triginta quinque milia quadringenti
NUM|2|24|omnes qui numerati sunt in castris Ephraim centum octo milia centum per turmas suas tertii proficiscentur
NUM|2|25|ad aquilonis partem castrametati sunt filii Dan quorum princeps fuit Ahiezer filius Amisaddai
NUM|2|26|cunctus exercitus pugnatorum eius qui numerati sunt sexaginta duo milia septingenti
NUM|2|27|iuxta eum fixere tentoria de tribu Aser quorum princeps fuit Phegihel filius Ochran
NUM|2|28|cunctus exercitus pugnatorum eius qui numerati sunt quadraginta milia et mille quingenti
NUM|2|29|de tribu filiorum Nepthalim princeps fuit Ahira filius Henan
NUM|2|30|cunctus exercitus pugnatorum eius quinquaginta tria milia quadringenti
NUM|2|31|omnes qui numerati sunt in castris Dan fuerunt centum quinquaginta septem milia sescenti et novissimi proficiscentur
NUM|2|32|hic numerus filiorum Israhel per domos cognationum suarum et turmas divisi exercitus sescenta tria milia quingenti quinquaginta
NUM|2|33|Levitae autem non sunt numerati inter filios Israhel sic enim praecepit Dominus Mosi
NUM|2|34|feceruntque filii Israhel iuxta omnia quae mandaverat Dominus castrametati sunt per turmas suas et profecti per familias ac domos patrum suorum
NUM|3|1|haec sunt generationes Aaron et Mosi in die qua locutus est Dominus ad Mosen in monte Sinai
NUM|3|2|et haec nomina filiorum Aaron primogenitus eius Nadab dein Abiu et Eleazar et Ithamar
NUM|3|3|haec nomina filiorum Aaron sacerdotum qui uncti sunt et quorum repletae et consecratae manus ut sacerdotio fungerentur
NUM|3|4|mortui sunt Nadab et Abiu cum offerrent ignem alienum in conspectu Domini in deserto Sinai absque liberis functique sunt sacerdotio Eleazar et Ithamar coram Aaron patre suo
NUM|3|5|locutus est Dominus ad Mosen dicens
NUM|3|6|adplica tribum Levi et fac stare in conspectu Aaron sacerdotis ut ministrent ei et excubent
NUM|3|7|et observent quicquid ad cultum pertinet multitudinis coram tabernaculo testimonii
NUM|3|8|et custodiant vasa tabernaculi servientes in ministerio eius
NUM|3|9|dabisque dono Levitas
NUM|3|10|Aaron et filiis eius quibus traditi sunt a filiis Israhel Aaron autem et filios eius constitues super cultum sacerdotii externus qui ad ministrandum accesserit morietur
NUM|3|11|locutusque est Dominus ad Mosen dicens
NUM|3|12|ego tuli Levitas a filiis Israhel pro omni primogenito qui aperit vulvam in filiis Israhel eruntque Levitae mei
NUM|3|13|meum est enim omne primogenitum ex quo percussi primogenitos in terra Aegypti sanctificavi mihi quicquid primum nascitur in Israhel ab homine usque ad pecus mei sunt ego Dominus
NUM|3|14|locutus est Dominus ad Mosen in deserto Sinai dicens
NUM|3|15|numera filios Levi per domos patrum suorum et familias omnem masculum ab uno mense et supra
NUM|3|16|numeravit Moses ut praeceperat Dominus
NUM|3|17|et inventi sunt filii Levi per nomina sua Gerson et Caath et Merari
NUM|3|18|filii Gerson Lebni et Semei
NUM|3|19|filii Caath Amram et Iessaar Hebron et Ozihel
NUM|3|20|filii Merari Mooli et Musi
NUM|3|21|de Gerson fuere familiae duae lebnitica et semeitica
NUM|3|22|quarum numeratus est populus sexus masculini ab uno mense et supra septem milia quingentorum
NUM|3|23|hii post tabernaculum metabuntur ad occidentem
NUM|3|24|sub principe Eliasaph filio Lahel
NUM|3|25|et habebunt excubias in tabernaculo foederis
NUM|3|26|ipsum tabernaculum et operimentum eius tentorium quod trahitur ante fores tecti foederis et cortinas atrii tentorium quoque quod adpenditur in introitu atrii tabernaculi et quicquid ad ritum altaris pertinet funes tabernaculi et omnia utensilia eius
NUM|3|27|cognatio Caath habebit populos Amramitas et Iessaaritas et Hebronitas et Ozihelitas hae sunt familiae Caathitarum recensitae per nomina sua
NUM|3|28|omnes generis masculini ab uno mense et supra octo milia sescenti habebunt excubias sanctuarii
NUM|3|29|et castrametabuntur ad meridianam plagam
NUM|3|30|princepsque eorum erit Elisaphan filius Ozihel
NUM|3|31|et custodient arcam mensamque et candelabrum altaria et vasa sanctuarii in quibus ministratur et velum cunctamque huiuscemodi supellectilem
NUM|3|32|princeps autem principum Levitarum Eleazar filius Aaron sacerdotis erit super excubitores custodiae sanctuarii
NUM|3|33|at vero de Merari erunt populi Moolitae et Musitae recensiti per nomina sua
NUM|3|34|omnes generis masculini ab uno mense et supra sex milia ducenti
NUM|3|35|princeps eorum Surihel filius Abiahihel in plaga septentrionali castrametabuntur
NUM|3|36|erunt sub custodia eorum tabulae tabernaculi et vectes et columnae ac bases earum et omnia quae ad cultum huiuscemodi pertinent
NUM|3|37|columnaeque atrii per circuitum cum basibus suis et paxilli cum funibus
NUM|3|38|castrametabuntur ante tabernaculum foederis id est ad orientalem plagam Moses et Aaron cum filiis suis habentes custodiam sanctuarii in medio filiorum Israhel quisquis alienus accesserit morietur
NUM|3|39|omnes Levitae quos numeraverunt Moses et Aaron iuxta praeceptum Domini per familias suas in genere masculino a mense uno et supra fuerunt viginti duo milia
NUM|3|40|et ait Dominus ad Mosen numera primogenitos sexus masculini de filiis Israhel a mense uno et supra et habebis summam eorum
NUM|3|41|tollesque Levitas mihi pro omni primogenito filiorum Israhel ego sum Dominus et pecora eorum pro universis primogenitis pecoris filiorum Israhel
NUM|3|42|recensuit Moses sicut praeceperat Dominus primogenitos filiorum Israhel
NUM|3|43|et fuerunt masculi per nomina sua a mense uno et supra viginti duo milia ducenti septuaginta tres
NUM|3|44|locutusque est Dominus ad Mosen
NUM|3|45|tolle Levitas pro primogenitis filiorum Israhel et pecora Levitarum pro pecoribus eorum eruntque Levitae mei ego sum Dominus
NUM|3|46|in pretio autem ducentorum septuaginta trium qui excedunt numerum Levitarum de primogenitis filiorum Israhel
NUM|3|47|accipies quinque siclos per singula capita ad mensuram sanctuarii siclus habet obolos viginti
NUM|3|48|dabisque pecuniam Aaron et filiis eius pretium eorum qui supra sunt
NUM|3|49|tulit igitur Moses pecuniam eorum qui fuerant amplius et quos redemerant a Levitis
NUM|3|50|pro primogenitis filiorum Israhel mille trecentorum sexaginta quinque siclorum iuxta pondus sanctuarii
NUM|3|51|et dedit eam Aaroni et filiis eius iuxta verbum quod praeceperat sibi Dominus
NUM|4|1|locutusque est Dominus ad Mosen et Aaron dicens
NUM|4|2|tolle summam filiorum Caath de medio Levitarum per domos et familias suas
NUM|4|3|a tricesimo anno et supra usque ad quinquagesimum annum omnium qui ingrediuntur ut stent et ministrent in tabernaculo foederis
NUM|4|4|hic est cultus filiorum Caath tabernaculum foederis et sanctum sanctorum
NUM|4|5|ingredientur Aaron et filii eius quando movenda sunt castra et deponent velum quod pendet ante fores involventque eo arcam testimonii
NUM|4|6|et operient rursum velamine ianthinarum pellium extendentque desuper pallium totum hyacinthinum et inducent vectes
NUM|4|7|mensam quoque propositionis involvent hyacinthino pallio et ponent cum ea turibula et mortariola cyatos et crateras ad liba fundenda panes semper in ea erunt
NUM|4|8|extendentque desuper pallium coccineum quod rursum operient velamento ianthinarum pellium et inducent vectes
NUM|4|9|sument et pallium hyacinthinum quo operient candelabrum cum lucernis et forcipibus suis et emunctoriis et cunctis vasis olei quae ad concinnandas lucernas necessaria sunt
NUM|4|10|et super omnia ponent operimentum ianthinarum pellium et inducent vectes
NUM|4|11|nec non et altare aureum involvent hyacinthino vestimento et extendent desuper operimentum ianthinarum pellium inducentque vectes
NUM|4|12|omnia vasa quibus ministratur in sanctuario involvent hyacinthino pallio et extendent desuper operimentum ianthinarum pellium inducentque vectes
NUM|4|13|sed et altare mundabunt cinere et involvent illud purpureo vestimento
NUM|4|14|ponentque cum eo omnia vasa quibus in ministerio eius utuntur id est ignium receptacula fuscinulas ac tridentes uncinos et vatilla cuncta vasa altaris operient simul velamine ianthinarum pellium et inducent vectes
NUM|4|15|cumque involverint Aaron et filii eius sanctuarium et omnia vasa eius in commotione castrorum tunc intrabunt filii Caath ut portent involuta et non tangant vasa sanctuarii ne moriantur ista sunt onera filiorum Caath in tabernaculo foederis
NUM|4|16|super quos erit Eleazar filius Aaron sacerdotis ad cuius pertinet curam oleum ad concinnandas lucernas et conpositionis incensum et sacrificium quod semper offertur et oleum unctionis et quicquid ad cultum tabernaculi pertinet omniumque vasorum quae in sanctuario sunt
NUM|4|17|locutusque est Dominus ad Mosen et Aaron dicens
NUM|4|18|nolite perdere populum Caath de medio Levitarum
NUM|4|19|sed hoc facite eis ut vivant et non moriantur si tetigerint sancta sanctorum Aaron et filii eius intrabunt ipsique disponent opera singulorum et divident quid portare quis debeat
NUM|4|20|alii nulla curiositate videant quae sunt in sanctuario priusquam involvantur alioquin morientur
NUM|4|21|locutus est Dominus ad Mosen dicens
NUM|4|22|tolle summam etiam filiorum Gerson per domos ac familias et cognationes suas
NUM|4|23|a triginta annis et supra usque ad annos quinquaginta numera omnes qui ingrediuntur et ministrant in tabernaculo foederis
NUM|4|24|hoc est officium familiae Gersonitarum
NUM|4|25|ut portent cortinas tabernaculi et tectum foederis operimentum aliud et super omnia velamen ianthinum tentoriumque quod pendet in introitu foederis tabernaculi
NUM|4|26|cortinas atrii et velum in introitu quod est ante tabernaculum omnia quae ad altare pertinent funiculos et vasa ministerii
NUM|4|27|iubente Aaron et filiis eius portabunt filii Gerson et scient singuli cui debeant oneri mancipari
NUM|4|28|hic est cultus familiae Gersonitarum in tabernaculo foederis eruntque sub manu Ithamar filii Aaron sacerdotis
NUM|4|29|filios quoque Merari per familias et domos patrum suorum recensebis
NUM|4|30|a triginta annis et supra usque ad annos quinquaginta omnes qui ingrediuntur ad officium ministerii sui et cultum foederis testimonii
NUM|4|31|haec sunt onera eorum portabunt tabulas tabernaculi et vectes eius columnas et bases earum
NUM|4|32|columnas quoque atrii per circuitum cum basibus et paxillis et funibus suis omnia vasa et supellectilem ad numerum accipient sicque portabunt
NUM|4|33|hoc est officium familiae Meraritarum et ministerium in tabernaculo foederis eruntque sub manu Ithamar filii Aaron sacerdotis
NUM|4|34|recensuerunt igitur Moses et Aaron et principes synagogae filios Caath per cognationes et domos patrum suorum
NUM|4|35|a triginta annis et supra usque ad annum quinquagesimum omnes qui ingrediuntur ad ministerium tabernaculi foederis
NUM|4|36|et inventi sunt duo milia septingenti quinquaginta
NUM|4|37|hic est numerus populi Caath qui intrat tabernaculum foederis hos numeravit Moses et Aaron iuxta sermonem Domini per manum Mosi
NUM|4|38|numerati sunt et filii Gerson per cognationes et domos patrum suorum
NUM|4|39|a triginta annis et supra usque ad annum quinquagesimum omnes qui ingrediuntur ut ministrent in tabernaculo foederis
NUM|4|40|et inventi sunt duo milia sescenti triginta
NUM|4|41|hic est populus Gersonitarum quos numeraverunt Moses et Aaron iuxta verbum Domini
NUM|4|42|numerati sunt et filii Merari per cognationes et domos patrum suorum
NUM|4|43|a triginta annis et supra usque ad annum quinquagesimum omnes qui ingrediuntur ad explendos ritus tabernaculi foederis
NUM|4|44|et inventi sunt tria milia ducenti
NUM|4|45|hic est numerus filiorum Merari quos recensuerunt Moses et Aaron iuxta imperium Domini per manum Mosi
NUM|4|46|omnes qui recensiti sunt de Levitis et quos fecit ad nomen Moses et Aaron et principes Israhel per cognationes et domos patrum suorum
NUM|4|47|a triginta annis et supra usque ad annum quinquagesimum ingredientes ad ministerium tabernaculi et onera portanda
NUM|4|48|fuerunt simul octo milia quingenti octoginta
NUM|4|49|iuxta verbum Domini recensuit eos Moses unumquemque iuxta officium et onera sua sicut praeceperat ei Dominus
NUM|5|1|locutusque est Dominus ad Mosen dicens
NUM|5|2|praecipe filiis Israhel ut eiciant de castris omnem leprosum et qui semine fluit pollutusque est super mortuo
NUM|5|3|tam masculum quam feminam eicite de castris ne contaminent ea cum habitaverim vobiscum
NUM|5|4|feceruntque ita filii Israhel et eiecerunt eos extra castra sicut locutus erat Dominus Mosi
NUM|5|5|locutus est Dominus ad Mosen dicens
NUM|5|6|loquere ad filios Israhel vir sive mulier cum fecerint ex omnibus peccatis quae solent hominibus accidere et per neglegentiam transgressi fuerint mandatum Domini atque deliquerint
NUM|5|7|confitebuntur peccatum suum et reddent ipsum caput quintamque partem desuper ei in quem peccaverint
NUM|5|8|sin autem non fuerit qui recipiat dabunt Domino et erit sacerdotis excepto ariete qui offertur pro expiatione ut sit placabilis hostia
NUM|5|9|omnes quoque primitiae quas offerunt filii Israhel ad sacerdotem pertinent
NUM|5|10|et quicquid in sanctuarium offertur a singulis et traditur manibus sacerdotis ipsius erit
NUM|5|11|locutus est Dominus ad Mosen dicens
NUM|5|12|loquere ad filios Israhel et dices ad eos vir cuius uxor erraverit maritumque contemnens
NUM|5|13|dormierit cum altero viro et hoc maritus deprehendere non quiverit sed latet adulterium et testibus argui non potest quia non est inventa in stupro
NUM|5|14|si spiritus zelotypiae concitaverit virum contra uxorem suam quae vel polluta est vel falsa suspicione appetitur
NUM|5|15|adducet eam ad sacerdotem et offeret oblationem pro illa decimam partem sati farinae hordiaciae non fundet super eam oleum nec inponet tus quia sacrificium zelotypiae est et oblatio investigans adulterium
NUM|5|16|offeret igitur eam sacerdos et statuet coram Domino
NUM|5|17|adsumetque aquam sanctam in vase fictili et pauxillum terrae de pavimento tabernaculi mittet in eam
NUM|5|18|cumque steterit mulier in conspectu Domini discoperiet caput eius et ponet super manus illius sacrificium recordationis et oblationem zelotypiae ipse autem tenebit aquas amarissimas in quibus cum execratione maledicta congessit
NUM|5|19|adiurabitque eam et dicet si non dormivit vir alienus tecum et si non polluta es deserto mariti toro non te nocebunt aquae istae amarissimae in quas maledicta congessi
NUM|5|20|sin autem declinasti a viro tuo atque polluta es et concubuisti cum altero
NUM|5|21|his maledictionibus subiacebis det te Dominus in maledictionem exemplumque cunctorum in populo suo putrescere faciat femur tuum et tumens uterus disrumpatur
NUM|5|22|ingrediantur aquae maledictae in ventrem tuum et utero tumescente putrescat femur et respondebit mulier amen amen
NUM|5|23|scribetque sacerdos in libello ista maledicta et delebit ea aquis amarissimis in quas maledicta congessit
NUM|5|24|et dabit ei bibere quas cum exhauserit
NUM|5|25|tollet sacerdos de manu eius sacrificium zelotypiae et elevabit illud coram Domino inponetque super altare ita dumtaxat ut prius
NUM|5|26|pugillum sacrificii tollat de eo quod offertur et incendat super altare et sic potum det mulieri aquas amarissimas
NUM|5|27|quas cum biberit si polluta est et contempto viro adulterii rea pertransibunt eam aquae maledictionis et inflato ventre conputrescet femur eritque mulier in maledictionem et in exemplum omni populo
NUM|5|28|quod si polluta non fuerit erit innoxia et faciet liberos
NUM|5|29|ista est lex zelotypiae si declinaverit mulier a viro suo et si polluta fuerit
NUM|5|30|maritusque zelotypiae spiritu concitatus adduxerit eam in conspectu Domini et fecerit ei sacerdos iuxta omnia quae scripta sunt
NUM|5|31|maritus absque culpa erit et illa recipiet iniquitatem suam
NUM|6|1|locutus est Dominus ad Mosen dicens
NUM|6|2|loquere ad filios Israhel et dices ad eos vir sive mulier cum fecerit votum ut sanctificentur et se voluerint Domino consecrare
NUM|6|3|vino et omni quod inebriare potest abstinebunt acetum ex vino et ex qualibet alia potione et quicquid de uva exprimitur non bibent uvas recentes siccasque non comedent
NUM|6|4|cunctis diebus quibus ex voto Domino consecrantur quicquid ex vinea esse potest ab uva passa usque ad acinum non comedent
NUM|6|5|omni tempore separationis suae novacula non transibit super caput eius usque ad conpletum diem quo Domino consecratur sanctus erit crescente caesarie capitis eius
NUM|6|6|omni tempore consecrationis suae super mortuum non ingredietur
NUM|6|7|nec super patris quidem et matris et fratris sororisque funere contaminabitur quia consecratio Dei sui super caput eius est
NUM|6|8|omnes dies separationis suae sanctus erit Domino
NUM|6|9|sin autem mortuus fuerit subito quispiam coram eo polluetur caput consecrationis eius quod radet ilico et in eadem die purgationis suae et rursum septima
NUM|6|10|in octavo autem die offeret duos turtures vel duos pullos columbae sacerdoti in introitu foederis testimonii
NUM|6|11|facietque sacerdos unum pro peccato et alterum in holocaustum et deprecabitur pro eo quia peccavit super mortuo sanctificabitque caput eius in die illo
NUM|6|12|et consecrabit Domino dies separationis illius offerens agnum anniculum pro peccato ita tamen ut dies priores irriti fiant quoniam polluta est sanctificatio eius
NUM|6|13|ista est lex consecrationis cum dies quos ex voto decreverat conplebuntur adducet eum ad ostium tabernaculi foederis
NUM|6|14|et offeret oblationem eius Domino agnum anniculum inmaculatum in holocaustum et ovem anniculam inmaculatam pro peccato et arietem inmaculatum hostiam pacificam
NUM|6|15|canistrum quoque panum azymorum qui conspersi sunt oleo et lagana absque fermento uncta oleo ac libamina singulorum
NUM|6|16|quae offeret sacerdos coram Domino et faciet tam pro peccato quam in holocaustum
NUM|6|17|arietem vero immolabit hostiam pacificam Domino offerens simul canistrum azymorum et libamenta quae ex more debentur
NUM|6|18|tunc radetur nazareus ante ostium tabernaculi foederis caesarie consecrationis suae tolletque capillos eius et ponet super ignem qui est subpositus sacrificio pacificorum
NUM|6|19|et armum coctum arietis tortamque absque fermento unam de canistro et laganum azymum unum et tradet in manibus nazarei postquam rasum fuerit caput eius
NUM|6|20|susceptaque rursum ab eo elevabit in conspectu Domini et sanctificata sacerdotis erunt sicut pectusculum quod separari iussum est et femur post haec potest bibere nazareus vinum
NUM|6|21|ista est lex nazarei cum voverit oblationem suam Domino tempore consecrationis suae exceptis his quae invenerit manus eius iuxta quod mente devoverat ita faciet ad perfectionem sanctificationis suae
NUM|6|22|locutus est Dominus ad Mosen dicens
NUM|6|23|loquere Aaron et filiis eius sic benedicetis filiis Israhel et dicetis eis
NUM|6|24|benedicat tibi Dominus et custodiat te
NUM|6|25|ostendat Dominus faciem suam tibi et misereatur tui
NUM|6|26|convertat Dominus vultum suum ad te et det tibi pacem
NUM|6|27|invocabunt nomen meum super filios Israhel et ego benedicam eis
NUM|7|1|factum est autem in die qua conplevit Moses tabernaculum et erexit illud unxitque et sanctificavit cum omnibus vasis suis altare similiter et vasa eius
NUM|7|2|obtulerunt principes Israhel et capita familiarum qui erant per singulas tribus praefecti eorum qui numerati fuerant
NUM|7|3|munera coram Domino sex plaustra tecta cum duodecim bubus unum plaustrum obtulere duo duces et unum bovem singuli obtuleruntque ea in conspectu tabernaculi
NUM|7|4|ait autem Dominus ad Mosen
NUM|7|5|suscipe ab eis ut serviant in ministerio tabernaculi et tradas ea Levitis iuxta ordinem ministerii sui
NUM|7|6|itaque cum suscepisset Moses plaustra et boves tradidit eos Levitis
NUM|7|7|duo plaustra et quattuor boves dedit filiis Gerson iuxta id quod habebant necessarium
NUM|7|8|quattuor alia plaustra et octo boves dedit filiis Merari secundum officia et cultum suum sub manu Ithamar filii Aaron sacerdotis
NUM|7|9|filiis autem Caath non dedit plaustra et boves quia in sanctuario serviunt et onera propriis portant umeris
NUM|7|10|igitur obtulerunt duces in dedicationem altaris die qua unctum est oblationem suam ante altare
NUM|7|11|dixitque Dominus ad Mosen singuli duces per singulos dies offerant munera in dedicationem altaris
NUM|7|12|primo die obtulit oblationem suam Naasson filius Aminadab de tribu Iuda
NUM|7|13|fueruntque in ea acetabulum argenteum pondo centum triginta siclorum fiala argentea habens septuaginta siclos iuxta pondus sanctuarii utrumque plenum simila conspersa oleo in sacrificium
NUM|7|14|mortariolum ex decem siclis aureis plenum incenso
NUM|7|15|bovem et arietem et agnum anniculum in holocaustum
NUM|7|16|hircumque pro peccato
NUM|7|17|et in sacrificio pacificorum boves duos arietes quinque hircos quinque agnos anniculos quinque haec est oblatio Naasson filii Aminadab
NUM|7|18|secundo die obtulit Nathanahel filius Suar dux de tribu Isachar
NUM|7|19|acetabulum argenteum adpendens centum triginta siclos fialam argenteam habentem septuaginta siclos iuxta pondus sanctuarii utrumque plenum simila conspersa oleo in sacrificium
NUM|7|20|mortariolum aureum habens decem siclos plenum incenso
NUM|7|21|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|22|hircumque pro peccato
NUM|7|23|et in sacrificio pacificorum boves duos arietes quinque hircos quinque agnos anniculos quinque haec fuit oblatio Nathanahel filii Suar
NUM|7|24|tertio die princeps filiorum Zabulon Heliab filius Helon
NUM|7|25|obtulit acetabulum argenteum adpendens centum triginta siclos fialam argenteam habentem septuaginta siclos ad pondus sanctuarii utrumque plenum simila conspersa oleo in sacrificium
NUM|7|26|mortariolum aureum adpendens decem siclos plenum incenso
NUM|7|27|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|28|hircumque pro peccato
NUM|7|29|et in sacrificio pacificorum boves duos arietes quinque hircos quinque agnos anniculos quinque haec est oblatio Heliab filii Helon
NUM|7|30|die quarto princeps filiorum Ruben Helisur filius Sedeur
NUM|7|31|obtulit acetabulum argenteum adpendens centum triginta siclos fialam argenteam habentem septuaginta siclos ad pondus sanctuarii utrumque plenum simila conspersa oleo in sacrificium
NUM|7|32|mortariolum aureum adpendens decem siclos plenum incenso
NUM|7|33|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|34|hircumque pro peccato
NUM|7|35|et in hostias pacificorum boves duos arietes quinque hircos quinque agnos anniculos quinque haec fuit oblatio Helisur filii Sedeur
NUM|7|36|die quinto princeps filiorum Symeon Salamihel filius Surisaddai
NUM|7|37|obtulit acetabulum argenteum adpendens centum triginta siclos fialam argenteam habentem septuaginta siclos ad pondus sanctuarii utrumque plenum simila conspersa oleo in sacrificium
NUM|7|38|mortariolum aureum adpendens decem siclos plenum incenso
NUM|7|39|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|40|hircumque pro peccato
NUM|7|41|et in hostias pacificorum boves duos arietes quinque hircos quinque agnos anniculos quinque haec fuit oblatio Salamihel filii Surisaddai
NUM|7|42|die sexto princeps filiorum Gad Heliasaph filius Duhel
NUM|7|43|obtulit acetabulum argenteum adpendens centum triginta siclos fialam argenteam habentem septuaginta siclos ad pondus sanctuarii utrumque plenum simila conspersa oleo in sacrificium
NUM|7|44|mortariolum aureum adpendens siclos decem plenum incenso
NUM|7|45|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|46|hircumque pro peccato
NUM|7|47|et in hostias pacificorum boves duos arietes quinque hircos quinque agnos anniculos quinque haec fuit oblatio Heliasaph filii Duhel
NUM|7|48|die septimo princeps filiorum Ephraim Helisama filius Ammiud
NUM|7|49|obtulit acetabulum argenteum adpendens centum triginta siclos fialam argenteam habentem septuaginta siclos ad pondus sanctuarii utrumque plenum simila conspersa oleo in sacrificium
NUM|7|50|mortariolum aureum adpendens decem siclos plenum incenso
NUM|7|51|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|52|hircumque pro peccato
NUM|7|53|et in hostias pacificas boves duos arietes quinque hircos quinque agnos anniculos quinque haec fuit oblatio Helisama filii Ammiud
NUM|7|54|die octavo princeps filiorum Manasse Gamalihel filius Phadassur
NUM|7|55|obtulit acetabulum argenteum adpendens centum triginta siclos fialam argenteam habentem septuaginta siclos ad pondus sanctuarii utrumque plenum simila conspersa oleo in sacrificium
NUM|7|56|mortariolum aureum adpendens decem siclos plenum incenso
NUM|7|57|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|58|hircumque pro peccato
NUM|7|59|et in hostias pacificorum boves duos arietes quinque hircos quinque agnos anniculos quinque haec fuit oblatio Gamalihel filii Phadassur
NUM|7|60|die nono princeps filiorum Beniamin Abidan filius Gedeonis
NUM|7|61|obtulit acetabulum argenteum adpendens centum triginta siclos fialam argenteam habentem septuaginta siclos ad pondus sanctuarii utrumque plenum simila conspersa oleo in sacrificium
NUM|7|62|mortariolum aureum adpendens decem siclos plenum incenso
NUM|7|63|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|64|hircumque pro peccato
NUM|7|65|et in hostias pacificorum boves duos arietes quinque hircos quinque agnos anniculos quinque haec fuit oblatio Abidan filii Gedeonis
NUM|7|66|die decimo princeps filiorum Dan Ahiezer filius Amisaddai
NUM|7|67|obtulit acetabulum argenteum adpendens centum triginta siclos fialam argenteam habentem septuaginta siclos ad pondus sanctuarii utrumque plenum simila conspersa oleo in sacrificium
NUM|7|68|mortariolum aureum adpendens decem siclos plenum incenso
NUM|7|69|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|70|hircumque pro peccato
NUM|7|71|et in hostias pacificorum boves duos arietes quinque hircos quinque agnos anniculos quinque haec fuit oblatio Ahiezer filii Amisaddai
NUM|7|72|die undecimo princeps filiorum Aser Phagaihel filius Ochran
NUM|7|73|obtulit acetabulum argenteum adpendens centum triginta siclos fialam argenteam habentem septuaginta siclos ad pondus sanctuarii utrumque plenum simila conspersa oleo in sacrificium
NUM|7|74|mortariolum aureum adpendens decem siclos plenum incenso
NUM|7|75|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|76|hircumque pro peccato
NUM|7|77|et in hostias pacificorum boves duos arietes quinque hircos quinque agnos anniculos quinque haec fuit oblatio Phagaihel filii Ochran
NUM|7|78|die duodecimo princeps filiorum Nepthalim Achira filius Henan
NUM|7|79|obtulit acetabulum argenteum adpendens centum triginta siclos fialam argenteam habentem septuaginta siclos ad pondus sanctuarii utrumque plenum simila conspersa oleo in sacrificium
NUM|7|80|mortariolum aureum adpendens decem siclos plenum incenso
NUM|7|81|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|82|hircumque pro peccato
NUM|7|83|et in hostias pacificorum boves duos arietes quinque hircos quinque agnos anniculos quinque haec fuit oblatio Achira filii Henan
NUM|7|84|haec in dedicatione altaris oblata sunt a principibus Israhel in die qua consecratum est acetabula argentea duodecim fialae argenteae duodecim mortariola aurea duodecim
NUM|7|85|ita ut centum triginta argenti siclos haberet unum acetabulum et septuaginta siclos una fiala id est in commune vasorum omnium ex argento sicli duo milia quadringenti pondere sanctuarii
NUM|7|86|mortariola aurea duodecim plena incenso denos siclos adpendentia pondere sanctuarii id est simul auri sicli centum viginti
NUM|7|87|boves de armento in holocaustum duodecim arietes duodecim agni anniculi duodecim et libamenta eorum hirci duodecim pro peccato
NUM|7|88|hostiae pacificorum boves viginti quattuor arietes sexaginta hirci sexaginta agni anniculi sexaginta haec oblata sunt in dedicatione altaris quando unctum est
NUM|7|89|cumque ingrederetur Moses tabernaculum foederis ut consuleret oraculum audiebat vocem loquentis ad se de propitiatorio quod erat super arcam testimonii inter duos cherubin unde et loquebatur ei
NUM|8|1|locutus est Dominus ad Mosen dicens
NUM|8|2|loquere Aaroni et dices ad eum cum posueris septem lucernas contra eam partem quam candelabrum respicit lucere debebunt
NUM|8|3|fecitque Aaron et inposuit lucernas super candelabrum ut praeceperat Dominus Mosi
NUM|8|4|haec autem erat factura candelabri ex auro ductili tam medius stipes quam cuncta ex utroque calamorum latera nascebantur iuxta exemplum quod ostendit Dominus Mosi ita operatus est candelabrum
NUM|8|5|et locutus est Dominus ad Mosen dicens
NUM|8|6|tolle Levitas de medio filiorum Israhel et purificabis eos
NUM|8|7|iuxta hunc ritum aspergantur aqua lustrationis et radant omnes pilos carnis suae cumque laverint vestimenta sua et mundati fuerint
NUM|8|8|tollant bovem de armentis et libamentum eius similam oleo conspersam bovem autem alterum de armento tu accipies pro peccato
NUM|8|9|et adplicabis Levitas coram tabernaculo foederis convocata omni multitudine filiorum Israhel
NUM|8|10|cumque Levitae fuerint coram Domino ponent filii Israhel manus suas super eos
NUM|8|11|et offeret Aaron Levitas munus in conspectu Domini a filiis Israhel ut serviant in ministerio eius
NUM|8|12|Levitae quoque ponent manus suas super capita boum e quibus unum facies pro peccato et alterum in holocaustum Domini ut depreceris pro eis
NUM|8|13|statuesque Levitas in conspectu Aaron et filiorum eius et consecrabis oblatos Domino
NUM|8|14|ac separabis de medio filiorum Israhel ut sint mei
NUM|8|15|et postea ingrediantur tabernaculum foederis ut serviant mihi sicque purificabis et consecrabis eos in oblationem Domini quoniam dono donati sunt mihi a filiis Israhel
NUM|8|16|pro primogenitis quae aperiunt omnem vulvam in Israhel accepi eos
NUM|8|17|mea sunt omnia primogenita filiorum Israhel tam ex hominibus quam ex iumentis ex die quo percussi omnem primogenitum in terra Aegypti sanctificavi eos mihi
NUM|8|18|et tuli Levitas pro cunctis primogenitis filiorum Israhel
NUM|8|19|tradidique eos dono Aaroni et filiis eius de medio populi ut serviant mihi pro Israhel in tabernaculo foederis et orent pro eis ne sit in populo plaga si ausi fuerint accedere ad sanctuarium
NUM|8|20|feceruntque Moses et Aaron et omnis multitudo filiorum Israhel super Levitas quae praeceperat Dominus Mosi
NUM|8|21|purificatique sunt et laverunt vestimenta sua elevavitque eos Aaron in conspectu Domini et oravit pro eis
NUM|8|22|ut purificati ingrederentur ad officia sua in tabernaculum foederis coram Aaron et filiis eius sicut praeceperat Dominus Mosi de Levitis ita factum est
NUM|8|23|locutus est Dominus ad Mosen dicens
NUM|8|24|haec est lex Levitarum a viginti quinque annis et supra ingredientur ut ministrent in tabernaculo foederis
NUM|8|25|cumque quinquagesimum annum aetatis impleverint servire cessabunt
NUM|8|26|eruntque ministri fratrum suorum in tabernaculo foederis ut custodiant quae sibi fuerint commendata opera autem ipsa non faciant sic dispones Levitas in custodiis suis
NUM|9|1|locutus est Dominus ad Mosen in deserto Sinai anno secundo postquam egressi sunt de terra Aegypti mense primo dicens
NUM|9|2|faciant filii Israhel phase in tempore suo
NUM|9|3|quartadecima die mensis huius ad vesperam iuxta omnes caerimonias et iustificationes eius
NUM|9|4|praecepitque Moses filiis Israhel ut facerent phase
NUM|9|5|qui fecerunt tempore suo quartadecima die mensis ad vesperam in monte Sinai iuxta omnia quae mandaverat Dominus Mosi fecerunt filii Israhel
NUM|9|6|ecce autem quidam inmundi super animam hominis qui non poterant facere pascha in die illo accedentes ad Mosen et Aaron
NUM|9|7|dixerunt eis inmundi sumus super animam hominis quare fraudamur ut non valeamus offerre oblationem Domino in tempore suo inter filios Israhel
NUM|9|8|quibus respondit Moses state ut consulam quid praecipiat Dominus de vobis
NUM|9|9|locutusque est Dominus ad Mosen dicens
NUM|9|10|loquere filiis Israhel homo qui fuerit inmundus super anima sive in via procul in gente vestra faciat phase Domino
NUM|9|11|mense secundo quartadecima die mensis ad vesperam cum azymis et lactucis agrestibus comedent illud
NUM|9|12|non relinquent ex eo quippiam usque mane et os eius non confringent omnem ritum phase observabunt
NUM|9|13|si quis autem et mundus est et in itinere non fuit et tamen non fecit phase exterminabitur anima illa de populis suis quia sacrificium Domino non obtulit tempore suo peccatum suum ipse portabit
NUM|9|14|peregrinus quoque et advena si fuerit apud vos faciet phase Domini iuxta caerimonias et iustificationes eius praeceptum idem erit apud vos tam advenae quam indigenae
NUM|9|15|igitur die qua erectum est tabernaculum operuit illud nubes a vespere autem super tentorium erat quasi species ignis usque mane
NUM|9|16|sic fiebat iugiter per diem operiebat illud nubes et per noctem quasi species ignis
NUM|9|17|cumque ablata fuisset nubes quae tabernaculum protegebat tunc proficiscebantur filii Israhel et in loco ubi stetisset nubes ibi castrametabantur
NUM|9|18|ad imperium Domini proficiscebantur et ad imperium illius figebant tabernaculum cunctis diebus quibus stabat nubes super tabernaculum manebant in eodem loco
NUM|9|19|et si evenisset ut multo tempore maneret super illud erant filii Israhel in excubiis Domini et non proficiscebantur
NUM|9|20|quotquot diebus fuisset nubes super tabernaculum ad imperium Domini erigebant tentoria et ad imperium illius deponebant
NUM|9|21|si fuisset nubes a vespere usque mane et statim diluculo tabernaculum reliquisset proficiscebantur et si post diem et noctem recessisset dissipabant tentoria
NUM|9|22|si biduo aut uno mense vel longiori tempore fuisset super tabernaculum manebant filii Israhel in eodem loco et non proficiscebantur statim autem ut recessisset movebant castra
NUM|9|23|per verbum Domini figebant tentoria et per verbum illius proficiscebantur erantque in excubiis Domini iuxta imperium eius per manum Mosi
NUM|10|1|locutus est Dominus ad Mosen dicens
NUM|10|2|fac tibi duas tubas argenteas ductiles quibus convocare possis multitudinem quando movenda sunt castra
NUM|10|3|cumque increpueris tubis congregabitur ad te omnis turba ad ostium foederis tabernaculi
NUM|10|4|si semel clangueris venient ad te principes et capita multitudinis Israhel
NUM|10|5|sin autem prolixior atque concisus clangor increpuerit movebunt castra primi qui sunt ad orientalem plagam
NUM|10|6|in secundo autem sonitu et pari ululatu tubae levabunt tentoria qui habitant ad meridiem et iuxta hunc modum reliqui facient ululantibus tubis in profectione
NUM|10|7|quando autem congregandus est populus simplex tubarum clangor erit et non concise ululabunt
NUM|10|8|filii Aaron sacerdotes clangent tubis eritque hoc legitimum sempiternum in generationibus vestris
NUM|10|9|si exieritis ad bellum de terra vestra contra hostes qui dimicant adversum vos clangetis ululantibus tubis et erit recordatio vestri coram Domino Deo vestro ut eruamini de manibus inimicorum vestrorum
NUM|10|10|si quando habebitis epulum et dies festos et kalendas canetis tubis super holocaustis et pacificis victimis ut sint vobis in recordationem Dei vestri ego Dominus Deus vester
NUM|10|11|anno secundo mense secundo vicesima die mensis elevata est nubes de tabernaculo foederis
NUM|10|12|profectique sunt filii Israhel per turmas suas de deserto Sinai et recubuit nubes in solitudine Pharan
NUM|10|13|moveruntque castra primi iuxta imperium Domini in manu Mosi
NUM|10|14|filii Iuda per turmas suas quorum princeps erat Naasson filius Aminadab
NUM|10|15|in tribu filiorum Isachar fuit princeps Nathanahel filius Suar
NUM|10|16|in tribu Zabulon erat princeps Heliab filius Helon
NUM|10|17|depositumque est tabernaculum quod portantes egressi sunt filii Gerson et Merari
NUM|10|18|profectique sunt et filii Ruben per turmas et ordinem suum quorum princeps erat Helisur filius Sedeur
NUM|10|19|in tribu autem filiorum Symeon princeps fuit Salamihel filius Surisaddai
NUM|10|20|porro in tribu Gad erat princeps Heliasaph filius Duhel
NUM|10|21|profectique sunt et Caathitae portantes sanctuarium tamdiu tabernaculum portabatur donec venirent ad erectionis locum
NUM|10|22|moverunt castra et filii Ephraim per turmas suas in quorum exercitu princeps erat Helisama filius Ammiud
NUM|10|23|in tribu autem filiorum Manasse princeps fuit Gamalihel filius Phadassur
NUM|10|24|et in tribu Beniamin dux Abidan filius Gedeonis
NUM|10|25|novissimi castrorum omnium profecti sunt filii Dan per turmas suas in quorum exercitu princeps fuit Ahiezer filius Amisaddai
NUM|10|26|in tribu autem filiorum Aser erat princeps Phagaihel filius Ochran
NUM|10|27|et in tribu filiorum Nepthalim princeps Achira filius Henan
NUM|10|28|haec sunt castra et profectiones filiorum Israhel per turmas suas quando egrediebantur
NUM|10|29|dixitque Moses Hobab filio Rahuhel Madianiti cognato suo proficiscimur ad locum quem Dominus daturus est nobis veni nobiscum ut benefaciamus tibi quia Dominus bona promisit Israheli
NUM|10|30|cui ille respondit non vadam tecum sed revertar in terram meam in qua natus sum
NUM|10|31|et ille noli inquit nos relinquere tu enim nosti in quibus locis per desertum castra ponere debeamus et eris ductor noster
NUM|10|32|cumque nobiscum veneris quicquid optimum fuerit ex opibus quas nobis traditurus est Dominus dabimus tibi
NUM|10|33|profecti sunt ergo de monte Domini via trium dierum arcaque foederis Domini praecedebat eos per dies tres providens castrorum locum
NUM|10|34|nubes quoque Domini super eos erat per diem cum incederent
NUM|10|35|cumque elevaretur arca dicebat Moses surge Domine et dissipentur inimici tui et fugiant qui oderunt te a facie tua
NUM|10|36|cum autem deponeretur aiebat revertere Domine ad multitudinem exercitus Israhel
NUM|11|1|interea ortum est murmur populi quasi dolentium pro labore contra Dominum quod cum audisset iratus est et accensus in eos ignis Domini devoravit extremam castrorum partem
NUM|11|2|cumque clamasset populus ad Mosen oravit Moses Dominum et absortus est ignis
NUM|11|3|vocavitque nomen loci illius Incensio eo quod succensus fuisset contra eos ignis Domini
NUM|11|4|vulgus quippe promiscuum quod ascenderat cum eis flagravit desiderio sedens et flens iunctis sibi pariter filiis Israhel et ait quis dabit nobis ad vescendum carnes
NUM|11|5|recordamur piscium quos comedebamus in Aegypto gratis in mentem nobis veniunt cucumeres et pepones porrique et cepae et alia
NUM|11|6|anima nostra arida est nihil aliud respiciunt oculi nostri nisi man
NUM|11|7|erat autem man quasi semen coriandri coloris bdellii
NUM|11|8|circuibatque populus et colligens illud frangebat mola sive terebat in mortario coquens in olla et faciens ex eo tortulas saporis quasi panis oleati
NUM|11|9|cumque descenderet nocte super castra ros descendebat pariter et man
NUM|11|10|audivit ergo Moses flentem populum per familias singulos per ostia tentorii sui iratusque est furor Domini valde sed et Mosi intoleranda res visa est
NUM|11|11|et ait ad Dominum cur adflixisti servum tuum quare non invenio gratiam coram te et cur inposuisti pondus universi populi huius super me
NUM|11|12|numquid ego concepi omnem hanc multitudinem vel genui eam ut dicas mihi porta eos in sinu tuo sicut portare solet nutrix infantulum et defer in terram pro qua iurasti patribus eorum
NUM|11|13|unde mihi carnes ut dem tantae multitudini flent contra me dicentes da nobis carnes ut comedamus
NUM|11|14|non possum solus sustinere omnem hunc populum quia gravis mihi est
NUM|11|15|sin aliter tibi videtur obsecro ut interficias me et inveniam gratiam in oculis tuis ne tantis adficiar malis
NUM|11|16|et dixit Dominus ad Mosen congrega mihi septuaginta viros de senibus Israhel quos tu nosti quod senes populi sint ac magistri et duces eos ad ostium tabernaculi foederis faciesque ibi stare tecum
NUM|11|17|ut descendam et loquar tibi et auferam de spiritu tuo tradamque eis ut sustentent tecum onus populi et non tu solus graveris
NUM|11|18|populo quoque dices sanctificamini cras comedetis carnes ego enim audivi vos dicere quis dabit nobis escas carnium bene nobis erat in Aegypto ut det vobis Dominus carnes et comedatis
NUM|11|19|non uno die nec duobus vel quinque aut decem nec viginti quidem
NUM|11|20|sed usque ad mensem dierum donec exeat per nares vestras et vertatur in nausiam eo quod reppuleritis Dominum qui in medio vestri est et fleveritis coram eo dicentes quare egressi sumus ex Aegypto
NUM|11|21|et ait Moses sescenta milia peditum huius populi sunt et tu dicis dabo eis esum carnium mense integro
NUM|11|22|numquid ovium et boum multitudo caedetur ut possit sufficere ad cibum vel omnes pisces maris in unum congregabuntur ut eos satient
NUM|11|23|cui respondit Dominus numquid manus Domini invalida est iam nunc videbis utrum meus sermo opere conpleatur
NUM|11|24|venit igitur Moses et narravit populo verba Domini congregans septuaginta viros de senibus Israhel quos stare fecit circa tabernaculum
NUM|11|25|descenditque Dominus per nubem et locutus est ad eum auferens de spiritu qui erat in Mosen et dans septuaginta viris cumque requievisset in eis spiritus prophetaverunt nec ultra cessarunt
NUM|11|26|remanserant autem in castris duo viri quorum unus vocabatur Heldad et alter Medad super quos requievit spiritus nam et ipsi descripti fuerant et non exierant ad tabernaculum
NUM|11|27|cumque prophetarent in castris cucurrit puer et nuntiavit Mosi dicens Heldad et Medad prophetant in castris
NUM|11|28|statim Iosue filius Nun minister Mosi et electus e pluribus ait domine mi Moses prohibe eos
NUM|11|29|at ille quid inquit aemularis pro me quis tribuat ut omnis populus prophetet et det eis Dominus spiritum suum
NUM|11|30|reversusque est Moses et maiores natu Israhel in castra
NUM|11|31|ventus autem egrediens a Domino arreptas trans mare coturnices detulit et dimisit in castra itinere quantum uno die confici potest ex omni parte castrorum per circuitum volabantque in aere duobus cubitis altitudine super terram
NUM|11|32|surgens ergo populus toto die illo et nocte ac die altero congregavit coturnicum qui parum decem choros et siccaverunt eas per gyrum castrorum
NUM|11|33|adhuc carnes erant in dentibus eorum nec defecerat huiuscemodi cibus et ecce furor Domini concitatus in populum percussit eum plaga magna nimis
NUM|11|34|vocatusque est ille locus sepulchra Concupiscentiae ibi enim sepelierunt populum qui desideraverat egressi autem de sepulchris Concupiscentiae venerunt in Aseroth et manserunt ibi
NUM|11|35|
NUM|12|1|locutaque est Maria et Aaron contra Mosen propter uxorem eius aethiopissam
NUM|12|2|et dixerunt num per solum Mosen locutus est Dominus nonne et nobis similiter est locutus quod cum audisset Dominus
NUM|12|3|erat enim Moses vir mitissimus super omnes homines qui morabantur in terra
NUM|12|4|statim locutus est ad eum et ad Aaron et Mariam egredimini vos tantum tres ad tabernaculum foederis cumque fuissent egressi
NUM|12|5|descendit Dominus in columna nubis et stetit in introitu tabernaculi vocans Aaron et Mariam qui cum issent
NUM|12|6|dixit ad eos audite sermones meos si quis fuerit inter vos propheta Domini in visione apparebo ei vel per somnium loquar ad illum
NUM|12|7|at non talis servus meus Moses qui in omni domo mea fidelissimus est
NUM|12|8|ore enim ad os loquor ei et palam non per enigmata et figuras Dominum videt quare igitur non timuistis detrahere servo meo Mosi
NUM|12|9|iratusque contra eos abiit
NUM|12|10|nubes quoque recessit quae erat super tabernaculum et ecce Maria apparuit candens lepra quasi nix cumque respexisset eam Aaron et vidisset perfusam lepra
NUM|12|11|ait ad Mosen obsecro domine mi ne inponas nobis hoc peccatum quod stulte commisimus
NUM|12|12|ne fiat haec quasi mortua et ut abortivum quod proicitur de vulva matris suae ecce iam medium carnis eius devoratum est lepra
NUM|12|13|clamavitque Moses ad Dominum dicens Deus obsecro sana eam
NUM|12|14|cui respondit Dominus si pater eius spuisset in faciem illius nonne debuerat saltem septem dierum rubore suffundi separetur septem diebus extra castra et postea revocabitur
NUM|12|15|exclusa est itaque Maria extra castra septem diebus et populus non est motus de loco illo donec revocata est Maria
NUM|12|16|
NUM|13|1|profectus est de Aseroth fixis tentoriis in deserto Pharan
NUM|13|2|ibi locutus est Dominus ad Mosen dicens
NUM|13|3|mitte viros qui considerent terram Chanaan quam daturus sum filiis Israhel singulos de singulis tribubus ex principibus
NUM|13|4|fecit Moses quod Dominus imperarat de deserto Pharan mittens principes viros quorum ista sunt nomina
NUM|13|5|de tribu Ruben Semmua filium Zecchur
NUM|13|6|de tribu Symeon Saphat filium Huri
NUM|13|7|de tribu Iuda Chaleb filium Iepphonne
NUM|13|8|de tribu Isachar Igal filium Ioseph
NUM|13|9|de tribu Ephraim Osee filium Nun
NUM|13|10|de tribu Beniamin Phalti filium Raphu
NUM|13|11|de tribu Zabulon Geddihel filium Sodi
NUM|13|12|de tribu Ioseph sceptri Manasse Gaddi filium Susi
NUM|13|13|de tribu Dan Ammihel filium Gemalli
NUM|13|14|de tribu Aser Sthur filium Michahel
NUM|13|15|de tribu Nepthali Naabbi filium Vaphsi
NUM|13|16|de tribu Gad Guhel filium Machi
NUM|13|17|haec sunt nomina virorum quos misit Moses ad considerandam terram vocavitque Osee filium Nun Iosue
NUM|13|18|misit ergo eos Moses ad considerandam terram Chanaan et dixit ad eos ascendite per meridianam plagam cumque veneritis ad montes
NUM|13|19|considerate terram qualis sit et populum qui habitator est eius utrum fortis sit an infirmus pauci numero an plures
NUM|13|20|ipsa terra bona an mala urbes quales muratae an absque muris
NUM|13|21|humus pinguis an sterilis nemorosa an absque arboribus confortamini et adferte nobis de fructibus terrae erat autem tempus quando iam praecoquae uvae vesci possunt
NUM|13|22|cumque ascendissent exploraverunt terram a deserto Sin usque Roob intrantibus Emath
NUM|13|23|ascenderuntque ad meridiem et venerunt in Hebron ubi erant Ahiman et Sisai et Tholmai filii Enach nam Hebron septem annis ante Tanim urbem Aegypti condita est
NUM|13|24|pergentesque usque ad torrentem Botri absciderunt palmitem cum uva sua quem portaverunt in vecte duo viri de malis quoque granatis et de ficis loci illius tulerunt
NUM|13|25|qui appellatus est Neelescol id est torrens Botri eo quod botrum inde portassent filii Israhel
NUM|13|26|reversique exploratores terrae post quadraginta dies omni regione circuita
NUM|13|27|venerunt ad Mosen et Aaron et ad omnem coetum filiorum Israhel in desertum Pharan quod est in Cades locutique eis et omni multitudini ostenderunt fructus terrae
NUM|13|28|et narraverunt dicentes venimus in terram ad quam misisti nos quae re vera fluit lacte et melle ut ex his fructibus cognosci potest
NUM|13|29|sed cultores fortissimos habet et urbes grandes atque muratas stirpem Enach vidimus ibi
NUM|13|30|Amalech habitat in meridie Hettheus et Iebuseus et Amorreus in montanis Chananeus vero moratur iuxta mare et circa fluenta Iordanis
NUM|13|31|inter haec Chaleb conpescens murmur populi qui oriebatur contra Mosen ait ascendamus et possideamus terram quoniam poterimus obtinere eam
NUM|13|32|alii vero qui fuerant cum eo dicebant nequaquam ad hunc populum valemus ascendere quia fortior nobis est
NUM|13|33|detraxeruntque terrae quam inspexerant apud filios Israhel dicentes terram quam lustravimus devorat habitatores suos populum quem aspeximus procerae staturae est
NUM|13|34|ibi vidimus monstra quaedam filiorum Enach de genere giganteo quibus conparati quasi lucustae videbamur
NUM|14|1|igitur vociferans omnis turba flevit nocte illa
NUM|14|2|et murmurati sunt contra Mosen et Aaron cuncti filii Israhel dicentes
NUM|14|3|utinam mortui essemus in Aegypto et non in hac vasta solitudine utinam pereamus et non inducat nos Dominus in terram istam ne cadamus gladio et uxores ac liberi nostri ducantur captivi nonne melius est reverti in Aegyptum
NUM|14|4|dixeruntque alter ad alterum constituamus nobis ducem et revertamur in Aegyptum
NUM|14|5|quo audito Moses et Aaron ceciderunt proni in terram coram omni multitudine filiorum Israhel
NUM|14|6|at vero Iosue filius Nun et Chaleb filius Iepphonne qui et ipsi lustraverant terram sciderunt vestimenta sua
NUM|14|7|et ad omnem multitudinem filiorum Israhel locuti sunt terram quam circuivimus valde bona est
NUM|14|8|si propitius fuerit Dominus inducet nos in eam et tradet humum lacte et melle manantem
NUM|14|9|nolite rebelles esse contra Dominum neque timeatis populum terrae huius quia sicut panem ita eos possumus devorare recessit ab illis omne praesidium Dominus nobiscum est nolite metuere
NUM|14|10|cumque clamaret omnis multitudo et lapidibus eos vellet opprimere apparuit gloria Domini super tectum foederis cunctis filiis Israhel
NUM|14|11|et dixit Dominus ad Mosen usquequo detrahet mihi populus iste quousque non credent mihi in omnibus signis quae feci coram eis
NUM|14|12|feriam igitur eos pestilentia atque consumam te autem faciam principem super gentem magnam et fortiorem quam haec est
NUM|14|13|et ait Moses ad Dominum ut audiant Aegyptii de quorum medio eduxisti populum istum
NUM|14|14|et habitatores terrae huius qui audierunt quod tu Domine in populo isto sis et facie videaris ad faciem et nubes tua protegat illos et in columna nubis praecedas eos per diem et in columna ignis per noctem
NUM|14|15|quod occideris tantam multitudinem quasi unum hominem et dicant
NUM|14|16|non poterat introducere populum in terram pro qua iuraverat idcirco occidit eos in solitudine
NUM|14|17|magnificetur ergo fortitudo Domini sicut iurasti dicens
NUM|14|18|Dominus patiens et multae misericordiae auferens iniquitatem et scelera nullumque innoxium derelinquens qui visitas peccata patrum in filios in tertiam et quartam generationem
NUM|14|19|dimitte obsecro peccatum populi tui huius secundum magnitudinem misericordiae tuae sicut propitius fuisti egredientibus de Aegypto usque ad locum istum
NUM|14|20|dixitque Dominus dimisi iuxta verbum tuum
NUM|14|21|vivo ego et implebitur gloria Domini universa terra
NUM|14|22|attamen omnes homines qui viderunt maiestatem meam et signa quae feci in Aegypto et in solitudine et temptaverunt me iam per decem vices nec oboedierunt voci meae
NUM|14|23|non videbunt terram pro qua iuravi patribus eorum nec quisquam ex illis qui detraxit mihi intuebitur eam
NUM|14|24|servum meum Chaleb qui plenus alio spiritu secutus est me inducam in terram hanc quam circuivit et semen eius possidebit eam
NUM|14|25|quoniam Amalechites et Chananeus habitant in vallibus cras movete castra et revertimini in solitudinem per viam maris Rubri
NUM|14|26|locutusque est Dominus ad Mosen et Aaron dicens
NUM|14|27|usquequo multitudo haec pessima murmurat contra me querellas filiorum Israhel audivi
NUM|14|28|dic ergo eis vivo ego ait Dominus sicut locuti estis audiente me sic faciam vobis
NUM|14|29|in solitudine hac iacebunt cadavera vestra omnes qui numerati estis a viginti annis et supra et murmurastis contra me
NUM|14|30|non intrabitis terram super quam levavi manum meam ut habitare vos facerem praeter Chaleb filium Iepphonne et Iosue filium Nun
NUM|14|31|parvulos autem vestros de quibus dixistis quod praedae hostibus forent introducam ut videant terram quae vobis displicuit
NUM|14|32|vestra cadavera iacebunt in solitudine
NUM|14|33|filii vestri erunt vagi in deserto annis quadraginta et portabunt fornicationem vestram donec consumantur cadavera patrum in deserto
NUM|14|34|iuxta numerum quadraginta dierum quibus considerastis terram annus pro die inputabitur et quadraginta annis recipietis iniquitates vestras et scietis ultionem meam
NUM|14|35|quoniam sicut locutus sum ita faciam omni multitudini huic pessimae quae consurrexit adversum me in solitudine hac deficiet et morietur
NUM|14|36|igitur omnes viri quos miserat Moses ad contemplandam terram et qui reversi murmurare fecerant contra eum omnem multitudinem detrahentes terrae quod esset mala
NUM|14|37|mortui sunt atque percussi in conspectu Domini
NUM|14|38|Iosue autem filius Nun et Chaleb filius Iepphonne vixerunt ex omnibus qui perrexerant ad considerandam terram
NUM|14|39|locutusque est Moses universa verba haec ad omnes filios Israhel et luxit populus nimis
NUM|14|40|et ecce mane primo surgentes ascenderunt verticem montis atque dixerunt parati sumus ascendere ad locum de quo Dominus locutus est quia peccavimus
NUM|14|41|quibus Moses cur inquit transgredimini verbum Domini quod vobis non cedet in prosperum
NUM|14|42|nolite ascendere non enim est Dominus vobiscum ne corruatis coram inimicis vestris
NUM|14|43|Amalechites et Chananeus ante vos sunt quorum gladio corruetis eo quod nolueritis adquiescere Domino nec erit Dominus vobiscum
NUM|14|44|at illi contenebrati ascenderunt in verticem montis arca autem testamenti Domini et Moses non recesserunt de castris
NUM|14|45|descenditque Amalechites et Chananeus qui habitabant in monte et percutiens eos atque concidens persecutus est usque Horma
NUM|15|1|locutus est Dominus ad Mosen dicens
NUM|15|2|loquere ad filios Israhel et dices ad eos cum ingressi fueritis terram habitationis vestrae quam ego dabo vobis
NUM|15|3|et feceritis oblationem Domino in holocaustum aut victimam vota solventes vel sponte offerentes munera aut in sollemnitatibus vestris adolentes odorem suavitatis Domino de bubus sive de ovibus
NUM|15|4|offeret quicumque immolaverit victimam sacrificium similae decimam partem oephi conspersae oleo quod mensuram habebit quartam partem hin
NUM|15|5|et vinum ad liba fundenda eiusdem mensurae dabit in holocausto sive in victima per agnos singulos
NUM|15|6|et arietis erit sacrificium similae duarum decimarum quae conspersa sit oleo tertiae partis hin
NUM|15|7|et vinum ad libamentum tertiae partis eiusdem mensurae offeret in odorem suavitatis Domino
NUM|15|8|quando vero de bubus feceris holocaustum aut hostiam ut impleas votum vel pacificas victimas
NUM|15|9|dabis per singulos boves similae tres decimas conspersae oleo quod habeat medium mensurae hin
NUM|15|10|et vinum ad liba fundenda eiusdem mensurae in oblationem suavissimi odoris Domino
NUM|15|11|sic facietis
NUM|15|12|per singulos boves et arietes et agnos et hedos
NUM|15|13|tam indigenae quam peregrini
NUM|15|14|eodem ritu offerent sacrificia
NUM|15|15|unum praeceptum erit atque iudicium tam vobis quam advenis terrae
NUM|15|16|locutus est Dominus ad Mosen dicens
NUM|15|17|loquere filiis Israhel et dices ad eos
NUM|15|18|cum veneritis in terram quam dabo vobis
NUM|15|19|et comederitis de panibus regionis illius separabitis primitias Domino
NUM|15|20|de cibis vestris sicut de areis primitias separatis
NUM|15|21|ita et de pulmentis dabitis primitiva Domino
NUM|15|22|quod si per ignorantiam praeterieritis quicquam horum quae locutus est Dominus ad Mosen
NUM|15|23|et mandavit per eum ad vos a die qua coepit iubere et ultra
NUM|15|24|oblitaque fuerit facere multitudo offeret vitulum de armento holocaustum in odorem suavissimum Domino et sacrificium eius ac liba ut caerimoniae postulant hircumque pro peccato
NUM|15|25|et rogabit sacerdos pro omni multitudine filiorum Israhel et dimittetur eis quoniam non sponte peccaverunt nihilominus offerentes incensum Domino pro se et pro peccato atque errore suo
NUM|15|26|et dimittetur universae plebi filiorum Israhel et advenis qui peregrinantur inter vos quoniam culpa est omnis populi per ignorantiam
NUM|15|27|quod si anima una nesciens peccaverit offeret capram anniculam pro peccato suo
NUM|15|28|et deprecabitur pro ea sacerdos quod inscia peccaverit coram Domino inpetrabitque ei veniam et dimittetur illi
NUM|15|29|tam indigenis quam advenis una lex erit omnium qui peccaverint ignorantes
NUM|15|30|anima vero quae per superbiam aliquid commiserit sive civis sit ille sive peregrinus quoniam adversum Dominum rebellis fuit peribit de populo suo
NUM|15|31|verbum enim Domini contempsit et praeceptum illius fecit irritum idcirco delebitur et portabit iniquitatem suam
NUM|15|32|factum est autem cum essent filii Israhel in solitudine et invenissent hominem colligentem ligna in die sabbati
NUM|15|33|obtulerunt eum Mosi et Aaron et universae multitudini
NUM|15|34|qui recluserunt eum in carcerem nescientes quid super eo facere deberent
NUM|15|35|dixitque Dominus ad Mosen morte moriatur homo iste obruat eum lapidibus omnis turba extra castra
NUM|15|36|cumque eduxissent eum foras obruerunt lapidibus et mortuus est sicut praeceperat Dominus
NUM|15|37|dixit quoque Dominus ad Mosen
NUM|15|38|loquere filiis Israhel et dices ad eos ut faciant sibi fimbrias per angulos palliorum ponentes in eis vittas hyacinthinas
NUM|15|39|quas cum viderint recordentur omnium mandatorum Domini nec sequantur cogitationes suas et oculos per res varias fornicantes
NUM|15|40|sed magis memores praeceptorum Domini faciant ea sintque sancti Deo suo
NUM|15|41|ego Dominus Deus vester qui eduxi vos de terra Aegypti ut essem vester Deus
NUM|16|1|ecce autem Core filius Isaar filii Caath filii Levi et Dathan atque Abiram filii Heliab Hon quoque filius Pheleth de filiis Ruben
NUM|16|2|surrexerunt contra Mosen aliique filiorum Israhel ducenti quinquaginta viri proceres synagogae et qui tempore concilii per nomina vocabantur
NUM|16|3|cumque stetissent adversum Mosen et Aaron dixerunt sufficiat vobis quia omnis multitudo sanctorum est et in ipsis est Dominus cur elevamini super populum Domini
NUM|16|4|quod cum audisset Moses cecidit pronus in faciem
NUM|16|5|locutusque ad Core et ad omnem multitudinem mane inquit notum faciet Dominus qui ad se pertineant et sanctos adplicabit sibi et quos elegerit adpropinquabunt ei
NUM|16|6|hoc igitur facite tollat unusquisque turibula sua tu Core et omne concilium tuum
NUM|16|7|et hausto cras igne ponite desuper thymiama coram Domino et quemcumque elegerit ipse erit sanctus multum erigimini filii Levi
NUM|16|8|dixitque rursum ad Core audite filii Levi
NUM|16|9|num parum vobis est quod separavit vos Deus Israhel ab omni populo et iunxit sibi ut serviretis ei in cultu tabernaculi et staretis coram frequentia populi et ministraretis ei
NUM|16|10|idcirco ad se fecit accedere te et omnes fratres tuos filios Levi ut vobis etiam sacerdotium vindicetis
NUM|16|11|et omnis globus tuus stet contra Dominum quid est enim Aaron ut murmuretis contra eum
NUM|16|12|misit ergo Moses ut vocaret Dathan et Abiram filios Heliab qui responderunt non venimus
NUM|16|13|numquid parum est tibi quod eduxisti nos de terra quae lacte et melle manabat ut occideres in deserto nisi et dominatus fueris nostri
NUM|16|14|re vera induxisti nos in terram quae fluit rivis lactis et mellis et dedisti nobis possessiones agrorum et vinearum an et oculos nostros vis eruere non venimus
NUM|16|15|iratusque Moses valde ait ad Dominum ne respicias sacrificia eorum tu scis quod ne asellum quidem umquam acceperim ab eis nec adflixerim quempiam eorum
NUM|16|16|dixitque ad Core tu et omnis congregatio tua state seorsum coram Domino et Aaron die crastino separatim
NUM|16|17|tollite singuli turibula vestra et ponite super ea incensum offerentes Domino ducenta quinquaginta turibula Aaron quoque teneat turibulum suum
NUM|16|18|quod cum fecissent stantibus Mosen et Aaron
NUM|16|19|et coacervassent adversum eos omnem multitudinem ad ostium tabernaculi apparuit cunctis gloria Domini
NUM|16|20|locutusque Dominus ad Mosen et Aaron ait
NUM|16|21|separamini de medio congregationis huius ut eos repente disperdam
NUM|16|22|qui ceciderunt proni in faciem atque dixerunt fortissime Deus spirituum universae carnis num uno peccante contra omnes tua ira desaeviet
NUM|16|23|et ait Dominus ad Mosen
NUM|16|24|praecipe universo populo ut separetur a tabernaculis Core et Dathan et Abiram
NUM|16|25|surrexitque Moses et abiit ad Dathan et Abiram et sequentibus eum senioribus Israhel
NUM|16|26|dixit ad turbam recedite a tabernaculis hominum impiorum et nolite tangere quae ad eos pertinent ne involvamini in peccatis eorum
NUM|16|27|cumque recessissent a tentoriis eorum per circuitum Dathan et Abiram egressi stabant in introitu papilionum suorum cum uxoribus et liberis omnique frequentia
NUM|16|28|et ait Moses in hoc scietis quod Dominus miserit me ut facerem universa quae cernitis et non ex proprio ea corde protulerim
NUM|16|29|si consueta hominum morte interierint et visitaverit eos plaga qua et ceteri visitari solent non misit me Dominus
NUM|16|30|sin autem novam rem fecerit Dominus ut aperiens terra os suum degluttiat eos et omnia quae ad illos pertinent descenderintque viventes in infernum scietis quod blasphemaverint Dominum
NUM|16|31|confestim igitur ut cessavit loqui disrupta est terra sub pedibus eorum
NUM|16|32|et aperiens os suum devoravit illos cum tabernaculis suis et universa substantia
NUM|16|33|descenderuntque vivi in infernum operti humo et perierunt de medio multitudinis
NUM|16|34|at vero omnis Israhel qui stabat per gyrum fugit ad clamorem pereuntium dicens ne forte et nos terra degluttiat
NUM|16|35|sed et ignis egressus a Domino interfecit ducentos quinquaginta viros qui offerebant incensum
NUM|16|36|locutusque est Dominus ad Mosen dicens
NUM|16|37|praecipe Eleazaro filio Aaron sacerdotis ut tollat turibula quae iacent in incendio et ignem huc illucque dispergat quoniam sanctificata sunt
NUM|16|38|in mortibus peccatorum producatque ea in lamminas et adfigat altari eo quod oblatum sit in eis incensum Domino et sanctificata sint ut cernant ea pro signo et monumento filii Israhel
NUM|16|39|tulit ergo Eleazar sacerdos turibula aenea in quibus obtulerant hii quos incendium devoravit et produxit ea in lamminas adfigens altari
NUM|16|40|ut haberent postea filii Israhel quibus commonerentur ne quis accedat alienigena et qui non est de semine Aaron ad offerendum incensum Domino ne patiatur sicut passus est Core et omnis congregatio eius loquente Domino ad Mosen
NUM|16|41|murmuravit autem omnis multitudo filiorum Israhel sequenti die contra Mosen et Aaron dicens vos interfecistis populum Domini
NUM|16|42|cumque oreretur seditio et tumultus incresceret
NUM|16|43|Moses et Aaron fugerunt ad tabernaculum foederis quod postquam ingressi sunt operuit nubes et apparuit gloria Domini
NUM|16|44|dixitque Dominus ad Mosen
NUM|16|45|recedite de medio huius multitudinis etiam nunc delebo eos cumque iacerent in terra
NUM|16|46|dixit Moses ad Aaron tolle turibulum et hausto igne de altari mitte incensum desuper pergens cito ad populum ut roges pro eis iam enim egressa est ira a Domino et plaga desaevit
NUM|16|47|quod cum fecisset Aaron et cucurrisset ad mediam multitudinem quam iam vastabat incendium obtulit thymiama
NUM|16|48|et stans inter mortuos ac viventes pro populo deprecatus est et plaga cessavit
NUM|16|49|fuerunt autem qui percussi sunt quattuordecim milia hominum et septingenti absque his qui perierant in seditione Core
NUM|16|50|reversusque est Aaron ad Mosen ad ostium tabernaculi foederis postquam quievit interitus
NUM|17|1|et locutus est Dominus ad Mosen dicens
NUM|17|2|loquere ad filios Israhel et accipe ab eis virgas singulas per cognationes suas a cunctis principibus tribuum virgas duodecim et uniuscuiusque nomen superscribes virgae suae
NUM|17|3|nomen autem Aaron erit in tribu Levi et una virga cunctas eorum familias continebit
NUM|17|4|ponesque eas in tabernaculo foederis coram testimonio ubi loquar ad te
NUM|17|5|quem ex his elegero germinabit virga eius et cohibebo a me querimonias filiorum Israhel quibus contra vos murmurant
NUM|17|6|locutusque est Moses ad filios Israhel et dederunt ei omnes principes virgas per singulas tribus fueruntque virgae duodecim absque virga Aaron
NUM|17|7|quas cum posuisset Moses coram Domino in tabernaculo testimonii
NUM|17|8|sequenti die regressus invenit germinasse virgam Aaron in domo Levi et turgentibus gemmis eruperant flores qui foliis dilatatis in amigdalas deformati sunt
NUM|17|9|protulit ergo Moses omnes virgas de conspectu Domini ad cunctos filios Israhel videruntque et receperunt singuli virgas suas
NUM|17|10|dixitque Dominus ad Mosen refer virgam Aaron in tabernaculum testimonii ut servetur ibi in signum rebellium filiorum et quiescant querellae eorum a me ne moriantur
NUM|17|11|fecitque Moses sicut praeceperat Dominus
NUM|17|12|dixerunt autem filii Israhel ad Mosen ecce consumpti sumus omnes perivimus
NUM|17|13|quicumque accedit ad tabernaculum Domini moritur num usque ad internicionem cuncti delendi sumus
NUM|18|1|dixitque Dominus ad Aaron tu et filii tui et domus patris tui tecum portabitis iniquitatem sanctuarii et tu et filii tui simul sustinebitis peccata sacerdotii vestri
NUM|18|2|sed et fratres tuos de tribu Levi et sceptro patris tui sume tecum praestoque sint et ministrent tibi tu autem et filii tui ministrabitis in tabernaculo testimonii
NUM|18|3|excubabuntque Levitae ad praecepta tua et ad cuncta opera tabernaculi ita dumtaxat ut ad vasa sanctuarii et altare non accedant ne et illi moriantur et vos pereatis simul
NUM|18|4|sint autem tecum et excubent in custodiis tabernaculi et in omnibus caerimoniis eius alienigena non miscebitur vobis
NUM|18|5|excubate in custodia sanctuarii et in ministerio altaris ne oriatur indignatio super filios Israhel
NUM|18|6|ego dedi vobis fratres vestros Levitas de medio filiorum Israhel et tradidi donum Domino ut serviant in ministeriis tabernaculi eius
NUM|18|7|tu autem et filii tui custodite sacerdotium vestrum et omnia quae ad cultum altaris pertinent et intra velum sunt per sacerdotes administrabuntur si quis externus accesserit occidetur
NUM|18|8|locutus est Dominus ad Aaron ecce dedi tibi custodiam primitiarum mearum omnia quae sanctificantur a filiis Israhel tibi tradidi et filiis tuis pro officio sacerdotali legitima sempiterna
NUM|18|9|haec ergo accipies de his quae sanctificantur et oblata sunt Domino omnis oblatio et sacrificium et quicquid pro peccato atque delicto redditur mihi et cedet in sancta sanctorum tuum erit et filiorum tuorum
NUM|18|10|in sanctuario comedes illud mares tantum edent ex eo quia consecratum est tibi
NUM|18|11|primitias autem quas voverint et obtulerint filii Israhel tibi dedi et filiis ac filiabus tuis iure perpetuo qui mundus est in domo tua vescetur eis
NUM|18|12|omnem medullam olei et vini ac frumenti quicquid offerunt primitiarum Domino tibi dedi
NUM|18|13|universa frugum initia quas gignit humus et Domino deportantur cedent in usus tuos qui mundus est in domo tua vescetur eis
NUM|18|14|omne quod ex voto reddiderint filii Israhel tuum erit
NUM|18|15|quicquid primum erumpet e vulva cunctae carnis quam offerunt Domino sive ex hominibus sive de pecoribus fuerit tui iuris erit ita dumtaxat ut pro hominis primogenito pretium accipias et omne animal quod inmundum est redimi facias
NUM|18|16|cuius redemptio erit post unum mensem siclis argenti quinque pondere sanctuarii siclus viginti obolos habet
NUM|18|17|primogenitum autem bovis et ovis et caprae non facies redimi quia sanctificata sunt Domino sanguinem tantum eorum fundes super altare et adipes adolebis in suavissimum odorem Domino
NUM|18|18|carnes vero in usum tuum cedent sicut pectusculum consecratum et armus dexter tua erunt
NUM|18|19|omnes primitias sanctuarii quas offerunt filii Israhel Domino tibi dedi et filiis ac filiabus tuis iure perpetuo pactum salis est sempiternum coram Domino tibi ac filiis tuis
NUM|18|20|dixitque Dominus ad Aaron in terra eorum nihil possidebitis nec habebitis partem inter eos ego pars et hereditas tua in medio filiorum Israhel
NUM|18|21|filiis autem Levi dedi omnes decimas Israhelis in possessionem pro ministerio quo serviunt mihi in tabernaculo foederis
NUM|18|22|ut non accedant ultra filii Israhel ad tabernaculum nec committant peccatum mortiferum
NUM|18|23|solis filiis Levi mihi in tabernaculo servientibus et portantibus peccata populi legitimum sempiternum erit in generationibus vestris nihil aliud possidebunt
NUM|18|24|decimarum oblatione contenti quas in usus eorum et necessaria separavi
NUM|18|25|locutusque est Dominus ad Mosen dicens
NUM|18|26|praecipe Levitis atque denuntia cum acceperitis a filiis Israhel decimas quas dedi vobis primitias earum offerte Domino id est decimam partem decimae
NUM|18|27|ut reputetur vobis in oblationem primitivorum tam de areis quam de torcularibus
NUM|18|28|et universis quorum accipitis primitias offerte Domino et date Aaron sacerdoti
NUM|18|29|omnia quae offertis ex decimis et in donaria Domini separatis optima et electa erunt
NUM|18|30|dicesque ad eos si praeclara et meliora quaeque obtuleritis ex decimis reputabitur vobis quasi de area et torculari dederitis primitias
NUM|18|31|et comedetis eas in omnibus locis vestris tam vos quam familiae vestrae quia pretium est pro ministerio quo servitis in tabernaculo testimonii
NUM|18|32|et non peccabitis super hoc egregia vobis et pinguia reservantes ne polluatis oblationes filiorum Israhel et moriamini
NUM|19|1|locutusque est Dominus ad Mosen et Aaron dicens
NUM|19|2|ista est religio victimae quam constituit Dominus praecipe filiis Israhel ut adducant ad te vaccam rufam aetatis integrae in qua nulla sit macula nec portaverit iugum
NUM|19|3|tradetisque eam Eleazaro sacerdoti qui eductam extra castra immolabit in conspectu omnium
NUM|19|4|et tinguens digitum in sanguine eius asperget contra fores tabernaculi septem vicibus
NUM|19|5|conburetque eam cunctis videntibus tam pelle et carnibus eius quam sanguine et fimo flammae traditis
NUM|19|6|lignum quoque cedrinum et hysopum coccumque bis tinctum sacerdos mittet in flammam quae vaccam vorat
NUM|19|7|et tunc demum lotis vestibus et corpore suo ingredietur in castra commaculatusque erit usque ad vesperam
NUM|19|8|sed et ille qui conbuserit eam lavabit vestimenta sua et corpus et inmundus erit usque ad vesperam
NUM|19|9|colliget autem vir mundus cineres vaccae et effundet eos extra castra in loco purissimo ut sint multitudini filiorum Israhel in custodiam et in aquam aspersionis quia pro peccato vacca conbusta est
NUM|19|10|cumque laverit qui vaccae portaverat cineres vestimenta sua inmundus erit usque ad vesperum habebunt hoc filii Israhel et advenae qui habitant inter eos sanctum iure perpetuo
NUM|19|11|qui tetigerit cadaver hominis et propter hoc septem diebus fuerit inmundus
NUM|19|12|aspergetur ex hac aqua die tertio et septimo et sic mundabitur si die tertio aspersus non fuerit septimo non poterit emundari
NUM|19|13|omnis qui tetigerit humanae animae morticinum et aspersus hac commixtione non fuerit polluet tabernaculum Domini et peribit ex Israhel quia aqua expiationis non est aspersus inmundus erit et manebit spurcitia eius super eum
NUM|19|14|ista est lex hominis qui moritur in tabernaculo omnes qui ingrediuntur tentorium illius et universa vasa quae ibi sunt polluta erunt septem diebus
NUM|19|15|vas quod non habuerit operculum nec ligaturam desuper inmundum erit
NUM|19|16|si quis in agro tetigerit cadaver occisi hominis aut per se mortui sive os illius vel sepulchrum inmundus erit septem diebus
NUM|19|17|tollent de cineribus conbustionis atque peccati et mittent aquas vivas super eos in vas
NUM|19|18|in quibus cum homo mundus tinxerit hysopum asperget eo omne tentorium et cunctam supellectilem et homines huiuscemodi contagione pollutos
NUM|19|19|atque hoc modo mundus lustrabit inmundum tertio et septimo die expiatusque die septimo lavabit et se et vestimenta sua et mundus erit ad vesperam
NUM|19|20|si quis hoc ritu non fuerit expiatus peribit anima illius de medio ecclesiae quia sanctuarium Domini polluit et non est aqua lustrationis aspersus
NUM|19|21|erit hoc praeceptum legitimum sempiternum ipse quoque qui aspergit aquas lavabit vestimenta sua omnis qui tetigerit aquas expiationis inmundus erit usque ad vesperam
NUM|19|22|quicquid tetigerit inmundus inmundum faciet et anima quae horum quippiam tetigerit inmunda erit usque ad vesperum
NUM|20|1|veneruntque filii Israhel et omnis multitudo in desertum Sin mense primo et mansit populus in Cades mortuaque est ibi Maria et sepulta in eodem loco
NUM|20|2|cumque indigeret aqua populus coierunt adversum Mosen et Aaron
NUM|20|3|et versi in seditionem dixerunt utinam perissemus inter fratres nostros coram Domino
NUM|20|4|cur eduxistis ecclesiam Domini in solitudinem ut et nos et nostra iumenta moriantur
NUM|20|5|quare nos fecistis ascendere de Aegypto et adduxistis in locum istum pessimum qui seri non potest qui nec ficum gignit nec vineas nec mala granata insuper et aquam non habet ad bibendum
NUM|20|6|ingressusque Moses et Aaron dimissa multitudine tabernaculum foederis corruerunt proni in terram et apparuit gloria Domini super eos
NUM|20|7|locutusque est Dominus ad Mosen dicens
NUM|20|8|tolle virgam et congrega populum tu et Aaron frater tuus et loquimini ad petram coram eis et illa dabit aquas cumque eduxeris aquam de petra bibet omnis multitudo et iumenta eius
NUM|20|9|tulit igitur Moses virgam quae erat in conspectu Domini sicut praeceperat ei
NUM|20|10|congregata multitudine ante petram dixitque eis audite rebelles et increduli num de petra hac vobis aquam poterimus eicere
NUM|20|11|cumque elevasset Moses manum percutiens virga bis silicem egressae sunt aquae largissimae ita ut et populus biberet et iumenta
NUM|20|12|dixitque Dominus ad Mosen et Aaron quia non credidistis mihi ut sanctificaretis me coram filiis Israhel non introducetis hos populos in terram quam dabo eis
NUM|20|13|haec est aqua Contradictionis ubi iurgati sunt filii Israhel contra Dominum et sanctificatus est in eis
NUM|20|14|misit interea nuntios Moses de Cades ad regem Edom qui dicerent haec mandat frater tuus Israhel nosti omnem laborem qui adprehendit nos
NUM|20|15|quomodo descenderint patres nostri in Aegyptum et habitaverimus ibi multo tempore adflixerintque nos Aegyptii et patres nostros
NUM|20|16|et quomodo clamaverimus ad Dominum et exaudierit nos miseritque angelum qui eduxerit nos de Aegypto ecce in urbe Cades quae est in extremis finibus tuis positi
NUM|20|17|obsecramus ut nobis transire liceat per terram tuam non ibimus per agros nec per vineas non bibemus aquas de puteis tuis sed gradiemur via publica nec ad dextram nec ad sinistram declinantes donec transeamus terminos tuos
NUM|20|18|cui respondit Edom non transibis per me alioquin armatus occurram tibi
NUM|20|19|dixeruntque filii Israhel per tritam gradiemur viam et si biberimus aquas tuas nos et pecora nostra dabimus quod iustum est nulla erit in pretio difficultas tantum velociter transeamus
NUM|20|20|at ille respondit non transibis statimque egressus est obvius cum infinita multitudine et manu forti
NUM|20|21|nec voluit adquiescere deprecanti ut concederet transitum per fines suos quam ob rem devertit ab eo Israhel
NUM|20|22|cumque castra movissent de Cades venerunt in montem Or qui est in finibus terrae Edom
NUM|20|23|ubi locutus est Dominus ad Mosen
NUM|20|24|pergat inquit Aaron ad populos suos non enim intrabit terram quam dedi filiis Israhel eo quod incredulus fuerit ori meo ad aquas Contradictionis
NUM|20|25|tolle Aaron et filium eius cum eo et duces eos in montem Or
NUM|20|26|cumque nudaveris patrem veste sua indues ea Eleazarum filium eius et Aaron colligetur et morietur ibi
NUM|20|27|fecit Moses ut praeceperat Dominus et ascenderunt in montem Or coram omni multitudine
NUM|20|28|cumque Aaron spoliasset vestibus suis induit eis Eleazarum filium eius
NUM|20|29|illo mortuo in montis supercilio descendit cum Eleazaro
NUM|20|30|omnis autem multitudo videns occubuisse Aaron flevit super eo triginta diebus per cunctas familias suas
NUM|21|1|quod cum audisset Chananeus rex Arad qui habitabat ad meridiem venisse scilicet Israhel per exploratorum viam pugnavit contra illum et victor existens duxit ex eo praedam
NUM|21|2|at Israhel voto se Domino obligans ait si tradideris populum istum in manu mea delebo urbes eius
NUM|21|3|exaudivitque Dominus preces Israhel et tradidit Chananeum quem ille interfecit subversis urbibus eius et vocavit nomen loci illius Horma id est anathema
NUM|21|4|profecti sunt autem et de monte Or per viam quae ducit ad mare Rubrum ut circumirent terram Edom et taedere coepit populum itineris ac laboris
NUM|21|5|locutusque contra Deum et Mosen ait cur eduxisti nos de Aegypto ut moreremur in solitudine deest panis non sunt aquae anima nostra iam nausiat super cibo isto levissimo
NUM|21|6|quam ob rem misit Dominus in populum ignitos serpentes ad quorum plagas et mortes plurimorum
NUM|21|7|venerunt ad Mosen atque dixerunt peccavimus quia locuti sumus contra Dominum et te ora ut tollat a nobis serpentes oravit Moses pro populo
NUM|21|8|et locutus est Dominus ad eum fac serpentem et pone eum pro signo qui percussus aspexerit eum vivet
NUM|21|9|fecit ergo Moses serpentem aeneum et posuit pro signo quem cum percussi aspicerent sanabantur
NUM|21|10|profectique filii Israhel castrametati sunt in Oboth
NUM|21|11|unde egressi fixere tentoria in Hieabarim in solitudine quae respicit Moab contra orientalem plagam
NUM|21|12|et inde moventes venerunt ad torrentem Zared
NUM|21|13|quem relinquentes castrametati sunt contra Arnon quae est in deserto et prominet in finibus Amorrei siquidem Arnon terminus est Moab dividens Moabitas et Amorreos
NUM|21|14|unde dicitur in libro bellorum Domini sicut fecit in mari Rubro sic faciet in torrentibus Arnon
NUM|21|15|scopuli torrentium inclinati sunt ut requiescerent in Ar et recumberent in finibus Moabitarum
NUM|21|16|ex eo loco apparuit puteus super quo locutus est Dominus ad Mosen congrega populum et dabo ei aquam
NUM|21|17|tunc cecinit Israhel carmen istud ascendat puteus concinebant
NUM|21|18|puteus quem foderunt principes et paraverunt duces multitudinis in datore legis et in baculis suis de solitudine Matthana
NUM|21|19|de Matthana Nahalihel de Nahalihel in Bamoth
NUM|21|20|de Bamoth vallis est in regione Moab in vertice Phasga et quod respicit contra desertum
NUM|21|21|misit autem Israhel nuntios ad Seon regem Amorreorum dicens
NUM|21|22|obsecro ut transire mihi liceat per terram tuam non declinabimus in agros et vineas non bibemus aquas ex puteis via regia gradiemur donec transeamus terminos tuos
NUM|21|23|qui concedere noluit ut transiret Israhel per fines suos quin potius exercitu congregato egressus est obviam in desertum et venit in Iasa pugnavitque contra eum
NUM|21|24|a quo percussus est in ore gladii et possessa est terra eius ab Arnon usque Iebboc et filios Ammon quia forti praesidio tenebantur termini Ammanitarum
NUM|21|25|tulit ergo Israhel omnes civitates eius et habitavit in urbibus Amorrei in Esebon scilicet et viculis eius
NUM|21|26|urbs Esebon fuit regis Seon Amorrei qui pugnavit contra regem Moab et tulit omnem terram quae dicionis illius fuerat usque Arnon
NUM|21|27|idcirco dicitur in proverbio venite in Esebon aedificetur et construatur civitas Seon
NUM|21|28|ignis egressus est de Esebon flamma de oppido Seon et devoravit Ar Moabitarum et habitatores excelsorum Arnon
NUM|21|29|vae tibi Moab peristi popule Chamos dedit filios eius in fugam et filias in captivitatem regi Amorreorum Seon
NUM|21|30|iugum ipsorum disperiit ab Esebon usque Dibon lassi pervenerunt in Nophe et usque Medaba
NUM|21|31|habitavit itaque Israhel in terra Amorrei
NUM|21|32|misitque Moses qui explorarent Iazer cuius ceperunt viculos et possederunt habitatores
NUM|21|33|verteruntque se et ascenderunt per viam Basan et occurrit eis Og rex Basan cum omni populo suo pugnaturus in Edrai
NUM|21|34|dixitque Dominus ad Mosen ne timeas eum quia in manu tua tradidi illum et omnem populum ac terram eius faciesque illi sicut fecisti Seon regi Amorreorum habitatori Esebon
NUM|21|35|percusserunt igitur et hunc cum filiis suis universumque populum eius usque ad internicionem et possederunt terram illius
NUM|22|1|profectique castrametati sunt in campestribus Moab ubi trans Iordanem Hierichus sita est
NUM|22|2|videns autem Balac filius Sepphor omnia quae fecerat Israhel Amorreo
NUM|22|3|et quod pertimuissent eum Moabitae et impetum eius ferre non possent
NUM|22|4|dixit ad maiores natu Madian ita delebit hic populus omnes qui in nostris finibus commorantur quomodo solet bos herbas usque ad radices carpere ipse erat eo tempore rex in Moab
NUM|22|5|misit ergo nuntios ad Balaam filium Beor ariolum qui habitabat super flumen terrae filiorum Ammon ut vocarent eum et dicerent ecce egressus est populus ex Aegypto qui operuit superficiem terrae sedens contra me
NUM|22|6|veni igitur et maledic populo huic quia fortior me est si quo modo possim percutere et eicere eum de terra mea novi enim quod benedictus sit cui benedixeris et maledictus in quem maledicta congesseris
NUM|22|7|perrexerunt seniores Moab et maiores natu Madian habentes divinationis pretium in manibus cumque venissent ad Balaam et narrassent ei omnia verba Balac
NUM|22|8|ille respondit manete hic nocte et respondebo quicquid mihi dixerit Dominus manentibus illis apud Balaam venit Deus et ait ad eum
NUM|22|9|quid sibi volunt homines isti apud te
NUM|22|10|respondit Balac filius Sepphor rex Moabitarum misit ad me
NUM|22|11|dicens ecce populus qui egressus est de Aegypto operuit superficiem terrae veni et maledic ei si quo modo possim pugnans abicere eum
NUM|22|12|dixitque Deus ad Balaam noli ire cum eis neque maledicas populo quia benedictus est
NUM|22|13|qui mane consurgens dixit ad principes ite in terram vestram quia prohibuit me Deus venire vobiscum
NUM|22|14|reversi principes dixerunt ad Balac noluit Balaam venire nobiscum
NUM|22|15|rursum ille multo plures et nobiliores quam ante miserat misit
NUM|22|16|qui cum venissent ad Balaam dixerunt sic dicit Balac filius Sepphor ne cuncteris venire ad me
NUM|22|17|paratum honorare te et quicquid volueris dare veni et maledic populo isti
NUM|22|18|respondit Balaam si dederit mihi Balac plenam domum suam argenti et auri non potero inmutare verbum Domini Dei mei ut vel plus vel minus loquar
NUM|22|19|obsecro ut hic maneatis etiam hac nocte et scire queam quid mihi rursum respondeat Dominus
NUM|22|20|venit ergo Deus ad Balaam nocte et ait ei si vocare te venerunt homines isti surge et vade cum eis ita dumtaxat ut quod tibi praecepero facias
NUM|22|21|surrexit Balaam mane et strata asina profectus est cum eis
NUM|22|22|et iratus est Deus stetitque angelus Domini in via contra Balaam qui sedebat asinae et duos pueros habebat secum
NUM|22|23|cernens asina angelum stantem in via evaginato gladio avertit se de itinere et ibat per agrum quam cum verberaret Balaam et vellet ad semitam reducere
NUM|22|24|stetit angelus in angustiis duarum maceriarum quibus vineae cingebantur
NUM|22|25|quem videns asina iunxit se parieti et adtrivit sedentis pedem at ille iterum verberabat
NUM|22|26|et nihilominus angelus ad locum angustum transiens ubi nec ad dextram nec ad sinistram poterat deviari obvius stetit
NUM|22|27|cumque vidisset asina stantem angelum concidit sub pedibus sedentis qui iratus vehementius caedebat fuste latera
NUM|22|28|aperuitque Dominus os asinae et locuta est quid feci tibi cur percutis me ecce iam tertio
NUM|22|29|respondit Balaam quia commeruisti et inlusisti mihi utinam haberem gladium ut te percuterem
NUM|22|30|dixit asina nonne animal tuum sum cui semper sedere consuesti usque in praesentem diem dic quid simile umquam fecerim tibi at ille ait numquam
NUM|22|31|protinus aperuit Dominus oculos Balaam et vidit angelum stantem in via evaginato gladio adoravitque eum pronus in terram
NUM|22|32|cui angelus cur inquit tertio verberas asinam tuam ego veni ut adversarer tibi quia perversa est via tua mihique contraria
NUM|22|33|et nisi asina declinasset de via dans locum resistenti te occidissem et illa viveret
NUM|22|34|dixit Balaam peccavi nesciens quod tu stares contra me et nunc si displicet tibi ut vadam revertar
NUM|22|35|ait angelus vade cum istis et cave ne aliud quam praecepero tibi loquaris ivit igitur cum principibus
NUM|22|36|quod cum audisset Balac egressus est in occursum eius in oppido Moabitarum quod situm est in extremis finibus Arnon
NUM|22|37|dixitque ad Balaam misi nuntios ut vocarent te cur non statim venisti ad me an quia mercedem adventui tuo reddere nequeo
NUM|22|38|cui ille respondit ecce adsum numquid loqui potero aliud nisi quod Deus posuerit in ore meo
NUM|22|39|perrexerunt ergo simul et venerunt in urbem quae in extremis regni eius finibus erat
NUM|22|40|cumque occidisset Balac boves et oves misit ad Balaam et principes qui cum eo erant munera
NUM|22|41|mane autem facto duxit eum ad excelsa Baal et intuitus est extremam partem populi
NUM|23|1|dixitque Balaam ad Balac aedifica mihi hic septem aras et para totidem vitulos eiusdemque numeri arietes
NUM|23|2|cumque fecisset iuxta sermonem Balaam inposuerunt simul vitulum et arietem super aram
NUM|23|3|dixitque Balaam ad Balac sta paulisper iuxta holocaustum tuum donec vadam si forte occurrat mihi Dominus et quodcumque imperaverit loquar tibi
NUM|23|4|cumque abisset velociter occurrit ei Deus locutusque ad eum Balaam septem inquit aras erexi et inposui vitulum et arietem desuper
NUM|23|5|Dominus autem posuit verbum in ore eius et ait revertere ad Balac et haec loqueris
NUM|23|6|reversus invenit stantem Balac iuxta holocaustum suum et omnes principes Moabitarum
NUM|23|7|adsumptaque parabola sua dixit de Aram adduxit me Balac rex Moabitarum de montibus orientis veni inquit et maledic Iacob propera et detestare Israhel
NUM|23|8|quomodo maledicam cui non maledixit Deus qua ratione detester quem Dominus non detestatur
NUM|23|9|de summis silicibus videbo eum et de collibus considerabo illum populus solus habitabit et inter gentes non reputabitur
NUM|23|10|quis dinumerare possit pulverem Iacob et nosse numerum stirpis Israhel moriatur anima mea morte iustorum et fiant novissima mea horum similia
NUM|23|11|dixitque Balac ad Balaam quid est hoc quod agis ut malediceres inimicis vocavi te et tu e contrario benedicis eis
NUM|23|12|cui ille respondit num aliud possum loqui nisi quod iusserit Dominus
NUM|23|13|dixit ergo Balac veni mecum in alterum locum unde partem Israhelis videas et totum videre non possis inde maledicito ei
NUM|23|14|cumque duxisset eum in locum sublimem super verticem montis Phasga aedificavit Balaam septem aras et inpositis supra vitulo atque ariete
NUM|23|15|dixit ad Balac sta hic iuxta holocaustum tuum donec ego pergam obvius
NUM|23|16|cui cum Dominus occurrisset posuissetque verbum in ore eius ait revertere ad Balac et haec loqueris ei
NUM|23|17|reversus invenit eum stantem iuxta holocaustum suum et principes Moabitarum cum eo ad quem Balac quid inquit locutus est Dominus
NUM|23|18|at ille adsumpta parabola sua ait sta Balac et ausculta audi fili Sepphor
NUM|23|19|non est Deus quasi homo ut mentiatur nec ut filius hominis ut mutetur dixit ergo et non faciet locutus est et non implebit
NUM|23|20|ad benedicendum adductus sum benedictionem prohibere non valeo
NUM|23|21|non est idolum in Iacob nec videtur simulacrum in Israhel Dominus Deus eius cum eo est et clangor victoriae regis in illo
NUM|23|22|Deus eduxit eum de Aegypto cuius fortitudo similis est rinocerotis
NUM|23|23|non est augurium in Iacob nec divinatio in Israhel temporibus suis dicetur Iacob et Israheli quid operatus sit Deus
NUM|23|24|ecce populus ut leaena consurget et quasi leo erigetur non accubabit donec devoret praedam et occisorum sanguinem bibat
NUM|23|25|dixitque Balac ad Balaam nec maledicas ei nec benedicas
NUM|23|26|et ille nonne ait dixi tibi quod quicquid mihi Deus imperaret hoc facerem
NUM|23|27|et ait Balac ad eum veni et ducam te ad alium locum si forte placeat Deo ut inde maledicas eis
NUM|23|28|cumque duxisset eum super verticem montis Phogor qui respicit solitudinem
NUM|23|29|dixit ei Balaam aedifica mihi hic septem aras et para totidem vitulos eiusdemque numeri arietes
NUM|23|30|fecit Balac ut Balaam dixerat inposuitque vitulos et arietes per singulas aras
NUM|24|1|cumque vidisset Balaam quod placeret Domino ut benediceret Israheli nequaquam abiit ut ante perrexerat ut augurium quaereret sed dirigens contra desertum vultum suum
NUM|24|2|et elevans oculos vidit Israhel in tentoriis commorantem per tribus suas et inruente in se spiritu Dei
NUM|24|3|adsumpta parabola ait dixit Balaam filius Beor dixit homo cuius obturatus est oculus
NUM|24|4|dixit auditor sermonum Dei qui visionem Omnipotentis intuitus est qui cadit et sic aperiuntur oculi eius
NUM|24|5|quam pulchra tabernacula tua Iacob et tentoria tua Israhel
NUM|24|6|ut valles nemorosae ut horti iuxta fluvios inrigui ut tabernacula quae fixit Dominus quasi cedri propter aquas
NUM|24|7|fluet aqua de situla eius et semen illius erit in aquas multas tolletur propter Agag rex eius et auferetur regnum illius
NUM|24|8|Deus eduxit illum de Aegypto cuius fortitudo similis est rinocerotis devorabunt gentes hostes illius ossaque eorum confringent et perforabunt sagittis
NUM|24|9|accubans dormivit ut leo et quasi leaena quam suscitare nullus audebit qui benedixerit tibi erit ipse benedictus qui maledixerit in maledictione reputabitur
NUM|24|10|iratusque Balac contra Balaam conplosis manibus ait ad maledicendum inimicis meis vocavi te quibus e contrario tertio benedixisti
NUM|24|11|revertere ad locum tuum decreveram quidem magnifice honorare te sed Dominus privavit te honore disposito
NUM|24|12|respondit Balaam ad Balac nonne nuntiis tuis quos misisti ad me dixi
NUM|24|13|si dederit mihi Balac plenam domum suam argenti et auri non potero praeterire sermonem Domini Dei mei ut vel boni quid vel mali proferam ex corde meo sed quicquid Dominus dixerit hoc loquar
NUM|24|14|verumtamen pergens ad populum meum dabo consilium quid populus tuus huic populo faciat extremo tempore
NUM|24|15|sumpta igitur parabola rursum ait dixit Balaam filius Beor dixit homo cuius obturatus est oculus
NUM|24|16|dixit auditor sermonum Dei qui novit doctrinam Altissimi et visiones Omnipotentis videt qui cadens apertos habet oculos
NUM|24|17|videbo eum sed non modo intuebor illum sed non prope orietur stella ex Iacob et consurget virga de Israhel et percutiet duces Moab vastabitque omnes filios Seth
NUM|24|18|et erit Idumea possessio eius hereditas Seir cedet inimicis suis Israhel vero fortiter aget
NUM|24|19|de Iacob erit qui dominetur et perdat reliquias civitatis
NUM|24|20|cumque vidisset Amalech adsumens parabolam ait principium gentium Amalech cuius extrema perdentur
NUM|24|21|vidit quoque Cineum et adsumpta parabola ait robustum est quidem habitaculum tuum sed si in petra posueris nidum tuum
NUM|24|22|et fueris electus de stirpe Cain quamdiu poteris permanere Assur enim capiet te
NUM|24|23|adsumptaque parabola iterum locutus est heu quis victurus est quando ista faciet Deus
NUM|24|24|venient in trieribus de Italia superabunt Assyrios vastabuntque Hebraeos et ad extremum etiam ipsi peribunt
NUM|24|25|surrexitque Balaam et reversus est in locum suum Balac quoque via qua venerat rediit
NUM|25|1|morabatur autem eo tempore Israhel in Setthim et fornicatus est populus cum filiabus Moab
NUM|25|2|quae vocaverunt eos ad sacrificia sua at illi comederunt et adoraverunt deos earum
NUM|25|3|initiatusque est Israhel Beelphegor et iratus Dominus
NUM|25|4|ait ad Mosen tolle cunctos principes populi et suspende eos contra solem in patibulis ut avertatur furor meus ab Israhel
NUM|25|5|dixitque Moses ad iudices Israhel occidat unusquisque proximos suos qui initiati sunt Beelphegor
NUM|25|6|et ecce unus de filiis Israhel intravit coram fratribus suis ad scortum madianitin vidente Mose et omni turba filiorum Israhel qui flebant ante fores tabernaculi
NUM|25|7|quod cum vidisset Finees filius Eleazari filii Aaron sacerdotis surrexit de medio multitudinis et arrepto pugione
NUM|25|8|ingressus est post virum israhelitem in lupanar et perfodit ambos simul virum scilicet et mulierem in locis genitalibus cessavitque plaga a filiis Israhel
NUM|25|9|et occisi sunt viginti quattuor milia homines
NUM|25|10|dixitque Dominus ad Mosen
NUM|25|11|Finees filius Eleazari filii Aaron sacerdotis avertit iram meam a filiis Israhel quia zelo meo commotus est contra eos ut non ipse delerem filios Israhel in zelo meo
NUM|25|12|idcirco loquere ad eos ecce do ei pacem foederis mei
NUM|25|13|et erit tam ipsi quam semini illius pactum sacerdotii sempiternum quia zelatus est pro Deo suo et expiavit scelus filiorum Israhel
NUM|25|14|erat autem nomen viri israhelitae qui occisus est cum Madianitide Zambri filius Salu dux de cognatione et tribu Symeonis
NUM|25|15|porro mulier madianitis quae pariter interfecta est vocabatur Chozbi filia Sur principis nobilissimi Madianitarum
NUM|25|16|locutusque est Dominus ad Mosen dicens
NUM|25|17|hostes vos sentiant Madianitae et percutite eos
NUM|25|18|quia et ipsi hostiliter egerunt contra vos et decepere insidiis per idolum Phogor et Chozbi filiam ducis Madian sororem suam quae percussa est in die plagae pro sacrilegio Phogor
NUM|26|1|postquam noxiorum sanguis effusus est dixit Dominus ad Mosen et Eleazarum filium Aaron sacerdotem
NUM|26|2|numerate omnem summam filiorum Israhel a viginti annis et supra per domos et cognationes suas cunctos qui possunt ad bella procedere
NUM|26|3|locuti sunt itaque Moses et Eleazar sacerdos in campestribus Moab super Iordanem contra Hierichum ad eos qui erant
NUM|26|4|a viginti annis et supra sicut Dominus imperarat quorum iste est numerus
NUM|26|5|Ruben primogenitus Israhel huius filius Enoch a quo familia Enochitarum et Phallu a quo familia Phalluitarum
NUM|26|6|et Esrom a quo familia Esromitarum et Charmi a quo familia Charmitarum
NUM|26|7|hae sunt familiae de stirpe Ruben quarum numerus inventus est quadraginta tria milia et septingenti triginta
NUM|26|8|filius Phallu Heliab
NUM|26|9|huius filii Namuhel et Dathan et Abiram isti sunt Dathan et Abiram principes populi qui surrexerunt contra Mosen et Aaron in seditione Core quando adversum Dominum rebellaverunt
NUM|26|10|et aperiens terra os suum devoravit Core morientibus plurimis quando conbusit ignis ducentos quinquaginta viros et factum est grande miraculum
NUM|26|11|ut Core pereunte filii illius non perirent
NUM|26|12|filii Symeon per cognationes suas Namuhel ab hoc familia Namuhelitarum Iamin ab hoc familia Iaminitarum Iachin ab hoc familia Iachinitarum
NUM|26|13|Zare ab hoc familia Zareitarum Saul ab hoc familia Saulitarum
NUM|26|14|hae sunt familiae de stirpe Symeon quarum omnis numerus fuit viginti duo milia ducentorum
NUM|26|15|filii Gad per cognationes suas Sephon ab hoc familia Sephonitarum Aggi ab hoc familia Aggitarum Suni ab hoc familia Sunitarum
NUM|26|16|Ozni ab hoc familia Oznitarum Heri ab hoc familia Heritarum
NUM|26|17|Arod ab hoc familia Aroditarum Arihel ab hoc familia Arihelitarum
NUM|26|18|istae sunt familiae Gad quarum omnis numerus fuit quadraginta milia quingentorum
NUM|26|19|filii Iuda Her et Onan qui ambo mortui sunt in terra Chanaan
NUM|26|20|fueruntque filii Iuda per cognationes suas Sela a quo familia Selanitarum Phares a quo familia Pharesitarum Zare a quo familia Zareitarum
NUM|26|21|porro filii Phares Esrom a quo familia Esromitarum et Amul a quo familia Amulitarum
NUM|26|22|istae sunt familiae Iuda quarum omnis numerus fuit septuaginta milia quingentorum
NUM|26|23|filii Isachar per cognationes suas Thola a quo familia Tholaitarum Phua a quo familia Phuaitarum
NUM|26|24|Iasub a quo familia Iasubitarum Semran a quo familia Semranitarum
NUM|26|25|hae sunt cognationes Isachar quarum numerus fuit sexaginta quattuor milia trecentorum
NUM|26|26|filii Zabulon per cognationes suas Sared a quo familia Sareditarum Helon a quo familia Helonitarum Ialel a quo familia Ialelitarum
NUM|26|27|hae sunt cognationes Zabulon quarum numerus fuit sexaginta milia quingentorum
NUM|26|28|filii Ioseph per cognationes suas Manasse et Ephraim
NUM|26|29|de Manasse ortus est Machir a quo familia Machiritarum Machir genuit Galaad a quo familia Galaaditarum
NUM|26|30|Galaad habuit filios Hiezer a quo familia Hiezeritarum et Elec a quo familia Elecarum
NUM|26|31|et Asrihel a quo familia Asrihelitarum et Sechem a quo familia Sechemitarum
NUM|26|32|et Semida a quo familia Semidatarum et Epher a quo familia Epheritarum
NUM|26|33|fuit autem Epher pater Salphaad qui filios non habebat sed tantum filias quarum ista sunt nomina Maala et Noa et Egla et Melcha et Thersa
NUM|26|34|hae sunt familiae Manasse et numerus earum quinquaginta duo milia septingentorum
NUM|26|35|filii autem Ephraim per cognationes suas fuerunt hii Suthala a quo familia Suthalitarum Becher a quo familia Becheritarum Tehen a quo familia Tehenitarum
NUM|26|36|porro filius Suthala fuit Heran a quo familia Heranitarum
NUM|26|37|hae sunt cognationes filiorum Ephraim quarum numerus triginta duo milia quingentorum
NUM|26|38|isti sunt filii Ioseph per familias suas filii Beniamin in cognationibus suis Bale a quo familia Baleitarum Azbel a quo familia Azbelitarum Ahiram a quo familia Ahiramitarum
NUM|26|39|Supham a quo familia Suphamitarum Hupham a quo familia Huphamitarum
NUM|26|40|filii Bale Hered et Noeman de Hered familia Hereditarum de Noeman familia Noemitarum
NUM|26|41|hii sunt filii Beniamin per cognationes suas quorum numerus quadraginta quinque milia sescentorum
NUM|26|42|filii Dan per cognationes suas Suham a quo familia Suhamitarum hae cognationes Dan per familias suas
NUM|26|43|omnes fuere Suhamitae quorum numerus erat sexaginta quattuor milia quadringentorum
NUM|26|44|filii Aser per cognationes suas Iemna a quo familia Iemnaitarum Iessui a quo familia Iessuitarum Brie a quo familia Brieitarum
NUM|26|45|filii Brie Haber a quo familia Haberitarum et Melchihel a quo familia Melchihelitarum
NUM|26|46|nomen autem filiae Aser fuit Sara
NUM|26|47|hae cognationes filiorum Aser et numerus eorum quinquaginta tria milia quadringentorum
NUM|26|48|filii Nepthalim per cognationes suas Iessihel a quo familia Iessihelitarum Guni a quo familia Gunitarum
NUM|26|49|Iesser a quo familia Iesseritarum Sellem a quo familia Sellemitarum
NUM|26|50|hae sunt cognationes filiorum Nepthalim per familias suas quorum numerus quadraginta quinque milia quadringentorum
NUM|26|51|ista est summa filiorum Israhel qui recensiti sunt sescenta milia et mille septingenti triginta
NUM|26|52|locutusque est Dominus ad Mosen dicens
NUM|26|53|istis dividetur terra iuxta numerum vocabulorum in possessiones suas
NUM|26|54|pluribus maiorem partem dabis et paucioribus minorem singulis sicut nunc recensiti sunt tradetur possessio
NUM|26|55|ita dumtaxat ut sors terram tribubus dividat et familiis
NUM|26|56|quicquid sorte contigerit hoc vel plures accipient vel pauciores
NUM|26|57|hic quoque est numerus filiorum Levi per familias suas Gerson a quo familia Gersonitarum Caath a quo familia Caathitarum Merari a quo familia Meraritarum
NUM|26|58|hae sunt familiae Levi familia Lobni familia Hebroni familia Mooli familia Musi familia Cori at vero Caath genuit Amram
NUM|26|59|qui habuit uxorem Iochabed filiam Levi quae nata est ei in Aegypto haec genuit viro suo Amram filios Aaron et Mosen et Mariam sororem eorum
NUM|26|60|de Aaron orti sunt Nadab et Abiu et Eleazar et Ithamar
NUM|26|61|quorum Nadab et Abiu mortui sunt cum obtulissent ignem alienum coram Domino
NUM|26|62|fueruntque omnes qui numerati sunt viginti tria milia generis masculini ab uno mense et supra quia non sunt recensiti inter filios Israhel nec eis cum ceteris data possessio
NUM|26|63|hic est numerus filiorum Israhel qui descripti sunt a Mosen et Eleazaro sacerdote in campestribus Moab supra Iordanem contra Hiericho
NUM|26|64|inter quos nullus fuit eorum qui ante numerati sunt a Mose et Aaron in deserto Sinai
NUM|26|65|praedixerat enim Dominus quod omnes morerentur in solitudine nullusque remansit ex eis nisi Chaleb filius Iepphonne et Iosue filius Nun
NUM|27|1|accesserunt autem filiae Salphaad filii Epher filii Galaad filii Machir filii Manasse qui fuit filius Ioseph quarum sunt nomina Maala et Noa et Egla et Melcha et Thersa
NUM|27|2|steteruntque coram Mosen et Eleazaro sacerdote et cunctis principibus populi ad ostium tabernaculi foederis atque dixerunt
NUM|27|3|pater noster mortuus est in deserto nec fuit in seditione quae concitata est contra Dominum sub Core sed in peccato suo mortuus est hic non habuit mares filios cur tollitur nomen illius de familia sua quia non habet filium date nobis possessionem inter cognatos patris nostri
NUM|27|4|rettulitque Moses causam earum ad iudicium Domini
NUM|27|5|qui dixit ad eum
NUM|27|6|iustam rem postulant filiae Salphaad da eis possessionem inter cognatos patris sui et ei in hereditate succedant
NUM|27|7|ad filios autem Israhel loqueris haec
NUM|27|8|homo cum mortuus fuerit absque filio ad filiam eius transibit hereditas
NUM|27|9|si filiam non habuerit habebit successores fratres suos
NUM|27|10|quod si et fratres non fuerint dabitis hereditatem fratribus patris eius
NUM|27|11|sin autem nec patruos habuerit dabitur hereditas his qui ei proximi sunt eritque hoc filiis Israhel sanctum lege perpetua sicut praecepit Dominus Mosi
NUM|27|12|dixit quoque Dominus ad Mosen ascende in montem istum Abarim et contemplare inde terram quam daturus sum filiis Israhel
NUM|27|13|cumque videris eam ibis et tu ad populum tuum sicut ivit frater tuus Aaron
NUM|27|14|quia offendistis me in deserto Sin in contradictione multitudinis nec sanctificare me voluistis coram ea super aquas hae sunt aquae Contradictionis in Cades deserti Sin
NUM|27|15|cui respondit Moses
NUM|27|16|provideat Dominus Deus spirituum omnis carnis hominem qui sit super multitudinem hanc
NUM|27|17|et possit exire et intrare ante eos et educere illos vel introducere ne sit populus Domini sicut oves absque pastore
NUM|27|18|dixitque Dominus ad eum tolle Iosue filium Nun virum in quo est spiritus et pone manum tuam super eum
NUM|27|19|qui stabit coram Eleazaro sacerdote et omni multitudine
NUM|27|20|et dabis ei praecepta cunctis videntibus et partem gloriae tuae ut audiat eum omnis synagoga filiorum Israhel
NUM|27|21|pro hoc si quid agendum erit Eleazar sacerdos consulet Dominum ad verbum eius egredietur et ingredietur ipse et omnes filii Israhel cum eo et cetera multitudo
NUM|27|22|fecit Moses ut praeceperat Dominus cumque tulisset Iosue statuit eum coram Eleazaro sacerdote et omni frequentia populi
NUM|27|23|et inpositis capiti eius manibus cuncta replicavit quae mandaverat Dominus
NUM|28|1|dixit quoque Dominus ad Mosen
NUM|28|2|praecipe filiis Israhel et dices ad eos oblationem meam et panes et incensum odoris suavissimi offerte per tempora sua
NUM|28|3|haec sunt sacrificia quae offerre debetis agnos anniculos inmaculatos duos cotidie in holocaustum sempiternum
NUM|28|4|unum offeretis mane et alterum ad vesperam
NUM|28|5|decimam partem oephi similae quae conspersa sit oleo purissimo et habeat quartam partem hin
NUM|28|6|holocaustum iuge est quod obtulistis in monte Sinai in odorem suavissimum incensi Domini
NUM|28|7|et libabitis vini quartam partem hin per agnos singulos in sanctuario Domini
NUM|28|8|alterumque agnum similiter offeretis ad vesperam iuxta omnem ritum sacrificii matutini et libamentorum eius oblationem suavissimi odoris Domino
NUM|28|9|die autem sabbati offeretis duos agnos anniculos inmaculatos et duas decimas similae oleo conspersae in sacrificio et liba
NUM|28|10|quae rite funduntur per singula sabbata in holocausto sempiterno
NUM|28|11|in kalendis autem id est in mensuum exordiis offeretis holocaustum Domino vitulos de armento duos arietem unum agnos anniculos septem inmaculatos
NUM|28|12|et tres decimas similae oleo conspersae in sacrificio per singulos vitulos et duas decimas similae oleo conspersae per singulos arietes
NUM|28|13|et decimam decimae similae ex oleo in sacrificio per agnos singulos holocaustum suavissimi odoris atque incensi est Domino
NUM|28|14|libamenta autem vini quae per singulas fundenda sunt victimas ista erunt media pars hin per vitulos singulos tertia per arietem quarta per agnum hoc erit holocaustum per omnes menses qui sibi anno vertente succedunt
NUM|28|15|hircus quoque offeretur Domino pro peccatis in holocaustum sempiternum cum libamentis suis
NUM|28|16|mense autem primo quartadecima die mensis phase Domini erit
NUM|28|17|et quintadecima die sollemnitas septem diebus vescentur azymis
NUM|28|18|quarum dies prima venerabilis et sancta erit omne opus servile non facietis in ea
NUM|28|19|offeretisque incensum holocaustum Domino vitulos de armento duos arietem unum agnos anniculos inmaculatos septem
NUM|28|20|et sacrificia singulorum ex simila quae conspersa sit oleo tres decimas per singulos vitulos et duas decimas per arietem
NUM|28|21|et decimam decimae per agnos singulos id est per septem agnos
NUM|28|22|et hircum pro peccato unum ut expietur pro vobis
NUM|28|23|praeter holocaustum matutinum quod semper offertis
NUM|28|24|ita facietis per singulos dies septem dierum in fomitem ignis et in odorem suavissimum Domino qui surget de holocausto et de libationibus singulorum
NUM|28|25|dies quoque septimus celeberrimus et sanctus erit vobis omne opus servile non facietis in eo
NUM|28|26|dies etiam primitivorum quando offertis novas fruges Domino expletis ebdomadibus venerabilis et sancta erit omne opus servile non facietis in ea
NUM|28|27|offeretisque holocaustum in odorem suavissimum Domino vitulos de armento duos arietem unum et agnos anniculos inmaculatos septem
NUM|28|28|atque in sacrificiis eorum similae oleo conspersae tres decimas per singulos vitulos per arietes duas
NUM|28|29|per agnos decimam decimae qui simul sunt agni septem hircum quoque
NUM|28|30|qui mactatur pro expiatione praeter holocaustum sempiternum et liba eius
NUM|28|31|inmaculata offeretis omnia cum libationibus suis
NUM|29|1|mensis etiam septimi prima dies venerabilis et sancta erit vobis omne opus servile non facietis in ea quia dies clangoris est et tubarum
NUM|29|2|offeretisque holocaustum in odorem suavissimum Domino vitulum de armento unum arietem unum agnos anniculos inmaculatos septem
NUM|29|3|et in sacrificiis eorum similae oleo conspersae tres decimas per singulos vitulos duas decimas per arietem
NUM|29|4|unam decimam per agnum qui simul sunt agni septem
NUM|29|5|et hircum pro peccato qui offertur in expiationem populi
NUM|29|6|praeter holocaustum kalendarum cum sacrificiis suis et holocaustum sempiternum cum libationibus solitis hisdem caerimoniis offeretis in odorem suavissimum incensum Domino
NUM|29|7|decima quoque dies mensis huius septimi erit vobis sancta atque venerabilis et adfligetis animas vestras omne opus servile non facietis in ea
NUM|29|8|offeretisque holocaustum Domino in odorem suavissimum vitulum de armento unum arietem unum agnos anniculos inmaculatos septem
NUM|29|9|et in sacrificiis eorum similae oleo conspersae tres decimas per vitulos singulos duas decimas per arietem
NUM|29|10|decimam decimae per agnos singulos qui sunt simul septem agni
NUM|29|11|et hircum pro peccato absque his quae offerri pro delicto solent in expiationem et holocaustum sempiternum in sacrificio et libaminibus eorum
NUM|29|12|quintadecima vero die mensis septimi quae vobis erit sancta atque venerabilis omne opus servile non facietis in ea sed celebrabitis sollemnitatem Domino septem diebus
NUM|29|13|offeretisque holocaustum in odorem suavissimum Domino vitulos de armento tredecim arietes duos agnos anniculos quattuordecim inmaculatos
NUM|29|14|et in libamentis eorum similae oleo conspersae tres decimas per vitulos singulos qui sunt simul vituli tredecim et duas decimas arieti uno id est simul arietibus duobus
NUM|29|15|et decimam decimae agnis singulis qui sunt simul agni quattuordecim
NUM|29|16|et hircum pro peccato absque holocausto sempiterno et sacrificio et libamine eius
NUM|29|17|in die altero offeres vitulos de armento duodecim arietes duos agnos anniculos inmaculatos quattuordecim
NUM|29|18|sacrificiaque et libamina singulorum per vitulos et arietes et agnos rite celebrabis
NUM|29|19|et hircum pro peccato absque holocausto sempiterno sacrificioque eius et libamine
NUM|29|20|die tertio offeres vitulos undecim arietes duos agnos anniculos inmaculatos quattuordecim
NUM|29|21|sacrificiaque et libamina singulorum per vitulos et arietes et agnos rite celebrabis
NUM|29|22|et hircum pro peccato absque holocausto sempiterno et sacrificio et libamine eius
NUM|29|23|die quarto offeres vitulos decem arietes duos agnos anniculos inmaculatos quattuordecim
NUM|29|24|sacrificiaque eorum et libamina singulorum per vitulos et arietes et agnos rite celebrabis
NUM|29|25|et hircum pro peccato absque holocausto sempiterno sacrificioque eius et libamine
NUM|29|26|die quinto offeres vitulos novem arietes duos agnos anniculos inmaculatos quattuordecim
NUM|29|27|sacrificiaque et libamina singulorum per vitulos et arietes et agnos rite celebrabis
NUM|29|28|et hircum pro peccato absque holocausto sempiterno sacrificioque eius et libamine
NUM|29|29|die sexto offeres vitulos octo arietes duos agnos anniculos inmaculatos quattuordecim
NUM|29|30|sacrificiaque et libamina singulorum per vitulos et arietes et agnos rite celebrabis
NUM|29|31|et hircum pro peccato absque holocausto sempiterno sacrificioque eius et libamine
NUM|29|32|die septimo offeres vitulos septem arietes duos agnos anniculos inmaculatos quattuordecim
NUM|29|33|sacrificiaque et libamina singulorum per vitulos et arietes et agnos rite celebrabis
NUM|29|34|et hircum pro peccato absque holocausto sempiterno sacrificioque eius et libamine
NUM|29|35|die octavo qui est celeberrimus omne opus servile non facietis
NUM|29|36|offerentes holocaustum in odorem suavissimum Domino vitulum unum arietem unum agnos anniculos inmaculatos septem
NUM|29|37|sacrificiaque et libamina singulorum per vitulos et arietes et agnos rite celebrabis
NUM|29|38|et hircum pro peccato absque holocausto sempiterno sacrificioque eius et libamine
NUM|29|39|haec offeretis Domino in sollemnitatibus vestris praeter vota et oblationes spontaneas in holocausto in sacrificio in libamine et in hostiis pacificis
NUM|30|1|narravitque Moses filiis Israhel omnia quae ei Dominus imperarat
NUM|30|2|et locutus est ad principes tribuum filiorum Israhel iste est sermo quem praecepit Dominus
NUM|30|3|si quis virorum votum Domino voverit aut se constrinxerit iuramento non faciet irritum verbum suum sed omne quod promisit implebit
NUM|30|4|mulier si quippiam voverit et se constrinxerit iuramento quae est in domo patris sui et in aetate adhuc puellari si cognoverit pater votum quod pollicita est et iuramentum quo obligavit animam suam et tacuerit voti rea erit
NUM|30|5|quicquid pollicita est et iuravit opere conplebit
NUM|30|6|sin autem statim ut audierit contradixerit pater et vota et iuramenta eius irrita erunt nec obnoxia tenebitur sponsioni eo quod contradixerit pater
NUM|30|7|si maritum habuerit et voverit aliquid et semel verbum de ore eius egrediens animam illius obligaverit iuramento
NUM|30|8|quo die audierit vir et non contradixerit voti rea erit reddet quodcumque promiserat
NUM|30|9|sin autem audiens statim contradixerit et irritas fecerit pollicitationes eius verbaque quibus obstrinxerat animam suam propitius ei erit Dominus
NUM|30|10|vidua et repudiata quicquid voverint reddent
NUM|30|11|uxor in domo viri cum se voto constrinxerit et iuramento
NUM|30|12|si audierit vir et tacuerit nec contradixerit sponsioni reddet quodcumque promiserat
NUM|30|13|sin autem extemplo contradixerit non tenebitur promissionis rea quia maritus contradixit et Dominus ei propitius erit
NUM|30|14|si voverit et iuramento se constrinxerit ut per ieiunium vel ceterarum rerum abstinentiam adfligat animam suam in arbitrio viri erit ut faciat sive non faciat
NUM|30|15|quod si audiens vir tacuerit et in alteram diem distulerit sententiam quicquid voverat atque promiserat reddet quia statim ut audivit tacuit
NUM|30|16|sin autem contradixerit postquam rescivit portabit ipse iniquitatem eius
NUM|30|17|istae sunt leges quas constituit Dominus Mosi inter virum et uxorem inter patrem et filiam quae in puellari adhuc aetate est vel quae manet in parentis domo
NUM|31|1|locutusque est Dominus ad Mosen dicens
NUM|31|2|ulciscere prius filios Israhel de Madianitis et sic colligeris ad populum tuum
NUM|31|3|statimque Moses armate inquit ex vobis viros ad pugnam qui possint ultionem Domini expetere de Madianitis
NUM|31|4|mille viri de singulis tribubus eligantur Israhel qui mittantur ad bellum
NUM|31|5|dederuntque millenos de cunctis tribubus id est duodecim milia expeditorum ad pugnam
NUM|31|6|quos misit Moses cum Finees filio Eleazari sacerdotis vasa quoque sancta et tubas ad clangendum tradidit ei
NUM|31|7|cumque pugnassent contra Madianitas atque vicissent omnes mares occiderunt
NUM|31|8|et reges eorum Evi et Recem et Sur et Ur et Rebe quinque principes gentis Balaam quoque filium Beor interfecerunt gladio
NUM|31|9|ceperuntque mulieres eorum et parvulos omniaque pecora et cunctam supellectilem quicquid habere potuerant depopulati sunt
NUM|31|10|tam urbes quam viculos et castella flamma consumpsit
NUM|31|11|et tulerunt praedam et universa quae ceperant tam ex hominibus quam ex iumentis
NUM|31|12|et adduxerunt ad Mosen et Eleazarum sacerdotem et ad omnem multitudinem filiorum Israhel reliqua etiam utensilia portaverunt ad castra in campestribus Moab iuxta Iordanem contra Hiericho
NUM|31|13|egressi sunt autem Moses et Eleazar sacerdos et omnes principes synagogae in occursum eorum extra castra
NUM|31|14|iratusque Moses principibus exercitus tribunis et centurionibus qui venerant de bello
NUM|31|15|ait cur feminas reservastis
NUM|31|16|nonne istae sunt quae deceperunt filios Israhel ad suggestionem Balaam et praevaricari vos fecerunt in Domino super peccato Phogor unde et percussus est populus
NUM|31|17|ergo cunctos interficite quicquid est generis masculini etiam in parvulis et mulieres quae noverunt viros in coitu iugulate
NUM|31|18|puellas autem et omnes feminas virgines reservate vobis
NUM|31|19|et manete extra castra septem diebus qui occiderit hominem vel occisum tetigerit lustrabitur die tertio et septimo
NUM|31|20|et de omni praeda sive vestimentum fuerit sive vas et aliquid in utensilia praeparatum de caprarum pellibus et pilis et ligno expiabitur
NUM|31|21|Eleazar quoque sacerdos ad viros exercitus qui pugnaverant sic locutus est hoc est praeceptum legis quod mandavit Dominus Mosi
NUM|31|22|aurum et argentum et aes et ferrum et stagnum et plumbum
NUM|31|23|et omne quod potest transire per flammas igne purgabitur quicquid autem ignem non potest sustinere aqua expiationis sanctificabitur
NUM|31|24|et lavabitis vestimenta vestra die septimo et purificati postea castra intrabitis
NUM|31|25|dixitque Dominus ad Mosen
NUM|31|26|tollite summam eorum quae capta sunt ab homine usque ad pecus tu et Eleazar sacerdos et principes vulgi
NUM|31|27|dividesque ex aequo praedam inter eos qui pugnaverunt et egressi sunt ad bellum et inter omnem reliquam multitudinem
NUM|31|28|et separabis partem Domino ab his qui pugnaverunt et fuerunt in bello unam animam de quingentis tam ex hominibus quam ex bubus et asinis et ovibus
NUM|31|29|et dabis eam Eleazaro sacerdoti quia primitiae Domini sunt
NUM|31|30|ex media quoque parte filiorum Israhel accipies quinquagesimum caput hominum et boum et asinorum et ovium cunctarumque animantium et dabis ea Levitis qui excubant in custodiis tabernaculi Domini
NUM|31|31|feceruntque Moses et Eleazar sicut praeceperat Dominus
NUM|31|32|fuit autem praeda quam exercitus ceperat ovium sescenta septuaginta quinque milia
NUM|31|33|boum septuaginta duo milia
NUM|31|34|asinorum sexaginta milia et mille
NUM|31|35|animae hominum sexus feminei quae non cognoverant viros triginta duo milia
NUM|31|36|dataque est media pars his qui in proelio fuerant ovium trecenta triginta septem milia quingenta
NUM|31|37|e quibus in partem Domini supputatae sunt oves sescentae septuaginta quinque
NUM|31|38|et de bubus triginta sex milibus boves septuaginta duo
NUM|31|39|de asinis triginta milibus quingentis asini sexaginta unus
NUM|31|40|de animabus hominum sedecim milibus cesserunt in partem Domini triginta duae animae
NUM|31|41|tradiditque Moses numerum primitiarum Domini Eleazaro sacerdoti sicut ei fuerat imperatum
NUM|31|42|ex media parte filiorum Israhel quam separaverat his qui in proelio fuerant
NUM|31|43|de media vero parte quae contigerat reliquae multitudini id est de ovium trecentis triginta septem milibus quingentis
NUM|31|44|et de bubus triginta sex milibus
NUM|31|45|et de asinis triginta milibus quingentis
NUM|31|46|et de hominibus sedecim milibus
NUM|31|47|tulit Moses quinquagesimum caput et dedit Levitis qui excubant in tabernaculo Domini sicut praeceperat Dominus
NUM|31|48|cumque accessissent principes exercitus ad Mosen et tribuni centurionesque dixerunt
NUM|31|49|nos servi tui recensuimus numerum pugnatorum quos habuimus sub manu nostra et ne unus quidem defuit
NUM|31|50|ob hanc causam offerimus in donariis Domini singuli quod in praeda auri potuimus invenire periscelides et armillas anulos et dextralia ac murenulas ut depreceris pro nobis Dominum
NUM|31|51|susceperuntque Moses et Eleazar sacerdos omne aurum in diversis speciebus
NUM|31|52|pondo sedecim milia septingentos quinquaginta siclos a tribunis et centurionibus
NUM|31|53|unusquisque enim quod in praeda rapuerat suum erat
NUM|31|54|et susceptum intulerunt in tabernaculum testimonii in monumentum filiorum Israhel coram Domino
NUM|32|1|filii autem Ruben et Gad habebant pecora multa et erat illis in iumentis infinita substantia cumque vidissent Iazer et Galaad aptas alendis animalibus
NUM|32|2|venerunt ad Mosen et ad Eleazarum sacerdotem et principes multitudinis atque dixerunt
NUM|32|3|Atharoth et Dibon et Iazer et Nemra Esbon et Eleale et Sabam et Nebo et Beon
NUM|32|4|terram quam percussit Dominus in conspectu filiorum Israhel regionis uberrimae est ad pastum animalium et nos servi tui habemus iumenta plurima
NUM|32|5|precamurque si invenimus gratiam coram te ut des nobis famulis tuis eam in possessionem ne facias nos transire Iordanem
NUM|32|6|quibus respondit Moses numquid fratres vestri ibunt ad pugnam et vos hic sedebitis
NUM|32|7|cur subvertitis mentes filiorum Israhel ne transire audeant in locum quem eis daturus est Dominus
NUM|32|8|nonne ita egerunt patres vestri quando misi de Cadesbarne ad explorandam terram
NUM|32|9|cumque venissent usque ad vallem Botri lustrata omni regione subverterunt cor filiorum Israhel ut non intrarent fines quos eis Dominus dedit
NUM|32|10|qui iratus iuravit dicens
NUM|32|11|si videbunt homines isti qui ascenderunt ex Aegypto a viginti annis et supra terram quam sub iuramento pollicitus sum Abraham Isaac et Iacob et noluerunt sequi me
NUM|32|12|praeter Chaleb filium Iepphonne Cenezeum et Iosue filium Nun isti impleverunt voluntatem meam
NUM|32|13|iratusque Dominus adversum Israhel circumduxit eum per desertum quadraginta annis donec consumeretur universa generatio quae fecerat malum in conspectu eius
NUM|32|14|et ecce inquit vos surrexistis pro patribus vestris incrementa et alumni hominum peccatorum ut augeretis furorem Domini contra Israhel
NUM|32|15|qui si nolueritis sequi eum in solitudine populum derelinquet et vos causa eritis necis omnium
NUM|32|16|at illi prope accedentes dixerunt caulas ovium fabricabimus et stabula iumentorum parvulis quoque nostris urbes munitas
NUM|32|17|nos autem ipsi armati et accincti pergemus ad proelium ante filios Israhel donec introducamus eos ad loca sua parvuli nostri et quicquid habere possumus erunt in urbibus muratis propter habitatorum insidias
NUM|32|18|non revertemur in domos nostras usquequo possideant filii Israhel hereditatem suam
NUM|32|19|nec quicquam quaeremus trans Iordanem quia iam habemus possessionem nostram in orientali eius plaga
NUM|32|20|quibus Moses ait si facitis quod promittitis expediti pergite coram Domino ad pugnam
NUM|32|21|et omnis vir bellator armatus Iordanem transeat donec subvertat Dominus inimicos suos
NUM|32|22|et subiciatur ei omnis terra tunc eritis inculpabiles et apud Dominum et apud Israhel et obtinebitis regiones quas vultis coram Domino
NUM|32|23|sin autem quod dicitis non feceritis nulli dubium quin peccetis in Dominum et scitote quoniam peccatum vestrum adprehendet vos
NUM|32|24|aedificate ergo urbes parvulis vestris et caulas ac stabula ovibus ac iumentis et quod polliciti estis implete
NUM|32|25|dixeruntque filii Gad et Ruben ad Mosen servi tui sumus faciemus quod iubet dominus noster
NUM|32|26|parvulos nostros et mulieres et pecora ac iumenta relinquemus in urbibus Galaad
NUM|32|27|nos autem famuli tui omnes expediti pergemus ad bellum sicut tu domine loqueris
NUM|32|28|praecepit ergo Moses Eleazaro sacerdoti et Iosue filio Nun et principibus familiarum per tribus Israhel et dixit ad eos
NUM|32|29|si transierint filii Gad et filii Ruben vobiscum Iordanem omnes armati ad bellum coram Domino et vobis fuerit terra subiecta date eis Galaad in possessionem
NUM|32|30|sin autem noluerint transire vobiscum in terram Chanaan inter vos habitandi accipiant loca
NUM|32|31|responderuntque filii Gad et filii Ruben sicut locutus est Dominus servis suis ita faciemus
NUM|32|32|ipsi armati pergemus coram Domino in terram Chanaan et possessionem iam suscepisse nos confitemur trans Iordanem
NUM|32|33|dedit itaque Moses filiis Gad et Ruben et dimidiae tribui Manasse filii Ioseph regnum Seon regis Amorrei et regnum Og regis Basan et terram eorum cum urbibus suis per circuitum
NUM|32|34|igitur extruxerunt filii Gad Dibon et Atharoth et Aroer
NUM|32|35|Etrothsophan et Iazer Iecbaa
NUM|32|36|et Bethnemra et Betharan urbes munitas et caulas pecoribus suis
NUM|32|37|filii vero Ruben aedificaverunt Esbon et Eleale et Cariathaim
NUM|32|38|et Nabo et Baalmeon versis nominibus Sabama quoque inponentes vocabula urbibus quas extruxerant
NUM|32|39|porro filii Machir filii Manasse perrexerunt in Galaad et vastaverunt eam interfecto Amorreo habitatore eius
NUM|32|40|dedit ergo Moses terram Galaad Machir filio Manasse qui habitavit in ea
NUM|32|41|Iair autem filius Manasse abiit et occupavit vicos eius quos appellavit Avothiair id est villas Iair
NUM|32|42|Nobe quoque perrexit et adprehendit Canath cum viculis suis vocavitque eam ex nomine suo Nobe
NUM|33|1|hae sunt mansiones filiorum Israhel qui egressi sunt de Aegypto per turmas suas in manu Mosi et Aaron
NUM|33|2|quas descripsit Moses iuxta castrorum loca quae Domini iussione mutabant
NUM|33|3|profecti igitur de Ramesse mense primo quintadecima die mensis primi altera die phase filii Israhel in manu excelsa videntibus cunctis Aegyptiis
NUM|33|4|et sepelientibus primogenitos quos percusserat Dominus nam et in diis eorum exercuerat ultionem
NUM|33|5|castrametati sunt in Soccoth
NUM|33|6|et de Soccoth venerunt in Aetham quae est in extremis finibus solitudinis
NUM|33|7|inde egressi venerunt contra Phiahiroth quae respicit Beelsephon et castrametati sunt ante Magdolum
NUM|33|8|profectique de Phiahiroth transierunt per medium mare in solitudinem et ambulantes tribus diebus per desertum Aetham castrametati sunt in Mara
NUM|33|9|profectique de Mara venerunt in Helim ubi erant duodecim fontes aquarum et palmae septuaginta ibique castrametati sunt
NUM|33|10|sed et inde egressi fixere tentoria super mare Rubrum profectique de mari Rubro
NUM|33|11|castrametati sunt in deserto Sin
NUM|33|12|unde egressi venerunt in Dephca
NUM|33|13|profectique de Dephca castrametati sunt in Alus
NUM|33|14|egressi de Alus Raphidim fixere tentoria ubi aqua populo defuit ad bibendum
NUM|33|15|profectique de Raphidim castrametati sunt in deserto Sinai
NUM|33|16|sed et de solitudine Sinai egressi venerunt ad sepulchra Concupiscentiae
NUM|33|17|profectique de sepulchris Concupiscentiae castrametati sunt in Aseroth
NUM|33|18|et de Aseroth venerunt in Rethma
NUM|33|19|profectique de Rethma castrametati sunt in Remmonphares
NUM|33|20|unde egressi venerunt in Lebna
NUM|33|21|et de Lebna castrametati sunt in Ressa
NUM|33|22|egressi de Ressa venerunt in Ceelatha
NUM|33|23|unde profecti castrametati sunt in monte Sepher
NUM|33|24|egressi de monte Sepher venerunt in Arada
NUM|33|25|inde proficiscentes castrametati sunt in Maceloth
NUM|33|26|profectique de Maceloth venerunt in Thaath
NUM|33|27|de Thaath castrametati sunt in Thare
NUM|33|28|unde egressi fixerunt tentoria in Methca
NUM|33|29|et de Methca castrametati sunt in Esmona
NUM|33|30|profectique de Esmona venerunt in Moseroth
NUM|33|31|et de Moseroth castrametati sunt in Baneiacan
NUM|33|32|egressique de Baneiacan venerunt in montem Gadgad
NUM|33|33|unde profecti castrametati sunt in Hietebatha
NUM|33|34|et de Hietebatha venerunt in Ebrona
NUM|33|35|egressique de Ebrona castrametati sunt in Asiongaber
NUM|33|36|inde profecti venerunt in desertum Sin haec est Cades
NUM|33|37|egressique de Cades castrametati sunt in monte Hor in extremis finibus terrae Edom
NUM|33|38|ascenditque Aaron sacerdos montem Hor iubente Domino et ibi mortuus est anno quadragesimo egressionis filiorum Israhel ex Aegypto mense quinto prima die mensis
NUM|33|39|cum esset annorum centum viginti trium
NUM|33|40|audivitque Chananeus rex Arad qui habitabat ad meridiem in terra Chanaan venisse filios Israhel
NUM|33|41|et profecti de monte Hor castrametati sunt in Salmona
NUM|33|42|unde egressi venerunt in Phinon
NUM|33|43|profectique de Phinon castrametati sunt in Oboth
NUM|33|44|et de Oboth venerunt in Ieabarim quae est in finibus Moabitarum
NUM|33|45|profectique de Ieabarim fixere tentoria in Dibongad
NUM|33|46|unde egressi castrametati sunt in Elmondeblathaim
NUM|33|47|egressi de Elmondeblathaim venerunt ad montes Abarim contra Nabo
NUM|33|48|profectique de montibus Abarim transierunt ad campestria Moab super Iordanem contra Hiericho
NUM|33|49|ibique castrametati sunt de Bethsimon usque ad Belsattim in planioribus locis Moabitarum
NUM|33|50|ubi locutus est Dominus ad Mosen
NUM|33|51|praecipe filiis Israhel et dic ad eos quando transieritis Iordanem intrantes terram Chanaan
NUM|33|52|disperdite cunctos habitatores regionis illius confringite titulos et statuas comminuite atque omnia excelsa vastate
NUM|33|53|mundantes terram et habitantes in ea ego enim dedi vobis illam in possessionem
NUM|33|54|quam dividetis vobis sorte pluribus dabitis latiorem et paucis angustiorem singulis ut sors ceciderit ita tribuetur hereditas per tribus et familias possessio dividetur
NUM|33|55|sin autem nolueritis interficere habitatores terrae qui remanserint erunt vobis quasi clavi in oculis et lanceae in lateribus et adversabuntur vobis in terra habitationis vestrae
NUM|33|56|et quicquid illis facere cogitaram vobis faciam
NUM|34|1|locutus est Dominus ad Mosen
NUM|34|2|praecipe filiis Israhel et dices ad eos cum ingressi fueritis terram Chanaan et in possessionem vobis sorte ceciderit his finibus terminabitur
NUM|34|3|pars meridiana incipiet a solitudine Sin quae est iuxta Edom et habebit terminos contra orientem mare Salsissimum
NUM|34|4|qui circumibunt australem plagam per ascensum Scorpionis ita ut transeant Senna et perveniant in meridiem usque ad Cadesbarne unde egredientur confinia ad villam nomine Addar et tendent usque Asemona
NUM|34|5|ibitque per gyrum terminus ab Asemona usque ad torrentem Aegypti et maris Magni litore finietur
NUM|34|6|plaga autem occidentalis a mari Magno incipiet et ipso fine cludetur
NUM|34|7|porro ad septentrionalem plagam a mari Magno termini incipient pervenientes usque ad montem Altissimum
NUM|34|8|a quo venies in Emath usque ad terminos Sedada
NUM|34|9|ibuntque confinia usque Zephrona et villam Henan hii erunt termini in parte aquilonis
NUM|34|10|inde metabuntur fines contra orientalem plagam de villa Henan usque Sephama
NUM|34|11|et de Sephama descendent termini in Rebla contra fontem inde pervenient contra orientem ad mare Chenereth
NUM|34|12|et tendent usque Iordanem et ad ultimum Salsissimo cludentur mari hanc habebitis terram per fines suos in circuitu
NUM|34|13|praecepitque Moses filiis Israhel dicens haec erit terra quam possidebitis sorte et quam iussit dari Dominus novem tribubus et dimidiae tribui
NUM|34|14|tribus enim filiorum Ruben per familias suas et tribus filiorum Gad iuxta cognationum numerum media quoque tribus Manasse
NUM|34|15|id est duae semis tribus acceperunt partem suam trans Iordanem contra Hiericho ad orientalem plagam
NUM|34|16|et ait Dominus ad Mosen
NUM|34|17|haec sunt nomina virorum qui terram vobis divident Eleazar sacerdos et Iosue filius Nun
NUM|34|18|et singuli principes de tribubus singulis
NUM|34|19|quorum ista sunt vocabula de tribu Iuda Chaleb filius Iepphonne
NUM|34|20|de tribu Symeon Samuhel filius Ammiud
NUM|34|21|de tribu Beniamin Helidad filius Chaselon
NUM|34|22|de tribu filiorum Dan Bocci filius Iogli
NUM|34|23|filiorum Ioseph de tribu Manasse Hannihel filius Ephod
NUM|34|24|de tribu Ephraim Camuhel filius Sephtan
NUM|34|25|de tribu Zabulon Elisaphan filius Pharnach
NUM|34|26|de tribu Isachar dux Faltihel filius Ozan
NUM|34|27|de tribu Aser Ahiud filius Salomi
NUM|34|28|de tribu Nepthali Phedahel filius Ameiud
NUM|34|29|hii sunt quibus praecepit Dominus ut dividerent filiis Israhel terram Chanaan
NUM|35|1|haec quoque locutus est Dominus ad Mosen in campestribus Moab super Iordanem contra Hiericho
NUM|35|2|praecipe filiis Israhel ut dent Levitis de possessionibus suis
NUM|35|3|urbes ad habitandum et suburbana earum per circuitum ut ipsi in oppidis maneant et suburbana sint pecoribus ac iumentis
NUM|35|4|quae a muris civitatum forinsecus per circuitum mille passuum spatio tendentur
NUM|35|5|contra orientem duo milia erunt cubiti et contra meridiem similiter duo milia ad mare quoque quod respicit occidentem eadem mensura erit et septentrionalis plaga aequali termino finietur eruntque urbes in medio et foris suburbana
NUM|35|6|de ipsis autem oppidis quae Levitis dabitis sex erunt in fugitivorum auxilia separata ut fugiat ad ea qui fuderit sanguinem exceptis his alia quadraginta duo oppida
NUM|35|7|id est simul quadraginta octo cum suburbanis suis
NUM|35|8|ipsaeque urbes quae dabuntur de possessionibus filiorum Israhel ab his qui plus habent plures auferentur et qui minus pauciores singuli iuxta mensuram hereditatis suae dabunt oppida Levitis
NUM|35|9|ait Dominus ad Mosen
NUM|35|10|loquere filiis Israhel et dices ad eos quando transgressi fueritis Iordanem in terram Chanaan
NUM|35|11|decernite quae urbes esse debeant in praesidia fugitivorum qui nolentes sanguinem fuderint
NUM|35|12|in quibus cum fuerit profugus cognatus occisi eum non poterit occidere donec stet in conspectu multitudinis et causa illius iudicetur
NUM|35|13|de ipsis autem urbibus quae ad fugitivorum subsidia separantur
NUM|35|14|tres erunt trans Iordanem et tres in terra Chanaan
NUM|35|15|tam filiis Israhel quam advenis atque peregrinis ut confugiat ad eas qui nolens sanguinem fuderit
NUM|35|16|si quis ferro percusserit et mortuus fuerit qui percussus est reus erit homicidii et ipse morietur
NUM|35|17|si lapidem iecerit et ictus occubuerit similiter punietur
NUM|35|18|si ligno percussus interierit percussoris sanguine vindicabitur
NUM|35|19|propinquus occisi homicidam interficiet statim ut adprehenderit eum percutiet
NUM|35|20|si per odium quis hominem inpulerit vel iecerit quippiam in eum per insidias
NUM|35|21|aut cum esset inimicus manu percusserit et ille mortuus fuerit percussor homicidii reus erit cognatus occisi statim ut invenerit eum iugulabit
NUM|35|22|quod si fortuito et absque odio
NUM|35|23|et inimicitiis quicquam horum fecerit
NUM|35|24|et hoc audiente populo fuerit conprobatum atque inter percussorem et propinquum sanguinis quaestio ventilata
NUM|35|25|liberabitur innocens de ultoris manu et reducetur per sententiam in urbem ad quam confugerat manebitque ibi donec sacerdos magnus qui oleo sancto unctus est moriatur
NUM|35|26|si interfector extra fines urbium quae exulibus deputatae sunt
NUM|35|27|fuerit inventus et percussus ab eo qui ultor est sanguinis absque noxa erit qui eum occiderit
NUM|35|28|debuerat enim profugus usque ad mortem pontificis in urbe residere postquam autem ille obierit homicida revertetur in terram suam
NUM|35|29|haec sempiterna erunt et legitima in cunctis habitationibus vestris
NUM|35|30|homicida sub testibus punietur ad unius testimonium nullus condemnabitur
NUM|35|31|non accipietis pretium ab eo qui reus est sanguinis statim et ipse morietur
NUM|35|32|exules et profugi ante mortem pontificis nullo modo in urbes suas reverti poterunt
NUM|35|33|ne polluatis terram habitationis vestrae quae insontium cruore maculatur nec aliter expiari potest nisi per eius sanguinem qui alterius sanguinem fuderit
NUM|35|34|atque ita emundabitur vestra possessio me commorante vobiscum ego enim sum Dominus qui habito inter filios Israhel
NUM|36|1|accesserunt autem et principes familiarum Galaad filii Machir filii Manasse de stirpe filiorum Ioseph locutique sunt Mosi coram principibus Israhel atque dixerunt
NUM|36|2|tibi domino nostro praecepit Dominus ut terram sorte divideres filiis Israhel et ut filiabus Salphaad fratris nostri dares possessionem debitam patri
NUM|36|3|quas si alterius tribus homines uxores acceperint sequetur possessio sua et translata ad aliam tribum de nostra hereditate minuetur
NUM|36|4|atque ita fiet ut cum iobeleus id est quinquagesimus annus remissionis advenerit confundatur sortium distributio et aliorum possessio ad alios transeat
NUM|36|5|respondit Moses filiis Israhel et Domino praecipiente ait recte tribus filiorum Ioseph locuta est
NUM|36|6|et haec lex super filiabus Salphaad a Domino promulgata est nubant quibus volunt tantum ut suae tribus hominibus
NUM|36|7|ne commisceatur possessio filiorum Israhel de tribu in tribum omnes enim viri ducent uxores de tribu et cognatione sua
NUM|36|8|et cunctae feminae maritos de eadem tribu accipient ut hereditas permaneat in familiis
NUM|36|9|nec sibi misceantur tribus sed ta maneant
NUM|36|10|ut a Domino separatae sunt feceruntque filiae Salphaad ut fuerat imperatum
NUM|36|11|et nupserunt Maala et Thersa et Egla et Melcha et Noa filiis patrui sui
NUM|36|12|de familia Manasse qui fuit filius Ioseph et possessio quae illis fuerat adtributa mansit in tribu et familia patris earum
NUM|36|13|haec sunt mandata atque iudicia quae praecepit Dominus per manum Mosi ad filios Israhel in campestribus Moab super Iordanem contra Hiericho
