2TIM|1|1|Paul, an apostle of Jesus Christ by the will of God, according to the promise of life which is in Christ Jesus,
2TIM|1|2|To Timothy, my dearly beloved son: Grace, mercy, and peace, from God the Father and Christ Jesus our Lord.
2TIM|1|3|I thank God, whom I serve from my forefathers with pure conscience, that without ceasing I have remembrance of thee in my prayers night and day;
2TIM|1|4|Greatly desiring to see thee, being mindful of thy tears, that I may be filled with joy;
2TIM|1|5|When I call to remembrance the unfeigned faith that is in thee, which dwelt first in thy grandmother Lois, and thy mother Eunice; and I am persuaded that in thee also.
2TIM|1|6|Wherefore I put thee in remembrance that thou stir up the gift of God, which is in thee by the putting on of my hands.
2TIM|1|7|For God hath not given us the spirit of fear; but of power, and of love, and of a sound mind.
2TIM|1|8|Be not thou therefore ashamed of the testimony of our Lord, nor of me his prisoner: but be thou partaker of the afflictions of the gospel according to the power of God;
2TIM|1|9|Who hath saved us, and called us with an holy calling, not according to our works, but according to his own purpose and grace, which was given us in Christ Jesus before the world began,
2TIM|1|10|But is now made manifest by the appearing of our Saviour Jesus Christ, who hath abolished death, and hath brought life and immortality to light through the gospel:
2TIM|1|11|Whereunto I am appointed a preacher, and an apostle, and a teacher of the Gentiles.
2TIM|1|12|For the which cause I also suffer these things: nevertheless I am not ashamed: for I know whom I have believed, and am persuaded that he is able to keep that which I have committed unto him against that day.
2TIM|1|13|Hold fast the form of sound words, which thou hast heard of me, in faith and love which is in Christ Jesus.
2TIM|1|14|That good thing which was committed unto thee keep by the Holy Ghost which dwelleth in us.
2TIM|1|15|This thou knowest, that all they which are in Asia be turned away from me; of whom are Phygellus and Hermogenes.
2TIM|1|16|The Lord give mercy unto the house of Onesiphorus; for he oft refreshed me, and was not ashamed of my chain:
2TIM|1|17|But, when he was in Rome, he sought me out very diligently, and found me.
2TIM|1|18|The Lord grant unto him that he may find mercy of the Lord in that day: and in how many things he ministered unto me at Ephesus, thou knowest very well.
2TIM|2|1|Thou therefore, my son, be strong in the grace that is in Christ Jesus.
2TIM|2|2|And the things that thou hast heard of me among many witnesses, the same commit thou to faithful men, who shall be able to teach others also.
2TIM|2|3|Thou therefore endure hardness, as a good soldier of Jesus Christ.
2TIM|2|4|No man that warreth entangleth himself with the affairs of this life; that he may please him who hath chosen him to be a soldier.
2TIM|2|5|And if a man also strive for masteries, yet is he not crowned, except he strive lawfully.
2TIM|2|6|The husbandman that laboureth must be first partaker of the fruits.
2TIM|2|7|Consider what I say; and the Lord give thee understanding in all things.
2TIM|2|8|Remember that Jesus Christ of the seed of David was raised from the dead according to my gospel:
2TIM|2|9|Wherein I suffer trouble, as an evil doer, even unto bonds; but the word of God is not bound.
2TIM|2|10|Therefore I endure all things for the elect's sakes, that they may also obtain the salvation which is in Christ Jesus with eternal glory.
2TIM|2|11|It is a faithful saying: For if we be dead with him, we shall also live with him:
2TIM|2|12|If we suffer, we shall also reign with him: if we deny him, he also will deny us:
2TIM|2|13|If we believe not, yet he abideth faithful: he cannot deny himself.
2TIM|2|14|Of these things put them in remembrance, charging them before the Lord that they strive not about words to no profit, but to the subverting of the hearers.
2TIM|2|15|Study to shew thyself approved unto God, a workman that needeth not to be ashamed, rightly dividing the word of truth.
2TIM|2|16|But shun profane and vain babblings: for they will increase unto more ungodliness.
2TIM|2|17|And their word will eat as doth a canker: of whom is Hymenaeus and Philetus;
2TIM|2|18|Who concerning the truth have erred, saying that the resurrection is past already; and overthrow the faith of some.
2TIM|2|19|Nevertheless the foundation of God standeth sure, having this seal, The Lord knoweth them that are his. And, Let every one that nameth the name of Christ depart from iniquity.
2TIM|2|20|But in a great house there are not only vessels of gold and of silver, but also of wood and of earth; and some to honour, and some to dishonour.
2TIM|2|21|If a man therefore purge himself from these, he shall be a vessel unto honour, sanctified, and meet for the master's use, and prepared unto every good work.
2TIM|2|22|Flee also youthful lusts: but follow righteousness, faith, charity, peace, with them that call on the Lord out of a pure heart.
2TIM|2|23|But foolish and unlearned questions avoid, knowing that they do gender strifes.
2TIM|2|24|And the servant of the Lord must not strive; but be gentle unto all men, apt to teach, patient,
2TIM|2|25|In meekness instructing those that oppose themselves; if God peradventure will give them repentance to the acknowledging of the truth;
2TIM|2|26|And that they may recover themselves out of the snare of the devil, who are taken captive by him at his will.
2TIM|3|1|This know also, that in the last days perilous times shall come.
2TIM|3|2|For men shall be lovers of their own selves, covetous, boasters, proud, blasphemers, disobedient to parents, unthankful, unholy,
2TIM|3|3|Without natural affection, trucebreakers, false accusers, incontinent, fierce, despisers of those that are good,
2TIM|3|4|Traitors, heady, highminded, lovers of pleasures more than lovers of God;
2TIM|3|5|Having a form of godliness, but denying the power thereof: from such turn away.
2TIM|3|6|For of this sort are they which creep into houses, and lead captive silly women laden with sins, led away with divers lusts,
2TIM|3|7|Ever learning, and never able to come to the knowledge of the truth.
2TIM|3|8|Now as Jannes and Jambres withstood Moses, so do these also resist the truth: men of corrupt minds, reprobate concerning the faith.
2TIM|3|9|But they shall proceed no further: for their folly shall be manifest unto all men, as their's also was.
2TIM|3|10|But thou hast fully known my doctrine, manner of life, purpose, faith, longsuffering, charity, patience,
2TIM|3|11|Persecutions, afflictions, which came unto me at Antioch, at Iconium, at Lystra; what persecutions I endured: but out of them all the Lord delivered me.
2TIM|3|12|Yea, and all that will live godly in Christ Jesus shall suffer persecution.
2TIM|3|13|But evil men and seducers shall wax worse and worse, deceiving, and being deceived.
2TIM|3|14|But continue thou in the things which thou hast learned and hast been assured of, knowing of whom thou hast learned them;
2TIM|3|15|And that from a child thou hast known the holy scriptures, which are able to make thee wise unto salvation through faith which is in Christ Jesus.
2TIM|3|16|All scripture is given by inspiration of God, and is profitable for doctrine, for reproof, for correction, for instruction in righteousness:
2TIM|3|17|That the man of God may be perfect, throughly furnished unto all good works.
2TIM|4|1|I charge thee therefore before God, and the Lord Jesus Christ, who shall judge the quick and the dead at his appearing and his kingdom;
2TIM|4|2|Preach the word; be instant in season, out of season; reprove, rebuke, exhort with all longsuffering and doctrine.
2TIM|4|3|For the time will come when they will not endure sound doctrine; but after their own lusts shall they heap to themselves teachers, having itching ears;
2TIM|4|4|And they shall turn away their ears from the truth, and shall be turned unto fables.
2TIM|4|5|But watch thou in all things, endure afflictions, do the work of an evangelist, make full proof of thy ministry.
2TIM|4|6|For I am now ready to be offered, and the time of my departure is at hand.
2TIM|4|7|I have fought a good fight, I have finished my course, I have kept the faith:
2TIM|4|8|Henceforth there is laid up for me a crown of righteousness, which the Lord, the righteous judge, shall give me at that day: and not to me only, but unto all them also that love his appearing.
2TIM|4|9|Do thy diligence to come shortly unto me:
2TIM|4|10|For Demas hath forsaken me, having loved this present world, and is departed unto Thessalonica; Crescens to Galatia, Titus unto Dalmatia.
2TIM|4|11|Only Luke is with me. Take Mark, and bring him with thee: for he is profitable to me for the ministry.
2TIM|4|12|And Tychicus have I sent to Ephesus.
2TIM|4|13|The cloke that I left at Troas with Carpus, when thou comest, bring with thee, and the books, but especially the parchments.
2TIM|4|14|Alexander the coppersmith did me much evil: the Lord reward him according to his works:
2TIM|4|15|Of whom be thou ware also; for he hath greatly withstood our words.
2TIM|4|16|At my first answer no man stood with me, but all men forsook me: I pray God that it may not be laid to their charge.
2TIM|4|17|Notwithstanding the Lord stood with me, and strengthened me; that by me the preaching might be fully known, and that all the Gentiles might hear: and I was delivered out of the mouth of the lion.
2TIM|4|18|And the Lord shall deliver me from every evil work, and will preserve me unto his heavenly kingdom: to whom be glory for ever and ever. Amen.
2TIM|4|19|Salute Prisca and Aquila, and the household of Onesiphorus.
2TIM|4|20|Erastus abode at Corinth: but Trophimus have I left at Miletum sick.
2TIM|4|21|Do thy diligence to come before winter. Eubulus greeteth thee, and Pudens, and Linus, and Claudia, and all the brethren.
2TIM|4|22|The Lord Jesus Christ be with thy spirit. Grace be with you. Amen.
