NEH|1|1|哈迦利亞 的兒子 尼希米 的言語如下： 亞達薛西 王二十年基斯流月，我在 書珊 城堡中。
NEH|1|2|那時，我有一個兄弟 哈拿尼 ，同幾個人從 猶大 來。我問他們那些被擄歸回、剩下殘存的 猶太 人和 耶路撒冷 的情況。
NEH|1|3|他們對我說：「那些被擄歸回剩下的餘民在 猶大 省那裏遭大難，受凌辱； 耶路撒冷 的城牆被拆毀，城門被火焚燒。」
NEH|1|4|我聽見這話，就坐下哭泣，悲哀幾日，在天上的上帝面前禁食祈禱，
NEH|1|5|說：「唉，耶和華－天上大而可畏的上帝，向愛你、守你誡命的人守約施慈愛的上帝啊，
NEH|1|6|願你睜眼看，側耳聽你僕人今日晝夜在你面前，為你眾僕人 以色列 人的祈禱，承認我們 以色列 人向你所犯的罪；我與我父家都犯了罪。
NEH|1|7|我們向你所行的非常敗壞，沒有遵守你吩咐你僕人 摩西 的誡命、律例、典章。
NEH|1|8|求你記念所吩咐你僕人 摩西 的話，說：『你們若犯罪，我就把你們分散在萬民中；
NEH|1|9|但你們若歸向我，謹守遵行我的誡命，你們被趕散的人雖在天涯，我也必從那裏將他們召集回來，帶到我所選擇立為我名居所的地方。』
NEH|1|10|他們是你的僕人和你的百姓，是你用大力和大能的手所救贖的。
NEH|1|11|唉，主啊，求你側耳聽你僕人的祈禱，聽喜愛敬畏你名眾僕人的祈禱，使你僕人今日亨通，在這人面前蒙恩。」 我是王的酒政。
NEH|2|1|亞達薛西 王二十年尼散月，酒擺在王面前 ，我拿起酒來奉給王。我在王面前從來沒有愁容。
NEH|2|2|王對我說：「你既沒有病，為甚麼面帶愁容呢？這不是別的，必是你心中愁煩。」於是我非常懼怕。
NEH|2|3|我對王說：「願王萬歲！我祖先墳墓所在的那城荒涼，城門被火焚燒，我豈能面無愁容呢？」
NEH|2|4|王對我說：「你想求甚麼？」於是我向天上的上帝祈禱。
NEH|2|5|我對王說：「王若以為好，僕人若在王面前蒙恩，求王差遣我往 猶大 ，到我祖先墳墓所在的那城去，我好重新建造。」
NEH|2|6|那時王后坐在王的旁邊，王對我說：「你要去多久？幾時回來？」王看這事為好，就派我去。我給王定了日期。
NEH|2|7|我又對王說：「王若以為好，求王賜我詔書，通知 河西 的省長准我經過，直到 猶大 ；
NEH|2|8|又賜詔書，通知管理王園林的 亞薩 ，叫他給我木材，作為殿的營樓之門、城牆，和我自己要住的房屋的橫梁。」王就允准我，因為我上帝施恩的手幫助我。
NEH|2|9|王派了軍官和騎兵護送我。我到了 河西 的省長那裏，將王的詔書交給他們。
NEH|2|10|和倫 人 參巴拉 和作臣僕的 亞捫 人 多比雅 ，聽見有人來為 以色列 人爭取利益，就很惱怒。
NEH|2|11|我到了 耶路撒冷 ，在那裏停留了三天。
NEH|2|12|夜間我和跟隨我的幾個人起來；但上帝感動我心要為 耶路撒冷 做的事，我並沒有告訴人。只有我自己騎的牲口，沒有別的牲口在我那裏。
NEH|2|13|當夜，我出了 谷門 ，往 野狗泉 去，到了 糞廠門 ，察看 耶路撒冷 的城牆，城牆被拆毀，城門被火焚燒。
NEH|2|14|我又往前，到了 泉門 ，又到 王池 ，但所騎的牲口沒有地方可以過去。
NEH|2|15|於是我夜間沿溪而上，察看城牆，又轉身進入 谷門 ，就回來了。
NEH|2|16|我往哪裏去，我做甚麼事，官長都不知道。我也沒有告訴 猶大 人、祭司、貴族、官長和其餘做工的人。
NEH|2|17|以後，我對他們說：「我們所遭的難， 耶路撒冷 怎樣荒涼，城門被火焚燒，你們都看見了。來吧，讓我們重建 耶路撒冷 的城牆，免得再受凌辱！」
NEH|2|18|我告訴他們我上帝施恩的手怎樣幫助我，以及王向我所說的話。他們就說：「我們起來建造吧！」於是他們使自己的手堅強，做這美好的工作。
NEH|2|19|但 和倫 人 參巴拉 、作臣僕的 亞捫 人 多比雅 和 阿拉伯 人 基善 聽見就嗤笑我們，藐視我們，說：「你們所做的這事是甚麼呢？要背叛王嗎？」
NEH|2|20|我回答他們的話，對他們說：「天上的上帝必使我們亨通。我們作他僕人的，要起來建造；你們卻在 耶路撒冷 無份、無權、無名號 。」
NEH|3|1|那時， 以利亞實 大祭司和他的弟兄眾祭司起來建立 羊門 ，將門分別為聖，安立門扇，直到 哈米亞樓 。他們又將它分別為聖，直到 哈楠業樓 。
NEH|3|2|在他旁邊建造的是 耶利哥 人。在他旁邊建造的是 音利 的兒子 撒刻 。
NEH|3|3|哈西拿 的子孫建立 魚門 ，架橫梁、安門扇，裝閂和鎖。
NEH|3|4|在他們旁邊修造的是 哈哥斯 的孫子， 烏利亞 的兒子 米利末 。在他們旁邊修造的是 米示薩別 的孫子， 比利迦 的兒子 米書蘭 。在他們旁邊修造的是 巴拿 的兒子 撒督 。
NEH|3|5|在他們旁邊修造的是 提哥亞 人；但是他們的貴族不用肩 扛他們主人的工作。
NEH|3|6|巴西亞 的兒子 耶何耶大 與 比所玳 的兒子 米書蘭 修造 古門 ，架橫梁，安門扇，裝閂和鎖。
NEH|3|7|在他們旁邊修造的是 基遍 人 米拉提 、 米倫 人 雅頓 、 基遍 人，和 河西 總督所管的 米斯巴 人。
NEH|3|8|在他旁邊修造的是 哈海雅 的兒子 烏薛 銀匠。在他旁邊修造的是做香料的 哈拿尼雅 。他們修復 耶路撒冷 ，直到 寬牆 。
NEH|3|9|在他們旁邊修造的是管理 耶路撒冷 城區的一半、 戶珥 的兒子 利法雅 。
NEH|3|10|在他們旁邊的是 哈路抹 的兒子 耶大雅 在自己房屋的對面修造。在他旁邊修造的是 哈沙尼 的兒子 哈突 。
NEH|3|11|哈琳 的兒子 瑪基雅 和 巴哈‧摩押 的兒子 哈述 修造下一段和 爐樓 。
NEH|3|12|在他旁邊修造的是管理 耶路撒冷 城區的另一半、 哈羅黑 的兒子 沙龍 和他的女兒們。
NEH|3|13|哈嫩 和 撒挪亞 的居民修造 谷門 ；他們立門，安門扇，裝閂和鎖，又修造城牆一千肘，直到 糞廠門 。
NEH|3|14|管理 伯‧哈基琳 區、 利甲 的兒子 瑪基雅 修造 糞廠門 ；他立門，安門扇，裝閂和鎖。
NEH|3|15|管理 米斯巴 區、 各‧荷西 的兒子 沙崙 修造 泉門 ；他立門，蓋門頂，安門扇，裝閂和鎖，又修造靠近王的花園 西羅亞池 的城牆，直到那從 大衛城 下來的臺階。
NEH|3|16|接續他修造的是管理 伯‧夙 區的一半、 押卜 的兒子 尼希米 ，直到 大衛 墳地的對面，又到人造池，到達勇士的房屋。
NEH|3|17|接續他修造的是 利未 人 巴尼 的兒子 利宏 。在他旁邊的是管理 基伊拉 區一半的 哈沙比雅 為本區修造。
NEH|3|18|接續他修造的是他們弟兄中管理 基伊拉 區的另一半、 希拿達 的兒子 賓內 。
NEH|3|19|在他旁邊的是管理 米斯巴 、 耶書亞 的兒子 以謝珥 修造武庫的上坡對面、城牆轉彎處的那一段。
NEH|3|20|接續他的是 薩拜 的兒子 巴錄 竭力修造下一段，從轉彎處，直到 以利亞實 大祭司的府門。
NEH|3|21|接續他的是 哈哥斯 的孫子， 烏利亞 的兒子 米利末 修造下一段，從 以利亞實 的府門，直到 以利亞實 府的盡頭。
NEH|3|22|接續他修造的是住平原的祭司。
NEH|3|23|接續他的是 便雅憫 與 哈述 在自己房屋的對面修造。接續他的是 亞難尼 的孫子， 瑪西雅 的兒子 亞撒利雅 在自己房屋的旁邊修造。
NEH|3|24|接續他的是 希拿達 的兒子 賓內 修造下一段，從 亞撒利雅 的房屋直到轉彎處，又到城角。
NEH|3|25|烏賽 的兒子 巴拉 修造轉彎處的對面和靠近護衛院、王宮上層凸出來的城樓。接續他的是 巴錄 的兒子 毗大雅 ，
NEH|3|26|（殿役住在 俄斐勒 ，直到朝東 水門 的對面和凸出來的城樓。）
NEH|3|27|接續他的是 提哥亞 人又修造一段，對著那凸出來的大城樓，直到 俄斐勒 的城牆。
NEH|3|28|從 馬門 往上，祭司各在自己房屋的對面修造。
NEH|3|29|接續他的是 音麥 的兒子 撒督 在自己房屋的對面修造。接續他修造的是 東門 的守衛、 示迦尼 的兒子 示瑪雅 。
NEH|3|30|接續他的是 示利米雅 的兒子 哈拿尼雅 和 薩拉 的第六個兒子 哈嫩 修造下一段。接續他的是 比利迦 的兒子 米書蘭 在自己房屋的對面修造。
NEH|3|31|接續他的是 瑪基雅 銀匠修造，直到殿役和商人的房屋，對著 集合門 ，直到角樓。
NEH|3|32|銀匠與商人在角樓和 羊門 之間修造。
NEH|4|1|參巴拉 聽見我們建造城牆就發怒，非常惱恨，並嗤笑 猶太 人。
NEH|4|2|他對他的弟兄和 撒瑪利亞 的軍兵說：「這些軟弱的 猶太 人做甚麼呢？要為自己重建嗎 ？要獻祭嗎？要一日完工嗎？要使土堆裏火燒過的石頭再有用嗎？」
NEH|4|3|亞捫 人 多比雅 在一旁說：「他們所修造的石牆，就是狐狸上去也必崩裂。」
NEH|4|4|我們的上帝啊，求你垂聽，因為我們被藐視。求你使他們的毀謗歸於他們自己頭上，使他們在被擄之地成為掠物。
NEH|4|5|不要遮掩他們的罪孽，不要使他們的罪惡從你面前塗去，因為他們在修造的人前面惹你發怒。
NEH|4|6|這樣，我們修造城牆，整個城牆就連接起來，到一半高，因為百姓一心做工。
NEH|4|7|參巴拉 、 多比雅 、 阿拉伯 人、 亞捫 人和 亞實突 人聽見 耶路撒冷 城牆正在修造，破裂的地方開始進行修補，就非常憤怒。
NEH|4|8|大家同謀要來攻打 耶路撒冷 ，使城混亂。
NEH|4|9|然而，我們向我們的上帝禱告，又因他們的緣故，就派人站崗，晝夜防備他們。
NEH|4|10|但 猶大 有話說： 「扛抬的人力氣衰弱， 瓦礫太多， 我們自己不可能 建造城牆。」
NEH|4|11|我們的敵人說：「趁他們不知道，看不見的時候，我們進入他們中間，殺了他們，使工作停止。」
NEH|4|12|那靠近敵人居住的 猶太 人十次從各處來見我們，說：「你們必須回到我們那裏。」
NEH|4|13|我叫百姓站在城牆後邊低窪的空處，使百姓各按宗族站著，拿刀、拿槍、拿弓。
NEH|4|14|我察看了，就起來對貴族、官長和其餘的百姓說：「不要怕他們！當記得主是大而可畏的。你們要為你們的弟兄、兒女、妻子、家園爭戰。」
NEH|4|15|仇敵聽見我們知道了他們的計謀，上帝也破壞他們的計謀，我們就都回到城牆那裏，各做各的工。
NEH|4|16|從那日起，我的僕人一半做工，一半拿槍、拿盾牌、拿弓、穿鎧甲，官長都站在 猶大 全家的後邊。
NEH|4|17|他們建造城牆；扛抬材料的人扛抬的時候，一手做工，一手拿兵器。
NEH|4|18|建造的人都腰間佩刀建造，吹角的人在我旁邊。
NEH|4|19|我對貴族、官長和其餘的百姓說：「這工程浩大，範圍遼闊，我們在城牆上彼此相離很遠。
NEH|4|20|你們一聽見角聲在哪裏，就聚集到我們那裏去。我們的上帝必為我們爭戰。」
NEH|4|21|於是，我們做這工程，一半的人拿槍，從天亮直到星宿出現的時候。
NEH|4|22|那時，我又對百姓說：「各人和他的僕人當在 耶路撒冷 過夜，好為我們夜間守衛，白晝做工。」
NEH|4|23|這樣，我和弟兄僕人，以及跟從我的衛兵都不脫衣服，各人打水時 也拿著自己的兵器。
NEH|5|1|百姓和他們的妻子大大呼號，埋怨他們的弟兄 猶太 人。
NEH|5|2|有的說：「我們和兒女人口眾多，必須得糧食吃，才能活下去。」
NEH|5|3|有的說：「我們典押了田地、葡萄園、房屋，才得糧食充飢。」
NEH|5|4|有的說：「我們借了錢付田地和葡萄園的稅給王。
NEH|5|5|現在，我們的身體與我們弟兄的身體是一樣的，我們的兒女與他們的兒女沒有差別。看哪，我們卻要迫使兒女作人的奴婢。我們有些女兒已被搶走了，我們卻無能為力，因為我們的田地和葡萄園已經歸了別人。」
NEH|5|6|我聽見他們的呼號和這些話，就非常憤怒。
NEH|5|7|我心裏作了決定，就斥責貴族和官長，對他們說：「你們各人借錢給弟兄，竟然索取利息！」於是我召開大會攻擊他們。
NEH|5|8|我對他們說：「我們已盡力贖回我們的弟兄，就是賣到列國的 猶太 人；你們還要賣弟兄，讓我們去買回來嗎？」他們就靜默不語，無話可答。
NEH|5|9|我又說：「你們做的這事不對！你們行事不是應該敬畏我們的上帝，免得列國我們的仇敵毀謗我們嗎？
NEH|5|10|我和我的弟兄僕人也要把銀錢糧食借給百姓，大家都當免除利息。
NEH|5|11|就在今日，你們要把他們的田地、葡萄園、橄欖園、房屋，以及向他們所取銀錢的利息 、糧食、新酒和新油都歸還他們。」
NEH|5|12|貴族和官長說：「我們必歸還，不再向他們索取，必照你所說的去做。」我就召了祭司來，叫貴族和官長起誓，必照這話去做。
NEH|5|13|我也抖著胸前的衣袋，說：「凡不實行這話的，願上帝照樣抖他離開他的家和他勞碌得來的，直到抖空了。」全會眾都說：「阿們！」又讚美耶和華。百姓就照著這話去做。
NEH|5|14|自從我奉派作 猶大 地省長的那日，就是從 亞達薛西 王二十年直到三十二年，共十二年之久，我與我弟兄都沒有吃省長的俸祿。
NEH|5|15|在我以前的省長加重百姓的負擔，向百姓索取糧食和酒，以及四十舍客勒銀子 ，甚至他們的僕人也轄制百姓，但我因敬畏上帝不這樣做。
NEH|5|16|我也努力修造城牆。我們並沒有購置田地，我所有的僕人也都聚集在那裏做工。
NEH|5|17|除了從四圍列國來的人以外，有 猶太 人和官長一百五十人與我同席。
NEH|5|18|每日預備一頭公牛，六隻肥羊，又為我預備飛禽；每十日一次多多預備各樣的酒。雖然如此，我並不索取省長的俸祿，因為這百姓負的勞役很重。
NEH|5|19|我的上帝啊，求你記念我為這百姓所做的一切，施恩於我。
NEH|6|1|參巴拉 、 多比雅 、 阿拉伯 人 基善 和我們其餘的仇敵聽見我已經建造了城牆，沒有破裂之處在其中，那時我還沒有在城門安門扇；
NEH|6|2|參巴拉 和 基善 就派人來見我，說：「請你來，我們在 阿挪 平原的村莊見面。」其實，他們想要害我。
NEH|6|3|於是我派使者到他們那裏，說：「我正在進行大的工程，不能下去。我怎麼能離開，下去見你們，而讓工程停頓呢？」
NEH|6|4|他們這樣派人來見我四次，我都用這話回答他們。
NEH|6|5|參巴拉 第五次同樣派僕人來見我，手裏拿著未封的信，
NEH|6|6|信上寫著：「列國中有風聲， 基善 也說，你和 猶太 人謀反，所以你建造城牆。據說，你要作他們的王，
NEH|6|7|並且你派先知在 耶路撒冷 指著你宣講說，『在 猶大 有王。』如今這些話必傳給王知，現在請你來，我們一起商議。」
NEH|6|8|我就派人到他那裏，說：「你所說的這些事，一概沒有，是你心裏捏造的。」
NEH|6|9|他們全都要使我們懼怕，說：「他們的手必軟弱，不能工作，以致不能完工。」現在，求你堅固我的手。
NEH|6|10|我到了 米希大別 的孫子， 第來雅 的兒子 示瑪雅 家裏；那時，他閉門不出。他說：「我們可以在上帝的殿裏，就在殿的中間會面，鎖住殿門，因為他們要來殺你，要在夜裏來殺你。」
NEH|6|11|我說：「像我這樣的人豈會逃跑呢？像我這樣的人豈能進入殿裏保全生命呢？我不進去！」
NEH|6|12|我看清楚了，看哪，上帝並沒有派他，是他自己說預言攻擊我，是 多比雅 和 參巴拉 收買了他；
NEH|6|13|收買他的目的是要叫我懼怕，依從他犯罪，留下一個壞名聲，好讓他們毀謗我。
NEH|6|14|我的上帝啊，求你記得 多比雅 、 參巴拉 、 挪亞底 女先知和其餘的先知，因他們行這些事，要叫我懼怕。
NEH|6|15|以祿月二十五日，城牆修完了，共修了五十二天。
NEH|6|16|我們所有的仇敵聽見了，四圍的列國就懼怕，愁眉不展，因為他們知道這工作得以完成，是出於我們的上帝。
NEH|6|17|而且，在那些日子， 猶大 的貴族屢次寄信給 多比雅 ， 多比雅 也回信給他們。
NEH|6|18|在 猶大 有許多人與 多比雅 結盟，因為他是 亞拉 的兒子 示迦尼 的女婿，並且他的兒子 約哈難 娶了 比利迦 的兒子 米書蘭 的女兒。
NEH|6|19|他們也在我面前說 多比雅 的好話，又把我的話傳給他。 多比雅 常寄信來，要叫我懼怕。
NEH|7|1|城牆修完，我安了門扇，門口的守衛、歌唱的和 利未 人都已派定。
NEH|7|2|我吩咐我的兄弟 哈拿尼 和城堡的官長 哈拿尼雅 管理 耶路撒冷 ，因為 哈拿尼雅 是一個忠信的人，敬畏上帝過於眾人。
NEH|7|3|我對他們說：「等到太陽熱的時候才可開 耶路撒冷 的城門；要派 耶路撒冷 的居民，各按班次在自己房屋的前面站崗。他們還在站崗的時候，就要關門上閂。」
NEH|7|4|城又寬又大，城中的百姓卻稀少，房屋也還沒有建造。
NEH|7|5|我的上帝感動我的心，我就召集貴族、官長和百姓，要登記家譜。我找到第一次上來之人的家譜，發現上面寫著：
NEH|7|6|這些是從被擄之地上來的省民， 巴比倫 王 尼布甲尼撒 把他們擄去，他們重返 耶路撒冷 和 猶大 ，各歸本城。
NEH|7|7|他們是同 所羅巴伯 、 耶書亞 、 尼希米 、 亞撒利雅 、 拉米 、 拿哈瑪尼 、 末底改 、 必珊 、 米斯毗列 、 比革瓦伊 、 尼宏 、 巴拿 一起回來的。 以色列 百姓的人數如下：
NEH|7|8|巴錄 的子孫二千一百七十二名；
NEH|7|9|示法提雅 的子孫三百七十二名；
NEH|7|10|亞拉 的子孫六百五十二名；
NEH|7|11|巴哈‧摩押 的後裔，就是 耶書亞 和 約押 的子孫二千八百一十八名；
NEH|7|12|以攔 的子孫一千二百五十四名；
NEH|7|13|薩土 的子孫八百四十五名；
NEH|7|14|薩改 的子孫七百六十名；
NEH|7|15|賓內 的子孫六百四十八名；
NEH|7|16|比拜 的子孫六百二十八名；
NEH|7|17|押甲 的子孫二千三百二十二名；
NEH|7|18|亞多尼干 的子孫六百六十七名；
NEH|7|19|比革瓦伊 的子孫二千零六十七名；
NEH|7|20|亞丁 的子孫六百五十五名；
NEH|7|21|亞特 的後裔，就是 希西家 的子孫九十八名；
NEH|7|22|哈順 的子孫三百二十八名；
NEH|7|23|比賽 的子孫三百二十四名；
NEH|7|24|哈拉 的子孫一百一十二名；
NEH|7|25|基遍 人九十五名；
NEH|7|26|伯利恆 人和 尼陀法 人共一百八十八名；
NEH|7|27|亞拿突 人一百二十八名；
NEH|7|28|伯‧亞斯瑪弗 人四十二名；
NEH|7|29|基列‧耶琳 人、 基非拉 人、 比錄 人共七百四十三名；
NEH|7|30|拉瑪 人和 迦巴 人共六百二十一名；
NEH|7|31|默瑪 人一百二十二名；
NEH|7|32|伯特利 人和 艾 人共一百二十三名；
NEH|7|33|別的 尼波 人五十二名；
NEH|7|34|另一個 以攔 子孫一千二百五十四名；
NEH|7|35|哈琳 的子孫三百二十名；
NEH|7|36|耶利哥 人三百四十五名；
NEH|7|37|羅德 人、 哈第 人、 阿挪 人共七百二十一名；
NEH|7|38|西拿 人三千九百三十名。
NEH|7|39|祭司： 耶書亞 家， 耶大雅 的子孫九百七十三名；
NEH|7|40|音麥 的子孫一千零五十二名；
NEH|7|41|巴施戶珥 的子孫一千二百四十七名；
NEH|7|42|哈琳 的子孫一千零一十七名。
NEH|7|43|利未 人： 何達威 的後裔，就是 耶書亞 和 甲篾 的子孫七十四名。
NEH|7|44|歌唱的： 亞薩 的子孫一百四十八名。
NEH|7|45|門口的守衛： 沙龍 的子孫、 亞特 的子孫、 達們 的子孫、 亞谷 的子孫、 哈底大 的子孫、 朔拜 的子孫，共一百三十八名。
NEH|7|46|殿役： 西哈 的子孫、 哈蘇巴 的子孫、 答巴俄 的子孫、
NEH|7|47|基綠 的子孫、 西亞 的子孫、 巴頓 的子孫、
NEH|7|48|利巴拿 的子孫、 哈迦巴 的子孫、 薩買 的子孫、
NEH|7|49|哈難 的子孫、 吉德 的子孫、 迦哈 的子孫、
NEH|7|50|利亞雅 的子孫、 利汛 的子孫、 尼哥大 的子孫、
NEH|7|51|迦散 的子孫、 烏撒 的子孫、 巴西亞 的子孫、
NEH|7|52|比賽 的子孫、 米烏寧 的子孫、 尼普心 的子孫、
NEH|7|53|巴卜 的子孫、 哈古巴 的子孫、 哈忽 的子孫、
NEH|7|54|巴洗律 的子孫、 米希大 的子孫、 哈沙 的子孫、
NEH|7|55|巴柯 的子孫、 西西拉 的子孫、 答瑪 的子孫、
NEH|7|56|尼細亞 的子孫、 哈提法 的子孫。
NEH|7|57|所羅門 僕人的後裔： 瑣太 的子孫、 瑣斐列 的子孫、 比路大 的子孫、
NEH|7|58|雅拉 的子孫、 達昆 的子孫、 吉德 的子孫、
NEH|7|59|示法提雅 的子孫、 哈替 的子孫、 玻黑列‧哈斯巴音 的子孫、 亞們 的子孫。
NEH|7|60|殿役和 所羅門 僕人的後裔共三百九十二名。
NEH|7|61|從 特‧米拉 、 特‧哈薩 、 基綠 、 亞頓 、 音麥 上來，不能證明他們的父系家族和後裔是否屬 以色列 的如下：
NEH|7|62|第萊雅 的子孫、 多比雅 的子孫、 尼哥大 的子孫，共六百四十二名。
NEH|7|63|祭司中， 哈巴雅 的子孫、 哈哥斯 的子孫、 巴西萊 的子孫， 巴西萊 因為娶了 基列 人 巴西萊 的女兒為妻，所以就以此為名。
NEH|7|64|這些人在族譜之中尋查自己的譜系，卻尋不著，因此算為不潔，不得作祭司。
NEH|7|65|省長對他們說，不可吃至聖的物，直到有會用烏陵和土明的祭司興起來。
NEH|7|66|全會眾共有四萬二千三百六十名。
NEH|7|67|此外，還有他們的僕婢七千三百三十七名，又有歌唱的男女二百四十五名。
NEH|7|68|他們有七百三十六匹馬，二百四十五匹騾子，
NEH|7|69|四百三十五匹駱駝，六千七百二十匹驢。
NEH|7|70|有些族長為工程捐助。省長捐入庫房中的有一千達利克 金子，五十個碗，五百三十件祭司的禮服。
NEH|7|71|有些族長捐入工程的庫房，有二萬達利克金子，二千二百彌那銀子。
NEH|7|72|其餘百姓所捐的有二萬達利克金子，二千彌那銀子，六十七件祭司的禮服。
NEH|7|73|於是祭司、 利未 人、門口的守衛、歌唱的、百姓中的一些人、殿役，並 以色列 眾人，都住在自己的城裏。 到了七月， 以色列 人住在自己的城裏。
NEH|8|1|那時，眾百姓如同一人聚集在 水門 前的廣場，請 以斯拉 文士將耶和華吩咐 以色列 的 摩西 的律法書帶來。
NEH|8|2|七月初一， 以斯拉 祭司將律法書帶到聽了能明白的男女會眾面前。
NEH|8|3|他在 水門 前的廣場，從清早到中午，在男女和能明白的人面前讀這律法書，眾百姓都側耳而聽。
NEH|8|4|以斯拉 文士站在為這事特製的木臺上。站在他旁邊的有 瑪他提雅 、 示瑪 、 亞奈雅 、 烏利亞 和 希勒家 ；站在他右邊的有 瑪西雅 ；站在他左邊的有 毗大雅 、 米沙利 、 瑪基雅 、 哈順 、 哈拔大拿 、 撒迦利亞 和 米書蘭 。
NEH|8|5|以斯拉 站在上面，在眾百姓眼前展開這書。他一展開，眾百姓都站起來。
NEH|8|6|以斯拉 稱頌耶和華至大的上帝，眾百姓都舉手應聲說：「阿們！阿們！」他們低頭，俯伏在地，敬拜耶和華。
NEH|8|7|耶書亞 、 巴尼 、 示利比 、 雅憫 、 亞谷 、 沙比太 、 荷第雅 、 瑪西雅 、 基利他 、 亞撒利雅 、 約撒拔 、 哈難 、 毗萊雅 和 利未 人使百姓明白律法；百姓都站在自己的地方。
NEH|8|8|他們清清楚楚地念上帝的律法書，講明意思，使百姓明白所念的。
NEH|8|9|尼希米 省長、 以斯拉 祭司文士，和教導百姓的 利未 人對眾百姓說：「今日是耶和華－你們上帝的聖日，不要悲哀，也不要哭泣。」這是因為眾百姓聽見律法書上的話都哭了。
NEH|8|10|尼希米 對他們說：「你們去吃肥美的，喝甘甜的，有不能預備的就分給他，因為今日是我們主的聖日。你們不要憂愁，因靠耶和華而得的喜樂是你們的力量。」
NEH|8|11|於是 利未 人叫眾百姓安靜，說：「安靜，因今日是聖日，不要憂愁。」
NEH|8|12|眾百姓去吃喝，也分給別人，都大大喜樂，因為他們明白所教導他們的話。
NEH|8|13|次日，眾百姓的族長、祭司和 利未 人都聚集到 以斯拉 文士那裏，要明白律法書上的話。
NEH|8|14|他們發現律法書上寫著，耶和華藉 摩西 吩咐 以色列 人要在七月的節期中住在棚裏，
NEH|8|15|並要在各城和 耶路撒冷 傳揚宣告說：「你們當出去，上山，把橄欖樹、野橄欖樹、番石榴樹、棕樹和各樣茂密樹的枝子取來，照著所寫的搭棚。」
NEH|8|16|於是百姓出去，取了樹枝來，各人在自己的房頂上、院子裏、上帝殿的院內、 水門 的廣場和 以法蓮門 的廣場搭棚。
NEH|8|17|從被擄之地歸回的全會眾就搭棚，住在棚裏。從 嫩 的兒子 約書亞 的時候直到這日， 以色列 人沒有這樣行。他們都大大喜樂。
NEH|8|18|從第一天直到末一天， 以斯拉 天天朗讀上帝的律法書。他們守節七日，第八日照例有嚴肅會。
NEH|9|1|這月二十四日， 以色列 人聚集禁食，他們披麻蒙灰。
NEH|9|2|以色列 的後裔與所有的外邦人分別出來，站著承認自己的罪和祖先的罪孽。
NEH|9|3|那日的四分之一，他們站在自己的地方念耶和華－他們上帝的律法書，又在那日的四分之一認罪，敬拜耶和華－他們的上帝。
NEH|9|4|耶書亞 、 巴尼 、 甲篾 、 示巴尼 、 布尼 、 示利比 、 巴尼 、 基拿尼 站在 利未 人的臺階上，大聲哀求耶和華－他們的上帝。
NEH|9|5|利未 人 耶書亞 、 甲篾 、 巴尼 、 哈沙尼 、 示利比 、 荷第雅 、 示巴尼 、 毗他希雅 說：「起來，稱頌耶和華－你們的上帝，永世無盡：『你榮耀之名是應當稱頌的，超乎一切稱頌和讚美。
NEH|9|6|「『你，惟獨你是耶和華！你造了天和天上的天，以及天上的萬象，地和地上的萬物，海和海中所有的；一切的生命全都是你賞賜的。天軍都敬拜你。
NEH|9|7|你是耶和華上帝，曾揀選 亞伯蘭 ，領他出 迦勒底 的 吾珥 ，給他改名叫 亞伯拉罕 。
NEH|9|8|你發現他在你面前心裏忠誠，就與他立約，要把 迦南 人、 赫 人、 亞摩利 人、 比利洗 人、 耶布斯 人、 革迦撒 人之地賜給他的後裔，並且你也實現了你的話，因為你是公義的。
NEH|9|9|「『你曾看見我們祖先在 埃及 所受的困苦，垂聽他們在 紅海 邊的哀求，
NEH|9|10|施行神蹟奇事在法老和他所有臣僕，以及他國中眾百姓身上，因為你知道他們向我們祖先行事狂傲。你也得了名聲，正如今日一樣。
NEH|9|11|你在我們祖先面前把海分開，使他們走過海中乾地，將追趕他們的人拋在深海，如石頭拋在大水中。
NEH|9|12|白晝你用雲柱引導他們，黑夜你用火柱照亮他們當行的路。
NEH|9|13|你降臨在 西奈山 ，從天上與他們說話，賜給他們正直的典章、真實的律法、美好的律例與誡命，
NEH|9|14|又使他們知道你的聖安息日，並藉你僕人 摩西 傳給他們誡命、律例、律法。
NEH|9|15|你從天上賜下糧食給他們充飢，使水從磐石流出給他們解渴。你吩咐他們進去，得你起誓應許要賜給他們的地。
NEH|9|16|「『但我們的祖先行事狂傲，硬著頸項不聽從你的誡命。
NEH|9|17|他們不肯順從，也不記念你在他們中間所行的奇事，竟硬著頸項，居心悖逆，自立領袖，要回 埃及 他們為奴之地 。但你是樂意饒恕人，有恩惠，有憐憫，不輕易發怒，有豐盛慈愛的上帝，並沒有丟棄他們。
NEH|9|18|他們雖然為自己鑄了一頭牛犢，說，這就是領你出 埃及 的神明，因而犯了褻瀆的大罪，
NEH|9|19|你還是有豐富的憐憫，不把他們丟棄在曠野。白晝，雲柱不離開他們，仍引導他們行路；黑夜，火柱仍照亮他們當行的路。
NEH|9|20|你賜下你良善的靈教導他們，沒有收回嗎哪不給他們吃，仍賜水給他們解渴。
NEH|9|21|在曠野四十年，你養育他們，他們一無所缺，衣服沒有穿破，腳也沒有腫。
NEH|9|22|你將列國和諸民族交給他們，把那些角落分給他們，他們就得了 西宏 之地，就是 希實本 王之地，和 巴珊 王 噩 之地。
NEH|9|23|你使他們的子孫多如天上的星，帶他們到你對他們祖先說要進去得為業之地。
NEH|9|24|這樣，這些子孫進去得了那地。你在他們面前制伏那地的居民 迦南 人，把 迦南 人和他們的君王，以及那地的民族，都交在他們手裏，讓他們任意處置。
NEH|9|25|他們得了堅固的城鎮、肥沃的土地，取了裝滿各樣美物的房屋、挖成的水井、葡萄園、橄欖園，以及許多果樹。他們就吃了，而且飽足，身體肥胖，因你的大恩活得快樂。
NEH|9|26|「『然而，他們不順從，竟背叛你，將你的律法丟在背後，又殺害那些勸他們回轉歸向你的眾先知，犯了褻瀆的大罪。
NEH|9|27|所以你將他們交在敵人的手中，敵人就折磨他們。他們遭難的時候哀求你，你就從天上垂聽，照你豐富的憐憫賜給他們拯救者，救他們脫離敵人的手。
NEH|9|28|但他們得享太平之後，又在你面前行惡，所以你丟棄他們，交在仇敵的手中，仇敵就轄制他們；然而他們轉回哀求你，你就從天上垂聽，屢次照你的憐憫拯救他們，
NEH|9|29|你警戒他們，要使他們歸順你的律法。他們卻行事狂傲，不聽從你的誡命，干犯你的典章，人若遵行就必因此存活。他們頑梗地扭轉肩頭，硬著頸項，不肯聽從。
NEH|9|30|但你多年寬容他們，又以你的靈藉眾先知勸戒他們，他們仍不側耳而聽，所以你將他們交在列邦民族的手中。
NEH|9|31|然而因你豐富的憐憫，你不全然滅絕他們，也不丟棄他們，因為你是有恩惠、有憐憫的上帝。
NEH|9|32|「『現在，我們的上帝啊，你是至大、至能、至可畏、守約施慈愛的上帝；我們的君王、官長、祭司、先知、祖先和你的眾百姓，從 亞述 諸王的時候直到今日所遭遇的一切苦難，求你不要看為小事。
NEH|9|33|在一切臨到我們的事上，你是公義的，因為你所行的是信實，我們所做的是邪惡。
NEH|9|34|我們的君王、官長、祭司、祖先都不遵守你的律法，不聽從你的誡命和你警戒他們的話。
NEH|9|35|他們在本國領受你大恩的時候，在你所賜給他們這廣大肥沃之地不事奉你，也不轉離他們的惡行。
NEH|9|36|看哪，我們今日成了奴僕！你賜給我們祖先享受土產和美物的地，看哪，我們在這地上竟作了奴僕！
NEH|9|37|這地許多的出產都歸了諸王，就是你因我們的罪派來轄制我們的。他們任意轄制我們的身體和牲畜，我們遭了大難。』」
NEH|9|38|因這一切，我們立確實的約，寫在冊上。我們的領袖、 利未 人和祭司都用了印。
NEH|10|1|用印的是 哈迦利亞 的兒子 尼希米 省長、 西底家 ；
NEH|10|2|還有 西萊雅 、 亞撒利雅 、 耶利米 、
NEH|10|3|巴施戶珥 、 亞瑪利雅 、 瑪基雅 、
NEH|10|4|哈突 、 示巴尼 、 瑪鹿 、
NEH|10|5|哈琳 、 米利末 、 俄巴底亞 、
NEH|10|6|但以理 、 近頓 、 巴錄 、
NEH|10|7|米書蘭 、 亞比雅 、 米雅民 、
NEH|10|8|瑪西亞 、 璧該 、 示瑪雅 等祭司；
NEH|10|9|又有 利未 人 亞散尼 的兒子 耶書亞 、 希拿達 的子孫 賓內 、 甲篾 ，
NEH|10|10|他們的弟兄 示巴尼 、 荷第雅 、 基利他 、 毗萊雅 、 哈難 、
NEH|10|11|米迦 、 利合 、 哈沙比雅 、
NEH|10|12|撒刻 、 示利比 、 示巴尼 、
NEH|10|13|荷第雅 、 巴尼 、 比尼努 ；
NEH|10|14|還有百姓中的領袖 巴錄 、 巴哈‧摩押 、 以攔 、 薩土 、 巴尼 、
NEH|10|15|布尼 、 押甲 、 比拜 、
NEH|10|16|亞多尼雅 、 比革瓦伊 、 亞丁 、
NEH|10|17|亞特 、 希西家 、 押朔 、
NEH|10|18|荷第雅 、 哈順 、 比賽 、
NEH|10|19|哈拉 、 亞拿突 、 尼拜 、
NEH|10|20|抹比押 、 米書蘭 、 希悉 、
NEH|10|21|米示薩別 、 撒督 、 押杜亞 、
NEH|10|22|毗拉提 、 哈難 、 亞奈雅 、
NEH|10|23|何細亞 、 哈拿尼雅 、 哈述 、
NEH|10|24|哈羅黑 、 毗利哈 、 朔百 、
NEH|10|25|利宏 、 哈沙拿 、 瑪西雅 、
NEH|10|26|亞希雅 、 哈難 、 亞難 、
NEH|10|27|瑪鹿 、 哈琳 、 巴拿 。
NEH|10|28|其餘的百姓、祭司、 利未 人、門口的守衛、歌唱的、殿役，所有與鄰邦民族分別出來、歸服上帝律法的，以及他們的妻子、兒女，凡有知識、能明白的，
NEH|10|29|都隨從他們貴族的弟兄發咒起誓，要遵行上帝藉他僕人 摩西 所賜的律法，謹守遵行耶和華－我們主的一切誡命、典章、律例。
NEH|10|30|我們不把我們的女兒嫁給這地的居民，也不為我們的兒子娶他們的女兒。
NEH|10|31|這地的民族若在安息日，或甚麼聖日，帶了貨物或糧食來賣，我們必不買。每逢第七年必不耕種，凡欠我們債的必不追討。
NEH|10|32|我們又為自己定例，每年各人捐獻三分之一舍客勒，作為我們上帝殿之用：
NEH|10|33|為供餅、常獻的素祭和燔祭，安息日、初一、節期所獻的祭和聖物， 以色列 的贖罪祭，以及我們上帝殿裏一切工作之用。
NEH|10|34|我們的祭司、 利未 人和百姓都抽籤，每年按父家定期將奉獻的木柴帶到我們上帝的殿裏，照著律法上所寫的，燒在耶和華－我們上帝的壇上。
NEH|10|35|每年我們又將地上初熟的土產和各樣樹上初熟的果子，都奉到耶和華的殿裏。
NEH|10|36|我們又照律法上所寫的，將我們頭胎的兒子和首生的牛羊都奉到我們上帝的殿，交給在上帝殿裏供職的祭司；
NEH|10|37|並將初熟麥子所磨的麵和舉祭、各樣樹上的果子、新酒與新油奉給祭司，收在我們上帝殿的庫房裏，又把我們土地所產的十分之一奉給 利未 人，因 利未 人在我們一切城鎮的土產中當取十分之一。
NEH|10|38|利未 人取十分之一的時候， 亞倫 的子孫中當有一個祭司與 利未 人同在。 利未 人也當從十分之一中取十分之一，奉到我們上帝的殿，收在庫房的倉裏。
NEH|10|39|因 以色列 人和 利未 人要把禮物，就是五穀、新酒和新油，帶到收存聖所器皿的倉裏，供職的祭司、門口的守衛、歌唱的都在那裏。我們絕不會不顧我們上帝的殿。
NEH|11|1|百姓的領袖住在 耶路撒冷 。其餘的百姓抽籤，每十人中選一人來住在聖城 耶路撒冷 ，另外九人住在別的城鎮。
NEH|11|2|凡甘心樂意住在 耶路撒冷 的，百姓都為他們祝福。
NEH|11|3|以色列 人、祭司、 利未 人、殿役和 所羅門 僕人的後裔都住在 猶大 的城鎮，各在自己城內的地業中。本省的領袖住在 耶路撒冷 的如下：
NEH|11|4|住在 耶路撒冷 的有一些 猶大 人和 便雅憫 人。 猶大 人中有 法勒斯 的子孫 亞他雅 ； 亞他雅 是 烏西雅 的兒子， 烏西雅 是 撒迦利雅 的兒子， 撒迦利雅 是 亞瑪利雅 的兒子， 亞瑪利雅 是 示法提雅 的兒子， 示法提雅 是 瑪勒列 的兒子；
NEH|11|5|又有 瑪西雅 ； 瑪西雅 是 巴錄 的兒子， 巴錄 是 谷‧何西 的兒子， 谷‧何西 是 哈賽雅 的兒子， 哈賽雅 是 亞大雅 的兒子， 亞大雅 是 約雅立 的兒子， 約雅立 是 撒迦利雅 的兒子， 撒迦利雅 是 示羅尼 的兒子；
NEH|11|6|住在 耶路撒冷 所有 法勒斯 的子孫共四百六十八名，都是勇士。
NEH|11|7|便雅憫 人中有 撒路 ； 撒路 是 米書蘭 的兒子， 米書蘭 是 約葉 的兒子， 約葉 是 毗大雅 的兒子， 毗大雅 是 哥賴雅 的兒子， 哥賴雅 是 瑪西雅 的兒子， 瑪西雅 是 以鐵 的兒子， 以鐵 是 耶篩亞 的兒子；
NEH|11|8|其次有 迦拜 、 撒來 ，共九百二十八名。
NEH|11|9|細基利 的兒子 約珥 是他們的長官； 哈西努亞 的兒子 猶大 是 耶路撒冷 的副長官。
NEH|11|10|祭司中有 約雅立 的兒子 耶大雅 ，又有 雅斤 ，
NEH|11|11|還有管理上帝殿的 西萊雅 ； 西萊雅 是 希勒家 的兒子， 希勒家 是 米書蘭 的兒子， 米書蘭 是 撒督 的兒子， 撒督 是 米拉約 的兒子， 米拉約 是 亞希突 的兒子；
NEH|11|12|還有他們的弟兄在殿裏供職的，共八百二十二名；又有 亞大雅 ； 亞大雅 是 耶羅罕 的兒子， 耶羅罕 是 毗拉利 的兒子， 毗拉利 是 暗洗 的兒子， 暗洗 是 撒迦利亞 的兒子， 撒迦利亞 是 巴施戶珥 的兒子， 巴施戶珥 是 瑪基雅 的兒子；
NEH|11|13|還有他的弟兄作族長的，共二百四十二名；又有 亞瑪帥 ； 亞瑪帥 是 亞薩列 的兒子， 亞薩列 是 亞哈賽 的兒子， 亞哈賽 是 米實利末 的兒子， 米實利末 是 音麥 的兒子；
NEH|11|14|還有他們的弟兄，大能的勇士共一百二十八名； 哈基多琳 的兒子 撒巴第業 是他們的長官。
NEH|11|15|利未 人中有 示瑪雅 ； 示瑪雅 是 哈述 的兒子， 哈述 是 押利甘 的兒子， 押利甘 是 哈沙比雅 的兒子， 哈沙比雅 是 布尼 的兒子；
NEH|11|16|又有 利未 人的族長 沙比太 和 約撒拔 管理上帝殿外面的事務；
NEH|11|17|祈禱的時候， 瑪他尼 是主禮，開始稱謝； 瑪他尼 是 米迦 的兒子， 米迦 是 撒底 的兒子， 撒底 是 亞薩 的兒子；又有 瑪他尼 弟兄中的 八布迦 為副；還有 押大 ； 押大 是 沙母亞 的兒子， 沙母亞 是 加拉 的兒子， 加拉 是 耶杜頓 的兒子；
NEH|11|18|在聖城所有的 利未 人共二百八十四名。
NEH|11|19|門口的守衛是 亞谷 和 達們 ，以及他們的弟兄，看守各門，共一百七十二名。
NEH|11|20|其餘的 以色列 人、祭司、 利未 人都住在 猶大 一切的城鎮，各在自己的地業中。
NEH|11|21|殿役卻住在 俄斐勒 ； 西哈 和 基斯帕 管理他們。
NEH|11|22|在 耶路撒冷 ， 利未 人的長官，管理上帝殿事務的是歌唱者 亞薩 的子孫 烏西 ； 烏西 是 巴尼 的兒子， 巴尼 是 哈沙比雅 的兒子， 哈沙比雅 是 瑪他尼 的兒子， 瑪他尼 是 米迦 的兒子。
NEH|11|23|王為歌唱者下命令，確定他們每日當辦的事 。
NEH|11|24|猶大 的兒子 謝拉 的子孫， 米示薩別 的兒子 毗他希雅 輔助王辦理百姓一切的事。
NEH|11|25|至於村莊和所屬的田地，有 猶大 人住在 基列‧亞巴 和所屬的鄉鎮 、 底本 和所屬的鄉鎮、 葉甲薛 和所屬的村莊、
NEH|11|26|耶書亞 、 摩拉大 、 伯‧帕列 、
NEH|11|27|哈薩‧書亞 、 別是巴 和所屬的鄉鎮、
NEH|11|28|洗革拉 、 米哥拿 和所屬的鄉鎮、
NEH|11|29|隱‧臨門 、 瑣拉 、 耶末 、
NEH|11|30|撒挪亞 、 亞杜蘭 和屬它們的村莊、 拉吉 和所屬的田地、 亞西加 和所屬的鄉鎮；他們所住的地方是從 別是巴 直到 欣嫩谷 。
NEH|11|31|便雅憫 人從 迦巴 起，住在 密抹 、 亞雅 、 伯特利 和所屬的鄉鎮、
NEH|11|32|亞拿突 、 挪伯 、 亞難雅 、
NEH|11|33|夏瑣 、 拉瑪 、 基他音 、
NEH|11|34|哈第 、 洗編 、 尼八拉 、
NEH|11|35|羅德 、 阿挪 、 革‧夏納欣 。
NEH|11|36|在 猶大 地區的 利未 人中，有些已歸屬 便雅憫 。
NEH|12|1|這些是同 撒拉鐵 的兒子 所羅巴伯 以及 耶書亞 一起上來的祭司和 利未 人： 西萊雅 、 耶利米 、 以斯拉 、
NEH|12|2|亞瑪利雅 、 瑪鹿 、 哈突 、
NEH|12|3|示迦尼 、 利宏 、 米利末 、
NEH|12|4|易多 、 近頓 、 亞比雅 、
NEH|12|5|米雅民 、 瑪底雅 、 璧迦 、
NEH|12|6|示瑪雅 、 約雅立 、 耶大雅 、
NEH|12|7|撒路 、 亞木 、 希勒家 、 耶大雅 ；這些人在 耶書亞 的時代作祭司和他們弟兄的領袖。
NEH|12|8|利未 人有 耶書亞 、 賓內 、 甲篾 、 示利比 、 猶大 、 瑪他尼 ； 瑪他尼 和他的弟兄負責讚美詩歌。
NEH|12|9|他們的弟兄 八布迦 和 烏尼 按照班次站在他們的對面。
NEH|12|10|耶書亞 生 約雅金 ， 約雅金 生 以利亞實 ， 以利亞實 生 耶何耶大 ，
NEH|12|11|耶何耶大 生 約拿單 ， 約拿單 生 押杜亞 。
NEH|12|12|在 約雅金 的時代，祭司作族長的， 西萊雅 族有 米拉雅 ， 耶利米 族有 哈拿尼雅 ，
NEH|12|13|以斯拉 族有 米書蘭 ， 亞瑪利雅 族有 約哈難 ，
NEH|12|14|米利古 族有 約拿單 ， 示巴尼 族有 約瑟 ，
NEH|12|15|哈琳 族有 押拿 ， 米拉約 族有 希勒愷 ，
NEH|12|16|易多 族有 撒迦利亞 ， 近頓 族有 米書蘭 ，
NEH|12|17|亞比雅 族有 細基利 ， 米拿民 族， 摩亞底 族有 毗勒太 ，
NEH|12|18|璧迦 族有 沙母亞 ， 示瑪雅 族有 約拿單 ，
NEH|12|19|約雅立 族有 瑪特乃 ， 耶大雅 族有 烏西 ，
NEH|12|20|撒來 族有 加萊 ， 亞木 族有 希伯 ，
NEH|12|21|希勒家 族有 哈沙比雅 ， 耶大雅 族有 拿坦業 。
NEH|12|22|在 以利亞實 、 耶何耶大 、 約哈難 、 押杜亞 的時代， 利未 人的族長都記在冊上，祭司也一樣，直到 波斯 王 大流士 在位的時候。
NEH|12|23|利未 人作族長的記在史籍上，一直記到 以利亞實 的兒子 約哈難 的時代。
NEH|12|24|利未 人的族長是 哈沙比雅 、 示利比 、 甲篾 的兒子 耶書亞 ，他們的弟兄站在他們的對面，照神人 大衛 的命令按著班次讚美稱謝。
NEH|12|25|瑪他尼 、 八布迦 、 俄巴底亞 、 米書蘭 、 達們 、 亞谷 是門口的守衛，在庫房的門口站崗。
NEH|12|26|這些人都在 約撒達 的孫子， 耶書亞 的兒子 約雅金 和 尼希米 省長，以及 以斯拉 祭司文士的時代供職。
NEH|12|27|為 耶路撒冷 城牆行奉獻禮的時候，眾人把各處的 利未 人召到 耶路撒冷 ，要以稱謝、歌唱、敲鈸、鼓瑟、彈琴，喜樂地行奉獻禮。
NEH|12|28|歌唱的人從 耶路撒冷 的周圍聚集，從 尼陀法 人的村莊、
NEH|12|29|伯‧吉甲 ，以及 迦巴 和 亞斯瑪弗 的田地而來；因為歌唱的人在 耶路撒冷 四圍為自己建立了村莊。
NEH|12|30|祭司和 利未 人就潔淨自己，也潔淨百姓，以及城門和城牆。
NEH|12|31|我帶 猶大 的領袖上城牆，把稱謝的人分為兩大隊，在城牆上往右邊的 糞廠門 行進，
NEH|12|32|在他們後面行進的有 何沙雅 與 猶大 一半的領袖，
NEH|12|33|又有 亞撒利雅 、 以斯拉 、 米書蘭 、
NEH|12|34|猶大 、 便雅憫 、 示瑪雅 、 耶利米 。
NEH|12|35|還有祭司的子孫，吹號的有 撒迦利亞 ； 撒迦利亞 是 約拿單 的兒子， 約拿單 是 示瑪雅 的兒子， 示瑪雅 是 瑪他尼 的兒子， 瑪他尼 是 米該亞 的兒子， 米該亞 是 撒刻 的兒子， 撒刻 是 亞薩 的兒子；
NEH|12|36|又有 撒迦利亞 的弟兄 示瑪雅 、 亞撒利 、 米拉萊 、 基拉萊 、 瑪艾 、 拿坦業 、 猶大 、 哈拿尼 ，各拿著神人 大衛 的樂器，由 以斯拉 文士在前面引領。
NEH|12|37|他們經過 泉門 往前，登 大衛城 的臺階，上城牆的斜坡，從 大衛 宮殿之上，直到朝東的 水門 。
NEH|12|38|第二隊稱謝的人要往反方向而行。我和一半的百姓在城牆上跟隨他們，從 爐樓 之上，直到 寬牆 ；
NEH|12|39|又過了 以法蓮門 、 古門 、 魚門 、 哈楠業樓 、 哈米亞樓 ，直到 羊門 ，就在 護衛門 站住。
NEH|12|40|於是，這兩隊稱謝的人連同我和一半跟隨我的官長，站在上帝的殿裏。
NEH|12|41|還有 以利亞金 、 瑪西雅 、 米拿民 、 米該亞 、 以利約乃 、 撒迦利亞 、 哈楠尼亞 等吹號的祭司；
NEH|12|42|又有 瑪西雅 、 示瑪雅 、 以利亞撒 、 烏西 、 約哈難 、 瑪基雅 、 以攔 和 以謝 。歌唱的大聲唱歌，有 伊斯拉希雅 作指揮。
NEH|12|43|那日，眾人獻上豐盛的祭物，並且歡樂，因為上帝使他們大大歡樂，連婦女帶孩童也都歡樂，甚至從遠處都可聽到 耶路撒冷 的歡聲。
NEH|12|44|當日，有些人受派管理庫房，把舉祭、初熟之物，和所取的十一奉獻，按各城的田地，照律法所定，歸給祭司和 利未 人的份，都收在庫房裏。 猶大 人因祭司和 利未 人供職就歡樂。
NEH|12|45|祭司和 利未 人遵守上帝所吩咐的，守潔淨禮。歌唱的和門口的守衛照著 大衛 和他兒子 所羅門 的命令也如此行。
NEH|12|46|古時，在 大衛 和 亞薩 的日子，有歌唱者的指揮，也有讚美稱謝上帝的詩歌。
NEH|12|47|在 所羅巴伯 和 尼希米 的時代， 以色列 眾人把歌唱者和門口的守衛每日當得的份供給他們，又把給 利未 人的分別出來； 利未 人又把給 亞倫 子孫的分別出來。
NEH|13|1|在那日，百姓聽到人朗讀 摩西 的律法書，發現書上寫著， 亞捫 人和 摩押 人永不可入上帝的會；
NEH|13|2|因為他們沒有拿食物和水來迎接 以色列 人，卻雇了 巴蘭 詛咒他們，但我們的上帝使那詛咒變為祝福。
NEH|13|3|以色列 人聽見這律法，就與所有不同族群的人分別出來。
NEH|13|4|在這之前，與 多比雅 結親的 以利亞實 祭司，受派管理我們上帝殿中的庫房，
NEH|13|5|為 多比雅 預備了一間大屋子，就是從前收存素祭、乳香、器皿，和照例供給 利未 人、歌唱者、門口守衛的五穀、新酒和新油的十分之一，以及歸祭司之舉祭的屋子。
NEH|13|6|當這一切事發生的時候，我不在 耶路撒冷 ，因為 巴比倫 王 亞達薛西 三十二年，我回到王那裏。過了多日，我又向王告假。
NEH|13|7|我來到 耶路撒冷 ，才知道 以利亞實 為 多比雅 所做、在上帝殿的院內為他預備屋子的那件惡事。
NEH|13|8|我非常憤怒，就把 多比雅 的一切家具都從屋子裏拋出去。
NEH|13|9|我又吩咐人潔淨這屋子，然後將上帝殿的器皿、素祭和乳香搬回那裏。
NEH|13|10|我發現 利未 人當得的份無人供給他們，甚至供職的 利未 人與歌唱的都各奔回自己的田地去了。
NEH|13|11|我就斥責官長說：「你們為何不顧上帝的殿呢？」於是我召集 利未 人，使他們在自己的崗位上供職。
NEH|13|12|猶大 眾人就把五穀、新酒和新油的十分之一送入庫房。
NEH|13|13|我派 示利米雅 祭司、 撒督 文士和 利未 人 毗大雅 作司庫管理庫房，副手是 哈難 ； 哈難 是 撒刻 的兒子， 撒刻 是 瑪他尼 的兒子；這些人都是忠實的，他們的職務是分派他們弟兄所當得的份。
NEH|13|14|我的上帝啊，求你因這事記念我，不要塗去我為上帝的殿與其中的禮儀所獻的忠心。
NEH|13|15|那些日子，我在 猶大 見有人在安息日踹醡酒池，搬運禾捆馱在驢上，又把酒、葡萄、無花果和各樣的擔子在安息日扛入 耶路撒冷 ，我就在他們賣食物的那日警戒他們。
NEH|13|16|有一些住在城裏的 推羅 人也把魚和各樣貨物運進來，甚至在 耶路撒冷 ，在安息日賣給 猶大 人。
NEH|13|17|我就斥責 猶大 的貴族，對他們說：「你們怎麼會做這惡事干犯安息日呢！
NEH|13|18|你們祖先豈不是這樣做，以致我們的上帝使一切災禍臨到我們和這城嗎？你們竟干犯安息日，使憤怒越發臨到 以色列 ！」
NEH|13|19|安息日前一日黃昏的時候，我吩咐人把 耶路撒冷 城門鎖上；我又吩咐，不過安息日不准開門。我也派幾個僕人在城門口站崗，免得有人在安息日挑擔子進城。
NEH|13|20|於是商人和販賣各樣貨物的人，有一兩次在 耶路撒冷 城外過夜。
NEH|13|21|我警告他們說：「你們為何在城牆前過夜呢？若再這樣，我必下手辦你們。」從此以後，他們在安息日就不再來了。
NEH|13|22|我吩咐 利未 人潔淨自己來守城門，使安息日分別為聖。我的上帝啊，求你因這事記念我，照你豐盛的慈愛憐憫我。
NEH|13|23|那些日子，我又看見 猶太 人娶了 亞實突 、 亞捫 和 摩押 的女子為妻。
NEH|13|24|他們的兒女，一半說 亞實突 話，或其他種族的方言，不會說 猶大 話。
NEH|13|25|我就斥責他們，詛咒他們，打了他們幾個人，拔下他們的鬍鬚，叫他們指著上帝起誓：「你們不可把自己的女兒嫁給外邦人的兒子，也不可為自己和兒子娶他們的女兒。
NEH|13|26|以色列 王 所羅門 不也在這樣的事上犯罪嗎？在許多國家中並沒有一位王像他，蒙他上帝喜愛，上帝立他作王治理全 以色列 。然而，連他也被外邦女子引誘犯罪。
NEH|13|27|我們豈能聽憑你們行這一切大惡，娶外邦女子干犯我們的上帝呢？」
NEH|13|28|以利亞實 大祭司的孫子， 耶何耶大 的一個兒子是 和倫 人 參巴拉 的女婿，我就把他從我這裏趕出去。
NEH|13|29|我的上帝啊，求你記得他們的罪，因為他們玷污了祭司的職分，違背祭司和 利未 人的約。
NEH|13|30|這樣，我潔淨他們，使他們脫離屬外邦人的一切；我又分派祭司和 利未 人的班次，使他們各盡其職，
NEH|13|31|按定期奉獻木柴和初熟的土產。我的上帝啊，求你記念我，施恩於我。
