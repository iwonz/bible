EXOD|1|1|These are the names of the sons of Israel who came to Egypt with Jacob, each with his household:
EXOD|1|2|Reuben, Simeon, Levi, and Judah,
EXOD|1|3|Issachar, Zebulun, and Benjamin,
EXOD|1|4|Dan and Naphtali, Gad and Asher.
EXOD|1|5|All the descendants of Jacob were seventy persons; Joseph was already in Egypt.
EXOD|1|6|Then Joseph died, and all his brothers and all that generation.
EXOD|1|7|But the people of Israel were fruitful and increased greatly; they multiplied and grew exceedingly strong, so that the land was filled with them.
EXOD|1|8|Now there arose a new king over Egypt, who did not know Joseph.
EXOD|1|9|And he said to his people, "Behold, the people of Israel are too many and too mighty for us.
EXOD|1|10|Come, let us deal shrewdly with them, lest they multiply, and, if war breaks out, they join our enemies and fight against us and escape from the land."
EXOD|1|11|Therefore they set taskmasters over them to afflict them with heavy burdens. They built for Pharaoh store cities, Pithom and Raamses.
EXOD|1|12|But the more they were oppressed, the more they multiplied and the more they spread abroad. And the Egyptians were in dread of the people of Israel.
EXOD|1|13|So they ruthlessly made the people of Israel work as slaves
EXOD|1|14|and made their lives bitter with hard service, in mortar and brick, and in all kinds of work in the field. In all their work they ruthlessly made them work as slaves.
EXOD|1|15|Then the king of Egypt said to the Hebrew midwives, one of whom was named Shiphrah and the other Puah,
EXOD|1|16|"When you serve as midwife to the Hebrew women and see them on the birthstool, if it is a son, you shall kill him, but if it is a daughter, she shall live."
EXOD|1|17|But the midwives feared God and did not do as the king of Egypt commanded them, but let the male children live.
EXOD|1|18|So the king of Egypt called the midwives and said to them, "Why have you done this, and let the male children live?"
EXOD|1|19|The midwives said to Pharaoh, "Because the Hebrew women are not like the Egyptian women, for they are vigorous and give birth before the midwife comes to them."
EXOD|1|20|So God dealt well with the midwives. And the people multiplied and grew very strong.
EXOD|1|21|And because the midwives feared God, he gave them families.
EXOD|1|22|Then Pharaoh commanded all his people, "Every son that is born to the Hebrews you shall cast into the Nile, but you shall let every daughter live."
EXOD|2|1|Now a man from the house of Levi went and took as his wife a Levite woman.
EXOD|2|2|The woman conceived and bore a son, and when she saw that he was a fine child, she hid him three months.
EXOD|2|3|When she could hide him no longer, she took for him a basket made of bulrushes and daubed it with bitumen and pitch. She put the child in it and placed it among the reeds by the river bank.
EXOD|2|4|And his sister stood at a distance to know what would be done to him.
EXOD|2|5|Now the daughter of Pharaoh came down to bathe at the river, while her young women walked beside the river. She saw the basket among the reeds and sent her servant woman, and she took it.
EXOD|2|6|When she opened it, she saw the child, and behold, the baby was crying. She took pity on him and said, "This is one of the Hebrews' children."
EXOD|2|7|Then his sister said to Pharaoh's daughter, "Shall I go and call you a nurse from the Hebrew women to nurse the child for you?"
EXOD|2|8|And Pharaoh's daughter said to her, "Go." So the girl went and called the child's mother.
EXOD|2|9|And Pharaoh's daughter said to her, "Take this child away and nurse him for me, and I will give you your wages." So the woman took the child and nursed him.
EXOD|2|10|When the child grew up, she brought him to Pharaoh's daughter, and he became her son. She named him Moses, "Because," she said, "I drew him out of the water."
EXOD|2|11|One day, when Moses had grown up, he went out to his people and looked on their burdens, and he saw an Egyptian beating a Hebrew, one of his people.
EXOD|2|12|He looked this way and that, and seeing no one, he struck down the Egyptian and hid him in the sand.
EXOD|2|13|When he went out the next day, behold, two Hebrews were struggling together. And he said to the man in the wrong, "Why do you strike your companion?"
EXOD|2|14|He answered, "Who made you a prince and a judge over us? Do you mean to kill me as you killed the Egyptian?" Then Moses was afraid, and thought, "Surely the thing is known."
EXOD|2|15|When Pharaoh heard of it, he sought to kill Moses. But Moses fled from Pharaoh and stayed in the land of Midian. And he sat down by a well.
EXOD|2|16|Now the priest of Midian had seven daughters, and they came and drew water and filled the troughs to water their father's flock.
EXOD|2|17|The shepherds came and drove them away, but Moses stood up and saved them, and watered their flock.
EXOD|2|18|When they came home to their father Reuel, he said, "How is it that you have come home so soon today?"
EXOD|2|19|They said, "An Egyptian delivered us out of the hand of the shepherds and even drew water for us and watered the flock."
EXOD|2|20|He said to his daughters, "Then where is he? Why have you left the man? Call him, that he may eat bread."
EXOD|2|21|And Moses was content to dwell with the man, and he gave Moses his daughter Zipporah.
EXOD|2|22|She gave birth to a son, and he called his name Gershom, for he said, "I have been a sojourner in a foreign land."
EXOD|2|23|During those many days the king of Egypt died, and the people of Israel groaned because of their slavery and cried out for help. Their cry for rescue from slavery came up to God.
EXOD|2|24|And God heard their groaning, and God remembered his covenant with Abraham, with Isaac, and with Jacob.
EXOD|2|25|God saw the people of Israel- and God knew.
EXOD|3|1|Now Moses was keeping the flock of his father-in-law, Jethro, the priest of Midian, and he led his flock to the west side of the wilderness and came to Horeb, the mountain of God.
EXOD|3|2|And the angel of the LORD appeared to him in a flame of fire out of the midst of a bush. He looked, and behold, the bush was burning, yet it was not consumed.
EXOD|3|3|And Moses said, "I will turn aside to see this great sight, why the bush is not burned."
EXOD|3|4|When the LORD saw that he turned aside to see, God called to him out of the bush, "Moses, Moses!" And he said, "Here I am."
EXOD|3|5|Then he said, "Do not come near; take your sandals off your feet, for the place on which you are standing is holy ground."
EXOD|3|6|And he said, "I am the God of your father, the God of Abraham, the God of Isaac, and the God of Jacob." And Moses hid his face, for he was afraid to look at God.
EXOD|3|7|Then the LORD said, "I have surely seen the affliction of my people who are in Egypt and have heard their cry because of their taskmasters. I know their sufferings,
EXOD|3|8|and I have come down to deliver them out of the hand of the Egyptians and to bring them up out of that land to a good and broad land, a land flowing with milk and honey, to the place of the Canaanites, the Hittites, the Amorites, the Perizzites, the Hivites, and the Jebusites.
EXOD|3|9|And now, behold, the cry of the people of Israel has come to me, and I have also seen the oppression with which the Egyptians oppress them.
EXOD|3|10|Come, I will send you to Pharaoh that you may bring my people, the children of Israel, out of Egypt."
EXOD|3|11|But Moses said to God, "Who am I that I should go to Pharaoh and bring the children of Israel out of Egypt?"
EXOD|3|12|He said, "But I will be with you, and this shall be the sign for you, that I have sent you: when you have brought the people out of Egypt, you shall serve God on this mountain."
EXOD|3|13|Then Moses said to God, "If I come to the people of Israel and say to them, 'The God of your fathers has sent me to you,' and they ask me, 'What is his name?' what shall I say to them?"
EXOD|3|14|God said to Moses, "I AM WHO I AM." And he said, "Say this to the people of Israel, 'I AM has sent me to you.'"
EXOD|3|15|God also said to Moses, "Say this to the people of Israel, 'The LORD, the God of your fathers, the God of Abraham, the God of Isaac, and the God of Jacob, has sent me to you.' This is my name forever, and thus I am to be remembered throughout all generations.
EXOD|3|16|Go and gather the elders of Israel together and say to them, 'The LORD, the God of your fathers, the God of Abraham, of Isaac, and of Jacob, has appeared to me, saying, "I have observed you and what has been done to you in Egypt,
EXOD|3|17|and I promise that I will bring you up out of the affliction of Egypt to the land of the Canaanites, the Hittites, the Amorites, the Perizzites, the Hivites, and the Jebusites, a land flowing with milk and honey."'
EXOD|3|18|And they will listen to your voice, and you and the elders of Israel shall go to the king of Egypt and say to him, 'The LORD, the God of the Hebrews, has met with us; and now, please let us go a three days' journey into the wilderness, that we may sacrifice to the LORD our God.'
EXOD|3|19|But I know that the king of Egypt will not let you go unless compelled by a mighty hand.
EXOD|3|20|So I will stretch out my hand and strike Egypt with all the wonders that I will do in it; after that he will let you go.
EXOD|3|21|And I will give this people favor in the sight of the Egyptians; and when you go, you shall not go empty,
EXOD|3|22|but each woman shall ask of her neighbor, and any woman who lives in her house, for silver and gold jewelry, and for clothing. You shall put them on your sons and on your daughters. So you shall plunder the Egyptians."
EXOD|4|1|Then Moses answered, "But behold, they will not believe me or listen to my voice, for they will say, 'The LORD did not appear to you.'"
EXOD|4|2|The LORD said to him, "What is that in your hand?" He said, "A staff."
EXOD|4|3|And he said, "Throw it on the ground." So he threw it on the ground, and it became a serpent, and Moses ran from it.
EXOD|4|4|But the LORD said to Moses, "Put out your hand and catch it by the tail"- so he put out his hand and caught it, and it became a staff in his hand-
EXOD|4|5|"that they may believe that the LORD, the God of their fathers, the God of Abraham, the God of Isaac, and the God of Jacob, has appeared to you."
EXOD|4|6|Again, the LORD said to him, "Put your hand inside your cloak." And he put his hand inside his cloak, and when he took it out, behold, his hand was leprous like snow.
EXOD|4|7|Then God said, "Put your hand back inside your cloak." So he put his hand back inside his cloak, and when he took it out, behold, it was restored like the rest of his flesh.
EXOD|4|8|"If they will not believe you," God said, "or listen to the first sign, they may believe the latter sign.
EXOD|4|9|If they will not believe even these two signs or listen to your voice, you shall take some water from the Nile and pour it on the dry ground, and the water that you shall take from the Nile will become blood on the dry ground."
EXOD|4|10|But Moses said to the LORD, "Oh, my Lord, I am not eloquent, either in the past or since you have spoken to your servant, but I am slow of speech and of tongue."
EXOD|4|11|Then the LORD said to him, "Who has made man's mouth? Who makes him mute, or deaf, or seeing, or blind? Is it not I, the LORD?
EXOD|4|12|Now therefore go, and I will be with your mouth and teach you what you shall speak."
EXOD|4|13|But he said, "Oh, my Lord, please send someone else."
EXOD|4|14|Then the anger of the LORD was kindled against Moses and he said, "Is there not Aaron, your brother, the Levite? I know that he can speak well. Behold, he is coming out to meet you, and when he sees you, he will be glad in his heart.
EXOD|4|15|You shall speak to him and put the words in his mouth, and I will be with your mouth and with his mouth and will teach you both what to do.
EXOD|4|16|He shall speak for you to the people, and he shall be your mouth, and you shall be as God to him.
EXOD|4|17|And take in your hand this staff, with which you shall do the signs."
EXOD|4|18|Moses went back to Jethro his father-in-law and said to him, "Please let me go back to my brothers in Egypt to see whether they are still alive." And Jethro said to Moses, "Go in peace."
EXOD|4|19|And the LORD said to Moses in Midian, "Go back to Egypt, for all the men who were seeking your life are dead."
EXOD|4|20|So Moses took his wife and his sons and had them ride on a donkey, and went back to the land of Egypt. And Moses took the staff of God in his hand.
EXOD|4|21|And the LORD said to Moses, "When you go back to Egypt, see that you do before Pharaoh all the miracles that I have put in your power. But I will harden his heart, so that he will not let the people go.
EXOD|4|22|Then you shall say to Pharaoh, 'Thus says the LORD, Israel is my firstborn son,
EXOD|4|23|and I say to you, "Let my son go that he may serve me." If you refuse to let him go, behold, I will kill your firstborn son.'"
EXOD|4|24|At a lodging place on the way the LORD met him and sought to put him to death.
EXOD|4|25|Then Zipporah took a flint and cut off her son's foreskin and touched Moses' feet with it and said, "Surely you are a bridegroom of blood to me!"
EXOD|4|26|So he let him alone. It was then that she said, "A bridegroom of blood," because of the circumcision.
EXOD|4|27|The LORD said to Aaron, "Go into the wilderness to meet Moses." So he went and met him at the mountain of God and kissed him.
EXOD|4|28|And Moses told Aaron all the words of the LORD with which he had sent him to speak, and all the signs that he had commanded him to do.
EXOD|4|29|Then Moses and Aaron went and gathered together all the elders of the people of Israel.
EXOD|4|30|Aaron spoke all the words that the LORD had spoken to Moses and did the signs in the sight of the people.
EXOD|4|31|And the people believed; and when they heard that the LORD had visited the people of Israel and that he had seen their affliction, they bowed their heads and worshiped.
EXOD|5|1|Afterward Moses and Aaron went and said to Pharaoh, "Thus says the LORD, the God of Israel, 'Let my people go, that they may hold a feast to me in the wilderness.'"
EXOD|5|2|But Pharaoh said, "Who is the LORD, that I should obey his voice and let Israel go? I do not know the LORD, and moreover, I will not let Israel go."
EXOD|5|3|Then they said, "The God of the Hebrews has met with us. Please let us go a three days' journey into the wilderness that we may sacrifice to the LORD our God, lest he fall upon us with pestilence or with the sword."
EXOD|5|4|But the king of Egypt said to them, "Moses and Aaron, why do you take the people away from their work? Get back to your burdens."
EXOD|5|5|And Pharaoh said, "Behold, the people of the land are now many, and you make them rest from their burdens!"
EXOD|5|6|The same day Pharaoh commanded the taskmasters of the people and their foremen,
EXOD|5|7|"You shall no longer give the people straw to make bricks, as in the past; let them go and gather straw for themselves.
EXOD|5|8|But the number of bricks that they made in the past you shall impose on them, you shall by no means reduce it, for they are idle. Therefore they cry, 'Let us go and offer sacrifice to our God.'
EXOD|5|9|Let heavier work be laid on the men that they may labor at it and pay no regard to lying words."
EXOD|5|10|So the taskmasters and the foremen of the people went out and said to the people, "Thus says Pharaoh, 'I will not give you straw.
EXOD|5|11|Go and get your straw yourselves wherever you can find it, but your work will not be reduced in the least.'"
EXOD|5|12|So the people were scattered throughout all the land of Egypt to gather stubble for straw.
EXOD|5|13|The taskmasters were urgent, saying, "Complete your work, your daily task each day, as when there was straw."
EXOD|5|14|And the foremen of the people of Israel, whom Pharaoh's taskmasters had set over them, were beaten and were asked, "Why have you not done all your task of making bricks today and yesterday, as in the past?"
EXOD|5|15|Then the foremen of the people of Israel came and cried to Pharaoh, "Why do you treat your servants like this?
EXOD|5|16|No straw is given to your servants, yet they say to us, 'Make bricks!' And behold, your servants are beaten; but the fault is in your own people."
EXOD|5|17|But he said, "You are idle, you are idle; that is why you say, 'Let us go and sacrifice to the LORD.'
EXOD|5|18|Go now and work. No straw will be given you, but you must still deliver the same number of bricks."
EXOD|5|19|The foremen of the people of Israel saw that they were in trouble when they said, "You shall by no means reduce your number of bricks, your daily task each day."
EXOD|5|20|They met Moses and Aaron, who were waiting for them, as they came out from Pharaoh;
EXOD|5|21|and they said to them, "The LORD look on you and judge, because you have made us stink in the sight of Pharaoh and his servants, and have put a sword in their hand to kill us."
EXOD|5|22|Then Moses turned to the LORD and said, "O LORD, why have you done evil to this people? Why did you ever send me?
EXOD|5|23|For since I came to Pharaoh to speak in your name, he has done evil to this people, and you have not delivered your people at all."
EXOD|6|1|But the LORD said to Moses, "Now you shall see what I will do to Pharaoh; for with a strong hand he will send them out, and with a strong hand he will drive them out of his land."
EXOD|6|2|God spoke to Moses and said to him, "I am the LORD.
EXOD|6|3|I appeared to Abraham, to Isaac, and to Jacob, as God Almighty, but by my name the LORD I did not make myself known to them.
EXOD|6|4|I also established my covenant with them to give them the land of Canaan, the land in which they lived as sojourners.
EXOD|6|5|Moreover, I have heard the groaning of the people of Israel whom the Egyptians hold as slaves, and I have remembered my covenant.
EXOD|6|6|Say therefore to the people of Israel, 'I am the LORD, and I will bring you out from under the burdens of the Egyptians, and I will deliver you from slavery to them, and I will redeem you with an outstretched arm and with great acts of judgment.
EXOD|6|7|I will take you to be my people, and I will be your God, and you shall know that I am the LORD your God, who has brought you out from under the burdens of the Egyptians.
EXOD|6|8|I will bring you into the land that I swore to give to Abraham, to Isaac, and to Jacob. I will give it to you for a possession. I am the LORD.'"
EXOD|6|9|Moses spoke thus to the people of Israel, but they did not listen to Moses, because of their broken spirit and harsh slavery.
EXOD|6|10|So the LORD said to Moses,
EXOD|6|11|"Go in, tell Pharaoh king of Egypt to let the people of Israel go out of his land."
EXOD|6|12|But Moses said to the LORD, "Behold, the people of Israel have not listened to me. How then shall Pharaoh listen to me, for I am of uncircumcised lips?"
EXOD|6|13|But the LORD spoke to Moses and Aaron and gave them a charge about the people of Israel and about Pharaoh king of Egypt: to bring the people of Israel out of the land of Egypt.
EXOD|6|14|These are the heads of their fathers' houses: the sons of Reuben, the firstborn of Israel: Hanoch, Pallu, Hezron, and Carmi; these are the clans of Reuben.
EXOD|6|15|The sons of Simeon: Jemuel, Jamin, Ohad, Jachin, Zohar, and Shaul, the son of a Canaanite woman; these are the clans of Simeon.
EXOD|6|16|These are the names of the sons of Levi according to their generations: Gershon, Kohath, and Merari, the years of the life of Levi being 137 years.
EXOD|6|17|The sons of Gershon: Libni and Shimei, by their clans.
EXOD|6|18|The sons of Kohath: Amram, Izhar, Hebron, and Uzziel, the years of the life of Kohath being 133 years.
EXOD|6|19|The sons of Merari: Mahli and Mushi. These are the clans of the Levites according to their generations.
EXOD|6|20|Amram took as his wife Jochebed his father's sister, and she bore him Aaron and Moses, the years of the life of Amram being 137 years.
EXOD|6|21|The sons of Izhar: Korah, Nepheg, and Zichri.
EXOD|6|22|The sons of Uzziel: Mishael, Elzaphan, and Sithri.
EXOD|6|23|Aaron took as his wife Elisheba, the daughter of Amminadab and the sister of Nahshon, and she bore him Nadab, Abihu, Eleazar, and Ithamar.
EXOD|6|24|The sons of Korah: Assir, Elkanah, and Abiasaph; these are the clans of the Korahites.
EXOD|6|25|Eleazar, Aaron's son, took as his wife one of the daughters of Putiel, and she bore him Phinehas. These are the heads of the fathers' houses of the Levites by their clans.
EXOD|6|26|These are the Aaron and Moses to whom the LORD said: "Bring out the people of Israel from the land of Egypt by their hosts."
EXOD|6|27|It was they who spoke to Pharaoh king of Egypt about bringing out the people of Israel from Egypt, this Moses and this Aaron.
EXOD|6|28|On the day when the LORD spoke to Moses in the land of Egypt,
EXOD|6|29|the LORD said to Moses, "I am the LORD; tell Pharaoh king of Egypt all that I say to you."
EXOD|6|30|But Moses said to the LORD, "Behold, I am of uncircumcised lips. How will Pharaoh listen to me?"
EXOD|7|1|And the LORD said to Moses, "See, I have made you like God to Pharaoh, and your brother Aaron shall be your prophet.
EXOD|7|2|You shall speak all that I command you, and your brother Aaron shall tell Pharaoh to let the people of Israel go out of his land.
EXOD|7|3|But I will harden Pharaoh's heart, and though I multiply my signs and wonders in the land of Egypt,
EXOD|7|4|Pharaoh will not listen to you. Then I will lay my hand on Egypt and bring my hosts, my people the children of Israel, out of the land of Egypt by great acts of judgment.
EXOD|7|5|The Egyptians shall know that I am the LORD, when I stretch out my hand against Egypt and bring out the people of Israel from among them."
EXOD|7|6|Moses and Aaron did so; they did just as the LORD commanded them.
EXOD|7|7|Now Moses was eighty years old, and Aaron eighty-three years old, when they spoke to Pharaoh.
EXOD|7|8|Then the LORD said to Moses and Aaron,
EXOD|7|9|"When Pharaoh says to you, 'Prove yourselves by working a miracle,' then you shall say to Aaron, 'Take your staff and cast it down before Pharaoh, that it may become a serpent.'"
EXOD|7|10|So Moses and Aaron went to Pharaoh and did just as the LORD commanded. Aaron cast down his staff before Pharaoh and his servants, and it became a serpent.
EXOD|7|11|Then Pharaoh summoned the wise men and the sorcerers, and they, the magicians of Egypt, also did the same by their secret arts.
EXOD|7|12|For each man cast down his staff, and they became serpents. But Aaron's staff swallowed up their staffs.
EXOD|7|13|Still Pharaoh's heart was hardened, and he would not listen to them, as the LORD had said.
EXOD|7|14|Then the LORD said to Moses, "Pharaoh's heart is hardened; he refuses to let the people go.
EXOD|7|15|Go to Pharaoh in the morning, as he is going out to the water. Stand on the bank of the Nile to meet him, and take in your hand the staff that turned into a serpent.
EXOD|7|16|And you shall say to him, 'The LORD, the God of the Hebrews, sent me to you, saying, "Let my people go, that they may serve me in the wilderness. But so far, you have not obeyed."
EXOD|7|17|Thus says the LORD, "By this you shall know that I am the LORD: behold, with the staff that is in my hand I will strike the water that is in the Nile, and it shall turn into blood.
EXOD|7|18|The fish in the Nile shall die, and the Nile will stink, and the Egyptians will grow weary of drinking water from the Nile."'"
EXOD|7|19|And the LORD said to Moses, "Say to Aaron, 'Take your staff and stretch out your hand over the waters of Egypt, over their rivers, their canals, and their ponds, and all their pools of water, so that they may become blood, and there shall be blood throughout all the land of Egypt, even in vessels of wood and in vessels of stone.'"
EXOD|7|20|Moses and Aaron did as the LORD commanded. In the sight of Pharaoh and in the sight of his servants he lifted up the staff and struck the water in the Nile, and all the water in the Nile turned into blood.
EXOD|7|21|And the fish in the Nile died, and the Nile stank, so that the Egyptians could not drink water from the Nile. There was blood throughout all the land of Egypt.
EXOD|7|22|But the magicians of Egypt did the same by their secret arts. So Pharaoh's heart remained hardened, and he would not listen to them, as the LORD had said.
EXOD|7|23|Pharaoh turned and went into his house, and he did not take even this to heart.
EXOD|7|24|And all the Egyptians dug along the Nile for water to drink, for they could not drink the water of the Nile.
EXOD|7|25|Seven full days passed after the LORD had struck the Nile.
EXOD|8|1|Then the LORD said to Moses, "Go in to Pharaoh and say to him,'Thus says the LORD, "Let my people go, that they may serve me.
EXOD|8|2|But if you refuse to let them go, behold, I will plague all your country with frogs.
EXOD|8|3|The Nile shall swarm with frogs that shall come up into your house and into your bedroom and on your bed and into the houses of your servants and your people, and into your ovens and your kneading bowls.
EXOD|8|4|The frogs shall come up on you and on your people and on all your servants."'"
EXOD|8|5|And the LORD said to Moses, "Say to Aaron, 'Stretch out your hand with your staff over the rivers, over the canals and over the pools, and make frogs come up on the land of Egypt!'"
EXOD|8|6|So Aaron stretched out his hand over the waters of Egypt, and the frogs came up and covered the land of Egypt.
EXOD|8|7|But the magicians did the same by their secret arts and made frogs come up on the land of Egypt.
EXOD|8|8|Then Pharaoh called Moses and Aaron and said, "Plead with the LORD to take away the frogs from me and from my people, and I will let the people go to sacrifice to the LORD."
EXOD|8|9|Moses said to Pharaoh, "Be pleased to command me when I am to plead for you and for your servants and for your people, that the frogs be cut off from you and your houses and be left only in the Nile."
EXOD|8|10|And he said, "Tomorrow." Moses said, "Be it as you say, so that you may know that there is no one like the LORD our God.
EXOD|8|11|The frogs shall go away from you and your houses and your servants and your people. They shall be left only in the Nile."
EXOD|8|12|So Moses and Aaron went out from Pharaoh, and Moses cried to the LORD about the frogs, as he had agreed with Pharaoh.
EXOD|8|13|And the LORD did according to the word of Moses. The frogs died out in the houses, the courtyards, and the fields.
EXOD|8|14|And they gathered them together in heaps, and the land stank.
EXOD|8|15|But when Pharaoh saw that there was a respite, he hardened his heart and would not listen to them, as the LORD had said.
EXOD|8|16|Then the LORD said to Moses, "Say to Aaron, 'Stretch out your staff and strike the dust of the earth, so that it may become gnats in all the land of Egypt.'"
EXOD|8|17|And they did so. Aaron stretched out his hand with his staff and struck the dust of the earth, and there were gnats on man and beast. All the dust of the earth became gnats in all the land of Egypt.
EXOD|8|18|The magicians tried by their secret arts to produce gnats, but they could not. So there were gnats on man and beast.
EXOD|8|19|Then the magicians said to Pharaoh, "This is the finger of God." But Pharaoh's heart was hardened, and he would not listen to them, as the LORD had said.
EXOD|8|20|Then the LORD said to Moses, "Rise up early in the morning and present yourself to Pharaoh, as he goes out to the water, and say to him, 'Thus says the LORD, "Let my people go, that they may serve me.
EXOD|8|21|Or else, if you will not let my people go, behold, I will send swarms of flies on you and your servants and your people, and into your houses. And the houses of the Egyptians shall be filled with swarms of flies, and also the ground on which they stand.
EXOD|8|22|But on that day I will set apart the land of Goshen, where my people dwell, so that no swarms of flies shall be there, that you may know that I am the LORD in the midst of the earth.
EXOD|8|23|Thus I will put a division between my people and your people. Tomorrow this sign shall happen."'"
EXOD|8|24|And the LORD did so. There came great swarms of flies into the house of Pharaoh and into his servants' houses. Throughout all the land of Egypt the land was ruined by the swarms of flies.
EXOD|8|25|Then Pharaoh called Moses and Aaron and said, "Go, sacrifice to your God within the land."
EXOD|8|26|But Moses said, "It would not be right to do so, for the offerings we shall sacrifice to the LORD our God are an abomination to the Egyptians. If we sacrifice offerings abominable to the Egyptians before their eyes, will they not stone us?
EXOD|8|27|We must go three days' journey into the wilderness and sacrifice to the LORD our God as he tells us."
EXOD|8|28|So Pharaoh said, "I will let you go to sacrifice to the LORD your God in the wilderness; only you must not go very far away. Plead for me."
EXOD|8|29|Then Moses said, "Behold, I am going out from you and I will plead with the LORD that the swarms of flies may depart from Pharaoh, from his servants, and from his people, tomorrow. Only let not Pharaoh cheat again by not letting the people go to sacrifice to the LORD."
EXOD|8|30|So Moses went out from Pharaoh and prayed to the LORD.
EXOD|8|31|And the LORD did as Moses asked, and removed the swarms of flies from Pharaoh, from his servants, and from his people; not one remained.
EXOD|8|32|But Pharaoh hardened his heart this time also, and did not let the people go.
EXOD|9|1|Then the LORD said to Moses, "Go in to Pharaoh and say to him, 'Thus says the LORD, the God of the Hebrews, "Let my people go, that they may serve me.
EXOD|9|2|For if you refuse to let them go and still hold them,
EXOD|9|3|behold, the hand of the LORD will fall with a very severe plague upon your livestock that are in the field, the horses, the donkeys, the camels, the herds, and the flocks.
EXOD|9|4|But the LORD will make a distinction between the livestock of Israel and the livestock of Egypt, so that nothing of all that belongs to the people of Israel shall die."'"
EXOD|9|5|And the LORD set a time, saying, "Tomorrow the LORD will do this thing in the land."
EXOD|9|6|And the next day the LORD did this thing. All the livestock of the Egyptians died, but not one of the livestock of the people of Israel died.
EXOD|9|7|And Pharaoh sent, and behold, not one of the livestock of Israel was dead. But the heart of Pharaoh was hardened, and he did not let the people go.
EXOD|9|8|And the LORD said to Moses and Aaron, "Take handfuls of soot from the kiln, and let Moses throw them in the air in the sight of Pharaoh.
EXOD|9|9|It shall become fine dust over all the land of Egypt, and become boils breaking out in sores on man and beast throughout all the land of Egypt."
EXOD|9|10|So they took soot from the kiln and stood before Pharaoh. And Moses threw it in the air, and it became boils breaking out in sores on man and beast.
EXOD|9|11|And the magicians could not stand before Moses because of the boils, for the boils came upon the magicians and upon all the Egyptians.
EXOD|9|12|But the LORD hardened the heart of Pharaoh, and he did not listen to them, as the LORD had spoken to Moses.
EXOD|9|13|Then the LORD said to Moses, "Rise up early in the morning and present yourself before Pharaoh and say to him, 'Thus says the LORD, the God of the Hebrews, "Let my people go, that they may serve me.
EXOD|9|14|For this time I will send all my plagues on you yourself, and on your servants and your people, so that you may know that there is none like me in all the earth.
EXOD|9|15|For by now I could have put out my hand and struck you and your people with pestilence, and you would have been cut off from the earth.
EXOD|9|16|But for this purpose I have raised you up, to show you my power, so that my name may be proclaimed in all the earth.
EXOD|9|17|You are still exalting yourself against my people and will not let them go.
EXOD|9|18|Behold, about this time tomorrow I will cause very heavy hail to fall, such as never has been in Egypt from the day it was founded until now.
EXOD|9|19|Now therefore send, get your livestock and all that you have in the field into safe shelter, for every man and beast that is in the field and is not brought home will die when the hail falls on them."'"
EXOD|9|20|Then whoever feared the word of the LORD among the servants of Pharaoh hurried his slaves and his livestock into the houses,
EXOD|9|21|but whoever did not pay attention to the word of the LORD left his slaves and his livestock in the field.
EXOD|9|22|Then the LORD said to Moses, "Stretch out your hand toward heaven, so that there may be hail in all the land of Egypt, on man and beast and every plant of the field, in the land of Egypt."
EXOD|9|23|Then Moses stretched out his staff toward heaven, and the LORD sent thunder and hail, and fire ran down to the earth. And the LORD rained hail upon the land of Egypt.
EXOD|9|24|There was hail and fire flashing continually in the midst of the hail, very heavy hail, such as had never been in all the land of Egypt since it became a nation.
EXOD|9|25|The hail struck down everything that was in the field in all the land of Egypt, both man and beast. And the hail struck down every plant of the field and broke every tree of the field.
EXOD|9|26|Only in the land of Goshen, where the people of Israel were, was there no hail.
EXOD|9|27|Then Pharaoh sent and called Moses and Aaron and said to them, "This time I have sinned; the LORD is in the right, and I and my people are in the wrong.
EXOD|9|28|Plead with the LORD, for there has been enough of God's thunder and hail. I will let you go, and you shall stay no longer."
EXOD|9|29|Moses said to him, "As soon as I have gone out of the city, I will stretch out my hands to the LORD. The thunder will cease, and there will be no more hail, so that you may know that the earth is the LORD's.
EXOD|9|30|But as for you and your servants, I know that you do not yet fear the LORD God."
EXOD|9|31|(The flax and the barley were struck down, for the barley was in the ear and the flax was in bud.
EXOD|9|32|But the wheat and the emmer were not struck down, for they are late in coming up.)
EXOD|9|33|So Moses went out of the city from Pharaoh and stretched out his hands to the LORD, and the thunder and the hail ceased, and the rain no longer poured upon the earth.
EXOD|9|34|But when Pharaoh saw that the rain and the hail and the thunder had ceased, he sinned yet again and hardened his heart, he and his servants.
EXOD|9|35|So the heart of Pharaoh was hardened, and he did not let the people of Israel go, just as the LORD had spoken through Moses.
EXOD|10|1|Then the LORD said to Moses, "Go in to Pharaoh, for I have hardened his heart and the heart of his servants, that I may show these signs of mine among them,
EXOD|10|2|and that you may tell in the hearing of your son and of your grandson how I have dealt harshly with the Egyptians and what signs I have done among them, that you may know that I am the LORD."
EXOD|10|3|So Moses and Aaron went in to Pharaoh and said to him, "Thus says the LORD, the God of the Hebrews, 'How long will you refuse to humble yourself before me? Let my people go, that they may serve me.
EXOD|10|4|For if you refuse to let my people go, behold, tomorrow I will bring locusts into your country,
EXOD|10|5|and they shall cover the face of the land, so that no one can see the land. And they shall eat what is left to you after the hail, and they shall eat every tree of yours that grows in the field,
EXOD|10|6|and they shall fill your houses and the houses of all your servants and of all the Egyptians, as neither your fathers nor your grandfathers have seen, from the day they came on earth to this day.'"Then he turned and went out from Pharaoh.
EXOD|10|7|Then Pharaoh's servants said to him, "How long shall this man be a snare to us? Let the men go, that they may serve the LORD their God. Do you not yet understand that Egypt is ruined?"
EXOD|10|8|So Moses and Aaron were brought back to Pharaoh. And he said to them, "Go, serve the LORD your God. But which ones are to go?"
EXOD|10|9|Moses said, "We will go with our young and our old. We will go with our sons and daughters and with our flocks and herds, for we must hold a feast to the LORD."
EXOD|10|10|But he said to them, "The LORD be with you, if ever I let you and your little ones go! Look, you have some evil purpose in mind.
EXOD|10|11|No! Go, the men among you, and serve the LORD, for that is what you are asking." And they were driven out from Pharaoh's presence.
EXOD|10|12|Then the LORD said to Moses, "Stretch out your hand over the land of Egypt for the locusts, so that they may come upon the land of Egypt and eat every plant in the land, all that the hail has left."
EXOD|10|13|So Moses stretched out his staff over the land of Egypt, and the LORD brought an east wind upon the land all that day and all that night. When it was morning, the east wind had brought the locusts.
EXOD|10|14|The locusts came up over all the land of Egypt and settled on the whole country of Egypt, such a dense swarm of locusts as had never been before, nor ever will be again.
EXOD|10|15|They covered the face of the whole land, so that the land was darkened, and they ate all the plants in the land and all the fruit of the trees that the hail had left. Not a green thing remained, neither tree nor plant of the field, through all the land of Egypt.
EXOD|10|16|Then Pharaoh hastily called Moses and Aaron and said, "I have sinned against the LORD your God, and against you.
EXOD|10|17|Now therefore, forgive my sin, please, only this once, and plead with the LORD your God only to remove this death from me."
EXOD|10|18|So he went out from Pharaoh and pleaded with the LORD.
EXOD|10|19|And the LORD turned the wind into a very strong west wind, which lifted the locusts and drove them into the Red Sea. Not a single locust was left in all the country of Egypt.
EXOD|10|20|But the LORD hardened Pharaoh's heart, and he did not let the people of Israel go.
EXOD|10|21|Then the LORD said to Moses, "Stretch out your hand toward heaven, that there may be darkness over the land of Egypt, a darkness to be felt."
EXOD|10|22|So Moses stretched out his hand toward heaven, and there was pitch darkness in all the land of Egypt three days.
EXOD|10|23|They did not see one another, nor did anyone rise from his place for three days, but all the people of Israel had light where they lived.
EXOD|10|24|Then Pharaoh called Moses and said, "Go, serve the LORD; your little ones also may go with you; only let your flocks and your herds remain behind."
EXOD|10|25|But Moses said, "You must also let us have sacrifices and burnt offerings, that we may sacrifice to the LORD our God.
EXOD|10|26|Our livestock also must go with us; not a hoof shall be left behind, for we must take of them to serve the LORD our God, and we do not know with what we must serve the LORD until we arrive there."
EXOD|10|27|But the LORD hardened Pharaoh's heart, and he would not let them go.
EXOD|10|28|Then Pharaoh said to him, "Get away from me; take care never to see my face again, for on the day you see my face you shall die."
EXOD|10|29|Moses said, "As you say! I will not see your face again."
EXOD|11|1|The LORD said to Moses, "Yet one plague more I will bring upon Pharaoh and upon Egypt. Afterward he will let you go from here. When he lets you go, he will drive you away completely.
EXOD|11|2|Speak now in the hearing of the people, that they ask, every man of his neighbor and every woman of her neighbor, for silver and gold jewelry."
EXOD|11|3|And the LORD gave the people favor in the sight of the Egyptians. Moreover, the man Moses was very great in the land of Egypt, in the sight of Pharaoh's servants and in the sight of the people.
EXOD|11|4|So Moses said, "Thus says the LORD: About midnight I will go out in the midst of Egypt,
EXOD|11|5|and every firstborn in the land of Egypt shall die, from the firstborn of Pharaoh who sits on his throne, even to the firstborn of the slave girl who is behind the hand mill, and all the firstborn of the cattle.
EXOD|11|6|There shall be a great cry throughout all the land of Egypt, such as there has never been, nor ever will be again.
EXOD|11|7|But not a dog shall growl against any of the people of Israel, either man or beast, that you may know that the LORD makes a distinction between Egypt and Israel.
EXOD|11|8|And all these your servants shall come down to me and bow down to me, saying, 'Get out, you and all the people who follow you.' And after that I will go out." And he went out from Pharaoh in hot anger.
EXOD|11|9|Then the LORD said to Moses, "Pharaoh will not listen to you, that my wonders may be multiplied in the land of Egypt."
EXOD|11|10|Moses and Aaron did all these wonders before Pharaoh, and the LORD hardened Pharaoh's heart, and he did not let the people of Israel go out of his land.
EXOD|12|1|The LORD said to Moses and Aaron in the land of Egypt,
EXOD|12|2|"This month shall be for you the beginning of months. It shall be the first month of the year for you.
EXOD|12|3|Tell all the congregation of Israel that on the tenth day of this month every man shall take a lamb according to their fathers' houses, a lamb for a household.
EXOD|12|4|And if the household is too small for a lamb, then he and his nearest neighbor shall take according to the number of persons; according to what each can eat you shall make your count for the lamb.
EXOD|12|5|Your lamb shall be without blemish, a male a year old. You may take it from the sheep or from the goats,
EXOD|12|6|and you shall keep it until the fourteenth day of this month, when the whole assembly of the congregation of Israel shall kill their lambs at twilight.
EXOD|12|7|"Then they shall take some of the blood and put it on the two doorposts and the lintel of the houses in which they eat it.
EXOD|12|8|They shall eat the flesh that night, roasted on the fire; with unleavened bread and bitter herbs they shall eat it.
EXOD|12|9|Do not eat any of it raw or boiled in water, but roasted, its head with its legs and its inner parts.
EXOD|12|10|And you shall let none of it remain until the morning; anything that remains until the morning you shall burn.
EXOD|12|11|In this manner you shall eat it: with your belt fastened, your sandals on your feet, and your staff in your hand. And you shall eat it in haste. It is the LORD's Passover.
EXOD|12|12|For I will pass through the land of Egypt that night, and I will strike all the firstborn in the land of Egypt, both man and beast; and on all the gods of Egypt I will execute judgments: I am the LORD.
EXOD|12|13|The blood shall be a sign for you, on the houses where you are. And when I see the blood, I will pass over you, and no plague will befall you to destroy you, when I strike the land of Egypt.
EXOD|12|14|"This day shall be for you a memorial day, and you shall keep it as a feast to the LORD; throughout your generations, as a statute forever, you shall keep it as a feast.
EXOD|12|15|Seven days you shall eat unleavened bread. On the first day you shall remove leaven out of your houses, for if anyone eats what is leavened, from the first day until the seventh day, that person shall be cut off from Israel.
EXOD|12|16|On the first day you shall hold a holy assembly, and on the seventh day a holy assembly. No work shall be done on those days. But what everyone needs to eat, that alone may be prepared by you.
EXOD|12|17|And you shall observe the Feast of Unleavened Bread, for on this very day I brought your hosts out of the land of Egypt. Therefore you shall observe this day, throughout your generations, as a statute forever.
EXOD|12|18|In the first month, from the fourteenth day of the month at evening, you shall eat unleavened bread until the twenty-first day of the month at evening.
EXOD|12|19|For seven days no leaven is to be found in your houses. If anyone eats what is leavened, that person will be cut off from the congregation of Israel, whether he is a sojourner or a native of the land.
EXOD|12|20|You shall eat nothing leavened; in all your dwelling places you shall eat unleavened bread."
EXOD|12|21|Then Moses called all the elders of Israel and said to them, "Go and select lambs for yourselves according to your clans, and kill the Passover lamb.
EXOD|12|22|Take a bunch of hyssop and dip it in the blood that is in the basin, and touch the lintel and the two doorposts with the blood that is in the basin. None of you shall go out of the door of his house until the morning.
EXOD|12|23|For the LORD will pass through to strike the Egyptians, and when he sees the blood on the lintel and on the two doorposts, the LORD will pass over the door and will not allow the destroyer to enter your houses to strike you.
EXOD|12|24|You shall observe this rite as a statute for you and for your sons forever.
EXOD|12|25|And when you come to the land that the LORD will give you, as he has promised, you shall keep this service.
EXOD|12|26|And when your children say to you, 'What do you mean by this service?'
EXOD|12|27|you shall say, 'It is the sacrifice of the LORD's Passover, for he passed over the houses of the people of Israel in Egypt, when he struck the Egyptians but spared our houses.'"And the people bowed their heads and worshiped.
EXOD|12|28|Then the people of Israel went and did so; as the LORD had commanded Moses and Aaron, so they did.
EXOD|12|29|At midnight the LORD struck down all the firstborn in the land of Egypt, from the firstborn of Pharaoh who sat on his throne to the firstborn of the captive who was in the dungeon, and all the firstborn of the livestock.
EXOD|12|30|And Pharaoh rose up in the night, he and all his servants and all the Egyptians. And there was a great cry in Egypt, for there was not a house where someone was not dead.
EXOD|12|31|Then he summoned Moses and Aaron by night and said, "Up, go out from among my people, both you and the people of Israel; and go, serve the LORD, as you have said.
EXOD|12|32|Take your flocks and your herds, as you have said, and be gone, and bless me also!"
EXOD|12|33|The Egyptians were urgent with the people to send them out of the land in haste. For they said, "We shall all be dead."
EXOD|12|34|So the people took their dough before it was leavened, their kneading bowls being bound up in their cloaks on their shoulders.
EXOD|12|35|The people of Israel had also done as Moses told them, for they had asked the Egyptians for silver and gold jewelry and for clothing.
EXOD|12|36|And the LORD had given the people favor in the sight of the Egyptians, so that they let them have what they asked. Thus they plundered the Egyptians.
EXOD|12|37|And the people of Israel journeyed from Rameses to Succoth, about six hundred thousand men on foot, besides women and children.
EXOD|12|38|A mixed multitude also went up with them, and very much livestock, both flocks and herds.
EXOD|12|39|And they baked unleavened cakes of the dough that they had brought out of Egypt, for it was not leavened, because they were thrust out of Egypt and could not wait, nor had they prepared any provisions for themselves.
EXOD|12|40|The time that the people of Israel lived in Egypt was 430 years.
EXOD|12|41|At the end of 430 years, on that very day, all the hosts of the LORD went out from the land of Egypt.
EXOD|12|42|It was a night of watching by the LORD, to bring them out of the land of Egypt; so this same night is a night of watching kept to the LORD by all the people of Israel throughout their generations.
EXOD|12|43|And the LORD said to Moses and Aaron, "This is the statute of the Passover: no foreigner shall eat of it,
EXOD|12|44|but every slave that is bought for money may eat of it after you have circumcised him.
EXOD|12|45|No foreigner or hired servant may eat of it.
EXOD|12|46|It shall be eaten in one house; you shall not take any of the flesh outside the house, and you shall not break any of its bones.
EXOD|12|47|All the congregation of Israel shall keep it.
EXOD|12|48|If a stranger shall sojourn with you and would keep the Passover to the LORD, let all his males be circumcised. Then he may come near and keep it; he shall be as a native of the land. But no uncircumcised person shall eat of it.
EXOD|12|49|There shall be one law for the native and for the stranger who sojourns among you."
EXOD|12|50|All the people of Israel did just as the LORD commanded Moses and Aaron.
EXOD|12|51|And on that very day the LORD brought the people of Israel out of the land of Egypt by their hosts.
EXOD|13|1|The LORD said to Moses,
EXOD|13|2|"Consecrate to me all the firstborn. Whatever is the first to open the womb among the people of Israel, both of man and of beast, is mine."
EXOD|13|3|Then Moses said to the people, "Remember this day in which you came out from Egypt, out of the house of slavery, for by strength of hand the LORD brought you out from this place. No leavened bread shall be eaten.
EXOD|13|4|Today, in the month of Abib, you are going out.
EXOD|13|5|And when the LORD brings you into the land of the Canaanites, the Hittites, the Amorites, the Hivites, and the Jebusites, which he swore to your fathers to give you, a land flowing with milk and honey, you shall keep this service in this month.
EXOD|13|6|Seven days you shall eat unleavened bread, and on the seventh day there shall be a feast to the LORD.
EXOD|13|7|Unleavened bread shall be eaten for seven days; no leavened bread shall be seen with you, and no leaven shall be seen with you in all your territory.
EXOD|13|8|You shall tell your son on that day, 'It is because of what the LORD did for me when I came out of Egypt.'
EXOD|13|9|And it shall be to you as a sign on your hand and as a memorial between your eyes, that the law of the LORD may be in your mouth. For with a strong hand the LORD has brought you out of Egypt.
EXOD|13|10|You shall therefore keep this statute at its appointed time from year to year.
EXOD|13|11|"When the LORD brings you into the land of the Canaanites, as he swore to you and your fathers, and shall give it to you,
EXOD|13|12|you shall set apart to the LORD all that first opens the womb. All the firstborn of your animals that are males shall be the LORD's.
EXOD|13|13|Every firstborn of a donkey you shall redeem with a lamb, or if you will not redeem it you shall break its neck. Every firstborn of man among your sons you shall redeem.
EXOD|13|14|And when in time to come your son asks you, 'What does this mean?' you shall say to him, 'By strength of hand the LORD brought us out of Egypt, from the house of slavery.
EXOD|13|15|For when Pharaoh stubbornly refused to let us go, the LORD killed all the firstborn in the land of Egypt, both the firstborn of man and the firstborn of animals. Therefore I sacrifice to the LORD all the males that first open the womb, but all the firstborn of my sons I redeem.'
EXOD|13|16|It shall be as a mark on your hand or frontlets between your eyes, for by a strong hand the LORD brought us out of Egypt."
EXOD|13|17|When Pharaoh let the people go, God did not lead them by way of the land of the Philistines, although that was near. For God said, "Lest the people change their minds when they see war and return to Egypt."
EXOD|13|18|But God led the people around by the way of the wilderness toward the Red Sea. And the people of Israel went up out of the land of Egypt equipped for battle.
EXOD|13|19|Moses took the bones of Joseph with him, for Joseph had made the sons of Israel solemnly swear, saying, "God will surely visit you, and you shall carry up my bones with you from here."
EXOD|13|20|And they moved on from Succoth and encamped at Etham, on the edge of the wilderness.
EXOD|13|21|And the LORD went before them by day in a pillar of cloud to lead them along the way, and by night in a pillar of fire to give them light, that they might travel by day and by night.
EXOD|13|22|The pillar of cloud by day and the pillar of fire by night did not depart from before the people.
EXOD|14|1|Then the LORD said to Moses,
EXOD|14|2|"Tell the people of Israel to turn back and encamp in front of Pihahiroth, between Migdol and the sea, in front of Baal-zephon; you shall encamp facing it, by the sea.
EXOD|14|3|For Pharaoh will say of the people of Israel, 'They are wandering in the land; the wilderness has shut them in.'
EXOD|14|4|And I will harden Pharaoh's heart, and he will pursue them, and I will get glory over Pharaoh and all his host, and the Egyptians shall know that I am the LORD." And they did so.
EXOD|14|5|When the king of Egypt was told that the people had fled, the mind of Pharaoh and his servants was changed toward the people, and they said, "What is this we have done, that we have let Israel go from serving us?"
EXOD|14|6|So he made ready his chariot and took his army with him,
EXOD|14|7|and took six hundred chosen chariots and all the other chariots of Egypt with officers over all of them.
EXOD|14|8|And the LORD hardened the heart of Pharaoh king of Egypt, and he pursued the people of Israel while the people of Israel were going out defiantly.
EXOD|14|9|The Egyptians pursued them, all Pharaoh's horses and chariots and his horsemen and his army, and overtook them encamped at the sea, by Pihahiroth, in front of Baal-zephon.
EXOD|14|10|When Pharaoh drew near, the people of Israel lifted up their eyes, and behold, the Egyptians were marching after them, and they feared greatly. And the people of Israel cried out to the LORD.
EXOD|14|11|They said to Moses, "Is it because there are no graves in Egypt that you have taken us away to die in the wilderness? What have you done to us in bringing us out of Egypt?
EXOD|14|12|Is not this what we said to you in Egypt, 'Leave us alone that we may serve the Egyptians'? For it would have been better for us to serve the Egyptians than to die in the wilderness."
EXOD|14|13|And Moses said to the people, "Fear not, stand firm, and see the salvation of the LORD, which he will work for you today. For the Egyptians whom you see today, you shall never see again.
EXOD|14|14|The LORD will fight for you, and you have only to be silent."
EXOD|14|15|The LORD said to Moses, "Why do you cry to me? Tell the people of Israel to go forward.
EXOD|14|16|Lift up your staff, and stretch out your hand over the sea and divide it, that the people of Israel may go through the sea on dry ground.
EXOD|14|17|And I will harden the hearts of the Egyptians so that they shall go in after them, and I will get glory over Pharaoh and all his host, his chariots, and his horsemen.
EXOD|14|18|And the Egyptians shall know that I am the LORD, when I have gotten glory over Pharaoh, his chariots, and his horsemen."
EXOD|14|19|Then the angel of God who was going before the host of Israel moved and went behind them, and the pillar of cloud moved from before them and stood behind them,
EXOD|14|20|coming between the host of Egypt and the host of Israel. And there was the cloud and the darkness. And it lit up the night without one coming near the other all night.
EXOD|14|21|Then Moses stretched out his hand over the sea, and the LORD drove the sea back by a strong east wind all night and made the sea dry land, and the waters were divided.
EXOD|14|22|And the people of Israel went into the midst of the sea on dry ground, the waters being a wall to them on their right hand and on their left.
EXOD|14|23|The Egyptians pursued and went in after them into the midst of the sea, all Pharaoh's horses, his chariots, and his horsemen.
EXOD|14|24|And in the morning watch the LORD in the pillar of fire and of cloud looked down on the Egyptian forces and threw the Egyptian forces into a panic,
EXOD|14|25|clogging their chariot wheels so that they drove heavily. And the Egyptians said, "Let us flee from before Israel, for the LORD fights for them against the Egyptians."
EXOD|14|26|Then the LORD said to Moses, "Stretch out your hand over the sea, that the water may come back upon the Egyptians, upon their chariots, and upon their horsemen."
EXOD|14|27|So Moses stretched out his hand over the sea, and the sea returned to its normal course when the morning appeared. And as the Egyptians fled into it, the LORD threw the Egyptians into the midst of the sea.
EXOD|14|28|The waters returned and covered the chariots and the horsemen; of all the host of Pharaoh that had followed them into the sea, not one of them remained.
EXOD|14|29|But the people of Israel walked on dry ground through the sea, the waters being a wall to them on their right hand and on their left.
EXOD|14|30|Thus the LORD saved Israel that day from the hand of the Egyptians, and Israel saw the Egyptians dead on the seashore.
EXOD|14|31|Israel saw the great power that the LORD used against the Egyptians, so the people feared the LORD, and they believed in the LORD and in his servant Moses.
EXOD|15|1|Then Moses and the people of Israel sang this song to the LORD, saying, "I will sing to the LORD, for he has triumphed gloriously; the horse and his rider he has thrown into the sea.
EXOD|15|2|The LORD is my strength and my song, and he has become my salvation; this is my God, and I will praise him, my father's God, and I will exalt him.
EXOD|15|3|The LORD is a man of war; the LORD is his name.
EXOD|15|4|"Pharaoh's chariots and his host he cast into the sea, and his chosen officers were sunk in the Red Sea.
EXOD|15|5|The floods covered them; they went down into the depths like a stone.
EXOD|15|6|Your right hand, O LORD, glorious in power, your right hand, O LORD, shatters the enemy.
EXOD|15|7|In the greatness of your majesty you overthrow your adversaries; you send out your fury; it consumes them like stubble.
EXOD|15|8|At the blast of your nostrils the waters piled up; the floods stood up in a heap; the deeps congealed in the heart of the sea.
EXOD|15|9|The enemy said, 'I will pursue, I will overtake, I will divide the spoil, my desire shall have its fill of them. I will draw my sword; my hand shall destroy them.'
EXOD|15|10|You blew with your wind; the sea covered them; they sank like lead in the mighty waters.
EXOD|15|11|"Who is like you, O LORD, among the gods? Who is like you, majestic in holiness, awesome in glorious deeds, doing wonders?
EXOD|15|12|You stretched out your right hand; the earth swallowed them.
EXOD|15|13|"You have led in your steadfast love the people whom you have redeemed; you have guided them by your strength to your holy abode.
EXOD|15|14|The peoples have heard; they tremble; pangs have seized the inhabitants of Philistia.
EXOD|15|15|Now are the chiefs of Edom dismayed; trembling seizes the leaders of Moab; all the inhabitants of Canaan have melted away.
EXOD|15|16|Terror and dread fall upon them; because of the greatness of your arm, they are still as a stone, till your people, O LORD, pass by, till the people pass by whom you have purchased.
EXOD|15|17|You will bring them in and plant them on your own mountain, the place, O LORD, which you have made for your abode, the sanctuary, O Lord, which your hands have established.
EXOD|15|18|The LORD will reign forever and ever."
EXOD|15|19|For when the horses of Pharaoh with his chariots and his horsemen went into the sea, the LORD brought back the waters of the sea upon them, but the people of Israel walked on dry ground in the midst of the sea.
EXOD|15|20|Then Miriam the prophetess, the sister of Aaron, took a tambourine in her hand, and all the women went out after her with tambourines and dancing.
EXOD|15|21|And Miriam sang to them: "Sing to the LORD, for he has triumphed gloriously; the horse and his rider he has thrown into the sea."
EXOD|15|22|Then Moses made Israel set out from the Red Sea, and they went into the wilderness of Shur. They went three days in the wilderness and found no water.
EXOD|15|23|When they came to Marah, they could not drink the water of Marah because it was bitter; therefore it was named Marah.
EXOD|15|24|And the people grumbled against Moses, saying, "What shall we drink?"
EXOD|15|25|And he cried to the LORD, and the LORD showed him a log, and he threw it into the water, and the water became sweet. There the LORD made for them a statute and a rule, and there he tested them,
EXOD|15|26|saying, "If you will diligently listen to the voice of the LORD your God, and do that which is right in his eyes, and give ear to his commandments and keep all his statutes, I will put none of the diseases on you that I put on the Egyptians, for I am the LORD, your healer."
EXOD|15|27|Then they came to Elim, where there were twelve springs of water and seventy palm trees, and they encamped there by the water.
EXOD|16|1|They set out from Elim, and all the congregation of the people of Israel came to the wilderness of Sin, which is between Elim and Sinai, on the fifteenth day of the second month after they had departed from the land of Egypt.
EXOD|16|2|And the whole congregation of the people of Israel grumbled against Moses and Aaron in the wilderness,
EXOD|16|3|and the people of Israel said to them, "Would that we had died by the hand of the LORD in the land of Egypt, when we sat by the meat pots and ate bread to the full, for you have brought us out into this wilderness to kill this whole assembly with hunger."
EXOD|16|4|Then the LORD said to Moses, "Behold, I am about to rain bread from heaven for you, and the people shall go out and gather a day's portion every day, that I may test them, whether they will walk in my law or not.
EXOD|16|5|On the sixth day, when they prepare what they bring in, it will be twice as much as they gather daily."
EXOD|16|6|So Moses and Aaron said to all the people of Israel, "At evening you shall know that it was the LORD who brought you out of the land of Egypt,
EXOD|16|7|and in the morning you shall see the glory of the LORD, because he has heard your grumbling against the LORD. For what are we, that you grumble against us?"
EXOD|16|8|And Moses said, "When the LORD gives you in the evening meat to eat and in the morning bread to the full, because the LORD has heard your grumbling that you grumble against him- what are we? Your grumbling is not against us but against the LORD."
EXOD|16|9|Then Moses said to Aaron, "Say to the whole congregation of the people of Israel, 'Come near before the LORD, for he has heard your grumbling.'"
EXOD|16|10|And as soon as Aaron spoke to the whole congregation of the people of Israel, they looked toward the wilderness, and behold, the glory of the LORD appeared in the cloud.
EXOD|16|11|And the LORD said to Moses,
EXOD|16|12|"I have heard the grumbling of the people of Israel. Say to them, 'At twilight you shall eat meat, and in the morning you shall be filled with bread. Then you shall know that I am the LORD your God.'"
EXOD|16|13|In the evening quail came up and covered the camp, and in the morning dew lay around the camp.
EXOD|16|14|And when the dew had gone up, there was on the face of the wilderness a fine, flake-like thing, fine as frost on the ground.
EXOD|16|15|When the people of Israel saw it, they said to one another, "What is it?" For they did not know what it was. And Moses said to them, "It is the bread that the LORD has given you to eat.
EXOD|16|16|This is what the LORD has commanded: 'Gather of it, each one of you, as much as he can eat. You shall each take an omer, according to the number of the persons that each of you has in his tent.'"
EXOD|16|17|And the people of Israel did so. They gathered, some more, some less.
EXOD|16|18|But when they measured it with an omer, whoever gathered much had nothing left over, and whoever gathered little had no lack. Each of them gathered as much as he could eat.
EXOD|16|19|And Moses said to them, "Let no one leave any of it over till the morning."
EXOD|16|20|But they did not listen to Moses. Some left part of it till the morning, and it bred worms and stank. And Moses was angry with them.
EXOD|16|21|Morning by morning they gathered it, each as much as he could eat; but when the sun grew hot, it melted.
EXOD|16|22|On the sixth day they gathered twice as much bread, two omers each. And when all the leaders of the congregation came and told Moses,
EXOD|16|23|he said to them, "This is what the LORD has commanded: 'Tomorrow is a day of solemn rest, a holy Sabbath to the LORD; bake what you will bake and boil what you will boil, and all that is left over lay aside to be kept till the morning.'"
EXOD|16|24|So they laid it aside till the morning, as Moses commanded them, and it did not stink, and there were no worms in it.
EXOD|16|25|Moses said, "Eat it today, for today is a Sabbath to the LORD; today you will not find it in the field.
EXOD|16|26|Six days you shall gather it, but on the seventh day, which is a Sabbath, there will be none."
EXOD|16|27|On the seventh day some of the people went out to gather, but they found none.
EXOD|16|28|And the LORD said to Moses, "How long will you refuse to keep my commandments and my laws?
EXOD|16|29|See! The LORD has given you the Sabbath; therefore on the sixth day he gives you bread for two days. Remain each of you in his place; let no one go out of his place on the seventh day."
EXOD|16|30|So the people rested on the seventh day.
EXOD|16|31|Now the house of Israel called its name manna. It was like coriander seed, white, and the taste of it was like wafers made with honey.
EXOD|16|32|Moses said, "This is what the LORD has commanded: 'Let an omer of it be kept throughout your generations, so that they may see the bread with which I fed you in the wilderness, when I brought you out of the land of Egypt.'"
EXOD|16|33|And Moses said to Aaron, "Take a jar, and put an omer of manna in it, and place it before the LORD to be kept throughout your generations."
EXOD|16|34|As the LORD commanded Moses, so Aaron placed it before the testimony to be kept.
EXOD|16|35|The people of Israel ate the manna forty years, till they came to a habitable land. They ate the manna till they came to the border of the land of Canaan.
EXOD|16|36|(An omer is the tenth part of an ephah.)
EXOD|17|1|All the congregation of the people of Israel moved on from the wilderness of Sin by stages, according to the commandment of the LORD, and camped at Rephidim, but there was no water for the people to drink.
EXOD|17|2|Therefore the people quarreled with Moses and said, "Give us water to drink." And Moses said to them, "Why do you quarrel with me? Why do you test the LORD?"
EXOD|17|3|But the people thirsted there for water, and the people grumbled against Moses and said, "Why did you bring us up out of Egypt, to kill us and our children and our livestock with thirst?"
EXOD|17|4|So Moses cried to the LORD, "What shall I do with this people? They are almost ready to stone me."
EXOD|17|5|And the LORD said to Moses, "Pass on before the people, taking with you some of the elders of Israel, and take in your hand the staff with which you struck the Nile, and go.
EXOD|17|6|Behold, I will stand before you there on the rock at Horeb, and you shall strike the rock, and water shall come out of it, and the people will drink." And Moses did so, in the sight of the elders of Israel.
EXOD|17|7|And he called the name of the place Massah and Meribah, because of the quarreling of the people of Israel, and because they tested the LORD by saying, "Is the LORD among us or not?"
EXOD|17|8|Then Amalek came and fought with Israel at Rephidim.
EXOD|17|9|So Moses said to Joshua, "Choose for us men, and go out and fight with Amalek. Tomorrow I will stand on the top of the hill with the staff of God in my hand."
EXOD|17|10|So Joshua did as Moses told him, and fought with Amalek, while Moses, Aaron, and Hur went up to the top of the hill.
EXOD|17|11|Whenever Moses held up his hand, Israel prevailed, and whenever he lowered his hand, Amalek prevailed.
EXOD|17|12|But Moses' hands grew weary, so they took a stone and put it under him, and he sat on it, while Aaron and Hur held up his hands, one on one side, and the other on the other side. So his hands were steady until the going down of the sun.
EXOD|17|13|And Joshua overwhelmed Amalek and his people with the sword.
EXOD|17|14|Then the LORD said to Moses, "Write this as a memorial in a book and recite it in the ears of Joshua, that I will utterly blot out the memory of Amalek from under heaven."
EXOD|17|15|And Moses built an altar and called the name of it, The LORD is my banner,
EXOD|17|16|saying, "A hand upon the throne of the LORD! The LORD will have war with Amalek from generation to generation."
EXOD|18|1|Jethro, the priest of Midian, Moses' father-in-law, heard of all that God had done for Moses and for Israel his people, how the LORD had brought Israel out of Egypt.
EXOD|18|2|Now Jethro, Moses' father-in-law, had taken Zipporah, Moses' wife, after he had sent her home,
EXOD|18|3|along with her two sons. The name of the one was Gershom (for he said, "I have been a sojourner in a foreign land"),
EXOD|18|4|and the name of the other, Eliezer (for he said, "The God of my father was my help, and delivered me from the sword of Pharaoh").
EXOD|18|5|Jethro, Moses' father-in-law, came with his sons and his wife to Moses in the wilderness where he was encamped at the mountain of God.
EXOD|18|6|And when he sent word to Moses, "I, your father-in-law Jethro, am coming to you with your wife and her two sons with her,"
EXOD|18|7|Moses went out to meet his father-in-law and bowed down and kissed him. And they asked each other of their welfare and went into the tent.
EXOD|18|8|Then Moses told his father-in-law all that the LORD had done to Pharaoh and to the Egyptians for Israel's sake, all the hardship that had come upon them in the way, and how the LORD had delivered them.
EXOD|18|9|And Jethro rejoiced for all the good that the LORD had done to Israel, in that he had delivered them out of the hand of the Egyptians.
EXOD|18|10|Jethro said, "Blessed be the LORD, who has delivered you out of the hand of the Egyptians and out of the hand of Pharaoh and has delivered the people from under the hand of the Egyptians.
EXOD|18|11|Now I know that the LORD is greater than all gods, because in this affair they dealt arrogantly with the people."
EXOD|18|12|And Jethro, Moses' father-in-law, brought a burnt offering and sacrifices to God; and Aaron came with all the elders of Israel to eat bread with Moses' father-in-law before God.
EXOD|18|13|The next day Moses sat to judge the people, and the people stood around Moses from morning till evening.
EXOD|18|14|When Moses' father-in-law saw all that he was doing for the people, he said, "What is this that you are doing for the people? Why do you sit alone, and all the people stand around you from morning till evening?"
EXOD|18|15|And Moses said to his father-in-law, "Because the people come to me to inquire of God;
EXOD|18|16|when they have a dispute, they come to me and I decide between one person and another, and I make them know the statutes of God and his laws."
EXOD|18|17|Moses' father-in-law said to him, "What you are doing is not good.
EXOD|18|18|You and the people with you will certainly wear yourselves out, for the thing is too heavy for you. You are not able to do it alone.
EXOD|18|19|Now obey my voice; I will give you advice, and God be with you! You shall represent the people before God and bring their cases to God,
EXOD|18|20|and you shall warn them about the statutes and the laws, and make them know the way in which they must walk and what they must do.
EXOD|18|21|Moreover, look for able men from all the people, men who fear God, who are trustworthy and hate a bribe, and place such men over the people as chiefs of thousands, of hundreds, of fifties, and of tens.
EXOD|18|22|And let them judge the people at all times. Every great matter they shall bring to you, but any small matter they shall decide themselves. So it will be easier for you, and they will bear the burden with you.
EXOD|18|23|If you do this, God will direct you, you will be able to endure, and all this people also will go to their place in peace."
EXOD|18|24|So Moses listened to the voice of his father-in-law and did all that he had said.
EXOD|18|25|Moses chose able men out of all Israel and made them heads over the people, chiefs of thousands, of hundreds, of fifties, and of tens.
EXOD|18|26|And they judged the people at all times. Any hard case they brought to Moses, but any small matter they decided themselves.
EXOD|18|27|Then Moses let his father-in-law depart, and he went away to his own country.
EXOD|19|1|On the third new moon after the people of Israel had gone out of the land of Egypt, on that day they came into the wilderness of Sinai.
EXOD|19|2|They set out from Rephidim and came into the wilderness of Sinai, and they encamped in the wilderness. There Israel encamped before the mountain,
EXOD|19|3|while Moses went up to God. The LORD called to him out of the mountain, saying, "Thus you shall say to the house of Jacob, and tell the people of Israel:
EXOD|19|4|You yourselves have seen what I did to the Egyptians, and how I bore you on eagles' wings and brought you to myself.
EXOD|19|5|Now therefore, if you will indeed obey my voice and keep my covenant, you shall be my treasured possession among all peoples, for all the earth is mine;
EXOD|19|6|and you shall be to me a kingdom of priests and a holy nation. These are the words that you shall speak to the people of Israel."
EXOD|19|7|So Moses came and called the elders of the people and set before them all these words that the LORD had commanded him.
EXOD|19|8|All the people answered together and said, "All that the LORD has spoken we will do." And Moses reported the words of the people to the LORD.
EXOD|19|9|And the LORD said to Moses. "Behold, I am coming to you in a thick cloud, that the people may hear when I speak with you, and may also believe you forever." When Moses told the words of the people to the LORD,
EXOD|19|10|the LORD said to Moses, "Go to the people and consecrate them today and tomorrow, and let them wash their garments
EXOD|19|11|and be ready for the third day. For on the third day the LORD will come down on Mount Sinai in the sight of all the people.
EXOD|19|12|And you shall set limits for the people all around, saying, 'Take care not to go up into the mountain or touch the edge of it. Whoever touches the mountain shall be put to death.
EXOD|19|13|No hand shall touch him, but he shall be stoned or shot; whether beast or man, he shall not live.' When the trumpet sounds a long blast, they shall come up to the mountain."
EXOD|19|14|So Moses went down from the mountain to the people and consecrated the people; and they washed their garments.
EXOD|19|15|And he said to the people, "Be ready for the third day; do not go near a woman."
EXOD|19|16|On the morning of the third day there were thunders and lightnings and a thick cloud on the mountain and a very loud trumpet blast, so that all the people in the camp trembled.
EXOD|19|17|Then Moses brought the people out of the camp to meet God, and they took their stand at the foot of the mountain.
EXOD|19|18|Now Mount Sinai was wrapped in smoke because the LORD had descended on it in fire. The smoke of it went up like the smoke of a kiln, and the whole mountain trembled greatly.
EXOD|19|19|And as the sound of the trumpet grew louder and louder, Moses spoke, and God answered him in thunder.
EXOD|19|20|The LORD came down on Mount Sinai, to the top of the mountain. And the LORD called Moses to the top of the mountain, and Moses went up.
EXOD|19|21|And the LORD said to Moses, "Go down and warn the people, lest they break through to the LORD to look and many of them perish.
EXOD|19|22|Also let the priests who come near to the LORD consecrate themselves, lest the LORD break out against them."
EXOD|19|23|And Moses said to the LORD, "The people cannot come up to Mount Sinai, for you yourself warned us, saying, 'Set limits around the mountain and consecrate it.'"
EXOD|19|24|And the LORD said to him, "Go down, and come up bringing Aaron with you. But do not let the priests and the people break through to come up to the LORD, lest he break out against them."
EXOD|19|25|So Moses went down to the people and told them.
EXOD|20|1|And God spoke all these words, saying,
EXOD|20|2|"I am the LORD your God, who brought you out of the land of Egypt, out of the house of slavery.
EXOD|20|3|"You shall have no other gods before me.
EXOD|20|4|"You shall not make for yourself a carved image, or any likeness of anything that is in heaven above, or that is in the earth beneath, or that is in the water under the earth.
EXOD|20|5|You shall not bow down to them or serve them, for I the LORD your God am a jealous God, visiting the iniquity of the fathers on the children to the third and the fourth generation of those who hate me,
EXOD|20|6|but showing steadfast love to thousands of those who love me and keep my commandments.
EXOD|20|7|"You shall not take the name of the LORD your God in vain, for the LORD will not hold him guiltless who takes his name in vain.
EXOD|20|8|"Remember the Sabbath day, to keep it holy.
EXOD|20|9|Six days you shall labor, and do all your work,
EXOD|20|10|but the seventh day is a Sabbath to the LORD your God. On it you shall not do any work, you, or your son, or your daughter, your male servant, or your female servant, or your livestock, or the sojourner who is within your gates.
EXOD|20|11|For in six days the LORD made heaven and earth, the sea, and all that is in them, and rested the seventh day. Therefore the LORD blessed the Sabbath day and made it holy.
EXOD|20|12|"Honor your father and your mother, that your days may be long in the land that the LORD your God is giving you.
EXOD|20|13|"You shall not murder.
EXOD|20|14|"You shall not commit adultery.
EXOD|20|15|"You shall not steal.
EXOD|20|16|"You shall not bear false witness against your neighbor.
EXOD|20|17|"You shall not covet your neighbor's house; you shall not covet your neighbor's wife, or his male servant, or his female servant, or his ox, or his donkey, or anything that is your neighbor's."
EXOD|20|18|Now when all the people saw the thunder and the flashes of lightning and the sound of the trumpet and the mountain smoking, the people were afraid and trembled, and they stood far off
EXOD|20|19|and said to Moses, "You speak to us, and we will listen; but do not let God speak to us, lest we die."
EXOD|20|20|Moses said to the people, "Do not fear, for God has come to test you, that the fear of him may be before you, that you may not sin."
EXOD|20|21|The people stood far off, while Moses drew near to the thick darkness where God was.
EXOD|20|22|And the LORD said to Moses, "Thus you shall say to the people of Israel: 'You have seen for yourselves that I have talked with you from heaven.
EXOD|20|23|You shall not make gods of silver to be with me, nor shall you make for yourselves gods of gold.
EXOD|20|24|An altar of earth you shall make for me and sacrifice on it your burnt offerings and your peace offerings, your sheep and your oxen. In every place where I cause my name to be remembered I will come to you and bless you.
EXOD|20|25|If you make me an altar of stone, you shall not build it of hewn stones, for if you wield your tool on it you profane it.
EXOD|20|26|And you shall not go up by steps to my altar, that your nakedness be not exposed on it.'
EXOD|21|1|"Now these are the rules that you shall set before them.
EXOD|21|2|When you buy a Hebrew slave, he shall serve six years, and in the seventh he shall go out free, for nothing.
EXOD|21|3|If he comes in single, he shall go out single; if he comes in married, then his wife shall go out with him.
EXOD|21|4|If his master gives him a wife and she bears him sons or daughters, the wife and her children shall be her master's, and he shall go out alone.
EXOD|21|5|But if the slave plainly says, 'I love my master, my wife, and my children; I will not go out free,'
EXOD|21|6|then his master shall bring him to God, and he shall bring him to the door or the doorpost. And his master shall bore his ear through with an awl, and he shall be his slave forever.
EXOD|21|7|"When a man sells his daughter as a slave, she shall not go out as the male slaves do.
EXOD|21|8|If she does not please her master, who has designated her for himself, then he shall let her be redeemed. He shall have no right to sell her to a foreign people, since he has broken faith with her.
EXOD|21|9|If he designates her for his son, he shall deal with her as with a daughter.
EXOD|21|10|If he takes another wife to himself, he shall not diminish her food, her clothing, or her marital rights.
EXOD|21|11|And if he does not do these three things for her, she shall go out for nothing, without payment of money.
EXOD|21|12|"Whoever strikes a man so that he dies shall be put to death.
EXOD|21|13|But if he did not lie in wait for him, but God let him fall into his hand, then I will appoint for you a place to which he may flee.
EXOD|21|14|But if a man willfully attacks another to kill him by cunning, you shall take him from my altar, that he may die.
EXOD|21|15|"Whoever strikes his father or his mother shall be put to death.
EXOD|21|16|"Whoever steals a man and sells him, and anyone found in possession of him, shall be put to death.
EXOD|21|17|"Whoever curses his father or his mother shall be put to death.
EXOD|21|18|"When men quarrel and one strikes the other with a stone or with his fist and the man does not die but takes to his bed,
EXOD|21|19|then if the man rises again and walks outdoors with his staff, he who struck him shall be clear; only he shall pay for the loss of his time, and shall have him thoroughly healed.
EXOD|21|20|"When a man strikes his slave, male or female, with a rod and the slave dies under his hand, he shall be avenged.
EXOD|21|21|But if the slave survives a day or two, he is not to be avenged, for the slave is his money.
EXOD|21|22|"When men strive together and hit a pregnant woman, so that her children come out, but there is no harm, the one who hit her shall surely be fined, as the woman's husband shall impose on him, and he shall pay as the judges determine.
EXOD|21|23|But if there is harm, then you shall pay life for life,
EXOD|21|24|eye for eye, tooth for tooth, hand for hand, foot for foot,
EXOD|21|25|burn for burn, wound for wound, stripe for stripe.
EXOD|21|26|"When a man strikes the eye of his slave, male or female, and destroys it, he shall let the slave go free because of his eye.
EXOD|21|27|If he knocks out the tooth of his slave, male or female, he shall let the slave go free because of his tooth.
EXOD|21|28|"When an ox gores a man or a woman to death, the ox shall be stoned, and its flesh shall not be eaten, but the owner of the ox shall not be liable.
EXOD|21|29|But if the ox has been accustomed to gore in the past, and its owner has been warned but has not kept it in, and it kills a man or a woman, the ox shall be stoned, and its owner also shall be put to death.
EXOD|21|30|If a ransom is imposed on him, then he shall give for the redemption of his life whatever is imposed on him.
EXOD|21|31|If it gores a man's son or daughter, he shall be dealt with according to this same rule.
EXOD|21|32|If the ox gores a slave, male or female, the owner shall give to their master thirty shekels of silver, and the ox shall be stoned.
EXOD|21|33|"When a man opens a pit, or when a man digs a pit and does not cover it, and an ox or a donkey falls into it,
EXOD|21|34|the owner of the pit shall make restoration. He shall give money to its owner, and the dead beast shall be his.
EXOD|21|35|"When one man's ox butts another's, so that it dies, then they shall sell the live ox and share its price, and the dead beast also they shall share.
EXOD|21|36|Or if it is known that the ox has been accustomed to gore in the past, and its owner has not kept it in, he shall repay ox for ox, and the dead beast shall be his.
EXOD|22|1|"If a man steals an ox or a sheep, and kills it or sells it, he shall repay five oxen for an ox, and four sheep for a sheep.
EXOD|22|2|"If a thief is found breaking in and is struck so that he dies, there shall be no bloodguilt for him,
EXOD|22|3|but if the sun has risen on him, there shall be bloodguilt for him. He shall surely pay. If he has nothing, then he shall be sold for his theft.
EXOD|22|4|If the stolen beast is found alive in his possession, whether it is an ox or a donkey or a sheep, he shall pay double.
EXOD|22|5|"If a man causes a field or vineyard to be grazed over, or lets his beast loose and it feeds in another man's field, he shall make restitution from the best in his own field and in his own vineyard.
EXOD|22|6|"If fire breaks out and catches in thorns so that the stacked grain or the standing grain or the field is consumed, he who started the fire shall make full restitution.
EXOD|22|7|"If a man gives to his neighbor money or goods to keep safe, and it is stolen from the man's house, then, if the thief is found, he shall pay double.
EXOD|22|8|If the thief is not found, the owner of the house shall come near to God to show whether or not he has put his hand to his neighbor's property.
EXOD|22|9|For every breach of trust, whether it is for an ox, for a donkey, for a sheep, for a cloak, or for any kind of lost thing, of which one says, 'This is it,' the case of both parties shall come before God. The one whom God condemns shall pay double to his neighbor.
EXOD|22|10|"If a man gives to his neighbor a donkey or an ox or a sheep or any beast to keep safe, and it dies or is injured or is driven away, without anyone seeing it,
EXOD|22|11|an oath by the LORD shall be between them both to see whether or not he has put his hand to his neighbor's property. The owner shall accept the oath, and he shall not make restitution.
EXOD|22|12|But if it is stolen from him, he shall make restitution to its owner.
EXOD|22|13|If it is torn by beasts, let him bring it as evidence. He shall not make restitution for what has been torn.
EXOD|22|14|"If a man borrows anything of his neighbor, and it is injured or dies, the owner not being with it, he shall make full restitution.
EXOD|22|15|If the owner was with it, he shall not make restitution; if it was hired, it came for its hiring fee.
EXOD|22|16|"If a man seduces a virgin who is not engaged to be married and lies with her, he shall give the bride-price for her and make her his wife.
EXOD|22|17|If her father utterly refuses to give her to him, he shall pay money equal to the bride-price for virgins.
EXOD|22|18|"You shall not permit a sorceress to live.
EXOD|22|19|"Whoever lies with an animal shall be put to death.
EXOD|22|20|"Whoever sacrifices to any god, other than the LORD alone, shall be devoted to destruction.
EXOD|22|21|"You shall not wrong a sojourner or oppress him, for you were sojourners in the land of Egypt.
EXOD|22|22|You shall not mistreat any widow or fatherless child.
EXOD|22|23|If you do mistreat them, and they cry out to me, I will surely hear their cry,
EXOD|22|24|and my wrath will burn, and I will kill you with the sword, and your wives shall become widows and your children fatherless.
EXOD|22|25|"If you lend money to any of my people with you who is poor, you shall not be like a moneylender to him, and you shall not exact interest from him.
EXOD|22|26|If ever you take your neighbor's cloak in pledge, you shall return it to him before the sun goes down,
EXOD|22|27|for that is his only covering, and it is his cloak for his body; in what else shall he sleep? And if he cries to me, I will hear, for I am compassionate.
EXOD|22|28|"You shall not revile God, nor curse a ruler of your people.
EXOD|22|29|"You shall not delay to offer from the fullness of your harvest and from the outflow of your presses. The firstborn of your sons you shall give to me.
EXOD|22|30|You shall do the same with your oxen and with your sheep: seven days it shall be with its mother; on the eighth day you shall give it to me.
EXOD|22|31|"You shall be consecrated to me. Therefore you shall not eat any flesh that is torn by beasts in the field; you shall throw it to the dogs.
EXOD|23|1|"You shall not spread a false report. You shall not join hands with a wicked man to be a malicious witness.
EXOD|23|2|You shall not fall in with the many to do evil, nor shall you bear witness in a lawsuit, siding with the many, so as to pervert justice,
EXOD|23|3|nor shall you be partial to a poor man in his lawsuit.
EXOD|23|4|"If you meet your enemy's ox or his donkey going astray, you shall bring it back to him.
EXOD|23|5|If you see the donkey of one who hates you lying down under its burden, you shall refrain from leaving him with it; you shall rescue it with him.
EXOD|23|6|"You shall not pervert the justice due to your poor in his lawsuit.
EXOD|23|7|Keep far from a false charge, and do not kill the innocent and righteous, for I will not acquit the wicked.
EXOD|23|8|And you shall take no bribe, for a bribe blinds the clear-sighted and subverts the cause of those who are in the right.
EXOD|23|9|"You shall not oppress a sojourner. You know the heart of a sojourner, for you were sojourners in the land of Egypt.
EXOD|23|10|"For six years you shall sow your land and gather in its yield,
EXOD|23|11|but the seventh year you shall let it rest and lie fallow, that the poor of your people may eat; and what they leave the beasts of the field may eat. You shall do likewise with your vineyard, and with your olive orchard.
EXOD|23|12|"Six days you shall do your work, but on the seventh day you shall rest; that your ox and your donkey may have rest, and the son of your servant woman, and the alien, may be refreshed.
EXOD|23|13|"Pay attention to all that I have said to you, and make no mention of the names of other gods, nor let it be heard on your lips.
EXOD|23|14|"Three times in the year you shall keep a feast to me.
EXOD|23|15|You shall keep the Feast of Unleavened Bread. As I commanded you, you shall eat unleavened bread for seven days at the appointed time in the month of Abib, for in it you came out of Egypt. None shall appear before me empty-handed.
EXOD|23|16|You shall keep the Feast of Harvest, of the firstfruits of your labor, of what you sow in the field. You shall keep the Feast of Ingathering at the end of the year, when you gather in from the field the fruit of your labor.
EXOD|23|17|Three times in the year shall all your males appear before the Lord GOD.
EXOD|23|18|"You shall not offer the blood of my sacrifice with anything leavened, or let the fat of my feast remain until the morning.
EXOD|23|19|"The best of the firstfruits of your ground you shall bring into the house of the LORD your God. "You shall not boil a young goat in its mother's milk.
EXOD|23|20|"Behold, I send an angel before you to guard you on the way and to bring you to the place that I have prepared.
EXOD|23|21|Pay careful attention to him and obey his voice; do not rebel against him, for he will not pardon your transgression, for my name is in him.
EXOD|23|22|"But if you carefully obey his voice and do all that I say, then I will be an enemy to your enemies and an adversary to your adversaries.
EXOD|23|23|"When my angel goes before you and brings you to the Amorites and the Hittites and the Perizzites and the Canaanites, the Hivites and the Jebusites, and I blot them out,
EXOD|23|24|you shall not bow down to their gods nor serve them, nor do as they do, but you shall utterly overthrow them and break their pillars in pieces.
EXOD|23|25|You shall serve the LORD your God, and he will bless your bread and your water, and I will take sickness away from among you.
EXOD|23|26|None shall miscarry or be barren in your land; I will fulfill the number of your days.
EXOD|23|27|I will send my terror before you and will throw into confusion all the people against whom you shall come, and I will make all your enemies turn their backs to you.
EXOD|23|28|And I will send hornets before you, which shall drive out the Hivites, the Canaanites, and the Hittites from before you.
EXOD|23|29|I will not drive them out from before you in one year, lest the land become desolate and the wild beasts multiply against you.
EXOD|23|30|Little by little I will drive them out from before you, until you have increased and possess the land.
EXOD|23|31|And I will set your border from the Red Sea to the Sea of the Philistines, and from the wilderness to the Euphrates, for I will give the inhabitants of the land into your hand, and you shall drive them out before you.
EXOD|23|32|You shall make no covenant with them and their gods.
EXOD|23|33|They shall not dwell in your land, lest they make you sin against me; for if you serve their gods, it will surely be a snare to you."
EXOD|24|1|Then he said to Moses, "Come up to the LORD, you and Aaron, Nadab, and Abihu, and seventy of the elders of Israel, and worship from afar.
EXOD|24|2|Moses alone shall come near to the LORD, but the others shall not come near, and the people shall not come up with him."
EXOD|24|3|Moses came and told the people all the words of the LORD and all the rules. And all the people answered with one voice and said, "All the words that the LORD has spoken we will do."
EXOD|24|4|And Moses wrote down all the words of the LORD. He rose early in the morning and built an altar at the foot of the mountain, and twelve pillars, according to the twelve tribes of Israel.
EXOD|24|5|And he sent young men of the people of Israel, who offered burnt offerings and sacrificed peace offerings of oxen to the LORD.
EXOD|24|6|And Moses took half of the blood and put it in basins, and half of the blood he threw against the altar.
EXOD|24|7|Then he took the Book of the Covenant and read it in the hearing of the people. And they said, "All that the LORD has spoken we will do, and we will be obedient."
EXOD|24|8|And Moses took the blood and threw it on the people and said, "Behold the blood of the covenant that the LORD has made with you in accordance with all these words."
EXOD|24|9|Then Moses and Aaron, Nadab, and Abihu, and seventy of the elders of Israel went up,
EXOD|24|10|and they saw the God of Israel. There was under his feet as it were a pavement of sapphire stone, like the very heaven for clearness.
EXOD|24|11|And he did not lay his hand on the chief men of the people of Israel; they beheld God, and ate and drank.
EXOD|24|12|The LORD said to Moses, "Come up to me on the mountain and wait there, that I may give you the tablets of stone, with the law and the commandment, which I have written for their instruction."
EXOD|24|13|So Moses rose with his assistant Joshua, and Moses went up into the mountain of God.
EXOD|24|14|And he said to the elders, "Wait here for us until we return to you. And behold, Aaron and Hur are with you. Whoever has a dispute, let him go to them."
EXOD|24|15|Then Moses went up on the mountain, and the cloud covered the mountain.
EXOD|24|16|The glory of the LORD dwelt on Mount Sinai, and the cloud covered it six days. And on the seventh day he called to Moses out of the midst of the cloud.
EXOD|24|17|Now the appearance of the glory of the LORD was like a devouring fire on the top of the mountain in the sight of the people of Israel.
EXOD|24|18|Moses entered the cloud and went up on the mountain. And Moses was on the mountain forty days and forty nights.
EXOD|25|1|The LORD said to Moses,
EXOD|25|2|"Speak to the people of Israel, that they take for me a contribution. From every man whose heart moves him you shall receive the contribution for me.
EXOD|25|3|And this is the contribution that you shall receive from them: gold, silver, and bronze,
EXOD|25|4|blue and purple and scarlet yarns and fine twined linen, goats' hair,
EXOD|25|5|tanned rams' skins, goatskins, acacia wood,
EXOD|25|6|oil for the lamps, spices for the anointing oil and for the fragrant incense,
EXOD|25|7|onyx stones, and stones for setting, for the ephod and for the breastpiece.
EXOD|25|8|And let them make me a sanctuary, that I may dwell in their midst.
EXOD|25|9|Exactly as I show you concerning the pattern of the tabernacle, and of all its furniture, so you shall make it.
EXOD|25|10|"They shall make an ark of acacia wood. Two cubits and a half shall be its length, a cubit and a half its breadth, and a cubit and a half its height.
EXOD|25|11|You shall overlay it with pure gold, inside and outside shall you overlay it, and you shall make on it a molding of gold around it.
EXOD|25|12|You shall cast four rings of gold for it and put them on its four feet, two rings on the one side of it, and two rings on the other side of it.
EXOD|25|13|You shall make poles of acacia wood and overlay them with gold.
EXOD|25|14|And you shall put the poles into the rings on the sides of the ark to carry the ark by them.
EXOD|25|15|The poles shall remain in the rings of the ark; they shall not be taken from it.
EXOD|25|16|And you shall put into the ark the testimony that I shall give you.
EXOD|25|17|"You shall make a mercy seat of pure gold. Two cubits and a half shall be its length, and a cubit and a half its breadth.
EXOD|25|18|And you shall make two cherubim of gold; of hammered work shall you make them, on the two ends of the mercy seat.
EXOD|25|19|Make one cherub on the one end, and one cherub on the other end. Of one piece with the mercy seat shall you make the cherubim on its two ends.
EXOD|25|20|The cherubim shall spread out their wings above, overshadowing the mercy seat with their wings, their faces one to another; toward the mercy seat shall the faces of the cherubim be.
EXOD|25|21|And you shall put the mercy seat on the top of the ark, and in the ark you shall put the testimony that I shall give you.
EXOD|25|22|There I will meet with you, and from above the mercy seat, from between the two cherubim that are on the ark of the testimony, I will speak with you about all that I will give you in commandment for the people of Israel.
EXOD|25|23|"You shall make a table of acacia wood. Two cubits shall be its length, a cubit its breadth, and a cubit and a half its height.
EXOD|25|24|You shall overlay it with pure gold and make a molding of gold around it.
EXOD|25|25|And you shall make a rim around it a handbreadth wide, and a molding of gold around the rim.
EXOD|25|26|And you shall make for it four rings of gold, and fasten the rings to the four corners at its four legs.
EXOD|25|27|Close to the frame the rings shall lie, as holders for the poles to carry the table.
EXOD|25|28|You shall make the poles of acacia wood, and overlay them with gold, and the table shall be carried with these.
EXOD|25|29|And you shall make its plates and dishes for incense, and its flagons and bowls with which to pour drink offerings; you shall make them of pure gold.
EXOD|25|30|And you shall set the bread of the Presence on the table before me regularly.
EXOD|25|31|"You shall make a lampstand of pure gold. The lampstand shall be made of hammered work: its base, its stem, its cups, its calyxes, and its flowers shall be of one piece with it.
EXOD|25|32|And there shall be six branches going out of its sides, three branches of the lampstand out of one side of it and three branches of the lampstand out of the other side of it;
EXOD|25|33|three cups made like almond blossoms, each with calyx and flower, on one branch, and three cups made like almond blossoms, each with calyx and flower, on the other branch- so for the six branches going out of the lampstand.
EXOD|25|34|And on the lampstand itself there shall be four cups made like almond blossoms, with their calyxes and flowers,
EXOD|25|35|and a calyx of one piece with it under each pair of the six branches going out from the lampstand.
EXOD|25|36|Their calyxes and their branches shall be of one piece with it, the whole of it a single piece of hammered work of pure gold.
EXOD|25|37|You shall make seven lamps for it. And the lamps shall be set up so as to give light on the space in front of it.
EXOD|25|38|Its tongs and their trays shall be of pure gold.
EXOD|25|39|It shall be made, with all these utensils, out of a talent of pure gold.
EXOD|25|40|And see that you make them after the pattern for them, which is being shown you on the mountain.
EXOD|26|1|"Moreover, you shall make the tabernacle with ten curtains of fine twined linen and blue and purple and scarlet yarns; you shall make them with cherubim skillfully worked into them.
EXOD|26|2|The length of each curtain shall be twenty-eight cubits, and the breadth of each curtain four cubits; all the curtains shall be the same size.
EXOD|26|3|Five curtains shall be coupled to one another, and the other five curtains shall be coupled to one another.
EXOD|26|4|And you shall make loops of blue on the edge of the outermost curtain in the first set. Likewise you shall make loops on the edge of the outermost curtain in the second set.
EXOD|26|5|Fifty loops you shall make on the one curtain, and fifty loops you shall make on the edge of the curtain that is in the second set; the loops shall be opposite one another.
EXOD|26|6|And you shall make fifty clasps of gold, and couple the curtains one to the other with the clasps, so that the tabernacle may be a single whole.
EXOD|26|7|"You shall also make curtains of goats' hair for a tent over the tabernacle; eleven curtains shall you make.
EXOD|26|8|The length of each curtain shall be thirty cubits, and the breadth of each curtain four cubits. The eleven curtains shall be the same size.
EXOD|26|9|You shall couple five curtains by themselves, and six curtains by themselves, and the sixth curtain you shall double over at the front of the tent.
EXOD|26|10|You shall make fifty loops on the edge of the curtain that is outermost in one set, and fifty loops on the edge of the curtain that is outermost in the second set.
EXOD|26|11|"You shall make fifty clasps of bronze, and put the clasps into the loops, and couple the tent together that it may be a single whole.
EXOD|26|12|And the part that remains of the curtains of the tent, the half curtain that remains, shall hang over the back of the tabernacle.
EXOD|26|13|And the extra that remains in the length of the curtains, the cubit on the one side, and the cubit on the other side, shall hang over the sides of the tabernacle, on this side and that side, to cover it.
EXOD|26|14|And you shall make for the tent a covering of tanned rams' skins and a covering of goatskins on top.
EXOD|26|15|"You shall make upright frames for the tabernacle of acacia wood.
EXOD|26|16|Ten cubits shall be the length of a frame, and a cubit and a half the breadth of each frame.
EXOD|26|17|There shall be two tenons in each frame, for fitting together. So shall you do for all the frames of the tabernacle.
EXOD|26|18|You shall make the frames for the tabernacle: twenty frames for the south side;
EXOD|26|19|and forty bases of silver you shall make under the twenty frames, two bases under one frame for its two tenons, and two bases under the next frame for its two tenons;
EXOD|26|20|and for the second side of the tabernacle, on the north side twenty frames,
EXOD|26|21|and their forty bases of silver, two bases under one frame, and two bases under the next frame.
EXOD|26|22|And for the rear of the tabernacle westward you shall make six frames.
EXOD|26|23|And you shall make two frames for corners of the tabernacle in the rear;
EXOD|26|24|they shall be separate beneath, but joined at the top, at the first ring. Thus shall it be with both of them; they shall form the two corners.
EXOD|26|25|And there shall be eight frames, with their bases of silver, sixteen bases; two bases under one frame, and two bases under another frame.
EXOD|26|26|"You shall make bars of acacia wood, five for the frames of the one side of the tabernacle,
EXOD|26|27|and five bars for the frames of the other side of the tabernacle, and five bars for the frames of the side of the tabernacle at the rear westward.
EXOD|26|28|The middle bar, halfway up the frames, shall run from end to end.
EXOD|26|29|You shall overlay the frames with gold and shall make their rings of gold for holders for the bars, and you shall overlay the bars with gold.
EXOD|26|30|Then you shall erect the tabernacle according to the plan for it that you were shown on the mountain.
EXOD|26|31|"And you shall make a veil of blue and purple and scarlet yarns and fine twined linen. It shall be made with cherubim skillfully worked into it.
EXOD|26|32|And you shall hang it on four pillars of acacia overlaid with gold, with hooks of gold, on four bases of silver.
EXOD|26|33|And you shall hang the veil from the clasps, and bring the ark of the testimony in there within the veil. And the veil shall separate for you the Holy Place from the Most Holy.
EXOD|26|34|You shall put the mercy seat on the ark of the testimony in the Most Holy Place.
EXOD|26|35|And you shall set the table outside the veil, and the lampstand on the south side of the tabernacle opposite the table, and you shall put the table on the north side.
EXOD|26|36|"You shall make a screen for the entrance of the tent, of blue and purple and scarlet yarns and fine twined linen, embroidered with needlework.
EXOD|26|37|And you shall make for the screen five pillars of acacia, and overlay them with gold. Their hooks shall be of gold, and you shall cast five bases of bronze for them.
EXOD|27|1|"You shall make the altar of acacia wood, five cubits long and five cubits broad. The altar shall be square, and its height shall be three cubits.
EXOD|27|2|And you shall make horns for it on its four corners; its horns shall be of one piece with it, and you shall overlay it with bronze.
EXOD|27|3|You shall make pots for it to receive its ashes, and shovels and basins and forks and fire pans. You shall make all its utensils of bronze.
EXOD|27|4|You shall also make for it a grating, a network of bronze, and on the net you shall make four bronze rings at its four corners.
EXOD|27|5|And you shall set it under the ledge of the altar so that the net extends halfway down the altar.
EXOD|27|6|And you shall make poles for the altar, poles of acacia wood, and overlay them with bronze.
EXOD|27|7|And the poles shall be put through the rings, so that the poles are on the two sides of the altar when it is carried.
EXOD|27|8|You shall make it hollow, with boards. As it has been shown you on the mountain, so shall it be made.
EXOD|27|9|"You shall make the court of the tabernacle. On the south side the court shall have hangings of fine twined linen a hundred cubits long for one side.
EXOD|27|10|Its twenty pillars and their twenty bases shall be of bronze, but the hooks of the pillars and their fillets shall be of silver.
EXOD|27|11|And likewise for its length on the north side there shall be hangings a hundred cubits long, its pillars twenty and their bases twenty, of bronze, but the hooks of the pillars and their fillets shall be of silver.
EXOD|27|12|And for the breadth of the court on the west side there shall be hangings for fifty cubits, with ten pillars and ten bases.
EXOD|27|13|The breadth of the court on the front to the east shall be fifty cubits.
EXOD|27|14|The hangings for the one side of the gate shall be fifteen cubits, with their three pillars and three bases.
EXOD|27|15|On the other side the hangings shall be fifteen cubits, with their three pillars and three bases.
EXOD|27|16|For the gate of the court there shall be a screen twenty cubits long, of blue and purple and scarlet yarns and fine twined linen, embroidered with needlework. It shall have four pillars and with them four bases.
EXOD|27|17|All the pillars around the court shall be filleted with silver. Their hooks shall be of silver, and their bases of bronze.
EXOD|27|18|The length of the court shall be a hundred cubits, the breadth fifty, and the height five cubits, with hangings of fine twined linen and bases of bronze.
EXOD|27|19|All the utensils of the tabernacle for every use, and all its pegs and all the pegs of the court, shall be of bronze.
EXOD|27|20|"You shall command the people of Israel that they bring to you pure beaten olive oil for the light, that a lamp may regularly be set up to burn.
EXOD|27|21|In the tent of meeting, outside the veil that is before the testimony, Aaron and his sons shall tend it from evening to morning before the LORD. It shall be a statute forever to be observed throughout their generations by the people of Israel.
EXOD|28|1|"Then bring near to you Aaron your brother, and his sons with him, from among the people of Israel, to serve me as priests- Aaron and Aaron's sons, Nadab and Abihu, Eleazar and Ithamar.
EXOD|28|2|And you shall make holy garments for Aaron your brother, for glory and for beauty.
EXOD|28|3|You shall speak to all the skillful, whom I have filled with a spirit of skill, that they make Aaron's garments to consecrate him for my priesthood.
EXOD|28|4|These are the garments that they shall make: a breastpiece, an ephod, a robe, a coat of checker work, a turban, and a sash. They shall make holy garments for Aaron your brother and his sons to serve me as priests.
EXOD|28|5|They shall receive gold, blue and purple and scarlet yarns, and fine twined linen.
EXOD|28|6|"And they shall make the ephod of gold, of blue and purple and scarlet yarns, and of fine twined linen, skillfully worked.
EXOD|28|7|It shall have two shoulder pieces attached to its two edges, so that it may be joined together.
EXOD|28|8|And the skillfully woven band on it shall be made like it and be of one piece with it, of gold, blue and purple and scarlet yarns, and fine twined linen.
EXOD|28|9|You shall take two onyx stones, and engrave on them the names of the sons of Israel,
EXOD|28|10|six of their names on the one stone, and the names of the remaining six on the other stone, in the order of their birth.
EXOD|28|11|As a jeweler engraves signets, so shall you engrave the two stones with the names of the sons of Israel. You shall enclose them in settings of gold filigree.
EXOD|28|12|And you shall set the two stones on the shoulder pieces of the ephod, as stones of remembrance for the sons of Israel. And Aaron shall bear their names before the LORD on his two shoulders for remembrance.
EXOD|28|13|You shall make settings of gold filigree,
EXOD|28|14|and two chains of pure gold, twisted like cords; and you shall attach the corded chains to the settings.
EXOD|28|15|"You shall make a breastpiece of judgment, in skilled work. In the style of the ephod you shall make it- of gold, blue and purple and scarlet yarns, and fine twined linen shall you make it.
EXOD|28|16|It shall be square and doubled, a span its length and a span its breadth.
EXOD|28|17|You shall set in it four rows of stones. A row of sardius, topaz, and carbuncle shall be the first row;
EXOD|28|18|and the second row an emerald, a sapphire, and a diamond;
EXOD|28|19|and the third row a jacinth, an agate, and an amethyst;
EXOD|28|20|and the fourth row a beryl, an onyx, and a jasper. They shall be set in gold filigree.
EXOD|28|21|There shall be twelve stones with their names according to the names of the sons of Israel. They shall be like signets, each engraved with its name, for the twelve tribes.
EXOD|28|22|You shall make for the breastpiece twisted chains like cords, of pure gold.
EXOD|28|23|And you shall make for the breastpiece two rings of gold, and put the two rings on the two edges of the breastpiece.
EXOD|28|24|And you shall put the two cords of gold in the two rings at the edges of the breastpiece.
EXOD|28|25|The two ends of the two cords you shall attach to the two settings of filigree, and so attach it in front to the shoulder pieces of the ephod.
EXOD|28|26|You shall make two rings of gold, and put them at the two ends of the breastpiece, on its inside edge next to the ephod.
EXOD|28|27|And you shall make two rings of gold, and attach them in front to the lower part of the two shoulder pieces of the ephod, at its seam above the skillfully woven band of the ephod.
EXOD|28|28|And they shall bind the breastpiece by its rings to the rings of the ephod with a lace of blue, so that it may lie on the skillfully woven band of the ephod, so that the breastpiece shall not come loose from the ephod.
EXOD|28|29|So Aaron shall bear the names of the sons of Israel in the breastpiece of judgment on his heart, when he goes into the Holy Place, to bring them to regular remembrance before the LORD.
EXOD|28|30|And in the breastpiece of judgment you shall put the Urim and the Thummim, and they shall be on Aaron's heart, when he goes in before the LORD. Thus Aaron shall bear the judgment of the people of Israel on his heart before the LORD regularly.
EXOD|28|31|"You shall make the robe of the ephod all of blue.
EXOD|28|32|It shall have an opening for the head in the middle of it, with a woven binding around the opening, like the opening in a garment, so that it may not tear.
EXOD|28|33|On its hem you shall make pomegranates of blue and purple and scarlet yarns, around its hem, with bells of gold between them,
EXOD|28|34|a golden bell and a pomegranate, a golden bell and a pomegranate, around the hem of the robe.
EXOD|28|35|And it shall be on Aaron when he ministers, and its sound shall be heard when he goes into the Holy Place before the LORD, and when he comes out, so that he does not die.
EXOD|28|36|"You shall make a plate of pure gold and engrave on it, like the engraving of a signet, 'Holy to the LORD.'
EXOD|28|37|And you shall fasten it on the turban by a cord of blue. It shall be on the front of the turban.
EXOD|28|38|It shall be on Aaron's forehead, and Aaron shall bear any guilt from the holy things that the people of Israel consecrate as their holy gifts. It shall regularly be on his forehead, that they may be accepted before the LORD.
EXOD|28|39|"You shall weave the coat in checker work of fine linen, and you shall make a turban of fine linen, and you shall make a sash embroidered with needlework.
EXOD|28|40|"For Aaron's sons you shall make coats and sashes and caps. You shall make them for glory and beauty.
EXOD|28|41|And you shall put them on Aaron your brother, and on his sons with him, and shall anoint them and ordain them and consecrate them, that they may serve me as priests.
EXOD|28|42|You shall make for them linen undergarments to cover their naked flesh. They shall reach from the hips to the thighs;
EXOD|28|43|and they shall be on Aaron and on his sons when they go into the tent of meeting or when they come near the altar to minister in the Holy Place, lest they bear guilt and die. This shall be a statute forever for him and for his offspring after him.
EXOD|29|1|"Now this is what you shall do to them to consecrate them, that they may serve me as priests. Take one bull of the herd and two rams without blemish,
EXOD|29|2|and unleavened bread, unleavened cakes mixed with oil, and unleavened wafers smeared with oil. You shall make them of fine wheat flour.
EXOD|29|3|You shall put them in one basket and bring them in the basket, and bring the bull and the two rams.
EXOD|29|4|You shall bring Aaron and his sons to the entrance of the tent of meeting and wash them with water.
EXOD|29|5|Then you shall take the garments, and put on Aaron the coat and the robe of the ephod, and the ephod, and the breastpiece, and gird him with the skillfully woven band of the ephod.
EXOD|29|6|And you shall set the turban on his head and put the holy crown on the turban.
EXOD|29|7|You shall take the anointing oil and pour it on his head and anoint him.
EXOD|29|8|Then you shall bring his sons and put coats on them,
EXOD|29|9|and you shall gird Aaron and his sons with sashes and bind caps on them. And the priesthood shall be theirs by a statute forever. Thus you shall ordain Aaron and his sons.
EXOD|29|10|"Then you shall bring the bull before the tent of meeting. Aaron and his sons shall lay their hands on the head of the bull.
EXOD|29|11|Then you shall kill the bull before the LORD at the entrance of the tent of meeting,
EXOD|29|12|and shall take part of the blood of the bull and put it on the horns of the altar with your finger, and the rest of the blood you shall pour out at the base of the altar.
EXOD|29|13|And you shall take all the fat that covers the entrails, and the long lobe of the liver, and the two kidneys with the fat that is on them, and burn them on the altar.
EXOD|29|14|But the flesh of the bull and its skin and its dung you shall burn with fire outside the camp; it is a sin offering.
EXOD|29|15|"Then you shall take one of the rams, and Aaron and his sons shall lay their hands on the head of the ram,
EXOD|29|16|and you shall kill the ram and shall take its blood and throw it against the sides of the altar.
EXOD|29|17|Then you shall cut the ram into pieces, and wash its entrails and its legs, and put them with its pieces and its head,
EXOD|29|18|and burn the whole ram on the altar. It is a burnt offering to the LORD. It is a pleasing aroma, a food offering to the LORD.
EXOD|29|19|"You shall take the other ram, and Aaron and his sons shall lay their hands on the head of the ram,
EXOD|29|20|and you shall kill the ram and take part of its blood and put it on the tip of the right ear of Aaron and on the tips of the right ears of his sons, and on the thumbs of their right hands and on the great toes of their right feet, and throw the rest of the blood against the sides of the altar.
EXOD|29|21|Then you shall take part of the blood that is on the altar, and of the anointing oil, and sprinkle it on Aaron and his garments, and on his sons and his sons' garments with him. He and his garments shall be holy, and his sons and his sons' garments with him.
EXOD|29|22|"You shall also take the fat from the ram and the fat tail and the fat that covers the entrails, and the long lobe of the liver and the two kidneys with the fat that is on them, and the right thigh (for it is a ram of ordination),
EXOD|29|23|and one loaf of bread and one cake of bread made with oil, and one wafer out of the basket of unleavened bread that is before the LORD.
EXOD|29|24|You shall put all these on the palms of Aaron and on the palms of his sons, and wave them for a wave offering before the LORD.
EXOD|29|25|Then you shall take them from their hands and burn them on the altar on top of the burnt offering, as a pleasing aroma before the LORD. It is a food offering to the LORD.
EXOD|29|26|"You shall take the breast of the ram of Aaron's ordination and wave it for a wave offering before the LORD, and it shall be your portion.
EXOD|29|27|And you shall consecrate the breast of the wave offering that is waved and the thigh of the priests' portion that is contributed from the ram of ordination, from what was Aaron's and his sons.
EXOD|29|28|It shall be for Aaron and his sons as a perpetual due from the people of Israel, for it is a contribution. It shall be a contribution from the people of Israel from their peace offerings, their contribution to the LORD.
EXOD|29|29|"The holy garments of Aaron shall be for his sons after him; they shall be anointed in them and ordained in them.
EXOD|29|30|The son who succeeds him as priest, who comes into the tent of meeting to minister in the Holy Place, shall wear them seven days.
EXOD|29|31|"You shall take the ram of ordination and boil its flesh in a holy place.
EXOD|29|32|And Aaron and his sons shall eat the flesh of the ram and the bread that is in the basket in the entrance of the tent of meeting.
EXOD|29|33|They shall eat those things with which atonement was made at their ordination and consecration, but an outsider shall not eat of them, because they are holy.
EXOD|29|34|And if any of the flesh for the ordination or of the bread remain until the morning, then you shall burn the remainder with fire. It shall not be eaten, because it is holy.
EXOD|29|35|"Thus you shall do to Aaron and to his sons, according to all that I have commanded you. Through seven days shall you ordain them,
EXOD|29|36|and every day you shall offer a bull as a sin offering for atonement. Also you shall purify the altar, when you make atonement for it, and shall anoint it to consecrate it.
EXOD|29|37|Seven days you shall make atonement for the altar and consecrate it, and the altar shall be most holy. Whatever touches the altar shall become holy.
EXOD|29|38|"Now this is what you shall offer on the altar: two lambs a year old day by day regularly.
EXOD|29|39|One lamb you shall offer in the morning, and the other lamb you shall offer at twilight.
EXOD|29|40|And with the first lamb a tenth seah of fine flour mingled with a fourth of a hin of beaten oil, and a fourth of a hin of wine for a drink offering.
EXOD|29|41|The other lamb you shall offer at twilight, and shall offer with it a grain offering and its drink offering, as in the morning, for a pleasing aroma, a food offering to the LORD.
EXOD|29|42|It shall be a regular burnt offering throughout your generations at the entrance of the tent of meeting before the LORD, where I will meet with you, to speak to you there.
EXOD|29|43|There I will meet with the people of Israel, and it shall be sanctified by my glory.
EXOD|29|44|I will consecrate the tent of meeting and the altar. Aaron also and his sons I will consecrate to serve me as priests.
EXOD|29|45|I will dwell among the people of Israel and will be their God.
EXOD|29|46|And they shall know that I am the LORD their God, who brought them out of the land of Egypt that I might dwell among them. I am the LORD their God.
EXOD|30|1|"You shall make an altar on which to burn incense; you shall make it of acacia wood.
EXOD|30|2|A cubit shall be its length, and a cubit its breadth. It shall be square, and two cubits shall be its height. Its horns shall be of one piece with it.
EXOD|30|3|You shall overlay it with pure gold, its top and around its sides and its horns. And you shall make a molding of gold around it.
EXOD|30|4|And you shall make two golden rings for it. Under its molding on two opposite sides of it you shall make them, and they shall be holders for poles with which to carry it.
EXOD|30|5|You shall make the poles of acacia wood and overlay them with gold.
EXOD|30|6|And you shall put it in front of the veil that is above the ark of the testimony, in front of the mercy seat that is above the testimony, where I will meet with you.
EXOD|30|7|And Aaron shall burn fragrant incense on it. Every morning when he dresses the lamps he shall burn it,
EXOD|30|8|and when Aaron sets up the lamps at twilight, he shall burn it, a regular incense offering before the LORD throughout your generations.
EXOD|30|9|You shall not offer unauthorized incense on it, or a burnt offering, or a grain offering, and you shall not pour a drink offering on it.
EXOD|30|10|Aaron shall make atonement on its horns once a year. With the blood of the sin offering of atonement he shall make atonement for it once in the year throughout your generations. It is most holy to the LORD."
EXOD|30|11|The LORD said to Moses,
EXOD|30|12|"When you take the census of the people of Israel, then each shall give a ransom for his life to the LORD when you number them, that there be no plague among them when you number them.
EXOD|30|13|Each one who is numbered in the census shall give this: half a shekel according to the shekel of the sanctuary (the shekel is twenty gerahs), half a shekel as an offering to the LORD.
EXOD|30|14|Everyone who is numbered in the census, from twenty years old and upward, shall give the LORD's offering.
EXOD|30|15|The rich shall not give more, and the poor shall not give less, than the half shekel, when you give the LORD's offering to make atonement for your lives.
EXOD|30|16|You shall take the atonement money from the people of Israel and shall give it for the service of the tent of meeting, that it may bring the people of Israel to remembrance before the LORD, so as to make atonement for your lives."
EXOD|30|17|The LORD said to Moses,
EXOD|30|18|"You shall also make a basin of bronze, with its stand of bronze, for washing. You shall put it between the tent of meeting and the altar, and you shall put water in it,
EXOD|30|19|with which Aaron and his sons shall wash their hands and their feet.
EXOD|30|20|When they go into the tent of meeting, or when they come near the altar to minister, to burn a food offering to the LORD, they shall wash with water, so that they may not die.
EXOD|30|21|They shall wash their hands and their feet, so that they may not die. It shall be a statute forever to them, even to him and to his offspring throughout their generations."
EXOD|30|22|The LORD said to Moses,
EXOD|30|23|"Take the finest spices: of liquid myrrh 500 shekels, and of sweet-smelling cinnamon half as much, that is, 250, and 250 of aromatic cane,
EXOD|30|24|and 500 of cassia, according to the shekel of the sanctuary, and a hin of olive oil.
EXOD|30|25|And you shall make of these a sacred anointing oil blended as by the perfumer; it shall be a holy anointing oil.
EXOD|30|26|With it you shall anoint the tent of meeting and the ark of the testimony,
EXOD|30|27|and the table and all its utensils, and the lampstand and its utensils, and the altar of incense,
EXOD|30|28|and the altar of burnt offering with all its utensils and the basin and its stand.
EXOD|30|29|You shall consecrate them, that they may be most holy. Whatever touches them will become holy.
EXOD|30|30|You shall anoint Aaron and his sons, and consecrate them, that they may serve me as priests.
EXOD|30|31|And you shall say to the people of Israel, 'This shall be my holy anointing oil throughout your generations.
EXOD|30|32|It shall not be poured on the body of an ordinary person, and you shall make no other like it in composition. It is holy, and it shall be holy to you.
EXOD|30|33|Whoever compounds any like it or whoever puts any of it on an outsider shall be cut off from his people.'"
EXOD|30|34|The LORD said to Moses, "Take sweet spices, stacte, and onycha, and galbanum, sweet spices with pure frankincense (of each shall there be an equal part),
EXOD|30|35|and make an incense blended as by the perfumer, seasoned with salt, pure and holy.
EXOD|30|36|You shall beat some of it very small, and put part of it before the testimony in the tent of meeting where I shall meet with you. It shall be most holy for you.
EXOD|30|37|And the incense that you shall make according to its composition, you shall not make for yourselves. It shall be for you holy to the LORD.
EXOD|30|38|Whoever makes any like it to use as perfume shall be cut off from his people."
EXOD|31|1|The LORD said to Moses,
EXOD|31|2|"See, I have called by name Bezalel the son of Uri, son of Hur, of the tribe of Judah,
EXOD|31|3|and I have filled him with the Spirit of God, with ability and intelligence, with knowledge and all craftsmanship,
EXOD|31|4|to devise artistic designs, to work in gold, silver, and bronze,
EXOD|31|5|in cutting stones for setting, and in carving wood, to work in every craft.
EXOD|31|6|And behold, I have appointed with him Oholiab, the son of Ahisamach, of the tribe of Dan. And I have given to all able men ability, that they may make all that I have commanded you:
EXOD|31|7|the tent of meeting, and the ark of the testimony, and the mercy seat that is on it, and all the furnishings of the tent,
EXOD|31|8|the table and its utensils, and the pure lampstand with all its utensils, and the altar of incense,
EXOD|31|9|and the altar of burnt offering with all its utensils, and the basin and its stand,
EXOD|31|10|and the finely worked garments, the holy garments for Aaron the priest and the garments of his sons, for their service as priests,
EXOD|31|11|and the anointing oil and the fragrant incense for the Holy Place. According to all that I have commanded you, they shall do."
EXOD|31|12|And the LORD said to Moses,
EXOD|31|13|"You are to speak to the people of Israel and say, 'Above all you shall keep my Sabbaths, for this is a sign between me and you throughout your generations, that you may know that I, the LORD, sanctify you.
EXOD|31|14|You shall keep the Sabbath, because it is holy for you. Everyone who profanes it shall be put to death. Whoever does any work on it, that soul shall be cut off from among his people.
EXOD|31|15|Six days shall work be done, but the seventh day is a Sabbath of solemn rest, holy to the LORD. Whoever does any work on the Sabbath day shall be put to death.
EXOD|31|16|Therefore the people of Israel shall keep the Sabbath, observing the Sabbath throughout their generations, as a covenant forever.
EXOD|31|17|It is a sign forever between me and the people of Israel that in six days the LORD made heaven and earth, and on the seventh day he rested and was refreshed.'"
EXOD|31|18|And he gave to Moses, when he had finished speaking with him on Mount Sinai, the two tablets of the testimony, tablets of stone, written with the finger of God.
EXOD|32|1|When the people saw that Moses delayed to come down from the mountain, the people gathered themselves together to Aaron and said to him, "Up, make us gods who shall go before us. As for this Moses, the man who brought us up out of the land of Egypt, we do not know what has become of him."
EXOD|32|2|So Aaron said to them, "Take off the rings of gold that are in the ears of your wives, your sons, and your daughters, and bring them to me."
EXOD|32|3|So all the people took off the rings of gold that were in their ears and brought them to Aaron.
EXOD|32|4|And he received the gold from their hand and fashioned it with a graving tool and made a golden calf. And they said, "These are your gods, O Israel, who brought you up out of the land of Egypt!"
EXOD|32|5|When Aaron saw this, he built an altar before it. And Aaron made proclamation and said, "Tomorrow shall be a feast to the LORD."
EXOD|32|6|And they rose up early the next day and offered burnt offerings and brought peace offerings. And the people sat down to eat and drink and rose up to play.
EXOD|32|7|And the LORD said to Moses, "Go down, for your people, whom you brought up out of the land of Egypt, have corrupted themselves.
EXOD|32|8|They have turned aside quickly out of the way that I commanded them. They have made for themselves a golden calf and have worshiped it and sacrificed to it and said, 'These are your gods, O Israel, who brought you up out of the land of Egypt!'"
EXOD|32|9|And the LORD said to Moses, "I have seen this people, and behold, it is a stiff-necked people.
EXOD|32|10|Now therefore let me alone, that my wrath may burn hot against them and I may consume them, in order that I may make a great nation of you."
EXOD|32|11|But Moses implored the LORD his God and said, "O LORD, why does your wrath burn hot against your people, whom you have brought out of the land of Egypt with great power and with a mighty hand?
EXOD|32|12|Why should the Egyptians say, 'With evil intent did he bring them out, to kill them in the mountains and to consume them from the face of the earth'? Turn from your burning anger and relent from this disaster against your people.
EXOD|32|13|Remember Abraham, Isaac, and Israel, your servants, to whom you swore by your own self, and said to them, 'I will multiply your offspring as the stars of heaven, and all this land that I have promised I will give to your offspring, and they shall inherit it forever.'"
EXOD|32|14|And the LORD relented from the disaster that he had spoken of bringing on his people.
EXOD|32|15|Then Moses turned and went down from the mountain with the two tablets of the testimony in his hand, tablets that were written on both sides; on the front and on the back they were written.
EXOD|32|16|The tablets were the work of God, and the writing was the writing of God, engraved on the tablets.
EXOD|32|17|When Joshua heard the noise of the people as they shouted, he said to Moses, "There is a noise of war in the camp."
EXOD|32|18|But he said, "It is not the sound of shouting for victory, or the sound of the cry of defeat, but the sound of singing that I hear."
EXOD|32|19|And as soon as he came near the camp and saw the calf and the dancing, Moses' anger burned hot, and he threw the tablets out of his hands and broke them at the foot of the mountain.
EXOD|32|20|He took the calf that they had made and burned it with fire and ground it to powder and scattered it on the water and made the people of Israel drink it.
EXOD|32|21|And Moses said to Aaron, "What did this people do to you that you have brought such a great sin upon them?"
EXOD|32|22|And Aaron said, "Let not the anger of my lord burn hot. You know the people, that they are set on evil.
EXOD|32|23|For they said to me, 'Make us gods who shall go before us. As for this Moses, the man who brought us up out of the land of Egypt, we do not know what has become of him.'
EXOD|32|24|So I said to them, 'Let any who have gold take it off.' So they gave it to me, and I threw it into the fire, and out came this calf."
EXOD|32|25|And when Moses saw that the people had broken loose (for Aaron had let them break loose, to the derision of their enemies),
EXOD|32|26|then Moses stood in the gate of the camp and said, "Who is on the LORD's side? Come to me." And all the sons of Levi gathered around him.
EXOD|32|27|And he said to them, "Thus says the LORD God of Israel, 'Put your sword on your side each of you, and go to and fro from gate to gate throughout the camp, and each of you kill his brother and his companion and his neighbor.'"
EXOD|32|28|And the sons of Levi did according to the word of Moses. And that day about three thousand men of the people fell.
EXOD|32|29|And Moses said, "Today you have been ordained for the service of the LORD, each one at the cost of his son and of his brother, so that he might bestow a blessing upon you this day."
EXOD|32|30|The next day Moses said to the people, "You have sinned a great sin. And now I will go up to the LORD; perhaps I can make atonement for your sin."
EXOD|32|31|So Moses returned to the LORD and said, "Alas, this people have sinned a great sin. They have made for themselves gods of gold.
EXOD|32|32|But now, if you will forgive their sin- but if not, please blot me out of your book that you have written."
EXOD|32|33|But the LORD said to Moses, "Whoever has sinned against me, I will blot out of my book.
EXOD|32|34|But now go, lead the people to the place about which I have spoken to you; behold, my angel shall go before you. Nevertheless, in the day when I visit, I will visit their sin upon them."
EXOD|32|35|Then the LORD sent a plague on the people, because they made the calf, the one that Aaron made.
EXOD|33|1|The LORD said to Moses, "Depart; go up from here, you and the people whom you have brought up out of the land of Egypt, to the land of which I swore to Abraham, Isaac, and Jacob, saying, 'To your offspring I will give it.'
EXOD|33|2|I will send an angel before you, and I will drive out the Canaanites, the Amorites, the Hittites, the Perizzites, the Hivites, and the Jebusites.
EXOD|33|3|Go up to a land flowing with milk and honey; but I will not go up among you, lest I consume you on the way, for you are a stiff-necked people."
EXOD|33|4|When the people heard this disastrous word, they mourned, and no one put on his ornaments.
EXOD|33|5|For the LORD had said to Moses, "Say to the people of Israel, 'You are a stiff-necked people; if for a single moment I should go up among you, I would consume you. So now take off your ornaments, that I may know what to do with you.'"
EXOD|33|6|Therefore the people of Israel stripped themselves of their ornaments, from Mount Horeb onward.
EXOD|33|7|Now Moses used to take the tent and pitch it outside the camp, far off from the camp, and he called it the tent of meeting. And everyone who sought the LORD would go out to the tent of meeting, which was outside the camp.
EXOD|33|8|Whenever Moses went out to the tent, all the people would rise up, and each would stand at his tent door, and watch Moses until he had gone into the tent.
EXOD|33|9|When Moses entered the tent, the pillar of cloud would descend and stand at the entrance of the tent, and the LORD would speak with Moses.
EXOD|33|10|And when all the people saw the pillar of cloud standing at the entrance of the tent, all the people would rise up and worship, each at his tent door.
EXOD|33|11|Thus the LORD used to speak to Moses face to face, as a man speaks to his friend. When Moses turned again into the camp, his assistant Joshua the son of Nun, a young man, would not depart from the tent.
EXOD|33|12|Moses said to the LORD, "See, you say to me, 'Bring up this people,' but you have not let me know whom you will send with me. Yet you have said, 'I know you by name, and you have also found favor in my sight.'
EXOD|33|13|Now therefore, if I have found favor in your sight, please show me now your ways, that I may know you in order to find favor in your sight. Consider too that this nation is your people."
EXOD|33|14|And he said, "My presence will go with you, and I will give you rest."
EXOD|33|15|And he said to him, "If your presence will not go with me, do not bring us up from here.
EXOD|33|16|For how shall it be known that I have found favor in your sight, I and your people? Is it not in your going with us, so that we are distinct, I and your people, from every other people on the face of the earth?"
EXOD|33|17|And the LORD said to Moses, "This very thing that you have spoken I will do, for you have found favor in my sight, and I know you by name."
EXOD|33|18|Moses said, "Please show me your glory."
EXOD|33|19|And he said, "I will make all my goodness pass before you and will proclaim before you my name 'The LORD.' And I will be gracious to whom I will be gracious, and will show mercy on whom I will show mercy.
EXOD|33|20|But," he said, "you cannot see my face, for man shall not see me and live."
EXOD|33|21|And the LORD said, "Behold, there is a place by me where you shall stand on the rock,
EXOD|33|22|and while my glory passes by I will put you in a cleft of the rock, and I will cover you with my hand until I have passed by.
EXOD|33|23|Then I will take away my hand, and you shall see my back, but my face shall not be seen."
EXOD|34|1|The LORD said to Moses, "Cut for yourself two tablets of stone like the first, and I will write on the tablets the words that were on the first tablets, which you broke.
EXOD|34|2|Be ready by the morning, and come up in the morning to Mount Sinai, and present yourself there to me on the top of the mountain.
EXOD|34|3|No one shall come up with you, and let no one be seen throughout all the mountain. Let no flocks or herds graze opposite that mountain."
EXOD|34|4|So Moses cut two tablets of stone like the first. And he rose early in the morning and went up on Mount Sinai, as the LORD had commanded him, and took in his hand two tablets of stone.
EXOD|34|5|The LORD descended in the cloud and stood with him there, and proclaimed the name of the LORD.
EXOD|34|6|The LORD passed before him and proclaimed, "The LORD, the LORD, a God merciful and gracious, slow to anger, and abounding in steadfast love and faithfulness,
EXOD|34|7|keeping steadfast love for thousands, forgiving iniquity and transgression and sin, but who will by no means clear the guilty, visiting the iniquity of the fathers on the children and the children's children, to the third and the fourth generation."
EXOD|34|8|And Moses quickly bowed his head toward the earth and worshiped.
EXOD|34|9|And he said, "If now I have found favor in your sight, O Lord, please let the Lord go in the midst of us, for it is a stiff-necked people, and pardon our iniquity and our sin, and take us for your inheritance."
EXOD|34|10|And he said, "Behold, I am making a covenant. Before all your people I will do marvels, such as have not been created in all the earth or in any nation. And all the people among whom you are shall see the work of the LORD, for it is an awesome thing that I will do with you.
EXOD|34|11|"Observe what I command you this day. Behold, I will drive out before you the Amorites, the Canaanites, the Hittites, the Perizzites, the Hivites, and the Jebusites.
EXOD|34|12|Take care, lest you make a covenant with the inhabitants of the land to which you go, lest it become a snare in your midst.
EXOD|34|13|You shall tear down their altars and break their pillars and cut down their Asherim
EXOD|34|14|(for you shall worship no other god, for the LORD, whose name is Jealous, is a jealous God),
EXOD|34|15|lest you make a covenant with the inhabitants of the land, and when they whore after their gods and sacrifice to their gods and you are invited, you eat of his sacrifice,
EXOD|34|16|and you take of their daughters for your sons, and their daughters whore after their gods and make your sons whore after their gods.
EXOD|34|17|"You shall not make for yourself any gods of cast metal.
EXOD|34|18|"You shall keep the Feast of Unleavened Bread. Seven days you shall eat unleavened bread, as I commanded you, at the time appointed in the month Abib, for in the month Abib you came out from Egypt.
EXOD|34|19|All that open the womb are mine, all your male livestock, the firstborn of cow and sheep.
EXOD|34|20|The firstborn of a donkey you shall redeem with a lamb, or if you will not redeem it you shall break its neck. All the firstborn of your sons you shall redeem. And none shall appear before me empty-handed.
EXOD|34|21|"Six days you shall work, but on the seventh day you shall rest. In plowing time and in harvest you shall rest.
EXOD|34|22|You shall observe the Feast of Weeks, the firstfruits of wheat harvest, and the Feast of Ingathering at the year's end.
EXOD|34|23|Three times in the year shall all your males appear before the LORD God, the God of Israel.
EXOD|34|24|For I will cast out nations before you and enlarge your borders; no one shall covet your land, when you go up to appear before the LORD your God three times in the year.
EXOD|34|25|"You shall not offer the blood of my sacrifice with anything leavened, or let the sacrifice of the Feast of the Passover remain until the morning.
EXOD|34|26|The best of the firstfruits of your ground you shall bring to the house of the LORD your God. You shall not boil a young goat in its mother's milk."
EXOD|34|27|And the LORD said to Moses, "Write these words, for in accordance with these words I have made a covenant with you and with Israel."
EXOD|34|28|So he was there with the LORD forty days and forty nights. He neither ate bread nor drank water. And he wrote on the tablets the words of the covenant, the ten commandments.
EXOD|34|29|When Moses came down from Mount Sinai, with the two tablets of the testimony in his hand as he came down from the mountain, Moses did not know that the skin of his face shone because he had been talking with God.
EXOD|34|30|Aaron and all the people of Israel saw Moses, and behold, the skin of his face shone, and they were afraid to come near him.
EXOD|34|31|But Moses called to them, and Aaron and all the leaders of the congregation returned to him, and Moses talked with them.
EXOD|34|32|Afterward all the people of Israel came near, and he commanded them all that the LORD had spoken with him in Mount Sinai.
EXOD|34|33|And when Moses had finished speaking with them, he put a veil over his face.
EXOD|34|34|Whenever Moses went in before the LORD to speak with him, he would remove the veil, until he came out. And when he came out and told the people of Israel what he was commanded,
EXOD|34|35|the people of Israel would see the face of Moses, that the skin of Moses' face was shining. And Moses would put the veil over his face again, until he went in to speak with him.
EXOD|35|1|Moses assembled all the congregation of the people of Israel and said to them, "These are the things that the LORD has commanded you to do.
EXOD|35|2|Six days work shall be done, but on the seventh day you shall have a Sabbath of solemn rest, holy to the LORD. Whoever does any work on it shall be put to death.
EXOD|35|3|You shall kindle no fire in all your dwelling places on the Sabbath day."
EXOD|35|4|Moses said to all the congregation of the people of Israel, "This is the thing that the LORD has commanded.
EXOD|35|5|Take from among you a contribution to the LORD. Whoever is of a generous heart, let him bring the LORD's contribution: gold, silver, and bronze;
EXOD|35|6|blue and purple and scarlet yarns and fine twined linen; goats' hair,
EXOD|35|7|tanned rams' skins, and goatskins; acacia wood,
EXOD|35|8|oil for the light, spices for the anointing oil and for the fragrant incense,
EXOD|35|9|and onyx stones and stones for setting, for the ephod and for the breastpiece.
EXOD|35|10|"Let every skillful craftsman among you come and make all that the LORD has commanded:
EXOD|35|11|the tabernacle, its tent and its covering, its hooks and its frames, its bars, its pillars, and its bases;
EXOD|35|12|the ark with its poles, the mercy seat, and the veil of the screen;
EXOD|35|13|the table with its poles and all its utensils, and the bread of the Presence;
EXOD|35|14|the lampstand also for the light, with its utensils and its lamps, and the oil for the light;
EXOD|35|15|and the altar of incense, with its poles, and the anointing oil and the fragrant incense, and the screen for the door, at the door of the tabernacle;
EXOD|35|16|the altar of burnt offering, with its grating of bronze, its poles, and all its utensils, the basin and its stand;
EXOD|35|17|the hangings of the court, its pillars and its bases, and the screen for the gate of the court;
EXOD|35|18|the pegs of the tabernacle and the pegs of the court, and their cords;
EXOD|35|19|the finely worked garments for ministering in the Holy Place, the holy garments for Aaron the priest, and the garments of his sons, for their service as priests."
EXOD|35|20|Then all the congregation of the people of Israel departed from the presence of Moses.
EXOD|35|21|And they came, everyone whose heart stirred him, and everyone whose spirit moved him, and brought the LORD's contribution to be used for the tent of meeting, and for all its service, and for the holy garments.
EXOD|35|22|So they came, both men and women. All who were of a willing heart brought brooches and earrings and signet rings and armlets, all sorts of gold objects, every man dedicating an offering of gold to the LORD.
EXOD|35|23|And every one who possessed blue or purple or scarlet yarns or fine linen or goats' hair or tanned rams' skins or goatskins brought them.
EXOD|35|24|Everyone who could make a contribution of silver or bronze brought it as the LORD's contribution. And every one who possessed acacia wood of any use in the work brought it.
EXOD|35|25|And every skillful woman spun with her hands, and they all brought what they had spun in blue and purple and scarlet yarns and fine twined linen.
EXOD|35|26|All the women whose hearts stirred them to use their skill spun the goats' hair.
EXOD|35|27|And the leaders brought onyx stones and stones to be set, for the ephod and for the breastpiece,
EXOD|35|28|and spices and oil for the light, and for the anointing oil, and for the fragrant incense.
EXOD|35|29|All the men and women, the people of Israel, whose heart moved them to bring anything for the work that the LORD had commanded by Moses to be done brought it as a freewill offering to the LORD.
EXOD|35|30|Then Moses said to the people of Israel, "See, the LORD has called by name Bezalel the son of Uri, son of Hur, of the tribe of Judah;
EXOD|35|31|and he has filled him with the Spirit of God, with skill, with intelligence, with knowledge, and with all craftsmanship,
EXOD|35|32|to devise artistic designs, to work in gold and silver and bronze,
EXOD|35|33|in cutting stones for setting, and in carving wood, for work in every skilled craft.
EXOD|35|34|And he has inspired him to teach, both him and Oholiab the son of Ahisamach of the tribe of Dan.
EXOD|35|35|He has filled them with skill to do every sort of work done by an engraver or by a designer or by an embroiderer in blue and purple and scarlet yarns and fine twined linen, or by a weaver- by any sort of workman or skilled designer.
EXOD|36|1|"Bezalel and Oholiab and every craftsman in whom the LORD has put skill and intelligence to know how to do any work in the construction of the sanctuary shall work in accordance with all that the LORD has commanded."
EXOD|36|2|And Moses called Bezalel and Oholiab and every craftsman in whose mind the LORD had put skill, everyone whose heart stirred him up to come to do the work.
EXOD|36|3|And they received from Moses all the contribution that the people of Israel had brought for doing the work on the sanctuary. They still kept bringing him freewill offerings every morning,
EXOD|36|4|so that all the craftsmen who were doing every sort of task on the sanctuary came, each from the task that he was doing,
EXOD|36|5|and said to Moses, "The people bring much more than enough for doing the work that the LORD has commanded us to do."
EXOD|36|6|So Moses gave command, and word was proclaimed throughout the camp, "Let no man or woman do anything more for the contribution for the sanctuary." So the people were restrained from bringing,
EXOD|36|7|for the material they had was sufficient to do all the work, and more.
EXOD|36|8|And all the craftsmen among the workmen made the tabernacle with ten curtains. They were made of fine twined linen and blue and purple and scarlet yarns, with cherubim skillfully worked.
EXOD|36|9|The length of each curtain was twenty-eight cubits, and the breadth of each curtain four cubits. All the curtains were the same size.
EXOD|36|10|He coupled five curtains to one another, and the other five curtains he coupled to one another.
EXOD|36|11|He made loops of blue on the edge of the outermost curtain of the first set. Likewise he made them on the edge of the outermost curtain of the second set.
EXOD|36|12|He made fifty loops on the one curtain, and he made fifty loops on the edge of the curtain that was in the second set. The loops were opposite one another.
EXOD|36|13|And he made fifty clasps of gold, and coupled the curtains one to the other with clasps. So the tabernacle was a single whole.
EXOD|36|14|He also made curtains of goats' hair for a tent over the tabernacle. He made eleven curtains.
EXOD|36|15|The length of each curtain was thirty cubits, and the breadth of each curtain four cubits. The eleven curtains were the same size.
EXOD|36|16|He coupled five curtains by themselves, and six curtains by themselves.
EXOD|36|17|And he made fifty loops on the edge of the outermost curtain of the one set, and fifty loops on the edge of the other connecting curtain.
EXOD|36|18|And he made fifty clasps of bronze to couple the tent together that it might be a single whole.
EXOD|36|19|And he made for the tent a covering of tanned rams' skins and goatskins.
EXOD|36|20|Then he made the upright frames for the tabernacle of acacia wood.
EXOD|36|21|Ten cubits was the length of a frame, and a cubit and a half the breadth of each frame.
EXOD|36|22|Each frame had two tenons for fitting together. He did this for all the frames of the tabernacle.
EXOD|36|23|The frames for the tabernacle he made thus: twenty frames for the south side.
EXOD|36|24|And he made forty bases of silver under the twenty frames, two bases under one frame for its two tenons, and two bases under the next frame for its two tenons.
EXOD|36|25|For the second side of the tabernacle, on the north side, he made twenty frames
EXOD|36|26|and their forty bases of silver, two bases under one frame and two bases under the next frame.
EXOD|36|27|For the rear of the tabernacle westward he made six frames.
EXOD|36|28|He made two frames for corners of the tabernacle in the rear.
EXOD|36|29|And they were separate beneath but joined at the top, at the first ring. He made two of them this way for the two corners.
EXOD|36|30|There were eight frames with their bases of silver: sixteen bases, under every frame two bases.
EXOD|36|31|He made bars of acacia wood, five for the frames of the one side of the tabernacle,
EXOD|36|32|and five bars for the frames of the other side of the tabernacle, and five bars for the frames of the tabernacle at the rear westward.
EXOD|36|33|And he made the middle bar to run from end to end halfway up the frames.
EXOD|36|34|And he overlaid the frames with gold, and made their rings of gold for holders for the bars, and overlaid the bars with gold.
EXOD|36|35|He made the veil of blue and purple and scarlet yarns and fine twined linen; with cherubim skillfully worked into it he made it.
EXOD|36|36|And for it he made four pillars of acacia and overlaid them with gold. Their hooks were of gold, and he cast for them four bases of silver.
EXOD|36|37|He also made a screen for the entrance of the tent, of blue and purple and scarlet yarns and fine twined linen, embroidered with needlework,
EXOD|36|38|and its five pillars with their hooks. He overlaid their capitals, and their fillets were of gold, but their five bases were of bronze.
EXOD|37|1|Bezalel made the ark of acacia wood. Two cubits and a half was its length, a cubit and a half its breadth, and a cubit and a half its height.
EXOD|37|2|And he overlaid it with pure gold inside and outside, and made a molding of gold around it.
EXOD|37|3|And he cast for it four rings of gold for its four feet, two rings on its one side and two rings on its other side.
EXOD|37|4|And he made poles of acacia wood and overlaid them with gold
EXOD|37|5|and put the poles into the rings on the sides of the ark to carry the ark.
EXOD|37|6|And he made a mercy seat of pure gold. Two cubits and a half was its length, and a cubit and a half its breadth.
EXOD|37|7|And he made two cherubim of gold. He made them of hammered work on the two ends of the mercy seat,
EXOD|37|8|one cherub on the one end, and one cherub on the other end. Of one piece with the mercy seat he made the cherubim on its two ends.
EXOD|37|9|The cherubim spread out their wings above, overshadowing the mercy seat with their wings, with their faces one to another; toward the mercy seat were the faces of the cherubim.
EXOD|37|10|He also made the table of acacia wood. Two cubits was its length, a cubit its breadth, and a cubit and a half its height.
EXOD|37|11|And he overlaid it with pure gold, and made a molding of gold around it.
EXOD|37|12|And he made a rim around it a handbreadth wide, and made a molding of gold around the rim.
EXOD|37|13|He cast for it four rings of gold and fastened the rings to the four corners at its four legs.
EXOD|37|14|Close to the frame were the rings, as holders for the poles to carry the table.
EXOD|37|15|He made the poles of acacia wood to carry the table, and overlaid them with gold.
EXOD|37|16|And he made the vessels of pure gold that were to be on the table, its plates and dishes for incense, and its bowls and flagons with which to pour drink offerings.
EXOD|37|17|He also made the lampstand of pure gold. He made the lampstand of hammered work. Its base, its stem, its cups, its calyxes, and its flowers were of one piece with it.
EXOD|37|18|And there were six branches going out of its sides, three branches of the lampstand out of one side of it and three branches of the lampstand out of the other side of it;
EXOD|37|19|three cups made like almond blossoms, each with calyx and flower, on one branch, and three cups made like almond blossoms, each with calyx and flower, on the other branch- so for the six branches going out of the lampstand.
EXOD|37|20|And on the lampstand itself were four cups made like almond blossoms, with their calyxes and flowers,
EXOD|37|21|and a calyx of one piece with it under each pair of the six branches going out of it.
EXOD|37|22|Their calyxes and their branches were of one piece with it. The whole of it was a single piece of hammered work of pure gold.
EXOD|37|23|And he made its seven lamps and its tongs and its trays of pure gold.
EXOD|37|24|He made it and all its utensils out of a talent of pure gold.
EXOD|37|25|He made the altar of incense of acacia wood. Its length was a cubit, and its breadth was a cubit. It was square, and two cubits was its height. Its horns were of one piece with it.
EXOD|37|26|He overlaid it with pure gold, its top and around its sides and its horns. And he made a molding of gold around it,
EXOD|37|27|and made two rings of gold on it under its molding, on two opposite sides of it, as holders for the poles with which to carry it.
EXOD|37|28|And he made the poles of acacia wood and overlaid them with gold.
EXOD|37|29|He made the holy anointing oil also, and the pure fragrant incense, blended as by the perfumer.
EXOD|38|1|He made the altar of burnt offering of acacia wood. Five cubits was its length, and five cubits its breadth. It was square, and three cubits was its height.
EXOD|38|2|He made horns for it on its four corners. Its horns were of one piece with it, and he overlaid it with bronze.
EXOD|38|3|And he made all the utensils of the altar, the pots, the shovels, the basins, the forks, and the fire pans. He made all its utensils of bronze.
EXOD|38|4|And he made for the altar a grating, a network of bronze, under its ledge, extending halfway down.
EXOD|38|5|He cast four rings on the four corners of the bronze grating as holders for the poles.
EXOD|38|6|He made the poles of acacia wood and overlaid them with bronze.
EXOD|38|7|And he put the poles through the rings on the sides of the altar to carry it with them. He made it hollow, with boards.
EXOD|38|8|He made the basin of bronze and its stand of bronze, from the mirrors of the ministering women who ministered in the entrance of the tent of meeting.
EXOD|38|9|And he made the court. For the south side the hangings of the court were of fine twined linen, a hundred cubits;
EXOD|38|10|their twenty pillars and their twenty bases were of bronze, but the hooks of the pillars and their fillets were of silver.
EXOD|38|11|And for the north side there were hangings of a hundred cubits, their twenty pillars, their twenty bases were of bronze, but the hooks of the pillars and their fillets were of silver.
EXOD|38|12|And for the west side were hangings of fifty cubits, their ten pillars, and their ten bases; the hooks of the pillars and their fillets were of silver.
EXOD|38|13|And for the front to the east, fifty cubits.
EXOD|38|14|The hangings for one side of the gate were fifteen cubits, with their three pillars and three bases.
EXOD|38|15|And so for the other side. On both sides of the gate of the court were hangings of fifteen cubits, with their three pillars and their three bases.
EXOD|38|16|All the hangings around the court were of fine twined linen.
EXOD|38|17|And the bases for the pillars were of bronze, but the hooks of the pillars and their fillets were of silver. The overlaying of their capitals was also of silver, and all the pillars of the court were filleted with silver.
EXOD|38|18|And the screen for the gate of the court was embroidered with needlework in blue and purple and scarlet yarns and fine twined linen. It was twenty cubits long and five cubits high in its breadth, corresponding to the hangings of the court.
EXOD|38|19|And their pillars were four in number. Their four bases were of bronze, their hooks of silver, and the overlaying of their capitals and their fillets of silver.
EXOD|38|20|And all the pegs for the tabernacle and for the court all around were of bronze.
EXOD|38|21|These are the records of the tabernacle, the tabernacle of the testimony, as they were recorded at the commandment of Moses, the responsibility of the Levites under the direction of Ithamar the son of Aaron the priest.
EXOD|38|22|Bezalel the son of Uri, son of Hur, of the tribe of Judah, made all that the LORD commanded Moses;
EXOD|38|23|and with him was Oholiab the son of Ahisamach, of the tribe of Dan, an engraver and designer and embroiderer in blue and purple and scarlet yarns and fine twined linen.
EXOD|38|24|All the gold that was used for the work, in all the construction of the sanctuary, the gold from the offering, was twenty-nine talents and 730 shekels, by the shekel of the sanctuary.
EXOD|38|25|The silver from those of the congregation who were recorded was a hundred talents and 1,775 shekels, by the shekel of the sanctuary:
EXOD|38|26|a beka a head (that is, half a shekel, by the shekel of the sanctuary), for everyone who was listed in the records, from twenty years old and upward, for 603,550 men.
EXOD|38|27|The hundred talents of silver were for casting the bases of the sanctuary and the bases of the veil; a hundred bases for the hundred talents, a talent a base.
EXOD|38|28|And of the 1,775 shekels he made hooks for the pillars and overlaid their capitals and made fillets for them.
EXOD|38|29|The bronze that was offered was seventy talents and 2,400 shekels;
EXOD|38|30|with it he made the bases for the entrance of the tent of meeting, the bronze altar and the bronze grating for it and all the utensils of the altar,
EXOD|38|31|the bases around the court, and the bases of the gate of the court, all the pegs of the tabernacle, and all the pegs around the court.
EXOD|39|1|From the blue and purple and scarlet yarns they made finely woven garments, for ministering in the Holy Place. They made the holy garments for Aaron, as the LORD had commanded Moses.
EXOD|39|2|He made the ephod of gold, blue and purple and scarlet yarns, and fine twined linen.
EXOD|39|3|And they hammered out gold leaf, and he cut it into threads to work into the blue and purple and the scarlet yarns, and into the fine twined linen, in skilled design.
EXOD|39|4|They made for the ephod attaching shoulder pieces, joined to it at its two edges.
EXOD|39|5|And the skillfully woven band on it was of one piece with it and made like it, of gold, blue and purple and scarlet yarns, and fine twined linen, as the LORD had commanded Moses.
EXOD|39|6|They made the onyx stones, enclosed in settings of gold filigree, and engraved like the engravings of a signet, according to the names of the sons of Israel.
EXOD|39|7|And he set them on the shoulder pieces of the ephod to be stones of remembrance for the sons of Israel, as the LORD had commanded Moses.
EXOD|39|8|He made the breastpiece, in skilled work, in the style of the ephod, of gold, blue and purple and scarlet yarns, and fine twined linen.
EXOD|39|9|It was square. They made the breastpiece doubled, a span its length and a span its breadth when doubled.
EXOD|39|10|And they set in it four rows of stones. A row of sardius, topaz, and carbuncle was the first row;
EXOD|39|11|and the second row, an emerald, a sapphire, and a diamond;
EXOD|39|12|and the third row, a jacinth, an agate, and an amethyst;
EXOD|39|13|and the fourth row, a beryl, an onyx, and a jasper. They were enclosed in settings of gold filigree.
EXOD|39|14|There were twelve stones with their names according to the names of the sons of Israel. They were like signets, each engraved with its name, for the twelve tribes.
EXOD|39|15|And they made on the breastpiece twisted chains like cords, of pure gold.
EXOD|39|16|And they made two settings of gold filigree and two gold rings, and put the two rings on the two edges of the breastpiece.
EXOD|39|17|And they put the two cords of gold in the two rings at the edges of the breastpiece.
EXOD|39|18|They attached the two ends of the two cords to the two settings of filigree. Thus they attached it in front to the shoulder pieces of the ephod.
EXOD|39|19|Then they made two rings of gold, and put them at the two ends of the breastpiece, on its inside edge next to the ephod.
EXOD|39|20|And they made two rings of gold, and attached them in front to the lower part of the two shoulder pieces of the ephod, at its seam above the skillfully woven band of the ephod.
EXOD|39|21|And they bound the breastpiece by its rings to the rings of the ephod with a lace of blue, so that it should lie on the skillfully woven band of the ephod, and that the breastpiece should not come loose from the ephod, as the LORD had commanded Moses.
EXOD|39|22|He also made the robe of the ephod woven all of blue,
EXOD|39|23|and the opening of the robe in it was like the opening in a garment, with a binding around the opening, so that it might not tear.
EXOD|39|24|On the hem of the robe they made pomegranates of blue and purple and scarlet yarns and fine twined linen.
EXOD|39|25|They also made bells of pure gold, and put the bells between the pomegranates all around the hem of the robe, between the pomegranates-
EXOD|39|26|a bell and a pomegranate, a bell and a pomegranate around the hem of the robe for ministering, as the LORD had commanded Moses.
EXOD|39|27|They also made the coats, woven of fine linen, for Aaron and his sons,
EXOD|39|28|and the turban of fine linen, and the caps of fine linen, and the linen undergarments of fine twined linen,
EXOD|39|29|and the sash of fine twined linen and of blue and purple and scarlet yarns, embroidered with needlework, as the LORD had commanded Moses.
EXOD|39|30|They made the plate of the holy crown of pure gold, and wrote on it an inscription, like the engraving of a signet, "Holy to the LORD."
EXOD|39|31|And they tied to it a cord of blue to fasten it on the turban above, as the LORD had commanded Moses.
EXOD|39|32|Thus all the work of the tabernacle of the tent of meeting was finished, and the people of Israel did according to all that the LORD had commanded Moses; so they did.
EXOD|39|33|Then they brought the tabernacle to Moses, the tent and all its utensils, its hooks, its frames, its bars, its pillars, and its bases;
EXOD|39|34|the covering of tanned rams' skins and goatskins, and the veil of the screen;
EXOD|39|35|the ark of the testimony with its poles and the mercy seat;
EXOD|39|36|the table with all its utensils, and the bread of the Presence;
EXOD|39|37|the lampstand of pure gold and its lamps with the lamps set and all its utensils, and the oil for the light;
EXOD|39|38|the golden altar, the anointing oil and the fragrant incense, and the screen for the entrance of the tent;
EXOD|39|39|the bronze altar, and its grating of bronze, its poles, and all its utensils; the basin and its stand;
EXOD|39|40|the hangings of the court, its pillars, and its bases, and the screen for the gate of the court, its cords, and its pegs; and all the utensils for the service of the tabernacle, for the tent of meeting;
EXOD|39|41|the finely worked garments for ministering in the Holy Place, the holy garments for Aaron the priest, and the garments of his sons for their service as priests.
EXOD|39|42|According to all that the LORD had commanded Moses, so the people of Israel had done all the work.
EXOD|39|43|And Moses saw all the work, and behold, they had done it; as the LORD had commanded, so had they done it. Then Moses blessed them.
EXOD|40|1|The LORD spoke to Moses, saying,
EXOD|40|2|"On the first day of the first month you shall erect the tabernacle of the tent of meeting.
EXOD|40|3|And you shall put in it the ark of the testimony, and you shall screen the ark with the veil.
EXOD|40|4|And you shall bring in the table and arrange it, and you shall bring in the lampstand and set up its lamps.
EXOD|40|5|And you shall put the golden altar for incense before the ark of the testimony, and set up the screen for the door of the tabernacle.
EXOD|40|6|You shall set the altar of burnt offering before the door of the tabernacle of the tent of meeting,
EXOD|40|7|and place the basin between the tent of meeting and the altar, and put water in it.
EXOD|40|8|And you shall set up the court all around, and hang up the screen for the gate of the court.
EXOD|40|9|"Then you shall take the anointing oil and anoint the tabernacle and all that is in it, and consecrate it and all its furniture, so that it may become holy.
EXOD|40|10|You shall also anoint the altar of burnt offering and all its utensils, and consecrate the altar, so that the altar may become most holy.
EXOD|40|11|You shall also anoint the basin and its stand, and consecrate it.
EXOD|40|12|Then you shall bring Aaron and his sons to the entrance of the tent of meeting and shall wash them with water
EXOD|40|13|and put on Aaron the holy garments. And you shall anoint him and consecrate him, that he may serve me as priest.
EXOD|40|14|You shall bring his sons also and put coats on them,
EXOD|40|15|and anoint them, as you anointed their father, that they may serve me as priests. And their anointing shall admit them to a perpetual priesthood throughout their generations."
EXOD|40|16|This Moses did; according to all that the LORD commanded him, so he did.
EXOD|40|17|In the first month in the second year, on the first day of the month, the tabernacle was erected.
EXOD|40|18|Moses erected the tabernacle. He laid its bases, and set up its frames, and put in its poles, and raised up its pillars.
EXOD|40|19|And he spread the tent over the tabernacle and put the covering of the tent over it, as the LORD had commanded Moses.
EXOD|40|20|He took the testimony and put it into the ark, and put the poles on the ark and set the mercy seat above on the ark.
EXOD|40|21|And he brought the ark into the tabernacle and set up the veil of the screen, and screened the ark of the testimony, as the LORD had commanded Moses.
EXOD|40|22|He put the table in the tent of meeting, on the north side of the tabernacle, outside the veil,
EXOD|40|23|and arranged the bread on it before the LORD, as the LORD had commanded Moses.
EXOD|40|24|He put the lampstand in the tent of meeting, opposite the table on the south side of the tabernacle,
EXOD|40|25|and set up the lamps before the LORD, as the LORD had commanded Moses.
EXOD|40|26|He put the golden altar in the tent of meeting before the veil,
EXOD|40|27|and burned fragrant incense on it, as the LORD had commanded Moses.
EXOD|40|28|He put in place the screen for the door of the tabernacle.
EXOD|40|29|And he set the altar of burnt offering at the entrance of the tabernacle of the tent of meeting, and offered on it the burnt offering and the grain offering, as the LORD had commanded Moses.
EXOD|40|30|He set the basin between the tent of meeting and the altar, and put water in it for washing,
EXOD|40|31|with which Moses and Aaron and his sons washed their hands and their feet.
EXOD|40|32|When they went into the tent of meeting, and when they approached the altar, they washed, as the LORD commanded Moses.
EXOD|40|33|And he erected the court around the tabernacle and the altar, and set up the screen of the gate of the court. So Moses finished the work.
EXOD|40|34|Then the cloud covered the tent of meeting, and the glory of the LORD filled the tabernacle.
EXOD|40|35|And Moses was not able to enter the tent of meeting because the cloud settled on it, and the glory of the LORD filled the tabernacle.
EXOD|40|36|Throughout all their journeys, whenever the cloud was taken up from over the tabernacle, the people of Israel would set out.
EXOD|40|37|But if the cloud was not taken up, then they did not set out till the day that it was taken up.
EXOD|40|38|For the cloud of the LORD was on the tabernacle by day, and fire was in it by night, in the sight of all the house of Israel throughout all their journeys.
