1CHR|1|1|Adam Seth Enos
1CHR|1|2|Cainan Malelehel Iared
1CHR|1|3|Enoch Matusale Lamech
1CHR|1|4|Noe Sem Ham et Iafeth
1CHR|1|5|filii Iafeth Gomer Magog Madai et Iavan Thubal Mosoch Thiras
1CHR|1|6|porro filii Gomer Aschenez et Rifath et Thogorma
1CHR|1|7|filii autem Iavan Elisa et Tharsis Cetthim et Dodanim
1CHR|1|8|filii Ham Chus et Mesraim Phut et Chanaan
1CHR|1|9|filii autem Chus Saba et Evila Sabatha et Rechma et Sabathaca porro filii Rechma Saba et Dadan
1CHR|1|10|Chus autem genuit Nemrod iste coepit esse potens in terra
1CHR|1|11|Mesraim vero genuit Ludim et Anamim et Laabim et Nepthuim
1CHR|1|12|Phethrosim quoque et Chasluim de quibus egressi sunt Philisthim et Capthurim
1CHR|1|13|Chanaan vero genuit Sidonem primogenitum et Heth
1CHR|1|14|Iebuseum quoque et Amorreum et Gergeseum
1CHR|1|15|Evheumque et Aruceum et Asineum
1CHR|1|16|Aradium quoque et Samareum et Ematheum
1CHR|1|17|filii Sem Aelam et Assur et Arfaxad et Lud et Aram et Us et Hul et Gothor et Mosoch
1CHR|1|18|Arfaxad autem genuit Sala qui et ipse genuit Heber
1CHR|1|19|porro Heber nati sunt duo filii nomen uni Phaleg quia in diebus eius divisa est terra et nomen fratris eius Iectan
1CHR|1|20|Iectan autem genuit Helmodad et Saleph et Asermoth et Iare
1CHR|1|21|Aduram quoque et Uzal et Decla
1CHR|1|22|Ebal etiam et Abimahel et Saba necnon
1CHR|1|23|et Ophir et Evila et Iobab omnes isti filii Iectan
1CHR|1|24|Sem Arfaxad Sale
1CHR|1|25|Heber Phaleg Raau
1CHR|1|26|Serug Nahor Thare
1CHR|1|27|Abram iste est Abraham
1CHR|1|28|filii autem Abraham Isaac et Ismahel
1CHR|1|29|et hae generationes eorum primogenitus Ismahelis Nabaioth et Cedar et Adbeel et Mabsam
1CHR|1|30|Masma et Duma Massa Adad et Thema
1CHR|1|31|Iathur Naphis Cedma hii sunt filii Ismahelis
1CHR|1|32|filii autem Cetthurae concubinae Abraham quos genuit Zamram Iecsan Madan Madian Iesboc Sue porro filii Iecsan Saba et Dadan
1CHR|1|33|filii autem Madian Epha et Apher et Enoch et Abida et Eldaa omnes hii filii Cetthurae
1CHR|1|34|generavit autem Abraham Isaac cuius fuerunt filii Esau et Israhel
1CHR|1|35|filii Esau Eliphaz Rauhel Iaus Ialam Core
1CHR|1|36|filii Eliphaz Theman Omer Sepphu Gethem Cenez Thamna Amalech
1CHR|1|37|filii Rauhel Naath Zara Samma Maza
1CHR|1|38|filii Seir Lothan Sobal Sebeon Ana Dison Eser Disan
1CHR|1|39|filii Lothan Horri Humam soror autem Lothan fuit Thamna
1CHR|1|40|filii Sobal Alian et Manaath et Ebal et Sepphi et Onam filii Sebeon Aia et Ana filii Ana Dison
1CHR|1|41|filii Dison Amaran et Eseban et Iethran et Charan
1CHR|1|42|filii Eser Balaan et Zaban et Iacan filii Dison Us et Aran
1CHR|1|43|isti sunt reges qui imperaverunt in terra Edom antequam esset rex super filios Israhel Bale filius Beor et nomen civitatis eius Denaba
1CHR|1|44|mortuus est autem Bale et regnavit pro eo Iobab filius Zare de Bosra
1CHR|1|45|cumque et Iobab fuisset mortuus regnavit pro eo Husam de terra Themanorum
1CHR|1|46|obiit quoque et Husam et regnavit pro eo Adad filius Badad qui percussit Madian in terra Moab et nomen civitatis eius Avith
1CHR|1|47|cumque et Adad fuisset mortuus regnavit pro eo Semla de Masreca
1CHR|1|48|sed et Semla mortuus est et regnavit pro eo Saul de Rooboth quae iuxta amnem sita est
1CHR|1|49|mortuo quoque Saul regnavit pro eo Baalanan filius Achobor
1CHR|1|50|sed et hic mortuus est et regnavit pro eo Adad cuius urbis fuit nomen Phou et appellata est uxor eius Mehetabel filia Matred filiae Mezaab
1CHR|1|51|Adad autem mortuo duces pro regibus in Edom esse coeperunt dux Thamna dux Alva dux Ietheth
1CHR|1|52|dux Oolibama dux Hela dux Phinon
1CHR|1|53|dux Cenez dux Theman dux Mabsar
1CHR|1|54|dux Magdihel dux Iram hii duces Edom
1CHR|2|1|filii autem Israhel Ruben Symeon Levi Iuda Isachar et Zabulon
1CHR|2|2|Dan Ioseph Beniamin Nepthali Gad Aser
1CHR|2|3|filii Iuda Her Aunan Sela tres nati sunt ei de filia Sue Chananitidis fuit autem Her primogenitus Iuda malus coram Domino et occidit eum
1CHR|2|4|Thamar autem nurus eius peperit ei Phares et Zara omnes ergo filii Iuda quinque
1CHR|2|5|filii autem Phares Esrom et Hamul
1CHR|2|6|filii quoque Zarae Zamri et Ethan et Eman Chalchal quoque et Darda simul quinque
1CHR|2|7|filii Carmi Achar qui turbavit Israhel et peccavit in furto anathematis
1CHR|2|8|filii Ethan Azarias
1CHR|2|9|filii autem Esrom qui nati sunt ei Ieremahel et Ram et Chalubi
1CHR|2|10|porro Ram genuit Aminadab Aminadab autem genuit Naasson principem filiorum Iuda
1CHR|2|11|Naasson quoque genuit Salma de quo ortus est Boez
1CHR|2|12|Boez vero genuit Obed qui et ipse genuit Isai
1CHR|2|13|Isai autem genuit primogenitum Heliab secundum Abinadab tertium Samaa
1CHR|2|14|quartum Nathanahel quintum Raddai
1CHR|2|15|sextum Asom septimum David
1CHR|2|16|quorum sorores fuerunt Sarvia et Abigail filii Sarviae Abisai Ioab et Asahel tres
1CHR|2|17|Abigail autem genuit Amasa cuius pater fuit Iether Ismahelites
1CHR|2|18|Chaleb vero filius Esrom accepit uxorem nomine Azuba de qua genuit Ierioth fueruntque filii eius Iesar et Sobab et Ardon
1CHR|2|19|cumque mortua fuisset Azuba accepit uxorem Chaleb Ephrath quae peperit ei Ur
1CHR|2|20|porro Ur genuit Uri et Uri genuit Beselehel
1CHR|2|21|post haec ingressus est Esrom ad filiam Machir patris Galaad et accepit eam cum esset annorum sexaginta quae peperit ei Segub
1CHR|2|22|sed et Segub genuit Iair et possedit viginti tres civitates in terra Galaad
1CHR|2|23|cepitque Gessur et Aram oppida Iair et Canath et viculos eius sexaginta civitatum omnes isti filii Machir patris Galaad
1CHR|2|24|cum autem mortuus esset Esrom ingressus est Chaleb ad Ephrata habuit quoque Esrom uxorem Abia quae peperit ei Assur patrem Thecue
1CHR|2|25|nati sunt autem filii Hieramehel primogeniti Esrom Ram primogenitus eius et Buna et Aran et Asom et Ahia
1CHR|2|26|duxit quoque uxorem alteram Hieramehel nomine Atara quae fuit mater Onam
1CHR|2|27|sed et filii Ram primogeniti Hieramehel fuerunt Moos et Iamin et Achar
1CHR|2|28|Onam autem habuit filios Semmei et Iada filii autem Semmei Nadab et Abisur
1CHR|2|29|nomen vero uxoris Abisur Abiail quae peperit Ahobban et Molid
1CHR|2|30|filii autem Nadab fuerunt Saled et Apphaim mortuus est autem Saled absque liberis
1CHR|2|31|filius vero Apphaim Iesi qui Iesi genuit Sesan porro Sesan genuit Oholi
1CHR|2|32|filii autem Iada fratris Semmei Iether et Ionathan sed et Iether mortuus est absque liberis
1CHR|2|33|porro Ionathan genuit Phaleth et Ziza isti fuerunt filii Hieramehel
1CHR|2|34|Sesan autem non habuit filios sed filias et servum aegyptium nomine Ieraa
1CHR|2|35|deditque ei filiam suam uxorem quae peperit ei Eththei
1CHR|2|36|Eththei autem genuit Nathan et Nathan genuit Zabad
1CHR|2|37|Zabad quoque genuit Ophlal et Ophlal genuit Obed
1CHR|2|38|Obed genuit Ieu Ieu genuit Azariam
1CHR|2|39|Azarias genuit Helles Helles genuit Elasa
1CHR|2|40|Elasa genuit Sisamoi Sisamoi genuit Sellum
1CHR|2|41|Sellum genuit Icamian Icamian genuit Elisama
1CHR|2|42|filii autem Chaleb fratris Hieramehel Mosa primogenitus eius ipse est pater Ziph et filii Maresa patris Hebron
1CHR|2|43|porro filii Hebron Core et Thapphu et Recem et Samma
1CHR|2|44|Samma autem genuit Raam patrem Iercaam et Recem genuit Semmei
1CHR|2|45|filius Semmei Maon et Maon pater Bethsur
1CHR|2|46|Epha autem concubina Chaleb peperit Arran et Musa et Gezez porro Arran genuit Gezez
1CHR|2|47|filii Iadai Regom et Iotham et Gesum et Phaleth et Epha et Saaph
1CHR|2|48|concubina Chaleb Maacha peperit Saber et Tharana
1CHR|2|49|genuit autem Saaph pater Madmena Sue patrem Machbena et patrem Gabaa filia vero Chaleb fuit Achsa
1CHR|2|50|hii erant filii Chaleb filii Ur primogeniti Ephrata Sobal pater Cariathiarim
1CHR|2|51|Salma pater Bethleem Ariph pater Bethgader
1CHR|2|52|fuerunt autem filii Sobal patris Cariathiarim qui videbat dimidium requietionum
1CHR|2|53|et de cognatione Cariathiarim Iethrei et Apphutei et Semathei et Maserei ex his egressi sunt Saraitae et Esthaolitae
1CHR|2|54|filii Salma Bethleem et Netophathi coronae domus Ioab et dimidium requietionis Sarai
1CHR|2|55|cognationes quoque scribarum habitantium in Iabis canentes atque resonantes et in tabernaculis commorantes hii sunt Cinei qui venerunt de calore patris domus Rechab
1CHR|3|1|David vero hos habuit filios qui ei nati sunt in Hebron primogenitum Amnon ex Achinaam Iezrahelitide secundum Danihel de Abigail Carmelitide
1CHR|3|2|tertium Absalom filium Maacha filiae Tholmei regis Gessur quartum Adoniam filium Aggith
1CHR|3|3|quintum Saphatiam ex Abital sextum Iethraam de Egla uxore sua
1CHR|3|4|sex ergo nati sunt ei in Hebron ubi regnavit septem annis et sex mensibus triginta autem et tribus annis regnavit in Hierusalem
1CHR|3|5|porro in Hierusalem nati sunt ei filii Samaa et Sobab et Nathan et Salomon quattuor de Bethsabee filia Amihel
1CHR|3|6|Iebaar quoque et Elisama
1CHR|3|7|et Eliphalet et Noge et Napheg et Iaphie
1CHR|3|8|necnon Elisama et Heliade et Eliphalet novem
1CHR|3|9|omnes hii filii David absque filiis concubinarum habuerunt sororem Thamar
1CHR|3|10|filius autem Salomonis Roboam cuius Abia filius genuit Asa de hoc quoque natus est Iosaphat
1CHR|3|11|pater Ioram qui Ioram genuit Ohoziam ex quo ortus est Ioas
1CHR|3|12|et huius Amasias filius genuit Azariam porro Azariae filius Ioatham
1CHR|3|13|procreavit Achaz patrem Ezechiae de quo natus est Manasses
1CHR|3|14|sed et Manasses genuit Amon patrem Iosiae
1CHR|3|15|filii autem Iosiae fuerunt primogenitus Iohanan secundus Ioacim tertius Sedecias quartus Sellum
1CHR|3|16|de Ioacim natus est Iechonias et Sedecias
1CHR|3|17|filii Iechoniae fuerunt Asir Salathihel
1CHR|3|18|Melchiram Phadaia Sennaser et Iecemia Sama et Nadabia
1CHR|3|19|de Phadaia orti sunt Zorobabel et Semei Zorobabel genuit Mosollam Ananiam et Salomith sororem eorum
1CHR|3|20|Asabamque et Ohol et Barachiam et Asadiam Iosabesed quinque
1CHR|3|21|filius autem Ananiae Phaltias pater Ieseiae cuius filius Raphaia huius quoque filius Arnam de quo natus est Obdia cuius filius fuit Sechenia
1CHR|3|22|filius Secheniae Semeia cuius filii Attus et Iegal et Baria et Naaria et Saphat sex numero
1CHR|3|23|filius Naariae Helioenai et Ezechias et Ezricam tres
1CHR|3|24|filii Helioenai Oduia et Heliasub et Pheleia et Accub et Iohanan et Dalaia et Anani septem
1CHR|4|1|filii Iuda Phares Esrom et Carmi et Ur et Subal
1CHR|4|2|Reaia vero filius Subal genuit Ieth de quo nati sunt Ahimai et Laed hae cognationes Sarathi
1CHR|4|3|ista quoque stirps Hetam Iezrahel et Iesema et Iedebos nomenque sororis eorum Asalelphuni
1CHR|4|4|Phunihel autem pater Gedor et Ezer pater Osa isti sunt filii Ur primogeniti Ephrata patris Bethleem
1CHR|4|5|Asur vero patris Thecue erant duae uxores Halaa et Naara
1CHR|4|6|peperit autem ei Naara Oozam et Epher et Themani et Asthari isti sunt filii Naara
1CHR|4|7|porro filii Halaa Sereth Isaar et Ethnan
1CHR|4|8|Cos autem genuit Anob et Sobaba et cognationem Aral filii Arum
1CHR|4|9|fuit autem Iabes inclitus prae fratribus suis et mater eius vocavit nomen illius Iabes dicens quia peperi eum in dolore
1CHR|4|10|invocavit vero Iabes Deum Israhel dicens si benedicens benedixeris mihi et dilataveris terminos meos et fuerit manus tua mecum et feceris me a malitia non opprimi et praestitit Deus quae precatus est
1CHR|4|11|Chaleb autem frater Suaa genuit Machir qui fuit pater Esthon
1CHR|4|12|porro Esthon genuit Bethrapha et Phesse et Thena patrem urbis Naas hii sunt viri Recha
1CHR|4|13|filii autem Cenez Othonihel et Saraia porro filii Othonihel Athath
1CHR|4|14|et Maonathi genuit Ophra Saraias autem genuit Ioab patrem vallis Artificum ibi quippe artifices erant
1CHR|4|15|filii vero Chaleb filii Iephonne Hir et Hela et Nahem filiique Hela et Cenez
1CHR|4|16|filii quoque Iallelel Ziph et Zipha Thiria et Asrahel
1CHR|4|17|et filii Ezra Iether et Mered et Epher et Ialon genuitque Mariam et Sammai et Iesba patrem Esthamo
1CHR|4|18|uxor quoque eius Iudaia peperit Iared patrem Gedor et Heber patrem Soccho et Hicuthihel patrem Zano hii autem filii Beththiae filiae Pharaonis quam accepit Mered
1CHR|4|19|et filii uxoris Odaiae sororis Naham patris Ceila Garmi et Esthamo qui fuit de Machathi
1CHR|4|20|filii quoque Simon Amnon et Rena filius Anan et Thilon et filii Iesi Zoeth et Benzoeth
1CHR|4|21|filii Sela filii Iuda Her pater Lecha et Laada pater Maresa et cognationes Domus operantium byssum in domo Iuramenti
1CHR|4|22|et Qui stare fecit solem virique Mendacii et Securus et Incendens qui principes fuerunt in Moab et qui reversi sunt in Leem haec autem verba vetera
1CHR|4|23|hii sunt figuli habitantes in plantationibus et in praesepibus apud regem in operibus eius commoratique sunt ibi
1CHR|4|24|filii Symeon Namuhel et Iamin Iarib Zara Saul
1CHR|4|25|Sellum filius eius Mabsam filius eius Masma filius eius
1CHR|4|26|filii Masma Amuhel filius eius Zacchur filius eius Semei filius eius
1CHR|4|27|filii Semei sedecim et filiae sex fratres autem eius non habuerunt filios multos et universa cognatio non potuit adaequare summam filiorum Iuda
1CHR|4|28|habitaverunt autem in Bersabee et Molada et Asarsual
1CHR|4|29|et in Ballaa et in Asom et in Tholad
1CHR|4|30|et in Bathuhel et in Orma et in Siceleg
1CHR|4|31|et in Bethmarchaboth et in Asarsusim et in Bethberai et in Saarim hae civitates eorum usque ad regem David
1CHR|4|32|villae quoque eorum Etham et Aen et Remmon et Thochen et Asan civitates quinque
1CHR|4|33|et universi viculi eorum per circuitum civitatum istarum usque ad Baal haec est habitatio eorum et sedum distributio
1CHR|4|34|Masobab quoque et Iemlech et Iosa filius Amasiae
1CHR|4|35|et Iohel et Ieu filius Iosabiae filii Saraiae filii Asihel
1CHR|4|36|et Helioenai et Iacoba et Isuaia et Asaia et Adihel et Isimihel et Banaia
1CHR|4|37|Ziza quoque filius Sephei filii Allon filii Idaia filii Semri filii Samaia
1CHR|4|38|isti sunt nominati principes in cognationibus suis et in domo adfinitatum suarum multiplicati sunt vehementer
1CHR|4|39|et profecti sunt ut ingrederentur in Gador usque ad orientem vallis et ut quaererent pascua gregibus suis
1CHR|4|40|inveneruntque pascuas uberes et valde bonas et terram latissimam et quietam et fertilem in qua ante habitaverunt de stirpe Ham
1CHR|4|41|hii ergo venerunt quos supra descripsimus nominatim in diebus Ezechiae regis Iuda et percusserunt tabernacula eorum et habitatores qui inventi fuerant ibi et deleverunt eos usque in praesentem diem habitaveruntque pro eis quoniam uberrimas ibidem pascuas reppererunt
1CHR|4|42|de filiis quoque Symeon abierunt in montem Seir viri quingenti habentes principes Phaltiam et Nahariam et Raphaiam et Ozihel filios Iesi
1CHR|4|43|et percusserunt reliquias quae evadere potuerant Amalechitarum et habitaverunt ibi pro eis usque ad diem hanc
1CHR|5|1|filii quoque Ruben primogeniti Israhel ipse quippe fuit primogenitus eius sed cum violasset torum patris sui data sunt primogenita eius filiis Ioseph filii Israhel et non est ille reputatus in primogenitum
1CHR|5|2|porro Iudas qui erat fortissimus inter fratres suos de stirpe eius principes germinati sunt primogenita autem reputata sunt Ioseph
1CHR|5|3|filii ergo Ruben primogeniti Israhel Enoch et Phallu Esrom et Charmi
1CHR|5|4|filii Iohel Samaia filius eius Gog filius eius Semei filius eius
1CHR|5|5|Micha filius eius Reeia filius eius Baal filius eius
1CHR|5|6|Beera filius eius quem captivum duxit Theglathphalnasar rex Assyriorum et fuit princeps in tribu Ruben
1CHR|5|7|fratres autem eius et universa cognatio quando numerabantur per familias suas habuerunt principes Ieihel et Zacchariam
1CHR|5|8|porro Bala filius Azaz filii Samma filii Iohel ipse habitavit in Aroer usque ad Nebo et Beelmeon
1CHR|5|9|contra orientalem quoque plagam habitavit usque ad introitum heremi et flumen Eufraten multum quippe iumentorum numerum possidebat in terra Galaad
1CHR|5|10|in diebus autem Saul proeliati sunt contra Agareos et interfecerunt illos habitaveruntque pro eis in tabernaculis eorum in omni plaga quae respicit ad orientem Galaad
1CHR|5|11|filii vero Gad e regione eorum habitaverunt in terra Basan usque Selcha
1CHR|5|12|Iohel in capite et Saphan secundus Ianai autem et Saphat in Basan
1CHR|5|13|fratres vero eorum secundum domos cognationum suarum Michahel et Mosollam et Sebe et Iori et Iachan et Zie et Heber septem
1CHR|5|14|hii filii Abiahil filii Uri filii Iaro filii Galaad filii Michahel filii Iesesi filii Ieddo filii Buz
1CHR|5|15|fratres quoque filii Abdihel filii Guni princeps domus in familiis suis
1CHR|5|16|et habitaverunt in Galaad et in Basan et in viculis eius et in cunctis suburbanis Saron usque ad terminos
1CHR|5|17|omnes hii numerati sunt in diebus Ioatham regis Iuda et in diebus Hieroboam regis Israhel
1CHR|5|18|filii Ruben et Gad et dimidiae tribus Manasse viri bellatores scuta portantes et gladios et tendentes arcum eruditique ad proelia quadraginta quattuor milia et septingenti sexaginta procedentes ad pugnam
1CHR|5|19|dimicaverunt contra Agarenos Iturei vero et Naphei et Nodab
1CHR|5|20|praebuerunt eis auxilium traditique sunt in manus eorum Agareni et universi qui fuerant cum eis quia Deum invocaverunt cum proeliarentur et exaudivit eos eo quod credidissent in eum
1CHR|5|21|ceperuntque omnia quae possederant camelorum quinquaginta milia et ovium ducenta quinquaginta milia asinos duo milia et animas hominum centum milia
1CHR|5|22|vulnerati autem multi corruerunt fuit enim bellum Domini habitaveruntque pro eis usque ad transmigrationem
1CHR|5|23|filii quoque dimidiae tribus Manasse possederunt terram a finibus Basan usque Baalhermon et Sanir et montem Hermon ingens quippe numerus erat
1CHR|5|24|et hii fuerunt principes domus cognationis eorum Epher et Iesi et Helihel Ezrihel et Hieremia et Odoia et Iedihel viri fortissimi et potentes et nominati duces in familiis suis
1CHR|5|25|reliquerunt autem Deum patrum suorum et fornicati sunt post deos populorum terrae quos abstulit Dominus coram eis
1CHR|5|26|et suscitavit Deus Israhel spiritum Ful regis Assyriorum et spiritum Theglathphalnasar regis Assur et transtulit Ruben et Gad et dimidium tribus Manasse et adduxit eos in Alae et Abor et Ara et fluvium Gozan usque ad diem hanc
1CHR|6|1|filii Levi Gersom Caath Merari
1CHR|6|2|filii Caath Amram Isaar Hebron et Ozihel
1CHR|6|3|filii Amram Aaron Moses et Maria filii Aaron Nadab et Abiu Eleazar et Ithamar
1CHR|6|4|Eleazar genuit Finees et Finees genuit Abisue
1CHR|6|5|Abisue vero genuit Bocci et Bocci genuit Ozi
1CHR|6|6|Ozi genuit Zaraiam et Zaraias genuit Meraioth
1CHR|6|7|porro Meraioth genuit Amariam et Amarias genuit Ahitob
1CHR|6|8|Ahitob genuit Sadoc Sadoc genuit Achimaas
1CHR|6|9|Achimaas genuit Azariam Azarias genuit Iohanan
1CHR|6|10|Iohanan genuit Azariam ipse est qui sacerdotio functus est in domo quam aedificavit Salomon in Hierusalem
1CHR|6|11|genuit autem Azarias Amariam et Amarias genuit Ahitob
1CHR|6|12|Ahitob genuit Sadoc et Sadoc genuit Sellum
1CHR|6|13|Sellum genuit Helciam et Helcias genuit Azariam
1CHR|6|14|Azarias genuit Saraiam et Saraias genuit Iosedec
1CHR|6|15|porro Iosedec egressus est quando transtulit Dominus Iudam et Hierusalem per manus Nabuchodonosor
1CHR|6|16|filii ergo Levi Gersom Caath et Merari
1CHR|6|17|et haec nomina filiorum Gersom Lobeni et Semei
1CHR|6|18|filii Caath Amram et Isaar et Hebron et Ozihel
1CHR|6|19|filii Merari Mooli et Musi hae autem cognationes Levi secundum familias eorum
1CHR|6|20|Gersom Lobeni filius eius Iaath filius eius Zamma filius eius
1CHR|6|21|Ioaa filius eius Addo filius eius Zara filius eius Iethrai filius eius
1CHR|6|22|filii Caath Aminadab filius eius Core filius eius Asir filius eius
1CHR|6|23|Helcana filius eius Abiasaph filius eius Asir filius eius
1CHR|6|24|Thaath filius eius Urihel filius eius Ozias filius eius Saul filius eius
1CHR|6|25|filii Helcana Amasai et Ahimoth
1CHR|6|26|Helcana filii Helcana Sophai filius eius Naath filius eius
1CHR|6|27|Heliab filius eius Hieroam filius eius Helcana filius eius
1CHR|6|28|filii Samuhel primogenitus Vasseni et Abia
1CHR|6|29|filii autem Merari Mooli Lobeni filius eius Semei filius eius Oza filius eius
1CHR|6|30|Samaa filius eius Aggia filius eius Asaia filius eius
1CHR|6|31|isti sunt quos constituit David super cantores domus Domini ex quo conlocata est arca
1CHR|6|32|et ministrabant coram tabernaculo testimonii canentes donec aedificaret Salomon domum Domini in Hierusalem stabant autem iuxta ordinem suum in ministerio
1CHR|6|33|hii vero sunt qui adsistebant cum filiis suis de filiis Caath Heman cantor filius Iohel filii Samuhel
1CHR|6|34|filii Helcana filii Hieroam filii Helihel filii Thou
1CHR|6|35|filii Suph filii Helcana filii Maath filii Amasai
1CHR|6|36|filii Helcana filii Iohel filii Azariae filii Sophoniae
1CHR|6|37|filii Thaath filii Asir filii Abiasaph filii Core
1CHR|6|38|filii Isaar filii Caath filii Levi filii Israhel
1CHR|6|39|et fratres eius Asaph qui stabat a dextris eius Asaph filius Barachiae filii Samaa
1CHR|6|40|filii Michahel filii Basiae filii Melchiae
1CHR|6|41|filii Athnai filii Zara filii Adaia
1CHR|6|42|filii Ethan filii Zamma filii Semei
1CHR|6|43|filii Ieth filii Gersom filii Levi
1CHR|6|44|filii autem Merari fratres eorum ad sinistram Ethan filius Cusi filii Abdi filii Maloch
1CHR|6|45|filii Asabiae filii Amasiae filii Helciae
1CHR|6|46|filii Amasai filii Bonni filii Somer
1CHR|6|47|filii Mooli filii Musi filii Merari filii Levi
1CHR|6|48|fratres quoque eorum Levitae qui ordinati sunt in cunctum ministerium tabernaculi domus Domini
1CHR|6|49|Aaron vero et filii eius adolebant incensum super altare holocausti et super altare thymiamatis in omne opus sancti sanctorum et ut precarentur pro Israhel iuxta omnia quae praecepit Moses servus Dei
1CHR|6|50|hii sunt autem filii Aaron Eleazar filius eius Finees filius eius Abisue filius eius
1CHR|6|51|Bocci filius eius Ozi filius eius Zaraia filius eius
1CHR|6|52|Meraioth filius eius Amaria filius eius Ahitob filius eius
1CHR|6|53|Sadoc filius eius Achimaas filius eius
1CHR|6|54|et haec habitacula eorum per vicos atque confinia filiorum scilicet Aaron iuxta cognationes Caathitarum ipsis enim sorte contigerat
1CHR|6|55|dederunt igitur eis Hebron in terra Iuda et suburbana eius per circuitum
1CHR|6|56|agros autem civitatis et villas Chaleb filio Iephonne
1CHR|6|57|porro filiis Aaron dederunt civitates ad confugiendum Hebron et Lobna et suburbana eius
1CHR|6|58|Iether quoque et Esthmo cum suburbanis suis sed et Helon et Dabir cum suburbanis suis
1CHR|6|59|Asan quoque et Bethsemes et suburbana eorum
1CHR|6|60|de tribu autem Beniamin Gabee et suburbana eius et Almath cum suburbanis suis Anathoth quoque cum suburbanis suis omnes civitates tredecim per cognationes suas
1CHR|6|61|filiis autem Caath residuis de cognatione sua dederunt ex dimidia tribu Manasse in possessionem urbes decem
1CHR|6|62|porro filiis Gersom per cognationes suas de tribu Isachar et de tribu Aser et de tribu Nepthali et de tribu Manasse in Basan urbes tredecim
1CHR|6|63|filiis autem Merari per cognationes suas de tribu Ruben et de tribu Gad et de tribu Zabulon dederunt sorte civitates duodecim
1CHR|6|64|dederunt quoque filii Israhel Levitis civitates et suburbana earum
1CHR|6|65|dederuntque per sortem ex tribu filiorum Iuda et ex tribu filiorum Symeon et ex tribu filiorum Beniamin urbes has quas vocaverunt nominibus suis
1CHR|6|66|et his qui erant ex cognatione filiorum Caath fueruntque civitates in terminis eorum de tribu Ephraim
1CHR|6|67|dederunt ergo eis urbes ad confugiendum Sychem cum suburbanis suis in monte Ephraim et Gazer cum suburbanis suis
1CHR|6|68|Hicmaam quoque cum suburbanis suis et Bethoron similiter
1CHR|6|69|necnon et Helon cum suburbanis suis et Gethremmon in eundem modum
1CHR|6|70|porro ex dimidia tribu Manasse Aner et suburbana eius Balaam et suburbana eius his videlicet qui de cognatione filiorum Caath reliqui erant
1CHR|6|71|filiis autem Gersom de cognatione dimidiae tribus Manasse Gaulon in Basan et suburbana eius et Astharoth cum suburbanis suis
1CHR|6|72|de tribu Isachar Cedes et suburbana eius et Dabereth cum suburbanis suis
1CHR|6|73|Ramoth quoque et suburbana illius et Anem cum suburbanis suis
1CHR|6|74|de tribu vero Aser Masal cum suburbanis suis et Abdon similiter
1CHR|6|75|Acac quoque et suburbana eius et Roob cum suburbanis suis
1CHR|6|76|porro de tribu Nepthali Cedes in Galilea et suburbana eius Amon cum suburbanis suis et Cariathaim et suburbana eius
1CHR|6|77|filiis autem Merari residuis de tribu Zabulon Remmono et suburbana eius et Thabor cum suburbanis suis
1CHR|6|78|trans Iordanem quoque ex adverso Hiericho contra orientem Iordanis de tribu Ruben Bosor in solitudine cum suburbanis suis et Iasa cum suburbanis suis
1CHR|6|79|Cademoth quoque et suburbana eius et Miphaath cum suburbanis suis
1CHR|6|80|necnon de tribu Gad Ramoth in Galaad et suburbana eius et Manaim cum suburbanis suis
1CHR|6|81|sed et Esbon cum suburbanis eius et Iezer cum suburbanis suis
1CHR|7|1|porro filii Isachar Thola et Phua Iasub et Samaron quattuor
1CHR|7|2|filii Thola Ozi et Raphaia et Ierihel et Iemai et Iebsem et Samuhel principes per domos cognationum suarum de stirpe Thola viri fortissimi numerati sunt in diebus David viginti duo milia sescenti
1CHR|7|3|filii Ozi Iezraia de quo nati sunt Michahel et Obadia et Iohel et Iesia quinque omnes principes
1CHR|7|4|cumque eis per familias et populos suos accincti ad proelium viri fortissimi triginta sex milia multas enim habuere uxores et filios
1CHR|7|5|fratresque eorum per omnem cognationem Isachar robustissimi ad pugnandum octoginta septem milia numerati sunt
1CHR|7|6|Beniamin Bale et Bochor et Iadihel tres
1CHR|7|7|filii Bale Esbon et Ozi et Ozihel et Ierimoth et Urai quinque principes familiarum et ad pugnandum robustissimi numerus autem eorum viginti duo milia et triginta quattuor
1CHR|7|8|porro filii Bochor Zamira et Ioas et Eliezer et Helioenai et Amri et Ierimoth et Abia et Anathoth et Almathan omnes hii filii Bochor
1CHR|7|9|numerati sunt autem per familias suas principes cognationum ad bella fortissimi viginti milia et ducenti
1CHR|7|10|porro filii Iadihel Balan filii autem Balan Hieus et Beniamin et Ahoth et Chanana et Iothan et Tharsis et Haisaar
1CHR|7|11|omnes hii filii Iadihel principes cognationum suarum viri fortissimi decem et septem milia et ducenti ad proelium procedentes
1CHR|7|12|Sephan quoque et Apham filii Hir et Asim filii Aer
1CHR|7|13|filii autem Nepthali Iasihel et Guni et Asar et Sellum filii Balaa
1CHR|7|14|porro filius Manasse Esrihel concubinaque eius syra peperit Machir patrem Galaad
1CHR|7|15|Machir autem accepit uxores filiis suis Happhim et Sepham et habuit sororem nomine Maacha nomen autem secundi Salphaad nataeque sunt Salphaad filiae
1CHR|7|16|et peperit Maacha uxor Machir filium vocavitque nomen eius Phares porro nomen fratris eius Sares et filii eius Ulam et Recem
1CHR|7|17|filius autem Ulam Badan hii sunt filii Galaad filii Machir filii Manasse
1CHR|7|18|soror autem eius Regina peperit virum Decorum et Abiezer et Moola
1CHR|7|19|erant autem filii Semida Ahin et Sechem et Leci et Aniam
1CHR|7|20|filii autem Ephraim Suthala Bareth filius eius Thaath filius eius Elada filius eius Thaath filius eius et huius filius Zabad
1CHR|7|21|et huius filius Suthala et huius filius Ezer et Elad occiderunt autem eos viri Geth indigenae quia descenderant ut invaderent possessiones eorum
1CHR|7|22|luxit igitur Ephraim pater eorum multis diebus et venerunt fratres eius ut consolarentur eum
1CHR|7|23|ingressusque est ad uxorem suam quae concepit et peperit filium et vocavit nomen eius Beria eo quod in malis domus eius ortus esset
1CHR|7|24|filia autem eius fuit Sara quae aedificavit Bethoron inferiorem et superiorem et Ozensara
1CHR|7|25|porro filius eius Rapha et Reseph et Thale de quo natus est Thaan
1CHR|7|26|qui genuit Laadan huius quoque filius Ammiud genuit Elisama
1CHR|7|27|de quo ortus est Nun qui habuit filium Iosue
1CHR|7|28|possessio autem eorum et habitatio Bethel cum filiabus suis et contra orientem Noran ad occidentalem plagam Gazer et filiae eius Sychem quoque cum filiabus suis usque Aza et filias eius
1CHR|7|29|iuxta filios quoque Manasse Bethsan et filias eius Thanach et filias eius Mageddo et filias eius Dor et filias eius in his habitaverunt filii Ioseph filii Israhel
1CHR|7|30|filii Aser Iomna et Iesua et Isui et Baria et Sara soror eorum
1CHR|7|31|filii autem Baria Heber et Melchihel ipse est pater Barzaith
1CHR|7|32|Heber autem genuit Iephlat et Somer et Otham et Suaa sororem eorum
1CHR|7|33|filii Iephlat Phosech et Chamaal et Asoth hii filii Iephlat
1CHR|7|34|porro filii Somer Ahi et Roaga et Iaba et Aram
1CHR|7|35|filii autem Helem fratris eius Supha et Iemna et Selles et Amal
1CHR|7|36|filii Supha Sue Arnaphed et Sual et Beri et Iamra
1CHR|7|37|Bosor et Od et Samma et Salusa et Iethran et Bera
1CHR|7|38|filii Iether Iephonne et Phaspha et Ara
1CHR|7|39|filii autem Olla Aree et Anihel et Resia
1CHR|7|40|omnes hii filii Aser principes cognationum electi atque fortissimi duces ducum numerus autem eorum aetatis quae apta esset ad bellum viginti sex milia
1CHR|8|1|Beniamin autem genuit Bale primogenitum suum Asbal secundum Ohora tertium
1CHR|8|2|Nuaha quartum et Rapha quintum
1CHR|8|3|fueruntque filii Bale Addaor et Gera et Abiud
1CHR|8|4|Abisue quoque et Neman et Ahoe
1CHR|8|5|sed et Gera et Sephuphan et Uram
1CHR|8|6|hii sunt filii Aod principes cognationum habitantium in Gabaa qui translati sunt in Manath
1CHR|8|7|Nooman autem et Achia et Gera ipse transtulit eos et genuit Oza et Ahiud
1CHR|8|8|porro Saarim genuit in regione Moab postquam dimisit Usim et Bara uxores suas
1CHR|8|9|genuit autem de Edes uxore sua Iobab et Sebia et Mosa et Molchom
1CHR|8|10|Iehus quoque et Sechia et Marma hii sunt filii eius principes in familiis suis
1CHR|8|11|Meusim vero genuit Abitob et Elphaal
1CHR|8|12|porro filii Elphaal Heber et Misaam et Samad hic aedificavit Ono et Lod et filias eius
1CHR|8|13|Bara autem et Samma principes cognationum habitantium in Aialon hii fugaverunt habitatores Geth
1CHR|8|14|et Haio et Sesac et Ierimoth
1CHR|8|15|et Zabadia et Arod et Eder
1CHR|8|16|Michahel quoque et Iespha et Ioaa filii Baria
1CHR|8|17|et Zabadia et Mosollam et Ezeci et Heber
1CHR|8|18|et Iesamari et Iezlia et Iobab filii Elphaal
1CHR|8|19|et Iacim et Zechri et Zabdi
1CHR|8|20|et Helioenai et Selethai et Helihel
1CHR|8|21|et Adaia et Baraia et Samarath filii Semei
1CHR|8|22|et Iesphan et Heber et Helihel
1CHR|8|23|et Abdon et Zechri et Hanan
1CHR|8|24|et Anania et Ailam et Anathothia
1CHR|8|25|et Iephdaia et Phanuhel filii Sesac
1CHR|8|26|et Samsari et Sooria et Otholia
1CHR|8|27|et Iersia et Helia et Zechri filii Ieroam
1CHR|8|28|hii patriarchae et cognationum principes qui habitaverunt in Hierusalem
1CHR|8|29|in Gabaon autem habitaverunt Abigabaon et nomen uxoris eius Maacha
1CHR|8|30|filiusque eius primogenitus Abdon et Sur et Cis et Baal et Nadab
1CHR|8|31|Gedor quoque et Ahio et Zacher
1CHR|8|32|et Macelloth genuit Samaa habitaveruntque ex adverso fratrum suorum in Hierusalem cum fratribus suis
1CHR|8|33|Ner autem genuit Cis et Cis genuit Saul porro Saul genuit Ionathan et Melchisuae et Abinadab et Esbaal
1CHR|8|34|filius autem Ionathan Meribbaal et Meribbaal genuit Micha
1CHR|8|35|filii Micha Phithon et Melech et Thara et Ahaz
1CHR|8|36|et Ahaz genuit Ioada et Ioada genuit Almoth et Azmoth et Zamari porro Zamari genuit Mosa
1CHR|8|37|et Mosa genuit Baana cuius filius fuit Rapha de quo ortus est Elasa qui genuit Asel
1CHR|8|38|porro Asel sex filii fuere his nominibus Ezricam Bochru Ismahel Saria Abadia Anan omnes hii filii Asel
1CHR|8|39|filii autem Esec fratris eius Ulam primogenitus et Us secundus et Eliphalet tertius
1CHR|8|40|fueruntque filii Ulam viri robustissimi et magno robore tendentes arcum et multos habentes filios ac nepotes usque ad centum quinquaginta omnes hii filii Beniamin
1CHR|9|1|universus ergo Israhel dinumeratus est et summa eorum scripta est in libro regum Israhel et Iuda translatique sunt in Babylonem propter delictum suum
1CHR|9|2|qui autem habitaverunt primi in possessionibus et in urbibus suis Israhel et sacerdotes Levitae et Nathinnei
1CHR|9|3|commorati sunt in Hierusalem de filiis Iuda et de filiis Beniamin de filiis quoque Ephraim et Manasse
1CHR|9|4|Othei filius Amiud filius Emri filii Omrai filii Bonni de filiis Phares filii Iuda
1CHR|9|5|et de Siloni Asaia primogenitus et filii eius
1CHR|9|6|de filiis autem Zara Ieuhel et fratres eorum sescenti nonaginta
1CHR|9|7|porro de filiis Beniamin Salo filius Mosollam filii Oduia filii Asana
1CHR|9|8|et Iobania filius Hieroam et Hela filius Ozi filii Mochori et Mosollam filius Saphatiae filii Rahuhel filii Iebaniae
1CHR|9|9|et fratres eorum per familias suas nongenti quinquaginta sex omnes hii principes cognationum per domos patrum suorum
1CHR|9|10|de sacerdotibus autem Iedaia Ioiarib et Iachin
1CHR|9|11|Azarias quoque filius Helciae filii Mosollam filii Sadoc filii Maraioth filii Ahitob pontifex domus Dei
1CHR|9|12|porro Adaias filius Hieroam filii Phasor filii Melchia et Masaia filius Adihel filii Iezra filii Mosollam filii Mosollamoth filii Emmer
1CHR|9|13|fratres quoque eorum principes per familias suas mille septingenti sexaginta fortissimi robore ad faciendum opus ministerii in domo Dei
1CHR|9|14|de Levitis autem Semeia filius Assub filii Ezricam filii Asebiu de filiis Merari
1CHR|9|15|Bacbacar quoque carpentarius et Galal et Mathania filius Micha filii Zechri filii Asaph
1CHR|9|16|et Obdia filius Semeiae filii Galal filii Idithun et Barachia filius Asa filii Helcana qui habitavit in atriis Netophathi
1CHR|9|17|ianitores autem Sellum et Acub et Telmon et Ahiman et frater eorum Sellum princeps
1CHR|9|18|usque ad illud tempus in porta Regis ad orientem observabant per vices suas de filiis Levi
1CHR|9|19|Sellum vero filius Core filii Abiasaph filii Core cum fratribus suis et domo patris sui hii sunt Coritae super opera ministerii custodes vestibulorum tabernaculi et familiae eorum per vices castrorum Domini custodientes introitum
1CHR|9|20|Finees autem filius Eleazar erat dux eorum coram Domino
1CHR|9|21|porro Zaccharias filius Mosollamia ianitor portae tabernaculi testimonii
1CHR|9|22|omnes hii electi in ostiarios per portas ducenti duodecim et descripti in villis propriis quos constituerunt David et Samuhel videns in fide sua
1CHR|9|23|tam ipsos quam filios eorum in ostiis domus Domini et in tabernaculo vicibus suis
1CHR|9|24|per quattuor ventos erant ostiarii id est ad orientem et ad occidentem ad aquilonem et ad austrum
1CHR|9|25|fratres autem eorum in viculis morabantur et veniebant in sabbatis suis de tempore usque ad tempus
1CHR|9|26|his quattuor Levitis creditus erat omnis numerus ianitorum et erant super exedras et thesauros domus Domini
1CHR|9|27|per gyrum quoque templi Domini morabantur in custodiis suis ut cum tempus fuisset ipsi mane aperirent fores
1CHR|9|28|de horum grege erant et super vasa ministerii ad numerum enim et inferebantur vasa et efferebantur
1CHR|9|29|de ipsis et qui credita habebant utensilia sanctuarii praeerant similae et vino et oleo et turi et aromatibus
1CHR|9|30|filii autem sacerdotum unguenta ex aromatibus conficiebant
1CHR|9|31|et Matthathias Levites primogenitus Sellum Coritae praefectus erat eorum quae in sartagine frigebantur
1CHR|9|32|porro de filiis Caath fratribus eorum super panes erant propositionis ut semper novos per singula sabbata praepararent
1CHR|9|33|hii sunt principes cantorum per familias Levitarum qui in exedris morabantur ita ut die et nocte iugiter suo ministerio deservirent
1CHR|9|34|capita Levitarum per familias suas principes manserunt in Hierusalem
1CHR|9|35|in Gabaon autem commorati sunt pater Gabaon Iaihel et nomen uxoris eius Maacha
1CHR|9|36|filius primogenitus eius Abdon et Sur et Cis et Baal et Ner et Nadab
1CHR|9|37|Gedor quoque et Ahio et Zaccharias et Macelloth
1CHR|9|38|porro Macelloth genuit Semmaam isti habitaverunt e regione fratrum suorum in Hierusalem cum fratribus suis
1CHR|9|39|Ner autem genuit Cis et Cis genuit Saul et Saul genuit Ionathan et Melchisuae et Abinadab et Esbaal
1CHR|9|40|filius autem Ionathan Meribbaal et Meribbaal genuit Micha
1CHR|9|41|porro filii Micha Phiton et Malech et Thara
1CHR|9|42|Ahaz autem genuit Iara et Iara genuit Alamath et Azmoth et Zamri et Zamri genuit Mosa
1CHR|9|43|Mosa vero genuit Baana cuius filius Raphaia genuit Elasa de quo ortus est Esel
1CHR|9|44|porro Esel sex filios habuit his nominibus Ezricam Bochru Ismahel Saria Obdia Anan hii filii Esel
1CHR|10|1|Philisthim autem pugnabant contra Israhel fugeruntque viri Israhel Palestinos et ceciderunt vulnerati in monte Gelboe
1CHR|10|2|cumque adpropinquassent Philisthei persequentes Saul et filios eius percusserunt Ionathan et Abinadab et Melchisuae filios Saul
1CHR|10|3|et adgravatum est proelium contra Saul inveneruntque eum sagittarii et vulneraverunt iaculis
1CHR|10|4|et dixit Saul ad armigerum suum evagina gladium tuum et interfice me ne forte veniant incircumcisi isti et inludant mihi noluit autem armiger eius hoc facere timore perterritus arripuit igitur Saul ensem et inruit in eum
1CHR|10|5|quod cum vidisset armiger eius videlicet mortuum esse Saul inruit etiam ipse in gladium suum et mortuus est
1CHR|10|6|interiit ergo Saul et tres filii eius et omnis domus illius pariter concidit
1CHR|10|7|quod cum vidissent viri Israhel qui habitabant in campestribus fugerunt et Saul ac filiis eius mortuis dereliquerunt urbes suas et huc illucque dispersi sunt veneruntque Philisthim et habitaverunt in eis
1CHR|10|8|die igitur altero detrahentes Philisthim spolia caesorum invenerunt Saul et filios eius iacentes in monte Gelboe
1CHR|10|9|cumque spoliassent eum et amputassent caput armisque nudassent miserunt in terram suam ut circumferretur et ostenderetur idolorum templis et populis
1CHR|10|10|arma autem eius consecraverunt in fano dei sui et caput adfixerunt in templo Dagon
1CHR|10|11|hoc cum audissent viri Iabesgalaad omnia scilicet quae Philisthim fecerunt super Saul
1CHR|10|12|consurrexerunt singuli virorum fortium et tulerunt cadavera Saul et filiorum eius adtuleruntque ea in Iabes et sepelierunt ossa eorum subter quercum quae erat in Iabes et ieiunaverunt septem diebus
1CHR|10|13|mortuus est ergo Saul propter iniquitates suas eo quod praevaricatus sit mandatum Domini quod praeceperat et non custodierit illud sed insuper etiam pythonissam consuluerit
1CHR|10|14|nec speraverit in Domino propter quod et interfecit eum et transtulit regnum eius ad David filium Isai
1CHR|11|1|congregatus est igitur omnis Israhel ad David in Hebron dicens os tuum sumus et caro tua
1CHR|11|2|heri quoque et nudius tertius cum adhuc regnaret Saul tu eras qui educebas et introducebas Israhel tibi enim dixit Dominus Deus tuus tu pasces populum meum Israhel et tu eris princeps super eum
1CHR|11|3|venerunt ergo omnes maiores natu Israhel ad regem in Hebron et iniit David cum eis foedus coram Domino unxeruntque eum regem super Israhel iuxta sermonem Domini quem locutus est in manu Samuhel
1CHR|11|4|abiit quoque David et omnis Israhel in Hierusalem haec est Iebus ubi erant Iebusei habitatores terrae
1CHR|11|5|dixeruntque qui habitabant in Iebus ad David non ingredieris huc porro David cepit arcem Sion quae est civitas David
1CHR|11|6|dixitque omnis qui percusserit Iebuseum in primis erit princeps et dux ascendit igitur primus Ioab filius Sarviae et factus est princeps
1CHR|11|7|habitavit autem David in arce et idcirco appellata est civitas David
1CHR|11|8|aedificavitque urbem in circuitu a Mello usque ad gyrum Ioab autem reliqua urbis extruxit
1CHR|11|9|proficiebatque David vadens et crescens et Dominus exercituum erat cum eo
1CHR|11|10|hii principes virorum fortium David qui adiuverunt eum ut rex fieret super omnem Israhel iuxta verbum Domini quod locutus est ad Israhel
1CHR|11|11|et iste numerus robustorum David Iesbaam filius Achamoni princeps inter triginta iste levavit hastam suam super trecentos vulneratos una vice
1CHR|11|12|et post eum Eleazar filius patrui eius Ahoites qui erat inter tres potentes
1CHR|11|13|iste fuit cum David in Aphesdommim quando Philisthim congregati sunt ad locum illum in proelium et erat ager regionis illius plenus hordeo fugeratque populus a facie Philisthinorum
1CHR|11|14|hic stetit in medio agri et defendit eum cumque percussisset Philistheos dedit Dominus salutem magnam populo suo
1CHR|11|15|descenderunt autem tres de triginta principibus ad petram in qua erat David ad speluncam Odollam quando Philisthim fuerant castrametati in valle Raphaim
1CHR|11|16|porro David erat in praesidio et statio Philisthinorum in Bethleem
1CHR|11|17|desideravit igitur David et dixit o si quis daret mihi aquam de cisterna Bethleem quae est in porta
1CHR|11|18|tres ergo isti per media castra Philisthinorum perrexerunt et hauserunt aquam de cisterna Bethleem quae erat in porta et adtulerunt ad David ut biberet qui noluit sed magis libavit illam Domino
1CHR|11|19|dicens absit ut in conspectu Dei mei hoc faciam et sanguinem virorum istorum bibam quia in periculo animarum suarum adtulerunt mihi aquam et ob hanc causam noluit bibere haec fecerunt tres robustissimi
1CHR|11|20|Abisai quoque frater Ioab ipse erat princeps trium et ipse levavit hastam suam contra trecentos vulneratos et ipse erat inter tres nominatissimus
1CHR|11|21|inter tres secundos inclitus et princeps eorum verumtamen usque ad tres primos non pervenerat
1CHR|11|22|Banaia filius Ioiadae viri robustissimi qui multa opera perpetrarat de Capsehel ipse percussit duos Arihel Moab et ipse descendit et interfecit leonem in media cisterna tempore nivis
1CHR|11|23|et ipse percussit virum aegyptium cuius statura erat quinque cubitorum et habebat lanceam ut liciatorium texentium descendit ergo ad eum cum virga et rapuit hastam quam tenebat manu et interfecit eum hasta sua
1CHR|11|24|haec fecit Banaia filius Ioiada qui erat inter tres robustos nominatissimus
1CHR|11|25|inter triginta primus verumtamen ad tres usque non pervenerat posuit autem eum David ad auriculam suam
1CHR|11|26|porro fortissimi in exercitu Asahel frater Ioab et Eleanan filius patrui eius de Bethleem
1CHR|11|27|Semmoth Arorites Helles Phallonites
1CHR|11|28|Iras filius Acces Thecuites Abiezer Anathothites
1CHR|11|29|Sobbochai Asothites Ilai Ahoites
1CHR|11|30|Marai Netophathites Heled filius Baana Netophathites
1CHR|11|31|Ethai filius Ribai de Gabaath filiorum Beniamin Banaia Pharathonites
1CHR|11|32|Uri de torrente Gaas Abial Arabathites Azmoth Bauramites Eliaba Salabonites
1CHR|11|33|filii Asom Gezonites Ionathan filius Sega Ararites
1CHR|11|34|Ahiam filius Sachar Ararites
1CHR|11|35|Eliphal filius Ur
1CHR|11|36|Apher Mechurathites Ahia Phellonites
1CHR|11|37|Asrai Carmelites Noorai filius Azbi
1CHR|11|38|Iohel frater Nathan Mabar filius Agarai
1CHR|11|39|Sellec Ammonites Noorai Berothites armiger Ioab filii Sarviae
1CHR|11|40|Iras Iethreus Gareb Iethreus
1CHR|11|41|Urias Ettheus Zabad filius Ooli
1CHR|11|42|Adina filius Seza Rubenites princeps Rubenitarum et cum eo triginta
1CHR|11|43|Hanan filius Maacha et Iosaphat Mathanites
1CHR|11|44|Ozias Astharothites Semma et Iaihel filii Hotam Aroerites
1CHR|11|45|Iedihel filius Samri et Ioha frater eius Thosaites
1CHR|11|46|Elihel Maumites et Ieribai et Iosaia filii Elnaem et Iethma Moabites Elihel et Obed et Iasihel de Masobia
1CHR|12|1|hii quoque venerunt ad David in Siceleg cum adhuc fugeret Saul filium Cis qui erant fortissimi et egregii pugnatores
1CHR|12|2|tendentes arcum et utraque manu fundis saxa iacientes et dirigentes sagittas de fratribus Saul ex Beniamin
1CHR|12|3|princeps Ahiezer et Ioas filii Sammaa Gabathites et Iazihel et Phallet filii Azmoth et Baracha et Ieu Anathothites
1CHR|12|4|Samaias quoque Gabaonites fortissimus inter triginta et super triginta Hieremias et Iezihel et Iohanan et Iezbad Gaderothites
1CHR|12|5|Eluzai et Ierimuth et Baalia et Samaria et Saphatia Aruphites
1CHR|12|6|Helcana et Iesia et Azrahel et Ioezer et Iesbaam de Careim
1CHR|12|7|Ioeela quoque et Zabadia filii Ieroam de Gedor
1CHR|12|8|sed et de Gaddi transfugerunt ad David cum lateret in deserto viri robustissimi et pugnatores optimi tenentes clypeum et hastam facies eorum quasi facies leonis et veloces quasi capreae in montibus
1CHR|12|9|Ezer princeps Obdias secundus Eliab tertius
1CHR|12|10|Masmana quartus Hieremias quintus
1CHR|12|11|Hetthi sextus Helihel septimus
1CHR|12|12|Iohanan octavus Helzebad nonus
1CHR|12|13|Hieremias decimus Bachannai undecimus
1CHR|12|14|hii de filiis Gad principes exercitus novissimus centum militibus praeerat et maximus mille
1CHR|12|15|isti sunt qui transierunt Iordanem mense primo quando inundare consuevit super ripas suas et omnes fugaverunt qui morabantur in vallibus ad orientalem plagam et occidentalem
1CHR|12|16|venerunt autem et de Beniamin et de Iuda ad praesidium in quo morabatur David
1CHR|12|17|egressusque est David obviam eis et ait si pacifice venistis ad me ut auxiliemini mihi cor meum iungatur vobis si autem insidiamini mihi pro adversariis meis cum ego iniquitatem in manibus non habeam videat Deus patrum nostrorum et iudicet
1CHR|12|18|spiritus vero induit Amessai principem inter triginta et ait tui sumus o David et tecum fili Isai pax pax tibi et pax adiutoribus tuis te enim adiuvat Deus tuus suscepit ergo eos David et constituit principes turmae
1CHR|12|19|porro de Manasse transfugerunt ad David quando veniebat cum Philisthim adversum Saul ut pugnaret et non dimicavit cum eis quia inito consilio remiserunt eum principes Philisthinorum dicentes periculo capitis nostri revertetur ad dominum suum Saul
1CHR|12|20|quando igitur reversus est in Siceleg transfugerunt ad eum de Manasse Ednas et Iozabad et Iedihel et Michahel et Iozabad et Heliu et Salathi principes milium in Manasse
1CHR|12|21|hii praebuerunt auxilium David adversum latrunculos omnes enim erant viri fortissimi et facti sunt principes in exercitu
1CHR|12|22|sed et per singulos dies veniebant ad David ad auxiliandum ei usque dum fieret grandis numerus quasi exercitus Dei
1CHR|12|23|iste quoque est numerus principum exercitus qui venerunt ad David cum esset in Hebron ut transferrent regnum Saul ad eum iuxta verbum Domini
1CHR|12|24|filii Iuda portantes clypeum et hastam sex milia octingenti expediti ad proelium
1CHR|12|25|de filiis Symeon virorum fortissimorum ad pugnandum septem milia centum
1CHR|12|26|de filiis Levi quattuor milia sescenti
1CHR|12|27|Ioiada quoque princeps de stirpe Aaron et cum eo tria milia septingenti
1CHR|12|28|Sadoc etiam puer egregiae indolis et domus patris eius principes viginti duo
1CHR|12|29|de filiis autem Beniamin fratribus Saul tria milia magna enim pars eorum adhuc sequebatur domum Saul
1CHR|12|30|porro de filiis Ephraim viginti milia octingenti fortissimi robore viri nominati in cognationibus suis
1CHR|12|31|et ex dimidia parte tribus Manasse decem et octo milia singuli per nomina sua venerunt ut constituerent regem David
1CHR|12|32|de filiis quoque Isachar viri eruditi qui norant singula tempora ad praecipiendum quid facere deberet Israhel principes ducenti omnis autem reliqua tribus eorum consilium sequebatur
1CHR|12|33|porro de Zabulon qui egrediebantur ad proelium et stabant in acie instructi armis bellicis quinquaginta milia venerunt in auxilium non in corde duplici
1CHR|12|34|et de Nepthali principes mille et cum eis instructa clypeo et hasta triginta septem milia
1CHR|12|35|de Dan etiam praeparata ad proelium viginti octo milia sescentorum
1CHR|12|36|et de Aser egredientes ad pugnam et in acie provocantes quadraginta milia
1CHR|12|37|trans Iordanem autem de filiis Ruben et Gad et dimidia parte tribus Manasse instructa armis bellicis centum viginti milia
1CHR|12|38|omnes isti viri bellatores et expediti ad pugnandum corde perfecto venerunt in Hebron ut constituerent regem David super universum Israhel sed et omnes reliqui ex Israhel uno corde erant ut rex fieret David
1CHR|12|39|fueruntque ibi apud David tribus diebus comedentes et bibentes praeparaverunt enim eis fratres sui
1CHR|12|40|sed et qui iuxta eos erant usque ad Isachar et Zabulon et Nepthalim adferebant panes in asinis et camelis et mulis et bubus ad vescendum farinam palatas uvam passam vinum oleum boves arietes ad omnem copiam gaudium quippe erat in Israhel
1CHR|13|1|iniit autem consilium David cum tribunis et centurionibus et universis principibus
1CHR|13|2|et ait ad omnem coetum Israhel si placet vobis et a Domino Deo nostro egreditur sermo quem loquor mittamus ad fratres nostros reliquos in universas regiones Israhel et ad sacerdotes et Levitas qui habitant in suburbanis urbium ut congregentur ad nos
1CHR|13|3|et reducamus arcam Dei nostri ad nos non enim requisivimus eam in diebus Saul
1CHR|13|4|et respondit universa multitudo ut ita fieret placuerat enim sermo omni populo
1CHR|13|5|congregavit ergo David cunctum Israhel a Sior Aegypti usque dum ingrediaris Emath ut adduceret arcam Dei de Cariathiarim
1CHR|13|6|et ascendit David et omnis vir Israhel ad collem Cariathiarim quae est in Iuda ut adferrent inde arcam Dei Domini sedentis super cherubin ubi invocatum est nomen eius
1CHR|13|7|inposueruntque arcam Dei super plaustrum novum de domo Aminadab Oza autem et fratres eius minabant plaustrum
1CHR|13|8|porro David et universus Israhel ludebant coram Deo omni virtute in canticis et in citharis et psalteriis et tympanis et cymbalis et tubis
1CHR|13|9|cum autem pervenissent ad aream Chidon tetendit Oza manum suam ut sustentaret arcam bos quippe lasciviens paululum inclinaverat eam
1CHR|13|10|iratus est itaque Dominus contra Ozam et percussit eum eo quod contigisset arcam et mortuus est ibi coram Deo
1CHR|13|11|contristatusque David eo quod divisisset Dominus Ozam vocavit locum illum Divisio Oza usque in praesentem diem
1CHR|13|12|et timuit Deum tunc temporis dicens quomodo possum ad me introducere arcam Dei
1CHR|13|13|et ob hanc causam non eam adduxit ad se hoc est in civitatem David sed avertit in domum Obededom Getthei
1CHR|13|14|mansit ergo arca Dei in domo Obededom tribus mensibus et benedixit Dominus domui eius et omnibus quae habebat
1CHR|14|1|misit quoque Hiram rex Tyri nuntios ad David et ligna cedrina et artifices parietum lignorumque ut aedificarent ei domum
1CHR|14|2|cognovitque David eo quod confirmasset eum Dominus in regem super Israhel et sublevatum esset regnum suum super populum eius Israhel
1CHR|14|3|accepit quoque David alias uxores in Hierusalem genuitque filios et filias
1CHR|14|4|et haec nomina eorum qui nati sunt ei in Hierusalem Sammu et Sobab Nathan et Salomon
1CHR|14|5|Iebar et Helisu et Eliphaleth
1CHR|14|6|Noga quoque et Napheg et Iaphiae
1CHR|14|7|Elisama et Baliada et Eliphaleth
1CHR|14|8|audientes autem Philisthim eo quod unctus esset David in regem super universum Israhel ascenderunt omnes ut quaererent eum quod cum audisset David egressus est obviam eis
1CHR|14|9|porro Philisthim venientes diffusi sunt in valle Raphaim
1CHR|14|10|consuluitque David Deum dicens si ascendam ad Philistheos si trades eos in manu mea et dixit ei Dominus ascende et tradam eos in manu tua
1CHR|14|11|cumque illi ascendissent in Baalpharasim percussit eos ibi David et dixit divisit Deus inimicos meos per manum meam sicuti dividuntur aquae et idcirco vocatum est nomen loci illius Baalpharasim
1CHR|14|12|dereliqueruntque ibi deos suos quos David iussit exuri
1CHR|14|13|alia etiam vice Philisthim inruerunt et diffusi sunt in valle
1CHR|14|14|consuluitque rursum David Deum et dixit ei Deus non ascendas post eos recede ab eis et venies contra illos ex adverso pirorum
1CHR|14|15|cumque audieris sonitum gradientis in cacumine pirorum tunc egredieris ad bellum egressus est enim Deus ante te ut percutiat castra Philisthim
1CHR|14|16|fecit ergo David sicut praeceperat ei Deus et percussit castra Philisthinorum de Gabaon usque Gazera
1CHR|14|17|divulgatumque est nomen David in universis regionibus et Dominus dedit pavorem eius super omnes gentes
1CHR|15|1|fecit quoque sibi domos in civitate David et aedificavit locum arcae Dei tetenditque ei tabernaculum
1CHR|15|2|tunc dixit David inlicitum est ut a quocumque portetur arca Dei nisi a Levitis quos elegit Dominus ad portandum eam et ad ministrandum sibi usque in aeternum
1CHR|15|3|congregavitque universum Israhel in Hierusalem ut adferretur arca Dei in locum suum quem praeparaverat ei
1CHR|15|4|necnon et filios Aaron et Levitas
1CHR|15|5|de filiis Caath Urihel princeps fuit et fratres eius centum viginti
1CHR|15|6|de filiis Merari Asaia princeps et fratres eius ducenti viginti
1CHR|15|7|de filiis Gersom Iohel princeps et fratres eius centum triginta
1CHR|15|8|de filiis Elisaphan Semeias princeps et fratres eius ducenti
1CHR|15|9|de filiis Hebron Elihel princeps et fratres eius octoginta
1CHR|15|10|de filiis Ozihel Aminadab princeps et fratres eius centum duodecim
1CHR|15|11|vocavitque David Sadoc et Abiathar sacerdotes et Levitas Urihel Asaiam Iohel Semeiam Elihel et Aminadab
1CHR|15|12|et dixit ad eos vos qui estis principes familiarum leviticarum sanctificamini cum fratribus vestris et adferte arcam Domini Dei Israhel ad locum qui ei praeparatus est
1CHR|15|13|ne ut a principio quia non eratis praesentes percussit nos Dominus sic et nunc fiat inlicitum quid nobis agentibus
1CHR|15|14|sanctificati sunt ergo sacerdotes et Levitae ut portarent arcam Domini Dei Israhel
1CHR|15|15|et tulerunt filii Levi arcam Dei sicut praeceperat Moses iuxta verbum Domini umeris suis in vectibus
1CHR|15|16|dixit quoque David principibus Levitarum ut constituerent de fratribus suis cantores in organis musicorum nablis videlicet et lyris et cymbalis ut resonaret in excelsum sonitus laetitiae
1CHR|15|17|constitueruntque Levitas Heman filium Iohel et de fratribus eius Asaph filium Barachiae de filiis vero Merari fratribus eorum Ethan filium Casaiae
1CHR|15|18|et cum eis fratres eorum in secundo ordine Zacchariam et Ben et Iazihel et Semiramoth et Iahihel et Ani Eliab et Banaiam et Maasiam et Matthathiam et Eliphalu et Macheniam et Obededom et Ieihel ianitores
1CHR|15|19|porro cantores Heman Asaph et Ethan in cymbalis aeneis concrepantes
1CHR|15|20|Zaccharias autem et Ozihel et Semiramoth et Iahihel et Ani et Eliab et Maasias et Banaias in nablis arcana cantabant
1CHR|15|21|porro Matthathias et Eliphalu et Machenias et Obededom et Ieihel et Ozaziu in citharis pro octava canebant epinikion
1CHR|15|22|Chonenias autem princeps Levitarum prophetiae praeerat ad praecinendam melodiam erat quippe valde sapiens
1CHR|15|23|et Barachias et Helcana ianitores arcae
1CHR|15|24|porro Sebenias et Iosaphat et Nathanahel et Amasai et Zaccharias et Banaias et Eliezer sacerdotes clangebant tubis coram arca Dei et Obededom et Ahias erant ianitores arcae
1CHR|15|25|igitur David et maiores natu Israhel et tribuni ierunt ad deportandam arcam foederis Domini de domo Obededom cum laetitia
1CHR|15|26|cumque adiuvisset Deus Levitas qui portabant arcam foederis Domini immolabantur septem tauri et septem arietes
1CHR|15|27|porro David erat indutus stola byssina et universi Levitae qui portabant arcam cantoresque et Chonenias princeps prophetiae inter cantores David autem indutus erat etiam ephod lineo
1CHR|15|28|universusque Israhel deducebant arcam foederis Domini in iubilo et sonitu bucinae et tubis et cymbalis et nablis et citharis concrepantes
1CHR|15|29|cumque pervenisset arca foederis Domini usque ad civitatem David Michol filia Saul prospiciens per fenestram vidit regem David saltantem atque ludentem et despexit eum in corde suo
1CHR|16|1|adtulerunt igitur arcam Dei et constituerunt eam in medio tabernaculi quod tetenderat ei David et obtulerunt holocausta et pacifica coram Deo
1CHR|16|2|cumque conplesset David offerens holocausta et pacifica benedixit populo in nomine Domini
1CHR|16|3|et divisit universis per singulos a viro usque ad mulierem tortam panis et partem assae carnis bubulae et frixam oleo similam
1CHR|16|4|constituitque coram arca Domini de Levitis qui ministrarent et recordarentur operum eius et glorificarent atque laudarent Dominum Deum Israhel
1CHR|16|5|Asaph principem et secundum eius Zacchariam porro Iahihel et Semiramoth et Ieihel et Matthathiam et Eliab et Banaiam et Obededom et Ieihel super organa psalterii et lyras Asaph autem ut cymbalis personaret
1CHR|16|6|Banaiam vero et Azihel sacerdotes canere tuba iugiter coram arca foederis Domini
1CHR|16|7|in illo die fecit David principem ad confitendum Domino Asaph et fratres eius
1CHR|16|8|confitemini Domino invocate nomen eius notas facite in populis adinventiones illius
1CHR|16|9|canite ei et psallite et narrate omnia mirabilia eius
1CHR|16|10|laudate nomen sanctum eius laetetur cor quaerentium Dominum
1CHR|16|11|quaerite Dominum et virtutem eius quaerite faciem eius semper
1CHR|16|12|recordamini mirabilium eius quae fecit signorum illius et iudiciorum oris eius
1CHR|16|13|semen Israhel servi eius filii Iacob electi illius
1CHR|16|14|ipse Dominus Deus noster in universa terra iudicia eius
1CHR|16|15|recordamini in sempiternum pacti eius sermonis quem praecepit in mille generationes
1CHR|16|16|quem pepigit cum Abraham et iuramenti illius cum Isaac
1CHR|16|17|et constituit illud Iacob in praeceptum et Israhel in pactum sempiternum
1CHR|16|18|dicens tibi dabo terram Chanaan funiculum hereditatis vestrae
1CHR|16|19|cum essent pauci numero parvi et coloni eius
1CHR|16|20|et transierunt de gente in gentem et de regno ad populum alterum
1CHR|16|21|non dimisit quemquam calumniari eos sed increpuit pro eis reges
1CHR|16|22|nolite tangere christos meos et in prophetis meis nolite malignari
1CHR|16|23|canite Domino omnis terra adnuntiate ex die in diem salutare eius
1CHR|16|24|narrate in gentibus gloriam eius in cunctis populis mirabilia illius
1CHR|16|25|quia magnus Dominus et laudabilis nimis et horribilis super omnes deos
1CHR|16|26|omnes enim dii populorum idola Dominus autem caelos fecit
1CHR|16|27|confessio et magnificentia coram eo fortitudo et gaudium in loco eius
1CHR|16|28|adferte Domino familiae populorum adferte Domino gloriam et imperium
1CHR|16|29|date Domino gloriam nomini eius levate sacrificium et venite in conspectu eius et adorate Dominum in decore sancto
1CHR|16|30|commoveatur a facie illius omnis terra ipse enim fundavit orbem inmobilem
1CHR|16|31|laetentur caeli et exultet terra et dicant in nationibus Dominus regnavit
1CHR|16|32|tonet mare et plenitudo eius exultent agri et omnia quae in eis sunt
1CHR|16|33|tunc laudabunt ligna saltus coram Domino quia venit iudicare terram
1CHR|16|34|confitemini Domino quoniam bonus quoniam in aeternum misericordia eius
1CHR|16|35|et dicite salva nos Deus salvator noster et congrega nos et erue de gentibus ut confiteamur nomini sancto tuo et exultemus in carminibus tuis
1CHR|16|36|benedictus Dominus Deus Israhel ab aeterno usque in aeternum et dicat omnis populus amen et hymnus Domino
1CHR|16|37|dereliquit itaque ibi coram arca foederis Domini Asaph et fratres eius ut ministrarent in conspectu arcae iugiter per singulos dies et vices suas
1CHR|16|38|porro Obededom et fratres eius sexaginta octo et Obededom filium Idithun et Osa constituit ianitores
1CHR|16|39|Sadoc autem sacerdotem et fratres illius sacerdotes coram tabernaculo Domini in excelso quod erat in Gabaon
1CHR|16|40|ut offerrent holocausta Domino super altare holocaustomatis iugiter mane et vespere iuxta omnia quae scripta sunt in lege Domini quam praecepit Israheli
1CHR|16|41|et post eum Heman et Idithun et reliquos electos unumquemque vocabulo suo ad confitendum Domino quoniam in aeternum misericordia eius
1CHR|16|42|Heman quoque et Idithun canentes tuba et quatientes cymbala et omnia musicorum organa ad canendum Deo filios autem Idithun fecit esse portarios
1CHR|16|43|reversusque est omnis populus in domum suam et David ut benediceret etiam domui suae
1CHR|17|1|cum autem habitaret David in domo sua dixit ad Nathan prophetam ecce ego habito in domo cedrina arca autem foederis Domini sub pellibus est
1CHR|17|2|et ait Nathan ad David omnia quae in corde tuo sunt fac Deus enim tecum est
1CHR|17|3|igitur nocte illa factus est sermo Dei ad Nathan dicens
1CHR|17|4|vade et loquere David servo meo haec dicit Dominus non aedificabis tu mihi domum ad habitandum
1CHR|17|5|neque enim mansi in domo ex eo tempore quo eduxi Israhel usque ad hanc diem sed fui semper mutans loca tabernaculi et in tentorio
1CHR|17|6|manens cum omni Israhel numquid locutus sum saltim uni iudicum Israhel quibus praeceperam ut pascerent populum meum et dixi quare non aedificastis mihi domum cedrinam
1CHR|17|7|nunc itaque sic loqueris ad servum meum David haec dicit Dominus exercituum ego tuli te cum in pascuis sequereris gregem ut esses dux populi mei Israhel
1CHR|17|8|et fui tecum quocumque perrexisti et interfeci omnes inimicos tuos coram te fecique tibi nomen quasi unius magnorum qui celebrantur in terra
1CHR|17|9|et dedi locum populo meo Israhel plantabitur et habitabit in eo et ultra non commovebitur nec filii iniquitatis adterent eos sicut a principio
1CHR|17|10|ex diebus quibus dedi iudices populo meo Israhel et humiliavi universos inimicos tuos adnuntio ergo tibi quod aedificaturus sit domum tibi Dominus
1CHR|17|11|cumque impleveris dies tuos ut vadas ad patres tuos suscitabo semen tuum post te quod erit de filiis tuis et stabiliam regnum eius
1CHR|17|12|ipse aedificabit mihi domum et firmabo solium eius usque in aeternum
1CHR|17|13|ego ero ei in patrem et ipse erit mihi in filium et misericordiam meam non auferam ab eo sicut abstuli ab eo qui ante te fuit
1CHR|17|14|et statuam eum in domo mea et in regno meo usque in sempiternum et thronus eius erit firmissimus in perpetuum
1CHR|17|15|iuxta omnia verba haec et iuxta universam visionem istam sic locutus est Nathan ad David
1CHR|17|16|cumque venisset rex David et sedisset coram Domino dixit quis ego sum Domine Deus et quae domus mea ut praestares mihi talia
1CHR|17|17|sed et hoc parum visum est in conspectu tuo ideoque locutus es super domum servi tui etiam in futurum et fecisti me spectabilem super omnes homines Domine Deus meus
1CHR|17|18|quid ultra addere potest David cum ita glorificaveris servum tuum et cognoveris eum
1CHR|17|19|Domine propter famulum tuum iuxta cor tuum fecisti omnem magnificentiam hanc et nota esse voluisti universa magnalia
1CHR|17|20|Domine non est similis tui et non est alius deus absque te ex omnibus quos audivimus auribus nostris
1CHR|17|21|quis autem est alius ut populus tuus Israhel gens una in terra ad quam perrexit Deus ut liberaret et faceret populum sibi et magnitudine sua atque terroribus eiceret nationes a facie eius quem de Aegypto liberarat
1CHR|17|22|et posuisti populum tuum Israhel tibi in populum usque in aeternum et tu Domine factus es Deus eius
1CHR|17|23|nunc igitur Domine sermo quem locutus es famulo tuo et super domum eius confirmetur in perpetuum et fac sicut locutus es
1CHR|17|24|permaneatque et magnificetur nomen tuum usque in sempiternum et dicatur Dominus exercituum Deus Israhel et domus David servi eius permanens coram eo
1CHR|17|25|tu enim Domine Deus meus revelasti auriculam servi tui ut aedificares ei domum et idcirco invenit servus tuus fiduciam ut oret coram te
1CHR|17|26|nunc ergo Domine tu es Deus et locutus es ad servum tuum tanta beneficia
1CHR|17|27|et coepisti benedicere domui servi tui ut sit semper coram te te enim Domine benedicente benedicta erit in perpetuum
1CHR|18|1|factum est autem post haec ut percuteret David Philisthim et humiliaret eos et tolleret Geth et filias eius de manu Philisthim
1CHR|18|2|percuteretque Moab et fierent Moabitae servi David offerentes ei munera
1CHR|18|3|eo tempore percussit David etiam Adadezer regem Suba regionis Emath quando perrexit ut dilataret imperium suum usque ad flumen Eufraten
1CHR|18|4|cepit ergo David mille quadrigas eius et septem milia equites ac viginti milia virorum peditum subnervavitque omnes equos curruum exceptis centum quadrigis quas reservavit sibi
1CHR|18|5|supervenit autem et Syrus damascenus ut auxilium praeberet Adadezer regi Suba sed et huius percussit David viginti duo milia virorum
1CHR|18|6|et posuit milites in Damasco ut Syria quoque serviret sibi et offerret munera adiuvitque eum Dominus in cunctis ad quae perrexerat
1CHR|18|7|tulit quoque David faretras aureas quas habuerant servi Adadezer et adtulit eas in Hierusalem
1CHR|18|8|necnon de Thebath et Chun urbibus Adadezer aeris plurimum de quo fecit Salomon mare aeneum et columnas et vasa aenea
1CHR|18|9|quod cum audisset Thou rex Emath percussisse videlicet David omnem exercitum Adadezer regis Suba
1CHR|18|10|misit Aduram filium suum ad regem David ut postularet ab eo pacem et congratularetur ei eo quod expugnasset et percussisset Adadezer adversarius quippe Thou erat Adadezer
1CHR|18|11|sed et omnia vasa aurea et argentea et aenea consecravit rex David Domino cum argento et auro quod tulerat ex universis gentibus tam de Idumea et Moab et filiis Ammon quam de Philisthim et Amalech
1CHR|18|12|Abisai vero filius Sarviae percussit Edom in valle Salinarum decem et octo milia
1CHR|18|13|et constituit in Edom praesidium ut serviret Idumea David salvavitque Dominus David in cunctis ad quae perrexerat
1CHR|18|14|regnavit ergo David super universum Israhel et faciebat iudicium atque iustitiam cuncto populo suo
1CHR|18|15|porro Ioab filius Sarviae erat super exercitum et Iosaphat filius Ahilud a commentariis
1CHR|18|16|Sadoc autem filius Ahitob et Ahimelech filius Abiathar sacerdotes et Susa scriba
1CHR|18|17|Banaias vero filius Ioiada super legiones Cherethi et Felethi porro filii David primi ad manum regis
1CHR|19|1|accidit autem ut moreretur Naas rex filiorum Ammon et regnaret filius eius pro eo
1CHR|19|2|dixitque David faciam misericordiam cum Hanon filio Naas praestitit enim pater eius mihi gratiam misitque David nuntios ad consolandum eum super morte patris sui qui cum pervenissent in terram filiorum Ammon ut consolarentur Hanon
1CHR|19|3|dixerunt principes filiorum Ammon ad Hanon tu forsitan putas quod David honoris causa in patrem tuum miserit qui consolentur te nec animadvertis quod ut explorent et investigent et scrutentur terram tuam venerint ad te servi eius
1CHR|19|4|igitur Hanon pueros David decalvavit et rasit et praecidit tunicas eorum a natibus usque ad pedes et dimisit eos
1CHR|19|5|qui cum abissent et hoc mandassent David misit in occursum eorum grandem enim contumeliam sustinuerant et praecepit ut manerent in Hiericho donec cresceret barba eorum et tunc reverterentur
1CHR|19|6|videntes autem filii Ammon quod iniuriam fecissent David tam Hanon quam reliquus populus miserunt mille talenta argenti ut conducerent sibi de Mesopotamia et de Syria Macha et de Suba currus et equites
1CHR|19|7|conduxeruntque triginta duo milia curruum et regem Macha cum populo eius qui cum venissent castrametati sunt e regione Medaba filii quoque Ammon congregati de urbibus suis venerunt ad bellum
1CHR|19|8|quod cum audisset David misit Ioab et omnem exercitum virorum fortium
1CHR|19|9|egressique filii Ammon direxerunt aciem iuxta portam civitatis reges autem qui ad auxilium venerant separatim in agro steterunt
1CHR|19|10|igitur Ioab intellegens bellum et ex adverso et post tergum contra se fieri elegit viros fortissimos de universo Israhel et perrexit contra Syrum
1CHR|19|11|reliquam autem partem populi dedit sub manu Abisai fratris sui et perrexerunt contra filios Ammon
1CHR|19|12|dixitque si vicerit me Syrus auxilio eris mihi sin autem superaverint te filii Ammon ero tibi in praesidium
1CHR|19|13|confortare et agamus viriliter pro populo nostro et pro urbibus Dei nostri Dominus autem quod in conspectu suo bonum est faciet
1CHR|19|14|perrexit ergo Ioab et populus qui cum eo erat contra Syrum ad proelium et fugavit eos
1CHR|19|15|porro filii Ammon videntes quod fugisset Syrus ipsi quoque fugerunt Abisai fratrem eius et ingressi sunt civitatem reversusque est etiam Ioab in Hierusalem
1CHR|19|16|videns autem Syrus quod cecidisset coram Israhel misit nuntios et adduxit Syrum qui erat trans Fluvium Sophach autem princeps militiae Adadezer erat dux eorum
1CHR|19|17|quod cum nuntiatum esset David congregavit universum Israhel et transivit Iordanem inruitque in eos et direxit ex adverso aciem illis contra pugnantibus
1CHR|19|18|fugit autem Syrus Israhel et interfecit David de Syris septem milia curruum et quadraginta milia peditum et Sophach exercitus principem
1CHR|19|19|videntes autem servi Adadezer se ab Israhel esse superatos transfugerunt ad David et servierunt ei noluitque ultra Syria auxilium praebere filiis Ammon
1CHR|20|1|factum est autem post anni circulum eo tempore quo solent reges ad bella procedere congregavit Ioab exercitum et robur militiae et vastavit terram filiorum Ammon perrexitque et obsedit Rabba porro David manebat in Hierusalem quando Ioab percussit Rabba et destruxit eam
1CHR|20|2|tulit autem David coronam Melchom de capite eius et invenit in ea auri pondo talentum et pretiosissimas gemmas fecitque sibi inde diadema manubias quoque urbis plurimas tulit
1CHR|20|3|populum autem qui erat in ea eduxit et fecit super eos tribulas et trahas et ferrata carpenta transire ita ut dissicarentur et contererentur sic fecit David cunctis urbibus filiorum Ammon et reversus est cum omni populo suo in Hierusalem
1CHR|20|4|post haec initum est bellum in Gazer adversus Philistheos in quo percussit Sobbochai Usathites Saphai de genere Raphaim et humiliavit eos
1CHR|20|5|aliud quoque bellum gestum est adversum Philistheos in quo percussit Adeodatus filius Saltus Lehemites fratrem Goliath Getthei cuius hastae lignum erat quasi liciatorium texentium
1CHR|20|6|sed et aliud bellum accidit in Geth in quo fuit homo longissimus habens digitos senos id est simul viginti quattuor qui et ipse de Rapha fuerat stirpe generatus
1CHR|20|7|hic blasphemavit Israhel et percussit eum Ionathan filius Sammaa fratris David hii sunt filii Rapha in Geth qui ceciderunt in manu David et servorum eius
1CHR|21|1|consurrexit autem Satan contra Israhel et incitavit David ut numeraret Israhel
1CHR|21|2|dixitque David ad Ioab et ad principes populi ite et numerate Israhel a Bersabee usque Dan et adferte mihi numerum ut sciam
1CHR|21|3|responditque Ioab augeat Dominus populum suum centuplum quam sunt nonne domine mi rex omnes servi tui sunt quare hoc quaerit dominus meus quod in peccatum reputetur Israheli
1CHR|21|4|sed sermo regis magis praevaluit egressusque est Ioab et circuivit universum Israhel et reversus est Hierusalem
1CHR|21|5|deditque David numerum eorum quos circumierat et inventus est omnis Israhel numerus mille milia et centum milia virorum educentium gladium de Iuda autem trecenta septuaginta milia bellatorum
1CHR|21|6|nam Levi et Beniamin non numeravit eo quod invitus exsequeretur regis imperium
1CHR|21|7|displicuit autem Deo quod iussum erat et percussit Israhel
1CHR|21|8|dixitque David ad Deum peccavi nimis ut hoc facerem obsecro aufer iniquitatem servi tui quia insipienter egi
1CHR|21|9|et locutus est Dominus ad Gad videntem David dicens
1CHR|21|10|vade et loquere ad David et dic haec dicit Dominus trium tibi optionem do unum quod volueris elige et faciam tibi
1CHR|21|11|cumque venisset Gad ad David dixit ei haec dicit Dominus elige quod volueris
1CHR|21|12|aut tribus annis pestilentiam aut tribus mensibus fugere te hostes tuos et gladium eorum non posse evadere aut tribus diebus gladium Domini et mortem versari in terra et angelum Domini interficere in universis finibus Israhel nunc igitur vide quid respondeam ei qui misit me
1CHR|21|13|et dixit David ad Gad ex omni parte me angustiae premunt sed melius mihi est ut incidam in manus Domini quia multae sunt miserationes eius quam in manus hominum
1CHR|21|14|misit ergo Dominus pestilentiam in Israhel et ceciderunt de Israhel septuaginta milia virorum
1CHR|21|15|misit quoque angelum in Hierusalem ut percuteret eam cumque percuteretur vidit Dominus et misertus est super magnitudinem mali et imperavit angelo qui percutiebat sufficit iam cesset manus tua porro angelus Domini stabat iuxta aream Ornan Iebusei
1CHR|21|16|levansque David oculos suos vidit angelum Domini stantem inter terram et caelum et evaginatum gladium in manu eius et versum contra Hierusalem et ceciderunt tam ipse quam maiores natu vestiti ciliciis et proni in terram
1CHR|21|17|dixitque David ad Deum nonne ego sum qui iussi ut numeraretur populus ego qui peccavi ego qui malum feci iste grex quid commeruit Domine Deus meus vertatur obsecro manus tua in me et in domum patris mei populus autem tuus non percutiatur
1CHR|21|18|angelus autem Domini praecepit Gad ut diceret David et ascenderet extrueretque altare Domino Deo in area Ornan Iebusei
1CHR|21|19|ascendit ergo David iuxta sermonem Gad quem locutus fuerat ex nomine Domini
1CHR|21|20|porro Ornan cum suspexisset et vidisset angelum quattuorque filii eius cum eo absconderunt se nam eo tempore terebat in area triticum
1CHR|21|21|igitur cum venisset David ad Ornan conspexit eum Ornan et processit ei obviam de area et adoravit illum pronus in terram
1CHR|21|22|dixitque ei David da mihi locum areae tuae ut aedificem in ea altare Domini ita ut quantum valet argenti accipias et cesset plaga a populo
1CHR|21|23|dixit autem Ornan ad David tolle et faciat dominus meus rex quodcumque ei placet sed et boves do in holocaustum et tribulas in ligna et triticum in sacrificium omnia libens praebeo
1CHR|21|24|dixitque ei rex David nequaquam ita fiet sed argentum dabo quantum valet neque enim tibi auferre debeo et sic offerre Domino holocausta gratuita
1CHR|21|25|dedit ergo David Ornan pro loco siclos auri iustissimi ponderis sescentos
1CHR|21|26|et aedificavit ibi altare Domino obtulitque holocausta et pacifica et invocavit Dominum et exaudivit eum in igne de caelo super altare holocausti
1CHR|21|27|praecepitque Dominus angelo et convertit gladium suum in vaginam
1CHR|21|28|protinus ergo David videns quod exaudisset eum Dominus in area Ornan Iebusei immolavit ibi victimas
1CHR|21|29|tabernaculum autem Domini quod fecerat Moses in deserto et altare holocaustorum ea tempestate erat in excelso Gabaon
1CHR|21|30|et non praevaluit David ire ad altare ut ibi obsecraret Deum nimio enim fuerat timore perterritus videns gladium angeli Domini
1CHR|22|1|dixitque David haec est domus Dei et hoc altare in holocaustum Israhel
1CHR|22|2|et praecepit ut congregarentur omnes proselyti de terra Israhel et constituit ex eis latomos ad caedendos lapides et poliendos ut aedificaretur domus Dei
1CHR|22|3|ferrum quoque plurimum ad clavos ianuarum et ad commissuras atque iuncturas praeparavit David et aeris pondus innumerabile
1CHR|22|4|ligna quoque cedrina non poterant aestimari quae Sidonii et Tyrii deportaverant ad David
1CHR|22|5|et dixit David Salomon filius meus puer parvulus est et delicatus domus autem quam aedificari volo Domino talis esse debet ut in cunctis regionibus nominetur praeparabo ergo ei necessaria et ob hanc causam ante mortem suam omnes paravit inpensas
1CHR|22|6|vocavitque Salomonem filium suum et praecepit ei ut aedificaret domum Domino Deo Israhel
1CHR|22|7|dixitque David ad Salomonem fili mi voluntatis meae fuit ut aedificarem domum nomini Domini Dei mei
1CHR|22|8|sed factus est ad me sermo Domini dicens multum sanguinem effudisti et plurima bella bellasti non poteris aedificare domum nomini meo tanto effuso sanguine coram me
1CHR|22|9|filius qui nascetur tibi et erit vir quietissimus faciam enim eum requiescere ab omnibus inimicis suis per circuitum et ob hanc causam pacificus vocabitur et pacem et otium dabo in Israhel cunctis diebus eius
1CHR|22|10|ipse aedificabit domum nomini meo et ipse erit mihi in filium et ego ero ei in patrem firmaboque solium regni eius super Israhel in aeternum
1CHR|22|11|nunc ergo fili mi sit Dominus tecum et prosperare et aedifica domum Domino Deo tuo sicut locutus est de te
1CHR|22|12|det quoque tibi Dominus prudentiam et sensum ut regere possis Israhel et custodire legem Domini Dei tui
1CHR|22|13|tunc enim proficere poteris si custodieris mandata et iudicia quae praecepit Dominus Mosi ut doceret Israhel confortare viriliter age ne timeas neque paveas
1CHR|22|14|ecce ego in paupertatula mea praeparavi inpensas domus Domini auri talenta centum milia et argenti mille milia talentorum aeris vero et ferri non est pondus vincitur enim numerus magnitudine ligna et lapides praeparavi ad universa inpendia
1CHR|22|15|habes quoque plurimos artifices latomos et cementarios artificesque lignorum et omnium artium ad faciendum opus prudentissimos
1CHR|22|16|in auro et argento aere et ferro cuius non est numerus surge igitur et fac et erit Dominus tecum
1CHR|22|17|praecepit quoque David cunctis principibus Israhel ut adiuvarent Salomonem filium suum
1CHR|22|18|cernitis inquiens quod Dominus Deus vester vobiscum sit et dederit vobis requiem per circuitum et tradiderit omnes inimicos in manu vestra et subiecta sit terra coram Domino et coram populo eius
1CHR|22|19|praebete igitur corda vestra et animas vestras ut quaeratis Dominum Deum vestrum et consurgite et aedificate sanctuarium Domino Deo ut introducatur arca foederis Domini et vasa Domino consecrata in domum quae aedificatur nomini Domini
1CHR|23|1|igitur David senex et plenus dierum regem constituit Salomonem filium suum super Israhel
1CHR|23|2|et congregavit omnes principes Israhel et sacerdotes atque Levitas
1CHR|23|3|numeratique sunt Levitae a triginta annis et supra et inventa sunt triginta octo milia virorum
1CHR|23|4|ex his electi sunt et distributi in ministerium domus Domini viginti quattuor milia praepositorum autem et iudicum sex milia
1CHR|23|5|porro quattuor milia ianitores et totidem psaltae canentes Domino in organis quae fecerat ad canendum
1CHR|23|6|et distribuit eos David per vices filiorum Levi Gersom videlicet et Caath et Merari
1CHR|23|7|Gersom Leedan et Semei
1CHR|23|8|filii Leedan princeps Ieihel et Zetham et Iohel tres
1CHR|23|9|filii Semei Salomith et Ozihel et Aran tres isti principes familiarum Leedan
1CHR|23|10|porro filii Semei Ieeth et Ziza et Iaus et Baria isti filii Semei quattuor
1CHR|23|11|erat autem Ieeth prior Ziza secundus porro Iaus et Baria non habuerunt plurimos filios et idcirco in una familia unaque domo conputati sunt
1CHR|23|12|filii Caath Amram et Isaar Hebron et Ozihel quattuor
1CHR|23|13|filii Amram Aaron et Moses separatusque est Aaron ut ministraret in sancto sanctorum ipse et filii eius in sempiternum et adoleret incensum Domino secundum ritum suum ac benediceret nomini eius in perpetuum
1CHR|23|14|Mosi quoque hominis Dei filii adnumerati sunt in tribu Levi
1CHR|23|15|filii Mosi Gersom et Eliezer
1CHR|23|16|filii Gersom Subuhel primus
1CHR|23|17|fuerunt autem filii Eliezer Roobia primus et non erant Eliezer filii alii porro filii Roobia multiplicati sunt nimis
1CHR|23|18|filii Isaar Salumith primus
1CHR|23|19|filii Hebron Ieriau primus Amarias secundus Iazihel tertius Iecmaam quartus
1CHR|23|20|filii Ozihel Micha primus Iesia secundus
1CHR|23|21|filii Merari Mooli et Musi filii Mooli Eleazar et Cis
1CHR|23|22|mortuus est autem Eleazar et non habuit filios sed filias acceperuntque eas filii Cis fratres earum
1CHR|23|23|filii Musi Mooli et Eder et Ierimuth tres
1CHR|23|24|hii filii Levi in cognationibus et familiis suis principes per vices et numerum capitum singulorum qui faciebant opera ministerii domus Domini a viginti annis et supra
1CHR|23|25|dixit enim David requiem dedit Dominus Deus Israhel populo suo et habitationem Hierusalem usque in aeternum
1CHR|23|26|nec erit officii Levitarum ut ultra portent tabernaculum et omnia vasa eius ad ministrandum
1CHR|23|27|iuxta praecepta quoque David novissima supputabitur numerus filiorum Levi a viginti annis et supra
1CHR|23|28|et erunt sub manu filiorum Aaron in cultum domus Domini in vestibulis et in exedris et in loco purificationis et in sanctuario et in universis operibus ministerii templi Domini
1CHR|23|29|sacerdotes autem super panes propositionis et ad similae sacrificium et ad lagana et azyma et sartaginem et ad ferventem similam et super omne pondus atque mensuram
1CHR|23|30|Levitae vero ut stent mane ad confitendum et canendum Domino similiterque ad vesperam
1CHR|23|31|tam in oblatione holocaustorum Domini quam in sabbatis et kalendis et sollemnitatibus reliquis iuxta numerum et caerimonias uniuscuiusque rei iugiter coram Domino
1CHR|23|32|et custodiant observationes tabernaculi foederis et ritum sanctuarii et observationem filiorum Aaron fratrum suorum ut ministrent in domo Domini
1CHR|24|1|porro filiis Aaron hae partitiones erunt filii Aaron Nadab et Abiu et Eleazar et Ithamar
1CHR|24|2|mortui sunt autem Nadab et Abiu ante patrem suum absque liberis sacerdotioque functus est Eleazar et Ithamar
1CHR|24|3|et divisit eos David id est Sadoc de filiis Eleazar et Ahimelech de filiis Ithamar secundum vices suas et ministerium
1CHR|24|4|inventique sunt multo plures filii Eleazar in principibus viris quam filii Ithamar divisit autem eis hoc est filiis Eleazar principes per familias sedecim et filiis Ithamar per familias et domos suas octo
1CHR|24|5|porro divisit utrasque inter se familias sortibus erant enim principes sanctuarii et principes Dei tam de filiis Eleazar quam de filiis Ithamar
1CHR|24|6|descripsitque eos Semeias filius Nathanahel scriba Levites coram rege et principibus et Sadoc sacerdote et Ahimelech filio Abiathar principibus quoque familiarum sacerdotalium et leviticarum unam domum quae ceteris praeerat Eleazar et alteram domum quae sub se habebat ceteros Ithamar
1CHR|24|7|exivit autem sors prima Ioiarib secunda Iedeiae
1CHR|24|8|tertia Arim quarta Seorim
1CHR|24|9|quinta Melchia sexta Maiman
1CHR|24|10|septima Accos octava Abia
1CHR|24|11|nona Hiesu decima Sechenia
1CHR|24|12|undecima Eliasib duodecima Iacim
1CHR|24|13|tertiadecima Oppa quartadecima Isbaal
1CHR|24|14|quintadecima Belga sextadecima Emmer
1CHR|24|15|septimadecima Ezir octavadecima Hapses
1CHR|24|16|nonadecima Phetheia vicesima Iezecel
1CHR|24|17|vicesima prima Iachin vicesima secunda Gamul
1CHR|24|18|vicesima tertia Dalaiau vicesima quarta Mazziau
1CHR|24|19|hae vices eorum secundum ministeria sua ut ingrediantur domum Domini et iuxta ritum suum sub manu Aaron patris eorum sicut praecepit Dominus Deus Israhel
1CHR|24|20|porro filiorum Levi qui reliqui fuerant de filiis Amram erat Subahel et filiis Subahel Iedeia
1CHR|24|21|de filiis quoque Roobiae princeps Iesias
1CHR|24|22|Isaaris vero Salemoth filiusque Salemoth Iaath
1CHR|24|23|filiusque eius Ieriahu Amarias secundus Iazihel tertius Iecmaam quartus
1CHR|24|24|filius Ozihel Micha filius Micha Samir
1CHR|24|25|frater Micha Iesia filiusque Iesiae Zaccharias
1CHR|24|26|filii Merari Mooli et Musi filius Ioziau Benno
1CHR|24|27|filius quoque Merari Oziau et Soem et Zacchur et Hebri
1CHR|24|28|porro Mooli filius Eleazar qui non habebat liberos
1CHR|24|29|filius vero Cis Ierahemel
1CHR|24|30|filii Musi Mooli Eder et Ierimoth isti filii Levi secundum domos familiarum suarum
1CHR|24|31|miseruntque et ipsi sortes contra fratres suos filios Aaron coram David rege et Sadoc et Ahimelech et principibus familiarum sacerdotalium et leviticarum tam maiores quam minores omnes sors aequaliter dividebat
1CHR|25|1|igitur David et magistratus exercitus secreverunt in ministerium filios Asaph et Heman et Idithun qui prophetarent in citharis et psalteriis et cymbalis secundum numerum suum dedicato sibi officio servientes
1CHR|25|2|de filiis Asaph Zacchur et Ioseph et Nathania et Asarela filii Asaph sub manu Asaph prophetantis iuxta regem
1CHR|25|3|porro Idithun filii Idithun Godolias Sori Iesaias et Sabias et Matthathias sex sub manu patris sui Idithun qui in cithara prophetabat super confitentes et laudantes Dominum
1CHR|25|4|Heman quoque filii Heman Bocciau Matthaniau Ozihel Subuhel et Ierimoth Ananias Anani Elietha Geddelthi et Romemthiezer et Iesbacasa Mellothi Othir Mazioth
1CHR|25|5|omnes isti filii Heman videntis regis in sermonibus Dei ut exaltaret cornu deditque Deus Heman filios quattuordecim et filias tres
1CHR|25|6|universi sub manu patris sui ad cantandum in templo Domini distributi erant in cymbalis et psalteriis et citharis in ministeria domus Domini iuxta regem Asaph videlicet et Idithun et Heman
1CHR|25|7|fuit autem numerus eorum cum fratribus suis qui erudiebant canticum Domini cuncti doctores ducenti octoginta octo
1CHR|25|8|miseruntque sortes per vices suas ex aequo tam maior quam minor doctus pariter et indoctus
1CHR|25|9|egressaque est sors prima Ioseph qui erat de Asaph secunda Godoliae ipsi et filiis eius et fratribus duodecim
1CHR|25|10|tertia Zacchur filiis et fratribus eius duodecim
1CHR|25|11|quarta Isari filiis et fratribus eius duodecim
1CHR|25|12|quinta Nathaniae filiis et fratribus eius duodecim
1CHR|25|13|sexta Bocciau filiis et fratribus eius duodecim
1CHR|25|14|septima Israhela filiis et fratribus eius duodecim
1CHR|25|15|octava Isaiae filiis et fratribus eius duodecim
1CHR|25|16|nona Matthaniae filiis et fratribus eius duodecim
1CHR|25|17|decima Semeiae filiis et fratribus eius duodecim
1CHR|25|18|undecima Ezrahel filiis et fratribus eius duodecim
1CHR|25|19|duodecima Asabiae filiis et fratribus eius duodecim
1CHR|25|20|tertiadecima Subahel filiis et fratribus eius duodecim
1CHR|25|21|quartadecima Matthathiae filiis et fratribus eius duodecim
1CHR|25|22|quintadecima Ierimoth filiis et fratribus eius duodecim
1CHR|25|23|sextadecima Ananiae filiis et fratribus eius duodecim
1CHR|25|24|septimadecima Iesbocasae filiis et fratribus eius duodecim
1CHR|25|25|octavadecima Anani filiis et fratribus eius duodecim
1CHR|25|26|nonadecima Mellothi filiis et fratribus eius duodecim
1CHR|25|27|vicesima Eliatha filiis et fratribus eius duodecim
1CHR|25|28|vicesima prima Othir filiis et fratribus eius duodecim
1CHR|25|29|vicesima secunda Godollathi filiis et fratribus eius duodecim
1CHR|25|30|vicesima tertia Maziuth filiis et fratribus eius duodecim
1CHR|25|31|vicesima quarta Romamthiezer filiis et fratribus eius duodecim
1CHR|26|1|divisiones autem ianitorum de Coritis Mesellemia filius Core de filiis Asaph
1CHR|26|2|filii Mesellemiae Zaccharias primogenitus Iadihel secundus Zabadias tertius Iathanahel quartus
1CHR|26|3|Ahilam quintus Iohanan sextus Helioenai septimus
1CHR|26|4|filii autem Obededom Semeias primogenitus Iozabad secundus Iohaa tertius Sachar quartus Nathanahel quintus
1CHR|26|5|Amihel sextus Isachar septimus Phollathi octavus quia benedixit illi Dominus
1CHR|26|6|Semeiae autem filio eius nati sunt filii praefecti familiarum suarum erant enim viri fortissimi
1CHR|26|7|filii ergo Semeiae Othni et Raphahel et Obedihel Zabad fratres eius viri fortissimi Heliu quoque et Samachias
1CHR|26|8|omnes hii de filiis Obededom ipsi et filii et fratres eorum fortissimi ad ministrandum sexaginta duo de Obededom
1CHR|26|9|porro Mesellamiae filii et fratres robustissimi decem et octo
1CHR|26|10|de Hosa autem id est de filiis Merari Semri princeps non enim habuerat primogenitum et idcirco posuerat eum pater eius in principem
1CHR|26|11|Helchias secundus Tabelias tertius Zaccharias quartus omnes hii filii et fratres Hosa tredecim
1CHR|26|12|hii divisi sunt in ianitores ut semper principes custodiarum sicut et fratres eorum ministrarent in domo Domini
1CHR|26|13|missae sunt autem sortes ex aequo et parvis et magnis per familias suas in unamquamque portarum
1CHR|26|14|cecidit igitur sors orientalis Selemiae porro Zacchariae filio eius viro prudentissimo et erudito sortito obtigit plaga septentrionalis
1CHR|26|15|Obededom vero et filiis eius ad austrum in qua parte domus erat seniorum concilium
1CHR|26|16|Sepphima et Hosa ad occidentem iuxta portam quae ducit ad viam ascensionis custodia contra custodiam
1CHR|26|17|ad orientem vero Levitae sex et ad aquilonem quattuor per diem atque ad meridiem similiter in die quattuor et ubi erat concilium bini et bini
1CHR|26|18|in cellulis quoque ianitorum ad occidentem quattuor in via binique per cellulas
1CHR|26|19|hae sunt divisiones ianitorum filiorum Core et Merari
1CHR|26|20|porro Achias erat super thesauros domus Dei ac vasa sanctorum
1CHR|26|21|filii Ledan filii Gersonni de Ledan principes familiarum Ledan et Gersonni Ieiheli
1CHR|26|22|filii Ieiheli Zathan et Iohel frater eius super thesauros domus Domini
1CHR|26|23|Amramitis et Isaaritis et Hebronitis et Ozihelitibus
1CHR|26|24|Subahel autem filius Gersom filii Mosi praepositus thesauris
1CHR|26|25|fratres quoque eius Eliezer cuius filius Raabia et huius filius Isaias et huius filius Ioram huius quoque filius Zechri sed et huius filius Selemith
1CHR|26|26|ipse Selemith et fratres eius super thesauros sanctorum quae sanctificavit David rex et principes familiarum et tribuni et centuriones et duces exercitus
1CHR|26|27|de bellis et manubiis proeliorum quae consecraverant ad instaurationem et supellectilem templi Domini
1CHR|26|28|haec autem universa sanctificavit Samuhel videns et Saul filius Cis et Abner filius Ner et Ioab filius Sarviae omnes qui sanctificaverunt ea per manum Salemith et fratrum eius
1CHR|26|29|Saaritis vero praeerat Chonenias et filii eius ad opera forinsecus super Israhel ad docendum et ad iudicandum eos
1CHR|26|30|porro de Hebronitis Asabias et fratres eius viri fortissimi mille septingenti praeerant Israheli trans Iordanem contra occidentem in cunctis operibus Domini et in ministerium regis
1CHR|26|31|Hebronitarum autem princeps fuit Hieria secundum familias et cognationes eorum quadragesimo anno regni David recensiti sunt et inventi viri fortissimi in Iazer Galaad
1CHR|26|32|fratresque eius robustioris aetatis duo milia septingenti principes familiarum praeposuit autem eos David rex Rubenitis et Gadditis et dimidio tribus Manasse in omne ministerium Dei et regis
1CHR|27|1|filii autem Israhel secundum numerum suum principes familiarum tribuni et centuriones et praefecti qui ministrabant regi iuxta turmas suas ingredientes et egredientes per singulos menses in anno viginti quattuor milibus singuli praeerant
1CHR|27|2|primae turmae in primo mense Isboam praeerat filius Zabdihel et sub eo viginti quattuor milia
1CHR|27|3|de filiis Phares princeps cunctorum principum in exercitu mense primo
1CHR|27|4|secundi mensis habebat turmam Dudi Ahohites et post se alterum nomine Macelloth qui regebat partem exercitus viginti quattuor milium
1CHR|27|5|dux quoque turmae tertiae in mense tertio erat Banaias filius Ioiadae sacerdos et in divisione sua viginti quattuor milia
1CHR|27|6|ipse est Banaias fortissimus inter triginta et super triginta praeerat autem turmae ipsius Amizabad filius eius
1CHR|27|7|quartus mense quarto Asahel frater Ioab et Zabadias filius eius post eum et in turma eius viginti quattuor milia
1CHR|27|8|quintus mense quinto princeps Samaoth Iezarites et in turma eius viginti quattuor milia
1CHR|27|9|sextus mense sexto Hira filius Acces Thecuites et in turma eius viginti quattuor milia
1CHR|27|10|septimus mense septimo Helles Phallonites de filiis Ephraim et in turma eius viginti quattuor milia
1CHR|27|11|octavus mense octavo Sobochai Asothites de stirpe Zarai et in turma eius viginti quattuor milia
1CHR|27|12|nonus mense nono Abiezer Anathothites de filiis Iemini et in turma eius viginti quattuor milia
1CHR|27|13|decimus mense decimo Marai et ipse Netophathites de stirpe Zarai et in turma eius viginti quattuor milia
1CHR|27|14|undecimus mense undecimo Banaias Pharathonites de filiis Ephraim et in turma eius viginti quattuor milia
1CHR|27|15|duodecimus mense duodecimo Holdai Netophathites de stirpe Gothonihel et in turma eius viginti quattuor milia
1CHR|27|16|porro tribubus praeerant Israhel Rubenitis dux Eliezer filius Zechri Symeonitis dux Saphatias filius Macha
1CHR|27|17|Levitis Asabias filius Camuhel Aaronitis Sadoc
1CHR|27|18|Iuda Heliu frater David Isachar Amri filius Michahel
1CHR|27|19|Zabulonitis Iesmaias filius Abdiae Nepthalitibus Ierimoth filius Ozihel
1CHR|27|20|filiis Ephraim Osee filius Ozaziu dimidio tribus Manasse Iohel filius Phadiae
1CHR|27|21|et dimidio tribus Manasse in Galaad Iaddo filius Zacchariae Beniamin autem Iasihel filius Abner
1CHR|27|22|Dan vero Ezrihel filius Hieroam hii principes filiorum Israhel
1CHR|27|23|noluit autem David numerare eos a viginti annis inferius quia dixerat Dominus ut multiplicaret Israhel quasi stellas caeli
1CHR|27|24|Ioab filius Sarviae coeperat numerare nec conplevit quia super hoc ira inruerat in Israhel et idcirco numerus eorum qui fuerant recensiti non est relatus in fastos regis David
1CHR|27|25|super thesauros autem regis fuit Azmoth filius Adihel his autem thesauris qui erant in urbibus et in vicis et in turribus praesidebat Ionathan filius Oziae
1CHR|27|26|operi autem rustico et agricolis qui exercebant terram praeerat Ezri filius Chelub
1CHR|27|27|vinearumque cultoribus Semeias Ramathites cellis autem vinariis Zabdias Aphonites
1CHR|27|28|nam super oliveta et ficeta quae erant in campestribus Balanan Gaderites super apothecas autem olei Ioas
1CHR|27|29|porro armentis quae pascebantur in Sarona praepositus fuit Setrai Saronites et super boves in vallibus Saphat filius Adli
1CHR|27|30|super camelos vero Ubil Ismahelites et super asinos Iadias Meronathites
1CHR|27|31|super oves quoque Iaziz Agarenus omnes hii principes substantiae regis David
1CHR|27|32|Ionathan autem patruus David consiliarius vir prudens et litteratus ipse et Iaihel filius Achamoni erant cum filiis regis
1CHR|27|33|Ahitophel etiam consiliarius regis et Husi Arachites amicus regis
1CHR|27|34|post Ahitophel fuit Ioiada filius Banaiae et Abiathar princeps autem exercitus regis erat Ioab
1CHR|28|1|convocavit igitur David omnes principes Israhel duces tribuum et praepositos turmarum qui ministrabant regi tribunos quoque et centuriones et qui praeerant substantiae et possessionibus regis filiosque suos cum eunuchis et potentes et robustissimos quosque in exercitu Hierusalem
1CHR|28|2|cumque surrexisset rex et stetisset ait audite me fratres mei et populus meus cogitavi ut aedificarem domum in qua requiesceret arca foederis Domini et scabillum pedum Dei nostri et ad aedificandum omnia praeparavi
1CHR|28|3|Deus autem dixit mihi non aedificabis domum nomini meo eo quod sis vir bellator et sanguinem fuderis
1CHR|28|4|sed elegit Dominus Deus Israhel me de universa domo patris mei ut essem rex super Israhel in sempiternum de Iuda enim elegit principes porro de domo Iuda domum patris mei et de filiis patris mei placuit ei ut me eligeret regem super cunctum Israhel
1CHR|28|5|sed et de filiis meis filios enim multos dedit mihi Dominus elegit Salomonem filium meum ut sederet in throno regni Domini super Israhel
1CHR|28|6|dixitque mihi Salomon filius tuus aedificabit domum meam et atria mea ipsum enim elegi mihi in filium et ego ero ei in patrem
1CHR|28|7|et firmabo regnum eius usque in aeternum si perseveraverit facere praecepta mea et iudicia sicut et hodie
1CHR|28|8|nunc igitur coram universo coetu Israhel audiente Deo nostro custodite et perquirite cuncta mandata Domini Dei nostri ut possideatis terram bonam et relinquatis eam filiis vestris post vos usque in sempiternum
1CHR|28|9|tu autem Salomon fili mi scito Deum patris tui et servi ei corde perfecto et animo voluntario omnia enim corda scrutatur Dominus et universas mentium cogitationes intellegit si quaesieris eum invenies si autem dereliqueris illum proiciet te in aeternum
1CHR|28|10|nunc ergo quia elegit te Dominus ut aedificares domum sanctuarii confortare et perfice
1CHR|28|11|dedit autem David Salomoni filio suo descriptionem porticus et templi et cellariorum et cenaculi et cubiculorum in adytis et domus propitiationis
1CHR|28|12|necnon et omnium quae cogitaverat atriorum et exedrarum per circuitum in thesauros domus Domini et in thesauros sanctorum
1CHR|28|13|divisionumque sacerdotalium et leviticarum in omnia opera domus Domini et in universa vasa ministerii templi Domini
1CHR|28|14|aurum in pondere per singula vasa ministerii argenti quoque pondus pro vasorum ad opera diversitate
1CHR|28|15|sed et ad candelabra aurea et ad lucernas eorum aurum pro mensura uniuscuiusque candelabri et lucernarum similiter et in candelabris argenteis et in lucernis eorum pro diversitate mensurae pondus argenti tradidit
1CHR|28|16|aurum quoque dedit in mensas propositionis pro diversitate mensarum similiter et argentum in alias mensas argenteas
1CHR|28|17|ad fuscinulas quoque et fialas et turibula ex auro purissimo et leunculos aureos pro qualitate mensurae pondus distribuit in leunculum et leunculum similiter et in leones argenteos diversum argenti pondus separavit
1CHR|28|18|altari autem in quo adoletur incensum aurum purissimum dedit ut ex ipso fieret similitudo quadrigae cherubin extendentium alas et velantium arcam foederis Domini
1CHR|28|19|omnia inquit venerunt scripta manu Domini ad me ut intellegerem universa opera exemplaris
1CHR|28|20|dixit quoque David Salomoni filio suo viriliter age et confortare et fac ne timeas et ne paveas Dominus enim Deus meus tecum erit et non dimittet te nec derelinquet donec perficias omne opus ministerii domus Domini
1CHR|28|21|ecce divisiones sacerdotum et Levitarum in omne ministerium domus Domini adsistunt tibi et parati sunt et noverunt tam principes quam populus facere omnia praecepta tua
1CHR|29|1|locutusque est David rex ad omnem ecclesiam Salomonem filium meum unum elegit Deus adhuc puerum et tenellum opus autem grande est neque enim homini praeparatur habitatio sed Deo
1CHR|29|2|ego autem totis viribus meis praeparavi inpensas domus Dei mei aurum ad vasa aurea et argentum in argentea aes in aenea ferrum in ferrea lignum ad lignea lapides onychinos et quasi stibinos et diversorum colorum omnem pretiosum lapidem et marmor parium abundantissime
1CHR|29|3|et super haec quae obtuli in domum Dei mei de peculio meo aurum et argentum do in templum Dei mei exceptis his quae paravi in aedem sanctam
1CHR|29|4|tria milia talenta auri de auro Ophir et septem milia talentorum argenti probatissimi ad deaurandos parietes templi
1CHR|29|5|ut ubicumque opus est aurum de auro et ubicumque opus est argentum argenti opera fiant per manus artificum et si quis sponte offert impleat manum suam hodie et offerat quod voluerit Domino
1CHR|29|6|polliciti sunt itaque principes familiarum et proceres tribuum Israhel tribuni quoque et centuriones et principes possessionum regis
1CHR|29|7|dederuntque in opera domus Dei auri talenta quinque milia et solidos decem milia argenti talenta decem milia et aeris talenta decem et octo milia ferri quoque centum milia talentorum
1CHR|29|8|et apud quemcumque inventi sunt lapides dederunt in thesaurum domus Domini per manum Ieihel Gersonitis
1CHR|29|9|laetatusque est populus cum vota sponte promitterent quia corde toto offerebant ea Domino sed et David rex laetatus est gaudio magno
1CHR|29|10|et benedixit Domino coram universa multitudine et ait benedictus es Domine Deus Israhel patris nostri ab aeterno in aeternum
1CHR|29|11|tua est Domine magnificentia et potentia et gloria atque victoria et tibi laus cuncta enim quae in caelo sunt et in terra tua sunt tuum Domine regnum et tu es super omnes principes
1CHR|29|12|tuae divitiae et tua est gloria tu dominaris omnium in manu tua virtus et potentia in manu tua magnitudo et imperium omnium
1CHR|29|13|nunc igitur Deus noster confitemur tibi et laudamus nomen tuum inclitum
1CHR|29|14|quis ego et quis populus meus ut possimus haec tibi universa promittere tua sunt omnia et quae de manu tua accepimus dedimus tibi
1CHR|29|15|peregrini enim sumus coram te et advenae sicut omnes patres nostri dies nostri quasi umbra super terram et nulla est mora
1CHR|29|16|Domine Deus noster omnis haec copia quam paravimus ut aedificaretur domus nomini sancto tuo de manu tua est et tua sunt omnia
1CHR|29|17|scio Deus meus quod probes corda et simplicitatem diligas unde et ego in simplicitate cordis mei laetus obtuli universa haec et populum tuum qui hic reppertus est vidi cum ingenti gaudio tibi offerre donaria
1CHR|29|18|Domine Deus Abraham et Isaac et Israhel patrum nostrorum custodi in aeternum hanc voluntatem cordis eorum et semper in venerationem tui mens ista permaneat
1CHR|29|19|Salomoni quoque filio meo da cor perfectum ut custodiat mandata tua testimonia tua caerimonias tuas et faciat universa et aedificet aedem cuius inpensas paravi
1CHR|29|20|praecepit autem David universae ecclesiae benedicite Domino Deo nostro et benedixit omnis ecclesia Domino Deo patrum suorum et inclinaverunt se et adoraverunt Deum et deinde regem
1CHR|29|21|immolaveruntque victimas Domino et obtulerunt holocausta die sequenti tauros mille arietes mille agnos mille cum libaminibus suis et universo ritu abundantissime in omnem Israhel
1CHR|29|22|et comederunt et biberunt coram Domino in die illo cum grandi laetitia et unxerunt secundo Salomonem filium David unxerunt autem Domino in principem et Sadoc in pontificem
1CHR|29|23|seditque Salomon super solium Domini in regem pro David patre suo et cunctis placuit et paruit illi omnis Israhel
1CHR|29|24|sed et universi principes et potentes et cuncti filii regis David dederunt manum et subiecti fuerunt Salomoni regi
1CHR|29|25|magnificavit ergo Dominus Salomonem super omnem Israhel et dedit illi gloriam regni qualem nullus habuit ante eum rex Israhel
1CHR|29|26|igitur David filius Isai regnavit super universum Israhel
1CHR|29|27|et dies quibus regnavit super Israhel fuerunt quadraginta anni in Hebron regnavit septem annis et in Hierusalem triginta tribus
1CHR|29|28|et mortuus est in senectute bona plenus dierum et divitiis et gloria regnavitque Salomon filius eius pro eo
1CHR|29|29|gesta autem David regis priora et novissima scripta sunt in libro Samuhel videntis et in libro Nathan prophetae atque in volumine Gad videntis
1CHR|29|30|universique regni eius et fortitudinis et temporum quae transierunt sub eo sive in Israhel sive in cunctis regnis terrarum
