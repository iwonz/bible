HAG|1|1|大流士 王第二年六月初一，耶和华的话藉 哈该 先知向 撒拉铁 的儿子 犹大 省长 所罗巴伯 和 约撒答 的儿子 约书亚 大祭司传讲，说：
HAG|1|2|“万军之耶和华如此说，这百姓说，建造耶和华殿的时候还没有到 。”
HAG|1|3|耶和华的话藉 哈该 先知传讲，说：
HAG|1|4|“这殿荒凉，你们自己还住天花板的房屋吗？
HAG|1|5|现在，万军之耶和华如此说，你们要省察自己的行为。
HAG|1|6|你们撒的种多，收的却少；你们吃，却不得饱；喝，却不得足；穿衣服，却不得暖；领工钱的，领了工钱却装入有破洞的袋中。
HAG|1|7|“万军之耶和华如此说，你们要省察自己的行为。
HAG|1|8|你们要上山取木料，建造这殿，我就因此喜乐，且得荣耀。这是耶和华说的。
HAG|1|9|你们盼望多得，看哪，所得的却少；你们收到家中，我就吹去。这是为什么呢？因为我的殿荒凉，你们各人却只为自己的房屋奔走。这是万军之耶和华说的。
HAG|1|10|所以，因你们的缘故 ，天不降甘露，地也不出土产。
HAG|1|11|我命令干旱临到土地、山冈、五谷、新酒、新油和地上的出产，也临到人和牲畜，以及一切人手劳碌得来的。”
HAG|1|12|那时， 撒拉铁 的儿子 所罗巴伯 、 约撒答 的儿子 约书亚 大祭司，和所有幸存的百姓都听从耶和华－他们上帝的话，就是 哈该 先知奉耶和华－他们上帝差遣所说的话；百姓在耶和华面前存敬畏的心。
HAG|1|13|耶和华的使者 哈该 奉耶和华差遣对百姓说：“我与你们同在。这是耶和华说的。”
HAG|1|14|耶和华激发 撒拉铁 的儿子 犹大 省长 所罗巴伯 、 约撒答 的儿子 约书亚 大祭司，和所有幸存百姓的心，他们就来为万军之耶和华－他们上帝的殿做工。
HAG|1|15|这是在 大流士 王第二年六月二十四日。
HAG|2|1|七月二十一日，耶和华的话藉 哈该 先知传讲，说：
HAG|2|2|“你要晓谕 撒拉铁 的儿子 犹大 省长 所罗巴伯 、 约撒答 的儿子 约书亚 大祭司，和所有幸存的百姓，说：
HAG|2|3|‘你们中间存留的，有谁见过这殿从前的荣耀呢？现在你们看如何？在你们眼中岂不是如同无有吗？
HAG|2|4|所罗巴伯 啊，现在，你当刚强！这是耶和华说的。 约撒答 的儿子 约书亚 大祭司啊，你当刚强！这是耶和华说的。这地的百姓啊，你们都当刚强做工，因为我与你们同在。这是万军之耶和华说的。
HAG|2|5|这是照着你们出 埃及 时我与你们立约的话。我的灵仍要住在你们中间，你们不必惧怕。
HAG|2|6|万军之耶和华如此说：过些时候，我必再一次震动天地、沧海与干地。
HAG|2|7|我必震动万国，万国的珍宝都必运来 ，我就使这殿充满荣耀。这是万军之耶和华说的。
HAG|2|8|银子是我的，金子也是我的。这是万军之耶和华说的。
HAG|2|9|这后来的殿的荣耀必大过先前的荣耀。这是万军之耶和华说的。在这地方我必赐平安。这是万军之耶和华说的。’”
HAG|2|10|大流士 王第二年九月二十四日，耶和华的话临到 哈该 先知，说：
HAG|2|11|“万军之耶和华如此说，你要向祭司请教律法，说：
HAG|2|12|‘看哪，若有人用衣服的边兜圣肉，这衣服的边接触了饼，或汤，或酒，或油，或别的食物，这些是否成为圣呢？’”祭司回答说：“不。”
HAG|2|13|哈该 又说：“若有人因摸尸体染了不洁净，然后接触任何东西，这东西就变为不洁净吗？”祭司回答说：“必不洁净。”
HAG|2|14|于是 哈该 说：“耶和华说，在我面前这民如此，这国也是如此；他们手里的各样工作都是如此；他们在那里所献的都不洁净。”
HAG|2|15|“现在，你们心里要想一想，从今日起，耶和华的殿还没有一块石头放在石头上的情况。
HAG|2|16|那时你们怎么了？ 有人来到二十斗的谷堆那里，却只得了十斗；有人来到酒池那里要取五十桶，却只得了二十桶。
HAG|2|17|我以焚风 、霉烂、冰雹攻击你们，和你们手上的各样工作，你们仍不归向我。这是耶和华说的。
HAG|2|18|你们心里要想一想，从今日起，就是从这九月二十四日起，从立耶和华殿根基的日子起，你们心里想一想：
HAG|2|19|仓里还有谷种吗？葡萄树、无花果树、石榴树、橄榄树虽没有结果子， 从今日起，我必赐福。”
HAG|2|20|这月二十四日，耶和华的话再次临到 哈该 ，说：
HAG|2|21|“你要告诉 犹大 省长 所罗巴伯 说，我必震动天地，
HAG|2|22|倾覆列国的宝座，除灭列邦列国的势力，并倾覆战车和坐在其上的。马和骑兵都必跌倒，各人被弟兄的刀所杀。
HAG|2|23|万军之耶和华说： 撒拉铁 的儿子我仆人 所罗巴伯 啊，这是耶和华说的，到那日，我必以你为印，因我拣选了你。这是万军之耶和华说的。”
