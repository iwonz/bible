PROV|1|1|The proverbs of Solomon son of David, king of Israel:
PROV|1|2|for attaining wisdom and discipline; for understanding words of insight;
PROV|1|3|for acquiring a disciplined and prudent life, doing what is right and just and fair;
PROV|1|4|for giving prudence to the simple, knowledge and discretion to the young-
PROV|1|5|let the wise listen and add to their learning, and let the discerning get guidance-
PROV|1|6|for understanding proverbs and parables, the sayings and riddles of the wise.
PROV|1|7|The fear of the Lord is the beginning of knowledge, but fools despise wisdom and discipline.
PROV|1|8|Listen, my son, to your father's instruction and do not forsake your mother's teaching.
PROV|1|9|They will be a garland to grace your head and a chain to adorn your neck.
PROV|1|10|My son, if sinners entice you, do not give in to them.
PROV|1|11|If they say, "Come along with us; let's lie in wait for someone's blood, let's waylay some harmless soul;
PROV|1|12|let's swallow them alive, like the grave, and whole, like those who go down to the pit;
PROV|1|13|we will get all sorts of valuable things and fill our houses with plunder;
PROV|1|14|throw in your lot with us, and we will share a common purse"-
PROV|1|15|my son, do not go along with them, do not set foot on their paths;
PROV|1|16|for their feet rush into sin, they are swift to shed blood.
PROV|1|17|How useless to spread a net in full view of all the birds!
PROV|1|18|These men lie in wait for their own blood; they waylay only themselves!
PROV|1|19|Such is the end of all who go after ill-gotten gain; it takes away the lives of those who get it.
PROV|1|20|Wisdom calls aloud in the street, she raises her voice in the public squares;
PROV|1|21|at the head of the noisy streets she cries out, in the gateways of the city she makes her speech:
PROV|1|22|"How long will you simple ones love your simple ways? How long will mockers delight in mockery and fools hate knowledge?
PROV|1|23|If you had responded to my rebuke, I would have poured out my heart to you and made my thoughts known to you.
PROV|1|24|But since you rejected me when I called and no one gave heed when I stretched out my hand,
PROV|1|25|since you ignored all my advice and would not accept my rebuke,
PROV|1|26|I in turn will laugh at your disaster; I will mock when calamity overtakes you-
PROV|1|27|when calamity overtakes you like a storm, when disaster sweeps over you like a whirlwind, when distress and trouble overwhelm you.
PROV|1|28|"Then they will call to me but I will not answer; they will look for me but will not find me.
PROV|1|29|Since they hated knowledge and did not choose to fear the LORD,
PROV|1|30|since they would not accept my advice and spurned my rebuke,
PROV|1|31|they will eat the fruit of their ways and be filled with the fruit of their schemes.
PROV|1|32|For the waywardness of the simple will kill them, and the complacency of fools will destroy them;
PROV|1|33|but whoever listens to me will live in safety and be at ease, without fear of harm."
PROV|2|1|My son, if you accept my words and store up my commands within you,
PROV|2|2|turning your ear to wisdom and applying your heart to understanding,
PROV|2|3|and if you call out for insight and cry aloud for understanding,
PROV|2|4|and if you look for it as for silver and search for it as for hidden treasure,
PROV|2|5|then you will understand the fear of the LORD and find the knowledge of God.
PROV|2|6|For the LORD gives wisdom, and from his mouth come knowledge and understanding.
PROV|2|7|He holds victory in store for the upright, he is a shield to those whose walk is blameless,
PROV|2|8|for he guards the course of the just and protects the way of his faithful ones.
PROV|2|9|Then you will understand what is right and just and fair-every good path.
PROV|2|10|For wisdom will enter your heart, and knowledge will be pleasant to your soul.
PROV|2|11|Discretion will protect you, and understanding will guard you.
PROV|2|12|Wisdom will save you from the ways of wicked men, from men whose words are perverse,
PROV|2|13|who leave the straight paths to walk in dark ways,
PROV|2|14|who delight in doing wrong and rejoice in the perverseness of evil,
PROV|2|15|whose paths are crooked and who are devious in their ways.
PROV|2|16|It will save you also from the adulteress, from the wayward wife with her seductive words,
PROV|2|17|who has left the partner of her youth and ignored the covenant she made before God.
PROV|2|18|For her house leads down to death and her paths to the spirits of the dead.
PROV|2|19|None who go to her return or attain the paths of life.
PROV|2|20|Thus you will walk in the ways of good men and keep to the paths of the righteous.
PROV|2|21|For the upright will live in the land, and the blameless will remain in it;
PROV|2|22|but the wicked will be cut off from the land, and the unfaithful will be torn from it.
PROV|3|1|My son, do not forget my teaching, but keep my commands in your heart,
PROV|3|2|for they will prolong your life many years and bring you prosperity.
PROV|3|3|Let love and faithfulness never leave you; bind them around your neck, write them on the tablet of your heart.
PROV|3|4|Then you will win favor and a good name in the sight of God and man.
PROV|3|5|Trust in the LORD with all your heart and lean not on your own understanding;
PROV|3|6|in all your ways acknowledge him, and he will make your paths straight.
PROV|3|7|Do not be wise in your own eyes; fear the LORD and shun evil.
PROV|3|8|This will bring health to your body and nourishment to your bones.
PROV|3|9|Honor the LORD with your wealth, with the firstfruits of all your crops;
PROV|3|10|then your barns will be filled to overflowing, and your vats will brim over with new wine.
PROV|3|11|My son, do not despise the LORD's discipline and do not resent his rebuke,
PROV|3|12|because the LORD disciplines those he loves, as a father the son he delights in.
PROV|3|13|Blessed is the man who finds wisdom, the man who gains understanding,
PROV|3|14|for she is more profitable than silver and yields better returns than gold.
PROV|3|15|She is more precious than rubies; nothing you desire can compare with her.
PROV|3|16|Long life is in her right hand; in her left hand are riches and honor.
PROV|3|17|Her ways are pleasant ways, and all her paths are peace.
PROV|3|18|She is a tree of life to those who embrace her; those who lay hold of her will be blessed.
PROV|3|19|By wisdom the LORD laid the earth's foundations, by understanding he set the heavens in place;
PROV|3|20|by his knowledge the deeps were divided, and the clouds let drop the dew.
PROV|3|21|My son, preserve sound judgment and discernment, do not let them out of your sight;
PROV|3|22|they will be life for you, an ornament to grace your neck.
PROV|3|23|Then you will go on your way in safety, and your foot will not stumble;
PROV|3|24|when you lie down, you will not be afraid; when you lie down, your sleep will be sweet.
PROV|3|25|Have no fear of sudden disaster or of the ruin that overtakes the wicked,
PROV|3|26|for the LORD will be your confidence and will keep your foot from being snared.
PROV|3|27|Do not withhold good from those who deserve it, when it is in your power to act.
PROV|3|28|Do not say to your neighbor, "Come back later; I'll give it tomorrow"- when you now have it with you.
PROV|3|29|Do not plot harm against your neighbor, who lives trustfully near you.
PROV|3|30|Do not accuse a man for no reason- when he has done you no harm.
PROV|3|31|Do not envy a violent man or choose any of his ways,
PROV|3|32|for the LORD detests a perverse man but takes the upright into his confidence.
PROV|3|33|The LORD's curse is on the house of the wicked, but he blesses the home of the righteous.
PROV|3|34|He mocks proud mockers but gives grace to the humble.
PROV|3|35|The wise inherit honor, but fools he holds up to shame.
PROV|4|1|Listen, my sons, to a father's instruction; pay attention and gain understanding.
PROV|4|2|I give you sound learning, so do not forsake my teaching.
PROV|4|3|When I was a boy in my father's house, still tender, and an only child of my mother,
PROV|4|4|he taught me and said, "Lay hold of my words with all your heart; keep my commands and you will live.
PROV|4|5|Get wisdom, get understanding; do not forget my words or swerve from them.
PROV|4|6|Do not forsake wisdom, and she will protect you; love her, and she will watch over you.
PROV|4|7|Wisdom is supreme; therefore get wisdom. Though it cost all you have, get understanding.
PROV|4|8|Esteem her, and she will exalt you; embrace her, and she will honor you.
PROV|4|9|She will set a garland of grace on your head and present you with a crown of splendor."
PROV|4|10|Listen, my son, accept what I say, and the years of your life will be many.
PROV|4|11|I guide you in the way of wisdom and lead you along straight paths.
PROV|4|12|When you walk, your steps will not be hampered; when you run, you will not stumble.
PROV|4|13|Hold on to instruction, do not let it go; guard it well, for it is your life.
PROV|4|14|Do not set foot on the path of the wicked or walk in the way of evil men.
PROV|4|15|Avoid it, do not travel on it; turn from it and go on your way.
PROV|4|16|For they cannot sleep till they do evil; they are robbed of slumber till they make someone fall.
PROV|4|17|They eat the bread of wickedness and drink the wine of violence.
PROV|4|18|The path of the righteous is like the first gleam of dawn, shining ever brighter till the full light of day.
PROV|4|19|But the way of the wicked is like deep darkness; they do not know what makes them stumble.
PROV|4|20|My son, pay attention to what I say; listen closely to my words.
PROV|4|21|Do not let them out of your sight, keep them within your heart;
PROV|4|22|for they are life to those who find them and health to a man's whole body.
PROV|4|23|Above all else, guard your heart, for it is the wellspring of life.
PROV|4|24|Put away perversity from your mouth; keep corrupt talk far from your lips.
PROV|4|25|Let your eyes look straight ahead, fix your gaze directly before you.
PROV|4|26|Make level paths for your feet and take only ways that are firm.
PROV|4|27|Do not swerve to the right or the left; keep your foot from evil.
PROV|5|1|My son, pay attention to my wisdom, listen well to my words of insight,
PROV|5|2|that you may maintain discretion and your lips may preserve knowledge.
PROV|5|3|For the lips of an adulteress drip honey, and her speech is smoother than oil;
PROV|5|4|but in the end she is bitter as gall, sharp as a double-edged sword.
PROV|5|5|Her feet go down to death; her steps lead straight to the grave.
PROV|5|6|She gives no thought to the way of life; her paths are crooked, but she knows it not.
PROV|5|7|Now then, my sons, listen to me; do not turn aside from what I say.
PROV|5|8|Keep to a path far from her, do not go near the door of her house,
PROV|5|9|lest you give your best strength to others and your years to one who is cruel,
PROV|5|10|lest strangers feast on your wealth and your toil enrich another man's house.
PROV|5|11|At the end of your life you will groan, when your flesh and body are spent.
PROV|5|12|You will say, "How I hated discipline! How my heart spurned correction!
PROV|5|13|I would not obey my teachers or listen to my instructors.
PROV|5|14|I have come to the brink of utter ruin in the midst of the whole assembly."
PROV|5|15|Drink water from your own cistern, running water from your own well.
PROV|5|16|Should your springs overflow in the streets, your streams of water in the public squares?
PROV|5|17|Let them be yours alone, never to be shared with strangers.
PROV|5|18|May your fountain be blessed, and may you rejoice in the wife of your youth.
PROV|5|19|A loving doe, a graceful deer- may her breasts satisfy you always, may you ever be captivated by her love.
PROV|5|20|Why be captivated, my son, by an adulteress? Why embrace the bosom of another man's wife?
PROV|5|21|For a man's ways are in full view of the LORD, and he examines all his paths.
PROV|5|22|The evil deeds of a wicked man ensnare him; the cords of his sin hold him fast.
PROV|5|23|He will die for lack of discipline, led astray by his own great folly.
PROV|6|1|My son, if you have put up security for your neighbor, if you have struck hands in pledge for another,
PROV|6|2|if you have been trapped by what you said, ensnared by the words of your mouth,
PROV|6|3|then do this, my son, to free yourself, since you have fallen into your neighbor's hands: Go and humble yourself; press your plea with your neighbor!
PROV|6|4|Allow no sleep to your eyes, no slumber to your eyelids.
PROV|6|5|Free yourself, like a gazelle from the hand of the hunter, like a bird from the snare of the fowler.
PROV|6|6|Go to the ant, you sluggard; consider its ways and be wise!
PROV|6|7|It has no commander, no overseer or ruler,
PROV|6|8|yet it stores its provisions in summer and gathers its food at harvest.
PROV|6|9|How long will you lie there, you sluggard? When will you get up from your sleep?
PROV|6|10|A little sleep, a little slumber, a little folding of the hands to rest-
PROV|6|11|and poverty will come on you like a bandit and scarcity like an armed man.
PROV|6|12|A scoundrel and villain, who goes about with a corrupt mouth,
PROV|6|13|who winks with his eye, signals with his feet and motions with his fingers,
PROV|6|14|who plots evil with deceit in his heart- he always stirs up dissension.
PROV|6|15|Therefore disaster will overtake him in an instant; he will suddenly be destroyed-without remedy.
PROV|6|16|There are six things the LORD hates, seven that are detestable to him:
PROV|6|17|haughty eyes, a lying tongue, hands that shed innocent blood,
PROV|6|18|a heart that devises wicked schemes, feet that are quick to rush into evil,
PROV|6|19|a false witness who pours out lies and a man who stirs up dissension among brothers.
PROV|6|20|My son, keep your father's commands and do not forsake your mother's teaching.
PROV|6|21|Bind them upon your heart forever; fasten them around your neck.
PROV|6|22|When you walk, they will guide you; when you sleep, they will watch over you; when you awake, they will speak to you.
PROV|6|23|For these commands are a lamp, this teaching is a light, and the corrections of discipline are the way to life,
PROV|6|24|keeping you from the immoral woman, from the smooth tongue of the wayward wife.
PROV|6|25|Do not lust in your heart after her beauty or let her captivate you with her eyes,
PROV|6|26|for the prostitute reduces you to a loaf of bread, and the adulteress preys upon your very life.
PROV|6|27|Can a man scoop fire into his lap without his clothes being burned?
PROV|6|28|Can a man walk on hot coals without his feet being scorched?
PROV|6|29|So is he who sleeps with another man's wife; no one who touches her will go unpunished.
PROV|6|30|Men do not despise a thief if he steals to satisfy his hunger when he is starving.
PROV|6|31|Yet if he is caught, he must pay sevenfold, though it costs him all the wealth of his house.
PROV|6|32|But a man who commits adultery lacks judgment; whoever does so destroys himself.
PROV|6|33|Blows and disgrace are his lot, and his shame will never be wiped away;
PROV|6|34|for jealousy arouses a husband's fury, and he will show no mercy when he takes revenge.
PROV|6|35|He will not accept any compensation; he will refuse the bribe, however great it is.
PROV|7|1|My son, keep my words and store up my commands within you.
PROV|7|2|Keep my commands and you will live; guard my teachings as the apple of your eye.
PROV|7|3|Bind them on your fingers; write them on the tablet of your heart.
PROV|7|4|Say to wisdom, "You are my sister," and call understanding your kinsman;
PROV|7|5|they will keep you from the adulteress, from the wayward wife with her seductive words.
PROV|7|6|At the window of my house I looked out through the lattice.
PROV|7|7|I saw among the simple, I noticed among the young men, a youth who lacked judgment.
PROV|7|8|He was going down the street near her corner, walking along in the direction of her house
PROV|7|9|at twilight, as the day was fading, as the dark of night set in.
PROV|7|10|Then out came a woman to meet him, dressed like a prostitute and with crafty intent.
PROV|7|11|(She is loud and defiant, her feet never stay at home;
PROV|7|12|now in the street, now in the squares, at every corner she lurks.)
PROV|7|13|She took hold of him and kissed him and with a brazen face she said:
PROV|7|14|"I have fellowship offerings at home; today I fulfilled my vows.
PROV|7|15|So I came out to meet you; I looked for you and have found you!
PROV|7|16|I have covered my bed with colored linens from Egypt.
PROV|7|17|I have perfumed my bed with myrrh, aloes and cinnamon.
PROV|7|18|Come, let's drink deep of love till morning; let's enjoy ourselves with love!
PROV|7|19|My husband is not at home; he has gone on a long journey.
PROV|7|20|He took his purse filled with money and will not be home till full moon."
PROV|7|21|With persuasive words she led him astray; she seduced him with her smooth talk.
PROV|7|22|All at once he followed her like an ox going to the slaughter, like a deer stepping into a noose
PROV|7|23|till an arrow pierces his liver, like a bird darting into a snare, little knowing it will cost him his life.
PROV|7|24|Now then, my sons, listen to me; pay attention to what I say.
PROV|7|25|Do not let your heart turn to her ways or stray into her paths.
PROV|7|26|Many are the victims she has brought down; her slain are a mighty throng.
PROV|7|27|Her house is a highway to the grave, leading down to the chambers of death.
PROV|8|1|Does not wisdom call out? Does not understanding raise her voice?
PROV|8|2|On the heights along the way, where the paths meet, she takes her stand;
PROV|8|3|beside the gates leading into the city, at the entrances, she cries aloud:
PROV|8|4|"To you, O men, I call out; I raise my voice to all mankind.
PROV|8|5|You who are simple, gain prudence; you who are foolish, gain understanding.
PROV|8|6|Listen, for I have worthy things to say; I open my lips to speak what is right.
PROV|8|7|My mouth speaks what is true, for my lips detest wickedness.
PROV|8|8|All the words of my mouth are just; none of them is crooked or perverse.
PROV|8|9|To the discerning all of them are right; they are faultless to those who have knowledge.
PROV|8|10|Choose my instruction instead of silver, knowledge rather than choice gold,
PROV|8|11|for wisdom is more precious than rubies, and nothing you desire can compare with her.
PROV|8|12|"I, wisdom, dwell together with prudence; I possess knowledge and discretion.
PROV|8|13|To fear the LORD is to hate evil; I hate pride and arrogance, evil behavior and perverse speech.
PROV|8|14|Counsel and sound judgment are mine; I have understanding and power.
PROV|8|15|By me kings reign and rulers make laws that are just;
PROV|8|16|by me princes govern, and all nobles who rule on earth.
PROV|8|17|I love those who love me, and those who seek me find me.
PROV|8|18|With me are riches and honor, enduring wealth and prosperity.
PROV|8|19|My fruit is better than fine gold; what I yield surpasses choice silver.
PROV|8|20|I walk in the way of righteousness, along the paths of justice,
PROV|8|21|bestowing wealth on those who love me and making their treasuries full.
PROV|8|22|"The LORD brought me forth as the first of his works,, before his deeds of old;
PROV|8|23|I was appointed from eternity, from the beginning, before the world began.
PROV|8|24|When there were no oceans, I was given birth, when there were no springs abounding with water;
PROV|8|25|before the mountains were settled in place, before the hills, I was given birth,
PROV|8|26|before he made the earth or its fields or any of the dust of the world.
PROV|8|27|I was there when he set the heavens in place, when he marked out the horizon on the face of the deep,
PROV|8|28|when he established the clouds above and fixed securely the fountains of the deep,
PROV|8|29|when he gave the sea its boundary so the waters would not overstep his command, and when he marked out the foundations of the earth.
PROV|8|30|Then I was the craftsman at his side. I was filled with delight day after day, rejoicing always in his presence,
PROV|8|31|rejoicing in his whole world and delighting in mankind.
PROV|8|32|"Now then, my sons, listen to me; blessed are those who keep my ways.
PROV|8|33|Listen to my instruction and be wise; do not ignore it.
PROV|8|34|Blessed is the man who listens to me, watching daily at my doors, waiting at my doorway.
PROV|8|35|For whoever finds me finds life and receives favor from the LORD.
PROV|8|36|But whoever fails to find me harms himself; all who hate me love death."
PROV|9|1|Wisdom has built her house; she has hewn out its seven pillars.
PROV|9|2|She has prepared her meat and mixed her wine; she has also set her table.
PROV|9|3|She has sent out her maids, and she calls from the highest point of the city.
PROV|9|4|"Let all who are simple come in here!" she says to those who lack judgment.
PROV|9|5|"Come, eat my food and drink the wine I have mixed.
PROV|9|6|Leave your simple ways and you will live; walk in the way of understanding.
PROV|9|7|"Whoever corrects a mocker invites insult; whoever rebukes a wicked man incurs abuse.
PROV|9|8|Do not rebuke a mocker or he will hate you; rebuke a wise man and he will love you.
PROV|9|9|Instruct a wise man and he will be wiser still; teach a righteous man and he will add to his learning.
PROV|9|10|"The fear of the LORD is the beginning of wisdom, and knowledge of the Holy One is understanding.
PROV|9|11|For through me your days will be many, and years will be added to your life.
PROV|9|12|If you are wise, your wisdom will reward you; if you are a mocker, you alone will suffer."
PROV|9|13|The woman Folly is loud; she is undisciplined and without knowledge.
PROV|9|14|She sits at the door of her house, on a seat at the highest point of the city,
PROV|9|15|calling out to those who pass by, who go straight on their way.
PROV|9|16|"Let all who are simple come in here!" she says to those who lack judgment.
PROV|9|17|"Stolen water is sweet; food eaten in secret is delicious!"
PROV|9|18|But little do they know that the dead are there, that her guests are in the depths of the grave.
PROV|10|1|The proverbs of Solomon: A wise son brings joy to his father, but a foolish son grief to his mother.
PROV|10|2|Ill-gotten treasures are of no value, but righteousness delivers from death.
PROV|10|3|The LORD does not let the righteous go hungry but he thwarts the craving of the wicked.
PROV|10|4|Lazy hands make a man poor, but diligent hands bring wealth.
PROV|10|5|He who gathers crops in summer is a wise son, but he who sleeps during harvest is a disgraceful son.
PROV|10|6|Blessings crown the head of the righteous, but violence overwhelms the mouth of the wicked.
PROV|10|7|The memory of the righteous will be a blessing, but the name of the wicked will rot.
PROV|10|8|The wise in heart accept commands, but a chattering fool comes to ruin.
PROV|10|9|The man of integrity walks securely, but he who takes crooked paths will be found out.
PROV|10|10|He who winks maliciously causes grief, and a chattering fool comes to ruin.
PROV|10|11|The mouth of the righteous is a fountain of life, but violence overwhelms the mouth of the wicked.
PROV|10|12|Hatred stirs up dissension, but love covers over all wrongs.
PROV|10|13|Wisdom is found on the lips of the discerning, but a rod is for the back of him who lacks judgment.
PROV|10|14|Wise men store up knowledge, but the mouth of a fool invites ruin.
PROV|10|15|The wealth of the rich is their fortified city, but poverty is the ruin of the poor.
PROV|10|16|The wages of the righteous bring them life, but the income of the wicked brings them punishment.
PROV|10|17|He who heeds discipline shows the way to life, but whoever ignores correction leads others astray.
PROV|10|18|He who conceals his hatred has lying lips, and whoever spreads slander is a fool.
PROV|10|19|When words are many, sin is not absent, but he who holds his tongue is wise.
PROV|10|20|The tongue of the righteous is choice silver, but the heart of the wicked is of little value.
PROV|10|21|The lips of the righteous nourish many, but fools die for lack of judgment.
PROV|10|22|The blessing of the LORD brings wealth, and he adds no trouble to it.
PROV|10|23|A fool finds pleasure in evil conduct, but a man of understanding delights in wisdom.
PROV|10|24|What the wicked dreads will overtake him; what the righteous desire will be granted.
PROV|10|25|When the storm has swept by, the wicked are gone, but the righteous stand firm forever.
PROV|10|26|As vinegar to the teeth and smoke to the eyes, so is a sluggard to those who send him.
PROV|10|27|The fear of the LORD adds length to life, but the years of the wicked are cut short.
PROV|10|28|The prospect of the righteous is joy, but the hopes of the wicked come to nothing.
PROV|10|29|The way of the LORD is a refuge for the righteous, but it is the ruin of those who do evil.
PROV|10|30|The righteous will never be uprooted, but the wicked will not remain in the land.
PROV|10|31|The mouth of the righteous brings forth wisdom, but a perverse tongue will be cut out.
PROV|10|32|The lips of the righteous know what is fitting, but the mouth of the wicked only what is perverse.
PROV|11|1|The LORD abhors dishonest scales, but accurate weights are his delight.
PROV|11|2|When pride comes, then comes disgrace, but with humility comes wisdom.
PROV|11|3|The integrity of the upright guides them, but the unfaithful are destroyed by their duplicity.
PROV|11|4|Wealth is worthless in the day of wrath, but righteousness delivers from death.
PROV|11|5|The righteousness of the blameless makes a straight way for them, but the wicked are brought down by their own wickedness.
PROV|11|6|The righteousness of the upright delivers them, but the unfaithful are trapped by evil desires.
PROV|11|7|When a wicked man dies, his hope perishes; all he expected from his power comes to nothing.
PROV|11|8|The righteous man is rescued from trouble, and it comes on the wicked instead.
PROV|11|9|With his mouth the godless destroys his neighbor, but through knowledge the righteous escape.
PROV|11|10|When the righteous prosper, the city rejoices; when the wicked perish, there are shouts of joy.
PROV|11|11|Through the blessing of the upright a city is exalted, but by the mouth of the wicked it is destroyed.
PROV|11|12|A man who lacks judgment derides his neighbor, but a man of understanding holds his tongue.
PROV|11|13|A gossip betrays a confidence, but a trustworthy man keeps a secret.
PROV|11|14|For lack of guidance a nation falls, but many advisers make victory sure.
PROV|11|15|He who puts up security for another will surely suffer, but whoever refuses to strike hands in pledge is safe.
PROV|11|16|A kindhearted woman gains respect, but ruthless men gain only wealth.
PROV|11|17|A kind man benefits himself, but a cruel man brings trouble on himself.
PROV|11|18|The wicked man earns deceptive wages, but he who sows righteousness reaps a sure reward.
PROV|11|19|The truly righteous man attains life, but he who pursues evil goes to his death.
PROV|11|20|The LORD detests men of perverse heart but he delights in those whose ways are blameless.
PROV|11|21|Be sure of this: The wicked will not go unpunished, but those who are righteous will go free.
PROV|11|22|Like a gold ring in a pig's snout is a beautiful woman who shows no discretion.
PROV|11|23|The desire of the righteous ends only in good, but the hope of the wicked only in wrath.
PROV|11|24|One man gives freely, yet gains even more; another withholds unduly, but comes to poverty.
PROV|11|25|A generous man will prosper; he who refreshes others will himself be refreshed.
PROV|11|26|People curse the man who hoards grain, but blessing crowns him who is willing to sell.
PROV|11|27|He who seeks good finds goodwill, but evil comes to him who searches for it.
PROV|11|28|Whoever trusts in his riches will fall, but the righteous will thrive like a green leaf.
PROV|11|29|He who brings trouble on his family will inherit only wind, and the fool will be servant to the wise.
PROV|11|30|The fruit of the righteous is a tree of life, and he who wins souls is wise.
PROV|11|31|If the righteous receive their due on earth, how much more the ungodly and the sinner!
PROV|12|1|Whoever loves discipline loves knowledge, but he who hates correction is stupid.
PROV|12|2|A good man obtains favor from the LORD, but the LORD condemns a crafty man.
PROV|12|3|A man cannot be established through wickedness, but the righteous cannot be uprooted.
PROV|12|4|A wife of noble character is her husband's crown, but a disgraceful wife is like decay in his bones.
PROV|12|5|The plans of the righteous are just, but the advice of the wicked is deceitful.
PROV|12|6|The words of the wicked lie in wait for blood, but the speech of the upright rescues them.
PROV|12|7|Wicked men are overthrown and are no more, but the house of the righteous stands firm.
PROV|12|8|A man is praised according to his wisdom, but men with warped minds are despised.
PROV|12|9|Better to be a nobody and yet have a servant than pretend to be somebody and have no food.
PROV|12|10|A righteous man cares for the needs of his animal, but the kindest acts of the wicked are cruel.
PROV|12|11|He who works his land will have abundant food, but he who chases fantasies lacks judgment.
PROV|12|12|The wicked desire the plunder of evil men, but the root of the righteous flourishes.
PROV|12|13|An evil man is trapped by his sinful talk, but a righteous man escapes trouble.
PROV|12|14|From the fruit of his lips a man is filled with good things as surely as the work of his hands rewards him.
PROV|12|15|The way of a fool seems right to him, but a wise man listens to advice.
PROV|12|16|A fool shows his annoyance at once, but a prudent man overlooks an insult.
PROV|12|17|A truthful witness gives honest testimony, but a false witness tells lies.
PROV|12|18|Reckless words pierce like a sword, but the tongue of the wise brings healing.
PROV|12|19|Truthful lips endure forever, but a lying tongue lasts only a moment.
PROV|12|20|There is deceit in the hearts of those who plot evil, but joy for those who promote peace.
PROV|12|21|No harm befalls the righteous, but the wicked have their fill of trouble.
PROV|12|22|The LORD detests lying lips, but he delights in men who are truthful.
PROV|12|23|A prudent man keeps his knowledge to himself, but the heart of fools blurts out folly.
PROV|12|24|Diligent hands will rule, but laziness ends in slave labor.
PROV|12|25|An anxious heart weighs a man down, but a kind word cheers him up.
PROV|12|26|A righteous man is cautious in friendship, but the way of the wicked leads them astray.
PROV|12|27|The lazy man does not roast his game, but the diligent man prizes his possessions.
PROV|12|28|In the way of righteousness there is life; along that path is immortality.
PROV|13|1|A wise son heeds his father's instruction, but a mocker does not listen to rebuke.
PROV|13|2|From the fruit of his lips a man enjoys good things, but the unfaithful have a craving for violence.
PROV|13|3|He who guards his lips guards his life, but he who speaks rashly will come to ruin.
PROV|13|4|The sluggard craves and gets nothing, but the desires of the diligent are fully satisfied.
PROV|13|5|The righteous hate what is false, but the wicked bring shame and disgrace.
PROV|13|6|Righteousness guards the man of integrity, but wickedness overthrows the sinner.
PROV|13|7|One man pretends to be rich, yet has nothing; another pretends to be poor, yet has great wealth.
PROV|13|8|A man's riches may ransom his life, but a poor man hears no threat.
PROV|13|9|The light of the righteous shines brightly, but the lamp of the wicked is snuffed out.
PROV|13|10|Pride only breeds quarrels, but wisdom is found in those who take advice.
PROV|13|11|Dishonest money dwindles away, but he who gathers money little by little makes it grow.
PROV|13|12|Hope deferred makes the heart sick, but a longing fulfilled is a tree of life.
PROV|13|13|He who scorns instruction will pay for it, but he who respects a command is rewarded.
PROV|13|14|The teaching of the wise is a fountain of life, turning a man from the snares of death.
PROV|13|15|Good understanding wins favor, but the way of the unfaithful is hard.
PROV|13|16|Every prudent man acts out of knowledge, but a fool exposes his folly.
PROV|13|17|A wicked messenger falls into trouble, but a trustworthy envoy brings healing.
PROV|13|18|He who ignores discipline comes to poverty and shame, but whoever heeds correction is honored.
PROV|13|19|A longing fulfilled is sweet to the soul, but fools detest turning from evil.
PROV|13|20|He who walks with the wise grows wise, but a companion of fools suffers harm.
PROV|13|21|Misfortune pursues the sinner, but prosperity is the reward of the righteous.
PROV|13|22|A good man leaves an inheritance for his children's children, but a sinner's wealth is stored up for the righteous.
PROV|13|23|A poor man's field may produce abundant food, but injustice sweeps it away.
PROV|13|24|He who spares the rod hates his son, but he who loves him is careful to discipline him.
PROV|13|25|The righteous eat to their hearts' content, but the stomach of the wicked goes hungry.
PROV|14|1|The wise woman builds her house, but with her own hands the foolish one tears hers down.
PROV|14|2|He whose walk is upright fears the LORD, but he whose ways are devious despises him.
PROV|14|3|A fool's talk brings a rod to his back, but the lips of the wise protect them.
PROV|14|4|Where there are no oxen, the manger is empty, but from the strength of an ox comes an abundant harvest.
PROV|14|5|A truthful witness does not deceive, but a false witness pours out lies.
PROV|14|6|The mocker seeks wisdom and finds none, but knowledge comes easily to the discerning.
PROV|14|7|Stay away from a foolish man, for you will not find knowledge on his lips.
PROV|14|8|The wisdom of the prudent is to give thought to their ways, but the folly of fools is deception.
PROV|14|9|Fools mock at making amends for sin, but goodwill is found among the upright.
PROV|14|10|Each heart knows its own bitterness, and no one else can share its joy.
PROV|14|11|The house of the wicked will be destroyed, but the tent of the upright will flourish.
PROV|14|12|There is a way that seems right to a man, but in the end it leads to death.
PROV|14|13|Even in laughter the heart may ache, and joy may end in grief.
PROV|14|14|The faithless will be fully repaid for their ways, and the good man rewarded for his.
PROV|14|15|A simple man believes anything, but a prudent man gives thought to his steps.
PROV|14|16|A wise man fears the LORD and shuns evil, but a fool is hotheaded and reckless.
PROV|14|17|A quick-tempered man does foolish things, and a crafty man is hated.
PROV|14|18|The simple inherit folly, but the prudent are crowned with knowledge.
PROV|14|19|Evil men will bow down in the presence of the good, and the wicked at the gates of the righteous.
PROV|14|20|The poor are shunned even by their neighbors, but the rich have many friends.
PROV|14|21|He who despises his neighbor sins, but blessed is he who is kind to the needy.
PROV|14|22|Do not those who plot evil go astray? But those who plan what is good find love and faithfulness.
PROV|14|23|All hard work brings a profit, but mere talk leads only to poverty.
PROV|14|24|The wealth of the wise is their crown, but the folly of fools yields folly.
PROV|14|25|A truthful witness saves lives, but a false witness is deceitful.
PROV|14|26|He who fears the LORD has a secure fortress, and for his children it will be a refuge.
PROV|14|27|The fear of the LORD is a fountain of life, turning a man from the snares of death.
PROV|14|28|A large population is a king's glory, but without subjects a prince is ruined.
PROV|14|29|A patient man has great understanding, but a quick-tempered man displays folly.
PROV|14|30|A heart at peace gives life to the body, but envy rots the bones.
PROV|14|31|He who oppresses the poor shows contempt for their Maker, but whoever is kind to the needy honors God.
PROV|14|32|When calamity comes, the wicked are brought down, but even in death the righteous have a refuge.
PROV|14|33|Wisdom reposes in the heart of the discerning and even among fools she lets herself be known.
PROV|14|34|Righteousness exalts a nation, but sin is a disgrace to any people.
PROV|14|35|A king delights in a wise servant, but a shameful servant incurs his wrath.
PROV|15|1|A gentle answer turns away wrath, but a harsh word stirs up anger.
PROV|15|2|The tongue of the wise commends knowledge, but the mouth of the fool gushes folly.
PROV|15|3|The eyes of the LORD are everywhere, keeping watch on the wicked and the good.
PROV|15|4|The tongue that brings healing is a tree of life, but a deceitful tongue crushes the spirit.
PROV|15|5|A fool spurns his father's discipline, but whoever heeds correction shows prudence.
PROV|15|6|The house of the righteous contains great treasure, but the income of the wicked brings them trouble.
PROV|15|7|The lips of the wise spread knowledge; not so the hearts of fools.
PROV|15|8|The LORD detests the sacrifice of the wicked, but the prayer of the upright pleases him.
PROV|15|9|The LORD detests the way of the wicked but he loves those who pursue righteousness.
PROV|15|10|Stern discipline awaits him who leaves the path; he who hates correction will die.
PROV|15|11|Death and Destruction lie open before the LORD - how much more the hearts of men!
PROV|15|12|A mocker resents correction; he will not consult the wise.
PROV|15|13|A happy heart makes the face cheerful, but heartache crushes the spirit.
PROV|15|14|The discerning heart seeks knowledge, but the mouth of a fool feeds on folly.
PROV|15|15|All the days of the oppressed are wretched, but the cheerful heart has a continual feast.
PROV|15|16|Better a little with the fear of the LORD than great wealth with turmoil.
PROV|15|17|Better a meal of vegetables where there is love than a fattened calf with hatred.
PROV|15|18|A hot-tempered man stirs up dissension, but a patient man calms a quarrel.
PROV|15|19|The way of the sluggard is blocked with thorns, but the path of the upright is a highway.
PROV|15|20|A wise son brings joy to his father, but a foolish man despises his mother.
PROV|15|21|Folly delights a man who lacks judgment, but a man of understanding keeps a straight course.
PROV|15|22|Plans fail for lack of counsel, but with many advisers they succeed.
PROV|15|23|A man finds joy in giving an apt reply- and how good is a timely word!
PROV|15|24|The path of life leads upward for the wise to keep him from going down to the grave.
PROV|15|25|The LORD tears down the proud man's house but he keeps the widow's boundaries intact.
PROV|15|26|The LORD detests the thoughts of the wicked, but those of the pure are pleasing to him.
PROV|15|27|A greedy man brings trouble to his family, but he who hates bribes will live.
PROV|15|28|The heart of the righteous weighs its answers, but the mouth of the wicked gushes evil.
PROV|15|29|The LORD is far from the wicked but he hears the prayer of the righteous.
PROV|15|30|A cheerful look brings joy to the heart, and good news gives health to the bones.
PROV|15|31|He who listens to a life-giving rebuke will be at home among the wise.
PROV|15|32|He who ignores discipline despises himself, but whoever heeds correction gains understanding.
PROV|15|33|The fear of the LORD teaches a man wisdom, and humility comes before honor.
PROV|16|1|To man belong the plans of the heart, but from the LORD comes the reply of the tongue.
PROV|16|2|All a man's ways seem innocent to him, but motives are weighed by the LORD.
PROV|16|3|Commit to the LORD whatever you do, and your plans will succeed.
PROV|16|4|The LORD works out everything for his own ends- even the wicked for a day of disaster.
PROV|16|5|The LORD detests all the proud of heart. Be sure of this: They will not go unpunished.
PROV|16|6|Through love and faithfulness sin is atoned for; through the fear of the LORD a man avoids evil.
PROV|16|7|When a man's ways are pleasing to the LORD, he makes even his enemies live at peace with him.
PROV|16|8|Better a little with righteousness than much gain with injustice.
PROV|16|9|In his heart a man plans his course, but the LORD determines his steps.
PROV|16|10|The lips of a king speak as an oracle, and his mouth should not betray justice.
PROV|16|11|Honest scales and balances are from the LORD; all the weights in the bag are of his making.
PROV|16|12|Kings detest wrongdoing, for a throne is established through righteousness.
PROV|16|13|Kings take pleasure in honest lips; they value a man who speaks the truth.
PROV|16|14|A king's wrath is a messenger of death, but a wise man will appease it.
PROV|16|15|When a king's face brightens, it means life; his favor is like a rain cloud in spring.
PROV|16|16|How much better to get wisdom than gold, to choose understanding rather than silver!
PROV|16|17|The highway of the upright avoids evil; he who guards his way guards his life.
PROV|16|18|Pride goes before destruction, a haughty spirit before a fall.
PROV|16|19|Better to be lowly in spirit and among the oppressed than to share plunder with the proud.
PROV|16|20|Whoever gives heed to instruction prospers, and blessed is he who trusts in the LORD.
PROV|16|21|The wise in heart are called discerning, and pleasant words promote instruction.
PROV|16|22|Understanding is a fountain of life to those who have it, but folly brings punishment to fools.
PROV|16|23|A wise man's heart guides his mouth, and his lips promote instruction.
PROV|16|24|Pleasant words are a honeycomb, sweet to the soul and healing to the bones.
PROV|16|25|There is a way that seems right to a man, but in the end it leads to death.
PROV|16|26|The laborer's appetite works for him; his hunger drives him on.
PROV|16|27|A scoundrel plots evil, and his speech is like a scorching fire.
PROV|16|28|A perverse man stirs up dissension, and a gossip separates close friends.
PROV|16|29|A violent man entices his neighbor and leads him down a path that is not good.
PROV|16|30|He who winks with his eye is plotting perversity; he who purses his lips is bent on evil.
PROV|16|31|Gray hair is a crown of splendor; it is attained by a righteous life.
PROV|16|32|Better a patient man than a warrior, a man who controls his temper than one who takes a city.
PROV|16|33|The lot is cast into the lap, but its every decision is from the LORD.
PROV|17|1|Better a dry crust with peace and quiet than a house full of feasting, with strife.
PROV|17|2|A wise servant will rule over a disgraceful son, and will share the inheritance as one of the brothers.
PROV|17|3|The crucible for silver and the furnace for gold, but the LORD tests the heart.
PROV|17|4|A wicked man listens to evil lips; a liar pays attention to a malicious tongue.
PROV|17|5|He who mocks the poor shows contempt for their Maker; whoever gloats over disaster will not go unpunished.
PROV|17|6|Children's children are a crown to the aged, and parents are the pride of their children.
PROV|17|7|Arrogant lips are unsuited to a fool- how much worse lying lips to a ruler!
PROV|17|8|A bribe is a charm to the one who gives it; wherever he turns, he succeeds.
PROV|17|9|He who covers over an offense promotes love, but whoever repeats the matter separates close friends.
PROV|17|10|A rebuke impresses a man of discernment more than a hundred lashes a fool.
PROV|17|11|An evil man is bent only on rebellion; a merciless official will be sent against him.
PROV|17|12|Better to meet a bear robbed of her cubs than a fool in his folly.
PROV|17|13|If a man pays back evil for good, evil will never leave his house.
PROV|17|14|Starting a quarrel is like breaching a dam; so drop the matter before a dispute breaks out.
PROV|17|15|Acquitting the guilty and condemning the innocent- the LORD detests them both.
PROV|17|16|Of what use is money in the hand of a fool, since he has no desire to get wisdom?
PROV|17|17|A friend loves at all times, and a brother is born for adversity.
PROV|17|18|A man lacking in judgment strikes hands in pledge and puts up security for his neighbor.
PROV|17|19|He who loves a quarrel loves sin; he who builds a high gate invites destruction.
PROV|17|20|A man of perverse heart does not prosper; he whose tongue is deceitful falls into trouble.
PROV|17|21|To have a fool for a son brings grief; there is no joy for the father of a fool.
PROV|17|22|A cheerful heart is good medicine, but a crushed spirit dries up the bones.
PROV|17|23|A wicked man accepts a bribe in secret to pervert the course of justice.
PROV|17|24|A discerning man keeps wisdom in view, but a fool's eyes wander to the ends of the earth.
PROV|17|25|A foolish son brings grief to his father and bitterness to the one who bore him.
PROV|17|26|It is not good to punish an innocent man, or to flog officials for their integrity.
PROV|17|27|A man of knowledge uses words with restraint, and a man of understanding is even-tempered.
PROV|17|28|Even a fool is thought wise if he keeps silent, and discerning if he holds his tongue.
PROV|18|1|An unfriendly man pursues selfish ends; he defies all sound judgment.
PROV|18|2|A fool finds no pleasure in understanding but delights in airing his own opinions.
PROV|18|3|When wickedness comes, so does contempt, and with shame comes disgrace.
PROV|18|4|The words of a man's mouth are deep waters, but the fountain of wisdom is a bubbling brook.
PROV|18|5|It is not good to be partial to the wicked or to deprive the innocent of justice.
PROV|18|6|A fool's lips bring him strife, and his mouth invites a beating.
PROV|18|7|A fool's mouth is his undoing, and his lips are a snare to his soul.
PROV|18|8|The words of a gossip are like choice morsels; they go down to a man's inmost parts.
PROV|18|9|One who is slack in his work is brother to one who destroys.
PROV|18|10|The name of the LORD is a strong tower; the righteous run to it and are safe.
PROV|18|11|The wealth of the rich is their fortified city; they imagine it an unscalable wall.
PROV|18|12|Before his downfall a man's heart is proud, but humility comes before honor.
PROV|18|13|He who answers before listening- that is his folly and his shame.
PROV|18|14|A man's spirit sustains him in sickness, but a crushed spirit who can bear?
PROV|18|15|The heart of the discerning acquires knowledge; the ears of the wise seek it out.
PROV|18|16|A gift opens the way for the giver and ushers him into the presence of the great.
PROV|18|17|The first to present his case seems right, till another comes forward and questions him.
PROV|18|18|Casting the lot settles disputes and keeps strong opponents apart.
PROV|18|19|An offended brother is more unyielding than a fortified city, and disputes are like the barred gates of a citadel.
PROV|18|20|From the fruit of his mouth a man's stomach is filled; with the harvest from his lips he is satisfied.
PROV|18|21|The tongue has the power of life and death, and those who love it will eat its fruit.
PROV|18|22|He who finds a wife finds what is good and receives favor from the LORD.
PROV|18|23|A poor man pleads for mercy, but a rich man answers harshly.
PROV|18|24|A man of many companions may come to ruin, but there is a friend who sticks closer than a brother.
PROV|19|1|Better a poor man whose walk is blameless than a fool whose lips are perverse.
PROV|19|2|It is not good to have zeal without knowledge, nor to be hasty and miss the way.
PROV|19|3|A man's own folly ruins his life, yet his heart rages against the LORD.
PROV|19|4|Wealth brings many friends, but a poor man's friend deserts him.
PROV|19|5|A false witness will not go unpunished, and he who pours out lies will not go free.
PROV|19|6|Many curry favor with a ruler, and everyone is the friend of a man who gives gifts.
PROV|19|7|A poor man is shunned by all his relatives- how much more do his friends avoid him! Though he pursues them with pleading, they are nowhere to be found.
PROV|19|8|He who gets wisdom loves his own soul; he who cherishes understanding prospers.
PROV|19|9|A false witness will not go unpunished, and he who pours out lies will perish.
PROV|19|10|It is not fitting for a fool to live in luxury- how much worse for a slave to rule over princes!
PROV|19|11|A man's wisdom gives him patience; it is to his glory to overlook an offense.
PROV|19|12|A king's rage is like the roar of a lion, but his favor is like dew on the grass.
PROV|19|13|A foolish son is his father's ruin, and a quarrelsome wife is like a constant dripping.
PROV|19|14|Houses and wealth are inherited from parents, but a prudent wife is from the LORD.
PROV|19|15|Laziness brings on deep sleep, and the shiftless man goes hungry.
PROV|19|16|He who obeys instructions guards his life, but he who is contemptuous of his ways will die.
PROV|19|17|He who is kind to the poor lends to the LORD, and he will reward him for what he has done.
PROV|19|18|Discipline your son, for in that there is hope; do not be a willing party to his death.
PROV|19|19|A hot-tempered man must pay the penalty; if you rescue him, you will have to do it again.
PROV|19|20|Listen to advice and accept instruction, and in the end you will be wise.
PROV|19|21|Many are the plans in a man's heart, but it is the LORD's purpose that prevails.
PROV|19|22|What a man desires is unfailing love; better to be poor than a liar.
PROV|19|23|The fear of the LORD leads to life: Then one rests content, untouched by trouble.
PROV|19|24|The sluggard buries his hand in the dish; he will not even bring it back to his mouth!
PROV|19|25|Flog a mocker, and the simple will learn prudence; rebuke a discerning man, and he will gain knowledge.
PROV|19|26|He who robs his father and drives out his mother is a son who brings shame and disgrace.
PROV|19|27|Stop listening to instruction, my son, and you will stray from the words of knowledge.
PROV|19|28|A corrupt witness mocks at justice, and the mouth of the wicked gulps down evil.
PROV|19|29|Penalties are prepared for mockers, and beatings for the backs of fools.
PROV|20|1|Wine is a mocker and beer a brawler; whoever is led astray by them is not wise.
PROV|20|2|A king's wrath is like the roar of a lion; he who angers him forfeits his life.
PROV|20|3|It is to a man's honor to avoid strife, but every fool is quick to quarrel.
PROV|20|4|A sluggard does not plow in season; so at harvest time he looks but finds nothing.
PROV|20|5|The purposes of a man's heart are deep waters, but a man of understanding draws them out.
PROV|20|6|Many a man claims to have unfailing love, but a faithful man who can find?
PROV|20|7|The righteous man leads a blameless life; blessed are his children after him.
PROV|20|8|When a king sits on his throne to judge, he winnows out all evil with his eyes.
PROV|20|9|Who can say, "I have kept my heart pure; I am clean and without sin"?
PROV|20|10|Differing weights and differing measures- the LORD detests them both.
PROV|20|11|Even a child is known by his actions, by whether his conduct is pure and right.
PROV|20|12|Ears that hear and eyes that see- the LORD has made them both.
PROV|20|13|Do not love sleep or you will grow poor; stay awake and you will have food to spare.
PROV|20|14|"It's no good, it's no good!" says the buyer; then off he goes and boasts about his purchase.
PROV|20|15|Gold there is, and rubies in abundance, but lips that speak knowledge are a rare jewel.
PROV|20|16|Take the garment of one who puts up security for a stranger; hold it in pledge if he does it for a wayward woman.
PROV|20|17|Food gained by fraud tastes sweet to a man, but he ends up with a mouth full of gravel.
PROV|20|18|Make plans by seeking advice; if you wage war, obtain guidance.
PROV|20|19|A gossip betrays a confidence; so avoid a man who talks too much.
PROV|20|20|If a man curses his father or mother, his lamp will be snuffed out in pitch darkness.
PROV|20|21|An inheritance quickly gained at the beginning will not be blessed at the end.
PROV|20|22|Do not say, "I'll pay you back for this wrong!" Wait for the LORD, and he will deliver you.
PROV|20|23|The LORD detests differing weights, and dishonest scales do not please him.
PROV|20|24|A man's steps are directed by the LORD. How then can anyone understand his own way?
PROV|20|25|It is a trap for a man to dedicate something rashly and only later to consider his vows.
PROV|20|26|A wise king winnows out the wicked; he drives the threshing wheel over them.
PROV|20|27|The lamp of the LORD searches the spirit of a man; it searches out his inmost being.
PROV|20|28|Love and faithfulness keep a king safe; through love his throne is made secure.
PROV|20|29|The glory of young men is their strength, gray hair the splendor of the old.
PROV|20|30|Blows and wounds cleanse away evil, and beatings purge the inmost being.
PROV|21|1|The king's heart is in the hand of the LORD; he directs it like a watercourse wherever he pleases.
PROV|21|2|All a man's ways seem right to him, but the LORD weighs the heart.
PROV|21|3|To do what is right and just is more acceptable to the LORD than sacrifice.
PROV|21|4|Haughty eyes and a proud heart, the lamp of the wicked, are sin!
PROV|21|5|The plans of the diligent lead to profit as surely as haste leads to poverty.
PROV|21|6|A fortune made by a lying tongue is a fleeting vapor and a deadly snare.
PROV|21|7|The violence of the wicked will drag them away, for they refuse to do what is right.
PROV|21|8|The way of the guilty is devious, but the conduct of the innocent is upright.
PROV|21|9|Better to live on a corner of the roof than share a house with a quarrelsome wife.
PROV|21|10|The wicked man craves evil; his neighbor gets no mercy from him.
PROV|21|11|When a mocker is punished, the simple gain wisdom; when a wise man is instructed, he gets knowledge.
PROV|21|12|The Righteous One takes note of the house of the wicked and brings the wicked to ruin.
PROV|21|13|If a man shuts his ears to the cry of the poor, he too will cry out and not be answered.
PROV|21|14|A gift given in secret soothes anger, and a bribe concealed in the cloak pacifies great wrath.
PROV|21|15|When justice is done, it brings joy to the righteous but terror to evildoers.
PROV|21|16|A man who strays from the path of understanding comes to rest in the company of the dead.
PROV|21|17|He who loves pleasure will become poor; whoever loves wine and oil will never be rich.
PROV|21|18|The wicked become a ransom for the righteous, and the unfaithful for the upright.
PROV|21|19|Better to live in a desert than with a quarrelsome and ill-tempered wife.
PROV|21|20|In the house of the wise are stores of choice food and oil, but a foolish man devours all he has.
PROV|21|21|He who pursues righteousness and love finds life, prosperity and honor.
PROV|21|22|A wise man attacks the city of the mighty and pulls down the stronghold in which they trust.
PROV|21|23|He who guards his mouth and his tongue keeps himself from calamity.
PROV|21|24|The proud and arrogant man-"Mocker" is his name; he behaves with overweening pride.
PROV|21|25|The sluggard's craving will be the death of him, because his hands refuse to work.
PROV|21|26|All day long he craves for more, but the righteous give without sparing.
PROV|21|27|The sacrifice of the wicked is detestable- how much more so when brought with evil intent!
PROV|21|28|A false witness will perish, and whoever listens to him will be destroyed forever.
PROV|21|29|A wicked man puts up a bold front, but an upright man gives thought to his ways.
PROV|21|30|There is no wisdom, no insight, no plan that can succeed against the LORD.
PROV|21|31|The horse is made ready for the day of battle, but victory rests with the LORD.
PROV|22|1|A good name is more desirable than great riches; to be esteemed is better than silver or gold.
PROV|22|2|Rich and poor have this in common: The LORD is the Maker of them all.
PROV|22|3|A prudent man sees danger and takes refuge, but the simple keep going and suffer for it.
PROV|22|4|Humility and the fear of the LORD bring wealth and honor and life.
PROV|22|5|In the paths of the wicked lie thorns and snares, but he who guards his soul stays far from them.
PROV|22|6|Train a child in the way he should go, and when he is old he will not turn from it.
PROV|22|7|The rich rule over the poor, and the borrower is servant to the lender.
PROV|22|8|He who sows wickedness reaps trouble, and the rod of his fury will be destroyed.
PROV|22|9|A generous man will himself be blessed, for he shares his food with the poor.
PROV|22|10|Drive out the mocker, and out goes strife; quarrels and insults are ended.
PROV|22|11|He who loves a pure heart and whose speech is gracious will have the king for his friend.
PROV|22|12|The eyes of the LORD keep watch over knowledge, but he frustrates the words of the unfaithful.
PROV|22|13|The sluggard says, "There is a lion outside!" or, "I will be murdered in the streets!"
PROV|22|14|The mouth of an adulteress is a deep pit; he who is under the LORD's wrath will fall into it.
PROV|22|15|Folly is bound up in the heart of a child, but the rod of discipline will drive it far from him.
PROV|22|16|He who oppresses the poor to increase his wealth and he who gives gifts to the rich-both come to poverty.
PROV|22|17|Pay attention and listen to the sayings of the wise; apply your heart to what I teach,
PROV|22|18|for it is pleasing when you keep them in your heart and have all of them ready on your lips.
PROV|22|19|So that your trust may be in the LORD, I teach you today, even you.
PROV|22|20|Have I not written thirty sayings for you, sayings of counsel and knowledge,
PROV|22|21|teaching you true and reliable words, so that you can give sound answers to him who sent you?
PROV|22|22|Do not exploit the poor because they are poor and do not crush the needy in court,
PROV|22|23|for the LORD will take up their case and will plunder those who plunder them.
PROV|22|24|Do not make friends with a hot-tempered man, do not associate with one easily angered,
PROV|22|25|or you may learn his ways and get yourself ensnared.
PROV|22|26|Do not be a man who strikes hands in pledge or puts up security for debts;
PROV|22|27|if you lack the means to pay, your very bed will be snatched from under you.
PROV|22|28|Do not move an ancient boundary stone set up by your forefathers.
PROV|22|29|Do you see a man skilled in his work? He will serve before kings; he will not serve before obscure men.
PROV|23|1|When you sit to dine with a ruler, note well what is before you,
PROV|23|2|and put a knife to your throat if you are given to gluttony.
PROV|23|3|Do not crave his delicacies, for that food is deceptive.
PROV|23|4|Do not wear yourself out to get rich; have the wisdom to show restraint.
PROV|23|5|Cast but a glance at riches, and they are gone, for they will surely sprout wings and fly off to the sky like an eagle.
PROV|23|6|Do not eat the food of a stingy man, do not crave his delicacies;
PROV|23|7|for he is the kind of man who is always thinking about the cost. "Eat and drink," he says to you, but his heart is not with you.
PROV|23|8|You will vomit up the little you have eaten and will have wasted your compliments.
PROV|23|9|Do not speak to a fool, for he will scorn the wisdom of your words.
PROV|23|10|Do not move an ancient boundary stone or encroach on the fields of the fatherless,
PROV|23|11|for their Defender is strong; he will take up their case against you.
PROV|23|12|Apply your heart to instruction and your ears to words of knowledge.
PROV|23|13|Do not withhold discipline from a child; if you punish him with the rod, he will not die.
PROV|23|14|Punish him with the rod and save his soul from death.
PROV|23|15|My son, if your heart is wise, then my heart will be glad;
PROV|23|16|my inmost being will rejoice when your lips speak what is right.
PROV|23|17|Do not let your heart envy sinners, but always be zealous for the fear of the LORD.
PROV|23|18|There is surely a future hope for you, and your hope will not be cut off.
PROV|23|19|Listen, my son, and be wise, and keep your heart on the right path.
PROV|23|20|Do not join those who drink too much wine or gorge themselves on meat,
PROV|23|21|for drunkards and gluttons become poor, and drowsiness clothes them in rags.
PROV|23|22|Listen to your father, who gave you life, and do not despise your mother when she is old.
PROV|23|23|Buy the truth and do not sell it; get wisdom, discipline and understanding.
PROV|23|24|The father of a righteous man has great joy; he who has a wise son delights in him.
PROV|23|25|May your father and mother be glad; may she who gave you birth rejoice!
PROV|23|26|My son, give me your heart and let your eyes keep to my ways,
PROV|23|27|for a prostitute is a deep pit and a wayward wife is a narrow well.
PROV|23|28|Like a bandit she lies in wait, and multiplies the unfaithful among men.
PROV|23|29|Who has woe? Who has sorrow? Who has strife? Who has complaints? Who has needless bruises? Who has bloodshot eyes?
PROV|23|30|Those who linger over wine, who go to sample bowls of mixed wine.
PROV|23|31|Do not gaze at wine when it is red, when it sparkles in the cup, when it goes down smoothly!
PROV|23|32|In the end it bites like a snake and poisons like a viper.
PROV|23|33|Your eyes will see strange sights and your mind imagine confusing things.
PROV|23|34|You will be like one sleeping on the high seas, lying on top of the rigging.
PROV|23|35|"They hit me," you will say, "but I'm not hurt! They beat me, but I don't feel it! When will I wake up so I can find another drink?"
PROV|24|1|Do not envy wicked men, do not desire their company;
PROV|24|2|for their hearts plot violence, and their lips talk about making trouble.
PROV|24|3|By wisdom a house is built, and through understanding it is established;
PROV|24|4|through knowledge its rooms are filled with rare and beautiful treasures.
PROV|24|5|A wise man has great power, and a man of knowledge increases strength;
PROV|24|6|for waging war you need guidance, and for victory many advisers.
PROV|24|7|Wisdom is too high for a fool; in the assembly at the gate he has nothing to say.
PROV|24|8|He who plots evil will be known as a schemer.
PROV|24|9|The schemes of folly are sin, and men detest a mocker.
PROV|24|10|If you falter in times of trouble, how small is your strength!
PROV|24|11|Rescue those being led away to death; hold back those staggering toward slaughter.
PROV|24|12|If you say, "But we knew nothing about this," does not he who weighs the heart perceive it? Does not he who guards your life know it? Will he not repay each person according to what he has done?
PROV|24|13|Eat honey, my son, for it is good; honey from the comb is sweet to your taste.
PROV|24|14|Know also that wisdom is sweet to your soul; if you find it, there is a future hope for you, and your hope will not be cut off.
PROV|24|15|Do not lie in wait like an outlaw against a righteous man's house, do not raid his dwelling place;
PROV|24|16|for though a righteous man falls seven times, he rises again, but the wicked are brought down by calamity.
PROV|24|17|Do not gloat when your enemy falls; when he stumbles, do not let your heart rejoice,
PROV|24|18|or the LORD will see and disapprove and turn his wrath away from him.
PROV|24|19|Do not fret because of evil men or be envious of the wicked,
PROV|24|20|for the evil man has no future hope, and the lamp of the wicked will be snuffed out.
PROV|24|21|Fear the LORD and the king, my son, and do not join with the rebellious,
PROV|24|22|for those two will send sudden destruction upon them, and who knows what calamities they can bring? Further Sayings of the Wise
PROV|24|23|These also are sayings of the wise: To show partiality in judging is not good:
PROV|24|24|Whoever says to the guilty, "You are innocent"- peoples will curse him and nations denounce him.
PROV|24|25|But it will go well with those who convict the guilty, and rich blessing will come upon them.
PROV|24|26|An honest answer is like a kiss on the lips.
PROV|24|27|Finish your outdoor work and get your fields ready; after that, build your house.
PROV|24|28|Do not testify against your neighbor without cause, or use your lips to deceive.
PROV|24|29|Do not say, "I'll do to him as he has done to me; I'll pay that man back for what he did."
PROV|24|30|I went past the field of the sluggard, past the vineyard of the man who lacks judgment;
PROV|24|31|thorns had come up everywhere, the ground was covered with weeds, and the stone wall was in ruins.
PROV|24|32|I applied my heart to what I observed and learned a lesson from what I saw:
PROV|24|33|A little sleep, a little slumber, a little folding of the hands to rest-
PROV|24|34|and poverty will come on you like a bandit and scarcity like an armed man.
PROV|25|1|These are more proverbs of Solomon, copied by the men of Hezekiah king of Judah:
PROV|25|2|It is the glory of God to conceal a matter; to search out a matter is the glory of kings.
PROV|25|3|As the heavens are high and the earth is deep, so the hearts of kings are unsearchable.
PROV|25|4|Remove the dross from the silver, and out comes material for the silversmith;
PROV|25|5|remove the wicked from the king's presence, and his throne will be established through righteousness.
PROV|25|6|Do not exalt yourself in the king's presence, and do not claim a place among great men;
PROV|25|7|it is better for him to say to you, "Come up here," than for him to humiliate you before a nobleman. What you have seen with your eyes
PROV|25|8|do not bring hastily to court, for what will you do in the end if your neighbor puts you to shame?
PROV|25|9|If you argue your case with a neighbor, do not betray another man's confidence,
PROV|25|10|or he who hears it may shame you and you will never lose your bad reputation.
PROV|25|11|A word aptly spoken is like apples of gold in settings of silver.
PROV|25|12|Like an earring of gold or an ornament of fine gold is a wise man's rebuke to a listening ear.
PROV|25|13|Like the coolness of snow at harvest time is a trustworthy messenger to those who send him; he refreshes the spirit of his masters.
PROV|25|14|Like clouds and wind without rain is a man who boasts of gifts he does not give.
PROV|25|15|Through patience a ruler can be persuaded, and a gentle tongue can break a bone.
PROV|25|16|If you find honey, eat just enough- too much of it, and you will vomit.
PROV|25|17|Seldom set foot in your neighbor's house- too much of you, and he will hate you.
PROV|25|18|Like a club or a sword or a sharp arrow is the man who gives false testimony against his neighbor.
PROV|25|19|Like a bad tooth or a lame foot is reliance on the unfaithful in times of trouble.
PROV|25|20|Like one who takes away a garment on a cold day, or like vinegar poured on soda, is one who sings songs to a heavy heart.
PROV|25|21|If your enemy is hungry, give him food to eat; if he is thirsty, give him water to drink.
PROV|25|22|In doing this, you will heap burning coals on his head, and the LORD will reward you.
PROV|25|23|As a north wind brings rain, so a sly tongue brings angry looks.
PROV|25|24|Better to live on a corner of the roof than share a house with a quarrelsome wife.
PROV|25|25|Like cold water to a weary soul is good news from a distant land.
PROV|25|26|Like a muddied spring or a polluted well is a righteous man who gives way to the wicked.
PROV|25|27|It is not good to eat too much honey, nor is it honorable to seek one's own honor.
PROV|25|28|Like a city whose walls are broken down is a man who lacks self-control.
PROV|26|1|Like snow in summer or rain in harvest, honor is not fitting for a fool.
PROV|26|2|Like a fluttering sparrow or a darting swallow, an undeserved curse does not come to rest.
PROV|26|3|A whip for the horse, a halter for the donkey, and a rod for the backs of fools!
PROV|26|4|Do not answer a fool according to his folly, or you will be like him yourself.
PROV|26|5|Answer a fool according to his folly, or he will be wise in his own eyes.
PROV|26|6|Like cutting off one's feet or drinking violence is the sending of a message by the hand of a fool.
PROV|26|7|Like a lame man's legs that hang limp is a proverb in the mouth of a fool.
PROV|26|8|Like tying a stone in a sling is the giving of honor to a fool.
PROV|26|9|Like a thornbush in a drunkard's hand is a proverb in the mouth of a fool.
PROV|26|10|Like an archer who wounds at random is he who hires a fool or any passer-by.
PROV|26|11|As a dog returns to its vomit, so a fool repeats his folly.
PROV|26|12|Do you see a man wise in his own eyes? There is more hope for a fool than for him.
PROV|26|13|The sluggard says, "There is a lion in the road, a fierce lion roaming the streets!"
PROV|26|14|As a door turns on its hinges, so a sluggard turns on his bed.
PROV|26|15|The sluggard buries his hand in the dish; he is too lazy to bring it back to his mouth.
PROV|26|16|The sluggard is wiser in his own eyes than seven men who answer discreetly.
PROV|26|17|Like one who seizes a dog by the ears is a passer-by who meddles in a quarrel not his own.
PROV|26|18|Like a madman shooting firebrands or deadly arrows
PROV|26|19|is a man who deceives his neighbor and says, "I was only joking!"
PROV|26|20|Without wood a fire goes out; without gossip a quarrel dies down.
PROV|26|21|As charcoal to embers and as wood to fire, so is a quarrelsome man for kindling strife.
PROV|26|22|The words of a gossip are like choice morsels; they go down to a man's inmost parts.
PROV|26|23|Like a coating of glaze over earthenware are fervent lips with an evil heart.
PROV|26|24|A malicious man disguises himself with his lips, but in his heart he harbors deceit.
PROV|26|25|Though his speech is charming, do not believe him, for seven abominations fill his heart.
PROV|26|26|His malice may be concealed by deception, but his wickedness will be exposed in the assembly.
PROV|26|27|If a man digs a pit, he will fall into it; if a man rolls a stone, it will roll back on him.
PROV|26|28|A lying tongue hates those it hurts, and a flattering mouth works ruin.
PROV|27|1|Do not boast about tomorrow, for you do not know what a day may bring forth.
PROV|27|2|Let another praise you, and not your own mouth; someone else, and not your own lips.
PROV|27|3|Stone is heavy and sand a burden, but provocation by a fool is heavier than both.
PROV|27|4|Anger is cruel and fury overwhelming, but who can stand before jealousy?
PROV|27|5|Better is open rebuke than hidden love.
PROV|27|6|Wounds from a friend can be trusted, but an enemy multiplies kisses.
PROV|27|7|He who is full loathes honey, but to the hungry even what is bitter tastes sweet.
PROV|27|8|Like a bird that strays from its nest is a man who strays from his home.
PROV|27|9|Perfume and incense bring joy to the heart, and the pleasantness of one's friend springs from his earnest counsel.
PROV|27|10|Do not forsake your friend and the friend of your father, and do not go to your brother's house when disaster strikes you- better a neighbor nearby than a brother far away.
PROV|27|11|Be wise, my son, and bring joy to my heart; then I can answer anyone who treats me with contempt.
PROV|27|12|The prudent see danger and take refuge, but the simple keep going and suffer for it.
PROV|27|13|Take the garment of one who puts up security for a stranger; hold it in pledge if he does it for a wayward woman.
PROV|27|14|If a man loudly blesses his neighbor early in the morning, it will be taken as a curse.
PROV|27|15|A quarrelsome wife is like a constant dripping on a rainy day;
PROV|27|16|restraining her is like restraining the wind or grasping oil with the hand.
PROV|27|17|As iron sharpens iron, so one man sharpens another.
PROV|27|18|He who tends a fig tree will eat its fruit, and he who looks after his master will be honored.
PROV|27|19|As water reflects a face, so a man's heart reflects the man.
PROV|27|20|Death and Destruction are never satisfied, and neither are the eyes of man.
PROV|27|21|The crucible for silver and the furnace for gold, but man is tested by the praise he receives.
PROV|27|22|Though you grind a fool in a mortar, grinding him like grain with a pestle, you will not remove his folly from him.
PROV|27|23|Be sure you know the condition of your flocks, give careful attention to your herds;
PROV|27|24|for riches do not endure forever, and a crown is not secure for all generations.
PROV|27|25|When the hay is removed and new growth appears and the grass from the hills is gathered in,
PROV|27|26|the lambs will provide you with clothing, and the goats with the price of a field.
PROV|27|27|You will have plenty of goats' milk to feed you and your family and to nourish your servant girls.
PROV|28|1|The wicked man flees though no one pursues, but the righteous are as bold as a lion.
PROV|28|2|When a country is rebellious, it has many rulers, but a man of understanding and knowledge maintains order.
PROV|28|3|A ruler who oppresses the poor is like a driving rain that leaves no crops.
PROV|28|4|Those who forsake the law praise the wicked, but those who keep the law resist them.
PROV|28|5|Evil men do not understand justice, but those who seek the LORD understand it fully.
PROV|28|6|Better a poor man whose walk is blameless than a rich man whose ways are perverse.
PROV|28|7|He who keeps the law is a discerning son, but a companion of gluttons disgraces his father.
PROV|28|8|He who increases his wealth by exorbitant interest amasses it for another, who will be kind to the poor.
PROV|28|9|If anyone turns a deaf ear to the law, even his prayers are detestable.
PROV|28|10|He who leads the upright along an evil path will fall into his own trap, but the blameless will receive a good inheritance.
PROV|28|11|A rich man may be wise in his own eyes, but a poor man who has discernment sees through him.
PROV|28|12|When the righteous triumph, there is great elation; but when the wicked rise to power, men go into hiding.
PROV|28|13|He who conceals his sins does not prosper, but whoever confesses and renounces them finds mercy.
PROV|28|14|Blessed is the man who always fears the LORD, but he who hardens his heart falls into trouble.
PROV|28|15|Like a roaring lion or a charging bear is a wicked man ruling over a helpless people.
PROV|28|16|A tyrannical ruler lacks judgment, but he who hates ill-gotten gain will enjoy a long life.
PROV|28|17|A man tormented by the guilt of murder will be a fugitive till death; let no one support him.
PROV|28|18|He whose walk is blameless is kept safe, but he whose ways are perverse will suddenly fall.
PROV|28|19|He who works his land will have abundant food, but the one who chases fantasies will have his fill of poverty.
PROV|28|20|A faithful man will be richly blessed, but one eager to get rich will not go unpunished.
PROV|28|21|To show partiality is not good- yet a man will do wrong for a piece of bread.
PROV|28|22|A stingy man is eager to get rich and is unaware that poverty awaits him.
PROV|28|23|He who rebukes a man will in the end gain more favor than he who has a flattering tongue.
PROV|28|24|He who robs his father or mother and says, "It's not wrong"- he is partner to him who destroys.
PROV|28|25|A greedy man stirs up dissension, but he who trusts in the LORD will prosper.
PROV|28|26|He who trusts in himself is a fool, but he who walks in wisdom is kept safe.
PROV|28|27|He who gives to the poor will lack nothing, but he who closes his eyes to them receives many curses.
PROV|28|28|When the wicked rise to power, people go into hiding; but when the wicked perish, the righteous thrive.
PROV|29|1|A man who remains stiff-necked after many rebukes will suddenly be destroyed-without remedy.
PROV|29|2|When the righteous thrive, the people rejoice; when the wicked rule, the people groan.
PROV|29|3|A man who loves wisdom brings joy to his father, but a companion of prostitutes squanders his wealth.
PROV|29|4|By justice a king gives a country stability, but one who is greedy for bribes tears it down.
PROV|29|5|Whoever flatters his neighbor is spreading a net for his feet.
PROV|29|6|An evil man is snared by his own sin, but a righteous one can sing and be glad.
PROV|29|7|The righteous care about justice for the poor, but the wicked have no such concern.
PROV|29|8|Mockers stir up a city, but wise men turn away anger.
PROV|29|9|If a wise man goes to court with a fool, the fool rages and scoffs, and there is no peace.
PROV|29|10|Bloodthirsty men hate a man of integrity and seek to kill the upright.
PROV|29|11|A fool gives full vent to his anger, but a wise man keeps himself under control.
PROV|29|12|If a ruler listens to lies, all his officials become wicked.
PROV|29|13|The poor man and the oppressor have this in common: The LORD gives sight to the eyes of both.
PROV|29|14|If a king judges the poor with fairness, his throne will always be secure.
PROV|29|15|The rod of correction imparts wisdom, but a child left to himself disgraces his mother.
PROV|29|16|When the wicked thrive, so does sin, but the righteous will see their downfall.
PROV|29|17|Discipline your son, and he will give you peace; he will bring delight to your soul.
PROV|29|18|Where there is no revelation, the people cast off restraint; but blessed is he who keeps the law.
PROV|29|19|A servant cannot be corrected by mere words; though he understands, he will not respond.
PROV|29|20|Do you see a man who speaks in haste? There is more hope for a fool than for him.
PROV|29|21|If a man pampers his servant from youth, he will bring grief in the end.
PROV|29|22|An angry man stirs up dissension, and a hot-tempered one commits many sins.
PROV|29|23|A man's pride brings him low, but a man of lowly spirit gains honor.
PROV|29|24|The accomplice of a thief is his own enemy; he is put under oath and dare not testify.
PROV|29|25|Fear of man will prove to be a snare, but whoever trusts in the LORD is kept safe.
PROV|29|26|Many seek an audience with a ruler, but it is from the LORD that man gets justice.
PROV|29|27|The righteous detest the dishonest; the wicked detest the upright.
PROV|30|1|The sayings of Agur son of Jakeh-an oracle: This man declared to Ithiel, to Ithiel and to Ucal:
PROV|30|2|"I am the most ignorant of men; I do not have a man's understanding.
PROV|30|3|I have not learned wisdom, nor have I knowledge of the Holy One.
PROV|30|4|Who has gone up to heaven and come down? Who has gathered up the wind in the hollow of his hands? Who has wrapped up the waters in his cloak? Who has established all the ends of the earth? What is his name, and the name of his son? Tell me if you know!
PROV|30|5|"Every word of God is flawless; he is a shield to those who take refuge in him.
PROV|30|6|Do not add to his words, or he will rebuke you and prove you a liar.
PROV|30|7|"Two things I ask of you, O LORD; do not refuse me before I die:
PROV|30|8|Keep falsehood and lies far from me; give me neither poverty nor riches, but give me only my daily bread.
PROV|30|9|Otherwise, I may have too much and disown you and say, 'Who is the LORD?' Or I may become poor and steal, and so dishonor the name of my God.
PROV|30|10|"Do not slander a servant to his master, or he will curse you, and you will pay for it.
PROV|30|11|"There are those who curse their fathers and do not bless their mothers;
PROV|30|12|those who are pure in their own eyes and yet are not cleansed of their filth;
PROV|30|13|those whose eyes are ever so haughty, whose glances are so disdainful;
PROV|30|14|those whose teeth are swords and whose jaws are set with knives to devour the poor from the earth, the needy from among mankind.
PROV|30|15|"The leech has two daughters. 'Give! Give!' they cry. "There are three things that are never satisfied, four that never say, 'Enough!':
PROV|30|16|the grave, the barren womb, land, which is never satisfied with water, and fire, which never says, 'Enough!'
PROV|30|17|"The eye that mocks a father, that scorns obedience to a mother, will be pecked out by the ravens of the valley, will be eaten by the vultures.
PROV|30|18|"There are three things that are too amazing for me, four that I do not understand:
PROV|30|19|the way of an eagle in the sky, the way of a snake on a rock, the way of a ship on the high seas, and the way of a man with a maiden.
PROV|30|20|"This is the way of an adulteress: She eats and wipes her mouth and says, 'I've done nothing wrong.'
PROV|30|21|"Under three things the earth trembles, under four it cannot bear up:
PROV|30|22|a servant who becomes king, a fool who is full of food,
PROV|30|23|an unloved woman who is married, and a maidservant who displaces her mistress.
PROV|30|24|"Four things on earth are small, yet they are extremely wise:
PROV|30|25|Ants are creatures of little strength, yet they store up their food in the summer;
PROV|30|26|coneys are creatures of little power, yet they make their home in the crags;
PROV|30|27|locusts have no king, yet they advance together in ranks;
PROV|30|28|a lizard can be caught with the hand, yet it is found in kings' palaces.
PROV|30|29|"There are three things that are stately in their stride, four that move with stately bearing:
PROV|30|30|a lion, mighty among beasts, who retreats before nothing;
PROV|30|31|a strutting rooster, a he-goat, and a king with his army around him.
PROV|30|32|"If you have played the fool and exalted yourself, or if you have planned evil, clap your hand over your mouth!
PROV|30|33|For as churning the milk produces butter, and as twisting the nose produces blood, so stirring up anger produces strife."
PROV|31|1|The sayings of King Lemuel-an oracle his mother taught him:
PROV|31|2|"O my son, O son of my womb, O son of my vows,
PROV|31|3|do not spend your strength on women, your vigor on those who ruin kings.
PROV|31|4|"It is not for kings, O Lemuel- not for kings to drink wine, not for rulers to crave beer,
PROV|31|5|lest they drink and forget what the law decrees, and deprive all the oppressed of their rights.
PROV|31|6|Give beer to those who are perishing, wine to those who are in anguish;
PROV|31|7|let them drink and forget their poverty and remember their misery no more.
PROV|31|8|"Speak up for those who cannot speak for themselves, for the rights of all who are destitute.
PROV|31|9|Speak up and judge fairly; defend the rights of the poor and needy." Epilogue: The Wife of Noble Character
PROV|31|10|A wife of noble character who can find? She is worth far more than rubies.
PROV|31|11|Her husband has full confidence in her and lacks nothing of value.
PROV|31|12|She brings him good, not harm, all the days of her life.
PROV|31|13|She selects wool and flax and works with eager hands.
PROV|31|14|She is like the merchant ships, bringing her food from afar.
PROV|31|15|She gets up while it is still dark; she provides food for her family and portions for her servant girls.
PROV|31|16|She considers a field and buys it; out of her earnings she plants a vineyard.
PROV|31|17|She sets about her work vigorously; her arms are strong for her tasks.
PROV|31|18|She sees that her trading is profitable, and her lamp does not go out at night.
PROV|31|19|In her hand she holds the distaff and grasps the spindle with her fingers.
PROV|31|20|She opens her arms to the poor and extends her hands to the needy.
PROV|31|21|When it snows, she has no fear for her household; for all of them are clothed in scarlet.
PROV|31|22|She makes coverings for her bed; she is clothed in fine linen and purple.
PROV|31|23|Her husband is respected at the city gate, where he takes his seat among the elders of the land.
PROV|31|24|She makes linen garments and sells them, and supplies the merchants with sashes.
PROV|31|25|She is clothed with strength and dignity; she can laugh at the days to come.
PROV|31|26|She speaks with wisdom, and faithful instruction is on her tongue.
PROV|31|27|She watches over the affairs of her household and does not eat the bread of idleness.
PROV|31|28|Her children arise and call her blessed; her husband also, and he praises her:
PROV|31|29|"Many women do noble things, but you surpass them all."
PROV|31|30|Charm is deceptive, and beauty is fleeting; but a woman who fears the LORD is to be praised.
PROV|31|31|Give her the reward she has earned, and let her works bring her praise at the city gate.
