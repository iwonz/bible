JOB|1|1|There was a man in the land of Uz, whose name was Job; and that man was perfect and upright, and one that feared God, and eschewed evil.
JOB|1|2|And there were born unto him seven sons and three daughters.
JOB|1|3|His substance also was seven thousand sheep, and three thousand camels, and five hundred yoke of oxen, and five hundred she asses, and a very great household; so that this man was the greatest of all the men of the east.
JOB|1|4|And his sons went and feasted in their houses, every one his day; and sent and called for their three sisters to eat and to drink with them.
JOB|1|5|And it was so, when the days of their feasting were gone about, that Job sent and sanctified them, and rose up early in the morning, and offered burnt offerings according to the number of them all: for Job said, It may be that my sons have sinned, and cursed God in their hearts. Thus did Job continually.
JOB|1|6|Now there was a day when the sons of God came to present themselves before the LORD, and Satan came also among them.
JOB|1|7|And the LORD said unto Satan, Whence comest thou? Then Satan answered the LORD, and said, From going to and fro in the earth, and from walking up and down in it.
JOB|1|8|And the LORD said unto Satan, Hast thou considered my servant Job, that there is none like him in the earth, a perfect and an upright man, one that feareth God, and escheweth evil?
JOB|1|9|Then Satan answered the LORD, and said, Doth Job fear God for nought?
JOB|1|10|Hast not thou made an hedge about him, and about his house, and about all that he hath on every side? thou hast blessed the work of his hands, and his substance is increased in the land.
JOB|1|11|But put forth thine hand now, and touch all that he hath, and he will curse thee to thy face.
JOB|1|12|And the LORD said unto Satan, Behold, all that he hath is in thy power; only upon himself put not forth thine hand. So Satan went forth from the presence of the LORD.
JOB|1|13|And there was a day when his sons and his daughters were eating and drinking wine in their eldest brother's house:
JOB|1|14|And there came a messenger unto Job, and said, The oxen were plowing, and the asses feeding beside them:
JOB|1|15|And the Sabeans fell upon them, and took them away; yea, they have slain the servants with the edge of the sword; and I only am escaped alone to tell thee.
JOB|1|16|While he was yet speaking, there came also another, and said, The fire of God is fallen from heaven, and hath burned up the sheep, and the servants, and consumed them; and I only am escaped alone to tell thee.
JOB|1|17|While he was yet speaking, there came also another, and said, The Chaldeans made out three bands, and fell upon the camels, and have carried them away, yea, and slain the servants with the edge of the sword; and I only am escaped alone to tell thee.
JOB|1|18|While he was yet speaking, there came also another, and said, Thy sons and thy daughters were eating and drinking wine in their eldest brother's house:
JOB|1|19|And, behold, there came a great wind from the wilderness, and smote the four corners of the house, and it fell upon the young men, and they are dead; and I only am escaped alone to tell thee.
JOB|1|20|Then Job arose, and rent his mantle, and shaved his head, and fell down upon the ground, and worshipped,
JOB|1|21|And said, Naked came I out of my mother's womb, and naked shall I return thither: the LORD gave, and the LORD hath taken away; blessed be the name of the LORD.
JOB|1|22|In all this Job sinned not, nor charged God foolishly.
JOB|2|1|Again there was a day when the sons of God came to present themselves before the LORD, and Satan came also among them to present himself before the LORD.
JOB|2|2|And the LORD said unto Satan, From whence comest thou? And Satan answered the LORD, and said, From going to and fro in the earth, and from walking up and down in it.
JOB|2|3|And the LORD said unto Satan, Hast thou considered my servant Job, that there is none like him in the earth, a perfect and an upright man, one that feareth God, and escheweth evil? and still he holdeth fast his integrity, although thou movedst me against him, to destroy him without cause.
JOB|2|4|And Satan answered the LORD, and said, Skin for skin, yea, all that a man hath will he give for his life.
JOB|2|5|But put forth thine hand now, and touch his bone and his flesh, and he will curse thee to thy face.
JOB|2|6|And the LORD said unto Satan, Behold, he is in thine hand; but save his life.
JOB|2|7|So went Satan forth from the presence of the LORD, and smote Job with sore boils from the sole of his foot unto his crown.
JOB|2|8|And he took him a potsherd to scrape himself withal; and he sat down among the ashes.
JOB|2|9|Then said his wife unto him, Dost thou still retain thine integrity? curse God, and die.
JOB|2|10|But he said unto her, Thou speakest as one of the foolish women speaketh. What? shall we receive good at the hand of God, and shall we not receive evil? In all this did not Job sin with his lips.
JOB|2|11|Now when Job's three friends heard of all this evil that was come upon him, they came every one from his own place; Eliphaz the Temanite, and Bildad the Shuhite, and Zophar the Naamathite: for they had made an appointment together to come to mourn with him and to comfort him.
JOB|2|12|And when they lifted up their eyes afar off, and knew him not, they lifted up their voice, and wept; and they rent every one his mantle, and sprinkled dust upon their heads toward heaven.
JOB|2|13|So they sat down with him upon the ground seven days and seven nights, and none spake a word unto him: for they saw that his grief was very great.
JOB|3|1|After this opened Job his mouth, and cursed his day.
JOB|3|2|And Job spake, and said,
JOB|3|3|Let the day perish wherein I was born, and the night in which it was said, There is a man child conceived.
JOB|3|4|Let that day be darkness; let not God regard it from above, neither let the light shine upon it.
JOB|3|5|Let darkness and the shadow of death stain it; let a cloud dwell upon it; let the blackness of the day terrify it.
JOB|3|6|As for that night, let darkness seize upon it; let it not be joined unto the days of the year, let it not come into the number of the months.
JOB|3|7|Lo, let that night be solitary, let no joyful voice come therein.
JOB|3|8|Let them curse it that curse the day, who are ready to raise up their mourning.
JOB|3|9|Let the stars of the twilight thereof be dark; let it look for light, but have none; neither let it see the dawning of the day:
JOB|3|10|Because it shut not up the doors of my mother's womb, nor hid sorrow from mine eyes.
JOB|3|11|Why died I not from the womb? why did I not give up the ghost when I came out of the belly?
JOB|3|12|Why did the knees prevent me? or why the breasts that I should suck?
JOB|3|13|For now should I have lain still and been quiet, I should have slept: then had I been at rest,
JOB|3|14|With kings and counsellors of the earth, which build desolate places for themselves;
JOB|3|15|Or with princes that had gold, who filled their houses with silver:
JOB|3|16|Or as an hidden untimely birth I had not been; as infants which never saw light.
JOB|3|17|There the wicked cease from troubling; and there the weary be at rest.
JOB|3|18|There the prisoners rest together; they hear not the voice of the oppressor.
JOB|3|19|The small and great are there; and the servant is free from his master.
JOB|3|20|Wherefore is light given to him that is in misery, and life unto the bitter in soul;
JOB|3|21|Which long for death, but it cometh not; and dig for it more than for hid treasures;
JOB|3|22|Which rejoice exceedingly, and are glad, when they can find the grave?
JOB|3|23|Why is light given to a man whose way is hid, and whom God hath hedged in?
JOB|3|24|For my sighing cometh before I eat, and my roarings are poured out like the waters.
JOB|3|25|For the thing which I greatly feared is come upon me, and that which I was afraid of is come unto me.
JOB|3|26|I was not in safety, neither had I rest, neither was I quiet; yet trouble came.
JOB|4|1|Then Eliphaz the Temanite answered and said,
JOB|4|2|If we assay to commune with thee, wilt thou be grieved? but who can withhold himself from speaking?
JOB|4|3|Behold, thou hast instructed many, and thou hast strengthened the weak hands.
JOB|4|4|Thy words have upholden him that was falling, and thou hast strengthened the feeble knees.
JOB|4|5|But now it is come upon thee, and thou faintest; it toucheth thee, and thou art troubled.
JOB|4|6|Is not this thy fear, thy confidence, thy hope, and the uprightness of thy ways?
JOB|4|7|Remember, I pray thee, who ever perished, being innocent? or where were the righteous cut off?
JOB|4|8|Even as I have seen, they that plow iniquity, and sow wickedness, reap the same.
JOB|4|9|By the blast of God they perish, and by the breath of his nostrils are they consumed.
JOB|4|10|The roaring of the lion, and the voice of the fierce lion, and the teeth of the young lions, are broken.
JOB|4|11|The old lion perisheth for lack of prey, and the stout lion's whelps are scattered abroad.
JOB|4|12|Now a thing was secretly brought to me, and mine ear received a little thereof.
JOB|4|13|In thoughts from the visions of the night, when deep sleep falleth on men,
JOB|4|14|Fear came upon me, and trembling, which made all my bones to shake.
JOB|4|15|Then a spirit passed before my face; the hair of my flesh stood up:
JOB|4|16|It stood still, but I could not discern the form thereof: an image was before mine eyes, there was silence, and I heard a voice, saying,
JOB|4|17|Shall mortal man be more just than God? shall a man be more pure than his maker?
JOB|4|18|Behold, he put no trust in his servants; and his angels he charged with folly:
JOB|4|19|How much less in them that dwell in houses of clay, whose foundation is in the dust, which are crushed before the moth?
JOB|4|20|They are destroyed from morning to evening: they perish for ever without any regarding it.
JOB|4|21|Doth not their excellency which is in them go away? they die, even without wisdom.
JOB|5|1|Call now, if there be any that will answer thee; and to which of the saints wilt thou turn?
JOB|5|2|For wrath killeth the foolish man, and envy slayeth the silly one.
JOB|5|3|I have seen the foolish taking root: but suddenly I cursed his habitation.
JOB|5|4|His children are far from safety, and they are crushed in the gate, neither is there any to deliver them.
JOB|5|5|Whose harvest the hungry eateth up, and taketh it even out of the thorns, and the robber swalloweth up their substance.
JOB|5|6|Although affliction cometh not forth of the dust, neither doth trouble spring out of the ground;
JOB|5|7|Yet man is born unto trouble, as the sparks fly upward.
JOB|5|8|I would seek unto God, and unto God would I commit my cause:
JOB|5|9|Which doeth great things and unsearchable; marvellous things without number:
JOB|5|10|Who giveth rain upon the earth, and sendeth waters upon the fields:
JOB|5|11|To set up on high those that be low; that those which mourn may be exalted to safety.
JOB|5|12|He disappointeth the devices of the crafty, so that their hands cannot perform their enterprise.
JOB|5|13|He taketh the wise in their own craftiness: and the counsel of the froward is carried headlong.
JOB|5|14|They meet with darkness in the day time, and grope in the noonday as in the night.
JOB|5|15|But he saveth the poor from the sword, from their mouth, and from the hand of the mighty.
JOB|5|16|So the poor hath hope, and iniquity stoppeth her mouth.
JOB|5|17|Behold, happy is the man whom God correcteth: therefore despise not thou the chastening of the Almighty:
JOB|5|18|For he maketh sore, and bindeth up: he woundeth, and his hands make whole.
JOB|5|19|He shall deliver thee in six troubles: yea, in seven there shall no evil touch thee.
JOB|5|20|In famine he shall redeem thee from death: and in war from the power of the sword.
JOB|5|21|Thou shalt be hid from the scourge of the tongue: neither shalt thou be afraid of destruction when it cometh.
JOB|5|22|At destruction and famine thou shalt laugh: neither shalt thou be afraid of the beasts of the earth.
JOB|5|23|For thou shalt be in league with the stones of the field: and the beasts of the field shall be at peace with thee.
JOB|5|24|And thou shalt know that thy tabernacle shall be in peace; and thou shalt visit thy habitation, and shalt not sin.
JOB|5|25|Thou shalt know also that thy seed shall be great, and thine offspring as the grass of the earth.
JOB|5|26|Thou shalt come to thy grave in a full age, like as a shock of corn cometh in in his season.
JOB|5|27|Lo this, we have searched it, so it is; hear it, and know thou it for thy good.
JOB|6|1|But Job answered and said,
JOB|6|2|Oh that my grief were throughly weighed, and my calamity laid in the balances together!
JOB|6|3|For now it would be heavier than the sand of the sea: therefore my words are swallowed up.
JOB|6|4|For the arrows of the Almighty are within me, the poison whereof drinketh up my spirit: the terrors of God do set themselves in array against me.
JOB|6|5|Doth the wild ass bray when he hath grass? or loweth the ox over his fodder?
JOB|6|6|Can that which is unsavoury be eaten without salt? or is there any taste in the white of an egg?
JOB|6|7|The things that my soul refused to touch are as my sorrowful meat.
JOB|6|8|Oh that I might have my request; and that God would grant me the thing that I long for!
JOB|6|9|Even that it would please God to destroy me; that he would let loose his hand, and cut me off!
JOB|6|10|Then should I yet have comfort; yea, I would harden myself in sorrow: let him not spare; for I have not concealed the words of the Holy One.
JOB|6|11|What is my strength, that I should hope? and what is mine end, that I should prolong my life?
JOB|6|12|Is my strength the strength of stones? or is my flesh of brass?
JOB|6|13|Is not my help in me? and is wisdom driven quite from me?
JOB|6|14|To him that is afflicted pity should be shewed from his friend; but he forsaketh the fear of the Almighty.
JOB|6|15|My brethren have dealt deceitfully as a brook, and as the stream of brooks they pass away;
JOB|6|16|Which are blackish by reason of the ice, and wherein the snow is hid:
JOB|6|17|What time they wax warm, they vanish: when it is hot, they are consumed out of their place.
JOB|6|18|The paths of their way are turned aside; they go to nothing, and perish.
JOB|6|19|The troops of Tema looked, the companies of Sheba waited for them.
JOB|6|20|They were confounded because they had hoped; they came thither, and were ashamed.
JOB|6|21|For now ye are nothing; ye see my casting down, and are afraid.
JOB|6|22|Did I say, Bring unto me? or, Give a reward for me of your substance?
JOB|6|23|Or, Deliver me from the enemy's hand? or, Redeem me from the hand of the mighty?
JOB|6|24|Teach me, and I will hold my tongue: and cause me to understand wherein I have erred.
JOB|6|25|How forcible are right words! but what doth your arguing reprove?
JOB|6|26|Do ye imagine to reprove words, and the speeches of one that is desperate, which are as wind?
JOB|6|27|Yea, ye overwhelm the fatherless, and ye dig a pit for your friend.
JOB|6|28|Now therefore be content, look upon me; for it is evident unto you if I lie.
JOB|6|29|Return, I pray you, let it not be iniquity; yea, return again, my righteousness is in it.
JOB|6|30|Is there iniquity in my tongue? cannot my taste discern perverse things?
JOB|7|1|Is there not an appointed time to man upon earth? are not his days also like the days of an hireling?
JOB|7|2|As a servant earnestly desireth the shadow, and as an hireling looketh for the reward of his work:
JOB|7|3|So am I made to possess months of vanity, and wearisome nights are appointed to me.
JOB|7|4|When I lie down, I say, When shall I arise, and the night be gone? and I am full of tossings to and fro unto the dawning of the day.
JOB|7|5|My flesh is clothed with worms and clods of dust; my skin is broken, and become loathsome.
JOB|7|6|My days are swifter than a weaver's shuttle, and are spent without hope.
JOB|7|7|O remember that my life is wind: mine eye shall no more see good.
JOB|7|8|The eye of him that hath seen me shall see me no more: thine eyes are upon me, and I am not.
JOB|7|9|As the cloud is consumed and vanisheth away: so he that goeth down to the grave shall come up no more.
JOB|7|10|He shall return no more to his house, neither shall his place know him any more.
JOB|7|11|Therefore I will not refrain my mouth; I will speak in the anguish of my spirit; I will complain in the bitterness of my soul.
JOB|7|12|Am I a sea, or a whale, that thou settest a watch over me?
JOB|7|13|When I say, My bed shall comfort me, my couch shall ease my complaints;
JOB|7|14|Then thou scarest me with dreams, and terrifiest me through visions:
JOB|7|15|So that my soul chooseth strangling, and death rather than my life.
JOB|7|16|I loathe it; I would not live alway: let me alone; for my days are vanity.
JOB|7|17|What is man, that thou shouldest magnify him? and that thou shouldest set thine heart upon him?
JOB|7|18|And that thou shouldest visit him every morning, and try him every moment?
JOB|7|19|How long wilt thou not depart from me, nor let me alone till I swallow down my spittle?
JOB|7|20|I have sinned; what shall I do unto thee, O thou preserver of men? why hast thou set me as a mark against thee, so that I am a burden to myself?
JOB|7|21|And why dost thou not pardon my transgression, and take away my iniquity? for now shall I sleep in the dust; and thou shalt seek me in the morning, but I shall not be.
JOB|8|1|Then answered Bildad the Shuhite, and said,
JOB|8|2|How long wilt thou speak these things? and how long shall the words of thy mouth be like a strong wind?
JOB|8|3|Doth God pervert judgment? or doth the Almighty pervert justice?
JOB|8|4|If thy children have sinned against him, and he have cast them away for their transgression;
JOB|8|5|If thou wouldest seek unto God betimes, and make thy supplication to the Almighty;
JOB|8|6|If thou wert pure and upright; surely now he would awake for thee, and make the habitation of thy righteousness prosperous.
JOB|8|7|Though thy beginning was small, yet thy latter end should greatly increase.
JOB|8|8|For enquire, I pray thee, of the former age, and prepare thyself to the search of their fathers:
JOB|8|9|(For we are but of yesterday, and know nothing, because our days upon earth are a shadow:)
JOB|8|10|Shall not they teach thee, and tell thee, and utter words out of their heart?
JOB|8|11|Can the rush grow up without mire? can the flag grow without water?
JOB|8|12|Whilst it is yet in his greenness, and not cut down, it withereth before any other herb.
JOB|8|13|So are the paths of all that forget God; and the hypocrite's hope shall perish:
JOB|8|14|Whose hope shall be cut off, and whose trust shall be a spider's web.
JOB|8|15|He shall lean upon his house, but it shall not stand: he shall hold it fast, but it shall not endure.
JOB|8|16|He is green before the sun, and his branch shooteth forth in his garden.
JOB|8|17|His roots are wrapped about the heap, and seeth the place of stones.
JOB|8|18|If he destroy him from his place, then it shall deny him, saying, I have not seen thee.
JOB|8|19|Behold, this is the joy of his way, and out of the earth shall others grow.
JOB|8|20|Behold, God will not cast away a perfect man, neither will he help the evil doers:
JOB|8|21|Till he fill thy mouth with laughing, and thy lips with rejoicing.
JOB|8|22|They that hate thee shall be clothed with shame; and the dwelling place of the wicked shall come to nought.
JOB|9|1|Then Job answered and said,
JOB|9|2|I know it is so of a truth: but how should man be just with God?
JOB|9|3|If he will contend with him, he cannot answer him one of a thousand.
JOB|9|4|He is wise in heart, and mighty in strength: who hath hardened himself against him, and hath prospered?
JOB|9|5|Which removeth the mountains, and they know not: which overturneth them in his anger.
JOB|9|6|Which shaketh the earth out of her place, and the pillars thereof tremble.
JOB|9|7|Which commandeth the sun, and it riseth not; and sealeth up the stars.
JOB|9|8|Which alone spreadeth out the heavens, and treadeth upon the waves of the sea.
JOB|9|9|Which maketh Arcturus, Orion, and Pleiades, and the chambers of the south.
JOB|9|10|Which doeth great things past finding out; yea, and wonders without number.
JOB|9|11|Lo, he goeth by me, and I see him not: he passeth on also, but I perceive him not.
JOB|9|12|Behold, he taketh away, who can hinder him? who will say unto him, What doest thou?
JOB|9|13|If God will not withdraw his anger, the proud helpers do stoop under him.
JOB|9|14|How much less shall I answer him, and choose out my words to reason with him?
JOB|9|15|Whom, though I were righteous, yet would I not answer, but I would make supplication to my judge.
JOB|9|16|If I had called, and he had answered me; yet would I not believe that he had hearkened unto my voice.
JOB|9|17|For he breaketh me with a tempest, and multiplieth my wounds without cause.
JOB|9|18|He will not suffer me to take my breath, but filleth me with bitterness.
JOB|9|19|If I speak of strength, lo, he is strong: and if of judgment, who shall set me a time to plead?
JOB|9|20|If I justify myself, mine own mouth shall condemn me: if I say, I am perfect, it shall also prove me perverse.
JOB|9|21|Though I were perfect, yet would I not know my soul: I would despise my life.
JOB|9|22|This is one thing, therefore I said it, He destroyeth the perfect and the wicked.
JOB|9|23|If the scourge slay suddenly, he will laugh at the trial of the innocent.
JOB|9|24|The earth is given into the hand of the wicked: he covereth the faces of the judges thereof; if not, where, and who is he?
JOB|9|25|Now my days are swifter than a post: they flee away, they see no good.
JOB|9|26|They are passed away as the swift ships: as the eagle that hasteth to the prey.
JOB|9|27|If I say, I will forget my complaint, I will leave off my heaviness, and comfort myself:
JOB|9|28|I am afraid of all my sorrows, I know that thou wilt not hold me innocent.
JOB|9|29|If I be wicked, why then labour I in vain?
JOB|9|30|If I wash myself with snow water, and make my hands never so clean;
JOB|9|31|Yet shalt thou plunge me in the ditch, and mine own clothes shall abhor me.
JOB|9|32|For he is not a man, as I am, that I should answer him, and we should come together in judgment.
JOB|9|33|Neither is there any daysman betwixt us, that might lay his hand upon us both.
JOB|9|34|Let him take his rod away from me, and let not his fear terrify me:
JOB|9|35|Then would I speak, and not fear him; but it is not so with me.
JOB|10|1|My soul is weary of my life; I will leave my complaint upon myself; I will speak in the bitterness of my soul.
JOB|10|2|I will say unto God, Do not condemn me; shew me wherefore thou contendest with me.
JOB|10|3|Is it good unto thee that thou shouldest oppress, that thou shouldest despise the work of thine hands, and shine upon the counsel of the wicked?
JOB|10|4|Hast thou eyes of flesh? or seest thou as man seeth?
JOB|10|5|Are thy days as the days of man? are thy years as man's days,
JOB|10|6|That thou enquirest after mine iniquity, and searchest after my sin?
JOB|10|7|Thou knowest that I am not wicked; and there is none that can deliver out of thine hand.
JOB|10|8|Thine hands have made me and fashioned me together round about; yet thou dost destroy me.
JOB|10|9|Remember, I beseech thee, that thou hast made me as the clay; and wilt thou bring me into dust again?
JOB|10|10|Hast thou not poured me out as milk, and curdled me like cheese?
JOB|10|11|Thou hast clothed me with skin and flesh, and hast fenced me with bones and sinews.
JOB|10|12|Thou hast granted me life and favour, and thy visitation hath preserved my spirit.
JOB|10|13|And these things hast thou hid in thine heart: I know that this is with thee.
JOB|10|14|If I sin, then thou markest me, and thou wilt not acquit me from mine iniquity.
JOB|10|15|If I be wicked, woe unto me; and if I be righteous, yet will I not lift up my head. I am full of confusion; therefore see thou mine affliction;
JOB|10|16|For it increaseth. Thou huntest me as a fierce lion: and again thou shewest thyself marvellous upon me.
JOB|10|17|Thou renewest thy witnesses against me, and increasest thine indignation upon me; changes and war are against me.
JOB|10|18|Wherefore then hast thou brought me forth out of the womb? Oh that I had given up the ghost, and no eye had seen me!
JOB|10|19|I should have been as though I had not been; I should have been carried from the womb to the grave.
JOB|10|20|Are not my days few? cease then, and let me alone, that I may take comfort a little,
JOB|10|21|Before I go whence I shall not return, even to the land of darkness and the shadow of death;
JOB|10|22|A land of darkness, as darkness itself; and of the shadow of death, without any order, and where the light is as darkness.
JOB|11|1|Then answered Zophar the Naamathite, and said,
JOB|11|2|Should not the multitude of words be answered? and should a man full of talk be justified?
JOB|11|3|Should thy lies make men hold their peace? and when thou mockest, shall no man make thee ashamed?
JOB|11|4|For thou hast said, My doctrine is pure, and I am clean in thine eyes.
JOB|11|5|But oh that God would speak, and open his lips against thee;
JOB|11|6|And that he would shew thee the secrets of wisdom, that they are double to that which is! Know therefore that God exacteth of thee less than thine iniquity deserveth.
JOB|11|7|Canst thou by searching find out God? canst thou find out the Almighty unto perfection?
JOB|11|8|It is as high as heaven; what canst thou do? deeper than hell; what canst thou know?
JOB|11|9|The measure thereof is longer than the earth, and broader than the sea.
JOB|11|10|If he cut off, and shut up, or gather together, then who can hinder him?
JOB|11|11|For he knoweth vain men: he seeth wickedness also; will he not then consider it?
JOB|11|12|For vain men would be wise, though man be born like a wild ass's colt.
JOB|11|13|If thou prepare thine heart, and stretch out thine hands toward him;
JOB|11|14|If iniquity be in thine hand, put it far away, and let not wickedness dwell in thy tabernacles.
JOB|11|15|For then shalt thou lift up thy face without spot; yea, thou shalt be stedfast, and shalt not fear:
JOB|11|16|Because thou shalt forget thy misery, and remember it as waters that pass away:
JOB|11|17|And thine age shall be clearer than the noonday: thou shalt shine forth, thou shalt be as the morning.
JOB|11|18|And thou shalt be secure, because there is hope; yea, thou shalt dig about thee, and thou shalt take thy rest in safety.
JOB|11|19|Also thou shalt lie down, and none shall make thee afraid; yea, many shall make suit unto thee.
JOB|11|20|But the eyes of the wicked shall fail, and they shall not escape, and their hope shall be as the giving up of the ghost.
JOB|12|1|And Job answered and said,
JOB|12|2|No doubt but ye are the people, and wisdom shall die with you.
JOB|12|3|But I have understanding as well as you; I am not inferior to you: yea, who knoweth not such things as these?
JOB|12|4|I am as one mocked of his neighbour, who calleth upon God, and he answereth him: the just upright man is laughed to scorn.
JOB|12|5|He that is ready to slip with his feet is as a lamp despised in the thought of him that is at ease.
JOB|12|6|The tabernacles of robbers prosper, and they that provoke God are secure; into whose hand God bringeth abundantly.
JOB|12|7|But ask now the beasts, and they shall teach thee; and the fowls of the air, and they shall tell thee:
JOB|12|8|Or speak to the earth, and it shall teach thee: and the fishes of the sea shall declare unto thee.
JOB|12|9|Who knoweth not in all these that the hand of the LORD hath wrought this?
JOB|12|10|In whose hand is the soul of every living thing, and the breath of all mankind.
JOB|12|11|Doth not the ear try words? and the mouth taste his meat?
JOB|12|12|With the ancient is wisdom; and in length of days understanding.
JOB|12|13|With him is wisdom and strength, he hath counsel and understanding.
JOB|12|14|Behold, he breaketh down, and it cannot be built again: he shutteth up a man, and there can be no opening.
JOB|12|15|Behold, he withholdeth the waters, and they dry up: also he sendeth them out, and they overturn the earth.
JOB|12|16|With him is strength and wisdom: the deceived and the deceiver are his.
JOB|12|17|He leadeth counsellors away spoiled, and maketh the judges fools.
JOB|12|18|He looseth the bond of kings, and girdeth their loins with a girdle.
JOB|12|19|He leadeth princes away spoiled, and overthroweth the mighty.
JOB|12|20|He removeth away the speech of the trusty, and taketh away the understanding of the aged.
JOB|12|21|He poureth contempt upon princes, and weakeneth the strength of the mighty.
JOB|12|22|He discovereth deep things out of darkness, and bringeth out to light the shadow of death.
JOB|12|23|He increaseth the nations, and destroyeth them: he enlargeth the nations, and straiteneth them again.
JOB|12|24|He taketh away the heart of the chief of the people of the earth, and causeth them to wander in a wilderness where there is no way.
JOB|12|25|They grope in the dark without light, and he maketh them to stagger like a drunken man.
JOB|13|1|Lo, mine eye hath seen all this, mine ear hath heard and understood it.
JOB|13|2|What ye know, the same do I know also: I am not inferior unto you.
JOB|13|3|Surely I would speak to the Almighty, and I desire to reason with God.
JOB|13|4|But ye are forgers of lies, ye are all physicians of no value.
JOB|13|5|O that ye would altogether hold your peace! and it should be your wisdom.
JOB|13|6|Hear now my reasoning, and hearken to the pleadings of my lips.
JOB|13|7|Will ye speak wickedly for God? and talk deceitfully for him?
JOB|13|8|Will ye accept his person? will ye contend for God?
JOB|13|9|Is it good that he should search you out? or as one man mocketh another, do ye so mock him?
JOB|13|10|He will surely reprove you, if ye do secretly accept persons.
JOB|13|11|Shall not his excellency make you afraid? and his dread fall upon you?
JOB|13|12|Your remembrances are like unto ashes, your bodies to bodies of clay.
JOB|13|13|Hold your peace, let me alone, that I may speak, and let come on me what will.
JOB|13|14|Wherefore do I take my flesh in my teeth, and put my life in mine hand?
JOB|13|15|Though he slay me, yet will I trust in him: but I will maintain mine own ways before him.
JOB|13|16|He also shall be my salvation: for an hypocrite shall not come before him.
JOB|13|17|Hear diligently my speech, and my declaration with your ears.
JOB|13|18|Behold now, I have ordered my cause; I know that I shall be justified.
JOB|13|19|Who is he that will plead with me? for now, if I hold my tongue, I shall give up the ghost.
JOB|13|20|Only do not two things unto me: then will I not hide myself from thee.
JOB|13|21|Withdraw thine hand far from me: and let not thy dread make me afraid.
JOB|13|22|Then call thou, and I will answer: or let me speak, and answer thou me.
JOB|13|23|How many are mine iniquities and sins? make me to know my transgression and my sin.
JOB|13|24|Wherefore hidest thou thy face, and holdest me for thine enemy?
JOB|13|25|Wilt thou break a leaf driven to and fro? and wilt thou pursue the dry stubble?
JOB|13|26|For thou writest bitter things against me, and makest me to possess the iniquities of my youth.
JOB|13|27|Thou puttest my feet also in the stocks, and lookest narrowly unto all my paths; thou settest a print upon the heels of my feet.
JOB|13|28|And he, as a rotten thing, consumeth, as a garment that is moth eaten.
JOB|14|1|Man that is born of a woman is of few days and full of trouble.
JOB|14|2|He cometh forth like a flower, and is cut down: he fleeth also as a shadow, and continueth not.
JOB|14|3|And doth thou open thine eyes upon such an one, and bringest me into judgment with thee?
JOB|14|4|Who can bring a clean thing out of an unclean? not one.
JOB|14|5|Seeing his days are determined, the number of his months are with thee, thou hast appointed his bounds that he cannot pass;
JOB|14|6|Turn from him, that he may rest, till he shall accomplish, as an hireling, his day.
JOB|14|7|For there is hope of a tree, if it be cut down, that it will sprout again, and that the tender branch thereof will not cease.
JOB|14|8|Though the root thereof wax old in the earth, and the stock thereof die in the ground;
JOB|14|9|Yet through the scent of water it will bud, and bring forth boughs like a plant.
JOB|14|10|But man dieth, and wasteth away: yea, man giveth up the ghost, and where is he?
JOB|14|11|As the waters fail from the sea, and the flood decayeth and drieth up:
JOB|14|12|So man lieth down, and riseth not: till the heavens be no more, they shall not awake, nor be raised out of their sleep.
JOB|14|13|O that thou wouldest hide me in the grave, that thou wouldest keep me secret, until thy wrath be past, that thou wouldest appoint me a set time, and remember me!
JOB|14|14|If a man die, shall he live again? all the days of my appointed time will I wait, till my change come.
JOB|14|15|Thou shalt call, and I will answer thee: thou wilt have a desire to the work of thine hands.
JOB|14|16|For now thou numberest my steps: dost thou not watch over my sin?
JOB|14|17|My transgression is sealed up in a bag, and thou sewest up mine iniquity.
JOB|14|18|And surely the mountains falling cometh to nought, and the rock is removed out of his place.
JOB|14|19|The waters wear the stones: thou washest away the things which grow out of the dust of the earth; and thou destroyest the hope of man.
JOB|14|20|Thou prevailest for ever against him, and he passeth: thou changest his countenance, and sendest him away.
JOB|14|21|His sons come to honour, and he knoweth it not; and they are brought low, but he perceiveth it not of them.
JOB|14|22|But his flesh upon him shall have pain, and his soul within him shall mourn.
JOB|15|1|Then answered Eliphaz the Temanite, and said,
JOB|15|2|Should a wise man utter vain knowledge, and fill his belly with the east wind?
JOB|15|3|Should he reason with unprofitable talk? or with speeches wherewith he can do no good?
JOB|15|4|Yea, thou castest off fear, and restrainest prayer before God.
JOB|15|5|For thy mouth uttereth thine iniquity, and thou choosest the tongue of the crafty.
JOB|15|6|Thine own mouth condemneth thee, and not I: yea, thine own lips testify against thee.
JOB|15|7|Art thou the first man that was born? or wast thou made before the hills?
JOB|15|8|Hast thou heard the secret of God? and dost thou restrain wisdom to thyself?
JOB|15|9|What knowest thou, that we know not? what understandest thou, which is not in us?
JOB|15|10|With us are both the grayheaded and very aged men, much elder than thy father.
JOB|15|11|Are the consolations of God small with thee? is there any secret thing with thee?
JOB|15|12|Why doth thine heart carry thee away? and what do thy eyes wink at,
JOB|15|13|That thou turnest thy spirit against God, and lettest such words go out of thy mouth?
JOB|15|14|What is man, that he should be clean? and he which is born of a woman, that he should be righteous?
JOB|15|15|Behold, he putteth no trust in his saints; yea, the heavens are not clean in his sight.
JOB|15|16|How much more abominable and filthy is man, which drinketh iniquity like water?
JOB|15|17|I will shew thee, hear me; and that which I have seen I will declare;
JOB|15|18|Which wise men have told from their fathers, and have not hid it:
JOB|15|19|Unto whom alone the earth was given, and no stranger passed among them.
JOB|15|20|The wicked man travaileth with pain all his days, and the number of years is hidden to the oppressor.
JOB|15|21|A dreadful sound is in his ears: in prosperity the destroyer shall come upon him.
JOB|15|22|He believeth not that he shall return out of darkness, and he is waited for of the sword.
JOB|15|23|He wandereth abroad for bread, saying, Where is it? he knoweth that the day of darkness is ready at his hand.
JOB|15|24|Trouble and anguish shall make him afraid; they shall prevail against him, as a king ready to the battle.
JOB|15|25|For he stretcheth out his hand against God, and strengtheneth himself against the Almighty.
JOB|15|26|He runneth upon him, even on his neck, upon the thick bosses of his bucklers:
JOB|15|27|Because he covereth his face with his fatness, and maketh collops of fat on his flanks.
JOB|15|28|And he dwelleth in desolate cities, and in houses which no man inhabiteth, which are ready to become heaps.
JOB|15|29|He shall not be rich, neither shall his substance continue, neither shall he prolong the perfection thereof upon the earth.
JOB|15|30|He shall not depart out of darkness; the flame shall dry up his branches, and by the breath of his mouth shall he go away.
JOB|15|31|Let not him that is deceived trust in vanity: for vanity shall be his recompence.
JOB|15|32|It shall be accomplished before his time, and his branch shall not be green.
JOB|15|33|He shall shake off his unripe grape as the vine, and shall cast off his flower as the olive.
JOB|15|34|For the congregation of hypocrites shall be desolate, and fire shall consume the tabernacles of bribery.
JOB|15|35|They conceive mischief, and bring forth vanity, and their belly prepareth deceit.
JOB|16|1|Then Job answered and said,
JOB|16|2|I have heard many such things: miserable comforters are ye all.
JOB|16|3|Shall vain words have an end? or what emboldeneth thee that thou answerest?
JOB|16|4|I also could speak as ye do: if your soul were in my soul's stead, I could heap up words against you, and shake mine head at you.
JOB|16|5|But I would strengthen you with my mouth, and the moving of my lips should asswage your grief.
JOB|16|6|Though I speak, my grief is not asswaged: and though I forbear, what am I eased?
JOB|16|7|But now he hath made me weary: thou hast made desolate all my company.
JOB|16|8|And thou hast filled me with wrinkles, which is a witness against me: and my leanness rising up in me beareth witness to my face.
JOB|16|9|He teareth me in his wrath, who hateth me: he gnasheth upon me with his teeth; mine enemy sharpeneth his eyes upon me.
JOB|16|10|They have gaped upon me with their mouth; they have smitten me upon the cheek reproachfully; they have gathered themselves together against me.
JOB|16|11|God hath delivered me to the ungodly, and turned me over into the hands of the wicked.
JOB|16|12|I was at ease, but he hath broken me asunder: he hath also taken me by my neck, and shaken me to pieces, and set me up for his mark.
JOB|16|13|His archers compass me round about, he cleaveth my reins asunder, and doth not spare; he poureth out my gall upon the ground.
JOB|16|14|He breaketh me with breach upon breach, he runneth upon me like a giant.
JOB|16|15|I have sewed sackcloth upon my skin, and defiled my horn in the dust.
JOB|16|16|My face is foul with weeping, and on my eyelids is the shadow of death;
JOB|16|17|Not for any injustice in mine hands: also my prayer is pure.
JOB|16|18|O earth, cover not thou my blood, and let my cry have no place.
JOB|16|19|Also now, behold, my witness is in heaven, and my record is on high.
JOB|16|20|My friends scorn me: but mine eye poureth out tears unto God.
JOB|16|21|O that one might plead for a man with God, as a man pleadeth for his neighbour!
JOB|16|22|When a few years are come, then I shall go the way whence I shall not return.
JOB|17|1|My breath is corrupt, my days are extinct, the graves are ready for me.
JOB|17|2|Are there not mockers with me? and doth not mine eye continue in their provocation?
JOB|17|3|Lay down now, put me in a surety with thee; who is he that will strike hands with me?
JOB|17|4|For thou hast hid their heart from understanding: therefore shalt thou not exalt them.
JOB|17|5|He that speaketh flattery to his friends, even the eyes of his children shall fail.
JOB|17|6|He hath made me also a byword of the people; and aforetime I was as a tabret.
JOB|17|7|Mine eye also is dim by reason of sorrow, and all my members are as a shadow.
JOB|17|8|Upright men shall be astonied at this, and the innocent shall stir up himself against the hypocrite.
JOB|17|9|The righteous also shall hold on his way, and he that hath clean hands shall be stronger and stronger.
JOB|17|10|But as for you all, do ye return, and come now: for I cannot find one wise man among you.
JOB|17|11|My days are past, my purposes are broken off, even the thoughts of my heart.
JOB|17|12|They change the night into day: the light is short because of darkness.
JOB|17|13|If I wait, the grave is mine house: I have made my bed in the darkness.
JOB|17|14|I have said to corruption, Thou art my father: to the worm, Thou art my mother, and my sister.
JOB|17|15|And where is now my hope? as for my hope, who shall see it?
JOB|17|16|They shall go down to the bars of the pit, when our rest together is in the dust.
JOB|18|1|Then answered Bildad the Shuhite, and said,
JOB|18|2|How long will it be ere ye make an end of words? mark, and afterwards we will speak.
JOB|18|3|Wherefore are we counted as beasts, and reputed vile in your sight?
JOB|18|4|He teareth himself in his anger: shall the earth be forsaken for thee? and shall the rock be removed out of his place?
JOB|18|5|Yea, the light of the wicked shall be put out, and the spark of his fire shall not shine.
JOB|18|6|The light shall be dark in his tabernacle, and his candle shall be put out with him.
JOB|18|7|The steps of his strength shall be straitened, and his own counsel shall cast him down.
JOB|18|8|For he is cast into a net by his own feet, and he walketh upon a snare.
JOB|18|9|The gin shall take him by the heel, and the robber shall prevail against him.
JOB|18|10|The snare is laid for him in the ground, and a trap for him in the way.
JOB|18|11|Terrors shall make him afraid on every side, and shall drive him to his feet.
JOB|18|12|His strength shall be hungerbitten, and destruction shall be ready at his side.
JOB|18|13|It shall devour the strength of his skin: even the firstborn of death shall devour his strength.
JOB|18|14|His confidence shall be rooted out of his tabernacle, and it shall bring him to the king of terrors.
JOB|18|15|It shall dwell in his tabernacle, because it is none of his: brimstone shall be scattered upon his habitation.
JOB|18|16|His roots shall be dried up beneath, and above shall his branch be cut off.
JOB|18|17|His remembrance shall perish from the earth, and he shall have no name in the street.
JOB|18|18|He shall be driven from light into darkness, and chased out of the world.
JOB|18|19|He shall neither have son nor nephew among his people, nor any remaining in his dwellings.
JOB|18|20|They that come after him shall be astonied at his day, as they that went before were affrighted.
JOB|18|21|Surely such are the dwellings of the wicked, and this is the place of him that knoweth not God.
JOB|19|1|Then Job answered and said,
JOB|19|2|How long will ye vex my soul, and break me in pieces with words?
JOB|19|3|These ten times have ye reproached me: ye are not ashamed that ye make yourselves strange to me.
JOB|19|4|And be it indeed that I have erred, mine error remaineth with myself.
JOB|19|5|If indeed ye will magnify yourselves against me, and plead against me my reproach:
JOB|19|6|Know now that God hath overthrown me, and hath compassed me with his net.
JOB|19|7|Behold, I cry out of wrong, but I am not heard: I cry aloud, but there is no judgment.
JOB|19|8|He hath fenced up my way that I cannot pass, and he hath set darkness in my paths.
JOB|19|9|He hath stripped me of my glory, and taken the crown from my head.
JOB|19|10|He hath destroyed me on every side, and I am gone: and mine hope hath he removed like a tree.
JOB|19|11|He hath also kindled his wrath against me, and he counteth me unto him as one of his enemies.
JOB|19|12|His troops come together, and raise up their way against me, and encamp round about my tabernacle.
JOB|19|13|He hath put my brethren far from me, and mine acquaintance are verily estranged from me.
JOB|19|14|My kinsfolk have failed, and my familiar friends have forgotten me.
JOB|19|15|They that dwell in mine house, and my maids, count me for a stranger: I am an alien in their sight.
JOB|19|16|I called my servant, and he gave me no answer; I intreated him with my mouth.
JOB|19|17|My breath is strange to my wife, though I intreated for the children's sake of mine own body.
JOB|19|18|Yea, young children despised me; I arose, and they spake against me.
JOB|19|19|All my inward friends abhorred me: and they whom I loved are turned against me.
JOB|19|20|My bone cleaveth to my skin and to my flesh, and I am escaped with the skin of my teeth.
JOB|19|21|Have pity upon me, have pity upon me, O ye my friends; for the hand of God hath touched me.
JOB|19|22|Why do ye persecute me as God, and are not satisfied with my flesh?
JOB|19|23|Oh that my words were now written! oh that they were printed in a book!
JOB|19|24|That they were graven with an iron pen and lead in the rock for ever!
JOB|19|25|For I know that my redeemer liveth, and that he shall stand at the latter day upon the earth:
JOB|19|26|And though after my skin worms destroy this body, yet in my flesh shall I see God:
JOB|19|27|Whom I shall see for myself, and mine eyes shall behold, and not another; though my reins be consumed within me.
JOB|19|28|But ye should say, Why persecute we him, seeing the root of the matter is found in me?
JOB|19|29|Be ye afraid of the sword: for wrath bringeth the punishments of the sword, that ye may know there is a judgment.
JOB|20|1|Then answered Zophar the Naamathite, and said,
JOB|20|2|Therefore do my thoughts cause me to answer, and for this I make haste.
JOB|20|3|I have heard the check of my reproach, and the spirit of my understanding causeth me to answer.
JOB|20|4|Knowest thou not this of old, since man was placed upon earth,
JOB|20|5|That the triumphing of the wicked is short, and the joy of the hypocrite but for a moment?
JOB|20|6|Though his excellency mount up to the heavens, and his head reach unto the clouds;
JOB|20|7|Yet he shall perish for ever like his own dung: they which have seen him shall say, Where is he?
JOB|20|8|He shall fly away as a dream, and shall not be found: yea, he shall be chased away as a vision of the night.
JOB|20|9|The eye also which saw him shall see him no more; neither shall his place any more behold him.
JOB|20|10|His children shall seek to please the poor, and his hands shall restore their goods.
JOB|20|11|His bones are full of the sin of his youth, which shall lie down with him in the dust.
JOB|20|12|Though wickedness be sweet in his mouth, though he hide it under his tongue;
JOB|20|13|Though he spare it, and forsake it not; but keep it still within his mouth:
JOB|20|14|Yet his meat in his bowels is turned, it is the gall of asps within him.
JOB|20|15|He hath swallowed down riches, and he shall vomit them up again: God shall cast them out of his belly.
JOB|20|16|He shall suck the poison of asps: the viper's tongue shall slay him.
JOB|20|17|He shall not see the rivers, the floods, the brooks of honey and butter.
JOB|20|18|That which he laboured for shall he restore, and shall not swallow it down: according to his substance shall the restitution be, and he shall not rejoice therein.
JOB|20|19|Because he hath oppressed and hath forsaken the poor; because he hath violently taken away an house which he builded not;
JOB|20|20|Surely he shall not feel quietness in his belly, he shall not save of that which he desired.
JOB|20|21|There shall none of his meat be left; therefore shall no man look for his goods.
JOB|20|22|In the fulness of his sufficiency he shall be in straits: every hand of the wicked shall come upon him.
JOB|20|23|When he is about to fill his belly, God shall cast the fury of his wrath upon him, and shall rain it upon him while he is eating.
JOB|20|24|He shall flee from the iron weapon, and the bow of steel shall strike him through.
JOB|20|25|It is drawn, and cometh out of the body; yea, the glittering sword cometh out of his gall: terrors are upon him.
JOB|20|26|All darkness shall be hid in his secret places: a fire not blown shall consume him; it shall go ill with him that is left in his tabernacle.
JOB|20|27|The heaven shall reveal his iniquity; and the earth shall rise up against him.
JOB|20|28|The increase of his house shall depart, and his goods shall flow away in the day of his wrath.
JOB|20|29|This is the portion of a wicked man from God, and the heritage appointed unto him by God.
JOB|21|1|But Job answered and said,
JOB|21|2|Hear diligently my speech, and let this be your consolations.
JOB|21|3|Suffer me that I may speak; and after that I have spoken, mock on.
JOB|21|4|As for me, is my complaint to man? and if it were so, why should not my spirit be troubled?
JOB|21|5|Mark me, and be astonished, and lay your hand upon your mouth.
JOB|21|6|Even when I remember I am afraid, and trembling taketh hold on my flesh.
JOB|21|7|Wherefore do the wicked live, become old, yea, are mighty in power?
JOB|21|8|Their seed is established in their sight with them, and their offspring before their eyes.
JOB|21|9|Their houses are safe from fear, neither is the rod of God upon them.
JOB|21|10|Their bull gendereth, and faileth not; their cow calveth, and casteth not her calf.
JOB|21|11|They send forth their little ones like a flock, and their children dance.
JOB|21|12|They take the timbrel and harp, and rejoice at the sound of the organ.
JOB|21|13|They spend their days in wealth, and in a moment go down to the grave.
JOB|21|14|Therefore they say unto God, Depart from us; for we desire not the knowledge of thy ways.
JOB|21|15|What is the Almighty, that we should serve him? and what profit should we have, if we pray unto him?
JOB|21|16|Lo, their good is not in their hand: the counsel of the wicked is far from me.
JOB|21|17|How oft is the candle of the wicked put out! and how oft cometh their destruction upon them! God distributeth sorrows in his anger.
JOB|21|18|They are as stubble before the wind, and as chaff that the storm carrieth away.
JOB|21|19|God layeth up his iniquity for his children: he rewardeth him, and he shall know it.
JOB|21|20|His eyes shall see his destruction, and he shall drink of the wrath of the Almighty.
JOB|21|21|For what pleasure hath he in his house after him, when the number of his months is cut off in the midst?
JOB|21|22|Shall any teach God knowledge? seeing he judgeth those that are high.
JOB|21|23|One dieth in his full strength, being wholly at ease and quiet.
JOB|21|24|His breasts are full of milk, and his bones are moistened with marrow.
JOB|21|25|And another dieth in the bitterness of his soul, and never eateth with pleasure.
JOB|21|26|They shall lie down alike in the dust, and the worms shall cover them.
JOB|21|27|Behold, I know your thoughts, and the devices which ye wrongfully imagine against me.
JOB|21|28|For ye say, Where is the house of the prince? and where are the dwelling places of the wicked?
JOB|21|29|Have ye not asked them that go by the way? and do ye not know their tokens,
JOB|21|30|That the wicked is reserved to the day of destruction? they shall be brought forth to the day of wrath.
JOB|21|31|Who shall declare his way to his face? and who shall repay him what he hath done?
JOB|21|32|Yet shall he be brought to the grave, and shall remain in the tomb.
JOB|21|33|The clods of the valley shall be sweet unto him, and every man shall draw after him, as there are innumerable before him.
JOB|21|34|How then comfort ye me in vain, seeing in your answers there remaineth falsehood?
JOB|22|1|Then Eliphaz the Temanite answered and said,
JOB|22|2|Can a man be profitable unto God, as he that is wise may be profitable unto himself?
JOB|22|3|Is it any pleasure to the Almighty, that thou art righteous? or is it gain to him, that thou makest thy ways perfect?
JOB|22|4|Will he reprove thee for fear of thee? will he enter with thee into judgment?
JOB|22|5|Is not thy wickedness great? and thine iniquities infinite?
JOB|22|6|For thou hast taken a pledge from thy brother for nought, and stripped the naked of their clothing.
JOB|22|7|Thou hast not given water to the weary to drink, and thou hast withholden bread from the hungry.
JOB|22|8|But as for the mighty man, he had the earth; and the honourable man dwelt in it.
JOB|22|9|Thou hast sent widows away empty, and the arms of the fatherless have been broken.
JOB|22|10|Therefore snares are round about thee, and sudden fear troubleth thee;
JOB|22|11|Or darkness, that thou canst not see; and abundance of waters cover thee.
JOB|22|12|Is not God in the height of heaven? and behold the height of the stars, how high they are!
JOB|22|13|And thou sayest, How doth God know? can he judge through the dark cloud?
JOB|22|14|Thick clouds are a covering to him, that he seeth not; and he walketh in the circuit of heaven.
JOB|22|15|Hast thou marked the old way which wicked men have trodden?
JOB|22|16|Which were cut down out of time, whose foundation was overflown with a flood:
JOB|22|17|Which said unto God, Depart from us: and what can the Almighty do for them?
JOB|22|18|Yet he filled their houses with good things: but the counsel of the wicked is far from me.
JOB|22|19|The righteous see it, and are glad: and the innocent laugh them to scorn.
JOB|22|20|Whereas our substance is not cut down, but the remnant of them the fire consumeth.
JOB|22|21|Acquaint now thyself with him, and be at peace: thereby good shall come unto thee.
JOB|22|22|Receive, I pray thee, the law from his mouth, and lay up his words in thine heart.
JOB|22|23|If thou return to the Almighty, thou shalt be built up, thou shalt put away iniquity far from thy tabernacles.
JOB|22|24|Then shalt thou lay up gold as dust, and the gold of Ophir as the stones of the brooks.
JOB|22|25|Yea, the Almighty shall be thy defence, and thou shalt have plenty of silver.
JOB|22|26|For then shalt thou have thy delight in the Almighty, and shalt lift up thy face unto God.
JOB|22|27|Thou shalt make thy prayer unto him, and he shall hear thee, and thou shalt pay thy vows.
JOB|22|28|Thou shalt also decree a thing, and it shall be established unto thee: and the light shall shine upon thy ways.
JOB|22|29|When men are cast down, then thou shalt say, There is lifting up; and he shall save the humble person.
JOB|22|30|He shall deliver the island of the innocent: and it is delivered by the pureness of thine hands.
JOB|23|1|Then Job answered and said,
JOB|23|2|Even to day is my complaint bitter: my stroke is heavier than my groaning.
JOB|23|3|Oh that I knew where I might find him! that I might come even to his seat!
JOB|23|4|I would order my cause before him, and fill my mouth with arguments.
JOB|23|5|I would know the words which he would answer me, and understand what he would say unto me.
JOB|23|6|Will he plead against me with his great power? No; but he would put strength in me.
JOB|23|7|There the righteous might dispute with him; so should I be delivered for ever from my judge.
JOB|23|8|Behold, I go forward, but he is not there; and backward, but I cannot perceive him:
JOB|23|9|On the left hand, where he doth work, but I cannot behold him: he hideth himself on the right hand, that I cannot see him:
JOB|23|10|But he knoweth the way that I take: when he hath tried me, I shall come forth as gold.
JOB|23|11|My foot hath held his steps, his way have I kept, and not declined.
JOB|23|12|Neither have I gone back from the commandment of his lips; I have esteemed the words of his mouth more than my necessary food.
JOB|23|13|But he is in one mind, and who can turn him? and what his soul desireth, even that he doeth.
JOB|23|14|For he performeth the thing that is appointed for me: and many such things are with him.
JOB|23|15|Therefore am I troubled at his presence: when I consider, I am afraid of him.
JOB|23|16|For God maketh my heart soft, and the Almighty troubleth me:
JOB|23|17|Because I was not cut off before the darkness, neither hath he covered the darkness from my face.
JOB|24|1|Why, seeing times are not hidden from the Almighty, do they that know him not see his days?
JOB|24|2|Some remove the landmarks; they violently take away flocks, and feed thereof.
JOB|24|3|They drive away the ass of the fatherless, they take the widow's ox for a pledge.
JOB|24|4|They turn the needy out of the way: the poor of the earth hide themselves together.
JOB|24|5|Behold, as wild asses in the desert, go they forth to their work; rising betimes for a prey: the wilderness yieldeth food for them and for their children.
JOB|24|6|They reap every one his corn in the field: and they gather the vintage of the wicked.
JOB|24|7|They cause the naked to lodge without clothing, that they have no covering in the cold.
JOB|24|8|They are wet with the showers of the mountains, and embrace the rock for want of a shelter.
JOB|24|9|They pluck the fatherless from the breast, and take a pledge of the poor.
JOB|24|10|They cause him to go naked without clothing, and they take away the sheaf from the hungry;
JOB|24|11|Which make oil within their walls, and tread their winepresses, and suffer thirst.
JOB|24|12|Men groan from out of the city, and the soul of the wounded crieth out: yet God layeth not folly to them.
JOB|24|13|They are of those that rebel against the light; they know not the ways thereof, nor abide in the paths thereof.
JOB|24|14|The murderer rising with the light killeth the poor and needy, and in the night is as a thief.
JOB|24|15|The eye also of the adulterer waiteth for the twilight, saying, No eye shall see me: and disguiseth his face.
JOB|24|16|In the dark they dig through houses, which they had marked for themselves in the daytime: they know not the light.
JOB|24|17|For the morning is to them even as the shadow of death: if one know them, they are in the terrors of the shadow of death.
JOB|24|18|He is swift as the waters; their portion is cursed in the earth: he beholdeth not the way of the vineyards.
JOB|24|19|Drought and heat consume the snow waters: so doth the grave those which have sinned.
JOB|24|20|The womb shall forget him; the worm shall feed sweetly on him; he shall be no more remembered; and wickedness shall be broken as a tree.
JOB|24|21|He evil entreateth the barren that beareth not: and doeth not good to the widow.
JOB|24|22|He draweth also the mighty with his power: he riseth up, and no man is sure of life.
JOB|24|23|Though it be given him to be in safety, whereon he resteth; yet his eyes are upon their ways.
JOB|24|24|They are exalted for a little while, but are gone and brought low; they are taken out of the way as all other, and cut off as the tops of the ears of corn.
JOB|24|25|And if it be not so now, who will make me a liar, and make my speech nothing worth?
JOB|25|1|Then answered Bildad the Shuhite, and said,
JOB|25|2|Dominion and fear are with him, he maketh peace in his high places.
JOB|25|3|Is there any number of his armies? and upon whom doth not his light arise?
JOB|25|4|How then can man be justified with God? or how can he be clean that is born of a woman?
JOB|25|5|Behold even to the moon, and it shineth not; yea, the stars are not pure in his sight.
JOB|25|6|How much less man, that is a worm? and the son of man, which is a worm?
JOB|26|1|But Job answered and said,
JOB|26|2|How hast thou helped him that is without power? how savest thou the arm that hath no strength?
JOB|26|3|How hast thou counselled him that hath no wisdom? and how hast thou plentifully declared the thing as it is?
JOB|26|4|To whom hast thou uttered words? and whose spirit came from thee?
JOB|26|5|Dead things are formed from under the waters, and the inhabitants thereof.
JOB|26|6|Hell is naked before him, and destruction hath no covering.
JOB|26|7|He stretcheth out the north over the empty place, and hangeth the earth upon nothing.
JOB|26|8|He bindeth up the waters in his thick clouds; and the cloud is not rent under them.
JOB|26|9|He holdeth back the face of his throne, and spreadeth his cloud upon it.
JOB|26|10|He hath compassed the waters with bounds, until the day and night come to an end.
JOB|26|11|The pillars of heaven tremble and are astonished at his reproof.
JOB|26|12|He divideth the sea with his power, and by his understanding he smiteth through the proud.
JOB|26|13|By his spirit he hath garnished the heavens; his hand hath formed the crooked serpent.
JOB|26|14|Lo, these are parts of his ways: but how little a portion is heard of him? but the thunder of his power who can understand?
JOB|27|1|Moreover Job continued his parable, and said,
JOB|27|2|As God liveth, who hath taken away my judgment; and the Almighty, who hath vexed my soul;
JOB|27|3|All the while my breath is in me, and the spirit of God is in my nostrils;
JOB|27|4|My lips shall not speak wickedness, nor my tongue utter deceit.
JOB|27|5|God forbid that I should justify you: till I die I will not remove mine integrity from me.
JOB|27|6|My righteousness I hold fast, and will not let it go: my heart shall not reproach me so long as I live.
JOB|27|7|Let mine enemy be as the wicked, and he that riseth up against me as the unrighteous.
JOB|27|8|For what is the hope of the hypocrite, though he hath gained, when God taketh away his soul?
JOB|27|9|Will God hear his cry when trouble cometh upon him?
JOB|27|10|Will he delight himself in the Almighty? will he always call upon God?
JOB|27|11|I will teach you by the hand of God: that which is with the Almighty will I not conceal.
JOB|27|12|Behold, all ye yourselves have seen it; why then are ye thus altogether vain?
JOB|27|13|This is the portion of a wicked man with God, and the heritage of oppressors, which they shall receive of the Almighty.
JOB|27|14|If his children be multiplied, it is for the sword: and his offspring shall not be satisfied with bread.
JOB|27|15|Those that remain of him shall be buried in death: and his widows shall not weep.
JOB|27|16|Though he heap up silver as the dust, and prepare raiment as the clay;
JOB|27|17|He may prepare it, but the just shall put it on, and the innocent shall divide the silver.
JOB|27|18|He buildeth his house as a moth, and as a booth that the keeper maketh.
JOB|27|19|The rich man shall lie down, but he shall not be gathered: he openeth his eyes, and he is not.
JOB|27|20|Terrors take hold on him as waters, a tempest stealeth him away in the night.
JOB|27|21|The east wind carrieth him away, and he departeth: and as a storm hurleth him out of his place.
JOB|27|22|For God shall cast upon him, and not spare: he would fain flee out of his hand.
JOB|27|23|Men shall clap their hands at him, and shall hiss him out of his place.
JOB|28|1|Surely there is a vein for the silver, and a place for gold where they fine it.
JOB|28|2|Iron is taken out of the earth, and brass is molten out of the stone.
JOB|28|3|He setteth an end to darkness, and searcheth out all perfection: the stones of darkness, and the shadow of death.
JOB|28|4|The flood breaketh out from the inhabitant; even the waters forgotten of the foot: they are dried up, they are gone away from men.
JOB|28|5|As for the earth, out of it cometh bread: and under it is turned up as it were fire.
JOB|28|6|The stones of it are the place of sapphires: and it hath dust of gold.
JOB|28|7|There is a path which no fowl knoweth, and which the vulture's eye hath not seen:
JOB|28|8|The lion's whelps have not trodden it, nor the fierce lion passed by it.
JOB|28|9|He putteth forth his hand upon the rock; he overturneth the mountains by the roots.
JOB|28|10|He cutteth out rivers among the rocks; and his eye seeth every precious thing.
JOB|28|11|He bindeth the floods from overflowing; and the thing that is hid bringeth he forth to light.
JOB|28|12|But where shall wisdom be found? and where is the place of understanding?
JOB|28|13|Man knoweth not the price thereof; neither is it found in the land of the living.
JOB|28|14|The depth saith, It is not in me: and the sea saith, It is not with me.
JOB|28|15|It cannot be gotten for gold, neither shall silver be weighed for the price thereof.
JOB|28|16|It cannot be valued with the gold of Ophir, with the precious onyx, or the sapphire.
JOB|28|17|The gold and the crystal cannot equal it: and the exchange of it shall not be for jewels of fine gold.
JOB|28|18|No mention shall be made of coral, or of pearls: for the price of wisdom is above rubies.
JOB|28|19|The topaz of Ethiopia shall not equal it, neither shall it be valued with pure gold.
JOB|28|20|Whence then cometh wisdom? and where is the place of understanding?
JOB|28|21|Seeing it is hid from the eyes of all living, and kept close from the fowls of the air.
JOB|28|22|Destruction and death say, We have heard the fame thereof with our ears.
JOB|28|23|God understandeth the way thereof, and he knoweth the place thereof.
JOB|28|24|For he looketh to the ends of the earth, and seeth under the whole heaven;
JOB|28|25|To make the weight for the winds; and he weigheth the waters by measure.
JOB|28|26|When he made a decree for the rain, and a way for the lightning of the thunder:
JOB|28|27|Then did he see it, and declare it; he prepared it, yea, and searched it out.
JOB|28|28|And unto man he said, Behold, the fear of the LORD, that is wisdom; and to depart from evil is understanding.
JOB|29|1|Moreover Job continued his parable, and said,
JOB|29|2|Oh that I were as in months past, as in the days when God preserved me;
JOB|29|3|When his candle shined upon my head, and when by his light I walked through darkness;
JOB|29|4|As I was in the days of my youth, when the secret of God was upon my tabernacle;
JOB|29|5|When the Almighty was yet with me, when my children were about me;
JOB|29|6|When I washed my steps with butter, and the rock poured me out rivers of oil;
JOB|29|7|When I went out to the gate through the city, when I prepared my seat in the street!
JOB|29|8|The young men saw me, and hid themselves: and the aged arose, and stood up.
JOB|29|9|The princes refrained talking, and laid their hand on their mouth.
JOB|29|10|The nobles held their peace, and their tongue cleaved to the roof of their mouth.
JOB|29|11|When the ear heard me, then it blessed me; and when the eye saw me, it gave witness to me:
JOB|29|12|Because I delivered the poor that cried, and the fatherless, and him that had none to help him.
JOB|29|13|The blessing of him that was ready to perish came upon me: and I caused the widow's heart to sing for joy.
JOB|29|14|I put on righteousness, and it clothed me: my judgment was as a robe and a diadem.
JOB|29|15|I was eyes to the blind, and feet was I to the lame.
JOB|29|16|I was a father to the poor: and the cause which I knew not I searched out.
JOB|29|17|And I brake the jaws of the wicked, and plucked the spoil out of his teeth.
JOB|29|18|Then I said, I shall die in my nest, and I shall multiply my days as the sand.
JOB|29|19|My root was spread out by the waters, and the dew lay all night upon my branch.
JOB|29|20|My glory was fresh in me, and my bow was renewed in my hand.
JOB|29|21|Unto me men gave ear, and waited, and kept silence at my counsel.
JOB|29|22|After my words they spake not again; and my speech dropped upon them.
JOB|29|23|And they waited for me as for the rain; and they opened their mouth wide as for the latter rain.
JOB|29|24|If I laughed on them, they believed it not; and the light of my countenance they cast not down.
JOB|29|25|I chose out their way, and sat chief, and dwelt as a king in the army, as one that comforteth the mourners.
JOB|30|1|But now they that are younger than I have me in derision, whose fathers I would have disdained to have set with the dogs of my flock.
JOB|30|2|Yea, whereto might the strength of their hands profit me, in whom old age was perished?
JOB|30|3|For want and famine they were solitary; fleeing into the wilderness in former time desolate and waste.
JOB|30|4|Who cut up mallows by the bushes, and juniper roots for their meat.
JOB|30|5|They were driven forth from among men, (they cried after them as after a thief;)
JOB|30|6|To dwell in the cliffs of the valleys, in caves of the earth, and in the rocks.
JOB|30|7|Among the bushes they brayed; under the nettles they were gathered together.
JOB|30|8|They were children of fools, yea, children of base men: they were viler than the earth.
JOB|30|9|And now am I their song, yea, I am their byword.
JOB|30|10|They abhor me, they flee far from me, and spare not to spit in my face.
JOB|30|11|Because he hath loosed my cord, and afflicted me, they have also let loose the bridle before me.
JOB|30|12|Upon my right hand rise the youth; they push away my feet, and they raise up against me the ways of their destruction.
JOB|30|13|They mar my path, they set forward my calamity, they have no helper.
JOB|30|14|They came upon me as a wide breaking in of waters: in the desolation they rolled themselves upon me.
JOB|30|15|Terrors are turned upon me: they pursue my soul as the wind: and my welfare passeth away as a cloud.
JOB|30|16|And now my soul is poured out upon me; the days of affliction have taken hold upon me.
JOB|30|17|My bones are pierced in me in the night season: and my sinews take no rest.
JOB|30|18|By the great force of my disease is my garment changed: it bindeth me about as the collar of my coat.
JOB|30|19|He hath cast me into the mire, and I am become like dust and ashes.
JOB|30|20|I cry unto thee, and thou dost not hear me: I stand up, and thou regardest me not.
JOB|30|21|Thou art become cruel to me: with thy strong hand thou opposest thyself against me.
JOB|30|22|Thou liftest me up to the wind; thou causest me to ride upon it, and dissolvest my substance.
JOB|30|23|For I know that thou wilt bring me to death, and to the house appointed for all living.
JOB|30|24|Howbeit he will not stretch out his hand to the grave, though they cry in his destruction.
JOB|30|25|Did not I weep for him that was in trouble? was not my soul grieved for the poor?
JOB|30|26|When I looked for good, then evil came unto me: and when I waited for light, there came darkness.
JOB|30|27|My bowels boiled, and rested not: the days of affliction prevented me.
JOB|30|28|I went mourning without the sun: I stood up, and I cried in the congregation.
JOB|30|29|I am a brother to dragons, and a companion to owls.
JOB|30|30|My skin is black upon me, and my bones are burned with heat.
JOB|30|31|My harp also is turned to mourning, and my organ into the voice of them that weep.
JOB|31|1|I made a covenant with mine eyes; why then should I think upon a maid?
JOB|31|2|For what portion of God is there from above? and what inheritance of the Almighty from on high?
JOB|31|3|Is not destruction to the wicked? and a strange punishment to the workers of iniquity?
JOB|31|4|Doth not he see my ways, and count all my steps?
JOB|31|5|If I have walked with vanity, or if my foot hath hasted to deceit;
JOB|31|6|Let me be weighed in an even balance that God may know mine integrity.
JOB|31|7|If my step hath turned out of the way, and mine heart walked after mine eyes, and if any blot hath cleaved to mine hands;
JOB|31|8|Then let me sow, and let another eat; yea, let my offspring be rooted out.
JOB|31|9|If mine heart have been deceived by a woman, or if I have laid wait at my neighbour's door;
JOB|31|10|Then let my wife grind unto another, and let others bow down upon her.
JOB|31|11|For this is an heinous crime; yea, it is an iniquity to be punished by the judges.
JOB|31|12|For it is a fire that consumeth to destruction, and would root out all mine increase.
JOB|31|13|If I did despise the cause of my manservant or of my maidservant, when they contended with me;
JOB|31|14|What then shall I do when God riseth up? and when he visiteth, what shall I answer him?
JOB|31|15|Did not he that made me in the womb make him? and did not one fashion us in the womb?
JOB|31|16|If I have withheld the poor from their desire, or have caused the eyes of the widow to fail;
JOB|31|17|Or have eaten my morsel myself alone, and the fatherless hath not eaten thereof;
JOB|31|18|(For from my youth he was brought up with me, as with a father, and I have guided her from my mother's womb;)
JOB|31|19|If I have seen any perish for want of clothing, or any poor without covering;
JOB|31|20|If his loins have not blessed me, and if he were not warmed with the fleece of my sheep;
JOB|31|21|If I have lifted up my hand against the fatherless, when I saw my help in the gate:
JOB|31|22|Then let mine arm fall from my shoulder blade, and mine arm be broken from the bone.
JOB|31|23|For destruction from God was a terror to me, and by reason of his highness I could not endure.
JOB|31|24|If I have made gold my hope, or have said to the fine gold, Thou art my confidence;
JOB|31|25|If I rejoice because my wealth was great, and because mine hand had gotten much;
JOB|31|26|If I beheld the sun when it shined, or the moon walking in brightness;
JOB|31|27|And my heart hath been secretly enticed, or my mouth hath kissed my hand:
JOB|31|28|This also were an iniquity to be punished by the judge: for I should have denied the God that is above.
JOB|31|29|If I rejoice at the destruction of him that hated me, or lifted up myself when evil found him:
JOB|31|30|Neither have I suffered my mouth to sin by wishing a curse to his soul.
JOB|31|31|If the men of my tabernacle said not, Oh that we had of his flesh! we cannot be satisfied.
JOB|31|32|The stranger did not lodge in the street: but I opened my doors to the traveller.
JOB|31|33|If I covered my transgressions as Adam, by hiding mine iniquity in my bosom:
JOB|31|34|Did I fear a great multitude, or did the contempt of families terrify me, that I kept silence, and went not out of the door?
JOB|31|35|Oh that one would hear me! behold, my desire is, that the Almighty would answer me, and that mine adversary had written a book.
JOB|31|36|Surely I would take it upon my shoulder, and bind it as a crown to me.
JOB|31|37|I would declare unto him the number of my steps; as a prince would I go near unto him.
JOB|31|38|If my land cry against me, or that the furrows likewise thereof complain;
JOB|31|39|If I have eaten the fruits thereof without money, or have caused the owners thereof to lose their life:
JOB|31|40|Let thistles grow instead of wheat, and cockle instead of barley. The words of Job are ended.
JOB|32|1|So these three men ceased to answer Job, because he was righteous in his own eyes.
JOB|32|2|Then was kindled the wrath of Elihu the son of Barachel the Buzite, of the kindred of Ram: against Job was his wrath kindled, because he justified himself rather than God.
JOB|32|3|Also against his three friends was his wrath kindled, because they had found no answer, and yet had condemned Job.
JOB|32|4|Now Elihu had waited till Job had spoken, because they were elder than he.
JOB|32|5|When Elihu saw that there was no answer in the mouth of these three men, then his wrath was kindled.
JOB|32|6|And Elihu the son of Barachel the Buzite answered and said, I am young, and ye are very old; wherefore I was afraid, and durst not shew you mine opinion.
JOB|32|7|I said, Days should speak, and multitude of years should teach wisdom.
JOB|32|8|But there is a spirit in man: and the inspiration of the Almighty giveth them understanding.
JOB|32|9|Great men are not always wise: neither do the aged understand judgment.
JOB|32|10|Therefore I said, Hearken to me; I also will shew mine opinion.
JOB|32|11|Behold, I waited for your words; I gave ear to your reasons, whilst ye searched out what to say.
JOB|32|12|Yea, I attended unto you, and, behold, there was none of you that convinced Job, or that answered his words:
JOB|32|13|Lest ye should say, We have found out wisdom: God thrusteth him down, not man.
JOB|32|14|Now he hath not directed his words against me: neither will I answer him with your speeches.
JOB|32|15|They were amazed, they answered no more: they left off speaking.
JOB|32|16|When I had waited, (for they spake not, but stood still, and answered no more;)
JOB|32|17|I said, I will answer also my part, I also will shew mine opinion.
JOB|32|18|For I am full of matter, the spirit within me constraineth me.
JOB|32|19|Behold, my belly is as wine which hath no vent; it is ready to burst like new bottles.
JOB|32|20|I will speak, that I may be refreshed: I will open my lips and answer.
JOB|32|21|Let me not, I pray you, accept any man's person, neither let me give flattering titles unto man.
JOB|32|22|For I know not to give flattering titles; in so doing my maker would soon take me away.
JOB|33|1|Wherefore, Job, I pray thee, hear my speeches, and hearken to all my words.
JOB|33|2|Behold, now I have opened my mouth, my tongue hath spoken in my mouth.
JOB|33|3|My words shall be of the uprightness of my heart: and my lips shall utter knowledge clearly.
JOB|33|4|The spirit of God hath made me, and the breath of the Almighty hath given me life.
JOB|33|5|If thou canst answer me, set thy words in order before me, stand up.
JOB|33|6|Behold, I am according to thy wish in God's stead: I also am formed out of the clay.
JOB|33|7|Behold, my terror shall not make thee afraid, neither shall my hand be heavy upon thee.
JOB|33|8|Surely thou hast spoken in mine hearing, and I have heard the voice of thy words, saying,
JOB|33|9|I am clean without transgression, I am innocent; neither is there iniquity in me.
JOB|33|10|Behold, he findeth occasions against me, he counteth me for his enemy,
JOB|33|11|He putteth my feet in the stocks, he marketh all my paths.
JOB|33|12|Behold, in this thou art not just: I will answer thee, that God is greater than man.
JOB|33|13|Why dost thou strive against him? for he giveth not account of any of his matters.
JOB|33|14|For God speaketh once, yea twice, yet man perceiveth it not.
JOB|33|15|In a dream, in a vision of the night, when deep sleep falleth upon men, in slumberings upon the bed;
JOB|33|16|Then he openeth the ears of men, and sealeth their instruction,
JOB|33|17|That he may withdraw man from his purpose, and hide pride from man.
JOB|33|18|He keepeth back his soul from the pit, and his life from perishing by the sword.
JOB|33|19|He is chastened also with pain upon his bed, and the multitude of his bones with strong pain:
JOB|33|20|So that his life abhorreth bread, and his soul dainty meat.
JOB|33|21|His flesh is consumed away, that it cannot be seen; and his bones that were not seen stick out.
JOB|33|22|Yea, his soul draweth near unto the grave, and his life to the destroyers.
JOB|33|23|If there be a messenger with him, an interpreter, one among a thousand, to shew unto man his uprightness:
JOB|33|24|Then he is gracious unto him, and saith, Deliver him from going down to the pit: I have found a ransom.
JOB|33|25|His flesh shall be fresher than a child's: he shall return to the days of his youth:
JOB|33|26|He shall pray unto God, and he will be favourable unto him: and he shall see his face with joy: for he will render unto man his righteousness.
JOB|33|27|He looketh upon men, and if any say, I have sinned, and perverted that which was right, and it profited me not;
JOB|33|28|He will deliver his soul from going into the pit, and his life shall see the light.
JOB|33|29|Lo, all these things worketh God oftentimes with man,
JOB|33|30|To bring back his soul from the pit, to be enlightened with the light of the living.
JOB|33|31|Mark well, O Job, hearken unto me: hold thy peace, and I will speak.
JOB|33|32|If thou hast anything to say, answer me: speak, for I desire to justify thee.
JOB|33|33|If not, hearken unto me: hold thy peace, and I shall teach thee wisdom.
JOB|34|1|Furthermore Elihu answered and said,
JOB|34|2|Hear my words, O ye wise men; and give ear unto me, ye that have knowledge.
JOB|34|3|For the ear trieth words, as the mouth tasteth meat.
JOB|34|4|Let us choose to us judgment: let us know among ourselves what is good.
JOB|34|5|For Job hath said, I am righteous: and God hath taken away my judgment.
JOB|34|6|Should I lie against my right? my wound is incurable without transgression.
JOB|34|7|What man is like Job, who drinketh up scorning like water?
JOB|34|8|Which goeth in company with the workers of iniquity, and walketh with wicked men.
JOB|34|9|For he hath said, It profiteth a man nothing that he should delight himself with God.
JOB|34|10|Therefore hearken unto me ye men of understanding: far be it from God, that he should do wickedness; and from the Almighty, that he should commit iniquity.
JOB|34|11|For the work of a man shall he render unto him, and cause every man to find according to his ways.
JOB|34|12|Yea, surely God will not do wickedly, neither will the Almighty pervert judgment.
JOB|34|13|Who hath given him a charge over the earth? or who hath disposed the whole world?
JOB|34|14|If he set his heart upon man, if he gather unto himself his spirit and his breath;
JOB|34|15|All flesh shall perish together, and man shall turn again unto dust.
JOB|34|16|If now thou hast understanding, hear this: hearken to the voice of my words.
JOB|34|17|Shall even he that hateth right govern? and wilt thou condemn him that is most just?
JOB|34|18|Is it fit to say to a king, Thou art wicked? and to princes, Ye are ungodly?
JOB|34|19|How much less to him that accepteth not the persons of princes, nor regardeth the rich more than the poor? for they all are the work of his hands.
JOB|34|20|In a moment shall they die, and the people shall be troubled at midnight, and pass away: and the mighty shall be taken away without hand.
JOB|34|21|For his eyes are upon the ways of man, and he seeth all his goings.
JOB|34|22|There is no darkness, nor shadow of death, where the workers of iniquity may hide themselves.
JOB|34|23|For he will not lay upon man more than right; that he should enter into judgment with God.
JOB|34|24|He shall break in pieces mighty men without number, and set others in their stead.
JOB|34|25|Therefore he knoweth their works, and he overturneth them in the night, so that they are destroyed.
JOB|34|26|He striketh them as wicked men in the open sight of others;
JOB|34|27|Because they turned back from him, and would not consider any of his ways:
JOB|34|28|So that they cause the cry of the poor to come unto him, and he heareth the cry of the afflicted.
JOB|34|29|When he giveth quietness, who then can make trouble? and when he hideth his face, who then can behold him? whether it be done against a nation, or against a man only:
JOB|34|30|That the hypocrite reign not, lest the people be ensnared.
JOB|34|31|Surely it is meet to be said unto God, I have borne chastisement, I will not offend any more:
JOB|34|32|That which I see not teach thou me: if I have done iniquity, I will do no more.
JOB|34|33|Should it be according to thy mind? he will recompense it, whether thou refuse, or whether thou choose; and not I: therefore speak what thou knowest.
JOB|34|34|Let men of understanding tell me, and let a wise man hearken unto me.
JOB|34|35|Job hath spoken without knowledge, and his words were without wisdom.
JOB|34|36|My desire is that Job may be tried unto the end because of his answers for wicked men.
JOB|34|37|For he addeth rebellion unto his sin, he clappeth his hands among us, and multiplieth his words against God.
JOB|35|1|Elihu spake moreover, and said,
JOB|35|2|Thinkest thou this to be right, that thou saidst, My righteousness is more than God's?
JOB|35|3|For thou saidst, What advantage will it be unto thee? and, What profit shall I have, if I be cleansed from my sin?
JOB|35|4|I will answer thee, and thy companions with thee.
JOB|35|5|Look unto the heavens, and see; and behold the clouds which are higher than thou.
JOB|35|6|If thou sinnest, what doest thou against him? or if thy transgressions be multiplied, what doest thou unto him?
JOB|35|7|If thou be righteous, what givest thou him? or what receiveth he of thine hand?
JOB|35|8|Thy wickedness may hurt a man as thou art; and thy righteousness may profit the son of man.
JOB|35|9|By reason of the multitude of oppressions they make the oppressed to cry: they cry out by reason of the arm of the mighty.
JOB|35|10|But none saith, Where is God my maker, who giveth songs in the night;
JOB|35|11|Who teacheth us more than the beasts of the earth, and maketh us wiser than the fowls of heaven?
JOB|35|12|There they cry, but none giveth answer, because of the pride of evil men.
JOB|35|13|Surely God will not hear vanity, neither will the Almighty regard it.
JOB|35|14|Although thou sayest thou shalt not see him, yet judgment is before him; therefore trust thou in him.
JOB|35|15|But now, because it is not so, he hath visited in his anger; yet he knoweth it not in great extremity:
JOB|35|16|Therefore doth Job open his mouth in vain; he multiplieth words without knowledge.
JOB|36|1|Elihu also proceeded, and said,
JOB|36|2|Suffer me a little, and I will shew thee that I have yet to speak on God's behalf.
JOB|36|3|I will fetch my knowledge from afar, and will ascribe righteousness to my Maker.
JOB|36|4|For truly my words shall not be false: he that is perfect in knowledge is with thee.
JOB|36|5|Behold, God is mighty, and despiseth not any: he is mighty in strength and wisdom.
JOB|36|6|He preserveth not the life of the wicked: but giveth right to the poor.
JOB|36|7|He withdraweth not his eyes from the righteous: but with kings are they on the throne; yea, he doth establish them for ever, and they are exalted.
JOB|36|8|And if they be bound in fetters, and be holden in cords of affliction;
JOB|36|9|Then he sheweth them their work, and their transgressions that they have exceeded.
JOB|36|10|He openeth also their ear to discipline, and commandeth that they return from iniquity.
JOB|36|11|If they obey and serve him, they shall spend their days in prosperity, and their years in pleasures.
JOB|36|12|But if they obey not, they shall perish by the sword, and they shall die without knowledge.
JOB|36|13|But the hypocrites in heart heap up wrath: they cry not when he bindeth them.
JOB|36|14|They die in youth, and their life is among the unclean.
JOB|36|15|He delivereth the poor in his affliction, and openeth their ears in oppression.
JOB|36|16|Even so would he have removed thee out of the strait into a broad place, where there is no straitness; and that which should be set on thy table should be full of fatness.
JOB|36|17|But thou hast fulfilled the judgment of the wicked: judgment and justice take hold on thee.
JOB|36|18|Because there is wrath, beware lest he take thee away with his stroke: then a great ransom cannot deliver thee.
JOB|36|19|Will he esteem thy riches? no, not gold, nor all the forces of strength.
JOB|36|20|Desire not the night, when people are cut off in their place.
JOB|36|21|Take heed, regard not iniquity: for this hast thou chosen rather than affliction.
JOB|36|22|Behold, God exalteth by his power: who teacheth like him?
JOB|36|23|Who hath enjoined him his way? or who can say, Thou hast wrought iniquity?
JOB|36|24|Remember that thou magnify his work, which men behold.
JOB|36|25|Every man may see it; man may behold it afar off.
JOB|36|26|Behold, God is great, and we know him not, neither can the number of his years be searched out.
JOB|36|27|For he maketh small the drops of water: they pour down rain according to the vapour thereof:
JOB|36|28|Which the clouds do drop and distil upon man abundantly.
JOB|36|29|Also can any understand the spreadings of the clouds, or the noise of his tabernacle?
JOB|36|30|Behold, he spreadeth his light upon it, and covereth the bottom of the sea.
JOB|36|31|For by them judgeth he the people; he giveth meat in abundance.
JOB|36|32|With clouds he covereth the light; and commandeth it not to shine by the cloud that cometh betwixt.
JOB|36|33|The noise thereof sheweth concerning it, the cattle also concerning the vapour.
JOB|37|1|At this also my heart trembleth, and is moved out of his place.
JOB|37|2|Hear attentively the noise of his voice, and the sound that goeth out of his mouth.
JOB|37|3|He directeth it under the whole heaven, and his lightning unto the ends of the earth.
JOB|37|4|After it a voice roareth: he thundereth with the voice of his excellency; and he will not stay them when his voice is heard.
JOB|37|5|God thundereth marvellously with his voice; great things doeth he, which we cannot comprehend.
JOB|37|6|For he saith to the snow, Be thou on the earth; likewise to the small rain, and to the great rain of his strength.
JOB|37|7|He sealeth up the hand of every man; that all men may know his work.
JOB|37|8|Then the beasts go into dens, and remain in their places.
JOB|37|9|Out of the south cometh the whirlwind: and cold out of the north.
JOB|37|10|By the breath of God frost is given: and the breadth of the waters is straitened.
JOB|37|11|Also by watering he wearieth the thick cloud: he scattereth his bright cloud:
JOB|37|12|And it is turned round about by his counsels: that they may do whatsoever he commandeth them upon the face of the world in the earth.
JOB|37|13|He causeth it to come, whether for correction, or for his land, or for mercy.
JOB|37|14|Hearken unto this, O Job: stand still, and consider the wondrous works of God.
JOB|37|15|Dost thou know when God disposed them, and caused the light of his cloud to shine?
JOB|37|16|Dost thou know the balancings of the clouds, the wondrous works of him which is perfect in knowledge?
JOB|37|17|How thy garments are warm, when he quieteth the earth by the south wind?
JOB|37|18|Hast thou with him spread out the sky, which is strong, and as a molten looking glass?
JOB|37|19|Teach us what we shall say unto him; for we cannot order our speech by reason of darkness.
JOB|37|20|Shall it be told him that I speak? if a man speak, surely he shall be swallowed up.
JOB|37|21|And now men see not the bright light which is in the clouds: but the wind passeth, and cleanseth them.
JOB|37|22|Fair weather cometh out of the north: with God is terrible majesty.
JOB|37|23|Touching the Almighty, we cannot find him out: he is excellent in power, and in judgment, and in plenty of justice: he will not afflict.
JOB|37|24|Men do therefore fear him: he respecteth not any that are wise of heart.
JOB|38|1|Then the LORD answered Job out of the whirlwind, and said,
JOB|38|2|Who is this that darkeneth counsel by words without knowledge?
JOB|38|3|Gird up now thy loins like a man; for I will demand of thee, and answer thou me.
JOB|38|4|Where wast thou when I laid the foundations of the earth? declare, if thou hast understanding.
JOB|38|5|Who hath laid the measures thereof, if thou knowest? or who hath stretched the line upon it?
JOB|38|6|Whereupon are the foundations thereof fastened? or who laid the corner stone thereof;
JOB|38|7|When the morning stars sang together, and all the sons of God shouted for joy?
JOB|38|8|Or who shut up the sea with doors, when it brake forth, as if it had issued out of the womb?
JOB|38|9|When I made the cloud the garment thereof, and thick darkness a swaddlingband for it,
JOB|38|10|And brake up for it my decreed place, and set bars and doors,
JOB|38|11|And said, Hitherto shalt thou come, but no further: and here shall thy proud waves be stayed?
JOB|38|12|Hast thou commanded the morning since thy days; and caused the dayspring to know his place;
JOB|38|13|That it might take hold of the ends of the earth, that the wicked might be shaken out of it?
JOB|38|14|It is turned as clay to the seal; and they stand as a garment.
JOB|38|15|And from the wicked their light is withholden, and the high arm shall be broken.
JOB|38|16|Hast thou entered into the springs of the sea? or hast thou walked in the search of the depth?
JOB|38|17|Have the gates of death been opened unto thee? or hast thou seen the doors of the shadow of death?
JOB|38|18|Hast thou perceived the breadth of the earth? declare if thou knowest it all.
JOB|38|19|Where is the way where light dwelleth? and as for darkness, where is the place thereof,
JOB|38|20|That thou shouldest take it to the bound thereof, and that thou shouldest know the paths to the house thereof?
JOB|38|21|Knowest thou it, because thou wast then born? or because the number of thy days is great?
JOB|38|22|Hast thou entered into the treasures of the snow? or hast thou seen the treasures of the hail,
JOB|38|23|Which I have reserved against the time of trouble, against the day of battle and war?
JOB|38|24|By what way is the light parted, which scattereth the east wind upon the earth?
JOB|38|25|Who hath divided a watercourse for the overflowing of waters, or a way for the lightning of thunder;
JOB|38|26|To cause it to rain on the earth, where no man is; on the wilderness, wherein there is no man;
JOB|38|27|To satisfy the desolate and waste ground; and to cause the bud of the tender herb to spring forth?
JOB|38|28|Hath the rain a father? or who hath begotten the drops of dew?
JOB|38|29|Out of whose womb came the ice? and the hoary frost of heaven, who hath gendered it?
JOB|38|30|The waters are hid as with a stone, and the face of the deep is frozen.
JOB|38|31|Canst thou bind the sweet influences of Pleiades, or loose the bands of Orion?
JOB|38|32|Canst thou bring forth Mazzaroth in his season? or canst thou guide Arcturus with his sons?
JOB|38|33|Knowest thou the ordinances of heaven? canst thou set the dominion thereof in the earth?
JOB|38|34|Canst thou lift up thy voice to the clouds, that abundance of waters may cover thee?
JOB|38|35|Canst thou send lightnings, that they may go and say unto thee, Here we are?
JOB|38|36|Who hath put wisdom in the inward parts? or who hath given understanding to the heart?
JOB|38|37|Who can number the clouds in wisdom? or who can stay the bottles of heaven,
JOB|38|38|When the dust groweth into hardness, and the clods cleave fast together?
JOB|38|39|Wilt thou hunt the prey for the lion? or fill the appetite of the young lions,
JOB|38|40|When they couch in their dens, and abide in the covert to lie in wait?
JOB|38|41|Who provideth for the raven his food? when his young ones cry unto God, they wander for lack of meat.
JOB|39|1|Knowest thou the time when the wild goats of the rock bring forth? or canst thou mark when the hinds do calve?
JOB|39|2|Canst thou number the months that they fulfil? or knowest thou the time when they bring forth?
JOB|39|3|They bow themselves, they bring forth their young ones, they cast out their sorrows.
JOB|39|4|Their young ones are in good liking, they grow up with corn; they go forth, and return not unto them.
JOB|39|5|Who hath sent out the wild ass free? or who hath loosed the bands of the wild ass?
JOB|39|6|Whose house I have made the wilderness, and the barren land his dwellings.
JOB|39|7|He scorneth the multitude of the city, neither regardeth he the crying of the driver.
JOB|39|8|The range of the mountains is his pasture, and he searcheth after every green thing.
JOB|39|9|Will the unicorn be willing to serve thee, or abide by thy crib?
JOB|39|10|Canst thou bind the unicorn with his band in the furrow? or will he harrow the valleys after thee?
JOB|39|11|Wilt thou trust him, because his strength is great? or wilt thou leave thy labour to him?
JOB|39|12|Wilt thou believe him, that he will bring home thy seed, and gather it into thy barn?
JOB|39|13|Gavest thou the goodly wings unto the peacocks? or wings and feathers unto the ostrich?
JOB|39|14|Which leaveth her eggs in the earth, and warmeth them in dust,
JOB|39|15|And forgetteth that the foot may crush them, or that the wild beast may break them.
JOB|39|16|She is hardened against her young ones, as though they were not her's: her labour is in vain without fear;
JOB|39|17|Because God hath deprived her of wisdom, neither hath he imparted to her understanding.
JOB|39|18|What time she lifteth up herself on high, she scorneth the horse and his rider.
JOB|39|19|Hast thou given the horse strength? hast thou clothed his neck with thunder?
JOB|39|20|Canst thou make him afraid as a grasshopper? the glory of his nostrils is terrible.
JOB|39|21|He paweth in the valley, and rejoiceth in his strength: he goeth on to meet the armed men.
JOB|39|22|He mocketh at fear, and is not affrighted; neither turneth he back from the sword.
JOB|39|23|The quiver rattleth against him, the glittering spear and the shield.
JOB|39|24|He swalloweth the ground with fierceness and rage: neither believeth he that it is the sound of the trumpet.
JOB|39|25|He saith among the trumpets, Ha, ha; and he smelleth the battle afar off, the thunder of the captains, and the shouting.
JOB|39|26|Doth the hawk fly by thy wisdom, and stretch her wings toward the south?
JOB|39|27|Doth the eagle mount up at thy command, and make her nest on high?
JOB|39|28|She dwelleth and abideth on the rock, upon the crag of the rock, and the strong place.
JOB|39|29|From thence she seeketh the prey, and her eyes behold afar off.
JOB|39|30|Her young ones also suck up blood: and where the slain are, there is she.
JOB|40|1|Moreover the LORD answered Job, and said,
JOB|40|2|Shall he that contendeth with the Almighty instruct him? he that reproveth God, let him answer it.
JOB|40|3|Then Job answered the LORD, and said,
JOB|40|4|Behold, I am vile; what shall I answer thee? I will lay mine hand upon my mouth.
JOB|40|5|Once have I spoken; but I will not answer: yea, twice; but I will proceed no further.
JOB|40|6|Then answered the LORD unto Job out of the whirlwind, and said,
JOB|40|7|Gird up thy loins now like a man: I will demand of thee, and declare thou unto me.
JOB|40|8|Wilt thou also disannul my judgment? wilt thou condemn me, that thou mayest be righteous?
JOB|40|9|Hast thou an arm like God? or canst thou thunder with a voice like him?
JOB|40|10|Deck thyself now with majesty and excellency; and array thyself with glory and beauty.
JOB|40|11|Cast abroad the rage of thy wrath: and behold every one that is proud, and abase him.
JOB|40|12|Look on every one that is proud, and bring him low; and tread down the wicked in their place.
JOB|40|13|Hide them in the dust together; and bind their faces in secret.
JOB|40|14|Then will I also confess unto thee that thine own right hand can save thee.
JOB|40|15|Behold now behemoth, which I made with thee; he eateth grass as an ox.
JOB|40|16|Lo now, his strength is in his loins, and his force is in the navel of his belly.
JOB|40|17|He moveth his tail like a cedar: the sinews of his stones are wrapped together.
JOB|40|18|His bones are as strong pieces of brass; his bones are like bars of iron.
JOB|40|19|He is the chief of the ways of God: he that made him can make his sword to approach unto him.
JOB|40|20|Surely the mountains bring him forth food, where all the beasts of the field play.
JOB|40|21|He lieth under the shady trees, in the covert of the reed, and fens.
JOB|40|22|The shady trees cover him with their shadow; the willows of the brook compass him about.
JOB|40|23|Behold, he drinketh up a river, and hasteth not: he trusteth that he can draw up Jordan into his mouth.
JOB|40|24|He taketh it with his eyes: his nose pierceth through snares.
JOB|41|1|Canst thou draw out leviathan with an hook? or his tongue with a cord which thou lettest down?
JOB|41|2|Canst thou put an hook into his nose? or bore his jaw through with a thorn?
JOB|41|3|Will he make many supplications unto thee? will he speak soft words unto thee?
JOB|41|4|Will he make a covenant with thee? wilt thou take him for a servant for ever?
JOB|41|5|Wilt thou play with him as with a bird? or wilt thou bind him for thy maidens?
JOB|41|6|Shall the companions make a banquet of him? shall they part him among the merchants?
JOB|41|7|Canst thou fill his skin with barbed irons? or his head with fish spears?
JOB|41|8|Lay thine hand upon him, remember the battle, do no more.
JOB|41|9|Behold, the hope of him is in vain: shall not one be cast down even at the sight of him?
JOB|41|10|None is so fierce that dare stir him up: who then is able to stand before me?
JOB|41|11|Who hath prevented me, that I should repay him? whatsoever is under the whole heaven is mine.
JOB|41|12|I will not conceal his parts, nor his power, nor his comely proportion.
JOB|41|13|Who can discover the face of his garment? or who can come to him with his double bridle?
JOB|41|14|Who can open the doors of his face? his teeth are terrible round about.
JOB|41|15|His scales are his pride, shut up together as with a close seal.
JOB|41|16|One is so near to another, that no air can come between them.
JOB|41|17|They are joined one to another, they stick together, that they cannot be sundered.
JOB|41|18|By his neesings a light doth shine, and his eyes are like the eyelids of the morning.
JOB|41|19|Out of his mouth go burning lamps, and sparks of fire leap out.
JOB|41|20|Out of his nostrils goeth smoke, as out of a seething pot or caldron.
JOB|41|21|His breath kindleth coals, and a flame goeth out of his mouth.
JOB|41|22|In his neck remaineth strength, and sorrow is turned into joy before him.
JOB|41|23|The flakes of his flesh are joined together: they are firm in themselves; they cannot be moved.
JOB|41|24|His heart is as firm as a stone; yea, as hard as a piece of the nether millstone.
JOB|41|25|When he raiseth up himself, the mighty are afraid: by reason of breakings they purify themselves.
JOB|41|26|The sword of him that layeth at him cannot hold: the spear, the dart, nor the habergeon.
JOB|41|27|He esteemeth iron as straw, and brass as rotten wood.
JOB|41|28|The arrow cannot make him flee: slingstones are turned with him into stubble.
JOB|41|29|Darts are counted as stubble: he laugheth at the shaking of a spear.
JOB|41|30|Sharp stones are under him: he spreadeth sharp pointed things upon the mire.
JOB|41|31|He maketh the deep to boil like a pot: he maketh the sea like a pot of ointment.
JOB|41|32|He maketh a path to shine after him; one would think the deep to be hoary.
JOB|41|33|Upon earth there is not his like, who is made without fear.
JOB|41|34|He beholdeth all high things: he is a king over all the children of pride.
JOB|42|1|Then Job answered the LORD, and said,
JOB|42|2|I know that thou canst do every thing, and that no thought can be withholden from thee.
JOB|42|3|Who is he that hideth counsel without knowledge? therefore have I uttered that I understood not; things too wonderful for me, which I knew not.
JOB|42|4|Hear, I beseech thee, and I will speak: I will demand of thee, and declare thou unto me.
JOB|42|5|I have heard of thee by the hearing of the ear: but now mine eye seeth thee.
JOB|42|6|Wherefore I abhor myself, and repent in dust and ashes.
JOB|42|7|And it was so, that after the LORD had spoken these words unto Job, the LORD said to Eliphaz the Temanite, My wrath is kindled against thee, and against thy two friends: for ye have not spoken of me the thing that is right, as my servant Job hath.
JOB|42|8|Therefore take unto you now seven bullocks and seven rams, and go to my servant Job, and offer up for yourselves a burnt offering; and my servant Job shall pray for you: for him will I accept: lest I deal with you after your folly, in that ye have not spoken of me the thing which is right, like my servant Job.
JOB|42|9|So Eliphaz the Temanite and Bildad the Shuhite and Zophar the Naamathite went, and did according as the LORD commanded them: the LORD also accepted Job.
JOB|42|10|And the LORD turned the captivity of Job, when he prayed for his friends: also the LORD gave Job twice as much as he had before.
JOB|42|11|Then came there unto him all his brethren, and all his sisters, and all they that had been of his acquaintance before, and did eat bread with him in his house: and they bemoaned him, and comforted him over all the evil that the LORD had brought upon him: every man also gave him a piece of money, and every one an earring of gold.
JOB|42|12|So the LORD blessed the latter end of Job more than his beginning: for he had fourteen thousand sheep, and six thousand camels, and a thousand yoke of oxen, and a thousand she asses.
JOB|42|13|He had also seven sons and three daughters.
JOB|42|14|And he called the name of the first, Jemima; and the name of the second, Kezia; and the name of the third, Kerenhappuch.
JOB|42|15|And in all the land were no women found so fair as the daughters of Job: and their father gave them inheritance among their brethren.
JOB|42|16|After this lived Job an hundred and forty years, and saw his sons, and his sons' sons, even four generations.
JOB|42|17|So Job died, being old and full of days.
