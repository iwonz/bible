JONAH|1|1|Et factum est verbum Domini ad Ionam filium Amathi dicens:
JONAH|1|2|" Surge et vade in Nineven civitatem grandem et praedica in ea, quia ascendit malitia eius coram me ".
JONAH|1|3|Et surrexit Ionas, ut fugeret in Tharsis a facie Domini; et descendit Ioppen et invenit navem euntem in Tharsis et dedit naulum eius et descendit in eam, ut iret cum eis in Tharsis a facie Domini.
JONAH|1|4|Dominus autem misit ventum magnum in mare, et facta est tempestas magna in mari, et navis periclitabatur conteri.
JONAH|1|5|Et timuerunt nautae et clamaverunt unusquisque ad deum suum et miserunt vasa, quae erant in navi, in mare, ut alleviaretur ab eis. Ionas autem descenderat ad interiora navis et, cum recubuisset, dormiebat sopore gravi.
JONAH|1|6|Et accessit ad eum gubernator et dixit ei: " Quid? Tu sopore deprimeris? Surge, invoca Deum tuum, si forte recogitet Deus de nobis, et non pereamus.
JONAH|1|7|Et dixit unusquisque ad collegam suum: " Venite, et mittamus sortes, ut sciamus quare hoc malum sit nobis ". Et miserunt sortes, et cecidit sors super Ionam.
JONAH|1|8|Et dixerunt ad eum: " Indica nobis cuius causa malum istud sit nobis. Quod est opus tuum, et unde venis? Quae terra tua, et ex quo populo es tu?.
JONAH|1|9|Et dixit ad eos: " Hebraeus ego sum et Dominum, Deum caeli, ego timeo, qui fecit mare et aridam ".
JONAH|1|10|Et timuerunt viri timore magno et dixerunt ad eum: " Quid hoc fecisti?. Cognoverant enim viri quod a facie Domini fugeret, quia indicaverat eis.
JONAH|1|11|Et dixerunt ad eum: " Quid faciemus tibi, ut conticescat mare a nobis?. Mare enim magis ac magis intumescebat.
JONAH|1|12|Et dixit ad eos: " Tollite me et mittite in mare, et cessabit mare a vobis; scio enim ego quoniam propter me tempestas haec grandis super vos.
JONAH|1|13|Et remigabant viri, ut reverterentur ad aridam; et non valebant, quia mare magis intumescebat super eos.
JONAH|1|14|Et clamaverunt ad Dominum et dixerunt: " Quaesumus, Domine, ne pereamus in anima viri istius, et ne des super nos sanguinem innocentem; quia tu, Domine, sicut voluisti, fecisti ".
JONAH|1|15|Et tulerunt Ionam et miserunt in mare; et stetit mare a fervore suo.
JONAH|1|16|Et timuerunt viri timore magno Dominum et immolaverunt hostias Domino et voverunt vota.
JONAH|2|1|Et praeparavit Dominus piscem grandem, ut deglutiret Ionam; et erat Ionas in ventre piscis tribus diebus et tribus noctibus.
JONAH|2|2|Et oravit Ionas ad Dominum Deum suum de ventre piscis
JONAH|2|3|et dixit: " Clamavi de tribulatione mea ad Dominum,et respondit mihi;de ventre inferi clamavi,et exaudisti vocem meam.
JONAH|2|4|Et proiecisti me in profundum in corde maris,et flumen circumdedit me;omnes gurgites tui et fluctus tuisuper me transierunt.
JONAH|2|5|Et ego dixi: "Abiectus suma conspectu oculorum tuorum;verumtamen rursus videbotemplum sanctum tuum".
JONAH|2|6|Circumdederunt me aquae usque ad guttur,abyssus vallavit me,iuncus alligatus est capiti meo.
JONAH|2|7|Ad extrema montium descendi,terrae vectes concluserunt me in aeternum,sed eduxisti de fovea vitam meam,Domine Deus meus.
JONAH|2|8|Cum angustiaretur in me anima mea,Domini recordatus sum,et venit ad te oratio mea,ad templum sanctum tuum.
JONAH|2|9|Qui colunt idola vana,pietatem suam derelinquunt;
JONAH|2|10|ego autem in voce laudisimmolabo tibi,quaecumque vovi, reddam;salus Domini est ".
JONAH|2|11|Et dixit Dominus pisci, et evomuit Ionam in aridam.
JONAH|3|1|Et factum est verbum Domini ad Ionam secundo dicens:
JONAH|3|2|" Surge, vade in Nineven civitatem magnam et praedica in ea praedicationem, quam ego loquor ad te ".
JONAH|3|3|Et surrexit Ionas et abiit in Nineven iuxta verbum Domini.Et Nineve erat civitas magna coram Deo, itinere trium dierum.
JONAH|3|4|Et coepit Ionas introire in civitatem itinere diei unius; et clamavit et dixit: " Adhuc quadraginta dies, et Nineve subvertetur ".
JONAH|3|5|Et crediderunt viri Ninevitae in Deo; et praedicaverunt ieiunium et vestiti sunt saccis a maiore usque ad minorem.
JONAH|3|6|Et pervenit verbum ad regem Nineve; et surrexit de solio suo et abiecit pallium suum a se et indutus est sacco et sedit in cinere.
JONAH|3|7|Et clamavit et dixit in Nineve decreto regis et principum eius dicens: " Homines et iumenta et boves et pecora non gustent quidquam nec pascantur et aquam non bibant;
JONAH|3|8|et operiantur saccis homines et iumenta et clament ad Deum in fortitudine, et convertatur vir a via sua mala et a violentia, quae est in manibus eorum.
JONAH|3|9|Quis scit si convertatur et ignoscat Deus et revertatur a furore irae suae, et non peribimus? ".
JONAH|3|10|Et vidit Deus opera eorum, quia conversi sunt de via sua mala; et misertus est Deus super malum, quod lo cutus fuerat ut faceret eis, etnon fecit.
JONAH|4|1|Et afflictus est Ionas afflictione magna et iratus est;
JONAH|4|2|et oravit ad Dominum et dixit: " Obsecro, Domine, numquid non hoc est verbum meum, cum adhuc essem in terra mea? Propter hoc praeoccupavi ut fugerem in Tharsis. Sciebam enim quia tu Deus clemens et misericors es, longanimis et multae miserationis et ignoscens super malitia.
JONAH|4|3|Et nunc, Domine, tolle, quaeso, animam meam a me, quia melior est mihi mors quam vita".
JONAH|4|4|Et dixit Dominus: " Putasne bene irasceris tu? ".
JONAH|4|5|Et egressus est Ionas de civitate et sedit contra orientem civitatis et fecit sibimet umbraculum ibi et sedebat subter illud in umbra, donec videret quid accideret in civitate.
JONAH|4|6|Et praeparavit Dominus Deus hederam, et ascendit super Ionam, ut esset umbra super caput eius et protegeret eum ab afflictione sua. Et laetatus est Ionas super hedera laetitia magna.
JONAH|4|7|Et paravit Deus vermem, cum surgeret aurora in crastinum, et percussit hederam, quae exaruit.
JONAH|4|8|Et, cum ortus fuisset sol, praecepit Deus vento orientali calido; et percussit sol super caput Ionae, et elanguit; et petivit animae suae, ut moreretur, et dixit: " Melius est mihi mori quam vivere "
JONAH|4|9|Et dixit Deus ad Ionam: " Putasne bene irasceris tu super hedera? ". Et dixit: " Bene irascor ego usque ad mortem ".
JONAH|4|10|Et dixit Dominus: " Tu doles super hederam, in qua non laborasti neque fecisti, ut cresceret, quae sub una nocte nata est et sub una nocte periit.
JONAH|4|11|Et ego non parcam Nineve civitati magnae, in qua sunt plus quam centum viginti milia hominum, qui nesciunt quid sit inter dexteram et sinistram suam, et iumenta multa? ".
