1THESS|1|1|保罗 、 西拉 、 提摩太 写信给 帖撒罗尼迦 在父上帝和主耶稣基督里的教会。愿恩惠、平安 归给你们！
1THESS|1|2|我们为你们众人常常感谢上帝，祷告的时候提到你们，
1THESS|1|3|在我们的父上帝面前，不住地记念你们因信心所做的工作，因爱心所受的劳苦，因盼望我们主耶稣基督所存的坚忍。
1THESS|1|4|上帝所爱的弟兄啊，我知道你们是蒙拣选的；
1THESS|1|5|因为我们的福音传到你们那里，不仅在言语，也在能力，也在圣灵和充足的确信。你们知道，我们在你们那里，为你们的缘故是怎样为人。
1THESS|1|6|你们成为效法我们，更效法主的人，因圣灵所激发的喜乐，在大患难中领受了真道，
1THESS|1|7|从此你们作了 马其顿 和 亚该亚 所有信主的人的榜样。
1THESS|1|8|因为主的道已经从你们那里传播出去，你们向上帝的信心不只在 马其顿 和 亚该亚 ，就是在各处也都传开了，所以不用我们说什么话。
1THESS|1|9|因为他们自己已经传讲我们是怎样进到你们那里，你们是怎样离弃偶像，归向上帝来服侍那又真又活的上帝，
1THESS|1|10|等候他儿子从天降临，就是上帝使他从死人中复活的那位救我们脱离将来愤怒的耶稣。
1THESS|2|1|弟兄们，你们自己知道我们来到你们那里并不是徒然的。
1THESS|2|2|我们从前在 腓立比 蒙难受辱，这是你们知道的，可是我们还是靠着上帝给我们的勇气，在强烈反对中把上帝的福音传给你们。
1THESS|2|3|我们的劝勉不是出于错误，也不是出于污秽，也不是用诡诈。
1THESS|2|4|但上帝既然认定我们经得起考验，把福音托付我们，我们就照着传讲，不是要讨人喜欢，而是要讨那考验我们的心的上帝喜欢。
1THESS|2|5|因为我们从来没有用过谄媚的话，这是你们知道的，也没有藏着贪心，这是上帝可以作证的。
1THESS|2|6|我们作为基督的使徒，虽然可以受人尊重，却没有向你们或向别人求荣耀，反而在你们当中心存温柔，如同母亲哺乳自己的孩子。
1THESS|2|7|
1THESS|2|8|既然我们这样爱你们，不但乐意将上帝的福音给你们，连自己的性命也乐意给你们，因为你们是我们所疼爱的。
1THESS|2|9|弟兄们，你们记念我们的辛苦劳碌，昼夜做工，传上帝的福音给你们，免得你们任何人受累。
1THESS|2|10|我们对你们信主的人是何等圣洁、正直、无可指责，这有你们作证，也有上帝作证。
1THESS|2|11|正如你们知道，我们待你们好像父亲待自己的儿女一样。
1THESS|2|12|我们劝勉你们，安慰你们，嘱咐你们，使你们行事对得起那召你们进他自己的国、得他荣耀的上帝。
1THESS|2|13|为此，我们也不断地感谢上帝，因为你们听见我们所传上帝的道的时候，你们领受了，不以为这是人的道，而以为这确实是上帝的道，而且在你们信主的人当中运行着。
1THESS|2|14|弟兄们，你们与 犹太 地区上帝的各教会，就是在基督耶稣里的各教会，有同样的遭遇，因为你们也受了同胞的迫害，像他们受了 犹太 人的迫害一样。
1THESS|2|15|这些 犹太 人不但杀了主耶稣和先知们，又把我们赶出去。他们令上帝不悦，且与众人为敌，
1THESS|2|16|阻挠我们传道给外邦人，使他们得救，以致常常恶贯满盈，但上帝的愤怒终于临到他们身上。
1THESS|2|17|弟兄们，我们被迫暂时与你们分离，身体离开，心却没有；我们极力想法子，渴望见你们的面。
1THESS|2|18|所以我们很想到你们那里去。我－ 保罗 有一两次要去，只是撒但阻挡了我们。
1THESS|2|19|当我们的主耶稣再来，我们站在他面前的时候，我们的盼望、喜乐和所夸的冠冕是什么呢？不正是你们吗？
1THESS|2|20|你们就是我们的荣耀和喜乐！
1THESS|3|1|既然我们不能再忍，就决定独自留在 雅典 ，
1THESS|3|2|于是差派我们在基督福音上作上帝同工的弟兄 提摩太 前去，在你们所信的道上坚固你们，劝勉你们，
1THESS|3|3|免得有人被这些患难动摇。因为你们自己知道，我们受患难原是命定的。
1THESS|3|4|我们在你们那里的时候，曾预先告诉你们，我们必受患难；你们知道，这果然发生了。
1THESS|3|5|为此，既然我不能再忍，就差派人去，要知道你们的信心如何，恐怕那诱惑人的果真诱惑了你们，以致我们的劳苦归于徒然。
1THESS|3|6|但是， 提摩太 刚从你们那里回来，将你们信心和爱心的好消息报给我们，又说你们常常记念我们，切切想见我们，如同我们想见你们一样。
1THESS|3|7|所以，弟兄们，我们在一切困苦患难中，因着你们的信心得到鼓励。
1THESS|3|8|如今你们若靠主站立得稳，我们就得生了。
1THESS|3|9|我们在上帝面前，因着你们满有喜乐。为这一切喜乐，我们能用怎样的感谢为你们报答上帝呢？
1THESS|3|10|我们昼夜切切祈求要见你们的面，来补足你们信心的不足。
1THESS|3|11|愿我们的父上帝自己和我们的主耶稣，为我们开路到你们那里去。
1THESS|3|12|又愿主使你们彼此相爱的心，和爱众人的心，都能增长，充足，如同我们爱你们一样，
1THESS|3|13|好坚固你们的心，使你们在我们的主耶稣同他众圣徒来临的时候，在我们父上帝面前，成为圣洁，无可指责。阿们！
1THESS|4|1|末了，弟兄们，我们靠着主耶稣求你们，劝你们，既然你们领受了我们的教导，知道该怎样行事为人，讨上帝的喜悦，其实你们也正这样行，我劝你们要更加努力。
1THESS|4|2|你们原知道，我们凭主耶稣传给你们什么命令。
1THESS|4|3|上帝的旨意就是要你们成为圣洁，远避淫行；
1THESS|4|4|要你们各人知道怎样用圣洁、尊贵控制自己的身体 ，
1THESS|4|5|不放纵私欲的邪情，像不认识上帝的外邦人。
1THESS|4|6|不准有人在这事上越轨，占他弟兄的便宜；因为这一类的事，主必报应，正如我预先对你们说过，又切切警告过你们的。
1THESS|4|7|上帝召我们本不是要我们沾染污秽，而是要我们圣洁。
1THESS|4|8|所以，那弃绝这教导的不是弃绝人，而是弃绝那把自己的圣灵赐给你们的上帝。
1THESS|4|9|有关弟兄间的手足之情，不用人写信给你们，因为你们自己蒙了上帝的教导要彼此相爱。
1THESS|4|10|你们向全 马其顿 的众弟兄固然是这样行，但我劝弟兄们要更加努力。
1THESS|4|11|要立志过安静的生活，管自己的事，亲手 做工，正如我们从前吩咐你们的，
1THESS|4|12|好使你们的行为能得外人的尊敬，同时也不依赖任何人。
1THESS|4|13|弟兄们，至于已睡了的人，我们不愿意你们不知道，恐怕你们忧伤，像那些没有指望的人一样。
1THESS|4|14|既然我们信耶稣死了，复活了，那些已经在耶稣里睡了的人，上帝也必将他们与耶稣一同带来。
1THESS|4|15|我们照主的话告诉你们一件事：我们这活着还存留到主来临的人，绝不会在那已经睡了的人之先。
1THESS|4|16|因为，召集令一发，天使长的呼声一叫，上帝的号角一吹，主必亲自从天降临；那在基督里死了的人必先复活，
1THESS|4|17|然后我们这些活着还存留的人必和他们一同被提到云里，在空中与主相会。这样，我们就要和主永远同在。
1THESS|4|18|所以，你们当用这些话彼此劝勉。
1THESS|5|1|弟兄们，关于那时候和日期，不用人写信给你们，
1THESS|5|2|因为你们自己明明知道，主的日子来到会像贼在夜间突然来到一样。
1THESS|5|3|人正说平安稳定的时候，灾祸忽然临到他们，如同阵痛临到怀胎的妇人一样，他们绝逃脱不了。
1THESS|5|4|弟兄们，你们并不在黑暗里，那日子不会像贼一样临到你们。
1THESS|5|5|你们都是光明之子，都是白昼之子；我们不属黑夜，也不属幽暗。
1THESS|5|6|所以，我们不要沉睡，像别人一样，总要警醒谨慎。
1THESS|5|7|因为睡了的人是在夜间睡，醉了的人是在夜间醉。
1THESS|5|8|但既然我们属于白昼，就应当谨慎，把信和爱当作护心镜遮胸，把得救的盼望当作头盔戴上。
1THESS|5|9|因为上帝不是预定我们受惩罚，而是预定我们藉着我们的主耶稣基督得救。
1THESS|5|10|他替我们死，让我们无论醒着、睡着，都与他同活。
1THESS|5|11|所以，你们该彼此劝勉，互相造就，正如你们素常做的。
1THESS|5|12|弟兄们，我们劝你们要敬重那些在你们中间劳苦的，就是在主里面督导你们、劝戒你们的人。
1THESS|5|13|又因他们所做的工作，要以爱心格外尊重他们。你们也要彼此和睦。
1THESS|5|14|弟兄们，我们劝你们，要警戒不守规矩的人，勉励灰心的人，扶助软弱的人，对众人要有耐心。
1THESS|5|15|你们要谨慎，无论是谁都不要以恶报恶，彼此间和对众人都要追求做好事。
1THESS|5|16|要常常喜乐，
1THESS|5|17|不住地祷告，
1THESS|5|18|凡事谢恩，因为这是上帝在基督耶稣里向你们所定的旨意。
1THESS|5|19|不要熄灭圣灵；
1THESS|5|20|不要藐视先知的讲论。
1THESS|5|21|但凡事要察验：美善的事要持守，
1THESS|5|22|各样恶事要禁戒。
1THESS|5|23|愿赐平安 的上帝亲自使你们完全成圣！愿你们的灵、魂、体得蒙保守，在我们的主耶稣基督来临的时候，完全无可指责。
1THESS|5|24|那召你们的本是信实的，他必成就这事。
1THESS|5|25|弟兄们，请也为 我们祷告。
1THESS|5|26|用圣洁的吻向众弟兄问安。
1THESS|5|27|我指着主嘱咐你们，要把这信宣读给众弟兄听。
1THESS|5|28|愿我们的主耶稣基督的恩惠与你们同在！
