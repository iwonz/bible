NUM|1|1|Locutusque est Dominus ad Moysen in deserto Sinai in ta bernaculo conventus, prima die mensis secundi, anno altero egressionis eorum ex Aegypto, dicens:
NUM|1|2|" Tollite summam universae congregationis filiorum Israel per cognationes et domos suas et nomina singulorum, quidquid sexus est masculini
NUM|1|3|a vicesimo anno et supra omnium ex Israel, qui possunt ad bella procedere, et numerabitis eos per turmas suas, tu et Aaron.
NUM|1|4|Eritque vobiscum vir per tribum, princeps domus patrum suorum,
NUM|1|5|quorum ista sunt nomina: de Ruben Elisur filius Sedeur;
NUM|1|6|de Simeon Salamiel filius Surisaddai;
NUM|1|7|de Iuda Naasson filius Aminadab;
NUM|1|8|de Issachar Nathanael filius Suar;
NUM|1|9|de Zabulon Eliab filius Helon.
NUM|1|10|Filiorum autem Ioseph: de Ephraim Elisama filius Ammiud; de Manasse Gamaliel filius Phadassur.
NUM|1|11|De Beniamin Abidan filius Gedeonis;
NUM|1|12|de Dan Ahiezer filius Ammisaddai;
NUM|1|13|de Aser Phegiel filius Ochran;
NUM|1|14|de Gad Eliasaph filius Deuel;
NUM|1|15|de Nephthali Ahira filius Enan ".
NUM|1|16|Hi viri nobilissimi congregationis principes tribuum patrum suorum et capita milium Israel.
NUM|1|17|Quos tulerunt Moyses et Aaron nominatim designatos
NUM|1|18|et omnem congregationem congregaverunt primo die mensis secundi recensentes eos per cognationes et domos patrum eorum, per nomina singulorum a vicesimo anno et supra per capita,
NUM|1|19|sicut praeceperat Dominus Moysi. Numeratique sunt in deserto Sinai.
NUM|1|20|De Ruben primogenito Israelis generationes per familias ac domos patrum suorum, per nomina capitum singulorum omne quod sexus est masculini a vicesimo anno et supra procedentium ad bellum.
NUM|1|21|Recensiti tribus Ruben quadraginta sex milia quingenti.
NUM|1|22|De filiis Simeon generationes per familias ac domos cognationum suarum recensiti sunt per nomina et capita singulorum omne quod sexus est masculini a vicesimo anno et supra procedentium ad bellum.
NUM|1|23|Recensiti tribus Simeon quinquaginta novem milia trecenti.
NUM|1|24|De filiis Gad generationes per familias ac domos cognationum suarum recensiti sunt per nomina singulorum a viginti annis et supra omnes, qui ad bella procederent,
NUM|1|25|quadraginta quinque milia sescenti quinquaginta.
NUM|1|26|De filiis Iudae generationes per familias ac domos cognationum suarum per nomina singulorum a vicesimo anno et supra omnes, qui poterant ad bella procedere,
NUM|1|27|recensiti sunt septuaginta quattuor milia sescenti.
NUM|1|28|De filiis Issachar generationes per familias ac domos cognationum suarum per nomina singulorum a vicesimo anno et supra omnes, qui ad bella procederent,
NUM|1|29|recensiti sunt quinquaginta quattuor milia quadringenti.
NUM|1|30|De filiis Zabulon generationes per familias ac domos cognationum suarum recensiti sunt per nomina singulorum a vicesimo anno et supra omnes, qui poterant ad bella procedere,
NUM|1|31|quinquaginta septem milia quadringenti.
NUM|1|32|De filiis Ioseph filiorum Ephraim generationes per familias ac domos cognationum suarum recensiti sunt per nomina singulorum a vicesimo anno et supra omnes, qui poterant ad bella procedere,
NUM|1|33|quadraginta milia quingenti.
NUM|1|34|Porro filiorum Manasse generationes per familias ac domos cognationum suarum recensiti sunt per nomina singulorum a viginti annis et supra omnes, qui poterant ad bella procedere,
NUM|1|35|triginta duo milia ducenti.
NUM|1|36|De filiis Beniamin generationes per familias ac domos cognationum suarum recensiti sunt nominibus singulorum a vicesimo anno et supra omnes, qui poterant ad bella procedere,
NUM|1|37|triginta quinque milia quadringenti.
NUM|1|38|De filiis Dan generationes per familias ac domos cognationum suarum recensiti sunt nominibus singulorum a vicesimo anno et supra omnes, qui poterant ad bella procedere,
NUM|1|39|sexaginta duo milia septingenti.
NUM|1|40|De filiis Aser generationes per familias ac domos cognationum suarum recensiti sunt per nomina singulorum a vicesimo anno et supra omnes, qui poterant ad bella procedere,
NUM|1|41|quadraginta milia et mille quingenti.
NUM|1|42|De filiis Nephthali generationes per familias ac domos cognationum suarum recensiti sunt nominibus singulorum a vicesimo anno et supra omnes, qui poterant ad bella procedere,
NUM|1|43|quinquaginta tria milia quadringenti.
NUM|1|44|Hi sunt quos numeraverunt Moyses et Aaron et duodecim principes Israel, singuli per domos patrum suorum.
NUM|1|45|Fueruntque omnis numerus filiorum Israel per domos patrum suorum a vicesimo anno et supra, qui poterant ad bella procedere,
NUM|1|46|sescenta tria milia virorum quingenti quinquaginta.
NUM|1|47|Levitae autem in tribu patrum suorum non sunt numerati cum eis.
NUM|1|48|Locutusque est Dominus ad Moysen dicens:
NUM|1|49|" Tribum Levi noli numerare neque pones summam eorum cum filiis Israel,
NUM|1|50|sed constitue eos super habitaculum testimonii et cuncta vasa eius et quidquid ad caeremonias pertinet. Ipsi portabunt habitaculum et omnia utensilia eius et erunt in ministerio ac per gyrum habitaculi metabuntur.
NUM|1|51|Cum proficiscendum fuerit, deponent Levitae habitaculum; cum castrametandum, erigent; quisquis externorum accesserit, occidetur.
NUM|1|52|Metabuntur autem castra filii Israel, unusquisque per turmas et cuneos atque exercitum suum.
NUM|1|53|Porro Levitae per gyrum habitaculi testimonii figent tentoria, ne fiat indignatio super congregationem filiorum Israel, et excubabunt in custodiis habitaculi testimonii ".
NUM|1|54|Fecerunt ergo filii Israel iuxta omnia, quae praeceperat Dominus Moysi.
NUM|2|1|Locutusque est Dominus ad Moysen et Aaron dicens:
NUM|2|2|" Singuli per turmas, signa atque vexilla et domos patrum suorum castrametabuntur filii Israel per gyrum tabernaculi conventus.
NUM|2|3|Ad orientem Iudas figet tentoria per turmas exercitus sui, fuitque princeps filiorum eius Naasson filius Aminadab;
NUM|2|4|et eius summa pugnantium septuaginta quattuor milia sescenti.
NUM|2|5|Iuxta eum castrametabuntur de tribu Issachar, quorum princeps fuit Nathanael filius Suar;
NUM|2|6|et omnis numerus pugnatorum eius quinquaginta quattuor milia quadringenti.
NUM|2|7|In tribu Zabulon princeps fuit Eliab filius Helon;
NUM|2|8|et numerus exercitus pugnatorum eius quinquaginta septem milia quadringenti.
NUM|2|9|Universi, qui in castris Iudae annumerati sunt, fuerunt centum octoginta sex milia quadringenti, et per turmas suas primi egredientur.
NUM|2|10|Vexillum castrorum Ruben ad meridianam plagam erit, secundum exercitus eorum; princeps Elisur filius Sedeur;
NUM|2|11|et cunctus exercitus pugnatorum eius, qui numerati sunt, quadraginta sex milia quingenti.
NUM|2|12|Iuxta eum castrametabuntur de tribu Simeon, quorum princeps fuit Salamiel filius Surisaddai;
NUM|2|13|et cunctus exercitus pugnatorum eius, qui numerati sunt, quinquaginta novem milia trecenti.
NUM|2|14|In tribu Gad princeps fuit Eliasaph filius Deuel;
NUM|2|15|et cunctus exercitus pugnatorum eius, qui numerati sunt, quadraginta quinque milia sescenti quinquaginta.
NUM|2|16|Omnes, qui recensiti sunt in castris Ruben, centum quinquaginta milia et mille quadringenti quinquaginta, per turmas suas in secundo loco proficiscentur.
NUM|2|17|Levabitur deinde tabernaculum conventus, castra Levitarum in medio castrorum, quomodo erigetur ita et deponetur; singuli per loca et vexilla sua proficiscentur.
NUM|2|18|Ad occidentalem plagam erit vexillum castrorum filiorum Ephraim per turmas suas, quorum princeps fuit Elisama filius Ammiud;
NUM|2|19|cunctus exercitus pugnatorum eius, qui numerati sunt, quadraginta milia quingenti.
NUM|2|20|Et cum eis tribus filiorum Manasse, quorum princeps fuit Gamaliel filius Phadassur;
NUM|2|21|cunctusque exercitus pugnatorum eius, qui numerati sunt, triginta duo milia ducenti.
NUM|2|22|In tribu filiorum Beniamin princeps fuit Abidan filius Gedeonis;
NUM|2|23|et cunctus exercitus pugnatorum eius, qui recensiti sunt, triginta quinque milia quadringenti.
NUM|2|24|Omnes, qui numerati sunt in castris Ephraim, centum octo milia centum, per turmas suas tertii proficiscentur.
NUM|2|25|Ad aquilonis partem stabit vexillum castrorum filiorum Dan secundum exercitus suos, quorum princeps fuit Ahiezer filius Ammisaddai;
NUM|2|26|cunctus exercitus pugnatorum eius, qui numerati sunt, sexaginta duo milia septingenti.
NUM|2|27|Iuxta eum figet tentoria tribus Aser, quorum princeps fuit Phegiel filius Ochran;
NUM|2|28|cunctus exercitus pugnatorum eius, qui numerati sunt, quadraginta milia et mille quingenti.
NUM|2|29|De tribu filiorum Nephthali princeps fuit Ahira filius Enan;
NUM|2|30|cunctus exercitus pugnatorum eius quinquaginta tria milia quadringenti.
NUM|2|31|Omnes, qui numerati sunt in castris Dan, fuerunt centum quinquaginta septem milia sescenti, et novissimi proficiscentur secundum vexilla sua ".
NUM|2|32|Hic numerus filiorum Israel, per domos patrum suorum omnes recensiti secundum exercitus suos, sescenta tria milia quingenti quinquaginta.
NUM|2|33|Levitae autem non sunt numerati inter filios Israel; sic enim praeceperat Dominus Moysi.
NUM|2|34|Feceruntque filii Israel iuxta omnia, quae mandaverat Dominus: castrametati sunt per vexilla sua et profecti per tribus ad domos patrum suorum.
NUM|3|1|Hae sunt generationes Aaron et Moysi in die, qua locutus est Dominus ad Moysen in monte Sinai.
NUM|3|2|Et haec nomina filiorum Aaron: primogenitus eius Nadab, deinde Abiu et Eleazar et Ithamar.
NUM|3|3|Haec nomina filiorum Aaron sacerdotum, qui uncti sunt et quorum repletae manus, ut sacerdotio fungerentur.
NUM|3|4|Mortui sunt enim Nadab et Abiu, cum offerrent ignem alienum in conspectu Domini in deserto Sinai, absque liberis; functique sunt sacerdotio Eleazar et Ithamar coram Aaron patre suo.
NUM|3|5|Locutusque est Dominus ad Moysen dicens:
NUM|3|6|" Applica tribum Levi et fac stare in conspectu Aaron sacerdotis, ut ministrent ei
NUM|3|7|et observent, quidquid ad eum pertinet et ad totam congregationem coram tabernaculo conventus, servientes in ministerio habitaculi,
NUM|3|8|et custodiant vasa tabernaculi conventus explentes officia filiorum Israel, servientes in ministerio habitaculi.
NUM|3|9|Dabisque dono Levitas Aaron et filiis eius, quibus traditi sunt a filiis Israel;
NUM|3|10|Aaron autem et filios eius constitues super cultum sacerdotii. Externus, qui ad ministrandum accesserit, morietur ".
NUM|3|11|Locutusque est Dominus ad Moysen dicens:
NUM|3|12|" Ecce ego tuli Levitas a filiis Israel pro omni primogenito, qui aperit vulvam in filiis Israel; eruntque Levitae mei.
NUM|3|13|Meum est enim omne primogenitum: ex quo percussi omnes primogenitos in terra Aegypti, sanctificavi mihi, quidquid primum nascitur in Israel ab homine usque ad pecus; mei sunt. Ego Dominus ".
NUM|3|14|Locutusque est Dominus ad Moysen in deserto Sinai dicens:
NUM|3|15|" Numera filios Levi per domos patrum suorum et familias omnem masculum ab uno mense et supra ".
NUM|3|16|Numeravit eos Moyses, ut praeceperat Dominus,
NUM|3|17|et inventi sunt filii Levi per nomina sua Gerson et Caath et Merari.
NUM|3|18|Haec sunt nomina filiorum Gerson secundum familias suas: Lobni et Semei;
NUM|3|19|filii Caath secundum familias suas: Amram et Isaar, Hebron et Oziel;
NUM|3|20|filii Merari secundum familias suas: Moholi et Musi. Hae sunt familiae Levi per domos patrum suorum.
NUM|3|21|De Gerson fuere familiae duae Lobnitica et Semeitica,
NUM|3|22|quarum numeratus est omnis populus sexus masculini ab uno mense et supra septem milia quingenti.
NUM|3|23|Hi post habitaculum metabantur ad occidentem
NUM|3|24|sub principe Eliasaph filio Lael;
NUM|3|25|et habebant excubias in tabernaculo conventus, ipsum habitaculum et tabernaculum, operimentum eius, velum, quod trahitur ante fores tabernaculi conventus,
NUM|3|26|et cortinas atrii, velum quoque, quod appenditur in introitu atrii, quod est circa habitaculum et circa altare, et funes ad omne opus eius.
NUM|3|27|Caath habet familias: Amramitas et Isaaritas et Hebronitas et Ozielitas; hae sunt familiae Caathitarum.
NUM|3|28|Omnes generis masculini ab uno mense et supra octo milia sescenti habebant excubias sanctuarii.
NUM|3|29|Familiae filiorum Caath castrametabantur ad latus habitaculi ad meridianam plagam,
NUM|3|30|princepsque eorum erat Elisaphan filius Oziel.
NUM|3|31|Et custodiebant arcam mensamque et candelabrum, altaria et vasa sanctuarii, in quibus ministratur, et velum cunctamque huiuscemodi supellectilem.
NUM|3|32|Princeps autem principum Levitarum Eleazar filius Aaron sacerdotis erat super excubitores custodiae sanctuarii.
NUM|3|33|At vero de Merari erant familiae Moholitae et Musitae.
NUM|3|34|Omnes generis masculini ab uno mense et supra sex milia ducenti;
NUM|3|35|princeps familiarum Merari Suriel filius Abihail. In plaga septentrionali ad latus habitaculi castrametabantur;
NUM|3|36|erant sub custodia eorum tabulae habitaculi et vectes et columnae ac bases earum et cuncta vasa eius et omnia, quae ad cultum huiuscemodi pertinent,
NUM|3|37|columnaeque atrii per circuitum cum basibus suis et paxilli cum funibus.
NUM|3|38|Castrametabantur ante habitaculum, ad orientalem plagam ante tabernaculum conventus ad orientem, Moyses et Aaron cum filiis suis habentes custodiam sanctuarii in medio filiorum Israel. Quisquis alienus accesserit, morietur.
NUM|3|39|Omnes Levitae, quos numeravit Moyses iuxta praeceptum Domini per familias suas in genere masculino a mense uno et supra, fuerunt viginti duo milia.
NUM|3|40|Et ait Dominus ad Moysen: " Numera omnes primogenitos sexus masculini de filiis Israel ab uno mense et supra et habebis summam eorum;
NUM|3|41|tollesque Levitas mihi pro omni primogenito filiorum Israel ­ ego sum Dominus ­ et pecora eorum pro universis primogenitis pecorum filiorum Israel ".
NUM|3|42|Recensuit Moyses, sicut praeceperat Dominus, omnes primogenitos filiorum Israel,
NUM|3|43|et fuerunt omnes masculi per nomina sua a mense uno et supra viginti duo milia ducenti septuaginta tres.
NUM|3|44|Locutusque est Dominus ad Moysen dicens:
NUM|3|45|" Tolle Levitas pro omnibus primogenitis filiorum Israel et pecora Levitarum pro pecoribus corum; eruntque Levitae mei. Ego sum Dominus.
NUM|3|46|In pretio autem ducentorum septuaginta trium, qui excedunt numerum Levitarum de primogenitis filiorum Israel,
NUM|3|47|accipies quinque siclos per singula capita, ad mensuram sanctuarii. Siclus habet viginti obolos.
NUM|3|48|Dabisque pecuniam Aaron et filiis eius pretium eorum, qui supra sunt ".
NUM|3|49|Tulit igitur Moyses pecuniam eorum, qui excesserant numerum eorum, qui redempti erant a Levitis;
NUM|3|50|a primogenitis filiorum Israel tulit pecuniam mille trecentorum sexaginta quinque siclorum iuxta pondus sanctuarii.
NUM|3|51|Et dedit eam Aaron et filiis eius iuxta verbum, quod praeceperat sibi Dominus.
NUM|4|1|Locutusque est Dominus ad Moysen et Aaron dicens:
NUM|4|2|" Tolle summam filiorum Caath de medio Levitarum per familias et domos suas
NUM|4|3|a tricesimo anno et supra usque ad quinquagesimum annum omnium, qui ingrediuntur, ut stent et ministrent in tabernaculo conventus.
NUM|4|4|Hic est cultus filiorum Caath in tabernaculo conventus: sanctum sanctorum.
NUM|4|5|Ingredientur Aaron et filii eius, quando movenda sunt castra, et deponent velum, quod pendet ante fores, involventque eo arcam testimonii;
NUM|4|6|et operient rursum velamine pellium delphini extendentque desuper pallium totum hyacinthinum et inducent vectes.
NUM|4|7|Mensam quoque propositionis involvent hyacinthino pallio et ponent cum ea acetabula et phialas, cyathos et crateras ad liba fundenda; panes semper in ea erunt.
NUM|4|8|Extendentque desuper pallium coccineum, quod rursum operient velamento pellium delphini et inducent vectes.
NUM|4|9|Sument et pallium hyacinthinum, quo operient candelabrum cum lucernis et forcipibus suis et emunctoriis et cunctis vasis olei, quae ad concinnandas lucernas necessaria sunt;
NUM|4|10|et super omnia ponent operimentum pellium delphini et ponent super feretrum.
NUM|4|11|Nec non et altare aureum involvent hyacinthino vestimento et extendent desuper operimentum pellium delphini et inducent vectes.
NUM|4|12|Omnia vasa, quibus ministratur in sanctuario, involvent hyacinthino pallio; et extendent desuper operimentum pellium delphini ponentque super feretrum.
NUM|4|13|Sed et altare mundabunt cinere et involvent illud purpureo vestimento;
NUM|4|14|ponentque super illud omnia vasa, quibus in ministerio eius utuntur, id est ignium receptacula, fuscinulas ac vatilla et pateras. Cuncta vasa altaris operient simul velamine pellium delphini et inducent vectes.
NUM|4|15|Cumque involverint Aaron et filii eius sanctuarium et omnia vasa eius in commotione castrorum, tunc intrabunt filii Caath, ut portent involuta, et non tangent sanctuarium, ne moriantur. Ista sunt onera filiorum Caath in tabernaculo conventus.
NUM|4|16|Ad curam Eleazari filii Aaron sacerdotis pertinet oleum ad concinnandas lucernas et gratissimum incensum et oblatio, quae semper offertur, et oleum unctionis et quidquid ad cultum habitaculi pertinet omniumque vasorum, quae in sanctuario sunt ".
NUM|4|17|Locutusque est Dominus ad Moysen et Aaron dicens:
NUM|4|18|" Nolite perdere populum Caath de medio Levitarum,
NUM|4|19|sed hoc facite eis, ut vivant et non moriantur, quando appropinquant ad sancta sanctorum: Aaron et filii eius intrabunt ipsique disponent opera singulorum et divident quid portare quis debeat.
NUM|4|20|Non intrabunt ad videndum, nec puncto quidem, sanctuarium; alioquin morientur ".
NUM|4|21|Locutusque est Dominus ad Moysen dicens:
NUM|4|22|" Tolle summam etiam filiorum Gerson per domos ac familias et cognationes suas;
NUM|4|23|a triginta annis et supra usque ad annos quinquaginta numera omnes, qui ingrediuntur et ministrant in tabernaculo conventus.
NUM|4|24|Hoc est officium familiarum Gersonitarum,
NUM|4|25|ut portent cortinas habitaculi, tabernaculum conventus, operimentum eius et super illud velamen delphini velumque, quod pendet in introitu tabernaculi conventus,
NUM|4|26|cortinas atrii et velum in introitu atrii, quod est circa habitaculum et altare, funiculos et vasa ministerii, omnia, quae facta sunt, ut eis laborent.
NUM|4|27|Iubente Aaron et filiis eius, portabunt filii Gerson, et scient singuli cui debeant oneri mancipari.
NUM|4|28|Hic est cultus familiarum Gersonitarum in tabernaculo conventus; eruntque sub manu Ithamar filii Aaron sacerdotis.
NUM|4|29|Filios quoque Merari per familias et domos patrum suorum recensebis
NUM|4|30|a triginta annis et supra usque ad annos quinquaginta, omnes, qui ingrediuntur ad officium ministerii sui et cultum tabernaculi conventus.
NUM|4|31|Haec sunt onera eorum: portabunt tabulas habitaculi et vectes eius, columnas ac bases earum,
NUM|4|32|columnas quoque atrii per circuitum cum basibus et paxillis et funibus suis; omnia vasa et supellectilem ad numerum accipient sicque portabunt.
NUM|4|33|Hoc est officium familiarum Meraritarum et ministerium in tabernaculo conventus; eruntque sub manu Ithamar filii Aaron sacerdotis ".
NUM|4|34|Recensuerunt igitur Moyses et Aaron et principes synagogae filios Caath per cognationes et domos patrum suorum
NUM|4|35|a triginta annis et supra usque ad annum quinquagesimum, omnes, qui ingrediuntur ad ministerium tabernaculi conventus;
NUM|4|36|et inventi sunt duo milia septingenti quinquaginta.
NUM|4|37|Hic est numerus familiarum Caath, qui ministrant in tabernaculo conventus: hos numeravit Moyses et Aaron iuxta sermonem Domini per manum Moysi.
NUM|4|38|Numerati sunt et filii Gerson per cognationes et domos patrum suorum
NUM|4|39|a triginta annis et supra usque ad quinquagesimum annum, omnes, qui ingrediuntur, ut ministrent in tabernaculo conventus;
NUM|4|40|et inventi sunt secundum familias et domus patrum suorum duo milia sescenti triginta.
NUM|4|41|Hic est numerus Gersonitarum, omnes, qui ministrant in tabernaculo conventus, quos numeraverunt Moy ses et Aaron iuxta verbum Domini.
NUM|4|42|Numeratae sunt et familiae filiorum Merari per cognationes et domos patrum suorum
NUM|4|43|a triginta annis et supra usque ad annum quinquagesimum, omnes, qui ingrediuntur ad explendos ritus tabernaculi conventus;
NUM|4|44|et inventi sunt tria milia ducenti.
NUM|4|45|Hic est numerus familiarum filiorum Merari, quos recensuerunt Moyses et Aaron iuxta imperium Domini per manum Moysi.
NUM|4|46|Omnes, qui recensiti sunt de Levitis et quos recenseri fecit ad nomen Moyses et Aaron et principes Israel per cognationes et domos patrum suorum
NUM|4|47|a triginta annis et supra usque ad annum quinquagesimum ingredientes ad ministerium tabernaculi et onera portanda in tabernaculo conventus,
NUM|4|48|fuerunt simul octo milia quingenti octoginta. 49 Iuxta verbum Domini per manum Moysi recensuit eos unumquemque iuxta officium et onera sua, sicut praeceperat ei Dominus.
NUM|5|1|Locutusque est Dominus ad Moysen dicens:
NUM|5|2|" Praecipe filiis Israel, ut eiciant de castris omnem leprosum et qui semine fluit pollutusque est super mortuo.
NUM|5|3|Tam masculum quam feminam eicite de castris, ne contaminent ea, cum habitaverim cum eis ".
NUM|5|4|Feceruntque ita filii Israel et eiecerunt eos extra castra, sicut locutus erat Dominus Moysi.
NUM|5|5|Locutusque est Dominus ad Moysen dicens:
NUM|5|6|" Loquere ad filios Israel: Vir sive mulier, cum fecerint ex omnibus peccatis, quae solent hominibus accidere, et fraude transgressi fuerint mandatum Domini, ille homo reus erit;
NUM|5|7|et confitebuntur peccatum suum et reddent ipsum caput quintamque partem desuper ei, in quem peccaverint.
NUM|5|8|Sin autem non fuerit qui recipiat, dabunt Domino, et erit sacerdotis, praeter arietem, qui offertur pro expiatione, ut sit placabilis hostia.
NUM|5|9|Omnis quoque praelibatio rerum sacrarum, quas offerunt filii Israel, ad sacerdotem pertinet;
NUM|5|10|et, quidquid in sanctuarium offertur a singulis et traditur manibus sacerdotis, ipsius erit ".
NUM|5|11|Locutusque est Dominus ad Moysen dicens:
NUM|5|12|" Loquere ad filios Israel et dices ad eos: Vir, cuius uxor erraverit maritumque decipiens
NUM|5|13|dormierit cum altero viro, et hoc maritus deprehendere non quiverit, sed latet quod impuram se reddiderit et testibus argui non potest, quia non est inventa in stupro,
NUM|5|14|si spiritus zelotypiae concitaverit virum contra uxorem suam, quae vel polluta est vel falsa suspicione appetitur,
NUM|5|15|adducet eam ad sacerdotem et offeret oblationem pro illa decimam partem ephi farinae hordeaceae. Non fundet super eam oleum nec imponet tus, quia sacrificium zelotypiae est et oblatio investigans adulterium.
NUM|5|16|Afferet igitur eam sacerdos et statuet coram Domino;
NUM|5|17|assumetque aquam sanctam in vase fictili et pauxillum terrae de pavimento habitaculi mittet in eam.
NUM|5|18|Cumque posuerit sacerdos mulierem in conspectu Domini, discooperiet caput eius et ponet super manus illius sacrificium recordationis, oblationem zelotypiae; ipse autem tenebit aquas amarissimas, in quibus cum exsecratione maledicta congessit.
NUM|5|19|Adiurabitque eam et dicet: "Si non dormivit vir alienus tecum, et si non declinasti a viro tuo et non polluta es, deserto mariti toro, non te nocebunt aquae istae amarissimae, in quas maledicta congessi.
NUM|5|20|Sin autem declinasti a viro tuo atque polluta es et concubuisti cum altero viro",
NUM|5|21|adiurabit eam sacerdos iuramento maledictionis: "Det te Dominus in maledictionem, iuramentum in medio populi tui; putrescere faciat femur tuum, et tumens uterus tuus disrumpatur;
NUM|5|22|ingrediantur aquae maledictae in ventrem tuum, et utero tumescente putrescat femur!". Et respondebit mulier: "Amen, amen".
NUM|5|23|Scribetque sacerdos in libello ista maledicta et delebit ea aquis amarissimis
NUM|5|24|et dabit ei bibere aquas amaras, in quas maledicta congessit, et ingredientur in eam aquae maledictionis, quae amarae fient;
NUM|5|25|tollet sacerdos de manu eius sacrificium zelotypiae et agitabit illud coram Domino imponetque illud super altare;
NUM|5|26|pugillum sacrificii tollat de eo, quod offertur in memoriale, et incendat super altare; et deinde potum det mulieri aquas amarissimas.
NUM|5|27|Quas cum biberit, si polluta est et, contempto viro, adulterii rea, pertransibunt eam aquae maledictionis et, inflato ventre, computrescet femur; eritque mulier in maledictionem omni populo eius.
NUM|5|28|Quod si polluta non fuerit sed munda, erit innoxia et faciet liberos ".
NUM|5|29|Ista est lex zelotypiae, si declinaverit mulier a viro suo et si polluta fuerit,
NUM|5|30|maritusque zelotypiae spiritu concitatus adduxerit eam in conspectu Domini, et fecerit ei sacerdos iuxta omnia, quae scripta sunt;
NUM|5|31|maritus absque culpa erit, et illa recipiet iniquitatem suam.
NUM|6|1|Locutusque est Dominus ad Moysen dicens:
NUM|6|2|" Loquere ad filios Israel et dices ad eos: Vir sive mulier cum fecerint votum, ut sanctificentur et se voluerint Domino consecrare,
NUM|6|3|a vino et omni quod inebriare potest abstinebunt; acetum ex vino et ex qualibet alia potione et, quidquid de uva exprimitur, non bibent; uvas recentes siccasque non comedent
NUM|6|4|cunctis diebus, quibus ex voto Domino consecrantur: quidquid ex vinea esse potest ab uva acerba usque ad pellicula non comedent.
NUM|6|5|Omni tempore separationis suae novacula non transibit per caput eius usque ad completum tempus, quo Domino consecratur; sanctus erit crescente caesarie capitis eius.
NUM|6|6|Omni tempore consecrationis suae ad mortuum non ingredietur;
NUM|6|7|nec super patris quidem et matris et fratris sororisque funere contaminabitur, quia consecratio Dei sui super caput eius est.
NUM|6|8|Omnibus diebus separationis suae sanctus erit Domino.
NUM|6|9|Sin autem mortuus fuerit subito quispiam coram eo, polluetur caput consecrationis eius; quod radet ilico in eadem die purgationis suae, id est die septima.
NUM|6|10|In octava autem die offeret duos turtures vel duos pullos columbae sacerdoti in introitu tabernaculi conventus,
NUM|6|11|facietque sacerdos unum pro peccato et alterum in holocaustum et expiabit pro eo, quia peccavit super mortuo, sanctificabitque caput eius in die illo
NUM|6|12|et consecrabit Domino dies separationis suae offerens agnum anniculum pro delicto; ita tamen, ut dies priores irriti fiant, quoniam polluta est consecratio eius.
NUM|6|13|Ista est lex consecrationis, cum dies, quos ex voto decreverat, complebuntur: adducent eum ad ostium tabernaculi conventus,
NUM|6|14|et offeret oblationem suam Domino agnum anniculum immaculatum in holocaustum et ovem anniculam immaculatam pro peccato et arietem immaculatum hostiam pacificam,
NUM|6|15|canistrum quoque panum azymorum, qui permixti sint oleo, et lagana absque fermento uncta oleo ac oblationem et libamina singulorum.
NUM|6|16|Quae offeret sacerdos coram Domino et faciet tam pro peccato quam in holocaustum;
NUM|6|17|arietem vero immolabit hostiam pacificam Domino offerens simul canistrum azymorum; facietque oblationem eius et libamenta.
NUM|6|18|Tunc radet nazaraeus ante ostium tabernaculi conventus caesariem consecrationis suae tolletque capillos suos et ponet super ignem, qui est suppositus sacrificio pacificorum,
NUM|6|19|et sumet sacerdos armum coctum arietis tortamque absque fermento unam de canistro et laganum azymum unum et tradet in manus nazaraei, postquam rasum fuerit caput eius;
NUM|6|20|et agitabit in conspectu Domini, et sanctificata sacerdotis erunt sicut pectusculum, quod agitari, et femur, quod praelevari iussum est. Post haec potest bibere nazaraeus vinum ".
NUM|6|21|Ista est lex nazaraei, cum voverit oblationem suam Domino tempore consecrationis suae, exceptis his, quae invenerit manus eius. Iuxta quod devoverat, ita faciet secundum legem consecrationis suae.
NUM|6|22|Locutusque est Dominus ad Moysen dicens:
NUM|6|23|" Loquere Aaron et filiis eius: Sic benedicetis filiis Israel et dicetis eis:
NUM|6|24|"Benedicat tibi Dominus et custodiat te!
NUM|6|25|Illuminet Dominus faciem suam super te et misereatur tui!
NUM|6|26|Convertat Dominus vultum suum ad te et det tibi pacem!".
NUM|6|27|Invocabuntque nomen meum super filios Israel, et ego benedicam eis ".
NUM|7|1|Factum est autem in die, qua complevit Moyses habitaculum et erexit illud unxitque et sanctificavit cum omnibus vasis suis, altare similiter et omnia vasa eius,
NUM|7|2|obtulerunt principes Israel et capita familiarum, qui erant per singulas tribus praefecti eorum, qui numerati fuerant,
NUM|7|3|munera coram Domino sex plaustra tecta cum duodecim bobus. Unum plaustrum obtulere duo duces et unum bovem singuli; obtuleruntque ea in conspectu habitaculi.
NUM|7|4|Ait autem Dominus ad Moysen:
NUM|7|5|" Suscipe ab eis, ut serviant in ministerio tabernaculi conventus, et trades ea Levitis iuxta ordinem ministerii sui ".
NUM|7|6|Itaque cum suscepisset Moyses plaustra et boves, tradidit eos Levitis.
NUM|7|7|Duo plaustra et quattuor boves dedit filiis Gerson, iuxta id quod habebant necessarium.
NUM|7|8|Quattuor alia plaustra et octo boves dedit filiis Merari, secundum offficia sua sub manu Ithamar filii Aaron sacerdotis.
NUM|7|9|Filiis autem Caath non dedit plaustra et boves, quia in sanctuario serviunt et onera propriis portant umeris.
NUM|7|10|Igitur obtulerunt duces in dedicationem altaris die, qua unctum est, oblationem suam ante altare.
NUM|7|11|Dixitque Dominus ad Moysen: " Singuli duces per singulos dies offerant munera in dedicationem altaris ".
NUM|7|12|Primo die obtulit oblationem suam Naasson filius Aminadab de tribu Iudae.
NUM|7|13|Fueruntque in ea scutula argentea pondo centum triginta siclorum, phiala argentea habens septuaginta siclos iuxta pondus sanctuarii, utraque plena simila conspersa oleo in sacrificium,
NUM|7|14|acetabulum ex decem siclis aureis plenum incenso,
NUM|7|15|bos de armento et aries et agnus anniculus in holocaustum
NUM|7|16|hircusque pro peccato;
NUM|7|17|et in sacrificio pacificorum boves duo, arietes quinque, hirci quinque, agni anniculi quinque: haec est oblatio Naasson filii Aminadab.
NUM|7|18|Secundo die obtulit Nathanael filius Suar dux de tribu Issachar
NUM|7|19|scutulam argenteam appendentem centum triginta siclos, phialam argenteam habentem septuaginta siclos iuxta pondus sanctuarii, utramque plenam simila conspersa oleo in sacrificium,
NUM|7|20|acetabulum aureum habens decem siclos plenum incenso,
NUM|7|21|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|22|hircumque pro peccato;
NUM|7|23|et in sacrificio pacificorum boves duos, arietes quinque, hircos quinque, agnos anniculos quinque: haec fuit oblatio Nathanael filii Suar.
NUM|7|24|Tertio die princeps filiorum Zabulon Eliab filius Helon
NUM|7|25|obtulit scutulam argenteam appendentem centum triginta siclos, phialam argenteam habentem septuaginta siclos ad pondus sanctuarii, utramque plenam simila conspersa oleo in sacrificium,
NUM|7|26|acetabulum aureum appendens decem siclos plenum incenso,
NUM|7|27|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|28|hircumque pro peccato;
NUM|7|29|et in sacrificio pacificorum boves duos, arietes quinque, hircos quinque, agnos anniculos quinque: haec est oblatio Eliab filii Helon.
NUM|7|30|Die quarto princeps filiorum Ruben Elisur filius Sedeur
NUM|7|31|obtulit scutulam argenteam appendentem centum triginta siclos, phialam argenteam habentem septuaginta siclos ad pondus sanctuarii, utramque plenam simila conspersa oleo in sacrificium,
NUM|7|32|acetabulum aureum appendens decem siclos plenum incenso,
NUM|7|33|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|34|hircumque pro peccato;
NUM|7|35|et in hostias pacificorum boves duos, arietes quinque, hircos quinque, agnos anniculos quinque: haec fuit oblatio Elisur filii Sedeur.
NUM|7|36|Die quinto princeps filiorum Simeon Salamiel filius Surisaddai
NUM|7|37|obtulit scutulam argenteam appendentem centum triginta siclos, phialam argenteam habentem septuaginta siclos ad pondus sanctuarii, utramque plenam simila conspersa oleo in sacrificium,
NUM|7|38|acetabulum aureum appendens decem siclos plenum incenso,
NUM|7|39|bovem de armento et arietem et agnum anniculum in holocaustum,
NUM|7|40|hircumque pro peccato;
NUM|7|41|et in hostias pacificorum boves duos, arietes quinque, hircos quinque, agnos anniculos quinque: haec fuit oblatio Salamiel filii Surisaddai.
NUM|7|42|Die sexto princeps filiorum Gad Eliasaph filius Deuel
NUM|7|43|obtulit scutulam argenteam appendentem centum triginta siclos, phialam argenteam habentem septuaginta siclos ad pondus sanctuarii, utramque plenam simila conspersa oleo in sacrificium,
NUM|7|44|acetabulum aureum appendens decem siclos plenum incenso,
NUM|7|45|bovem de armento et arietem et agnum anniculum in holocaustum,
NUM|7|46|hircumque pro peccato;
NUM|7|47|et in hostias pacificorum boves duos, arietes quinque, hircos quinque, agnos anniculos quinque: haec fuit oblatio Eliasaph filii Deuel.
NUM|7|48|Die septimo princeps filiorum Ephraim Elisama filius Ammiud
NUM|7|49|obtulit scutulam argenteam appendentem centum triginta siclos, phialam argenteam habentem septuaginta siclos ad pondus sanctuarii, utramque plenam simila conspersa oleo in sacrificium,
NUM|7|50|acetabulum aureum appendens decem siclos plenum incenso,
NUM|7|51|bovem de armento et arietem et agnum anniculum in holocaustum,
NUM|7|52|hircumque pro peccato;
NUM|7|53|et in hostias pacificorum boves duos, arietes quinque, hircos quinque, agnos anniculos quinque: haec fuit oblatio Elisama filii Ammiud.
NUM|7|54|Die octavo princeps filiorum Manasse Gamaliel filius Phadassur
NUM|7|55|obtulit scutulam argenteam appendentem centum triginta siclos, phialam argenteam habentem septuaginta siclos ad pondus sanctuarii, utramque plenam simila conspersa oleo in sacrificium,
NUM|7|56|acetabulum aureum appendens decem siclos plenum incenso,
NUM|7|57|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|58|hircumque pro peccato;
NUM|7|59|et in hostias pacificorum boves duos, arietes quinque, hircos quinque, agnos anniculos quinque: haec fuit oblatio Gamaliel filii Phadassur.
NUM|7|60|Die nono princeps filiorum Beniamin Abidan filius Gedeonis
NUM|7|61|obtulit scutulam argenteam appendentem centum triginta siclos, phialam argenteam habentem septuaginta siclos ad pondus sanctuarii, utramque plenam simila conspersa oleo in sacrificium,
NUM|7|62|et acetabulum aureum appendens decem siclos plenum incenso,
NUM|7|63|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|64|hircumque pro peccato;
NUM|7|65|et in hostias pacificorum boves duos, arietes quinque, hircos quinque, agnos anniculos quinque: haec fuit oblatio Abidan filii Gedeonis.
NUM|7|66|Die decimo princeps filiorum Dan Ahiezer filius Ammisaddai
NUM|7|67|obtulit scutulam argenteam appendentem centum triginta siclos, phialam argenteam habentem septuaginta siclos ad pondus sanctuarii, utramque plenam simila conspersa oleo in sacrificium,
NUM|7|68|acetabulum aureum appendens decem siclos plenum incenso,
NUM|7|69|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|70|hircumque pro peccato;
NUM|7|71|et in hostias pacificorum boves duos, arietes quinque, hircos quinque, agnos anniculos quinque: haec fuit oblatio Ahiezer filii Ammisaddai.
NUM|7|72|Die undecimo princeps filiorum Aser Phegiel filius Ochran
NUM|7|73|obtulit scutulam argenteam appendentem centum triginta siclos, phialam argenteam habentem septuaginta siclos ad pondus sanctuarii, utramque plenam simila conspersa oleo in sacrificium,
NUM|7|74|acetabulum aureum appendens decem siclos plenum incenso,
NUM|7|75|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|76|hircumque pro peccato;
NUM|7|77|et in hostias pacificorum boves duos, arietes quinque, hircos quinque, agnos anniculos quinque: haec fuit oblatio Phegiel filii Ochran.
NUM|7|78|Die duodecimo princeps filiorum Nephthali Ahira filius Enan
NUM|7|79|obtulit scutulam argenteam appendentem centum triginta siclos, phialam argenteam habentem septuaginta siclos ad pondus sanctuarii, utramque plenam simila oleo conspersa in sacrificium,
NUM|7|80|acetabulum aureum appendens decem siclos plenum incenso,
NUM|7|81|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|82|hircumque pro peccato;
NUM|7|83|et in hostias pacificorum boves duos, arietes quinque, hircos quinque, agnos anniculos quinque: haec fuit oblatio Ahira filii Enan.
NUM|7|84|Haec in dedicatione altaris oblata sunt a principibus Israel in die, qua consecratum est: scutulae argenteae duodecim, phialae argenteae duodecim, acetabula duodecim,
NUM|7|85|ita ut centum triginta siclos argenti haberet una scutella, et septuaginta siclos haberet una phiala, id est in commune vasorum omnium ex argento sicli duo milia quadringenti pondere sanctuarii;
NUM|7|86|acetabula aurea duodecim plena incenso denos siclos appendentia pondere sanctuarii, id est simul auri sicli centum viginti;
NUM|7|87|omnes boves de armento in holocaustum duodecim, arietes duodecim, agni anniculi duodecim et libamenta eorum; hirci duodecim pro peccato.
NUM|7|88|In hostias pacificorum omnes boves viginti quattuor, arietes sexaginta, hirci sexaginta, agni anniculi sexaginta: haec oblata sunt in dedicatione altaris, quando unctum est.
NUM|7|89|Cumque ingrederetur Moyses tabernaculum testimonii, ut consuleret oraculum, audiebat vocem loquentis ad se de propitiatorio, quod erat super arcam testimonii inter duos cherubim, unde et loquebatur ei.
NUM|8|1|Locutusque est Dominus ad Moysen dicens:
NUM|8|2|" Loquere Aa ron et dices ad eum: Cum posueris lucernas, contra eam partem, quam candelabrum respicit, lucere debebunt septem lucernae ".
NUM|8|3|Fecitque sic Aaron et posuit lucernas super candelabrum, ut praeceperat Dominus Moysi.
NUM|8|4|Haec autem erat factura candelabri: ex auro ductili, tam medius stipes quam flores eius. Iuxta exemplum, quod ostendit Dominus Moysi, ita operatus est candelabrum.
NUM|8|5|Et locutus est Dominus ad Moysen dicens:
NUM|8|6|" Tolle Levitas de medio filiorum Israel et purificabis eos
NUM|8|7|iuxta hunc ritum. Aspergantur aqua lustrationis et radant omnes pilos carnis suae, lavabunt vestimenta sua et mundabunt se.
NUM|8|8|Tollent bovem de armentis et oblationem eius similam oleo conspersam; bovem autem alterum de armento tu accipies pro peccato
NUM|8|9|et applicabis Levitas coram tabernaculo conventus, convocata omni multitudine filiorum Israel.
NUM|8|10|Cumque Levitae fuerint coram Domino, ponent filii Israel manus suas super eos,
NUM|8|11|et agitabit Aaron Levitas munus in conspectu Domini a filiis Israel, ut serviant in ministerio eius.
NUM|8|12|Levitae quoque ponent manus suas super capita boum, e quibus unum facies pro peccato et alterum in holocaustum Domini, ut expies eos.
NUM|8|13|Statuesque Levitas in conspectu Aaron et filiorum eius et agitabis eos Domino
NUM|8|14|ac separabis de medio filiorum Israel, ut sint mei;
NUM|8|15|et postea ingredientur, ut serviant tabernaculo conventus.Sicque purificabis et agitabis eos,
NUM|8|16|quoniam dono donati sunt mihi e medio filiorum Israel; pro primogenitis, quae aperiunt omnem vulvam in Israel, accepi eos.
NUM|8|17|Mea sunt enim omnia primogenita filiorum Israel, tam ex hominibus quam ex iumentis. Ex die, quo percussi omne primogenitum in terra Aegypti, sanctificavi eos mihi.
NUM|8|18|Et tuli Levitas pro cunctis primogenitis filiorum Israel
NUM|8|19|tradidique eos dono Aaron et filiis eius de medio filiorum Israel, ut serviant mihi pro Israel in tabernaculo conventus et expient pro eis, ne sit in populo plaga, si ausi fuerint accedere ad sanctuarium ".
NUM|8|20|Feceruntque Moyses et Aaron et omnis congregatio filiorum Israel super Levitis, quae praeceperat Dominus Moysi.
NUM|8|21|Purificatique sunt et laverunt vestimenta sua, agitavitque eos Aaron in conspectu Domini et expiavit eos, ut purificati
NUM|8|22|ingrederentur ad officia sua in tabernaculo conventus coram Aaron et filiis eius; sicut praeceperat Dominus Moysi de Levitis, ita factum est.
NUM|8|23|Locutusque est Dominus ad Moysen dicens:
NUM|8|24|" Haec est lex Levitarum: a viginti quinque annis et supra ingredientur, ut ministrent in tabernaculo conventus;
NUM|8|25|cumque quinquagesimum annum aetatis impleverint, servire cessabunt
NUM|8|26|eruntque ministri fratrum suorum in tabernaculo conventus, ut custodiant, quae sibi fuerint commendata; opera autem ipsa non faciant. Sic dispones Levitis in custodiis suis ".
NUM|9|1|Locutus est Dominus ad Moy sen in deserto Sinai anno secun do, postquam egressi sunt de terra Aegypti, mense primo dicens:
NUM|9|2|" Faciant filii Israel Pascha in tempore suo
NUM|9|3|quarta decima die mensis huius ad vesperam iuxta omnia praecepta et iustificationes eius ".
NUM|9|4|Praecepitque Moyses filiis Israel, ut facerent Pascha.
NUM|9|5|Qui fecerunt tempore suo quarta decima die mensis ad vesperam in deserto Sinai; iuxta omnia, quae mandaverat Dominus Moysi, fecerunt filii Israel.
NUM|9|6|Ecce autem quidam immundi super animam hominis, qui non poterant facere Pascha in die illo, accedentes ad Moysen et Aaron
NUM|9|7|dixerunt ei: " Immundi sumus super animam hominis; quare fraudamur, ut non valeamus oblationem offerre Domino in tempore suo inter filios Israel? ".
NUM|9|8|Quibus respondit Moyses: " State, ut consulam quid praecipiat Dominus de vobis ".
NUM|9|9|Locutusque est Dominus ad Moysen dicens:
NUM|9|10|" Loquere filiis Israel: Homo, qui fuerit immundus super anima, sive in via procul in gente vestra, faciat Pascha Domino
NUM|9|11|in mense secundo quarta decima die mensis ad vesperam; cum azymis et lactucis agrestibus comedent illud,
NUM|9|12|non relinquent ex eo quippiam usque mane et os eius non confringent: omnem ritum Pascha observabunt.
NUM|9|13|Si quis autem et mundus est et in itinere non fuit et tamen non fecit Pascha, exterminabitur anima illa de populis suis, quia sacrificium Domino non obtulit tempore suo: peccatum suum ipse portabit.
NUM|9|14|Peregrinus quoque et advena, si fuerint apud vos, facient Pascha Domino iuxta praecepta et iustificationes eius; praeceptum idem erit apud vos tam advenae quam indigenae ".
NUM|9|15|Igitur die, qua erectum est habitaculum, operuit nubes habitaculum, tabernaculum testimonii; a vespere autem super habitaculum erat quasi species ignis usque mane.
NUM|9|16|Sic fiebat iugiter: per diem operiebat illud nubes, et per noctem quasi species ignis.
NUM|9|17|Cumque ablata fuisset nubes, quae tabernaculum protegebat, tunc proficiscebantur filii Israel; et in loco, ubi stetisset nubes, ibi castrametabantur.
NUM|9|18|Ad imperium Domini proficiscebantur et ad imperium illius castrametabantur. Cunctis diebus, quibus stabat nubes super habitaculum, manebant in eodem loco.
NUM|9|19|Et si evenisset ut multo tempore maneret super illud, erant filii Israel in excubiis Domini et non proficiscebantur;
NUM|9|20|si diebus paucis fuisset nubes super habitaculum, ad imperium Domini erigebant tentoria et ad imperium illius deponebant.
NUM|9|21|Si fuisset nubes a vespere usque mane et statim diluculo habitaculum reliquisset, proficiscebantur; et si post diem et noctem recessisset, dissipabant tentoria.
NUM|9|22|Si vero biduo aut uno mense vel longiore tempore fuisset super habitaculum, manebant filii Israel in eodem loco et non proficiscebantur. Statim autem ut recessisset, movebant castra.
NUM|9|23|Per verbum Domini figebant tentoria et per verbum illius proficiscebantur; erantque in excubiis Domini iuxta imperium eius per manum Moysi.
NUM|10|1|Locutusque est Dominus ad Moysen dicens:
NUM|10|2|" Fac tibi duas tubas argenteas ductiles, quibus convocare possis congregationem, quando movenda sunt castra.
NUM|10|3|Cumque increpueris tubis, congregabitur ad te omnis turba ad ostium tabernaculi conventus.
NUM|10|4|Si semel clangueris, venient ad te principes et capita congregationis Israel;
NUM|10|5|si autem prolixior clangor increpuerit, movebunt castra primi, qui sunt ad orientalem plagam;
NUM|10|6|in secundo autem sonitu et pari ululatu tubae levabunt tentoria, qui habitant ad meridiem, et iuxta hunc modum reliqui facient, ululantibus tubis in profectionem.
NUM|10|7|Quando autem congregandus est populus, simplex tubarum clangor erit, et non ululabunt.
NUM|10|8|Filii autem Aaron sacerdotes clangent tubis. Eritque hoc vobis legitimum sempiternum in generationibus vestris.
NUM|10|9|Si exieritis ad bellum in terra vestra contra hostes, qui dimicant adversum vos, clangetis ululantibus tubis; et erit recordatio vestri coram Domino Deo vestro, ut eruamini de manibus inimicorum vestrorum.
NUM|10|10|Si quando habebitis epulum et dies festos et calendas, canetis tubis super holocaustis vestris et pacificis victimis, ut sint vobis in recordationem Dei vestri. Ego Dominus Deus vester ".
NUM|10|11|Anno secundo, mense secundo, vicesima die mensis elevata est nubes de habitaculo testimonii;
NUM|10|12|profectique sunt filii Israel per migrationes suas de deserto Sinai, et recubuit nubes in solitudine Pharan.
NUM|10|13|Moveruntque castra prima vice, iuxta imperium Domini in manu Moysi.
NUM|10|14|Elevatum est primum vexillum castrorum filiorum Iudae per turmas suas, quorum princeps erat Naasson filius Aminadab;
NUM|10|15|et super turmam tribus filiorum Issachar fuit princeps Nathanael filius Suar;
NUM|10|16|et super turmam tribus Zabulon erat princeps Eliab filius Helon.
NUM|10|17|Depositumque est habitaculum, quod portantes egressi sunt filii Gerson et Merari.
NUM|10|18|Profectum est vexillum castrorum filiorum Ruben per turmas suas, et super turbam suam princeps erat Elisur filius Sedeur.
NUM|10|19|Super turmam autem tribus filiorum Simeon princeps fuit Salamiel filius Surisaddai.
NUM|10|20|Porro super turmam tribus filiorum Gad erat princeps Eliasaph filius Deuel.
NUM|10|21|Profectique sunt et Caathitae portantes sanctuarium. Et erectum est habitaculum, antequam venirent.
NUM|10|22|Elevatum est vexillum castrorum filiorum Ephraim per turmas suas, in quorum exercitu princeps erat Elisama filius Ammiud.
NUM|10|23|Et super turmam tribus filiorum Manasse princeps fuit Gamaliel filius Phadassur;
NUM|10|24|et super turmam tribus filiorum Beniamin erat dux Abidan filius Gedeonis.
NUM|10|25|Novissime elevatum est vexillum castrorum filiorum Dan per turmas suas, in quorum exercitu princeps fuit Ahiezer filius Ammisaddai.
NUM|10|26|Et super turmam tribus filiorum Aser erat princeps Phegiel filius Ochran;
NUM|10|27|et super turmam tribus filiorum Nephthali princeps fuit Ahira filius Enan.
NUM|10|28|Hae sunt profectiones filiorum Israel per turmas suas, quando egrediebantur.
NUM|10|29|Dixitque Moyses Hobab filio Raguel Madianitae cognato suo: " Proficiscimur ad locum, quem Dominus daturus est nobis; veni nobiscum, ut benefaciamus tibi, quia Dominus bona promisit Israeli ".
NUM|10|30|Cui ille respondit: " Non vadam tecum, sed revertar in terram meam, in qua natus sum ".
NUM|10|31|Et ille: " Noli, inquit, nos relinquere; tu enim nosti in quibus locis per desertum castra ponere debeamus, et eris ductor noster.
NUM|10|32|Cumque nobiscum veneris, quidquid optimum fuerit ex opibus, quas nobis traditurus est Dominus, dabimus tibi ".
NUM|10|33|Profecti sunt ergo de monte Domini viam trium dierum; arcaque foederis Domini praecedebat eos per dies tres providens castrorum locum.
NUM|10|34|Nubes quoque Domini super eos erat per diem, cum incederent.
NUM|10|35|Cumque elevaretur arca, dicebat Moyses: " Surge, Domine, et dissipentur inimici tui; et fugiant, qui oderunt te, a facie tua ".
NUM|10|36|Cum autem deponeretur, aiebat: " Revertere, Domine, ad multitudinem exercitus Israel ".
NUM|11|1|Ortum est murmur populi, quasi dolentium pro labore, contra Dominum. Quod cum audisset Dominus, iratus est, et accensus in eos ignis Domini devoravit extremam castrorum partem.
NUM|11|2|Cumque clamasset populus ad Moysen, oravit Moyses ad Dominum, et absorptus est ignis.
NUM|11|3|Vocaverunt nomen loci illius Tabera, eo quod incensus fuisset contra eos ignis Domini.
NUM|11|4|Vulgus autem promiscuum, quod erat in medio eius, flagravit desiderio, et sedentes fleverunt pariter filii Israel et dixerunt: " Quis dabit nobis ad vescendum carnes?
NUM|11|5|Recordamur piscium, quos comedebamus in Aegypto gratis; in mentem nobis veniunt cucumeres et pepones porrique et cepae et alia.
NUM|11|6|Guttur nostrum aridum est; nihil aliud respiciunt oculi nostri nisi man ".
NUM|11|7|Erat autem man quasi semen coriandri aspectus bdellii.
NUM|11|8|Circuibatque populus et colligens illud frangebat mola sive terebat in mortario coquens in olla et faciens ex eo tortulas saporis quasi panis oleati.
NUM|11|9|Cumque descenderet nocte super castra ros, descendebat pariter et man.
NUM|11|10|Audivit ergo Moyses flentem populum per familias, singulos per ostia tentorii sui. Iratusque est furor Domini valde; quod Moysi intoleranda res visa est,
NUM|11|11|et ait ad Dominum: " Cur afflixisti servum tuum? Quare non invenio gratiam coram te? Et cur imposuisti pondus universi populi huius super me?
NUM|11|12|Numquid ego concepi omnem hunc populum vel genui eum, ut dicas mihi: "Porta eum in sinu tuo, sicut portare solet nutrix infantulum, et defer in terram, pro qua iurasti patribus eorum?".
NUM|11|13|Unde mihi carnes, ut dem universo populo isti? Flent contra me dicentes: "Da nobis carnes, ut comedamus!".
NUM|11|14|Non possum ego solus sustinere omnem hunc populum, quia nimis gravis est mihi.
NUM|11|15|Si hoc modo agis mecum, obsecro ut interficias me, si inveni gratiam in oculis tuis, ne videam amplius mala mea! ".
NUM|11|16|Et dixit Dominus ad Moysen: " Congrega mihi septuaginta viros de senibus Israel, quos tu nosti quod senes populi sint ac magistri, et duces eos ad ostium tabernaculi conventus, stabuntque ibi tecum.
NUM|11|17|Et descendam et loquar tibi et auferam de spiritu tuo tradamque eis, ut sustentent tecum onus populi, et non tu solus graveris.
NUM|11|18|Populo quoque dices: Sanctificamini, cras comedetis carnes; ego enim audivi vos flere: "Quis dabit nobis escas carnium? Bene nobis erat in Aegypto". Et dabit vobis Dominus carnes, et comedetis
NUM|11|19|non uno die nec duobus vel quinque aut decem nec viginti quidem,
NUM|11|20|sed usque ad mensem dierum, donec exeat per nares vestras et vertatur in nauseam, eo quod reppuleritis Dominum, qui in medio vestri est, et fleveritis coram eo dicentes: "Quare egressi sumus ex Aegypto?" ".
NUM|11|21|Et ait Moyses: " Populus, in cuius medio sum, sescenta milia peditum sunt, et tu dicis: "Dabo eis esum carnium mense integro!".
NUM|11|22|Numquid ovium et boum multitudo caedetur, ut possit sufficere ad cibum? Vel omnes pisces maris in unum congregabuntur, ut eos satient? ".
NUM|11|23|Cui respondit Dominus: " Numquid manus Domini abbreviata est? Iam nunc videbis utrum meus sermo opere compleatur an non ".
NUM|11|24|Venit igitur Moyses et narravit populo verba Domini congregans septuaginta viros de senibus Israel, quos stare fecit circa tabernaculum.
NUM|11|25|Descenditque Dominus per nubem et locutus est ad eum auferens de spiritu, qui erat in Moyse, et dans septuaginta viris senibus. Cumque requievisset in eis spiritus, prophetaverunt nec ultra fecerunt.
NUM|11|26|Remanserant autem in castris duo viri, quorum unus vocabatur Eldad et alter Medad, super quos requievit spiritus; nam et ipsi descripti fuerant et non exierant ad tabernaculum. Cumque prophetarent in castris,
NUM|11|27|cucurrit puer et nuntiavit Moysi dicens: " Eldad et Medad prophetant in castris ".
NUM|11|28|Statim Iosue filius Nun minister Moysi et electus eius a iuventute sua ait: " Domine mi Moyses, prohibe eos! ".
NUM|11|29|At ille: " Quid, inquit, aemularis pro me? Quis tribuat, ut omnis populus prophetet, et det eis Dominus spiritum suum? ".
NUM|11|30|Reversusque est Moyses et maiores natu Israel in castra.
NUM|11|31|Ventus autem egrediens a Domino arreptas trans mare coturnices detulit et demisit in castra itinere, quantum uno die confici potest, ex omni parte castrorum per circuitum; volabantque in aere duobus cubitis altitudine super terram.
NUM|11|32|Surgens ergo populus toto die illo et nocte ac die altero congregavit coturnicum, qui parum, decem choros; et extenderunt eas per gyrum castrorum.
NUM|11|33|Adhuc carnes erant in dentibus eorum, nec defecerat huiuscemodi cibus, et ecce furor Domini concitatus in populum percussit eum plaga magna nimis.
NUM|11|34|Vocatusque est ille locus Cibrottaava; ibi enim sepelierunt populum, qui desideraverat.
NUM|11|35|Egressi autem de Cibrottaava, venerunt in Aseroth et manserunt ibi.
NUM|12|1|Locutaque est Maria et Aaron contra Moysen propter uxorem eius Aethiopissam
NUM|12|2|et dixerunt: " Num per solum Moysen locutus est Dominus? Nonne et per nos similiter est locutus? ". Quod cum audisset Dominus
NUM|12|3|­ erat enim Moyses vir humillimus super omnes homines, qui morabantur in terra ­
NUM|12|4|statim locutus est ad eum et ad Aaron et Mariam: " Egredimini vos tantum tres ad tabernaculum conventus ". Cumque fuissent egressi,
NUM|12|5|descendit Dominus in columna nubis et stetit in introitu tabernaculi vocans Aaron et Mariam. Qui cum issent,
NUM|12|6|dixit ad eos:" Audite sermones meos!Si quis fuerit inter vos propheta Domini,in visione apparebo eivel per somnium loquar ad illum.
NUM|12|7|At non talis servus meus Moyses,qui in omni domo mea fidelissimus est!
NUM|12|8|Ore enim ad os loquor ei,et palam et non per aenigmata et figurasDominum videt!Quare ergo non timuistis detrahereservo meo Moysi? ".
NUM|12|9|Iratusque contra eos abiit,
NUM|12|10|nubes quoque recessit, quae erat super tabernaculum; et ecce Maria apparuit candens lepra quasi nix.Cumque respexisset eam Aaron et vidisset perfusam lepra,
NUM|12|11|ait ad Moysen: " Obsecro, domine mi, ne imponas nobis hoc peccatum, quod stulte commisimus,
NUM|12|12|ne fiat haec quasi mortua et ut abortivum, quod proicitur de vulva matris suae; ecce iam medium carnis eius devoratum est a lepra ".
NUM|12|13|Clamavitque Moyses ad Dominum dicens: " Deus, obsecro, sana eam! ".
NUM|12|14|Cui respondit Dominus: " Si pater eius spuisset in faciem illius, nonne debuerat saltem septem diebus rubore suffundi? Separetur septem diebus extra castra et postea revocabitur ".
NUM|12|15|Exclusa est itaque Maria extra castra septem diebus, et populus non est motus de loco illo, donec revocata est Maria.
NUM|12|16|Profectusque est populus de Aseroth, fixis tentoriis in deserto Pharan.
NUM|13|1|Ibi locutus est Dominus ad Moysen dicens:
NUM|13|2|" Mitte vi ros, qui considerent terram Chanaan, quam daturus sum filiis Israel, singulos de singulis tribubus ex principibus ".
NUM|13|3|Fecit Moyses quod Dominus imperaverat, de deserto Pharan mittens principes viros, quorum ista sunt nomina:
NUM|13|4|de tribu Ruben Sammua filium Zacchur,
NUM|13|5|de tribu Simeon Saphat filium Hori,
NUM|13|6|de tribu Iudae Chaleb filium Iephonne,
NUM|13|7|de tribu Issachar Igal filium Ioseph,
NUM|13|8|de tribu Ephraim Osee filium Nun,
NUM|13|9|de tribu Beniamin Phalti filium Raphu,
NUM|13|10|de tribu Zabulon Geddiel filium Sodi,
NUM|13|11|de tribu Ioseph, tribu Manasse, Gaddi filium Susi,
NUM|13|12|de tribu Dan Ammiel filium Gemalli,
NUM|13|13|de tribu Aser Sthur filium Michael,
NUM|13|14|de tribu Nephthali Nahabi filium Vaphsi,
NUM|13|15|de tribu Gad Guel filium Machi.
NUM|13|16|Haec sunt nomina virorum, quos misit Moyses ad considerandam terram. Vocavitque Osee filium Nun Iosue.
NUM|13|17|Misit ergo eos Moyses ad considerandam terram Chanaan et dixit ad eos: " Ascendite per Nageb. Cumque veneritis ad montes,
NUM|13|18|considerate terram, qualis sit, et populum, qui habitator est eius, utrum fortis sit an infirmus, si pauci numero an plures;
NUM|13|19|ipsa terra bona an mala, urbes quales, absque muris an muratae;
NUM|13|20|humus pinguis an sterilis, nemorosa an absque arboribus. Confortamini et afferte nobis de fructibus terrae ". Erat autem tempus, quando iam praecoquae uvae vesci possunt.
NUM|13|21|Cumque ascendissent, exploraverunt terram a deserto Sin usque Rohob in introitu Emath.
NUM|13|22|Ascenderuntque ad Nageb et venerunt in Hebron, ubi erant Ahiman et Sesai et Tholmai filii Enac. Nam Hebron septem annis ante Tanim urbem Aegypti condita est.
NUM|13|23|Pergentesque usque ad Nehelescol absciderunt palmitem cum uva sua, quem portaverunt in vecte duo viri. De malis quoque granatis et de ficis loci illius tulerunt,
NUM|13|24|qui appellatus est Nehelescol, eo quod botrum portassent inde filii Israel.
NUM|13|25|Reversique exploratores terrae post quadraginta dies, omni regione circuita,
NUM|13|26|venerunt ad Moysen et Aaron et ad omnem coetum filiorum Israel in desertum Pharan, quod est in Cades. Locutique eis et omni congregationi ostenderunt fructus terrae
NUM|13|27|et narraverunt dicentes: " Venimus in terram, ad quam misisti nos, quae re vera fluit lacte et melle, ut ex his fructibus cognosci potest.
NUM|13|28|Sed cultores fortissimos habet et urbes grandes atque muratas. Stirpem Enac vidimus ibi;
NUM|13|29|Amalec habitat in Nageb, Hetthaeus et Iebusaeus et Amorraeus in montanis, Chananaeus vero moratur iuxta mare et circa fluenta Iordanis ".
NUM|13|30|Inter haec Chaleb compescens murmur populi, qui oriebatur contra Moysen, ait: " Ascendamus et possideamus terram, quoniam poterimus obtinere eam ".
NUM|13|31|Alii vero, qui fuerant cum eo, dicebant: " Nequaquam ad hunc populum valemus ascendere, quia fortior nobis est ".
NUM|13|32|Detraxeruntque terrae, quam inspexerant, apud filios Israel dicentes: " Terra, quam lustravimus, devorat habitatores suos; populus, quem aspeximus, procerae staturae est;
NUM|13|33|ibi vidimus gigantes, filios Enac de genere giganteo, quibus comparati quasi locustae videbamur ".
NUM|14|1|Igitur vociferans omnis tur ba flevit nocte illa,
NUM|14|2|et mur murati sunt contra Moysen et Aaron cuncti filii Israel dicentes: " Utinam mortui essemus in Aegypto vel in hac vasta solitudine!
NUM|14|3|Cur inducit nos Dominus in terram istam, ut cadamus gladio, et uxores ac liberi nostri ducantur captivi? Nonne melius est reverti in Aegyptum? ".
NUM|14|4|Dixeruntque alter ad alterum: " Constituamus nobis ducem et revertamur in Aegyptum! ".
NUM|14|5|Quo audito, Moyses et Aaron ceciderunt proni in terram coram omni congregatione filiorum Israel.
NUM|14|6|At vero Iosue filius Nun et Chaleb filius Iephonne, qui et ipsi lustraverant terram, sciderunt vestimenta sua
NUM|14|7|et ad omnem congregationem filiorum Israel locuti sunt: " Terra, quam circuivimus, valde bona est.
NUM|14|8|Si propitius fuerit Dominus, inducet nos in eam et tradet humum lacte et melle manantem.
NUM|14|9|Nolite rebelles esse contra Dominum neque timeatis populum terrae huius, quia sicut panem ita eos possumus devorare. Recessit ab eis omne praesidium; Dominus nobiscum est, nolite metuere ".
NUM|14|10|Cumque clamaret omnis congregatio et lapidibus eos vellet opprimere, apparuit gloria Domini super tabernaculum conventus cunctis filiis Israel,
NUM|14|11|et dixit Dominus ad Moysen: " Usquequo detrahet mihi populus iste? Quousque non credent mihi in omnibus signis, quae feci coram eis?
NUM|14|12|Feriam igitur eos pestilentia atque consumam; te autem faciam in gentem magnam et fortiorem quam haec est ".
NUM|14|13|Et ait Moyses ad Dominum:? Audient Aegyptii, de quorum medio eduxisti populum istum in virtute tua,
NUM|14|14|et dicent ad habitatores terrae huius, quia audierunt quod tu, Domine, in populo isto sis et facie videaris ad faciem, et nubes tua protegat illos, et in columna nubis praecedas eos per diem et in columna ignis per noctem.
NUM|14|15|Et occidisti hunc populum quasi unum hominem, et dicent gentes, quae audierunt auditum tuum:
NUM|14|16|"Non poterat Dominus introducere populum in terram, pro qua iuraverat, idcirco occidit eos in solitudine!".
NUM|14|17|Magnificetur ergo fortitudo Domini, sicut iurasti dicens:
NUM|14|18|"Dominus patiens et multae misericordiae, auferens iniquitatem et scelera nullumque innoxium derelinquens, qui visitas peccata patrum in filios in tertiam et quartam generationem".
NUM|14|19|Dimitte obsecro peccatum populi huius secundum magnitudinem misericordiae tuae, sicut propitius fuisti populo huic de Aegypto usque ad locum istum ".
NUM|14|20|Dixitque Dominus: " Dimisi iuxta verbum tuum.
NUM|14|21|Vivo ego, et implebit gloria Domini universam terram!
NUM|14|22|Attamen omnes homines, qui viderunt maiestatem meam et signa, quae feci in Aegypto et in solitudine, et tentaverunt me iam per decem vices nec oboedierunt voci meae,
NUM|14|23|non videbunt terram, pro qua iuravi patribus eorum; nec quisquam ex illis, qui detraxit mihi, intuebitur eam.
NUM|14|24|Servum meum Chaleb, qui plenus alio spiritu secutus est me, inducam in terram hanc, quam circuivit, et semen eius possidebit eam.
NUM|14|25|Quoniam Amalecites et Chananaeus habitant in vallibus, cras movete castra et revertimini in solitudinem per viam maris Rubri ".
NUM|14|26|Locutusque est Dominus ad Moysen et Aaron dicens:
NUM|14|27|" Usquequo congregatio haec pessima murmurat contra me? Querelas filiorum Israel audivi.
NUM|14|28|Dic ergo eis: Vivo ego, ait Dominus, sicut locuti estis, audiente me, sic faciam vobis!
NUM|14|29|In solitudine hac iacebunt cadavera vestra. Omnes, qui numerati estis a viginti annis et supra et murmurastis contra me,
NUM|14|30|non intrabitis terram, super quam levavi manum meam, ut habitare vos facerem, praeter Chaleb filium Iephonne et Iosue filium Nun.
NUM|14|31|Parvulos autem vestros, de quibus dixistis quod praedae hostibus forent, introducam, ut videant terram, quae vobis displicuit.
NUM|14|32|Vestra cadavera iacebunt in solitudine hac;
NUM|14|33|filii vestri erunt pastores in deserto annis quadraginta et portabunt fornicationem vestram, donec consumantur cadavera vestra in deserto.
NUM|14|34|Iuxta numerum quadraginta dierum, quibus considerastis terram ­ annus pro die imputabitur ­ quadraginta annis portabitis iniquitates vestras et scietis ultionem meam.
NUM|14|35|Ego Dominus locutus sum, ita faciam omni congregationi huic pessimae, quae consurrexit adversum me: in solitudine hac deficiet et morietur ".
NUM|14|36|Igitur omnes viri, quos miserat Moyses ad contemplandam terram et qui reversi murmurare fecerant contra eum omnem congregationem detrahentes terrae quod esset mala,
NUM|14|37|mortui sunt atque percussi in conspectu Domini.
NUM|14|38|Iosue autem filius Nun et Chaleb filius Iephonne vixerunt ex omnibus, qui perrexerant ad considerandam terram.
NUM|14|39|Locutusque est Moyses universa verba haec ad omnes filios Israel, et luxit populus nimis.
NUM|14|40|Et ecce mane primo surgentes ascenderunt verticem montis atque dixerunt: " Parati sumus ascendere ad locum, de quo Dominus locutus est, quia peccavimus ".
NUM|14|41|Quibus Moyses: " Cur, inquit, transgredimini verbum Domini, quod vobis non cedet in prosperum?
NUM|14|42|Nolite ascendere, non enim est Dominus vobiscum, ne corruatis coram inimicis vestris!
NUM|14|43|Amalecites et Chananaeus ante vos sunt, quorum gladio corruetis, eo quod nolueritis acquiescere Domino, nec erit Dominus vobiscum ".
NUM|14|44|At illi contenebrati ascenderunt in verticem montis; arca autem foederis Domini et Moyses non recesserunt de castris.
NUM|14|45|Descenditque Amalecites et Chananaeus, qui habitabat in monte, et percutiens eos atque concidens persecutus est eos usque Horma.
NUM|15|1|Locutus est Dominus ad Moysen dicens:
NUM|15|2|" Loquere ad filios Israel et dices ad eos: Cum ingressi fueritis terram habitationis vestrae, quam ego dabo vobis,
NUM|15|3|et feceritis oblationem Domino in holocaustum aut victimam vota solventes vel sponte offerentes munera aut in sollemnitatibus vestris adolentes odorem suavitatis Domino de bobus sive de ovibus,
NUM|15|4|offeret, quicumque immolaverit victimam, sacrificium similae decimam partem ephi conspersae oleo, quod mensuram habebit quartam partem hin,
NUM|15|5|et vinum ad liba fundenda eiusdem mensurae dabit in holocaustum sive in victimam per agnos singulos.
NUM|15|6|Per arietes erit sacrificium similae duarum decimarum, quae conspersa sit oleo tertiae partis hin;
NUM|15|7|et vinum ad libamentum tertiae partis eiusdem mensurae offeret in odorem suavitatis Domino.
NUM|15|8|Quando vero de bobus feceris holocaustum aut hostiam, ut impleas votum vel pacificas victimas,
NUM|15|9|dabis per singulos boves similae tres decimas conspersae oleo, quod habeat medium mensurae hin,
NUM|15|10|et vinum ad liba fundenda eiusdem mensurae in oblationem suavissimi odoris Domino.
NUM|15|11|Sic facies per singulos boves et arietes et agnos et capras.
NUM|15|12|Secundum numerum victimarum quas offeretis, ita facietis singulis secundum numerum earum.
NUM|15|13|Omnis indigena eodem ritu offeret sacrificium ignis in odorem suavitatis Domino.
NUM|15|14|Et omnis peregrinus, qui habitat vobiscum vel qui commoratur in medio vestri in omnibus generationibus vestris, offeret sacrificium ignis in odorem suavitatis Domino eodem modo sicut et vos.
NUM|15|15|Unum praeceptum erit tam vobis quam advenis pro omnibus generationibus vestris coram Domino.
NUM|15|16|Una lex erit atque unum iudicium tam vobis quam advenis, qui vobiscum commorantur ".
NUM|15|17|Locutus est Dominus ad Moysen dicens:
NUM|15|18|" Loquere filiis Israel et dices ad eos: Cum veneritis in terram, quam dabo vobis,
NUM|15|19|et comederitis de panibus regionis illius, separabitis donaria Domino
NUM|15|20|de pulmento placentam. Sicut de areis donaria separatis,
NUM|15|21|ita et de pulmentis dabitis ea Domino.
NUM|15|22|Quod si per ignorantiam praeterieritis quidquam horum, quae locutus est Dominus ad Moysen
NUM|15|23|et mandavit per eum ad vos a die, qua coepit iubere et ultra ad generationes vestras,
NUM|15|24|si longe ab oculis congregationis, offeret congregatio vitulum de armento, holocaustum in odorem placabilem Domino et oblationem ac liba eius, ut caeremoniae postulant, hircumque pro peccato.
NUM|15|25|Et expiabit sacerdos pro omni congregatione filiorum Israel, et dimittetur eis, quoniam non sponte peccaverunt, nihilominus offerentes sacrificium ignis Domino pro se et pro peccato atque errore suo.
NUM|15|26|Et dimittetur universae plebi filiorum Israel et advenis, qui peregrinantur inter eos, quoniam culpa est omnis populi per ignorantiam.
NUM|15|27|Quod si anima una nesciens peccaverit, offeret capram anniculam pro peccato suo.
NUM|15|28|Et expiabit pro ea sacerdos, quod inscia peccaverit coram Domino; expiabit pro ea, et dimittetur illi.
NUM|15|29|Tam indigenis quam advenis una lex erit omnium, qui peccaverint ignorantes.
NUM|15|30|Anima vero, quae per superbiam aliquid commiserit, sive civis sit ille sive peregrinus, quoniam adversus Dominum rebellis fuit, peribit de populo suo.
NUM|15|31|Verbum enim Domini contempsit et praeceptum illius fecit irritum; idcirco delebitur et portabit iniquitatem suam ".
NUM|15|32|Factum est autem, cum essent filii Israel in solitudine et invenissent hominem colligentem ligna in die sabbati,
NUM|15|33|obtulerunt eum Moysi et Aaron et universae congregationi,
NUM|15|34|qui recluserunt eum in carcerem nescientes quid super eo facere deberent.
NUM|15|35|Dixitque Dominus ad Moysen: " Morte moriatur homo iste; obruat eum lapidibus omnis turba extra castra ".
NUM|15|36|Cumque eduxissent eum foras, obruerunt lapidibus; et mortuus est, sicut praeceperat Dominus.
NUM|15|37|Dixit quoque Dominus ad Moysen:
NUM|15|38|" Loquere filiis Israel et dices ad eos, ut faciant sibi fimbrias per angulos palliorum ponentes in eis vittas hyacinthinas.
NUM|15|39|Quas cum videbitis, recordabimini omnium mandatorum Domini eaque facietis nec sequamini cogitationes vestras et oculos per res varias fornicantes,
NUM|15|40|sed magis memores omnium praeceptorum meorum faciatis ea sitisque sancti Deo vestro.
NUM|15|41|Ego Dominus Deus vester, qui eduxi vos de terra Aegypti, ut essem Deus vester. Ego Dominus Deus vester ".
NUM|16|1|Ecce autem Core filius Isaar filii Caath filii Levi et Dathan atque Abiram filii Eliab, Hon quoque filius Pheleth de filiis Ruben
NUM|16|2|surrexerunt contra Moysen aliique filiorum Israel ducenti quinquaginta viri proceres synagogae vocati ad concilium, viri famosi.
NUM|16|3|Cumque stetissent adversum Moysen et Aaron, dixerunt: " Sufficiat vobis quia omnis congregatio sanctorum est, et in ipsis est Dominus! Cur elevamini super congregationem Domini? ".
NUM|16|4|Quod cum audisset Moyses, cecidit pronus in faciem
NUM|16|5|locutusque ad Core et ad omne concilium: " Mane, inquit, notum faciet Dominus qui ad se pertineant et qui sint sancti, et sanctos applicabit sibi; et, quos elegerit, appropinquare sibi faciet.
NUM|16|6|Hoc igitur facite: tollat unusquisque turibulum suum, tu, Core, et omne concilium tuum;
NUM|16|7|et hausto cras igne, ponite desuper thymiama coram Domino; et, quemcumque elegerit, ipse erit sanctus. Sufficiat vobis, filii Levi! ".
NUM|16|8|Dixitque rursum ad Core: " Audite, filii Levi.
NUM|16|9|Num parum vobis est quod separavit vos Deus Israel ab omni congregatione et iunxit sibi, ut serviretis ei in cultu habitaculi Domini et staretis coram frequentia populi et ministraretis pro ea?
NUM|16|10|Idcirco ad se fecit accedere te et omnes fratres tuos filios Levi, ut vobis etiam sacerdotium vindicetis,
NUM|16|11|et omne concilium tuum stet contra Dominum? Quid est enim Aaron, ut murmuretis contra eum? ".
NUM|16|12|Misit ergo Moyses, ut vocaret Dathan et Abiram filios Eliab, qui responderunt: " Non venimus!
NUM|16|13|Numquid parum est tibi quod eduxisti nos de terra, quae lacte et melle manabat, ut occideres in deserto, nisi et dominatus fueris nostri?
NUM|16|14|Revera non induxisti nos in terram, quae fluit rivis lactis et mellis, nec dedisti nobis possessiones agrorum et vinearum! An et oculos illorum hominum vis eruere? Non venimus! ".
NUM|16|15|Iratusque Moyses valde ait ad Dominum: " Ne respicias sacrificia eorum; tu scis quod ne asellum quidem umquam acceperim ab eis nec afflixerim quempiam eorum ".
NUM|16|16|Dixitque ad Core: " Tu et omne concilium tuum state seorsum coram Domino, et Aaron die crastino separatim.
NUM|16|17|Tollite singuli turibula vestra et ponite super ea incensum offerentes Domino ducenta quinquaginta turibula; tu et Aaron teneatis unusquisque turibulum suum ".
NUM|16|18|Quod cum fecissent, stantibus Moyse et Aaron,
NUM|16|19|et coacervasset Core adversum eos omne concilium ad ostium tabernaculi conventus, apparuit cunctis gloria Dornini.
NUM|16|20|Locutusque Dominus ad Moysen et Aaron ait:
NUM|16|21|" Separamini de medio congregationis huius, ut eos repente disperdam ".
NUM|16|22|Qui ceciderunt proni in faciem atque dixerunt: " Deus, Deus spirituum universae carnis; num, uno peccante, contra omnes ira tua desaeviet? ".
NUM|16|23|Et ait Dominus ad Moysen:
NUM|16|24|" Praecipe universo populo, ut separetur ab habitaculis Core et Dathan et Abiram ".
NUM|16|25|Surrexitque Moyses et abiit ad Dathan et Abiram et, sequentibus eum senioribus Israel,
NUM|16|26|dixit ad turbam: " Recedite ab habitaculis hominum impiorum et nolite tangere, quae ad eos pertinent, ne involvamini in peccatis eorum ".
NUM|16|27|Cumque recessissent a tentoriis eorum per circuitum, Dathan et Abiram egressi stabant in introitu papilionum suorum cum uxoribus et filiis et parvulis.
NUM|16|28|Et ait Moyses: " In hoc scietis quod Dominus miserit me, ut facerem universa, quae cernitis, et non ex proprio ea corde protulerim:
NUM|16|29|si consueta hominum morte interierint, et visitaverit eos plaga, qua et ceteri visitari solent, non misit me Dominus.
NUM|16|30|Sin autem novam rem fecerit Dominus, ut aperiens terra os suum deglutiat eos et omnia, quae ad illos pertinent, descenderintque viventes in infernum, scietis quod blasphemaverint Dominum ".
NUM|16|31|Confestim igitur, ut cessavit loqui, dirupta est terra sub pedibus eorum
NUM|16|32|et aperiens os suum devoravit illos cum domibus suis et omnibus hominibus Core et universa substantia eorum;
NUM|16|33|descenderuntque vivi in infernum operti humo et perierunt de medio congregationis.
NUM|16|34|At vero omnis Israel, qui stabat per gyrum, fugit ad clamorem pereuntium dicens: " Ne forte et nos terra deglutiat ".
NUM|16|35|Sed et ignis egressus a Domino interfecit ducentos quinquaginta viros, qui offerebant incensum.
NUM|17|1|Locutusque est Dominus ad Moysen dicens:
NUM|17|2|" Praecipe Eleazaro filio Aaron sacerdoti, ut tollat turibula, quae iacent in incendio, et ignem huc illucque dispergat, quoniam sanctificata sunt
NUM|17|3|in mortibus peccatorum; producatque ea in laminas et affigat altari, eo quod attulerunt ea Domino, et sanctificata sunt, ut sint pro signo filiis Israel ".
NUM|17|4|Tulit ergo Eleazar sacerdos turibula aenea, in quibus obtulerant hi, quos incendium devoravit, et produxit ea in laminas affigens altari,
NUM|17|5|ut haberent postea filii Israel, quibus commonerentur, ne quis accedat alienigena et, qui non est de semine Aaron, ad offerendum incensum Domino, ne patiatur sicut passus est Core et omnis congregatio eius, loquente Domino ad Moysen.
NUM|17|6|Murmuravit autem omnis congregatio filiorum Israel sequenti die contra Moysen et Aaron dicens: " Vos interfecistis populum Domini ".
NUM|17|7|Cumque oriretur seditio contra Moysen et Aaron, converterunt se ad tabernaculum conventus; quod operuit nubes, et apparuit gloria Domini.
NUM|17|8|Moyses et Aaron venerunt ante tabernaculum conventus.
NUM|17|9|Dixitque Dominus ad Moysen:
NUM|17|10|" Recedite de medio congregationis huius, nam extemplo delebo eos ". Et ceciderunt in faciem suam.
NUM|17|11|Dixit Moyses ad Aaron: " Tolle turibulum et, hausto igne de altari, mitte incensum desuper pergens cito ad populum, ut expies pro eis; iam enim egressa est ira a Domino, et plaga desaevit ".
NUM|17|12|Quod cum fecisset Aaron et cucurrisset ad mediam congregationem, quam iam vastabat plaga, obtulit thymiama et expiavit pro populo;
NUM|17|13|et stetit inter mortuos ac viventes, et plaga cessavit.
NUM|17|14|Fuerunt autem, qui percussi sunt, quattuordecim milia hominum et septingenti, absque his, qui perierant in seditione Core.
NUM|17|15|Reversusque est Aaron ad Moysen ad ostium tabernaculi conventus, postquam quievit interitus.
NUM|17|16|Et locutus est Dominus ad Moysen dicens:
NUM|17|17|" Loquere ad filios Israel et accipe ab eis virgas singulas per cognationes suas, a cunctis principibus tribuum virgas duodecim, et uniuscuiusque nomen superscribes virgae suae.
NUM|17|18|Nomen autem Aaron scribes in virga Levi, et una virga cunctas seorsum familias continebit.
NUM|17|19|Ponesque eas in tabernaculo conventus coram testimonio, ubi conveniam cum vobis.
NUM|17|20|Quem ex his elegero, germinabit virga eius; et cohibebo a me querimonias filiorum Israel, quibus contra vos murmurant ".
NUM|17|21|Locutusque est Moyses ad filios Israel, et dederunt ei omnes principes virgas per singulas tribus; fueruntque virgae duodecim, et virga Aaron in medio earum.
NUM|17|22|Quas cum posuisset Moyses coram Domino in tabernaculo testimonii,
NUM|17|23|sequenti die regressus invenit germinasse virgam Aaron in domo Levi; et turgentibus gemmis eruperant flores, qui, foliis dilatatis, in amygdalas deformati sunt.
NUM|17|24|Protulit ergo Moyses omnes virgas de conspectu Domini ad cunctos filios Israel; videruntque et receperunt singuli virgas suas.
NUM|17|25|Dixitque Dominus ad Moysen: " Refer virgam Aaron coram testimonio, ut servetur ibi in signum rebellium filiorum Israel, et quiescant querelae eorum a me, ne moriantur ".
NUM|17|26|Fecitque Moyses, sicut praeceperat Dominus.
NUM|17|27|Dixerunt autem filii Israel ad Moysen: " Ecce consumpti sumus, perimus, omnes perimus!
NUM|17|28|Quicumque accedit ad habitaculum Domini, moritur. Num usque ad internecionem cuncti delendi sumus? ".
NUM|18|1|Dixitque Dominus ad Aaron: " Tu et filii tui et domus patris tui tecum portabitis iniquitatem sanctuarii; et tu et filii tui simul sustinebitis peccata sacerdotii vestri.
NUM|18|2|Sed et fratres tuos de tribu Levi, tribum patris tui sume tecum, praestoque sint et ministrent tibi; tu autem et filii tui ministrabitis in tabernaculo testimonii.
NUM|18|3|Excubabuntque Levitae ad praecepta tua et ad cuncta opera tabernaculi, ita dumtaxat ut ad vasa sanctuarii et ad altare non accedant, ne et illi moriantur, et vos pereatis simul.
NUM|18|4|Sint autem tecum et excubent in custodiis tabernaculi conventus et in omni ministerio eius; alienigena non miscebitur vobis.
NUM|18|5|Excubate in ministerio sanctuarii et in ministerio altaris, ne oriatur amplius indignatio super filios Israel.
NUM|18|6|Ego sumpsi fratres vestros Levitas de medio filiorum Israel et tradidi donum Domino, ut serviant in ministeriis tabernaculi conventus.
NUM|18|7|Tu autem et filii tui custodite sacerdotium vestrum et omnia, quae ad cultum altaris pertinent et intra velum sunt, administrabitis. Ministerium do vobis sacerdotium in donum; si quis externus accesserit, occidetur ".
NUM|18|8|Locutusque est Dominus ad Aaron: " Ecce dedi tibi custodiam praelibationum mearum. Omnia, quae sanctificantur a filiis Israel, tradidi tibi et filiis tuis pro officio sacerdotali, legitima sempiterna.
NUM|18|9|Haec ergo accipies de sanctis sanctorum, exceptis his, quae comburuntur: omnis oblatio et sacrificium pro peccato atque delicto, quod redditur mihi, sanctum sanctorum tuum erit et filiorum tuorum.
NUM|18|10|In sanctuario comedes illud; mares tantum edent ex eo, quia consecratum est tibi.
NUM|18|11|Praelibationem donorum, quae elevando obtulerint filii Israel, tibi dedi et filiis tuis ac filiabus tuis iure perpetuo: qui mundus est in domo tua, vescetur eis.
NUM|18|12|Omnem medullam olei et vini ac frumenti quidquid offerunt primitiarum Domino, tibi dedi.
NUM|18|13|Universa frugum initia, quas gignit humus et Domino deportantur, cedent in usus tuos: qui mundus est in domo tua, vescetur eis.
NUM|18|14|Omne, quod ex voto reddiderint filii Israel, tuum erit.
NUM|18|15|Quidquid primum erumpit e vulva cunctae carnis, quod offerunt Domino, sive ex hominibus sive de pecoribus fuerit, tui iuris erit; ita dumtaxat, ut hominis primogenitum et omne animal, quod immundum est, redimi facias.
NUM|18|16|Cuius redemptio erit post unum mensem siclis argenti quinque pondere sanctuarii. Siclus viginti obolos habet.
NUM|18|17|Primogenitum autem bovis vel ovis vel caprae non facies redimi, quia sanctificata sunt Domino; sanguinem tantum eorum fundes super altare et adipes adolebis in suavissimum odorem Domino.
NUM|18|18|Carnes vero eorum in usum tuum cedent, sicut pectusculum elevatum et armus dexter tua erunt.
NUM|18|19|Omnes praelibationes sanctas, quas offerunt filii Israel Domino, tibi dedi et filiis ac filiabus tuis iure perpetuo: pactum salis est sempiternum coram Domino tibi ac filiis tuis ".
NUM|18|20|Dixitque Dominus ad Aaron: " In terra eorum nihil possidebitis nec habebitis partem inter eos: Ego pars et hereditas tua in medio filiorum Israel.
NUM|18|21|Filiis autem Levi dedi omnes decimas Israelis in possessionem pro ministerio, quo serviunt mihi in tabernaculo conventus,
NUM|18|22|ut non accedant ultra filii Israel ad tabernaculum conventus nec committant peccatum mortiferum.
NUM|18|23|Solis filiis Levi mihi in tabernaculo conventus servientibus et portantibus peccata populi; legitimum sempiternum erit in generationibus vestris, et in medio filiorum Israel nihil aliud possidebunt.
NUM|18|24|Decimas, quas filii Israel in praelibationem elevant Domino, dedi Levitis in possessionem. Propterea dixi eis: In medio filiorum Israel non habebitis possessionem ".
NUM|18|25|Locutusque est Dominus ad Moysen dicens:
NUM|18|26|" Praecipe Levitis atque denuntia: Cum acceperitis a filiis Israel decimas, quas dedi vobis, praelibationem earum elevabitis Domino, id est decimam partem decimae,
NUM|18|27|ut reputetur vobis in praelibationem tam de areis quam de torcularibus.
NUM|18|28|Sic de universis, quorum accipitis primitias a filiis Israel, elevate Domino: date Aaron sacerdoti.
NUM|18|29|Omnia, quae offeretis ex decimis, in donaria Domini separabitis: optima et electa erunt.
NUM|18|30|Dicesque ad eos: Si praeclara et meliora quaeque obtuleritis ex decimis, reputabitur vobis quasi de area et torculari dederitis fructus;
NUM|18|31|et comedetis eas in omnibus locis vestris, tam vos quam familiae vestrae, quia pretium est pro ministerio, quo servitis in tabernaculo conventus.
NUM|18|32|Et non peccabitis super hoc egregia vobis et pinguia reservantes, ne polluatis oblationes filiorum Israel et moriamini ".
NUM|19|1|Locutusque est Dominus ad Moysen et Aaron dicens:
NUM|19|2|" Ista est religio legis, quam constituit Dominus. Praecipe filiis Israel, ut adducant ad te vaccam rufam aetatis integrae, in qua nulla sit macula, nec portaverit iugum.
NUM|19|3|Tradetisque eam Eleazaro sacerdoti, quae educta extra castra mactabitur in conspectu eius;
NUM|19|4|et tinguens digitum in sanguine eius asperget contra fores tabernaculi conventus septem vicibus,
NUM|19|5|combureturque in conspectu eius, tam pelle et carnibus eius quam sanguine et fimo flammae traditis.
NUM|19|6|Lignum quoque cedrinum et hyssopum coccumque sacerdos mittet in flammam, quae vaccam vorat.
NUM|19|7|Et tunc demum, lotis vestibus et corpore suo, ingredietur in castra commaculatusque erit usque ad vesperum.
NUM|19|8|Sed et ille, qui combusserit eam, lavabit vestimenta sua et corpus, et immundus erit usque ad vesperum.
NUM|19|9|Colliget autem vir mundus cineres vaccae et effundet eos extra castra in loco purissimo, ut sint congregationi filiorum Israel in custodiam pro aqua aspersionis.
NUM|19|10|Cumque laverit, qui vaccae portaverat cineres, vestimenta sua, immundus erit usque ad vesperum. Habebunt hoc filii Israel et advenae, qui habitant inter eos, sanctum iure perpetuo.
NUM|19|11|Qui tetigerit cadaver hominis et propter hoc septem diebus fuerit immundus,
NUM|19|12|aspergetur ex hac aqua die tertio et septimo et sic mundabitur. Si die tertio aspersus non fuerit, septimo non erit mundus.
NUM|19|13|Omnis, qui tetigerit humanae animae morticinum et aspersus hac commixtione non fuerit, polluet habitaculum Domini et peribit ex Israel, quia aqua expiationis non est aspersus: immundus erit, et manebit spurcitia eius super eum.
NUM|19|14|Ista est lex hominis, qui moritur in tabernaculo: omnes, qui ingrediuntur tentorium illius, et universa vasa, quae ibi sunt, polluta erunt septem diebus.
NUM|19|15|Vas, quod non habuerit operculum nec ligaturam desuper, immundum erit.
NUM|19|16|Si quis in agro tetigerit cadaver hominis gladio occisi aut per se mortui sive os illius vel sepulcrum, immundus erit septem diebus.
NUM|19|17|Tollentque de cineribus combustionis peccati et mittent aquas vivas super eos in vas;
NUM|19|18|in quibus cum homo mundus tinxerit hyssopum, asperget ex eo omne tentorium et cunctam supellectilem et homines, qui ibi fuerint, et super eum, qui tetigerit ossa vel occisum hominem aut per se mortuum aut sepultum.
NUM|19|19|Atque hoc modo mundus lustrabit immundum tertio et septimo die; expiatusque die septimo lavabit et se et vestimenta sua et mundus erit ad vesperum.
NUM|19|20|Si quis hoc ritu non fuerit expiatus, peribit anima illius de medio ecclesiae, quia sanctuarium Domini polluit et non est aqua lustrationis aspersus; immundus est.
NUM|19|21|Erit vobis praeceptum legitimum sempiternum. Ipse quoque, qui aspergit aqua lustrali, lavabit vestimenta sua; omnis, qui tetigerit aquas expiationis, immundus erit usque ad vesperum.
NUM|19|22|Quidquid tetigerit immundus, immundum erit, et anima, quae horum quippiam tetigerit, immunda erit usque ad vesperum ".
NUM|20|1|Veneruntque filii Israel et omnis congregatio in de sertum Sin mense primo, et mansit populus in Cades. Mortuaque est ibi Maria et sepulta in eodem loco.
NUM|20|2|Cumque indigeret aqua populus, convenerunt adversum Moysen et Aaron
NUM|20|3|et versi in seditionem dixerunt: " Utinam perissemus inter fratres nostros coram Domino!
NUM|20|4|Cur eduxistis ecclesiam Domini in solitudinem, ut et nos et nostra iumenta moriamur?
NUM|20|5|Quare nos fecistis ascendere de Aegypto et adduxistis in locum istum pessimum, qui seri non potest, qui nec ficum gignit nec vineas nec malogranata, insuper et aquam non habet ad bibendum? ".
NUM|20|6|Venitque Moyses et Aaron, relicta congregatione, ad introitum tabernaculi conventus corrueruntque proni in terram, et apparuit gloria Domini super eos.
NUM|20|7|Locutusque est Dominus ad Moysen dicens:
NUM|20|8|" Tolle virgam et congrega populum, tu et Aaron frater tuus; et loquimini ad petram coram eis, et illa dabit aquas. Cumque eduxeris aquam de petra, potabis congregationem et iumenta eius ".
NUM|20|9|Tulit igitur Moyses virgam, quae erat in conspectu Domini, sicut praeceperat ei.
NUM|20|10|Et congregaverunt Moyses et Aaron populum ante petram, dixitque eis: " Audite, rebelles; num de petra hac vobis aquam poterimus eicere? ".
NUM|20|11|Cumque elevasset Moyses manum percutiens virga bis silicem, egressae sunt aquae largissimae, ita ut populus biberet et iumenta.
NUM|20|12|Dixitque Dominus ad Moysen et Aaron: " Quia non credidistis mihi, ut sanctificaretis me coram filiis Israel, non introducetis hos populos in terram, quam dabo eis ".
NUM|20|13|Hae sunt aquae Meriba, ubi iurgati sunt filii Israel contra Dominum, et sanctificatus est in eis.
NUM|20|14|Misit nuntios Moyses de Cades ad regem Edom, qui dicerent: " Haec mandat frater tuus Israel: Nosti omnem laborem, qui apprehendit nos,
NUM|20|15|quomodo descenderint patres nostri in Aegyptum, et habitaverimus ibi multo tempore, afflixerintque nos Aegyptii et patres nostros,
NUM|20|16|et quomodo clamaverimus ad Dominum, et exaudierit nos miseritque angelum, qui eduxerit nos de Aegypto. Ecce nos in urbe Cades, quae est in extremis finibus tuis, positi
NUM|20|17|obsecramus, ut nobis transire liceat per terram tuam: non ibimus per agros nec per vineas, non bibemus aquas de puteis tuis; sed gradiemur via regia, nec ad dexteram nec ad sinistram declinantes, donec transeamus terminos tuos ".
NUM|20|18|Cui respondit Edom: " Non transibis per me, alioquin armatus occurram tibi ".
NUM|20|19|Dixeruntque filii Israel: " Per tritam gradiemur viam et, si biberimus aquas tuas ego et pecora mea, dabo, quod iustum est: nulla erit in pretio difficultas; tantum velociter transeamus ".
NUM|20|20|At ille respondit: " Non transibis! ". Statimque egressus est obvius cum infinita multitudine et manu forti
NUM|20|21|nec voluit acquiescere Israeli, ut concederet transitum per fines suos; quam ob rem divertit ab eo Israel.
NUM|20|22|Cumque castra movissent de Cades, venerunt in montem Hor,
NUM|20|23|ubi locutus est Dominus ad Moysen et Aaron in monte Hor, qui est in finibus terrae Edom:
NUM|20|24|" Congregabitur, inquit, Aaron ad populum suum. Non enim intrabit terram, quam dedi filiis Israel, eo quod rebelles fuistis ori meo ad aquas Meriba.
NUM|20|25|Tolle Aaron et Eleazarum filium eius cum eo et duces eos in montem Hor.
NUM|20|26|Cumque nudaveris patrem veste sua, indues ea Eleazarum filium eius: Aaron colligetur et morietur ibi ".
NUM|20|27|Fecit Moyses, ut praeceperat Dominus, et ascenderunt in montem Hor coram omni congregatione.
NUM|20|28|Cumque Aaron spoliasset vestibus suis, induit eis Eleazarum filium eius. Illo mortuo in montis supercilio, descendit cum Eleazaro.
NUM|20|29|Omnis autem congregatio videns occubuisse Aaron flevit super eo triginta diebus tota domus Israel.
NUM|21|1|Quod cum audisset Chana naeus rex Arad, qui habita bat in Nageb, venisse scilicet Israel per viam Atarim, pugnavit contra illum et duxit ex eo captivos.
NUM|21|2|At Israel voto se Domino obligans ait: " Si tradideris populum istum in manu mea, delebo urbes eius ".
NUM|21|3|Exaudivitque Dominus preces Israel et tradidit Chananaeum, quem ille interfecit, subversis urbibus eius, et vocavit nomen loci illius Horma.
NUM|21|4|Profecti sunt autem et de monte Hor per viam, quae ducit ad mare Rubrum, ut circumirent terram Edom. Et taedere coepit populum itineris.
NUM|21|5|Locutusque contra Deum et Moysen ait: " Cur eduxisti nos de Aegypto, ut moreremur in solitudine? Deest panis, non sunt aquae; anima nostra iam nauseat super cibo isto levissimo ".
NUM|21|6|Quam ob rem misit Dominus in populum ignitos serpentes, qui mordebant populum, et mortuus est populus multus ex Israel.
NUM|21|7|Et venerunt ad Moysen atque dixerunt: " Peccavimus, quia locuti sumus contra Dominum et te; ora, ut tollat a nobis serpentes ". Oravitque Moyses pro populo.
NUM|21|8|Et locutus est Dominus ad eum: " Fac serpentem ignitum et pone eum pro signo: qui percussus aspexerit eum, vivet ".
NUM|21|9|Fecit ergo Moyses serpentem aeneum et posuit eum pro signo; quem cum percussi aspicerent, sanabantur.
NUM|21|10|Profectique filii Israel castrametati sunt in Oboth,
NUM|21|11|unde egressi fixere tentoria in Ieabarim, in solitudine, quae respicit Moab contra orientalem plagam.
NUM|21|12|Et inde moventes venerunt ad torrentem Zared;
NUM|21|13|quem relinquentes castrametati sunt ultra Arnon, qui est in deserto, quod prominet de finibus Amorraei. Siquidem Arnon terminus est Moab dividens Moabitas et Amorraeos.
NUM|21|14|Unde dicitur in libro bellorum Domini:" Vaheb in Suphaet torrentes Arnon.
NUM|21|15|Scopuli torrentium inclinati suntin habitationem Aret recumbunt in finibus Moabitarum ".
NUM|21|16|Ex eo loco in Beer. Hic est puteus, super quo locutus est Dominus ad Moysen: " Congrega populum, et dabo ei aquam ".
NUM|21|17|Tunc cecinit Israel carmen istud:" Ascendat puteus. Concinite ei.
NUM|21|18|Puteus, quem foderunt principeset paraverunt duces populiin sceptris et in baculis suis ".De solitudine in Matthana;
NUM|21|19|de Matthana in Nahaliel; de Nahaliel in Bamoth;
NUM|21|20|de Bamoth in vallem, quae est in regione Moab in vertice Phasga, qui respicit contra desertum.
NUM|21|21|Misit autem Israel nuntios ad Sehon regem Amorraeorum dicens:
NUM|21|22|" Obsecro, ut transire mihi liceat per terram tuam: non declinabimus in agros et vineas, non bibemus aquas ex puteis. Via regia gradiemur, donec transeamus terminos tuos ".
NUM|21|23|Qui concedere noluit, ut transiret Israel per fines suos; quin potius, populo congregato, egressus est obviam in desertum et venit in Iasa pugnavitque contra Israel.
NUM|21|24|A quo percussus est in ore gladii, et possessa est terra eius ab Arnon usque Iaboc et filios Ammon; quia forti praesidio tenebantur termini Ammonitarum.
NUM|21|25|Tulit ergo Israel omnes civitates eius et habitavit in urbibus Amorraei, in Hesebon scilicet et viculis eius.
NUM|21|26|Hesebon enim erat urbs Sehon regis Amorraei, qui pugnavit contra primum regem Moab et tulit omnem terram, quae dicionis illius fuerat usque Arnon.
NUM|21|27|Idcirco dicitur in proverbio:" Venite in Hesebon!Aedificetur et construatur civitas Sehon!
NUM|21|28|Ignis egressus est de Hesebon,flamma de oppido Sehonet devoravit Ar Moabitarumet deglutivit excelsa Arnon.
NUM|21|29|Vae tibi, Moab;peristi, popule Chamos!Dedit filios eius in fugamet filias in captivitatemregi Amorraeorum Sehon.
NUM|21|30|Iecimus sagittas in eos,disperiit Hesebon usque Dibon.Vastavimus usque Nopheet usque Medaba ".
NUM|21|31|Habitavit itaque Israel in terra Amorraei.
NUM|21|32|Misitque Moyses, qui explorarent Iazer, cuius ceperunt viculos et expulerunt Amorraeos, qui erant ibi.
NUM|21|33|Verteruntque se et ascenderunt per viam Basan, et occurrit eis Og rex Basan cum omni populo suo pugnaturus in Edrai.
NUM|21|34|Dixitque Dominus ad Moysen: " Ne timeas eum, quia in manu tua tradidi illum et omnem populum ac terram eius, faciesque illi, sicut fecisti Sehon regi Amorraeorum habitatori Hesebon ".
NUM|21|35|Percusserunt igitur et hunc cum filiis suis universumque populum eius usque ad internecionem; et possederunt terram illius.
NUM|22|1|Profectique castrametati sunt filii Israel in campestri bus Moab, ubi trans Iordanem Iericho sita est.
NUM|22|2|Videns autem Balac filius Sephor omnia, quae fecerat Israel Amorraeo,
NUM|22|3|valde metuit Moab populum, quia multus erat. Et cum pertimeret Moab filios Israel,
NUM|22|4|dixit ad maiores natu Madian: " Nunc carpet haec congregatio omnem regionem per circuitum, quomodo solet bos herbas campi carpere ".Balac filius Sephor erat eo tempore rex in Moab.
NUM|22|5|Misit ergo nuntios ad Balaam filium Beor in Phethor, quae est super flumen in terra filiorum Ammau, ut vocarent eum et dicerent: " Ecce egressus est populus ex Aegypto, qui operuit superficiem terrae sedens contra me.
NUM|22|6|Veni igitur et maledic populo huic, quia fortior me est; si quo modo possim percutere et eicere eum de terra mea. Novi enim quod benedictus sit, cui benedixeris, et maledictus, in quem maledicta congesseris ".
NUM|22|7|Perrexeruntque seniores Moab et maiores natu Madian habentes divinationis pretium in manibus. Cumque venissent ad Balaam et narrassent ei omnia verba Balac,
NUM|22|8|ille respondit: " Manete hic nocte, et respondebo quidquid mihi dixerit Dominus ". Manentibus illis apud Balaam,
NUM|22|9|venit Deus et ait ad eum: " Quid sibi volunt homines isti apud te? ".
NUM|22|10|Respondit: " Balac filius Sephor rex Moabitarum misit ad me
NUM|22|11|dicens: "Ecce populus, qui egressus est de Aegypto, operuit superficiem terrae; veni et maledic ei pro me, si quo modo possim pugnans abigere eum".
NUM|22|12|Dixitque Deus ad Balaam: "Noli ire cum eis neque maledicas populo, quia benedictus est ".
NUM|22|13|Qui mane consurgens dixit ad principes: " Ite in terram vestram, quia prohibuit me Dominus venire vobiscum ".
NUM|22|14|Reversi principes dixerunt ad Balac: " Noluit Balaam venire nobiscum ".
NUM|22|15|Rursum ille multo plures et nobiliores, quam ante miserat, misit.
NUM|22|16|Qui cum venissent ad Balaam, dixerunt: " Sic dicit Balac filius Sephor: "Ne cuncteris venire ad me;
NUM|22|17|paratus sum honorare te et, quidquid volueris, dabo tibi. Veni et maledic pro me populo isti" ".
NUM|22|18|Respondit Balaam: " Si dederit mihi Balac plenam domum suam argenti et auri, non potero transgredi verbum Domini Dei mei, ut vel plus vel minus loquar.
NUM|22|19|Obsecro, ut hic maneatis etiam hac nocte, et scire queam quid mihi rursum respondeat Dominus ".
NUM|22|20|Venit ergo Deus ad Balaam nocte et ait ei: " Si vocare te venerunt homines isti, surge et vade cum eis, ita dumtaxat, ut, quod tibi praecepero, facias ".
NUM|22|21|Surrexit Balaam mane et, strata asina sua, profectus est cum eis.
NUM|22|22|Et iratus est Deus, cum profectus esset; stetitque angelus Domini in via contra Balaam, ut adversaretur ei, qui insidebat asinae et duos pueros habebat secum.
NUM|22|23|Cernens asina angelum Domini stantem in via, evaginato gladio in manu sua, avertit se de itinere et ibat per agrum. Quam cum verberaret Balaam et vellet ad semitam reducere,
NUM|22|24|stetit angelus Domini in angustiis duarum maceriarum, quibus vineae cingebantur.
NUM|22|25|Quem videns asina iunxit se parieti et attrivit sedentis pedem. At ille iterum verberabat eam;
NUM|22|26|et angelus Domini iterum transiens ad locum angustum, ubi nec ad dexteram nec ad sinistram poterat deviare, obvius stetit.
NUM|22|27|Cumque vidisset asina stantem angelum Domini, concidit sub pedibus sedentis; qui iratus vehementius caedebat fuste latera eius.
NUM|22|28|Aperuitque Dominus os asinae, et locuta est: " Quid feci tibi? Cur percutis me ecce iam tertio? ".
NUM|22|29|Respondit Balaam: " Quia illusisti mihi. Utinam haberem gladium, ut te interficerem! ".
NUM|22|30|Dixit asina: " Nonne animal tuum sum, cui semper sedere consuevisti usque in praesentem diem? Dic quid simile umquam fecerim tibi ". At ille ait: " Numquam ".
NUM|22|31|Protinus aperuit Dominus oculos Balaam, et vidit angelum Domini stantem in via, evaginato gladio in manu eius; adoravitque eum pronus in terram.
NUM|22|32|Cui angelus Domini: " Cur, inquit, tertio verberas asinam tuam? Ego veni, ut adversarer tibi, quia perversa est via tua mihique contraria.
NUM|22|33|Et videns me asina declinavit ter a me; nisi declinasset, te occidissem et illam vivam reliquissem ".
NUM|22|34|Dixit Balaam: " Peccavi nesciens quod tu stares contra me in via; et nunc, si displicet tibi, revertar ".
NUM|22|35|Ait angelus Domini: " Vade cum istis et cave, ne aliud, quam praecepero tibi, loquaris ". Ivit igitur cum principibus Balac.
NUM|22|36|Quod cum audisset Balac, venisse scilicet Balaam, egressus est in occursum eius in Irmoab, quod situm est in extremis finibus Arnon;
NUM|22|37|dixitque ad Balaam: " Nonne misi nuntios, ut vocarem te? Cur non statim venisti ad me? An quia honorare te nequeo? ".
NUM|22|38|Cui ille respondit: " Ecce adsum; numquid loqui potero aliud, nisi quod Deus posuerit in ore meo? ".
NUM|22|39|Perrexerunt ergo simul et venerunt in Cariathusoth.
NUM|22|40|Cumque occidisset Balac boves et oves, misit ad Balaam et principes, qui cum eo erant.
NUM|22|41|Mane autem facto, duxit eum ad excelsa Baal et intuitus est extremam partem populi.
NUM|23|1|Dixitque Balaam ad Balac: " Aedifica mihi hic septem aras et para totidem vitulos eiusdemque numeri arietes ".
NUM|23|2|Cumque fecisset iuxta sermonem Balaam, imposuerunt vitulum et arietem super aram.
NUM|23|3|Dixitque Balaam ad Balac: " Sta paulisper iuxta holocaustum tuum, donec vadam, si forte occurrat mihi Dominus; et, quodcumque imperaverit, loquar tibi ". Cumque abiisset in collem nudum,
NUM|23|4|occurrit illi Deus. Locutusque ad eum Balaam: " Septem, inquit, aras erexi et imposui vitulum et arietem desuper ".
NUM|23|5|Dominus autem posuit verbum in ore eius et ait: " Revertere ad Balac et haec loqueris ".
NUM|23|6|Reversus invenit stantem Balac iuxta holocaustum suum et omnes principes Moabitarum;
NUM|23|7|assumptaque parabola sua, dixit:" De Aram adduxit me Balac,rex Moabitarum de montibus orientis:"Veni, inquit, et maledic pro me Iacob;propera et detestare Israel!".
NUM|23|8|Quomodo maledicam, cui non maledixit Deus?Qua ratione detester, quem Dominus non detestatur?
NUM|23|9|De summis silicibus video eumet de collibus considero illum:populus solus habitabitet inter gentes non reputabitur.
NUM|23|10|Et quis dinumerare possit pulverem Iacobet quis numeravit arenam Israel?Moriatur anima mea morte iustorum,et fiant novissima mea horum similia ".
NUM|23|11|Dixitque Balac ad Balaam: " Quid est hoc, quod agis? Ut malediceres inimicis meis, vocavi te, et tu e contrario benedicis eis! ".
NUM|23|12|Cui ille respondit: " Num aliud possum loqui, nisi quod iusserit Dominus? ".
NUM|23|13|Dixit ergo Balac: " Veni mecum in alterum locum, unde partem Israel videas et totum videre non possis; inde maledicito ei ".
NUM|23|14|Cumque duxisset eum in campum speculatorum super verticem montis Phasga, aedificavit septem aras imposuitque supra vitulum atque arietem.
NUM|23|15|Et dixit Balaam ad Balac: " Sta hic iuxta holocaustum tuum, donec ego obvius pergam ".
NUM|23|16|Cui cum Dominus occurrisset posuissetque verbum in ore eius, ait: " Revertere ad Balac et haec loqueris ei ".
NUM|23|17|Reversus invenit eum stantem iuxta holocaustum suum et principes Moabitarum cum eo. Ad quem Balac: " Quid, inquit, locutus est Dominus? ".
NUM|23|18|At ille, assumpta parabola sua, ait:" Surge, Balac, et ausculta;audi, fili Sephor.
NUM|23|19|Non est Deus quasi homo, ut mentiatur,nec ut filius hominis, ut mutetur.Numquid dixit et non faciet?Locutus est et non implebit?
NUM|23|20|Ad benedicendum adductus sum,benedictionem prohibere non valeo.
NUM|23|21|Non conspicitur malum in Iacob,nec videtur calamitas in Israel.Dominus Deus eius cum eo est,et clangor regis in illo.
NUM|23|22|Deus eduxit illum de Aegypto,sicut cornua bubali est ei.
NUM|23|23|Non est augurium in Iacob,nec divinatio in Israel.Temporibus suis dicetur Iacob et Israeliquid operatus sit Deus.
NUM|23|24|Ecce populus ut leaena consurget,et quasi leo erigetur;non accubabit, donec devoret praedamet occisorum sanguinem bibat ".
NUM|23|25|Dixitque Balac ad Balaam: " Nec maledicas ei, nec benedicas! ".
NUM|23|26|Et ille ait: " Nonne dixi tibi quod, quidquid mihi Dominus imperaret, hoc facerem? ".
NUM|23|27|Et ait Balac ad eum: " Veni, et ducam te ad alîum locum, si forte placeat Deo, ut inde maledicas ei ".
NUM|23|28|Cumque duxisset eum super verticem montis Phegor, qui respicit solitudinem,
NUM|23|29|dixit ei Balaam: " Aedifica mihi hic septem aras et para totidem vitulos eiusdemque numeri arietes ".
NUM|23|30|Fecit Balac, ut Balaam dixerat, imposuitque vitulos et arietes per singulas aras.
NUM|24|1|Cumque vidisset Balaam quod placeret Domino, ut be nediceret Israeli, nequaquam abiit, ut ante perrexerat, ut augurium quaereret; sed dirigens contra desertum vultum suum
NUM|24|2|et elevans oculos vidit Israel commorantem per tribus suas et, irruente in se spiritu Dei,
NUM|24|3|assumpta parabola sua, ait:" Dixit Balaam filius Beor,dixit homo, cuius apertus est oculus,
NUM|24|4|dixit auditor sermonum Dei,qui visionem Omnipotentis intuitus est,qui cadit, et sic aperiuntur oculi eius.
NUM|24|5|Quam pulchra tabernacula tua, Iacob,et tentoria tua, Israel!
NUM|24|6|Ut valles dilatantur,ut horti iuxta fluvios irrigui,ut aloe, quam plantavit Dominus,quasi cedri prope aquas.
NUM|24|7|Fluet aqua de situlis eius,et semen illius erit in aquis multis. Extolletur super Agag rex eius,et elevabitur regnum illius.
NUM|24|8|Deus eduxit illum de Aegypto,sicut cornua bubali est ei.Devorabit gentes, hostes suos,ossaque eorum confringetet perforabit sagittis.
NUM|24|9|Accubans dormit ut leo,et quasi leaena, quis suscitare illum audebit?Qui benedixerit tibi, erit et ipse benedictus;qui maledixerit tibi, maledictus erit! ".
NUM|24|10|Iratusque Balac contra Balaam, complosis manibus, ait: " Ad maledicendum inimicis meis vocavi te, quibus iam tertio benedixisti!
NUM|24|11|Revertere nunc ad locum tuum! Decreveram quidem magnifice honorare te, sed Dominus privavit te honore disposito ".
NUM|24|12|Respondit Balaam ad Balac: " Nonne iam nuntiis tuis, quos misisti ad me, dixi:
NUM|24|13|Si dederit mihi Balac plenam domum suam argenti et auri, non potero praeterire sermonem Domini, ut vel boni quid vel mali proferam ex corde meo, sed, quidquid Dominus dixerit, hoc loquar?
NUM|24|14|Et nunc, pergens ad populum meum dabo consilium, quid populus hic populo tuo faciat extremo tempore ".
NUM|24|15|Sumpta igitur parabola sua, rursum ait:" Dixit Balaam filius Beor,dixit homo, cuius apertus est oculus,
NUM|24|16|dixit auditor sermonum Dei,qui novit doctrinam Altissimiet visiones Omnipotentis videt,qui cadens apertos habet oculos.
NUM|24|17|Video eum, sed non modo;intueor illum, sed non prope.Oritur stella ex Iacob,et consurgit virga de Israel;et percutit tempora Moabet verticem omnium filiorum Seth.
NUM|24|18|Et erit Idumaea possessio eius,et hereditas eius Seir, inimicus eius; Israel vero fortiter aget.
NUM|24|19|De Iacob erit, qui domineturet perdat reliquias civitatis ".
NUM|24|20|Cumque vidisset Amalec, assumens parabolam suam ait:" Principium gentium Amalec,cuius extrema perdentur ".
NUM|24|21|Vidit quoque Cinaeum et, assumpta parabola sua, ait:" Robustum quidem est habitaculum tuum,et in petra positus nidus tuus.
NUM|24|22|Erit in combustionem Cain,donec Assur capiat te ".
NUM|24|23|Assumptaque parabola sua, iterum locutus est:" Heu! Quis vivet,quando ista faciet Deus?
NUM|24|24|Venient naves de Cetthim,superabunt Assyrios vastabuntque Heber;et ad extremum etiam ipsi peribunt ".Surrexitque Balaam et reversus est in locum suum; Balac quoque via, qua venerat, rediit.
NUM|25|1|Morabatur autem Israel in Settim, et incepit populus fornicari cum filiabus Moab,
NUM|25|2|quae vocaverunt populum ad sacrificia deorum suorum. Et illi comederunt et adoraverunt deos earum;
NUM|25|3|et adhaesit Israel Baalphegor. Et iratus Dominus
NUM|25|4|ait ad Moysen: " Tolle cunctos principes populi et suspende eos coram Domino contra solem in patibulis, ut avertatur furor meus ab Israel ".
NUM|25|5|Dixitque Moyses ad iudices Israel: " Occidat unusquisque proximos suos, qui adhaeserunt Baalphegor ".
NUM|25|6|Et ecce unus de filiis Israel intravit coram fratribus suis ad Madianitin, vidente Moyse et omni turba filiorum Israel, qui flebant ante fores tabernaculi conventus.
NUM|25|7|Quod cum vidisset Phinees filius Eleazari filii Aaron sacerdotis, surrexit de medio congregationis et, arrepta lancea,
NUM|25|8|ingressus est post virum Israelitem in cubiculum et perfodit ambos simul, virum scilicet et mulierem, in locis genitalibus; cessavitque plaga a filiis Israel.
NUM|25|9|Et occisi sunt viginti quattuor milia hominum.
NUM|25|10|Dixitque Dominus ad Moysen:
NUM|25|11|" Phinees filius Eleazari filii Aaron sacerdotis avertit iram meam a filiis Israel, quia zelo meo commotus est in medio eorum, ut non ipse delerem filios Israel in zelo meo.
NUM|25|12|Idcirco loquere ad eum: Ecce do ei pacem foederis mei,
NUM|25|13|et erit tam ipsi quam semini eius pactum sacerdotii sempiternum, quia zelatus est pro Deo suo et expiavit scelus filiorum Israel ".
NUM|25|14|Erat autem nomen viri Israelitae, qui occisus est cum Madianitide, Zamri filius Salu dux de cognatione et tribu Simeonis;
NUM|25|15|porro mulier Madianitis, quae pariter interfecta est, vocabatur Cozbi filia Sur principis tribus in Madian.
NUM|25|16|Locutusque est Dominus ad Moysen dicens:
NUM|25|17|" Pugnate contra Madianitas et percutite eos,
NUM|25|18|quia ipsi hostiliter egerunt contra vos et decepere insidiis per idolum Phegor et in negotio Cozbi filiae ducis Madian sororis eorum, quae percussa est in die plagae pro sacrilegio Phegor ".
NUM|26|1|Post hanc plagam dixit Do minus ad Moysen et Eleaza rum filium Aaron sacerdotem:
NUM|26|2|" Numerate summam totius congregationis filiorum Israel a viginti annis et supra per domos et cognationes suas, cunctos, qui possunt ad bella procedere ".
NUM|26|3|Locuti sunt itaque Moyses et Eleazar sacerdos in campestribus Moab super Iordanem contra Iericho ad eos, qui erant
NUM|26|4|a viginti annis et supra, sicut Dominus imperaverat Moysi.Filiorum Israel, qui egressi sunt de terra Aegypti, iste est numerus.
NUM|26|5|Ruben primogenitus Israel. Huius filius Henoch, a quo familia Henochitarum, et Phallu, a quo familia Phalluitarum,
NUM|26|6|et Hesron, a quo familia Hesronitarum, et Charmi, a quo familia Charmitarum.
NUM|26|7|Hae sunt familiae de stirpe Ruben, quarum numerus inventus est quadraginta tria milia et septingenti triginta.
NUM|26|8|Filius Phallu: Eliab.
NUM|26|9|Huius filii: Namuel et Dathan et Abiram. Isti sunt Dathan et Abiram principes populi, qui surrexerunt contra Moysen et Aaron in seditione Core, quando adversus Dominum rebellaverunt,
NUM|26|10|et aperiens terra os suum devoravit eos et Core, morientibus plurimis, quando combussit ignis ducentos quinquaginta viros; et facti sunt in signum.
NUM|26|11|Core pereunte, filii illius non perierunt.
NUM|26|12|Filii Simeon per cognationes suas: Namuel, ab hoc familia Namuelitarum; Iamin, ab hoc familia Iaminitarum; Iachin, ab hoc familia Iachinitarum;
NUM|26|13|Zara, ab hoc familia Zaraitarum; Saul, ab hoc familia Saulitarum.
NUM|26|14|Hae sunt familiae de stirpe Simeon, quarum omnis numerus fuit viginti duo milia ducenti.
NUM|26|15|Filii Gad per cognationes suas: Sephon, ab hoc familia Sephonitarum; Haggi, ab hoc familia Haggitarum; Suni, ab hoc familia Sunitarum;
NUM|26|16|Ozni, ab hoc familia Oznitarum; Heri, ab hoc familia Heritarum;
NUM|26|17|Arodi, ab hoc familia Aroditarum; Areli, ab hoc familia Arelitarum.
NUM|26|18|Istae sunt familiae Gad, quarum omnis numerus fuit quadraginta milia quingenti.
NUM|26|19|Filii Iudae Her et Onan, qui ambo mortui sunt in terra Chanaan.
NUM|26|20|Fueruntque filii Iudae per cognationes suas: Sela, a quo familia Selanitarum; Phares, a quo familia Pharesitarum; Zara, a quo familia Zaraitarum.
NUM|26|21|Porro filii Phares: Esrom, a quo familia Esromitarum; et Hamul, a quo familia Hamulitarum.
NUM|26|22|Istae sunt familiae Iudae, quarum omnis numerus fuit septuaginta sex milia quingenti.
NUM|26|23|Filii Issachar per cognationes suas: Thola, a quo familia Tholaitarum; Phua, a quo familia Phuaitarum;
NUM|26|24|Iasub, a quo familia Iasubitarum; Semron, a quo familia Semronitarum.
NUM|26|25|Hae sunt cognationes Issachar, quarum numerus fuit sexaginta quattuor milia trecenti.
NUM|26|26|Filii Zabulon per cognationes suas: Sared, a quo familia Sareditarum; Elon, a quo familia Elonitarum; Iahelel, a quo familia Iahelelitarum.
NUM|26|27|Hae sunt cognationes Zabulon, quarum numerus fuit sexaginta milia quingenti.
NUM|26|28|Filii Ioseph per cognationes suas: Manasse et Ephraim.
NUM|26|29|De Manasse ortus est Machir, a quo familia Machiritarum; Machir genuit Galaad, a quo familia Galaaditarum.
NUM|26|30|Galaad habuit filios: Iezer, a quo familia Iezeritarum; et Helec, a quo familia Helecitarum;
NUM|26|31|et Asriel, a quo familia Asrielitarum; et Sechem, a quo familia Sechemitarum;
NUM|26|32|et Semida, a quo familia Semidaitarum; et Hepher, a quo familia Hepheritarum.
NUM|26|33|Fuit autem Hepher pater Salphaad, qui filios non habebat sed tantum filias, quarum ista sunt nomina: Maala et Noa et Hegla et Melcha et Thersa.
NUM|26|34|Hae sunt familiae Manasse, et numerus earum quinquaginta duo milia septingenti.
NUM|26|35|Filii autem Ephraim per cognationes suas fuerunt hi: Suthala, a quo familia Suthalaitarum; Becher, a quo familia Becheritarum; Thehen, a quo familia Thehenitarum.
NUM|26|36|Porro filius Suthala fuit Heran, a quo familia Heranitarum.
NUM|26|37|Hae sunt cognationes filiorum Ephraim, quarum numerus fuit triginta duo milia quingenti. Isti sunt filii Ioseph per familias suas.
NUM|26|38|Filii Beniamin in cognationibus suis: Bela, a quo familia Belaitarum; Asbel, a quo familia Asbelitarum; Ahiram, a quo familia Ahiramitarum;
NUM|26|39|Supham, a quo familia Suphamitarum; Hupham, a quo familia Huphamitarum.
NUM|26|40|Filii Bela: Ared et Naaman; de Ared familia Areditarum, de Naaman familia Naamanitarum.
NUM|26|41|Hi sunt filii Beniamin per cognationes suas, quorum numerus fuit quadraginta quinque milia sescenti.
NUM|26|42|Filii Dan per cognationes suas: Suham, a quo familia Suhamitarum. Hae sunt cognationes Dan per familias suas:
NUM|26|43|omnes fuere Suhamitae, quorum numerus erat sexaginta quattuor milia quadringenti.
NUM|26|44|Filii Aser per cognationes suas: Iemna, a quo familia Iemnaitarum; Isui, a quo familia Isuitarum; Beria, a quo familia Beriaitarum.
NUM|26|45|Filii Beria: Heber, a quo familia Heberitarum, et Melchiel a quo familia Melchielitarum.
NUM|26|46|Nomen autem filiae Aser fuit Sara.
NUM|26|47|Hae cognationes filiorum Aser, et numerus eorum quinquaginta tria milia quadringenti.
NUM|26|48|Filii Nephthali per cognationes suas: Iasiel, a quo familia Iasielitarum; Guni, a quo familia Gunitarum;
NUM|26|49|Ieser, a quo familia Ieseritarum; Sellem, a quo familia Sellemitarum.
NUM|26|50|Hae sunt cognationes filiorum Nephthali per familias suas, quorum numerus quadraginta quinque milia quadringenti.
NUM|26|51|Ista est summa filiorum Israel qui recensiti sunt: sescenta milia et mille septingenti triginta.
NUM|26|52|Locutusque est Dominus ad Moysen dicens:
NUM|26|53|" Istis dividetur terra iuxta numerum vocabulorum in possessiones suas.
NUM|26|54|Pluribus maiorem partem dabis et paucioribus minorem: singulis, sicut nunc recensiti sunt, tradetur possessio;
NUM|26|55|ita dumtaxat, ut sors terram dividat. Secundum numerum tribuum patrum suorum hereditabunt.
NUM|26|56|Quidquid sorte contigerit, hoc vel plures accipiant vel pauciores.
NUM|26|57|Hic quoque est numerus filiorum Levi per familias suas: Gerson, a quo familia Gersonitarum; Caath, a quo familia Caathitarum; Merari, a quo familia Meraritarum.
NUM|26|58|Hae sunt familiae Levi: familia Lobni, familia Hebroni, familia Moholi, familia Musi, familia Core. At vero Caath genuit Amram,
NUM|26|59|qui habuit uxorem Iochabed filiam Levi, quae nata est ei in Aegypto. Haec genuit Amram viro suo filios, Aaron et Moysen et Mariam sororem eorum.
NUM|26|60|De Aaron orti sunt Nadab et Abiu et Eleazar et Ithamar,
NUM|26|61|quorum Nadab et Abiu mortui sunt, cum obtulissent ignem alienum coram Domino.
NUM|26|62|Fueruntque omnes, qui numerati sunt, viginti tria milia generis masculini ab uno mense et supra; quia non sunt recensiti inter filios Israel, nec eis cum ceteris data possessio est.
NUM|26|63|Hic est numerus filiorum Israel, qui descripti sunt a Moyse et Eleazaro sacerdote in campestribus Moab supra Iordanem contra Iericho;
NUM|26|64|inter quos nullus fuit eorum, qui ante numerati sunt a Moyse et Aaron in deserto Sinai:
NUM|26|65|praedixerat enim Dominus quod omnes morerentur in solitudine; nullusque remansit ex eis, nisi Chaleb filius Iephonne et Iosue filius Nun.
NUM|27|1|Accesserunt autem filiae Sal phaad filii Hepher filii Ga laad filii Machir filii Manasse, e cognationibus Manasse, qui fuit filius Ioseph, quarum sunt nomina: Maala et Noa et Hegla et Melcha et Thersa.
NUM|27|2|Steteruntque coram Moyse et Eleazaro sacerdote et principibus et cuncta congregatione ad ostium tabernaculi conventus atque dixerunt:
NUM|27|3|" Pater noster mortuus est in deserto, nec fuit in seditione, quae concitata est contra Dominum sub Core, sed in peccato suo mortuus est; hic non habuit mares filios.
NUM|27|4|Cur tollitur nomen illius de familia sua, quia non habuit filium? Date nobis possessionem inter fratres patris nostri ".
NUM|27|5|Rettulitque Moyses causam earum ad iudicium Domini,
NUM|27|6|qui dixit ad eum:
NUM|27|7|" Iustam rem postulant filiae Salphaad. Da eis possessionem inter fratres patris sui, et ei in hereditatem succedant.
NUM|27|8|Ad filios autem Israel loqueris haec: Homo cum mortuus fuerit absque filio, ad filiam eius transibit hereditas;
NUM|27|9|si filiam non habuerit, habebit successores fratres suos.
NUM|27|10|Quod si et fratres non fuerint, dabitis hereditatem fratribus patris eius.
NUM|27|11|Sin autem nec patruos habuerit, dabitur hereditas illi, qui ei proximus est e cognatione sua; possidebitque eam. Eritque hoc filiis Israel sanctum lege perpetua, sicut praecepit Dominus Moysi ".
NUM|27|12|Dixit quoque Dominus ad Moysen: " Ascende in montem istum Abarim et contemplare inde terram, quam daturus sum filiis Israel.
NUM|27|13|Cumque videris eam, ibis et tu ad populum tuum, sicut ivit frater tuus Aaron,
NUM|27|14|quia offendistis me in deserto Sin in contradictione congregationis, nec sanctificare me voluistis coram ea super aquas ". Hae sunt aquae Meribathcades deserti Sin.
NUM|27|15|Cui respondit Moyses:
NUM|27|16|" Provideat Dominus, Deus spirituum omnis carnis, hominem, qui sit super congregationem hanc
NUM|27|17|et possit exire et intrare ante eos et educere eos vel introducere, ne sit populus Domini sicut oves absque pastore ".
NUM|27|18|Dixitque Dominus ad eum: " Tolle Iosue filium Nun, virum in quo est spiritus; et pone manum tuam super eum,
NUM|27|19|quem statues coram Eleazaro sacerdote et omni congregatione et dabis ei praecepta, cunctis videntibus,
NUM|27|20|et partem gloriae tuae, ut audiat eum omnis synagoga filiorum Israel.
NUM|27|21|Stabit coram Eleazaro sacerdote, qui pro eo iudicium Urim consulet Dominum. Ad verbum eius egredietur et ingredietur ipse et omnes filii Israel cum eo, cuncta congregatio ".
NUM|27|22|Fecit Moyses, ut praeceperat Dominus. Cumque tulisset Iosue, statuit eum coram Eleazaro sacerdote et omni frequentia populi;
NUM|27|23|et, impositis capiti eius manibus, constituit eum, sicut mandaverat Dominus per manum Moysi.
NUM|28|1|Dixit quoque Dominus ad Moysen:
NUM|28|2|" Praecipe filiis Is rael et dices ad eos: Oblationem meam et panem meum, sacrificium ignis in odorem suavissimum offerte per tempora sua.
NUM|28|3|Hoc est sacrificium ignis, quod offerre debetis: agnos anniculos immaculatos duos cotidie in holocaustum sempiternum;
NUM|28|4|unum offeretis mane et alterum ad vesperam;
NUM|28|5|decimam partem ephi similae in oblationem, quae conspersa sit oleo purissimo et habeat quartam partem hin.
NUM|28|6|Holocaustum iuge est, quod obtulistis in monte Sinai in odorem suavissimum, sacrificium ignis Domino;
NUM|28|7|et libabitis vini quartam partem hin per agnos singulos; in sanctuario effundetis libamen potus inebriantis Domino.
NUM|28|8|Alterumque agnum similiter offeretis ad vesperam, iuxta ritum sacrificii matutini: sacrificium ignis in odorem suavissimum Domino.
NUM|28|9|Die autem sabbati offeretis duos agnos anniculos immaculatos et duas decimas similae oleo conspersae et libamentum eius.
NUM|28|10|Est holocaustum sabbati per singula sabbata, praeter holocaustum sempiternum et libamentum eius.
NUM|28|11|In calendis autem offeretis holocaustum Domino vitulos de armento duos, arietem unum, agnos anniculos septem immaculatos
NUM|28|12|et tres decimas similae oleo conspersae in oblatione per singulos vitulos et duas decimas similae oleo conspersae per singulos arietes,
NUM|28|13|et decimam unam similae oleo conspersae in oblatione per agnos singulos: holocaustum in odorem suavissimum, sacrificium ignis Domino.
NUM|28|14|Libamenta autem eorum ista erunt: media pars hin vini per singulos vitulos, tertia per arietem, quarta per agnum. Hoc erit holocaustum per omnes menses, qui sibi anno vertente succedunt.
NUM|28|15|Hircus quoque offeretur Domino pro peccato, praeter holocaustum sempiternum cum libamentis suis.
NUM|28|16|Mense autem primo, quarta decima die mensis Pascha Domini erit,
NUM|28|17|et quinta decima die sollemnitas. Septem diebus vescemini azymis,
NUM|28|18|quarum die prima conventus sanctus erit; omne opus servile non facietis in ea.
NUM|28|19|Offeretisque sacrificium ignis, holocaustum Domino: vitulos de armento duos, arietem unum, agnos anniculos immaculatos septem;
NUM|28|20|et oblationem singulorum ex simila, quae conspersa sit oleo, tres decimas per singulos vitulos et duas decimas per arietem
NUM|28|21|et decimam unam per agnos singulos, id est per septem agnos;
NUM|28|22|et hircum pro peccato unum, ut expietur pro vobis,
NUM|28|23|praeter holocaustum matutinum, quod semper offeretis.
NUM|28|24|Ita facietis per singulos dies septem dierum: panem, sacrificium ignis in odorem suavissimum Domino praeter holocaustum iuge et libationem eius.
NUM|28|25|Die quoque septimo conventus sanctus erit vobis; omne opus servile non facietis in eo.
NUM|28|26|Die etiam primitivorum, quando offeretis oblationem novam Domino, in sollemnitate Hebdomadarum, conventus sanctus erit vobis; omne opus servile non facietis in ea.
NUM|28|27|Offeretisque holocaustum in odorem suavissimum Domino: vitulos de armento duos, arietem unum et agnos anniculos immaculatos septem,
NUM|28|28|atque in oblatione eorum similae oleo conspersae, tres decimas per singulos vitulos, per arietem duas,
NUM|28|29|per agnos decimam unam, qui simul sunt agni septem;
NUM|28|30|hircum quoque, qui mactatur pro expiatione,
NUM|28|31|praeter holocaustum sempiternum et oblationem eius. Immaculata offeretis omnia cum libationibus suis.
NUM|29|1|Mensis etiam septimi prima die conventus sanctus erit vo bis; omne opus servile non facietis in ea, quia dies clangoris est et tubarum.
NUM|29|2|Offeretisque holocaustum in odorem suavissimum Domino: vitulum de armento unum, arietem unum et agnos anniculos immaculatos septem;
NUM|29|3|et in oblationibus eorum similae oleo conspersae tres decimas per vitulum, duas decimas per arietem,
NUM|29|4|unam decimam per agnum, qui simul sunt agni septem;
NUM|29|5|et hircum pro peccato, qui offertur in expiationem vestram,
NUM|29|6|praeter holocaustum calendarum cum oblatione et holocaustum sempiternum cum oblatione et libationibus solitis in odorem suavissimum, sacrificium ignis Domino.
NUM|29|7|Decima quoque die mensis huius septimi erit vobis conventus sanctus, et affligetis animas vestras; omne opus servile non facietis.
NUM|29|8|Offeretisque holocaustum Domino in odorem suavissimum: vitulum de armento unum, arietem unum, agnos anniculos immaculatos septem;
NUM|29|9|et in oblatione eorum similae oleo conspersae tres decimas per vitulum, duas decimas per arietem,
NUM|29|10|decimam unam per agnos singulos, qui sunt simul septem agni;
NUM|29|11|et hircum pro peccato, absque his, quae offerri pro delicto solent in expiationem et holocaustum sempiternum cum oblatione et libaminibus eorum.
NUM|29|12|Quinta decima vero die mensis septimi conventus sanctus erit; omne opus servile non facietis in ea, sed celebrabitis sollemnitatem Domino septem diebus
NUM|29|13|offeretisque holocaustum in odorem suavissimum Domino: vitulos de armento tredecim, arietes duos, agnos anniculos immaculatos quattuordecim;
NUM|29|14|et in oblatione eorum similae oleo conspersae tres decimas per vitulos singulos, qui sunt simul vituli tredecim, et duas decimas arieti uno, id est simul arietibus duobus,
NUM|29|15|et decimam unam agnis singulis, qui sunt simul agni quattuordecim;
NUM|29|16|et hircum pro peccato absque holocausto sempiterno et oblatione et libamine eius.
NUM|29|17|In die altero offeretis vitulos de armento duodecim, arietes duos, agnos anniculos immaculatos quattuordecim;
NUM|29|18|oblationemque et libamina singulorum per vitulos et arietes et agnos iuxta numerum eorum rite celebrabitis,
NUM|29|19|et hircum pro peccato absque holocausto sempiterno oblationeque et libamine eorum.
NUM|29|20|Die tertio offeretis vitulos undecim, arietes duos, agnos anniculos imma culatos quattuordecim,
NUM|29|21|oblationem et libamina singulorum per vitulos et arietes et agnos iuxta numerum eorum rite celebrabitis,
NUM|29|22|et hircum pro peccato absque holocausto sempiterno oblationeque et libamine eius.
NUM|29|23|Die quarto offeretis vitulos decem, arietes duos, agnos anniculos immaculatos quattuordecim,
NUM|29|24|oblationem et libamina singulorum per vitulos et arietes et agnos iuxta numerum eorum rite celebrabitis,
NUM|29|25|et hircum pro peccato absque holocausto sempiterno, oblatione eius et libamine.
NUM|29|26|Die quinto offeretis vitulos novem, arietes duos, agnos anniculos immaculatos quattuordecim,
NUM|29|27|oblationem et libamina singulorum per vitulos et arietes et agnos iuxta numerum eorum rite celebrabitis,
NUM|29|28|et hircum pro peccato absque holocausto sempiterno, oblatione eius et libamine.
NUM|29|29|Die sexto offeretis vitulos octo, arietes duos, agnos anniculos immaculatos quattuordecim,
NUM|29|30|oblationem et libamina singulorum per vitulos et arietes et agnos iuxta numerum eorum rite celebrabitis,
NUM|29|31|et hircum pro peccato absque holocausto sempiterno, oblatione eius et libamine.
NUM|29|32|Die septimo offeretis vitulos septem et arietes duos, agnos anniculos immaculatos quattuordecim,
NUM|29|33|oblationem et libamina singulorum per vitulos et arietes et agnos iuxta numerum eorum rite celebrabitis,
NUM|29|34|et hircum pro peccato absque holocausto sempiterno, oblatione eius et libamine.
NUM|29|35|Die octavo erit conventus sollemnis, omne opus servile non facietis
NUM|29|36|offerentes holocaustum in odorem suavissimum Domino: vitulum unum, arietem unum, agnos anniculos immaculatos septem,
NUM|29|37|oblationem et libamina singulorum per vitulum et arietem et agnos iuxta numerum eorum rite celebrabitis,
NUM|29|38|et hircum pro peccato absque holocausto sempiterno, oblatione eius et libamine.
NUM|29|39|Haec offeretis Domino in sollemnitatibus vestris, praeter vota et oblationes spontaneas in holocaustis, in oblationibus, in libaminibus et in hostiis pacificis ".
NUM|30|1|Narravitque Moyses filiis Israel omnia, quae ei Dominus imperarat,
NUM|30|2|et locutus est ad principes tribuum filiorum Israel: " Iste est sermo, quem praecepit Dominus:
NUM|30|3|Si quis virorum votum Domino voverit aut se constrinxerit iuramento, non faciet irritum verbum suum, sed omne, quod promisit, implebit.
NUM|30|4|Mulier, si quippiam voverit Domino aut se constrinxerit iuramento, quae est in domo patris sui et in aetate adhuc puellari,
NUM|30|5|si cognoverit pater votum, quod pollicita est, aut iuramentum, quo ligavit animam suam, et tacuerit, voti rea erit; quidquid pollicita est aut iuravit, opere complebit.
NUM|30|6|Sin autem, quo die audierit contradixerit pater, et vota et iuramenta eius irrita erunt; et propitius erit ei Dominus, eo quod contradixerit pater.
NUM|30|7|Si maritum habuerit et voverit aliquid, aut semel de ore eius verbum egrediens animam eius ligaverit iuramento,
NUM|30|8|quo die audierit vir eius et non contradixerit, voti rea erit reddetque, quodcumque promiserat.
NUM|30|9|Sin autem, quo die audierit contradixerit, irritas facit pollicitationes eius verbaque, quibus obstrinxerat animam suam; et propitius erit ei Dominus.
NUM|30|10|Vidua et repudiata, quidquid voverint, reddent.
NUM|30|11|Uxor in domo viri cum se voto constrinxerit aut iuramento,
NUM|30|12|si audierit vir et tacuerit nec contradixerit sponsioni, reddet, quodcumque promiserat.
NUM|30|13|Sin autem extemplo contradixerit, non tenebitur promissionis rea, quia maritus contradixit, et Dominus ei propitius erit.
NUM|30|14|Si voverit aut iuramento se constrinxerit, ut per ieiunium affligat animam suam, in arbitrio viri erit, ut faciat sive non faciat.
NUM|30|15|Quod si audiens vir tacuerit et de die in diem distulerit sententiam, quidquid voverat atque promiserat, reddet, quia, quo die audierat, tacuit.
NUM|30|16|Sin autem contradixerit, postquam rescivit, portabit ipse iniquitatem eius ".
NUM|30|17|Istae sunt leges, quas constituit Dominus Moysi inter virum et uxorem, inter patrem et filiam, quae in puellari adhuc aetate manet in parentis domo.
NUM|31|1|Locutusque est Dominus ad Moysen dicens:
NUM|31|2|" Ulciscere filios Israel de Madianitis et sic colligeris ad populum tuum ".
NUM|31|3|Statimque Moyses: " Armate, inquit, ex vobis viros ad pugnam, qui possint ultionem Domini expetere de Madianitis.
NUM|31|4|Mille viri de singulis tribubus eligantur ex Israel, qui mittantur ad bellum ".
NUM|31|5|Dederuntque millenos de singulis tribubus, id est duodecim milia expeditorum ad pugnam,
NUM|31|6|quos misit Moyses cum Phinees filio Eleazari sacerdotis. Vasa quoque sancta et tubas ad clangendum tradidit ei.
NUM|31|7|Cumque pugnassent contra Madianitas, sicut praeceperat Dominus Moysi, omnes mares occiderunt
NUM|31|8|et reges eorum Evi et Recem et Sur et Hur et Rebe, quinque principes gentis, Balaam quoque filium Beor interfecerunt gladio;
NUM|31|9|ceperuntque mulieres eorum et parvulos. Omniaque pecora et cunctam supellectilem, quidquid habere potuerant, depopulati sunt:
NUM|31|10|tam urbes quam viculos et castra flamma consumpsit;
NUM|31|11|et tulerunt praedam et universa, quae ceperant, tam ex hominibus quam ex iumentis,
NUM|31|12|et adduxerunt captivos, spolia et praedam ad Moysen et Eleazarum sacerdotem et ad omnem congregationem filiorum Israel ad castra in campestribus Moab iuxta Iordanem contra Iericho.
NUM|31|13|Egressi sunt autem Moyses et Eleazar sacerdos et omnes principes synagogae in occursum eorum extra castra.
NUM|31|14|Iratusque Moyses principibus exercitus, tribunis et centurionibus, qui venerant de bello,
NUM|31|15|ait: " Cur omnes feminas reservastis?
NUM|31|16|Nonne istae sunt, quae deceperunt filios Israel ad suggestionem Balaam et praevaricari vos fecerunt in Dominum super peccato Phegor, unde et percussus est populus Domini?
NUM|31|17|Ergo cunctos interficite parvulos generis masculini et omnes mulieres, quae noverunt viros in coitu, iugulate;
NUM|31|18|puellas autem et omnes feminas virgines reservate vobis.
NUM|31|19|Et vos manete extra castra septem diebus; qui occiderit hominem vel occisum tetigerit, lustrabitur die tertio et septimo, vos et captivi vestri.
NUM|31|20|Et de omni praeda, sive vestimentum fuerit sive aliquid in utensilia praeparatum de caprarum pellibus et pilis et ligno, lustrabitis ".
NUM|31|21|Eleazar quoque sacerdos ad viros exercitus, qui pugnaverant, sic locutus est: " Hoc est praeceptum legis, quod mandavit Dominus Moysi:
NUM|31|22|Aurum et argentum et aes et ferrum et stannum et plumbum,
NUM|31|23|omne, quod potest transire per flammas, igne purgabitur; quidquid autem ignem non potest sustinere, aqua expiationis sanctificabitur.
NUM|31|24|Et lavabitis vestimenta vestra die septimo, et purificati postea castra intrabitis ".
NUM|31|25|Dixit quoque Dominus ad Moysen:
NUM|31|26|" Tollite summam eorum, quae capta sunt, ab homine usque ad pecus, tu et Eleazar sacerdos et principes familiarum;
NUM|31|27|dividesque ex aequo praedam inter eos, qui pugnaverunt egressique sunt ad bellum, et inter omnem congregationem.
NUM|31|28|Et separabis partem Domino ab his, qui pugnaverunt et fuerunt in bello, unam animam de quingentis tam ex hominibus quam ex bobus et asinis et ovibus
NUM|31|29|et dabis eam Eleazaro sacerdoti, quia praelibatio Domini sunt.
NUM|31|30|Ex media quoque parte filiorum Israel accipies quinquagesimum caput hominum et boum et asinorum et ovium cunctorum animantium et dabis ea Levitis, qui excubant in custodiis habitaculi Domini ".
NUM|31|31|Feceruntque Moyses et Eleazar sacerdos, sicut praeceperat Dominus.
NUM|31|32|Fuit autem praeda, quae supererat, quam exercitus ceperat, ovium sescenta septuaginta quinque milia,
NUM|31|33|boum septuaginta duo milia,
NUM|31|34|asinorum sexaginta milia et mille,
NUM|31|35|animae hominum sexus feminei, quae non cognoverant viros, triginta duo milia.
NUM|31|36|Dataque est media pars his, qui in proelio fuerant, ovium trecenta triginta septem milia quingentae,
NUM|31|37|e quibus in partem Domini supputatae sunt oves sescentae septuaginta quinque,
NUM|31|38|et de bobus triginta sex milibus, boves septuaginta et duo,
NUM|31|39|de asinis triginta milibus quingentis, asini sexaginta unus,
NUM|31|40|de animabus hominum sedecim milibus, cesserunt in partem Domini triginta duae animae.
NUM|31|41|Tradiditque Moyses tributum praelibationis Domini Eleazaro sacerdoti, sicut fuerat ei imperatum.
NUM|31|42|Ex media vero parte filiorum Israel, quam separaverat a parte eorum, qui in proelio fuerant,
NUM|31|43|de hac media parte, quae contigerat congregationi, id est de ovibus trecentis triginta septem milibus quingentis
NUM|31|44|et de bobus triginta sex milibus
NUM|31|45|et de asinis triginta milibus quingentis
NUM|31|46|et de hominibus sedecim milibus,
NUM|31|47|tulit Moyses quinquagesimum caput et dedit Levitis, qui excubabant in habitaculo Domini, sicut praeceperat Dominus.
NUM|31|48|Cumque accessissent principes exercitus ad Moysen, tribuni centurionesque, dixerunt:
NUM|31|49|" Nos servi tui recensuimus numerum pugnatorum, quos habuimus sub manu nostra, et ne unus quidem defuit.
NUM|31|50|Ob hanc causam offerimus in donariis Domini singuli, quod auri potuimus invenire, periscelidas et armillas, anulos et inaures ac muraenulas, ad placandum pro nobis Dominum ".
NUM|31|51|Susceperuntque Moyses et Eleazar sacerdos aurum in diversis speciebus;
NUM|31|52|omne aurum, quod elevaverunt Domino, pondo sedecim milia septingentos quinquaginta siclos, a tribunis et centurionibus.
NUM|31|53|Unusquisque enim, quod in praeda rapuerat, suum erat.
NUM|31|54|Et susceptum intulerunt in tabernaculum conventus in monumentum filiorum Israel coram Domino.
NUM|32|1|Filii autem Ruben et Gad habebant pecora multa, et erat illis in iumentis infinita substantia. Cumque vidissent Iazer et Galaad aptas animalibus alendis terras,
NUM|32|2|venerunt ad Moysen et ad Eleazarum sacerdotem et principes congregationis atque dixerunt:
NUM|32|3|" Ataroth et Dibon et Iazer et Nemra, Hesebon et Eleale et Sabam et Nabo et Beon,
NUM|32|4|terra, quam percussit Dominus in conspectu congregationis Israel, regio uberrima est ad pastum animalium, et nos servi tui habemus iumenta plurima ".
NUM|32|5|Dixeruntque: " Si invenimus gratiam coram te, detur haec terra famulis tuis in possessionem, nec facias nos transire Iordanem ".
NUM|32|6|Quibus respondit Moyses: " Numquid fratres vestri ibunt ad pugnam, et vos hic sedebitis?
NUM|32|7|Cur subvertitis mentes filiorum Israel, ne transire audeant in terram, quam eis daturus est Dominus?
NUM|32|8|Nonne ita egerunt patres vestri, quando misi de Cadesbarne ad explorandam terram?
NUM|32|9|Cumque venissent usque ad Nehelescol, lustrata omni regione, subverterunt cor filiorum Israel, ut non intrarent terram, quam eis Dominus dedit.
NUM|32|10|Qui iratus iuravit dicens:
NUM|32|11|"Non videbunt homines isti, qui ascenderunt ex Aegypto, a viginti annis et supra, terram, quam sub iuramento pollicitus sum Abraham, Isaac et Iacob; nam noluerunt sequi me,
NUM|32|12|praeter Chaleb filium Iephonne Cenezaeum et Iosue filium Nun: isti secuti sunt Dominum!".
NUM|32|13|Iratusque Dominus adversum Israel circumduxit eum per desertum quadraginta annis, donec consumeretur universa generatio, quae fecerat malum in conspectu eius.
NUM|32|14|Et ecce, inquit, vos surrexistis pro patribus vestris progenies hominum peccatorum, ut augeretis furorem irae Domini contra Israel.
NUM|32|15|Quod si nolueritis sequi eum, in solitudine iterum populum hunc circumducet, et vos causa eritis necis omnium ".
NUM|32|16|At illi prope accedentes dixerunt: " Caulas ovium fabricabimus pro iumentis nostris, parvulis quoque nostris urbes;
NUM|32|17|nos autem ipsi armati et accincti pergemus ad proelium ante filios Israel, donec introducamus eos ad loca sua. Parvuli nostri erunt in urbibus muratis propter habitatorum insidias.
NUM|32|18|Non revertemur in domos nostras usque dum possideant filii Israel hereditatem suam;
NUM|32|19|nec quidquam quaeremus trans Iordanem et ultra, quia iam habemus nostram hereditatem in orientali eius plaga ".
NUM|32|20|Quibus Moyses ait: " Si feceritis quod promittitis, si expediti perrexeritis coram Domino ad pugnam,
NUM|32|21|et omnis vir bellator armatus Iordanem transierit, donec expulerit Dominus inimicos suos ante se,
NUM|32|22|et subiecta ei omni terra redieritis in terram hanc, tunc eritis inculpabiles apud Dominum et apud Israel et obtinebitis terram hanc in hereditatem coram Domino.
NUM|32|23|Sin autem, quod dicitis, non feceritis, nulli dubium est quin peccetis in Dominum; et scitote quoniam peccatum vestrum apprehendet vos.
NUM|32|24|Aedificate ergo urbes parvulis vestris et caulas ovibus et, quod polliciti estis, implete ".
NUM|32|25|Dixeruntque filii Gad et Ruben ad Moysen: " Servi tui sumus, faciemus, quod iubet dominus noster:
NUM|32|26|parvulos nostros, mulieres, pecora ac iumenta remanebunt ibi in urbibus Galaad;
NUM|32|27|famuli autem tui, omnes expediti pergent coram Domino ad bellum, sicut tu, domine, loqueris ".
NUM|32|28|Praecepit ergo Moyses Eleazaro sacerdoti et Iosue filio Nun et principibus familiarum per tribus filiorum Israel et dixit ad eos:
NUM|32|29|" Si transierint filii Gad et filii Ruben vobiscum Iordanem omnes armati ad bellum coram Domino, et vobis fuerit terra subiecta, date eis Galaad in possessionem.
NUM|32|30|Sin autem noluerint transire armati vobiscum in terram Chanaan, inter vos habitandi accipiant loca ".
NUM|32|31|Responderuntque filii Gad et filii Ruben: " Sicut locutus est Dominus servis suis, ita faciemus.
NUM|32|32|Ipsi armati pergemus coram Domino in terram Chanaan; et possidebimus hereditatem nostram trans Iordanem ".
NUM|32|33|Dedit itaque Moyses filiis Gad et Ruben et dimidiae tribui Manasse filii Ioseph regnum Sehon regis Amorraei et regnum Og regis Basan, terram cum urbibus suis et terminis, urbes terrae per circuitum.
NUM|32|34|Igitur exstruxerunt filii Gad Dibon et Ataroth et Aroer
NUM|32|35|et Atrothsophan et Iazer et Iegbaa
NUM|32|36|et Bethnemra et Betharan, urbes munitas, et caulas pecoribus suis.
NUM|32|37|Filii vero Ruben aedificaverunt Hesebon et Eleale et Cariathaim
NUM|32|38|et Nabo et Baalmeon, versis nominibus, Sabama quoque, imponentes vocabula urbibus, quas exstruxerant.
NUM|32|39|Porro filii Machir filii Manasse perrexerunt in Galaad et ceperunt eam, expulso Amorraeo habitatore eius.
NUM|32|40|Dedit ergo Moyses terram Galaad Machir filio Manasse, qui habitavit in ea.
NUM|32|41|Iair autem filius Manasse abiit et occupavit vicos eius, quos appellavit Havoth Iair (id est villas Iair).
NUM|32|42|Nobe quoque perrexit et apprehendit Canath cum viculis suis vocavitque eam ex nomine suo Nobe.
NUM|33|1|Hae sunt mansiones filiorum Israel, qui egressi sunt de Ae gypto per turmas suas in manu Moysi et Aaron,
NUM|33|2|quas descripsit Moyses iuxta castrorum loca, quae Domini iussione mutabant.
NUM|33|3|Profecti igitur de Ramesse mense primo, quinta decima die mensis primi, altera die Paschae, filii Israel in manu excelsa, videntibus cunctis Aegyptiis
NUM|33|4|et sepelientibus primogenitos, quos percusserat Dominus, nam et in diis eorum exercuerat ultionem,
NUM|33|5|castrametati sunt in Succoth.
NUM|33|6|Et de Succoth venerunt in Etham, quae est in extremis finibus solitudinis.
NUM|33|7|Inde egressi venerunt contra Phihahiroth, quae respicit Beelsephon, et castrametati sunt ante Magdolum.
NUM|33|8|Profectique de Phihahiroth transierunt per medium mare in solitudinem, et ambulantes tribus diebus per desertum Etham castrametati sunt in Mara.
NUM|33|9|Profectique de Mara venerunt in Elim, ubi erant duodecim fontes aquarum et palmae septuaginta; ibique castrametati sunt.
NUM|33|10|Sed et inde egressi fixerunt tentoria super mare Rubrum. Profectique de mari Rubro
NUM|33|11|castrametati sunt in deserto Sin;
NUM|33|12|unde egressi venerunt in Daphca.
NUM|33|13|Profectique de Daphca castrametati sunt in Alus.
NUM|33|14|Egressique de Alus in Raphidim fixere tentoria, ubi populo defuit aqua ad bibendum;
NUM|33|15|profectique de Raphidim castrametati sunt in deserto Sinai.
NUM|33|16|Sed et de solitudine Sinai egressi venerunt ad Cibrottaava;
NUM|33|17|profectique de Cibrottaava castrametati sunt in Aseroth.
NUM|33|18|Et de Aseroth venerunt in Rethma;
NUM|33|19|profectique de Rethma castrametati sunt in Remmonphares.
NUM|33|20|Unde egressi venerunt in Lebna;
NUM|33|21|de Lebna castrametati sunt in Ressa;
NUM|33|22|egressique de Ressa venerunt in Ceelatha,
NUM|33|23|unde profecti castrametati sunt in monte Sepher.
NUM|33|24|Egressi de monte Sepher venerunt in Arada;
NUM|33|25|inde proficiscentes castrametati sunt in Maceloth;
NUM|33|26|profectique de Maceloth venerunt in Thahath;
NUM|33|27|de Thahath castrametati sunt in Thare.
NUM|33|28|Unde egressi fixere tentoria in Methca
NUM|33|29|et de Methca castrametati sunt in Hesmona;
NUM|33|30|profectique de Hesmona venerunt in Moseroth.
NUM|33|31|Et de Moseroth castrametati sunt in Beneiacan;
NUM|33|32|profectique de Beneiacan venerunt in montem Gadgad;
NUM|33|33|unde profecti castrametati sunt in Ietebatha.
NUM|33|34|Et de Ietebatha venerunt in Ebrona;
NUM|33|35|egressique de Ebrona castrametati sunt in Asiongaber.
NUM|33|36|Inde profecti venerunt in desertum Sin, hoc est Cades.
NUM|33|37|Egressique de Cades castrametati sunt in monte Hor in extremis finibus terrae Edom.
NUM|33|38|Ascenditque Aaron sacerdos in montem Hor, iubente Domino, et ibi mortuus est anno quadragesimo egressionis filiorum Israel ex Aegypto, mense quinto, prima die mensis,
NUM|33|39|cum esset annorum centum viginti trium.
NUM|33|40|Audivitque Chananaeus rex Arad, qui habitabat in Nageb, in terra Chanaan, venisse filios Israel.
NUM|33|41|Et profecti de monte Hor castrametati sunt in Salmona;
NUM|33|42|unde egressi venerunt in Phinon.
NUM|33|43|Profectique de Phinon castrametati sunt in Oboth;
NUM|33|44|et de Oboth venerunt in Ieabarim, quae est in finibus Moabitarum.
NUM|33|45|Profectique de Ieabarim fixere tentoria in Dibongad;
NUM|33|46|unde egressi castrametati sunt in Elmondeblathaim.
NUM|33|47|Egressique de Elmondeblathaim venerunt ad montes Abarim contra Nabo.
NUM|33|48|Profectique de montibus Abarim transierunt ad campestria Moab supra Iordanem contra Iericho;
NUM|33|49|ibique castrametati sunt de Bethiesimoth usque ad Abelsettim in campestribus Moab.
NUM|33|50|Ubi locutus est Dominus ad Moysen:
NUM|33|51|" Praecipe filiis Israel et dic ad eos: Quando transieritis Iordanem intrantes terram Chanaan,
NUM|33|52|disperdite cunctos habitatores terrae ante vos, confringite omnes imagines eorum et omnes statuas comminuite atque omnia excelsa vastate.
NUM|33|53|Possidebitis terram et habitabitis in ea. Ego enim dedi vobis illam in possessionem,
NUM|33|54|quam dividetis inter tribus vestras. Maiori dabitis latiorem et minori angustiorem; singulis, ut sors ceciderit, ita tribuetur hereditas; per tribus et familias possessio dividetur.
NUM|33|55|Sin autem nolueritis expellere habitatores terrae, qui remanserint, erunt vobis quasi spinae in oculis vestris et sudes in lateribus, et adversabuntur vobis in terra habitationis vestrae;
NUM|33|56|et, quidquid illis cogitaveram facere, vobis faciam ".
NUM|34|1|Locutusque est Dominus ad Moysen dicens:
NUM|34|2|" Praecipe fi liis Israel et dices ad eos: Cum ingressi fueritis terram hanc Chanaan, et in possessionem vobis sorte ceciderit, his finibus terminabitur.
NUM|34|3|Pars meridiana incipiet a solitudine Sin, quae est iuxta Edom, et habebit terminos contra orientem mare Salsissimum.
NUM|34|4|Qui circuibunt australem plagam per ascensum Acrabbim (id est Scorpionum), ita ut transeant in Sin et perveniant ad meridiem Cadesbarne, unde egredientur ad Asaraddar et tendent usque ad Asemona.
NUM|34|5|Ibitque per gyrum terminus ab Asemona usque ad torrentem Aegypti, et maris Magni litore finietur.
NUM|34|6|Plaga autem occidentalis a mari Magno incipiet et ipso fine claudetur.
NUM|34|7|Porro ad septentrionalem plagam a mari Magno termini incipient pervenientes usque ad montem Hor,
NUM|34|8|a quo venient in introitum Emath usque ad terminos Sedada.
NUM|34|9|Ibuntque confinia usque ad Zephrona et Asarenon. Hi erunt termini in parte aquilonis.
NUM|34|10|Inde metabuntur fines contra orientalem plagam de Asarenon usque Sephama;
NUM|34|11|et de Sephama descendent termini in Rebla ad orientem Ain; inde descendent et pervenient ad latus maris Chenereth in oriente
NUM|34|12|et tendent usque ad Iordanem, et ad ultimum Salsissimo claudentur mari.Hanc habebitis terram per fines suos in circuitu ".
NUM|34|13|Praecepitque Moyses filiis Israel dicens: " Haec erit terra, quam possidebitis sorte et quam iussit Dominus dari novem tribubus et dimidiae tribui.
NUM|34|14|Tribus enim filiorum Ruben per familias suas et tribus filiorum Gad iuxta cognationum numerum media quoque tribus Manasse,
NUM|34|15|id est duae semis tribus, acceperunt partem suam trans Iordanem contra Iericho ad orientalem plagam ".
NUM|34|16|Et ait Dominus ad Moysen:
NUM|34|17|" Haec sunt nomina virorum, qui terram vobis divident: Eleazar sacerdos et Iosue filius Nun
NUM|34|18|et singuli principes de tribubus singulis,
NUM|34|19|quorum ista sunt vocabula: de tribu Iudae Chaleb filius Iephonne;
NUM|34|20|de tribu Simeon Samuel filius Ammiud;
NUM|34|21|de tribu Beniamin Elidad filius Chaselon;
NUM|34|22|de tribu filiorum Dan Bocci filius Iogli.
NUM|34|23|Filiorum Ioseph: de tribu Manasse Hanniel filius Ephod,
NUM|34|24|de tribu Ephraim Camuel filius Sephtan.
NUM|34|25|De tribu Zabulon Elisaphan filius Pharnach;
NUM|34|26|de tribu Issachar dux Phaltiel filius Ozan;
NUM|34|27|de tribu Aser Ahiud filius Salomi;
NUM|34|28|de tribu Nephthali Phedael filius Ammiud ".
NUM|34|29|Hi sunt, quibus praecepit Dominus, ut dividerent filiis Israel terram Chanaan.
NUM|35|1|Haec quoque locutus est Do minus ad Moysen in campe stribus Moab supra Iordanem contra Iericho:
NUM|35|2|" Praecipe filiis Israel, ut dent Levitis de possessionibus suis urbes ad habitandum et suburbana earum per circuitum,
NUM|35|3|ut ipsi in oppidis maneant, et suburbana sint pecoribus ac substantiae et omnibus animalibus eorum;
NUM|35|4|quae a muris civitatum forinsecus per circuitum mille cubitos spatio tendentur.
NUM|35|5|Et mensurabitis extra civitatem contra orientem duo milia cubitorum, et contra meridiem similiter duo milia, ad mare quoque, quod respicit ad occidentem, eadem mensura erit, et septentrionalis plaga aequali termino finietur; eruntque urbes in medio et foris suburbana.
NUM|35|6|De ipsis autem oppidis, quae Levitis dabitis, sex erunt in fugitivorum auxilia separata, ut fugiat ad ea, qui nesciens fuderit sanguinem; et, exceptis his, alia quadraginta duo oppida dabitis,
NUM|35|7|id est simul quadraginta octo cum suburbanis suis.
NUM|35|8|Ipsaeque urbes, quas dabitis de possessionibus filiorum Israel, ab his, qui plus habent, plures auferetis, et, qui minus, pauciores; singuli iuxta mensuram hereditatis suae dabunt oppida Levitis ".
NUM|35|9|Ait Dominus ad Moysen:
NUM|35|10|" Loquere filiis Israel et dices ad eos: Quando transgressi fueritis Iordanem in terram Chanaan,
NUM|35|11|eligetis urbes, quae esse debeant in praesidia fugitivorum, qui nolentes sanguinem fuderint;
NUM|35|12|erunt vobis urbes refugii contra ultorem, et occisor non morietur, donec stet in conspectu congregationis, et causa illius iudicetur.
NUM|35|13|De ipsis autem sex urbibus, quae ad fugitivorum subsidia separantur,
NUM|35|14|tres erunt trans Iordanem et tres in terra Chanaan,
NUM|35|15|tam filiis Israel quam advenis atque peregrinis, ut confugiat ad eas sex, qui nolens sanguinem fuderit.
NUM|35|16|Si quis ferro percusserit, et mortuus fuerit, qui percussus est, reus erit homicidii et ipse morietur.
NUM|35|17|Si lapidem mortiferum iecerit, et ictus occiderit, similiter punietur.
NUM|35|18|Si ligno mortifero percusserit eum et interfecerit, homicida est; ipse morte punietur.
NUM|35|19|Ultor sanguinis homicidam interficiet: statim ut apprehenderit eum, interficiet.
NUM|35|20|Si per odium quis hominem impulerit vel iecerit quippiam in eum per insidias
NUM|35|21|aut, cum esset inimicus, manu percusserit, et ille mortuus fuerit, percussor homicidii reus erit: ultor sanguinis statim ut invenerit eum, iugulabit.
NUM|35|22|Quod si fortuitu et absque odio eum percusserit vel quidpiam in eum iecerit absque insidiis,
NUM|35|23|vel quemlibet lapidem mortiferum in eum devolverit, cum eum non vidisset, et ille mortuus est, quamvis eum non oderit nec quaesierit ei malum,
NUM|35|24|iudicabit congregatio inter percussorem et ultorem sanguinis secundum has regulas
NUM|35|25|et liberabit occisorem de manu ultoris sanguinis et reducet in civitatem refugii, ad quam confugerat, manebitque ibi, donec sacerdos magnus, qui oleo sancto unctus est, moriatur.
NUM|35|26|Si interfector extra fines civitatis refugii, in quam confugerat, exierit,
NUM|35|27|et invenerit eum ultor sanguinis ibi et interfecerit, absque noxa erit, qui eum occiderit;
NUM|35|28|debuerat enim profugus usque ad mortem pontificis in civitate refugii residere. Postquam autem ille obierit, homicida revertetur in terram suam.
NUM|35|29|Haec erunt vobis in legitima iudicii pro generationibus vestris, in cunctis habitationibus vestris.
NUM|35|30|Homicida sub testibus occidetur; ad unius testimonium nullus ad mortem condemnabitur.
NUM|35|31|Non accipietis pretium pro eo, qui reus est sanguinis, sed morietur.
NUM|35|32|Neque accipietis pretium, ut fugiat in civitatem refugii sui, ut revertatur et habitet in terra ante mortem sacerdotis.
NUM|35|33|Non polluetis terram habitationis vestrae, quia sanguis polluit terram, nec aliter expiari potest nisi per eius sanguinem, qui alterius sanguinem fuderit.
NUM|35|34|Non maculabitis terram habitationis vestrae, me commorante vobiscum. Ego enim sum Dominus, qui habito inter filios Israel ".
NUM|36|1|Accesserunt autem et princi pes familiarum tribus filio rum Galaad filii Machir filii Manasse de stirpe filiorum Ioseph; locutique sunt Moysi coram principibus familiarum Israel
NUM|36|2|atque dixerunt: " Tibi domino nostro praecepit Dominus, ut terram sorte divideres filiis Israel et ut filiabus Salphaad fratris nostri dares hereditatem debitam patri;
NUM|36|3|quas si alterius tribus homines uxores acceperint, sequetur possessio sua, et translata ad aliam tribum de nostra hereditate minuetur.
NUM|36|4|Atque ita fiet, ut cum iobeleus advenerit, addetur possessio earum possessioni tribus, ad quam pertinent, et a possessione tribus patrum nostrorum auferetur ".
NUM|36|5|Respondit Moyses filiis Israel et, Domino praecipiente, ait: " Recte tribus filiorum Ioseph locuta est,
NUM|36|6|et haec lex super filiabus Salphaad a Domino promulgata est: Nubant, quibus volunt, tantum ut suae tribus hominibus,
NUM|36|7|ne commisceatur possessio filiorum Israel de tribu in tribum; filii Israel adhaerebunt possessioni tribus patrum suorum,
NUM|36|8|et cunctae filiae heredes e filiis Israel maritos e cognatione tribus patrum suorum accipient, ut hereditas permaneat in familiis,
NUM|36|9|nec commisceatur possessio de tribu in tribum alteram, sed filii Israel adhaerebunt possessioni tribuum suarum ".
NUM|36|10|Sicut mandavit Dominus Moysi, sic fecerunt filiae Salphaad
NUM|36|11|et nupserunt Maala et Thersa et Hegla et Melcha et Noa filiis patruorum suorum
NUM|36|12|de familiis Manasse, qui fuit filius Ioseph; et possessio, quae illis fuerat attributa, mansit in tribu et familia patris earum.
NUM|36|13|Haec sunt mandata atque iudicia, quae mandavit Dominus per manum Moysi ad filios Israel in campestribus Moab supra Iordanem contra Iericho.
