2PET|1|1|Simon Petrus servus et apo stolus Iesu Christi his, qui coae qualem nobis sortiti sunt fidem in iustitia Dei nostri et salvatoris Iesu Christi:
2PET|1|2|gratia vobis et pax multiplicetur in cognitione Dei et Iesu Domini nostri.
2PET|1|3|Quomodo omnia nobis divinae virtutis suae ad vitam et pietatem donatae per cognitionem eius, qui vocavit nos propria gloria et virtute,
2PET|1|4|per quae pretiosa et maxima nobis promissa donata sunt, ut per haec efficiamini divinae consortes naturae, fugientes eam, quae in mundo est in concupiscentia, corruptionem;
2PET|1|5|et propter hoc ipsum curam omnem subinferentes ministrate in fide vestra virtutem, in virtute autem scientiam,
2PET|1|6|in scientia autem continentiam, in continentia autem patientiam, in patientia autem pietatem,
2PET|1|7|in pietate autem amorem fraternitatis, in amore autem fraternitatis caritatem.
2PET|1|8|Haec enim vobis, cum adsint et abundent, non vacuos nec sine fructu vos constituunt in Domini nostri Iesu Christi cognitionem;
2PET|1|9|cui enim non praesto sunt haec, caecus est et nihil procul cernens, oblivionem accipiens purgationis veterum suorum delictorum.
2PET|1|10|Quapropter, fratres, magis satagite, ut firmam vestram vocationem et electionem faciatis. Haec enim facientes non offendetis aliquando;
2PET|1|11|sic enim abundanter ministrabitur vobis introitus in aeternum regnum Domini nostri et salvatoris Iesu Christi.
2PET|1|12|Propter quod incipiam vos semper commonere de his, et quidem scientes et confirmatos in praesenti veritate.
2PET|1|13|Iustum autem arbitror, quamdiu sum in hoc tabernaculo, suscitare vos in commonitione,
2PET|1|14|certus quod velox est depositio tabernaculi mei, secundum quod et Dominus noster Iesus Christus significavit mihi;
2PET|1|15|dabo autem operam et frequenter habere vos post obitum meum, ut horum memoriam faciatis.
2PET|1|16|Non enim captiosas fabulas secuti notam fecimus vobis Domini nostri Iesu Christi virtutem et adventum, sed speculatores facti illius magnitudinis.
2PET|1|17|Accipiens enim a Deo Patre honorem et gloriam, voce prolata ad eum huiuscemodi a magnifica gloria: " Filius meus, dilectus meus hic est, in quo ego mihi complacui ";
2PET|1|18|et hanc vocem nos audivimus de caelo prolatam, cum essemus cum ipso in monte sancto.
2PET|1|19|Et habemus firmiorem propheticum sermonem, cui bene facitis attendentes quasi lucernae lucenti in caliginoso loco, donec dies illucescat, et lucifer oriatur in cordibus vestris,
2PET|1|20|hoc primum intellegentes quod omnis prophetia Scripturae propria interpretatione non fit;
2PET|1|21|non enim voluntate humana prolata est prophetia aliquando, sed a Spiritu Sancto ducti locuti sunt a Deo homines.
2PET|2|1|Fuerunt vero et pseudopro phetae in populo, sicut et in vo bis erunt magistri mendaces, qui introducent sectas perditionis et eum, qui emit eos, Dominatorem negantes superducent sibi celerem perditionem.
2PET|2|2|Et multi sequentur eorum luxurias, propter quos via veritatis blasphemabitur;
2PET|2|3|et in avaritia fictis verbis de vobis negotiabuntur. Quibus iudicium iam olim non cessat, et perditio eorum non dormitat.
2PET|2|4|Si enim Deus angelis peccantibus non pepercit, sed rudentibus inferni detractos in tartarum tradidit in iudicium reservatos:
2PET|2|5|et originali mundo non pepercit, sed octavum Noe iustitiae praeconem custodivit diluvium mundo impiorum inducens;
2PET|2|6|et civitates Sodomae et Gomorrae in cinerem redigens eversione damnavit, exemplum ponens eorum, quae sunt impiis futura:
2PET|2|7|et iustum Lot oppressum a nefandorum luxuria conversationis eruit:
2PET|2|8|aspectu enim et auditu iustus habitans apud eos, de die in diem animam iustam iniquis operibus cruciabat.
2PET|2|9|Novit Dominus pios de tentatione eripere, iniquos vero in diem iudicii puniendos reservare,
2PET|2|10|maxime autem eos, qui post carnem in concupiscentia immunditiae ambulant dominationemque contemnunt.Audaces, superbi, glorias non metuunt blasphemantes,
2PET|2|11|ubi angeli fortitudine et virtute cum sint maiores, non portant adversum illas coram Domino iudicium blasphemiae.
2PET|2|12|Hi vero, velut irrationabilia animalia naturaliter genita in captionem et in corruptionem, in his, quae ignorant, blasphemantes, in corruptione sua et corrumpentur
2PET|2|13|inviti percipientes mercedem iniustitiae; voluptatem existimantes diei delicias, coinquinationes et maculae deliciis affluentes, in voluptatibus suis luxuriantes vobiscum,
2PET|2|14|oculos habentes plenos adulterae et incessabiles delicti, pellicientes animas instabiles, cor exercitatum avaritiae habentes, maledictionis filii;
2PET|2|15|derelinquentes rectam viam erraverunt, secuti viam Balaam ex Bosor, qui mercedem iniquitatis amavit,
2PET|2|16|correptionem vero habuit suae praevaricationis; subiugale mutum in hominis voce loquens prohibuit prophetae insipientiam.
2PET|2|17|Hi sunt fontes sine aqua, et nebulae turbine exagitatae, quibus caligo tenebrarum reservatur.
2PET|2|18|Superba enim vanitatis loquentes pelliciunt in concupiscentiis carnis luxuriis illos, qui paululum effugiunt eos, qui in errore conversantur,
2PET|2|19|libertatem illis promittentes, cum ipsi servi sint corruptionis; a quo enim quis superatus est, huius servus est.
2PET|2|20|Si enim refugientes coinquinationes mundi in cognitione Domini nostri et Salvatoris Iesu Christi his rursus implicati superantur, facta sunt eis posteriora deteriora prioribus.
2PET|2|21|Melius enim erat illis non cognoscere viam iustitiae, quam post agnitionem retrorsum converti ab eo, quod illis traditum est, sancto mandato.
2PET|2|22|Contigit enim eis illud veri proverbii: Canis reversus ad suum vomitum ",et " Sus lota in volutabro luti ".
2PET|3|1|Hanc vobis, carissimi, iam se cundam scribo epistulam, in quibus excito vestram in commonitione sinceram mentem,
2PET|3|2|ut memores sitis eorum, quae praedicta sunt verborum a sanctis prophetis, et ab apostolis traditi vobis praecepti Domini et Salvatoris;
2PET|3|3|hoc primum scientes, quod venient in novissimis diebus in illusione illudentes, iuxta proprias concupiscentias suas ambulantes,
2PET|3|4|dicentes: " Ubi est promissio adventus eius? Ex quo enim patres dormierunt, omnia sic perseverant ab initio creaturae ".
2PET|3|5|Latet enim eos hoc volentes, quod caeli erant prius, et terra de aqua et per aquam consistens Dei verbo,
2PET|3|6|per quae ille tunc mundus aqua inundatus periit;
2PET|3|7|caeli autem, qui nunc sunt, et terra eodem verbo repositi sunt igni, servati in diem iudicii et perditionis impiorum hominum.
2PET|3|8|Unum vero hoc non lateat vos, carissimi, quia unus dies apud Dominum sicut mille anni, et mille anni sicut dies unus.
2PET|3|9|Non tardat Dominus promissionem, sicut quidam tarditatem existimant, sed patienter agit in vos nolens aliquos perire, sed omnes ad paenitentiam reverti.
2PET|3|10|Adveniet autem dies Domini ut fur, in qua caeli magno impetu transient, elementa vero calore solventur, et terra et opera, quae in ea invenientur.
2PET|3|11|Cum haec omnia ita dissolvenda sint, quales oportet esse vos in sanctis conversationibus et pietatibus,
2PET|3|12|exspectantes et properantes adventum diei Dei, propter quam caeli ardentes solventur, et elementa ignis ardore tabescent!
2PET|3|13|Novos vero caelos et terram novam secundum promissum ipsius exspectamus, in quibus iustitia habitat.
2PET|3|14|Propter quod, carissimi, haec exspectantes satagite immaculati et inviolati ei inveniri in pace;
2PET|3|15|et Domini nostri longanimitatem, salutem arbitramini, sicut et carissimus frater noster Paulus secundum datam sibi sapientiam scripsit vobis,
2PET|3|16|sicut et in omnibus epistulis loquens in eis de his; in quibus sunt quaedam difficilia intellectu, quae indocti et instabiles depravant, sicut et ceteras Scripturas, ad suam ipsorum perditionem.
2PET|3|17|Vos igitur, dilecti, praescientes custodite, ne iniquorum errore simul abducti excidatis a propria firmitate;
2PET|3|18|crescite vero in gratia et in cognitione Domini nostri et Salvatoris Iesu Christi. Ipsi gloria et nunc et in diem aeternitatis. Amen.
