JAS|1|1|Iacobus, Dei et Domini Iesu Christi servus, duodecim tribu bus, quae sunt in dispersione, salutem.
JAS|1|2|Omne gaudium existimate, fratres mei, cum in tentationibus variis incideritis,
JAS|1|3|scientes quod probatio fidei vestrae patientiam operatur;
JAS|1|4|patientia autem opus perfectum habeat, ut sitis perfecti et integri, in nullo deficientes.
JAS|1|5|Si quis autem vestrum indiget sapientia, postulet a Deo, qui dat omnibus affluenter et non improperat, et dabitur ei.
JAS|1|6|Postulet autem in fide nihil haesitans; qui enim haesitat, similis est fluctui maris, qui a vento movetur et circumfertur.
JAS|1|7|Non ergo aestimet homo ille quod accipiat aliquid a Domino,
JAS|1|8|vir duplex animo, inconstans in omnibus viis suis.
JAS|1|9|Glorietur autem frater humilis in exaltatione sua,
JAS|1|10|dives autem in humilitate sua, quoniam sicut flos feni transibit.
JAS|1|11|Exortus est enim sol cum ardore et arefecit fenum, et flos eius decidit, et decor vultus eius deperiit; ita et dives in itineribus suis marcescet.
JAS|1|12|Beatus vir, qui suffert tentationem, quia, cum probatus fuerit, accipiet coronam vitae, quam repromisit Deus diligentibus se.
JAS|1|13|Nemo, cum tentatur, dicat: " A Deo tentor "; Deus enim non tentatur malis, ipse autem neminem tentat.
JAS|1|14|Unusquisque vero tentatur a concupiscentia sua abstractus et illectus;
JAS|1|15|dein concupiscentia, cum conceperit, parit peccatum; peccatum vero, cum consummatum fuerit, generat mortem.
JAS|1|16|Nolite errare, fratres mei dilectissimi.
JAS|1|17|Omne datum optimum et omne donum perfectum de sursum est, descendens a Patre luminum, apud quem non est transmutatio nec vicissitudinis obumbratio.
JAS|1|18|Voluntarie genuit nos verbo veritatis, ut simus primitiae quaedam creaturae eius.
JAS|1|19|Scitis, fratres mei dilecti. Sit autem omnis homo velox ad audiendum, tardus autem ad loquendum et tardus ad iram;
JAS|1|20|ira enim viri iustitiam Dei non operatur.
JAS|1|21|Propter quod abicientes omnem immunditiam et abundantiam malitiae, in mansuetudine suscipite insitum verbum, quod potest salvare animas vestras.
JAS|1|22|Estote autem factores verbi et non auditores tantum fallentes vosmetipsos.
JAS|1|23|Quia si quis auditor est verbi et non factor, hic comparabitur viro consideranti vultum nativitatis suae in speculo;
JAS|1|24|consideravit enim se et abiit, et statim oblitus est qualis fuerit.
JAS|1|25|Qui autem perspexerit in lege perfecta libertatis et permanserit, non auditor obliviosus factus sed factor operis, hic beatus in facto suo erit.
JAS|1|26|Si quis putat se religiosum esse, non freno circumducens linguam suam sed seducens cor suum, huius vana est religio.
JAS|1|27|Religio munda et immaculata apud Deum et Patrem haec est: visitare pupillos et viduas in tribulatione eorum, immaculatum se custodire ab hoc saeculo.
JAS|2|1|Fratres mei, nolite in persona rum acceptione habere fidem Domini nostri Iesu Christi gloriae.
JAS|2|2|Etenim, si introierit in synagogam vestram vir aureum anulum habens in veste candida, introierit autem et pauper in sordido habitu,
JAS|2|3|et intendatis in eum, qui indutus est veste praeclara, et dixeritis: " Tu sede hic bene ", pauperi autem dicatis: " Tu sta illic aut sede sub scabello meo ";
JAS|2|4|nonne iudicatis apud vosmetipsos et facti estis iudices cogitationum iniquarum?
JAS|2|5|Audite, fratres mei dilectissimi. Nonne Deus elegit, qui pauperes sunt mundo, divites in fide et heredes regni, quod repromisit diligentibus se?
JAS|2|6|Vos autem exhonorastis pauperem. Nonne divites opprimunt vos et ipsi trahunt vos ad iudicia?
JAS|2|7|Nonne ipsi blasphemant bonum nomen, quod invocatum est super vos?
JAS|2|8|Si tamen legem perficitis regalem secundum Scripturam: " Diliges proximum tuum sicut teipsum ", bene facitis;
JAS|2|9|si autem personas accipitis, peccatum operamini, redarguti a lege quasi transgressores.
JAS|2|10|Quicumque autem totam legem servaverit, offendat autem in uno, factus est omnium reus.
JAS|2|11|Qui enim dixit: " Non moechaberis ", dixit et: " Non occides "; quod si non moecharis, occidis autem, factus es transgressor legis.
JAS|2|12|Sic loquimini et sic facite sicut per legem libertatis iudicandi.
JAS|2|13|Iudicium enim sine misericordia illi, qui non fecit misericordiam; superexsultat misericordia iudicio.
JAS|2|14|Quid proderit, fratres mei, si fidem quis dicat se habere, opera autem non habeat? Numquid poterit fides salvare eum?
JAS|2|15|Si frater aut soror nudi sunt et indigent victu cotidiano,
JAS|2|16|dicat autem aliquis de vobis illis: " Ite in pace, calefacimini et saturamini ", non dederitis autem eis, quae necessaria sunt corporis, quid proderit?
JAS|2|17|Sic et fides, si non habeat opera, mortua est in semetipsa.
JAS|2|18|Sed dicet quis: " Tu fidem habes, et ego opera habeo ". Ostende mihi fidem tuam sine operibus, et ego tibi ostendam ex operibus meis fidem.
JAS|2|19|Tu credis quoniam unus est Deus? Bene facis; et daemones credunt et contremiscunt!
JAS|2|20|Vis autem scire, o homo inanis, quoniam fides sine operibus otiosa est?
JAS|2|21|Abraham, pater noster, nonne ex operibus iustificatus est offerens Isaac filium suum super altare?
JAS|2|22|Vides quoniam fides cooperabatur operibus illius, et ex operibus fides consummata est;
JAS|2|23|et suppleta est Scriptura dicens: " Credidit Abraham Deo, et reputatum est illi ad iustitiam ", et amicus Dei appellatus est.
JAS|2|24|Videtis quoniam ex operibus iustificatur homo et non ex fide tantum.
JAS|2|25|Similiter autem et Rahab, meretrix nonne ex operibus iustificata est suscipiens nuntios et alia via eiciens?
JAS|2|26|Sicut enim corpus sine spiritu emortuum est, ita et fides sine operibus mortua est.
JAS|3|1|Nolite plures magistri fieri, fra tres mei, scientes quoniam maius iudicium accipiemus.
JAS|3|2|In multis enim offendimus omnes. Si quis in verbo non offendit, hic perfectus est vir, potens etiam freno circumducere totum corpus.
JAS|3|3|Si autem equorum frenos in ora mittimus ad oboediendum nobis, et omne corpus illorum circumferimus.
JAS|3|4|Ecce et naves, cum tam magnae sint et a ventis validis minentur, circumferuntur a minimo gubernaculo, ubi impetus dirigentis voluerit;
JAS|3|5|ita et lingua modicum quidem membrum est et magna exsultat. Ecce quantus ignis quam magnam silvam incendit!
JAS|3|6|Et lingua ignis est, universitas iniquitatis; lingua constituitur in membris nostris, quae maculat totum corpus et inflammat rotam nativitatis et inflammatur a gehenna.
JAS|3|7|Omnis enim natura et bestiarum et volucrum et serpentium et etiam cetorum domatur et domita est a natura humana;
JAS|3|8|linguam autem nullus hominum domare potest, inquietum malum, plena veneno mortifero.
JAS|3|9|In ipsa benedicimus Dominum et Patrem et in ipsa maledicimus homines, qui ad similitudinem Dei facti sunt;
JAS|3|10|ex ipso ore procedit benedictio et maledictio. Non oportet, fratres mei, haec ita fieri.
JAS|3|11|Numquid fons de eodem foramine emanat dulcem et amaram aquam?
JAS|3|12|Numquid potest, fratres mei, ficus olivas facere, aut vitis ficus? Neque salsa dulcem potest facere aquam.
JAS|3|13|Quis sapiens et disciplinatus inter vos? Ostendat ex bona conversatione operationem suam in mansuetudine sapientiae.
JAS|3|14|Quod si zelum amarum habetis et contentiones in cordibus vestris, nolite gloriari et mendaces esse adversus veritatem.
JAS|3|15|Non est ista sapientia desursum descendens, sed terrena, animalis, diabolica;
JAS|3|16|ubi enim zelus et contentio, ibi inconstantia et omne opus pravum.
JAS|3|17|Quae autem desursum est sapientia primum quidem pudica est, deinde pacifica, modesta, suadibilis, plena misericordia et fructibus bonis, non iudicans, sine simulatione;
JAS|3|18|fructus autem iustitiae in pace seminatur facientibus pacem.
JAS|4|1|Unde bella et unde lites in vobis? Nonne hinc, ex concupi scentiis vestris, quae militant in membris vestris?
JAS|4|2|Concupiscitis et non habetis; occiditis et zelatis et non potestis adipisci; litigatis et belligeratis. Non habetis, propter quod non postulatis;
JAS|4|3|petitis et non accipitis, eo quod male petitis, ut in concupiscentiis vestris insumatis.
JAS|4|4|Adulteri, nescitis quia amicitia huius mundi inimica est Dei?Quicumque ergo voluerit amicus esse saeculi huius, inimicus Dei constituitur.
JAS|4|5|Aut putatis quia inaniter Scriptura dicat: " Ad invidiam concupiscit Spiritus, qui inhabitat in nobis? ".
JAS|4|6|Maiorem autem dat gratiam; propter quod dicit: Deus superbis resistit,humilibus autem dat gratiam ".
JAS|4|7|Subicimini igitur Deo; resistite autem Diabolo, et fugiet a vobis.
JAS|4|8|Appropiate Deo, et appropinquabit vobis. Emundate manus, peccatores; et purificate corda, duplices animo.
JAS|4|9|Miseri estote et lugete et plorate; risus vester in luctum convertatur, et gaudium in maerorem.
JAS|4|10|Humiliamini in conspectu Domini, et exaltabit vos.
JAS|4|11|Nolite detrahere alterutrum, fratres; qui detrahit fratri, aut qui iudicat fratrem suum, detrahit legi et iudicat legem; si autem iudicas legem, non es factor legis sed iudex.
JAS|4|12|Unus est legislator et iudex, qui potest salvare et perdere; tu autem quis es, qui iudicas proximum?
JAS|4|13|Age nunc, qui dicitis: " Hodie aut crastino ibimus in illam civitatem et faciemus quidem ibi annum et mercabimur et lucrum faciemus ";
JAS|4|14|qui ignoratis, quae erit in crastinum vita vestra! Vapor enim estis ad modicum parens, deinceps exterminatur;
JAS|4|15|pro eo ut dicatis: " Si Dominus voluerit, et vivemus et faciemus hoc aut illud ".
JAS|4|16|Nunc autem gloriamini in superbiis vestris; omnis gloriatio talis maligna est.
JAS|4|17|Scienti igitur bonum facere et non facienti, peccatum est illi!
JAS|5|1|Age nunc, divites, plorate ulu lantes in miseriis, quae adve nient vobis.
JAS|5|2|Divitiae vestrae putrefactae sunt, et vestimenta vestra a tineis comesta sunt,
JAS|5|3|aurum et argentum vestrum aeruginavit, et aerugo eorum in testimonium vobis erit et manducabit carnes vestras sicut ignis: thesaurizastis in novissimis diebus.
JAS|5|4|Ecce merces operariorum, qui messuerunt regiones vestras, quae fraudata est a vobis, clamat, et clamores eorum, qui messuerunt, in aures Domini Sabaoth introierunt.
JAS|5|5|Epulati estis super terram et in luxuriis fuistis, enutristis corda vestra in die occisionis.
JAS|5|6|Addixistis, occidistis iustum. Non resistit vobis.
JAS|5|7|Patientes igitur estote, fratres, usque ad adventum Domini. Ecce agricola exspectat pretiosum fructum terrae, patienter ferens, donec accipiat imbrem temporaneum et serotinum.
JAS|5|8|Patientes estote, et vos, confirmate corda vestra, quoniam adventus Domini appropinquavit.
JAS|5|9|Nolite ingemiscere, fratres, in alterutrum, ut non iudicemini; ecce iudex ante ianuam assistit.
JAS|5|10|Exemplum accipite, fratres, laboris et patientiae prophetas, qui locuti sunt in nomine Domini.
JAS|5|11|Ecce beatificamus eos, qui sustinuerunt; sufferentiam Iob audistis et finem Domini vidistis, quoniam misericors est Dominus et miserator.
JAS|5|12|Ante omnia autem, fratres mei, nolite iurare neque per caelum neque per terram, neque aliud quodcumque iuramentum; sit autem vestrum " Est " est, et " Non " non, uti non sub iudicio decidatis.
JAS|5|13|Tristatur aliquis vestrum? Oret. Aequo animo est? Psallat.
JAS|5|14|Infirmatur quis in vobis? Advocet presbyteros ecclesiae, et orent super eum, unguentes eum oleo in nomine Domini.
JAS|5|15|Et oratio fidei salvabit infirmum, et allevabit eum Dominus; et si peccata operatus fuerit, dimittentur ei.
JAS|5|16|Confitemini ergo alterutrum peccata et orate pro invicem, ut sanemini. Multum enim valet deprecatio iusti operans.
JAS|5|17|Elias homo erat similis nobis passibilis et oratione oravit, ut non plueret, et non pluit super terram annos tres et menses sex;
JAS|5|18|et rursum oravit, et caelum dedit pluviam, et terra germinavit fructum suum.
JAS|5|19|Fratres mei, si quis ex vobis erraverit a veritate, et converterit quis eum,
JAS|5|20|scire debet quoniam, qui converti fecerit peccatorem ab errore viae eius, salvabit animam suam a morte et operiet multitudinem peccatorum.
