1TIM|1|1|Paul, an apostle of Christ Jesus by command of God our Savior and of Christ Jesus our hope,
1TIM|1|2|To Timothy, my true child in the faith: Grace, mercy, and peace from God the Father and Christ Jesus our Lord.
1TIM|1|3|As I urged you when I was going to Macedonia, remain at Ephesus that you may charge certain persons not to teach any different doctrine,
1TIM|1|4|nor to devote themselves to myths and endless genealogies, which promote speculations rather than the stewardship from God that is by faith.
1TIM|1|5|The aim of our charge is love that issues from a pure heart and a good conscience and a sincere faith.
1TIM|1|6|Certain persons, by swerving from these, have wandered away into vain discussion,
1TIM|1|7|desiring to be teachers of the law, without understanding either what they are saying or the things about which they make confident assertions.
1TIM|1|8|Now we know that the law is good, if one uses it lawfully,
1TIM|1|9|understanding this, that the law is not laid down for the just but for the lawless and disobedient, for the ungodly and sinners, for the unholy and profane, for those who strike their fathers and mothers, for murderers,
1TIM|1|10|the sexually immoral, men who practice homosexuality, enslavers, liars, perjurers, and whatever else is contrary to sound doctrine,
1TIM|1|11|in accordance with the glorious gospel of the blessed God with which I have been entrusted.
1TIM|1|12|I thank him who has given me strength, Christ Jesus our Lord, because he judged me faithful, appointing me to his service,
1TIM|1|13|though formerly I was a blasphemer, persecutor, and insolent opponent. But I received mercy because I had acted ignorantly in unbelief,
1TIM|1|14|and the grace of our Lord overflowed for me with the faith and love that are in Christ Jesus.
1TIM|1|15|The saying is trustworthy and deserving of full acceptance, that Christ Jesus came into the world to save sinners, of whom I am the foremost.
1TIM|1|16|But I received mercy for this reason, that in me, as the foremost, Jesus Christ might display his perfect patience as an example to those who were to believe in him for eternal life.
1TIM|1|17|To the King of ages, immortal, invisible, the only God, be honor and glory forever and ever. Amen.
1TIM|1|18|This charge I entrust to you, Timothy, my child, in accordance with the prophecies previously made about you, that by them you may wage the good warfare,
1TIM|1|19|holding faith and a good conscience. By rejecting this, some have made shipwreck of their faith,
1TIM|1|20|among whom are Hymenaeus and Alexander, whom I have handed over to Satan that they may learn not to blaspheme.
1TIM|2|1|First of all, then, I urge that supplications, prayers, intercessions, and thanksgivings be made for all people,
1TIM|2|2|for kings and all who are in high positions, that we may lead a peaceful and quiet life, godly and dignified in every way.
1TIM|2|3|This is good, and it is pleasing in the sight of God our Savior,
1TIM|2|4|who desires all people to be saved and to come to the knowledge of the truth.
1TIM|2|5|For there is one God, and there is one mediator between God and men, the man Christ Jesus,
1TIM|2|6|who gave himself as a ransom for all, which is the testimony given at the proper time.
1TIM|2|7|For this I was appointed a preacher and an apostle (I am telling the truth, I am not lying), a teacher of the Gentiles in faith and truth.
1TIM|2|8|I desire then that in every place the men should pray, lifting holy hands without anger or quarreling;
1TIM|2|9|likewise also that women should adorn themselves in respectable apparel, with modesty and self-control, not with braided hair and gold or pearls or costly attire,
1TIM|2|10|but with what is proper for women who profess godliness- with good works.
1TIM|2|11|Let a woman learn quietly with all submissiveness.
1TIM|2|12|I do not permit a woman to teach or to exercise authority over a man; rather, she is to remain quiet.
1TIM|2|13|For Adam was formed first, then Eve;
1TIM|2|14|and Adam was not deceived, but the woman was deceived and became a transgressor.
1TIM|2|15|Yet she will be saved through childbearing- if they continue in faith and love and holiness, with self-control.
1TIM|3|1|The saying is trustworthy: If anyone aspires to the office of overseer, he desires a noble task.
1TIM|3|2|Therefore an overseer must be above reproach, the husband of one wife, sober-minded, self-controlled, respectable, hospitable, able to teach,
1TIM|3|3|not a drunkard, not violent but gentle, not quarrelsome, not a lover of money.
1TIM|3|4|He must manage his own household well, with all dignity keeping his children submissive,
1TIM|3|5|for if someone does not know how to manage his own household, how will he care for God's church?
1TIM|3|6|He must not be a recent convert, or he may become puffed up with conceit and fall into the condemnation of the devil.
1TIM|3|7|Moreover, he must be well thought of by outsiders, so that he may not fall into disgrace, into a snare of the devil.
1TIM|3|8|Deacons likewise must be dignified, not double-tongued, not addicted to much wine, not greedy for dishonest gain.
1TIM|3|9|They must hold the mystery of the faith with a clear conscience.
1TIM|3|10|And let them also be tested first; then let them serve as deacons if they prove themselves blameless.
1TIM|3|11|Their wives likewise must be dignified, not slanderers, but sober-minded, faithful in all things.
1TIM|3|12|Let deacons each be the husband of one wife, managing their children and their own households well.
1TIM|3|13|For those who serve well as deacons gain a good standing for themselves and also great confidence in the faith that is in Christ Jesus.
1TIM|3|14|I hope to come to you soon, but I am writing these things to you so that,
1TIM|3|15|if I delay, you may know how one ought to behave in the household of God, which is the church of the living God, a pillar and buttress of truth.
1TIM|3|16|Great indeed, we confess, is the mystery of godliness: He was manifested in the flesh, vindicated by the Spirit, seen by angels, proclaimed among the nations, believed on in the world, taken up in glory.
1TIM|4|1|Now the Spirit expressly says that in later times some will depart from the faith by devoting themselves to deceitful spirits and teachings of demons,
1TIM|4|2|through the insincerity of liars whose consciences are seared,
1TIM|4|3|who forbid marriage and require abstinence from foods that God created to be received with thanksgiving by those who believe and know the truth.
1TIM|4|4|For everything created by God is good, and nothing is to be rejected if it is received with thanksgiving,
1TIM|4|5|for it is made holy by the word of God and prayer.
1TIM|4|6|If you put these things before the brothers, you will be a good servant of Christ Jesus, being trained in the words of the faith and of the good doctrine that you have followed.
1TIM|4|7|Have nothing to do with irreverent, silly myths. Rather train yourself for godliness;
1TIM|4|8|for while bodily training is of some value, godliness is of value in every way, as it holds promise for the present life and also for the life to come.
1TIM|4|9|The saying is trustworthy and deserving of full acceptance.
1TIM|4|10|For to this end we toil and strive, because we have our hope set on the living God, who is the Savior of all people, especially of those who believe.
1TIM|4|11|Command and teach these things.
1TIM|4|12|Let no one despise you for your youth, but set the believers an example in speech, in conduct, in love, in faith, in purity.
1TIM|4|13|Until I come, devote yourself to the public reading of Scripture, to exhortation, to teaching.
1TIM|4|14|Do not neglect the gift you have, which was given you by prophecy when the council of elders laid their hands on you.
1TIM|4|15|Practice these things, devote yourself to them, so that all may see your progress.
1TIM|4|16|Keep a close watch on yourself and on the teaching. Persist in this, for by so doing you will save both yourself and your hearers.
1TIM|5|1|Do not rebuke an older man but encourage him as you would a father. Treat younger men like brothers,
1TIM|5|2|older women like mothers, younger women like sisters, in all purity.
1TIM|5|3|Honor widows who are truly widows.
1TIM|5|4|But if a widow has children or grandchildren, let them first learn to show godliness to their own household and to make some return to their parents, for this is pleasing in the sight of God.
1TIM|5|5|She who is truly a widow, left all alone, has set her hope on God and continues in supplications and prayers night and day,
1TIM|5|6|but she who is self-indulgent is dead even while she lives.
1TIM|5|7|Command these things as well, so that they may be without reproach.
1TIM|5|8|But if anyone does not provide for his relatives, and especially for members of his household, he has denied the faith and is worse than an unbeliever.
1TIM|5|9|Let a widow be enrolled if she is not less than sixty years of age, having been the wife of one husband,
1TIM|5|10|and having a reputation for good works: if she has brought up children, has shown hospitality, has washed the feet of the saints, has cared for the afflicted, and has devoted herself to every good work.
1TIM|5|11|But refuse to enroll younger widows, for when their passions draw them away from Christ, they desire to marry
1TIM|5|12|and so incur condemnation for having abandoned their former faith.
1TIM|5|13|Besides that, they learn to be idlers, going about from house to house, and not only idlers, but also gossips and busybodies, saying what they should not.
1TIM|5|14|So I would have younger widows marry, bear children, manage their households, and give the adversary no occasion for slander.
1TIM|5|15|For some have already strayed after Satan.
1TIM|5|16|If any believing woman has relatives who are widows, let her care for them. Let the church not be burdened, so that it may care for those who are really widows.
1TIM|5|17|Let the elders who rule well be considered worthy of double honor, especially those who labor in preaching and teaching.
1TIM|5|18|For the Scripture says, "You shall not muzzle an ox when it treads out the grain," and, "The laborer deserves his wages."
1TIM|5|19|Do not admit a charge against an elder except on the evidence of two or three witnesses.
1TIM|5|20|As for those who persist in sin, rebuke them in the presence of all, so that the rest may stand in fear.
1TIM|5|21|In the presence of God and of Christ Jesus and of the elect angels I charge you to keep these rules without prejudging, doing nothing from partiality.
1TIM|5|22|Do not be hasty in the laying on of hands, nor take part in the sins of others; keep yourself pure.
1TIM|5|23|(No longer drink only water, but use a little wine for the sake of your stomach and your frequent ailments.)
1TIM|5|24|The sins of some men are conspicuous, going before them to judgment, but the sins of others appear later.
1TIM|5|25|So also good works are conspicuous, and even those that are not cannot remain hidden.
1TIM|6|1|Let all who are under a yoke as slaves regard their own masters as worthy of all honor, so that the name of God and the teaching may not be reviled.
1TIM|6|2|Those who have believing masters must not be disrespectful on the ground that they are brothers; rather they must serve all the better since those who benefit by their good service are believers and beloved. Teach and urge these things.
1TIM|6|3|If anyone teaches a different doctrine and does not agree with the sound words of our Lord Jesus Christ and the teaching that accords with godliness,
1TIM|6|4|he is puffed up with conceit and understands nothing. He has an unhealthy craving for controversy and for quarrels about words, which produce envy, dissension, slander, evil suspicions,
1TIM|6|5|and constant friction among people who are depraved in mind and deprived of the truth, imagining that godliness is a means of gain.
1TIM|6|6|Now there is great gain in godliness with contentment,
1TIM|6|7|for we brought nothing into the world, and we cannot take anything out of the world.
1TIM|6|8|But if we have food and clothing, with these we will be content.
1TIM|6|9|But those who desire to be rich fall into temptation, into a snare, into many senseless and harmful desires that plunge people into ruin and destruction.
1TIM|6|10|For the love of money is a root of all kinds of evils. It is through this craving that some have wandered away from the faith and pierced themselves with many pangs.
1TIM|6|11|But as for you, O man of God, flee these things. Pursue righteousness, godliness, faith, love, steadfastness, gentleness.
1TIM|6|12|Fight the good fight of the faith. Take hold of the eternal life to which you were called and about which you made the good confession in the presence of many witnesses.
1TIM|6|13|I charge you in the presence of God, who gives life to all things, and of Christ Jesus, who in his testimony before Pontius Pilate made the good confession,
1TIM|6|14|to keep the commandment unstained and free from reproach until the appearing of our Lord Jesus Christ,
1TIM|6|15|which he will display at the proper time- he who is the blessed and only Sovereign, the King of kings and Lord of lords,
1TIM|6|16|who alone has immortality, who dwells in unapproachable light, whom no one has ever seen or can see. To him be honor and eternal dominion. Amen.
1TIM|6|17|As for the rich in this present age, charge them not to be haughty, nor to set their hopes on the uncertainty of riches, but on God, who richly provides us with everything to enjoy.
1TIM|6|18|They are to do good, to be rich in good works, to be generous and ready to share,
1TIM|6|19|thus storing up treasure for themselves as a good foundation for the future, so that they may take hold of that which is truly life.
1TIM|6|20|O Timothy, guard the deposit entrusted to you. Avoid the irreverent babble and contradictions of what is falsely called "knowledge,"
1TIM|6|21|for by professing it some have swerved from the faith. Grace be with you.
