PHLM|1|1|為基督耶穌被囚的 保羅 ，同弟兄 提摩太 ，寫信給我們所親愛的同工 腓利門 、
PHLM|1|2|亞腓亞 姊妹，和我們的戰友 亞基布 ，以及在你家裏的教會。
PHLM|1|3|願恩惠、平安 從我們的父上帝和主耶穌基督歸給你們！
PHLM|1|4|我在禱告中記念你的時候，常為你感謝我的上帝，
PHLM|1|5|因聽說你對眾聖徒的愛心，和你對主耶穌的信心。
PHLM|1|6|願你與人分享信心的時候，能產生功效，讓人知道我們 所行的各樣善事都是為基督做的。
PHLM|1|7|弟兄啊，由於你的愛心，我得到極大的快樂和安慰，因為眾聖徒的心從你得到舒暢。
PHLM|1|8|雖然我靠著基督能放膽吩咐你做該做的事，
PHLM|1|9|可是像我這上了年紀的 保羅 ，現在又是為基督耶穌被囚的，寧可憑著愛心求你，
PHLM|1|10|就是為我在捆鎖中所生的兒子 阿尼西謀 求你。
PHLM|1|11|從前他與你沒有益處，但如今與你我都有益處。
PHLM|1|12|我現在打發他回到你那裏去，他是我心肝。
PHLM|1|13|我本來有意將他留下，在我為福音所受的捆鎖中替你伺候我。
PHLM|1|14|但不知道你的意見，我不願意這樣做，好使你的善行不是出於勉強，而是出於自願。
PHLM|1|15|他暫時離開你，也許是要讓你永遠得著他，
PHLM|1|16|不再是奴隸，而是高過奴隸，是親愛的弟兄；對我確實如此，何況對你呢！無論在肉身或在主裏更是如此。
PHLM|1|17|所以，你若以我為同伴，就接納他，如同接納我一樣。
PHLM|1|18|他若虧負你，或欠你甚麼，都算在我的賬上吧，
PHLM|1|19|我必償還。這是我— 保羅 親筆寫的。我並不用對你說，甚至你自己也虧欠我呢！
PHLM|1|20|弟兄啊，希望你使我在主裏因你得益處，讓我的心在基督裏得到舒暢。
PHLM|1|21|我寫信給你，深信你必順服，知道你所要做的，必過於我所說的。
PHLM|1|22|此外，還請給我預備住處，因為我盼望藉著你們的禱告，必蒙恩回到你們那裏去。
PHLM|1|23|為基督耶穌與我一同坐監的 以巴弗 問候你。
PHLM|1|24|我的同工 馬可 、 亞里達古 、 底馬 、 路加 也都問候你。
PHLM|1|25|願 主耶穌基督的恩與你們的靈同在。
