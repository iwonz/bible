HAB|1|1|哈巴谷 先知所看見的默示。
HAB|1|2|耶和華啊，我呼求， 你不應允，要到幾時呢？ 我向你呼喊「暴力！」 你還不拯救？
HAB|1|3|你為何使我看見罪孽？ 你為何坐視奸惡呢？ 毀滅和兇暴在我面前， 爭執與紛爭不斷發生。
HAB|1|4|因此律法無效， 公理從未彰顯。 因惡人圍困義人， 所以公理遭受扭曲。
HAB|1|5|你們要向列國觀看 ，注意看， 要驚奇，再驚奇！ 因為在你們的日子，有一件事發生 ， 儘管有人說了，你們還是不信。
HAB|1|6|看哪，我必興起 迦勒底 人， 就是那殘忍暴躁之民，通行遍地， 霸佔不屬自己的住處。
HAB|1|7|他威武可畏， 審判與威權都由他而出。
HAB|1|8|他的馬比豹更快， 比晚上 的野狼更猛。 他的戰馬跳躍， 他的戰馬從遠方而來 ； 他們飛跑，如鷹急速抓食，
HAB|1|9|都為施行殘暴而來， 他們的臉面向東 ， 聚集俘虜，多如塵沙。
HAB|1|10|他譏誚列王， 嘲諷領袖， 嗤笑一切堡壘， 堆土攻取它。
HAB|1|11|那時，他如風猛然掃過， 他背叛，顯為有罪； 他以自己的力量為神明。
HAB|1|12|耶和華－我的上帝，我的聖者啊， 你不是從亙古就有嗎？ 我們必不致死。 耶和華啊，你派他為要行審判； 磐石啊，你立他為要懲治人。
HAB|1|13|你的眼目清潔， 不看邪惡，也不看奸惡， 為何你卻看著人行詭詐呢？ 惡人吞滅比自己公義的人， 為何你保持沉默呢？
HAB|1|14|你為何使人如海中的魚， 又如無人管轄的爬行動物呢？
HAB|1|15|他用鉤子把他們全拉上來， 用羅網捕獲他們， 拉漁網聚集他們。 因此，他歡喜快樂，
HAB|1|16|向羅網獻祭， 向漁網燒香； 因為他藉此得豐盛的收穫 與肥美的食物。
HAB|1|17|但他豈可因此屢屢倒空羅網 ， 時常殺戮列國的人，毫不顧惜呢？
HAB|2|1|我要站在我的瞭望臺， 立在城樓 上觀看， 看耶和華要對我說甚麼， 我可用甚麼話向他訴冤。
HAB|2|2|耶和華回答我，說： 將這默示清楚地寫在看板上， 使人容易朗讀 。
HAB|2|3|因為這默示有一定日期， 論及終局，絕不落空。 它雖然耽延，你要等候； 因為它必臨到，不再遲延。
HAB|2|4|看哪，惡人自高自大，心不正直； 惟義人必因他的信得生 。
HAB|2|5|他因酒詭詐、 狂傲、不安於位； 他張開喉嚨 ，好像陰間， 如死亡不能知足， 他聚集萬國， 招聚萬民全歸自己。
HAB|2|6|這些人豈不都要提起詩歌和俗語，嘲諷他說： 禍哉！你增添不屬自己的財物， 靠押金發財，要到幾時呢？
HAB|2|7|咬傷你的 豈不忽然興起， 擾害你的豈不突然崛起， 你就成為他們的擄物嗎？
HAB|2|8|因你搶奪許多國家， 流人的血，向土地、城鎮和全城的居民施行殘暴， 各國殘存之民都必搶奪你。
HAB|2|9|禍哉！那為本家積蓄不義之財、 在高處搭窩、指望得免災禍的人！
HAB|2|10|你圖謀剪除許多民族，犯了罪， 使自己的家蒙羞，自害己命。
HAB|2|11|牆裏的石頭要呼叫， 屋內的棟梁必應聲。
HAB|2|12|禍哉！那以鮮血建城、 以罪孽造鎮的人！
HAB|2|13|看哪，這不都是 出於萬軍之耶和華嗎？ 萬民勞碌得來的被火焚燒， 萬族辛苦建造的，歸於虛空。
HAB|2|14|全地都必認識耶和華的榮耀， 好像水充滿海洋一般。
HAB|2|15|禍哉！那給鄰舍酒喝，加上毒物 ， 使人喝醉，為要看見他們下體的人！
HAB|2|16|你滿受羞辱，不得榮耀； 你也喝吧，顯明你是未受割禮的 ！ 耶和華右手的杯必傳到你那裏， 你的榮耀就變為羞辱。
HAB|2|17|黎巴嫩 所受的殘暴必淹沒你， 野獸所遭遇的毀滅使你驚嚇 ； 因你流人的血， 向土地、城鎮和全城的居民施行殘暴。
HAB|2|18|偶像有甚麼益處呢？ 製造者雕刻它， 鑄成偶像，作虛假的教師； 製造者倚靠的是自己所做的啞巴偶像。
HAB|2|19|禍哉！那對木頭說「醒起」， 對啞巴石頭說「起來」的人！ 偶像豈能教導人呢？ 看哪，它以金銀包裹，其中並無氣息。
HAB|2|20|惟耶和華在他的聖殿中， 全地都當在他面前肅靜。
HAB|3|1|哈巴谷 先知的禱告，調用流離歌。
HAB|3|2|耶和華啊，我聽見你的名聲； 耶和華啊，我懼怕你的作為。 求你在這些年間 復興你的作為， 在這些年間將它顯明出來 ； 在發怒的時候以憐憫為念。
HAB|3|3|上帝從 提幔 而來， 聖者從 巴蘭山 臨到； 他的榮光遮蔽諸天， 頌讚遍滿全地。
HAB|3|4|他的輝煌如同日光， 從他手裏發出光芒， 那裏 隱藏他的能力。
HAB|3|5|在他前面有瘟疫流行， 在他腳下有熱症發出。
HAB|3|6|他站立，震動 大地， 他觀看，震動列國。 永久的山崩裂， 長存的嶺塌陷， 他的作為與古時一樣。
HAB|3|7|我見 古珊 的帳棚遭難， 米甸 地的幔子動搖。
HAB|3|8|耶和華啊，你豈是向江河發怒， 向江河生氣， 向海洋發烈怒嗎？ 你騎在馬上， 坐在得勝的戰車上，
HAB|3|9|你的弓全然顯露 ， 箭是發誓的言語 ； 你以江河分開大地。
HAB|3|10|山嶺見你，無不戰抖； 大水氾濫而過， 深淵發聲， 洶湧翻騰 。
HAB|3|11|因你的箭射出光芒， 你的槍閃出光耀， 日月都停在原處。
HAB|3|12|你發怒遍行大地， 以怒氣責打列國，如打穀一般。
HAB|3|13|你出來拯救你的百姓， 拯救你的受膏者； 你打破惡人之家的頭， 暴露其根基，直到頸項 。
HAB|3|14|你以其戈矛刺透他戰士的頭； 他們如旋風將我 颳散， 他們喜愛暗中吞吃困苦的人。
HAB|3|15|你騎馬踐踏海， 踐踏洶湧的大水。
HAB|3|16|我聽見這聲音，身體戰兢， 嘴唇發顫， 骨中朽爛， 在所立之處戰兢 ； 但我安靜等候 災難之日臨到那上來侵犯我們的民 。
HAB|3|17|雖然無花果樹不發旺， 葡萄樹不結果， 橄欖樹也不收成， 田地不出糧食， 圈中絕了羊， 棚內也沒有牛；
HAB|3|18|然而，我要因耶和華歡欣， 因救我的上帝喜樂。
HAB|3|19|主耶和華是我的力量， 他使我的腳快如母鹿， 又使我穩行在高處。 這歌交給聖詠團長，用絲弦的樂器。
