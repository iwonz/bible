ESTH|1|1|Now in the days of Ahasuerus, the Ahasuerus who reigned from India to Ethiopia over 127 provinces,
ESTH|1|2|in those days when King Ahasuerus sat on his royal throne in Susa, the capital,
ESTH|1|3|in the third year of his reign he gave a feast for all his officials and servants. The army of Persia and Media and the nobles and governors of the provinces were before him,
ESTH|1|4|while he showed the riches of his royal glory and the splendor and pomp of his greatness for many days, 180 days.
ESTH|1|5|And when these days were completed, the king gave for all the people present in Susa, the citadel, both great and small, a feast lasting for seven days in the court of the garden of the king's palace.
ESTH|1|6|There were white cotton curtains and violet hangings fastened with cords of fine linen and purple to silver rods and marble pillars, and also couches of gold and silver on a mosaic pavement of porphyry, marble, mother-of-pearl and precious stones.
ESTH|1|7|Drinks were served in golden vessels, vessels of different kinds, and the royal wine was lavished according to the bounty of the king.
ESTH|1|8|And drinking was according to this edict: "There is no compulsion." For the king had given orders to all the staff of his palace to do as each man desired.
ESTH|1|9|Queen Vashti also gave a feast for the women in the palace that belonged to King Ahasuerus.
ESTH|1|10|On the seventh day, when the heart of the king was merry with wine, he commanded Mehuman, Biztha, Harbona, Bigtha and Abagtha, Zethar and Carkas, the seven eunuchs who served in the presence of King Ahasuerus,
ESTH|1|11|to bring Queen Vashti before the king with her royal crown, in order to show the peoples and the princes her beauty, for she was lovely to look at.
ESTH|1|12|But Queen Vashti refused to come at the king's command delivered by the eunuchs. At this the king became enraged, and his anger burned within him.
ESTH|1|13|Then the king said to the wise men who knew the times (for this was the king's procedure toward all who were versed in law and judgment,
ESTH|1|14|the men next to him being Carshena, Shethar, Admatha, Tarshish, Meres, Marsena, and Memucan, the seven princes of Persia and Media, who saw the king's face, and sat first in the kingdom):
ESTH|1|15|"According to the law, what is to be done to Queen Vashti, because she has not performed the command of King Ahasuerus delivered by the eunuchs?"
ESTH|1|16|Then Memucan said in the presence of the king and the officials, "Not only against the king has Queen Vashti done wrong, but also against all the officials and all the peoples who are in all the provinces of King Ahasuerus.
ESTH|1|17|For the queen's behavior will be made known to all women, causing them to look at their husbands with contempt, since they will say, 'King Ahasuerus commanded Queen Vashti to be brought before him, and she did not come.'
ESTH|1|18|This very day the noble women of Persia and Media who have heard of the queen's behavior will say the same to all the king's officials, and there will be contempt and wrath in plenty.
ESTH|1|19|If it please the king, let a royal order go out from him, and let it be written among the laws of the Persians and the Medes so that it may not be repealed, that Vashti is never again to come before King Ahasuerus. And let the king give her royal position to another who is better than she.
ESTH|1|20|So when the decree made by the king is proclaimed throughout all his kingdom, for it is vast, all women will give honor to their husbands, high and low alike."
ESTH|1|21|This advice pleased the king and the princes, and the king did as Memucan proposed.
ESTH|1|22|He sent letters to all the royal provinces, to every province in its own script and to every people in its own language, that every man be master in his own household and speak according to the language of his people.
ESTH|2|1|After these things, when the anger of King Ahasuerus had abated, he remembered Vashti and what she had done and what had been decreed against her.
ESTH|2|2|Then the king's young men who attended him said, "Let beautiful young virgins be sought out for the king.
ESTH|2|3|And let the king appoint officers in all the provinces of his kingdom to gather all the beautiful young virgins to the harem in Susa the capital, under custody of Hegai, the king's eunuch, who is in charge of the women. Let their cosmetics be given them.
ESTH|2|4|And let the young woman who pleases the king be queen instead of Vashti." This pleased the king, and he did so.
ESTH|2|5|Now there was a Jew in Susa the citadel whose name was Mordecai, the son of Jair, son of Shimei, son of Kish, a Benjaminite,
ESTH|2|6|who had been carried away from Jerusalem among the captives carried away with Jeconiah king of Judah, whom Nebuchadnezzar king of Babylon had carried away.
ESTH|2|7|He was bringing up Hadassah, that is Esther, the daughter of his uncle, for she had neither father nor mother. The young woman had a beautiful figure and was lovely to look at, and when her father and her mother died, Mordecai took her as his own daughter.
ESTH|2|8|So when the king's order and his edict were proclaimed, and when many young women were gathered in Susa the citadel in custody of Hegai, Esther also was taken into the king's palace and put in custody of Hegai, who had charge of the women.
ESTH|2|9|And the young woman pleased him and won his favor. And he quickly provided her with her cosmetics and her portion of food, and with seven chosen young women from the king's palace, and advanced her and her young women to the best place in the harem.
ESTH|2|10|Esther had not made known her people or kindred, for Mordecai had commanded her not to make it known.
ESTH|2|11|And every day Mordecai walked in front of the court of the harem to learn how Esther was and what was happening to her.
ESTH|2|12|Now when the turn came for each young woman to go in to King Ahasuerus, after being twelve months under the regulations for the women, since this was the regular period of their beautifying, six months with oil of myrrh and six months with spices and ointments for women-
ESTH|2|13|when the young woman went in to the king in this way, she was given whatever she desired to take with her from the harem to the king's palace.
ESTH|2|14|In the evening she would go in, and in the morning she would return to the second harem in custody of Shaashgaz, the king's eunuch, who was in charge of the concubines. She would not go in to the king again, unless the king delighted in her and she was summoned by name.
ESTH|2|15|When the turn came for Esther the daughter of Abihail the uncle of Mordecai, who had taken her as his own daughter, to go in to the king, she asked for nothing except what Hegai the king's eunuch, who had charge of the women, advised. Now Esther was winning favor in the eyes of all who saw her.
ESTH|2|16|And when Esther was taken to King Ahasuerus into his royal palace in the tenth month, which is the month of Tebeth, in the seventh year of his reign,
ESTH|2|17|the king loved Esther more than all the women, and she won grace and favor in his sight more than all the virgins, so that he set the royal crown on her head and made her queen instead of Vashti.
ESTH|2|18|Then the king gave a great feast for all his officials and servants; it was Esther's feast. He also granted a remission of taxes to the provinces and gave gifts with royal generosity.
ESTH|2|19|Now when the virgins were gathered together the second time, Mordecai was sitting at the king's gate.
ESTH|2|20|Esther had not made known her kindred or her people, as Mordecai had commanded her, for Esther obeyed Mordecai just as when she was brought up by him.
ESTH|2|21|In those days, as Mordecai was sitting at the king's gate, Bigthan and Teresh, two of the king's eunuchs, who guarded the threshold, became angry and sought to lay hands on King Ahasuerus.
ESTH|2|22|And this came to the knowledge of Mordecai, and he told it to Queen Esther, and Esther told the king in the name of Mordecai.
ESTH|2|23|When the affair was investigated and found to be so, the men were both hanged on the gallows. And it was recorded in the book of the chronicles in the presence of the king.
ESTH|3|1|After these things King Ahasuerus promoted Haman the Agagite, the son of Hammedatha, and advanced him and set his throne above all the officials who were with him.
ESTH|3|2|And all the king's servants who were at the king's gate bowed down and paid homage to Haman, for the king had so commanded concerning him. But Mordecai did not bow down or pay homage.
ESTH|3|3|Then the king's servants who were at the king's gate said to Mordecai, "Why do you transgress the king's command?"
ESTH|3|4|And when they spoke to him day after day and he would not listen to them, they told Haman, in order to see whether Mordecai's words would stand, for he had told them that he was a Jew.
ESTH|3|5|And when Haman saw that Mordecai did not bow down or pay homage to him, Haman was filled with fury.
ESTH|3|6|But he disdained to lay hands on Mordecai alone. So, as they had made known to him the people of Mordecai, Haman sought to destroy all the Jews, the people of Mordecai, throughout the whole kingdom of Ahasuerus.
ESTH|3|7|In the first month, which is the month of Nisan, in the twelfth year of King Ahasuerus, they cast Pur (that is, they cast lots) before Haman day after day; and they cast it month after month till the twelfth month, which is the month of Adar.
ESTH|3|8|Then Haman said to King Ahasuerus, "There is a certain people scattered abroad and dispersed among the peoples in all the provinces of your kingdom. Their laws are different from those of every other people, and they do not keep the king's laws, so that it is not to the king's profit to tolerate them.
ESTH|3|9|If it please the king, let it be decreed that they be destroyed, and I will pay 10,000 talents of silver into the hands of those who have charge of the king's business, that they may put it into the king's treasuries."
ESTH|3|10|So the king took his signet ring from his hand and gave it to Haman the Agagite, the son of Hammedatha, the enemy of the Jews.
ESTH|3|11|And the king said to Haman, "The money is given to you, the people also, to do with them as it seems good to you."
ESTH|3|12|Then the king's scribes were summoned on the thirteenth day of the first month, and an edict, according to all that Haman commanded, was written to the king's satraps and to the governors over all the provinces and to the officials of all the peoples, to every province in its own script and every people in its own language. It was written in the name of King Ahasuerus and sealed with the king's signet ring.
ESTH|3|13|Letters were sent by couriers to all the king's provinces with instruction to destroy, to kill, and to annihilate all Jews, young and old, women and children, in one day, the thirteenth day of the twelfth month, which is the month of Adar, and to plunder their goods.
ESTH|3|14|A copy of the document was to be issued as a decree in every province by proclamation to all the peoples to be ready for that day.
ESTH|3|15|The couriers went out hurriedly by order of the king, and the decree was issued in Susa the citadel. And the king and Haman sat down to drink, but the city of Susa was thrown into confusion.
ESTH|4|1|When Mordecai learned all that had been done, Mordecai tore his clothes and put on sackcloth and ashes, and went out into the midst of the city, and he cried out with a loud and bitter cry.
ESTH|4|2|He went up to the entrance of the king's gate, for no one was allowed to enter the king's gate clothed in sackcloth.
ESTH|4|3|And in every province, wherever the king's command and his decree reached, there was great mourning among the Jews, with fasting and weeping and lamenting, and many of them lay in sackcloth and ashes.
ESTH|4|4|When Esther's young women and her eunuchs came and told her, the queen was deeply distressed. She sent garments to clothe Mordecai, so that he might take off his sackcloth, but he would not accept them.
ESTH|4|5|Then Esther called for Hathach, one of the king's eunuchs, who had been appointed to attend her, and ordered him to go to Mordecai to learn what this was and why it was.
ESTH|4|6|Hathach went out to Mordecai in the open square of the city in front of the king's gate,
ESTH|4|7|and Mordecai told him all that had happened to him, and the exact sum of money that Haman had promised to pay into the king's treasuries for the destruction of the Jews.
ESTH|4|8|Mordecai also gave him a copy of the written decree issued in Susa for their destruction, that he might show it to Esther and explain it to her and command her to go to the king to beg his favor and plead with him on behalf of her people.
ESTH|4|9|And Hathach went and told Esther what Mordecai had said.
ESTH|4|10|Then Esther spoke to Hathach and commanded him to go to Mordecai and say,
ESTH|4|11|"All the king's servants and the people of the king's provinces know that if any man or woman goes to the king inside the inner court without being called, there is but one law- to be put to death, except the one to whom the king holds out the golden scepter so that he may live. But as for me, I have not been called to come in to the king these thirty days."
ESTH|4|12|And they told Mordecai what Esther had said.
ESTH|4|13|Then Mordecai told them to reply to Esther, "Do not think to yourself that in the king's palace you will escape any more than all the other Jews.
ESTH|4|14|For if you keep silent at this time, relief and deliverance will rise for the Jews from another place, but you and your father's house will perish. And who knows whether you have not come to the kingdom for such a time as this?"
ESTH|4|15|Then Esther told them to reply to Mordecai,
ESTH|4|16|"Go, gather all the Jews to be found in Susa, and hold a fast on my behalf, and do not eat or drink for three days, night or day. I and my young women will also fast as you do. Then I will go to the king, though it is against the law, and if I perish, I perish."
ESTH|4|17|Mordecai then went away and did everything as Esther had ordered him.
ESTH|5|1|On the third day Esther put on her royal robes and stood in the inner court of the king's palace, in front of the king's quarters, while the king was sitting on his royal throne inside the throne room opposite the entrance to the palace.
ESTH|5|2|And when the king saw Queen Esther standing in the court, she won favor in his sight, and he held out to Esther the golden scepter that was in his hand. Then Esther approached and touched the tip of the scepter.
ESTH|5|3|And the king said to her, "What is it, Queen Esther? What is your request? It shall be given you, even to the half of my kingdom."
ESTH|5|4|And Esther said, "If it please the king, let the king and Haman come today to a feast that I have prepared for the king."
ESTH|5|5|Then the king said, "Bring Haman quickly, so that we may do as Esther has asked." So the king and Haman came to the feast that Esther had prepared.
ESTH|5|6|And as they were drinking wine after the feast, the king said to Esther, "What is your wish? It shall be granted you. And what is your request? Even to the half of my kingdom, it shall be fulfilled."
ESTH|5|7|Then Esther answered, "My wish and my request is:
ESTH|5|8|If I have found favor in the sight of the king, and if it please the king to grant my wish and fulfill my request, let the king and Haman come to the feast that I will prepare for them, and tomorrow I will do as the king has said."
ESTH|5|9|And Haman went out that day joyful and glad of heart. But when Haman saw Mordecai in the king's gate, that he neither rose nor trembled before him, he was filled with wrath against Mordecai.
ESTH|5|10|Nevertheless, Haman restrained himself and went home, and he sent and brought his friends and his wife Zeresh.
ESTH|5|11|And Haman recounted to them the splendor of his riches, the number of his sons, all the promotions with which the king had honored him, and how he had advanced him above the officials and the servants of the king.
ESTH|5|12|Then Haman said, "Even Queen Esther let no one but me come with the king to the feast she prepared. And tomorrow also I am invited by her together with the king.
ESTH|5|13|Yet all this is worth nothing to me, so long as I see Mordecai the Jew sitting at the king's gate."
ESTH|5|14|Then his wife Zeresh and all his friends said to him, "Let a gallows fifty cubits high be made, and in the morning tell the king to have Mordecai hanged upon it. Then go joyfully with the king to the feast." This idea pleased Haman, and he had the gallows made.
ESTH|6|1|On that night the king could not sleep. And he gave orders to bring the book of memorable deeds, the chronicles, and they were read before the king.
ESTH|6|2|And it was found written how Mordecai had told about Bigthana and Teresh, two of the king's eunuchs, who guarded the threshold, and who had sought to lay hands on King Ahasuerus.
ESTH|6|3|And the king said, "What honor or distinction has been bestowed on Mordecai for this?" The king's young men who attended him said, "Nothing has been done for him."
ESTH|6|4|And the king said, "Who is in the court?" Now Haman had just entered the outer court of the king's palace to speak to the king about having Mordecai hanged on the gallows that he had prepared for him.
ESTH|6|5|And the king's young men told him, "Haman is there, standing in the court." And the king said, "Let him come in."
ESTH|6|6|So Haman came in, and the king said to him, "What should be done to the man whom the king delights to honor?" And Haman said to himself, "Whom would the king delight to honor more than me?"
ESTH|6|7|And Haman said to the king, "For the man whom the king delights to honor,
ESTH|6|8|let royal robes be brought, which the king has worn, and the horse that the king has ridden, and on whose head a royal crown is set.
ESTH|6|9|And let the robes and the horse be handed over to one of the king's most noble officials. Let them dress the man whom the king delights to honor, and let them lead him on the horse through the square of the city, proclaiming before him: 'Thus shall it be done to the man whom the king delights to honor.'"
ESTH|6|10|Then the king said to Haman, "Hurry; take the robes and the horse, as you have said, and do so to Mordecai the Jew who sits at the king's gate. Leave out nothing that you have mentioned."
ESTH|6|11|So Haman took the robes and the horse, and he dressed Mordecai and led him through the square of the city, proclaiming before him, "Thus shall it be done to the man whom the king delights to honor."
ESTH|6|12|Then Mordecai returned to the king's gate. But Haman hurried to his house, mourning and with his head covered.
ESTH|6|13|And Haman told his wife Zeresh and all his friends everything that had happened to him. Then his wise men and his wife Zeresh said to him, "If Mordecai, before whom you have begun to fall, is of the Jewish people, you will not overcome him but will surely fall before him."
ESTH|6|14|While they were yet talking with him, the king's eunuchs arrived and hurried to bring Haman to the feast that Esther had prepared.
ESTH|7|1|So the king and Haman went in to feast with Queen Esther.
ESTH|7|2|And on the second day, as they were drinking wine after the feast, the king again said to Esther, "What is your wish, Queen Esther? It shall be granted you. And what is your request? Even to the half of my kingdom, it shall be fulfilled."
ESTH|7|3|Then Queen Esther answered, "If I have found favor in your sight, O king, and if it please the king, let my life be granted me for my wish, and my people for my request.
ESTH|7|4|For we have been sold, I and my people, to be destroyed, to be killed, and to be annihilated. If we had been sold merely as slaves, men and women, I would have been silent, for our affliction is not to be compared with the loss to the king."
ESTH|7|5|Then King Ahasuerus said to Queen Esther, "Who is he, and where is he, who has dared to do this?"
ESTH|7|6|And Esther said, "A foe and enemy! This wicked Haman!" Then Haman was terrified before the king and the queen.
ESTH|7|7|And the king arose in his wrath from the wine-drinking and went into the palace garden, but Haman stayed to beg for his life from Queen Esther, for he saw that harm was determined against him by the king.
ESTH|7|8|And the king returned from the palace garden to the place where they were drinking wine, as Haman was falling on the couch where Esther was. And the king said, "Will he even assault the queen in my presence, in my own house?" As the word left the mouth of the king, they covered Haman's face.
ESTH|7|9|Then Harbona, one of the eunuchs in attendance on the king, said, "Moreover, the gallows that Haman has prepared for Mordecai, whose word saved the king, is standing at Haman's house, fifty cubits high."
ESTH|7|10|And the king said, "Hang him on that." So they hanged Haman on the gallows that he had prepared for Mordecai. Then the wrath of the king abated.
ESTH|8|1|On that day King Ahasuerus gave to Queen Esther the house of Haman, the enemy of the Jews. And Mordecai came before the king, for Esther had told what he was to her.
ESTH|8|2|And the king took off his signet ring, which he had taken from Haman, and gave it to Mordecai. And Esther set Mordecai over the house of Haman.
ESTH|8|3|Then Esther spoke again to the king. She fell at his feet and wept and pleaded with him to avert the evil plan of Haman the Agagite and the plot that he had devised against the Jews.
ESTH|8|4|When the king held out the golden scepter to Esther,
ESTH|8|5|Esther rose and stood before the king. And she said, "If it please the king, and if I have found favor in his sight, and if the thing seems right before the king, and I am pleasing in his eyes, let an order be written to revoke the letters devised by Haman the Agagite, the son of Hammedatha, which he wrote to destroy the Jews who are in all the provinces of the king.
ESTH|8|6|For how can I bear to see the calamity that is coming to my people? Or how can I bear to see the destruction of my kindred?"
ESTH|8|7|Then King Ahasuerus said to Queen Esther and to Mordecai the Jew, "Behold, I have given Esther the house of Haman, and they have hanged him on the gallows, because he intended to lay hands on the Jews.
ESTH|8|8|But you may write as you please with regard to the Jews, in the name of the king, and seal it with the king's ring, for an edict written in the name of the king and sealed with the king's ring cannot be revoked."
ESTH|8|9|The king's scribes were summoned at that time, in the third month, which is the month of Sivan, on the twenty-third day. And an edict was written, according to all that Mordecai commanded concerning the Jews, to the satraps and the governors and the officials of the provinces from India to Ethiopia, 127 provinces, to each province in its own script and to each people in its own language, and also to the Jews in their script and their language.
ESTH|8|10|And he wrote in the name of King Ahasuerus and sealed it with the king's signet ring. Then he sent the letters by mounted couriers riding on swift horses that were used in the king's service, bred from the royal stud,
ESTH|8|11|saying that the king allowed the Jews who were in every city to gather and defend their lives, to destroy, to kill, and to annihilate any armed force of any people or province that might attack them, children and women included, and to plunder their goods,
ESTH|8|12|on one day throughout all the provinces of King Ahasuerus, on the thirteenth day of the twelfth month, which is the month of Adar.
ESTH|8|13|A copy of what was written was to be issued as a decree in every province, being publicly displayed to all peoples, and the Jews were to be ready on that day to take vengeance on their enemies.
ESTH|8|14|So the couriers, mounted on their swift horses that were used in the king's service, rode out hurriedly, urged by the king's command. And the decree was issued in Susa the citadel.
ESTH|8|15|Then Mordecai went out from the presence of the king in royal robes of blue and white, with a great golden crown and a robe of fine linen and purple, and the city of Susa shouted and rejoiced.
ESTH|8|16|The Jews had light and gladness and joy and honor.
ESTH|8|17|And in every province and in every city, wherever the king's command and his edict reached, there was gladness and joy among the Jews, a feast and a holiday. And many from the peoples of the country declared themselves Jews, for fear of the Jews had fallen on them.
ESTH|9|1|Now in the twelfth month, which is the month of Adar, on the thirteenth day of the same, when the king's command and edict were about to be carried out, on the very day when the enemies of the Jews hoped to gain the mastery over them, the reverse occurred: the Jews gained mastery over those who hated them.
ESTH|9|2|The Jews gathered in their cities throughout all the provinces of King Ahasuerus to lay hands on those who sought their harm. And no one could stand against them, for the fear of them had fallen on all peoples.
ESTH|9|3|All the officials of the provinces and the satraps and the governors and the royal agents also helped the Jews, for the fear of Mordecai had fallen on them.
ESTH|9|4|For Mordecai was great in the king's house, and his fame spread throughout all the provinces, for the man Mordecai grew more and more powerful.
ESTH|9|5|The Jews struck all their enemies with the sword, killing and destroying them, and did as they pleased to those who hated them.
ESTH|9|6|In Susa the citadel itself the Jews killed and destroyed 500 men,
ESTH|9|7|and also killed Parshandatha and Dalphon and Aspatha
ESTH|9|8|and Poratha and Adalia and Aridatha
ESTH|9|9|and Parmashta and Arisai and Aridai and Vaizatha,
ESTH|9|10|the ten sons of Haman the son of Hammedatha, the enemy of the Jews, but they laid no hand on the plunder.
ESTH|9|11|That very day the number of those killed in Susa the citadel was reported to the king.
ESTH|9|12|And the king said to Queen Esther, "In Susa the citadel the Jews have killed and destroyed 500 men and also the ten sons of Haman. What then have they done in the rest of the king's provinces! Now what is your wish? It shall be granted you. And what further is your request? It shall be fulfilled."
ESTH|9|13|And Esther said, "If it please the king, let the Jews who are in Susa be allowed tomorrow also to do according to this day's edict. And let the ten sons of Haman be hanged on the gallows."
ESTH|9|14|So the king commanded this to be done. A decree was issued in Susa, and the ten sons of Haman were hanged.
ESTH|9|15|The Jews who were in Susa gathered also on the fourteenth day of the month of Adar and they killed 300 men in Susa, but they laid no hands on the plunder.
ESTH|9|16|Now the rest of the Jews who were in the king's provinces also gathered to defend their lives, and got relief from their enemies and killed 75,000 of those who hated them, but they laid no hands on the plunder.
ESTH|9|17|This was on the thirteenth day of the month of Adar, and on the fourteenth day they rested and made that a day of feasting and gladness.
ESTH|9|18|But the Jews who were in Susa gathered on the thirteenth day and on the fourteenth, and rested on the fifteenth day, making that a day of feasting and gladness.
ESTH|9|19|Therefore the Jews of the villages, who live in the rural towns, hold the fourteenth day of the month of Adar as a day for gladness and feasting, as a holiday, and as a day on which they send gifts of food to one another.
ESTH|9|20|And Mordecai recorded these things and sent letters to all the Jews who were in all the provinces of King Ahasuerus, both near and far,
ESTH|9|21|obliging them to keep the fourteenth day of the month Adar and also the fifteenth day of the same, year by year,
ESTH|9|22|as the days on which the Jews got relief from their enemies, and as the month that had been turned for them from sorrow into gladness and from mourning into a holiday; that they should make them days of feasting and gladness, days for sending gifts of food to one another and gifts to the poor.
ESTH|9|23|So the Jews accepted what they had started to do, and what Mordecai had written to them.
ESTH|9|24|For Haman the Agagite, the son of Hammedatha, the enemy of all the Jews, had plotted against the Jews to destroy them, and had cast Pur (that is, cast lots), to crush and to destroy them.
ESTH|9|25|But when it came before the king, he gave orders in writing that his evil plan that he had devised against the Jews should return on his own head, and that he and his sons should be hanged on the gallows.
ESTH|9|26|Therefore they called these days Purim, after the term Pur. Therefore, because of all that was written in this letter, and of what they had faced in this matter, and of what had happened to them,
ESTH|9|27|the Jews firmly obligated themselves and their offspring and all who joined them, that without fail they would keep these two days according to what was written and at the time appointed every year,
ESTH|9|28|that these days should be remembered and kept throughout every generation, in every clan, province, and city, and that these days of Purim should never fall into disuse among the Jews, nor should the commemoration of these days cease among their descendants.
ESTH|9|29|Then Queen Esther, the daughter of Abihail, and Mordecai the Jew gave full written authority, confirming this second letter about Purim.
ESTH|9|30|Letters were sent to all the Jews, to the 127 provinces of the kingdom of Ahasuerus, in words of peace and truth,
ESTH|9|31|that these days of Purim should be observed at their appointed seasons, as Mordecai the Jew and Queen Esther obligated them, and as they had obligated themselves and their offspring, with regard to their fasts and their lamenting.
ESTH|9|32|The command of Queen Esther confirmed these practices of Purim, and it was recorded in writing.
ESTH|10|1|King Ahasuerus imposed tax on the land and on the coastlands of the sea.
ESTH|10|2|And all the acts of his power and might, and the full account of the high honor of Mordecai, to which the king advanced him, are they not written in the Book of the Chronicles of the kings of Media and Persia?
ESTH|10|3|For Mordecai the Jew was second in rank to King Ahasuerus, and he was great among the Jews and popular with the multitude of his brothers, for he sought the welfare of his people and spoke peace to all his people.
