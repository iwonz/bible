EZEK|1|1|Et factum est in tricesimo anno, in quarto mense, in quinta men sis, cum essem in medio captivorum iuxta fluvium Chobar, aperti sunt caeli, et vidi visiones Dei.
EZEK|1|2|In quinta mensis, ipse est annus quintus transmigrationis regis Ioachin,
EZEK|1|3|factum est verbum Domini ad Ezechielem filium Buzi, sacerdotem, in terra Chaldaeorum secus flumen Chobar, et facta est super eum ibi manus Domini.
EZEK|1|4|Et vidi: et ecce ventus turbinis veniebat ab aquilone et nubes magna et ignis conglobatus, et splendor in circuitu eius, et de medio eius quasi species electri, id est de medio ignis;
EZEK|1|5|et ex medio eius similitudo quattuor animalium, et hic aspectus eorum: similitudo hominis erat eis.
EZEK|1|6|Quattuor facies uni et quattuor pennae uni;
EZEK|1|7|pedes eorum pedes recti, et planta pedis eorum quasi planta pedis vituli, et scintillabant quasi aspectus aeris candentis.
EZEK|1|8|Et manus hominis erant sub pennis eorum in quattuor partibus. Facies autem et pennae illorum quattuor:
EZEK|1|9|iunctae erant pennae eorum altera ad alteram; non revertebantur, cum incederent, sed unumquodque ante faciem suam gradiebatur.
EZEK|1|10|Similitudo autem vultus eorum: facies hominis et facies leonis a dextris ipsorum quattuor, facies autem bovis a sinistris ipsorum quattuor et facies aquilae ipsorum quattuor.
EZEK|1|11|Et pennae eorum extentae desuper; duae pennae singulorum iungebantur, et duae tegebant corpora eorum.
EZEK|1|12|Et unumquodque coram facie sua ambulabat: ubi erat impetus spiritus, illuc gradiebantur nec revertebantur, cum ambularent.
EZEK|1|13|Et in medio animalium, aspectus quasi carbonum ignis ardentium, quasi aspectus lampadarum discurrentium in medio animalium; et splendor erat ignis, et de igne fulgur egrediens.
EZEK|1|14|Et animalia ibant et revertebantur in similitudinem fulguris coruscantis.
EZEK|1|15|Cumque aspicerem animalia, apparuit rota una super terram iuxta singula animalia.
EZEK|1|16|Et aspectus rotarum et opus earum quasi species chrysolithi, et una similitudo ipsarum quattuor; et aspectus earum et opera, quasi sit rota in medio rotae.
EZEK|1|17|Per quattuor partes earum euntes ibant et non revertebantur, cum ambularent.
EZEK|1|18|Canthis autem earum erat altitudo et horribilis aspectus; et canthi earum erant oculis pleni in circuitu ipsarum quattuor.
EZEK|1|19|Cumque ambularent animalia, ambulabant pariter et rotae iuxta ea; et cum elevarentur animalia de terra, elevabantur simul et rotae.
EZEK|1|20|Quocumque impellebat spiritus ut irent, ibant, et rotae pariter levabantur sequentes eum; spiritus enim animalium erat in rotis.
EZEK|1|21|Cum euntibus ibant et cum stantibus stabant; et cum elevatis a terra pariter elevabantur, et rotae sequentes ea, quia spiritus animalium erat in rotis.
EZEK|1|22|Et similitudo super capita animalium firmamenti quasi aspectus crystalli horribilis et extenti super capita eorum desuper.
EZEK|1|23|Sub firmamento autem pennae eorum rectae altera ad alteram; unumquodque duabus alis velabat corpus suum.
EZEK|1|24|Et audiebam sonum alarum quasi sonum aquarum multarum, quasi sonum Omnipotentis: cum ambularent, erat strepitus vehemens ut sonus castrorum; cumque starent, demittebantur pennae eorum.
EZEK|1|25|Nam cum fieret vox supra firmamentum, quod erat super caput eorum, stabant et submittebant alas suas.
EZEK|1|26|Et super firmamentum, quod erat imminens capiti eorum, quasi aspectus lapidis sapphiri similitudo throni; et super similitudinem throni similitudo quasi aspectus hominis desuper.
EZEK|1|27|Et vidi quasi speciem electri, velut aspectum ignis per circuitum ab aspectu lumborum eius et desuper; et ab aspectu lumborum eius usque deorsum vidi quasi speciem ignis splendentis in circuitu.
EZEK|1|28|Velut aspectus arcus, cum fuerit in nube in die pluviae: sic erat aspectus splendoris per gyrum. Haec visio similitudinis gloriae Domini. Et vidi et cecidi in faciem meam et audivi vocem loquentis.
EZEK|2|1|Et dixit ad me: " Fili hominis, sta super pedes tuos, et loquar tecum ".
EZEK|2|2|Et ingressus est in me spiritus, postquam locutus est mihi et statuit me supra pedes meos, et audivi loquentem ad me
EZEK|2|3|et dicentem: " Fili hominis, mitto ego te ad filios Israel, ad gentes apostatrices, quae recesserunt a me; ipsi et patres eorum praevaricati sunt in me usque ad diem hanc.
EZEK|2|4|Et filii dura facie et obstinato corde sunt, ad quos ego mitto te; et dices ad eos: Haec dicit Dominus Deus.
EZEK|2|5|Ipsi sive audiant, sive contemnant - quoniam domus exasperans est - sciant tamen quia propheta fuerit in medio eorum.
EZEK|2|6|Tu ergo, fili hominis, ne timeas eos neque sermones eorum metuas, etsi cardui et spinae te circumdant, et cum scorpionibus habitas. Verba eorum ne timeas et vultus eorum ne formides, quia domus exasperans est.
EZEK|2|7|Loqueris ergo verba mea ad eos, sive audiant, sive contemnant, quoniam exasperantes sunt.
EZEK|2|8|Tu autem, fili hominis, audi, quaecumque loquor ad te, et noli esse exasperans, sicut domus exasperatrix est; aperi os tuum et comede, quaecumque ego do tibi ".
EZEK|2|9|Et vidi: et ecce manus missa ad me, in qua erat involutus liber; et expandit illum coram me, qui erat scriptus intus et foris, et scriptae erant in eo lamentationes et gemitus et vae.
EZEK|3|1|Et dixit ad me: " Fili hominis, quodcumque inveneris, comede; comede volumen istud et vadens loquere ad filios Israel ".
EZEK|3|2|Et aperui os meum, et cibavit me volumine illo
EZEK|3|3|et dixit ad me: " Fili hominis, venter tuus comedet, et viscera tua complebuntur volumine isto, quod ego do tibi ". Et comedi illud, et factum est in ore meo sicut mel dulce.
EZEK|3|4|Et dixit ad me: " Fili hominis, vade ad domum Israel et loqueris verba mea ad eos.
EZEK|3|5|Non enim ad populum profundi sermonis et ignotae linguae tu mitteris, ad domum Israel;
EZEK|3|6|neque ad populos multos profundi sermonis et ignotae linguae, quorum non possis audire sermones; et si ad illos mittereris, ipsi audirent te.
EZEK|3|7|Domus autem Israel nolunt audire te, quia nolunt audire me; omnis quippe domus Israel dura fronte est et obstinato corde.
EZEK|3|8|Ecce dedi faciem tuam valentiorem faciebus eorum et frontem tuam duriorem frontibus eorum;
EZEK|3|9|ut adamantem et duriorem silice dedi faciem tuam: ne timeas eos neque metuas a facie eorum, quia domus exasperans est ".
EZEK|3|10|Et dixit ad me: " Fili hominis, omnes sermones meos, quos loquor ad te, assume in corde tuo et auribus tuis audi.
EZEK|3|11|Et vade, ingredere ad transmigrationem, ad filios populi tui, et loqueris ad eos et dices eis: Haec dicit Dominus Deus; sive audiant, sive contemnant ".
EZEK|3|12|Et assumpsit me spiritus, et audivi post me vocem commotionis magnae, cum elevaretur gloria Domini de loco suo;
EZEK|3|13|et vocem alarum animalium percutientium alteram ad alteram et vocem rotarum sequentium animalia et vocem commotionis magnae.
EZEK|3|14|Spiritus quoque levavit me et assumpsit me; et abii amarus in indignatione spiritus mei: manus enim Domini erat super me gravis.
EZEK|3|15|Et veni ad transmigrationem, ad Telabib, ad eos, qui habitabant iuxta flumen Chobar; et sedi, ubi illi sedebant, et mansi ibi septem diebus obstupefactus in medio eorum.
EZEK|3|16|Cum autem pertransissent septem dies, factum est verbum Domini ad me dicens:
EZEK|3|17|" Fili hominis, speculatorem dedi te domui Israel; et audies de ore meo verbum et commonebis eos ex me.
EZEK|3|18|Si, dicente me ad impium: Morte morieris, non commonueris eum neque locutus fueris ei, ut avertatur a via sua impia et vivat, ipse impius in iniquitate sua morietur, sanguinem autem eius de manu tua requiram.
EZEK|3|19|Si autem tu commonueris impium, et ille non fuerit conversus ab impietate sua et a via sua impia, ipse quidem in iniquitate sua morietur, tu autem animam tuam liberasti.
EZEK|3|20|Sed et si conversus iustus a iustitia sua, fecerit iniquitatem, ponam offendiculum coram eo; ipse morietur, quia non commonuisti eum: in peccato suo morietur, et non erunt in memoria iustitiae eius, quas fecit; sanguinem vero eius de manu tua requiram.
EZEK|3|21|Si autem tu commonueris iustum, ut non peccet iustus, et ille non peccaverit, vivens vivet, quia commonuisti eum et tu animam tuam liberasti.
EZEK|3|22|Et facta est super me manus Domini, et dixit ad me: " Surgens egredere in campum, et ibi loquar tecum ".
EZEK|3|23|Et surgens egressus sum in campum, et ecce ibi gloria Domini stabat quasi gloria, quam vidi iuxta fluvium Chobar, et cecidi in faciem meam.
EZEK|3|24|Et ingressus est in me spiritus et statuit me super pedes meos et locutus est mihi et dixit ad me: " Ingredere et includere in medio domus tuae.
EZEK|3|25|Et tu, fili hominis, ecce data sunt super te vincula, et ligabunt te in eis, et non egredieris in medio eorum;
EZEK|3|26|et linguam tuam adhaerere faciam palato tuo, et eris mutus nec quasi vir obiurgans, quia domus exasperans est.
EZEK|3|27|Cum autem locutus fuero tibi, aperiam os tuum, et dices ad eos: Haec dicit Dominus Deus. Qui audit, audiat; et, qui contemnit, contemnat, quia domus exasperans est ".
EZEK|4|1|" Et tu, fili hominis, sume tibi laterem et pones eum coram te et describes in eo civitatem Ierusalem.
EZEK|4|2|Et ordinabis adversus eam obsidionem et aedificabis munitiones et comportabis aggerem et dabis contra eam castra et pones arietes in gyro.
EZEK|4|3|Et tu sume tibi sartaginem ferream et pones eam in murum ferreum inter te et inter civitatem; et obfirmabis faciem tuam ad eam, et erit in obsidionem, et circumdabis eam: signum est domui Israel.
EZEK|4|4|Et tu recumbes super latus tuum sinistrum et pones iniquitates domus Israel super eo; numero dierum, quibus recumbes super illud, assumes iniquitatem eorum.
EZEK|4|5|Ego autem dedi tibi annos iniquitatis eorum numero dierum trecentos et nonaginta dies, et portabis iniquitatem domus Israel.
EZEK|4|6|Et cum compleveris haec, recumbes super latus tuum dextrum secundo et assumes iniquitatem domus Iudae quadraginta diebus; diem pro anno, diem, inquam, pro anno dedi tibi.
EZEK|4|7|Et ad obsidionem Ierusalem convertes faciem tuam, et brachium tuum erit exsertum, et prophetabis adversus eam.
EZEK|4|8|Ecce circumdedi te vinculis, et non te convertes a latere tuo in latus aliud, donec compleas dies obsidionis tuae.
EZEK|4|9|Et tu sume tibi frumentum et hordeum et fabam et lentem et milium et far et mittes ea in vas unum et facies tibi panes numero dierum, quibus recumbes super latus tuum: trecentis et nonaginta diebus comedes illud.
EZEK|4|10|Cibus autem tuus, quo vesceris, erit in pondere viginti stateres in die; a tempore usque ad tempus comedes illud.
EZEK|4|11|Et aquam in mensura bibes, sextam partem hin; a tempore usque ad tempus bibes illud.
EZEK|4|12|Et quasi subcinericium hordeaceum comedes illud; et stercore, quod egreditur de homine, coques illud in oculis eorum".
EZEK|4|13|Et dixit Dominus: " Sic comedent filii Israel panem suum pollutum inter gentes, ad quas eiciam eos ".
EZEK|4|14|Et dixi: " Heu, Domine Deus, ecce anima mea non est polluta, et morticinum et laceratum a bestiis non comedi ab infantia mea usque nunc, et non est ingressa in os meum caro immunda ".
EZEK|4|15|Et dixit ad me: " Ecce dedi tibi fimum boum pro stercoribus humanis, et facies panem tuum in eo ".
EZEK|4|16|Et dixit ad me: " Fili hominis, ecce ego conteram baculum panis in Ierusalem, et comedent panem in pondere et in sollicitudine et aquam in mensura et in desolatione bibent,
EZEK|4|17|ut, deficientibus pane et aqua, desoletur unusquisque cum fratre suo, et contabescant in iniquitatibus suis.
EZEK|5|1|Et tu, fili hominis, sume tibi gladium acutum radentem pilos et assumes eum et duces per caput tuum et per barbam tuam et assumes tibi stateram ponderis et divides eos.
EZEK|5|2|Tertiam partem igne combures in medio civitatis, post completionem dierum obsidionis; et assumens tertiam partem, concides gladio in circuitu eius; tertiam vero aliam disperges in ventum, et gladium nudabo post eos.
EZEK|5|3|Et sumes inde parvum numerum et ligabis eos in summitate pallii tui;
EZEK|5|4|et ex eis rursum tolles et proicies eos in medio ignis et combures eos igne; ex eo egredietur ignis. Et dices ad omnem domum Israel:
EZEK|5|5|Haec dicit Dominus Deus: Ista est Ierusalem! In medio gentium posui eam et in circuitu eius terras.
EZEK|5|6|Et contempsit iudicia mea, ut plus esset impia quam gentes, et praecepta mea ultra quam terrae, quae in circuitu eius sunt: iudicia enim mea proiecerunt et in praeceptis meis non ambulaverunt.
EZEK|5|7|Idcirco haec dicit Dominus Deus: Quia tumultuati estis magis quam gentes, quae in circuitu vestro sunt, et in praeceptis meis non ambulastis et iudicia mea non fecistis et iuxta iudicia gentium, quae in circuitu vestro sunt, non estis operati,
EZEK|5|8|ideo haec dicit Dominus Deus: Ecce ego ad te et ipse ego faciam in medio tui iudicia in oculis gentium
EZEK|5|9|et faciam in te, quae non feci et quibus similia ultra non faciam, propter omnes abominationes tuas.
EZEK|5|10|Ideo patres comedent filios in medio tui, et filii comedent patres suos, et faciam in te iudicia et ventilabo universas reliquias tuas in omnem ventum.
EZEK|5|11|Idcirco vivo ego, dicit Dominus Deus, vere pro eo quod sanctum meum violasti in omnibus offensionibus tuis et in omnibus abominationibus tuis, ego quoque radam, et non parcet oculus meus, et non miserebor.
EZEK|5|12|Tertia tui pars peste morietur et fame consumetur in medio tui, et tertia tui pars in gladio cadet in circuitu tuo, tertiam vero partem tuam in omnem ventum dispergam et gladium evaginabo post eos.
EZEK|5|13|Et complebo furorem meum et requiescere faciam indignationem meam in eis et consolabor; et scient quia ego Dominus locutus sum in zelo meo, cum implevero indignationem meam in eis.
EZEK|5|14|Et dabo te in desertum et in opprobrium in gentibus, quae in circuitu tuo sunt, in conspectu omnis praetereuntis;
EZEK|5|15|et eris opprobrium et blasphemia, exemplum et stupor in gentibus, quae in circuitu tuo sunt, cum fecero in te iudicia in furore et in indignatione et in castigationibus irae.
EZEK|5|16|Ego Dominus locutus sum. Quando misero sagittas famis pessimas in vos, quae erunt mortiferae, et quas mittam, ut destruam vos, et famem congregabo super vos et conteram vobis baculum panis;
EZEK|5|17|et immittam in vos famem et bestias pessimas, et absque liberis facient te, et pestilentia et sanguis transibunt per te, et gladium inducam super te. Ego Dominus locutus sum ".
EZEK|6|1|Et factus est sermo Domini ad me dicens:
EZEK|6|2|" Fili hominis, pone faciem tuam ad montes Israel et prophetabis ad eos
EZEK|6|3|et dices: Montes Israel, audite verbum Domini Dei. Haec dicit Dominus Deus montibus et collibus, voraginibus et vallibus: Ecce ego inducam super vos gladium et destruam excelsa vestra;
EZEK|6|4|et demoliar aras vestras, et confringentur delubra vestra, et deiciam interfectos vestros ante idola vestra.
EZEK|6|5|Et dabo cadavera filiorum Israel ante faciem simulacrorum vestrorum et dispergam ossa vestra circum aras vestras;
EZEK|6|6|in omnibus habitationibus vestris urbes desertae erunt, et excelsa demolientur, ut dissipentur et intereant arae vestrae, et confringantur et cessent idola vestra, et conterantur delubra vestra, et deleantur opera vestra.
EZEK|6|7|Et cadet interfectus in medio vestri, et scietis quia ego Dominus.
EZEK|6|8|Et relinquam in vobis eos, qui fugerint gladium in gentibus, cum dispersero vos in terris;
EZEK|6|9|et recordabuntur mei liberati vestri in gentibus, ad quas captivi ducti sunt, quia contrivi cor eorum fornicans et recedens a me, et oculos eorum fornicantes post idola sua; et displicebunt sibimet super malis, quae fecerunt in universis abominationibus suis,
EZEK|6|10|et scient quia ego Dominus non frustra locutus sum, ut facerem eis malum hoc.
EZEK|6|11|Haec dicit Dominus Deus: Plaude manu tua et percute pede tuo et dic: Heu ad omnes abominationes malas domus Israel, quia gladio, fame et peste ruituri sunt!
EZEK|6|12|Qui longe est, peste morietur; qui autem prope, gladio corruet; et, qui relictus fuerit et obsessus, fame morietur, et complebo indignationem meam in eis.
EZEK|6|13|Et scietis quia ego Dominus, cum fuerint interfecti eorum in medio idolorum suorum, in circuitu ararum suarum, in omni colle excelso, in cunctis summitatibus montium et subtus omne lignum nemorosum et subtus universam quercum frondosam, locum ubi obtulerunt tura redolentia universis idolis suis.
EZEK|6|14|Et extendam manum meam super eos et faciam terram desolatam et destitutam a deserto usque Rebla in omnibus habitationibus eorum, et scient quia ego Dominus ".
EZEK|7|1|Et factus est sermo Domini ad me dicens:
EZEK|7|2|" Et tu, fili hominis, loquere. Haec dicit Dominus Deus terrae Israel: Finis venit, finis super quattuor plagas terrae;
EZEK|7|3|nunc finis super te, et immittam furorem meum in te et iudicabo te iuxta vias tuas et ponam super te omnes abominationes tuas.
EZEK|7|4|Et non parcet oculus meus super te, et non miserebor, sed vias tuas ponam super te, et abominationes tuae in medio tui erunt, et scietis quia ego Dominus.
EZEK|7|5|Haec dicit Dominus Deus: Afflictio super afflictionem ecce venit.
EZEK|7|6|Finis venit, venit finis; evigilavit adversum te, ecce venit.
EZEK|7|7|Venit contractio super te, qui habitas in terra; venit tempus, prope est dies turbationis et non iubilationis in montibus.
EZEK|7|8|Nunc de propinquo effundam iram meam super te et complebo furorem meum in te et iudicabo te iuxta vias tuas et imponam tibi omnia scelera tua;
EZEK|7|9|et non parcet oculus meus, nec miserebor, sed vias tuas imponam tibi, et abominationes tuae in medio tui erunt, et scietis quia ego sum Dominus percutiens.
EZEK|7|10|Ecce dies, ecce venit; egressa est contractio, floruit iniustitia, germinavit superbia;
EZEK|7|11|violentia surrexit, ut esset virga impietatis: non ex eis et non ex pompa eorum neque ex sonitu eorum; et non erit requies in eis.
EZEK|7|12|Venit tempus, appropinquavit dies: qui emit, non laetetur; et, qui vendit, non lugeat, quia ira super omnem pompam eius.
EZEK|7|13|Quia, qui vendit, ad id quod vendidit non revertetur, cum adhuc sit in viventibus vita eorum. Visio enim ad omnem pompam eius non regredietur, et unusquisque in iniquitate sua vitam suam non confortabit.
EZEK|7|14|Canite tuba, praeparentur omnia, sed non est qui vadat ad proelium; ira enim mea super universam pompam eius.
EZEK|7|15|Gladius foris, pestis et fames intrinsecus. Qui in agro est, gladio morietur; et, qui in civitate, fame et pestilentia devorabuntur.
EZEK|7|16|Et salvabuntur, qui fugerint ex eis, et erunt in montibus quasi columbae convallium omnes gementes, unusquisque in iniquitate sua.
EZEK|7|17|Omnes manus dissolventur, et omnia genua fluent aquis.
EZEK|7|18|Et accingent se ciliciis, et operiet eos formido; et in omni facie confusio, et in universis capitibus eorum calvitium.
EZEK|7|19|Argentum suum foras proicient, et aurum eorum in immunditiam erit; argentum eorum et aurum eorum non valebit liberare eos in die furoris Domini; animam suam non saturabunt, et ventres eorum non implebuntur, quia scandalum iniquitatis eorum factum est,
EZEK|7|20|et ornamentum monilium suorum in superbiam posuerunt et imagines abominationum suarum et simulacrorum fecerunt ex eo; propter hoc dedi eis illud in immunditiam.
EZEK|7|21|Et dabo illud in manus alienorum ad diripiendum et impiis terrae in praedam, et contaminabunt illud.
EZEK|7|22|Et avertam faciem meam ab eis, et violabunt thesaurum meum absconditum; et introibunt in illud praedones et contaminabunt illud
EZEK|7|23|et facient ex illo catenas; quoniam terra plena est iudicio sanguinum, et civitas plena iniquitate.
EZEK|7|24|Et adducam pessimos de gentibus, et possidebunt domos eorum; et quiescere faciam superbiam potentium, et possidebunt sanctuaria eorum.
EZEK|7|25|Angustia superveniente, requirent pacem, et non erit.
EZEK|7|26|Calamitas super calamitatem veniet, et auditus super auditum; et quaerent visionem de propheta, et lex peribit a sacerdote, et consilium a senioribus.
EZEK|7|27|Rex lugebit, et princeps induetur horrore, et manus populi terrae conturbabuntur. Secundum viam eorum faciam eis et secundum iudicia eorum iudicabo eos, et scient quia ego Dominus ".
EZEK|8|1|Et factum est in anno sexto, in sexto mense, in quinta mensis, ego sedebam in domo mea, et senes Iudae sedebant coram me, et cecidit super me ibi manus Domini Dei,
EZEK|8|2|et vidi: et ecce similitudo quasi aspectus viri, ab aspectu lumborum eius et deorsum ignis, et a lumbis eius et sursum quasi aspectus splendoris ut visio electri.
EZEK|8|3|Emisit similitudinem manus et apprehendit me in cincinno capitis mei; et elevavit me spiritus inter terram et caelum et adduxit in Ierusalem, in visionibus Dei, iuxta ostium interius, quod respiciebat aquilonem, ubi erat statutum idolum zeli ad provocandam aemulationem.
EZEK|8|4|Et ecce ibi gloria Dei Israel secundum visionem, quam videram in campo;
EZEK|8|5|et dixit ad me: " Fili hominis, leva oculos tuos ad viam aquilonis ". Et levavi oculos meos ad viam aquilonis, et ecce ab aquilone portae altaris hoc idolum zeli in introitu.
EZEK|8|6|Et dixit ad me: " Fili hominis, putasne vides tu, quid isti faciunt, abominationes magnas, quas domus Israel facit hic, ut procul recedam a sanctuario meo? Et adhuc conversus videbis abominationes maiores ".
EZEK|8|7|Et duxit me ad ostium atrii, et vidi: et ecce foramen unum in pariete.
EZEK|8|8|Et dixit ad me: "Fili hominis, fode parietem"; et cum perfodissem parietem, apparuit ostium unum.
EZEK|8|9|Et dixit ad me: " Ingredere et vide abominationes pessimas, quas isti faciunt hic ".
EZEK|8|10|Et ingressus vidi: et ecce omnis similitudo reptilium et animalium abominatio et universa idola domus Israel depicta erant in pariete in circuitu per totum;
EZEK|8|11|et septuaginta viri de senioribus domus Israel, et Iezonias filius Saphan stabat in medio eorum stantium ante picturas, et unusquisque habebat turibulum in manu sua, et vapor nebulae de ture consurgebat.
EZEK|8|12|Et dixit ad me: " Certe vides, fili hominis, quae seniores domus Israel faciunt in tenebris, unusquisque in cubiculo simulacri sui; dicunt enim: Non videt Dominus nos, dereliquit Dominus terram"".
EZEK|8|13|Et dixit ad me: " Adhuc videbis abominationes maiores, quas isti faciunt ".
EZEK|8|14|Et duxit me ad ostium portae domus Domini, quod respiciebat ad aquilonem, et ecce ibi mulieres sedebant plangentes Thammuz.
EZEK|8|15|Et dixit ad me: "Certe vidisti, fili hominis; adhuc videbis abominationes maiores his ".
EZEK|8|16|Et introduxit me in atrium domus Domini interius, et ecce in ostio templi Domini, inter vestibulum et altare, quasi viginti quinque viri dorsa habentes contra templum Domini et facies ad orientem, et adorabant ad ortum solis.
EZEK|8|17|Et dixit ad me: " Certe vidisti, fili hominis; numquid parum est hoc domui Iudae, ut facerent abominationes istas, quas fecerunt hic, quia replentes terram iniquitate iterum irritaverunt me et ecce applicant ramum ad nares suas.
EZEK|8|18|Ergo et ego faciam in furore: non parcet oculus meus, nec miserebor et, cum clamaverint ad aures meas voce magna, non exaudiam eos ".
EZEK|9|1|Et clamavit in auribus meis voce magna dicens: " Appro pinquaverunt visitationes urbis, et unusquisque vas interfectionis habet in manu sua ".
EZEK|9|2|Et ecce sex viri veniebant de via portae superioris, quae respicit ad aquilonem, et uniuscuiusque vas interitus in manu eius; vir quoque unus in medio eorum vestitus lineis, et atramentarium scriptoris ad renes eius; et ingressi sunt et steterunt iuxta altare aereum.
EZEK|9|3|Et gloria Dei Israel elevata est de cherub, super quem erat, ad limen domus; et vocavit virum, qui indutus erat lineis et atramentarium scriptoris habebat in lumbis suis.
EZEK|9|4|Et dixit Dominus ad eum: " Transi per mediam civitatem in medio Ierusalem et signa thau super frontes virorum gementium et dolentium super cunctis abominationibus, quae fiunt in medio eius ".
EZEK|9|5|Et illis dixit, audiente me: " Transite per civitatem sequentes eum et percutite; non parcat oculus vester, neque misereamini:
EZEK|9|6|senem, adulescentulum et virginem et parvulum et mulieres interficite usque ad internecionem; omnem autem, super quem videritis thau, ne occidatis, et a sanctuario meo incipite ". Coeperunt ergo a viris senioribus, qui erant ante faciem domus.
EZEK|9|7|Et dixit ad eos: "Contaminate domum et implete atria interfectis. Egredimini ". Et egressi sunt et percutiebant eos, qui erant in civitate.
EZEK|9|8|Et caede completa, remansi ego ruique super faciem meam et clamans aio: Heu, Domine Deus! Ergone disperdes omnes reliquias Israel, effundens furorem tuum super Ierusalem? ".
EZEK|9|9|Et dixit ad me: " Iniquitas domus Israel et Iudae magna est nimis valde; et repleta est terra sanguinibus, et civitas repleta est iniustitia. Dixerunt enim: "Dereliquit Dominus terram, et Dominus non videt";
EZEK|9|10|igitur et meus non parcet oculus, neque miserebor: viam eorum super caput eorum reddam ".
EZEK|9|11|Et ecce vir, qui indutus erat lineis, qui habebat atramentarium in lumbis suis, respondit verbum dicens: " Feci, sicut praecepisti mihi ".
EZEK|10|1|Et vidi: et ecce super fir mamentum, quod erat super caput cherubim, quasi lapis sapphirus, quasi species similitudinis solii apparuit super ea.
EZEK|10|2|Et dixit ad virum, qui indutus erat lineis, et ait: " Ingredere in medio rotarum, quae sunt subtus cherub, et imple manus tuas prunis ignis, quae sunt inter cherubim, et effunde super civitatem ". Ingressusque est in conspectu meo.
EZEK|10|3|Cherubim autem stabant a dextris domus, cum ingrederetur vir, et nubes implevit atrium interius.
EZEK|10|4|Et elevata est gloria Domini desuper cherub ad limen domus, et repleta est domus nube, et atrium repletum est splendore gloriae Domini.
EZEK|10|5|Et sonitus alarum cherubim audiebatur usque ad atrium exterius, quasi vox Dei omnipotentis loquentis.
EZEK|10|6|Cumque praecepisset viro, qui indutus erat lineis, dicens: " Sume ignem de medio rotarum, de medio cherubim ", ingressus ille stetit iuxta rotam;
EZEK|10|7|et extendit cherub manum de medio cherubim ad ignem, qui erat inter cherubim, et sumpsit et dedit in manus eius, qui indutus erat lineis; qui accipiens egressus est.
EZEK|10|8|Et apparuit in cherubim similitudo manus hominis subtus pennas eorum,
EZEK|10|9|et vidi: et ecce quattuor rotae iuxta cherubim; rota una iuxta cherub unum, et rota alia iuxta cherub unum, species autem rotarum erat quasi species lapidis chrysolithi,
EZEK|10|10|et aspectus earum similitudo una illis quattuor, quasi sit rota in medio rotae.
EZEK|10|11|Cumque ambularent in quattuor partes, gradiebantur et non convertebantur ambulantes, sed ad locum, ad quem ire declinabat quae prima erat, sequebantur et ceterae nec convertebantur, cum ambularent.
EZEK|10|12|Et omne corpus eorum et terga et manus et pennae et rotae plena erant oculis in circuitu illis quattuor;
EZEK|10|13|et rotae istae vocatae sunt Volubiles, audiente me.
EZEK|10|14|Quattuor autem facies habebat unumquodque: facies prima facies cherub, et facies secunda facies hominis, et tertia facies leonis, et quarta facies aquilae.
EZEK|10|15|Et elevati sunt cherubim: ipsum est animal, quod videram iuxta fluvium Chobar.
EZEK|10|16|Cumque ambularent, cherubim ibant pariter, et rotae iuxta ea; et cum elevarent cherubim alas suas, ut exaltarentur de terra, non convertebantur rotae, sed et ipsae iuxta erant.
EZEK|10|17|Stantibus illis, stabant et cum elevatis elevabantur; spiritus enim animalium erat in eis.
EZEK|10|18|Et egressa est gloria Domini a limine templi et stetit super cherubim;
EZEK|10|19|et elevantes cherubim alas suas exaltata sunt a terra coram me, et, illis egredientibus, rotae quoque subsecutae sunt; et stetit in introitu portae domus Domini orientalis, et gloria Dei Israel erat super eos.
EZEK|10|20|Ipsum est animal, quod vidi subter Deum Israel iuxta fluvium Chobar, et intellexi quia cherubim essent.
EZEK|10|21|Quattuor per quattuor vultus unicuique, et quattuor alae unicuique, et similitudo manus hominis sub alis eorum;
EZEK|10|22|et similitudo vultuum eorum, ipsi vultus quorum aspectum videram iuxta fluvium Chobar. Et singuli ante faciem suam gradiebantur.
EZEK|11|1|Et elevavit me spiritus et duxit me ad portam domus Domini orientalem, quae respicit solis ortum; et ecce in introitu portae viginti quinque viri, et vidi in medio eorum Iezoniam filium Azur et Pheltiam filium Banaiae, principes populi.
EZEK|11|2|Dixitque ad me: " Fili hominis, hi sunt viri, qui cogitant iniquitatem et tractant consilium pessimum in urbe ista
EZEK|11|3|dicentes: "Nonne dudum aedificatae sunt domus? Haec est lebes, nos autem carnes".
EZEK|11|4|Idcirco vaticinare de eis; vaticinare, fili hominis ".
EZEK|11|5|Et irruit in me spiritus Domini et dixit ad me: " Loquere. Haec dicit Dominus: Sic locuti estis, domus Israel, et cogitationes cordis vestri ego novi.
EZEK|11|6|Plurimos occidistis in urbe hac et implestis vias eius interfectis.
EZEK|11|7|Propterea haec dicit Dominus Deus: Interfecti vestri, quos posuistis in medio eius, hi sunt carnes, et haec est lebes, et educam vos de medio eius.
EZEK|11|8|Gladium metuitis, et gladium inducam super vos, ait Dominus Deus.
EZEK|11|9|Et eiciam vos de medio eius daboque vos in manu hostium et faciam in vobis iudicia.
EZEK|11|10|Gladio cadetis, in finibus Israel iudicabo vos, et scietis quia ego Dominus.
EZEK|11|11|Haec non erit vobis in lebetem, et vos non eritis in medio eius in carnes: in finibus Israel iudicabo vos;
EZEK|11|12|et scietis quia ego Dominus, qui in praeceptis meis non ambulastis et iudicia mea non fecistis, sed iuxta iudicia gentium, quae in circuitu vestro sunt, estis operati ".
EZEK|11|13|Et factum est cum prophetarem, Pheltias filius Banaiae mortuus est; et cecidi in faciem meam, clamans voce magna, et dixi: " Heu, Domine Deus, consummationem tu facis reliquiarum Israel! ".
EZEK|11|14|Et factum est verbum Domini ad me dicens:
EZEK|11|15|" Fili hominis, fratres tui, fratres tui, viri propinqui tui et omnis domus Israel, universi, quibus dixerunt habitatores Ierusalem: "Longe sunt a Domino; nobis data est terra in possessionem".
EZEK|11|16|Propterea haec dicit Dominus Deus: Quia longe feci eos in gentibus et quia dispersi eos in terris, ero eis in sanctificationem modicam in terris, ad quas venerunt.
EZEK|11|17|Propterea loquere: Haec dicit Dominus Deus: Congregabo vos de populis et adunabo de terris, in quibus dispersi estis, daboque vobis humum Israel.
EZEK|11|18|Et ingredientur illuc et auferent omnes offensiones cunctasque abominationes eius de illa.
EZEK|11|19|Et dabo eis cor aliud et spiritum novum tribuam in visceribus eorum; et auferam cor lapideum de carne eorum et dabo eis cor carneum,
EZEK|11|20|ut in praeceptis meis ambulent et iudicia mea custodiant faciantque ea et sint mihi in populum, et ego sim eis in Deum.
EZEK|11|21|Quorum cor post offendicula et abominationes suas ambulat, horum viam in capite suo ponam ", dicit Dominus Deus.
EZEK|11|22|Et elevaverunt cherubim alas suas, et rotae cum eis, et gloria Dei Israel erat super eos;
EZEK|11|23|et ascendit gloria Domini de medio civitatis stetitque super montem, qui est ad orientem urbis.
EZEK|11|24|Et spiritus levavit me adduxitque in Chaldaeam ad transmigrationem in visione in spiritu Dei; et sublata est a me visio, quam videram.
EZEK|11|25|Et locutus sum ad transmigrationem omnia verba Domini, quae ostenderat mihi.
EZEK|12|1|Et factus est sermo Domini ad me dicens:
EZEK|12|2|" Fili hominis, in medio domus exasperantis tu habitas, qui oculos habent ad videndum et non vident, et aures ad audiendum et non audiunt, quia domus exasperans est.
EZEK|12|3|Tu ergo, fili hominis, fac tibi vasa transmigrationis et transmigrabis per diem coram eis; transmigrabis autem de loco tuo ad locum alterum in conspectu eorum, si forte aspiciant, quia domus exasperans est.
EZEK|12|4|Et efferes foras vasa tua quasi vasa transmigrantis per diem in conspectu eorum; tu autem egredieris vespere coram eis, sicut egreditur migrans.
EZEK|12|5|Ante oculos eorum perfode tibi parietem et efferes per eum;
EZEK|12|6|in conspectu eorum in umeris portabis, in caligine efferes: faciem tuam velabis et non videbis terram, quia portentum dedi te domui Israel ".
EZEK|12|7|Feci ergo, sicut praeceperat mihi Dominus: vasa mea protuli quasi vasa transmigrantis per diem et vespere perfodi mihi parietem manu; et in caligine extuli in umeris portans in conspectu eorum.
EZEK|12|8|Et factus est sermo Domini ad me mane dicens:
EZEK|12|9|" Fili hominis, numquid non dixerunt ad te domus Israel, domus exasperans: "Quid tu facis?".
EZEK|12|10|Dic ad eos: Haec dicit Dominus Deus: Super ducem onus istud, qui est in Ierusalem, et super omnem domum Israel, quae est in medio eius.
EZEK|12|11|Dic: Ego portentum vestrum. Quomodo feci, sic fiet illis: in transmigrationem et in captivitatem ibunt.
EZEK|12|12|Et dux, qui est in medio eorum, in umeris portabit, in caligine, et egredietur; parietem perfodient, ut transitus fiat per eum; faciem suam operiet, ut non videat oculo terram.
EZEK|12|13|Et extendam rete meum super illum, et capietur in tendicula mea; et adducam eum in Babylonem in terram Chaldaeorum, et ipsam non videbit ibique morietur.
EZEK|12|14|Et omnes, qui circa eum sunt, praesidium eius et agmina eius, dispergam in omnem ventum; et gladium evaginabo post eos.
EZEK|12|15|Et scient quia ego Dominus, quando dispersero illos in gentibus et disseminavero eos in terris.
EZEK|12|16|Et relinquam ex eis viros paucos a gladio et fame et pestilentia, ut narrent omnia scelera eorum in gentibus, ad quas ingredientur, et scient quia ego Dominus ".
EZEK|12|17|Et factus est sermo Domini ad me dicens:
EZEK|12|18|" Fili hominis, panem tuum in conturbatione comede; sed et aquam tuam in trepidatione et sollicitudine bibe.
EZEK|12|19|Et dices ad populum terrae: Haec dicit Dominus Deus ad eos, qui habitant in Ierusalem in terra Israel: Panem suum in sollicitudine comedent et aquam suam in desolatione bibent, quia desolabitur terra a plenitudine sua propter violentiam omnium, qui habitant in ea;
EZEK|12|20|et civitates, quae nunc habitantur, desolatae erunt, terraque deserta, et scietis quia ego Dominus ".
EZEK|12|21|Et factus est sermo Domini ad me dicens:
EZEK|12|22|" Fili hominis, quod est proverbium istud vobis in terra Israel dicentibus: "In longum differentur dies, et peribit omnis visio"?
EZEK|12|23|Ideo dic ad eos: Haec dicit Dominus Deus: Quiescere faciam proverbium istud, neque vulgo dicetur ultra in Israel; et loquere ad eos quod appropinquaverint dies et sermo omnis visionis.
EZEK|12|24|Non enim erit ultra omnis visio vana neque divinatio ambigua in medio filiorum Israel,
EZEK|12|25|quia ego Dominus loquar; quodcumque locutus fuero verbum, et fiet: non prolongabitur amplius, sed in diebus vestris, domus exasperans, loquar verbum et faciam illud ", dicit Dominus Deus.
EZEK|12|26|Et factus est sermo Domini ad me dicens:
EZEK|12|27|" Fili hominis, ecce domus Israel dicentium: "Visio, quam hic videt, in dies multos et in tempora longa iste prophetat";
EZEK|12|28|propterea dic ad eos: Haec dicit Dominus Deus: Non differetur ultra omnis sermo meus; verbum, quod locutus fuero, complebitur ", dicit Dominus Deus.
EZEK|13|1|Et factus est sermo Domini ad me dicens:
EZEK|13|2|" Fili hominis, vaticinare ad prophetas Israel, qui prophetant; et dices prophetantibus de corde suo: Audite verbum Domini.
EZEK|13|3|Haec dicit Dominus Deus: Vae prophetis insipientibus, qui sequuntur spiritum suum et nihil vident!
EZEK|13|4|Quasi vulpes in ruinis prophetae tui, Israel, facti sunt.
EZEK|13|5|Non ascendistis confractiones neque opposuistis murum pro domo Israel, ut staretis in proelio in die Domini.
EZEK|13|6|Vident vana et divinant mendacium dicentes: "Ait Dominus", cum Dominus non miserit eos; et exspectant, ut confirmet sermonem.
EZEK|13|7|Numquid non visionem cassam vidistis et divinationem mendacem locuti estis, et dicitis: "Ait Dominus", cum ego non sim locutus?
EZEK|13|8|Propterea haec dicit Dominus Deus: Quia locuti estis vana et vidistis mendacium, ideo ecce ego ad vos, ait Dominus Deus;
EZEK|13|9|et erit manus mea super prophetas, qui vident vana et divinant mendacium: in consilio populi mei non erunt et in scriptura domus Israel non scribentur nec in terram Israel ingredientur, et scietis quia ego Dominus Deus.
EZEK|13|10|Eo quod deceperint populum meum dicentes: "Pax", et non est pax; et ipse aedificabat parietem, illi autem liniebant eum calce.
EZEK|13|11|Dic ad eos, qui liniunt calce, quod casurus sit; erit enim imber inundans, et dabo lapides grandinis desuper irruentes et ventum procellae dissipantem.
EZEK|13|12|Siquidem ecce cecidit paries; numquid non dicetur vobis: "Ubi est litura, quam levistis?".
EZEK|13|13|Propterea haec dicit Dominus Deus: Et erumpere faciam spiritum tempestatum in indignatione mea, et imber inundans in furore meo erit, et lapides grandinis in ira in consumptionem;
EZEK|13|14|et destruam parietem, quem levistis calce, et adaequabo eum terrae, et revelabitur fundamentum eius, et cadet, et consumemini in medio eius et scietis quia ego sum Dominus.
EZEK|13|15|Et complebo indignationem meam in pariete et in his, qui leverunt eum calce, dicamque vobis: Non est paries, et non sunt qui leverunt eum;
EZEK|13|16|prophetae Israel, qui prophetant ad Ierusalem et vident ei visionem pacis, et non est pax, ait Dominus Deus.
EZEK|13|17|Et tu, fili hominis, pone faciem tuam contra filias populi tui, quae prophetant de corde suo, et vaticinare super eas
EZEK|13|18|et dic: Haec dicit Dominus Deus: Vae, quae consuunt fascias pro omni articulo manus et faciunt velamina pro capite omnis staturae ad capiendas animas! Numquid capietis animas de populo meo et vivificabitis animas vobis?
EZEK|13|19|Et violastis me ad populum meum pro pugillo hordei et fragmento panis, ut interficeretis animas, quae mori non deberent, et vivificastis animas, quae non deberent vivere, mentientes populo meo credenti mendaciis.
EZEK|13|20|Propter hoc haec dicit Dominus Deus: Ecce ego ad fascias vestras, quibus vos capitis animas quasi volatilia, et disrumpam eas de brachiis vestris; et dimittam animas, quas vos cepistis, animas quasi volatilia,
EZEK|13|21|et disrumpam velamina vestra et liberabo populum meum de manu vestra, neque erunt ultra in manibus vestris ad praedandum, et scietis quia ego Dominus.
EZEK|13|22|Pro eo quod maerere fecistis cor iusti mendaciter, quem ego non contristavi, et confortastis manus impii, ut non reverteretur a via sua mala et viveret,
EZEK|13|23|propterea vana non videbitis et divinationes non divinabitis amplius, et eruam populum meum de manu vestra, et scietis quia ego Dominus ".
EZEK|14|1|Et venerunt ad me viri seniorum Israel et sederunt coram me.
EZEK|14|2|Et factus est sermo Domini ad me dicens:
EZEK|14|3|" Fili hominis, viri isti posuerunt idola sua in cordibus suis et scandalum iniquitatis suae statuerunt contra faciem suam; numquid interrogatus respondebo eis?
EZEK|14|4|Propter hoc loquere eis et dices ad eos: Haec dicit Dominus Deus: Omnis homo de domo Israel, qui posuerit idola sua in corde suo et scandalum iniquitatis suae statuerit contra faciem suam et venerit ad prophetam interrogans per eum me, ego Dominus respondebo ei per me pro multitudine idolorum suorum,
EZEK|14|5|ut capiam domum Israel in corde suo, quo recesserunt a me in cunctis idolis suis.
EZEK|14|6|Propterea dic ad domum Israel: Haec dicit Dominus Deus: Convertimini et recedite ab idolis vestris et ab universis contaminationibus vestris avertite facies vestras.
EZEK|14|7|Quia omnis homo de domo Israel et de advenis, quicumque advena fuerit in Israel, si alienatus fuerit a me et posuerit idola sua in corde suo et scandalum iniquitatis suae statuerit contra faciem suam et venerit ad prophetam, ut interroget per eum me, ego Dominus respondebo ei per me;
EZEK|14|8|et ponam faciem meam contra hominem illum et faciam eum in exemplum et in proberbium et disperdam eum de medio populi mei, et scietis quia ego Dominus.
EZEK|14|9|Et propheta cum erraverit et locutus fuerit verbum, ego Dominus decepi prophetam illum et extendam manum meam contra eum et delebo eum de medio populi mei Israel.
EZEK|14|10|Et portabunt iniquitatem suam: sicut iniquitas interrogantis, sic et iniquitas prophetae erit,
EZEK|14|11|ut non erret ultra domus Israel a me neque polluatur in universis praevaricationibus suis, sed sit mihi in populum, et ego sim eis in Deum, ait Dominus Deus.
EZEK|14|12|Et factus est sermo Domini ad me dicens:
EZEK|14|13|" Fili hominis, terra cum peccaverit mihi, ut praevaricetur praevaricans, extendam manum meam super eam et conteram virgam panis eius et immittam in eam famem et interficiam de ea hominem et iumentum;
EZEK|14|14|et si fuerint tres viri isti in medio eius, Noe, Danel et Iob, ipsi iustitia sua liberabunt animas suas, ait Dominus Deus.
EZEK|14|15|Quod si et bestias pessimas induxero super terram, ut absque liberis faciant eam, et fuerit deserta, in qua nullus pertranseat propter bestias,
EZEK|14|16|tres viri isti si fuerint in ea, vivo ego, dicit Dominus Deus, quia nec filios nec filias liberabunt, sed ipsi soli liberabuntur, terra autem desolabitur.
EZEK|14|17|Vel si gladium induxero super terram illam et dixero gladio: Transi per terram, et interfecero de ea hominem et iumentum,
EZEK|14|18|et tres viri isti fuerint in medio eius, vivo ego, dicit Dominus Deus, non liberabunt filios neque filias, sed ipsi soli liberabuntur.
EZEK|14|19|Vel si pestilentiam immisero super terram illam et effudero indignationem meam super eam in sanguine, ut auferam ex ea hominem et iumentum,
EZEK|14|20|et Noe et Danel et Iob fuerint in medio eius, vivo ego, dicit Dominus Deus, quia filium et filiam non liberabunt, sed ipsi iustitia sua liberabunt animas suas.
EZEK|14|21|Quoniam haec dicit Dominus Deus: Quod si et quattuor iudicia mea pessima, gladium et famem et bestias malas et pestilentiam misero in Ierusalem, ut interficiam de ea hominem et pecus,
EZEK|14|22|tamen relinquetur in ea salvatio educentium filios et filias: ecce ipsi egredientur ad vos, et videbitis viam eorum et opera eorum et consolabimini super malo, quod induxi in Ierusalem in omnibus, quae importavi super eam.
EZEK|14|23|Et consolabuntur vos, cum videritis viam eorum et opera eorum, et cognoscetis quod non frustra fecerim omnia, quae feci in ea ", ait Dominus Deus.
EZEK|15|1|Et factus est sermo Domini ad me dicens:
EZEK|15|2|" Fili hominis, quid habet lignum vitisprae omnibus lignis sarmentorum,quae sunt inter ligna silvarum?
EZEK|15|3|Numquid tolletur de ea lignum,ut fiat opus,aut fabricabitur de ea paxillus,ut dependeat in eo quodcumque vas?
EZEK|15|4|Ecce igni datum est in escam,utramque partem eius consumpsit ignis,et medietas eius adusta est;numquid utile erit ad opus?
EZEK|15|5|Etiam cum esset integrum,non erat aptum ad opus;quanto magis cum ignis illud devoraverit et combusserit,nihil ex eo fiet operis.
EZEK|15|6|Propterea haec dicit Dominus Deus:Quomodo lignum vitis inter ligna silvarum,quod dedi igni ad devorandum,sic tradam habitatores Ierusalem.
EZEK|15|7|Et ponam faciem meam in eos:de igne egressi sunt,et ignis consumet eos.Et scietis quia ego Dominus,cum posuero faciem meam in eos
EZEK|15|8|et dedero terram inviam et desolatam,eo quod praevaricatores exstiterint ",dicit Dominus Deus.
EZEK|16|1|Et factus est sermo Domini ad me dicens:
EZEK|16|2|" Fili hominis, notas fac Ierusalem abominationes suas
EZEK|16|3|et dices: Haec dicit Dominus Deus ad Ierusalem: Radix tua et generatio tua de terra Chanaan, pater tuus Amorraeus et mater tua Hetthaea.
EZEK|16|4|Et quando nata es, in die ortus tui non est praecisus umbilicus tuus, et in aqua non es lota in emundationem nec sale salita nec involuta pannis.
EZEK|16|5|Non pepercit super te oculus, ut faceret tibi unum de his, miseratus tui, sed proiecta es super faciem terrae in abiectione animae tuae in die, qua nata es.
EZEK|16|6|Praeteriens autem te, vidi te palpitare in sanguine tuo et dixi tibi, cum esses in sanguine tuo: Vive. Dixi, inquam, tibi: In sanguine tuo vive.
EZEK|16|7|Crescentem quasi germen agri dedi te, et crevisti et grandis effecta es et pervenisti ad mundum muliebrem: ubera tua intumuerunt, et pilus tuus germinavit; sed eras nuda et confusione plena.
EZEK|16|8|Et transivi per te et vidi te; et ecce tempus tuum, tempus amantium. Et expandi amictum meum super te et operui ignominiam tuam; et iuravi tibi et ingressus sum pactum tecum, ait Dominus Deus, et facta es mea.
EZEK|16|9|Et lavi te aqua et emundavi sanguinem tuum ex te et unxi te oleo;
EZEK|16|10|et vestivi te discoloribus et calceavi te calceis corii delphini et cinxi te bysso et indui te serico.
EZEK|16|11|Et ornavi te ornamento et dedi armillas in manibus tuis et torquem circa collum tuum;
EZEK|16|12|et dedi inaurem super os tuum et circulos auribus tuis et coronam decoris in capite tuo.
EZEK|16|13|Et ornata es auro et argento et vestita es bysso et serico et multicoloribus. Similam et mel et oleum comedisti et decora facta es vehementer nimis et apta ad regnum.
EZEK|16|14|Et egressum est nomen tuum in gentes propter speciem tuam, quia perfecta eras in decore meo, quem posueram super te, dicit Dominus Deus.
EZEK|16|15|Et habens fiduciam in pulchritudine tua fornicata es in nomine tuo et exposuisti fornicationem tuam omni transeunti, quisquis fuerit.
EZEK|16|16|Et sumens de vestimentis tuis fecisti tibi excelsa variegata et fornicata es super eis, sicut non est factum neque futurum est.
EZEK|16|17|Et tulisti vasa decoris tui de auro meo atque argento meo, quae dedi tibi, et fecisti tibi imagines masculinas et fornicata es in eis.
EZEK|16|18|Et sumpsisti vestimenta tua multicoloria et operuisti illas et oleum meum et thymiama meum posuisti coram eis.
EZEK|16|19|Et panem meum, quem dedi tibi, similam et oleum et mel, quibus enutrivi te, posuisti in conspectu eorum in odorem suavitatis, et factum est, ait Dominus Deus.
EZEK|16|20|Et tulisti filios tuos et filias tuas, quas generasti mihi, et immolasti eis ad devorandum. Numquid parva est fornicatio tua?
EZEK|16|21|Immolasti filios meos et dedisti illos consecrans eis.
EZEK|16|22|Et post omnes abominationes tuas et fornicationes non es recordata dierum adulescentiae tuae, quando eras nuda et confusione plena, palpitans in sanguine tuo.
EZEK|16|23|Et accidit post omnem malitiam tuam - vae, vae tibi!, ait Dominus Deus
EZEK|16|24|et aedificasti tibi fornicem et fecisti tibi excelsum in cunctis plateis;
EZEK|16|25|ad omne caput viae aedificasti locum elevatum tuum et abominabilem fecisti decorem tuum et divisisti pedes tuos omni transeunti et multiplicasti fornicationes tuas.
EZEK|16|26|Et fornicata es cum filiis Aegypti vicinis tuis magnorum membrorum et multiplicasti fornicationem tuam ad irritandum me.
EZEK|16|27|Ecce ego extendi manum meam super te et imminui portionem tuam et dedi te in animam odientium te, filiarum Palaestinarum, quae erubescunt in via tua scelerata.
EZEK|16|28|Et fornicata es in filiis Assyriorum, eo quod necdum fueris expleta; et, postquam fornicata es, nec sic es satiata.
EZEK|16|29|Et multiplicasti fornicationem tuam usque ad terram mercatorum Chaldaeam, et nec sic satiata es.
EZEK|16|30|In quo mundabo cor tuum, ait Dominus Deus, cum faceres omnia haec opera mulieris meretricis et procacis?
EZEK|16|31|Quia fabricasti fornicem tuum in capite omnis viae et excelsum tuum fecisti in omni platea; nec facta es quasi meretrix, quia sprevisti pretium.
EZEK|16|32|Mulier adultera loco viri sui accipit alienos.
EZEK|16|33|Omnibus meretricibus dantur mercedes, tu autem dedisti mercedes cunctis amatoribus tuis et donabas eis, ut intrarent ad te undique ad fornicandum tecum.
EZEK|16|34|Factumque in te est contra consuetudinem mulierum in fornicationibus tuis, et post te non sunt fornicati; in eo enim quod dedisti mercedes et mercedes non accepisti, factum est in te contrarium.
EZEK|16|35|Propterea, meretrix, audi verbum Domini.
EZEK|16|36|Haec dicit Dominus Deus: Quia effusum est aes tuum, et revelata est ignominia tua in fornicationibus tuis ad amatores tuos et ad omnia idola abominabilia tua, in sanguine filiorum tuorum, quos dedisti eis,
EZEK|16|37|ideo ecce ego congregabo omnes amatores tuos, quibus iucunda fuisti, et omnes, quos dilexisti, cum universis, quos oderas; et congregabo eos super te undique et nudabo ignominiam tuam coram eis, et videbunt omnem turpitudinem tuam.
EZEK|16|38|Et iudicabo te iudiciis adulterarum et effundentium sanguinem et dabo te in sanguinem furoris et zeli.
EZEK|16|39|Et dabo te in manus eorum, et destruent fornicem tuum et demolientur excelsa tua et denudabunt te vestimentis tuis et auferent vasa decoris tui et derelinquent te nudam plenamque ignominia.
EZEK|16|40|Et convocabunt contra te congregationem et lapidabunt te lapidibus et trucidabunt te gladiis suis.
EZEK|16|41|Et comburent domos tuas igni et facient in te iudicia in oculis mulierum plurimarum; et faciam ut desinas fornicari, et mercedes ultra non dabis.
EZEK|16|42|Et satiabo indignationem meam in te, et auferetur zelus meus a te; et quiescam nec irascar amplius.
EZEK|16|43|Eo quod non fueris recordata dierum adulescentiae tuae et provocasti me in omnibus his, propterea et ego vias tuas in capite tuo dabo, ait Dominus Deus, et non feci iuxta scelera tua in omnibus abominationibus tuis.
EZEK|16|44|Ecce omnis, qui dicit vulgo proverbium in te, assumet illud dicens: Sicut mater, ita et filia eius".
EZEK|16|45|Filia matris tuae es tu, quae sprevit virum suum et filios suos; et soror sororum tuarum es tu, quae spreverunt viros suos et filios suos. Mater vestra Hetthaea, et pater vester Amorraeus.
EZEK|16|46|Et soror tua maior Samaria, ipsa et filiae eius, quae habitat ad sinistram tuam; soror autem tua minor te, quae habitat a dextris tuis, Sodoma et filiae eius.
EZEK|16|47|Sed nec in viis earum ambulasti neque secundum scelera earum fecisti; quasi parum fuisset, sceleratiora fecisti illis in omnibus viis tuis.
EZEK|16|48|Vivo ego, dicit Dominus Deus, non fecit Sodoma soror tua, ipsa et filiae eius, sicut fecisti tu et filiae tuae.
EZEK|16|49|Ecce haec fuit iniquitas Sodomae, sororis tuae: superbia, saturitas panis et securum otium erat ei et filiabus eius, et manum egeni et pauperis non sustentabant;
EZEK|16|50|et elevatae sunt et fecerunt abominationes coram me, et abstuli eas, sicut vidisti.
EZEK|16|51|Et Samaria dimidium peccatorum tuorum non peccavit, sed vicisti eas sceleribus tuis et iustificasti sorores tuas in omnibus abominationibus tuis, quas operata es.
EZEK|16|52|Ergo et tu porta confusionem tuam, quae absolvisti sorores tuas peccatis tuis, sceleratius agens quam illae; iustificatae sunt enim a te. Ergo et tu confundere et porta ignominiam tuam, quae iustificasti sorores tuas.
EZEK|16|53|Et convertam sortem earum, sortem Sodomorum cum filiabus suis et sortem Samariae et filiarum eius; et convertam sortem tuam in medio earum,
EZEK|16|54|ut portes ignominiam tuam et confundaris in omnibus, quae fecisti consolans eas.
EZEK|16|55|Et soror tua Sodoma et filiae eius revertentur ad pristinum statum suum, et Samaria et filiae eius revertentur ad pristinum statum suum, et tu et filiae tuae revertimini ad pristinum statum vestrum.
EZEK|16|56|Nonne fuit Sodoma, soror tua, in fabulam in ore tuo in die superbiae tuae,
EZEK|16|57|antequam revelaretur malitia tua, sicut hoc tempore tu es in opprobrium filiarum Syriae et cunctarum in circuitu tuo filiarum Palaestinarum, quae ambiunt te per gyrum?
EZEK|16|58|Scelus tuum et ignominiam tuam tu portabis, ait Dominus.
EZEK|16|59|Quia haec dicit Dominus Deus: Et faciam tibi, sicut fecisti, qui despexisti iuramentum, ut irritum faceres pactum.
EZEK|16|60|Et recordabor ego pacti mei tecum in diebus adulescentiae tuae et suscitabo tibi pactum sempiternum.
EZEK|16|61|Et recordaberis viarum tuarum et confunderis, cum receperis sorores tuas te maiores cum minoribus tuis, et dabo eas tibi in filias sed non ex pacto tuo.
EZEK|16|62|Et suscitabo ego pactum meum tecum, et scies quia ego Dominus,
EZEK|16|63|ut recorderis et confundaris, et non sit tibi ultra aperire os prae confusione tua, cum placatus fuero tibi in omnibus, quae fecisti ", ait Dominus Deus.
EZEK|17|1|Et factum est verbum Do mini ad me dicens:
EZEK|17|2|"Fili ho minis, propone aenigma et narra parabolam ad domum Israel
EZEK|17|3|et dices:Haec dicit Dominus Deus:Aquila grandismagnarum alarum,longo pennarum ductu,plena plumis et varietate,venit ad Libanumet tulit cacumen cedri;
EZEK|17|4|summitatem frondium eius avellitet transportavit eam in terram Chanaan,in urbem negotiatorum posuit illam.
EZEK|17|5|Et tulit de semine terraeet posuit illud in terra pro semine,super aquas multas,quasi salicem posuit illud,
EZEK|17|6|ut germinaret et cresceret in vineam latioremhumili statura,respicientibus ramis eius ad illam,et radices eius sub illa essent.Facta est ergo vineaet fructificavit in palmiteset emisit propagines.
EZEK|17|7|Et fuit aquila altera grandis,magnis alismultisque plumis;et ecce vinea ista,quasi mittens radices suas ad eam,palmites suos extendit ad illam,ut irrigaret eam abundantiusquam areolae, in quibus erat plantata.
EZEK|17|8|In terra bonasuper aquas multasplantata est,ut faciat frondeset portet fructumet sit in vineam grandem.
EZEK|17|9|Dic: Haec dicit Dominus Deus:Ergone prosperabitur?Nonne radices eius evelletet fructum eius distringet,et marcescent omnia recentia germina eius, et arescet?Et non opus erit brachio grandi neque populo multo,ut evellat eam radicitus.
EZEK|17|10|Ecce plantata est; ergone prosperabitur?Nonne, cum tetigerit eam ventus urens,siccabituret in areis, in quibus germinaverat, arescet? ".
EZEK|17|11|Et factum est verbum Domini ad me dicens:
EZEK|17|12|" Dic ad domum exasperantem: Nescitis quid ista significent? Dic: Ecce venit rex Babylonis Ierusalem et assumpsit regem et principes eius et adduxit eos ad semetipsum in Babylonem;
EZEK|17|13|et tulit de semine regni pepigitque cum eo foedus et accepit ab eo iusiurandum, sed et fortes terrae sustulit,
EZEK|17|14|ut esset regnum humile et non elevaretur, sed custodiret pactum eius et servaret illud.
EZEK|17|15|Qui recedens ab eo, misit nuntios ad Aegyptum, ut daret sibi equos et populum multum. Numquid prosperabitur vel consequetur salutem, qui fecit haec? Et, qui dissolvit pactum, numquid effugiet?
EZEK|17|16|Vivo ego, dicit Dominus Deus, quoniam in loco regis, qui constituit eum regem, cuius fecit irritum iuramentum et solvit pactum, quod habebat cum eo, in medio Babylonis morietur.
EZEK|17|17|Et non in exercitu grandi neque in populo multo adiuvabit eum pharao in proelio, in iactu aggeris et in exstructione munitionum, ut interficiat animas multas.
EZEK|17|18|Spreverat enim iuramentum, ut solveret foedus, et ecce dedit manum suam et, cum omnia haec fecerit, non effugiet.
EZEK|17|19|Propterea haec dicit Dominus Deus: Vivo ego, quoniam iuramentum meum, quod sprevit, et foedus meum, quod praevaricatus est, ponam in caput eius
EZEK|17|20|et expandam super eum rete meum, et comprehendetur tendicula mea, et adducam eum in Babylonem et iudicabo illum ibi in praevaricatione, qua praevaricatus est in me.
EZEK|17|21|Et omnes electi eius in universo agmine suo gladio cadent; residui autem in omnem ventum dispergentur, et scietis quia ego Dominus locutus sum.
EZEK|17|22|Haec dicit Dominus Deus:Et sumam ego de cacumine cedri sublimis et ponam;de vertice ramorum eius tenerum distringamet plantabo super montem excelsum et eminentem.
EZEK|17|23|In monte sublimi Israel plantabo illud;et erumpet in germen et faciet fructumet erit in cedrum magnam;et habitabunt sub ea omnes volucres,et universum volatile sub umbra frondium eius nidificabit.
EZEK|17|24|Et scient omnia ligna regionisquia ego Dominushumiliavi lignum sublimeet exaltavi lignum humileet siccavi lignum virideet frondere feci lignum aridum.Ego Dominus locutus sum et feci ".
EZEK|18|1|Et factus est sermo Domini ad me dicens:
EZEK|18|2|"Quid est vo bis quod vulgo dicitis proverbium istud in terra Israel dicentes:Patres comederunt uvam acerbam,et dentes filiorum obstupescunt"?
EZEK|18|3|Vivo ego, dicit Dominus Deus, non dicetis ultra hoc proverbium in Israel.
EZEK|18|4|Ecce omnes animae meae sunt: ut anima patris, ita et anima filii mea est; anima, quae peccaverit, ipsa morietur.
EZEK|18|5|Et vir, si fuerit iustus et fecerit iudicium et iustitiam,
EZEK|18|6|in montibus non comederit et oculos suos non levaverit ad idola domus Israel et uxorem proximi sui non violaverit et ad mulierem menstruatam non accesserit
EZEK|18|7|et hominem non afflixerit, pignus debitori reddiderit, per vim nihil rapuerit, panem suum esurienti dederit et nudum operuerit vestimento,
EZEK|18|8|ad usuram non commodaverit et fenus non acceperit, ab iniquitate averterit manum suam, iudicium verum fecerit inter virum et virum,
EZEK|18|9|in praeceptis meis ambulaverit et iudicia mea custodierit, ut faciat veritatem, hic iustus est, vita vivet, ait Dominus Deus.
EZEK|18|10|Quod si genuerit filium latronem, effundentem sanguinem et facientem unum de istis,
EZEK|18|11|cum ipse haec omnia non fecerit, et etiam in montibus comedentem et uxorem proximi sui polluentem,
EZEK|18|12|egenum et pauperem affligentem, rapientem rapinas, pignus non reddentem et ad idola levantem oculos suos, abominationem facientem,
EZEK|18|13|ad usuram dantem et fenus accipientem, numquid vivet? Non vivet. Cum universa detestanda haec fecerit, morte morietur; sanguis eius in ipso erit.
EZEK|18|14|Quod si genuerit filium, qui videns omnia peccata patris sui, quae fecit, timuerit et non fecerit simile eis:
EZEK|18|15|super montes non comederit et oculos suos non levaverit ad idola domus Israel et uxorem proximi sui non violaverit
EZEK|18|16|et virum non afflixerit, pignus non retinuerit et rapinam non rapuerit, panem suum esurienti dederit et nudum operuerit vestimento,
EZEK|18|17|ab iniuria averterit manum suam, usuram et fenus non acceperit, iudicia mea fecerit, in praeceptis meis ambulaverit, hic non morietur in iniquitate patris sui, sed vita vivet.
EZEK|18|18|Pater eius, quia calumniatus est et fecit rapinas nec bonum operatus est in medio populi sui, ecce mortuus est in iniquitate sua.
EZEK|18|19|Et dicitis: "Quare non portavit filius iniquitatem patris?". Videlicet, quia filius iudicium et iustitiam operatus est, omnia praecepta mea custodivit et fecit illa, vivet vita.
EZEK|18|20|Anima, quae peccaverit, ipsa morietur; filius non portabit iniquitatem patris, et pater non portabit iniquitatem filii. Iustitia iusti super eum erit, et impietas impii erit super eum.
EZEK|18|21|Si autem impius egerit paenitentiam ab omnibus peccatis suis, quae operatus est, et custodierit universa praecepta mea et fecerit iudicium et iustitiam, vita vivet, non morietur.
EZEK|18|22|Omnes iniquitates eius, quas operatus est, non memorabuntur ei; in iustitia sua, quam operatus est, vivet.
EZEK|18|23|Numquid voluntatis meae est mors impii, dicit Dominus Deus, et non ut convertatur a viis suis et vivat?
EZEK|18|24|Si autem averterit se iustus a iustitia sua et fecerit iniquitatem secundum omnes abominationes, quas operari solet impius, numquid vivet? Omnes iustitiae eius, quas fecerat, non recordabuntur; in praevaricatione, qua praevaricatus est, et in peccato suo, quod peccavit, in ipsis morietur.
EZEK|18|25|Et dixistis: "Non est aequa via Domini". Audite ergo, domus Israel: Numquid via mea non est aequa, et non magis viae vestrae pravae sunt?
EZEK|18|26|Cum enim averterit se iustus a iustitia sua et fecerit iniquitatem, morietur; in iniustitia, quam operatus est, morietur.
EZEK|18|27|Et cum averterit se impius ab impietate sua, quam operatus est, et fecerit iudicium et iustitiam, ipse animam suam vivificabit;
EZEK|18|28|considerans enim et avertens se ab omnibus iniquitatibus suis, quas operatus est, vita vivet, non morietur.
EZEK|18|29|Et dicunt domus Israel: "Non est aequa via Domini". Numquid viae meae non sunt aequae, domus Israel, et non magis viae vestrae pravae?
EZEK|18|30|Idcirco unumquemque iuxta vias suas iudicabo, domus Israel, ait Dominus Deus. Convertimini et agite paenitentiam ab omnibus iniquitatibus vestris, et non erit vobis in scandalum iniquitatis.
EZEK|18|31|Proicite a vobis omnes praevaricationes vestras, in quibus praevaricati estis, et facite vobis cor novum et spiritum novum. Et quare moriemini, domus Israel?
EZEK|18|32|Quia nolo mortem morientis, dicit Dominus Deus. Revertimini et vivite.
EZEK|19|1|Et tu, assume planctum super principes Israel
EZEK|19|2|et dices:Qualis erat mater tua leaenainter leones!Cubavit in medio leunculorum,enutrivit catulos suos.
EZEK|19|3|Et educavit unum de leunculis suis;leo factus estet didicit capere praedam,homines devoravit.
EZEK|19|4|Et convocaverunt contra eum gentes,in fovea earum captus est;et adduxerunt eum in circulisin terram Aegypti.
EZEK|19|5|Quae cum vidisset quoniam exspectaverat,et perierat spes eius,tulit alium de leunculis suis,leonem constituit eum.
EZEK|19|6|Qui incedebat inter leones,factus est leoet didicit praedam capere,homines devoravit;
EZEK|19|7|et fregit arces eorumet civitates eorum vastavit.Et obstupuit terra et plenitudo eiusa voce rugitus illius.
EZEK|19|8|Et convenerunt adversum eum gentesundique de provinciiset expanderunt super eum rete suum,in fovea earum captus est.
EZEK|19|9|Et miserunt eum in caveam in circuliset adduxerunt eum ad regem Babylonis;qui misit eum in carcerem,ne audiretur vox eius ultrasuper montes Israel.
EZEK|19|10|Mater tua vineae assimilabatursuper aquam plantata.Fructus eius et frondes eius creveruntex aquis multis;
EZEK|19|11|et factae sunt ei virgae solidaein sceptra dominantium,et exaltata est statura eiususque in nubes,et apparuit in altitudine sua,in multitudine palmitum suorum.
EZEK|19|12|Et evulsa est in irain terramque proiecta,et ventus urens siccavit fructum eius;abrepta et arefacta est virga roboris eius,ignis comedit eam.
EZEK|19|13|Et nunc transplantata est in desertum,in terra invia et sitienti.
EZEK|19|14|Et egressus est ignis de virga ramorum eius,qui fructum eius comedit;et non fuit in ea virga fortis,sceptrum regni ".Planctus est, et erit in planctum.
EZEK|20|1|Et factum est in anno sep timo, in quinto mense, in de cima mensis, venerunt viri de senioribus Israel, ut interrogarent Dominum, et sederunt coram me.
EZEK|20|2|Et factus est sermo Domini ad me dicens:
EZEK|20|3|" Fili hominis, loquere senioribus Israel et dices ad eos: Haec dicit Dominus Deus: Num ad interrogandum me vos venistis? Vivo ego, quia non respondebo vobis, ait Dominus Deus.
EZEK|20|4|Numquid iudicabis eos, numquid iudicabis, fili hominis? Abominationes patrum eorum ostende eis.
EZEK|20|5|Et dices ad eos: Haec dicit Dominus Deus: In die qua elegi Israel et levavi manum meam pro stirpe domus Iacob et apparui eis in terra Aegypti et levavi manum meam pro eis dicens: Ego Dominus Deus vester;
EZEK|20|6|in die illa levavi manum meam pro eis, ut educerem eos de terra Aegypti in terram, quam provideram eis fluentem lacte et melle, quae est egregia inter omnes terras.
EZEK|20|7|Et dixi ad eos: Unusquisque abominationes oculorum suorum abiciat, et in idolis Aegypti nolite pollui: ego Dominus Deus vester.
EZEK|20|8|Et irritaverunt me nolueruntque me audire; unusquisque abominationes oculorum suorum non proiecit, nec idola Aegypti reliquerunt. Et dixi, ut effunderem indignationem meam super eos et consummarem iram meam in eis in medio terrae Aegypti.
EZEK|20|9|Et feci propter nomen meum, ut non violaretur coram gentibus, in quarum medio erant, et inter quas apparui eis, ut educerem eos de terra Aegypti.
EZEK|20|10|Eduxi ergo eos de terra Aegypti et duxi in desertum.
EZEK|20|11|Et dedi eis praecepta mea et iudicia mea ostendi eis, quae faciat homo et vivat in eis.
EZEK|20|12|Insuper et sabbata mea dedi eis, ut essent signum inter me et eos, et scirent quia ego Dominus sanctificans eos.
EZEK|20|13|Et irritaverunt me domus Israel in deserto: in praeceptis meis non ambulaverunt et iudicia mea proiecerunt, quae faciens homo vivet in eis, et sabbata mea violaverunt vehementer. Dixi ergo, ut effunderem furorem meum super eos in deserto et consumerem eos.
EZEK|20|14|Et feci propter nomen meum, ne violaretur coram gentibus, de quibus eduxi eos in conspectu earum.
EZEK|20|15|Attamen ego levavi quoque manum meam super eos in deserto, ne inducerem eos in terram, quam dedi eis fluentem lacte et melle, praecipuam terrarum omnium;
EZEK|20|16|quia iudicia mea proiecerunt et in praeceptis meis non ambulaverunt et sabbata mea violaverunt, post idola enim sua cor eorum gradiebatur.
EZEK|20|17|Et pepercit oculus meus super eos, ut non interficerem eos; nec consumpsi eos in deserto.
EZEK|20|18|Dixi autem ad filios eorum in solitudine: In praeceptis patrum vestrorum nolite incedere nec iudicia eorum custodiatis nec in idolis eorum polluamini.
EZEK|20|19|Ego Dominus Deus vester. In praeceptis meis ambulate et iudicia mea custodite et facite ea
EZEK|20|20|et sabbata mea sanctificate, ut sint signum inter me et vos, et sciatur quia ego Dominus Deus vester.
EZEK|20|21|Et exacerbaverunt me filii; in praeceptis meis non ambulaverunt et iudicia mea non custodierunt, ut facerent ea, quae cum fecerit homo, vivet in eis, et sabbata mea violaverunt. Et comminatus sum, ut effunderem furorem meum super eos et consummarem iram meam in eis in deserto.
EZEK|20|22|Averti autem manum meam et feci propter nomen meum, ut non violaretur coram gentibus, de quibus eduxi eos in oculis earum.
EZEK|20|23|Iterum levavi manum meam in eos in solitudine, ut dispergerem illos in nationes et ventilarem in terras,
EZEK|20|24|eo quod iudicia mea non fecissent et praecepta mea reprobassent et sabbata mea violassent et post idola patrum suorum fuissent oculi eorum.
EZEK|20|25|Ergo et ego dedi eis praecepta non bona et iudicia, in quibus non vivent;
EZEK|20|26|et pollui eos in muneribus suis, cum offerrent omne, quod aperit vulvam, ut horrorem eis incuterem, et sciant quia ego Dominus.
EZEK|20|27|Quam ob rem loquere ad domum Israel, fili hominis, et dices ad eos: Haec dicit Dominus Deus: Adhuc et in hoc blasphemaverunt me patres vestri, cum sprevissent me contemnentes,
EZEK|20|28|et induxissem eos in terram, super quam levavi manum meam, ut darem eis. Viderunt omnem collem excelsum et omne lignum nemorosum et immolaverunt ibi victimas suas et dederunt ibi irritationem oblationis suae et posuerunt ibi odorem suavitatis suae et libaverunt libationes suas.
EZEK|20|29|Et dixi ad eos: Quid est excelsum, ad quod vos ingredimini? Et vocatum est nomen eius Excelsum usque ad hanc diem.
EZEK|20|30|Propterea dic ad domum Israel: Haec dicit Dominus Deus: Certe in via patrum vestrorum vos polluimini et post offendicula eorum vos fornicamini
EZEK|20|31|et in oblatione donorum vestrorum, cum traducitis filios vestros per ignem; vos polluimini in omnibus idolis vestris usque hodie, et ego respondebo vobis, domus Israel? Vivo ego, dicit Dominus Deus, quia non respondebo vobis.
EZEK|20|32|Neque cogitatio mentis vestrae fiet dicentium: "Erimus sicut gentes et sicut cognationes terrarum, ut colamus ligna et lapides".
EZEK|20|33|Vivo ego, dicit Dominus Deus, quoniam in manu forti et brachio extento et in furore effuso regnabo super vos.
EZEK|20|34|Et educam vos de populis et congregabo vos de terris, in quibus dispersi estis; in manu valida et brachio extento et in furore effuso.
EZEK|20|35|Et adducam vos in desertum populorum et iudicio contendam vobiscum ibi facie ad faciem.
EZEK|20|36|Sicut iudicio contendi adversum patres vestros in deserto terrae Aegypti, sic iudicio contendam vobiscum, dicit Dominus Deus,
EZEK|20|37|et transire vos faciam sub baculo meo et inducam vos in vinculis foederis.
EZEK|20|38|Et segregabo de vobis transgressores et impios et de terra incolatus eorum educam eos, et terram Israel non ingredientur, et scietis quia ego Dominus.
EZEK|20|39|Et vos, domus Israel, haec dicit Dominus Deus: Singuli post idola vestra ambulate et servite eis. Sed postea nonne audietis me et nomen meum sanctum non polluetis ultra in muneribus vestris et in idolis vestris?
EZEK|20|40|In monte enim sancto meo, in monte excelso Israel, ait Dominus Deus, ibi serviet mihi omnis domus Israel: omnes, inquam, in terra, in qua placebunt mihi; et ibi quaeram donaria vestra et primitias oblationum vestrarum in omnibus sanctificationibus vestris.
EZEK|20|41|In odorem suavitatis suscipiam vos, cum eduxero vos de populis et congregavero vos de terris, in quas dispersi estis, et sanctificabor in vobis in oculis nationum.
EZEK|20|42|Et scietis quia ego Dominus, cum induxero vos ad terram Israel, in terram, pro qua levavi manum meam, ut darem eam patribus vestris.
EZEK|20|43|Et recordabimini ibi viarum vestrarum et omnium scelerum vestrorum, quibus polluti estis, et displicebitis vobis in conspectu vestro in omnibus malitiis vestris, quas fecistis.
EZEK|20|44|Et scietis quia ego Dominus, cum benefecero vobis propter nomen meum, non secundum vias vestras malas neque secundum scelera vestra pessima, domus Israel ", ait Dominus Deus.
EZEK|21|1|Et factus est sermo Domini ad me dicens:
EZEK|21|2|" Fili hominis, pone faciem tuam contra meridiem et stilla ad austrum et propheta ad saltum agri Nageb.
EZEK|21|3|Et dices saltui Nageb: Audi verbum Domini. Haec dicit Dominus Deus: Ecce ego succendam in te ignem, et comburet in te omne lignum viride et omne lignum aridum; non exstinguetur flamma succensionis, et comburetur in ea omnis facies ab austro usque ad aquilonem.
EZEK|21|4|Et videbit universa caro quia ego Domínus succendi eam, nec exstinguetur.
EZEK|21|5|Et dixi: " Heu, Domine Deus! Ipsi dicunt de me: "Numquid non per parabolas loquitur iste?" ".
EZEK|21|6|Et factus est sermo Domini ad me dicens:
EZEK|21|7|" Fili hominis, pone faciem tuam ad Ierusalem et stilla ad sanctuaria et propheta contra humum Israel.
EZEK|21|8|Et dices terrae Israel: Haec dicit Dominus Deus: Ecce ego ad te, et eiciam gladium meum de vagina sua et occidam in te iustum et impium.
EZEK|21|9|Pro eo autem quod occidi in te iustum et impium, idcirco egredietur gladius meus de vagina sua ad omnem carnem, ab austro ad aquilonem,
EZEK|21|10|ut sciat omnis caro quia ego Dominus eduxi gladium meum de vagina sua irrevocabilem.
EZEK|21|11|Et tu, fili hominis, ingemisce in contritione lumborum et in amaritudinibus ingemisce coram eis.
EZEK|21|12|Cumque dixerint ad te: "Quare tu gemis?", dices: Pro auditu quia venit et tabescet omne cor, et dissolventur universae manus, et infirmabitur omnis spiritus, et per cuncta genua fluent aquae; ecce venit et fiet ", ait Dominus Deus.
EZEK|21|13|Et factus est sermo Domini ad me dicens:
EZEK|21|14|" Fili hominis, propheta et dices: Haec dicit Dominus Deus: Loquere:Gladius, gladius exacutus estet etiam limatus;
EZEK|21|15|ut caedat victimas exacutus est,ut splendeat limatus est.
EZEK|21|16|Et datus est ad levigandum,ut teneatur manu.Iste exacutus est gladius et iste limatus,ut sit in manu interficientis.
EZEK|21|17|Clama et ulula, fili hominis,quia hic directus est in populum meum,hic in cunctos duces Israel,qui gladio traditi sunt cum populo meo.
EZEK|21|18|Idcirco plaude super femur,quia probatio est,dicit Dominus Deus.
EZEK|21|19|Tu ergo, fili hominis,propheta et percute manu ad manum.Et duplicetur gladius,ac triplicetur gladius interfectorum: hic est gladius occisionis magnae,qui eos circumdat,
EZEK|21|20|ut cor tabescat,et multiplicentur corruentes.In omnibus portis eorumdedi occisionem gladii:eheu, facti acuti et limati ad fulgendum,politi ad caedem!
EZEK|21|21|"Exacuere, vade ad dexteram sive ad sinistram,quocumque acies tuae sunt destinatae".
EZEK|21|22|Quin et ego plaudam manu ad manumet saturabo indignationem meam,ego Dominus locutus sum ".
EZEK|21|23|Et factus est sermo Domini ad me dicens:
EZEK|21|24|"Et tu, fili hominis, pone tibi duas vias, ut veniat gladius regis Babylonis: de terra una egrediantur ambae; et indicem statue, in capite viae civitatis statue.
EZEK|21|25|Viam pones, quo veniat gladius, ad Rabba filiorum Ammon et ad Iudam in Ierusalem munitissimam.
EZEK|21|26|Stat enim rex Babylonis in bivio in capite duarum viarum, divinationem quaerens, commiscens sagittas; interrogat teraphim, iecur consulit.
EZEK|21|27|Ad dexteram eius facta est divinatio super Ierusalem, ut ponat arietes, ut aperiat os ad caedem, ut elevet vocem in ululatu, ut ponat arietes contra portas, ut comportet aggerem, ut aedificet munitiones.
EZEK|21|28|Eritque quasi consulens frustra oraculum in oculis eorum, et iuramenta sanctissima sunt eis; ipse autem in memoriam revocabit iniquitatem ad capiendum.
EZEK|21|29|Idcirco haec dicit Dominus Deus: Pro eo quod in memoriam revocastis iniquitatem vestram, et revelatae sunt praevaricationes vestrae, et apparuerunt peccata vestra in omnibus operibus vestris; pro eo, inquam, quod in memoriam revocati estis, manu capiemini.
EZEK|21|30|Tu autem, profane, impie dux Israel, cuius venit dies in tempore iniquitatis finitae -
EZEK|21|31|haec dicit Dominus Deus - auferatur cidaris, tollatur corona; hoc non erit amplius. Humile sublevetur, et sublime humilietur.
EZEK|21|32|Ruinam, ruinam, ruinam ponam illud; et hoc non fiet, donec veniat, cuius est iudicium, et tradam ei.
EZEK|21|33|Et tu, fili hominis, propheta et dic: Haec dicit Dominus Deus ad filios Ammon et ad opprobrium eorum; et dices: Gladius, gladius est evaginatus ad occidendum, limatus ad consumendum, ut fulgeat,
EZEK|21|34|cum tibi videntur vana, et divinantur mendacia, ut ponatur gladius ad colla profanorum impiorum, quorum venit dies in tempore iniquitatis finitae.
EZEK|21|35|Revertatur ad vaginam suam. In loco, in quo creatus es, in terra nativitatis tuae iudicabo te.
EZEK|21|36|Et effundam super te indignationem meam, in igne furoris mei sufflabo in te; daboque te in manus hominum insipientium et fabricantium interitum.
EZEK|21|37|Igni eris cibus, sanguis tuus erit in medio terrae; oblivioni traderis, quia ego Dominus locutus sum ".
EZEK|22|1|Et factum est verbum Do mini ad me dicens:
EZEK|22|2|" Et tu, fili hominis, num iudicas, num iudicas civitatem sanguinum?
EZEK|22|3|Et ostendes ei omnes abominationes suas et dices: Haec dicit Dominus Deus: Civitas effundens sanguinem in medio sui, ut veniat tempus eius et, quae fecit idola contra semetipsam, ut pollueretur.
EZEK|22|4|In sanguine tuo, qui a te effusus est, deliquisti; et in idolis tuis, quae fecisti, polluta es; et appropinquare fecisti dies tuos et adduxisti tempus annorum tuorum. Propterea dedi te opprobrium gentibus et irrisionem universis terris.
EZEK|22|5|Quae iuxta sunt et quae procul a te, triumphabunt de te, sordibus famosa, grandis tumultu.
EZEK|22|6|Ecce principes Israel singuli pro brachio suo fuerunt in te ad effundendum sanguinem.
EZEK|22|7|Pater et mater contempti sunt in te, advena oppressus est in medio tui, pupillum et viduam afflixerunt apud te.
EZEK|22|8|Sanctuaria mea sprevisti et sabbata mea profanasti.
EZEK|22|9|Viri detractores fuerunt in te ad effundendum sanguinem et super montes comederunt in te; scelus operati sunt in medio tui.
EZEK|22|10|Verecundiora patris discooperuerunt in te, immunditiam menstruatae humiliaverunt in te;
EZEK|22|11|et unus in uxorem proximi sui operatus est abominationem, et alter nurum suam polluit nefarie; frater sororem suam, filiam patris sui, oppressit in te.
EZEK|22|12|Munera acceperunt apud te ad effundendum sanguinem, usuram et fenus accepisti et avare proximos tuos calumniabaris meique oblita es, ait Dominus Deus.
EZEK|22|13|Ecce complosi manus meas super lucrum tuum, quod fecisti, et super sanguinem, qui effusus est in medio tui.
EZEK|22|14|Numquid sustinebit cor tuum, aut praevalebunt manus tuae in diebus, quos ego faciam tibi? Ego Dominus locutus sum et faciam;
EZEK|22|15|et dispergam te in nationes et ventilabo te in terras et deficere faciam immunditiam tuam a te:
EZEK|22|16|et profanabo me in te in conspectu gentium, et scies quia ego Dominus.
EZEK|22|17|Et factum est verbum Domini ad me dicens:
EZEK|22|18|" Fili hominis, versa est mihi domus Israel in scoriam; omnes isti argentum et aes et stannum et ferrum et plumbum in medio fornacis, scoria facti sunt.
EZEK|22|19|Propterea haec dicit Dominus Deus: Eo quod versi estis omnes in scoriam, propterea ecce ego congregabo vos in medio Ierusalem
EZEK|22|20|congregatione argenti et aeris et ferri et plumbi et stanni in medio fornacis, ut succendatur in ea ignis ad conflandum: sic congregabo in furore meo et in ira mea et ponam et conflabo vos
EZEK|22|21|et congregabo vos et succendam vos in igne furoris mei, et conflabimini in medio eius.
EZEK|22|22|Ut conflatur argentum in medio fornacis, sic conflabimini in medio eius; et scietis quia ego Dominus effuderim indignationem meam super vos.
EZEK|22|23|Et factum est verbum Domini ad me dicens:
EZEK|22|24|" Fili hominis, dic ei: Tu es terra, super quam non cecidit pluvia neque imber in die furoris,
EZEK|22|25|cuius duces in medio eius sicut leo rugiens capiensque praedam: animas devoraverunt, opes et pretium acceperunt, viduas eius multiplicaverunt in medio illius.
EZEK|22|26|Sacerdotes eius contempserunt legem meam et polluerunt sanctuaria mea, inter sanctum et profanum non habuerunt distantiam et inter pollutum et mundum non docuerunt distinguere et a sabbatis meis averterunt oculos suos, et coinquinabar in medio eorum.
EZEK|22|27|Principes eius in medio illius quasi lupi rapientes praedam ad effundendum sanguinem et perdendas animas et avare sectanda lucra.
EZEK|22|28|Prophetae autem eius liniebant eis omnia calce, videntes vana et divinantes eis mendacium, dicentes: "Haec dicit Dominus Deus", cum Dominus non sit locutus.
EZEK|22|29|Populus terrae calumniabatur calumniam et rapiebat violenter; egenum et pauperem affligebant et advenam opprimebant absque iudicio.
EZEK|22|30|Et quaesivi de eis virum, qui interponeret saepem et staret in confractione contra me pro terra, ne dissiparem eam, et non inveni.
EZEK|22|31|Et effudi super eos indignationem meam, in igne irae meae consumpsi eos, viam eorum in caput eorum reddidi ", ait Dominus Deus.
EZEK|23|1|Et factus est sermo Domini ad me dicens:
EZEK|23|2|" Fili hominis, duae mulieres filiae matris unius fuerunt
EZEK|23|3|et fornicatae sunt in Aegypto, in adulescentia sua fornicatae sunt; ibi subacta sunt ubera earum, et tactae sunt mammae virginitatis earum.
EZEK|23|4|Nomina autem earum Oolla maior et Ooliba soror eius; et habui eas, et pepererunt filios et filias: porro earum nomina Samaria Oolla et Ierusalem Ooliba.
EZEK|23|5|Fornicata est igitur Oolla discedens a me; et insanivit in amatores suos, in Assyrios: bellatores
EZEK|23|6|vestitos hyacintho, principes et magistratus, iuvenes desiderabiles universi, equites ascensores equorum.
EZEK|23|7|Et dedit fornicationes suas ad eos electos filiorum Assyriae universos; et apud omnes, in quos insanivit, in omnibus idolis eorum polluta est.
EZEK|23|8|Insuper et fornicationes suas, quas habuerat in Aegypto, non reliquit; nam et illi dormierunt cum ea in adulescentia eius, et illi tetigerant ubera virginitatis eius et effuderant fornicationem suam super eam.
EZEK|23|9|Propterea tradidi eam in manus amatorum suorum, in manus filiorum Assyriae, in quos insanivit;
EZEK|23|10|ipsi discooperuerunt ignominiam eius, filios et filias illius tulerunt et ipsam occiderunt gladio; et facta est famosa mulieribus, et iudicia perpetrarunt in ea.
EZEK|23|11|Quod cum vidisset soror eius Ooliba, plus quam illa insanivit libidine et fornicatione sua super fornicationem sororis suae.
EZEK|23|12|In filios Assyriorum amore exarsit: duces et magistratus, bellatores indutos veste pretiosa, equites, qui vectabantur equis, adulescentes cuncti desiderabiles.
EZEK|23|13|Et vidi quod polluta esset: via una ambarum;
EZEK|23|14|et auxit fornicationes suas. Cumque vidisset viros depictos in pariete, imagines Chaldaeorum expressas sinopide,
EZEK|23|15|et accinctos balteis renes, et tiaras defluentes in capitibus eorum; aspectus essedariorum omnibus, similitudo filiorum Babylonis, quorum patria Chaldaea.
EZEK|23|16|Et insanivit super eos concupiscentia oculorum suorum et misit nuntios ad eos in Chaldaeam.
EZEK|23|17|Cumque venissent ad eam filii Babylonis ad cubile amoris, polluerunt eam stupris suis; et, cum polluta esset ab eis, recessit anima eius ab illis.
EZEK|23|18|Cum manifestasset fornicationes suas et discooperuisset ignominiam suam, recessit anima mea ab ea, sicut recesserat anima mea a sorore eius.
EZEK|23|19|Multiplicavit autem fornicationes suas, recordans dies adulescentiae suae, quibus fornicata est in terra Aegypti;
EZEK|23|20|et insanivit libidine in amatores suos, quorum membra sunt ut membra asinorum, et sicut fluxus equorum fluxus eorum.
EZEK|23|21|Et desiderasti scelus adulescentiae tuae, quando subacta sunt in Aegypto ubera tua, et tactae mammae pubertatis tuae.
EZEK|23|22|Propterea, Ooliba, haec dicit Dominus Deus: Ecce ego suscitabo amatores tuos contra te, de quibus recessit anima tua; et congregabo eos adversum te in circuitu,
EZEK|23|23|filios Babylonis et universos Chaldaeos, Phacud et Sue et Cue, omnes filios Assyriorum cum eis, iuvenes desiderabiles, duces et magistratus universos, essedarios et nominatos, ascensores equorum omnes.
EZEK|23|24|Et venient super te instructi curru et rota, cum multitudine populorum; scuto et clipeo et galea armabuntur contra te undique, et dabo coram eis iudicium, et iudicabunt te iudiciis suis.
EZEK|23|25|Et ponam zelum meum in te, quem exercent tecum in furore: nasum tuum et aures tuas praecident et, quae remanserint de te, gladio concident; ipsi filios tuos et filias tuas capient, et novissimum tuum devorabitur igni.
EZEK|23|26|Et denudabunt te vestimentis tuis et tollent vasa gloriae tuae;
EZEK|23|27|et cessare faciam scelus tuum de te et fornicationem tuam de terra Aegypti, nec levabis oculos tuos ad eos et Aegypti non recordaberis amplius.
EZEK|23|28|Quia haec dicit Dominus Deus: Ecce ego tradam te in manu eorum, quos odisti, in manu, de quibus recessit anima tua;
EZEK|23|29|et agent tecum in odio et tollent omnes labores tuos et dimittent te nudam et ignominia plenam, et revelabitur ignominia fornicationum tuarum, scelus tuum et fornicationes tuae.
EZEK|23|30|Fecerunt haec tibi, quia fornicata es post gentes, inter quas polluta es in idolis earum.
EZEK|23|31|In via sororis tuae ambulasti, et dabo calicem eius in manu tua.
EZEK|23|32|Haec dicit Dominus Deus:Calicem sororis tuae bibesprofundum et latumC eris in derisum et in subsannationem C:est capacissimus.
EZEK|23|33|Ebrietate et dolore repleberis,calice stuporis et horroris,calice sororis tuae Samariae,
EZEK|23|34|et bibes illum et epotabis usque ad faeces;et fragmenta eius rodeset ubera tua lacerabis,quia ego locutus sum ",ait Dominus Deus.
EZEK|23|35|Propterea haec dicit Dominus Deus: " Quia oblita es mei et proiecisti me post tergum tuum, tu quoque porta scelus tuum et fornicationes tuas ".
EZEK|23|36|Et ait Dominus ad me: " Fili hominis, numquid iudicas Oollam et Oolibam? Annuntia ergo eis scelera earum.
EZEK|23|37|Quia adulteratae sunt, et sanguis in manibus earum, et cum idolis suis fornicatae sunt; insuper et filios suos, quos genuerunt mihi, obtulerunt eis ad devorandum.
EZEK|23|38|Sed et hoc fecerunt mihi: polluerunt sanctuarium meum in die illa et sabbata mea profanaverunt.
EZEK|23|39|Cumque immolarent filios suos idolis suis et ingrederentur sanctuarium meum in die illa, ut polluerent illud, ecce haec fecerunt in medio domus meae.
EZEK|23|40|Quin et miserunt ad viros venientes de longe, ad quos nuntius missus erat; itaque ecce venerunt. Quibus te lavisti et circumlevisti stibio oculos tuos et ornata es mundo muliebri;
EZEK|23|41|sedisti in lecto pulcherrimo, et mensa ornata est ante te, thymiama meum et unguentum meum posuisti super eam.
EZEK|23|42|Et vox multitudinis exsultantis erat apud eam et apud viros multitudo hominum, qui adducebantur de deserto; et posuerunt armillas in manibus earum et coronas speciosas in capitibus earum.
EZEK|23|43|Et dixi de ea, quae attrita est in adulteriis: Nunc fornicabitur in fornicatione sua etiam haec.
EZEK|23|44|Et ingressi sunt ad eam quasi ad mulierem meretricem; sic ingrediebantur ad Oollam et ad Oolibam, mulieres nefarias.
EZEK|23|45|Viri ergo iusti sunt; hi iudicabunt eas iudicio adulterarum et iudicio effundentium sanguinem, quia adulterae sunt, et sanguis in manibus earum.
EZEK|23|46|Haec enim dicit Dominus Deus: " Adduc ad eas congregationem et trade eas in terrorem et in rapinam;
EZEK|23|47|et lapidentur lapidibus congregationis et confodiantur gladiis eorum; filios et filias earum interficiant et domos earum igne succendant.
EZEK|23|48|Et auferam scelus de terra, et discent omnes mulieres, ne faciant secundum scelus vestrum;
EZEK|23|49|et dabunt scelus vestrum super vos, et peccata idolorum vestrorum portabitis et scietis quia ego Dominus Deus ".
EZEK|24|1|Et factum est verbum Do mini ad me in anno nono, in mense decimo, decima mensis, dicens:
EZEK|24|2|"Fili hominis, scribe tibi nomen diei huius, in qua aggressus est rex Babylonis adversum Ierusalem hodie.
EZEK|24|3|Et dices per proverbium ad domum irritatricem parabolam et loqueris ad eos: Haec dicit Dominus Deus:Pone ollam; pone, inquam,et mitte in ea aquam.
EZEK|24|4|Congere frusta eius in ea,omnem partem bonam, femur et armum,electis ossibus imple eam,
EZEK|24|5|pinguissimum pecus assume.Compone quoque struem lignorum sub ea;effervescant frusta eius,et coque ossa illius in medio eius.
EZEK|24|6|Propterea haec dicit Dominus Deus:Vae civitati sanguinum,ollae, cuius rubigo in ea est,et rubigo eius non exivit de ea!Per partes et per partes suas eice ex ea,neque cadat super eam sors.
EZEK|24|7|Sanguis enim eius in medio eius est,super limpidissimam petram effudit illum;non effudit illum super terram,ut possit operiri pulvere;
EZEK|24|8|ut superducerem indignationem meamet vindicta ulciscerer,dedi sanguinem eiussuper petram limpidissimam, ne operiretur.
EZEK|24|9|Propterea haec dicit Dominus Deus:Vae civitati sanguinum,cuius ego grandem faciam pyram!
EZEK|24|10|Congere ligna, succende ignem,coque carnes usque ad consumptionemet effunde ius,et ossa comburentur.
EZEK|24|11|Relinque quoque eam super prunas vacuam,ut incalescat, et ardescat aes eius,et confletur in medio eius inquinamentum eius,et consumatur rubigo eius.
EZEK|24|12|Multo labore sudatum est,et non exibit de ea nimia rubigo eius,neque per ignem.
EZEK|24|13|Immunditia tua execrabilis, quia mundare te volui, et non es mundata a sordibus tuis; sed nec mundaberis prius, donec quiescere faciam indignationem meam in te.
EZEK|24|14|Ego Dominus locutus sum; veniet et faciam: non indulgebo nec parcam nec placabor. Iuxta vias tuas et iuxta opera tua iudicabo te ", dicit Dominus.
EZEK|24|15|Et factum est verbum Domini ad me dicens:
EZEK|24|16|" Fili hominis, ecce ego tollo a te delicias oculorum tuorum in plaga, et non planges neque plorabis, neque fluent lacrimae tuae.
EZEK|24|17|Ingemisce tacens, mortuorum luctum non facies, corona tua circumligata sit tibi, et calceamenta tua pones in pedibus tuis nec amictu ora velabis nec cibos lugentium comedes ".
EZEK|24|18|Locutus sum ergo ad populum mane, et mortua est uxor mea vespere; fecique mane, sicut praeceperat mihi.
EZEK|24|19|Et dixit ad me populus: " Quare non indicas nobis, quid ista significent, quae tu facis? ".
EZEK|24|20|Et dixi ad eos: " Sermo Domini factus est ad me dicens:
EZEK|24|21|Loquere domui Israel: Haec dicit Dominus Deus: Ecce ego polluam sanctuarium meum, superbiam roboris vestri et delicias oculorum vestrorum et sollicitudinem animae vestrae. Filii vestri et filiae, quas reliquistis, gladio cadent.
EZEK|24|22|Et facietis, sicut feci: ora amictu non velabitis et cibos lugentium non comedetis,
EZEK|24|23|coronas habebitis in capitibus vestris et calceamenta in pedibus, non plangetis neque flebitis, sed tabescetis in iniquitatibus vestris, et unusquisque gemet ad fratrem suum.
EZEK|24|24|Eritque Ezechiel vobis in portentum: iuxta omnia, quae fecit, facietis, cum venerit istud, et scietis quia ego Dominus Deus.
EZEK|24|25|Et tu, fili hominis, ecce in die, quo tollam ab eis fortitudinem eorum et gaudium magnificentiae et delicias oculorum eorum et desiderium animae eorum, filios et filias eorum;
EZEK|24|26|in die illa, cum venerit fugiens ad te, ut annuntiet tibi,
EZEK|24|27|in die, inquam, illa aperietur os tuum cum eo, qui fugit; et loqueris et non silebis ultra erisque eis in portentum, et scient quia ego Dominus.
EZEK|25|1|Et factus est sermo Domini ad me dicens:
EZEK|25|2|" Fili hominis, pone faciem tuam contra filios Ammon et propheta de eis
EZEK|25|3|et dices filiis Ammon: Audite verbum Domini Dei.Haec dicit Dominus Deus: Pro eo quod dixisti: "Euge!" super sanctuarium meum, quia pollutum est, et super terram Israel, quoniam desolata est, et super domum Iudae, quoniam ducti sunt in captivitatem,
EZEK|25|4|idcirco ego tradam te filiis orientalibus in hereditatem, et collocabunt castra sua in te et ponent in te tentoria sua; ipsi comedent fruges tuas, et ipsi bibent lac tuum.
EZEK|25|5|Daboque Rabba in pascua camelorum et filios Ammon in cubile pecorum, et scietis quia ego Dominus.
EZEK|25|6|Quia haec dicit Dominus Deus: Pro eo quod plausisti manu et percussisti pede et gavisa es ex toto affectu super terram Israel,
EZEK|25|7|idcirco ecce ego extendam manum meam super te et tradam te in direptionem gentium et interficiam te de populis et perdam de terris et conteram, et scies quia ego Dominus.
EZEK|25|8|Haec dicit Dominus Deus: Pro eo quod dixerunt Moab et Seir: "Ecce sicut omnes gentes domus Iudae!",
EZEK|25|9|idcirco ecce ego aperiam latus Moab privans eam civitatibus, civitatibus, inquam, eius, a finibus eius, decore terrae: Bethiesimoth et Baalmeon et Cariathaim;
EZEK|25|10|filiis orientis cum filiis Ammon dabo eam in hereditatem, ut non sit memoria ultra filiorum Ammon in gentibus.
EZEK|25|11|Et in Moab faciam iudicia, et scient quia ego Dominus.
EZEK|25|12|Haec dicit Dominus Deus: Pro eo quod fecit Idumaea ultionem, ut se vindicaret de domo Iudae, peccavitque delinquens et vindictam expetivit de eis,
EZEK|25|13|idcirco haec dicit Dominus Deus: Extendam manum meam super Idumaeam et auferam de ea hominem et iumentum et faciam eam desertum; de Theman et usque Dedan gladio cadent.
EZEK|25|14|Et dabo ultionem meam super Idumaeam per manum populi mei Israel, et facient in Edom iuxta iram meam et furorem meum, et scient vindictam meam, dicit Dominus Deus.
EZEK|25|15|Haec dicit Dominus Deus: Pro eo quod fecerunt Palaestini in vindicta et ulti se sunt toto animo interficientes et implentes inimicitias sempiternas,
EZEK|25|16|propterea haec dicit Dominus Deus: Ecce ego extendam manum meam super Palaestinos et interficiam Cherethaeos et perdam reliquias maritimae regionis;
EZEK|25|17|faciamque in eis ultiones magnas, arguens in furore, et scient quia ego Dominus, cum dedero vindictam meam super eos ".
EZEK|26|1|Et factum est in undecimo anno, prima mensis, factus est sermo Domini ad me dicens:
EZEK|26|2|"Fili hominis, pro eo quod dixit Tyrus de Ierusalem:Euge, confracta estporta populorum!Conversa est ad me;quae erat plena, deserta est",
EZEK|26|3|propterea haec dicit Dominus Deus:Ecce ego super te, Tyre,et ascendere faciam ad te gentes multas,sicut ascendit mare fluctuans;
EZEK|26|4|et dissipabunt muros Tyriet destruent turres eius,et radam pulverem eius de ea,et dabo eam in limpidissimam petram.
EZEK|26|5|Siccatio sagenarumerit in medio maris,quia ego locutus sum,ait Dominus Deus;et erit in direptionem gentibus.
EZEK|26|6|Filiae quoque eius, quae sunt in agro,gladio interficientur,et scient quia ego Dominus.
EZEK|26|7|Quia haec dicit Dominus Deus:Ecce ego adducam ad TyrumNabuchodonosor, regem Babylonis,ab aquilone, regem regum,cum equis et curribus et equitibuset coetu populoque magno.
EZEK|26|8|Filias tuas, quae sunt in agro,gladio interficiet,et circumdabit te munitionibuset comportabit aggerem in gyroet levabit contra te clipeum
EZEK|26|9|et vineas et arietes temperabit in muros tuoset turres tuas destruet in armatura sua.
EZEK|26|10|Inundatione equorum eiusoperiet te pulvis eorum,a sonitu equitumet rotarum et curruummovebuntur muri tui,dum ingressus fuerit portas tuasquasi per introitus urbis dissipatae.
EZEK|26|11|Ungulis equorum suorumconculcabit omnes plateas tuas,populum tuum gladio caedet,et columnae tuae fortissimaein terram corruent.
EZEK|26|12|Vastabunt opes tuas,diripient negotiationes tuaset destruent muros tuoset domos tuas praeclaras subvertentet lapides tuos et ligna tua et pulverem tuumin medio aquarum ponent.
EZEK|26|13|Et quiescere faciam tumultum canticorum tuorum,et sonitus cithararum tuarum non audietur amplius,
EZEK|26|14|et dabo te in limpidissimam petram;siccatio sagenarum eris,nec aedificaberis ultra,quia ego locutus sum,dicit Dominus Deus.
EZEK|26|15|Haec dicit Dominus Deus Tyro: Numquid non a sonitu ruinae tuae et gemitu interfectorum tuorum, cum occisi fuerint in medio tui, commovebuntur insulae?
EZEK|26|16|Et descendent de sedibus suis omnes principes maris et auferent pallia sua et vestimenta sua varia abicient; et induentur stupore, in terra sedebunt et attoniti et tremefacti stupebunt super te.
EZEK|26|17|Et assumentes super te lamentum dicent tibi:Quomodo peristi, quae habitas in mari,urbs inclita,quae fuisti fortis in maricum habitatoribus tuis,quos formidabant universi!
EZEK|26|18|Nunc stupebunt navesin die ruinae tuae,et turbabuntur insulae in mariob exitum tuum".
EZEK|26|19|Quia haec dicit Dominus Deus: Cum dedero te urbem desolatam sicut civitates, quae non habitantur, et adduxero super te abyssum, et operuerint te aquae multae,
EZEK|26|20|detraham te cum his, qui descendunt in lacum, ad populum pristinum et collocabo te in profundis terrae sicut ruinas a saeculo cum his, qui descendunt in lacum, ut non habiteris et consistas in terra viventium;
EZEK|26|21|in nihilum redigam te, et non eris et requisita non invenieris ultra in sempiternum ", dicit Dominus Deus.
EZEK|27|1|Et factum est verbum Do mini ad me dicens:
EZEK|27|2|"Tu er go, fili hominis, assume super Tyrum lamentum
EZEK|27|3|et dices Tyro, quae habitat in introitu maris, negotiatrici populorum ad insulas multas: Haec dicit Dominus Deus:O Tyre, tu dixisti: "Perfecti decoris ego sum!".
EZEK|27|4|In corde maris fines tui;qui te aedificaverunt, impleverunt decorem tuum.
EZEK|27|5|Abietibus de Sanir exstruxerunttibi omnia tabulata;cedrum de libano tulerunt,ut facerent tibi malum;
EZEK|27|6|quercus de Basandolaverunt in remos tuoset transtra tua fecerunt ex eboreet cupressis de insulis Cetthim.
EZEK|27|7|Byssus varia texta de Aegyptoerat tibi in velum,ut poneretur in malo,hyacinthus et purpura de insulis Elisafacta sunt operimentum tuum.
EZEK|27|8|Habitatores Sidonis et Aradiifuerunt remiges tui;sapientes tui, Tyre,facti sunt nautae tui.
EZEK|27|9|Senes Gibli et prudentes eius fuerunt in te,ut sarcirent rimas tuas.Omnes naves maris et nautae earumfuerunt in te, ut mercarentur merces tuas.
EZEK|27|10|Persae et Lud et Phuterant in exercitu tuo,viri bellatores tui.Clipeum et galeam suspenderunt in te;ipsi dederunt tibi splendorem.
EZEK|27|11|Filii Aradii cum exercitu tuo erant super muros tuos in circuitu, et Gammadii erant in turribus tuis. Clipeos suos suspenderunt in muris tuis per gyrum; ipsi compleverunt pulchritudinem tuam.
EZEK|27|12|Tharsis negotiatrix tua propter multitudinem cunctarum divitiarum; argentum, ferrum, stannum plumbumque dederunt pro mercibus tuis.
EZEK|27|13|Iavan, Thubal et Mosoch ipsi institores tui; mancipia et vasa aerea adduxerunt tibi in commutationem populo tuo.
EZEK|27|14|De domo Thogorma equos et equites et mulos adduxerunt pro mercibus tuis ad forum tuum;
EZEK|27|15|filii Rhodi negotiatores tui; insulae multae negotiatio manus tuae: dentes eburneos et ebenina reddiderunt tibi ut tributum.
EZEK|27|16|Edom negotiator tuus propter multitudinem operum tuorum; carbunculum, purpuram et scutulata et byssum et corallia et rubinum attulerunt pro mercibus tuis.
EZEK|27|17|Iuda et terra Israel ipsi institores tui; frumentum primum, balsamum et mel et oleum et resinam attulerunt tibi in commutationem.
EZEK|27|18|Damascenus negotiator tuus propter multitudinem operum tuorum, propter multitudinem diversarum opum; vinum de Helbon et lanam de Sahar
EZEK|27|19|et vinum de Uzal pro mercibus tuis dederunt; ferrum fabrefactum, cassia et calamus in commutatione tua erat.
EZEK|27|20|Dedan institores tui in tapetibus ad equitandum.
EZEK|27|21|Arabia et universi principes Cedar ipsi negotiatores manus tuae; cum agnis et arietibus et haedis, cum quibus erant negotiatores tui.
EZEK|27|22|Venditores Saba et Regma, ipsi negotiatores tui, universa prima aromata et omnem lapidem pretiosum et aurum dederunt pro mercibus tuis.
EZEK|27|23|Charran et Chenne et Eden negotiatores tui; Saba, Assyria et Chelmad venditores tui.
EZEK|27|24|Ipsi negotiatores tui cum vestibus splendidis, involucris hyacinthinis et polymitis texturisque discoloribus, funibus obvolutis et cedris in negotiationibus tuis.
EZEK|27|25|Naves Tharsis, principes tuiin negotiatione tua;et repleta es et glorificata nimisin corde maris.
EZEK|27|26|In aquis multis adduxerunt teremiges tui;ventus auster contrivit tein corde maris.
EZEK|27|27|Divitiae tuae et thesauri tui et multiplices merces tuae,nautae tui et gubernatores tui,resarcientes rimas tuas et commutantes merces tuas,omnes quoque viri bellatores tui,qui sunt in te,cum universa multitudine tua,quae est in medio tui,cadent in corde marisin die ruinae tuae.
EZEK|27|28|A sonitu clamoris gubernatorum tuorumconturbabuntur litora.
EZEK|27|29|Et descendent de navibus suisomnes, qui tenebant remum;nautae et universi gubernatores marisin terra stabunt.
EZEK|27|30|Et eiulabunt super te voce magnaet clamabunt amare;et superiacient pulverem capitibus suis,in cinere volutabuntur.
EZEK|27|31|Et radent super te calvitiumet accingentur ciliciiset plorabunt te in amaritudine animaeploratu amarissimo;
EZEK|27|32|et assument super te congementes carmen lugubreet plangent te:Quae est ut Tyrus, quae obmutuitin medio maris?
EZEK|27|33|Cum venissent merces tuae de mari, satiasti populos multos;in multitudine divitiarum tuarum et mercium tuarumditasti reges terrae.
EZEK|27|34|Nunc contrita es a mariin profundis aquarum.Opes tuae et omnis multitudo tua,quae erat in medio tui,ceciderunt.
EZEK|27|35|Universi habitatores insularumobstupuerunt super te,et reges earum horrore formidarunt vultu conturbato;
EZEK|27|36|negotiatores in populis sibilaverunt super te.In horrorem facta eset non eris usque in perpetuum" ".
EZEK|28|1|Et factus est sermo Domini ad me dicens:
EZEK|28|2|" Fili hominis, dic principi Tyri: Haec dicit Dominus Deus:Eo quod elevatum est cor tuum,et dixisti: "Deus ego sumet in cathedra deorum sedeoin corde maris!",cum sis homo et non Deus,et dedisti cor tuum quasi cor Dei.
EZEK|28|3|Ecce sapientior es tu Danel,omne secretum non est absconditum a te,
EZEK|28|4|in sapientia et prudentia tuafecisti tibi opeset acquisisti aurum et argentumin thesauris tuis;
EZEK|28|5|in multitudine sapientiae tuae et in negotiatione tuamultiplicasti tibi opes,et elevatum est cor tuum in opibus tuis.
EZEK|28|6|Propterea haec dicit Dominus Deus: Eo quod fecisti cor tuum quasi cor Dei,
EZEK|28|7|idcirco ecce ego adducam super tealienos violentissimos gentium;et nudabunt gladios suos super pulchritudinem sapientiae tuaeet polluent splendorem tuum.
EZEK|28|8|In fossam detrahent te, et morierisinteritu occisorum in corde maris.
EZEK|28|9|Numquid dicens loqueris: "Deus ego sum!"coram interficientibus te,cum sis homo et non Deusin manu occidentium te?
EZEK|28|10|Morte incircumcisorum morierisin manu alienorum,quia ego locutus sum ",ait Dominus Deus.
EZEK|28|11|Et factus est sermo Domini ad me dicens: " Fili hominis, leva planctum super regem Tyri
EZEK|28|12|et dices ei: Haec dicit Dominus Deus:Tu signaculum perfectum,plenus sapientia et perfectus decore;
EZEK|28|13|in deliciis paradisi Dei fuisti,omnis lapis pretiosus operimentum tuum:sardius, topazius et iaspis,chrysolithus et onyx et beryllus,sapphirus et carbunculus et smaragdus,aurum opus caelaturae in te;in die, qua conditus es, praeparata sunt.
EZEK|28|14|Cum cherub extento et protegente te posui te,in monte sancto Dei fuisti,in medio lapidum ignitorum ambulasti,
EZEK|28|15|perfectus in viis tuisa die conditionis tuae,donec inventa est iniquitas in te.
EZEK|28|16|In multitudine negotiationis tuae repleta sunt interiora tuainiquitate, et peccasti.Et eieci te de monte Dei,et perdidit te cherub protegensde medio lapidum ignitorum.
EZEK|28|17|Elevatum est cor tuum in decore tuo;perdidisti sapientiam tuam propter splendorem tuum:in terram proieci te,ante faciem regum dedi te, ut cernerent te.
EZEK|28|18|In multitudine iniquitatum tuarumet iniquitate negotiationis tuaepolluisti sanctuaria tua;producam ergo ignem de medio tui,qui comedat te,et dabo te in cinerem super terramin conspectu omnium videntium te.
EZEK|28|19|Omnes, qui viderint te, in gentibusobstupescent super te;in horrorem factus eset non eris in perpetuum ".
EZEK|28|20|Et factus est sermo Domini ad me dicens:
EZEK|28|21|" Fili hominis, pone faciem tuam contra Sidonem et propheta de ea
EZEK|28|22|et dices: Haec dicit Dominus Deus:Ecce ego ad te, Sidon,et glorificabor in medio tui,et scient quia ego Dominus,cum fecero in ea iudiciaet sanctificatus fuero in ea.
EZEK|28|23|Et immittam ei pestilentiamet sanguinem in plateis eius,et corruent interfecti in medio eius gladio per circuitum,et scient quia ego Dominus.
EZEK|28|24|Et non erit ultra domui Israel stimulus amaritudinis et spina dolorem inferens undique per circuitum eorum, qui adversantur eis, et scient quia ego Dominus Deus.
EZEK|28|25|Haec dicit Dominus Deus: Quando congregavero domum Israel de populis, in quibus dispersi sunt, sanctificabor in eis coram gentibus, et habitabunt in terra sua, quam dedi servo meo Iacob;
EZEK|28|26|et habitabunt in ea securi et aedificabunt domos plantabuntque vineas et habitabunt confidenter, cum fecero iudicia in omnibus, qui adversantur eis per circuitum, et scient quia ego Dominus Deus eorum ".
EZEK|29|1|In anno decimo, in decimo mense, duodecima mensis, factum est verbum Domini ad me dicens:
EZEK|29|2|" Fili hominis, pone faciem tuam contra pharaonem, regem Aegypti, et prophetabis de eo et de Aegypto universa.
EZEK|29|3|Loquere et dices: Haec dicit Dominus Deus:Ecce ego ad te, pharao,rex Aegypti,draco magne, qui cubasin medio fluminum tuorumet dicis: "Meus est fluvius,et ego feci memetipsum!".
EZEK|29|4|Et ponam uncos in maxillis tuiset agglutinabo pisces fluminum tuorum squamis tuiset extraham te de medio fluminum tuorum,et universi pisces tui squamis tuis adhaerebunt.
EZEK|29|5|Et proiciam te in desertumet omnes pisces fluminum tuorum.Super faciem terrae cades;non colligeris neque congregaberis.Bestiis terrae et volatilibus caelidedi te ad devorandum.
EZEK|29|6|Et scient omnes habitatores Aegyptiquia ego Dominus,pro eo quod fuisti baculus arundineusdomui Israel:
EZEK|29|7|quando apprehenderunt te manu,confractus es et lacerasti omnem umerum eorumet, innitentibus eis super te,comminutus eset dissolvisti omnes lumbos eorum.
EZEK|29|8|Propterea haec dicit Dominus Deus: Ecce ego adducam super te gladium et interficiam de te hominem et iumentum;
EZEK|29|9|et erit terra Aegypti in desertum et solitudinem, et scient quia ego Dominus. Pro eo quod dixeris: "Fluvius meus est, et ego feci!",
EZEK|29|10|idcirco ecce ego ad te et ad flumina tua, daboque terram Aegypti in solitudines, gladio dissipatam a Magdolo ad Syenen et usque ad terminos Chus.
EZEK|29|11|Non pertransibit eam pes hominis, neque pes iumenti gradietur in ea, et non habitabitur quadraginta annis;
EZEK|29|12|daboque terram Aegypti desertam in medio terrarum desertarum, et civitates eius in medio urbium subversarum erunt desolatae quadraginta annis, et dispergam Aegyptios in nationes et ventilabo eos in terras.
EZEK|29|13|Quia haec dicit Dominus Deus: Post finem quadraginta annorum congregabo Aegyptios de populis, in quibus dispersi fuerunt,
EZEK|29|14|et convertam sortem Aegypti et collocabo eos in terra Phatures, in terra nativitatis suae; et erunt ibi in regnum humile.
EZEK|29|15|Inter regna cetera erit humillima et non elevabitur ultra super nationes, et imminuam eos, ne imperent gentibus.
EZEK|29|16|Neque erunt ultra domui Israel in confidentiam, in memoriam revocans iniquitatem, cum sequerentur eos, et scient quia ego Dominus Deus ".
EZEK|29|17|Et factum est in vicesimo et septimo anno, in primo, in una mensis, factum est verbum Domini ad me dicens:
EZEK|29|18|" Fili hominis, Nabuchodonosor, rex Babylonis, servire fecit exercitum suum servitute magna adversus Tyrum; omne caput decalvatum et omnis umerus attritus est, et merces non est reddita ei neque exercitui eius de Tyro pro servitute, qua servivit adversum eam.
EZEK|29|19|Propterea haec dicit Dominus Deus: Ecce ego dabo Nabuchodonosor, regi Babylonis, terram Aegypti, et accipiet opes eius et depraedabitur manubias eius et diripiet spolia eius, et erit merces exercitui illius,
EZEK|29|20|ut stipendium eius, pro quo servivit adversum eam. Dedi ei terram Aegypti pro eo quod laboraverunt mihi, ait Dominus Deus.
EZEK|29|21|In die illo germinare faciam cornu domui Israel, et tibi dabo apertum os in medio eorum, et scient quoniam ego Dominus ".
EZEK|30|1|Et factum est verbum Do mini ad me dicens:
EZEK|30|2|" Fili ho minis, propheta et dic: Haec dicit Dominus Deus:Ululate, vae diei,
EZEK|30|3|quia iuxta est dies,et appropinquat dies Domini,dies nubis; tempus gentium erit.
EZEK|30|4|Et veniet gladius in Aegyptum,et erit pavor in Chus,cum ceciderint vulnerati in Aegypto,et ablatae fuerint opes illius,et destructa fundamenta eius.
EZEK|30|5|Chus et Phut et Lud et omne vulgus promiscuumet Chub et filii terrae foederiscum eis gladio cadent.
EZEK|30|6|Haec dicit Dominus Deus:Et corruent fulcientes Aegyptum,et destruetur superbia potentiae eius;a Magdolo usque ad Syenen gladio cadent in ea,ait Dominus Deus.
EZEK|30|7|Et dissipabuntur in medio terrarum desolatarum, et urbes eius in medio civitatum desertarum erunt;
EZEK|30|8|et scient quia ego Dominus, cum dedero ignem in Aegyptum, et attriti fuerint omnes auxiliatores eius.
EZEK|30|9|In die illa egredientur nuntii a facie mea in navibus ad conterendam confidentiam Chus, et erit pavor in eis in die Aegypti, quia veniet.
EZEK|30|10|Haec dicit Dominus Deus: Cessare faciam pompam Aegypti in manu Nabuchodonosor, regis Babylonis.
EZEK|30|11|Ipse et populus eius cum eo violentissimi gentium adducentur ad disperdendam terram; et evaginabunt gladios suos super Aegyptum et implebunt terram interfectis.
EZEK|30|12|Et faciam alveos fluminum aridos et tradam terram in manu pessimorum et dissipabo terram et plenitudinem eius in manu alienorum. Ego Dominus locutus sum.
EZEK|30|13|Haec dicit Dominus Deus:Et disperdam simulacraet cessare faciam idola de Memphi,et dux de terra Aegyptinon erit amplius,et dabo terrorem in terra Aegypti.
EZEK|30|14|Et disperdam terram Phatureset dabo ignem in Taniet faciam iudicia in No.
EZEK|30|15|Et effundam indignationem meam super Sin, robur Aegypti, et interficiam multitudinem No.
EZEK|30|16|Et dabo ignem in Aegypto; quasi parturiens dolebit Sin, et in No scissura erit, et contra Memphin hostes plena die.
EZEK|30|17|Iuvenes Heliopoleos et Bubasti gladio cadent, et ipsae captivae ducentur.
EZEK|30|18|Et in Taphnis nigrescet dies, cum contrivero ibi sceptra Aegypti, et defecerit in ea superbia potentiae eius; ipsam nubes operiet, filiae autem eius in captivitatem ducentur.
EZEK|30|19|Et faciam iudicia in Aegypto, et scient quia ego Dominus ".
EZEK|30|20|Et factum est in undecimo anno, in primo, in septima mensis, factum est verbum Domini ad me dicens:
EZEK|30|21|" Fili hominis, brachium pharaonis, regis Aegypti, confregi, et ecce non est obvolutum, ut restitueretur ei sanitas, ut ligaretur pannis et farciretur linteolis, ut recepto robore posset tenere gladium.
EZEK|30|22|Propterea haec dicit Dominus Deus: Ecce ego ad pharaonem, regem Aegypti, et comminuam brachium eius forte sed confractum et deiciam gladium de manu eius
EZEK|30|23|et dispergam Aegyptum in gentibus et ventilabo eos in terris.
EZEK|30|24|Et confortabo brachia regis Babylonis daboque gladium meum in manu eius; et confringam brachia pharaonis, et gemet gemitibus sicut transfixus coram facie eius.
EZEK|30|25|Et confortabo brachia regis Babylonis, et brachia pharaonis concident; et scient quia ego Dominus, cum dedero gladium meum in manu regis Babylonis, et extenderit eum super terram Aegypti.
EZEK|30|26|Et dispergam Aegyptum in nationes et ventilabo eos in terras, et scient quia ego Dominus ".
EZEK|31|1|Et factum est in anno unde cimo, in tertio, una mensis, factum est verbum Domini ad me dicens:
EZEK|31|2|" Fili hominis, dic pharaoni, regi Aegypti, et pompae eius:Cui similis factus es in magnitudine tua?
EZEK|31|3|Ecce abies, quasi cedrus in Libano,pulcher ramis et frondibus nemorosusexcelsusque altitudine,et inter nubes elevatum est cacumen eius;
EZEK|31|4|aquae nutrierunt illum,abyssus exaltavit eum,flumina eius manabantin circuitu radicum eius,et rivos suos emisitad universa ligna campi.
EZEK|31|5|Propterea elevata est altitudo eiussuper omnia ligna campi,et multiplicata sunt arbusta eius,et elevati sunt rami eiuspropter aquas multas.
EZEK|31|6|Cumque extendisset umbram suam,in ramis eius fecerunt nidosomnia volatilia caeli,et sub frondibus eius genueruntomnes bestiae campi,et sub umbra illius habitabatuniversa multitudo gentium;
EZEK|31|7|eratque pulcherrimus in magnitudine suaet in dilatatione arbustorum suorum,erat enim radix illiusiuxta aquas multas.
EZEK|31|8|Cedri non fuerunt pares illiin paradiso Dei;abietes non adaequaveruntramos eius,et platani non fueruntaequae frondibus illius;omne lignum paradisi Deinon est assimilatum illi et pulchritudini eius,
EZEK|31|9|quoniam speciosum feci eumet multis condensisque frondibus:et aemulata sunt eum omnia ligna Eden,quae erant in paradiso Dei.
EZEK|31|10|Propterea haec dicit Dominus Deus: Pro eo quod sublimatus est in altitudine et dedit summitatem suam usque in nubes, et elevatum est cor eius in altitudine sua,
EZEK|31|11|tradam eum in manu potentis principis gentium; faciens faciet ei: iuxta impietatem eius eieci eum.
EZEK|31|12|Et succident illum alieni, violentissimi nationum; et proicient eum super montes, et in cunctis convallibus corruent rami eius, et confringentur arbusta eius in universis voraginibus terrae, et recedent de umbra eius omnes populi terrae et relinquent eum.
EZEK|31|13|Super ruinam eius habitabuntomnia volatilia caeli,et in ramis eius eruntuniversae bestiae campi,
EZEK|31|14|ne eleventur in altitudine suaomnia ligna aquarum neque ponantsublimitatem suam inter nubes necstent apud eas in sublimitate suaomnia, quae irrigantur aquis, quiaomnes traditi sunt in mortemad inferiora terrae,in medio filiorum hominum,ad eos, qui descendunt in lacum.
EZEK|31|15|Haec dicit Dominus Deus: In die, quando descendit ad inferos, induxi luctum, operui propter eum abyssum et prohibui flumina eius et coercui aquas multas; obscuravi super eum Libanum, et omnia ligna agri concussa sunt.
EZEK|31|16|A sonitu ruinae eius commovi gentes, cum deducerem eum ad infernum cum his, qui descendebant in lacum; et consolata sunt in inferioribus terrae omnia ligna Eden, egregia atque praeclara in Libano, universa, quae irrigabantur aquis.
EZEK|31|17|Nam et ipsi cum eo descenderunt ad infernum ad interfectos gladio et auxiliatores eius, qui sederant sub umbra eius in medio nationum.
EZEK|31|18|Cui assimilatus es, o inclite atque sublimis inter ligna Eden? Et ecce deductus es cum lignis Eden ad inferiora terrae; in medio incircumcisorum dormies cum his, qui interfecti sunt gladio. Ipse est pharao et omnis pompa eius ", dicit Dominus Deus.
EZEK|32|1|Et factum est duodecimo anno, in mense duodecimo, in una mensis, factum est verbum Domini ad me dicens:
EZEK|32|2|" Fili hominis, assume lamentum super pharaonem, regem Aegypti, et dices ad eum:Leo gentium peristi,et eras sicut draco in mari;et bulliebas in fluminibus tuiset conturbabas aquas pedibus tuiset turbida faciebas flumina earum.
EZEK|32|3|Haec dicit Dominus Deus:Expandam super te rete meumin coetu populorum multorum,et extrahent te in sagena mea;
EZEK|32|4|et proiciam te in terram,super faciem agri abiciam teet habitare faciam super te omnia volatilia caeliet saturabo de te bestias universae terrae;
EZEK|32|5|et dabo carnes tuas super monteset implebo valles sanie tua.
EZEK|32|6|Et irrigabo terram paedoresanguinis tui super montes,et voragines implebuntur ex te;
EZEK|32|7|et operiam, cum exstinctus fueris, caelumet nigrescere faciam stellas eius:solem nube tegam,et luna non dabit lumen suum;
EZEK|32|8|omnia luminaria caelimaerere faciam super teet dabo tenebras super terram tuam,dicit Dominus Deus.
EZEK|32|9|Et commovebo cor populorum multorum, cum induxero contritionem tuam in gentibus super terras, quas nescis.
EZEK|32|10|Et stupescere faciam super te populos multos, et reges eorum horrore nimio formidabunt super te, cum volare coeperit gladius meus coram facie eorum, et obstupescet tremefactus unusquisque pro anima sua in die ruinae tuae.
EZEK|32|11|Quia haec dicit Dominus Deus: Gladius regis Babylonis veniet tibi,
EZEK|32|12|in gladiis fortium deiciam multitudinem tuam;violentissimae gentium omnium haeet vastabunt superbiam Aegypti,et dissipabitur omnis pompa eius.
EZEK|32|13|Et perdam omnia iumenta eius,quae erant super aquas plurimas,et non conturbabit eas pes hominis ultra,neque ungula iumentorum turbabit eas;
EZEK|32|14|tunc purissimas reddam aquas eorumet flumina eorum quasi oleum adducam,ait Dominus Deus.
EZEK|32|15|Cum dedero terram Aegypti desolatam,deseretur autem terra a plenitudine sua, quando percussero omnes habitatores eius,scient quia ego Dominus.
EZEK|32|16|Planctus est, et plangent eum; filiae gentium plangent eum, super Aegyptum et super omnem pompam eius plangent eum ", ait Dominus Deus.
EZEK|32|17|Et factum est in duodecimo anno, in quinta decima mensis, factum est verbum Domini ad me dicens:
EZEK|32|18|" Fili hominis, cane lugubre super pompam Aegypti et detrahe eam, ipsam et filias gentium robustarum ad inferiora terrae cum his, qui descendunt in lacum.
EZEK|32|19|Quo pulchrior es?Descende et dormi cum incircumcisis.
EZEK|32|20|In medio interfectorum gladio cadent; gladius datus est, attraxerunt eam et omnes populos eius.
EZEK|32|21|Loquentur ei potentissimi robustorum de medio inferni, cum auxiliatoribus eius descenderunt:Tacent incircumcisi interfecti gladio!".
EZEK|32|22|Ibi Assyria et omnis multitudo eius, in circuitu illius sepulcra eius, omnes interfecti, qui ceciderunt gladio;
EZEK|32|23|quorum data sunt sepulcra in profundissimis laci, et facta est multitudo eius per gyrum sepulcri eius; universi interfecti, cadentes gladio, qui dederant quondam formidinem in terra viventium.
EZEK|32|24|Ibi Elam et omnis pompa eius per gyrum sepulcri sui; omnes hi interfecti ruentesque gladio, qui descenderunt incircumcisi ad inferiora terrae, qui dederant quondam formidinem suam in terra viventium et sustulerunt ignominiam suam cum his, qui descendunt in lacum.
EZEK|32|25|In medio interfectorum posuerunt cubile eius, in omni pompa eius, in circuitu eius sepulcra illius, omnes hi incircumcisi interfectique gladio; dederant enim terrorem suum in terra viventium et sustulerunt ignominiam suam cum his, qui descendunt in lacum, in medio interfectorum positi sunt.
EZEK|32|26|Ibi Mosoch, Thubal et omnis pompa eius, in circuitu illius sepulcra eius, omnes hi incircumcisi interfectique gladio, quia dederunt formidinem suam in terra viventium;
EZEK|32|27|et non dormient cum fortibus, qui ceciderunt a saeculo et descenderunt ad infernum cum armis suis et posuerunt gladios suos sub capitibus suis, et fuerunt scuta eorum super ossa eorum, quia terror fortium erat in terra viventium.
EZEK|32|28|Et tu ergo in medio incircumcisorum contereris et dormies cum interfectis gladio.
EZEK|32|29|Ibi Idumaea, reges eius et omnes duces eius, qui dati sunt in robore suo cum interfectis gladio et qui cum incircumcisis dormiunt et cum his, qui descenderunt in lacum.
EZEK|32|30|Ibi principes aquilonis omnes et universi Sidonii, qui deducti sunt cum interfectis in terrore suo, in sua fortitudine confusi; qui dormiunt incircumcisi cum interfectis gladio et sustulerunt confusionem suam cum his, qui descendunt in lacum.
EZEK|32|31|Videbit eos pharao et consolabitur super universa pompa sua. Interfecti sunt gladio pharaonis et omnis exercitus eius, ait Dominus Deus,
EZEK|32|32|quia dedi terrorem meum in terra viventium; et prostratus est in medio incircumcisorum cum interfectis gladio pharaonis et omnis pompa eius ", ait Dominus Deus.
EZEK|33|1|Et factum est verbum Do mini ad me dicens:
EZEK|33|2|" Fili ho minis, loquere ad filios populi tui et dices ad eos: Terra, cum induxero super eam gladium, et tulerit populus terrae virum unum de finibus suis et constituerit eum sibi speculatorem,
EZEK|33|3|et ille viderit gladium venientem super terram et cecinerit bucina et annuntiaverit populo;
EZEK|33|4|audiens autem quisquis ille est sonum bucinae, non se observaverit, veneritque gladius et tulerit eum: sanguis ipsius super caput eius erit;
EZEK|33|5|sonum bucinae audivit et non se observavit, sanguis eius in ipso erit. Si autem se custodierit, animam suam salvavit.
EZEK|33|6|Quod si speculator viderit gladium venientem et non insonuerit bucina, et populus non se custodierit; veneritque gladius et tulerit de eis animam: ille quidem in iniquitate sua captus est, sanguinem autem eius de manu speculatoris requiram.
EZEK|33|7|Te autem, fili hominis, speculatorem dedi domui Israel. Audiens ergo ex ore meo sermonem, commonebis eos ex me.
EZEK|33|8|Si, me dicente ad impium: Impie, morte morieris, non fueris locutus, ut se custodiat impius a via sua, ipse impius in iniquitate sua morietur, sanguinem autem eius de manu tua requiram.
EZEK|33|9|Si autem commonueris impium, ut a viis suis convertatur, et ille non fuerit conversus a via sua, ipse in iniquitate sua morietur, porro tu animam tuam liberasti.
EZEK|33|10|Tu ergo, fili hominis, dic ad domum Israel: Sic locuti estis, dicentes: Iniquitates nostrae et peccata nostra super nos sunt, et in ipsis nos tabescimus; quomodo ergo vivere poterimus?".
EZEK|33|11|Dic ad eos: Vivo ego, dicit Dominus Deus; nolo mortem impii, sed ut revertatur impius a via sua et vivat. Convertimini, convertimini a viis vestris pessimis; et quare moriemini, domus Israel?
EZEK|33|12|Tu itaque, fili hominis, dic ad filios populi tui: Iustitia iusti non liberabit eum in quacumque die praevaricatus fuerit; et impietas impii non nocebit ei in quacumque die conversus fuerit ab impietate sua; et iustus non poterit vivere in iustitia sua in quacumque die peccaverit.
EZEK|33|13|Etiamsi dixero iusto quod vita vivat, et, confisus in iustitia sua, fecerit iniquitatem, omnes iustitiae eius oblivioni tradentur, et in iniquitate sua, quam operatus est, in ipsa morietur.
EZEK|33|14|Sin autem dixero impio: Morte morieris, et egerit paenitentiam a peccato suo feceritque iudicium et iustitiam,
EZEK|33|15|pignus restituerit ille impius rapinamque reddiderit, in mandatis vitae ambulaverit nec fecerit quidquam iniustum, vita vivet et non morietur;
EZEK|33|16|omnia peccata eius, quae peccavit, non imputabuntur ei: iudicium et iustitiam fecit, vita vivet.
EZEK|33|17|Et dicunt filii populi tui: "Non est aequa via Domini"; et ipsorum via iniqua est.
EZEK|33|18|Cum enim recesserit iustus a iustitia sua feceritque iniquitates, morietur in eis;
EZEK|33|19|et cum recesserit impius ab impietate sua feceritque iudicium et iustitiam, vivet in eis.
EZEK|33|20|Et dicitis: "Non est recta via Domini". Unumquemque iuxta vias suas iudicabo de vobis, domus Israel ".
EZEK|33|21|Et factum est in duodecimo anno, in decimo, in quinta mensis transmigrationis nostrae, venit ad me, qui fugerat de Ierusalem, dicens: " Vastata est civitas ".
EZEK|33|22|Manus autem Domini facta fuerat ad me vespere, antequam veniret qui fugerat; aperuitque os meum, donec veniret ad me mane, et, aperto ore meo, non silui amplius.
EZEK|33|23|Et factum est verbum Domini ad me dicens:
EZEK|33|24|" Fili hominis, qui habitant in ruinosis his super humum Israel, loquentes aiunt: "Unus erat Abraham et hereditate possedit terram; nos autem multi, nobis data est terra in possessionem".
EZEK|33|25|Idcirco dices ad eos: Haec dicit Dominus Deus: Qui in sanguine comeditis et oculos vestros levatis ad idola vestra et sanguinem funditis, numquid terram hereditate possidebitis?
EZEK|33|26|Stetistis in gladiis vestris, fecistis abominationes, et unusquisque uxorem proximi sui polluit, et terram hereditate possidebitis?
EZEK|33|27|Haec dices ad eos: Sic dicit Dominus Deus: Vivo ego, qui in ruinosis habitant, gladio cadent; et, qui in agro est, bestiis tradetur ad devorandum; qui autem in praesidiis et in speluncis sunt, peste morientur.
EZEK|33|28|Et dabo terram in solitudinem et desertum, et deficiet superba fortitudo eius, et desolabuntur montes Israel, ita ut nullus sit qui per eos transeat;
EZEK|33|29|et scient quia ego Dominus, cum dedero terram desolatam et desertam propter universas abominationes suas, quas operati sunt.
EZEK|33|30|Et tu, fili hominis, filii populi tui, qui loquuntur de te iuxta parietes et in ostiis domorum et dicunt unus ad alterum, vir ad fratrem suum, loquentes: "Venite et audite, qui sit sermo egrediens a Domino".
EZEK|33|31|Et veniunt ad te quasi si conveniat populus, et sedent coram te populus meus; et audiunt sermones tuos et non faciunt eos, quia quasi amatores loquuntur, et avaritiam suam sequitur cor eorum.
EZEK|33|32|Et es eis quasi carmen amatorum, quod suavi voce et cum dulci chordarum sono canitur, et audiunt verba tua et non faciunt ea.
EZEK|33|33|Et cum venerit, quod praedictum est - ecce enim venit - tunc scient quod prophetes fuerit inter eos ".
EZEK|34|1|Et factum est verbum Do mini ad me dicens:
EZEK|34|2|" Fili ho minis, propheta de pastoribus Israel, propheta et dices pastoribus: Haec dicit Dominus Deus: Vae pastoribus Israel, qui pascebant semetipsos! Nonne greges pascuntur a pastoribus?
EZEK|34|3|Lac comedebatis et lana operiebamini et, quod crassum erat, occidebatis, gregem autem non pascebatis;
EZEK|34|4|quod infirmum fuit, non consolidastis et, quod aegrotum, non sanastis; quod fractum est, non alligastis et, quod eiectum est, non reduxistis et, quod perierat, non quaesistis et super forte imperabatis cum violentia.
EZEK|34|5|Et dispersae sunt oves meae, eo quod non esset pastor; et factae sunt in devorationem omnium bestiarum agri et dispersae sunt.
EZEK|34|6|Erraverunt greges mei in cunctis montibus et in universo colle excelso, et super omnem faciem terrae dispersi sunt greges mei; et non erat qui requireret, non erat qui requireret.
EZEK|34|7|Propterea, pastores, audite verbum Domini:
EZEK|34|8|Vivo ego, dicit Dominus Deus, pro eo quod factus est grex meus in rapinam et oves meae in devorationem omnium bestiarum agri, eo quod non esset pastor, neque enim quaesierunt pastores mei gregem meum, sed pascebant pastores semetipsos et gregem meum non pascebant,
EZEK|34|9|propterea, pastores, audite verbum Domini.
EZEK|34|10|Haec dicit Dominus Deus: Ecce ego ipse super pastores requiram gregem meum de manu eorum et cessare eos faciam, ut ultra non pascant gregem nec pascant amplius pastores semetipsos; et liberabo gregem meum de ore eorum, et non erit ultra eis in escam.
EZEK|34|11|Quia haec dicit Dominus Deus: Ecce ego ipse requiram oves meas et visitabo eas.
EZEK|34|12|Sicut visitat pastor gregem suum in die, quando fuerit in medio ovium suarum dissipatarum, sic visitabo oves meas et liberabo eas de omnibus locis, in quibus dispersae fuerant in die nubis et caliginis.
EZEK|34|13|Et educam eas de populis et congregabo eas de terris et inducam eas in terram suam et pascam eas in montibus Israel, in rivis et in cunctis sedibus terrae.
EZEK|34|14|In pascuis uberrimis pascam eas, et in montibus excelsis Israel erunt pascua earum; ibi requiescent in herbis virentibus et in pascuis pinguibus pascentur super montes Israel.
EZEK|34|15|Ego pascam oves meas et ego eas accubare faciam, dicit Dominus Deus.
EZEK|34|16|Quod perierat, requiram et, quod eiectum erat, reducam et, quod confractum fuerat, alligabo et, quod infirmum erat, consolidabo et, quod pingue et forte, custodiam et pascam illas in iudicio.
EZEK|34|17|Vos autem, grex meus, haec dicit Dominus Deus: Ecce ego iudico inter pecus et pecus, inter arietes et hircos.
EZEK|34|18|Nonne satis vobis erat pascuam bonam depasci? Insuper et reliquias pascuarum vestrarum conculcastis pedibus vestris et, cum purissimam aquam biberetis, reliquam pedibus vestris turbabatis;
EZEK|34|19|et oves meae his, quae conculcata pedibus vestris fuerant, pascebantur et, quae pedes vestri turbaverant, haec bibebant.
EZEK|34|20|Propterea haec dicit Dominus Deus ad eos: Ecce ego ipse iudico inter pecus pingue et macilentum;
EZEK|34|21|pro eo quod lateribus et umeris impingebatis et cornibus vestris ventilabatis omnia infirma pecora, donec dispergerentur foras,
EZEK|34|22|salvabo gregem meum, et non erit ultra in rapinam, et iudicabo inter pecus et pecus.
EZEK|34|23|Et suscitabo super eas pastorem unum, qui pascat eas, servum meum David; ipse pascet eas et ipse erit eis in pastorem.
EZEK|34|24|Ego autem Dominus ero eis in Deum, et servus meus David princeps in medio eorum. Ego Dominus locutus sum.
EZEK|34|25|Et faciam cum eis pactum pacis et cessare faciam bestias pessimas de terra, et habitabunt in deserto securi et dormient in saltibus;
EZEK|34|26|et ponam eos et, quae sunt in circuitu collis mei, benedictionem et deducam imbrem in tempore suo: pluviae benedictionis erunt.
EZEK|34|27|Et dabit lignum agri fructum suum, et terra dabit germen suum, et erunt in terra sua absque timore et scient quia ego Dominus, cum contrivero vectes iugi eorum et eruero eos de manu imperantium sibi.
EZEK|34|28|Et non erunt ultra in rapinam gentibus, neque bestiae terrae devorabunt eos, sed habitabunt confidenter absque ullo terrore.
EZEK|34|29|Et suscitabo eis germen nominatum, et non erunt ultra imminuti fame in terra neque portabunt ultra opprobrium gentium;
EZEK|34|30|et scient quia ego Dominus Deus eorum cum eis, et ipsi populus meus domus Israel, ait Dominus Deus.
EZEK|34|31|Vos autem grex meus, grex pascuae meae vos, et ego Dominus Deus vester, dicit Dominus Deus.
EZEK|35|1|Et factus est sermo Domini ad me dicens:
EZEK|35|2|" Fili hominis, pone faciem tuam adversum montem Seir et propheta de eo et dices illi:
EZEK|35|3|Haec dicit Dominus Deus:Ecce ego ad te, mons Seir;et extendam manum meam super teet dabo te desolatum atque desertum.
EZEK|35|4|Urbes tuas demoliar,et tu desertus eriset scies quia ego Dominus.
EZEK|35|5|Eo quod fueris inimicus sempiternus et concluseris filios Israel in manus gladii in tempore afflictionis eorum, in tempore poenae extremae;
EZEK|35|6|propterea, vivo ego, dicit Dominus Deus, sanguini tradam te, et sanguis te persequetur et, cum sanguinem non oderis, sanguis persequetur te.
EZEK|35|7|Et dabo montem Seir desolatum atque desertum et auferam de eo euntem et redeuntem
EZEK|35|8|et implebo montes eius occisorum suorum, in collibus tuis et in vallibus tuis, atque in omnibus torrentibus tuis interfecti gladio cadent.
EZEK|35|9|In solitudines sempiternas tradam te, et civitates tuae non habitabuntur, et scietis quoniam ego Dominus.
EZEK|35|10|Eo quod dixeris: "Duae gentes et duae terrae meae erunt, et hereditate possidebo eas!", cum Dominus esset ibi;
EZEK|35|11|propterea, vivo ego, dicit Dominus Deus, faciam iuxta iram tuam et secundum zelum tuum, quem fecisti odio habens eos, et notus efficiar in eis, cum te iudicavero.
EZEK|35|12|Et scies quia ego Dominus audivi universa opprobria tua, quae locutus es de montibus Israel dicens: "Deserti nobis ad devorandum dati sunt!".
EZEK|35|13|Et insurrexistis super me ore vestro et vociferati estis vobis adversum me verba vestra; ego audivi.
EZEK|35|14|Haec dicit Dominus Deus: Laetante universa terra, in solitudinem te redigam;
EZEK|35|15|sicuti gavisus es super hereditatem domus Israel, eo quod fuerit dissipata, sic faciam tibi: dissipatus eris, mons Seir, et Idumaea omnis, et scient quia ego Dominus.
EZEK|36|1|Tu autem, fili hominis, pro pheta super montes Israel et dices: Montes Israel, audite verbum Domini.
EZEK|36|2|Haec dicit Dominus Deus: Eo quod dixerit inimicus de vobis: "Euge, altitudines sempiternae in hereditatem datae sunt nobis";
EZEK|36|3|propterea vaticinare et dic: Haec dicit Dominus Deus: Pro eo quod desolati estis, et inhiaverunt vobis per circuitum, ut fieretis in hereditatem reliquis gentibus, et ascendistis super labium linguae et opprobrium populi;
EZEK|36|4|propterea, montes Israel, audite verbum Domini Dei: Haec dicit Dominus Deus montibus et collibus, torrentibus vallibusque et desertis dissipatis et urbibus derelictis, quae depopulatae sunt et subsannatae a reliquis gentibus per circuitum;
EZEK|36|5|propterea haec dicit Dominus Deus: In igne zeli mei locutus sum de reliquis gentibus et de Idumaea universa, quae dederunt terram meam sibi in hereditatem cum gaudio et toto corde et ex animo maligno, ut pascua eius depraedarentur.
EZEK|36|6|Idcirco vaticinare super humum Israel et dices montibus et collibus, torrentibus et vallibus: Haec dicit Dominus Deus: Ecce ego in zelo meo et in furore meo locutus sum, eo quod confusionem gentium sustinueritis;
EZEK|36|7|idcirco haec dicit Dominus Deus: Ego levavi manum meam: gentes, quae in circuitu vestro sunt, ipsae confusionem suam portabunt;
EZEK|36|8|vos autem, montes Israel, ramos vestros germinabitis et fructum vestrum afferetis populo meo Israel, prope est enim ut veniat.
EZEK|36|9|Quia ecce ego ad vos et convertar ad vos, et arabimini et accipietis sementem;
EZEK|36|10|et multiplicabo in vobis homines, omnem domum Israel, et habitabuntur civitates, et ruinosa instaurabuntur.
EZEK|36|11|Et replebo vos hominibus et iumentis, et multiplicabuntur et crescent; et habitari vos faciam, sicut a principio bonisque donabo maioribus quam habuistis ab initio, et scietis quia ego Dominus.
EZEK|36|12|Et adducam super vos homines, populum meum Israel, et hereditate possidebunt te, et eris eis in hereditatem et non addes ultra ut eos facias absque liberis.
EZEK|36|13|Haec dicit Dominus Deus: Pro eo quod dicunt de vobis: "Devoratrix hominum es et faciens gentem tuam absque liberis";
EZEK|36|14|propterea homines non comedes amplius et gentem tuam non facies ultra absque liberis, ait Dominus Deus.
EZEK|36|15|Nec auditam faciam in te amplius ignominiam gentium, et opprobrium populorum nequaquam portabis ultra et gentem tuam non facies amplius absque liberis ", ait Dominus Deus.
EZEK|36|16|Et factum est verbum Domini ad me dicens:
EZEK|36|17|" Fili hominis, domus Israel habitaverunt in humo sua et polluerunt eam in viis suis et in operibus suis; iuxta immunditiam menstruatae facta est via eorum coram me.
EZEK|36|18|Et effudi indignationem meam super eos pro sanguine, quem fuderunt super terram, et in idolis suis polluerunt eam.
EZEK|36|19|Et dispersi eos in gentes, et ventilati sunt in terras; iuxta vias eorum et iuxta opera eorum iudicavi eos.
EZEK|36|20|Et ingressi sunt ad gentes, ad quas introierunt, et polluerunt nomen sanctum meum, cum diceretur de eis: "Populus Domini iste est, et de terra eius egressi sunt".
EZEK|36|21|Et peperci nomini meo sancto, quod polluerat domus Israel in gentibus, ad quas ingressi sunt.
EZEK|36|22|Idcirco dices domui Israel: Haec dicit Domihus Deus: Non propter vos ego faciam, domus Israel, sed propter nomen sanctum meum, quod polluistis in gentibus, ad quas intrastis;
EZEK|36|23|et sanctificabo nomen meum magnum, quod pollutum est inter gentes, quod polluistis in medio earum, ut sciant gentes quia ego Dominus, ait Dominus Deus, cum sanctificatus fuero in vobis coram eis.
EZEK|36|24|Tollam quippe vos de gentibus et congregabo vos de universis terris et adducam vos in terram vestram;
EZEK|36|25|et effundam super vos aquam mundam, et mundabimini ab omnibus inquinamentis vestris, et ab universis idolis vestris mundabo vos.
EZEK|36|26|Et dabo vobis cor novum et spiritum novum ponam in medio vestri et auferam cor lapideum de carne vestra et dabo vobis cor carneum;
EZEK|36|27|et spiritum meum ponam in medio vestri et faciam, ut in praeceptis meis ambuletis et iudicia mea custodiatis et operemini.
EZEK|36|28|Et habitabitis in terra, quam dedi patribus vestris, et eritis mihi in populum, et ego ero vobis in Deum.
EZEK|36|29|Et salvabo vos ex universis inquinamentis vestris et vocabo frumentum et multiplicabo illud et non imponam vobis famem.
EZEK|36|30|Et multiplicabo fructum ligni et genimina agri, ut non portetis ultra opprobrium famis in gentibus.
EZEK|36|31|Et recordabimini viarum vestrarum pessimarum operumque non bonorum, et displicebunt vobis iniquitates vestrae et scelera vestra.
EZEK|36|32|Non propter vos ego faciam, ait Dominus Deus, notum sit vobis; confundimini et erubescite super viis vestris, domus Israel.
EZEK|36|33|Haec dicit Dominus Deus: In die, qua mundavero vos ex omnibus iniquitatibus vestris et inhabitari fecero urbes et instauravero ruinosa,
EZEK|36|34|et terra deserta fuerit exculta, quae quondam erat desolata in oculis omnis viatoris,
EZEK|36|35|dicent: "Terra illa inculta facta est ut hortus Eden, et civitates desertae et destitutae atque destructae munitae inhabitantur".
EZEK|36|36|Et scient gentes, quaecumque derelictae fuerint in circuitu vestro, quia ego Dominus aedificavi dissipata plantavique inculta; ego Dominus locutus sum et facio.
EZEK|36|37|Haec dicit Dominus Deus: Adhuc in hoc exorabor a domo Israel, ut faciam eis: multiplicabo eos sicut gregem hominum,
EZEK|36|38|ut gregem sanctum, ut gregem Ierusalem in sollemnitatibus eius; sic erunt civitates desertae plenae gregibus hominum, et scient quia ego Dominus ".
EZEK|37|1|Facta est super me manus Domini et eduxit me in spiri tu Domini et posuit me in medio campi, qui erat plenus ossibus,
EZEK|37|2|et circumduxit me per ea in gyro: erant autem multa valde super faciem campi siccaque vehementer.
EZEK|37|3|Et dixit ad me: " Fili hominis, putasne vivent ossa ista? ". Et dixi: " Domine, tu nosti ".
EZEK|37|4|Et dixit ad me: " Vaticinare super ossa ista et dices eis: Ossa arida, audite verbum Domini.
EZEK|37|5|Haec dicit Dominus Deus ossibus his: Ecce ego intromittam in vos spiritum, et vivetis,
EZEK|37|6|et dabo super vos nervos et succrescere faciam super vos carnes et superextendam in vobis cutem et dabo vobis spiritum, et vivetis et scietis quia ego Dominus ".
EZEK|37|7|Et prophetavi, sicut praeceperat mihi. Factus est autem sonitus, prophetante me, et ecce commotio; et accesserunt ossa ad ossa, unumquodque ad iuncturam suam.
EZEK|37|8|Et vidi: et ecce super ea nervi et carnes ascenderunt, et extenta est in eis cutis desuper, sed spiritum non habebant.
EZEK|37|9|Et dixit ad me: " Vaticinare ad spiritum; vaticinare, fili hominis, et dices ad spiritum: Haec dicit Dominus Deus: A quattuor ventis veni, spiritus, et insuffla super interfectos istos, ut reviviscant ".
EZEK|37|10|Et prophetavi, sicut praeceperat mihi, et ingressus est in ea spiritus; et vixerunt steteruntque super pedes suos, exercitus grandis nimis valde.
EZEK|37|11|Et dixit ad me: " Fili hominis, ossa haec universa domus Israel est. Ipsi dicunt: "Aruerunt ossa nostra, et periit spes nostra, et abscissi sumus".
EZEK|37|12|Propterea vaticinare et dices ad eos: Haec dicit Dominus Deus: Ecce ego aperiam tumulos vestros et educam vos de sepulcris vestris, populus meus, et inducam vos in terram Israel;
EZEK|37|13|et scietis quia ego Dominus, cum aperuero sepulcra vestra et eduxero vos de tumulis vestris, populus meus.
EZEK|37|14|Et dabo spiritum meum in vobis, et vivetis, et collocabo vos super humum vestram, et scietis quia ego Dominus. Locutus sum et facio ", ait Dominus Deus.
EZEK|37|15|Et factus est sermo Domini ad me dicens:
EZEK|37|16|" Et tu, fili hominis, sume tibi lignum unum et scribe super illud: Iudae et filiis Israel sociis eius. Et tolle lignum alterum et scribe super illud: Ioseph, lignum Ephraim, et cunctae domui Israel sociis eius.
EZEK|37|17|Et adiunge illa unum ad alterum tibi in lignum unum; et erunt in unionem in manu tua.
EZEK|37|18|Cum autem dixerint ad te filii populi tui loquentes: "Nonne indicas nobis, quid in his tibi velis?",
EZEK|37|19|loqueris ad eos: Haec dicit Dominus Deus: Ecce ego assumam lignum Ioseph, quod est in manu Ephraim, et tribus Israel, quae iunctae sunt ei, et dabo eas pariter cum ligno Iudae et faciam eas in lignum unum, et erunt unum in manu mea.
EZEK|37|20|Erunt autem ligna, super quae scripseris, in manu tua in oculis eorum,
EZEK|37|21|et dices ad eos: Haec dicit Dominus Deus: Ecce ego assumam filios Israel de medio nationum, ad quas abierunt, et congregabo eos undique et adducam eos ad humum suam
EZEK|37|22|et faciam eos in gentem unam in terra, in montibus Israel; et rex unus erit omnibus imperans, et non erunt ultra duae gentes nec dividentur amplius in duo regna.
EZEK|37|23|Neque polluentur ultra in idolis suis et abominationibus suis et in cunctis iniquitatibus suis, et salvos eos faciam de universis aversionibus suis, quibus peccaverunt, et mundabo eos, et erunt mihi populus, et ego ero eis Deus.
EZEK|37|24|Et servus meus David rex super eos, et pastor unus erit omnium eorum; in iudiciis meis ambulabunt et mandata mea custodient et facient ea.
EZEK|37|25|Et habitabunt super terram, quam dedi servo meo Iacob, in qua habitaverunt patres vestri; et habitabunt super eam, ipsi et filii eorum et filii filiorum eorum usque in sempiternum, et David servus meus princeps eorum in perpetuum.
EZEK|37|26|Et percutiam illis foedus pacis, pactum sempiternum erit eis, et fundabo eos et multiplicabo; et dabo sanctuarium meum in medio eorum in perpetuum,
EZEK|37|27|et erit habitaculum meum in eis, et ero eis Deus, et ipsi erunt mihi populus;
EZEK|37|28|et scient gentes quia ego Dominus sanctificator Israel, cum fuerit sanctuarium meum in medio eorum in perpetuum ".
EZEK|38|1|Et factus est sermo Domini ad me dicens:
EZEK|38|2|" Fili hominis, pone faciem tuam contra Gog, in terra Magog, principem summum Mosoch et Thubal, et vaticinare de eo
EZEK|38|3|et dices: Haec dicit Dominus Deus: Ecce ego ad te, Gog, principem summum Mosoch et Thubal,
EZEK|38|4|et circumagam te et ponam uncos in maxillis tuis et educam te et omnem exercitum tuum, equos et equites vestitos perfecte universos, multitudinem magnam cum scuto et clipeo arripientes gladium.
EZEK|38|5|Persae, Chus et Phut cum eis, omnes scutati et galeati;
EZEK|38|6|Gomer et universa agmina eius, domus Thogorma de extremo aquilone et totum robur eius, populi multi tecum.
EZEK|38|7|Praepara et instrue te et omnem multitudinem tuam, quae coacervata est ad te, et esto mihi in custodiam.
EZEK|38|8|Post dies multos evocaberis; in novissimo annorum venies ad terram, quae reversa est a gladio, congregata est de populis multis ad montes Israel, qui fuerunt deserti iugiter: haec de populis educta est, et habitant in ea confidenter universi.
EZEK|38|9|Ascendens autem quasi tempestas venies, quasi nubes, ut operias terram, tu et omnia agmina tua et populi multi tecum.
EZEK|38|10|Haec dicit Dominus Deus: In die illa ascendent sermones super cor tuum, et cogitabis cogitationem pessimam
EZEK|38|11|et dices: "Ascendam ad terram absque muro, veniam ad quiescentes habitantesque secure; hi omnes habitant sine muro, vectes et portae non sunt eis";
EZEK|38|12|ut diripias spolia et capias praedam, ut inferas manum tuam super deserta iterum inhabitata et super populum, qui est congregatus ex gentibus, qui acquisivit pecora et substantiam et habitat in umbilico terrae.
EZEK|38|13|Saba et Dedan et negotiatores Tharsis et omnes principes eius dicent tibi: "Numquid ad sumenda spolia tu venis? Numquid ad diripiendam praedam congregasti multitudinem tuam, ut tollas argentum et aurum, auferas pecora atque substantiam et diripias manubias infinitas?".
EZEK|38|14|Propterea vaticinare, fili hominis, et dices ad Gog: Haec dicit Dominus Deus: Numquid non in die illo, cum habitaverit populus meus Israel confidenter, consurges?
EZEK|38|15|Et venies de loco tuo ab extremo aquilone, tu et populi multi tecum, ascensores equorum universi, coetus magnus et exercitus vehemens.
EZEK|38|16|Et ascendes super populum meum Israel quasi nubes, ut operias terram. In novissimis diebus erit, et adducam te super terram meam, ut sciant gentes me, cum sanctificatus fuero in te in oculis eorum, o Gog.
EZEK|38|17|Haec dicit Dominus Deus: Tu ergo ille es, de quo locutus sum in diebus antiquis in manu servorum meorum prophetarum Israel, qui prophetaverunt in diebus illis per annos, ut adducerem te super eos.
EZEK|38|18|Et erit in die illa, in die adventus Gog super terram Israel, ait Dominus Deus, ascendet indignatio mea in furore meo.
EZEK|38|19|Et in zelo meo, in igne irae meae locutus sum: In die illa erit commotio magna super terram Israel,
EZEK|38|20|et commovebuntur a facie mea pisces maris et volucres caeli et bestiae agri et omne reptile, quod movetur super humum, cunctique homines, qui sunt super faciem terrae; et subvertentur montes, et cadent rupes, et omnis murus in terram corruet.
EZEK|38|21|Et convocabo adversus eum in cunctis montibus meis gladium, ait Dominus Deus; gladius uniuscuiusque in fratrem suum dirigetur.
EZEK|38|22|Et iudicabo eum peste et sanguine et imbre vehementi et lapidibus grandinis; ignem et sulphur pluam super eum et super exercitum eius et super populos multos, qui sunt cum eo,
EZEK|38|23|et magnificabor et sanctificabor et notus ero in oculis multarum gentium, et scient quia ego Dominus.
EZEK|39|1|Tu autem, fili hominis, va ticinare adversum Gog et dices: Haec dicit Dominus Deus: Ecce ego super te, Gog, principem summum Mosoch e Thubal;
EZEK|39|2|et circumagam te et seducam te et ascendere faciam de extremo aquilone et adducam te super montes Israel.
EZEK|39|3|Et percutiam arcum tuum in manu sinistra tua et sagittas tuas de manu dextera tua deiciam.
EZEK|39|4|Super montes Israel cades, tu et omnia agmina tua et populi, qui sunt tecum; feris avibus, omni volatili et bestiis terrae dedi te devorandum:
EZEK|39|5|super faciem agri cades, quia ego locutus sum, ait Dominus Deus.
EZEK|39|6|Et emittam ignem in Magog et in his, qui habitant in insulis confidenter, et scient quia ego Dominus.
EZEK|39|7|Et nomen sanctum meum notum faciam in medio populi mei Israel et non polluam nomen sanctum meum amplius, et scient gentes quia ego Dominus, sanctus in Israel.
EZEK|39|8|Ecce venit et fit, ait Dominus Deus; haec est dies, de qua locutus sum.
EZEK|39|9|Et egredientur habitatores de civitatibus Israel et succendent et comburent arma, clipeum et scutum, arcum et sagittas et baculos, manus et contos, et succendent ea igne septem annis.
EZEK|39|10|Et non portabunt ligna de campis neque succident de saltibus, quoniam arma succendent igne et depraedabuntur eos, quibus praedae fuerant, et diripient vastatores suos, ait Dominus Deus.
EZEK|39|11|Et erit, in die illa dabo Gog locum nominatum sepulcrum in Israel, vallem viatorum ad orientem maris, quae oppilat viam praetereuntibus; et sepelient ibi Gog et omnem multitudinem eius, et vocabitur vallis Multitudinis Gog.
EZEK|39|12|Et sepelient eos domus Israel, ut mundent terram septem mensibus;
EZEK|39|13|sepeliet autem eum omnis populus terrae, et erit eis nominata dies, in qua glorificatus sum, ait Dominus Deus.
EZEK|39|14|Et viros iugiter constituent lustrantes terram, qui sepeliant eos, qui remanserant super faciem terrae, ut emundent eam; post menses autem septem quaerere incipient
EZEK|39|15|et circuibunt peragrantes terram; cumque viderint os hominis, statuent iuxta illud titulum, donec sepeliant illud pollinctores in valle Multitudinis Gog.
EZEK|39|16|Nomen quoque civitatis Amona, et mundabunt terram.
EZEK|39|17|Tu ergo, fili hominis, haec dicit Dominus Deus, dic volucri, universis avibus cunctisque bestiis agri: Convenite, properate, concurrite undique ad victimam meam, quam ego immolo vobis, victimam grandem super montes Israel, ut comedatis carnes et bibatis sanguinem.
EZEK|39|18|Carnes fortium comedetis et sanguinem principum terrae bibetis: arietes, agni et hirci taurique saginati de Basan sunt omnes;
EZEK|39|19|et comedetis adipem in saturitatem et bibetis sanguinem in ebrietatem de victima, quam ego immolabo vobis.
EZEK|39|20|Et saturabimini super mensam meam de equo et de iugali currus, de forti et de universis viris bellatoribus, ait Dominus Deus.
EZEK|39|21|Et ponam gloriam meam in gentibus, et videbunt omnes gentes iudicium meum, quod fecerim, et manum meam, quam posuerim super eos;
EZEK|39|22|et scient domus Israel quia ego Dominus Deus eorum a die illa et deinceps,
EZEK|39|23|et scient gentes quoniam in iniquitate sua capta sit domus Israel, eo quod reliquerint me, et absconderim faciem meam ab eis et tradiderim eos in manus hostium suorum, et ceciderint in gladio universi.
EZEK|39|24|Iuxta immunditiam eorum et scelera eorum feci eis et abscondi faciem meam ab illis.
EZEK|39|25|Propterea haec dicit Dominus Deus: Nunc restituam Iacob et miserebor omnis domus Israel et assumam zelum pro nomine sancto meo.
EZEK|39|26|Et portabunt confusionem suam et omnem praevaricationem, quam praevaricati sunt in me, cum habitaverint in terra sua confidenter; et nemo erit qui exterreat.
EZEK|39|27|Et reduxero eos de populis et congregavero de terris inimicorum suorum et sanctificatus fuero in eis in oculis gentium plurimarum,
EZEK|39|28|et scient quia ego Dominus Deus eorum, eo quod transtulerim eos in nationes et congregaverim eos super terram suam et non dereliquerim quemquam ex eis ibi.
EZEK|39|29|Et non abscondam ultra faciem meam ab eis, eo quod effuderim spiritum meum super domum Israel ", ait Dominus Deus.
EZEK|40|1|In vicesimo et quinto anno transmigrationis nostrae, in exordio anni, decima mensis, quarto decimo anno, postquam percussa est civitas, in ipsa hac die facta est super me manus Domini et adduxit me illuc.
EZEK|40|2|In visionibus Dei adduxit me in terram Israel et posuit me super montem excelsum nimis, super quem erat quasi aedificium civitatis ad austrum.
EZEK|40|3|Et introduxit me illuc; et ecce vir, cuius erat species quasi species aeris, et funiculus lineus in manu eius, et calamus mensurae in manu eius, stabat autem in porta.
EZEK|40|4|Et locutus est ad me idem vir: " Fili hominis, vide oculis tuis et auribus tuis audi et pone cor tuum in omnia, quae ego ostendam tibi, quia ut ostendantur tibi, adductus es huc; annuntia omnia, quae tu vides, domui Israel ".
EZEK|40|5|Et ecce murus forinsecus in circuitu domus undique, et in manu viri calamus mensurae sex cubitorum, qui habebant cubitum et palmum; et mensus est latitudinem aedificii calamo uno, altitudinem quoque calamo uno.
EZEK|40|6|Et venit ad portam, quae respiciebat viam orientalem, et ascendit per gradus eius et mensus est limen portae calamo uno latitudinem
EZEK|40|7|et cubiculum uno calamo in longum et uno calamo in latum et inter cubicula quinque cubitos et limen portae iuxta vestibulum portae intrinsecus calamo uno.
EZEK|40|8|Et mensus est vestibulum portae
EZEK|40|9|octo cubitorum et postem eius duobus cubitis; vestibulum autem portae erat intrinsecus.
EZEK|40|10|Porro cubicula portae ad viam orientalem, tria hinc et tria inde, mensura una trium et mensura una postium ex utraque parte.
EZEK|40|11|Et mensus est latitudinem ostii portae decem cubitorum et longitudinem portae tredecim cubitorum,
EZEK|40|12|et saeptum ante cubicula cubiti unius utrimque; cubicula autem sex cubitorum erant hinc et inde.
EZEK|40|13|Et mensus est portam a tecto cubiculi usque ad tectum eius a contra, latitudinem viginti et quinque cubitorum, ostium contra ostium,
EZEK|40|14|()
EZEK|40|15|et a facie ingressus portae usque ad faciem vestibuli portae intrinsecus, quinquaginta cubitos.
EZEK|40|16|Et erant fenestrae marginatae in cubiculis et in postibus intra portam undique per circuitum; similiter autem erant et in vestibulo fenestrae per gyrum intrinsecus, et ante postes pictura palmarum.
EZEK|40|17|Et eduxit me ad atrium exterius, et ecce exedrae et pavimentum stratum lapide in atrio per circuitum, triginta exedrae in circuitu pavimenti;
EZEK|40|18|et pavimentum ad latus portarum secundum longitudinem portarum; hoc erat pavimentum inferius.
EZEK|40|19|Et mensus est latitudinem a facie portae inferioris usque ad frontem portae interioris extrinsecus, centum cubitos. Sic oriens. Et sic aquilo.
EZEK|40|20|Portam quoque, quae respiciebat viam aquilonis atrii exterioris, mensus est, tam in longitudine quam in latitudine;
EZEK|40|21|et cubicula eius, tria hinc et tria inde, et postes eius et vestibulum eius secundum mensuram portae prioris; quinquaginta cubitorum longitudo eius et latitudo viginti quinque cubitorum.
EZEK|40|22|Et fenestrae vestibuli eius et sculpturae palmarum secundum mensuram portae, quae respiciebat ad orientem; et septem graduum erat ascensus eius, et vestibulum intrinsecus.
EZEK|40|23|Et porta atrii interioris contra portam aquilonis sicut in porta orientali; et mensus est a porta usque ad portam centum cubitos.
EZEK|40|24|Et duxit me ad viam australem, et ecce porta, quae respiciebat ad austrum; et mensus est postes eius et vestibulum eius iuxta mensuras superiores.
EZEK|40|25|Et fenestrae eius et vestibuli in circuitu sicut fenestrae ceterae; quinquaginta cubitorum longitudo erat et latitudo viginti quinque cubitorum.
EZEK|40|26|Et in gradibus septem ascendebatur ad eam, et vestibulum erat intrinsecus, et caelatae palmae erant, una hinc et altera inde, in postibus eius.
EZEK|40|27|Et porta erat atrio interiori in via australi, et mensus est a porta usque ad portam in via australi centum cubitos.
EZEK|40|28|Et introduxit me in atrium interius per portam australem et mensus est portam iuxta mensuras superiores;
EZEK|40|29|cubicula eius et postes eius, et vestibulum eius eisdem mensuris; et fenestrae erant ei et vestibulo eius in circuitu. Quinquaginta cubitorum longitudo erat et latitudo viginti quinque cubitorum.
EZEK|40|30|()
EZEK|40|31|Et vestibulum eius respiciebat ad atrium exterius, et palmae in postibus eius, et octo gradus erant, quibus ascendebatur ad eam.
EZEK|40|32|Et introduxit me in atrium interius per viam orientalem et mensus est portam secundum mensuras superiores;
EZEK|40|33|cubicula eius et postes eius et vestibulum eius sicut supra; et fenestrae erant ei et vestibulo eius in circuitu. Longitudo erat quinquaginta cubitorum et latitudo viginti quinque cubitorum.
EZEK|40|34|Et vestibulum eius respiciebat ad atrium exterius, et palmae caelatae in postibus eius hinc et inde et in octo gradibus ascensus eius.
EZEK|40|35|Et introduxit me ad portam, quae respiciebat ad aquilonem, et mensus est secundum mensuras superiores
EZEK|40|36|cubicula eius et postes eius et vestibulum eius; et fenestrae ei erant per circuitum. Longitudo quinquaginta cubitorum erat et latitudo viginti quinque cubitorum.
EZEK|40|37|Et vestibulum eius respiciebat ad atrium exterius, et caelatura palmarum in postibus illius hinc et inde et in octo gradibus ascensus eius.
EZEK|40|38|Et erat exedra, cuius ostium in vestibulo portae; ibi lavabunt holocaustum.
EZEK|40|39|Et in vestibulo portae duae mensae hinc et duae mensae inde, ut mactetur super eas holocaustum et pro peccato et pro delicto.
EZEK|40|40|Et ad latus extra vestibulum ad ostium portae, quae respicit ad aquilonem, duae mensae; et ad la tus alterum vestibuli portae duae mensae.
EZEK|40|41|Quattuor mensae hinc et quattuor mensae inde ad latus portae: octo mensae erant, super quas mactabunt.
EZEK|40|42|Quattuor autem mensae ad holocaustum de lapidibus quadris exstructae longitudine cubiti unius et dimidii et latitudine cubiti unius et dimidii et altitudine cubiti unius, super ista ponant vasa, quibus mactetur holocaustum et victima,
EZEK|40|43|et labia palmi unius reflexa intrinsecus per circuitum; super mensas autem carnes oblationis.
EZEK|40|44|Et extra portam interiorem exedrae duae, in atrio interiori; una erat in latere portae respicientis ad aquilonem, et facies eius contra viam australem, et una ex latere portae australis, quae respiciebat ad viam aquilonis.
EZEK|40|45|Et dixit ad me: " Haec est exedra, quae respicit viam meridianam; sacerdotum erit, qui excubant in custodiis templi.
EZEK|40|46|Porro exedra, quae respicit ad viam aquilonis, sacerdotum erit, qui excubant ad ministerium altaris: isti sunt filii Sadoc, qui accedunt de filiis Levi ad Dominum, ut ministrent ei ".
EZEK|40|47|Et mensus est atrium longitudine centum cubitorum et latitudine centum cubitorum per quadrum. Altare autem erat ante faciem templi.
EZEK|40|48|Et introduxit me in vestibulum templi; et mensus est postes vestibuli quinque cubitis hinc et quinque cubitis inde et latitudinem portae quattuordecim cubitorum et latera portae trium cubitorum hinc et trium cubitorum inde;
EZEK|40|49|longitudinem autem vestibuli viginti cubitorum et latitudinem duodecim cubitorum, et decem gradibus ascendebatur ad illud, et columnae erant in postibus, una hinc et altera inde.
EZEK|41|1|Et introduxit me in templum et mensus est postes: sex cu bitos latitudinis hinc et sex cubitos latitudinis inde.
EZEK|41|2|Et latitudo portae decem cubitorum erat, et latera portae quinque cubitis hinc et quinque cubitis inde; et mensus est longitudinem eius quadraginta cubitorum et latitudinem viginti cubitorum.
EZEK|41|3|Et introgressus intrinsecus, mensus est in poste portae duos cubitos et portam sex cubitorum et latitudinem laterum portae septem cubitorum hinc et septem cubitorum inde.
EZEK|41|4|Et mensus est longitudinem eius viginti cubitorum et latitudinem viginti cubitorum versus faciem templi. Et dixit ad me: " Hoc est Sanctum sanctorum ".
EZEK|41|5|Et mensus est parietem domus sex cubitorum et latitudinem aedificii adiacentis quattuor cubitorum undique per circuitum domus;
EZEK|41|6|cubicula autem adiacentia, cubiculum super cubiculum, in tribus tabulatis. Et erant margines eminentes in pariete domus pro cubiculis adiacentibus per circuitum, ut essent fulcra, neque essent fulcra intra parietem domus,
EZEK|41|7|et latitudo ambitus sursum ascendens iuxta cubicula adiacentia, quia circumdata erat domus usque sursum circa domum; idcirco amplificata erat domus usque sursum, et de inferiore tabulato ascendebatur ad superius per medium.
EZEK|41|8|Et vidi in domo altitudinem per circuitum, fundamenta aedificii adiacentis mensura calami pleni, id est sex cubitorum, in altitudine.
EZEK|41|9|Et latitudo parietis aedificii adiacentis forinsecus erat quinque cubitorum. Et area vacua inter cubicula domui adiacentia,
EZEK|41|10|et inter exedras habebat latitudinem viginti cubitorum in circuitu domus undique.
EZEK|41|11|Et ostia aedificii adiacentis ad aream vacuam, ostium unum ad viam aquilonis et ostium unum ad viam australem; et latitudo muri areae vacuae quinque cubitorum in circuitu.
EZEK|41|12|Et aedificium, quod erat ex adverso areae separatae versumque ad viam respicientem ad mare, latitudinis septuaginta cubitorum; paries autem aedificii quinque cubitorum latitudinis per circuitum et longitudo eius nonaginta cubitorum.
EZEK|41|13|Et mensus est domus longitudinem centum cubitorum et areae separatae et aedificii et parietum eius longitudinem centum cubitorum;
EZEK|41|14|latitudinem autem faciei domus et areae separatae contra orientem centum cubitorum.
EZEK|41|15|Et mensus est longitudinem aedificii ex adverso areae separatae ad dorsum et parietum eius ex utraque parte centum cubitorum. Et templum interius et vestibulum exterius
EZEK|41|16|strata erant ligno, et fenestrae marginatae et margines in circuitu triplices contra limen erant strato ligno per gyrum in circuitu, et a terra usque ad fenestras - et fenestrae poterant claudi - usque ad superiora ostii;
EZEK|41|17|et usque ad domum interiorem et forinsecus et per omnem parietem in circuitu, intrinsecus et forinsecus, ad mensuram
EZEK|41|18|fabrefacti cherubim et palmae, et palma inter cherub et cherub; duasque facies habebat cherub,
EZEK|41|19|faciem hominis versam ad palmam ex hac parte et faciem leonis versam ad palmam ex alia parte: expressi per omnem domum in circuitu.
EZEK|41|20|De terra usque ad superiora portae cherubim et palmae caelatae erant. In pariete templi
EZEK|41|21|postes portae quadruplices, et coram sanctuario aspectus quasi aspectus
EZEK|41|22|altaris lignei trium cubitorum altitudo, et longitudo eius duorum cubitorum, et anguli eius et bases eius et parietes eius lignei. Et locutus est ad me: " Haec est mensa coram Domino ".
EZEK|41|23|Et duo ostia erant templo et sanctuario
EZEK|41|24|duo ostia. Ostiis erant duae valvae versatiles usque ad parietem, valvae duae ostio uni et valvae duae ostio alteri.
EZEK|41|25|Et caelati erant in ipsis ostiis templi cherubim et sculpturae palmarum, sicut in parietibus quoque expressi erant; et tectum ligneum erat in vestibuli fronte forinsecus.
EZEK|41|26|Et fenestrae marginatae et similitudo palmarum hinc atque inde in lateribus vestibuli et in cubiculis adiacentibus domus.
EZEK|42|1|Et eduxit me in atrium ex terius per viam ducentem ad aquilonem; et duxit me ad exedram, quae erat contra aream separatam, et contra aedem ad aquilonem.
EZEK|42|2|Longitudo erat centum cubitorum in latere aquilonis et latitudo quinquaginta cubitorum.
EZEK|42|3|Contra viginti cubitos atrii interioris et contra pavimentum stratum lapide atrii exterioris elevabatur pars iuxta partem in tribus gradibus.
EZEK|42|4|Et ante exedras deambulatio decem cubitorum latitudinis, ad interiora respiciens, longitudinis centum cubitorum; et ostia eorum ad aquilonem.
EZEK|42|5|Exedrae superiores angustiores erant, quia gradus auferebant eis spatium, prae inferioribus et mediis aedificii.
EZEK|42|6|Tristega enim erant et non habebant columnas, sicut erant columnae exteriorum; sic ergo in gradibus de inferioribus, et de mediis a terra surgebat aedificium.
EZEK|42|7|Et murus exterior secundum exedras erat in via atrii exterioris ante exedras, longitudo eius quinquaginta cubitorum,
EZEK|42|8|quia longitudo erat exedrarum atrii exterioris quinquaginta cubitorum, quae erant ante faciem illarum, totum erat centum cubitorum.
EZEK|42|9|Et erat subter exedras has introitus ab oriente ingredientibus in ea de atrio exteriori
EZEK|42|10|in capite muri atrii. Contra viam meridianam in facie areae separatae, et erant exedrae ante aedificium,
EZEK|42|11|et via ante faciem earum iuxta similitudinem exedrarum, quae erant in via aquilonis; secundum longitudinem earum et latitudinem earum, sic et omnes exitus earum et dispositiones et ostia earum.
EZEK|42|12|Et ad ostia exedrarum, quae erant in via respiciente ad notum, ostium in capite viae, quae via erat ante murum protegentem per viam orientalem ingredientibus.
EZEK|42|13|Et dixit ad me: "Exedrae aquilonis et exedrae austri, quae sunt ante aream separatam, hae sunt exedrae sanctae, in quibus vescuntur sacerdotes, qui appropinquant ad Dominum sancta sanctorum: ibi ponent sancta sanctorum et oblationem et pro peccato et pro delicto, locus enim sanctus est.
EZEK|42|14|Cum autem ingressi fuerint sacerdotes, non egredientur de sanctis in atrium exterius, sed ibi reponent vestimenta sua, in quibus ministrant, quia sancta sunt; vestienturque vestimentis aliis et sic procedent ad locum populi ".
EZEK|42|15|Cumque complesset mensuras interioris areae domus, eduxit me per viam portae, quae respiciebat ad viam orientalem, et mensus est ibi undique per circuitum.
EZEK|42|16|Mensus est autem contra ventum orientalem calamo mensurae quingentos calamos in calamo mensurae per circuitum.
EZEK|42|17|Et mensus est contra ventum aquilonis quingentos calamos in calamo mensurae per gyrum.
EZEK|42|18|Et ad ventum australem mensus est quingentos calamos in calamo mensurae per circuitum.
EZEK|42|19|Et conversus ad ventum occidentalem mensus est quingentos calamos in calamo mensurae.
EZEK|42|20|Per quattuor ventos mensus est illud; murus ei erat undique per circuitum longitudine quingentorum cubitorum et latitudine quingentorum cubitorum, dividens inter sanctuarium et locum profanum.
EZEK|43|1|Et duxit me ad portam, quae respiciebat ad viam orientalem,
EZEK|43|2|et ecce gloria Dei Israel ingrediebatur per viam orientalem, et vox erat ei quasi vox aquarum multarum, et terra splendebat a maiestate eius.
EZEK|43|3|Et vidi visionem secundum speciem, quam videram, quando venit, ut disperderet civitatem, et species secundum aspectum, quem videram iuxta fluvium Chobar; et cecidi super faciem meam.
EZEK|43|4|Et maiestas Domini ingressa est templum per viam portae, quae respiciebat ad orientem.
EZEK|43|5|Et levavit me spiritus et introduxit me in atrium interius; et ecce repleta erat gloria Domini domus.
EZEK|43|6|Et audivi loquentem ad me de domo, cum vir staret iuxta me,
EZEK|43|7|et dixit ad me: " Fili hominis, locus solii mei et locus vestigiorum pedum meorum, ubi habitabo in medio filiorum Israel in aeternum; et non polluent ultra domus Israel nomen sanctum meum, ipsi et reges eorum, in fornicationibus suis et in cadaveribus regum suorum in morte eorum,
EZEK|43|8|qui fabricati sunt limen suum iuxta limen meum et postes suos iuxta postes meos, et paries erat inter me et eos, et polluerunt nomen sanctum meum in abominationibus, quas fecerunt; propter quod consumpsi eos in ira mea.
EZEK|43|9|Nunc ergo repellant procul fornicationem suam et cadavera regum suorum a me, et habitabo in medio eorum semper.
EZEK|43|10|Tu autem, fili hominis, ostende domui Israel templum, et confundantur ab iniquitatibus suis et metiantur fabricam.
EZEK|43|11|Et si erubuerint ex omnibus, quae fecerunt, describe domum et supellectilem eius, exitus et introitus, et omnem figuram eius et universa praecepta eius et omnes leges eius ostende eis et scribes oculis eorum, ut custodiant omnem figuram eius et omnia praecepta illius et faciant ea.
EZEK|43|12|Ista est lex domus in summitate montis: omnes fines eius in circuitu sanctum sanctorum sunt; haec est ergo lex domus ".
EZEK|43|13|Istae autem mensurae altaris in cubitis, cubitus habebat cubitum et palmum; fossae in circuitu eius erat cubitus in altitudine et cubitus in latitudine; et saepto eius ad marginem eius in circuitu palmus unus. Haec autem erat altitudo altaris:
EZEK|43|14|de fossa terrae usque ad crepidinem inferiorem duo cubiti, et latitudo cubiti unius; et a crepidine minore usque ad crepidinem maiorem quattuor cubiti, et latitudo unius cubiti.
EZEK|43|15|Ipse autem focus quattuor cubitorum, et a foco usque sursum cornua quattuor.
EZEK|43|16|Et focus duodecim cubitorum in longitudine per duodecim cubitos latitudinis, quadrangulatum aequis lateribus.
EZEK|43|17|Et crepido quattuordecim cubitorum longitudinis per quattuordecim cubitos latitudinis in quattuor angulis eius; et saeptum in circuitu eius dimidii cubiti, et fossa eius unius cubiti per circuitum; gradus autem eius versi ad orientem.
EZEK|43|18|Et dixit ad me: " Fili hominis, haec dicit Dominus Deus: Hi sunt ritus altaris: in qua die fuerit fabricatum, ut offeratur super illud holocaustum, et effundatur sanguis,
EZEK|43|19|dabis sacerdotibus levitis, qui sunt de semine Sadoc, qui accedunt ad me, ait Dominus Deus, ut ministrent mihi, vitulum de armento pro peccato.
EZEK|43|20|Et assumens de sanguine eius, pones super quattuor cornua eius et super quattuor angulos crepidinis et super saeptum in circuitu et mundabis illud et expiabis.
EZEK|43|21|Et tolles vitulum, qui oblatus fuerit pro peccato, et combures illum in destinato loco domus extra sanctuarium.
EZEK|43|22|Et in die secunda offeres hircum caprarum immaculatum pro peccato, et expiabunt altare, sicut expiaverunt in vitulo.
EZEK|43|23|Cumque compleveris expians illud, offeres vitulum de armento immaculatum et arietem de grege immaculatum;
EZEK|43|24|et offeres eos in conspectu Domini, et mittent sacerdotes super eos sal et offerent eos holocaustum Domino.
EZEK|43|25|Septem diebus facies hircum pro peccato cotidie, et vitulum de armento et arietem de pecoribus immaculatos offerent.
EZEK|43|26|Septem diebus expiabunt altare et mundabunt illud et consecrabunt illud.
EZEK|43|27|Expletis autem diebus, in die octava et ultra facient sacerdotes super altare holocausta vestra et pacifica, et placatus ero vobis ", ait Dominus Deus.
EZEK|44|1|Et convertit me ad viam portae sanctuarii exterioris, quae respiciebat ad orientem, et erat clausa;
EZEK|44|2|et dixit Dominus ad me: " Porta haec clausa erit; non aperietur, et vir non transibit per eam, quoniam Dominus, Deus Israel, ingressus est per eam, eritque clausa.
EZEK|44|3|Princeps, ut princeps ipse sedebit in ea, ut comedat panem coram Domino; per viam vestibuli portae ingredietur et per eandem viam egredietur ".
EZEK|44|4|Et adduxit me per viam portae aquilonis in conspectum domus; et vidi: et ecce implevit gloria Domini domum Domini, et cecidi in faciem meam.
EZEK|44|5|Et dixit ad me Dominus: " Fili hominis, pone cor tuum et vide oculis tuis et auribus tuis audi omnia, quae ego loquor ad te de universis caeremoniis domus Domini et de cunctis legibus eius; et pones cor tuum in introitu templi et in omni exitu sanctuarii
EZEK|44|6|et dices ad exasperantem me domum Israel: Haec dicit Dominus Deus: Sufficiant vobis omnes abominationes vestrae, domus Israel,
EZEK|44|7|eo quod induxistis alienigenas incircumcisos corde et incircumcisos carne, ut essent in sanctuario meo et polluerent domum meam, cum offertis panem meum, adipem et sanguinem; et dissolvistis pactum meum in omnibus abominationibus vestris
EZEK|44|8|et non explevistis ministerium sanctorum meorum et posuistis illos ministrantes mihi in sanctuario meo. Propterea
EZEK|44|9|haec dicit Dominus Deus: Omnis alienigena incircumcisus corde et incircumcisus carne non ingredietur sanctuarium meum, omnis alienigena, qui est in medio filiorum Israel.
EZEK|44|10|Sed Levitae, qui longe recesserint a me in errore filiorum Israel, qui erraverunt a me post idola sua, portabunt iniquitatem suam
EZEK|44|11|et erunt in sanctuario meo aeditui et ianitores portarum domus et ministri domus: ipsi mactabunt holocausta et victimas populo et ipsi stabunt in conspectu eorum, ut ministrent eis.
EZEK|44|12|Pro eo quod ministraverunt illis in conspectu idolorum suorum et facti sunt domui Israel in offendiculum iniquitatis, idcirco levavi manum meam super eos, dicit Dominus Deus; portabunt iniquitatem suam.
EZEK|44|13|Et non appropinquabunt ad me, ut sacerdotio fungantur mihi, neque accedent ad omnia sancta mea, ad sanctissima, sed portabunt confusionem suam et abominationes suas, quas fecerunt.
EZEK|44|14|Et faciam eos ministros in omni ministerio domus et in universis, quae facienda sunt in ea.
EZEK|44|15|Sacerdotes autem levitae filii Sadoc, qui custodierunt caeremonias sanctuarii mei, cum errarent filii Israel a me, ipsi accedent ad me, ut ministrent mihi, et stabunt in conspectu meo, ut offerant mihi adipem et sanguinem, ait Dominus Deus.
EZEK|44|16|Ipsi ingredientur sanctuarium meum et ipsi accedent ad mensam meam, ut serviant mihi et custodiant ministerium meum.
EZEK|44|17|Cumque ingredientur portas atrii interioris, vestibus lineis induentur, nec ascendet super eos quidquam laneum, quando ministrant in portis atrii interioris et in domo.
EZEK|44|18|Vittae lineae erunt in capitibus eorum, et feminalia linea erunt in lumbis eorum, et non accingentur in sudore.
EZEK|44|19|Cumque egredientur atrium exterius ad populum, exuent se vestimenta sua, in quibus ministraverunt, et reponent ea in exedris sanctis et vestient se vestimentis aliis et non sanctificabunt populum in vestibus suis.
EZEK|44|20|Caput autem suum non radent neque comam nutrient, sed tondentes attondent capita sua.
EZEK|44|21|Et vinum non bibet omnis sacerdos, quando ingressurus est atrium interius.
EZEK|44|22|Et viduam et repudiatam non accipient sibi uxores sed virgines de semine domus Israel; sed et viduam, quae fuerit vidua a sacerdote, accipient.
EZEK|44|23|Et populum meum docebunt quid sit inter sanctum et profanum et inter mundum et immundum ostendent eis.
EZEK|44|24|Et cum fuerit controversia, stabunt ad iudicandum et in iudiciis meis iudicabunt; leges meas et praecepta mea in omnibus sollemnitatibus meis custodient et sabbata mea sanctificabunt.
EZEK|44|25|Et ad mortuum hominem non ingredientur, ne polluantur, nisi ad patrem et matrem et filium et filiam et fratrem et sororem, quae virum non habuit: in quibus contaminabuntur.
EZEK|44|26|Et postquam fuerit emundatus, septem dies numerabuntur ei,
EZEK|44|27|et in die introitus sui in sanctuarium ad atrium interius, ut ministret mihi in sanctuario, offeret pro peccato suo, ait Dominus Deus.
EZEK|44|28|Et erit eis in hereditatem: ego hereditas eorum; et possessionem non dabitis eis in Israel: ego enim possessio eorum.
EZEK|44|29|Oblationem et pro peccato et pro delicto ipsi comedent, et omne anathema in Israel ipsorum erit;
EZEK|44|30|et primitiva omnium primogenitorum et omnia libamenta ex omnibus, quae offertis, sacerdotum erunt; et primitiva farinae vestrae dabitis sacerdoti, ut reponat benedictionem domui tuae.
EZEK|44|31|Omne morticinum et captum a bestia de avibus et de pecoribus non comedent sacerdotes.
EZEK|45|1|Cumque coeperitis terram dividere sortito, separate oblationem Domino sanctificatum de terra, longitudine viginti quinque milia et latitudine viginti milia: sanctificatum erit in omni termino suo per circuitum;
EZEK|45|2|ex quo sanctuarium obtinebit quingentos per quingentos, quadrifariam per circuitum, et quinquaginta cubitos pascua eius per gyrum.
EZEK|45|3|Et a mensura ista mensurabis longitudinem viginti quinque milium et latitudinem decem milium, et in ipso erit templum, Sanctum sanctorum.
EZEK|45|4|Sanctificatum de terra erit sacerdotibus ministris sanctuarii, qui accedunt ad ministerium Domini; et erit eis locus in domos et in pascua pecoribus.
EZEK|45|5|Viginti quinque autem milia longitudinis et decem milia latitudinis erunt Levitis, qui ministrant domui; ipsis in possessionem, civitates ad habitandum.
EZEK|45|6|Et possessionem civitatis dabitis quinque milia latitudinis et longitudinis viginti quinque milia, iuxta oblationem sacram; omni domui Israel erit.
EZEK|45|7|Principi quoque ex utraque parte oblationis sacrae et possessionis civitatis, secundum oblationem sacram et possessionem urbis, a latere maris usque ad mare et a latere orientis versus orientem, longitudinem autem iuxta unamquamque partium, a termino occidentali usque ad terminum orientalem.
EZEK|45|8|Haec terra erit ei possessio in Israel, et non depopulabuntur ultra principes mei populum meum; sed terram dabunt domui Israel secundum tribus eorum.
EZEK|45|9|Haec dicit Dominus Deus: Sufficiat vobis, principes Israel; violentiam et rapinas omittite et iudicium et iustitiam facite; auferte exactiones vestras a populo meo, ait Dominus Deus.
EZEK|45|10|Statera iusta et ephi iustum et batus iustus sit vobis;
EZEK|45|11|ephi et batus aequalia et unius mensurae sint, ut capiat decimam partem homer batus, et decimam partem homer ephi: iuxta mensuram homer sit aequa libratio eorum.
EZEK|45|12|Siclus autem viginti gera habeat; quinque sicli sint quinque, et decem sicli sint decem, et quinquaginta sint vobis mina.
EZEK|45|13|Haec est oblatio, quam offeratis: sextam partem ephi de gomor frumenti et sextam partem ephi de gomor hordei.
EZEK|45|14|Praeceptum quoque de oleo - batus est mensura olei C: decimam partem bati offeratis de choro - decem bati homer faciunt, quia decem bati implent chorum C.
EZEK|45|15|Et pecus unum de grege ducentorum, de pascuis irriguis Israel, in oblationem et in holocaustum et in pacifica ad expiandum pro eis, ait Dominus Deus.
EZEK|45|16|Omnis populus terrae tenebitur ad hanc oblationem principi in Israel;
EZEK|45|17|et super principem erunt holocausta et oblationes et libamina in diebus festis et in calendis et in sabbatis et in universis sollemnitatibus domus Israel; ipse faciet pro peccato et oblationem et holocaustum et pacifica ad expiandum pro domo Israel.
EZEK|45|18|Haec dicit Dominus Deus: In primo mense, una mensis, sumes vitulum de armento immaculatum et expiabis sanctuarium.
EZEK|45|19|Et tollet sacerdos de sanguine hostiae pro peccato et ponet in postibus domus et in quattuor angulis crepidinis altaris et in postibus portae atrii interioris.
EZEK|45|20|Et sic facies in septima mensis pro unoquoque, qui ignoravit et errore deceptus est, et expiabitis pro domo.
EZEK|45|21|In primo mense, quarta decima die mensis, erit vobis Paschae sollemnitas; septem diebus azyma comedentur.
EZEK|45|22|Et faciet princeps in die illa pro se et pro universo populo terrae vitulum pro peccato;
EZEK|45|23|et in septem dierum sollemnitate faciet holocaustum Domino septem vitulos et septem arietes immaculatos cotidie septem diebus et pro peccato hircum caprarum cotidie;
EZEK|45|24|et oblationem ephi per vitulum et ephi per arietem faciet et olei hin per singula ephi.
EZEK|45|25|Septimo mense, quinta decima die mensis, in sollemnitate faciet, sicut supra dicta sunt, per septem dies, tam pro peccato quam pro holocausto et in oblatione et in oleo.
EZEK|46|1|Haec dixit Dominus Deus: Porta atrii interioris, quae respicit ad orientem, erit clausa sex diebus, in quibus opus fit; die autem sabbati aperietur, sed et in die calendarum aperietur,
EZEK|46|2|et intrabit princeps per viam vestibuli portae deforis et stabit in poste portae, et facient sacerdotes holocaustum eius et pacifica eius, et adorabit super limen portae et egredietur; porta autem non claudetur usque ad vesperam.
EZEK|46|3|Et adorabit populus terrae ad ostium portae illius in sabbatis et in calendis coram Domino.
EZEK|46|4|Holocaustum autem hoc offeret princeps Domino: in die sabbati sex agnos immaculatos et arietem immaculatum
EZEK|46|5|et oblationem ephi per arietem, per agnos autem oblationem, quantum dederit manus eius, et olei hin per singula ephi;
EZEK|46|6|in die autem calendarum vitulum de armento immaculatum et sex agni et aries immaculati erunt
EZEK|46|7|et ephi per vitulum, ephi quoque per arietem faciet oblationem, per agnos autem sicut invenerit manus eius, et olei hin per singula ephi.
EZEK|46|8|Cumque ingressurus est princeps, per viam vestibuli portae ingrediatur et per eandem viam exeat.
EZEK|46|9|Et cum intrabit populus terrae in conspectu Domini in sollemnitatibus, qui ingreditur per portam aquilonis, ut adoret, egrediatur per viam portae meridianae; porro qui ingreditur per viam portae meridianae, egrediatur per viam portae aquilonis: non revertetur per viam portae, per quam ingressus est, sed e regione illius egredietur.
EZEK|46|10|Princeps autem in medio eorum cum ingredientibus ingredietur et cum egredientibus egredietur.
EZEK|46|11|Et in diebus festis et in sollemnitatibus erit oblatio ephi per vitulum et ephi per arietem, per agnos autem erit oblatio, quantum invenerit manus eius, et olei hin per singula ephi.
EZEK|46|12|Cum autem fecerit princeps spontaneum holocaustum aut pacifica voluntaria Domino, aperietur ei porta, quae respicit ad orientem, et faciet holocaustum suum et pacifica sua, sicut facere solet in die sabbati, et egredietur, claudeturque porta, postquam exierit.
EZEK|46|13|Et agnum anniculum immaculatum facies holocaustum cotidie Domino; semper mane facies illud.
EZEK|46|14|Et oblationem facies super eo mane mane sextam partem ephi, et de oleo tertiam partem hin, ut conspergatur simila; oblatio Domino, legitimum iuge atque perpetuum.
EZEK|46|15|Facient agnum et oblationem et oleum mane mane, holocaustum sempiternum.
EZEK|46|16|Haec dixit Dominus Deus: Si dederit princeps donum alicui de filiis suis de hereditate sua, filiorum suorum erit; possidebunt illud hereditarie.
EZEK|46|17|Si autem dederit legatum de hereditate sua uni servorum suorum, erit illius usque ad annum remissionis et revertetur ad principem; sola hereditas filiorum eius illorum erit.
EZEK|46|18|Et non accipiet princeps de hereditate populi, ut expellat eos de possessione eorum, sed de possessione sua hereditatem dabit filiis suis, ut non dispergatur populus meus unusquisque a possessione sua ".
EZEK|46|19|Et introduxit me per ingressum, qui erat ex latere portae, in exedras sacras sacerdotum, quae respiciebant ad aquilonem, et erat ibi locus in extrema parte vergens ad occidentem;
EZEK|46|20|et dixit ad me: " Iste est locus, ubi coquent sacerdotes pro delicto et pro peccato, ubi coquent oblationem, ut non efferant in atrium exterius, et sanctificetur populus ".
EZEK|46|21|Et eduxit me in atrium exterius et circumduxit me per quattuor angulos atrii, et ecce atriola singula per angulos atrii.
EZEK|46|22|In quattuor angulis atrii atriola inclusa quadraginta cubitorum per longum et triginta per latum: mensurae unius quattuor erant.
EZEK|46|23|Et paries per circuitum ambiens quattuor atriola, et culinae fabricatae erant subter parietes per gyrum.
EZEK|46|24|Et dixit ad me: "Hae sunt domus culinarum, in quibus coquent ministri domus Domini victimas populi ".
EZEK|47|1|Et convertit me ad portam domus, et ecce aquae egre diebantur subter limen domus ad orientem; facies enim domus respiciebat ad orientem, aquae autem descendebant a latere templi dextro a meridie altaris.
EZEK|47|2|Et eduxit me per viam portae aquilonis et convertit me ad viam foras ad portam exteriorem, quae respiciebat ad orientem; et ecce aquae exeuntes a latere dextro.
EZEK|47|3|Cum egrederetur vir ad orientem, qui habebat funiculum in manu sua, mensus est mille cubitos et traduxit me per aquam usque ad talos.
EZEK|47|4|Rursumque mensus est mille et traduxit me per aquam usque ad genua.
EZEK|47|5|Et mensus est mille et traduxit me per aquam usque ad renes. Et mensus est mille; torrens, quem non potui pertransire, quoniam intumuerant aquae, aquae ad natandum; torrens, qui non poterat transvadari.
EZEK|47|6|Et dixit ad me: " Certe vidisti, fili hominis "; et duxit me et convertit ad ripam torrentis.
EZEK|47|7|Cumque me convertissem, ecce in ripa torrentis ligna multa nimis ex utraque parte;
EZEK|47|8|et ait ad me: " Aquae istae, quae egrediuntur ad regionem orientalem et descendunt ad Arabam, intrabunt mare, aquas salsas, et sanabuntur aquae:
EZEK|47|9|et omnis anima vivens, quae movetur, quocumque venerit torrens, vivet, et erunt pisces multi satis, postquam venerint illuc aquae istae, et sanabuntur et vivent omnia, ad quae venerit torrens.
EZEK|47|10|Et stabunt super mare piscatores; ab Engaddi usque ad Engallim siccatio sagenarum erit; plurimae species erunt piscium eius, sicut pisces maris Magni, multitudinis nimiae.
EZEK|47|11|Palustria autem eius et stagna non sanabuntur, quia in salinas dabuntur.
EZEK|47|12|Et super torrentem orietur in ripis eius ex utraque parte omne lignum pomiferum; non defluet folium ex eo, et non deficiet fructus eius: per singulos menses afferet primitiva, quia aquae eius de sanctuario egredientur, et erunt fructus eius in cibum, et folia eius ad medicinam.
EZEK|47|13|Haec dicit Dominus Deus: Hic est terminus, in quo possidebitis terram in duodecim tribubus Israel, quia Ioseph duplicem funiculum habet;
EZEK|47|14|possidebitis autem eam, singuli aeque ut frater suus, super quam levavi manum meam, ut darem patribus vestris; et cadet terra haec vobis in possessionem.
EZEK|47|15|Hic est autem terminus terrae: ad plagam septentrionalem a mari Magno via Hethalon ad introitum Emath,
EZEK|47|16|Sedada, Berotha, Sabarim, quae est inter terminum Damasci et confinium Emath, usque ad Asarenon, quae est iuxta terminum Auran;
EZEK|47|17|erit ergo terminus a mari usque ad Asarenon, cum fines Damasci et fines Emath sint in aquilone; haec est plaga septentrionalis.
EZEK|47|18|Porro plaga orientalis de loco inter Auran et inter Damascum et in medio inter Galaad et terram Israel, Iordanis disterminans usque ad mare orientale, usque Thamar; haec est plaga orientalis.
EZEK|47|19|Plaga autem australis meridiana a Thamar usque ad aquas Meribathcades et torrentem usque ad mare Magnum; haec est plaga ad meridiem australis.
EZEK|47|20|Et plaga maris, mare Magnum a confinio per directum, donec venias Emath; haec est plaga maris.
EZEK|47|21|Et dividetis terram istam vobis per tribus Israel
EZEK|47|22|et mittetis eam in hereditatem, vobis et advenis, qui accesserint ad vos, qui genuerint filios in medio vestrum, et erunt vobis sicut indigenae inter filios Israel: vobiscum divident possessionem in medio tribuum Israel;
EZEK|47|23|in tribu autem quacumque fuerit advena, ibi dabitis possessionem illi, ait Dominus Deus.
EZEK|48|1|Et haec nomina tribuum: in finibus aquilonis iuxta viam Hethalon ad introitum Emath, Asarenon - fines Damasci ad aquilonem iuxta Emath - erit a plaga orientali usque ad mare, Dan pars una.
EZEK|48|2|Et iuxta terminum Dan a plaga orientali usque ad plagam maris, Aser una.
EZEK|48|3|Et iuxta terminum Aser a plaga orientali usque ad plagam maris, Nephthali una.
EZEK|48|4|Et iuxta terminum Nephthali a plaga orientali usque ad plagam maris, Manasse una.
EZEK|48|5|Et iuxta terminum Manasse a plaga orientali usque ad plagam maris, Ephraim una.
EZEK|48|6|Et iuxta terminum Ephraim a plaga orientali usque ad plagam maris, Ruben una.
EZEK|48|7|Et iuxta terminum Ruben a plaga orientali usque ad plagam maris, Iudae una.
EZEK|48|8|Et iuxta terminum Iudae a plaga orientali usque ad plagam maris oblatio, quam separabitis viginti quinque milibus latitudinis et longitudinis, sicuti singulae partes a plaga orientali usque ad plagam maris; et erit sanctuarium in medio eius.
EZEK|48|9|Oblatio, quam separabitis Domino, longitudo viginti quinque milibus et latitudo viginti milibus.
EZEK|48|10|His autem est oblatio sacra: sacerdotibus, ad aquilonem viginti quinque milia et ad mare latitudinis decem milia et ad orientem latitudinis decem milia et ad meridiem longitudinis viginti quinque milia; et erit sanctuarium Domini in medio eius.
EZEK|48|11|Sacerdotibus consecratis erit, filiis Sadoc, qui custodierunt caeremonias meas et non erraverunt, cum errarent filii Israel, sicut erraverunt Levitae.
EZEK|48|12|Et erit eis oblatio de oblatione terrae sanctum sanctorum iuxta terminum Levitarum;
EZEK|48|13|sed et Levitis similiter secundum fines sacerdotum, viginti quinque milia longitudinis et latitudinis decem milia, totum in longitudine viginti et quinque milia et in latitudine viginti milia;
EZEK|48|14|et non venumdabunt ex eo neque mutabunt, neque transferetur oblatio terrae, quia sanctificata est Domino.
EZEK|48|15|Quinque milia autem, quae supersunt in latitudine per viginti quinque milia, profana erunt urbi in habitaculum et in pascua, et erit civitas in medio eius.
EZEK|48|16|Et hae mensurae eius: ad plagam septentrionalem quingenti et quattuor milia et ad plagam meridianam quingenti et quattuor milia et ad plagam orientalem quingenti et quattuor milia et ad plagam occidentalem quingenti et quattuor milia.
EZEK|48|17|Erunt autem pascua civitatis ad aquilonem ducenti quinquaginta et ad meridiem ducenti quinquaginta et ad orientem ducenti quinquaginta et ad mare ducenti quinquaginta.
EZEK|48|18|Quod autem reliquum fuerit in longitudine iuxta oblationem sacram, decem milia ad orientem et decem milia ad occidentem, erunt iuxta oblationem sacram, et erunt fruges eius in panem his, qui serviunt civitati.
EZEK|48|19|Servientes autem civitati operabuntur ex omnibus tribubus Israel.
EZEK|48|20|Tota oblatio viginti quinque milium, per viginti quinque milia: in quadrum; separabitis oblationem sacram una cum possessione civitatis.
EZEK|48|21|Quod autem reliquum fuerit, principis erit, ex utraque parte oblationis sacrae et possessionis civitatis, e regione viginti quinque milium oblationis usque ad terminum orientalem, sed et ad mare e regione viginti quinque milium usque ad terminum maris secundum partes tribuum, principis erit. Et erit oblatio sacra et sanctuarium templi in medio eius,
EZEK|48|22|segregata a possessione Levitarum et a possessione civitatis in medio partium principis: inter terminum Iudae et inter terminum Beniamin erit possessio principis.
EZEK|48|23|Et reliquis tribubus: a plaga orientali usque ad plagam occidentalem, Beniamin una.
EZEK|48|24|Et iuxta terminum Beniamin a plaga orientali usque ad plagam occidentalem, Simeon una.
EZEK|48|25|Et iuxta terminum Simeonis a plaga orientali usque ad plagam occidentalem, Issachar una.
EZEK|48|26|Et iuxta terminum Issachar a plaga orientali usque ad plagam occidentalem, Zabulon una.
EZEK|48|27|Et iuxta terminum Zabulon a plaga orientali usque ad plagam maris, Gad una.
EZEK|48|28|Et iuxta terminum Gad ad plagam austri in meridiem, erit finis de Thamar usque ad aquas Meribathcades, ad torrentem usque ad mare Magnum.
EZEK|48|29|Haec est terra, quam mittetis in sortem tribubus Israel, et hae partitiones earum, ait Dominus Deus.
EZEK|48|30|Et hi egressus civitatis: a plaga septentrionali, cuius mensura quingenti et quattuor milia,
EZEK|48|31|portae civitatis in nominibus tribuum Israel: portae tres a septentrione, porta Ruben una, porta Iudae una, porta Levi una.
EZEK|48|32|Et ad plagam orientalem quingentorum et quattuor milium, portae tres: porta Ioseph una, porta Beniamin una, porta Dan una.
EZEK|48|33|Et ad plagam meridianam, cuius mensura quingenti et quattuor milia, portae tres: porta Simeonis una, porta Issachar una, porta Zabulon una.
EZEK|48|34|Et ad plagam occidentalem quingentorum et quattuor milium, portae tres: porta Gad una, porta Aser una, porta Nephthali una.
EZEK|48|35|Per circuitum decem et octo milia, et nomen civitatis ex illa die: Dominus ibidem ".
