PHLM|1|1|Павло, в'язень Христа Ісуса, та брат Тимофій, улюбленому Филимонові й співробітникові нашому,
PHLM|1|2|і сестрі любій Апфії, і співвойовникові нашому Архипові, і Церкві домашній твоїй:
PHLM|1|3|благодать вам і мир від Бога Отця нашого й Господа Ісуса Христа!
PHLM|1|4|Я завсіди дякую Богові моєму, коли тебе згадую в молитвах своїх.
PHLM|1|5|Бо я чув про любов твою й віру, яку маєш до Господа Ісуса, і до всіх святих,
PHLM|1|6|щоб спільність віри твоєї діяльна була в пізнанні всякого добра, що в нас для Христа.
PHLM|1|7|Бо ми маємо радість велику й потіху в любові твоїй, серця бо святих заспокоїв ти, брате.
PHLM|1|8|Через це, хоч я маю велику відвагу в Христі подавати накази тобі про потрібне,
PHLM|1|9|але більше з любови благаю я, як Павло, старий, тепер же ще й в'язень Христа Ісуса.
PHLM|1|10|Благаю тебе про сина свого, про Онисима, що його породив я в кайданах своїх.
PHLM|1|11|Колись то для тебе він був непотрібний, тепер же для тебе й для мене він дуже потрібний.
PHLM|1|12|Тобі я вертаю його, того, хто є неначе серце моє.
PHLM|1|13|Я хотів був тримати його при собі, щоб він замість тебе мені послужив у кайданах за Євангелію,
PHLM|1|14|та без волі твоєї нічого робити не хотів я, щоб твій добрий учинок не був ніби вимушений, але добровільний.
PHLM|1|15|Бо може для того він був розлучився на час, щоб навіки прийняв ти його,
PHLM|1|16|і вже не як раба, але вище від раба, як брата улюбленого, особливо для мене, а тим більше для тебе, і за тілом, і в Господі.
PHLM|1|17|Отож, коли маєш за друга мене, то прийми його, як мене.
PHLM|1|18|Коли ж він чим скривдив тебе або винен тобі, полічи це мені.
PHLM|1|19|Я, Павло, написав це рукою своєю: Я віддам, щоб тобі не казати, що ти навіть самого себе мені винен.
PHLM|1|20|Так, брате, нехай я одержу те, що від тебе прохаю в Господі. Заспокой моє серце в Христі!
PHLM|1|21|Пересвідчений я про слухняність твою, і тобі написав оце, відаючи, що ти зробиш і більше, ніж я говорю.
PHLM|1|22|А разом мені приготуй і помешкання, бо надіюся я, що за ваші молитви я буду дарований вам.
PHLM|1|23|Вітає тебе Епафрас, мій співв'язень у Христі Ісусі,
PHLM|1|24|Марко, Аристарх, Димас, Лука, мої співробітники.
PHLM|1|25|Благодать Господа Ісуса Христа з вашим духом! Амінь.
