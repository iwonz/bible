JUDE|1|1|Иуда, раб Иисуса Христа, брат Иакова, призванным, которые освящены Богом Отцем и сохранены Иисусом Христом:
JUDE|1|2|милость вам и мир и любовь да умножатся.
JUDE|1|3|Возлюбленные! имея все усердие писать вам об общем спасении, я почел за нужное написать вам увещание – подвизаться за веру, однажды преданную святым.
JUDE|1|4|Ибо вкрались некоторые люди, издревле предназначенные к сему осуждению, нечестивые, обращающие благодать Бога нашего в [повод к] распутству и отвергающиеся единого Владыки Бога и Господа нашего Иисуса Христа.
JUDE|1|5|Я хочу напомнить вам, уже знающим это, что Господь, избавив народ из земли Египетской, потом неверовавших погубил,
JUDE|1|6|и ангелов, не сохранивших своего достоинства, но оставивших свое жилище, соблюдает в вечных узах, под мраком, на суд великого дня.
JUDE|1|7|Как Содом и Гоморра и окрестные города, подобно им блудодействовавшие и ходившие за иною плотию, подвергшись казни огня вечного, поставлены в пример, –
JUDE|1|8|так точно будет и с сими мечтателями, которые оскверняют плоть, отвергают начальства и злословят высокие власти.
JUDE|1|9|Михаил Архангел, когда говорил с диаволом, споря о Моисеевом теле, не смел произнести укоризненного суда, но сказал: "да запретит тебе Господь".
JUDE|1|10|А сии злословят то, чего не знают; что же по природе, как бессловесные животные, знают, тем растлевают себя.
JUDE|1|11|Горе им, потому что идут путем Каиновым, предаются обольщению мзды, как Валаам, и в упорстве погибают, как Корей.
JUDE|1|12|Таковые бывают соблазном на ваших вечерях любви; пиршествуя с вами, без страха утучняют себя. Это безводные облака, носимые ветром; осенние деревья, бесплодные, дважды умершие, исторгнутые;
JUDE|1|13|свирепые морские волны, пенящиеся срамотами своими; звезды блуждающие, которым блюдется мрак тьмы на веки.
JUDE|1|14|О них пророчествовал и Енох, седьмый от Адама, говоря: "се, идет Господь со тьмами святых Ангелов Своих –
JUDE|1|15|сотворить суд над всеми и обличить всех между ними нечестивых во всех делах, которые произвело их нечестие, и во всех жестоких словах, которые произносили на Него нечестивые грешники".
JUDE|1|16|Это ропотники, ничем не довольные, поступающие по своим похотям (нечестиво и беззаконно); уста их произносят надутые слова; они оказывают лицеприятие для корысти.
JUDE|1|17|Но вы, возлюбленные, помните предсказанное Апостолами Господа нашего Иисуса Христа.
JUDE|1|18|Они говорили вам, что в последнее время появятся ругатели, поступающие по своим нечестивым похотям.
JUDE|1|19|Это люди, отделяющие себя (от единства веры), душевные, не имеющие духа.
JUDE|1|20|А вы, возлюбленные, назидая себя на святейшей вере вашей, молясь Духом Святым,
JUDE|1|21|сохраняйте себя в любви Божией, ожидая милости от Господа нашего Иисуса Христа, для вечной жизни.
JUDE|1|22|И к одним будьте милостивы, с рассмотрением,
JUDE|1|23|а других страхом спасайте, исторгая из огня, обличайте же со страхом, гнушаясь даже одеждою, которая осквернена плотью.
JUDE|1|24|Могущему же соблюсти вас от падения и поставить пред славою Своею непорочными в радости,
JUDE|1|25|Единому Премудрому Богу, Спасителю нашему чрез Иисуса Христа Господа нашего, слава и величие, сила и власть прежде всех веков, ныне и во все веки. Аминь.
