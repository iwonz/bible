MIC|1|1|當 猶大 王 約坦 、 亞哈斯 、 希西家 在位的時候，耶和華的話臨到 摩利沙 人 彌迦 ，他見到有關 撒瑪利亞 和 耶路撒冷 的異象。
MIC|1|2|萬民哪，你們都要聽！ 地和其上所有的，要留心聽！ 主耶和華要從他的聖殿 指證你們的不是。
MIC|1|3|看哪，耶和華從他的居所出來， 降臨步行地之高處。
MIC|1|4|眾山在他底下熔化， 諸谷崩裂， 如蠟熔在火中， 如水沖下山坡。
MIC|1|5|這都是因 雅各 的罪過， 因 以色列 家的罪惡。 雅各 的罪過在哪裏呢？ 豈不是在 撒瑪利亞 嗎？ 猶大 的丘壇在哪裏呢？ 豈不是在 耶路撒冷 嗎？
MIC|1|6|因此，我必使 撒瑪利亞 變為田野的廢墟， 用以栽植葡萄； 我必把它的石頭倒在山谷， 掀開它的地基。
MIC|1|7|城裏一切雕刻的偶像必被打碎， 行淫的賞金全被火燒， 我要毀滅它的一切偶像； 因為從妓女的賞金積聚而來的， 它們仍歸為妓女的賞金。
MIC|1|8|為此我要大聲哀號， 赤身赤腳行走； 我要呼號如野狗， 哀鳴如鴕鳥。
MIC|1|9|因為 撒瑪利亞 的創傷無法醫治， 蔓延到 猶大 ， 到了我百姓的城門， 直達 耶路撒冷 。
MIC|1|10|不要在 迦特 宣揚 這事， 千萬不要哭泣； 要在 伯‧亞弗拉 翻滾於灰塵 中。
MIC|1|11|沙斐 的居民哪，要赤身羞愧地經過， 撒南 的居民不敢出門， 伯‧以薛 哀哭，不再支持你們。
MIC|1|12|瑪律 的居民心甚憂急，切望得著福氣， 因為災禍已從耶和華那裏臨到 耶路撒冷 的城門。
MIC|1|13|拉吉 的居民哪，要用快馬 套車； 錫安 的罪由你而起， 以色列 的罪過在你那裏顯出。
MIC|1|14|因此，你要將送別禮送到 摩利設‧迦特 ； 亞革悉 的眾家族必用詭詐 待 以色列 諸王。
MIC|1|15|瑪利沙 的居民哪， 我必使搶奪者來到你這裏； 以色列 的貴族 必來到 亞杜蘭 。
MIC|1|16|猶大 啊，為了你所喜愛的兒女， 你要剪髮，剃光頭， 要使你的頭光禿，如同禿鷹， 因為他們被擄去離開你了。
MIC|2|1|禍哉，那些在床上圖謀罪孽、籌劃惡事的人！ 天一亮，他們因手中有能力就去行惡。
MIC|2|2|他們看上田地就佔據， 貪圖房屋便奪取； 他們欺壓戶主和他的家庭， 霸佔人和他的產業。
MIC|2|3|所以耶和華如此說： 看哪，我籌劃災禍降與這家族； 這災禍在你們頸項上無法解脫， 你們也不能昂首而行， 因為這是災禍的時刻。
MIC|2|4|到那日，必有人為你們唱詩歌， 用悲哀的哀歌哀號，說： 「我們全然敗落， 我百姓的產業易主了！ 耶和華竟然使它離開我， 我們的田地為悖逆的人所瓜分了！」
MIC|2|5|因此，你必無人能在耶和華的會中 抽籤拉繩 。
MIC|2|6|他們傳講說：「不可傳講； 人都不可傳講這些事， 羞辱不會臨到我們。」
MIC|2|7|雅各 家啊，可這麼說嗎 ？ 耶和華沒有耐心嗎？ 這些事是他所行的嗎？ 我的言語豈不是與行動正直的人有益嗎？
MIC|2|8|然而，近來我的百姓興起如仇敵。 你們剝去那些安然行路、不願打仗之人身上的外衣，
MIC|2|9|把我百姓中的婦人從安樂家中趕出， 又將我的榮耀從她們孩子身上永遠奪去。
MIC|2|10|起來，走吧！ 這裏並非安歇之處； 因為不潔淨帶來毀壞， 且是大大的毀壞。
MIC|2|11|若有人心存虛假，用謊言說 ： 「我向你們傳講可得清酒和烈酒 」， 那人就必作這百姓的傳講者。
MIC|2|12|雅各 家啊，我定要聚集你們， 定要召集 以色列 的餘民， 把他們安置在一處，如 波斯拉 的羊， 又如草場上的羊群， 人數眾多，大大喧嘩。
MIC|2|13|開路的在他們前面上去， 直闖過城門，從城門出去； 他們的王在前面行， 耶和華在他們的前頭。
MIC|3|1|於是我說： 雅各 的領袖， 以色列 家的官長啊， 你們要聽！ 你們豈不知道公平嗎？
MIC|3|2|你們惡善好惡， 剝我百姓 身上的皮， 從他們的骨頭上剔肉，
MIC|3|3|你們吃我百姓的肉， 剝他們的皮， 打斷他們的骨頭， 如切塊 下鍋， 如釜中的肉。
MIC|3|4|到了遭災的時候，這些人要哀求耶和華， 他卻不應允他們。 那時，因他們所行的惡， 他必轉臉離開他們。
MIC|3|5|論到使我百姓走入歧途的先知， 他們牙齒有所嚼，就呼喊說：「平安！」 誰不給他們吃，就揚言攻擊他， 耶和華如此說：
MIC|3|6|你們因此必遭遇黑夜，看不到異象； 遭遇幽暗，無法占卜。 太陽必向先知沉落， 白晝轉為黑暗。
MIC|3|7|先見必抱愧， 占卜的必蒙羞， 他們全都摀著鬍鬚， 因為上帝不應允他們。
MIC|3|8|至於我，我藉耶和華的靈， 滿有能力、公平和勇氣， 可向 雅各 述說他的過犯， 向 以色列 指出他的罪惡。
MIC|3|9|當聽這話， 雅各 家的領袖， 以色列 家的官長啊！ 你們厭棄公平， 在一切事上屈枉正直；
MIC|3|10|以血建立 錫安 ， 以罪孽建造 耶路撒冷 。
MIC|3|11|城裏的領袖為賄賂行審判， 祭司為酬勞施訓誨， 先知為銀錢行占卜； 他們卻倚賴耶和華，說： 「耶和華不是在我們中間嗎？ 災禍必不臨到我們。」
MIC|3|12|因此，為你們的緣故， 錫安 要被耕種像一塊田地， 耶路撒冷 要變為廢墟， 這殿的山必如叢林的高處。
MIC|4|1|末後的日子， 耶和華殿的山必堅立， 超乎諸山，高舉過於萬嶺； 萬民都要流歸這山。
MIC|4|2|必有許多民族前往，說： 「來吧，我們登耶和華的山， 到 雅各 上帝的殿。 他必將他的道指教我們， 我們也要行他的路。」 因為教誨必出於 錫安 ， 耶和華的言語必出於 耶路撒冷 。
MIC|4|3|他必在許多民族中施行審判， 為遠方強盛的國斷定是非。 他們要將刀打成犁頭， 把槍打成鐮刀。 這國不舉刀攻擊那國， 他們也不再學習戰事。
MIC|4|4|人人都要坐在自己的葡萄樹 和無花果樹下， 無人使他們驚嚇； 這是萬軍之耶和華親口說的。
MIC|4|5|萬民都奉自己神明的名行事， 我們卻要奉耶和華－我們上帝的名而行， 直到永永遠遠。
MIC|4|6|耶和華說：在那日， 我必聚集瘸腿的， 召集被趕逐的， 以及我所懲治的人。
MIC|4|7|我要使瘸腿的成為餘民， 使被趕到遠方的成為強盛之國。 耶和華要在 錫安山 作王治理他們， 從今直到永遠。
MIC|4|8|你， 以得臺 ， 錫安 的山岡啊， 先前的權柄必歸給你， 耶路撒冷 的國權必將歸還。
MIC|4|9|現在，你為何大聲呼喊呢？ 你中間沒有君王， 你的謀士滅絕， 以致疼痛抓住你， 如臨產的婦人嗎？
MIC|4|10|錫安 哪，你要疼痛生產， 彷彿臨產的婦人； 因你必從城裏出來，住在田野； 你要到 巴比倫 去， 在那裏，你要蒙解救， 在那裏，耶和華必救贖你 脫離仇敵的手掌。
MIC|4|11|現在，許多國家聚集攻擊你，說： 「讓 錫安 被玷污！ 讓我們親眼看到！」
MIC|4|12|他們卻不知道耶和華的意念， 也不明白他的籌算， 他聚集他們， 像把禾捆聚到禾場。
MIC|4|13|錫安 哪，起來踹穀吧！ 我必使你的角成為鐵， 使你的蹄成為銅。 你必打碎許多民族， 將他們的財寶獻給耶和華， 將他們的財富獻給全地的主。
MIC|5|1|成群的民 哪，現在要聚集成隊； 仇敵前來圍攻我們， 要用杖擊打 以色列 領袖的臉頰。
MIC|5|2|伯利恆 的 以法他 啊， 你在 猶大 諸城中雖小， 將來必有一位從你那裏出來， 在 以色列 中為我作掌權者； 他的根源自亙古，從太初就有。
MIC|5|3|因此，耶和華要將 以色列 人交給敵人， 直到臨產的婦人生下孩子； 那時，他其餘的弟兄 必回到 以色列 人那裏。
MIC|5|4|他必倚靠耶和華的大能， 倚靠耶和華－他上帝之名的威嚴， 站立並牧養， 使他們安然居住； 因為現在他必尊大， 直到地極。
MIC|5|5|這位就是和平 。 當 亞述 侵入我們領土， 踐踏我們宮殿時， 我們就立七個牧者， 八個領袖攻擊它。
MIC|5|6|他們要用刀劍毀壞 亞述 地 和 寧錄 地的關口 。 當 亞述 侵入我們領土， 踐踏我們邊境時， 他必拯救我們。
MIC|5|7|雅各 的餘民 必在許多民族中， 如從耶和華降下的露水， 又如甘霖降在草上； 他們不倚靠人， 也不仰賴世人。
MIC|5|8|雅各 的餘民必在列國中， 在許多民族中， 如林間百獸中的獅子， 又如少壯獅子在羊群中； 他若經過就必踐踏撕裂， 無人搭救。
MIC|5|9|願你的手舉起，高過敵人！ 願你的仇敵都被剪除！
MIC|5|10|耶和華說：到那日， 我必從你中間剪除馬匹， 毀壞戰車；
MIC|5|11|除滅你國中的城鎮， 拆毀你一切的堡壘；
MIC|5|12|除掉你手中的邪術， 你那裏不再有占卜的人。
MIC|5|13|我必從你中間除滅雕刻的偶像和柱像， 你就不再跪拜自己手所造的；
MIC|5|14|我必從你中間拔除 亞舍拉 ， 毀滅你的城鎮；
MIC|5|15|我必在怒氣和憤怒中 報應那不聽從我的列國。
MIC|6|1|當聽耶和華說的話： 起來，向山嶺爭辯， 使岡陵聽見你的聲音。
MIC|6|2|山嶺啊，要聽耶和華的指控！ 大地永久的根基啊，要聽！ 因耶和華控告他的百姓， 與 以色列 爭辯。
MIC|6|3|「我的百姓啊，我向你做了甚麼呢？ 我在甚麼事上使你厭煩？ 你回答我吧！
MIC|6|4|我曾將你從 埃及 地領出來， 從為奴之家救贖你， 我差遣 摩西 、 亞倫 和 米利暗 在你前面帶領。
MIC|6|5|我的百姓啊，當記念從前 摩押 王 巴勒 如何籌算， 比珥 的兒子 巴蘭 如何回應他， 當記念從 什亭 到 吉甲 所發生的事， 好使你們明白耶和華公義的作為。」
MIC|6|6|「我朝見耶和華， 在至高上帝面前跪拜，當獻上甚麼呢？ 難道獻一歲的牛犢為燔祭來朝見他嗎？
MIC|6|7|耶和華豈喜悅千千的公羊， 或是萬萬的油河嗎？ 我豈可為自己的過犯獻我的長子， 為自己的罪惡獻我所親生的嗎？」
MIC|6|8|世人哪，耶和華已指示你何為善。 他向你所要的是甚麼呢？ 只要你行公義，好憐憫， 存謙卑的心與你的上帝同行。
MIC|6|9|耶和華向這城呼叫 ─看重你的名是真智慧 ─ 你們當聽懲罰 和派定懲罰的人 。
MIC|6|10|惡人家中不是仍有不義之財 和惹人生氣的變小了的伊法嗎？
MIC|6|11|我若用不公道的天平 和袋中詭詐的法碼， 豈可算為清白呢？
MIC|6|12|城裏的有錢人遍行殘暴， 其中的居民說謊話， 口中的舌頭盡是詭詐。
MIC|6|13|因此，我也擊打你，使你受傷 ， 因你的罪惡使你受驚駭。
MIC|6|14|你要吃，卻吃不飽， 你的肚子仍是空空。 你必被挪去，不得逃脫； 如有逃脫的，我必交給刀劍。
MIC|6|15|你撒種，卻不得收割； 踹橄欖，卻不得油抹身； 有新酒，卻不得酒喝。
MIC|6|16|因為你遵守 暗利 的規條， 行 亞哈 家一切所行的， 順從他們的計謀； 因此，我必使你荒涼， 使你的居民遭人嗤笑， 你們也必擔當我百姓的羞辱。
MIC|7|1|我有禍了！我好像夏日收割後的果子， 又如收成之後剩餘的葡萄， 沒有一掛可吃的， 也沒有我心所渴想初熟的無花果。
MIC|7|2|地上的虔誠人滅盡了， 人世間已無正直的人； 他們都埋伏，為要流人的血， 用羅網獵取自己的弟兄。
MIC|7|3|他們雙手善於作惡， 君王和審判官都索取賄賂； 位高的人吐出心中的慾望， 彼此勾結 。
MIC|7|4|他們當中最好的，不過像蒺藜； 最正直的，不過如荊棘籬笆。 你守候的日子，懲罰已經來到， 他們必擾亂不安。
MIC|7|5|不可倚賴鄰舍， 不可信靠密友； 甚至對躺在你懷中的妻子 也要守住你的口。
MIC|7|6|因為兒子藐視父親， 女兒抵擋母親， 媳婦抗拒婆婆， 人的仇敵就是自己家裏的人。
MIC|7|7|至於我，我要仰望耶和華， 等候那救我的上帝； 我的上帝必應允我。
MIC|7|8|我的仇敵啊，不要向我誇耀。 我雖跌倒，仍要起來； 雖坐在黑暗裏，耶和華卻作我的光。
MIC|7|9|我要承受耶和華的惱怒， 直到他為我辯護，為我伸冤， 因我得罪了他； 他要領我進入光明， 我必得見他的公義。
MIC|7|10|那時我的仇敵看見這事就羞愧， 他曾對我說：「耶和華－你的上帝在哪裏？」 我必親眼見他遭報， 現在，他必被踐踏，如同街上的泥土。
MIC|7|11|你的城牆重修的日子到了！ 到那日，邊界必擴展。
MIC|7|12|到那日，人必從 亞述 ， 從 埃及 的城鎮， 從 埃及 到 大河 ， 從這海到那海， 從這山到那山， 都歸到你這裏。
MIC|7|13|然而，因居民的緣故， 為了他們行事的結果， 這地必然荒涼。
MIC|7|14|求你在 迦密 的樹林中， 以你的杖牧放你獨居的民， 你產業中的羊群； 願他們像古時一樣， 牧放在 巴珊 和 基列 。
MIC|7|15|我要顯奇事給他們看， 好像出 埃及 地的時候一樣。
MIC|7|16|列國看見，雖大有勢力仍覺慚愧； 他們必用手摀口，掩耳不聽。
MIC|7|17|他們要舔土如蛇， 又如地上爬行的動物， 戰戰兢兢離開他們的營寨； 他們必畏懼耶和華─我們的上帝， 也必因你而害怕。
MIC|7|18|有哪一個神明像你，赦免罪孽， 饒恕他產業中餘民的罪過？ 他不永遠懷怒，喜愛施恩。
MIC|7|19|他 必轉回憐憫我們， 把我們的罪孽踏在腳下。 你必將他們 一切的罪投於深海。
MIC|7|20|你必按古時向我們列祖起誓的話， 以信實待 雅各 ， 向 亞伯拉罕 施慈愛。
