ROM|1|1|Павло, раб Ісуса Христа, покликаний апостол, вибраний для звіщання Євангелії Божої,
ROM|1|2|яке Він перед тим приобіцяв через Своїх пророків у святих Писаннях,
ROM|1|3|про Сина Свого, що тілом був із насіння Давидового,
ROM|1|4|і об'явився Сином Божим у силі, за духом святости, через воскресення з мертвих, про Ісуса Христа, Господа нашого,
ROM|1|5|що через Нього прийняли ми благодать і апостольство на послух віри через Ім'я Його між усіма народами,
ROM|1|6|між якими й ви, покликані Ісуса Христа,
ROM|1|7|усім, хто знаходиться в Римі, улюбленим Божим, вибраним святим, благодать вам та мир від Бога, Отця нашого, і Господа Ісуса Христа!
ROM|1|8|Отже, насамперед дякую Богові моєму через Ісуса Христа за всіх вас, що віра ваша звіщається по всьому світові.
ROM|1|9|Бо свідок мені Бог, Якому служу духом своїм у звіщанні Євангелії Його Сина, що я безперестанно згадую про вас,
ROM|1|10|і в молитвах своїх завжди молюся, щоб воля Божа щасливо попровадила мене коли прийти до вас.
ROM|1|11|Бо прагну вас бачити, щоб подати вам якого дара духовного для зміцнення вас,
ROM|1|12|цебто потішитись разом між вами спільною вірою і вашою, і моєю.
ROM|1|13|Не хочу ж, щоб ви не знали, браття, що багато разів мав я замір прийти до вас, але мені перешкоджувано аж досі, щоб мати який плід і в вас, як і в інших народів.
ROM|1|14|А гелленам і чужоземцям, розумним і немудрим я боржник.
ROM|1|15|Отже, щодо мене, я готовий і вам, хто знаходиться в Римі, звіщати Євангелію.
ROM|1|16|Бо я не соромлюсь Євангелії, бож вона сила Божа на спасіння кожному, хто вірує, перше ж юдеєві, а потім гелленові.
ROM|1|17|Правда бо Божа з'являється в ній з віри в віру, як написано: А праведний житиме вірою.
ROM|1|18|Бо гнів Божий з'являється з неба на всяку безбожність і неправду людей, що правду гамують неправдою,
ROM|1|19|тому, що те, що можна знати про Бога, явне для них, бо їм Бог об'явив.
ROM|1|20|Бо Його невидиме від створення світу, власне Його вічна сила й Божество, думанням про твори стає видиме. Так що нема їм виправдання,
ROM|1|21|бо, пізнавши Бога, не прославляли Його, як Бога, і не дякували, але знікчемніли своїми думками, і запаморочилось нерозумне їхнє серце.
ROM|1|22|Називаючи себе мудрими, вони потуманіли,
ROM|1|23|і славу нетлінного Бога змінили на подобу образа тлінної людини, і птахів, і чотириногих, і гадів.
ROM|1|24|Тому то й видав їх Бог у пожадливостях їхніх сердець на нечистість, щоб вони самі знеславляли тіла свої.
ROM|1|25|Вони Божу правду замінили на неправду, і честь віддавали, і служили створінню більш, як Творцеві, що благословенний навіки, амінь.
ROM|1|26|Через це Бог їх видав на пожадливість ганебну, бо їхні жінки замінили природне єднання на протиприродне.
ROM|1|27|Так само й чоловіки, позоставивши природне єднання з жіночою статтю, розпалилися своєю пожадливістю один до одного, і чоловіки з чоловіками сором чинили. І вони прийняли в собі відплату, відповідну їхньому блудові.
ROM|1|28|А що вони не вважали за потрібне мати Бога в пізнанні, видав їх Бог на розум перевернений, щоб чинили непристойне.
ROM|1|29|Вони повні всякої неправди, лукавства, зажерливости, злоби, повні заздрости, убивства, суперечки, омани, лихих звичаїв,
ROM|1|30|обмовники, наклепники, богоненавидники, напасники, чваньки, пишні, винахідники зла, неслухняні батькам,
ROM|1|31|нерозумні, зрадники, нелюбовні, немилостиві.
ROM|1|32|Вони знають присуд Божий, що ті, хто чинить таке, варті смерти, а проте не тільки самі чинять, але й хвалять тих, хто робить таке.
ROM|2|1|Ось тому без виправдання ти, кожний чоловіче, що судиш, бо в чому осуджуєш іншого, сам себе осуджуєш, бо чиниш те саме й ти, що судиш.
ROM|2|2|А ми знаємо, що суд Божий поправді на тих, хто чинить таке.
ROM|2|3|Чи ти думаєш, чоловіче, судячи тих, хто чинить таке, а сам робиш таке саме, що ти втечеш від суду Божого?
ROM|2|4|Або погорджуєш багатством Його добрости, лагідности та довготерпіння, не знаючи, що Божа добрість провадить тебе до покаяння?
ROM|2|5|Та через жорстокість свою й нерозкаяність серця збираєш собі гнів на день гніву та об'явлення справедливого суду Бога,
ROM|2|6|що кожному віддасть за його вчинками:
ROM|2|7|тим, хто витривалістю в добрім ділі шукає слави, і чести, і нетління, життя вічне,
ROM|2|8|а сварливим та тим, хто противиться правді, але кориться неправді, лютість та гнів.
ROM|2|9|Недоля та утиск на всяку душу людини, хто чинить зле, юдея ж перше та геллена,
ROM|2|10|а слава, і честь, і мир усякому, хто чинить добре, юдеєві ж перше та гелленові.
ROM|2|11|Бо не дивиться Бог на обличчя!
ROM|2|12|Котрі бо згрішили без Закону, без Закону й загинуть, а котрі згрішили в Законі, приймуть суд за Законом.
ROM|2|13|Бо не слухачі Закону справедливі перед Богом, але виконавці Закону виправдані будуть.
ROM|2|14|Бо коли погани, що не мають Закону, з природи чинять законне, вони, не мавши Закону, самі собі Закон,
ROM|2|15|що виявляють діло Закону, написане в серцях своїх, як свідчить їм сумління та їхні думки, що то осуджують, то виправдують одна одну,
ROM|2|16|дня, коли Бог, згідно з моїм благовістям, буде судити таємні речі людей через Ісуса Христа.
ROM|2|17|Ось ти звешся юдеєм, і спираєшся на Закона, і хвалишся Богом,
ROM|2|18|і знаєш волю Його, і розумієш, що краще, навчившись із Закону,
ROM|2|19|і маєш певність, що ти провідник для сліпих, світло для тих, хто знаходиться в темряві,
ROM|2|20|виховник нерозумним, учитель дітям, що ти маєш зразок знання й правди в Законі.
ROM|2|21|Отож, ти, що іншого навчаєш, себе самого не вчиш! Проповідуєш не красти, а сам крадеш!
ROM|2|22|Наказуючи не чинити перелюбу, чиниш перелюб! Гидуючи ідолами, чиниш святокрадство!
ROM|2|23|Ти, що хвалишся Законом, зневажаєш Бога переступом Закону!
ROM|2|24|Бо через вас зневажається Боже Ймення в поган, як написано.
ROM|2|25|Обрізання корисне, коли виконуєш Закона; а коли ти переступник Закону, то обрізання твоє стало необрізанням.
ROM|2|26|Отож, коли необрізаний зберігає постанови Закону, то чи не порахується його необрізання за обрізання?
ROM|2|27|І необрізаний з природи, виконуючи Закона, чи не осудить тебе, переступника Закону з Писанням і обрізанням?
ROM|2|28|Бо не той юдей, що є ним назовні, і не то обрізання, що назовні на тілі,
ROM|2|29|але той, що є юдей потаємно, духово, і обрізання серця духом, а не за буквою; і йому похвала не від людей, а від Бога.
ROM|3|1|Отож, що має більшого юдей, або яка користь від обрізання?
ROM|3|2|Багато, на всякий спосіб, а насамперед, що їм довірені були Слова Божі.
ROM|3|3|Бо що ж, що не вірували деякі? Чи ж їхнє недовірство знищить вірність Божу?
ROM|3|4|Зовсім ні! Бож Бог правдивий, а кожна людина неправдива, як написано: Щоб був Ти виправданий у словах Своїх, і переміг, коли будеш судитися.
ROM|3|5|А коли наша неправда виставляє правду Божу, то що скажемо? Чи ж Бог несправедливий, коли гнів виявляє? Говорю по-людському.
ROM|3|6|Зовсім ні! Бож як Бог судитиме світ?
ROM|3|7|Бо коли Божа правда через мою неправду збільшилась на славу Йому, пощо судити ще й мене, як грішника?
ROM|3|8|І чи не так, як нас лають, і як деякі говорять, ніби ми кажемо: Робімо зле, щоб вийшло добре? Справедливий осуд на таких!
ROM|3|9|То що ж? Маємо перевагу? Анітрохи! Бож ми перед тим довели, що юдеї й геллени усі під гріхом,
ROM|3|10|як написано: Нема праведного ані одного;
ROM|3|11|нема, хто розумів би; немає, хто Бога шукав би,
ROM|3|12|усі повідступали, разом стали непотрібні, нема доброчинця, нема ні одного!
ROM|3|13|Гріб відкритий їхнє горло, язиком своїм кажуть неправду, отрута зміїна на їхніх губах,
ROM|3|14|уста їхні повні прокляття й гіркоти!
ROM|3|15|Швидкі їхні ноги, щоб кров проливати,
ROM|3|16|руїна та злидні на їхніх дорогах,
ROM|3|17|а дороги миру вони не пізнали!
ROM|3|18|Нема страху Божого перед очима їхніми...
ROM|3|19|А ми знаємо, що скільки говорить Закон, він говорить до тих, хто під Законом, щоб замкнути всякі уста, і щоб став увесь світ винний Богові.
ROM|3|20|Бо жадне тіло ділами Закону не виправдається перед Ним, Законом бо гріх пізнається.
ROM|3|21|А тепер, без Закону, правда Божа з'явилась, про яку свідчать Закон і Пророки.
ROM|3|22|А Божа правда через віру в Ісуса Христа в усіх і на всіх, хто вірує, бо різниці немає,
ROM|3|23|бо всі згрішили, і позбавлені Божої слави,
ROM|3|24|але дарма виправдуються Його благодаттю, через відкуплення, що в Ісусі Христі,
ROM|3|25|що Його Бог дав у жертву примирення в крові Його через віру, щоб виявити Свою правду через відпущення давніше вчинених гріхів,
ROM|3|26|за довготерпіння Божого, щоб виявити Свою правду за теперішнього часу, щоб бути Йому праведним, і виправдувати того, хто вірує в Ісуса.
ROM|3|27|Тож де похвальба? Виключена. Яким законом? Законом діл? Ні, але законом віри.
ROM|3|28|Отож, ми визнаємо, що людина виправдується вірою, без діл Закону.
ROM|3|29|Хіба ж Бог тільки для юдеїв, а не й для поган? Так, і для поган,
ROM|3|30|бо є один тільки Бог, що виправдає обрізання з віри й необрізання через віру.
ROM|3|31|Тож чи не нищимо ми Закона вірою? Зовсім ні, але зміцнюємо Закона.
ROM|4|1|Що ж, скажемо, знайшов Авраам, наш отець за тілом?
ROM|4|2|Бо коли Авраам виправдався ділами, то він має похвалу, та не в Бога.
ROM|4|3|Що бо Писання говорить? Увірував Авраам Богові, і це йому залічено в праведність.
ROM|4|4|А заплата виконавцеві не рахується з милости, але з обов'язку.
ROM|4|5|А тому, хто не виконує, але вірує в Того, Хто виправдує нечестивого, віра його порахується в праведність.
ROM|4|6|Як і Давид називає блаженною людину, якій рахує Бог праведність без діл:
ROM|4|7|Блаженні, кому прощені беззаконня, і кому прикриті гріхи.
ROM|4|8|Блаженна людина, якій Господь не порахує гріха!
ROM|4|9|Чи ж це блаженство з обрізання чи з необрізання? Бо говоримо, що віра залічена Авраамові в праведність.
ROM|4|10|Як же залічена? Як був в обрізанні, чи в необрізанні? Не в обрізанні, але в необрізанні!
ROM|4|11|І прийняв він ознаку обрізання, печать праведности через віру, що її в необрізанні мав, щоб йому бути отцем усіх віруючих, хоч були необрізані, щоб і їм залічено праведність,
ROM|4|12|і отцем обрізаних, не тільки тих, хто з обрізання, але й тих, хто ходить по слідах віри, що її в необрізанні мав наш отець Авраам.
ROM|4|13|Бо обітницю Авраамові чи його насінню, що бути йому спадкоємцем світу, дано не Законом, але праведністю віри.
ROM|4|14|Бо коли спадкоємці ті, хто з Закону, то спорожніла віра й знівечилась обітниця.
ROM|4|15|Бо Закон чинить гнів; де ж немає Закону, немає й переступу.
ROM|4|16|Через це з віри, щоб було з милости, щоб обітниця певна була всім нащадкам, не тільки тому, хто з Закону, але й тому, хто з віри Авраама, що отець усім нам,
ROM|4|17|як написано: Отцем багатьох народів Я поставив тебе, перед Богом, Якому він вірив, Який оживляє мертвих і кличе неіснуюче, як існуюче.
ROM|4|18|Він проти надії увірував у надії, що стане батьком багатьох народів, за сказаним: Таке численне буде насіння твоє!
ROM|4|19|І не знеміг він у вірі, і не вважав свого тіла за вже омертвіле, бувши майже сторічним, ні утроби Сариної за змертвілу,
ROM|4|20|і не мав сумніву в обітницю Божу через недовірство, але зміцнився в вірі, і віддав славу Богові,
ROM|4|21|і був зовсім певний, що Він має силу й виконати те, що обіцяв.
ROM|4|22|Тому й залічено це йому в праведність.
ROM|4|23|Та не написано за нього одного, що залічено йому,
ROM|4|24|а за нас, залічиться й нам, що віруємо в Того, Хто воскресив із мертвих Ісуса, Господа нашого,
ROM|4|25|що був виданий за наші гріхи, і воскрес для виправдання нашого.
ROM|5|1|Отож, виправдавшись вірою, майте мир із Богом через Господа нашого Ісуса Христа,
ROM|5|2|через Якого ми вірою одержали доступ до тієї благодаті, що в ній стоїмо, і хвалимось надією слави Божої.
ROM|5|3|І не тільки нею, але й хвалимося в утисках, знаючи, що утиски приносять терпеливість,
ROM|5|4|а терпеливість досвід, а досвід надію,
ROM|5|5|а надія не засоромить, бо любов Божа вилилася в наші серця Святим Духом, даним нам.
ROM|5|6|Бо Христос, коли ми були ще недужі, своєї пори помер за нечестивих.
ROM|5|7|Бо навряд чи помре хто за праведника, ще бо за доброго може хто й відважиться вмерти.
ROM|5|8|А Бог доводить Свою любов до нас тим, що Христос умер за нас, коли ми були ще грішниками.
ROM|5|9|Тож тим більше спасемося Ним від гніву тепер, коли кров'ю Його ми виправдані.
ROM|5|10|Бо коли ми, бувши ворогами, примирилися з Богом через смерть Сина Його, то тим більше, примирившися, спасемося життям Його.
ROM|5|11|І не тільки це, але й хвалимося в Бозі через Господа нашого Ісуса Христа, що через Нього одержали ми тепер примирення.
ROM|5|12|Тому то, як через одного чоловіка ввійшов до світу гріх, а гріхом смерть, так прийшла й смерть у всіх людей через те, що всі згрішили.
ROM|5|13|Гріх бо був у світі й до Закону, але гріх не ставиться в провину, коли немає Закону.
ROM|5|14|Та смерть панувала від Адама аж до Мойсея і над тими, хто не згрішив, подібно переступу Адама, який є образ майбутнього.
ROM|5|15|Але не такий дар благодаті, як переступ. Бо коли за переступ одного померло багато, то тим більш благодать Божа й дар через благодать однієї Людини, Ісуса Христа, щедро спливли на багатьох.
ROM|5|16|І дар не такий, як те, що сталось від одного, що згрішив; бо суд за один прогріх на осуд, а дар благодаті на виправдання від багатьох прогріхів.
ROM|5|17|Бо коли за переступ одного смерть панувала через одного, то тим більше ті, хто приймає рясноту благодаті й дар праведности, запанують у житті через одного Ісуса Христа.
ROM|5|18|Ось тому, як через переступ одного на всіх людей прийшов осуд, так і через праведність Одного прийшло виправдання для життя на всіх людей.
ROM|5|19|Бо як через непослух одного чоловіка багато-хто стали грішними, так і через послух Одного багато-хто стануть праведними.
ROM|5|20|Закон же прийшов, щоб збільшився переступ. А де збільшився гріх, там зарясніла благодать,
ROM|5|21|щоб, як гріх панував через смерть, так само й благодать запанувала через праведність для життя вічного Ісусом Христом, Господом нашим.
ROM|6|1|Що ж скажемо? Позостанемся в гріху, щоб благодать примножилась? Зовсім ні!
ROM|6|2|Ми, що вмерли для гріха, як ще будемо жити в нім?
ROM|6|3|Чи ви не знаєте, що ми всі, хто христився у Христа Ісуса, у смерть Його христилися?
ROM|6|4|Отож, ми поховані з Ним хрищенням у смерть, щоб, як воскрес Христос із мертвих славою Отця, так щоб і ми стали ходити в обновленні життя.
ROM|6|5|Бо коли ми з'єдналися подобою смерти Його, то з'єднаємось і подобою воскресення,
ROM|6|6|знаючи те, що наш давній чоловік розп'ятий із Ним, щоб знищилось тіло гріховне, щоб не бути нам більше рабами гріха,
ROM|6|7|бо хто вмер, той звільнивсь від гріха!
ROM|6|8|А коли ми померли з Христом, то віруємо, що й жити з Ним будемо,
ROM|6|9|знаючи, що Христос, воскреснувши з мертвих, уже більш не вмирає, смерть над Ним не панує вже більше!
ROM|6|10|Бо що вмер Він, то один раз умер для гріха, а що живе, то для Бога живе.
ROM|6|11|Так само ж і ви вважайте себе за мертвих для гріха й за живих для Бога в Христі Ісусі, Господі нашім.
ROM|6|12|Тож нехай не панує гріх у смертельному вашому тілі, щоб вам слухатись його пожадливостей,
ROM|6|13|і не віддавайте членів своїх гріхові за знаряддя неправедности, але віддавайте себе Богові, як ожилих із мертвих, а члени ваші Богові за знаряддя праведности.
ROM|6|14|Бо хай гріх не панує над вами, ви бо не під Законом, а під благодаттю.
ROM|6|15|Що ж? Чи будемо грішити, бо ми не під Законом, а під благодаттю? Зовсім ні!
ROM|6|16|Хіба ви не знаєте, що кому віддаєте себе за рабів на послух, то ви й раби того, кого слухаєтесь, або гріха на смерть, або послуху на праведність?
ROM|6|17|Тож дяка Богові, що ви, бувши рабами гріха, від серця послухались того роду науки, якому ви себе віддали.
ROM|6|18|А звільнившися від гріха, стали рабами праведности.
ROM|6|19|Говорю я по-людському, через неміч вашого тіла. Бо як ви віддавали були члени ваші за рабів нечистості й беззаконню на беззаконня, так тепер віддайте члени ваші за рабів праведности на освячення.
ROM|6|20|Бо коли були ви рабами гріха, то були вільні від праведности.
ROM|6|21|Який же плід ви мали тоді? Такі речі, що ними соромитесь тепер, бо кінець їх то смерть.
ROM|6|22|А тепер, звільнившися від гріха й ставши рабами Богові, маєте плід ваш на освячення, а кінець життя вічне.
ROM|6|23|Бо заплата за гріх смерть, а дар Божий вічне життя в Христі Ісусі, Господі нашім!
ROM|7|1|Чи ви не знаєте, браття, бо говорю тим, хто знає Закона, що Закон панує над людиною, поки вона живе?
ROM|7|2|Бо заміжня жінка, поки живе чоловік, прив'язана до нього Законом; а коли помре чоловік, вона звільняється від закону чоловіка.
ROM|7|3|Тому то, поки живе чоловік, вона буде вважатися перелюбницею, якщо стане дружиною іншому чоловікові; коли ж чоловік помре, вона вільна від Закону, і не буде перелюбницею, якщо стане за дружину іншому чоловікові.
ROM|7|4|Так, мої браття, і ви вмерли для Закону через тіло Христове, щоб належати вам іншому, Воскреслому з мертвих, щоб приносити плід Богові.
ROM|7|5|Бо коли ми жили за тілом, то пристрасті гріховні, що походять від Закону, діяли в наших членах, щоб приносити плід смерти.
ROM|7|6|А тепер ми звільнились від Закону, умерши для того, чим були зв'язані, щоб служити нам обновленням духа, а не старістю букви.
ROM|7|7|Що ж скажемо? Чи Закон то гріх? Зовсім ні! Але я не пізнав гріха, як тільки через Закон, бо я не знав би пожадливости, коли б Закон не наказував: Не пожадай.
ROM|7|8|Але гріх, узявши привід від заповіді, зробив у мені всяку пожадливість, бо без Закону гріх мертвий.
ROM|7|9|А я колись жив без Закону, але, коли прийшла заповідь, то гріх ожив,
ROM|7|10|а я вмер; і сталася мені та заповідь, що для життя, на смерть,
ROM|7|11|бо гріх, узявши причину від заповіді, звів мене, і нею вмертвив.
ROM|7|12|Тому то Закон святий, і заповідь свята, і праведна, і добра.
ROM|7|13|Тож чи добре стало мені смертю? Зовсім ні! Але гріх, щоб стати гріхом, приніс мені смерть добром, щоб гріх став міцно грішний через заповідь.
ROM|7|14|Бо ми знаємо, що Закон духовний, а я тілесний, проданий під гріх.
ROM|7|15|Бо що я виконую, не розумію; я бо чиню не те, що хочу, але що ненавиджу, те я роблю.
ROM|7|16|А коли роблю те, чого я не хочу, то згоджуюсь із Законом, що він добрий,
ROM|7|17|а тому вже не я це виконую, але гріх, що живе в мені.
ROM|7|18|Знаю бо, що не живе в мені, цебто в тілі моїм, добре; бо бажання лежить у мені, але щоб виконати добре, того не знаходжу.
ROM|7|19|Бо не роблю я доброго, що хочу, але зле, чого не хочу, це чиню.
ROM|7|20|Коли ж я роблю те, чого не хочу, то вже не я це виконую, але гріх, що живе в мені.
ROM|7|21|Тож знаходжу закона, коли хочу робити добро, що зло лежить у мені.
ROM|7|22|Бо маю задоволення в Законі Божому за внутрішнім чоловіком,
ROM|7|23|та бачу інший закон у членах своїх, що воює проти закону мого розуму, і полонить мене законом гріховним, що знаходиться в членах моїх.
ROM|7|24|Нещасна я людина! Хто мене визволить від тіла цієї смерти?
ROM|7|25|Дякую Богові через Ісуса Христа, Господа нашого. Тому то я сам служу розумом Законові Божому, але тілом закону гріховному...
ROM|8|1|Тож немає тепер жадного осуду тим, хто ходить у Христі Ісусі не за тілом, а за духом,
ROM|8|2|бо закон духа життя в Христі Ісусі визволив мене від закону гріха й смерти.
ROM|8|3|Бо що було неможливе для Закону, у чому був він безсилий тілом, Бог послав Сина Свого в подобі гріховного тіла, і за гріх осудив гріх у тілі,
ROM|8|4|щоб виконалось виправдання Закону на нас, що ходимо не за тілом, а за духом.
ROM|8|5|Бо ті, хто ходить за тілом, думають про тілесне, а хто за духом про духовне.
ROM|8|6|Бо думка тілесна то смерть, а думка духовна життя та мир,
ROM|8|7|думка бо тілесна ворожнеча на Бога, бо не кориться Законові Божому, та й не може.
ROM|8|8|І ті, хто ходить за тілом, не можуть догодити Богові.
ROM|8|9|А ви не в тілі, але в дусі, бо Дух Божий живе в вас. А коли хто не має Христового Духа, той не Його.
ROM|8|10|А коли Христос у вас, то хоч тіло мертве через гріх, але дух живий через праведність.
ROM|8|11|А коли живе в вас Дух Того, Хто воскресив Ісуса з мертвих, то Той, хто підняв Христа з мертвих, оживить і смертельні тіла ваші через Свого Духа, що живе в вас.
ROM|8|12|Тому то, браття, ми не боржники тіла, щоб жити за тілом;
ROM|8|13|бо коли живете за тілом, то маєте вмерти, а коли духом умертвляєте тілесні вчинки, то будете жити.
ROM|8|14|Бо всі, хто водиться Духом Божим, вони сини Божі;
ROM|8|15|бо не взяли ви духа неволі знов на страх, але взяли ви Духа синівства, що через Нього кличемо: Авва, Отче!
ROM|8|16|Сам Цей Дух свідчить разом із духом нашим, що ми діти Божі.
ROM|8|17|А коли діти, то й спадкоємці, спадкоємці ж Божі, а співспадкоємці Христові, коли тільки разом із Ним ми терпимо, щоб разом із Ним і прославитись.
ROM|8|18|Бо я думаю, що страждання теперішнього часу нічого не варті супроти тієї слави, що має з'явитися в нас.
ROM|8|19|Бо чекання створіння очікує з'явлення синів Божих,
ROM|8|20|бо створіння покорилось марноті не добровільно, але через того, хто скорив його, в надії,
ROM|8|21|що й саме створіння визволиться від неволі тління на волю слави синів Божих.
ROM|8|22|Бо знаємо, що все створіння разом зідхає й разом мучиться аж досі.
ROM|8|23|Але не тільки воно, але й ми самі, маючи зачаток Духа, і ми самі в собі зідхаємо, очікуючи синівства, відкуплення нашого тіла.
ROM|8|24|Надією бо ми спаслися. Надія ж, коли бачить, не є надія, бо хто що бачить, чому б того й надіявся?
ROM|8|25|А коли сподіваємось, чого не бачимо, то очікуємо того з терпеливістю.
ROM|8|26|Так само ж і Дух допомагає нам у наших немочах; бо ми не знаємо, про що маємо молитись, як належить, але Сам Дух заступається за нас невимовними зідханнями.
ROM|8|27|А Той, Хто досліджує серця, знає, яка думка Духа, бо з волі Божої заступається за святих.
ROM|8|28|І знаємо, що тим, хто любить Бога, хто покликаний Його постановою, усе допомагає на добре.
ROM|8|29|Бо кого Він передбачив, тих і призначив, щоб були подібні до образу Сина Його, щоб Він був перворідним поміж багатьма братами.
ROM|8|30|А кого Він призначив, тих і покликав, а кого покликав, тих і виправдав, а кого виправдав, тих і прославив.
ROM|8|31|Що ж скажем на це? Коли за нас Бог, то хто проти нас?
ROM|8|32|Той же, Хто Сина Свого не пожалів, але видав Його за всіх нас, як же не дав би Він нам із Ним і всього?
ROM|8|33|Хто оскаржувати буде Божих вибранців? Бог Той, що виправдує.
ROM|8|34|Хто ж той, що засуджує? Христос Ісус є Той, що вмер, надто й воскрес, Він праворуч Бога, і Він і заступається за нас.
ROM|8|35|Хто нас розлучить від любови Христової? Чи недоля, чи утиск, чи переслідування, чи голод, чи нагота, чи небезпека, чи меч?
ROM|8|36|Як написано: За Тебе нас цілий день умертвляють, нас уважають за овець, приречених на заколення.
ROM|8|37|Але в цьому всьому ми перемагаємо Тим, Хто нас полюбив.
ROM|8|38|Бо я пересвідчився, що ні смерть, ні життя, ні Анголи, ні влади, ні теперішнє, ні майбутнє, ні сили,
ROM|8|39|ні вишина, ні глибина, ані інше яке створіння не зможе відлучити нас від любови Божої, яка в Христі Ісусі, Господі нашім!
ROM|9|1|Кажу правду в Христі, не обманюю, як свідчить мені моє сумління через Духа Святого,
ROM|9|2|що маю велику скорботу й невпинну муку для серця свого!
ROM|9|3|Бо я бажав би сам бути відлучений від Христа замість братів моїх, рідних мені тілом;
ROM|9|4|вони ізраїльтяни, що їм належить синівство, і слава, і заповіти, і законодавство, і Богослужба, і обітниці,
ROM|9|5|що їхні й отці, і від них же тілом Христос, що Він над усіма Бог, благословенний, навіки, амінь.
ROM|9|6|Не так, щоб Слово Боже не збулося. Бо не всі ті ізраїльтяни, хто від Ізраїля,
ROM|9|7|і не всі діти Авраамові, хто від насіння його, але: в Ісаку буде насіння тобі.
ROM|9|8|Цебто, не тілесні діти то діти Божі, але діти обітниці признаються за насіння.
ROM|9|9|А слово обітниці таке: На той час прийду, і буде син у Сари.
ROM|9|10|І не тільки це, але й Ревекка зачала дітей від одного ложа отця нашого Ісака,
ROM|9|11|бо коли вони ще не народились, і нічого доброго чи злого не вчинили, щоб позосталась постанова Божа у вибранні
ROM|9|12|не від учинків, але від Того, Хто кличе, сказано їй: Більший служитиме меншому,
ROM|9|13|як і написано: Полюбив Я Якова, а Ісава зненавидів.
ROM|9|14|Що ж скажемо? Може в Бога неправда? Зовсім ні!
ROM|9|15|Бо Він каже Мойсеєві: Помилую, кого хочу помилувати, і змилосерджуся, над ким хочу змилосердитись.
ROM|9|16|Отож, не залежить це ні від того, хто хоче, ні від того, хто біжить, але від Бога, що милує.
ROM|9|17|Бо Писання говорить фараонові: Власне на те Я поставив тебе, щоб на тобі показати Свою силу, і щоб звістилось по цілій землі Моє Ймення.
ROM|9|18|Отож, кого хоче Він милує, і кого хоче ожорсточує.
ROM|9|19|А ти скажеш мені: Чого ж іще Він докоряє, бо хто може противитись волі Його?
ROM|9|20|Отже, хто ти, чоловіче, що ти сперечаєшся з Богом? Чи скаже твориво творцеві: Пощо ти зробив мене так?
ROM|9|21|Чи ганчар не має влади над глиною, щоб із того самого місива зробити одну посудину на честь, а одну на нечесть?
ROM|9|22|Тож Бог, бажаючи показати гнів і виявити могутність Свою, щадив із великим терпінням посудини гніву, що готові були на погибіль,
ROM|9|23|і щоб виявити багатство слави Своєї на посудинах милосердя, що їх приготував на славу,
ROM|9|24|на нас, що їх і покликав не тільки від юдеїв, але й від поган.
ROM|9|25|Як і в Осії Він говорить: Назву Своїм народом не людей Моїх, і не улюблену улюбленою,
ROM|9|26|і на місці, де сказано їм: Ви не Мій народ, там названі будуть синами Бога Живого!
ROM|9|27|А Ісая взиває про Ізраїля: Коли б число синів Ізраїлевих було, як морський пісок, то тільки останок спасеться,
ROM|9|28|бо вирок закінчений та скорочений учинить Господь на землі!
ROM|9|29|І як Ісая віщував: Коли б Господь Саваот не лишив нам насіння, то ми стали б, як Содом, і подібні були б до Гоморри!
ROM|9|30|Що ж скажемо? Що погани, які не шукали праведности, досягли праведности, тієї праведности, що від віри,
ROM|9|31|а Ізраїль, що шукав Закона праведности, не досяг Закону праведности.
ROM|9|32|Чому? Бо шукали не з віри, але якби з учинків Закону; вони бо спіткнулись об камінь спотикання,
ROM|9|33|як написано: Ось Я кладу на Сіоні камінь спотикання та скелю спокуси, і кожен, хто вірує в Нього, не посоромиться!
ROM|10|1|Браття, бажання мого серця й молитва до Бога за Ізраїля на спасіння.
ROM|10|2|Бо я свідчу їм, що вони мають ревність про Бога, але не за розумом.
ROM|10|3|Вони бо, не розуміючи праведности Божої, і силкуючись поставити власну праведність, не покорились праведності Божій.
ROM|10|4|Бо кінець Закону Христос на праведність кожному, хто вірує.
ROM|10|5|Мойсей бо пише про праведність, що від Закону, що людина, яка його виконує, буде ним жити.
ROM|10|6|А про праведність, що від віри, говорить так: Не кажи в своїм серці: Хто вийде на небо? цебто звести додолу Христа,
ROM|10|7|або: Хто зійде в безодню? цебто вивести з мертвих Христа.
ROM|10|8|Але що каже ще? Близько тебе слово, в устах твоїх і в серці твоїм, цебто слово віри, що його проповідуємо.
ROM|10|9|Бо коли ти устами своїми визнаватимеш Ісуса за Господа, і будеш вірувати в своїм серці, що Бог воскресив Його з мертвих, то спасешся,
ROM|10|10|бо серцем віруємо для праведности, а устами ісповідуємо для спасіння.
ROM|10|11|Каже бо Писання: Кожен, хто вірує в Нього, не буде засоромлений.
ROM|10|12|Бо нема різниці поміж юдеєм та гелленом, бо той же Господь є Господом усіх, багатий для всіх, хто кличе Його.
ROM|10|13|Бо кожен, хто покличе Господнє Ім'я, буде спасений.
ROM|10|14|Але як покличуть Того, в Кого не ввірували? А як увірують у Того, що про Нього не чули? А як почують без проповідника?
ROM|10|15|І як будуть проповідувати, коли не будуть послані? Як написано: Які гарні ноги благовісників миру, благовісників добра.
ROM|10|16|Але не всі послухались Євангелії. Бо Ісая каже: Господи, хто повірив тому, що почув був від нас?
ROM|10|17|Тож віра від слухання, а слухання через Слово Христове.
ROM|10|18|Та кажу: Чи не чули вони? Отож: По всій землі їхній голос пішов, і їхні слова в кінці світу!
ROM|10|19|Але кажу: Чи Ізраїль не знав? Перший Мойсей говорить: Я викличу заздрість у вас ненародом, роздражню вас нерозумним народом.
ROM|10|20|А Ісая сміливо говорить: Знайшли Мене ті, хто Мене не шукав, відкрився Я тим, хто не питався про Мене!
ROM|10|21|А про Ізраїля каже: Я руки Свої цілий день простягав до людей неслухняних і суперечних!
ROM|11|1|Отож я питаю: Чи ж Бог відкинув народа Свого? Зовсім ні! Бо й я ізраїльтянин, із насіння Авраамового, Веніяминового племени.
ROM|11|2|Не відкинув Бог народа Свого, що його перше знав. Чи ви не знаєте, що говорить Писання, де про Іллю, як він скаржиться Богові на Ізраїля, кажучи:
ROM|11|3|Господи, вони повбивали пророків Твоїх, і Твої жертівники поруйнували, і лишився я сам, і шукають моєї душі.
ROM|11|4|Та що каже йому Божа відповідь: Я для Себе зоставив сім тисяч мужа, що перед Ваалом колін не схилили.
ROM|11|5|Також і теперішнього часу залишився останок за вибором благодаті.
ROM|11|6|А коли за благодаттю, то не з учинків, інакше благодать не була б благодаттю. А коли з учинків, то це більше не благодать, інакше вчинок не є вже вчинок.
ROM|11|7|Що ж? Чого Ізраїль шукає, того не одержав, та одержали вибрані, а останні затверділи,
ROM|11|8|як написано: Бог дав їм духа засипання, очі, щоб не бачили, і вуха, щоб не чули, аж до сьогоднішнього дня.
ROM|11|9|А Давид каже: Нехай станеться стіл їхній за сітку й за пастку, і на спокусу, та їм на заплату;
ROM|11|10|нехай потемніють їхні очі, щоб не бачили, хай назавжди зігнеться хребет їхній!
ROM|11|11|Тож питаю: Чи ж спіткнулись вони, щоб упасти? Зовсім ні! Але з їхнього занепаду спасіння поганам, щоб викликати заздрість у них.
ROM|11|12|А коли їхній занепад багатство для світу, а їхнє упокорення багатство поганам, скільки ж більш повнота їхня?
ROM|11|13|Кажу бо я вам, поганам: через те, що я апостол поганів, я хвалю свою службу,
ROM|11|14|може як викличу заздрість у своїх за тілом, і спасу декого з них.
ROM|11|15|Коли ж відкинення їх то примирення світу, то що їхнє прийняття, як не життя з мертвих?
ROM|11|16|А коли святий первісток, то й тісто святе; а коли святий корінь, то й віття святе.
ROM|11|17|Коли ж деякі з галузок відломилися, а ти, бувши дике оливне дерево, прищепився між них і став спільником товщу оливного кореня,
ROM|11|18|то не вихваляйся перед галузками; а коли вихваляєшся, то знай, що не ти носиш кореня, але корінь тебе.
ROM|11|19|Отже скажеш: Галузки відломилися, щоб я прищепився.
ROM|11|20|Добре. Вони відломились невірством, а ти тримаєшся вірою; не величайся, але бійся.
ROM|11|21|Бо коли Бог природних галузок не пожалував, то Він і тебе не пожалує!
ROM|11|22|Отже, бач добрість і суворість Божу, на відпалих суворість, а на тебе добрість Божа, коли перебудеш у добрості, коли ж ні, то й ти будеш відтятий.
ROM|11|23|Та й вони, коли не зостануться в невірстві, прищепляться, бо має Бог силу їх знов прищепити.
ROM|11|24|Бо коли ти відтятий з оливки, дикої з природи, і проти природи защеплений до доброї оливки, то скільки ж більше ті, що природні, прищепляться до своєї власної оливки?
ROM|11|25|Бо не хочу я, браття, щоб ви не знали цієї таємниці, щоб не були ви високої думки про себе, що жорстокість сталась Ізраїлеві почасти, аж поки не ввійде повне число поган,
ROM|11|26|і так увесь Ізраїль спасеться, як написано: Прийде з Сіону Спаситель, і відверне безбожність від Якова,
ROM|11|27|і це заповіт їм від Мене, коли відійму гріхи їхні!
ROM|11|28|Тож вони за Євангелією вороги ради вас, а за вибором улюблені ради отців.
ROM|11|29|Бо дари й покликання Божі невідмінні.
ROM|11|30|Бо як і ви були колись неслухняні Богові, а тепер помилувані через їхній непослух,
ROM|11|31|так і вони тепер спротивились для помилування вас, щоб і самі були помилувані.
ROM|11|32|Бо замкнув Бог усіх у непослух, щоб помилувати всіх.
ROM|11|33|О глибино багатства, і премудрости, і знання Божого! Які недовідомі присуди Його, і недосліджені дороги Його!
ROM|11|34|Бо хто розум Господній пізнав? Або хто був дорадник Йому?
ROM|11|35|Або хто давніш Йому дав, і йому буде віддано?
ROM|11|36|Бо все з Нього, через Нього і для Нього! Йому слава навіки. Амінь.
ROM|12|1|Тож благаю вас, браття, через Боже милосердя, повіддавайте ваші тіла на жертву живу, святу, приємну Богові, як розумну службу вашу,
ROM|12|2|і не стосуйтесь до віку цього, але перемініться відновою вашого розуму, щоб пізнати вам, що то є воля Божа, добро, приємність та досконалість.
ROM|12|3|Через дану мені благодать кажу кожному з вас не думати про себе більш, ніж належить думати, але думати скромно, у міру віри, як кожному Бог наділив.
ROM|12|4|Бо як в однім тілі маємо багато членів, а всі члени мають не однакове діяння,
ROM|12|5|так багато нас є одне тіло в Христі, а зосібна ми один одному члени.
ROM|12|6|І ми маємо різні дари, згідно з благодаттю, даною нам: коли пророцтво то виконуй його в міру віри,
ROM|12|7|а коли служіння будь на служіння, коли вчитель на навчання,
ROM|12|8|коли втішитель на потішання, хто подає у простоті, хто головує то з пильністю, хто милосердствує то з привітністю!
ROM|12|9|Любов нехай буде нелицемірна; ненавидьте зло та туліться до доброго!
ROM|12|10|Любіть один одного братньою любов'ю; випереджайте один одного пошаною!
ROM|12|11|У ревності не лінуйтеся, духом палайте, служіть Господеві,
ROM|12|12|тіштесь надією, утиски терпіть, перебувайте в молитві,
ROM|12|13|беріть уділ у потребах святих, будьте гостинні до чужинців!
ROM|12|14|Благословляйте тих, хто вас переслідує; благословляйте, а не проклинайте!
ROM|12|15|Тіштеся з тими, хто тішиться, і плачте з отими, хто плаче!
ROM|12|16|Думайте між собою однаково; не величайтеся, але наслідуйте слухняних; не вважайте за мудрих себе!
ROM|12|17|Не платіть нікому злом за зло, дбайте про добре перед усіма людьми!
ROM|12|18|Коли можливо, якщо це залежить від вас, живіть у мирі зо всіма людьми!
ROM|12|19|Не мстіться самі, улюблені, але дайте місце гніву Божому, бо написано: Мені помста належить, Я відплачу, говорить Господь.
ROM|12|20|Отож, як твій ворог голодний, нагодуй його; як він прагне, напій його, бо, роблячи це, ти згортаєш розпалене вугілля йому на голову.
ROM|12|21|Не будь переможений злом, але перемагай зло добром!
ROM|13|1|Нехай кожна людина кориться вищій владі, бо немає влади, як не від Бога, і влади існуючі встановлені від Бога.
ROM|13|2|Тому той, хто противиться владі, противиться Божій постанові; а ті, хто противиться, самі візьмуть осуд на себе.
ROM|13|3|Бо володарі пострах не на добрі діла, а на злі. Хочеш не боятися влади? Роби добро, і матимеш похвалу від неї,
ROM|13|4|бо володар Божий слуга, тобі на добро. А як чиниш ти зле, то бійся, бо недармо він носить меча, він бо Божий слуга, месник у гніві злочинцеві!
ROM|13|5|Тому треба коритися не тільки ради страху кари, але й ради сумління.
ROM|13|6|Через це ви й податки даєте, бо вони служителі Божі, саме тим завжди зайняті.
ROM|13|7|Тож віддайте належне усім: кому податок податок, кому мито мито, кому страх страх, кому честь честь.
ROM|13|8|Не будьте винні нікому нічого, крім того, щоб любити один одного. Бо хто іншого любить, той виконав Закона.
ROM|13|9|Бо заповіді: Не чини перелюбу, Не вбивай, Не кради, Не свідкуй неправдиво, Не пожадай й які інші, вони містяться всі в цьому слові: Люби свого ближнього, як самого себе!
ROM|13|10|Любов не чинить зла ближньому, тож любов виконання Закону.
ROM|13|11|І це тому, що знаєте час, що пора нам уже пробудитись від сну. Бо тепер спасіння ближче до нас, аніж тоді, коли ми ввірували.
ROM|13|12|Ніч минула, а день наблизився, тож відкиньмо вчинки темряви й зодягнімось у зброю світла.
ROM|13|13|Як удень, поступаймо доброчесно, не в гульні та п'янстві, не в перелюбі та розпусті, не в сварні та заздрощах,
ROM|13|14|але зодягніться Господом Ісусом Христом, а догодження тілу не обертайте на пожадливість!
ROM|14|1|Слабого в вірі приймайте, але не для суперечок про погляди.
ROM|14|2|Один бо вірує, що можна їсти все, а немічний споживає ярину.
ROM|14|3|Хто їсть, нехай не погорджує тим, хто не їсть. А хто не їсть, нехай не осуджує того, хто їсть, Бог бо прийняв його.
ROM|14|4|Ти хто такий, що судиш чужого раба? Він для пана свого стоїть або падає; але він устоїть, бо має Бог силу поставити його.
ROM|14|5|Один вирізнює день від дня, інший же про кожен день судить однаково. Нехай кожен за власною думкою тримається свого переконання.
ROM|14|6|Хто вважає на день, для Господа вважає, а хто не вважає на день, для Господа не вважає. Хто їсть, для Господа їсть, бо дякує Богові. А хто не їсть, для Господа не їсть, і дякує Богові.
ROM|14|7|Бо ніхто з нас не живе сам для себе, і не вмирає ніхто сам для себе.
ROM|14|8|Бо коли живемо для Господа живемо, і коли вмираємо для Господа вмираємо. І чи живемо, чи вмираємо ми Господні!
ROM|14|9|Бо Христос на те й умер, і ожив, щоб панувати і над мертвими, і над живими.
ROM|14|10|А ти нащо осуджуєш брата свого? Чи чого ти погорджуєш братом своїм? Бо всі станемо перед судним престолом Божим.
ROM|14|11|Бо написано: Я живу, каже Господь, і схилиться кожне коліно передо Мною, і визнає Бога кожен язик!
ROM|14|12|Тому кожен із нас сам за себе дасть відповідь Богові.
ROM|14|13|Отож, не будемо більше осуджувати один одного, але краще судіть про те, щоб не давати братові спотикання та спокуси.
ROM|14|14|Я знаю, і пересвідчений у Господі Ісусі, що нема нічого нечистого в самому собі; тільки коли хто вважає що за нечисте, тому воно нечисте.
ROM|14|15|Коли ж через поживу сумує твій брат, то вже не за любов'ю поводишся ти, не губи своєю поживою того, за кого Христос був умер.
ROM|14|16|Нехай ваше добре не зневажається.
ROM|14|17|Бо Царство Боже не пожива й питво, але праведність, і мир, і радість у Дусі Святім.
ROM|14|18|Хто цим служить Христові, той Богові милий і шанований поміж людьми.
ROM|14|19|Отож, пильнуймо про мир, та про те, що на збудування один одного!
ROM|14|20|Не руйнуй діла Божого ради поживи, усе бо чисте, але зле людині, що їсть на спотикання.
ROM|14|21|Добре не їсти м'яса, ані пити вина, ані робити такого, від чого брат твій гіршиться, або спокушується, або слабне.
ROM|14|22|Ти маєш віру? Май її сам про себе перед Богом. Блаженний той, хто не осуджує самого себе за те, про що випробовується!
ROM|14|23|А хто має сумнів, коли їсть, буде осуджений, бо не робить із віри, а що не від віри, те гріх.
ROM|15|1|Ми, сильні, повинні нести слабості безсилих, а не собі догоджати.
ROM|15|2|Кожен із нас нехай догоджає ближньому на добро для збудування.
ROM|15|3|Бо й Христос не Собі догоджав, але як написано: Зневаги тих, хто Тебе зневажає, упали на Мене.
ROM|15|4|А все, що давніше написане, написане нам на науку, щоб терпінням і потіхою з Писання ми мали надію.
ROM|15|5|А Бог терпеливости й потіхи нехай дасть вам бути однодумними між собою за Христом Ісусом,
ROM|15|6|щоб ви однодушно, одними устами славили Бога й Отця Господа нашого Ісуса Христа.
ROM|15|7|Приймайте тому один одного, як і Христос прийняв нас до Божої слави.
ROM|15|8|Кажу ж, що Христос для обрізаних став за служку ради Божої правди, щоб отцям потвердити обітниці,
ROM|15|9|а для поган щоб славили Бога за милосердя, як написано: Тому я хвалитиму Тебе, Господи, серед поган, і Ім'я Твоє буду виспівувати!
ROM|15|10|І ще каже: Тіштесь, погани, з народом Його!
ROM|15|11|І ще: Хваліть, усі погани, Господа, виславляйте Його, усі люди!
ROM|15|12|І ще каже Ісая: Буде корінь Єссеїв, що постане, щоб панувати над поганами, погани на Нього надіятись будуть!
ROM|15|13|Бог же надії нехай вас наповнить усякою радістю й миром у вірі, щоб ви збагатились надією, силою Духа Святого!
ROM|15|14|І я про вас сам пересвідчений, браття мої, що й самі ви повні добрости, наповнені всяким знанням, і можете й один одного навчати.
ROM|15|15|А писав я вам почасти трохи сміліше, якби вам нагадуючи благодаттю, що дана мені від Бога,
ROM|15|16|щоб був я слугою Христа Ісуса між поганами, і виконував святу службу Євангелії Божої, щоб приношення поган стало приємне й освячене Духом Святим.
ROM|15|17|Тож маю я чим похвалитись у Христі Ісусі, щодо Божих речей,
ROM|15|18|бо не смію казати того, чого не зробив через мене Христос на послух поган, словом і чином,
ROM|15|19|силою ознак і чудес, силою Духа Божого, так що я поширив Євангелію Христову від Єрусалиму й околиць аж до Ілліріка.
ROM|15|20|При тому пильнував я звіщати Євангелію не там, де Христове Ім'я було знане, щоб не будувати на основі чужій,
ROM|15|21|але як написано: Кому не звіщалось про Нього, побачать, і ті, хто не чув, зрозуміють!
ROM|15|22|Тому часто я мав перешкоди, щоб прибути до вас.
ROM|15|23|А тепер, не маючи більше місця в країнах оцих, але з давніх літ мавши бажання прибути до вас,
ROM|15|24|коли тільки піду до Еспанії, прибуду до вас. Бо маю надію, як буду проходити, побачити вас, і що ви проведете мене туди, коли перше почасти матиму я задоволення з вами побути.
ROM|15|25|А тепер я йду до Єрусалиму послужити святим,
ROM|15|26|бо Македонія й Ахая визнали за добре подати деяку поміч незаможним святим, що в Єрусалимі живуть.
ROM|15|27|Бо визнали за добре, та й боржники вони їхні. Бо коли погани стали спільниками в їх духовнім, то повинні й у тілеснім послужити їм.
ROM|15|28|Як це докінчу та достачу їм плід цей, тоді через ваше місто я піду до Еспанії.
ROM|15|29|І знаю, що коли прийду до вас, то прийду в повноті Христового благословення.
ROM|15|30|Благаю ж вас, браття, Господом нашим Ісусом Христом і любов'ю Духа, помагайте мені в молитвах за мене до Бога,
ROM|15|31|щоб мені визволитися від неслухняних в Юдеї, і щоб служба моя в Єрусалимі була приємна святим,
ROM|15|32|щоб із волі Божої з радістю прийти до вас і відпочити з вами!
ROM|15|33|А Бог миру нехай буде зо всіма вами. Амінь.
ROM|16|1|Поручаю ж вам сестру нашу Фіву, служебницю Церкви в Кенхреях,
ROM|16|2|щоб ви прийняли її в Господі, як личить святим, і допомагайте їй, у якій речі буде вона чого потребувати від вас, бо й вона опікунка була багатьом і самому мені.
ROM|16|3|Вітайте Прискиллу й Акилу, співробітників моїх у Христі Ісусі,
ROM|16|4|що голови свої за душу мою клали, яким не я сам дякую, але й усі Церкви з поган, і їхню домашню Церкву.
ROM|16|5|Вітайте улюбленого мого Епенета, він первісток Ахаї для Христа.
ROM|16|6|Вітайте Марію, що напрацювалася багато для вас.
ROM|16|7|Вітайте Андроніка й Юнія, родичів моїх і співв'язнів моїх, що славні вони між апостолами, що й у Христі були перше мене.
ROM|16|8|Вітайте Амплія, мого улюбленого в Господі.
ROM|16|9|Вітайте Урбана, співробітника нашого в Христі, і улюбленого мого Стахія.
ROM|16|10|Вітайте Апеллеса, випробуваного в Христі. Вітайте Аристовулових.
ROM|16|11|Вітайте мого родича Іродіона. Вітайте Наркисових, що в Господі.
ROM|16|12|Вітайте Трифену й Трифосу, що працюють у Господі. Вітайте улюблену Персиду, що багато попрацювала в Господі.
ROM|16|13|Вітайте вибраного в Господі Руфа, і матір його та мою.
ROM|16|14|Вітайте Асинкрита, Флегонта, Єрма, Патрова, Єрмія і братів, що з ними.
ROM|16|15|Вітайте Філолога та Юлію, Нірея й сестру його, і Олімпіяна, і всіх святих, що з ними.
ROM|16|16|Вітайте один одного святим поцілунком. Вітають вас усі Церкви Христові!
ROM|16|17|Благаю ж вас, браття, щоб ви остерігалися тих, хто чинить розділення й згіршення проти науки, якої ви навчилися, і уникайте їх,
ROM|16|18|бо такі не служать Господеві нашому Ісусу Христу, але власному череву; вони добрими та гарними словами зводять серця простодушних.
ROM|16|19|Ваша ж слухняність дійшла до всіх. І я тішусь за вас, але хочу, щоб були ви мудрі в доброму, а прості в злому.
ROM|16|20|А Бог миру потопче незабаром сатану під ваші ноги. Благодать Господа нашого Ісуса Христа нехай буде з вами! Амінь.
ROM|16|21|Вітає вас мій співробітник Тимофій, і Лукій, і Ясон, і Сосипатр, мої родичі.
ROM|16|22|Вітаю вас у Господі й я, Тертій, що цього листа написав.
ROM|16|23|Вітає вас Гай, гостинний для мене й цілої Церкви. Вітає вас міський доморядник Ераст і брат Кварт.
ROM|16|24|Благодать Господа нашого Ісуса Христа нехай буде зо всіма вами! Амінь.
ROM|16|25|А Тому, хто може поставити вас міцно згідно з моєю Євангелією й проповіддю Ісуса Христа, за об'явленням таємниці, що від вічних часів була замовчана,
ROM|16|26|а тепер виявлена, і через пророцькі писання, з наказу вічного Бога, на послух вірі по всіх народах провіщена,
ROM|16|27|єдиному мудрому Богові, через Ісуса Христа, слава навіки! Амінь.
