2COR|1|1|Paul, an apostle of Jesus Christ by the will of God, and Timothy our brother, unto the church of God which is at Corinth, with all the saints which are in all Achaia:
2COR|1|2|Grace be to you and peace from God our Father, and from the Lord Jesus Christ.
2COR|1|3|Blessed be God, even the Father of our Lord Jesus Christ, the Father of mercies, and the God of all comfort;
2COR|1|4|Who comforteth us in all our tribulation, that we may be able to comfort them which are in any trouble, by the comfort wherewith we ourselves are comforted of God.
2COR|1|5|For as the sufferings of Christ abound in us, so our consolation also aboundeth by Christ.
2COR|1|6|And whether we be afflicted, it is for your consolation and salvation, which is effectual in the enduring of the same sufferings which we also suffer: or whether we be comforted, it is for your consolation and salvation.
2COR|1|7|And our hope of you is stedfast, knowing, that as ye are partakers of the sufferings, so shall ye be also of the consolation.
2COR|1|8|For we would not, brethren, have you ignorant of our trouble which came to us in Asia, that we were pressed out of measure, above strength, insomuch that we despaired even of life:
2COR|1|9|But we had the sentence of death in ourselves, that we should not trust in ourselves, but in God which raiseth the dead:
2COR|1|10|Who delivered us from so great a death, and doth deliver: in whom we trust that he will yet deliver us;
2COR|1|11|Ye also helping together by prayer for us, that for the gift bestowed upon us by the means of many persons thanks may be given by many on our behalf.
2COR|1|12|For our rejoicing is this, the testimony of our conscience, that in simplicity and godly sincerity, not with fleshly wisdom, but by the grace of God, we have had our conversation in the world, and more abundantly to you-ward.
2COR|1|13|For we write none other things unto you, than what ye read or acknowledge; and I trust ye shall acknowledge even to the end;
2COR|1|14|As also ye have acknowledged us in part, that we are your rejoicing, even as ye also are our's in the day of the Lord Jesus.
2COR|1|15|And in this confidence I was minded to come unto you before, that ye might have a second benefit;
2COR|1|16|And to pass by you into Macedonia, and to come again out of Macedonia unto you, and of you to be brought on my way toward Judaea.
2COR|1|17|When I therefore was thus minded, did I use lightness? or the things that I purpose, do I purpose according to the flesh, that with me there should be yea yea, and nay nay?
2COR|1|18|But as God is true, our word toward you was not yea and nay.
2COR|1|19|For the Son of God, Jesus Christ, who was preached among you by us, even by me and Silvanus and Timotheus, was not yea and nay, but in him was yea.
2COR|1|20|For all the promises of God in him are yea, and in him Amen, unto the glory of God by us.
2COR|1|21|Now he which stablisheth us with you in Christ, and hath anointed us, is God;
2COR|1|22|Who hath also sealed us, and given the earnest of the Spirit in our hearts.
2COR|1|23|Moreover I call God for a record upon my soul, that to spare you I came not as yet unto Corinth.
2COR|1|24|Not for that we have dominion over your faith, but are helpers of your joy: for by faith ye stand.
2COR|2|1|But I determined this with myself, that I would not come again to you in heaviness.
2COR|2|2|For if I make you sorry, who is he then that maketh me glad, but the same which is made sorry by me?
2COR|2|3|And I wrote this same unto you, lest, when I came, I should have sorrow from them of whom I ought to rejoice; having confidence in you all, that my joy is the joy of you all.
2COR|2|4|For out of much affliction and anguish of heart I wrote unto you with many tears; not that ye should be grieved, but that ye might know the love which I have more abundantly unto you.
2COR|2|5|But if any have caused grief, he hath not grieved me, but in part: that I may not overcharge you all.
2COR|2|6|Sufficient to such a man is this punishment, which was inflicted of many.
2COR|2|7|So that contrariwise ye ought rather to forgive him, and comfort him, lest perhaps such a one should be swallowed up with overmuch sorrow.
2COR|2|8|Wherefore I beseech you that ye would confirm your love toward him.
2COR|2|9|For to this end also did I write, that I might know the proof of you, whether ye be obedient in all things.
2COR|2|10|To whom ye forgive any thing, I forgive also: for if I forgave any thing, to whom I forgave it, for your sakes forgave I it in the person of Christ;
2COR|2|11|Lest Satan should get an advantage of us: for we are not ignorant of his devices.
2COR|2|12|Furthermore, when I came to Troas to preach Christ's gospel, and a door was opened unto me of the Lord,
2COR|2|13|I had no rest in my spirit, because I found not Titus my brother: but taking my leave of them, I went from thence into Macedonia.
2COR|2|14|Now thanks be unto God, which always causeth us to triumph in Christ, and maketh manifest the savour of his knowledge by us in every place.
2COR|2|15|For we are unto God a sweet savour of Christ, in them that are saved, and in them that perish:
2COR|2|16|To the one we are the savour of death unto death; and to the other the savour of life unto life. And who is sufficient for these things?
2COR|2|17|For we are not as many, which corrupt the word of God: but as of sincerity, but as of God, in the sight of God speak we in Christ.
2COR|3|1|Do we begin again to commend ourselves? or need we, as some others, epistles of commendation to you, or letters of commendation from you?
2COR|3|2|Ye are our epistle written in our hearts, known and read of all men:
2COR|3|3|Forasmuch as ye are manifestly declared to be the epistle of Christ ministered by us, written not with ink, but with the Spirit of the living God; not in tables of stone, but in fleshy tables of the heart.
2COR|3|4|And such trust have we through Christ to God-ward:
2COR|3|5|Not that we are sufficient of ourselves to think any thing as of ourselves; but our sufficiency is of God;
2COR|3|6|Who also hath made us able ministers of the new testament; not of the letter, but of the spirit: for the letter killeth, but the spirit giveth life.
2COR|3|7|But if the ministration of death, written and engraven in stones, was glorious, so that the children of Israel could not stedfastly behold the face of Moses for the glory of his countenance; which glory was to be done away:
2COR|3|8|How shall not the ministration of the spirit be rather glorious?
2COR|3|9|For if the ministration of condemnation be glory, much more doth the ministration of righteousness exceed in glory.
2COR|3|10|For even that which was made glorious had no glory in this respect, by reason of the glory that excelleth.
2COR|3|11|For if that which is done away was glorious, much more that which remaineth is glorious.
2COR|3|12|Seeing then that we have such hope, we use great plainness of speech:
2COR|3|13|And not as Moses, which put a vail over his face, that the children of Israel could not stedfastly look to the end of that which is abolished:
2COR|3|14|But their minds were blinded: for until this day remaineth the same vail untaken away in the reading of the old testament; which vail is done away in Christ.
2COR|3|15|But even unto this day, when Moses is read, the vail is upon their heart.
2COR|3|16|Nevertheless when it shall turn to the Lord, the vail shall be taken away.
2COR|3|17|Now the Lord is that Spirit: and where the Spirit of the Lord is, there is liberty.
2COR|3|18|But we all, with open face beholding as in a glass the glory of the Lord, are changed into the same image from glory to glory, even as by the Spirit of the Lord.
2COR|4|1|Therefore seeing we have this ministry, as we have received mercy, we faint not;
2COR|4|2|But have renounced the hidden things of dishonesty, not walking in craftiness, nor handling the word of God deceitfully; but by manifestation of the truth commending ourselves to every man's conscience in the sight of God.
2COR|4|3|But if our gospel be hid, it is hid to them that are lost:
2COR|4|4|In whom the god of this world hath blinded the minds of them which believe not, lest the light of the glorious gospel of Christ, who is the image of God, should shine unto them.
2COR|4|5|For we preach not ourselves, but Christ Jesus the Lord; and ourselves your servants for Jesus' sake.
2COR|4|6|For God, who commanded the light to shine out of darkness, hath shined in our hearts, to give the light of the knowledge of the glory of God in the face of Jesus Christ.
2COR|4|7|But we have this treasure in earthen vessels, that the excellency of the power may be of God, and not of us.
2COR|4|8|We are troubled on every side, yet not distressed; we are perplexed, but not in despair;
2COR|4|9|Persecuted, but not forsaken; cast down, but not destroyed;
2COR|4|10|Always bearing about in the body the dying of the Lord Jesus, that the life also of Jesus might be made manifest in our body.
2COR|4|11|For we which live are alway delivered unto death for Jesus' sake, that the life also of Jesus might be made manifest in our mortal flesh.
2COR|4|12|So then death worketh in us, but life in you.
2COR|4|13|We having the same spirit of faith, according as it is written, I believed, and therefore have I spoken; we also believe, and therefore speak;
2COR|4|14|Knowing that he which raised up the Lord Jesus shall raise up us also by Jesus, and shall present us with you.
2COR|4|15|For all things are for your sakes, that the abundant grace might through the thanksgiving of many redound to the glory of God.
2COR|4|16|For which cause we faint not; but though our outward man perish, yet the inward man is renewed day by day.
2COR|4|17|For our light affliction, which is but for a moment, worketh for us a far more exceeding and eternal weight of glory;
2COR|4|18|While we look not at the things which are seen, but at the things which are not seen: for the things which are seen are temporal; but the things which are not seen are eternal.
2COR|5|1|For we know that if our earthly house of this tabernacle were dissolved, we have a building of God, an house not made with hands, eternal in the heavens.
2COR|5|2|For in this we groan, earnestly desiring to be clothed upon with our house which is from heaven:
2COR|5|3|If so be that being clothed we shall not be found naked.
2COR|5|4|For we that are in this tabernacle do groan, being burdened: not for that we would be unclothed, but clothed upon, that mortality might be swallowed up of life.
2COR|5|5|Now he that hath wrought us for the selfsame thing is God, who also hath given unto us the earnest of the Spirit.
2COR|5|6|Therefore we are always confident, knowing that, whilst we are at home in the body, we are absent from the Lord:
2COR|5|7|(For we walk by faith, not by sight:)
2COR|5|8|We are confident, I say, and willing rather to be absent from the body, and to be present with the Lord.
2COR|5|9|Wherefore we labour, that, whether present or absent, we may be accepted of him.
2COR|5|10|For we must all appear before the judgment seat of Christ; that every one may receive the things done in his body, according to that he hath done, whether it be good or bad.
2COR|5|11|Knowing therefore the terror of the Lord, we persuade men; but we are made manifest unto God; and I trust also are made manifest in your consciences.
2COR|5|12|For we commend not ourselves again unto you, but give you occasion to glory on our behalf, that ye may have somewhat to answer them which glory in appearance, and not in heart.
2COR|5|13|For whether we be beside ourselves, it is to God: or whether we be sober, it is for your cause.
2COR|5|14|For the love of Christ constraineth us; because we thus judge, that if one died for all, then were all dead:
2COR|5|15|And that he died for all, that they which live should not henceforth live unto themselves, but unto him which died for them, and rose again.
2COR|5|16|Wherefore henceforth know we no man after the flesh: yea, though we have known Christ after the flesh, yet now henceforth know we him no more.
2COR|5|17|Therefore if any man be in Christ, he is a new creature: old things are passed away; behold, all things are become new.
2COR|5|18|And all things are of God, who hath reconciled us to himself by Jesus Christ, and hath given to us the ministry of reconciliation;
2COR|5|19|To wit, that God was in Christ, reconciling the world unto himself, not imputing their trespasses unto them; and hath committed unto us the word of reconciliation.
2COR|5|20|Now then we are ambassadors for Christ, as though God did beseech you by us: we pray you in Christ's stead, be ye reconciled to God.
2COR|5|21|For he hath made him to be sin for us, who knew no sin; that we might be made the righteousness of God in him.
2COR|6|1|We then, as workers together with him, beseech you also that ye receive not the grace of God in vain.
2COR|6|2|(For he saith, I have heard thee in a time accepted, and in the day of salvation have I succoured thee: behold, now is the accepted time; behold, now is the day of salvation.)
2COR|6|3|Giving no offence in any thing, that the ministry be not blamed:
2COR|6|4|But in all things approving ourselves as the ministers of God, in much patience, in afflictions, in necessities, in distresses,
2COR|6|5|In stripes, in imprisonments, in tumults, in labours, in watchings, in fastings;
2COR|6|6|By pureness, by knowledge, by longsuffering, by kindness, by the Holy Ghost, by love unfeigned,
2COR|6|7|By the word of truth, by the power of God, by the armour of righteousness on the right hand and on the left,
2COR|6|8|By honour and dishonour, by evil report and good report: as deceivers, and yet true;
2COR|6|9|As unknown, and yet well known; as dying, and, behold, we live; as chastened, and not killed;
2COR|6|10|As sorrowful, yet alway rejoicing; as poor, yet making many rich; as having nothing, and yet possessing all things.
2COR|6|11|O ye Corinthians, our mouth is open unto you, our heart is enlarged.
2COR|6|12|Ye are not straitened in us, but ye are straitened in your own bowels.
2COR|6|13|Now for a recompence in the same, (I speak as unto my children,) be ye also enlarged.
2COR|6|14|Be ye not unequally yoked together with unbelievers: for what fellowship hath righteousness with unrighteousness? and what communion hath light with darkness?
2COR|6|15|And what concord hath Christ with Belial? or what part hath he that believeth with an infidel?
2COR|6|16|And what agreement hath the temple of God with idols? for ye are the temple of the living God; as God hath said, I will dwell in them, and walk in them; and I will be their God, and they shall be my people.
2COR|6|17|Wherefore come out from among them, and be ye separate, saith the Lord, and touch not the unclean thing; and I will receive you.
2COR|6|18|And will be a Father unto you, and ye shall be my sons and daughters, saith the Lord Almighty.
2COR|7|1|Having therefore these promises, dearly beloved, let us cleanse ourselves from all filthiness of the flesh and spirit, perfecting holiness in the fear of God.
2COR|7|2|Receive us; we have wronged no man, we have corrupted no man, we have defrauded no man.
2COR|7|3|I speak not this to condemn you: for I have said before, that ye are in our hearts to die and live with you.
2COR|7|4|Great is my boldness of speech toward you, great is my glorying of you: I am filled with comfort, I am exceeding joyful in all our tribulation.
2COR|7|5|For, when we were come into Macedonia, our flesh had no rest, but we were troubled on every side; without were fightings, within were fears.
2COR|7|6|Nevertheless God, that comforteth those that are cast down, comforted us by the coming of Titus;
2COR|7|7|And not by his coming only, but by the consolation wherewith he was comforted in you, when he told us your earnest desire, your mourning, your fervent mind toward me; so that I rejoiced the more.
2COR|7|8|For though I made you sorry with a letter, I do not repent, though I did repent: for I perceive that the same epistle hath made you sorry, though it were but for a season.
2COR|7|9|Now I rejoice, not that ye were made sorry, but that ye sorrowed to repentance: for ye were made sorry after a godly manner, that ye might receive damage by us in nothing.
2COR|7|10|For godly sorrow worketh repentance to salvation not to be repented of: but the sorrow of the world worketh death.
2COR|7|11|For behold this selfsame thing, that ye sorrowed after a godly sort, what carefulness it wrought in you, yea, what clearing of yourselves, yea, what indignation, yea, what fear, yea, what vehement desire, yea, what zeal, yea, what revenge! In all things ye have approved yourselves to be clear in this matter.
2COR|7|12|Wherefore, though I wrote unto you, I did it not for his cause that had done the wrong, nor for his cause that suffered wrong, but that our care for you in the sight of God might appear unto you.
2COR|7|13|Therefore we were comforted in your comfort: yea, and exceedingly the more joyed we for the joy of Titus, because his spirit was refreshed by you all.
2COR|7|14|For if I have boasted any thing to him of you, I am not ashamed; but as we spake all things to you in truth, even so our boasting, which I made before Titus, is found a truth.
2COR|7|15|And his inward affection is more abundant toward you, whilst he remembereth the obedience of you all, how with fear and trembling ye received him.
2COR|7|16|I rejoice therefore that I have confidence in you in all things.
2COR|8|1|Moreover, brethren, we do you to wit of the grace of God bestowed on the churches of Macedonia;
2COR|8|2|How that in a great trial of affliction the abundance of their joy and their deep poverty abounded unto the riches of their liberality.
2COR|8|3|For to their power, I bear record, yea, and beyond their power they were willing of themselves;
2COR|8|4|Praying us with much intreaty that we would receive the gift, and take upon us the fellowship of the ministering to the saints.
2COR|8|5|And this they did, not as we hoped, but first gave their own selves to the Lord, and unto us by the will of God.
2COR|8|6|Insomuch that we desired Titus, that as he had begun, so he would also finish in you the same grace also.
2COR|8|7|Therefore, as ye abound in every thing, in faith, and utterance, and knowledge, and in all diligence, and in your love to us, see that ye abound in this grace also.
2COR|8|8|I speak not by commandment, but by occasion of the forwardness of others, and to prove the sincerity of your love.
2COR|8|9|For ye know the grace of our Lord Jesus Christ, that, though he was rich, yet for your sakes he became poor, that ye through his poverty might be rich.
2COR|8|10|And herein I give my advice: for this is expedient for you, who have begun before, not only to do, but also to be forward a year ago.
2COR|8|11|Now therefore perform the doing of it; that as there was a readiness to will, so there may be a performance also out of that which ye have.
2COR|8|12|For if there be first a willing mind, it is accepted according to that a man hath, and not according to that he hath not.
2COR|8|13|For I mean not that other men be eased, and ye burdened:
2COR|8|14|But by an equality, that now at this time your abundance may be a supply for their want, that their abundance also may be a supply for your want: that there may be equality:
2COR|8|15|As it is written, He that had gathered much had nothing over; and he that had gathered little had no lack.
2COR|8|16|But thanks be to God, which put the same earnest care into the heart of Titus for you.
2COR|8|17|For indeed he accepted the exhortation; but being more forward, of his own accord he went unto you.
2COR|8|18|And we have sent with him the brother, whose praise is in the gospel throughout all the churches;
2COR|8|19|And not that only, but who was also chosen of the churches to travel with us with this grace, which is administered by us to the glory of the same Lord, and declaration of your ready mind:
2COR|8|20|Avoiding this, that no man should blame us in this abundance which is administered by us:
2COR|8|21|Providing for honest things, not only in the sight of the Lord, but also in the sight of men.
2COR|8|22|And we have sent with them our brother, whom we have oftentimes proved diligent in many things, but now much more diligent, upon the great confidence which I have in you.
2COR|8|23|Whether any do enquire of Titus, he is my partner and fellowhelper concerning you: or our brethren be enquired of, they are the messengers of the churches, and the glory of Christ.
2COR|8|24|Wherefore shew ye to them, and before the churches, the proof of your love, and of our boasting on your behalf.
2COR|9|1|For as touching the ministering to the saints, it is superfluous for me to write to you:
2COR|9|2|For I know the forwardness of your mind, for which I boast of you to them of Macedonia, that Achaia was ready a year ago; and your zeal hath provoked very many.
2COR|9|3|Yet have I sent the brethren, lest our boasting of you should be in vain in this behalf; that, as I said, ye may be ready:
2COR|9|4|Lest haply if they of Macedonia come with me, and find you unprepared, we (that we say not, ye) should be ashamed in this same confident boasting.
2COR|9|5|Therefore I thought it necessary to exhort the brethren, that they would go before unto you, and make up beforehand your bounty, whereof ye had notice before, that the same might be ready, as a matter of bounty, and not as of covetousness.
2COR|9|6|But this I say, He which soweth sparingly shall reap also sparingly; and he which soweth bountifully shall reap also bountifully.
2COR|9|7|Every man according as he purposeth in his heart, so let him give; not grudgingly, or of necessity: for God loveth a cheerful giver.
2COR|9|8|And God is able to make all grace abound toward you; that ye, always having all sufficiency in all things, may abound to every good work:
2COR|9|9|(As it is written, He hath dispersed abroad; he hath given to the poor: his righteousness remaineth for ever.
2COR|9|10|Now he that ministereth seed to the sower both minister bread for your food, and multiply your seed sown, and increase the fruits of your righteousness;)
2COR|9|11|Being enriched in every thing to all bountifulness, which causeth through us thanksgiving to God.
2COR|9|12|For the administration of this service not only supplieth the want of the saints, but is abundant also by many thanksgivings unto God;
2COR|9|13|Whiles by the experiment of this ministration they glorify God for your professed subjection unto the gospel of Christ, and for your liberal distribution unto them, and unto all men;
2COR|9|14|And by their prayer for you, which long after you for the exceeding grace of God in you.
2COR|9|15|Thanks be unto God for his unspeakable gift.
2COR|10|1|Now I Paul myself beseech you by the meekness and gentleness of Christ, who in presence am base among you, but being absent am bold toward you:
2COR|10|2|But I beseech you, that I may not be bold when I am present with that confidence, wherewith I think to be bold against some, which think of us as if we walked according to the flesh.
2COR|10|3|For though we walk in the flesh, we do not war after the flesh:
2COR|10|4|(For the weapons of our warfare are not carnal, but mighty through God to the pulling down of strong holds;)
2COR|10|5|Casting down imaginations, and every high thing that exalteth itself against the knowledge of God, and bringing into captivity every thought to the obedience of Christ;
2COR|10|6|And having in a readiness to revenge all disobedience, when your obedience is fulfilled.
2COR|10|7|Do ye look on things after the outward appearance? If any man trust to himself that he is Christ's, let him of himself think this again, that, as he is Christ's, even so are we Christ's.
2COR|10|8|For though I should boast somewhat more of our authority, which the Lord hath given us for edification, and not for your destruction, I should not be ashamed:
2COR|10|9|That I may not seem as if I would terrify you by letters.
2COR|10|10|For his letters, say they, are weighty and powerful; but his bodily presence is weak, and his speech contemptible.
2COR|10|11|Let such an one think this, that, such as we are in word by letters when we are absent, such will we be also in deed when we are present.
2COR|10|12|For we dare not make ourselves of the number, or compare ourselves with some that commend themselves: but they measuring themselves by themselves, and comparing themselves among themselves, are not wise.
2COR|10|13|But we will not boast of things without our measure, but according to the measure of the rule which God hath distributed to us, a measure to reach even unto you.
2COR|10|14|For we stretch not ourselves beyond our measure, as though we reached not unto you: for we are come as far as to you also in preaching the gospel of Christ:
2COR|10|15|Not boasting of things without our measure, that is, of other men's labours; but having hope, when your faith is increased, that we shall be enlarged by you according to our rule abundantly,
2COR|10|16|To preach the gospel in the regions beyond you, and not to boast in another man's line of things made ready to our hand.
2COR|10|17|But he that glorieth, let him glory in the Lord.
2COR|10|18|For not he that commendeth himself is approved, but whom the Lord commendeth.
2COR|11|1|Would to God ye could bear with me a little in my folly: and indeed bear with me.
2COR|11|2|For I am jealous over you with godly jealousy: for I have espoused you to one husband, that I may present you as a chaste virgin to Christ.
2COR|11|3|But I fear, lest by any means, as the serpent beguiled Eve through his subtilty, so your minds should be corrupted from the simplicity that is in Christ.
2COR|11|4|For if he that cometh preacheth another Jesus, whom we have not preached, or if ye receive another spirit, which ye have not received, or another gospel, which ye have not accepted, ye might well bear with him.
2COR|11|5|For I suppose I was not a whit behind the very chiefest apostles.
2COR|11|6|But though I be rude in speech, yet not in knowledge; but we have been throughly made manifest among you in all things.
2COR|11|7|Have I committed an offence in abasing myself that ye might be exalted, because I have preached to you the gospel of God freely?
2COR|11|8|I robbed other churches, taking wages of them, to do you service.
2COR|11|9|And when I was present with you, and wanted, I was chargeable to no man: for that which was lacking to me the brethren which came from Macedonia supplied: and in all things I have kept myself from being burdensome unto you, and so will I keep myself.
2COR|11|10|As the truth of Christ is in me, no man shall stop me of this boasting in the regions of Achaia.
2COR|11|11|Wherefore? because I love you not? God knoweth.
2COR|11|12|But what I do, that I will do, that I may cut off occasion from them which desire occasion; that wherein they glory, they may be found even as we.
2COR|11|13|For such are false apostles, deceitful workers, transforming themselves into the apostles of Christ.
2COR|11|14|And no marvel; for Satan himself is transformed into an angel of light.
2COR|11|15|Therefore it is no great thing if his ministers also be transformed as the ministers of righteousness; whose end shall be according to their works.
2COR|11|16|I say again, Let no man think me a fool; if otherwise, yet as a fool receive me, that I may boast myself a little.
2COR|11|17|That which I speak, I speak it not after the Lord, but as it were foolishly, in this confidence of boasting.
2COR|11|18|Seeing that many glory after the flesh, I will glory also.
2COR|11|19|For ye suffer fools gladly, seeing ye yourselves are wise.
2COR|11|20|For ye suffer, if a man bring you into bondage, if a man devour you, if a man take of you, if a man exalt himself, if a man smite you on the face.
2COR|11|21|I speak as concerning reproach, as though we had been weak. Howbeit whereinsoever any is bold, (I speak foolishly,) I am bold also.
2COR|11|22|Are they Hebrews? so am I. Are they Israelites? so am I. Are they the seed of Abraham? so am I.
2COR|11|23|Are they ministers of Christ? (I speak as a fool) I am more; in labours more abundant, in stripes above measure, in prisons more frequent, in deaths oft.
2COR|11|24|Of the Jews five times received I forty stripes save one.
2COR|11|25|Thrice was I beaten with rods, once was I stoned, thrice I suffered shipwreck, a night and a day I have been in the deep;
2COR|11|26|In journeyings often, in perils of waters, in perils of robbers, in perils by mine own countrymen, in perils by the heathen, in perils in the city, in perils in the wilderness, in perils in the sea, in perils among false brethren;
2COR|11|27|In weariness and painfulness, in watchings often, in hunger and thirst, in fastings often, in cold and nakedness.
2COR|11|28|Beside those things that are without, that which cometh upon me daily, the care of all the churches.
2COR|11|29|Who is weak, and I am not weak? who is offended, and I burn not?
2COR|11|30|If I must needs glory, I will glory of the things which concern mine infirmities.
2COR|11|31|The God and Father of our Lord Jesus Christ, which is blessed for evermore, knoweth that I lie not.
2COR|11|32|In Damascus the governor under Aretas the king kept the city of the Damascenes with a garrison, desirous to apprehend me:
2COR|11|33|And through a window in a basket was I let down by the wall, and escaped his hands.
2COR|12|1|It is not expedient for me doubtless to glory. I will come to visions and revelations of the Lord.
2COR|12|2|I knew a man in Christ above fourteen years ago, (whether in the body, I cannot tell; or whether out of the body, I cannot tell: God knoweth;) such an one caught up to the third heaven.
2COR|12|3|And I knew such a man, (whether in the body, or out of the body, I cannot tell: God knoweth;)
2COR|12|4|How that he was caught up into paradise, and heard unspeakable words, which it is not lawful for a man to utter.
2COR|12|5|Of such an one will I glory: yet of myself I will not glory, but in mine infirmities.
2COR|12|6|For though I would desire to glory, I shall not be a fool; for I will say the truth: but now I forbear, lest any man should think of me above that which he seeth me to be, or that he heareth of me.
2COR|12|7|And lest I should be exalted above measure through the abundance of the revelations, there was given to me a thorn in the flesh, the messenger of Satan to buffet me, lest I should be exalted above measure.
2COR|12|8|For this thing I besought the Lord thrice, that it might depart from me.
2COR|12|9|And he said unto me, My grace is sufficient for thee: for my strength is made perfect in weakness. Most gladly therefore will I rather glory in my infirmities, that the power of Christ may rest upon me.
2COR|12|10|Therefore I take pleasure in infirmities, in reproaches, in necessities, in persecutions, in distresses for Christ's sake: for when I am weak, then am I strong.
2COR|12|11|I am become a fool in glorying; ye have compelled me: for I ought to have been commended of you: for in nothing am I behind the very chiefest apostles, though I be nothing.
2COR|12|12|Truly the signs of an apostle were wrought among you in all patience, in signs, and wonders, and mighty deeds.
2COR|12|13|For what is it wherein ye were inferior to other churches, except it be that I myself was not burdensome to you? forgive me this wrong.
2COR|12|14|Behold, the third time I am ready to come to you; and I will not be burdensome to you: for I seek not your's but you: for the children ought not to lay up for the parents, but the parents for the children.
2COR|12|15|And I will very gladly spend and be spent for you; though the more abundantly I love you, the less I be loved.
2COR|12|16|But be it so, I did not burden you: nevertheless, being crafty, I caught you with guile.
2COR|12|17|Did I make a gain of you by any of them whom I sent unto you?
2COR|12|18|I desired Titus, and with him I sent a brother. Did Titus make a gain of you? walked we not in the same spirit? walked we not in the same steps?
2COR|12|19|Again, think ye that we excuse ourselves unto you? we speak before God in Christ: but we do all things, dearly beloved, for your edifying.
2COR|12|20|For I fear, lest, when I come, I shall not find you such as I would, and that I shall be found unto you such as ye would not: lest there be debates, envyings, wraths, strifes, backbitings, whisperings, swellings, tumults:
2COR|12|21|And lest, when I come again, my God will humble me among you, and that I shall bewail many which have sinned already, and have not repented of the uncleanness and fornication and lasciviousness which they have committed.
2COR|13|1|This is the third time I am coming to you. In the mouth of two or three witnesses shall every word be established.
2COR|13|2|I told you before, and foretell you, as if I were present, the second time; and being absent now I write to them which heretofore have sinned, and to all other, that, if I come again, I will not spare:
2COR|13|3|Since ye seek a proof of Christ speaking in me, which to you-ward is not weak, but is mighty in you.
2COR|13|4|For though he was crucified through weakness, yet he liveth by the power of God. For we also are weak in him, but we shall live with him by the power of God toward you.
2COR|13|5|Examine yourselves, whether ye be in the faith; prove your own selves. Know ye not your own selves, how that Jesus Christ is in you, except ye be reprobates?
2COR|13|6|But I trust that ye shall know that we are not reprobates.
2COR|13|7|Now I pray to God that ye do no evil; not that we should appear approved, but that ye should do that which is honest, though we be as reprobates.
2COR|13|8|For we can do nothing against the truth, but for the truth.
2COR|13|9|For we are glad, when we are weak, and ye are strong: and this also we wish, even your perfection.
2COR|13|10|Therefore I write these things being absent, lest being present I should use sharpness, according to the power which the Lord hath given me to edification, and not to destruction.
2COR|13|11|Finally, brethren, farewell. Be perfect, be of good comfort, be of one mind, live in peace; and the God of love and peace shall be with you.
2COR|13|12|Greet one another with an holy kiss.
2COR|13|13|All the saints salute you.
2COR|13|14|The grace of the Lord Jesus Christ, and the love of God, and the communion of the Holy Ghost, be with you all. Amen.
