JAS|1|1|Иаков, раб Бога и Господа Иисуса Христа, двенадцати коленам, находящимся в рассеянии, – радоваться.
JAS|1|2|С великою радостью принимайте, братия мои, когда впадаете в различные искушения,
JAS|1|3|зная, что испытание вашей веры производит терпение;
JAS|1|4|терпение же должно иметь совершенное действие, чтобы вы были совершенны во всей полноте, без всякого недостатка.
JAS|1|5|Если же у кого из вас недостает мудрости, да просит у Бога, дающего всем просто и без упреков, – и дастся ему.
JAS|1|6|Но да просит с верою, нимало не сомневаясь, потому что сомневающийся подобен морской волне, ветром поднимаемой и развеваемой.
JAS|1|7|Да не думает такой человек получить что–нибудь от Господа.
JAS|1|8|Человек с двоящимися мыслями не тверд во всех путях своих.
JAS|1|9|Да хвалится брат униженный высотою своею,
JAS|1|10|а богатый – унижением своим, потому что он прейдет, как цвет на траве.
JAS|1|11|Восходит солнце, [настает] зной, и зноем иссушает траву, цвет ее опадает, исчезает красота вида ее; так увядает и богатый в путях своих.
JAS|1|12|Блажен человек, который переносит искушение, потому что, быв испытан, он получит венец жизни, который обещал Господь любящим Его.
JAS|1|13|В искушении никто не говори: Бог меня искушает; потому что Бог не искушается злом и Сам не искушает никого,
JAS|1|14|но каждый искушается, увлекаясь и обольщаясь собственною похотью;
JAS|1|15|похоть же, зачав, рождает грех, а сделанный грех рождает смерть.
JAS|1|16|Не обманывайтесь, братия мои возлюбленные.
JAS|1|17|Всякое даяние доброе и всякий дар совершенный нисходит свыше, от Отца светов, у Которого нет изменения и ни тени перемены.
JAS|1|18|Восхотев, родил Он нас словом истины, чтобы нам быть некоторым начатком Его созданий.
JAS|1|19|Итак, братия мои возлюбленные, всякий человек да будет скор на слышание, медлен на слова, медлен на гнев,
JAS|1|20|ибо гнев человека не творит правды Божией.
JAS|1|21|Посему, отложив всякую нечистоту и остаток злобы, в кротости примите насаждаемое слово, могущее спасти ваши души.
JAS|1|22|Будьте же исполнители слова, а не слышатели только, обманывающие самих себя.
JAS|1|23|Ибо, кто слушает слово и не исполняет, тот подобен человеку, рассматривающему природные черты лица своего в зеркале:
JAS|1|24|он посмотрел на себя, отошел и тотчас забыл, каков он.
JAS|1|25|Но кто вникнет в закон совершенный, [закон] свободы, и пребудет в нем, тот, будучи не слушателем забывчивым, но исполнителем дела, блажен будет в своем действии.
JAS|1|26|Если кто из вас думает, что он благочестив, и не обуздывает своего языка, но обольщает свое сердце, у того пустое благочестие.
JAS|1|27|Чистое и непорочное благочестие пред Богом и Отцем есть то, чтобы призирать сирот и вдов в их скорбях и хранить себя неоскверненным от мира.
JAS|2|1|Братия мои! имейте веру в Иисуса Христа нашего Господа славы, не взирая на лица.
JAS|2|2|Ибо, если в собрание ваше войдет человек с золотым перстнем, в богатой одежде, войдет же и бедный в скудной одежде,
JAS|2|3|и вы, смотря на одетого в богатую одежду, скажете ему: тебе хорошо сесть здесь, а бедному скажете: ты стань там, или садись здесь, у ног моих, –
JAS|2|4|то не пересуживаете ли вы в себе и не становитесь ли судьями с худыми мыслями?
JAS|2|5|Послушайте, братия мои возлюбленные: не бедных ли мира избрал Бог быть богатыми верою и наследниками Царствия, которое Он обещал любящим Его?
JAS|2|6|А вы презрели бедного. Не богатые ли притесняют вас, и не они ли влекут вас в суды?
JAS|2|7|Не они ли бесславят доброе имя, которым вы называетесь?
JAS|2|8|Если вы исполняете закон царский, по Писанию: возлюби ближнего твоего, как себя самого, – хорошо делаете.
JAS|2|9|Но если поступаете с лицеприятием, то грех делаете, и перед законом оказываетесь преступниками.
JAS|2|10|Кто соблюдает весь закон и согрешит в одном чем–нибудь, тот становится виновным во всем.
JAS|2|11|Ибо Тот же, Кто сказал: не прелюбодействуй, сказал и: не убей; посему, если ты не прелюбодействуешь, но убьешь, то ты также преступник закона.
JAS|2|12|Так говорите и так поступайте, как имеющие быть судимы по закону свободы.
JAS|2|13|Ибо суд без милости не оказавшему милости; милость превозносится над судом.
JAS|2|14|Что пользы, братия мои, если кто говорит, что он имеет веру, а дел не имеет? может ли эта вера спасти его?
JAS|2|15|Если брат или сестра наги и не имеют дневного пропитания,
JAS|2|16|а кто–нибудь из вас скажет им: "идите с миром, грейтесь и питайтесь", но не даст им потребного для тела: что пользы?
JAS|2|17|Так и вера, если не имеет дел, мертва сама по себе.
JAS|2|18|Но скажет кто–нибудь: "ты имеешь веру, а я имею дела": покажи мне веру твою без дел твоих, а я покажу тебе веру мою из дел моих.
JAS|2|19|Ты веруешь, что Бог един: хорошо делаешь; и бесы веруют, и трепещут.
JAS|2|20|Но хочешь ли знать, неосновательный человек, что вера без дел мертва?
JAS|2|21|Не делами ли оправдался Авраам, отец наш, возложив на жертвенник Исаака, сына своего?
JAS|2|22|Видишь ли, что вера содействовала делам его, и делами вера достигла совершенства?
JAS|2|23|И исполнилось слово Писания: "веровал Авраам Богу, и это вменилось ему в праведность, и он наречен другом Божиим".
JAS|2|24|Видите ли, что человек оправдывается делами, а не верою только?
JAS|2|25|Подобно и Раав блудница не делами ли оправдалась, приняв соглядатаев и отпустив их другим путем?
JAS|2|26|Ибо, как тело без духа мертво, так и вера без дел мертва.
JAS|3|1|Братия мои! не многие делайтесь учителями, зная, что мы подвергнемся большему осуждению,
JAS|3|2|ибо все мы много согрешаем. Кто не согрешает в слове, тот человек совершенный, могущий обуздать и все тело.
JAS|3|3|Вот, мы влагаем удила в рот коням, чтобы они повиновались нам, и управляем всем телом их.
JAS|3|4|Вот, и корабли, как ни велики они и как ни сильными ветрами носятся, небольшим рулем направляются, куда хочет кормчий;
JAS|3|5|так и язык – небольшой член, но много делает. Посмотри, небольшой огонь как много вещества зажигает!
JAS|3|6|И язык – огонь, прикраса неправды; язык в таком положении находится между членами нашими, что оскверняет все тело и воспаляет круг жизни, будучи сам воспаляем от геенны.
JAS|3|7|Ибо всякое естество зверей и птиц, пресмыкающихся и морских животных укрощается и укрощено естеством человеческим,
JAS|3|8|а язык укротить никто из людей не может: это – неудержимое зло; он исполнен смертоносного яда.
JAS|3|9|Им благословляем Бога и Отца, и им проклинаем человеков, сотворенных по подобию Божию.
JAS|3|10|Из тех же уст исходит благословение и проклятие: не должно, братия мои, сему так быть.
JAS|3|11|Течет ли из одного отверстия источника сладкая и горькая [вода]?
JAS|3|12|Не может, братия мои, смоковница приносить маслины или виноградная лоза смоквы. Также и один источник не [может] изливать соленую и сладкую воду.
JAS|3|13|Мудр ли и разумен кто из вас, докажи это на самом деле добрым поведением с мудрою кротостью.
JAS|3|14|Но если в вашем сердце вы имеете горькую зависть и сварливость, то не хвалитесь и не лгите на истину.
JAS|3|15|Это не есть мудрость, нисходящая свыше, но земная, душевная, бесовская,
JAS|3|16|ибо где зависть и сварливость, там неустройство и все худое.
JAS|3|17|Но мудрость, сходящая свыше, во–первых, чиста, потом мирна, скромна, послушлива, полна милосердия и добрых плодов, беспристрастна и нелицемерна.
JAS|3|18|Плод же правды в мире сеется у тех, которые хранят мир.
JAS|4|1|Откуда у вас вражды и распри? не отсюда ли, от вожделений ваших, воюющих в членах ваших?
JAS|4|2|Желаете – и не имеете; убиваете и завидуете – и не можете достигнуть; препираетесь и враждуете – и не имеете, потому что не просите.
JAS|4|3|Просите, и не получаете, потому что просите не на добро, а чтобы употребить для ваших вожделений.
JAS|4|4|Прелюбодеи и прелюбодейцы! не знаете ли, что дружба с миром есть вражда против Бога? Итак, кто хочет быть другом миру, тот становится врагом Богу.
JAS|4|5|Или вы думаете, что напрасно говорит Писание: "до ревности любит дух, живущий в нас"?
JAS|4|6|Но тем большую дает благодать; посему и сказано: Бог гордым противится, а смиренным дает благодать.
JAS|4|7|Итак покоритесь Богу; противостаньте диаволу, и убежит от вас.
JAS|4|8|Приблизьтесь к Богу, и приблизится к вам; очистите руки, грешники, исправьте сердца, двоедушные.
JAS|4|9|Сокрушайтесь, плачьте и рыдайте; смех ваш да обратится в плач, и радость – в печаль.
JAS|4|10|Смиритесь пред Господом, и вознесет вас.
JAS|4|11|Не злословьте друг друга, братия: кто злословит брата или судит брата своего, того злословит закон и судит закон; а если ты судишь закон, то ты не исполнитель закона, но судья.
JAS|4|12|Един Законодатель и Судия, могущий спасти и погубить; а ты кто, который судишь другого?
JAS|4|13|Теперь послушайте вы, говорящие: "сегодня или завтра отправимся в такой–то город, и проживем там один год, и будем торговать и получать прибыль";
JAS|4|14|вы, которые не знаете, что случится завтра: ибо что такое жизнь ваша? пар, являющийся на малое время, а потом исчезающий.
JAS|4|15|Вместо того, чтобы вам говорить: "если угодно будет Господу и живы будем, то сделаем то или другое", –
JAS|4|16|вы, по своей надменности, тщеславитесь: всякое такое тщеславие есть зло.
JAS|4|17|Итак, кто разумеет делать добро и не делает, тому грех.
JAS|5|1|Послушайте вы, богатые: плачьте и рыдайте о бедствиях ваших, находящих на вас.
JAS|5|2|Богатство ваше сгнило, и одежды ваши изъедены молью.
JAS|5|3|Золото ваше и серебро изоржавело, и ржавчина их будет свидетельством против вас и съест плоть вашу, как огонь: вы собрали себе сокровище на последние дни.
JAS|5|4|Вот, плата, удержанная вами у работников, пожавших поля ваши, вопиет, и вопли жнецов дошли до слуха Господа Саваофа.
JAS|5|5|Вы роскошествовали на земле и наслаждались; напитали сердца ваши, как бы на день заклания.
JAS|5|6|Вы осудили, убили Праведника; Он не противился вам.
JAS|5|7|Итак, братия, будьте долготерпеливы до пришествия Господня. Вот, земледелец ждет драгоценного плода от земли и для него терпит долго, пока получит дождь ранний и поздний.
JAS|5|8|Долготерпите и вы, укрепите сердца ваши, потому что пришествие Господне приближается.
JAS|5|9|Не сетуйте, братия, друг на друга, чтобы не быть осужденными: вот, Судия стоит у дверей.
JAS|5|10|В пример злострадания и долготерпения возьмите, братия мои, пророков, которые говорили именем Господним.
JAS|5|11|Вот, мы ублажаем тех, которые терпели. Вы слышали о терпении Иова и видели конец [оного] от Господа, ибо Господь весьма милосерд и сострадателен.
JAS|5|12|Прежде же всего, братия мои, не клянитесь ни небом, ни землею, и никакою другою клятвою, но да будет у вас: "да, да" и "нет, нет", дабы вам не подпасть осуждению.
JAS|5|13|Злостраждет ли кто из вас, пусть молится. Весел ли кто, пусть поет псалмы.
JAS|5|14|Болен ли кто из вас, пусть призовет пресвитеров Церкви, и пусть помолятся над ним, помазав его елеем во имя Господне.
JAS|5|15|И молитва веры исцелит болящего, и восставит его Господь; и если он соделал грехи, простятся ему.
JAS|5|16|Признавайтесь друг пред другом в проступках и молитесь друг за друга, чтобы исцелиться: много может усиленная молитва праведного.
JAS|5|17|Илия был человек, подобный нам, и молитвою помолился, чтобы не было дождя: и не было дождя на землю три года и шесть месяцев.
JAS|5|18|И опять помолился: и небо дало дождь, и земля произрастила плод свой.
JAS|5|19|Братия! если кто из вас уклонится от истины, и обратит кто его,
JAS|5|20|пусть тот знает, что обративший грешника от ложного пути его спасет душу от смерти и покроет множество грехов.
