2SAM|1|1|扫罗 死后， 大卫 击杀 亚玛力 人回来，在 洗革拉 住了两天。
2SAM|1|2|第三天，看哪，有一人从 扫罗 的营里出来，衣服撕裂，头蒙灰尘，到 大卫 面前伏地叩拜。
2SAM|1|3|大卫 对他说：“你从哪里来？”他说：“我从 以色列 的营里逃来。”
2SAM|1|4|大卫 又对他说：“事情怎么样？请你告诉我。”他说：“士兵从阵上逃跑，也有许多士兵仆倒死亡， 扫罗 和他儿子 约拿单 也死了。”
2SAM|1|5|大卫 问报信的青年说：“你怎么知道 扫罗 和他儿子 约拿单 死了呢？”
2SAM|1|6|报信的青年说：“我恰巧到 基利波山 ，看哪， 扫罗 靠在自己的枪上，看哪，有战车、骑兵紧紧地追他。
2SAM|1|7|他回头看见我，就呼叫我。我说：‘我在这里。’
2SAM|1|8|他问我说：‘你是什么人？’我说：‘我是 亚玛力 人。’
2SAM|1|9|他对我说：‘请你站到我这里来，把我杀死，因为我非常痛苦，只剩下一口气。’
2SAM|1|10|我就站到他那里，杀了他，因为我知道他一倒下就活不了。然后，我把他头上的冠冕和臂上的镯子拿到我主这里来。”
2SAM|1|11|大卫 就抓着自己的衣服，把衣服撕裂，所有跟随他的人也都如此。
2SAM|1|12|他们为 扫罗 和他儿子 约拿单 ，以及耶和华的百姓和 以色列 家的人悲哀哭泣，禁食到晚上，因为他们都倒在刀下。
2SAM|1|13|大卫 问报信的青年说：“你是哪里人？”他说：“我是一个寄居者的儿子，是 亚玛力 人。”
2SAM|1|14|大卫 对他说：“你动手杀害耶和华的受膏者，怎么不畏惧呢？”
2SAM|1|15|大卫 叫了一个仆人来，说：“来，杀了他！”仆人击杀他，他就死了。
2SAM|1|16|大卫 对他说：“你的血归到你自己头上，因为你亲口作证控诉自己，说：‘我杀了耶和华的受膏者。’”
2SAM|1|17|大卫 作了这首哀歌，哀悼 扫罗 和他儿子 约拿单 ，
2SAM|1|18|并吩咐人把这首“弓歌”教导 犹大 人，看哪，它写在《雅煞珥书》上：
2SAM|1|19|以色列 啊，尊荣者在你的高处被杀！ 大英雄竟然仆倒！
2SAM|1|20|不要在 迦特 报告， 不要在 亚实基伦 街上传扬， 免得 非利士 的女子欢喜， 免得未受割礼之人的女子欢乐。
2SAM|1|21|基利波山 哪，愿你那里没有雨，没有露！ 愿你的田地无土产可作供物！ 因为英雄的盾牌在那里受辱， 扫罗 的盾牌没有抹油。
2SAM|1|22|在被杀者的血前， 在勇士的脂肪前， 约拿单 的弓绝不退缩， 扫罗 的刀断不虚回。
2SAM|1|23|扫罗 和 约拿单 生时相悦相爱， 死时也不分离。 他们比鹰更快， 比狮子还强。
2SAM|1|24|以色列 的女子啊，当为 扫罗 哭泣！ 他曾使你们穿朱红色的美衣， 使你们衣服有黄金的妆饰。
2SAM|1|25|英雄竟然在阵上仆倒！ 约拿单 竟然在你的高处被杀！
2SAM|1|26|我兄 约拿单 哪，我为你悲伤！ 我甚喜爱你！ 你对我的爱何等奇妙， 过于妇女的爱情。
2SAM|1|27|英雄竟然仆倒！ 兵器竟然废弃！
2SAM|2|1|此后， 大卫 求问耶和华说：“我可以上 犹大 的一个城去吗？”耶和华对他说：“可以上去。” 大卫 说：“我上哪一个城去呢？”耶和华说：“ 希伯仑 。”
2SAM|2|2|于是 大卫 和他的两个妻子，一个是 耶斯列 人 亚希暖 ，一个是作过 迦密 人 拿八 妻子的 亚比该 ，都上那里去了。
2SAM|2|3|大卫 也把跟随他的人和他们各人的眷属一同带上去，住在 希伯仑 的城镇中。
2SAM|2|4|犹大 人来，在那里膏 大卫 作 犹大 家的王。 有人告诉 大卫 说：“埋葬 扫罗 的是 基列 的 雅比 人。”
2SAM|2|5|大卫 就派使者到 基列 的 雅比 人那里，对他们说：“愿耶和华赐福给你们！因为你们忠心对待你们的主 扫罗 ，埋葬了他。
2SAM|2|6|你们既做了这事，愿耶和华以慈爱和信实待你们，我也要为此厚待你们。
2SAM|2|7|现在，你们的主 扫罗 死了， 犹大 家也已经膏我作他们的王，你们的手要坚强，要作英勇的人。”
2SAM|2|8|扫罗 军队的元帅， 尼珥 的儿子 押尼珥 ，曾将 扫罗 的儿子 伊施．波设 带过河，到 玛哈念 ，
2SAM|2|9|立他作王，治理 基列 、 亚书利 、 耶斯列 、 以法莲 、 便雅悯 和 以色列 众人。
2SAM|2|10|扫罗 的儿子 伊施．波设 登基的时候年四十岁，作 以色列 王二年，但是 犹大 家却随从 大卫 。
2SAM|2|11|大卫 在 希伯仑 作 犹大 家的王，共七年六个月。
2SAM|2|12|尼珥 的儿子 押尼珥 和 扫罗 的儿子 伊施．波设 的仆人从 玛哈念 出来，往 基遍 去。
2SAM|2|13|洗鲁雅 的儿子 约押 和 大卫 的仆人也出来，在 基遍 池旁与他们相遇；一队坐在池的这边，一队坐在池的那边。
2SAM|2|14|押尼珥 对 约押 说：“让年轻人起来，在我们面前较量一下吧！” 约押 说：“让他们起来吧。”
2SAM|2|15|他们就起来，点了人数过来：属 扫罗 儿子 伊施．波设 的有 便雅悯 人十二名， 大卫 的仆人也有十二名。
2SAM|2|16|每人抓住对方的头，用刀刺对方的肋旁，一同仆倒。所以，那地叫做 希利甲．哈素林 ，就在 基遍 。
2SAM|2|17|那日战况激烈， 押尼珥 和 以色列 人败在 大卫 的仆人面前。
2SAM|2|18|在那里有 洗鲁雅 的三个儿子： 约押 、 亚比筛 、 亚撒黑 。 亚撒黑 的脚快如野地里的羚羊；
2SAM|2|19|亚撒黑 追赶 押尼珥 ，直追赶他不偏左右。
2SAM|2|20|押尼珥 回头说：“ 亚撒黑 ，是你吗？”他说：“是我。”
2SAM|2|21|押尼珥 对他说：“你转左或转右，去抓一个年轻人，剥去他的战衣吧。” 亚撒黑 却不肯转开而不追赶他。
2SAM|2|22|押尼珥 又对 亚撒黑 说：“转开，不要再追我了！我何必把你击杀在地上呢？我若杀了你，怎么有脸见你哥哥 约押 呢？”
2SAM|2|23|亚撒黑 仍不肯转开， 押尼珥 就用回马枪 刺入他的肚腹，甚至枪从背后穿出， 亚撒黑 就仆倒在那里，当场死了。众人赶到 亚撒黑 仆倒而死的地方，就都站住。
2SAM|2|24|约押 和 亚比筛 追赶 押尼珥 。日落的时候，他们到了通往 基遍 旷野的路旁， 基亚 对面的 亚玛山 。
2SAM|2|25|便雅悯 人聚集在 押尼珥 后面，成为一队，站在一座山顶上。
2SAM|2|26|押尼珥 呼叫 约押 说：“刀剑岂可永远吞噬呢？你岂不知，结局必是痛苦的吗？你要等到何时才叫百姓回去，不追赶他们的弟兄呢？”
2SAM|2|27|约押 说：“我指着永生的上帝起誓：你若没有这么说，百姓就必继续追赶弟兄，直到早晨 。”
2SAM|2|28|于是 约押 吹角，众百姓就站住，不再追赶 以色列 人，也不再打仗了。
2SAM|2|29|押尼珥 和他的人整夜行过 亚拉巴 。他们过了 约旦河 ，走过 毕伦 ，到了 玛哈念 。
2SAM|2|30|约押 追赶 押尼珥 回来，聚集众百姓， 大卫 的仆人中缺少了十九个人和 亚撒黑 。
2SAM|2|31|但 大卫 的仆人杀了 押尼珥 的人， 便雅悯 人三百六十名。
2SAM|2|32|他们把 亚撒黑 送到 伯利恒 ，葬在他父亲的坟墓里。 约押 和他的人走了一整夜，天亮的时候他们才到 希伯仑 。
2SAM|3|1|扫罗 家和 大卫 家争战许久。 大卫 家日见强盛， 扫罗 家却日见衰弱。
2SAM|3|2|大卫 在 希伯仑 生了几个儿子：长子 暗嫩 是 耶斯列 人 亚希暖 所生的；
2SAM|3|3|次子 基利押 是作过 迦密 人 拿八 的妻子 亚比该 所生的；三子 押沙龙 是 基述 王 达买 的女儿 玛迦 所生的；
2SAM|3|4|四子 亚多尼雅 是 哈及 所生的；五子 示法提雅 是 亚比她 所生的；
2SAM|3|5|六子 以特念 是 大卫 的妻子 以格拉 所生的。 大卫 这六个儿子都是在 希伯仑 生的。
2SAM|3|6|扫罗 家和 大卫 家争战的时候， 押尼珥 在 扫罗 家大有权势。
2SAM|3|7|扫罗 有一妃子，名叫 利斯巴 ，是 爱亚 的女儿。一日， 伊施．波设 对 押尼珥 说：“你为什么与我父的妃子同寝呢？”
2SAM|3|8|押尼珥 因 伊施．波设 的话非常生气，说：“我岂是狗的头，向着 犹大 呢？我今日忠心对待你父 扫罗 的家和他的弟兄、朋友，不将你交在 大卫 手里，今日你竟为这妇人责备我吗？
2SAM|3|9|愿上帝重重惩罚 押尼珥 ！我要照着耶和华起誓应许 大卫 的话为他成就，
2SAM|3|10|废去 扫罗 家的国度，建立 大卫 的王位，使他治理 以色列 和 犹大 ，从 但 直到 别是巴 。”
2SAM|3|11|伊施．波设 惧怕 押尼珥 ，一句话也不能回答。
2SAM|3|12|押尼珥 派使者到 大卫 所在的地方 ，说：“这地归谁呢？”又说：“你与我立约，看哪，我必帮助你，使全 以色列 都拥护你。”
2SAM|3|13|大卫 说：“好！我与你立约。但有一件事我要求你，你来见我面的时候，除非把 扫罗 的女儿 米甲 带来，就不必来见我的面了。”
2SAM|3|14|大卫 派使者到 扫罗 的儿子 伊施．波设 那里，说：“你要把我的妻子 米甲 归还我；她是我从前用一百 非利士 人的包皮所聘定的。”
2SAM|3|15|伊施．波设 就派人去，把 米甲 从 拉亿 的儿子，她丈夫 帕铁 那里带来。
2SAM|3|16|米甲 的丈夫跟着她，一面走一面哭，直跟到 巴户琳 。 押尼珥 对他说：“你回去吧！” 帕铁 就回去了。
2SAM|3|17|押尼珥 与 以色列 长老商议，说：“从前你们企盼 大卫 作王治理你们，
2SAM|3|18|现在你们可以这样做了。因为耶和华曾论到 大卫 说：‘我必藉我仆人 大卫 的手，救我民 以色列 脱离 非利士 人和众仇敌的手。’”
2SAM|3|19|押尼珥 也说给 便雅悯 人听。 押尼珥 又到 希伯仑 ，把 以色列 人和 便雅悯 全家所看为好的，说给 大卫 听。
2SAM|3|20|押尼珥 带着二十个人来到 希伯仑大卫 那里， 大卫 就为 押尼珥 和他带来的人摆设宴席。
2SAM|3|21|押尼珥 对 大卫 说：“我要起身去召集全 以色列 ，来到我主我王这里，与你立约，你就可以照你的心愿作王，统治一切。”于是 大卫 送走 押尼珥 ，他就平安地去了。
2SAM|3|22|看哪， 大卫 的仆人和 约押 突击回来，带回许多掠物。那时 押尼珥 不在 希伯仑大卫 那里，因 大卫 已经送他走，他也平安地去了。
2SAM|3|23|约押 和跟随他的全军到了，有人告诉 约押 说：“ 尼珥 的儿子 押尼珥 来到王这里，王送走他，他也平安地去了。”
2SAM|3|24|约押 到王那里，说：“你这是做什么呢？看哪， 押尼珥 来到你这里，你为何送他走，让他去了呢？
2SAM|3|25|你知道， 尼珥 的儿子 押尼珥 来，是要骗你，要打听你的出入，知道你一切所行的事。”
2SAM|3|26|约押 从 大卫 那里出来，派些使者去追 押尼珥 ，从 西拉井 那里带他回来， 大卫 却不知道。
2SAM|3|27|押尼珥 回到 希伯仑 ， 约押 领他到城门中间，要与他私下交谈，就在那里刺穿了他的肚腹。他就死了，因为他流了 约押 兄弟 亚撒黑 的血。
2SAM|3|28|这事以后， 大卫 听见了，说：“流 尼珥 儿子 押尼珥 的血，我和我的国在耶和华面前永远是无辜的。
2SAM|3|29|愿这血归到 约押 头上和他父的全家；又愿 约押 家不断有患漏症的，长痲疯 的，架柺杖而行的 ，仆倒在刀下的，缺乏食物的。”
2SAM|3|30|约押 和他弟弟 亚比筛 杀了 押尼珥 ，是因为在 基遍 战争的时候， 押尼珥 杀了他们的弟弟 亚撒黑 。
2SAM|3|31|大卫 对 约押 和跟随他的众百姓说：“你们当撕裂衣服，腰束麻布，在 押尼珥 前面哀哭。” 大卫 王也跟在棺木后面。
2SAM|3|32|他们把 押尼珥 葬在 希伯仑 。王在 押尼珥 的墓旁放声大哭，众百姓也都哭了。
2SAM|3|33|王为 押尼珥 举哀，说： 押尼珥 怎么会像愚顽人一样地死呢？
2SAM|3|34|你手未曾被捆绑，脚未曾被脚镣锁住。 你仆倒，如仆倒在凶恶之子手下一样。 于是众百姓又为 押尼珥 哀哭。
2SAM|3|35|白天的时候，众百姓来劝 大卫 吃饭，但 大卫 起誓说：“我若在太阳未下山以前吃饭，或吃任何东西，愿上帝重重惩罚我！”
2SAM|3|36|众百姓知道了就看为好。凡王所做的，众百姓都看为好。
2SAM|3|37|那日， 以色列 众百姓才知道杀 尼珥 的儿子 押尼珥 并非出于王意。
2SAM|3|38|王对臣仆说：“你们岂不知今日在 以色列 中倒了一个作元帅的大人物吗？
2SAM|3|39|我虽然受膏为王，今日还是软弱。 洗鲁雅 的两个儿子，这些人比我强硬。愿耶和华照着恶人所行的恶报应他。”
2SAM|4|1|扫罗 的儿子 伊施．波设 听见 押尼珥 死在 希伯仑 ，手就发软，全 以色列 也都惊惶。
2SAM|4|2|扫罗 的儿子 伊施．波设 有两个军官，一个叫 巴拿 ，第二个叫 利甲 ，都是 便雅悯 支派 比录 人 临门 的儿子；因为 比录 也算是属于 便雅悯 的。
2SAM|4|3|比录 人先前逃到 基他音 ，在那里寄居，直到今日。
2SAM|4|4|扫罗 的儿子 约拿单 有一个儿子，名叫 米非波设 ，是瘸腿的。 扫罗 和 约拿单 的消息从 耶斯列 传来的时候，他才五岁。他的奶妈抱着他逃跑；因为跑得太急，孩子掉在地上，腿就瘸了。
2SAM|4|5|比录 人 临门 的两个儿子 利甲 和 巴拿 出去，天正热的时候到了 伊施．波设 的家。那时， 伊施．波设 在睡午觉。
2SAM|4|6|妇人进到房子中间，要取麦子。 利甲 和他的哥哥 巴拿 刺穿了 伊施．波设 的肚腹，然后逃跑了。
2SAM|4|7|他们进到房子的时候， 伊施．波设 正躺在卧房的床上，他们就把他杀死，割了他的首级，拿着首级在 亚拉巴 的路上走了一整夜。
2SAM|4|8|他们把 伊施．波设 的首级拿到 希伯仑 大卫 那里，对王说：“王的仇敌 扫罗 曾寻索你的性命。看哪，这是他儿子 伊施．波设 的首级；耶和华今日为我主我王在 扫罗 和他后裔身上报了仇。”
2SAM|4|9|大卫 回答 比录 人 临门 的儿子 利甲 和他哥哥 巴拿 说：“我指着救我性命脱离一切苦难、永生的耶和华起誓：
2SAM|4|10|从前有人告诉我说：‘看哪， 扫罗 死了。’他自以为报好消息，我就拿住他，把他杀在 洗革拉 ，作为他报消息的赏赐。
2SAM|4|11|更何况恶人把义人杀在他家的床上，我岂不从你们手中追讨他的血，从地上除灭你们吗？”
2SAM|4|12|于是 大卫 吩咐仆人把他们杀了，砍断他们的手脚，挂在 希伯仑 的池旁。然后，他们把 伊施．波设 的首级葬在 希伯仑押尼珥 的坟墓里。
2SAM|5|1|以色列 众支派来到 希伯仑 见 大卫 ，说：“看哪，我们是你的骨肉。
2SAM|5|2|从前 扫罗 作我们王的时候，率领 以色列 人出入的是你。耶和华也曾对你说：‘你必牧养我的百姓 以色列 ，你必作 以色列 的君王。’”
2SAM|5|3|于是 以色列 的众长老都来到 希伯仑 见王 。 大卫 在 希伯仑 ，在耶和华面前与他们立约，他们就膏 大卫 作 以色列 的王。
2SAM|5|4|大卫 登基的时候年三十岁，作王四十年。
2SAM|5|5|他在 希伯仑 作 犹大 王七年六个月，在 耶路撒冷 作 以色列 和 犹大 王三十三年。
2SAM|5|6|王和他的人到了 耶路撒冷 ，要攻打住那地方的 耶布斯 人。 耶布斯 人对 大卫 说：“你必不能进到这里，就是盲人、瘸子都可以把你击退。”就是说：“ 大卫 绝不能进到这里。”
2SAM|5|7|然而 大卫 攻取了 锡安 的堡垒，就是 大卫 的城。
2SAM|5|8|当日， 大卫 说：“谁攻打 耶布斯 人，就要从水道上去，攻打我心里所恨恶的 瘸子、盲人。”因此有人说：“盲人和瘸子不得进殿里去。”
2SAM|5|9|大卫 住在堡垒里，给它起名叫 大卫城 。 大卫 又从 米罗 往内，周围建筑。
2SAM|5|10|大卫 日见强大，耶和华－万军之上帝与他同在。
2SAM|5|11|推罗 王 希兰 派使者把香柏木运到 大卫 那里，又派木匠和石匠给 大卫 建造宫殿。
2SAM|5|12|大卫 知道耶和华坚立他作 以色列 王，又为自己百姓 以色列 的缘故，使他的国兴盛。
2SAM|5|13|大卫 离开 希伯仑 之后，在 耶路撒冷 又立后妃，又生儿女。
2SAM|5|14|在 耶路撒冷 所生的孩子的名字是 沙母亚 、 朔罢 、 拿单 、 所罗门 、
2SAM|5|15|益辖 、 以利书亚 、 尼斐 、 雅非亚 、
2SAM|5|16|以利沙玛 、 以利雅大 、 以利法列 。
2SAM|5|17|非利士 人听见 大卫 受膏作 以色列 王， 非利士 众人就上来寻索 大卫 。 大卫 听见了，就下到堡垒去。
2SAM|5|18|非利士 人来了，散布在 利乏音谷 。
2SAM|5|19|大卫 求问耶和华说：“我可以上去攻打 非利士 人吗？你将他们交在我手里吗？”耶和华对 大卫 说：“你可以上去，我必将 非利士 人交在你手里。”
2SAM|5|20|大卫 来到 巴力．毗拉心 ，在那里击败了 非利士 人。他说：“耶和华在我面前冲破敌人，如水冲破一样。”因此他称那地方为 巴力．毗拉心 。
2SAM|5|21|非利士 人把偶像抛弃在那里， 大卫 和他的人拿去了。
2SAM|5|22|非利士 人又上来，散布在 利乏音谷 。
2SAM|5|23|大卫 求问耶和华；耶和华说：“不要直上，要绕到他们后头，从桑树林对面攻打他们。
2SAM|5|24|你听见桑树梢上有脚步的声音，就要急速前去，因为那时耶和华已经出去，在你前头攻打 非利士 人的军队了。”
2SAM|5|25|大卫 就遵照耶和华所吩咐的去做，攻打 非利士 人，从 迦巴 直到 基色 。
2SAM|6|1|大卫 又聚集 以色列 中所有挑选的人，共三万名。
2SAM|6|2|大卫 起身，和跟随他的众百姓前往，要从 巴拉．犹大 那里将上帝的约柜接上来；这约柜是以坐在二基路伯上万军之耶和华的名所命名的。
2SAM|6|3|他们将上帝的约柜从山冈上 亚比拿达 的家里抬出来，放在新车上； 亚比拿达 的儿子 乌撒 和 亚希约 赶这新车。
2SAM|6|4|他们将上帝的约柜从山冈上 亚比拿达 家里抬出来 ， 亚希约 在约柜前行走。
2SAM|6|5|大卫 和 以色列 全家在耶和华面前，随着松木制造的各样乐器 和琴、瑟、鼓、钹、锣跳舞。
2SAM|6|6|到了 拿艮 的禾场，因为牛失前蹄 ， 乌撒 就伸手扶住上帝的约柜。
2SAM|6|7|耶和华的怒气向 乌撒 发作；上帝因这冒犯在那里击打他，他就死在那里，在上帝的约柜旁。
2SAM|6|8|大卫 因耶和华突然冲出撞死 乌撒 就生气，称那地方为 毗列斯．乌撒 ，直到今日。
2SAM|6|9|那日， 大卫 惧怕耶和华，说：“耶和华的约柜怎可到我这里来呢？”
2SAM|6|10|于是 大卫 不愿将耶和华的约柜接进 大卫城 他自己的地方，却转送到 迦特 人 俄别．以东 的家中。
2SAM|6|11|耶和华的约柜停在 迦特 人 俄别．以东 家中三个月，耶和华赐福给 俄别．以东 和他的全家。
2SAM|6|12|有人告诉 大卫 王说：“耶和华因约柜的缘故赐福给 俄别．以东 的家和一切属他的。” 大卫 就去，欢欢喜喜地将上帝的约柜从 俄别．以东 家中接上来，到 大卫城 里。
2SAM|6|13|抬耶和华约柜的人走了六步， 大卫 就献牛与肥畜为祭。
2SAM|6|14|大卫 穿着细麻布以弗得，在耶和华面前极力跳舞。
2SAM|6|15|这样， 大卫 和 以色列 全家欢呼吹角，将耶和华的约柜接了上来。
2SAM|6|16|耶和华的约柜进 大卫城 的时候， 扫罗 的女儿 米甲 从窗户里往外观看，见 大卫 王在耶和华面前踊跃跳舞，心里就轻视他。
2SAM|6|17|众人将耶和华的约柜请进去，安放在所预备的地方，就是 大卫 为它搭的帐幕中。 大卫 在耶和华面前献燔祭和平安祭。
2SAM|6|18|大卫 献完了燔祭和平安祭，就奉万军之耶和华的名祝福百姓，
2SAM|6|19|并且分给 以色列 众人，所有的百姓，无论男女，每人一个饼，一个枣子饼 ，一个葡萄饼。众人就各自回家去了。
2SAM|6|20|大卫 回去要为家里的人祝福， 扫罗 的女儿 米甲 出来迎接他，说：“ 以色列 王今日有好大的荣耀啊！他今日在臣仆的使女眼前露体，如同一个无赖赤身露体一样，”
2SAM|6|21|大卫 对 米甲 说：“这是在耶和华面前的。耶和华已拣选我，在你父和你父的全家之上，立我作耶和华百姓 以色列 的君王，所以我在耶和华面前跳舞，
2SAM|6|22|我也必更加卑微，自己看为低贱 。至于你所说的那些使女，她们反而尊重我。”
2SAM|6|23|扫罗 的女儿 米甲 ，直到死的那日没有孩子。
2SAM|7|1|王住在自己宫中，耶和华使他平静，不被四围的仇敌扰乱。
2SAM|7|2|王对 拿单 先知说：“你看，我住在香柏木的宫中，上帝的约柜却停在幔子里。”
2SAM|7|3|拿单 对王说：“你可以完全照你的心意去做，因为耶和华与你同在。”
2SAM|7|4|当夜耶和华的话临到 拿单 ，说：
2SAM|7|5|“你去对我仆人 大卫 说：‘耶和华如此说：你要建造殿宇给我居住吗？
2SAM|7|6|自从我领 以色列 人从 埃及 上来，直到今日，我未曾住过殿宇，却在会幕和帐幕中行走。
2SAM|7|7|凡我同 以色列 人所走的地方，我何曾向 以色列 任何一个领袖 ，就是我吩咐牧养我百姓 以色列 的，说过这话：你们为何不给我建造香柏木的殿宇呢？’
2SAM|7|8|现在，你要对我仆人 大卫这样 说：‘万军之耶和华如此说：我从羊圈中将你召来，叫你不再牧放羊群，立你作我百姓 以色列 的君王。
2SAM|7|9|你无论往哪里去，我都与你同在，剪除你所有的仇敌。我必使你得大名，好像世上伟人的名一样。
2SAM|7|10|我必为我百姓 以色列 选定一个地方，栽植他们，使他们住自己的地方，不再受搅扰；凶恶之子也不像从前那样苦待他们，
2SAM|7|11|并不像我命令士师治理我百姓 以色列 的日子。我必使你平静，不受任何仇敌搅扰，并且耶和华应许你，耶和华必为你建立家室。
2SAM|7|12|当你寿数满足、与你祖先同睡的时候，我必使你身所生的后裔接续你；我也必坚定他的国。
2SAM|7|13|他必为我的名建造殿宇，我必坚定他国度的王位，直到永远。
2SAM|7|14|我要作他的父，他要作我的子；他若犯了罪，我必用人的杖，用世人的鞭责罚他。
2SAM|7|15|但我的慈爱仍不离开他，像离开在你面前所废的 扫罗 一样。
2SAM|7|16|你的家和你的国必在你 面前永远坚立，你的王位也必坚定，直到永远。’”
2SAM|7|17|拿单 就按这一切话，照这一切异象告诉 大卫 。
2SAM|7|18|于是 大卫 王进去，坐在耶和华面前，说：“主耶和华啊，我是谁，我的家算什么，你竟带领我到这地步呢？
2SAM|7|19|主耶和华啊，这在你眼中还看为小，你又说到你仆人的家将来的情况。主耶和华啊，这岂是人的常理吗？
2SAM|7|20|大卫 还有什么可以对你说呢？主耶和华啊，你是知道你仆人的。
2SAM|7|21|你行这一切大事，使你的仆人明白，是因你应许的缘故，也照着你的心意。
2SAM|7|22|因此，主耶和华啊，你本为大；照我们耳中一切所听见的，没有可比你的，除你以外再没有上帝。
2SAM|7|23|谁像你的百姓 以色列 呢？上帝亲自去救赎世上的一国 ，作自己的子民，显出他的大名；为了你的地，从列国和他们的神明中，在你亲自从埃及赎出来的子民面前，为自己行了大而可畏的事 。
2SAM|7|24|你曾坚立你的百姓 以色列 作你的子民，直到永远；你－耶和华也作他们的上帝。
2SAM|7|25|现在，耶和华上帝啊，你所应许仆人和仆人家的话，求你坚定，直到永远；求你照你所说的而行。
2SAM|7|26|愿人永远尊你的名为大，说：‘万军之耶和华是治理 以色列 的上帝。’这样，你仆人 大卫 的家必在你面前坚立。
2SAM|7|27|万军之耶和华－ 以色列 的上帝啊，因你启示你的仆人说：‘我必为你建立家室’，所以仆人大胆向你如此祈祷。
2SAM|7|28|现在，主耶和华啊，惟有你是上帝！你的话是真实的，你也应许将这福气赐给仆人。
2SAM|7|29|现在，求你赐福给你仆人的家，可以永存在你面前。主耶和华啊，因为这是你所应许的。愿你的福分永远赐给你仆人的家，使之蒙福！”
2SAM|8|1|此后， 大卫 攻打 非利士 人，制伏了他们。 大卫 从 非利士 人手中夺取了京城的治理权 。
2SAM|8|2|他又攻打 摩押 人，使他们躺卧在地上，用绳来量，量二绳的杀了，量一绳的活着。 摩押 人就臣服 大卫 ，向他进贡。
2SAM|8|3|利合 的儿子 琐巴 王 哈大底谢 往 幼发拉底河 去，要夺回他的国权， 大卫 就攻打他，
2SAM|8|4|俘掳了他的骑兵一千七百人，步兵二万人。 大卫 把所有战马的蹄筋砍断，只留下一百辆战车。
2SAM|8|5|大马士革 的 亚兰 人来帮助 琐巴 王 哈大底谢 ， 大卫 杀了 亚兰 人二万二千。
2SAM|8|6|于是 大卫 在 大马士革 的 亚兰 设立军营， 亚兰 人就臣服 大卫 ，向他进贡。 大卫 无论往哪里去，耶和华都使他得胜。
2SAM|8|7|大卫夺了 哈大底谢 臣仆拥有的金盾牌，带到 耶路撒冷 。
2SAM|8|8|大卫 王又从 哈大底谢 的 比他 和 比罗他 二城夺取了许多的铜。
2SAM|8|9|哈马 王 陀以 听见 大卫 击败 哈大底谢 的全军，
2SAM|8|10|就派他儿子 约兰 到 大卫 王那里，向他请安，为他祝福，因他与 哈大底谢 争战，并且击败了他；原来 哈大底谢 与 陀以 常常争战。 约兰 手里带了金银铜的器皿来。
2SAM|8|11|大卫 王把这些器皿分别为圣，连同他制伏各国所分别为圣的金银，献给耶和华，
2SAM|8|12|就是从 亚兰 、 摩押 、 亚扪 人、 非利士 人、 亚玛力 人，以及从 利合 的儿子 琐巴 王 哈大底谢 所掠之物。
2SAM|8|13|大卫 得了名声。当他回来的时候，在 盐谷 击杀了一万八千 以东 人。
2SAM|8|14|大卫 在 以东 设立军营；他在全 以东 设立军营， 以东 人就都臣服他。 大卫 无论往哪里去，耶和华都使他得胜。
2SAM|8|15|大卫 作全 以色列 的王，又向众百姓秉公行义。
2SAM|8|16|洗鲁雅 的儿子 约押 作元帅； 亚希律 的儿子 约沙法 作史官；
2SAM|8|17|亚希突 的儿子 撒督 和 亚比亚他 的儿子 亚希米勒 作祭司； 西莱雅 作书记；
2SAM|8|18|耶何耶大 的儿子 比拿雅 管辖 基利提 人和 比利提 人。 大卫 的众子都作祭司。
2SAM|9|1|大卫 说：“ 扫罗 家还有剩下的人没有？我要因 约拿单 的缘故向他施恩。”
2SAM|9|2|扫罗 家有一个仆人名叫 洗巴 ，有人叫他来到 大卫 那里。王对他说：“你是 洗巴 吗？”他说：“仆人是。”
2SAM|9|3|王说：“ 扫罗 家还有没有剩下的人？我要照上帝的慈爱恩待他。” 洗巴 对王说：“还有 约拿单 的一个儿子，双腿是瘸的。”
2SAM|9|4|王对他说：“他在哪里？” 洗巴 对王说：“看哪，他在 罗．底巴 ， 亚米利 的儿子 玛吉 家里。”
2SAM|9|5|于是 大卫 王派人去，从 罗．底巴 ， 亚米利 的儿子 玛吉 家里召了他来。
2SAM|9|6|扫罗 的孙子， 约拿单 的儿子 米非波设 来到 大卫 那里，脸伏于地叩拜。 大卫 说：“ 米非波设 ！” 米非波设 说：“看哪，仆人在此。”
2SAM|9|7|大卫 对他说：“你不要惧怕，我必因你父亲 约拿单 的缘故向你施恩，把你祖父 扫罗 的一切田地都归还你，你也可以常与我同席吃饭。”
2SAM|9|8|米非波设 叩拜，说：“你的仆人算什么，不过如死狗一般，竟蒙你这样眷顾！”
2SAM|9|9|王召了 扫罗 的仆人 洗巴 来，对他说：“我已把属 扫罗 和他的一切家产都赐给你主人的儿子了。
2SAM|9|10|你，你的众子和仆人要为你主人的儿子耕种田地，把所收获的拿来供他食用；你主人的儿子 米非波设 却要常与我同席吃饭。” 洗巴 有十五个儿子和二十个仆人。
2SAM|9|11|洗巴 对王说：“凡我主我王吩咐仆人的，仆人都必遵行。”于是 米非波设 与王 同席吃饭，如王的儿子一样。
2SAM|9|12|米非波设 有一个小儿子，名叫 米迦 。凡住在 洗巴 家里的人都作了 米非波设 的仆人。
2SAM|9|13|米非波设 住在 耶路撒冷 ，常与王同席吃饭。他两腿都是瘸的。
2SAM|10|1|此后， 亚扪 人的王死了，他儿子 哈嫩 接续他作王。
2SAM|10|2|大卫 说：“ 哈嫩 的父亲 拿辖 怎样向我施恩，我也要怎样向 哈嫩 施恩。”于是 大卫 派臣仆为他的父亲安慰他。当 大卫 的臣仆到了 亚扪 人的境内，
2SAM|10|3|亚扪 人的领袖对他们的主 哈嫩 说：“ 大卫 派人来安慰你，你看他是要尊敬你父亲吗？ 大卫 派臣仆到你这里，不是为了要窥探侦察，而倾覆这城吗？”
2SAM|10|4|哈嫩 就抓住 大卫 的臣仆，把他们的胡须剃去一半，又割断他们下半截的袍子，露出下体，然后放了他们。
2SAM|10|5|有人告诉 大卫 ，他就派人去迎接他们，因为这些人觉得很羞耻。王说：“可以住在 耶利哥 ，等到胡须长出来再回来。”
2SAM|10|6|亚扪 人看到 大卫 憎恶他们，就派人去雇用 伯．利合 的 亚兰 人和 琐巴 的 亚兰 人，步兵二万，以及 玛迦 王的人一千、 陀伯 人一万二千。
2SAM|10|7|大卫 听见了，就派 约押 和所有勇猛的军队出去。
2SAM|10|8|亚扪 人出来，在城门前摆阵； 琐巴 与 利合 的 亚兰 人、 陀伯 人，以及 玛迦 人另外在郊野摆阵。
2SAM|10|9|约押 看见战阵对着他前后摆列，就把从 以色列 所有精兵中挑选出来的，摆阵迎战 亚兰 人。
2SAM|10|10|他把其余的兵交在他兄弟 亚比筛 手里， 亚比筛 就摆阵迎战 亚扪 人。
2SAM|10|11|约押 对 亚比筛说：“ 亚兰 人若强过我，你就来帮助我； 亚扪 人若强过你，我就去帮助你。
2SAM|10|12|你要刚强，我们要为自己的百姓，为我们上帝的城镇奋勇。愿耶和华照他所看为好的去做！”
2SAM|10|13|于是， 约押 和跟随他的士兵前进攻打 亚兰 人； 亚兰 人在他面前逃跑。
2SAM|10|14|亚扪 人见 亚兰 人逃跑，他们也在 亚比筛 面前逃跑进城。 约押 就离开 亚扪 人，回 耶路撒冷 去了。
2SAM|10|15|亚兰 人见自己被 以色列 打败，就集合起来。
2SAM|10|16|哈大底谢 派人去，把 大河 那边的 亚兰 人调来；他们到了 希兰 ，由 哈大底谢 的将军 朔法 在他们前面率领。
2SAM|10|17|有人告诉 大卫 ，他就聚集 以色列 众人过 约旦河 ，来到 希兰 。 亚兰 人迎着 大卫 摆阵，与他打仗。
2SAM|10|18|亚兰 人在 以色列 人面前逃跑。 大卫 杀了 亚兰 七百辆战车的士兵，四万骑兵 ，又击杀 亚兰 的将军 朔法 ，他就死在那里。
2SAM|10|19|哈大底谢 属下的诸王见自己被 以色列 打败，就与 以色列 讲和，臣服他们。于是 亚兰 人害怕，不再帮助 亚扪 人了。
2SAM|11|1|过了一年，正是诸王出战的时候， 大卫 派 约押 率领臣仆和 以色列 众人出去。他们打败 亚扪 人，围攻 拉巴 。 大卫 仍然留在 耶路撒冷 。
2SAM|11|2|黄昏的时候， 大卫 从床上起来，在王宫的平顶上散步。他从平顶上看见一个妇人沐浴，这妇人容貌非常美丽。
2SAM|11|3|大卫 派人打听那妇人是谁。有人说：“她不是 以连 的女儿， 赫 人 乌利亚 的妻子 拔示巴 吗？”
2SAM|11|4|大卫 派使者去把妇人接来；她来到大卫那里，那时她的月经刚洁净， 大卫 与她同寝。她就回家去了。
2SAM|11|5|那妇人怀了孕，派人去告诉 大卫 说：“我怀孕了。”
2SAM|11|6|大卫 派人告诉 约押 ：“你派 赫 人 乌利亚 到我这里来。” 约押 就派 乌利亚 到 大卫 那里。
2SAM|11|7|乌利亚 来到 大卫那里， 大卫 问 约押 好，也问士兵好，又问战争的情况。
2SAM|11|8|大卫 对 乌利亚 说：“下到你家去，洗洗脚吧！” 乌利亚 出了王宫，随后王送他一份礼物。
2SAM|11|9|乌利亚 却和他主人所有的仆人一同睡在王宫门口，没有下到他家去。
2SAM|11|10|有人告诉 大卫 说：“ 乌利亚 没有下到他的家。” 大卫 就对 乌利亚 说：“你不是从远路上来吗？为什么不下到你家去呢？”
2SAM|11|11|乌利亚 对 大卫 说：“约柜， 以色列 和 犹大 都留在棚里，我主 约押 和我主的仆人都在田野安营，我岂可回家吃喝，与妻子同房呢？我指着王和王的性命起誓：‘我绝不做这事！’”
2SAM|11|12|大卫 对 乌利亚 说：“你今日仍留在这里，明日我打发你去。”于是 乌利亚 那日留在 耶路撒冷 。次日，
2SAM|11|13|大卫 召了 乌利亚 来，叫他在自己面前吃喝，使他喝醉。黄昏的时候， 乌利亚 出去，躺卧在自己的床上；与他主的仆人在一起，并没有下到他的家去。
2SAM|11|14|早晨， 大卫 写信给 约押 ，交 乌利亚 亲手带去。
2SAM|11|15|他在信内写着说：“要派 乌利亚 到战争激烈的前线去，然后你们撤退离开他，使他被击杀而死。”
2SAM|11|16|约押 侦察城的时候，知道敌人哪里有勇士，就派 乌利亚 到那地方。
2SAM|11|17|城里的人出来和 约押 打仗， 大卫 的仆人中有几个士兵被杀， 赫 人 乌利亚 也死了。
2SAM|11|18|于是， 约押 派人去将战争的一切事奏告 大卫 ，
2SAM|11|19|又吩咐使者说：“你把战争的一切事对王说完了，
2SAM|11|20|王若发怒，对你说：‘你们打仗为什么挨近城呢？岂不知敌人会从城墙上射箭吗？
2SAM|11|21|从前击杀 耶路比设 的儿子 亚比米勒 的是谁呢？岂不是一个妇人从城墙上抛下一块上磨石来，打在他身上，他就死在 提备斯 吗？你们为什么挨近城墙呢？’你就说：‘你的仆人 赫 人 乌利亚 也死了。’”
2SAM|11|22|使者就去，照着 约押 所吩咐的一切话来奏告 大卫 。
2SAM|11|23|使者对 大卫 说：“敌人强过我们，出到郊外攻打我们，我们把他们赶回到城门口。
2SAM|11|24|弓箭手从城墙上射你的仆人，射死几个王的仆人，你的仆人 赫 人 乌利亚 也死了。”
2SAM|11|25|大卫 向使者说：“你对 约押 这样说：‘不要为这事难过，因为刀剑可能吞灭这人或那人。你只管竭力攻城，将城倾覆。’你要勉励 约押 。”
2SAM|11|26|乌利亚 的妻听见丈夫 乌利亚 死了，就为丈夫哀哭。
2SAM|11|27|居丧的日子过了， 大卫 派人把她接到宫里，她就作了 大卫 的妻子，给 大卫 生了一个儿子。但 大卫 做的这事，耶和华的眼中看为恶。
2SAM|12|1|耶和华差遣 拿单 到 大卫 那里。 拿单 到了他那里，对他说：“在一座城里有两个人，一个是富翁，一个是穷人。
2SAM|12|2|富翁有极多的牛群羊群；
2SAM|12|3|穷人除了所买来养活的一只小母羊之外，一无所有。小羊在他家里和他儿女一同长大，吃他所吃的，喝他所喝的，睡在他怀中，在他看来如同女儿一样。
2SAM|12|4|有一客人来到这富翁那里，富翁舍不得从自己的牛群羊群中取一只招待来到他那里的旅客，却取了穷人的小母羊，招待来到他那里的人。”
2SAM|12|5|大卫 就非常恼怒那人，对 拿单 说：“我指着永生的耶和华起誓，做这事的人该死！
2SAM|12|6|他必须偿还小母羊四倍，因为他做这事，没有怜悯的心。”
2SAM|12|7|拿单 对 大卫 说：“你就是那人！耶和华－ 以色列 的上帝如此说：‘我膏你作 以色列 的王，我救你脱离 扫罗 的手；
2SAM|12|8|我将你主人的家业赐给你，将你主人的妃嫔交在你怀里，又将 以色列 和 犹大 家赐给你；若还嫌少，我也会如此这般加倍赐给你。
2SAM|12|9|你为什么藐视耶和华的命令，做他眼中看为恶的事呢？你用刀击杀 赫 人 乌利亚 ，又娶了他的妻子为妻，借 亚扪 人的刀杀死他。
2SAM|12|10|现在刀剑必永不离开你的家，因你藐视我，娶了 赫 人 乌利亚 的妻子为妻。’
2SAM|12|11|耶和华如此说：‘看哪，我必从你家中兴起灾祸攻击你；我必在你眼前把你的妃嫔赐给你身边的人，他要在光天化日下与你的妃嫔同寝。
2SAM|12|12|你在暗中做那事，我却要在 以色列 众人面前，在日光之下做这事。’”
2SAM|12|13|大卫 对 拿单 说：“我得罪耶和华了！” 拿单 说：“耶和华已经除去你的罪，你必不至于死。
2SAM|12|14|只是在这事上，你大大藐视耶和华 ，因此，你生的孩子必定要死。”
2SAM|12|15|拿单 就回家去了。 耶和华击打 乌利亚 的妻子为 大卫 生的孩子，他就得了重病。
2SAM|12|16|大卫 为这孩子恳求上帝。 大卫 刻苦禁食，到里面去，躺在地上过夜。
2SAM|12|17|他家中的老臣来到他旁边，要把他从地上扶起来，他却不肯，也不同他们吃饭。
2SAM|12|18|到第七日，孩子死了。 大卫 的臣仆不敢告诉他孩子死了，因他们说：“看哪，孩子还活着的时候，我们劝他，他尚且不听我们的话，我们怎么能告诉他孩子死了，让他做出不好的事呢？”
2SAM|12|19|大卫 见臣仆彼此低声说话，就知道孩子死了。他问臣仆说：“孩子死了吗？”他们说：“死了。”
2SAM|12|20|大卫 就从地上起来，沐浴，抹膏，换了衣服，进耶和华的殿敬拜。然后他回宫，吩咐人为他摆饭，他就吃了。
2SAM|12|21|臣仆对他说：“你所做的是什么事呢？孩子活着的时候，你为他禁食哭泣；孩子死了，你却起来吃饭。”
2SAM|12|22|大卫 说：“孩子还活着，我禁食哭泣，因为我想，或许耶和华怜悯我，会让孩子活下来。
2SAM|12|23|现在孩子死了，我何必禁食呢？我能使他回来吗？我必往他那里去，他却不能回到我这里来。”
2SAM|12|24|大卫 安慰他的妻子 拔示巴 ，与她同房，她就生了儿子，给他起名叫 所罗门 。耶和华喜爱他，
2SAM|12|25|就藉 拿单 先知赐他一个名字，叫 耶底底亚 ；这是为了耶和华的缘故。
2SAM|12|26|约押 攻打 亚扪 人的 拉巴 ，攻占了京城。
2SAM|12|27|约押 派使者到 大卫 那里，说：“我攻打 拉巴 ， 也攻占了水城。
2SAM|12|28|现在你要召集其余的军兵，安营围攻这城，攻占它，免得我攻占这城，人就以我的名叫这城。”
2SAM|12|29|于是 大卫 召集全军，往 拉巴 去攻城，就攻占了它。
2SAM|12|30|他也夺了 米勒公 头上所戴的冠冕，其上的金子重一他连得，又嵌着宝石。这冠冕就戴在 大卫 头上。 大卫 又从城里夺了许多财物，
2SAM|12|31|把城里的百姓拉出来，叫他们用锯，用铁耙，用铁斧做工，派他们在砖窑中服役； 大卫 待 亚扪 各城的居民都是如此。于是， 大卫 和全军都回 耶路撒冷 去了。
2SAM|13|1|后来发生了一件事。 大卫 的儿子 押沙龙 有一个美貌的妹妹，名叫 她玛 。 大卫 的儿子 暗嫩 爱上了她。
2SAM|13|2|暗嫩 为他妹妹 她玛 苦恋成疾，因为 她玛 还是处女， 暗嫩 眼看难以向她行事。
2SAM|13|3|暗嫩 有一个密友，名叫 约拿达 ，是 大卫 长兄 示米亚 的儿子。这 约拿达 为人极其狡猾。
2SAM|13|4|他对 暗嫩 说：“王的儿子啊，你何不告诉我，为何你一天比一天憔悴呢？” 暗嫩 对他说：“我爱上了我兄弟 押沙龙 的妹妹 她玛 。”
2SAM|13|5|约拿达 对他说：“你躺在床上装病，等你父亲来看你，就对他说：‘请让我妹妹 她玛 来，给我东西吃，在我眼前预备食物，使我可以看见，好从她手里接过来吃。’”
2SAM|13|6|于是 暗嫩 躺着装病，王来看他。 暗嫩 对王说：“请让我妹妹 她玛 来，在我眼前为我做两个饼，我好从她手里接过来吃。”
2SAM|13|7|大卫 就派人去宫里，到 她玛 那里，说：“你到你哥哥 暗嫩 的屋里去，为他预备食物。”
2SAM|13|8|她玛 就到她哥哥 暗嫩 的屋里，那时 暗嫩 正躺着。 她玛 拿了面团揉面，在他眼前做饼，把饼烤熟了。
2SAM|13|9|她玛 拿了锅子，在他面前把饼倒出来，他却不肯吃。 暗嫩 说：“每一个人都离开我，出去吧！”众人就都离开他，出去了。
2SAM|13|10|暗嫩 对 她玛 说：“你把食物拿进卧房，我好从你手里接过来吃。” 她玛 就把所做的饼拿进卧房，到她哥哥 暗嫩 那里。
2SAM|13|11|她玛 上前去给他吃，他就拉住 她玛 ，对她说：“我妹妹，你来与我同寝。”
2SAM|13|12|她玛 对他说：“哥哥，不可以！不要玷辱我！ 以色列 中不可以这样做，你不要做这丑事！
2SAM|13|13|我蒙受耻辱，该往那里去呢？至于你，你在 以色列 中也成了一个愚顽人。现在你可以求王，他必不禁止我归你。”
2SAM|13|14|但 暗嫩 不肯听她的话，因他比她更有力，就玷辱她，与她同寝。
2SAM|13|15|随后， 暗嫩 极其恨她，恨她的心比先前爱她的心更甚，就对她说：“你起来，去吧！”
2SAM|13|16|她玛 对 暗嫩 说：“不要这样！你赶我出去的这恶比你刚才向我所做的更严重！”但 暗嫩 不肯听她，
2SAM|13|17|就叫伺候自己的仆人来，说：“把这女子从我这里赶出去！她一出去，你就闩上门。”
2SAM|13|18|那时 她玛 穿着彩衣，因为没有出嫁的公主都穿这样的外袍。 暗嫩 的仆人把她赶出去，她一出去，仆人就闩上门。
2SAM|13|19|她玛 把灰尘撒在头上，撕裂所穿的彩衣，以手抱头，一面走一面哭喊。
2SAM|13|20|她胞兄 押沙龙 对她说：“你哥哥 暗嫩 与你亲近了吗？妹妹，现在暂且不要作声，他是你的哥哥，不要把这事放在心上。” 她玛 就孤孤单单地住在她胞兄 押沙龙 的家里。
2SAM|13|21|大卫 王听见这一切的事，就非常愤怒。
2SAM|13|22|押沙龙 却不和 暗嫩 说好说歹；因为 暗嫩 玷辱他妹妹 她玛 ，所以 押沙龙 恨恶他。
2SAM|13|23|过了二年，有人在靠近 以法莲 的 巴力．夏琐 为 押沙龙 剪羊毛。 押沙龙 请了王所有的儿子来。
2SAM|13|24|押沙龙 来到王那里，说：“看哪，有人正为你的仆人剪羊毛，请王和王的臣仆与你的仆人同去。”
2SAM|13|25|王对 押沙龙 说：“不，我儿，我们不必都去，免得成了你的负担。” 押沙龙 再三请王，王仍是不肯去，只为他祝福。
2SAM|13|26|押沙龙 说：“王若不去，请让我哥哥 暗嫩 与我们同去。”王对他说：“为何要他与你同去呢？”
2SAM|13|27|押沙龙 再三求王，王就派 暗嫩 和王所有的儿子与他同去。
2SAM|13|28|押沙龙 吩咐仆人说：“你们注意， 暗嫩 开怀畅饮的时候，我对你们说击杀 暗嫩 ，你们就杀他。不要惧怕，这不是我吩咐你们的吗？你们要刚强，作勇士！”
2SAM|13|29|押沙龙 的仆人就照 押沙龙 所吩咐的，向 暗嫩 行了。王所有的儿子都起来，各人骑上骡子逃跑了。
2SAM|13|30|他们还在路上，就有风声传到 大卫 那里，说：“ 押沙龙 击杀了王所有的儿子，没有留下一个。”
2SAM|13|31|王就起来，撕裂衣服，躺在地上。王的臣仆全都撕裂衣服，站在旁边。
2SAM|13|32|大卫 的长兄 示米亚 的儿子 约拿达 说：“我主，不要以为他们把所有的年轻人，就是王的儿子都杀了，只有 暗嫩 一个人死了。自从 暗嫩 玷辱了 押沙龙 的妹妹 她玛 那日， 押沙龙 已经决定这事了。
2SAM|13|33|现在，我主我王，不要把这事放在心上，以为王所有的儿子都死了。其实，只有 暗嫩 一人死了。”
2SAM|13|34|押沙龙 逃跑了。守望的年轻人举目观看，看哪，有许多人从 何罗念 山坡的路上来。
2SAM|13|35|约拿达 对王说：“看哪，王的儿子都来了，正如你仆人所说的，事情就这样发生了。”
2SAM|13|36|话刚说完，看哪，王的儿子都到了，放声大哭。王和他的众臣仆也都号啕痛哭。
2SAM|13|37|押沙龙 逃到 亚米忽 的儿子 基述 王 达买 那里去了。 大卫 天天为他儿子悲哀。
2SAM|13|38|押沙龙 逃到 基述 去了，在那里住了三年。
2SAM|13|39|王想要出去对付 押沙龙 的心化解了 ，因为王对 暗嫩 之死这事已经得了安慰。
2SAM|14|1|洗鲁雅 的儿子 约押 知道王心里想念 押沙龙 。
2SAM|14|2|他派人往 提哥亚 去，从那里叫了一个有智慧的妇人来，对她说：“请你装作居丧的人，穿上丧服，不用膏抹身，装作为死者悲哀多日的妇人。
2SAM|14|3|你到王那里，对王如此如此说。”于是 约押 把当说的话放在她口中。
2SAM|14|4|提哥亚 妇人到王面前 ，脸伏于地叩拜，说：“王啊，求你拯救！”
2SAM|14|5|王对她说：“你有什么事呢？”她说：“我实在是个寡妇，我丈夫死了。
2SAM|14|6|婢女有两个儿子，二人在田间打架，没有人从中劝解，一个击杀另一个，把他打死了。
2SAM|14|7|看哪，全家族都起来攻击婢女，说：‘把那打死兄弟的交出来，我们好处死他，为他所打死的兄弟偿命，灭绝那承受家业的。’这样，他们要把我剩下的炭火灭尽，不给我丈夫留名或留后在地面上。”
2SAM|14|8|王对妇人说：“你回家去吧！我必为你下个命令。”
2SAM|14|9|提哥亚 妇人又对王说：“我主我王，愿这罪孽归我和我的父家，与王和王的位无关。”
2SAM|14|10|王说：“有人说话难为你，你就带他到我这里来，他必不再搅扰你。”
2SAM|14|11|妇人说：“愿王对耶和华－你的上帝发誓，不许报血仇的人施行毁灭，免得他们灭绝我的儿子。”王说：“我指着永生的耶和华起誓：你的儿子连一根头发也不致落在地上。”
2SAM|14|12|妇人说：“求我主我王容许婢女再说一句话。”王说：“你说吧！”
2SAM|14|13|妇人说：“王为何起意做这事，要害上帝的百姓呢？王不使那逃亡的人回来，王说这话就证实自己错了！
2SAM|14|14|我们都必死，如同水泼在地上，不能收回。上帝不会让人不死，但仍设法 使逃亡的人不致成为赶出、回不来的人。
2SAM|14|15|现在我来将这话告诉我主我王，是因百姓使我惧怕。婢女想：‘不如告诉王，或者王会成就使女所求的。
2SAM|14|16|人要把我和我儿子从上帝的地业上一同除灭，王必应允救使女脱离他的手。’
2SAM|14|17|婢女想：‘我主我王的话必安慰我’；因为我主我王能辨别是非，如同上帝的使者一样。惟愿耶和华－你的上帝与你同在！”
2SAM|14|18|王回答妇人说：“我问你一句话，你一点也不可瞒我。”妇人说：“我主我王，请说。”
2SAM|14|19|王说：“这一切莫非是 约押 的手指使你的吗？”妇人回答说：“我敢在我主我王面前起誓：我主我王所说的一切不偏左右，这是王的仆人 约押 吩咐我的，这一切话是他放在婢女口中的。
2SAM|14|20|王的仆人 约押 做这事，为要扭转局面。我主的智慧却如上帝使者的智慧，能知地上一切的事。”
2SAM|14|21|王对 约押 说：“看哪，我应允这事。你去，把那年轻人 押沙龙 带回来。”
2SAM|14|22|约押 脸伏于地叩拜，为王祝福，说：“王既应允仆人这件事，仆人今日知道在我主我王眼前蒙恩宠了。”
2SAM|14|23|于是 约押 起身往 基述 去，把 押沙龙 带回 耶路撒冷 。
2SAM|14|24|王说：“让他回自己的家去，不要来见我的面。” 押沙龙 就回自己的家去，没有见王的面。
2SAM|14|25|全 以色列 中，无人像 押沙龙 那样俊美，得人称赞，从脚底到头顶毫无瑕疵。
2SAM|14|26|他的头发很重，每到年底剪发一次，所剪下来的，按王的秤称一称，重二百舍客勒。
2SAM|14|27|押沙龙 生了三个儿子，一个女儿。女儿名叫 她玛 ，是个容貌美丽的女子。
2SAM|14|28|押沙龙 住在 耶路撒冷 ，足足有二年没有见王的面。
2SAM|14|29|押沙龙 派人去叫 约押 来，要托他到王那里去， 约押 却不肯来。 押沙龙 第二次派人去叫他，他仍不肯来。
2SAM|14|30|于是 押沙龙 对仆人说：“你们看， 约押 有一块田靠近我的田，其中有大麦，你们去放火把它烧了。” 押沙龙 的仆人就去放火烧了那田。
2SAM|14|31|于是 约押 起来，到了 押沙龙 家里，对他说：“你的仆人为何放火烧我的田呢？”
2SAM|14|32|押沙龙 对 约押 说：“看哪，我派人去请你来，好托你到王那里去，说：‘我为何从 基述 回来呢？我仍在那里比较好。’现在让我去见王的面；我若有罪孽，就任凭王杀了我吧。”
2SAM|14|33|于是 约押 到王那里，奏告王，王就叫 押沙龙 来。 押沙龙 到王那里，在王面前脸伏于地，王就亲吻 押沙龙 。
2SAM|15|1|此后， 押沙龙 为自己预备车马，又派五十人在他前头奔跑。
2SAM|15|2|押沙龙 常常早晨起来，站在城门的路旁，任何人有争讼要去求王判决， 押沙龙 就叫他过来，说：“你是哪一城的人？”他说：“仆人是 以色列 某支派的人。”
2SAM|15|3|押沙龙 就对他说：“看，你的案件合情合理，无奈王没有委派人听你申诉。”
2SAM|15|4|押沙龙 又说：“恨不得我作这地的审判官！ 凡有争讼的人可以到我这里来，我必秉公判断。”
2SAM|15|5|若有人近前来要拜 押沙龙 ， 押沙龙 就伸手拉住他，亲吻他。
2SAM|15|6|以色列 中，凡到王那里求判决的， 押沙龙 都这么做。这样， 押沙龙 暗中赢得了 以色列 人的心。
2SAM|15|7|过了四年 ， 押沙龙 对王说：“求你准我往 希伯仑 去，还我向耶和华所许的愿。
2SAM|15|8|因为仆人住在 亚兰 的 基述 时，曾许愿说：‘耶和华若使我再回 耶路撒冷 ，我必事奉他 。’”
2SAM|15|9|王对他说：“你平安地去吧！” 押沙龙 就动身，往 希伯仑 去了。
2SAM|15|10|押沙龙 派密使走遍 以色列 各支派，说：“你们一听见角声就说：‘ 押沙龙 在 希伯仑 作王了！’”
2SAM|15|11|押沙龙 在 耶路撒冷 请了二百人与他同去，都是诚心诚意去的，一点也不知道实情。
2SAM|15|12|押沙龙 献祭的时候，派人去把 大卫 的谋士， 基罗 人 亚希多弗 从他本城 基罗 请来 。于是叛乱越发强大，因为随从 押沙龙 的百姓日渐增多。
2SAM|15|13|报信的人来到 大卫 那里，说：“ 以色列 人的心都归向 押沙龙 了！”
2SAM|15|14|大卫 就对 耶路撒冷 所有跟随他的臣仆说：“起来，我们逃吧！否则，我们来不及逃避 押沙龙 。要快点离开，免得他很快追上我们，加害于我们，用刀击杀城里的人。”
2SAM|15|15|王的臣仆对王说：“我主我王所决定的一切，看哪，仆人都愿遵行。”
2SAM|15|16|于是王出去了，他的全家都跟随他，但留下十个妃嫔看守宫殿。
2SAM|15|17|王出去，众百姓都跟随他；到了最后一座屋子 ，他们就停下来。
2SAM|15|18|王的众臣仆都在他旁边过去。 基利提 人、 比利提 人，和从 迦特 跟随王来的六百个 迦特 人，也都在王面前过去。
2SAM|15|19|王对 迦特 人 以太 说：“你是外邦人，从你本地逃来的，为什么与我们同去呢？你回去留在新王那里吧！
2SAM|15|20|你昨天才到，我今日怎好叫你与我们一同流亡，而我却要到处飘流呢？回去吧，你带你的弟兄回去吧！愿主用慈爱信实待你 。”
2SAM|15|21|以太 回答王说：“我指着永生的耶和华起誓，又敢在王面前起誓：无论生死，王在哪里，你的仆人也必在哪里。”
2SAM|15|22|大卫 对 以太 说：“去，过去吧！”于是 迦特 人 以太 带着所有跟随他的人和孩子过去了。
2SAM|15|23|众百姓过去时，当地的人全都放声大哭。王过了 汲沦溪 ，众百姓就往旷野的路上去了。
2SAM|15|24|看哪， 撒督 和所有抬上帝约柜的 利未 人也一同来了。他们将上帝的约柜放下， 亚比亚他 上来 ，直到众百姓从城里出来走过去为止。
2SAM|15|25|王对 撒督 说：“你将上帝的约柜请回城去。我若在耶和华眼前蒙恩，他必使我回来，再见到约柜和他的居所。
2SAM|15|26|倘若他说：‘我不喜爱你’；我在这里，就照他眼中看为好的待我！”
2SAM|15|27|王对 撒督 祭司说：“你不是先见吗？你可以平安地回城，你儿子 亚希玛斯 和 亚比亚他 的儿子 约拿单 ，你们二人的儿子可以与你们同去。
2SAM|15|28|看，我在旷野的渡口那里等，直到你们来报信给我。”
2SAM|15|29|于是 撒督 和 亚比亚他 将上帝的约柜请回 耶路撒冷 ，他们就留在那里。
2SAM|15|30|大卫 蒙头赤脚走上 橄榄山 的斜坡，一面上一面哭。所有跟随他的百姓也都各自蒙头哭着上去；
2SAM|15|31|有人告诉 大卫 说 ：“ 亚希多弗 也在叛党之中，随从 押沙龙 。” 大卫 说：“耶和华啊，求你使 亚希多弗 的计谋变为愚拙！”
2SAM|15|32|大卫 到了山顶，敬拜上帝的地方，看哪， 亚基 人 户筛 衣服撕裂，头蒙灰尘来迎见他。
2SAM|15|33|大卫 对他说：“你若与我一同过去，必拖累我；
2SAM|15|34|你若回城去，对 押沙龙 说：‘王啊，我愿作你的仆人。我向来作你父亲的仆人，现在我也愿意作你的仆人。’你就可以为我破坏 亚希多弗 的计谋。
2SAM|15|35|撒督 和 亚比亚他 二位祭司岂不都在你那里吗？你在王宫里听见什么，就要告诉 撒督 和 亚比亚他 二位祭司。
2SAM|15|36|看哪， 撒督 的儿子 亚希玛斯 ， 亚比亚他 的儿子 约拿单 ，也跟二位祭司在那里。凡你们所听见的事，可以托这二人来向我报告。”
2SAM|15|37|于是， 大卫 的朋友 户筛 进了城， 押沙龙 也进了 耶路撒冷 。
2SAM|16|1|大卫 刚过山顶，看哪， 米非波设 的仆人 洗巴 拉着装好鞍子的两匹驴，驴上驮着二百个面饼，一百个葡萄饼，一百个夏天的果饼，一皮袋酒来迎接他。
2SAM|16|2|王对 洗巴 说：“你的这些东西是什么意思呢？” 洗巴 说：“驴是给王的家眷骑的，面饼和夏天的果饼是给年轻人吃的，酒是给在旷野疲乏的人喝的。”
2SAM|16|3|王说：“你主人的儿子在哪里呢？” 洗巴 对王说：“看哪，他留在 耶路撒冷 ，因他说：‘ 以色列 家今日必将我父的国归还我。’”
2SAM|16|4|王对 洗巴 说：“看哪，凡属 米非波设 的都是你的了。” 洗巴 说：“我叩拜我主我王，愿我在你眼前蒙恩宠。”
2SAM|16|5|大卫 王到了 巴户琳 ，看哪，有一个人从那里出来，是 扫罗 家族中 基拉 的儿子，名叫 示每 。他一面走一面咒骂，
2SAM|16|6|又向 大卫 王和王的众臣仆扔石头；众百姓和勇士都在王的左右。
2SAM|16|7|示每 这样咒骂说：“你这好流人血的，你这无赖，滚吧！滚吧！
2SAM|16|8|你流了 扫罗 全家的血，接续他作王，耶和华把这罪归在你身上。耶和华将这国交在你儿子 押沙龙 的手中。看哪，你咎由自取，因为你是好流人血的人。”
2SAM|16|9|洗鲁雅 的儿子 亚比筛 对王说：“这死狗为何咒骂我主我王呢？让我过去，割下他的头来。”
2SAM|16|10|王说：“ 洗鲁雅 的儿子，我与你们有何相干呢？他这样咒骂是因耶和华吩咐他：‘你要咒骂 大卫 。’如此，谁敢说：‘你为什么这样做呢？’”
2SAM|16|11|大卫 又对 亚比筛 和众臣仆说：“看哪，我亲生的儿子尚且寻索我的性命，何况现在这 便雅悯 人呢？由他咒骂吧！因为这是耶和华吩咐他的。
2SAM|16|12|或者耶和华见我遭难 ，因我今日被这人咒骂而向我施恩。”
2SAM|16|13|于是 大卫 和他的人在路上走。 示每 走在 大卫 对面的山坡，一面走一面咒骂，又向他扔石头，扬起尘土。
2SAM|16|14|王和跟随他的众百姓来了，非常疲乏，就在那里歇息。
2SAM|16|15|押沙龙 和 以色列 众百姓来到 耶路撒冷 ， 亚希多弗 也与他同来。
2SAM|16|16|大卫 的朋友 亚基 人 户筛 来到 押沙龙 那里，对他说：“愿王万岁！愿王万岁！”
2SAM|16|17|押沙龙 对 户筛 说：“你这样做是忠诚对待你的朋友吗？为什么不与你的朋友同去呢？”
2SAM|16|18|户筛 对 押沙龙 说：“不，谁是耶和华和这百姓，以及 以色列 众人所拣选的，我必归顺他，留在他那里。
2SAM|16|19|再者，我当服事谁呢？岂不是前王的儿子吗？我怎样服事你父亲，也必照样服事你。”
2SAM|16|20|押沙龙 对 亚希多弗 说：“你们出个主意，我们该怎么做？”
2SAM|16|21|亚希多弗 对 押沙龙 说：“你父亲所留下看守宫殿的妃嫔，你可以与她们亲近。 以色列 众人听见你敢惹你父亲憎恶你，凡归顺你人的手就更坚强了。”
2SAM|16|22|于是他们为 押沙龙 在屋顶上支搭帐棚， 押沙龙 就在 以色列 众人眼前，与他父亲的妃嫔亲近。
2SAM|16|23|那时 亚希多弗 所出的主意好像人从上帝求问得来的话一样；他给 大卫 ，给 押沙龙 所出的一切主意，都是这样。
2SAM|17|1|亚希多弗 对 押沙龙 说：“请让我挑选一万二千人，今夜起身追赶 大卫 。
2SAM|17|2|我必趁他疲乏手软的时候追上他，使他惊惶。跟随他的众百姓必都逃跑，我就只杀王一个人。
2SAM|17|3|我必使众百姓都归顺你，正如众人归顺你所追杀的人一样 ，众百姓就都平安无事了。”
2SAM|17|4|这话在 押沙龙 和 以色列 众长老的眼中都看为好。
2SAM|17|5|押沙龙 说：“把 亚基 人 户筛 也召来，我们也要听他怎么说。”
2SAM|17|6|户筛 到了 押沙龙 那里， 押沙龙 向他说：“ 亚希多弗 说了这样的话，我们要照他的话做吗？若不可，你就说吧！”
2SAM|17|7|户筛 对 押沙龙 说：“ 亚希多弗 这次所出的主意不好。”
2SAM|17|8|户筛 又说：“你知道，你父亲和他的人都是勇士，他们心里恼怒，如同田野中失去小熊的母熊一样；而且你父亲是个战士，必不和百姓一同住宿。
2SAM|17|9|看哪，他现今或藏在一个坑中或在别处，若我们 有人首先被杀，听见的必说：‘跟随 押沙龙 的百姓被杀了。’
2SAM|17|10|虽有勇士胆大如狮子，他的心也必定融化，因为全 以色列 都知道你父亲是英雄，跟随他的人都是勇士。
2SAM|17|11|依我之计，要把如同海边的沙那样多的 以色列 众人，从 但 直到 别是巴 ，聚集到你这里来，由你亲自率领他们出战。
2SAM|17|12|我们到他那里，在任何地方遇见他，就突然临到他，如同露水滴在泥土上。这样，他和所有跟随他的人，一个也不留。
2SAM|17|13|他若撤退到一座城， 以色列 众人必带绳子去那城，把城拉到河里，甚至连一块小石子也找不到。”
2SAM|17|14|押沙龙 和 以色列 众人都说：“ 亚基 人 户筛 的计谋比 亚希多弗 的更好！”这是因为耶和华定意破坏 亚希多弗 的良谋，为的是耶和华要降祸给 押沙龙 。
2SAM|17|15|户筛 对 撒督 和 亚比亚他 二位祭司说：“ 亚希多弗 为 押沙龙 和 以色列 的长老出的主意是如此如此，我出的主意是如此如此。
2SAM|17|16|现在你们要急速派人去告诉 大卫 说：‘今夜不可在旷野的渡口住宿，务要过河，免得王和所有跟随他的百姓都被吞灭。’”
2SAM|17|17|约拿单 和 亚希玛斯 在 隐．罗结 等候，不敢进城，恐怕被人看见。有一个婢女出来，把这话告诉他们，他们就去报信给 大卫 王。
2SAM|17|18|然而有一个僮仆看见他们，就去告诉 押沙龙 。他们二人急忙离开，跑到 巴户琳 一个人的家里。那人院中有一口井，他们就下到那里。
2SAM|17|19|那家的妇人用盖盖上井口，又在上头铺上碎麦，事情就没有泄漏。
2SAM|17|20|押沙龙 的仆人来到妇人的家，说：“ 亚希玛斯 和 约拿单 在哪里？”妇人对他们说：“他们过了河了。”仆人搜寻，却找不着，就回 耶路撒冷 去了。
2SAM|17|21|他们走后，二人从井里上来，去告诉 大卫 王。他们对 大卫 说：“ 亚希多弗 出这样的主意要害你，你们起来，快快过河。”
2SAM|17|22|于是 大卫 和所有跟随他的百姓都起来，过 约旦河 。到了天亮，无一人不过 约旦河 的。
2SAM|17|23|亚希多弗 见他的计谋不被接纳，就备上驴，动身归回本城，到了自己的家。他留下遗嘱给他的家，就上吊死了，葬在他父亲的坟墓里。
2SAM|17|24|大卫 到了 玛哈念 ， 押沙龙 和跟随他的 以色列 众人也都过了 约旦河 。
2SAM|17|25|押沙龙 立 亚玛撒 作元帅，取代 约押 。 亚玛撒 是 以实玛利 人 以特拉 的儿子。 以特拉 曾与 拿辖 的女儿 亚比该 亲近；这 亚比该 与 约押 的母亲 洗鲁雅 是姊妹。
2SAM|17|26|押沙龙 和 以色列 人安营在 基列 地。
2SAM|17|27|大卫 到了 玛哈念 ， 亚扪 族的 拉巴 人 拿辖 的儿子 朔比 ， 罗．底巴 人 亚米利 的儿子 玛吉 ，来自 罗基琳 的 基列 人 巴西莱 ，
2SAM|17|28|带着被褥、盆、瓦器，还有小麦、大麦、麦面、烤熟的谷穗、豆子、红豆、炒豆、
2SAM|17|29|蜂蜜、奶油、绵羊、奶饼，供给 大卫 和跟随他的人吃，因为他们想：“百姓在旷野中，必定又饥渴又疲乏。”
2SAM|18|1|大卫 数点跟随他的百姓，立千夫长、百夫长率领他们。
2SAM|18|2|大卫 把军兵分为三队 ：三分之一在 约押 手下，三分之一在 洗鲁雅 的儿子 约押 弟弟 亚比筛 手下，三分之一在 迦特 人 以太 手下。王对军兵说：“我必与你们一同出战。”
2SAM|18|3|军兵却说：“你不可出战。若是我们逃跑，敌人不会把心放在我们身上；我们阵亡一半，敌人也不会把心放在我们身上。但现在你一人抵过我们万人，所以你最好留在城里支援我们。”
2SAM|18|4|王对他们说：“你们看怎样好，我就怎样做。”于是王站在城门旁，所有的军兵成百成千地挨次出战去了。
2SAM|18|5|王嘱咐 约押 、 亚比筛 、 以太 说：“你们要为我的缘故宽待那年轻人 押沙龙 。”王为 押沙龙 的事嘱咐众将领的话，所有的军兵都听见了。
2SAM|18|6|军兵出到田野迎战 以色列 ，在 以法莲 的树林里交战。
2SAM|18|7|在那里， 以色列 百姓败在 大卫 的臣仆面前。那日在那里阵亡的很多，共有二万人。
2SAM|18|8|战争蔓延到整个地面，那日被树林吞噬的军兵比被刀剑吞噬的更多。
2SAM|18|9|押沙龙 刚好遇见了 大卫 的臣仆。 押沙龙 骑着骡子，从大橡树密枝底下经过，他的头被橡树夹住，悬挂在空中 ，所骑的骡子就离他去了。
2SAM|18|10|有个人看见，就告诉 约押 说：“看哪，我看见 押沙龙 挂在橡树上了。”
2SAM|18|11|约押 对报信的人说：“看哪，你既看见了，为什么不当场把他击杀在地呢？我必赏你十个银子和一条带子。”
2SAM|18|12|那人对 约押 说：“即使我手里得了一千银子，也不敢伸手害王的儿子，因为我们听见王嘱咐你、 亚比筛 、 以太 说：‘你们要谨慎，不可害那年轻人 押沙龙 。’
2SAM|18|13|我若冒着生命危险做这傻事 ，无论何事都瞒不过王，你自己也必远远站在一旁。”
2SAM|18|14|约押 说：“我不能在你面前这样耗下去！” 约押 手拿三枝短枪，趁 押沙龙 在橡树上 还活着，就刺透他的心。
2SAM|18|15|给 约押 拿兵器的十个青年围着 押沙龙 ，击杀他，将他杀死。
2SAM|18|16|约押 吹角，军兵就回来，不去追赶 以色列 人，因为 约押 制止了军兵。
2SAM|18|17|他们拿下 押沙龙 ，把他丢在树林中一个大坑里，上头堆起一大堆石头。 以色列 众人都逃跑，各回自己的帐棚去了。
2SAM|18|18|押沙龙 活着的时候，曾在 王谷 立了一根柱子，因他说：“我没有儿子为我留名。”他就以自己的名字称那柱子为 押沙龙碑 ，直到今日。
2SAM|18|19|撒督 的儿子 亚希玛斯 说：“让我跑去报信给王，耶和华已经为王伸冤，使他脱离仇敌的手了。”
2SAM|18|20|约押 对他说：“你今日不可作报信的人，改日再去报信；因为今日王的儿子死了，所以你不可去报信。”
2SAM|18|21|约押 对 古实 人说：“你去把你所看见的告诉王。” 古实 人向 约押 叩拜后，就跑去了。
2SAM|18|22|撒督 的儿子 亚希玛斯 又对 约押 说：“无论怎样，让我随着 古实 人跑去吧！” 约押 说：“我儿，你报这信息，既不得赏赐，何必要跑去呢？”
2SAM|18|23|他说：“无论怎样，我要跑去。” 约押 对他说：“你跑去吧！” 亚希玛斯 就从平原的路往前跑，越过了 古实 人。
2SAM|18|24|大卫 正坐在内外城门之间。守望的人上到城墙，在城门的顶上举目观看，看哪，有一个人独自跑来。
2SAM|18|25|守望的人就大声告诉王。王说：“他若独自来，必是报口信的。”那人跑得越来越近了。
2SAM|18|26|守望的人又见一人跑来，就对守城门的人喊说：“看哪，又有一人独自跑来。”王说：“这也是报信的。”
2SAM|18|27|守望的人说：“我看前面那人的跑法，好像 撒督 的儿子 亚希玛斯 的跑法。”王说：“他是个好人，是来报好消息的。”
2SAM|18|28|亚希玛斯 向王呼叫说：“平安了！”他就脸伏于地向王叩拜，说：“耶和华－你的上帝是应当称颂的，他已把些那举手攻击我主我王的人交出来了。”
2SAM|18|29|王说：“年轻人 押沙龙 平安吗？” 亚希玛斯 说：“ 约押 派王的仆人，就是你的仆人时，我看见一阵大骚动，却不知道是什么事。”
2SAM|18|30|王说：“你退去，站在这里。”他就退去，站着。
2SAM|18|31|看哪， 古实 人也来到，说：“有信息报给我主我王！耶和华今日为你伸冤，使你脱离一切起来攻击你之人的手。”
2SAM|18|32|王对 古实 人说：“年轻人 押沙龙 平安吗？” 古实 人说：“愿我主我王的仇敌，和一切起来恶意要害你的人，都像那年轻人一样。”
2SAM|18|33|王战抖，就上城门的楼房去痛哭，一面走一面说：“我儿 押沙龙 啊！我儿，我儿 押沙龙 啊！我恨不得替你死， 押沙龙 啊，我儿！我儿！”
2SAM|19|1|有人告诉 约押 ：“看哪，王为 押沙龙 悲哀哭泣。”
2SAM|19|2|那日众军兵听说王为他儿子悲伤，他们得胜的日子变成悲哀了。
2SAM|19|3|那日军兵暗暗地进城，如同战场上逃跑、羞愧的士兵一般。
2SAM|19|4|王蒙着脸，大声哭号说：“我儿 押沙龙 啊！ 押沙龙 ，我儿，我儿啊！”
2SAM|19|5|约押 进了宫到王那里，说：“你今日使你众臣仆的脸面羞愧了！他们今日救了你的性命和你儿女妻妾的性命，
2SAM|19|6|你却爱那些恨你的人，恨那些爱你的人。今日你摆明了不以将帅、臣仆为念。我今日看得出，若 押沙龙 活着，我们今日全都死了，你就高兴了。
2SAM|19|7|现在你要起来，出去安慰你臣仆的心。我指着耶和华起誓：你若不出去，今夜必没有一人跟你在一起了。这祸患比你从幼年到如今所遭受的更严重！”
2SAM|19|8|于是王起来，坐在城门口。有人告诉众军兵说：“看哪，王坐在城门口。”众军兵就都到王的面前。 那时， 以色列 人已经逃跑，各回自己的帐棚去了。
2SAM|19|9|以色列 众支派的百姓都议论纷纷，说：“王曾救我们脱离仇敌的手，又救我们脱离 非利士 人的手，现在他为了 押沙龙 逃离这地了。
2SAM|19|10|我们所膏治理我们的 押沙龙 已经阵亡。现在你们为什么沉默，不请王回来呢？”
2SAM|19|11|大卫 王派人到 撒督 和 亚比亚他 二位祭司那里，说：“你们当向 犹大 长老说：‘ 以色列 众人已经有话到了王那里 ，你们为什么最后才请王回宫呢？
2SAM|19|12|你们是我的弟兄，是我的骨肉，为什么最后才请王回来呢？’
2SAM|19|13|你们要对 亚玛撒 说：‘你不是我的骨肉吗？我若不立你在我面前取代 约押 永久作元帅，愿上帝重重惩罚我！’”
2SAM|19|14|这样，他挽回了 犹大 众人的心，如同一人。他们就派人到王那里，说：“请王和王的众臣仆回来。”
2SAM|19|15|王回来了，到 约旦河 。 犹大 人来到 吉甲 ，去迎接王，请王过 约旦河 。
2SAM|19|16|来自 巴户琳 的 便雅悯 人 基拉 的儿子 示每 急忙与 犹大 人一同下去迎接 大卫 王。
2SAM|19|17|跟从 示每 的有一千个 便雅悯 人，还有 扫罗 家的仆人 洗巴 和他十五个儿子、二十个随从仆人，他们都赶紧过 约旦河 到王的面前。
2SAM|19|18|渡船就渡王的家眷过河 ，照王看为好的去做。 王过 约旦河 的时候， 基拉 的儿子 示每 俯伏在王面前，
2SAM|19|19|对王说：“我主我王离开 耶路撒冷 的那日，仆人行了悖逆的事，现在求我主不要因此加罪于仆人，不要记得，也不要放在心上。
2SAM|19|20|仆人明知自己有罪，看哪， 约瑟 全家之中，今日我首先下来迎接我主我王。”
2SAM|19|21|洗鲁雅 的儿子 亚比筛 回答说：“ 示每 既然咒骂耶和华的受膏者，不应当为这缘故处死他吗？”
2SAM|19|22|大卫 说：“ 洗鲁雅 的儿子，我与你们有何相干，你们今日要跟我作对吗？今日在 以色列 中岂可把任何人处死呢？我岂不知今日我是 以色列 的王吗？”
2SAM|19|23|于是王对 示每 说：“你必不死。”王就向他起誓。
2SAM|19|24|扫罗 的孙子 米非波设 也下去迎接王。他自从王离开的那一日，直到王平安回 耶路撒冷 的日子，没有修脚，没有剃胡须，也没有洗衣服。
2SAM|19|25|他来迎接王的时候 ，王对他说：“ 米非波设 ，你为什么没有与我同去呢？”
2SAM|19|26|他说：“我主我王啊，我的仆人欺骗了我。那日仆人想要备驴骑上，与王同去，因为仆人是瘸腿的。
2SAM|19|27|他却在我主我王面前毁谤仆人。然而我主我王如同上帝的使者一样，你看怎样好，就怎样做吧！
2SAM|19|28|因为我祖全家的人，在我主我王面前不过是该死的人，王却使仆人列在王的席上吃饭的人当中，我现在还有什么权利能向王请求呢？”
2SAM|19|29|王对他说：“你何必再提你的事呢？我说，你与 洗巴 要平分土地。”
2SAM|19|30|米非波设 对王说：“我主我王既然平安地回宫，甚至让 洗巴 全都拿去也没关系。”
2SAM|19|31|基列 人 巴西莱 从 罗基琳 下来，要护送王过 约旦河 ，就跟王一同过 约旦河 。
2SAM|19|32|巴西莱 年纪老迈，已经八十岁了。王住在 玛哈念 的时候，他拿食物来供给王，因他是个大富翁。
2SAM|19|33|王对 巴西莱 说：“你与我一同渡过去，我要在 耶路撒冷 我的身边奉养你。”
2SAM|19|34|巴西莱 对王说：“我还能活多少年日，可以与王一同上 耶路撒冷 呢？
2SAM|19|35|今日我已八十岁了，还能辨别美丑吗？仆人还能尝出饮食的滋味吗？还能听男女歌唱的声音吗？仆人何必拖累我主我王呢？
2SAM|19|36|仆人护送王过 约旦河 只是一件小事，王何必用这样的赏赐来报答我呢？
2SAM|19|37|请让我回去，死在我本城，葬在我父母的墓旁。看哪，这里有 金罕 作王的仆人，让他同我主我王过去，你看怎样好，就怎样对待他吧。”
2SAM|19|38|王说：“ 金罕 可以与我一同过去，我必照你看为好的待他。你要我做的，我都会为你做。”
2SAM|19|39|于是众百姓过了 约旦河 ，王也过去了。王亲吻 巴西莱 ，为他祝福， 巴西莱 就回自己的地方去了。
2SAM|19|40|王渡过去 ，到了 吉甲 ， 金罕 也跟他过去。 犹大 众百姓和 以色列 百姓的一半也都送王过去。
2SAM|19|41|看哪， 以色列 众人来到王那里，对王说：“我们的弟兄 犹大 人为什么暗暗地送王和王的家眷，以及所有跟随王的人，过 约旦河 呢？”
2SAM|19|42|犹大 众人回答 以色列 人说：“因为王与我们是亲属，你们为何因这事发怒呢？我们靠王吃了什么呢？王真正给了我们什么赏赐呢？”
2SAM|19|43|以色列 人回答 犹大 人说：“我们与王有十倍的关系，就是在 大卫 身上，我们也比你们更有权利 。你们为何藐视我们呢？我们不是最先提议请王回来的吗？”但 犹大 人的话比 以色列 人的话更强硬。
2SAM|20|1|在那里恰巧有一个无赖，名叫 示巴 ，是 便雅悯 人 比基利 的儿子。他吹角，说： “我们与 大卫 无份， 与 耶西 的儿子无关。 以色列 啊，各回自己的帐棚去吧！”
2SAM|20|2|于是 以色列 众人都离弃 大卫 去跟随 比基利 的儿子 示巴 ，但 犹大 人从 约旦河 直到 耶路撒冷 ，都紧紧跟随他们的王。
2SAM|20|3|大卫 王来到 耶路撒冷 ，进了宫，就把从前留下看守宫殿的十个妃嫔软禁在冷宫，养活她们，却不与她们亲近。她们被关起来，活着如同寡妇，直到死的日子。
2SAM|20|4|王对 亚玛撒 说：“你要在三日之内召集 犹大 人到我这里来，你自己也要留在这里。”
2SAM|20|5|亚玛撒 就去召集 犹大 人，不过他却耽延，过了王所定的期限。
2SAM|20|6|大卫 对 亚比筛 说：“现在 比基利 的儿子 示巴 对我们的危害恐怕比 押沙龙 更大。你要带领你主的一些仆人追赶他，免得他得了坚固的城镇，在我们眼前逃脱 。”
2SAM|20|7|约押 的人和 基利提 人、 比利提 人，以及所有的勇士都跟着 亚比筛 ，从 耶路撒冷 出去追赶 比基利 的儿子 示巴 。
2SAM|20|8|他们到了 基遍 的大石头那里， 亚玛撒 来迎接他们。那时 约押 穿着战衣，腰束佩刀的带子，刀在鞘内。 约押 前行时，刀从鞘内掉出来。
2SAM|20|9|约押 对 亚玛撒 说：“我的弟兄，你平安吗？”他就用右手抓住 亚玛撒 的胡子，要亲吻他。
2SAM|20|10|亚玛撒 没有防备 约押 手里拿着的刀； 约押 用刀刺入他的肚腹，他的肠子流在地上， 约押 没有再刺，他就死了。 约押 和他弟弟 亚比筛 往前追赶 比基利 的儿子 示巴 。
2SAM|20|11|有 约押 的一个仆人站在 亚玛撒 尸体的旁边，说：“谁喜爱 约押 ，谁归顺 大卫 ，就当跟随 约押 。”
2SAM|20|12|亚玛撒 浑身是血，躺在路中间。那人见众百姓都站住，就把 亚玛撒 的尸体从路上移到田间，把衣服盖在他身上，因为他看见众人经过时都站住。
2SAM|20|13|尸体从路上移走之后，众人就都跟随 约押 去追赶 比基利 的儿子 示巴 。
2SAM|20|14|示巴 走遍 以色列 各支派，直到 伯．玛迦 的 亚比拉 ；所有精选的人 都聚集跟随他。
2SAM|20|15|跟随 约押 的众百姓到了 伯．玛迦 的 亚比拉 ，围困 示巴 ，对着城建土堆，与城郭相对。他们猛撞城墙，要使城倒塌。
2SAM|20|16|一个有智慧的妇人从城上呼叫：“听啊，听啊，请你们告诉 约押 ：‘近前来到这里，我好与你说话。’”
2SAM|20|17|约押 就近前到她那里，妇人对他说：“你是 约押 吗？”他说：“我是。”妇人对他说：“请你听使女的话。” 约押 说：“我正在听。”
2SAM|20|18|妇人说：“古时有话说，当在 亚比拉 求问，事情就可以解决。
2SAM|20|19|我在 以色列 中是和平、忠诚的。你现在想要毁坏这城， 以色列 的根源 ，为何你要吞灭耶和华的产业呢？”
2SAM|20|20|约押 回答说：“不，我绝不吞灭和毁坏！
2SAM|20|21|话不是这么说的，只是因为有一个 以法莲 山区的人，就是 比基利 的儿子名叫 示巴 ，他举手攻击 大卫 王；你们只要把他一人交出来，我就离城而去。”妇人对 约押 说：“看哪，他的首级必从城墙上丢给你。”
2SAM|20|22|妇人凭她的智慧去劝众百姓，他们就割下 比基利 的儿子 示巴 的首级，丢给 约押 。 约押 吹角，众人就离城散开，各回自己的帐棚去了。 约押 回 耶路撒冷 ，到王那里。
2SAM|20|23|约押 统管 以色列 全军； 耶何耶大 的儿子 比拿雅 统管 基利提 人和 比利提 人；
2SAM|20|24|亚多兰 管理劳役的人； 亚希律 的儿子 约沙法 作史官；
2SAM|20|25|示法 作书记； 撒督 和 亚比亚他 作祭司；
2SAM|20|26|睚珥 人 以拉 也作 大卫 的祭司。
2SAM|21|1|大卫 在位年间有饥荒，一连三年， 大卫 求问耶和华，耶和华说：“ 扫罗 和他家犯了流人血之罪，因为他杀死了 基遍 人。”
2SAM|21|2|大卫 王召了 基遍 人来，跟他们说话。 基遍 人不是 以色列 人，而是 亚摩利 人中所剩下的人。 以色列 人曾向他们起誓， 扫罗 却为 以色列 人和 犹大 人大发热心，追杀他们，为了要消灭他们。
2SAM|21|3|大卫 对 基遍 人说：“我当为你们做什么呢？要用什么赎这罪，使你们为耶和华的产业祝福呢？”
2SAM|21|4|基遍 人对他说：“我们和 扫罗 以及他家的事与金银无关，也不要因我们的缘故杀任何 以色列 人。” 大卫 说：“你们怎样说，我就为你们怎样做。”
2SAM|21|5|他们对王说：“那谋害我们、要消灭我们、使我们不得住 以色列 境内的人，
2SAM|21|6|请把他的子孙七人交给我们，我们好在耶和华面前，把他们悬挂在 基比亚 ，就是耶和华拣选 扫罗 的地方。”王说：“我必交给你们。”
2SAM|21|7|王顾惜 扫罗 的孙子， 约拿单 的儿子 米非波设 ，因为在 大卫 和 扫罗 的儿子 约拿单 之间，有指着耶和华的誓言。
2SAM|21|8|王却把 爱亚 的女儿 利斯巴 为 扫罗 所生的两个儿子 亚摩尼 和 米非波设 ，以及 扫罗 的女儿 米拉 为 米何拉 人 巴西莱 儿子 亚得列 所生的五个儿子
2SAM|21|9|交在 基遍 人的手里。 基遍 人在耶和华面前把他们悬挂在山上，这七人就一起死了。他们被杀的时候正是收割的头几天，就是开始收割大麦的时候。
2SAM|21|10|爱亚 的女儿 利斯巴 用麻布铺在磐石上搭棚，从收割的开始直到天降雨在尸体上，她白日不许空中的飞鸟落在尸体上，夜间不让田野的走兽前来。
2SAM|21|11|有人把 扫罗 的妃子 爱亚 女儿 利斯巴 所做的事告诉 大卫 。
2SAM|21|12|大卫 就去，从 基列 的 雅比 人那里把 扫罗 和他儿子 约拿单 的骸骨搬来。先前 非利士 人在 基利波 杀了 扫罗 ，把尸体悬挂在 伯．珊 的广场上，后来 基列 的 雅比 人把尸体偷走。
2SAM|21|13|大卫 把 扫罗 和他儿子 约拿单 的骸骨从那里搬上来，又收殓了被悬挂的那些人的骸骨。
2SAM|21|14|他们将 扫罗 和他儿子 约拿单 的骸骨葬在 便雅悯 的 洗拉 ，在 扫罗 父亲 基士 的坟墓里。他们遵照王所吩咐的一切做了。此后上帝垂听了为那地的祈求。
2SAM|21|15|非利士 人与 以色列 人打仗。 大卫 带领仆人下去，与 非利士 人交战， 大卫 就疲乏了。
2SAM|21|16|巨人族的后裔 以实．比诺 说要杀 大卫 ；他的铜枪重三百舍客勒，腰间又佩着新刀 。
2SAM|21|17|但 洗鲁雅 的儿子 亚比筛 帮助 大卫 攻击 非利士 人，杀死了他。当日， 大卫 的人向 大卫 起誓说：“你不可再与我们一同出战，免得 以色列 的灯熄灭了。”
2SAM|21|18|后来，在 歌伯 又与 非利士 人打仗，那时 户沙 人 西比该 杀了巨人族的后裔 撒弗 。
2SAM|21|19|他们又在 歌伯 与 非利士 人打仗， 伯利恒 人 雅雷 的儿子 伊勒哈难 杀了 迦特 人 歌利亚 ；这人的枪杆粗如织布机的轴。
2SAM|21|20|又有一次，他们在 迦特 打仗。那里有一个身材高大的人，双手各有六根手指，双脚各有六根脚趾，共有二十四根；他也是巨人族的后裔。
2SAM|21|21|他向 以色列 骂阵， 大卫 的哥哥 示米亚 的儿子 约拿单 就杀了他。
2SAM|21|22|这四个人是 迦特 巨人族的后裔，都仆倒在 大卫 和他仆人的手下。
2SAM|22|1|当耶和华救 大卫 脱离所有仇敌和 扫罗 之手的日子，他用这诗的歌词向耶和华说话。
2SAM|22|2|他说： 耶和华是我的岩石、我的山寨、我的救主、
2SAM|22|3|我的上帝、我的磐石、我所投靠的。 他是我的盾牌，是拯救我的角， 是我的碉堡，是我的避难所， 是我的救主，救我脱离凶暴的。
2SAM|22|4|我要求告当赞美的耶和华， 我必从仇敌手中被救出来。
2SAM|22|5|死亡的波浪环绕我， 毁灭的急流惊吓我，
2SAM|22|6|阴间的绳索缠绕我， 死亡的圈套临到我。
2SAM|22|7|我在急难中求告耶和华， 向我的上帝呼求。 他从殿中听了我的声音； 我的呼求进入他的耳中。
2SAM|22|8|那时，因他发怒地就摇撼震动； 天的根基也战抖摇撼。
2SAM|22|9|他的鼻孔冒烟上腾； 他的口发火焚烧，连煤炭也烧着了。
2SAM|22|10|他使天下垂，亲自降临； 黑云在他脚下。
2SAM|22|11|他乘坐基路伯飞行， 在风的翅膀上显现。
2SAM|22|12|他以黑暗和聚集的水、 天空的密云为四围的行宫。
2SAM|22|13|因他发出光辉， 火炭都烧着了。
2SAM|22|14|耶和华在天上打雷； 至高者发出声音。
2SAM|22|15|他射出箭来，使仇敌四散； 发出闪电，击溃他们。
2SAM|22|16|耶和华的斥责一发，鼻孔的气一出， 海底就显现，大地的根基也暴露。
2SAM|22|17|他从高天伸手抓住我， 把我从大水中拉上来。
2SAM|22|18|他救我脱离我的强敌， 脱离那些恨我的人， 因为他们比我强盛。
2SAM|22|19|我遭遇灾难的日子，他们来攻击我； 但耶和华是我的倚靠。
2SAM|22|20|他领我到宽阔之处， 他救拔我，因他喜爱我。
2SAM|22|21|耶和华必按我的公义报答我， 按我手中的清洁赏赐我。
2SAM|22|22|因为我遵守耶和华的道， 未曾作恶离开我的上帝。
2SAM|22|23|他的一切典章在我面前， 他的律例我也未曾丢弃。
2SAM|22|24|我在他面前作了完全人， 我也持守自己远离罪孽。
2SAM|22|25|所以耶和华按我的公义， 在他眼前按我的清洁赏赐我。
2SAM|22|26|慈爱的人，你以慈爱待他； 完全的人，你以完善待他；
2SAM|22|27|清洁的人，你以清洁待他； 歪曲的人，你以弯曲待他。
2SAM|22|28|困苦的百姓，你必拯救； 但你的眼目察看高傲的人，使他们降卑。
2SAM|22|29|耶和华啊，你是我的灯； 耶和华必照明我的黑暗。
2SAM|22|30|我藉着你冲入敌军， 藉着我的上帝跳过城墙。
2SAM|22|31|至于上帝，他的道是完全的； 耶和华的话是纯净的。 凡投靠他的，他就作他们的盾牌。
2SAM|22|32|除了耶和华，谁是上帝呢？ 除了我们的上帝，谁是磐石呢？
2SAM|22|33|上帝是我坚固的保障， 他为我开完全的路。
2SAM|22|34|他使我的脚快如母鹿， 使我站稳在高处。
2SAM|22|35|他教导我的手能争战， 我的膀臂能开铜造的弓。
2SAM|22|36|你赐救恩给我作盾牌， 你的庇护 使我为大。
2SAM|22|37|你使我脚步宽阔， 我的脚踝未曾滑跌。
2SAM|22|38|我追赶我的仇敌，消灭他们； 若不将他们灭绝，我总不归回。
2SAM|22|39|我灭绝了他们， 打伤了他们，使他们站不起来； 他们都倒在我的脚下。
2SAM|22|40|你曾以力量束我的腰，使我能争战； 也曾使那起来攻击我的，都服在我以下。
2SAM|22|41|你又使我的仇敌在我面前转身逃跑， 使我能歼灭那恨我的人。
2SAM|22|42|他们仰望，却无人拯救； 就是呼求耶和华，他也不应允。
2SAM|22|43|我捣碎他们，如同地上的灰尘； 践踏压碎他们，如同街上的泥土。
2SAM|22|44|你救我脱离我百姓 的纷争， 保护我作列国的元首； 我素不认识的百姓必事奉我。
2SAM|22|45|外邦人要向我投降， 一听见我的名声就必顺从我。
2SAM|22|46|外邦人要丧胆， 战战兢兢地出营寨。
2SAM|22|47|耶和华永远活着。 愿我的磐石被称颂， 愿上帝－救我的磐石受尊崇。
2SAM|22|48|这位上帝为我伸冤， 使万民服在我以下。
2SAM|22|49|他救我脱离仇敌， 又把我举起，高过那些起来攻击我的人， 救我脱离残暴的人。
2SAM|22|50|耶和华啊，因此我要在列国中称谢你， 歌颂你的名。
2SAM|22|51|耶和华赐极大的救恩给他所立的王， 施慈爱给他的受膏者， 就是给 大卫 和他的后裔，直到永远！
2SAM|23|1|以下是 大卫 末了的话： “ 耶西 的儿子 大卫 的话， 得居高位的， 雅各 的上帝所膏的， 以色列 所喜爱的诗人的话。
2SAM|23|2|耶和华的灵藉着我说话， 他的言语在我的舌头上。
2SAM|23|3|以色列 的上帝说， 以色列 的磐石向我说： ‘那以公义治理人， 以敬畏上帝来治理的，
2SAM|23|4|他必像晨光， 如无云清晨的日出， 如雨后的光辉， 在嫩草地上。’
2SAM|23|5|我的家在上帝面前不是如此吗？ 上帝与我立永远的约， 这约既全备又稳妥。 我的一切救恩和我一切所想望的， 他岂不成全吗？
2SAM|23|6|但无赖全都像被丢弃的荆棘； 它们不能用手去拿；
2SAM|23|7|碰它们的人必须用铁器和枪杆， 它们必在那里被火烧尽。”
2SAM|23|8|大卫 勇士的名字如下： 哈革摩尼 人 约设．巴设 ，他是三勇士之首；他又名叫 伊斯尼 人 亚底挪 ，曾一次就杀了八百人 。
2SAM|23|9|跟随 大卫 的三勇士中，其次是 亚何亚 人 朵多 的儿子 以利亚撒 。从前 非利士 人聚集要打仗，他们向 非利士 人骂阵。 以色列 人上去的时候，
2SAM|23|10|他起来击杀 非利士 人，直到手臂疲乏，手粘住刀把。那日耶和华大获全胜，百姓跟在 以利亚撒 后面只顾夺取掠物。
2SAM|23|11|再其次是 哈拉 人 亚基 的儿子 沙玛 。一次， 非利士 人聚集在 利希 ，在一块长满红豆的田里，百姓在 非利士 人面前逃跑。
2SAM|23|12|沙玛 却站在那田的中间，防守那田，击败了 非利士 人。耶和华大获全胜。
2SAM|23|13|开始收割的时候，三个 侍卫 下到 亚杜兰洞 ，到 大卫 那里。 非利士 的军兵在 利乏音谷 安营。
2SAM|23|14|那时 大卫 在山寨， 非利士 人的驻军在 伯利恒 。
2SAM|23|15|大卫 渴想着说：“但愿有人从 伯利恒 城门旁的井里打水来给我喝！”
2SAM|23|16|这三个勇士就闯过 非利士 人的军营，从 伯利恒 城门旁的井里打水，拿来给 大卫 喝。他却不肯喝，将水浇在耶和华面前，
2SAM|23|17|说：“耶和华啊，我绝不做这事！这三个人冒生命的危险，这不是他们的血吗？” 大卫 不肯喝这水。这是三个勇士所做的事。
2SAM|23|18|洗鲁雅 的儿子， 约押 的兄弟 亚比筛 是这三个勇士的领袖；他曾举枪杀了三百人，就在三个勇士中得了名。
2SAM|23|19|他在这三个 勇士中是最有名望的，所以作他们的领袖，只是不及前三个勇士。
2SAM|23|20|耶何耶大 的儿子 比拿雅 是来自 甲薛 的勇士，曾行了大事。他杀了 摩押 人 亚利伊勒 的两个儿子，又在下雪的时候下到坑里去，杀了一只狮子。
2SAM|23|21|他又杀了一个魁梧的 埃及 人； 埃及 人手里拿着枪。 比拿雅 只拿着棍子下到他那里去，从 埃及 人手里夺过枪来，用那枪杀死了他。
2SAM|23|22|这些是 耶何耶大 的儿子 比拿雅 所做的事，就在三个勇士里得了名。
2SAM|23|23|他比那三十个勇士 更有名望，只是不及前三个勇士。 大卫 立他作护卫长。
2SAM|23|24|三十个勇士中有 约押 的兄弟 亚撒黑 ， 伯利恒 人 朵多 的儿子 伊勒哈难 ，
2SAM|23|25|哈律 人 沙玛 ， 哈律 人 以利加 ，
2SAM|23|26|帕勒提 人 希利斯 ， 提哥亚 人 益吉 的儿子 以拉 ，
2SAM|23|27|亚拿突 人 亚比以谢 ， 户沙 人 米本乃 ，
2SAM|23|28|亚何亚 人 撒们 ， 尼陀法 人 玛哈莱 ，
2SAM|23|29|尼陀法 人 巴拿 的儿子 希立 ， 便雅悯 族 基比亚 人 利拜 的儿子 以太 ，
2SAM|23|30|比拉顿 人 比拿雅 ， 迦实溪 人 希太 ，
2SAM|23|31|亚拉巴 人 亚比．亚本 ， 巴鲁米 人 押斯玛弗 ，
2SAM|23|32|沙本 人 以利雅哈巴 ， 雅善 儿子中的 约拿单 ，
2SAM|23|33|哈拉 人 沙玛 ， 哈拉 人 沙拉 的儿子 亚希暗 ，
2SAM|23|34|玛迦 人 亚哈拜 的儿子 以利法列 ， 基罗 人 亚希多弗 的儿子 以连 ，
2SAM|23|35|迦密 人 希斯莱 ， 亚巴 人 帕莱 ，
2SAM|23|36|琐巴 人 拿单 的儿子 以甲 ， 迦得 人 巴尼 ，
2SAM|23|37|亚扪 人 洗勒 ， 比录 人 拿哈莱 ，是给 洗鲁雅 的儿子 约押 拿兵器的，
2SAM|23|38|以帖 人 以拉 ， 以帖 人 迦立 ，
2SAM|23|39|赫 人 乌利亚 ，共三十七人。
2SAM|24|1|耶和华的怒气又向 以色列 发作，激起 大卫 来对付他们，说：“去，数点 以色列 人和 犹大 人。”
2SAM|24|2|大卫 对跟随他的 约押 元帅说：“你来回走遍 以色列 众支派，从 但 直到 别是巴 ，数点百姓，我好知道百姓的数目。”
2SAM|24|3|约押 对王说：“愿耶和华－你的上帝使百姓的数目增加百倍，使我主我王亲眼得见。我主我王何必要做这事呢？”
2SAM|24|4|但王坚持他对 约押 和众军官的命令。 约押 和众军官就从王面前出去，数点 以色列 的百姓。
2SAM|24|5|他们过 约旦河 ，在 迦得谷 中、城的右边 亚罗珥 安营，与 雅谢 相对。
2SAM|24|6|他们来到 基列 ，到了 他停．合示 地 ，又来到 但．雅安 ，绕到 西顿 。
2SAM|24|7|他们来到 推罗 的堡垒，以及 希未 人和 迦南 人的各城，又出来，到 犹大尼革夫 的 别是巴 。
2SAM|24|8|他们来回走遍全地，过了九个月又二十天，就回到 耶路撒冷 。
2SAM|24|9|约押 向王报告百姓的总数： 以色列 拿刀的勇士有八十万； 犹大 有五十万人。
2SAM|24|10|大卫 数点百姓以后，心中自责。大卫向耶和华说：“我做这事大大有罪了。耶和华啊，现在求你除掉仆人的罪孽，因我所做的非常愚昧。”
2SAM|24|11|大卫 早晨起来，耶和华的话临到 迦得 先知，就是 大卫 的先见，说：
2SAM|24|12|“你去告诉 大卫 ：‘耶和华如此说：我向你提出三样，随你选择一样，我好降给你。’”
2SAM|24|13|于是 迦得 来到 大卫 那里告诉他，问他：“你要国中有七 年的饥荒呢？或是你在敌人面前逃跑，被追赶三个月呢？或是在你国中有三日的瘟疫呢？现在你要考虑思量，我怎样去回覆那差我来的。”
2SAM|24|14|大卫 对 迦得 说：“我很为难。我们宁愿落在耶和华的手里，因为他有丰盛的怜悯；我不愿落在人的手里。”
2SAM|24|15|于是，耶和华降瘟疫给 以色列 。自早晨到所定的时候，从 但 直到 别是巴 ，百姓中死了七万人。
2SAM|24|16|天使向 耶路撒冷 伸手要毁灭这城的时候，耶和华改变心意，不降那灾难，就对那在百姓中施行毁灭的天使说：“够了！住手吧！”耶和华的使者正在 耶布斯 人 亚劳拿 的禾场那里。
2SAM|24|17|大卫 看见那在百姓中施行毁灭的天使，就向耶和华说：“看哪，我犯了罪，行了恶，但这群羊做了什么呢？愿你的手攻击我和我的父家。”
2SAM|24|18|当日， 迦得 来到 大卫 那里，对他说：“你上去，在 耶布斯 人 亚劳拿 的禾场上为耶和华立一座坛。”
2SAM|24|19|大卫 就照着 迦得 的话，照着耶和华所吩咐的上去了。
2SAM|24|20|亚劳拿 观看，看见王和臣仆向他走过来。 亚劳拿 就出去，脸伏于地，向王下拜。
2SAM|24|21|亚劳拿 说：“我主我王为何来到仆人这里呢？” 大卫 说：“我要买你这禾场，为耶和华筑一座坛，使瘟疫在百姓中停止。”
2SAM|24|22|亚劳拿 对 大卫 说：“我主我王，你眼中看为好，就拿去献祭。看，这里有牛可以作燔祭，有打粮的器具和套牛的轭可以当作柴。
2SAM|24|23|王啊，这一切， 亚劳拿 都献给王。” 亚劳拿 又对王说：“愿耶和华－你的上帝悦纳你。”
2SAM|24|24|王对 亚劳拿 说：“不，我一定要按价钱向你买；我不能用白白得来的东西作燔祭献给耶和华－我的上帝。” 大卫 就用五十舍客勒银子买了那禾场与牛。
2SAM|24|25|大卫 在那里为耶和华筑了一座坛，献燔祭和平安祭。耶和华垂听了为那地的祈求，瘟疫就在 以色列 中停止了。
