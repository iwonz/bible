EZEK|1|1|In the thirtieth year, in the fourth month, on the fifth day of the month, as I was among the exiles by the Chebar canal, the heavens were opened, and I saw visions of God.
EZEK|1|2|On the fifth day of the month (it was the fifth year of the exile of King Jehoiachin),
EZEK|1|3|the word of the LORD came to Ezekiel the priest, the son of Buzi, in the land of the Chaldeans by the Chebar canal, and the hand of the LORD was upon him there.
EZEK|1|4|As I looked, behold, a stormy wind came out of the north, and a great cloud, with brightness around it, and fire flashing forth continually, and in the midst of the fire, as it were gleaming metal.
EZEK|1|5|And from the midst of it came the likeness of four living creatures. And this was their appearance: they had a human likeness,
EZEK|1|6|but each had four faces, and each of them had four wings.
EZEK|1|7|Their legs were straight, and the soles of their feet were like the sole of a calf's foot. And they sparkled like burnished bronze.
EZEK|1|8|Under their wings on their four sides they had human hands. And the four had their faces and their wings thus:
EZEK|1|9|their wings touched one another. Each one of them went straight forward, without turning as they went.
EZEK|1|10|As for the likeness of their faces, each had a human face. The four had the face of a lion on the right side, the four had the face of an ox on the left side, and the four had the face of an eagle.
EZEK|1|11|Such were their faces. And their wings were spread out above. Each creature had two wings, each of which touched the wing of another, while two covered their bodies.
EZEK|1|12|And each went straight forward. Wherever the spirit would go, they went, without turning as they went.
EZEK|1|13|As for the likeness of the living creatures, their appearance was like burning coals of fire, like the appearance of torches moving to and fro among the living creatures. And the fire was bright, and out of the fire went forth lightning.
EZEK|1|14|And the living creatures darted to and fro, like the appearance of a flash of lightning.
EZEK|1|15|Now as I looked at the living creatures, I saw a wheel on the earth beside the living creatures, one for each of the four of them.
EZEK|1|16|As for the appearance of the wheels and their construction: their appearance was like the gleaming of beryl. And the four had the same likeness, their appearance and construction being as it were a wheel within a wheel.
EZEK|1|17|When they went, they went in any of their four directions without turning as they went.
EZEK|1|18|And their rims were tall and awesome, and the rims of all four were full of eyes all around.
EZEK|1|19|And when the living creatures went, the wheels went beside them; and when the living creatures rose from the earth, the wheels rose.
EZEK|1|20|Wherever the spirit wanted to go, they went, and the wheels rose along with them, for the spirit of the living creatures was in the wheels.
EZEK|1|21|When those went, these went; and when those stood, these stood; and when those rose from the earth, the wheels rose along with them, for the spirit of the living creatures was in the wheels.
EZEK|1|22|Over the heads of the living creatures there was the likeness of an expanse, shining like awe-inspiring crystal, spread out above their heads.
EZEK|1|23|And under the expanse their wings were stretched out straight, one toward another. And each creature had two wings covering its body.
EZEK|1|24|And when they went, I heard the sound of their wings like the sound of many waters, like the sound of the Almighty, a sound of tumult like the sound of an army. When they stood still, they let down their wings.
EZEK|1|25|And there came a voice from above the expanse over their heads. When they stood still, they let down their wings.
EZEK|1|26|And above the expanse over their heads there was the likeness of a throne, in appearance like sapphire; and seated above the likeness of a throne was a likeness with a human appearance.
EZEK|1|27|And upward from what had the appearance of his waist I saw as it were gleaming metal, like the appearance of fire enclosed all around. And downward from what had the appearance of his waist I saw as it were the appearance of fire, and there was brightness around him.
EZEK|1|28|Like the appearance of the bow that is in the cloud on the day of rain, so was the appearance of the brightness all around. Such was the appearance of the likeness of the glory of the LORD. And when I saw it, I fell on my face, and I heard the voice of one speaking.
EZEK|2|1|And he said to me, "Son of man, stand on your feet, and I will speak with you."
EZEK|2|2|And as he spoke to me, the Spirit entered into me and set me on my feet, and I heard him speaking to me.
EZEK|2|3|And he said to me, "Son of man, I send you to the people of Israel, to nations of rebels, who have rebelled against me. They and their fathers have transgressed against me to this very day.
EZEK|2|4|The descendants also are impudent and stubborn: I send you to them, and you shall say to them, 'Thus says the Lord GOD.'
EZEK|2|5|And whether they hear or refuse to hear (for they are a rebellious house) they will know that a prophet has been among them.
EZEK|2|6|And you, son of man, be not afraid of them, nor be afraid of their words, though briers and thorns are with you and you sit on scorpions. Be not afraid of their words, nor be dismayed at their looks, for they are a rebellious house.
EZEK|2|7|And you shall speak my words to them, whether they hear or refuse to hear, for they are a rebellious house.
EZEK|2|8|"But you, son of man, hear what I say to you. Be not rebellious like that rebellious house; open your mouth and eat what I give you."
EZEK|2|9|And when I looked, behold, a hand was stretched out to me, and behold, a scroll of a book was in it.
EZEK|2|10|And he spread it before me. And it had writing on the front and on the back, and there were written on it words of lamentation and mourning and woe.
EZEK|3|1|And he said to me, "Son of man, eat whatever you find here. Eat this scroll, and go, speak to the house of Israel."
EZEK|3|2|So I opened my mouth, and he gave me this scroll to eat.
EZEK|3|3|And he said to me, "Son of man, feed your belly with this scroll that I give you and fill your stomach with it." Then I ate it, and it was in my mouth as sweet as honey.
EZEK|3|4|And he said to me, "Son of man, go to the house of Israel and speak with my words to them.
EZEK|3|5|For you are not sent to a people of foreign speech and a hard language, but to the house of Israel-
EZEK|3|6|not to many peoples of foreign speech and a hard language, whose words you cannot understand. Surely, if I sent you to such, they would listen to you.
EZEK|3|7|But the house of Israel will not be willing to listen to you, for they are not willing to listen to me. Because all the house of Israel have a hard forehead and a stubborn heart.
EZEK|3|8|Behold, I have made your face as hard as their faces, and your forehead as hard as their foreheads.
EZEK|3|9|Like emery harder than flint have I made your forehead. Fear them not, nor be dismayed at their looks, for they are a rebellious house."
EZEK|3|10|Moreover, he said to me, "Son of man, all my words that I shall speak to you receive in your heart, and hear with your ears.
EZEK|3|11|And go to the exiles, to your people, and speak to them and say to them, 'Thus says the Lord GOD,' whether they hear or refuse to hear."
EZEK|3|12|Then the Spirit lifted me up, and I heard behind me the voice of a great earthquake: "Blessed be the glory of the LORD from its place!"
EZEK|3|13|It was the sound of the wings of the living creatures as they touched one another, and the sound of the wheels beside them, and the sound of a great earthquake.
EZEK|3|14|The Spirit lifted me up and took me away, and I went in bitterness in the heat of my spirit, the hand of the LORD being strong upon me.
EZEK|3|15|And I came to the exiles at Tel-abib, who were dwelling by the Chebar canal, and I sat where they were dwelling. And I sat there overwhelmed among them seven days.
EZEK|3|16|And at the end of seven days, the word of the LORD came to me:
EZEK|3|17|"Son of man, I have made you a watchman for the house of Israel. Whenever you hear a word from my mouth, you shall give them warning from me.
EZEK|3|18|If I say to the wicked, 'You shall surely die,' and you give him no warning, nor speak to warn the wicked from his wicked way, in order to save his life, that wicked person shall die for his iniquity, but his blood I will require at your hand.
EZEK|3|19|But if you warn the wicked, and he does not turn from his wickedness, or from his wicked way, he shall die for his iniquity, but you will have delivered your soul.
EZEK|3|20|Again, if a righteous person turns from his righteousness and commits injustice, and I lay a stumbling block before him, he shall die. Because you have not warned him, he shall die for his sin, and his righteous deeds that he has done shall not be remembered, but his blood I will require at your hand.
EZEK|3|21|But if you warn the righteous person not to sin, and he does not sin, he shall surely live, because he took warning, and you will have delivered your soul."
EZEK|3|22|And the hand of the LORD was upon me there. And he said to me, "Arise, go out into the valley, and there I will speak with you."
EZEK|3|23|So I arose and went out into the valley, and behold, the glory of the LORD stood there, like the glory that I had seen by the Chebar canal, and I fell on my face.
EZEK|3|24|But the Spirit entered into me and set me on my feet, and he spoke with me and said to me, "Go, shut yourself within your house.
EZEK|3|25|And you, O son of man, behold, cords will be placed upon you, and you shall be bound with them, so that you cannot go out among the people.
EZEK|3|26|And I will make your tongue cling to the roof of your mouth, so that you shall be mute and unable to reprove them, for they are a rebellious house.
EZEK|3|27|But when I speak with you, I will open your mouth, and you shall say to them, 'Thus says the Lord GOD.' He who will hear, let him hear; and he who will refuse to hear, let him refuse, for they are a rebellious house.
EZEK|4|1|"And you, son of man, take a brick and lay it before you, and engrave on it a city, even Jerusalem.
EZEK|4|2|And put siegeworks against it, and build a siege wall against it, and cast up a mound against it. Set camps also against it, and plant battering rams against it all around.
EZEK|4|3|And you, take an iron griddle, and place it as an iron wall between you and the city; and set your face toward it, and let it be in a state of siege, and press the siege against it. This is a sign for the house of Israel.
EZEK|4|4|"Then lie on your left side, and place the punishment of the house of Israel upon it. For the number of the days that you lie on it, you shall bear their punishment.
EZEK|4|5|For I assign to you a number of days, 390 days, equal to the number of the years of their punishment. So long shall you bear the punishment of the house of Israel.
EZEK|4|6|And when you have completed these, you shall lie down a second time, but on your right side, and bear the punishment of the house of Judah. Forty days I assign you, a day for each year.
EZEK|4|7|And you shall set your face toward the siege of Jerusalem, with your arm bared, and you shall prophesy against the city.
EZEK|4|8|And behold, I will place cords upon you, so that you cannot turn from one side to the other, till you have completed the days of your siege.
EZEK|4|9|"And you, take wheat and barley, beans and lentils, millet and emmer, and put them into a single vessel and make your bread from them. During the number of days that you lie on your side, 390 days, you shall eat it.
EZEK|4|10|And your food that you eat shall be by weight, twenty shekels a day; from day to day you shall eat it.
EZEK|4|11|And water you shall drink by measure, the sixth part of a hin; from day to day you shall drink.
EZEK|4|12|And you shall eat it as a barley cake, baking it in their sight on human dung."
EZEK|4|13|And the LORD said, "Thus shall the people of Israel eat their bread unclean, among the nations where I will drive them."
EZEK|4|14|Then I said, "Ah, Lord GOD! Behold, I have never defiled myself. From my youth up till now I have never eaten what died of itself or was torn by beasts, nor has tainted meat come into my mouth."
EZEK|4|15|Then he said to me, "See, I assign to you cow's dung instead of human dung, on which you may prepare your bread."
EZEK|4|16|Moreover, he said to me, "Son of man, behold, I will break the supply of bread in Jerusalem. They shall eat bread by weight and with anxiety, and they shall drink water by measure and in dismay.
EZEK|4|17|I will do this that they may lack bread and water, and look at one another in dismay, and rot away because of their punishment.
EZEK|5|1|"And you, O son of man, take a sharp sword. Use it as a barber's razor and pass it over your head and your beard. Then take balances for weighing and divide the hair.
EZEK|5|2|A third part you shall burn in the fire in the midst of the city, when the days of the siege are completed. And a third part you shall take and strike with the sword all around the city. And a third part you shall scatter to the wind, and I will unsheathe the sword after them.
EZEK|5|3|And you shall take from these a small number and bind them in the skirts of your robe.
EZEK|5|4|And of these again you shall take some and cast them into the midst of the fire and burn them in the fire. From there a fire will come out into all the house of Israel.
EZEK|5|5|"Thus says the Lord GOD: This is Jerusalem. I have set her in the center of the nations, with countries all around her.
EZEK|5|6|And she has rebelled against my rules by doing wickedness more than the nations, and against my statutes more than the countries all around her; for they have rejected my rules and have not walked in my statutes.
EZEK|5|7|Therefore thus says the Lord GOD: Because you are more turbulent than the nations that are all around you, and have not walked in my statutes or obeyed my rules, and have not even acted according to the rules of the nations that are all around you,
EZEK|5|8|therefore thus says the Lord GOD: Behold, I, even I, am against you. And I will execute judgments in your midst in the sight of the nations.
EZEK|5|9|And because of all your abominations I will do with you what I have never yet done, and the like of which I will never do again.
EZEK|5|10|Therefore fathers shall eat their sons in your midst, and sons shall eat their fathers. And I will execute judgments on you, and any of you who survive I will scatter to all the winds.
EZEK|5|11|Therefore, as I live, declares the Lord GOD, surely, because you have defiled my sanctuary with all your detestable things and with all your abominations, therefore I will withdraw. My eye will not spare, and I will have no pity.
EZEK|5|12|A third part of you shall die of pestilence and be consumed with famine in your midst; a third part shall fall by the sword all around you; and a third part I will scatter to all the winds and will unsheathe the sword after them.
EZEK|5|13|"Thus shall my anger spend itself, and I will vent my fury upon them and satisfy myself. And they shall know that I am the LORD- that I have spoken in my jealousy- when I spend my fury upon them.
EZEK|5|14|Moreover, I will make you a desolation and an object of reproach among the nations all around you and in the sight of all who pass by.
EZEK|5|15|You shall be a reproach and a taunt, a warning and a horror, to the nations all around you, when I execute judgments on you in anger and fury, and with furious rebukes- I am the LORD, I have spoken-
EZEK|5|16|when I send against you the deadly arrows of famine, arrows for destruction, which I will send to destroy you, and when I bring more and more famine upon you and break your supply of bread.
EZEK|5|17|I will send famine and wild beasts against you, and they will rob you of your children. Pestilence and blood shall pass through you, and I will bring the sword upon you. I am the LORD; I have spoken."
EZEK|6|1|The word of the LORD came to me:
EZEK|6|2|"Son of man, set your face toward the mountains of Israel, and prophesy against them,
EZEK|6|3|and say, You mountains of Israel, hear the word of the Lord GOD! Thus says the Lord GOD to the mountains and the hills, to the ravines and the valleys: Behold, I, even I, will bring a sword upon you, and I will destroy your high places.
EZEK|6|4|Your altars shall become desolate, and your incense altars shall be broken, and I will cast down your slain before your idols.
EZEK|6|5|And I will lay the dead bodies of the people of Israel before their idols, and I will scatter your bones around your altars.
EZEK|6|6|Wherever you dwell, the cities shall be waste and the high places ruined, so that your altars will be waste and ruined, your idols broken and destroyed, your incense altars cut down, and your works wiped out.
EZEK|6|7|And the slain shall fall in your midst, and you shall know that I am the LORD.
EZEK|6|8|"Yet I will leave some of you alive. When you have among the nations some who escape the sword, and when you are scattered through the countries,
EZEK|6|9|then those of you who escape will remember me among the nations where they are carried captive, how I have been broken over their whoring heart that has departed from me and over their eyes that go whoring after their idols. And they will be loathsome in their own sight for the evils that they have committed, for all their abominations.
EZEK|6|10|And they shall know that I am the LORD. I have not said in vain that I would do this evil to them."
EZEK|6|11|Thus says the Lord GOD: "Clap your hands and stamp your foot and say, Alas, because of all the evil abominations of the house of Israel, for they shall fall by the sword, by famine, and by pestilence.
EZEK|6|12|He who is far off shall die of pestilence, and he who is near shall fall by the sword, and he who is left and is preserved shall die of famine. Thus I will spend my fury upon them.
EZEK|6|13|And you shall know that I am the LORD, when their slain lie among their idols around their altars, on every high hill, on all the mountaintops, under every green tree, and under every leafy oak, wherever they offered pleasing aroma to all their idols.
EZEK|6|14|And I will stretch out my hand against them and make the land desolate and waste, in all their dwelling places, from the wilderness to Riblah. Then they will know that I am the LORD."
EZEK|7|1|The word of the LORD came to me:
EZEK|7|2|"And you, O son of man, thus says the Lord GOD to the land of Israel: An end! The end has come upon the four corners of the land.
EZEK|7|3|Now the end is upon you, and I will send my anger upon you; I will judge you according to your ways, and I will punish you for all your abominations.
EZEK|7|4|And my eye will not spare you, nor will I have pity, but I will punish you for your ways, while your abominations are in your midst. Then you will know that I am the LORD.
EZEK|7|5|"Thus says the Lord GOD: Disaster after disaster! Behold, it comes.
EZEK|7|6|An end has come; the end has come; it has awakened against you. Behold, it comes.
EZEK|7|7|Your doom has come to you, O inhabitant of the land. The time has come; the day is near, a day of tumult, and not of joyful shouting on the mountains.
EZEK|7|8|Now I will soon pour out my wrath upon you, and spend my anger against you, and judge you according to your ways, and I will punish you for all your abominations.
EZEK|7|9|And my eye will not spare, nor will I have pity. I will punish you according to your ways, while your abominations are in your midst. Then you will know that I am the LORD, who strikes.
EZEK|7|10|"Behold, the day! Behold, it comes! Your doom has come; the rod has blossomed; pride has budded.
EZEK|7|11|Violence has grown up into a rod of wickedness. None of them shall remain, nor their abundance, nor their wealth; neither shall there be preeminence among them.
EZEK|7|12|The time has come; the day has arrived. Let not the buyer rejoice, nor the seller mourn, for wrath is upon all their multitude.
EZEK|7|13|For the seller shall not return to what he has sold, while they live. For the vision concerns all their multitude; it shall not turn back; and because of his iniquity, none can maintain his life.
EZEK|7|14|"They have blown the trumpet and made everything ready, but none goes to battle, for my wrath is upon all their multitude.
EZEK|7|15|The sword is without; pestilence and famine are within. He who is in the field dies by the sword, and him who is in the city famine and pestilence devour.
EZEK|7|16|And if any survivors escape, they will be on the mountains, like doves of the valleys, all of them moaning, each one over his iniquity.
EZEK|7|17|All hands are feeble, and all knees turn to water.
EZEK|7|18|They put on sackcloth, and horror covers them. Shame is on all faces, and baldness on all their heads.
EZEK|7|19|They cast their silver into the streets, and their gold is like an unclean thing. Their silver and gold are not able to deliver them in the day of the wrath of the LORD. They cannot satisfy their hunger or fill their stomachs with it. For it was the stumbling block of their iniquity.
EZEK|7|20|His beautiful ornament they used for pride, and they made their abominable images and their detestable things of it. Therefore I make it an unclean thing to them.
EZEK|7|21|And I will give it into the hands of foreigners for prey, and to the wicked of the earth for spoil, and they shall profane it.
EZEK|7|22|I will turn my face from them, and they shall profane my treasured place. Robbers shall enter and profane it.
EZEK|7|23|"Forge a chain! For the land is full of bloody crimes and the city is full of violence.
EZEK|7|24|I will bring the worst of the nations to take possession of their houses. I will put an end to the pride of the strong, and their holy places shall be profaned.
EZEK|7|25|When anguish comes, they will seek peace, but there shall be none.
EZEK|7|26|Disaster comes upon disaster; rumor follows rumor. They seek a vision from the prophet, while the law perishes from the priest and counsel from the elders.
EZEK|7|27|The king mourns, the prince is wrapped in despair, and the hands of the people of the land are paralyzed by terror. According to their way I will do to them, and according to their judgments I will judge them, and they shall know that I am the LORD."
EZEK|8|1|In the sixth year, in the sixth month, on the fifth day of the month, as I sat in my house, with the elders of Judah sitting before me, the hand of the Lord GOD fell upon me there.
EZEK|8|2|Then I looked, and behold, a form that had the appearance of a man. Below what appeared to be his waist was fire, and above his waist was something like the appearance of brightness, like gleaming metal.
EZEK|8|3|He put out the form of a hand and took me by a lock of my head, and the Spirit lifted me up between earth and heaven and brought me in visions of God to Jerusalem, to the entrance of the gateway of the inner court that faces north, where was the seat of the image of jealousy, which provokes to jealousy.
EZEK|8|4|And behold, the glory of the God of Israel was there, like the vision that I saw in the valley.
EZEK|8|5|Then he said to me, "Son of man, lift up your eyes now toward the north." So I lifted up my eyes toward the north, and behold, north of the altar gate, in the entrance, was this image of jealousy.
EZEK|8|6|And he said to me, "Son of man, do you see what they are doing, the great abominations that the house of Israel are committing here, to drive me far from my sanctuary? But you will see still greater abominations."
EZEK|8|7|And he brought me to the entrance of the court, and when I looked, behold, there was a hole in the wall.
EZEK|8|8|Then he said to me, "Son of man, dig in the wall." So I dug in the wall, and behold, there was an entrance.
EZEK|8|9|And he said to me, "Go in, and see the vile abominations that they are committing here."
EZEK|8|10|So I went in and saw. And there, engraved on the wall all around, was every form of creeping things and loathsome beasts, and all the idols of the house of Israel.
EZEK|8|11|And before them stood seventy men of the elders of the house of Israel, with Jaazaniah the son of Shaphan standing among them. Each had his censer in his hand, and the smoke of the cloud of incense went up.
EZEK|8|12|Then he said to me, "Son of man, have you seen what the elders of the house of Israel are doing in the dark, each in his room of pictures? For they say, 'The LORD does not see us, the LORD has forsaken the land.'"
EZEK|8|13|He said also to me, "You will see still greater abominations that they commit."
EZEK|8|14|Then he brought me to the entrance of the north gate of the house of the LORD, and behold, there sat women weeping for Tammuz.
EZEK|8|15|Then he said to me, "Have you seen this, O son of man? You will see still greater abominations than these."
EZEK|8|16|And he brought me into the inner court of the house of the LORD. And behold, at the entrance of the temple of the LORD, between the porch and the altar, were about twenty-five men, with their backs to the temple of the LORD, and their faces toward the east, worshiping the sun toward the east.
EZEK|8|17|Then he said to me, "Have you seen this, O son of man? Is it too light a thing for the house of Judah to commit the abominations that they commit here, that they should fill the land with violence and provoke me still further to anger? Behold, they put the branch to their nose.
EZEK|8|18|Therefore I will act in wrath. My eye will not spare, nor will I have pity. And though they cry in my ears with a loud voice, I will not hear them."
EZEK|9|1|Then he cried in my ears with a loud voice, saying, "Bring near the executioners of the city, each with his destroying weapon in his hand."
EZEK|9|2|And behold, six men came from the direction of the upper gate, which faces north, each with his weapon for slaughter in his hand, and with them was a man clothed in linen, with a writing case at his waist. And they went in and stood beside the bronze altar.
EZEK|9|3|Now the glory of the God of Israel had gone up from the cherub on which it rested to the threshold of the house. And he called to the man clothed in linen, who had the writing case at his waist.
EZEK|9|4|And the LORD said to him, "Pass through the city, through Jerusalem, and put a mark on the foreheads of the men who sigh and groan over all the abominations that are committed in it."
EZEK|9|5|And to the others he said in my hearing, "Pass through the city after him, and strike. Your eye shall not spare, and you shall show no pity.
EZEK|9|6|Kill old men outright, young men and maidens, little children and women, but touch no one on whom is the mark. And begin at my sanctuary." So they began with the elders who were before the house.
EZEK|9|7|Then he said to them, "Defile the house, and fill the courts with the slain. Go out." So they went out and struck in the city.
EZEK|9|8|And while they were striking, and I was left alone, I fell upon my face, and cried, "Ah, Lord GOD! Will you destroy all the remnant of Israel in the outpouring of your wrath on Jerusalem?"
EZEK|9|9|Then he said to me, "The guilt of the house of Israel and Judah is exceedingly great. The land is full of blood, and the city full of injustice. For they say, 'The LORD has forsaken the land, and the LORD does not see.'
EZEK|9|10|As for me, my eye will not spare, nor will I have pity; I will bring their deeds upon their heads."
EZEK|9|11|And behold, the man clothed in linen, with the writing case at his waist, brought back word, saying, "I have done as you commanded me."
EZEK|10|1|Then I looked, and behold, on the expanse that was over the heads of the cherubim there appeared above them something like a sapphire, in appearance like a throne.
EZEK|10|2|And he said to the man clothed in linen, "Go in among the whirling wheels underneath the cherubim. Fill your hands with burning coals from between the cherubim, and scatter them over the city." And he went in before my eyes.
EZEK|10|3|Now the cherubim were standing on the south side of the house, when the man went in, and a cloud filled the inner court.
EZEK|10|4|And the glory of the LORD went up from the cherub to the threshold of the house, and the house was filled with the cloud, and the court was filled with the brightness of the glory of the LORD.
EZEK|10|5|And the sound of the wings of the cherubim was heard as far as the outer court, like the voice of God Almighty when he speaks.
EZEK|10|6|And when he commanded the man clothed in linen, "Take fire from between the whirling wheels, from between the cherubim," he went in and stood beside a wheel.
EZEK|10|7|And a cherub stretched out his hand from between the cherubim to the fire that was between the cherubim, and took some of it and put it into the hands of the man clothed in linen, who took it and went out.
EZEK|10|8|The cherubim appeared to have the form of a human hand under their wings.
EZEK|10|9|And I looked, and behold, there were four wheels beside the cherubim, one beside each cherub, and the appearance of the wheels was like sparkling beryl.
EZEK|10|10|And as for their appearance, the four had the same likeness, as if a wheel were within a wheel.
EZEK|10|11|When they went, they went in any of their four directions without turning as they went, but in whatever direction the front wheel faced, the others followed without turning as they went.
EZEK|10|12|And their whole body, their rims, and their spokes, their wings, and the wheels were full of eyes all around- the wheels that the four of them had.
EZEK|10|13|As for the wheels, they were called in my hearing "the whirling wheels."
EZEK|10|14|And every one had four faces: the first face was the face of the cherub, and the second face was a human face, and the third the face of a lion, and the fourth the face of an eagle.
EZEK|10|15|And the cherubim mounted up. These were the living creatures that I saw by the Chebar canal.
EZEK|10|16|And when the cherubim went, the wheels went beside them. And when the cherubim lifted up their wings to mount up from the earth, the wheels did not turn from beside them.
EZEK|10|17|When they stood still, these stood still, and when they mounted up, these mounted up with them, for the spirit of the living creatures was in them.
EZEK|10|18|Then the glory of the LORD went out from the threshold of the house, and stood over the cherubim.
EZEK|10|19|And the cherubim lifted up their wings and mounted up from the earth before my eyes as they went out, with the wheels beside them. And they stood at the entrance of the east gate of the house of the LORD, and the glory of the God of Israel was over them.
EZEK|10|20|These were the living creatures that I saw underneath the God of Israel by the Chebar canal; and I knew that they were cherubim.
EZEK|10|21|Each had four faces, and each four wings, and underneath their wings the likeness of human hands.
EZEK|10|22|And as for the likeness of their faces, they were the same faces whose appearance I had seen by the Chebar canal. Each one of them went straight forward.
EZEK|11|1|The Spirit lifted me up and brought me to the east gate of the house of the LORD, which faces east. And behold, at the entrance of the gateway there were twenty-five men. And I saw among them Jaazaniah the son of Azzur, and Pelatiah the son of Benaiah, princes of the people.
EZEK|11|2|And he said to me, "Son of man, these are the men who devise iniquity and who give wicked counsel in this city;
EZEK|11|3|who say, 'The time is not near to build houses. This city is the cauldron, and we are the meat.'
EZEK|11|4|Therefore prophesy against them, prophesy, O son of man."
EZEK|11|5|And the Spirit of the LORD fell upon me, and he said to me, "Say, Thus says the LORD: So you think, O house of Israel. For I know the things that come into your mind.
EZEK|11|6|You have multiplied your slain in this city and have filled its streets with the slain.
EZEK|11|7|Therefore thus says the Lord GOD: Your slain whom you have laid in the midst of it, they are the meat, and this city is the cauldron, but you shall be brought out of the midst of it.
EZEK|11|8|You have feared the sword, and I will bring the sword upon you, declares the Lord GOD.
EZEK|11|9|And I will bring you out of the midst of it, and give you into the hands of foreigners, and execute judgments upon you.
EZEK|11|10|You shall fall by the sword. I will judge you at the border of Israel, and you shall know that I am the LORD.
EZEK|11|11|This city shall not be your cauldron, nor shall you be the meat in the midst of it. I will judge you at the border of Israel,
EZEK|11|12|and you shall know that I am the LORD. For you have not walked in my statutes, nor obeyed my rules, but have acted according to the rules of the nations that are around you."
EZEK|11|13|And it came to pass, while I was prophesying, that Pelatiah the son of Benaiah died. Then I fell down on my face and cried out with a loud voice and said, "Ah, Lord GOD! Will you make a full end of the remnant of Israel?"
EZEK|11|14|And the word of the LORD came to me:
EZEK|11|15|"Son of man, your brothers, even your brothers, your kinsmen, the whole house of Israel, all of them, are those of whom the inhabitants of Jerusalem have said, 'Go far from the LORD; to us this land is given for a possession.'
EZEK|11|16|Therefore say, 'Thus says the Lord GOD: Though I removed them far off among the nations, and though I scattered them among the countries, yet I have been a sanctuary to them for a while in the countries where they have gone.'
EZEK|11|17|Therefore say, 'Thus says the Lord GOD: I will gather you from the peoples and assemble you out of the countries where you have been scattered, and I will give you the land of Israel.'
EZEK|11|18|And when they come there, they will remove from it all its detestable things and all its abominations.
EZEK|11|19|And I will give them one heart, and a new spirit I will put within them. I will remove the heart of stone from their flesh and give them a heart of flesh,
EZEK|11|20|that they may walk in my statutes and keep my rules and obey them. And they shall be my people, and I will be their God.
EZEK|11|21|But as for those whose heart goes after their detestable things and their abominations, I will bring their deeds upon their own heads, declares the Lord GOD."
EZEK|11|22|Then the cherubim lifted up their wings, with the wheels beside them, and the glory of the God of Israel was over them.
EZEK|11|23|And the glory of the LORD went up from the midst of the city and stood on the mountain that is on the east side of the city.
EZEK|11|24|And the Spirit lifted me up and brought me in the vision by the Spirit of God into Chaldea, to the exiles. Then the vision that I had seen went up from me.
EZEK|11|25|And I told the exiles all the things that the LORD had shown me.
EZEK|12|1|The word of the LORD came to me:
EZEK|12|2|"Son of man, you dwell in the midst of a rebellious house, who have eyes to see, but see not, who have ears to hear, but hear not, for they are a rebellious house.
EZEK|12|3|As for you, son of man, prepare for yourself an exile's baggage, and go into exile by day in their sight. You shall go like an exile from your place to another place in their sight. Perhaps they will understand, though they are a rebellious house.
EZEK|12|4|You shall bring out your baggage by day in their sight, as baggage for exile, and you shall go out yourself at evening in their sight, as those do who must go into exile.
EZEK|12|5|In their sight dig through the wall, and bring your baggage out through it.
EZEK|12|6|In their sight you shall lift the baggage upon your shoulder and carry it out at dusk. You shall cover your face that you may not see the land, for I have made you a sign for the house of Israel."
EZEK|12|7|And I did as I was commanded. I brought out my baggage by day, as baggage for exile, and in the evening I dug through the wall with my own hands. I brought out my baggage at dusk, carrying it on my shoulder in their sight.
EZEK|12|8|In the morning the word of the LORD came to me:
EZEK|12|9|"Son of man, has not the house of Israel, the rebellious house, said to you, 'What are you doing?'
EZEK|12|10|Say to them, 'Thus says the Lord GOD: This oracle concerns the prince in Jerusalem and all the house of Israel who are in it.'
EZEK|12|11|Say, 'I am a sign for you: as I have done, so shall it be done to them. They shall go into exile, into captivity.'
EZEK|12|12|And the prince who is among them shall lift his baggage upon his shoulder at dusk, and shall go out. They shall dig through the wall to bring him out through it. He shall cover his face, that he may not see the land with his eyes.
EZEK|12|13|And I will spread my net over him, and he shall be taken in my snare. And I will bring him to Babylon, the land of the Chaldeans, yet he shall not see it, and he shall die there.
EZEK|12|14|And I will scatter toward every wind all who are around him, his helpers and all his troops, and I will unsheathe the sword after them.
EZEK|12|15|And they shall know that I am the LORD, when I disperse them among the nations and scatter them among the countries.
EZEK|12|16|But I will let a few of them escape from the sword, from famine and pestilence, that they may declare all their abominations among the nations where they go, and may know that I am the LORD."
EZEK|12|17|And the word of the LORD came to me:
EZEK|12|18|"Son of man, eat your bread with quaking, and drink water with trembling and with anxiety.
EZEK|12|19|And say to the people of the land, Thus says the Lord GOD concerning the inhabitants of Jerusalem in the land of Israel: They shall eat their bread with anxiety, and drink water in dismay. In this way her land will be stripped of all it contains, on account of the violence of all those who dwell in it.
EZEK|12|20|And the inhabited cities shall be laid waste, and the land shall become a desolation; and you shall know that I am the LORD."
EZEK|12|21|And the word of the LORD came to me:
EZEK|12|22|"Son of man, what is this proverb that you have about the land of Israel, saying, 'The days grow long, and every vision comes to nothing'?
EZEK|12|23|Tell them therefore, 'Thus says the Lord GOD: I will put an end to this proverb, and they shall no more use it as a proverb in Israel.' But say to them, The days are near, and the fulfillment of every vision.
EZEK|12|24|For there shall be no more any false vision or flattering divination within the house of Israel.
EZEK|12|25|For I am the LORD; I will speak the word that I will speak, and it will be performed. It will no longer be delayed, but in your days, O rebellious house, I will speak the word and perform it, declares the Lord GOD."
EZEK|12|26|And the word of the LORD came to me:
EZEK|12|27|"Son of man, behold, they of the house of Israel say, 'The vision that he sees is for many days from now, and he prophesies of times far off.'
EZEK|12|28|Therefore say to them, Thus says the Lord GOD: None of my words will be delayed any longer, but the word that I speak will be performed, declares the Lord GOD."
EZEK|13|1|The word of the LORD came to me:
EZEK|13|2|"Son of man, prophesy against the prophets of Israel, who are prophesying, and say to those who prophesy from their own hearts: 'Hear the word of the LORD!'
EZEK|13|3|Thus says the Lord GOD, Woe to the foolish prophets who follow their own spirit, and have seen nothing!
EZEK|13|4|Your prophets have been like jackals among ruins, O Israel.
EZEK|13|5|You have not gone up into the breaches, or built up a wall for the house of Israel, that it might stand in battle in the day of the LORD.
EZEK|13|6|They have seen false visions and lying divinations. They say, 'Declares the LORD,' when the LORD has not sent them, and yet they expect him to fulfill their word.
EZEK|13|7|Have you not seen a false vision and uttered a lying divination, whenever you have said, 'Declares the LORD,' although I have not spoken?"
EZEK|13|8|Therefore thus says the Lord GOD: "Because you have uttered falsehood and seen lying visions, therefore behold, I am against you, declares the Lord GOD.
EZEK|13|9|My hand will be against the prophets who see false visions and who give lying divinations. They shall not be in the council of my people, nor be enrolled in the register of the house of Israel, nor shall they enter the land of Israel. And you shall know that I am the Lord GOD.
EZEK|13|10|Precisely because they have misled my people, saying, 'Peace,' when there is no peace, and because, when the people build a wall, these prophets smear it with whitewash,
EZEK|13|11|say to those who smear it with whitewash that it shall fall! There will be a deluge of rain, and you, O great hailstones, will fall, and a stormy wind break out.
EZEK|13|12|And when the wall falls, will it not be said to you, 'Where is the coating with which you smeared it?'
EZEK|13|13|Therefore thus says the Lord GOD: I will make a stormy wind break out in my wrath, and there shall be a deluge of rain in my anger, and great hailstones in wrath to make a full end.
EZEK|13|14|And I will break down the wall that you have smeared with whitewash, and bring it down to the ground, so that its foundation will be laid bare. When it falls, you shall perish in the midst of it, and you shall know that I am the LORD.
EZEK|13|15|Thus will I spend my wrath upon the wall and upon those who have smeared it with whitewash, and I will say to you, The wall is no more, nor those who smeared it,
EZEK|13|16|the prophets of Israel who prophesied concerning Jerusalem and saw visions of peace for her, when there was no peace, declares the Lord GOD.
EZEK|13|17|"And you, son of man, set your face against the daughters of your people, who prophesy out of their own minds. Prophesy against them
EZEK|13|18|and say, Thus says the Lord GOD: Woe to the women who sew magic bands upon all wrists, and make veils for the heads of persons of every stature, in the hunt for souls! Will you hunt down souls belonging to my people and keep your own souls alive?
EZEK|13|19|You have profaned me among my people for handfuls of barley and for pieces of bread, putting to death souls who should not die and keeping alive souls who should not live, by your lying to my people, who listen to lies.
EZEK|13|20|"Therefore thus says the Lord GOD: Behold, I am against your magic bands with which you hunt the souls like birds, and I will tear them from your arms, and I will let the souls whom you hunt go free, the souls like birds.
EZEK|13|21|Your veils also I will tear off and deliver my people out of your hand, and they shall be no more in your hand as prey, and you shall know that I am the LORD.
EZEK|13|22|Because you have disheartened the righteous falsely, although I have not grieved him, and you have encouraged the wicked, that he should not turn from his evil way to save his life,
EZEK|13|23|therefore you shall no more see false visions nor practice divination. I will deliver my people out of your hand. And you shall know that I am the LORD."
EZEK|14|1|Then certain of the elders of Israel came to me and sat before me.
EZEK|14|2|And the word of the LORD came to me:
EZEK|14|3|"Son of man, these men have taken their idols into their hearts, and set the stumbling block of their iniquity before their faces. Should I indeed let myself be consulted by them?
EZEK|14|4|Therefore speak to them and say to them, Thus says the Lord GOD: Any one of the house of Israel who takes his idols into his heart and sets the stumbling block of his iniquity before his face, and yet comes to the prophet, I the LORD will answer him as he comes with the multitude of his idols,
EZEK|14|5|that I may lay hold of the hearts of the house of Israel, who are all estranged from me through their idols.
EZEK|14|6|"Therefore say to the house of Israel, Thus says the Lord GOD: Repent and turn away from your idols, and turn away your faces from all your abominations.
EZEK|14|7|For any one of the house of Israel, or of the strangers who sojourn in Israel, who separates himself from me, taking his idols into his heart and putting the stumbling block of his iniquity before his face, and yet comes to a prophet to consult me through him, I the LORD will answer him myself.
EZEK|14|8|And I will set my face against that man; I will make him a sign and a byword and cut him off from the midst of my people, and you shall know that I am the LORD.
EZEK|14|9|And if the prophet is deceived and speaks a word, I, the LORD, have deceived that prophet, and I will stretch out my hand against him and will destroy him from the midst of my people Israel.
EZEK|14|10|And they shall bear their punishment- the punishment of the prophet and the punishment of the inquirer shall be alike-
EZEK|14|11|that the house of Israel may no more go astray from me, nor defile themselves anymore with all their transgressions, but that they may be my people and I may be their God, declares the Lord GOD."
EZEK|14|12|And the word of the LORD came to me:
EZEK|14|13|"Son of man, when a land sins against me by acting faithlessly, and I stretch out my hand against it and break its supply of bread and send famine upon it, and cut off from it man and beast,
EZEK|14|14|even if these three men, Noah, Daniel, and Job, were in it, they would deliver but their own lives by their righteousness, declares the Lord GOD.
EZEK|14|15|"If I cause wild beasts to pass through the land, and they ravage it, and it be made desolate, so that no one may pass through because of the beasts,
EZEK|14|16|even if these three men were in it, as I live, declares the Lord GOD, they would deliver neither sons nor daughters. They alone would be delivered, but the land would be desolate.
EZEK|14|17|"Or if I bring a sword upon that land and say, Let a sword pass through the land, and I cut off from it man and beast,
EZEK|14|18|though these three men were in it, as I live, declares the Lord GOD, they would deliver neither sons nor daughters, but they alone would be delivered.
EZEK|14|19|"Or if I send a pestilence into that land and pour out my wrath upon it with blood, to cut off from it man and beast,
EZEK|14|20|even if Noah, Daniel, and Job were in it, as I live, declares the Lord GOD, they would deliver neither son nor daughter. They would deliver but their own lives by their righteousness.
EZEK|14|21|"For thus says the Lord GOD: How much more when I send upon Jerusalem my four disastrous acts of judgment, sword, famine, wild beasts, and pestilence, to cut off from it man and beast!
EZEK|14|22|But behold, some survivors will be left in it, sons and daughters who will be brought out; behold, when they come out to you, and you see their ways and their deeds, you will be consoled for the disaster that I have brought upon Jerusalem, for all that I have brought upon it.
EZEK|14|23|They will console you, when you see their ways and their deeds, and you shall know that I have not done without cause all that I have done in it, declares the Lord GOD."
EZEK|15|1|And the word of the LORD came to me:
EZEK|15|2|"Son of man, how does the wood of the vine surpass any wood, the vine branch that is among the trees of the forest?
EZEK|15|3|Is wood taken from it to make anything? Do people take a peg from it to hang any vessel on it?
EZEK|15|4|Behold, it is given to the fire for fuel. When the fire has consumed both ends of it, and the middle of it is charred, is it useful for anything?
EZEK|15|5|Behold, when it was whole, it was used for nothing. How much less, when the fire has consumed it and it is charred, can it ever be used for anything!
EZEK|15|6|Therefore thus says the Lord GOD: Like the wood of the vine among the trees of the forest, which I have given to the fire for fuel, so have I given up the inhabitants of Jerusalem.
EZEK|15|7|And I will set my face against them. Though they escape from the fire, the fire shall yet consume them, and you will know that I am the LORD, when I set my face against them.
EZEK|15|8|And I will make the land desolate, because they have acted faithlessly, declares the Lord GOD."
EZEK|16|1|Again the word of the LORD came to me:
EZEK|16|2|"Son of man, make known to Jerusalem her abominations,
EZEK|16|3|and say, Thus says the Lord GOD to Jerusalem: Your origin and your birth are of the land of the Canaanites; your father was an Amorite and your mother a Hittite.
EZEK|16|4|And as for your birth, on the day you were born your cord was not cut, nor were you washed with water to cleanse you, nor rubbed with salt, nor wrapped in swaddling cloths.
EZEK|16|5|No eye pitied you, to do any of these things to you out of compassion for you, but you were cast out on the open field, for you were abhorred, on the day that you were born.
EZEK|16|6|"And when I passed by you and saw you wallowing in your blood, I said to you in your blood, 'Live!' I said to you in your blood, 'Live!'
EZEK|16|7|I made you flourish like a plant of the field. And you grew up and became tall and arrived at full adornment. Your breasts were formed, and your hair had grown; yet you were naked and bare.
EZEK|16|8|"When I passed by you again and saw you, behold, you were at the age for love, and I spread the corner of my garment over you and covered your nakedness; I made my vow to you and entered into a covenant with you, declares the Lord GOD, and you became mine.
EZEK|16|9|Then I bathed you with water and washed off your blood from you and anointed you with oil.
EZEK|16|10|I clothed you also with embroidered cloth and shod you with fine leather. I wrapped you in fine linen and covered you with silk.
EZEK|16|11|And I adorned you with ornaments and put bracelets on your wrists and a chain on your neck.
EZEK|16|12|And I put a ring on your nose and earrings in your ears and a beautiful crown on your head.
EZEK|16|13|Thus you were adorned with gold and silver, and your clothing was of fine linen and silk and embroidered cloth. You ate fine flour and honey and oil. You grew exceedingly beautiful and advanced to royalty.
EZEK|16|14|And your renown went forth among the nations because of your beauty, for it was perfect through the splendor that I had bestowed on you, declares the Lord GOD.
EZEK|16|15|"But you trusted in your beauty and played the whore because of your renown and lavished your whorings on any passerby; your beauty became his.
EZEK|16|16|You took some of your garments and made for yourself colorful shrines, and on them played the whore. The like has never been, nor ever shall be.
EZEK|16|17|You also took your beautiful jewels of my gold and of my silver, which I had given you, and made for yourself images of men, and with them played the whore.
EZEK|16|18|And you took your embroidered garments to cover them, and set my oil and my incense before them.
EZEK|16|19|Also my bread that I gave you- I fed you with fine flour and oil and honey- you set before them for a pleasing aroma; and so it was, declares the Lord GOD.
EZEK|16|20|And you took your sons and your daughters, whom you had borne to me, and these you sacrificed to them to be devoured. Were your whorings so small a matter
EZEK|16|21|that you slaughtered my children and delivered them up as an offering by fire to them?
EZEK|16|22|And in all your abominations and your whorings you did not remember the days of your youth, when you were naked and bare, wallowing in your blood.
EZEK|16|23|"And after all your wickedness (woe, woe to you! declares the Lord GOD),
EZEK|16|24|you built yourself a vaulted chamber and made yourself a lofty place in every square.
EZEK|16|25|At the head of every street you built your lofty place and made your beauty an abomination, offering yourself to any passerby and multiplying your whoring.
EZEK|16|26|You also played the whore with the Egyptians, your lustful neighbors, multiplying your whoring, to provoke me to anger.
EZEK|16|27|Behold, therefore, I stretched out my hand against you and diminished your allotted portion and delivered you to the greed of your enemies, the daughters of the Philistines, who were ashamed of your lewd behavior.
EZEK|16|28|You played the whore also with the Assyrians, because you were not satisfied; yes, you played the whore with them, and still you were not satisfied.
EZEK|16|29|You multiplied your whoring also with the trading land of Chaldea, and even with this you were not satisfied.
EZEK|16|30|"How lovesick is your heart, declares the Lord GOD, because you did all these things, the deeds of a brazen prostitute,
EZEK|16|31|building your vaulted chamber at the head of every street, and making your lofty place in every square. Yet you were not like a prostitute, because you scorned payment.
EZEK|16|32|Adulterous wife, who receives strangers instead of her husband!
EZEK|16|33|Men give gifts to all prostitutes, but you gave your gifts to all your lovers, bribing them to come to you from every side with your whorings.
EZEK|16|34|So you were different from other women in your whorings. No one solicited you to play the whore, and you gave payment, while no payment was given to you; therefore you were different.
EZEK|16|35|"Therefore, O prostitute, hear the word of the LORD:
EZEK|16|36|Thus says the Lord GOD, Because your lust was poured out and your nakedness uncovered in your whorings with your lovers, and with all your abominable idols, and because of the blood of your children that you gave to them,
EZEK|16|37|therefore, behold, I will gather all your lovers with whom you took pleasure, all those you loved and all those you hated. I will gather them against you from every side and will uncover your nakedness to them, that they may see all your nakedness.
EZEK|16|38|And I will judge you as women who commit adultery and shed blood are judged, and bring upon you the blood of wrath and jealousy.
EZEK|16|39|And I will give you into their hands, and they shall throw down your vaulted chamber and break down your lofty places. They shall strip you of your clothes and take your beautiful jewels and leave you naked and bare.
EZEK|16|40|They shall bring up a crowd against you, and they shall stone you and cut you to pieces with their swords.
EZEK|16|41|And they shall burn your houses and execute judgments upon you in the sight of many women. I will make you stop playing the whore, and you shall also give payment no more.
EZEK|16|42|So will I satisfy my wrath on you, and my jealousy shall depart from you. I will be calm and will no more be angry.
EZEK|16|43|Because you have not remembered the days of your youth, but have enraged me with all these things, therefore, behold, I have returned your deeds upon your head, declares the Lord GOD. "Have you not committed lewdness in addition to all your abominations?
EZEK|16|44|"Behold, everyone who uses proverbs will use this proverb about you: 'Like mother, like daughter.'
EZEK|16|45|You are the daughter of your mother, who loathed her husband and her children; and you are the sister of your sisters, who loathed their husbands and their children. Your mother was a Hittite and your father an Amorite.
EZEK|16|46|And your elder sister is Samaria, who lived with her daughters to the north of you; and your younger sister, who lived to the south of you, is Sodom with her daughters.
EZEK|16|47|Not only did you walk in their ways and do according to their abominations; within a very little time you were more corrupt than they in all your ways.
EZEK|16|48|As I live, declares the Lord GOD, your sister Sodom and her daughters have not done as you and your daughters have done.
EZEK|16|49|Behold, this was the guilt of your sister Sodom: she and her daughters had pride, excess of food, and prosperous ease, but did not aid the poor and needy.
EZEK|16|50|They were haughty and did an abomination before me. So I removed them, when I saw it.
EZEK|16|51|Samaria has not committed half your sins. You have committed more abominations than they, and have made your sisters appear righteous by all the abominations that you have committed.
EZEK|16|52|Bear your disgrace, you also, for you have intervened on behalf of your sisters. Because of your sins in which you acted more abominably than they, they are more in the right than you. So be ashamed, you also, and bear your disgrace, for you have made your sisters appear righteous.
EZEK|16|53|"I will restore their fortunes, both the fortunes of Sodom and her daughters, and the fortunes of Samaria and her daughters, and I will restore your own fortunes in their midst,
EZEK|16|54|that you may bear your disgrace and be ashamed of all that you have done, becoming a consolation to them.
EZEK|16|55|As for your sisters, Sodom and her daughters shall return to their former state, and Samaria and her daughters shall return to their former state, and you and your daughters shall return to your former state.
EZEK|16|56|Was not your sister Sodom a byword in your mouth in the day of your pride,
EZEK|16|57|before your wickedness was uncovered? Now you have become an object of reproach for the daughters of Syria and all those around her, and for the daughters of the Philistines, those all around who despise you.
EZEK|16|58|You bear the penalty of your lewdness and your abominations, declares the LORD.
EZEK|16|59|"For thus says the Lord GOD: I will deal with you as you have done, you who have despised the oath in breaking the covenant,
EZEK|16|60|yet I will remember my covenant with you in the days of your youth, and I will establish for you an everlasting covenant.
EZEK|16|61|Then you will remember your ways and be ashamed when you take your sisters, both your elder and your younger, and I give them to you as daughters, but not on account of the covenant with you.
EZEK|16|62|I will establish my covenant with you, and you shall know that I am the LORD,
EZEK|16|63|that you may remember and be confounded, and never open your mouth again because of your shame, when I atone for you for all that you have done, declares the Lord GOD."
EZEK|17|1|The word of the LORD came to me:
EZEK|17|2|"Son of man, propound a riddle, and speak a parable to the house of Israel;
EZEK|17|3|say, Thus says the Lord GOD: A great eagle with great wings and long pinions, rich in plumage of many colors, came to Lebanon and took the top of the cedar.
EZEK|17|4|He broke off the topmost of its young twigs and carried it to a land of trade and set it in a city of merchants.
EZEK|17|5|Then he took of the seed of the land and planted it in fertile soil. He placed it beside abundant waters. He set it like a willow twig,
EZEK|17|6|and it sprouted and became a low spreading vine, and its branches turned toward him, and its roots remained where it stood. So it became a vine and produced branches and put out boughs.
EZEK|17|7|"And there was another great eagle with great wings and much plumage, and behold, this vine bent its roots toward him and shot forth its branches toward him from the bed where it was planted, that he might water it.
EZEK|17|8|It had been planted on good soil by abundant waters, that it might produce branches and bear fruit and become a noble vine.
EZEK|17|9|"Say, Thus says the Lord GOD: Will it thrive? Will he not pull up its roots and cut off its fruit, so that it withers, so that all its fresh sprouting leaves wither? It will not take a strong arm or many people to pull it from its roots.
EZEK|17|10|Behold, it is planted; will it thrive? Will it not utterly wither when the east wind strikes it- wither away on the bed where it sprouted?"
EZEK|17|11|Then the word of the LORD came to me:
EZEK|17|12|"Say now to the rebellious house, Do you not know what these things mean? Tell them, behold, the king of Babylon came to Jerusalem, and took her king and her princes and brought them to him to Babylon.
EZEK|17|13|And he took one of the royal offspring and made a covenant with him, putting him under oath (the chief men of the land he had taken away),
EZEK|17|14|that the kingdom might be humble and not lift itself up, and keep his covenant that it might stand.
EZEK|17|15|But he rebelled against him by sending his ambassadors to Egypt, that they might give him horses and a large army. Will he thrive? Can one escape who does such things? Can he break the covenant and yet escape?
EZEK|17|16|"As I live, declares the Lord GOD, surely in the place where the king dwells who made him king, whose oath he despised, and whose covenant with him he broke, in Babylon he shall die.
EZEK|17|17|Pharaoh with his mighty army and great company will not help him in war, when mounds are cast up and siege walls built to cut off many lives.
EZEK|17|18|He despised the oath in breaking the covenant, and behold, he gave his hand and did all these things; he shall not escape.
EZEK|17|19|Therefore thus says the Lord GOD: As I live, surely it is my oath that he despised, and my covenant that he broke. I will return it upon his head.
EZEK|17|20|I will spread my net over him, and he shall be taken in my snare, and I will bring him to Babylon and enter into judgment with him there for the treachery he has committed against me.
EZEK|17|21|And all the pick of his troops shall fall by the sword, and the survivors shall be scattered to every wind, and you shall know that I am the LORD; I have spoken."
EZEK|17|22|Thus says the Lord GOD: "I myself will take a sprig from the lofty top of the cedar and will set it out. I will break off from the topmost of its young twigs a tender one, and I myself will plant it on a high and lofty mountain.
EZEK|17|23|On the mountain height of Israel will I plant it, that it may bear branches and produce fruit and become a noble cedar. And under it will dwell every kind of bird; in the shade of its branches birds of every sort will nest.
EZEK|17|24|And all the trees of the field shall know that I am the LORD; I bring low the high tree, and make high the low tree, dry up the green tree, and make the dry tree flourish. I am the LORD; I have spoken, and I will do it."
EZEK|18|1|The word of the LORD came to me:
EZEK|18|2|"What do you mean by repeating this proverb concerning the land of Israel, 'The fathers have eaten sour grapes, and the children's teeth are set on edge'?
EZEK|18|3|As I live, declares the Lord GOD, this proverb shall no more be used by you in Israel.
EZEK|18|4|Behold, all souls are mine; the soul of the father as well as the soul of the son is mine: the soul who sins shall die.
EZEK|18|5|"If a man is righteous and does what is just and right-
EZEK|18|6|if he does not eat upon the mountains or lift up his eyes to the idols of the house of Israel, does not defile his neighbor's wife or approach a woman in her time of menstrual impurity,
EZEK|18|7|does not oppress anyone, but restores to the debtor his pledge, commits no robbery, gives his bread to the hungry and covers the naked with a garment,
EZEK|18|8|does not lend at interest or take any profit, withholds his hand from injustice, executes true justice between man and man,
EZEK|18|9|walks in my statutes, and keeps my rules by acting faithfully- he is righteous; he shall surely live, declares the Lord GOD.
EZEK|18|10|"If he fathers a son who is violent, a shedder of blood, who does any of these things
EZEK|18|11|(though he himself did none of these things), who even eats upon the mountains, defiles his neighbor's wife,
EZEK|18|12|oppresses the poor and needy, commits robbery, does not restore the pledge, lifts up his eyes to the idols, commits abomination,
EZEK|18|13|lends at interest, and takes profit; shall he then live? He shall not live. He has done all these abominations; he shall surely die; his blood shall be upon himself.
EZEK|18|14|"Now suppose this man fathers a son who sees all the sins that his father has done; he sees, and does not do likewise:
EZEK|18|15|he does not eat upon the mountains or lift up his eyes to the idols of the house of Israel, does not defile his neighbor's wife,
EZEK|18|16|does not oppress anyone, exacts no pledge, commits no robbery, but gives his bread to the hungry and covers the naked with a garment,
EZEK|18|17|withholds his hand from iniquity, takes no interest or profit, obeys my rules, and walks in my statutes; he shall not die for his father's iniquity; he shall surely live.
EZEK|18|18|As for his father, because he practiced extortion, robbed his brother, and did what is not good among his people, behold, he shall die for his iniquity.
EZEK|18|19|"Yet you say, 'Why should not the son suffer for the iniquity of the father?' When the son has done what is just and right, and has been careful to observe all my statutes, he shall surely live.
EZEK|18|20|The soul who sins shall die. The son shall not suffer for the iniquity of the father, nor the father suffer for the iniquity of the son. The righteousness of the righteous shall be upon himself, and the wickedness of the wicked shall be upon himself.
EZEK|18|21|"But if a wicked person turns away from all his sins that he has committed and keeps all my statutes and does what is just and right, he shall surely live; he shall not die.
EZEK|18|22|None of the transgressions that he has committed shall be remembered against him; for the righteousness that he has done he shall live.
EZEK|18|23|Have I any pleasure in the death of the wicked, declares the Lord GOD, and not rather that he should turn from his way and live?
EZEK|18|24|But when a righteous person turns away from his righteousness and does injustice and does the same abominations that the wicked person does, shall he live? None of the righteous deeds that he has done shall be remembered; for the treachery of which he is guilty and the sin he has committed, for them he shall die.
EZEK|18|25|"Yet you say, 'The way of the Lord is not just.' Hear now, O house of Israel: Is my way not just? Is it not your ways that are not just?
EZEK|18|26|When a righteous person turns away from his righteousness and does injustice, he shall die for it; for the injustice that he has done he shall die.
EZEK|18|27|Again, when a wicked person turns away from the wickedness he has committed and does what is just and right, he shall save his life.
EZEK|18|28|Because he considered and turned away from all the transgressions that he had committed, he shall surely live; he shall not die.
EZEK|18|29|Yet the house of Israel says, 'The way of the Lord is not just.' O house of Israel, are my ways not just? Is it not your ways that are not just?
EZEK|18|30|"Therefore I will judge you, O house of Israel, every one according to his ways, declares the Lord GOD. Repent and turn from all your transgressions, lest iniquity be your ruin.
EZEK|18|31|Cast away from you all the transgressions that you have committed, and make yourselves a new heart and a new spirit! Why will you die, O house of Israel?
EZEK|18|32|For I have no pleasure in the death of anyone, declares the Lord GOD; so turn, and live."
EZEK|19|1|And you, take up a lamentation for the princes of Israel,
EZEK|19|2|and say: What was your mother? A lioness! Among lions she crouched; in the midst of young lions she reared her cubs.
EZEK|19|3|And she brought up one of her cubs; he became a young lion, and he learned to catch prey; he devoured men.
EZEK|19|4|The nations heard about him; he was caught in their pit, and they brought him with hooks to the land of Egypt.
EZEK|19|5|When she saw that she waited in vain, that her hope was lost, she took another of her cubs and made him a young lion.
EZEK|19|6|He prowled among the lions; he became a young lion, and he learned to catch prey; he devoured men,
EZEK|19|7|and seized their widows. He laid waste their cities, and the land was appalled and all who were in it at the sound of his roaring.
EZEK|19|8|Then the nations set against him from provinces on every side; they spread their net over him; he was taken in their pit.
EZEK|19|9|With hooks they put him in a cage and brought him to the king of Babylon; they brought him into custody, that his voice should no more be heard on the mountains of Israel.
EZEK|19|10|Your mother was like a vine in a vineyard planted by the water, fruitful and full of branches by reason of abundant water.
EZEK|19|11|Its strong stems became rulers' scepters; it towered aloft among the thick boughs; it was seen in its height with the mass of its branches.
EZEK|19|12|But the vine was plucked up in fury, cast down to the ground; the east wind dried up its fruit; they were stripped off and withered. As for its strong stem, fire consumed it.
EZEK|19|13|Now it is planted in the wilderness, in a dry and thirsty land.
EZEK|19|14|And fire has gone out from the stem of its shoots, has consumed its fruit, so that there remains in it no strong stem, no scepter for ruling. This is a lamentation and has become a lamentation.
EZEK|20|1|In the seventh year, in the fifth month, on the tenth day of the month, certain of the elders of Israel came to inquire of the LORD, and sat before me.
EZEK|20|2|And the word of the LORD came to me:
EZEK|20|3|"Son of man, speak to the elders of Israel, and say to them, Thus says the Lord GOD, Is it to inquire of me that you come? As I live, declares the Lord GOD, I will not be inquired of by you.
EZEK|20|4|Will you judge them, son of man, will you judge them? Let them know the abominations of their fathers,
EZEK|20|5|and say to them, Thus says the Lord GOD: On the day when I chose Israel, I swore to the offspring of the house of Jacob, making myself known to them in the land of Egypt; I swore to them, saying, I am the LORD your God.
EZEK|20|6|On that day I swore to them that I would bring them out of the land of Egypt into a land that I had searched out for them, a land flowing with milk and honey, the most glorious of all lands.
EZEK|20|7|And I said to them, Cast away the detestable things your eyes feast on, every one of you, and do not defile yourselves with the idols of Egypt; I am the LORD your God.
EZEK|20|8|But they rebelled against me and were not willing to listen to me. None of them cast away the detestable things their eyes feasted on, nor did they forsake the idols of Egypt. "Then I said I would pour out my wrath upon them and spend my anger against them in the midst of the land of Egypt.
EZEK|20|9|But I acted for the sake of my name, that it should not be profaned in the sight of the nations among whom they lived, in whose sight I made myself known to them in bringing them out of the land of Egypt.
EZEK|20|10|So I led them out of the land of Egypt and brought them into the wilderness.
EZEK|20|11|I gave them my statutes and made known to them my rules, by which, if a person does them, he shall live.
EZEK|20|12|Moreover, I gave them my Sabbaths, as a sign between me and them, that they might know that I am the LORD who sanctifies them.
EZEK|20|13|But the house of Israel rebelled against me in the wilderness. They did not walk in my statutes but rejected my rules, by which, if a person does them, he shall live; and my Sabbaths they greatly profaned. "Then I said I would pour out my wrath upon them in the wilderness, to make a full end of them.
EZEK|20|14|But I acted for the sake of my name, that it should not be profaned in the sight of the nations, in whose sight I had brought them out.
EZEK|20|15|Moreover, I swore to them in the wilderness that I would not bring them into the land that I had given them, a land flowing with milk and honey, the most glorious of all lands,
EZEK|20|16|because they rejected my rules and did not walk in my statutes, and profaned my Sabbaths; for their heart went after their idols.
EZEK|20|17|Nevertheless, my eye spared them, and I did not destroy them or make a full end of them in the wilderness.
EZEK|20|18|"And I said to their children in the wilderness, Do not walk in the statutes of your fathers, nor keep their rules, nor defile yourselves with their idols.
EZEK|20|19|I am the LORD your God; walk in my statutes, and be careful to obey my rules,
EZEK|20|20|and keep my Sabbaths holy that they may be a sign between me and you, that you may know that I am the LORD your God.
EZEK|20|21|But the children rebelled against me. They did not walk in my statutes and were not careful to obey my rules, by which, if a person does them, he shall live; they profaned my Sabbaths. "Then I said I would pour out my wrath upon them and spend my anger against them in the wilderness.
EZEK|20|22|But I withheld my hand and acted for the sake of my name, that it should not be profaned in the sight of the nations, in whose sight I had brought them out.
EZEK|20|23|Moreover, I swore to them in the wilderness that I would scatter them among the nations and disperse them through the countries,
EZEK|20|24|because they had not obeyed my rules, but had rejected my statutes and profaned my Sabbaths, and their eyes were set on their fathers' idols.
EZEK|20|25|Moreover, I gave them statutes that were not good and rules by which they could not have life,
EZEK|20|26|and I defiled them through their very gifts in their offering up all their firstborn, that I might devastate them. I did it that they might know that I am the LORD.
EZEK|20|27|"Therefore, son of man, speak to the house of Israel and say to them, Thus says the Lord GOD: In this also your fathers blasphemed me, by dealing treacherously with me.
EZEK|20|28|For when I had brought them into the land that I swore to give them, then wherever they saw any high hill or any leafy tree, there they offered their sacrifices and there they presented the provocation of their offering; there they sent up their pleasing aromas, and there they poured out their drink offerings.
EZEK|20|29|(I said to them, What is the high place to which you go? So its name is called Bamah to this day.)
EZEK|20|30|"Therefore say to the house of Israel, Thus says the Lord GOD: Will you defile yourselves after the manner of your fathers and go whoring after their detestable things?
EZEK|20|31|When you present your gifts and offer up your children in fire, you defile yourselves with all your idols to this day. And shall I be inquired of by you, O house of Israel? As I live, declares the Lord GOD, I will not be inquired of by you.
EZEK|20|32|"What is in your mind shall never happen- the thought, 'Let us be like the nations, like the tribes of the countries, and worship wood and stone.'
EZEK|20|33|"As I live, declares the Lord GOD, surely with a mighty hand and an outstretched arm and with wrath poured out I will be king over you.
EZEK|20|34|I will bring you out from the peoples and gather you out of the countries where you are scattered, with a mighty hand and an outstretched arm, and with wrath poured out.
EZEK|20|35|And I will bring you into the wilderness of the peoples, and there I will enter into judgment with you face to face.
EZEK|20|36|As I entered into judgment with your fathers in the wilderness of the land of Egypt, so I will enter into judgment with you, declares the Lord GOD.
EZEK|20|37|I will make you pass under the rod, and I will bring you into the bond of the covenant.
EZEK|20|38|I will purge out the rebels from among you, and those who transgress against me. I will bring them out of the land where they sojourn, but they shall not enter the land of Israel. Then you will know that I am the LORD.
EZEK|20|39|"As for you, O house of Israel, thus says the Lord GOD: Go serve every one of you his idols, now and hereafter, if you will not listen to me; but my holy name you shall no more profane with your gifts and your idols.
EZEK|20|40|"For on my holy mountain, the mountain height of Israel, declares the Lord GOD, there all the house of Israel, all of them, shall serve me in the land. There I will accept them, and there I will require your contributions and the choicest of your gifts, with all your sacred offerings.
EZEK|20|41|As a pleasing aroma I will accept you, when I bring you out from the peoples and gather you out of the countries where you have been scattered. And I will manifest my holiness among you in the sight of the nations.
EZEK|20|42|And you shall know that I am the LORD, when I bring you into the land of Israel, the country that I swore to give to your fathers.
EZEK|20|43|And there you shall remember your ways and all your deeds with which you have defiled yourselves, and you shall loathe yourselves for all the evils that you have committed.
EZEK|20|44|And you shall know that I am the LORD, when I deal with you for my name's sake, not according to your evil ways, nor according to your corrupt deeds, O house of Israel, declares the Lord GOD."
EZEK|20|45|And the word of the LORD came to me:
EZEK|20|46|"Son of man, set your face toward the southland; preach against the south, and prophesy against the forest land in the Negeb.
EZEK|20|47|Say to the forest of the Negeb, Hear the word of the LORD: Thus says the Lord GOD, Behold, I will kindle a fire in you, and it shall devour every green tree in you and every dry tree. The blazing flame shall not be quenched, and all faces from south to north shall be scorched by it.
EZEK|20|48|All flesh shall see that I the LORD have kindled it; it shall not be quenched."
EZEK|20|49|Then I said, "Ah, Lord GOD! They are saying of me, 'Is he not a maker of parables?'"
EZEK|21|1|The word of the LORD came to me:
EZEK|21|2|"Son of man, set your face toward Jerusalem and preach against the sanctuaries. Prophesy against the land of Israel
EZEK|21|3|and say to the land of Israel, Thus says the LORD: Behold, I am against you and will draw my sword from its sheath and will cut off from you both righteous and wicked.
EZEK|21|4|Because I will cut off from you both righteous and wicked, therefore my sword shall be drawn from its sheath against all flesh from south to north.
EZEK|21|5|And all flesh shall know that I am the LORD. I have drawn my sword from its sheath; it shall not be sheathed again.
EZEK|21|6|"As for you, son of man, groan; with breaking heart and bitter grief, groan before their eyes.
EZEK|21|7|And when they say to you, 'Why do you groan?' you shall say, 'Because of the news that it is coming. Every heart will melt, and all hands will be feeble; every spirit will faint, and all knees will be weak as water. Behold, it is coming, and it will be fulfilled,'"declares the Lord GOD.
EZEK|21|8|And the word of the LORD came to me:
EZEK|21|9|"Son of man, prophesy and say, Thus says the Lord; Say: "A sword, a sword is sharpened and also polished,
EZEK|21|10|sharpened for slaughter, polished to flash like lightning! (Or shall we rejoice? You have despised the rod, my son, with everything of wood.)
EZEK|21|11|So the sword is given to be polished, that it may be grasped in the hand. It is sharpened and polished to be given into the hand of the slayer.
EZEK|21|12|Cry out and wail, son of man, for it is against my people. It is against all the princes of Israel. They are delivered over to the sword with my people. Strike therefore upon your thigh.
EZEK|21|13|For it will not be a testing- what could it do if you despise the rod?" declares the Lord GOD.
EZEK|21|14|"As for you, son of man, prophesy. Clap your hands and let the sword come down twice, yes, three times, the sword for those to be slain. It is the sword for the great slaughter, which surrounds them,
EZEK|21|15|that their hearts may melt, and many stumble. At all their gates I have given the glittering sword. Ah, it is made like lightning; it is taken up for slaughter.
EZEK|21|16|Cut sharply to the right; set yourself to the left, wherever your face is directed.
EZEK|21|17|I also will clap my hands, and I will satisfy my fury; I the LORD have spoken."
EZEK|21|18|The word of the LORD came to me again:
EZEK|21|19|"As for you, son of man, mark two ways for the sword of the king of Babylon to come. Both of them shall come from the same land. And make a signpost; make it at the head of the way to a city.
EZEK|21|20|Mark a way for the sword to come to Rabbah of the Ammonites and to Judah, into Jerusalem the fortified.
EZEK|21|21|For the king of Babylon stands at the parting of the way, at the head of the two ways, to use divination. He shakes the arrows; he consults the teraphim; he looks at the liver.
EZEK|21|22|Into his right hand comes the divination for Jerusalem, to set battering rams, to open the mouth with murder, to lift up the voice with shouting, to set battering rams against the gates, to cast up mounds, to build siege towers.
EZEK|21|23|But to them it will seem like a false divination. They have sworn solemn oaths, but he brings their guilt to remembrance, that they may be taken.
EZEK|21|24|"Therefore thus says the Lord GOD: Because you have made your guilt to be remembered, in that your transgressions are uncovered, so that in all your deeds your sins appear- because you have come to remembrance, you shall be taken in hand.
EZEK|21|25|And you, O profane wicked one, prince of Israel, whose day has come, the time of your final punishment,
EZEK|21|26|thus says the Lord GOD: Remove the turban and take off the crown. Things shall not remain as they are. Exalt that which is low, and bring low that which is exalted.
EZEK|21|27|A ruin, ruin, ruin I will make it. This also shall not be, until he comes, the one to whom judgment belongs, and I will give it to him.
EZEK|21|28|"And you, son of man, prophesy, and say, Thus says the Lord GOD concerning the Ammonites and concerning their reproach; say, A sword, a sword is drawn for the slaughter. It is polished to consume and to flash like lightning-
EZEK|21|29|while they see for you false visions, while they divine lies for you- to place you on the necks of the profane wicked, whose day has come, the time of their final punishment.
EZEK|21|30|Return it to its sheath. In the place where you were created, in the land of your origin, I will judge you.
EZEK|21|31|And I will pour out my indignation upon you; I will blow upon you with the fire of my wrath, and I will deliver you into the hands of brutish men, skillful to destroy.
EZEK|21|32|You shall be fuel for the fire. Your blood shall be in the midst of the land. You shall be no more remembered, for I the LORD have spoken."
EZEK|22|1|And the word of the LORD came to me, saying,
EZEK|22|2|"And you, son of man, will you judge, will you judge the bloody city? Then declare to her all her abominations.
EZEK|22|3|You shall say, Thus says the Lord GOD: A city that sheds blood in her midst, so that her time may come, and that makes idols to defile herself!
EZEK|22|4|You have become guilty by the blood that you have shed, and defiled by the idols that you have made, and you have brought your days near, the appointed time of your years has come. Therefore I have made you a reproach to the nations, and a mockery to all the countries.
EZEK|22|5|Those who are near and those who are far from you will mock you; your name is defiled; you are full of tumult.
EZEK|22|6|"Behold, the princes of Israel in you, every one according to his power, have been bent on shedding blood.
EZEK|22|7|Father and mother are treated with contempt in you; the sojourner suffers extortion in your midst; the fatherless and the widow are wronged in you.
EZEK|22|8|You have despised my holy things and profaned my Sabbaths.
EZEK|22|9|There are men in you who slander to shed blood, and people in you who eat on the mountains; they commit lewdness in your midst.
EZEK|22|10|In you men uncover their fathers' nakedness; in you they violate women who are unclean in their menstrual impurity.
EZEK|22|11|One commits abomination with his neighbor's wife; another lewdly defiles his daughter-in-law; another in you violates his sister, his father's daughter.
EZEK|22|12|In you they take bribes to shed blood; you take interest and profit and make gain of your neighbors by extortion; but me you have forgotten, declares the Lord GOD.
EZEK|22|13|"Behold, I strike my hand at the dishonest gain that you have made, and at the blood that has been in your midst.
EZEK|22|14|Can your courage endure, or can your hands be strong, in the days that I shall deal with you? I the LORD have spoken, and I will do it.
EZEK|22|15|I will scatter you among the nations and disperse you through the countries, and I will consume your uncleanness out of you.
EZEK|22|16|And you shall be profaned by your own doing in the sight of the nations, and you shall know that I am the LORD."
EZEK|22|17|And the word of the LORD came to me:
EZEK|22|18|"Son of man, the house of Israel has become dross to me; all of them are bronze and tin and iron and lead in the furnace; they are dross of silver.
EZEK|22|19|Therefore thus says the Lord GOD: Because you have all become dross, therefore, behold, I will gather you into the midst of Jerusalem.
EZEK|22|20|As one gathers silver and bronze and iron and lead and tin into a furnace, to blow the fire on it in order to melt it, so I will gather you in my anger and in my wrath, and I will put you in and melt you.
EZEK|22|21|I will gather you and blow on you with the fire of my wrath, and you shall be melted in the midst of it.
EZEK|22|22|As silver is melted in a furnace, so you shall be melted in the midst of it, and you shall know that I am the LORD; I have poured out my wrath upon you."
EZEK|22|23|And the word of the LORD came to me:
EZEK|22|24|"Son of man, say to her, You are a land that is not cleansed or rained upon in the day of indignation.
EZEK|22|25|The conspiracy of her prophets in her midst is like a roaring lion tearing the prey; they have devoured human lives; they have taken treasure and precious things; they have made many widows in her midst.
EZEK|22|26|Her priests have done violence to my law and have profaned my holy things. They have made no distinction between the holy and the common, neither have they taught the difference between the unclean and the clean, and they have disregarded my Sabbaths, so that I am profaned among them.
EZEK|22|27|Her princes in her midst are like wolves tearing the prey, shedding blood, destroying lives to get dishonest gain.
EZEK|22|28|And her prophets have smeared whitewash for them, seeing false visions and divining lies for them, saying, 'Thus says the Lord GOD,' when the LORD has not spoken.
EZEK|22|29|The people of the land have practiced extortion and committed robbery. They have oppressed the poor and needy, and have extorted from the sojourner without justice.
EZEK|22|30|And I sought for a man among them who should build up the wall and stand in the breach before me for the land, that I should not destroy it, but I found none.
EZEK|22|31|Therefore I have poured out my indignation upon them. I have consumed them with the fire of my wrath. I have returned their way upon their heads, declares the Lord GOD."
EZEK|23|1|The word of the LORD came to me:
EZEK|23|2|"Son of man, there were two women, the daughters of one mother.
EZEK|23|3|They played the whore in Egypt; they played the whore in their youth; there their breasts were pressed and their virgin bosoms handled.
EZEK|23|4|Oholah was the name of the elder and Oholibah the name of her sister. They became mine, and they bore sons and daughters. As for their names, Oholah is Samaria, and Oholibah is Jerusalem.
EZEK|23|5|"Oholah played the whore while she was mine, and she lusted after her lovers the Assyrians, warriors
EZEK|23|6|clothed in purple, governors and commanders, all of them desirable young men, horsemen riding on horses.
EZEK|23|7|She bestowed her whoring upon them, the choicest men of Assyria all of them, and she defiled herself with all the idols of everyone after whom she lusted.
EZEK|23|8|She did not give up her whoring that she had begun in Egypt; for in her youth men had lain with her and handled her virgin bosom and poured out their whoring lust upon her.
EZEK|23|9|Therefore I delivered her into the hands of her lovers, into the hands of the Assyrians, after whom she lusted.
EZEK|23|10|These uncovered her nakedness; they seized her sons and her daughters; and as for her, they killed her with the sword; and she became a byword among women, when judgment had been executed on her.
EZEK|23|11|"Her sister Oholibah saw this, and she became more corrupt than her sister in her lust and in her whoring, which was worse than that of her sister.
EZEK|23|12|She lusted after the Assyrians, governors and commanders, warriors clothed in full armor, horsemen riding on horses, all of them desirable young men.
EZEK|23|13|And I saw that she was defiled; they both took the same way.
EZEK|23|14|But she carried her whoring further. She saw men portrayed on the wall, the images of the Chaldeans portrayed in vermilion,
EZEK|23|15|wearing belts on their waists, with flowing turbans on their heads, all of them having the appearance of officers, a likeness of Bab ylonians whose native land was Chaldea.
EZEK|23|16|When she saw them, she lusted after them and sent messengers to them in Chaldea.
EZEK|23|17|And the Babylonians came to her into the bed of love, and they defiled her with their whoring lust. And after she was defiled by them, she turned from them in disgust.
EZEK|23|18|When she carried on her whoring so openly and flaunted her nakedness, I turned in disgust from her, as I had turned in disgust from her sister.
EZEK|23|19|Yet she increased her whoring, remembering the days of her youth, when she played the whore in the land of Egypt
EZEK|23|20|and lusted after her paramours there, whose members were like those of donkeys, and whose issue was like that of horses.
EZEK|23|21|Thus you longed for the lewdness of your youth, when the Egyptians handled your bosom and pressed your young breasts."
EZEK|23|22|Therefore, O Oholibah, thus says the Lord GOD: "Behold, I will stir up against you your lovers from whom you turned in disgust, and I will bring them against you from every side:
EZEK|23|23|the Babylonians and all the Chaldeans, Pekod and Shoa and Koa, and all the Assyrians with them, desirable young men, governors and commanders all of them, officers and men of renown, all of them riding on horses.
EZEK|23|24|And they shall come against you from the north with chariots and wagons and a host of peoples. They shall set themselves against you on every side with buckler, shield, and helmet; and I will commit the judgment to them, and they shall judge you according to their judgments.
EZEK|23|25|And I will direct my jealousy against you, that they may deal with you in fury. They shall cut off your nose and your ears, and your survivors shall fall by the sword. They shall seize your sons and your daughters, and your survivors shall be devoured by fire.
EZEK|23|26|They shall also strip you of your clothes and take away your beautiful jewels.
EZEK|23|27|Thus I will put an end to your lewdness and your whoring begun in the land of Egypt, so that you shall not lift up your eyes to them or remember Egypt anymore.
EZEK|23|28|"For thus says the Lord GOD: Behold, I will deliver you into the hands of those whom you hate, into the hands of those from whom you turned in disgust,
EZEK|23|29|and they shall deal with you in hatred and take away all the fruit of your labor and leave you naked and bare, and the nakedness of your whoring shall be uncovered. Your lewdness and your whoring
EZEK|23|30|have brought this upon you, because you played the whore with the nations and defiled yourself with their idols.
EZEK|23|31|You have gone the way of your sister; therefore I will give her cup into your hand.
EZEK|23|32|Thus says the Lord GOD: "You shall drink your sister's cup that is deep and large; you shall be laughed at and held in derision, for it contains much;
EZEK|23|33|you will be filled with drunkenness and sorrow. A cup of horror and desolation, the cup of your sister Samaria;
EZEK|23|34|you shall drink it and drain it out, and gnaw its shards, and tear your breasts; for I have spoken, declares the Lord GOD.
EZEK|23|35|Therefore thus says the Lord GOD: Because you have forgotten me and cast me behind your back, you yourself must bear the consequences of your lewdness and whoring."
EZEK|23|36|The LORD said to me: "Son of man, will you judge Oholah and Oholibah? Declare to them their abominations.
EZEK|23|37|For they have committed adultery, and blood is on their hands. With their idols they have committed adultery, and they have even offered up to them for food the children whom they had borne to me.
EZEK|23|38|Moreover, this they have done to me: they have defiled my sanctuary on the same day and profaned my Sabbaths.
EZEK|23|39|For when they had slaughtered their children in sacrifice to their idols, on the same day they came into my sanctuary to profane it. And behold, this is what they did in my house.
EZEK|23|40|They even sent for men to come from far, to whom a messenger was sent; and behold, they came. For them you bathed yourself, painted your eyes, and adorned yourself with ornaments.
EZEK|23|41|You sat on a stately couch, with a table spread before it on which you had placed my incense and my oil.
EZEK|23|42|The sound of a carefree multitude was with her; and with men of the common sort drunkards were brought from the wilderness; and they put bracelets on the hands of the women, and beautiful crowns on their heads.
EZEK|23|43|"Then I said of her who was worn out by adultery, Now they will continue to use her for a whore, even her!
EZEK|23|44|For they have gone in to her, as men go in to a prostitute. Thus they went in to Oholah and to Oholibah, lewd women!
EZEK|23|45|But righteous men shall pass judgment on them with the sentence of adulteresses, and with the sentence of women who shed blood, because they are adulteresses, and blood is on their hands."
EZEK|23|46|For thus says the Lord GOD: "Bring up a vast host against them, and make them an object of terror and a plunder.
EZEK|23|47|And the host shall stone them and cut them down with their swords. They shall kill their sons and their daughters, and burn up their houses.
EZEK|23|48|Thus will I put an end to lewdness in the land, that all women may take warning and not commit lewdness as you have done.
EZEK|23|49|And they shall return your lewdness upon you, and you shall bear the penalty for your sinful idolatry, and you shall know that I am the Lord GOD."
EZEK|24|1|In the ninth year, in the tenth month, on the tenth day of the month, the word of the LORD came to me:
EZEK|24|2|"Son of man, write down the name of this day, this very day. The king of Babylon has laid siege to Jerusalem this very day.
EZEK|24|3|And utter a parable to the rebellious house and say to them, Thus says the Lord GOD: "Set on the pot, set it on; pour in water also;
EZEK|24|4|put in it the pieces of meat, all the good pieces, the thigh and the shoulder; fill it with choice bones.
EZEK|24|5|Take the choicest one of the flock; pile the logs under it; boil it well; seethe also its bones in it.
EZEK|24|6|"Therefore thus says the Lord GOD: Woe to the bloody city, to the pot whose corrosion is in it, and whose corrosion has not gone out of it! Take out of it piece after piece, without making any choice.
EZEK|24|7|For the blood she has shed is in her midst; she put it on the bare rock; she did not pour it out on the ground to cover it with dust.
EZEK|24|8|To rouse my wrath, to take vengeance, I have set on the bare rock the blood she has shed, that it may not be covered.
EZEK|24|9|Therefore thus says the Lord GOD: Woe to the bloody city! I also will make the pile great.
EZEK|24|10|Heap on the logs, kindle the fire, boil the meat well, mix in the spices, and let the bones be burned up.
EZEK|24|11|Then set it empty upon the coals, that it may become hot, and its copper may burn, that its uncleanness may be melted in it, its corrosion consumed.
EZEK|24|12|She has wearied herself with toil; its abundant corrosion does not go out of it. Into the fire with its corrosion!
EZEK|24|13|On account of your unclean lewdness, because I would have cleansed you and you were not cleansed from your uncleanness, you shall not be cleansed anymore till I have satisfied my fury upon you.
EZEK|24|14|I am the LORD. I have spoken; it shall come to pass; I will do it. I will not go back; I will not spare; I will not relent; according to your ways and your deeds you will be judged, declares the Lord GOD."
EZEK|24|15|The word of the LORD came to me:
EZEK|24|16|"Son of man, behold, I am about to take the delight of your eyes away from you at a stroke; yet you shall not mourn or weep, nor shall your tears run down.
EZEK|24|17|Sigh, but not aloud; make no mourning for the dead. Bind on your turban, and put your shoes on your feet; do not cover your lips, nor eat the bread of men."
EZEK|24|18|So I spoke to the people in the morning, and at evening my wife died. And on the next morning I did as I was commanded.
EZEK|24|19|And the people said to me, "Will you not tell us what these things mean for us, that you are acting thus?"
EZEK|24|20|Then I said to them, "The word of the LORD came to me:
EZEK|24|21|'Say to the house of Israel, Thus says the Lord GOD: Behold, I will profane my sanctuary, the pride of your power, the delight of your eyes, and the yearning of your soul, and your sons and your daughters whom you left behind shall fall by the sword.
EZEK|24|22|And you shall do as I have done; you shall not cover your lips, nor eat the bread of men.
EZEK|24|23|Your turbans shall be on your heads and your shoes on your feet; you shall not mourn or weep, but you shall rot away in your iniquities and groan to one another.
EZEK|24|24|Thus shall Ezekiel be to you a sign; according to all that he has done you shall do. When this comes, then you will know that I am the Lord GOD.'
EZEK|24|25|"As for you, son of man, surely on the day when I take from them their stronghold, their joy and glory, the delight of their eyes and their soul's desire, and also their sons and daughters,
EZEK|24|26|on that day a fugitive will come to you to report to you the news.
EZEK|24|27|On that day your mouth will be opened to the fugitive, and you shall speak and be no longer mute. So you will be a sign to them, and they will know that I am the LORD."
EZEK|25|1|The word of the LORD came to me:
EZEK|25|2|"Son of man, set your face toward the Ammonites and prophesy against them.
EZEK|25|3|Say to the Ammonites, Hear the word of the Lord GOD: Thus says the Lord GOD, Because you said, 'Aha!' over my sanctuary when it was profaned, and over the land of Israel when it was made desolate, and over the house of Judah when they went into exile,
EZEK|25|4|therefore behold, I am handing you over to the people of the East for a possession, and they shall set their encampments among you and make their dwellings in your midst. They shall eat your fruit, and they shall drink your milk.
EZEK|25|5|I will make Rabbah a pasture for camels and Ammon a fold for flocks. Then you will know that I am the LORD.
EZEK|25|6|For thus says the Lord GOD: Because you have clapped your hands and stamped your feet and rejoiced with all the malice within your soul against the land of Israel,
EZEK|25|7|therefore, behold, I have stretched out my hand against you, and will hand you over as plunder to the nations. And I will cut you off from the peoples and will make you perish out of the countries; I will destroy you. Then you will know that I am the LORD.
EZEK|25|8|"Thus says the Lord GOD: Because Moab and Seir said, 'Behold, the house of Judah is like all the other nations,'
EZEK|25|9|therefore I will lay open the flank of Moab from the cities, from its cities on its frontier, the glory of the country, Bethjeshimoth, Baal-meon, and Kiriathaim.
EZEK|25|10|I will give it along with the Ammonites to the people of the East as a possession, that the Ammonites may be remembered no more among the nations,
EZEK|25|11|and I will execute judgments upon Moab. Then they will know that I am the LORD.
EZEK|25|12|"Thus says the Lord GOD: Because Edom acted revengefully against the house of Judah and has grievously offended in taking vengeance on them,
EZEK|25|13|therefore thus says the Lord GOD, I will stretch out my hand against Edom and cut off from it man and beast. And I will make it desolate; from Teman even to Dedan they shall fall by the sword.
EZEK|25|14|And I will lay my vengeance upon Edom by the hand of my people Israel, and they shall do in Edom according to my anger and according to my wrath, and they shall know my vengeance, declares the Lord GOD.
EZEK|25|15|"Thus says the Lord GOD: Because the Philistines acted revengefully and took vengeance with malice of soul to destroy in never-ending enmity,
EZEK|25|16|therefore thus says the Lord GOD, Behold, I will stretch out my hand against the Philistines, and I will cut off the Cherethites and destroy the rest of the seacoast.
EZEK|25|17|I will execute great vengeance on them with wrathful rebukes. Then they will know that I am the LORD, when I lay my vengeance upon them."
EZEK|26|1|In the eleventh year, on the first day of the month, the word of the LORD came to me:
EZEK|26|2|"Son of man, because Tyre said concerning Jerusalem, 'Aha, the gate of the peoples is broken; it has swung open to me. I shall be replenished, now that she is laid waste,'
EZEK|26|3|therefore thus says the Lord GOD: Behold, I am against you, O Tyre, and will bring up many nations against you, as the sea brings up its waves.
EZEK|26|4|They shall destroy the walls of Tyre and break down her towers, and I will scrape her soil from her and make her a bare rock.
EZEK|26|5|She shall be in the midst of the sea a place for the spreading of nets, for I have spoken, declares the Lord GOD. And she shall become plunder for the nations,
EZEK|26|6|and her daughters on the mainland shall be killed by the sword. Then they will know that I am the LORD.
EZEK|26|7|"For thus says the Lord GOD: Behold, I will bring against Tyre from the north Nebuchadnezzar king of Babylon, king of kings, with horses and chariots, and with horsemen and a host of many soldiers.
EZEK|26|8|He will kill with the sword your daughters on the mainland. He will set up a siege wall against you and throw up a mound against you, and raise a roof of shields against you.
EZEK|26|9|He will direct the shock of his battering rams against your walls, and with his axes he will break down your towers.
EZEK|26|10|His horses will be so many that their dust will cover you. Your walls will shake at the noise of the horsemen and wagons and chariots, when he enters your gates as men enter a city that has been breached.
EZEK|26|11|With the hoofs of his horses he will trample all your streets. He will kill your people with the sword, and your mighty pillars will fall to the ground.
EZEK|26|12|They will plunder your riches and loot your merchandise. They will break down your walls and destroy your pleasant houses. Your stones and timber and soil they will cast into the midst of the waters.
EZEK|26|13|And I will stop the music of your songs, and the sound of your lyres shall be heard no more.
EZEK|26|14|I will make you a bare rock. You shall be a place for the spreading of nets. You shall never be rebuilt, for I am the LORD; I have spoken, declares the Lord GOD.
EZEK|26|15|"Thus says the Lord GOD to Tyre: Will not the coastlands shake at the sound of your fall, when the wounded groan, when slaughter is made in your midst?
EZEK|26|16|Then all the princes of the sea will step down from their thrones and remove their robes and strip off their embroidered garments. They will clothe themselves with trembling; they will sit on the ground and tremble every moment and be appalled at you.
EZEK|26|17|And they will raise a lamentation over you and say to you, "' How you have perished, you who were inhabited from the seas, O city renowned, who was mighty on the sea; she and her inhabitants imposed their terror on all her inhabitants!
EZEK|26|18|Now the coastlands tremble on the day of your fall, and the coastlands that are on the sea are dismayed at your passing.'
EZEK|26|19|"For thus says the Lord GOD: When I make you a city laid waste, like the cities that are not inhabited, when I bring up the deep over you, and the great waters cover you,
EZEK|26|20|then I will make you go down with those who go down to the pit, to the people of old, and I will make you to dwell in the world below, among ruins from of old, with those who go down to the pit, so that you will not be inhabited; but I will set beauty in the land of the living.
EZEK|26|21|I will bring you to a dreadful end, and you shall be no more. Though you be sought for, you will never be found again, declares the Lord GOD."
EZEK|27|1|The word of the LORD came to me:
EZEK|27|2|"Now you, son of man, raise a lamentation over Tyre,
EZEK|27|3|and say to Tyre, who dwells at the entrances to the sea, merchant of the peoples to many coastlands, thus says the Lord GOD: "O Tyre, you have said, 'I am perfect in beauty.'
EZEK|27|4|Your borders are in the heart of the seas; your builders made perfect your beauty.
EZEK|27|5|They made all your planks of fir trees from Senir; they took a cedar from Lebanon to make a mast for you.
EZEK|27|6|Of oaks of Bashan they made your oars; they made your deck of pines from the coasts of Cyprus, inlaid with ivory.
EZEK|27|7|Of fine embroidered linen from Egypt was your sail, serving as your banner; blue and purple from the coasts of Elishah was your awning.
EZEK|27|8|The inhabitants of Sidon and Arvad were your rowers; your skilled men, O Tyre, were in you; they were your pilots.
EZEK|27|9|The elders of Gebal and her skilled men were in you, caulking your seams; all the ships of the sea with their mariners were in you to barter for your wares.
EZEK|27|10|"Persia and Lud and Put were in your army as your men of war. They hung the shield and helmet in you; they gave you splendor.
EZEK|27|11|Men of Arvad and Helech were on your walls all around, and men of Gamad were in your towers. They hung their shields on your walls all around; they made perfect your beauty.
EZEK|27|12|"Tarshish did business with you because of your great wealth of every kind; silver, iron, tin, and lead they exchanged for your wares.
EZEK|27|13|Javan, Tubal, and Meshech traded with you; they exchanged human beings and vessels of bronze for your merchandise.
EZEK|27|14|From Beth-togarmah they exchanged horses, war horses, and mules for your wares.
EZEK|27|15|The men of Dedan traded with you. Many coastlands were your own special markets; they brought you in payment ivory tusks and ebony.
EZEK|27|16|Syria did business with you because of your abundant goods; they exchanged for your wares emeralds, purple, embroidered work, fine linen, coral, and ruby.
EZEK|27|17|Judah and the land of Israel traded with you; they exchanged for your merchandise wheat of Minnith, meal, honey, oil, and balm.
EZEK|27|18|Damascus did business with you for your abundant goods, because of your great wealth of every kind; wine of Helbon and wool of Sahar
EZEK|27|19|and casks of wine from Uzal they exchanged for your wares; wrought iron, cassia, and calamus were bartered for your merchandise.
EZEK|27|20|Dedan traded with you in saddlecloths for riding.
EZEK|27|21|Arabia and all the princes of Kedar were your favored dealers in lambs, rams, and goats; in these they did business with you.
EZEK|27|22|The traders of Sheba and Raamah traded with you; they exchanged for your wares the best of all kinds of spices and all precious stones and gold.
EZEK|27|23|Haran, Canneh, Eden, traders of Sheba, Asshur, and Chilmad traded with you.
EZEK|27|24|In your market these traded with you in choice garments, in clothes of blue and embroidered work, and in carpets of colored material, bound with cords and made secure.
EZEK|27|25|The ships of Tarshish traveled for you with your merchandise. So you were filled and heavily laden in the heart of the seas.
EZEK|27|26|"Your rowers have brought you out into the high seas. The east wind has wrecked you in the heart of the seas.
EZEK|27|27|Your riches, your wares, your merchandise, your mariners and your pilots, your caulkers, your dealers in merchandise, and all your men of war who are in you, with all your crew that is in your midst, sink into the heart of the seas on the day of your fall.
EZEK|27|28|At the sound of the cry of your pilots the countryside shakes,
EZEK|27|29|and down from their ships come all who handle the oar. The mariners and all the pilots of the sea stand on the land
EZEK|27|30|and shout aloud over you and cry out bitterly. They cast dust on their heads and wallow in ashes;
EZEK|27|31|they make themselves bald for you and put sackcloth on their waist, and they weep over you in bitterness of soul, with bitter mourning.
EZEK|27|32|In their wailing they raise a lamentation for you and lament over you: 'Who is like Tyre, like one destroyed in the midst of the sea?
EZEK|27|33|When your wares came from the seas, you satisfied many peoples; with your abundant wealth and merchandise you enriched the kings of the earth.
EZEK|27|34|Now you are wrecked by the seas, in the depths of the waters; your merchandise and all your crew in your midst have sunk with you.
EZEK|27|35|All the inhabitants of the coastlands are appalled at you, and the hair of their kings bristles with horror; their faces are convulsed.
EZEK|27|36|The merchants among the peoples hiss at you; you have come to a dreadful end and shall be no more forever.'"
EZEK|28|1|The word of the LORD came to me:
EZEK|28|2|"Son of man, say to the prince of Tyre, Thus says the Lord GOD: "Because your heart is proud, and you have said, 'I am a god, I sit in the seat of the gods, in the heart of the seas,' yet you are but a man, and no god, though you make your heart like the heart of a god-
EZEK|28|3|you are indeed wiser than Daniel; no secret is hidden from you;
EZEK|28|4|by your wisdom and your understanding you have made wealth for yourself, and have gathered gold and silver into your treasuries;
EZEK|28|5|by your great wisdom in your trade you have increased your wealth, and your heart has become proud in your wealth-
EZEK|28|6|therefore thus says the Lord GOD: Because you make your heart like the heart of a god,
EZEK|28|7|therefore, behold, I will bring foreigners upon you, the most ruthless of the nations; and they shall draw their swords against the beauty of your wisdom and defile your splendor.
EZEK|28|8|They shall thrust you down into the pit, and you shall die the death of the slain in the heart of the seas.
EZEK|28|9|Will you still say, 'I am a god,' in the presence of those who kill you, though you are but a man, and no god, in the hands of those who slay you?
EZEK|28|10|You shall die the death of the uncircumcised by the hand of foreigners; for I have spoken, declares the Lord GOD."
EZEK|28|11|Moreover, the word of the LORD came to me:
EZEK|28|12|"Son of man, raise a lamentation over the king of Tyre, and say to him, Thus says the Lord GOD: "You were the signet of perfection, full of wisdom and perfect in beauty.
EZEK|28|13|You were in Eden, the garden of God; every precious stone was your covering, sardius, topaz, and diamond, beryl, onyx, and jasper, sapphire, emerald, and carbuncle; and crafted in gold were your settings and your engravings. On the day that you were created they were prepared.
EZEK|28|14|You were an anointed guardian cherub. I placed you; you were on the holy mountain of God; in the midst of the stones of fire you walked.
EZEK|28|15|You were blameless in your ways from the day you were created, till unrighteousness was found in you.
EZEK|28|16|In the abundance of your trade you were filled with violence in your midst, and you sinned; so I cast you as a profane thing from the mountain of God, and I destroyed you, O guardian cherub, from the midst of the stones of fire.
EZEK|28|17|Your heart was proud because of your beauty; you corrupted your wisdom for the sake of your splendor. I cast you to the ground; I exposed you before kings, to feast their eyes on you.
EZEK|28|18|By the multitude of your iniquities, in the unrighteousness of your trade you profaned your sanctuaries; so I brought fire out from your midst; it consumed you, and I turned you to ashes on the earth in the sight of all who saw you.
EZEK|28|19|All who know you among the peoples are appalled at you; you have come to a dreadful end and shall be no more forever."
EZEK|28|20|The word of the LORD came to me:
EZEK|28|21|"Son of man, set your face toward Sidon, and prophesy against her
EZEK|28|22|and say, Thus says the Lord GOD: "Behold, I am against you, O Sidon, and I will manifest my glory in your midst. And they shall know that I am the LORD when I execute judgments in her and manifest my holiness in her;
EZEK|28|23|for I will send pestilence into her, and blood into her streets; and the slain shall fall in her midst, by the sword that is against her on every side. Then they will know that I am the LORD.
EZEK|28|24|"And for the house of Israel there shall be no more a brier to prick or a thorn to hurt them among all their neighbors who have treated them with contempt. Then they will know that I am the Lord GOD.
EZEK|28|25|"Thus says the Lord GOD: When I gather the house of Israel from the peoples among whom they are scattered, and manifest my holiness in them in the sight of the nations, then they shall dwell in their own land that I gave to my servant Jacob.
EZEK|28|26|And they shall dwell securely in it, and they shall build houses and plant vineyards. They shall dwell securely, when I execute judgments upon all their neighbors who have treated them with contempt. Then they will know that I am the LORD their God."
EZEK|29|1|In the tenth year, in the tenth month, on the twelfth day of the month, the word of the LORD came to me:
EZEK|29|2|"Son of man, set your face against Pharaoh king of Egypt, and prophesy against him and against all Egypt;
EZEK|29|3|speak, and say, Thus says the Lord GOD: "Behold, I am against you, Pharaoh king of Egypt, the great dragon that lies in the midst of his streams, that says, 'My Nile is my own; I made it for myself.'
EZEK|29|4|I will put hooks in your jaws, and make the fish of your streams stick to your scales; and I will draw you up out of the midst of your streams, with all the fish of your streams that stick to your scales.
EZEK|29|5|And I will cast you out into the wilderness, you and all the fish of your streams; you shall fall on the open field, and not be brought together or gathered. To the beasts of the earth and to the birds of the heavens I give you as food.
EZEK|29|6|Then all the inhabitants of Egypt shall know that I am the LORD. "Because you have been a staff of reed to the house of Israel;
EZEK|29|7|when they grasped you with the hand, you broke and tore all their shoulders; and when they leaned on you, you broke and made all their loins to shake.
EZEK|29|8|Therefore thus says the Lord GOD: Behold, I will bring a sword upon you, and will cut off from you man and beast,
EZEK|29|9|and the land of Egypt shall be a desolation and a waste. Then they will know that I am the LORD. "Because you said, 'The Nile is mine, and I made it,'
EZEK|29|10|therefore, behold, I am against you and against your streams, and I will make the land of Egypt an utter waste and desolation, from Migdol to Syene, as far as the border of Cush.
EZEK|29|11|No foot of man shall pass through it, and no foot of beast shall pass through it; it shall be uninhabited forty years.
EZEK|29|12|And I will make the land of Egypt a desolation in the midst of desolated countries, and her cities shall be a desolation forty years among cities that are laid waste. I will scatter the Egyptians among the nations, and disperse them through the countries.
EZEK|29|13|"For thus says the Lord GOD: At the end of forty years I will gather the Egyptians from the peoples among whom they were scattered,
EZEK|29|14|and I will restore the fortunes of Egypt and bring them back to the land of Pathros, the land of their origin, and there they shall be a lowly kingdom.
EZEK|29|15|It shall be the most lowly of the kingdoms, and never again exalt itself above the nations. And I will make them so small that they will never again rule over the nations.
EZEK|29|16|And it shall never again be the reliance of the house of Israel, recalling their iniquity, when they turn to them for aid. Then they will know that I am the Lord GOD."
EZEK|29|17|In the twenty-seventh year, in the first month, on the first day of the month, the word of the LORD came to me:
EZEK|29|18|"Son of man, Nebuchadnezzar king of Babylon made his army labor hard against Tyre. Every head was made bald, and every shoulder was rubbed bare, yet neither he nor his army got anything from Tyre to pay for the labor that he had performed against her.
EZEK|29|19|Therefore thus says the Lord GOD: Behold, I will give the land of Egypt to Nebuchadnezzar king of Babylon; and he shall carry off its wealth and despoil it and plunder it; and it shall be the wages for his army.
EZEK|29|20|I have given him the land of Egypt as his payment for which he labored, because they worked for me, declares the Lord GOD.
EZEK|29|21|"On that day I will cause a horn to spring up for the house of Israel, and I will open your lips among them. Then they will know that I am the LORD."
EZEK|30|1|The word of the LORD came to me:
EZEK|30|2|"Son of man, prophesy, and say, Thus says the Lord GOD: "Wail, 'Alas for the day!'
EZEK|30|3|For the day is near, the day of the LORD is near; it will be a day of clouds, a time of doom for the nations.
EZEK|30|4|A sword shall come upon Egypt, and anguish shall be in Cush, when the slain fall in Egypt, and her wealth is carried away, and her foundations are torn down.
EZEK|30|5|Cush, and Put, and Lud, and all Arabia, and Libya, and the people of the land that is in league, shall fall with them by the sword.
EZEK|30|6|"Thus says the LORD: Those who support Egypt shall fall, and her proud might shall come down; from Migdol to Syene they shall fall within her by the sword, declares the Lord GOD.
EZEK|30|7|And they shall be desolated in the midst of desolated countries, and their cities shall be in the midst of cities that are laid waste.
EZEK|30|8|Then they will know that I am the LORD, when I have set fire to Egypt, and all her helpers are broken.
EZEK|30|9|"On that day messengers shall go out from me in ships to terrify the unsuspecting people of Cush, and anguish shall come upon them on the day of Egypt's doom; for, behold, it comes!
EZEK|30|10|"Thus says the Lord GOD: "I will put an end to the wealth of Egypt, by the hand of Nebuchadnezzar king of Babylon.
EZEK|30|11|He and his people with him, the most ruthless of nations, shall be brought in to destroy the land, and they shall draw their swords against Egypt and fill the land with the slain.
EZEK|30|12|And I will dry up the Nile and will sell the land into the hand of evildoers; I will bring desolation upon the land and everything in it, by the hand of foreigners; I am the LORD; I have spoken.
EZEK|30|13|"Thus says the Lord GOD: "I will destroy the idols and put an end to the images in Memphis; there shall no longer be a prince from the land of Egypt; so I will put fear in the land of Egypt.
EZEK|30|14|I will make Pathros a desolation and will set fire to Zoan and will execute judgments on Thebes.
EZEK|30|15|And I will pour out my wrath on Pelusium, the stronghold of Egypt, and cut off the multitude of Thebes.
EZEK|30|16|And I will set fire to Egypt; Pelusium shall be in great agony; Thebes shall be breached, and Memphis shall face enemies by day.
EZEK|30|17|The young men of On and of Pibeseth shall fall by the sword, and the women shall go into captivity.
EZEK|30|18|At Tehaphnehes the day shall be dark, when I break there the yoke bars of Egypt, and her proud might shall come to an end in her; she shall be covered by a cloud, and her daughters shall go into captivity.
EZEK|30|19|Thus I will execute judgments on Egypt. Then they will know that I am the LORD."
EZEK|30|20|In the eleventh year, in the first month, on the seventh day of the month, the word of the LORD came to me:
EZEK|30|21|"Son of man, I have broken the arm of Pharaoh king of Egypt, and behold, it has not been bound up, to heal it by binding it with a bandage, so that it may become strong to wield the sword.
EZEK|30|22|Therefore thus says the Lord GOD: Behold, I am against Pharaoh king of Egypt and will break his arms, both the strong arm and the one that was broken, and I will make the sword fall from his hand.
EZEK|30|23|I will scatter the Egyptians among the nations and disperse them through the countries.
EZEK|30|24|And I will strengthen the arms of the king of Babylon and put my sword in his hand, but I will break the arms of Pharaoh, and he will groan before him like a man mortally wounded.
EZEK|30|25|I will strengthen the arms of the king of Babylon, but the arms of Pharaoh shall fall. Then they shall know that I am the LORD, when I put my sword into the hand of the king of Babylon and he stretches it out against the land of Egypt.
EZEK|30|26|And I will scatter the Egyptians among the nations and disperse them throughout the countries. Then they will know that I am the LORD."
EZEK|31|1|In the eleventh year, in the third month, on the first day of the month, the word of the LORD came to me:
EZEK|31|2|"Son of man, say to Pharaoh king of Egypt and to his multitude: "Whom are you like in your greatness?
EZEK|31|3|Behold, Assyria was a cedar in Lebanon, with beautiful branches and forest shade, and of towering height, its top among the clouds.
EZEK|31|4|The waters nourished it; the deep made it grow tall, making its rivers flow around the place of its planting, sending forth its streams to all the trees of the field.
EZEK|31|5|So it towered high above all the trees of the field; its boughs grew large and its branches long from abundant water in its shoots.
EZEK|31|6|All the birds of the heavens made their nests in its boughs; under its branches all the beasts of the field gave birth to their young, and under its shadow lived all great nations.
EZEK|31|7|It was beautiful in its greatness, in the length of its branches; for its roots went down to abundant waters.
EZEK|31|8|The cedars in the garden of God could not rival it, nor the fir trees equal its boughs; neither were the plane trees like its branches; no tree in the garden of God was its equal in beauty.
EZEK|31|9|I made it beautiful in the mass of its branches, and all the trees of Eden envied it, that were in the garden of God.
EZEK|31|10|"Therefore thus says the Lord GOD: Because it towered high and set its top among the clouds, and its heart was proud of its height,
EZEK|31|11|I will give it into the hand of a mighty one of the nations. He shall surely deal with it as its wickedness deserves. I have cast it out.
EZEK|31|12|Foreigners, the most ruthless of nations, have cut it down and left it. On the mountains and in all the valleys its branches have fallen, and its boughs have been broken in all the ravines of the land, and all the peoples of the earth have gone away from its shadow and left it.
EZEK|31|13|On its fallen trunk dwell all the birds of the heavens, and on its branches are all the beasts of the field.
EZEK|31|14|All this is in order that no trees by the waters may grow to towering height or set their tops among the clouds, and that no trees that drink water may reach up to them in height. For they are all given over to death, to the world below, among the children of man, with those who go down to the pit.
EZEK|31|15|"Thus says the Lord GOD: On the day the cedar went down to Sheol I caused mourning; I closed the deep over it, and restrained its rivers, and many waters were stopped. I clothed Lebanon in gloom for it, and all the trees of the field fainted because of it.
EZEK|31|16|I made the nations quake at the sound of its fall, when I cast it down to Sheol with those who go down to the pit. And all the trees of Eden, the choice and best of Lebanon, all that drink water, were comforted in the world below.
EZEK|31|17|They also went down to Sheol with it, to those who are slain by the sword; yes, those who were its arm, who lived under its shadow among the nations.
EZEK|31|18|"Whom are you thus like in glory and in greatness among the trees of Eden? You shall be brought down with the trees of Eden to the world below. You shall lie among the uncircumcised, with those who are slain by the sword. "This is Pharaoh and all his multitude, declares the Lord GOD."
EZEK|32|1|In the twelfth year, in the twelfth month, on the first day of the month, the word of the LORD came to me:
EZEK|32|2|"Son of man, raise a lamentation over Pharaoh king of Egypt and say to him: "You consider yourself a lion of the nations, but you are like a dragon in the seas; you burst forth in your rivers, trouble the waters with your feet, and foul their rivers.
EZEK|32|3|Thus says the Lord GOD: I will throw my net over you with a host of many peoples, and they will haul you up in my dragnet.
EZEK|32|4|And I will cast you on the ground; on the open field I will fling you, and will cause all the birds of the heavens to settle on you, and I will gorge the beasts of the whole earth with you.
EZEK|32|5|I will strew your flesh upon the mountains and fill the valleys with your carcass.
EZEK|32|6|I will drench the land even to the mountains with your flowing blood, and the ravines will be full of you.
EZEK|32|7|When I blot you out, I will cover the heavens and make their stars dark; I will cover the sun with a cloud, and the moon shall not give its light.
EZEK|32|8|All the bright lights of heaven will I make dark over you, and put darkness on your land, declares the Lord GOD.
EZEK|32|9|"I will trouble the hearts of many peoples, when I bring your destruction among the nations, into the countries that you have not known.
EZEK|32|10|I will make many peoples appalled at you, and the hair of their kings shall bristle with horror because of you, when I brandish my sword before them. They shall tremble every moment, every one for his own life, on the day of your downfall.
EZEK|32|11|"For thus says the Lord GOD: The sword of the king of Babylon shall come upon you.
EZEK|32|12|I will cause your multitude to fall by the swords of mighty ones, all of them most ruthless of nations. "They shall bring to ruin the pride of Egypt, and all its multitude shall perish.
EZEK|32|13|I will destroy all its beasts from beside many waters; and no foot of man shall trouble them anymore, nor shall the hoofs of beasts trouble them.
EZEK|32|14|Then I will make their waters clear, and cause their rivers to run like oil, declares the Lord GOD.
EZEK|32|15|When I make the land of Egypt desolate, and when the land is desolate of all that fills it, when I strike down all who dwell in it, then they will know that I am the LORD.
EZEK|32|16|This is a lamentation that shall be chanted; the daughters of the nations shall chant it; over Egypt, and over all her multitude, shall they chant it, declares the Lord GOD."
EZEK|32|17|In the twelfth year, in the twelfth month, on the fifteenth day of the month, the word of the LORD came to me:
EZEK|32|18|"Son of man, wail over the multitude of Egypt, and send them down, her and the daughters of majestic nations, to the world below, to those who have gone down to the pit:
EZEK|32|19|'Whom do you surpass in beauty? Go down and be laid to rest with the uncircumcised.'
EZEK|32|20|They shall fall amid those who are slain by the sword. Egypt is delivered to the sword; drag her away, and all her multitudes.
EZEK|32|21|The mighty chiefs shall speak of them, with their helpers, out of the midst of Sheol: 'They have come down, they lie still, the uncircumcised, slain by the sword.'
EZEK|32|22|"Assyria is there, and all her company, its graves all around it, all of them slain, fallen by the sword,
EZEK|32|23|whose graves are set in the uttermost parts of the pit; and her company is all around her grave, all of them slain, fallen by the sword, who spread terror in the land of the living.
EZEK|32|24|"Elam is there, and all her multitude around her grave; all of them slain, fallen by the sword, who went down uncircumcised into the world below, who spread their terror in the land of the living; and they bear their shame with those who go down to the pit.
EZEK|32|25|They have made her a bed among the slain with all her multitude, her graves all around it, all of them uncircumcised, slain by the sword; for terror of them was spread in the land of the living, and they bear their shame with those who go down to the pit; they are placed among the slain.
EZEK|32|26|"Meshech-Tubal is there, and all her multitude, her graves all around it, all of them uncircumcised, slain by the sword; for they spread their terror in the land of the living.
EZEK|32|27|And they do not lie with the mighty, the fallen from among the uncircumcised, who went down to Sheol with their weapons of war, whose swords were laid under their heads, and whose iniquities are upon their bones; for the terror of the mighty men was in the land of the living.
EZEK|32|28|But as for you, you shall be broken and lie among the uncircumcised, with those who are slain by the sword.
EZEK|32|29|"Edom is there, her kings and all her princes, who for all their might are laid with those who are killed by the sword; they lie with the uncircumcised, with those who go down to the pit.
EZEK|32|30|"The princes of the north are there, all of them, and all the Sidonians, who have gone down in shame with the slain, for all the terror that they caused by their might; they lie uncircumcised with those who are slain by the sword, and bear their shame with those who go down to the pit.
EZEK|32|31|"When Pharaoh sees them, he will be comforted for all his multitude, Pharaoh and all his army, slain by the sword, declares the Lord GOD.
EZEK|32|32|For I spread terror in the land of the living; and he shall be laid to rest among the uncircumcised, with those who are slain by the sword, Pharaoh and all his multitude, declares the Lord GOD."
EZEK|33|1|The word of the LORD came to me:
EZEK|33|2|"Son of man, speak to your people and say to them, If I bring the sword upon a land, and the people of the land take a man from among them, and make him their watchman,
EZEK|33|3|and if he sees the sword coming upon the land and blows the trumpet and warns the people,
EZEK|33|4|then if anyone who hears the sound of the trumpet does not take warning, and the sword comes and takes him away, his blood shall be upon his own head.
EZEK|33|5|He heard the sound of the trumpet and did not take warning; his blood shall be upon himself. But if he had taken warning, he would have saved his life.
EZEK|33|6|But if the watchman sees the sword coming and does not blow the trumpet, so that the people are not warned, and the sword comes and takes any one of them, that person is taken away in his iniquity, but his blood I will require at the watchman's hand.
EZEK|33|7|"So you, son of man, I have made a watchman for the house of Israel. Whenever you hear a word from my mouth, you shall give them warning from me.
EZEK|33|8|If I say to the wicked, O wicked one, you shall surely die, and you do not speak to warn the wicked to turn from his way, that wicked person shall die in his iniquity, but his blood I will require at your hand.
EZEK|33|9|But if you warn the wicked to turn from his way, and he does not turn from his way, that person shall die in his iniquity, but you will have delivered your soul.
EZEK|33|10|"And you, son of man, say to the house of Israel, Thus have you said: 'Surely our transgressions and our sins are upon us, and we rot away because of them. How then can we live?'
EZEK|33|11|Say to them, As I live, declares the Lord GOD, I have no pleasure in the death of the wicked, but that the wicked turn from his way and live; turn back, turn back from your evil ways, for why will you die, O house of Israel?
EZEK|33|12|"And you, son of man, say to your people, The righteousness of the righteous shall not deliver him when he transgresses, and as for the wickedness of the wicked, he shall not fall by it when he turns from his wickedness, and the righteous shall not be able to live by his righteousness when he sins.
EZEK|33|13|Though I say to the righteous that he shall surely live, yet if he trusts in his righteousness and does injustice, none of his righteous deeds shall be remembered, but in his injustice that he has done he shall die.
EZEK|33|14|Again, though I say to the wicked, 'You shall surely die,' yet if he turns from his sin and does what is just and right,
EZEK|33|15|if the wicked restores the pledge, gives back what he has taken by robbery, and walks in the statutes of life, not doing injustice, he shall surely live; he shall not die.
EZEK|33|16|None of the sins that he has committed shall be remembered against him. He has done what is just and right; he shall surely live.
EZEK|33|17|"Yet your people say, 'The way of the Lord is not just,' when it is their own way that is not just.
EZEK|33|18|When the righteous turns from his righteousness and does injustice, he shall die for it.
EZEK|33|19|And when the wicked turns from his wickedness and does what is just and right, he shall live by them.
EZEK|33|20|Yet you say, 'The way of the Lord is not just.' O house of Israel, I will judge each of you according to his ways."
EZEK|33|21|In the twelfth year of our exile, in the tenth month, on the fifth day of the month, a fugitive from Jerusalem came to me and said, "The city has been struck down."
EZEK|33|22|Now the hand of the LORD had been upon me the evening before the fugitive came; and he had opened my mouth by the time the man came to me in the morning, so my mouth was opened, and I was no longer mute.
EZEK|33|23|The word of the LORD came to me:
EZEK|33|24|"Son of man, the inhabitants of these waste places in the land of Israel keep saying, 'Abraham was only one man, yet he got possession of the land; but we are many; the land is surely given us to possess.'
EZEK|33|25|Therefore say to them, Thus says the Lord GOD: You eat flesh with the blood and lift up your eyes to your idols and shed blood; shall you then possess the land?
EZEK|33|26|You rely on the sword, you commit abominations, and each of you defiles his neighbor's wife; shall you then possess the land?
EZEK|33|27|Say this to them, Thus says the Lord GOD: As I live, surely those who are in the waste places shall fall by the sword, and whoever is in the open field I will give to the beasts to be devoured, and those who are in strongholds and in caves shall die by pestilence.
EZEK|33|28|And I will make the land a desolation and a waste, and her proud might shall come to an end, and the mountains of Israel shall be so desolate that none will pass through.
EZEK|33|29|Then they will know that I am the LORD, when I have made the land a desolation and a waste because of all their abominations that they have committed.
EZEK|33|30|"As for you, son of man, your people who talk together about you by the walls and at the doors of the houses, say to one another, each to his brother, 'Come, and hear what the word is that comes from the LORD.'
EZEK|33|31|And they come to you as people come, and they sit before you as my people, and they hear what you say but they will not do it; for with lustful talk in their mouths they act; their heart is set on their gain.
EZEK|33|32|And behold, you are to them like one who sings lustful songs with a beautiful voice and plays well on an instrument, for they hear what you say, but they will not do it.
EZEK|33|33|When this comes- and come it will!- then they will know that a prophet has been among them."
EZEK|34|1|The word of the LORD came to me:
EZEK|34|2|"Son of man, prophesy against the shepherds of Israel; prophesy, and say to them, even to the shepherds, Thus says the Lord GOD: Ah, shepherds of Israel who have been feeding yourselves! Should not shepherds feed the sheep?
EZEK|34|3|You eat the fat, you clothe yourselves with the wool, you slaughter the fat ones, but you do not feed the sheep.
EZEK|34|4|The weak you have not strengthened, the sick you have not healed, the injured you have not bound up, the strayed you have not brought back, the lost you have not sought, and with force and harshness you have ruled them.
EZEK|34|5|So they were scattered, because there was no shepherd, and they became food for all the wild beasts.
EZEK|34|6|My sheep were scattered; they wandered over all the mountains and on every high hill. My sheep were scattered over all the face of the earth, with none to search or seek for them.
EZEK|34|7|"Therefore, you shepherds, hear the word of the LORD:
EZEK|34|8|As I live, declares the Lord GOD, surely because my sheep have become a prey, and my sheep have become food for all the wild beasts, since there was no shepherd, and because my shepherds have not searched for my sheep, but the shepherds have fed themselves, and have not fed my sheep,
EZEK|34|9|therefore, you shepherds, hear the word of the LORD:
EZEK|34|10|Thus says the Lord GOD, Behold, I am against the shepherds, and I will require my sheep at their hand and put a stop to their feeding the sheep. No longer shall the shepherds feed themselves. I will rescue my sheep from their mouths, that they may not be food for them.
EZEK|34|11|"For thus says the Lord GOD: Behold, I, I myself will search for my sheep and will seek them out.
EZEK|34|12|As a shepherd seeks out his flock when he is among his sheep that have been scattered, so will I seek out my sheep, and I will rescue them from all places where they have been scattered on a day of clouds and thick darkness.
EZEK|34|13|And I will bring them out from the peoples and gather them from the countries, and will bring them into their own land. And I will feed them on the mountains of Israel, by the ravines, and in all the inhabited places of the country.
EZEK|34|14|I will feed them with good pasture, and on the mountain heights of Israel shall be their grazing land. There they shall lie down in good grazing land, and on rich pasture they shall feed on the mountains of Israel.
EZEK|34|15|I myself will be the shepherd of my sheep, and I myself will make them lie down, declares the Lord GOD.
EZEK|34|16|I will seek the lost, and I will bring back the strayed, and I will bind up the injured, and I will strengthen the weak, and the fat and the strong I will destroy. I will feed them in justice.
EZEK|34|17|"As for you, my flock, thus says the Lord GOD: Behold, I judge between sheep and sheep, between rams and male goats.
EZEK|34|18|Is it not enough for you to feed on the good pasture, that you must tread down with your feet the rest of your pasture; and to drink of clear water, that you must muddy the rest of the water with your feet?
EZEK|34|19|And must my sheep eat what you have trodden with your feet, and drink what you have muddied with your feet?
EZEK|34|20|"Therefore, thus says the Lord GOD to them: Behold, I, I myself will judge between the fat sheep and the lean sheep.
EZEK|34|21|Because you push with side and shoulder, and thrust at all the weak with your horns, till you have scattered them abroad,
EZEK|34|22|I will rescue my flock; they shall no longer be a prey. And I will judge between sheep and sheep.
EZEK|34|23|And I will set up over them one shepherd, my servant David, and he shall feed them: he shall feed them and be their shepherd.
EZEK|34|24|And I, the LORD, will be their God, and my servant David shall be prince among them. I am the LORD; I have spoken.
EZEK|34|25|"I will make with them a covenant of peace and banish wild beasts from the land, so that they may dwell securely in the wilderness and sleep in the woods.
EZEK|34|26|And I will make them and the places all around my hill a blessing, and I will send down the showers in their season; they shall be showers of blessing.
EZEK|34|27|And the trees of the field shall yield their fruit, and the earth shall yield its increase, and they shall be secure in their land. And they shall know that I am the LORD, when I break the bars of their yoke, and deliver them from the hand of those who enslaved them.
EZEK|34|28|They shall no more be a prey to the nations, nor shall the beasts of the land devour them. They shall dwell securely, and none shall make them afraid.
EZEK|34|29|And I will provide for them renowned plantations so that they shall no more be consumed with hunger in the land, and no longer suffer the reproach of the nations.
EZEK|34|30|And they shall know that I am the LORD their God with them, and that they, the house of Israel, are my people, declares the Lord GOD.
EZEK|34|31|And you are my sheep, human sheep of my pasture, and I am your God, declares the Lord GOD."
EZEK|35|1|The word of the LORD came to me:
EZEK|35|2|"Son of man, set your face against Mount Seir, and prophesy against it,
EZEK|35|3|and say to it, Thus says the Lord GOD: Behold, I am against you, Mount Seir, and I will stretch out my hand against you, and I will make you a desolation and a waste.
EZEK|35|4|I will lay your cities waste, and you shall become a desolation, and you shall know that I am the LORD.
EZEK|35|5|Because you cherished perpetual enmity and gave over the people of Israel to the power of the sword at the time of their calamity, at the time of their final punishment,
EZEK|35|6|therefore, as I live, declares the Lord GOD, I will prepare you for blood, and blood shall pursue you; because you did not hate bloodshed, therefore blood shall pursue you.
EZEK|35|7|I will make Mount Seir a waste and a desolation, and I will cut off from it all who come and go.
EZEK|35|8|And I will fill its mountains with the slain. On your hills and in your valleys and in all your ravines those slain with the sword shall fall.
EZEK|35|9|I will make you a perpetual desolation, and your cities shall not be inhabited. Then you will know that I am the LORD.
EZEK|35|10|"Because you said, 'These two nations and these two countries shall be mine, and we will take possession of them'- although the LORD was there-
EZEK|35|11|therefore, as I live, declares the Lord GOD, I will deal with you according to the anger and envy that you showed because of your hatred against them. And I will make myself known among them, when I judge you.
EZEK|35|12|And you shall know that I am the LORD. "I have heard all the revilings that you uttered against the mountains of Israel, saying, 'They are laid desolate; they are given us to devour.'
EZEK|35|13|And you magnified yourselves against me with your mouth, and multiplied your words against me; I heard it.
EZEK|35|14|Thus says the Lord GOD: While the whole earth rejoices, I will make you desolate.
EZEK|35|15|As you rejoiced over the inheritance of the house of Israel, because it was desolate, so I will deal with you; you shall be desolate, Mount Seir, and all Edom, all of it. Then they will know that I am the LORD.
EZEK|36|1|"And you, son of man, prophesy to the mountains of Israel, and say, O mountains of Israel, hear the word of the LORD.
EZEK|36|2|Thus says the Lord GOD: Because the enemy said of you, 'Aha!' and, 'The ancient heights have become our possession,'
EZEK|36|3|therefore prophesy, and say, Thus says the Lord GOD: Precisely because they made you desolate and crushed you from all sides, so that you became the possession of the rest of the nations, and you became the talk and evil gossip of the people,
EZEK|36|4|therefore, O mountains of Israel, hear the word of the Lord GOD: Thus says the Lord GOD to the mountains and the hills, the ravines and the valleys, the desolate wastes and the deserted cities, which have become a prey and derision to the rest of the nations all around,
EZEK|36|5|therefore thus says the Lord GOD: Surely I have spoken in my hot jealousy against the rest of the nations and against all Edom, who gave my land to themselves as a possession with wholehearted joy and utter contempt, that they might make its pasturelands a prey.
EZEK|36|6|Therefore prophesy concerning the land of Israel, and say to the mountains and hills, to the ravines and valleys, Thus says the Lord GOD: Behold, I have spoken in my jealous wrath, because you have suffered the reproach of the nations.
EZEK|36|7|Therefore thus says the Lord GOD: I swear that the nations that are all around you shall themselves suffer reproach.
EZEK|36|8|"But you, O mountains of Israel, shall shoot forth your branches and yield your fruit to my people Israel, for they will soon come home.
EZEK|36|9|For behold, I am for you, and I will turn to you, and you shall be tilled and sown.
EZEK|36|10|And I will multiply people on you, the whole house of Israel, all of it. The cities shall be inhabited and the waste places rebuilt.
EZEK|36|11|And I will multiply on you man and beast, and they shall multiply and be fruitful. And I will cause you to be inhabited as in your former times, and will do more good to you than ever before. Then you will know that I am the LORD.
EZEK|36|12|I will let people walk on you, even my people Israel. And they shall possess you, and you shall be their inheritance, and you shall no longer bereave them of children.
EZEK|36|13|Thus says the Lord GOD: Because they say to you, 'You devour people, and you bereave your nation of children,'
EZEK|36|14|therefore you shall no longer devour people and no longer bereave your nation of children, declares the Lord GOD.
EZEK|36|15|And I will not let you hear anymore the reproach of the nations, and you shall no longer bear the disgrace of the peoples and no longer cause your nation to stumble, declares the Lord GOD."
EZEK|36|16|The word of the LORD came to me:
EZEK|36|17|"Son of man, when the house of Israel lived in their own land, they defiled it by their ways and their deeds. Their ways before me were like the uncleanness of a woman in her menstrual impurity.
EZEK|36|18|So I poured out my wrath upon them for the blood that they had shed in the land, for the idols with which they had defiled it.
EZEK|36|19|I scattered them among the nations, and they were dispersed through the countries. In accordance with their ways and their deeds I judged them.
EZEK|36|20|But when they came to the nations, wherever they came, they profaned my holy name, in that people said of them, 'These are the people of the LORD, and yet they had to go out of his land.'
EZEK|36|21|But I had concern for my holy name, which the house of Israel had profaned among the nations to which they came.
EZEK|36|22|"Therefore say to the house of Israel, Thus says the Lord GOD: It is not for your sake, O house of Israel, that I am about to act, but for the sake of my holy name, which you have profaned among the nations to which you came.
EZEK|36|23|And I will vindicate the holiness of my great name, which has been profaned among the nations, and which you have profaned among them. And the nations will know that I am the LORD, declares the Lord GOD, when through you I vindicate my holiness before their eyes.
EZEK|36|24|I will take you from the nations and gather you from all the countries and bring you into your own land.
EZEK|36|25|I will sprinkle clean water on you, and you shall be clean from all your uncleannesses, and from all your idols I will cleanse you.
EZEK|36|26|And I will give you a new heart, and a new spirit I will put within you. And I will remove the heart of stone from your flesh and give you a heart of flesh.
EZEK|36|27|And I will put my Spirit within you, and cause you to walk in my statutes and be careful to obey my rules.
EZEK|36|28|You shall dwell in the land that I gave to your fathers, and you shall be my people, and I will be your God.
EZEK|36|29|And I will deliver you from all your uncleannesses. And I will summon the grain and make it abundant and lay no famine upon you.
EZEK|36|30|I will make the fruit of the tree and the increase of the field abundant, that you may never again suffer the disgrace of famine among the nations.
EZEK|36|31|Then you will remember your evil ways, and your deeds that were not good, and you will loathe yourselves for your iniquities and your abominations.
EZEK|36|32|It is not for your sake that I will act, declares the Lord GOD; let that be known to you. Be ashamed and confounded for your ways, O house of Israel.
EZEK|36|33|"Thus says the Lord GOD: On the day that I cleanse you from all your iniquities, I will cause the cities to be inhabited, and the waste places shall be rebuilt.
EZEK|36|34|And the land that was desolate shall be tilled, instead of being the desolation that it was in the sight of all who passed by.
EZEK|36|35|And they will say, 'This land that was desolate has become like the garden of Eden, and the waste and desolate and ruined cities are now fortified and inhabited.'
EZEK|36|36|Then the nations that are left all around you shall know that I am the LORD; I have rebuilt the ruined places and replanted that which was desolate. I am the LORD; I have spoken, and I will do it.
EZEK|36|37|"Thus says the Lord GOD: This also I will let the house of Israel ask me to do for them: to increase their people like a flock.
EZEK|36|38|Like the flock for sacrifices, like the flock at Jerusalem during her appointed feasts, so shall the waste cities be filled with flocks of people. Then they will know that I am the LORD."
EZEK|37|1|The hand of the LORD was upon me, and he brought me out in the Spirit of the LORD and set me down in the middle of the valley; it was full of bones.
EZEK|37|2|And he led me around among them, and behold, there were very many on the surface of the valley, and behold, they were very dry.
EZEK|37|3|And he said to me, "Son of man, can these bones live?" And I answered, "O Lord GOD, you know."
EZEK|37|4|Then he said to me, "Prophesy over these bones, and say to them, O dry bones, hear the word of the LORD.
EZEK|37|5|Thus says the Lord GOD to these bones: Behold, I will cause breath to enter you, and you shall live.
EZEK|37|6|And I will lay sinews upon you, and will cause flesh to come upon you, and cover you with skin, and put breath in you, and you shall live, and you shall know that I am the LORD."
EZEK|37|7|So I prophesied as I was commanded. And as I prophesied, there was a sound, and behold, a rattling, and the bones came together, bone to its bone.
EZEK|37|8|And I looked, and behold, there were sinews on them, and flesh had come upon them, and skin had covered them. But there was no breath in them.
EZEK|37|9|Then he said to me, "Prophesy to the breath; prophesy, son of man, and say to the breath, Thus says the Lord GOD: Come from the four winds, O breath, and breathe on these slain, that they may live."
EZEK|37|10|So I prophesied as he commanded me, and the breath came into them, and they lived and stood on their feet, an exceedingly great army.
EZEK|37|11|Then he said to me, "Son of man, these bones are the whole house of Israel. Behold, they say, 'Our bones are dried up, and our hope is lost; we are clean cut off.'
EZEK|37|12|Therefore prophesy, and say to them, Thus says the Lord GOD: Behold, I will open your graves and raise you from your graves, O my people. And I will bring you into the land of Israel.
EZEK|37|13|And you shall know that I am the LORD, when I open your graves, and raise you from your graves, O my people.
EZEK|37|14|And I will put my Spirit within you, and you shall live, and I will place you in your own land. Then you shall know that I am the LORD; I have spoken, and I will do it, declares the LORD."
EZEK|37|15|The word of the LORD came to me:
EZEK|37|16|"Son of man, take a stick and write on it, 'For Judah, and the people of Israel associated with him'; then take another stick and write on it, 'For Joseph (the stick of Ephraim) and all the house of Israel associated with him.'
EZEK|37|17|And join them one to another into one stick, that they may become one in your hand.
EZEK|37|18|And when your people say to you, 'Will you not tell us what you mean by these?'
EZEK|37|19|say to them, Thus says the Lord GOD: Behold, I am about to take the stick of Joseph (that is in the hand of Ephraim) and the tribes of Israel associated with him. And I will join with it the stick of Judah, and make them one stick, that they may be one in my hand.
EZEK|37|20|When the sticks on which you write are in your hand before their eyes,
EZEK|37|21|then say to them, Thus says the Lord GOD: Behold, I will take the people of Israel from the nations among which they have gone, and will gather them from all around, and bring them to their own land.
EZEK|37|22|And I will make them one nation in the land, on the mountains of Israel. And one king shall be king over them all, and they shall be no longer two nations, and no longer divided into two kingdoms.
EZEK|37|23|They shall not defile themselves anymore with their idols and their detestable things, or with any of their transgressions. But I will save them from all the backslidings in which they have sinned, and will cleanse them; and they shall be my people, and I will be their God.
EZEK|37|24|"My servant David shall be king over them, and they shall all have one shepherd. They shall walk in my rules and be careful to obey my statutes.
EZEK|37|25|They shall dwell in the land that I gave to my servant Jacob, where your fathers lived. They and their children and their children's children shall dwell there forever, and David my servant shall be their prince forever.
EZEK|37|26|I will make a covenant of peace with them. It shall be an everlasting covenant with them. And I will set them in their land and multiply them, and will set my sanctuary in their midst forevermore.
EZEK|37|27|My dwelling place shall be with them, and I will be their God, and they shall be my people.
EZEK|37|28|Then the nations will know that I am the LORD who sanctifies Israel, when my sanctuary is in their midst forevermore."
EZEK|38|1|The word of the LORD came to me:
EZEK|38|2|"Son of man, set your face toward Gog, of the land of Magog, the chief prince of Meshech and Tubal, and prophesy against him
EZEK|38|3|and say, Thus says the Lord GOD: Behold, I am against you, O Gog, chief prince of Meshech and Tubal.
EZEK|38|4|And I will turn you about and put hooks into your jaws, and I will bring you out, and all your army, horses and horsemen, all of them clothed in full armor, a great host, all of them with buckler and shield, wielding swords.
EZEK|38|5|Persia, Cush, and Put are with them, all of them with shield and helmet;
EZEK|38|6|Gomer and all his hordes; Beth-togarmah from the uttermost parts of the north with all his hordes- many peoples are with you.
EZEK|38|7|"Be ready and keep ready, you and all your hosts that are assembled about you, and be a guard for them.
EZEK|38|8|After many days you will be mustered. In the latter years you will go against the land that is restored from war, the land whose people were gathered from many peoples upon the mountains of Israel, which had been a continual waste. Its people were brought out from the peoples and now dwell securely, all of them.
EZEK|38|9|You will advance, coming on like a storm. You will be like a cloud covering the land, you and all your hordes, and many peoples with you.
EZEK|38|10|"Thus says the Lord GOD: On that day, thoughts will come into your mind, and you will devise an evil scheme
EZEK|38|11|and say, 'I will go up against the land of unwalled villages. I will fall upon the quiet people who dwell securely, all of them dwelling without walls, and having no bars or gates,'
EZEK|38|12|to seize spoil and carry off plunder, to turn your hand against the waste places that are now inhabited, and the people who were gathered from the nations, who have acquired livestock and goods, who dwell at the center of the earth.
EZEK|38|13|Sheba and Dedan and the merchants of Tarshish and all its leaders will say to you, 'Have you come to seize spoil? Have you assembled your hosts to carry off plunder, to carry away silver and gold, to take away livestock and goods, to seize great spoil?'
EZEK|38|14|"Therefore, son of man, prophesy, and say to Gog, Thus says the Lord GOD: On that day when my people Israel are dwelling securely, will you not know it?
EZEK|38|15|You will come from your place out of the uttermost parts of the north, you and many peoples with you, all of them riding on horses, a great host, a mighty army.
EZEK|38|16|You will come up against my people Israel, like a cloud covering the land. In the latter days I will bring you against my land, that the nations may know me, when through you, O Gog, I vindicate my holiness before their eyes.
EZEK|38|17|"Thus says the Lord GOD: Are you he of whom I spoke in former days by my servants the prophets of Israel, who in those days prophesied for years that I would bring you against them?
EZEK|38|18|But on that day, the day that Gog shall come against the land of Israel, declares the Lord GOD, my wrath will be roused in my anger.
EZEK|38|19|For in my jealousy and in my blazing wrath I declare, On that day there shall be a great earthquake in the land of Israel.
EZEK|38|20|The fish of the sea and the birds of the heavens and the beasts of the field and all creeping things that creep on the ground, and all the people who are on the face of the earth, shall quake at my presence. And the mountains shall be thrown down, and the cliffs shall fall, and every wall shall tumble to the ground.
EZEK|38|21|I will summon a sword against Gog on all my mountains, declares the Lord GOD. Every man's sword will be against his brother.
EZEK|38|22|With pestilence and bloodshed I will enter into judgment with him, and I will rain upon him and his hordes and the many peoples who are with him torrential rains and hailstones, fire and sulfur.
EZEK|38|23|So I will show my greatness and my holiness and make myself known in the eyes of many nations. Then they will know that I am the LORD.
EZEK|39|1|"And you, son of man, prophesy against Gog and say, Thus says the Lord GOD: Behold, I am against you, O Gog, chief prince of Meshech and Tubal.
EZEK|39|2|And I will turn you about and drive you forward, and bring you up from the uttermost parts of the north, and lead you against the mountains of Israel.
EZEK|39|3|Then I will strike your bow from your left hand, and will make your arrows drop out of your right hand.
EZEK|39|4|You shall fall on the mountains of Israel, you and all your hordes and the peoples who are with you. I will give you to birds of prey of every sort and to the beasts of the field to be devoured.
EZEK|39|5|You shall fall in the open field, for I have spoken, declares the Lord GOD.
EZEK|39|6|I will send fire on Magog and on those who dwell securely in the coastlands, and they shall know that I am the LORD.
EZEK|39|7|"And my holy name I will make known in the midst of my people Israel, and I will not let my holy name be profaned anymore. And the nations shall know that I am the LORD, the Holy One in Israel.
EZEK|39|8|Behold, it is coming and it will be brought about, declares the Lord GOD. That is the day of which I have spoken.
EZEK|39|9|"Then those who dwell in the cities of Israel will go out and make fires of the weapons and burn them, shields and bucklers, bow and arrows, clubs and spears; and they will make fires of them for seven years,
EZEK|39|10|so that they will not need to take wood out of the field or cut down any out of the forests, for they will make their fires of the weapons. They will seize the spoil of those who despoiled them, and plunder those who plundered them, declares the Lord GOD.
EZEK|39|11|"On that day I will give to Gog a place for burial in Israel, the Valley of the Travelers, east of the sea. It will block the travelers, for there Gog and all his multitude will be buried. It will be called the Valley of Hamon-gog.
EZEK|39|12|For seven months the house of Israel will be burying them, in order to cleanse the land.
EZEK|39|13|All the people of the land will bury them, and it will bring them renown on the day that I show my glory, declares the Lord GOD.
EZEK|39|14|They will set apart men to travel through the land regularly and bury those travelers remaining on the face of the land, so as to cleanse it. At the end of seven months they will make their search.
EZEK|39|15|And when these travel through the land and anyone sees a human bone, then he shall set up a sign by it, till the buriers have buried it in the Valley of Hamon-gog.
EZEK|39|16|(Hamonah is also the name of the city.) Thus shall they cleanse the land.
EZEK|39|17|"As for you, son of man, thus says the Lord GOD: Speak to the birds of every sort and to all beasts of the field, 'Assemble and come, gather from all around to the sacrificial feast that I am preparing for you, a great sacrificial feast on the mountains of Israel, and you shall eat flesh and drink blood.
EZEK|39|18|You shall eat the flesh of the mighty, and drink the blood of the princes of the earth- of rams, of lambs, and of he-goats, of bulls, all of them fat beasts of Bashan.
EZEK|39|19|And you shall eat fat till you are filled, and drink blood till you are drunk, at the sacrificial feast that I am preparing for you.
EZEK|39|20|And you shall be filled at my table with horses and charioteers, with mighty men and all kinds of warriors,' declares the Lord GOD.
EZEK|39|21|"And I will set my glory among the nations, and all the nations shall see my judgment that I have executed, and my hand that I have laid on them.
EZEK|39|22|The house of Israel shall know that I am the LORD their God, from that day forward.
EZEK|39|23|And the nations shall know that the house of Israel went into captivity for their iniquity, because they dealt so treacherously with me that I hid my face from them and gave them into the hand of their adversaries, and they all fell by the sword.
EZEK|39|24|I dealt with them according to their uncleanness and their transgressions, and hid my face from them.
EZEK|39|25|"Therefore thus says the Lord GOD: Now I will restore the fortunes of Jacob and have mercy on the whole house of Israel, and I will be jealous for my holy name.
EZEK|39|26|They shall forget their shame and all the treachery they have practiced against me, when they dwell securely in their land with none to make them afraid,
EZEK|39|27|when I have brought them back from the peoples and gathered them from their enemies' lands, and through them have vindicated my holiness in the sight of many nations.
EZEK|39|28|Then they shall know that I am the LORD their God, because I sent them into exile among the nations and then assembled them into their own land. I will leave none of them remaining among the nations anymore.
EZEK|39|29|And I will not hide my face anymore from them, when I pour out my Spirit upon the house of Israel, declares the Lord GOD."
EZEK|40|1|In the twenty-fifth year of our exile, at the beginning of the year, on the tenth day of the month, in the fourteenth year after the city was struck down, on that very day, the hand of the LORD was upon me, and he brought me to the city.
EZEK|40|2|In visions of God he brought me to the land of Israel, and set me down on a very high mountain, on which was a structure like a city to the south.
EZEK|40|3|When he brought me there, behold, there was a man whose appearance was like bronze, with a linen cord and a measuring reed in his hand. And he was standing in the gateway.
EZEK|40|4|And the man said to me, "Son of man, look with your eyes, and hear with your ears, and set your heart upon all that I shall show you, for you were brought here in order that I might show it to you. Declare all that you see to the house of Israel."
EZEK|40|5|And behold, there was a wall all around the outside of the temple area, and the length of the measuring reed in the man's hand was six long cubits, each being a cubit and a handbreadth in length. So he measured the thickness of the wall, one reed; and the height, one reed.
EZEK|40|6|Then he went into the gateway facing east, going up its steps, and measured the threshold of the gate, one reed deep.
EZEK|40|7|And the side rooms, one reed long and one reed broad; and the space between the side rooms, five cubits; and the threshold of the gate by the vestibule of the gate at the inner end, one reed.
EZEK|40|8|Then he measured the vestibule of the gateway, on the inside, one reed.
EZEK|40|9|Then he measured the vestibule of the gateway, eight cubits; and its jambs, two cubits; and the vestibule of the gate was at the inner end.
EZEK|40|10|And there were three side rooms on either side of the east gate. The three were of the same size, and the jambs on either side were of the same size.
EZEK|40|11|Then he measured the width of the opening of the gateway, ten cubits; and the length of the gateway, thirteen cubits.
EZEK|40|12|There was a barrier before the side rooms, one cubit on either side. And the side rooms were six cubits on either side.
EZEK|40|13|Then he measured the gate from the ceiling of the one side room to the ceiling of the other, a breadth of twenty-five cubits; the openings faced each other.
EZEK|40|14|He measured also the vestibule, twenty cubits. And around the vestibule of the gateway was the court.
EZEK|40|15|From the front of the gate at the entrance to the front of the inner vestibule of the gate was fifty cubits.
EZEK|40|16|And the gateway had windows all around, narrowing inwards toward the side rooms and toward their jambs, and likewise the vestibule had windows all around inside, and on the jambs were palm trees.
EZEK|40|17|Then he brought me into the outer court. And behold, there were chambers and a pavement, all around the court. Thirty chambers faced the pavement.
EZEK|40|18|And the pavement ran along the side of the gates, corresponding to the length of the gates. This was the lower pavement.
EZEK|40|19|Then he measured the distance from the inner front of the lower gate to the outer front of the inner court, a hundred cubits on the east side and on the north side.
EZEK|40|20|As for the gate that faced toward the north, belonging to the outer court, he measured its length and its breadth.
EZEK|40|21|Its side rooms, three on either side, and its jambs and its vestibule were of the same size as those of the first gate. Its length was fifty cubits, and its breadth twenty-five cubits.
EZEK|40|22|And its windows, its vestibule, and its palm trees were of the same size as those of the gate that faced toward the east. And by seven steps people would go up to it, and find its vestibule before them.
EZEK|40|23|And opposite the gate on the north, as on the east, was a gate to the inner court. And he measured from gate to gate, a hundred cubits.
EZEK|40|24|And he led me toward the south, and behold, there was a gate on the south. And he measured its jambs and its vestibule; they had the same size as the others.
EZEK|40|25|Both it and its vestibule had windows all around, like the windows of the others. Its length was fifty cubits, and its breadth twenty-five cubits.
EZEK|40|26|And there were seven steps leading up to it, and its vestibule was before them, and it had palm trees on its jambs, one on either side.
EZEK|40|27|And there was a gate on the south of the inner court. And he measured from gate to gate toward the south, a hundred cubits.
EZEK|40|28|Then he brought me to the inner court through the south gate, and he measured the south gate. It was of the same size as the others.
EZEK|40|29|Its side rooms, its jambs, and its vestibule were of the same size as the others, and both it and its vestibule had windows all around. Its length was fifty cubits, and its breadth twenty-five cubits.
EZEK|40|30|And there were vestibules all around, twenty-five cubits long and five cubits broad.
EZEK|40|31|Its vestibule faced the outer court, and palm trees were on its jambs, and its stairway had eight steps.
EZEK|40|32|Then he brought me to the inner court on the east side, and he measured the gate. It was of the same size as the others.
EZEK|40|33|Its side rooms, its jambs, and its vestibule were of the same size as the others, and both it and its vestibule had windows all around. Its length was fifty cubits, and its breadth twenty-five cubits.
EZEK|40|34|Its vestibule faced the outer court, and it had palm trees on its jambs, on either side, and its stairway had eight steps.
EZEK|40|35|Then he brought me to the north gate, and he measured it. It had the same size as the others.
EZEK|40|36|Its side rooms, its jambs, and its vestibule were of the same size as the others, and it had windows all around. Its length was fifty cubits, and its breadth twenty-five cubits.
EZEK|40|37|Its vestibule faced the outer court, and it had palm trees on its jambs, on either side, and its stairway had eight steps.
EZEK|40|38|There was a chamber with its door in the vestibule of the gate, where the burnt offering was to be washed.
EZEK|40|39|And in the vestibule of the gate were two tables on either side, on which the burnt offering and the sin offering and the guilt offering were to be slaughtered.
EZEK|40|40|And off to the side, on the outside as one goes up to the entrance of the north gate, were two tables; and off to the other side of the vestibule of the gate were two tables.
EZEK|40|41|Four tables were on either side of the gate, eight tables, on which to slaughter.
EZEK|40|42|And there were four tables of hewn stone for the burnt offering, a cubit and a half long, and a cubit and a half broad, and one cubit high, on which the instruments were to be laid with which the burnt offerings and the sacrifices were slaughtered.
EZEK|40|43|And hooks, a handbreadth long, were fastened all around within. And on the tables the flesh of the offering was to be laid.
EZEK|40|44|On the outside of the inner gateway there were two chambers in the inner court, one at the side of the north gate facing south, the other at the side of the south gate facing north.
EZEK|40|45|And he said to me, This chamber that faces south is for the priests who have charge of the temple,
EZEK|40|46|and the chamber that faces north is for the priests who have charge of the altar. These are the sons of Zadok, who alone among the sons of Levi may come near to the LORD to minister to him.
EZEK|40|47|And he measured the court, a hundred cubits long and a hundred cubits broad, a square. And the altar was in front of the temple.
EZEK|40|48|Then he brought me to the vestibule of the temple and measured the jambs of the vestibule, five cubits on either side. And the breadth of the gate was fourteen cubits, and the sidewalls of the gate were three cubits on either side.
EZEK|40|49|The length of the vestibule was twenty cubits, and the breadth twelve cubits, and people would go up to it by ten steps. And there were pillars beside the jambs, one on either side.
EZEK|41|1|Then he brought me to the nave and measured the jambs. On each side six cubits was the breadth of the jambs.
EZEK|41|2|And the breadth of the entrance was ten cubits, and the sidewalls of the entrance were five cubits on either side. And he measured the length of the nave, forty cubits, and its breadth, twenty cubits.
EZEK|41|3|Then he went into the inner room and measured the jambs of the entrance, two cubits; and the entrance, six cubits; and the sidewalls on either side of the entrance, seven cubits.
EZEK|41|4|And he measured the length of the room, twenty cubits, and its breadth, twenty cubits, across the nave. And he said to me, "This is the Most Holy Place."
EZEK|41|5|Then he measured the wall of the temple, six cubits thick, and the breadth of the side chambers, four cubits, all around the temple.
EZEK|41|6|And the side chambers were in three stories, one over another, thirty in each story. There were offsets all around the wall of the temple to serve as supports for the side chambers, so that they should not be supported by the wall of the temple.
EZEK|41|7|And it became broader as it wound upward to the side chambers, because the temple was enclosed upward all around the temple. Thus the temple had a broad area upwards, and so one went up from the lowest story to the top story through the middle story.
EZEK|41|8|I saw also that the temple had a raised platform all around; the foundations of the side chambers measured a full reed of six long cubits.
EZEK|41|9|The thickness of the outer wall of the side chambers was five cubits. The free space between the side chambers of the temple and the
EZEK|41|10|other chambers was a breadth of twenty cubits all around the temple on every side.
EZEK|41|11|And the doors of the side chambers opened on the free space, one door toward the north, and another door toward the south. And the breadth of the free space was five cubits all around.
EZEK|41|12|The building that was facing the separate yard on the west side was seventy cubits broad, and the wall of the building was five cubits thick all around, and its length ninety cubits.
EZEK|41|13|Then he measured the temple, a hundred cubits long; and the yard and the building with its walls, a hundred cubits long;
EZEK|41|14|also the breadth of the east front of the temple and the yard, a hundred cubits.
EZEK|41|15|Then he measured the length of the building facing the yard that was at the back and its galleries on either side, a hundred cubits. The inside of the nave and the vestibules of the court,
EZEK|41|16|the thresholds and the narrow windows and the galleries all around the three of them, opposite the threshold, were paneled with wood all around, from the floor up to the windows (now the windows were covered),
EZEK|41|17|to the space above the door, even to the inner room, and on the outside. And on all the walls all around, inside and outside, was a measured pattern.
EZEK|41|18|It was carved of cherubim and palm trees, a palm tree between cherub and cherub. Every cherub had two faces:
EZEK|41|19|a human face toward the palm tree on the one side, and the face of a young lion toward the palm tree on the other side. They were carved on the whole temple all around.
EZEK|41|20|From the floor to above the door, cherubim and palm trees were carved; similarly the wall of the nave.
EZEK|41|21|The doorposts of the nave were squared, and in front of the Holy Place was something resembling
EZEK|41|22|an altar of wood, three cubits high, two cubits long, and two cubits broad. Its corners, its base, and its walls were of wood. He said to me, "This is the table that is before the LORD."
EZEK|41|23|The nave and the Holy Place had each a double door.
EZEK|41|24|The double doors had two leaves apiece, two swinging leaves for each door.
EZEK|41|25|And on the doors of the nave were carved cherubim and palm trees, such as were carved on the walls. And there was a canopy of wood in front of the vestibule outside.
EZEK|41|26|And there were narrow windows and palm trees on either side, on the sidewalls of the vestibule, the side chambers of the temple, and the canopies.
EZEK|42|1|Then he led me out into the outer court, toward the north, and he brought me to the chambers that were opposite the separate yard and opposite the building on the north.
EZEK|42|2|The length of the building whose door faced north was a hundred cubits, and the breadth fifty cubits.
EZEK|42|3|Facing the twenty cubits that belonged to the inner court, and facing the pavement that belonged to the outer court, was gallery against gallery in three stories.
EZEK|42|4|And before the chambers was a passage inward, ten cubits wide and a hundred cubits long, and their doors were on the north.
EZEK|42|5|Now the upper chambers were narrower, for the galleries took more away from them than from the lower and middle chambers of the building.
EZEK|42|6|For they were in three stories, and they had no pillars like the pillars of the courts. Thus the upper chambers were set back from the ground more than the lower and the middle ones.
EZEK|42|7|And there was a wall outside parallel to the chambers, toward the outer court, opposite the chambers, fifty cubits long.
EZEK|42|8|For the chambers on the outer court were fifty cubits long, while those opposite the nave were a hundred cubits long.
EZEK|42|9|Below these chambers was an entrance on the east side, as one enters them from the outer court.
EZEK|42|10|In the thickness of the wall of the court, on the south also, opposite the yard and opposite the building, there were chambers
EZEK|42|11|with a passage in front of them. They were similar to the chambers on the north, of the same length and breadth, with the same exits and arrangements and doors,
EZEK|42|12|as were the entrances of the chambers on the south. There was an entrance at the beginning of the passage, the passage before the corresponding wall on the east as one enters them.
EZEK|42|13|Then he said to me, "The north chambers and the south chambers opposite the yard are the holy chambers, where the priests who approach the LORD shall eat the most holy offerings. There they shall put the most holy offerings- the grain offering, the sin offering, and the guilt offering, for the place is holy.
EZEK|42|14|When the priests enter the Holy Place, they shall not go out of it into the outer court without laying there the garments in which they minister, for these are holy. They shall put on other garments before they go near to that which is for the people."
EZEK|42|15|Now when he had finished measuring the interior of the temple area, he led me out by the gate that faced east, and measured the temple area all around.
EZEK|42|16|He measured the east side with the measuring reed, 500 cubits by the measuring reed all around.
EZEK|42|17|He measured the north side, 500 cubits by the measuring reed all around.
EZEK|42|18|He measured the south side, 500 cubits by the measuring reed.
EZEK|42|19|Then he turned to the west side and measured, 500 cubits by the measuring reed.
EZEK|42|20|He measured it on the four sides. It had a wall around it, 500 cubits long and 500 cubits broad, to make a separation between the holy and the common.
EZEK|43|1|Then he led me to the gate, the gate facing east.
EZEK|43|2|And behold, the glory of the God of Israel was coming from the east. And the sound of his coming was like the sound of many waters, and the earth shone with his glory.
EZEK|43|3|And the vision I saw was just like the vision that I had seen when he came to destroy the city, and just like the vision that I had seen by the Chebar canal. And I fell on my face.
EZEK|43|4|As the glory of the LORD entered the temple by the gate facing east,
EZEK|43|5|the Spirit lifted me up and brought me into the inner court; and behold, the glory of the LORD filled the temple.
EZEK|43|6|While the man was standing beside me, I heard one speaking to me out of the temple,
EZEK|43|7|and he said to me, "Son of man, this is the place of my throne and the place of the soles of my feet, where I will dwell in the midst of the people of Israel forever. And the house of Israel shall no more defile my holy name, neither they, nor their kings, by their whoring and by the dead bodies of their kings at their high places,
EZEK|43|8|by setting their threshold by my threshold and their doorposts beside my doorposts, with only a wall between me and them. They have defiled my holy name by their abominations that they have committed, so I have consumed them in my anger.
EZEK|43|9|Now let them put away their whoring and the dead bodies of their kings far from me, and I will dwell in their midst forever.
EZEK|43|10|"As for you, son of man, describe to the house of Israel the temple, that they may be ashamed of their iniquities; and they shall measure the plan.
EZEK|43|11|And if they are ashamed of all that they have done, make known to them the design of the temple, its arrangement, its exits and its entrances, that is, its whole design; and make known to them as well all its statutes and its whole design and all its laws, and write it down in their sight, so that they may observe all its laws and all its statutes and carry them out.
EZEK|43|12|This is the law of the temple: the whole territory on the top of the mountain all around shall be most holy. Behold, this is the law of the temple.
EZEK|43|13|"These are the measurements of the altar by cubits (the cubit being a cubit and a handbreadth): its base shall be one cubit high and one cubit broad, with a rim of one span around its edge. And this shall be the height of the altar:
EZEK|43|14|from the base on the ground to the lower ledge, two cubits, with a breadth of one cubit; and from the smaller ledge to the larger ledge, four cubits, with a breadth of one cubit;
EZEK|43|15|and the altar hearth, four cubits; and from the altar hearth projecting upward, four horns.
EZEK|43|16|The altar hearth shall be square, twelve cubits long by twelve broad.
EZEK|43|17|The ledge also shall be square, fourteen cubits long by fourteen broad, with a rim around it half a cubit broad, and its base one cubit all around. The steps of the altar shall face east."
EZEK|43|18|And he said to me, "Son of man, thus says the Lord GOD: These are the ordinances for the altar: On the day when it is erected for offering burnt offerings upon it and for throwing blood against it,
EZEK|43|19|you shall give to the Levitical priests of the family of Zadok, who draw near to me to minister to me, declares the Lord GOD, a bull from the herd for a sin offering.
EZEK|43|20|And you shall take some of its blood and put it on the four horns of the altar and on the four corners of the ledge and upon the rim all around. Thus you shall purify the altar and make atonement for it.
EZEK|43|21|You shall also take the bull of the sin offering, and it shall be burned in the appointed place belonging to the temple, outside the sacred area.
EZEK|43|22|And on the second day you shall offer a male goat without blemish for a sin offering; and the altar shall be purified, as it was purified with the bull.
EZEK|43|23|When you have finished purifying it, you shall offer a bull from the herd without blemish and a ram from the flock without blemish.
EZEK|43|24|You shall present them before the LORD, and the priests shall sprinkle salt on them and offer them up as a burnt offering to the LORD.
EZEK|43|25|For seven days you shall provide daily a male goat for a sin offering; also, a bull from the herd and a ram from the flock, without blemish, shall be provided.
EZEK|43|26|Seven days shall they make atonement for the altar and cleanse it, and so consecrate it.
EZEK|43|27|And when they have completed these days, then from the eighth day onward the priests shall offer on the altar your burnt offerings and your peace offerings, and I will accept you, declares the Lord GOD."
EZEK|44|1|Then he brought me back to the outer gate of the sanctuary, which faces east. And it was shut.
EZEK|44|2|And the LORD said to me, "This gate shall remain shut; it shall not be opened, and no one shall enter by it, for the LORD, the God of Israel, has entered by it. Therefore it shall remain shut.
EZEK|44|3|Only the prince may sit in it to eat bread before the LORD. He shall enter by way of the vestibule of the gate, and shall go out by the same way."
EZEK|44|4|Then he brought me by way of the north gate to the front of the temple, and I looked, and behold, the glory of the LORD filled the temple of the LORD. And I fell on my face.
EZEK|44|5|And the LORD said to me, "Son of man, mark well, see with your eyes, and hear with your ears all that I shall tell you concerning all the statutes of the temple of the LORD and all its laws. And mark well the entrance to the temple and all the exits from the sanctuary.
EZEK|44|6|And say to the rebellious house, to the house of Israel, Thus says the Lord GOD: O house of Israel, enough of all your abominations,
EZEK|44|7|in admitting foreigners, uncircumcised in heart and flesh, to be in my sanctuary, profaning my temple, when you offer to me my food, the fat and the blood. You have broken my covenant, in addition to all your abominations.
EZEK|44|8|And you have not kept charge of my holy things, but you have set others to keep my charge for you in my sanctuary.
EZEK|44|9|"Thus says the Lord GOD: No foreigner, uncircumcised in heart and flesh, of all the foreigners who are among the people of Israel, shall enter my sanctuary.
EZEK|44|10|But the Levites who went far from me, going astray from me after their idols when Israel went astray, shall bear their punishment.
EZEK|44|11|They shall be ministers in my sanctuary, having oversight at the gates of the temple and ministering in the temple. They shall slaughter the burnt offering and the sacrifice for the people, and they shall stand before the people, to minister to them.
EZEK|44|12|Because they ministered to them before their idols and became a stumbling block of iniquity to the house of Israel, therefore I have sworn concerning them, declares the Lord GOD, and they shall bear their punishment.
EZEK|44|13|They shall not come near to me, to serve me as priest, nor come near any of my holy things and the things that are most holy, but they shall bear their shame and the abominations that they have committed.
EZEK|44|14|Yet I will appoint them to keep charge of the temple, to do all its service and all that is to be done in it.
EZEK|44|15|"But the Levitical priests, the sons of Zadok, who kept the charge of my sanctuary when the people of Israel went astray from me, shall come near to me to minister to me. And they shall stand before me to offer me the fat and the blood, declares the Lord GOD.
EZEK|44|16|They shall enter my sanctuary, and they shall approach my table, to minister to me, and they shall keep my charge.
EZEK|44|17|When they enter the gates of the inner court, they shall wear linen garments. They shall have nothing of wool on them, while they minister at the gates of the inner court, and within.
EZEK|44|18|They shall have linen turbans on their heads, and linen undergarments around their waists. They shall not bind themselves with anything that causes sweat.
EZEK|44|19|And when they go out into the outer court to the people, they shall put off the garments in which they have been ministering and lay them in the holy chambers. And they shall put on other garments, lest they communicate holiness to the people with their garments.
EZEK|44|20|They shall not shave their heads or let their locks grow long; they shall surely trim the hair of their heads.
EZEK|44|21|No priest shall drink wine when he enters the inner court.
EZEK|44|22|They shall not marry a widow or a divorced woman, but only virgins of the offspring of the house of Israel, or a widow who is the widow of a priest.
EZEK|44|23|They shall teach my people the difference between the holy and the common, and show them how to distinguish between the unclean and the clean.
EZEK|44|24|In a dispute, they shall act as judges, and they shall judge it according to my judgments. They shall keep my laws and my statutes in all my appointed feasts, and they shall keep my Sabbaths holy.
EZEK|44|25|They shall not defile themselves by going near to a dead person. However, for father or mother, for son or daughter, for brother or unmarried sister they may defile themselves.
EZEK|44|26|After he has become clean, they shall count seven days for him.
EZEK|44|27|And on the day that he goes into the Holy Place, into the inner court, to minister in the Holy Place, he shall offer his sin offering, declares the Lord GOD.
EZEK|44|28|"This shall be their inheritance: I am their inheritance: and you shall give them no possession in Israel; I am their possession.
EZEK|44|29|They shall eat the grain offering, the sin offering, and the guilt offering, and every devoted thing in Israel shall be theirs.
EZEK|44|30|And the first of all the firstfruits of all kinds, and every offering of all kinds from all your offerings, shall belong to the priests. You shall also give to the priests the first of your dough, that a blessing may rest on your house.
EZEK|44|31|The priests shall not eat of anything, whether bird or beast, that has died of itself or is torn by wild animals.
EZEK|45|1|"When you allot the land as an inheritance, you shall set apart for the LORD a portion of the land as a holy district, 25,000 cubits long and 20,000 cubits broad. It shall be holy throughout its whole extent.
EZEK|45|2|Of this a square plot of 500 by 500 cubits shall be for the sanctuary, with fifty cubits for an open space around it.
EZEK|45|3|And from this measured district you shall measure off a section 25,000 cubits long and 10,000 broad, in which shall be the sanctuary, the Most Holy Place.
EZEK|45|4|It shall be the holy portion of the land. It shall be for the priests, who minister in the sanctuary and approach the LORD to minister to him, and it shall be a place for their houses and a holy place for the sanctuary.
EZEK|45|5|Another section, 25,000 cubits long and 10,000 cubits broad, shall be for the Levites who minister at the temple, as their possession for cities to live in.
EZEK|45|6|"Alongside the portion set apart as the holy district you shall assign for the property of the city an area 5,000 cubits broad and 25,000 cubits long. It shall belong to the whole house of Israel.
EZEK|45|7|"And to the prince shall belong the land on both sides of the holy district and the property of the city, alongside the holy district and the property of the city, on the west and on the east, corresponding in length to one of the tribal portions, and extending from the western to the eastern boundary
EZEK|45|8|of the land. It is to be his property in Israel. And my princes shall no more oppress my people, but they shall let the house of Israel have the land according to their tribes.
EZEK|45|9|"Thus says the Lord GOD: Enough, O princes of Israel! Put away violence and oppression, and execute justice and righteousness. Cease your evictions of my people, declares the Lord GOD.
EZEK|45|10|"You shall have just balances, a just ephah, and a just bath.
EZEK|45|11|The ephah and the bath shall be of the same measure, the bath containing one tenth of a homer, and the ephah one tenth of a homer; the homer shall be the standard measure.
EZEK|45|12|The shekel shall be twenty gerahs; twenty shekels plus twenty-five shekels plus fifteen shekels shall be your mina.
EZEK|45|13|"This is the offering that you shall make: one sixth of an ephah from each homer of wheat, and one sixth of an ephah from each homer of barley,
EZEK|45|14|and as the fixed portion of oil, measured in baths, one tenth of a bath from each cor (the cor, like the homer, contains ten baths).
EZEK|45|15|And one sheep from every flock of two hundred, from the watering places of Israel for grain offering, burnt offering, and peace offerings, to make atonement for them, declares the Lord GOD.
EZEK|45|16|All the people of the land shall be obliged to give this offering to the prince in Israel.
EZEK|45|17|It shall be the prince's duty to furnish the burnt offerings, grain offerings, and drink offerings, at the feasts, the new moons, and the Sabbaths, all the appointed feasts of the house of Israel: he shall provide the sin offerings, grain offerings, burnt offerings, and peace offerings, to make atonement on behalf of the house of Israel.
EZEK|45|18|"Thus says the Lord GOD: In the first month, on the first day of the month, you shall take a bull from the herd without blemish, and purify the sanctuary.
EZEK|45|19|The priest shall take some of the blood of the sin offering and put it on the doorposts of the temple, the four corners of the ledge of the altar, and the posts of the gate of the inner court.
EZEK|45|20|You shall do the same on the seventh day of the month for anyone who has sinned through error or ignorance; so you shall make atonement for the temple.
EZEK|45|21|"In the first month, on the fourteenth day of the month, you shall celebrate the Feast of the Passover, and for seven days unleavened bread shall be eaten.
EZEK|45|22|On that day the prince shall provide for himself and all the people of the land a young bull for a sin offering.
EZEK|45|23|And on the seven days of the festival he shall provide as a burnt offering to the LORD seven young bulls and seven rams without blemish, on each of the seven days; and a male goat daily for a sin offering.
EZEK|45|24|And he shall provide as a grain offering an ephah for each bull, an ephah for each ram, and a hin of oil to each ephah.
EZEK|45|25|In the seventh month, on the fifteenth day of the month and for the seven days of the feast, he shall make the same provision for sin offerings, burnt offerings, and grain offerings, and for the oil.
EZEK|46|1|"Thus says the Lord GOD: The gate of the inner court that faces east shall be shut on the six working days, but on the Sabbath day it shall be opened, and on the day of the new moon it shall be opened.
EZEK|46|2|The prince shall enter by the vestibule of the gate from outside, and shall take his stand by the post of the gate. The priests shall offer his burnt offering and his peace offerings, and he shall worship at the threshold of the gate. Then he shall go out, but the gate shall not be shut until evening.
EZEK|46|3|The people of the land shall bow down at the entrance of that gate before the LORD on the Sabbaths and on the new moons.
EZEK|46|4|The burnt offering that the prince offers to the LORD on the Sabbath day shall be six lambs without blemish and a ram without blemish.
EZEK|46|5|And the grain offering with the ram shall be an ephah, and the grain offering with the lambs shall be as much as he is able, together with a hin of oil to each ephah.
EZEK|46|6|On the day of the new moon he shall offer a bull from the herd without blemish, and six lambs and a ram, which shall be without blemish.
EZEK|46|7|As a grain offering he shall provide an ephah with the bull and an ephah with the ram, and with the lambs as much as he is able, together with a hin of oil to each ephah.
EZEK|46|8|When the prince enters, he shall enter by the vestibule of the gate, and he shall go out by the same way.
EZEK|46|9|"When the people of the land come before the LORD at the appointed feasts, he who enters by the north gate to worship shall go out by the south gate, and he who enters by the south gate shall go out by the north gate: no one shall return by way of the gate by which he entered, but each shall go out straight ahead.
EZEK|46|10|When they enter, the prince shall enter with them, and when they go out, he shall go out.
EZEK|46|11|"At the feasts and the appointed festivals, the grain offering with a young bull shall be an ephah, and with a ram an ephah, and with the lambs as much as one is able to give, together with a hin of oil to an ephah.
EZEK|46|12|When the prince provides a freewill offering, either a burnt offering or peace offerings as a freewill offering to the LORD, the gate facing east shall be opened for him. And he shall offer his burnt offering or his peace offerings as he does on the Sabbath day. Then he shall go out, and after he has gone out the gate shall be shut.
EZEK|46|13|"You shall provide a lamb a year old without blemish for a burnt offering to the LORD daily; morning by morning you shall provide it.
EZEK|46|14|And you shall provide a grain offering with it morning by morning, one sixth of an ephah, and one third of a hin of oil to moisten the flour, as a grain offering to the LORD. This is a perpetual statute.
EZEK|46|15|Thus the lamb and the meal offering and the oil shall be provided, morning by morning, for a regular burnt offering.
EZEK|46|16|"Thus says the Lord GOD: If the prince makes a gift to any of his sons as his inheritance, it shall belong to his sons. It is their property by inheritance.
EZEK|46|17|But if he makes a gift out of his inheritance to one of his servants, it shall be his to the year of liberty. Then it shall revert to the prince; surely it is his inheritance- it shall belong to his sons.
EZEK|46|18|The prince shall not take any of the inheritance of the people, thrusting them out of their property. He shall give his sons their inheritance out of his own property, so that none of my people shall be scattered from his property."
EZEK|46|19|Then he brought me through the entrance, which was at the side of the gate, to the north row of the holy chambers for the priests, and behold, a place was there at the extreme western end of them.
EZEK|46|20|And he said to me, "This is the place where the priests shall boil the guilt offering and the sin offering, and where they shall bake the grain offering, in order not to bring them out into the outer court and so communicate holiness to the people."
EZEK|46|21|Then he brought me out to the outer court and led me around to the four corners of the court. And behold, in each corner of the court there was another court-
EZEK|46|22|in the four corners of the court were small courts, forty cubits long and thirty broad; the four were of the same size.
EZEK|46|23|On the inside, around each of the four courts was a row of masonry, with hearths made at the bottom of the rows all around.
EZEK|46|24|Then he said to me, "These are the kitchens where those who minister at the temple shall boil the sacrifices of the people."
EZEK|47|1|Then he brought me back to the door of the temple, and behold, water was issuing from below the threshold of the temple toward the east (for the temple faced east). The water was flowing down from below the south end of the threshold of the temple, south of the altar.
EZEK|47|2|Then he brought me out by way of the north gate and led me around on the outside to the outer gate that faces toward the east; and behold, the water was trickling out on the south side.
EZEK|47|3|Going on eastward with a measuring line in his hand, the man measured a thousand cubits, and then led me through the water, and it was ankle-deep.
EZEK|47|4|Again he measured a thousand, and led me through the water, and it was knee-deep. Again he measured a thousand, and led me through the water, and it was waist-deep.
EZEK|47|5|Again he measured a thousand, and it was a river that I could not pass through, for the water had risen. It was deep enough to swim in, a river that could not be passed through.
EZEK|47|6|And he said to me, "Son of man, have you seen this?" Then he led me back to the bank of the river.
EZEK|47|7|As I went back, I saw on the bank of the river very many trees on the one side and on the other.
EZEK|47|8|And he said to me, "This water flows toward the eastern region and goes down into the Arabah, and enters the sea; when the water flows into the sea, the water will become fresh.
EZEK|47|9|And wherever the river goes, every living creature that swarms will live, and there will be very many fish. For this water goes there, that the waters of the sea may become fresh; so everything will live where the river goes.
EZEK|47|10|Fishermen will stand beside the sea. From Engedi to En-eglaim it will be a place for the spreading of nets. Its fish will be of very many kinds, like the fish of the Great Sea.
EZEK|47|11|But its swamps and marshes will not become fresh; they are to be left for salt.
EZEK|47|12|And on the banks, on both sides of the river, there will grow all kinds of trees for food. Their leaves will not wither, nor their fruit fail, but they will bear fresh fruit every month, because the water for them flows from the sanctuary. Their fruit will be for food, and their leaves for healing."
EZEK|47|13|Thus says the Lord GOD: "This is the boundary by which you shall divide the land for inheritance among the twelve tribes of Israel. Joseph shall have two portions.
EZEK|47|14|And you shall divide equally what I swore to give to your fathers. This land shall fall to you as your inheritance.
EZEK|47|15|"This shall be the boundary of the land: On the north side, from the Great Sea by way of Hethlon to Lebo-hamath, and on to Zedad,
EZEK|47|16|Berothah, Sibraim (which lies on the border between Damascus and Hamath), as far as Hazer-hatticon, which is on the border of Hauran.
EZEK|47|17|So the boundary shall run from the sea to Hazar-enan, which is on the northern border of Damascus, with the border of Hamath to the north. This shall be the north side.
EZEK|47|18|"On the east side, the boundary shall run between Hauran and Da mascus; along the Jordan between Gilead and the land of Israel; to the eastern sea and as far as Tamar. This shall be the east side.
EZEK|47|19|"On the south side, it shall run from Tamar as far as the waters of Meribah-kadesh, from there along the Brook of Egypt to the Great Sea. This shall be the south side.
EZEK|47|20|"On the west side, the Great Sea shall be the boundary to a point opposite Lebo-hamath. This shall be the west side.
EZEK|47|21|"So you shall divide this land among you according to the tribes of Israel.
EZEK|47|22|You shall allot it as an inheritance for yourselves and for the sojourners who reside among you and have had children among you. They shall be to you as native-born children of Israel. With you they shall be allotted an inheritance among the tribes of Israel.
EZEK|47|23|In whatever tribe the sojourner resides, there you shall assign him his inheritance, declares the Lord GOD.
EZEK|48|1|"These are the names of the tribes: Beginning at the northern extreme, beside the way of Hethlon to Lebo-hamath, as far as Hazar-enan (which is on the northern border of Damascus over against Hamath), and extending from the east side to the west, Dan, one portion.
EZEK|48|2|Adjoining the territory of Dan, from the east side to the west, Asher, one portion.
EZEK|48|3|Adjoining the territory of Asher, from the east side to the west, Naphtali, one portion.
EZEK|48|4|Adjoining the territory of Naphtali, from the east side to the west, Manasseh, one portion.
EZEK|48|5|Adjoining the territory of Manasseh, from the east side to the west, Ephraim, one portion.
EZEK|48|6|Adjoining the territory of Ephraim, from the east side to the west, Reuben, one portion.
EZEK|48|7|Adjoining the territory of Reuben, from the east side to the west, Judah, one portion.
EZEK|48|8|"Adjoining the territory of Judah, from the east side to the west, shall be the portion which you shall set apart, 25,000 cubits in breadth, and in length equal to one of the tribal portions, from the east side to the west, with the sanctuary in the midst of it.
EZEK|48|9|The portion that you shall set apart for the LORD shall be 25,000 cubits in length, and 20,000 in breadth.
EZEK|48|10|These shall be the allotments of the holy portion: the priests shall have an allotment measuring 25,000 cubits on the northern side, 10,000 cubits in breadth on the western side, 10,000 in breadth on the eastern side, and 25,000 in length on the southern side, with the sanctuary of the LORD in the midst of it.
EZEK|48|11|This shall be for the consecrated priests, the sons of Zadok, who kept my charge, who did not go astray when the people of Israel went astray, as the Levites did.
EZEK|48|12|And it shall belong to them as a special portion from the holy portion of the land, a most holy place, adjoining the territory of the Levites.
EZEK|48|13|And alongside the territory of the priests, the Levites shall have an allotment 25,000 cubits in length and 10,000 in breadth. The whole length shall be 25,000 cubits and the breadth 20,000.
EZEK|48|14|They shall not sell or exchange any of it. They shall not alienate this choice portion of the land, for it is holy to the LORD.
EZEK|48|15|"The remainder, 5,000 cubits in breadth and 25,000 in length, shall be for common use for the city, for dwellings and for open country. In the midst of it shall be the city,
EZEK|48|16|and these shall be its measurements: the north side 4,500 cubits, the south side 4,500, the east side 4,500, and the west side 4,500.
EZEK|48|17|And the city shall have open land: on the north 250 cubits, on the south 250, on the east 250, and on the west 250.
EZEK|48|18|The remainder of the length alongside the holy portion shall be 10,000 cubits to the east, and 10,000 to the west, and it shall be alongside the holy portion. Its produce shall be food for the workers of the city.
EZEK|48|19|And the workers of the city, from all the tribes of Israel, shall till it.
EZEK|48|20|The whole portion that you shall set apart shall be 25,000 cubits square, that is, the holy portion together with the property of the city.
EZEK|48|21|"What remains on both sides of the holy portion and of the property of the city shall belong to the prince. Extending from the 25,000 cubits of the holy portion to the east border, and westward from the 25,000 cubits to the west border, parallel to the tribal portions, it shall belong to the prince. The holy portion with the sanctuary of the temple shall be in its midst.
EZEK|48|22|It shall be separate from the property of the Levites and the property of the city, which are in the midst of that which belongs to the prince. The portion of the prince shall lie between the territory of Judah and the territory of Benjamin.
EZEK|48|23|"As for the rest of the tribes: from the east side to the west, Benjamin, one portion.
EZEK|48|24|Adjoining the territory of Benjamin, from the east side to the west, Simeon, one portion.
EZEK|48|25|Adjoining the territory of Simeon, from the east side to the west, Issachar, one portion.
EZEK|48|26|Adjoining the territory of Issachar, from the east side to the west, Zebulun, one portion.
EZEK|48|27|Adjoining the territory of Zebulun, from the east side to the west, Gad, one portion.
EZEK|48|28|And adjoining the territory of Gad to the south, the boundary shall run from Tamar to the waters of Meribah-kadesh, from there along the Brook of Egypt to the Great Sea.
EZEK|48|29|This is the land that you shall allot as an inheritance among the tribes of Israel, and these are their portions, declares the Lord GOD.
EZEK|48|30|"These shall be the exits of the city: On the north side, which is to be 4,500 cubits by measure,
EZEK|48|31|three gates, the gate of Reuben, the gate of Judah, and the gate of Levi, the gates of the city being named after the tribes of Israel.
EZEK|48|32|On the east side, which is to be 4,500 cubits, three gates, the gate of Joseph, the gate of Benjamin, and the gate of Dan.
EZEK|48|33|On the south side, which is to be 4,500 cubits by measure, three gates, the gate of Simeon, the gate of Issachar, and the gate of Zebulun.
EZEK|48|34|On the west side, which is to be 4,500 cubits, three gates, the gate of Gad, the gate of Asher, and the gate of Naphtali.
EZEK|48|35|The circumference of the city shall be 18,000 cubits. And the name of the city from that time on shall be, The LORD is there."
