ZEPH|1|1|Слово Господнє, що було до Софонії, сина Куші, сина Ґедалії, сина Амарії, сина Єзекії, за днів Йосії, Амонового сина, Юдиного царя.
ZEPH|1|2|Забираючи, все заберу з-над поверхні землі, промовляє Господь.
ZEPH|1|3|Заберу Я людину й худобу, заберу птаство небесне і риби морські, і спокуси з безбожними, і витну людину з поверхні землі, промовляє Господь.
ZEPH|1|4|І руку Свою простягну Я на Юду і на всіх мешканців Єрусалиму, і вигублю з місця оцього останок Ваала, імення жерців зо священиками,
ZEPH|1|5|і тих, хто вклоняється на дахах світилам небесним, і тих, хто вклоняється, хто присягає Господом, і хто присягає царем своїм,
ZEPH|1|6|і тих, хто відступає від Господа, і хто не шукає Господа, і не звертається до Нього.
ZEPH|1|7|Замовчи перед Господом Богом, бо близький день Господній, бо жертву Господь приготовив, посвятив Своїх покликаних.
ZEPH|1|8|І станеться в день Господньої жертви, і навіщу Я князів, і синів царя, і всіх, хто зодягає одежу чужинну.
ZEPH|1|9|І навіщу Я кожного, хто перескакує через поріг того дня, тих, хто наповнює дім свого пана насиллям й оманою.
ZEPH|1|10|І буде в дні тому, говорить Господь, голос крику із Рибної брами, і завивання із Міста Нового, і велика руїна із пагірків.
ZEPH|1|11|Ридайте, мешканці Махтешу, бо понищений буде ввесь купецький народ, будуть вигублені всі, хто важить срібло.
ZEPH|1|12|І станеться часу того, і перешукаю Я з лямпами Єрусалим, і навіщу Я тих мужів, які задубіли на дріжджах своїх, що говорять у серці своєму: Господь не вчинить добра, і лиха не зробить.
ZEPH|1|13|І здобиччю стане все їхнє багатство, а їхні доми за спустошення, і будуть вони будувати доми, але в них не сидітимуть, і виноградники будуть садити, та вина їхнього не питимуть.
ZEPH|1|14|Близький день Господній великий, він близький й дуже швидко настане. Ось голос Господнього дня, тоді гірко кричатиме навіть хоробрий!
ZEPH|1|15|День гніву цей день, день смутку й насилля, день збурення та зруйнування, день темноти та темряви, день хмари й імли,
ZEPH|1|16|день сурмлення й окрику проти укріплених міст та проти високих міських заборолів.
ZEPH|1|17|І буду чинити Я утиск людині, і будуть ходити вони, як сліпі, бо згрішили вони проти Господа. І виллється кров їхня, немов той пісок, а їхнє тіло, як гній.
ZEPH|1|18|Спасти їх не зможе в день гніву Господнього ні їхнє срібло, ані золото їхнє, і огнем Його заздрощів буде поїджена ціла земля, бо скінчення тільки приспішене зробить зо всіми мешканцями Краю цього.
ZEPH|2|1|Посоромтеся та застидайтесь, народе без сорому,
ZEPH|2|2|поки народиться установлене, мине день, як полова! поки не прийде на вас лютість гніву Господнього, поки не прийде на вас день Господнього гніву!
ZEPH|2|3|Шукайте Господа, всі покірні землі, хто виконує право Його! Шукайте правди, шукайте смирення, може будете сховані ви в день Господнього гніву!
ZEPH|2|4|Бо покинута буде Азза, а Ашкелон опустошенням стане, Ашдод опівдня його виженуть, а Екрон буде вирваний.
ZEPH|2|5|Горе мешканцям довкілля морського, народові критському! Слово Господнє на вас, хананеї, краю филистимлян, Я тебе вигублю так, що не буде мешканця!
ZEPH|2|6|І буде довкілля морське пасовищами, повними ям пастухів та кошар для отари,
ZEPH|2|7|і буде оце побережжя останкові дому Юдиного, на них пасти будуть, у домах Ашкелону ввечорі будуть лягати, бо їх відвідає Господь, їхній Бог, і Він їхню долю приверне.
ZEPH|2|8|Чув Я ганьбу Моавову й образи Аммонових синів, які ображали народ Мій і чванилися над границею їхньою.
ZEPH|2|9|Тому як живий Я! говорить Господь Саваот, Бог Ізраїлів, стане Моав як Содом, а Аммонові сини як Гоморра: землею тернини, і солончаком, і навіки спустошенням! Пограбує їх решта народу Мого, а залишок люду Мого їх посяде.
ZEPH|2|10|Оце їм за їхню пиху, бо вони ображали й чванилися проти народу Господа Саваота.
ZEPH|2|11|Господь буде грізний проти них, бо Він знищить всіх богів землі, і вклонятися будуть Йому кожен з місця свого, усі острови тих народів.
ZEPH|2|12|Також ви, етіопляни, побиті мечем Моїм будете.
ZEPH|2|13|І на північ простягне Він руку Свою, та й погубить Ашшура, і Ніневію учинить спустошенням, суходолом, мов ту пустелю.
ZEPH|2|14|І будуть лежати серед неї стада, усяка польова звірина, і пелікан, і їжак будуть ночувати на мистецьких прикрасах її, сова буде кричати в вікні, на порозі ворона, бо віддерто кедрину його.
ZEPH|2|15|Оце оте радісне місто, що безпечно живе, що говорить у серці своєму: Я, і немає вже більше нікого! Як стало воно опустошенням, леговищем для звірини! Кожен, хто буде проходить повз нього, засвище, своєю рукою махне!
ZEPH|3|1|Горе місту тому ворохобному та занечищеному, місту насильникові!
ZEPH|3|2|Не слухається воно голосу, не приймає картання, не складає надії на Господа, до Бога свого не зближається.
ZEPH|3|3|Його зверхники посеред нього то леви ревучі, його судді вечірні вовки, які не лишають до ранку нічого.
ZEPH|3|4|Пророки його чванькуваті, зрадливі, його священики зневажають святиню, ламають Закона.
ZEPH|3|5|Серед нього Господь справедливий, Він кривди не чинить, щоранку дає Своє право на соняшне світло, не бракне його, але кривдник не відає сорому.
ZEPH|3|6|Народи Я вигубив, попустошені їхні заборола, Я вулиці їхні зруйнував, і нема перехожого, їхні міста поруйновані, так що немає й людини, немає й мешканця!
ZEPH|3|7|Я йому говорив: Тільки будеш боятись Мене, тільки приймеш картання, і не витяте буде мешкання його, усе, що про нього Я постановив, та вони ревно псули всі чини свої!
ZEPH|3|8|Тому то чекайте Мене, промовляє Господь, на той день, коли встану, як свідок, бо право Моє позбирати народи, згромадити царства, щоб вилити на них Свою лють, увесь жар Свого гніву, бо огнем Моїх заздрощів буде поглинута ціла земля!
ZEPH|3|9|Бо тоді уста чисті народам Я дам, щоб усі вони кликали Ймення Господнє, щоб раменом одним послужити Йому.
ZEPH|3|10|З другого боку річок Етіопії Моїх поклонників, Моїх розпорошених дарунком Мені принесуть.
ZEPH|3|11|Того дня ти не будеш соромитись всіма своїми ділами, якими грішив проти Мене, бо тоді Я відкину з твоєї середини тих, хто радіє твоєю пишнотою, і ти високо більш не стоятимеш вже на святій Моїй горі.
ZEPH|3|12|І серед тебе зоставлю убогий й нужденний народ, і будуть шукати пристановища в Іменні Господнім вони.
ZEPH|3|13|Останок Ізраїлів кривди не буде робити, і не будуть казати неправди, і облудний язик в їхніх устах не знайдеться, бо пастися будуть вони та вилежуватись, і не буде такого, хто б їх настрашив.
ZEPH|3|14|Співай, дочко Сіону! Втішайся, Ізраїлю! Радій та втішайся всім серцем, дочко Єрусалиму!
ZEPH|3|15|Відкинув Господь твої присуди, усунув у кут твого ворога! Серед тебе Господь, цар Ізраїлів, уже ти не будеш боятися зла!
ZEPH|3|16|Того дня буде сказане Єрусалимові: Не бійся! Сіонові: Нехай не опустяться руки твої!
ZEPH|3|17|Господь, Бог твій, серед тебе, Велет спасе! Він у радості буде втішатись тобою, обновить любов Свою, зо співом втішатися буде тобою!
ZEPH|3|18|Тих, що сумують за святами, Я позбираю, від тебе вони, тягарем над ними був сором.
ZEPH|3|19|Ось Я вчиню зо всіма мучителями твоїми кінець того часу, і спасу кульгаве, і позбираю розігнане, і зроблю їх хвалою та йменням у цілому Краї їхнього сорому.
ZEPH|3|20|Того часу спроваджу Я вас, і того часу Я вас позбираю, бо на ймення й на славу віддам вас поміж усіх народів землі, коли долю верну вам на ваших очах, промовляє Господь.
