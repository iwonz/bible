JUDG|1|1|Post mortem Iosue consulue runt filii Israel Dominum dicen tes: " Quis nostrum primus ascendet ad Chananaeum ad pugnandum contra eum? ".
JUDG|1|2|Dixitque Dominus: " Iudas ascendet: ecce tradidi terram in manus eius ".
JUDG|1|3|Et ait Iudas Simeoni fratri suo: " Ascende mecum in sorte mea, et pugnemus contra Chananaeum, et ego pergam tecum in sorte tua ". Et abiit cum eo Simeon.
JUDG|1|4|Ascenditque Iudas, et tradidit Dominus Chananaeum ac Pherezaeum in manus eorum, et percusserunt in Bezec decem milia virorum.
JUDG|1|5|Inveneruntque Adonibezec in Bezec et pugnaverunt contra eum ac percusserunt Chananaeum et Pherezaeum.
JUDG|1|6|Fugit autem Adonibezec, quem persecuti comprehenderunt, caesis pollicibus manuum eius ac pedum.
JUDG|1|7|Dixitque Adonibezec: " Septuaginta reges, amputatis manuum ac pedum pollicibus, colligebant sub mensa mea ciborum reliquias. Sicut feci, ita reddidit mihi Deus ". Adduxeruntque eum in Ierusalem, et ibi mortuus est.
JUDG|1|8|Oppugnantes ergo filii Iudae Ierusalem ceperunt eam; et percusserunt in ore gladii tradentes incendio civitatem.
JUDG|1|9|Et postea descendentes pugnaverunt contra Chananaeum, qui habitabat in montanis et in Nageb et in Sephela.
JUDG|1|10|Pergensque Iuda contra Chananaeum, qui habitabat in Hebron, cui nomen fuit antiquitus Cariatharbe, percussit Sesai et Ahiman et Tholmai.
JUDG|1|11|Atque inde profectus abiit ad habitatores Dabir, cuius nomen vetus erat Cariathsepher (id est civitas Litterarum).
JUDG|1|12|Dixitque Chaleb: " Qui percusserit Cariathsepher et ceperit eam, dabo ei Axam filiam meam uxorem ".
JUDG|1|13|Cumque cepisset eam Othoniel filius Cenez frater Chaleb minor, dedit ei Axam filiam suam coniugem.
JUDG|1|14|Quae cum veniret, incitavit eum, ut peteret a patre suo agrum. Demisit ergo se de asino, et dixit ei Chaleb: " Quid habes? ".
JUDG|1|15|At illa respondit: " Da mihi benedictionem; quia terram arentem dedisti mihi, da et irriguam aquis ". Dedit ergo ei Chaleb irriguum superius et irriguum inferius.
JUDG|1|16|Filii autem Hobab Cinaei cognati Moysi ascenderunt de civitate Palmarum cum filiis Iudae in desertum Iudae, quod est ad meridiem Arad, et habitaverunt cum Amalecitis.
JUDG|1|17|Abiit autem Iudas cum Simeone fratre suo et percusserunt simul Chananaeum, qui habitabat in Sephath, et percusserunt urbem anathemate. Vocatumque est nomen eius Horma (id est Anathema).
JUDG|1|18|Cepitque Iudas Gazam cum finibus suis et Ascalonem atque Accaron cum terminis suis.
JUDG|1|19|Fuitque Dominus cum Iuda, et montana possedit; nec potuit expellere habitatores vallis, quia falcatis curribus abundabant.
JUDG|1|20|Dederuntque Chaleb Hebron, sicut dixerat Moyses, qui expulit ex ea tres filios Enac.
JUDG|1|21|Iebusaeum autem habitatorem Ierusalem non expulerunt filii Beniamin, habitavitque Iebusaeus cum filiis Beniamin in Ierusalem usque in praesentem diem.
JUDG|1|22|Domus quoque Ioseph ascendit Bethel, fuitque Dominus cum eis.
JUDG|1|23|Nam, cum explorarent urbem, quae prius Luza vocabatur,
JUDG|1|24|viderunt custodes hominem egredientem de civitate dixeruntque ad eum: " Ostende nobis introitum civitatis, et faciemus tecum misericordiam ".
JUDG|1|25|Qui cum ostendisset eis, percusserunt urbem in ore gladii; hominem autem illum et omnem cognationem eius dimiserunt.
JUDG|1|26|Qui dimissus abiit in terram Hetthim et aedificavit ibi civitatem vocavitque eam Luzam, quae ita appellatur usque in praesentem diem.
JUDG|1|27|Manasses quoque non occupavit Bethsan et Thanach cum viculis suis nec expulit habitatores Dor et Ieblaam et Mageddo cum viculis suis; mansitque Chananaeus in terra hac.
JUDG|1|28|Postquam autem confortatus est Israel, fecit eos tributarios et expellere noluit.
JUDG|1|29|Ephraim etiam non expulit Chananaeum, qui habitabat in Gazer, sed habitavit Chananaeus in medio eius in Gazer.
JUDG|1|30|Zabulon non expulit habitatores Cetron et Naalol, sed habitavit Chananaeus in medio eius factusque est ei tributarius.
JUDG|1|31|Aser quoque non expulit habitatores Achcho et Sidonis, Ahalab et Achazib et Helba et Aphec et Rohob;
JUDG|1|32|habitavitque Aser in medio Chananaei habitatoris illius terrae, quia non expulit eum.
JUDG|1|33|Nephthali non expulit habitatores Bethsames et Bethanath et habitavit inter Chananaeum habitatorem terrae, fueruntque ei Bethsamitae et Bethanitae tributarii.
JUDG|1|34|Artavitque Amorraeus filios Dan in montem nec dedit eis locum, ut ad planiora descenderent.
JUDG|1|35|Habitavitque Amorraeus in Hathares, in Aialon et Salebim; et aggravata est manus domus Ioseph, factusque est ei tributarius.
JUDG|1|36|Fuit autem terminus Amorraei ab ascensu Acrabbim ad Petram et superiora loca.
JUDG|2|1|Ascenditque angelus Domini de Galgalis in Bochim et ait: " Eduxi vos de Aegypto et introduxi in terram, pro qua iuravi patribus vestris et pollicitus sum, ut non facerem irritum pactum meum vobiscum in sempiternum,
JUDG|2|2|ita dumtaxat ut non feriretis foedus cum habitatoribus terrae huius, sed aras eorum subverteretis. Et noluistis audire vocem meam. Cur hoc fecistis?
JUDG|2|3|Quam ob rem nolui expellere eos a facie vestra, ut sint vobis in laqueum, et dii eorum in ruinam ".
JUDG|2|4|Cumque loqueretur angelus Domini verba haec ad omnes filios Israel, elevaverunt vocem suam et fleverunt.
JUDG|2|5|Et vocatum est nomen loci illius Bochim (id est locus Flentium); immolaveruntque ibi hostias Domino.
JUDG|2|6|Dimisit ergo Iosue populum, et abierunt filii Israel unusquisque in possessionem suam, ut obtinerent terram.
JUDG|2|7|Servieruntque Domino cunctis diebus Iosue et seniorum, qui longo post eum vixerunt tempore et viderant universum opus magnum Domini, quod fecerat cum Israel.
JUDG|2|8|Mortuus est autem Iosue filius Nun famulus Domini centum et decem annorum;
JUDG|2|9|et sepelierunt eum in finibus possessionis suae in Thamnathsare in monte Ephraim a septentrionali plaga montis Gaas.
JUDG|2|10|Omnisque illa generatio congregata est ad patres suos, et surrexerunt alii post illam, qui non noverant Dominum et opus, quod fecerat cum Israel.
JUDG|2|11|Feceruntque filii Israel malum in conspectu Domini et servierunt Baalim
JUDG|2|12|ac dimiserunt Dominum, Deum patrum suorum, qui eduxerat eos de terra Aegypti, et secuti sunt deos alienos, de diis populorum, qui habitabant in circuitu eorum, et adoraverunt eos et ad iracundiam concitaverunt Dominum
JUDG|2|13|dimittentes eum et servientes Baal et Astharoth.
JUDG|2|14|Iratusque Dominus contra Israel tradidit eos in manibus diripientium, qui diripuerunt eos, et vendidit eos hostibus, qui habitabant per gyrum, nec potuerunt resistere adversariis suis;
JUDG|2|15|sed, quocumque pergere voluissent, manus Domini erat super eos ad malum, sicut locutus est et iuravit eis, et vehementer afflicti sunt.
JUDG|2|16|Suscitavitque Dominus iudices, qui liberarent eos de vastantium manibus;
JUDG|2|17|sed nec illos audire voluerunt fornicantes cum diis alienis et adorantes eos. Cito deseruerunt viam, per quam ingressi fuerant patres eorum audientes mandata Domini, et omnia fecere contraria.
JUDG|2|18|Cumque Dominus iudices suscitaret eis, erat Dominus cum iudice et liberabat eos de manu hostium eorum toto tempore iudicis, quia flectebatur misericordia et audiebat gemitus afflictorum.
JUDG|2|19|Postquam autem mortuus esset iudex, revertebantur et multo faciebant peiora quam fecerant patres sui, sequentes deos alienos, servientes eis et adorantes illos: non dimiserunt opera sua et viam durissimam, per quam ambulare consueverant.
JUDG|2|20|Iratusque est furor Domini in Israel et ait: " Quia irritum fecit gens ista pactum meum, quod pepigeram cum patribus eorum, et vocem meam audire contempsit,
JUDG|2|21|et ego non expellam gentes, quas dimisit Iosue et mortuus est;
JUDG|2|22|ut in ipsis experiar Israel, utrum custodiant viam Domini et ambulent in ea, sicut custodierunt patres eorum, an non ".
JUDG|2|23|Dimisit ergo Dominus has nationes et cito expellere noluit nec tradidit in manibus Iosue.
JUDG|3|1|Hae sunt gentes, quas Dominus dereliquit, ut erudiret in eis Is raelem, omnes, qui non noverant bella Chananaeorum,
JUDG|3|2|ut discerent certare cum hostibus generationes filiorum Israel, quae non habebant consuetudinem proeliandi:
JUDG|3|3|quinque satrapae Philisthinorum omnisque Chananaeus et Sidonius atque Hevaeus, qui habitabat in monte Libano de monte Baalhermon usque ad introitum Emath.
JUDG|3|4|Dimisitque eos, ut in ipsis experiretur Israelem, utrum audiret mandata Domini, quae praeceperat patribus eorum per manum Moysi, an non.
JUDG|3|5|Itaque filii Israel habitaverunt in medio Chananaei et Hetthaei et Amorraei et Pherezaei et Hevaei et Iebusaei
JUDG|3|6|et duxerunt uxores filias eorum, ipsique filias suas eorum filiis tradiderunt, et servierunt diis eorum.
JUDG|3|7|Feceruntque filii Israel malum in conspectu Domini et obliti sunt Domini Dei sui servientes Baalim et Astharoth.
JUDG|3|8|Iratusque Dominus contra Israel tradidit eos in manus Chusanrasathaim regis Mesopotamiae, servieruntque ei octo annis.
JUDG|3|9|Et clamaverunt ad Dominum, qui suscitavit eis salvatorem et liberavit eos, Othoniel videlicet filium Cenez fratrem Chaleb minorem.
JUDG|3|10|Fuitque in eo spiritus Domini, et iudicavit Israelem egressusque est ad pugnam; et tradidit Dominus in manu eius Chusanrasathaim regem Mesopotamiae, et praevaluit adversus eum.
JUDG|3|11|Quievitque terra quadraginta annis, et mortuus est Othoniel filius Cenez.
JUDG|3|12|Addiderunt autem filii Israel facere malum in conspectu Domini, qui confortavit adversum eos Eglon regem Moab, quia fecerunt malum in conspectu Domini.
JUDG|3|13|Et copulavit sibi Eglon filios Ammon et Amalec abiitque et percussit Israel atque possedit urbem Palmarum.
JUDG|3|14|Servieruntque filii Israel Eglon regi Moab decem et octo annis.
JUDG|3|15|Et clamaverunt filii Israel ad Dominum, qui suscitavit eis salvatorem Aod filium Gera de Beniamin, qui sinistra manu utebatur pro dextera. Miseruntque filii Israel per illum munera Eglon regi Moab.
JUDG|3|16|Fecitque Aod sibi gladium ancipitem longitudinis palmae manus et accinctus est eo subter vestem in dextro femore
JUDG|3|17|obtulitque munera Eglon regi Moab. Erat autem Eglon crassus nimis.
JUDG|3|18|Cumque obtulisset ei munera, dimisit socios, qui illa portaverant;
JUDG|3|19|et reversus de Galgalis, ubi erant idola, dixit ad regem: " Verbum secretum habeo ad te, o rex ". Et ille imperavit silentium; egressique sunt omnes, qui circa eum erant.
JUDG|3|20|Aod autem ingressus erat ad eum, cum sederet in aestivo cenaculo, quod ipsi soli erat, dixitque: " Verbum Dei habeo ad te ". Qui statim surrexit de throno.
JUDG|3|21|Extenditque Aod manum sinistram et tulit sicam de dextro femore suo infixitque eam in ventre eius
JUDG|3|22|tam valide, ut capulus ferrum sequeretur in vulnere ac pinguissimo adipe stringeretur. Nec eduxit gladium, sed ita, ut percusserat, reliquit in corpore; statimque per secreta naturae alvi stercora proruperunt.
JUDG|3|23|Aod autem egressus in atrium clausit ostium cenaculi post se et obfirmavit sera.
JUDG|3|24|Egresso illo, servi regis venerunt et, cum viderent clausas fores cenaculi, dixerunt: " Certe purgat alvum in aestivo cubiculo ".
JUDG|3|25|Exspectantesque diu, donec erubescerent, et videntes quod nullus aperiret, tulerunt clavem et aperientes invenerunt dominum suum iacentem in terra mortuum.
JUDG|3|26|Aod autem, dum illi cunctarentur, effugerat et pertransiit locum idolorum, unde reversus fuerat, venitque in Seira.
JUDG|3|27|Et statim insonuit bucina in monte Ephraim; descenderuntque cum eo filii Israel, ipso in fronte gradiente.
JUDG|3|28|Qui dixit ad eos: " Sequimini me; tradidit enim Dominus inimicos vestros Moabitas in manus vestras ". Descenderuntque post eum et occupaverunt vada Iordanis, quae transmittunt in Moab, et non dimiserunt transire quemquam,
JUDG|3|29|sed percusserunt Moabitas in tempore illo circiter decem milia, omnes robustos et fortes viros. Nullus eorum evadere potuit.
JUDG|3|30|Humiliatusque est Moab die illo sub manu Israel; et quievit terra octoginta annis.
JUDG|3|31|Post hunc fuit Samgar filius Anath, qui percussit de Philisthim sescentos viros stimulo boum; et ipse quoque salvum fecit Israel.
JUDG|4|1|Addideruntque filii Israel facere malum in conspectu Domini post mortem Aod,
JUDG|4|2|et tradidit illos Dominus in manu Iabin regis Chanaan, qui regnavit in Asor. Habuitque ducem exercitus sui nomine Sisaram: ipse autem habitabat in Haroseth gentium.
JUDG|4|3|Clamaveruntque filii Israel ad Dominum; nongentos enim habebat falcatos currus et per viginti annos vehementer oppresserat eos.
JUDG|4|4|Erat autem Debora prophetis, uxor Lapidoth, quae iudicabat Israel in illo tempore.
JUDG|4|5|Et sedebat sub palma Deborae inter Rama et Bethel in monte Ephraim; ascendebantque ad eam filii Israel in iudicium.
JUDG|4|6|Quae misit et vocavit Barac filium Abinoem de Cedes Nephthali dixitque ad eum: " Praecepit tibi Dominus, Deus Israel: Vade et duc exercitum in montem Thabor tollesque tecum decem milia pugnatorum de filiis Nephthali et de filiis Zabulon.
JUDG|4|7|Ego autem ducam ad te in loco torrentis Cison Sisaram principem exercitus Iabin et currus eius atque omnem multitudinem et tradam eum in manu tua ".
JUDG|4|8|Dixitque ad eam Barac: " Si venis mecum, vadam; si nolueris venire mecum, non pergam ".
JUDG|4|9|Quae dixit ad eum: " Ibo quidem tecum; sed in hac via non erit tibi gloria, quia in manu mulieris tradet Dominus Sisaram ".Surrexit itaque Debora et perrexit cum Barac in Cedes.
JUDG|4|10|Qui, accitis Zabulon et Nephthali in Cedes, ascendit cum decem milibus pugnatorum habens Deboram in comitatu suo.
JUDG|4|11|Haber autem Cinaeus recesserat a ceteris Cinaeis fratribus suis filiis Hobab cognati Moysi et tetendit tabernaculum usque ad quercum in Saananim iuxta Cedes.
JUDG|4|12|Nuntiatumque est Sisarae quod ascendisset Barac filius Abinoem in montem Thabor,
JUDG|4|13|et congregavit omnes nongentos falcatos currus omnemque exercitum, qui cum eo erat, de Haroseth gentium ad torrentem Cison.
JUDG|4|14|Dixitque Debora ad Barac: " Surge: haec est enim dies, in qua tradidit Dominus Sisaram in manus tuas. En ipse ductor est tuus ". Descendit itaque Barac de monte Thabor, et decem milia pugnatorum cum eo.
JUDG|4|15|Perterruitque Dominus Sisaram et omnes currus eius universamque multitudinem in ore gladii ad conspectum Barac, in tantum ut Sisara de curru desiliens pedibus fugeret,
JUDG|4|16|et Barac persequeretur fugientes currus et exercitum usque ad Haroseth gentium, et omnis hostium multitudo usque ad internecionem caderet.
JUDG|4|17|Sisara autem fugiens pervenit ad tentorium Iahel uxoris Haber Cinaei; erat enim pax inter Iabin regem Asor et domum Haber Cinaei.
JUDG|4|18|Egressa igitur Iahel in occursum Sisarae dixit ad eum: " Intra ad me, domine mi; intra, ne timeas ". Qui ingressus tabernaculum eius et opertus ab ea panno,
JUDG|4|19|dixit ad eam: " Da mihi, obsecro, paululum aquae, quia sitio ". Quae aperuit utrem lactis et dedit ei bibere et operuit illum.
JUDG|4|20|Dixitque Sisara ad eam: " Sta ante ostium tabernaculi et, cum venerit aliquis interrogans te et dicens: "Numquid hic est aliquis?", respondebis: Nullus est" ".
JUDG|4|21|Tulit porro Iahel uxor Haber clavum tabernaculi assumens pariter malleum; et ingressa abscondite et cum silentio, posuit supra tempus capitis eius clavum, percussumque malleo defixit in cerebrum usque ad terram; qui soporem morti socians defecit et mortuus est.
JUDG|4|22|Et ecce Barac sequens Sisaram veniebat; egressaque Iahel in occursum eius dixit ei: " Veni, et ostendam tibi virum, quem quaeris ". Qui cum intrasset ad eam, vidit Sisaram iacentem mortuum et clavum infixum in tempore eius.
JUDG|4|23|Humiliavit ergo Deus in die illo Iabin regem Chanaan coram filiis Israel,
JUDG|4|24|qui crescebant cotidie et forti manu opprimebant Iabin regem Chanaan, donec delerent eum.
JUDG|5|1|Cecineruntque Debora et Barac filius Abinoem in die illo dicen tes:
JUDG|5|2|" Quia comae excussae sunt in Israel,cum sponte se obtulit populus,benedicite Domino!
JUDG|5|3|Audite, reges, percipite auribus, principes;ego sum, ego sum, quae Domino canam,psallam Domino, Deo Israel!
JUDG|5|4|Domine, cum exires de Seir,incederes de regione Edom,terra mota est, caelique stillaverunt, ac nubes stillaverunt aquis;
JUDG|5|5|montes fluxerunt a facie Domini Sinai,a facie Domini, Dei Israel.
JUDG|5|6|In diebus Samgar filii Anath,in diebus Iahel quieverunt semitae; et, qui ingrediebantur per eas,ambulaverunt per calles devios.
JUDG|5|7|Cessaverunt fortes in Israel et quieverunt,donec surgeres, Debora,surgeres mater in Israel.
JUDG|5|8|Elegerunt deos novos;tunc erat pugna in portis.Clipeus et hasta non apparueruntin quadraginta milibus Israel.
JUDG|5|9|Cor meum diligit principes Israel.Qui sponte obtulistis vos in populo, benedicite Domino!
JUDG|5|10|Qui ascenditis super nitentes asinaset sedetis super tapetiaet ambulatis in via, loquimini.
JUDG|5|11|Ad vocem eorum,qui distribuunt aquas ad canales,ibi narrant iustitias Domini,iustitias fortitudinis eius in Israel:tunc descendit populus Domini ad portas.
JUDG|5|12|Surge, surge, Debora;surge, surge et loquere canticum!Surge, Barac, et apprehende captivos tuos,fili Abinoem!
JUDG|5|13|Tunc descenderunt reliquiae ad inclitos,populus Domini descendit pro eo in fortibus.
JUDG|5|14|Ex Ephraim venerunt principes in vallempost te, Beniamin, in populis tuis.De Machir principes descenderunt, et de Zabulon, qui tenent sceptrum, praefecti.
JUDG|5|15|Duces Issachar fuere cum Debora;sic Barac in vallem missus cum peditibus suis.In pagis Ruben magna consilia cordis.
JUDG|5|16|Quare sedebas inter caulas,ut audires sibilos tibiae apud greges?Pagis Ruben magnae investigationes cordis.
JUDG|5|17|Galaad trans Iordanem quiescebat;et Dan cur peregrinus vacabat navibus?Aser habitabat in litore mariset in portibus morabatur.
JUDG|5|18|Zabulon vero obtulit animam suam morti,et Nephthali super excelsa regionis.
JUDG|5|19|Venerunt reges et pugnaverunt,pugnaverunt reges Chanaanin Thanach iuxta aquas Mageddo, praedam argenti non tulere!
JUDG|5|20|De caelo dimicaverunt stellae,cursu suo adversus Sisaram pugnaverunt.
JUDG|5|21|Torrens Cison traxit cadavera eorum,torrens proeliorum, torrens Cison; incede, anima mea, fortiter.
JUDG|5|22|Tunc calcaverunt ungulae equorumin cursu praecipiti fortium suorum.
JUDG|5|23|Maledicite, Meroz, dixit angelus Domini,maledicite habitatoribus eius,quia non venerunt ad auxilium Domini,in adiutorium Domini in fortibus.
JUDG|5|24|Benedicta prae mulieribus Iahel uxor Haber Cinaei,prae mulieribus tabernaculi benedicatur!
JUDG|5|25|Aquam petenti lac deditet in phiala principum obtulit butyrum.
JUDG|5|26|Sinistram manum misit ad clavumet dextram ad fabrorum malleum:percussitque Sisaram quaerens in capite vulneri locumet tempus valide perforans.
JUDG|5|27|Inter pedes eius ruit, cecidit, iacebat;inter pedes eius ruit, cecidit;ubi ruit, ibi iacebat exanimis.
JUDG|5|28|Per fenestram prospiciens eiulabatmater Sisarae per cancellos:Cur moratur regredi currus eius? Quare tardant rotae quadrigarum illius?".
JUDG|5|29|Una sapientior ceteris uxoribus respondit ei,et ipsa sibi repetit verba illius:
JUDG|5|30|"Certo nunc dividunt inventa spolia, unam, duas feminas singulis viris;duas vestes diversorum colorumSisarae in praedam;unam, duas texturas discolorescollo meo in praedam".
JUDG|5|31|Sic pereant omnes inimici tui, Domine!Qui autem diligunt eum, rutilent,sicut sol in ortu suo splendet ".
JUDG|5|32|Quievitque terra per quadraginta annos.
JUDG|6|1|Fecerunt autem filii Israel malum in conspectu Domini, qui tradidit eos in manu Madian septem annis.
JUDG|6|2|Et oppressi sunt valde ab eis. Feceruntque sibi antra et speluncas in montibus et tutissima loca.
JUDG|6|3|Cumque sevisset Israel, ascendebat Madian et Amalec ceterique orientalium nationum
JUDG|6|4|et apud eos figentes tentoria, sicut erant in herbis, cuncta vastabant usque ad introitum Gazae nihilque omnino ad vitam pertinens relinquebant in Israel, non oves, non boves, non asinos.
JUDG|6|5|Ipsi enim et universi greges eorum veniebant cum tabernaculis suis et, instar locustarum, universa complebant, innumera multitudo hominum et camelorum, quidquid tetigerant devastantes.
JUDG|6|6|Humiliatusque est Israel valde in conspectu Madian.
JUDG|6|7|Et clamavit ad Dominum postulans auxilium contra Madianitas.
JUDG|6|8|Qui misit ad eos virum prophetam, et locutus est: " Haec dicit Dominus, Deus Israel: Ego vos feci conscendere de Aegypto et eduxi vos de domo servitutis
JUDG|6|9|et liberavi de manu Aegyptiorum et omnium inimicorum, qui affligebant vos, eiecique eos ad introitum vestrum et tradidi vobis terram eorum.
JUDG|6|10|Et dixi: Ego Dominus Deus vester, ne timeatis deos Amorraeorum, in quorum terra habitatis. Et noluistis audire vocem meam ".
JUDG|6|11|Venit autem angelus Domini et sedit sub quercu, quae erat in Ephra et pertinebat ad Ioas de familia Abiezer. Cumque Gedeon filius eius excuteret atque purgaret frumenta in torculari, ut absconderet a Madian,
JUDG|6|12|apparuit ei angelus Domini et ait: " Dominus tecum, vir fortis! ".
JUDG|6|13|Dixitque ei Gedeon: " Obsecro, domine mi, si Dominus nobiscum est, cur apprehenderunt nos haec omnia? Ubi sunt omnia mirabilia eius, quae narraverunt patres nostri atque dixerunt: "De Aegypto eduxit nos Dominus"? Nunc autem dereliquit nos Dominus et tradidit in manu Madian ".
JUDG|6|14|Respexitque ad eum Dominus et ait: " Vade in hac fortitudine tua et liberabis Israel de manu Madian; scito quod miserim te ".
JUDG|6|15|Qui respondens ait: " Obsecro, Domine, in quo liberabo Israel? Ecce familia mea infima est in Manasse, et ego minimus in domo patris mei ".
JUDG|6|16|Dixitque ei Dominus: " Ego ero tecum, et percuties Madian quasi unum virum ".
JUDG|6|17|Et ille: " Si inveni, inquit, gratiam coram te, da mihi signum quod tu sis, qui loquaris ad me;
JUDG|6|18|ne recedas hinc, donec revertar ad te portans oblationem et offerens tibi ". Qui respondit: " Ego praestolabor adventum tuum ".
JUDG|6|19|Ingressus est itaque Gedeon et coxit haedum et de farinae ephi azymos panes; carnesque ponens in canistro et ius carnium mittens in ollam tulit omnia sub quercum et obtulit ei.
JUDG|6|20|Cui dixit angelus Dei: " Tolle carnes et panes azymos et pone super petram illam et ius desuper funde ". Cumque fecisset ita,
JUDG|6|21|extendit angelus Domini summitatem virgae, quam tenebat in manu, et tetigit carnes et azymos panes, ascenditque ignis de petra et carnes azymosque panes consumpsit. Angelus autem Domini evanuit ex oculis eius.
JUDG|6|22|Vidensque Gedeon quod esset angelus Domini ait: "Heu mihi, Domine Deus, quia vidi angelum Domini facie ad faciem! ".
JUDG|6|23|Dixitque ei Dominus: " Pax tecum, ne timeas, non morieris! ".
JUDG|6|24|Aedificavit ergo ibi Gedeon altare Domino vocavitque illud: " Dominus pax "; usque in praesentem diem adhuc est in Ephra filiorum Abiezer.
JUDG|6|25|Nocte illa dixit Dominus ad eum: " Tolle taurum patris tui, alterum taurum scilicet annorum septem, destruesque aram Baal, quae est patris tui, et palum, qui iuxta aram est, succide;
JUDG|6|26|et aedificabis altare Domino Deo tuo in summitate petrae huius secundum ordinem; tollesque taurum secundum et offeres holocaustum super struem lignorum pali, quem succideris ".
JUDG|6|27|Assumptis igitur Gedeon decem viris de servis suis, fecit, sicut praeceperat Dominus; timens autem domum patris sui et homines illius civitatis per diem facere noluit, sed omnia nocte complevit.
JUDG|6|28|Cumque surrexissent viri oppidi eius mane, viderunt destructam aram Baal palumque succisum et taurum alterum impositum super altare, quod tunc aedificatum erat.
JUDG|6|29|Dixeruntque ad invicem: " Quis hoc fecit? ". Cumque perquirerent auctorem facti, dictum est: " Gedeon filius Ioas fecit haec omnia ".
JUDG|6|30|Et dixerunt ad Ioas: " Produc filium tuum, ut moriatur, quia destruxit aram Baal et succidit palum ".
JUDG|6|31|Respondit Ioas omnibus, qui circumdabant eum: " Numquid certare vultis pro Baal et salvare eum? Qui certabit pro Baal, morietur usque mane. Si Deus est, certet pro seipso contra eum, qui destruxit aram eius ".
JUDG|6|32|Ex illo die vocatus est Gedeon Ierobbaal, eo quod dicebatur: " Certet contra eum Baal, quia destruxit altare eius ".
JUDG|6|33|Igitur omnis Madian et Amalec et orientales populi congregati sunt simul et transeuntes Iordanem castrametati sunt in valle Iezrahel.
JUDG|6|34|Spiritus autem Domini induit Gedeon, qui clangens bucina convocavit domum Abiezer, ut sequeretur.
JUDG|6|35|Misitque nuntios in universum Manassen, qui et ipse secutus est eum; et alios nuntios in Aser et Zabulon et Nephthali, qui occurrerunt ei.
JUDG|6|36|Dixitque Gedeon ad Deum: " Si salvum facis per manum meam Israel, sicut locutus es,
JUDG|6|37|ponam vellus lanae in area: si ros in solo vellere fuerit, et in omni terra siccitas, sciam quod per manum meam, sicut locutus es, liberabis Israel ".
JUDG|6|38|Factumque est ita. Et de nocte consurgens, expresso vellere concham rore complevit.
JUDG|6|39|Dixitque rursus ad Deum: " Ne irascatur furor tuus contra me, si adhuc semel tentavero signum quaerens in vellere. Oro, ut solum vellus siccum sit, et omnis terra rore madens ".
JUDG|6|40|Fecitque Deus nocte illa, ut postulaverat; et fuit siccitas in solo vellere, et ros in omni terra.
JUDG|7|1|Igitur Ierobbaal, qui et Gedeon, de nocte consurgens et omnis populus cum eo castrame tati sunt ad fontem, qui vocatur Harad. Erant autem castra Madian in valle ad septentrionalem plagam collis Moreh.
JUDG|7|2|Dixitque Dominus ad Gedeon: " Maior tecum est populus, quam ut tradatur Madian in manus eius, ne glorietur contra me Israel et dicat: "Meis viribus liberatus sum".
JUDG|7|3|Loquere ad populum et, cunctis audientibus, praedica: "Qui formidolosus et timidus est, revertatur et recedat de monte Gelboe" ". Et reversa sunt ex populo viginti duo milia virorum; et tantum decem milia remanserunt.
JUDG|7|4|Dixitque Dominus ad Gedeon: " Adhuc populus multus est; duc eos ad aquas, et ibi probabo illos, et, de quo dixero tibi ut tecum vadat, ipse pergat; quem ire prohibuero, revertatur ".
JUDG|7|5|Cumque deduxisset populum ad aquas, dixit Dominus ad Gedeon: " Qui lingua lambuerint aquas, sicut solent canes lambere, separabis eos seorsum; qui autem curvatis genibus biberint, in altera parte erunt ".
JUDG|7|6|Fuit itaque numerus eorum, qui manu ad os proiciente aquas lambuerant, trecenti viri; omnis autem reliqua multitudo flexo poplite biberat.
JUDG|7|7|Et ait Dominus ad Gedeon: " In trecentis viris, qui lambuerunt aquas, liberabo vos et tradam Madian in manu tua; omnis autem reliqua multitudo revertatur in locum suum ".
JUDG|7|8|Sumptis itaque pro numero cibariis et tubis, omnem reliquam multitudinem abire praecepit ad tabernacula sua et ipse trecentos viros tenuit. Castra autem Madian erant subter eum in valle.
JUDG|7|9|Eadem nocte dixit Dominus ad eum: " Surge et descende in castra, quia tradidi ea in manu tua.
JUDG|7|10|Sin autem ire formidas, descendat tecum Phara puer tuus.
JUDG|7|11|Et, cum audieris quid loquantur, tunc confortabuntur manus tuae, et securior ad hostium castra descendes ". Descendit ergo ipse et Phara puer eius in partem castrorum, ubi erant armatorum vigiliae.
JUDG|7|12|Madian autem et Amalec et omnes orientales populi fusi iacebant in valle ut locustarum multitudo; cameli quoque innumerabiles erant sicut arena, quae iacet in litoribus maris.
JUDG|7|13|Cumque venisset Gedeon, narrabat aliquis somnium proximo suo et dicebat: " Ecce vidi somnium, et videbatur mihi quasi subcinericius panis ex hordeo volvi et in Madian castra descendere; cumque pervenisset ad tabernaculum, percussit illud atque subvertit et terrae funditus coaequavit ".
JUDG|7|14|Respondit is, cui loquebatur: "Non est hoc aliud nisi gladius Gedeonis filii Ioas viri Israelitae; tradidit Deus in manu eius Madian et omnia castra eius ".
JUDG|7|15|Cumque audisset Gedeon somnium et interpretationem eius, adoravit et reversus ad castra Israel ait: " Surgite, tradidit enim Dominus in manus vestras castra Madian ".
JUDG|7|16|Divisitque trecentos viros in tres partes et dedit tubas in manibus eorum lagoenasque vacuas ac lampades in medio lagoenarum
JUDG|7|17|et dixit ad eos: " Quod me facere videritis, hoc facite; ingrediar extremam partem castrorum, et, quod fecero, sectamini.
JUDG|7|18|Quando personaverit tuba in manu mea et omnium eorum, qui mecum sunt, vos quoque per castrorum circuitum clangite et conclamate: "Domino et Gedeoni!" ".
JUDG|7|19|Ingressusque est Gedeon et trecenti viri, qui erant cum eo, extremam partem castrorum, incipientibus vigiliis noctis mediae, cum eo ipso tempore custodes mutati essent, et coeperunt bucinis clangere et conterere lagoenas.
JUDG|7|20|Cumque in tribus personarent turmis et hydrias confregissent, tenuerunt sinistris manibus lampades et dextris sonantes tubas clamaveruntque: " Gladius Domino et Gedeoni! ",
JUDG|7|21|stantes singuli in loco suo per circuitum castrorum hostilium. Omnia itaque castra turbata sunt, et vociferantes ululantesque fugerunt.
JUDG|7|22|Et insistebant trecenti viri bucinis personantes. Immisitque Dominus gladium in omnibus castris, et mutua se caede truncabant fugientes usque Bethsetta, Sareda et crepidinem Abelmehula in Tebbath.
JUDG|7|23|Convocati autem viri Israel de Nephthali et Aser et omni Manasse persequebantur Madian.
JUDG|7|24|Misitque Gedeon nuntios in omnem montem Ephraim dicens: " Descendite in occursum Madian et occupate aquas usque Bethbera atque Iordanem ". Omnis Ephraim praeoccupavit aquas usque Bethbera atque Iordanem.
JUDG|7|25|Apprehensosque duos principes Madian Oreb et Zeb interfecit Oreb in Petra Oreb, Zeb vero in Torculari Zeb; et persecuti sunt Madian capita Oreb et Zeb portantes ad Gedeon trans fluenta Iordanis.
JUDG|8|1|Dixeruntque ad eum viri Ephraim: " Quid est hoc quod nobis facere voluisti, ut non nos vocares, cum ad pugnam pergeres contra Madian? ", iurgantes fortiter et prope vim inferentes.
JUDG|8|2|Quibus ille respondit: " Quid enim tale facere potui, quale vos fecistis? Nonne melior est racemus Ephraim vindemiis Abiezer?
JUDG|8|3|In manus vestras Deus tradidit principes Madian Oreb et Zeb. Quid tale facere potui, quale vos fecistis? ". Quod cum locutus esset, requievit spiritus eorum, quo tumebant contra eum.
JUDG|8|4|Cumque venisset Gedeon ad Iordanem, transivit eum cum trecentis viris, qui secum erant et prae lassitudine fugientes persequi vix poterant.
JUDG|8|5|Dixitque ad viros Succoth: "Date, obsecro, panes populo, qui mecum est, quia valde defecerunt, et ego persequor Zebee et Salmana reges Madian ".
JUDG|8|6|Responderunt principes Succoth: " Forsitan palmae manuum Zebee et Salmana in manu tua sunt, ut demus exercitui tuo panes? ".
JUDG|8|7|Quibus ille ait: " Cum ergo tradiderit Dominus Zebee et Salmana in manus meas, triturabo carnes vestras cum spinis deserti et tribulis ".
JUDG|8|8|Et inde conscendens venit in Phanuel locutusque est ad viros eius loci similia. Cui et illi responderunt, sicut responderant viri Succoth.
JUDG|8|9|Dixit itaque et eis: "Cum reversus fuero in pace, destruam turrim hanc".
JUDG|8|10|Zebee autem et Salmana requiescebant in Carcar cum omni exercitu suo, quasi quindecim milia viri, qui remanserant ex omnibus turmis orientalium populorum, caesis centum viginti milibus bellatorum educentium gladium.
JUDG|8|11|Ascendensque Gedeon per viam eorum, qui in tabernaculis morabantur ad orientalem partem Nobe et Iegbaa, percussit castra hostium, qui securi erant et nihil adversi suspicabantur.
JUDG|8|12|Fugeruntque Zebee et Salmana. Persequens Gedeon comprehendit duos reges Madian Zebee et Salmana, turbato omni exercitu eorum.
JUDG|8|13|Revertensque Gedeon filius Ioas de bello per ascensum Hares,
JUDG|8|14|apprehendit puerum de viris Succoth interrogavitque eum nomina principum et seniorum Succoth, qui scripsit ei septuaginta septem viros.
JUDG|8|15|Venitque ad viros Succoth et dixit eis: "En Zebee et Salmana, super quibus exprobrastis mihi dicentes: "Forsitan manus Zebee et Salmana in manibus tuis sunt, ut demus viris tuis, qui lassi sunt, panes?" ".
JUDG|8|16|Tulit ergo seniores civitatis et spinas deserti ac tribulos; et trituravit cum eis viros Succoth.
JUDG|8|17|Turrim quoque Phanuel subvertit, occisis habitatoribus civitatis.
JUDG|8|18|Dixitque ad Zebee et Salmana: " Quales fuerunt viri, quos occidistis in Thabor? ". Qui responderunt: " Similes tui, et unusquisque ex eis quasi filius regis ".
JUDG|8|19|Quibus ille ait: " Fratres mei fuerunt, filii matris meae. Vivit Dominus, si servassetis eos, non vos occiderem! ".
JUDG|8|20|Dixitque Iether primogenito suo: " Surge et interfice eos! ". Qui non eduxit gladium; timebat enim, quia adhuc puer erat.
JUDG|8|21|Dixeruntque Zebee et Salmana: " Tu surge et irrue in nos, quia iuxta aetatem robur est hominis ". Surrexit Gedeon et interfecit Zebee et Salmana et tulit lunulas, quibus colla camelorum eorum decorata erant.
JUDG|8|22|Dixeruntque viri Israel ad Gedeon: " Dominare nostri, tu et filius tuus et filius filii tui, quia liberasti nos de manu Madian ".
JUDG|8|23|Quibus ille ait: " Non dominabor vestri, nec dominabitur in vos filius meus, sed dominabitur Dominus ".
JUDG|8|24|Dixitque ad eos: " Unam petitionem postulo a vobis: date mihi unusquisque anulum ex praeda sua ". Anulos enim aureos Ismaelitae habere consuerant.
JUDG|8|25|Qui responderunt: " Libentissime dabimus ". Expandentesque super terram pallium proiecerunt in eo unusquisque anulum de praeda sua.
JUDG|8|26|Et fuit pondus postulatorum anulorum mille septingenti auri sicli absque lunulis et inauribus et vestibus purpureis, quibus Madian reges uti soliti erant, et praeter torques camelorum.
JUDG|8|27|Fecitque ex eo Gedeon ephod et posuit illud in civitate sua Ephra. Fornicatusque est omnis Israel in eo, et factum est Gedeoni et omni domui eius in ruinam.
JUDG|8|28|Humiliatus est autem Madian coram filiis Israel, nec potuerunt ultra elevare cervices, sed quievit terra per quadraginta annos, quibus Gedeon vivebat.
JUDG|8|29|Abiit itaque Ierobbaal filius Ioas et habitavit in domo sua;
JUDG|8|30|habuitque Gedeon septuaginta filios, qui egressi sunt de femore eius, eo quod multas haberet uxores.
JUDG|8|31|Concubina quoque illius, quam habebat in Sichem, genuit ei filium, cui ipse nomen imposuit Abimelech.
JUDG|8|32|Mortuusque est Gedeon filius Ioas in senectute bona et sepultus est in sepulcro Ioas patris sui in Ephra filiorum Abiezer.
JUDG|8|33|Postquam autem mortuus est Gedeon, aversi sunt filii Israel et fornicati cum Baalim posuerunt sibi Baalberith in deum.
JUDG|8|34|Nec recordati sunt Domini Dei sui, qui eruit eos de manu omnium inimicorum suorum per circuitum,
JUDG|8|35|nec fecerunt misericordiam cum domo Ierobbaal Gedeon iuxta omnia bona, quae fecerat Israeli.
JUDG|9|1|Abiit autem Abimelech filius Ierobbaal in Sichem ad fratres matris suae et locutus est ad eos et ad omnem cognationem familiae matris suae dicens:
JUDG|9|2|" Loquimini ad omnes viros Sichem: "Quid vobis est melius, ut dominentur vestri septuaginta viri, omnes filii Ierobbaal, an ut dominetur vobis unus vir? Simulque considerate quod os vestrum et caro vestra sum" ".
JUDG|9|3|Locutique sunt fratres matris eius de eo ad omnes viros Sichem universos sermones istos et inclinaverunt cor eorum post Abimelech dicentes: " Frater noster est ".
JUDG|9|4|Dederuntque illi septuaginta pondo argenti de fano Baalberith; qui conduxit sibi ex eo viros inopes et vagos, secutique sunt eum.
JUDG|9|5|Et venit in domum patris sui Ephra et occidit fratres suos filios Ierobbaal septuaginta viros super lapidem unum. Remansitque Ioatham filius Ierobbaal minimus, quia absconditus erat.
JUDG|9|6|Congregati sunt autem omnes viri Sichem et universae domus Mello abieruntque et constituerunt regem Abimelech iuxta quercum, quae stabat in Sichem.
JUDG|9|7|Quod cum nuntiatum esset Ioatham, ivit et stetit in vertice montis Garizim elevataque voce clamavit et dixit: " Audite me, viri Sichem, ut audiat vos Deus.
JUDG|9|8|Ierunt ligna, ut ungerent super se regem, dixeruntque olivae: "Impera nobis".
JUDG|9|9|Quae respondit: "Numquid possum deserere pinguedinem meam, qua et dii honorantur et homines, et venire, ut super ligna movear?".
JUDG|9|10|Dixeruntque ligna ad arborem ficum: "Veni et super nos regnum accipe".
JUDG|9|11|Quae respondit eis: "Numquid possum deserere dulcedinem meam fructusque suavissimos et ire, ut super cetera ligna movear?".
JUDG|9|12|Locuta quoque sunt ligna ad vitem: "Veni et impera nobis".
JUDG|9|13|Quae respondit: "Numquid possum deserere vinum meum, quod laetificat deos et homines, et super ligna cetera commoveri?".
JUDG|9|14|Dixeruntque omnia ligna ad rhamnum: "Veni et impera super nos".
JUDG|9|15|Quae respondit eis: "Si vere me regem vobis constituitis, venite et sub mea umbra requiescite; sin autem non vultis, egrediatur ignis de rhamno et devoret cedros Libani!".
JUDG|9|16|Nunc igitur, si recte et absque peccato constituistis super vos regem Abimelech et bene egistis cum Ierobbaal et cum domo eius et reddidistis vicem beneficiis eius,
JUDG|9|17|qui pugnavit pro vobis et animam suam dedit periculis, ut erueret vos de manu Madian,
JUDG|9|18|qui nunc surrexistis contra domum patris mei et interfecistis filios eius septuaginta viros super unum lapidem et constituistis regem Abimelech filium ancillae eius super habitatores Sichem, eo quod frater vester sit;
JUDG|9|19|si ergo recte et absque vitio egistis cum Ierobbaal et domo eius hodie, laetamini in Abimelech, et ille laetetur in vobis.
JUDG|9|20|Sin autem perverse, egrediatur ignis ex Abimelech et consumat habitatores Sichem et domum Mello, egrediaturque ignis de viris Sichem et de domo Mello et devoret Abimelech! ".
JUDG|9|21|Quae cum Ioatham dixisset, fugit et abiit in Bera habitavitque ibi metu Abimelech fratris sui.
JUDG|9|22|Regnavit itaque Abimelech super Israel tribus annis.
JUDG|9|23|Misitque Deus spiritum pessimum inter Abimelech et habitatores Sichem, qui rebellaverunt contra eum,
JUDG|9|24|ut scelus interfectionis septuaginta filiorum Ierobbaal et effusio sanguinis eorum veniret super Abimelech fratrem suum et in viros Sichimorum, qui eum adiuverant.
JUDG|9|25|Posueruntque insidias adversus eum in montium summitate et exercebant latrocinia agentes praedas de omnibus praetereuntibus. Nuntiatumque est Abimelech.
JUDG|9|26|Venit autem Gaal filius Ebed cum fratribus suis et transivit in Sichimam, et confisi sunt habitatores Sichem in eo.
JUDG|9|27|Egressi in agros vindemiaverunt vineas uvasque calcaverunt et, factis cantantium choris, ingressi sunt fanum dei sui et inter epulas et pocula maledicebant Abimelech,
JUDG|9|28|clamante Gaal filio Ebed: " Quis est Abimelech, et quae est Sichem, ut serviamus ei? Numquid non est filius Ierobbaal et Zebul praefectus eius? Servite viris Hemmor patris Sichem! Cur serviemus ei?
JUDG|9|29|Utinam daret aliquis populum istum sub manu mea, ut auferrem de medio Abimelech et dicerem ei: Congrega exercitus multitudinem et veni ".
JUDG|9|30|Zebul princeps civitatis, auditis sermonibus Gaal filii Ebed, iratus est valde
JUDG|9|31|et misit clam ad Abimelech nuntios dicens: " Ecce Gaal filius Ebed venit in Sichimam cum fratribus suis et excitant adversum te civitatem.
JUDG|9|32|Surge itaque nocte cum populo, qui tecum est, et latita in agro.
JUDG|9|33|Et primo mane, oriente sole, irrue super civitatem; illo autem egrediente adversum te cum populo suo, fac ei, quod potueris ".
JUDG|9|34|Surrexit itaque Abimelech cum omni exercitu suo nocte et tetendit insidias iuxta Sichimam in quattuor locis.
JUDG|9|35|Egressusque est Gaal filius Ebed et stetit in introitu portae civitatis; surrexit autem Abimelech et omnis exercitus cum eo de insidiarum loco.
JUDG|9|36|Cumque vidisset populum Gaal, dixit ad Zebul: " Ecce de montibus multitudo descendit ". Cui ille respondit: " Umbras montium vides quasi homines ".
JUDG|9|37|Rursumque Gaal ait: " Ecce populus de Umbilico terrae descendit, et unus cuneus venit per viam Quercus Augurum ".
JUDG|9|38|Cui dixit Zebul: " Ubi est nunc os tuum, quo loquebaris: "Quis est Abimelech, ut serviamus ei?". Nonne iste est populus, quem despiciebas? Egredere et pugna contra eum ".
JUDG|9|39|Abiit ergo Gaal, spectante Sichimorum populo, et pugnavit contra Abimelech.
JUDG|9|40|Qui persecutus est eum fugientem, cecideruntque ex parte eius plurimi usque ad portam civitatis.
JUDG|9|41|Et Abimelech sedit in Aruma; Zebul autem Gaal et fratres eius expulit de urbe nec in ea passus est commorari.
JUDG|9|42|Sequenti ergo die egressus est populus in campum. Quod cum nuntiatum esset Abimelech,
JUDG|9|43|tulit exercitum suum et divisit in tres turmas tendens insidias in agris. Vidensque quod egrederetur populus de civitate, surrexit et percussit eos.
JUDG|9|44|Irruensque cum cuneo suo obsedit ingressum portae civitatis; duae autem turmae palantes per campum adversarios percusserunt.
JUDG|9|45|Porro Abimelech omni illo die oppugnabat urbem, quam cepit, interfectis habitatoribus eius ipsaque destructa, ita ut sal in ea dispergeret.
JUDG|9|46|Quod cum audissent, qui habitabant in turre Sichimorum, ingressi sunt cryptam fani Elberith (id est dei Foederis).
JUDG|9|47|Abimelech quoque audiens omnes viros turris Sichimorum pariter conglobatos,
JUDG|9|48|ascendit in montem Selmon cum omni populo suo et, arrepta securi, praecidit arboris ramum impositumque ferens umero dixit ad socios: " Quod me viditis facere, cito facite ".
JUDG|9|49|Igitur certatim ramos de arboribus praecidentes sequebantur ducem, quos circumdantes cryptae succenderunt; atque ita factum est, ut fumo et igne omnes homines necarentur, circiter mille viri pariter ac mulieres, habitatores turris Sichem.
JUDG|9|50|Abimelech autem inde proficiscens venit ad oppidum Thebes, quod obsidebat et cepit.
JUDG|9|51|Erat autem turris fortis in media civitate, ad quam confugerant viri simul ac mulieres et omnes cives civitatis, clausa firmissime ianua, et super turris tectum stantes per propugnacula.
JUDG|9|52|Accedensque Abimelech iuxta turrim pugnabat fortiter et appropinquans ostio ignem supponere nitebatur.
JUDG|9|53|Et ecce una mulier superiorem molam desuper iaciens illisit capiti Abimelech et confregit cerebrum eius.
JUDG|9|54|Qui vocavit cito armigerum suum et ait ad eum: " Evagina gladium tuum et percute me, ne forte dicatur quod a femina interfectus sim ". Qui transfodit eum.
JUDG|9|55|Illoque mortuo, omnes viri Israel hoc videntes reversi sunt in sedes suas.
JUDG|9|56|Et reddidit Deus malum, quod fecerat Abimelech contra patrem suum, interfectis septuaginta fratribus suis.
JUDG|9|57|Sichimitis quoque, quod operati erant, retributum est, et venit super eos maledictio Ioatham filii Ierobbaal.
JUDG|10|1|Post Abimelech surrexit dux ad salvandum Israel Thola fi lius Phua filii Dodo, vir de Issachar, qui habitavit in Samir montis Ephraim.
JUDG|10|2|Et iudicavit Israel viginti et tribus annis mortuusque ac sepultus est in Samir.
JUDG|10|3|Huic successit Iair Galaadites, qui iudicavit Israel per viginti et duos annos
JUDG|10|4|habens triginta filios sedentes super triginta pullos asinarum, et ipsis erant triginta civitates, quae appellatae sunt Havoth Iair (id est villae Iair) usque in praesentem diem, in terra Galaad.
JUDG|10|5|Mortuusque est Iair ac sepultus in Camon.
JUDG|10|6|Filii autem Israel peccatis veteribus iungentes nova fecerunt malum in conspectu Domini et servierunt Baalim et Astharoth et diis Syriae ac Sidonis et Moab et filiorum Ammon et Philisthim; dimiseruntque Dominum et non colebant eum.
JUDG|10|7|Contra quos iratus tradidit eos in manu Philisthim et filiorum Ammon.
JUDG|10|8|Afflictique sunt et vehementer oppressi per annos decem et octo omnes filii Israel, qui habitabant trans Iordanem in terra Amorraei in Galaad;
JUDG|10|9|in tantum ut filii Ammon Iordanem transirent ad pugnandum etiam contra Iudam et Beniamin et domum Ephraim; afflictusque est Israel nimis.
JUDG|10|10|Et clamantes filii Israel ad Dominum dixerunt: " Peccavimus tibi, quia dereliquimus Deum nostrum et servivimus Baalim ".
JUDG|10|11|Quibus locutus est Dominus: " Numquid non Aegyptii et Amorraei filiique Ammon et Philisthim,
JUDG|10|12|Sidonii quoque et Amalec et Madian oppresserunt vos, et clamastis ad me, et erui vos de manu eorum?
JUDG|10|13|Et tamen reliquistis me et coluistis deos alienos; idcirco non addam ut ultra vos liberem.
JUDG|10|14|Ite et invocate deos, quos elegistis: ipsi vos liberent in tempore angustiae! ".
JUDG|10|15|Dixeruntque filii Israel ad Dominum: "Peccavimus; redde tu nobis, quidquid tibi placet, tantum nunc libera nos ".
JUDG|10|16|Quae dicentes omnia de finibus suis alienorum deorum idola proiecerunt et servierunt Domino, qui doluit super miseriis Israel.
JUDG|10|17|Itaque filii Ammon convocati in Galaad fixere tentoria; contra quos congregati filii Israel in Maspha castrametati sunt.
JUDG|10|18|Dixeruntque populus, principes Galaad, singuli ad proximos suos: " Qui primus contra filios Ammon coeperit dimicare, erit dux omnium habitatorum Galaad ".
JUDG|11|1|Fuit Iephte Galaadites vir fortissimus, filius meretricis mulieris, quem genuit Galaad.
JUDG|11|2|Habuit autem Galaad uxorem, de qua suscepit filios, qui, postquam creverant, eiecerunt Iephte dicentes: " Heres in domo patris nostri esse non poteris, quia de altera matre generatus es ".
JUDG|11|3|Quos ille fugiens atque devitans habitavit in terra Tob; congregatique sunt ad eum viri inopes et exierunt cum eo.
JUDG|11|4|In illis diebus pugnabant filii Ammon contra Israel.
JUDG|11|5|Quibus acriter instantibus, perrexerunt maiores natu de Galaad, ut tollerent in auxilium sui Iephte de terra Tob.
JUDG|11|6|Dixeruntque ad eum: " Veni et esto princeps noster, et pugnemus contra filios Ammon ".
JUDG|11|7|Quibus ille respondit: " Nonne vos estis, qui odistis me et eiecistis de domo patris mei? Et nunc venistis ad me necessitate compulsi ".
JUDG|11|8|Dixeruntque principes Galaad ad Iephte: " Ob hanc igitur causam nunc ad te venimus, ut proficiscaris nobiscum et pugnes contra filios Ammon sisque dux omnium, qui habitant in Galaad ".
JUDG|11|9|Iephte quoque dixit eis: " Si revocatis me, ut pugnem pro vobis contra filios Ammon, tradideritque eos Dominus in manus meas, ego ero princeps vester ".
JUDG|11|10|Qui responderunt ei: " Dominus, qui haec audit, ipse mediator ac testis est quod secundum verbum tuum faciemus ".
JUDG|11|11|Abiit itaque Iephte cum principibus Galaad, fecitque eum omnis populus principem sui. Locutusque est Iephte omnes sermones suos coram Domino in Maspha.
JUDG|11|12|Et misit Iephte nuntios ad regem filiorum Ammon, qui ex persona sua dicerent: " Quid mihi et tibi est, quia venisti contra me, ut invaderes terram meam? ".
JUDG|11|13|Quibus ille respondit: " Quia tulit Israel terram meam, quando ascendit de Aegypto, a finibus Arnon usque Iaboc atque Iordanem; nunc igitur cum pace redde mihi eam ".
JUDG|11|14|Rursumque Iephte nuntios misit et imperavit eis, ut dicerent regi Ammon:
JUDG|11|15|" Haec dicit Iephte: Non tulit Israel terram Moab nec terram filiorum Ammon.
JUDG|11|16|Sed, quando de Aegypto conscenderunt, ambulavit Israel per solitudinem usque ad mare Rubrum et venit in Cades;
JUDG|11|17|misitque nuntios ad regem Edom dicens: "Dimitte, ut transeam per terram tuam". Qui noluit acquiescere precibus eius. Misit quoque et ad regem Moab, qui et ipse transitum praebere contempsit. Mansit itaque Israel in Cades
JUDG|11|18|et pertransiens desertum circuivit ex latere terram Edom et terram Moab venitque contra orientalem plagam terrae Moab et castrametatus est trans Arnon nec voluit intrare terminos Moab; Arnon quippe confinium est terrae Moab.
JUDG|11|19|Misit itaque Israel nuntios ad Sehon regem Amorraeorum, regem Hesebon, et dixit ei: "Dimitte, ut transeam per terram tuam usque ad locum meum".
JUDG|11|20|Qui et ipse Israel verbis diffidens non dimisit eum transire per terminos suos, sed, omni populo suo congregato, egressus est contra eum in Iasa et fortiter resistebat.
JUDG|11|21|Tradiditque eum Dominus in manu Israel cum omni exercitu suo, qui percussit eum et possedit omnem terram Amorraei habitatoris regionis illius,
JUDG|11|22|universos fines eius de Arnon usque Iaboc et de solitudine usque ad Iordanem.
JUDG|11|23|Dominus ergo, Deus Israel, subvertit Amorraeum coram populo suo Israel; et tu nunc vis possidere terram eius?
JUDG|11|24|Nonne ea, quae tibi Chamos deus tuus in possessionem dat, tibi iure debentur? Quae autem Dominus Deus noster victor obtinuit, in nostram cedunt possessionem.
JUDG|11|25|Num quid melior es Balac filio Sephor rege Moab? Numquid iurgatus est contra Israel et pugnavit contra eum?
JUDG|11|26|Quando habitabat in Hesebon et viculis eius et in Aroer et villis illius et in cunctis civitatibus iuxta Arnon per trecentos annos, quare tanto tempore nihil super hac repetitione tentastis?
JUDG|11|27|Igitur non ego pecco in te, sed tu contra me male agis indicens mihi bella non iusta. Iudicet Dominus arbiter huius diei inter filios Israel et inter filios Ammon ".
JUDG|11|28|Noluitque acquiescere rex filiorum Ammon verbis Iephte, quae per nuntios mandaverat.
JUDG|11|29|Factus est ergo super Iephte spiritus Domini, et pertransiens Galaad et Manasse venit in Maspha Galaad et inde ad filios Ammon.
JUDG|11|30|Votum autem vovit Domino dicens: " Si tradideris filios Ammon in manus meas,
JUDG|11|31|quicumque primus fuerit egressus de foribus domus meae mihique occurrerit revertenti cum pace a filiis Ammon, eum holocaustum offeram Domino ".
JUDG|11|32|Transivitque Iephte ad filios Ammon, ut pugnaret contra eos; quos tradidit Dominus in manus eius.
JUDG|11|33|Percussitque eos ab Aroer usque dum venias in Mennith viginti civitates et usque ad Abelcharmim plaga magna nimis; humiliatique sunt filii Ammon a filiis Israel.
JUDG|11|34|Revertenti autem Iephte in Maspha domum suam occurrit unigenita filia cum tympanis et choris: non enim habebat alios liberos.
JUDG|11|35|Qua visa, scidit vestimenta sua et ait: " Heu, filia mi, incurvans incurvasti me! Et tu es in eis, qui me perturbant! Aperui enim os meum ad Dominum et aliud facere non potero ".
JUDG|11|36|Cui illa respondit: " Pater mi, si aperuisti os tuum ad Dominum, fac mihi, quodcumque pollicitus es, concessa tibi a Domino ultione atque victoria de hostibus tuis filiis Ammon ".
JUDG|11|37|Dixitque ad patrem: " Hoc solum mihi praesta, quod deprecor: Dimitte me, ut duobus mensibus circumeam montes et plangam virginitatem meam cum sodalibus meis ".
JUDG|11|38|Cui ille respondit: " Vade! ". Et dimisit eam duobus mensibus. Cumque abisset cum sodalibus suis, flebat virginitatem suam in montibus.
JUDG|11|39|Expletisque duobus mensibus, reversa est ad patrem suum; et fecit ei, sicut voverat, quae non cognoverat virum. Exinde mos increbuit in Israel, et consuetudo servata est,
JUDG|11|40|ut post anni circulum conveniant in unum filiae Israel et plangant filiam Iephte Galaaditae diebus quattuor.
JUDG|12|1|Ecce autem convocatus vir Ephraim transiit contra aqui lonem, et dixerunt ad Iephte: " Quare vadens ad pugnam contra filios Ammon vocare nos noluisti, ut pergeremus tecum? Igitur incendemus domum tuam super te.
JUDG|12|2|Quibus ille respondit: " Disceptatio erat mihi et populo meo contra filios Ammon vehemens, vocavique vos, ut mihi praeberetis auxilium, et facere noluistis.
JUDG|12|3|Quod cernens posui in manibus meis animam meam transivique ad filios Ammon, et tradidit eos Dominus in manus meas. Quid commerui, ut hodie adversum me consurgatis in proelium? ".
JUDG|12|4|Vocatis itaque ad se cunctis viris Galaad, pugnabat contra Ephraim. Percusseruntque viri Galaad Ephraim, quia dixerat: " Fugitivi de Ephraim estis; Galaad habitat in medio Ephraim et Manasse ".
JUDG|12|5|Occupaveruntque Galaaditae vada Iordanis, per quae Ephraim reversurus erat. Cumque venisset ad ea de Ephraim numero fugiens atque dixisset: " Obsecro, ut me transire permittatis ", dicebant ei Galaaditae: " Numquid Ephrathaeus es? ". Quo dicente: " Non sum ",
JUDG|12|6|interrogabant eum: " Dic ergo: Scibboleth " (quod interpretatur Spica). Qui respondebat: " Sibboleth ", illud recte exprimere non valens. Statimque apprehensum iugulabant in ipso Iordanis transitu. Et ceciderunt in illo tempore de Ephraim quadraginta duo milia.
JUDG|12|7|Iudicavitque Iephte Galaadites Israel sex annis et mortuus est ac sepultus in civitate sua in Galaad.
JUDG|12|8|Post hunc iudicavit Israel Abesan de Bethlehem.
JUDG|12|9|Qui habuit triginta filios et totidem filias emittens foras maritis dedit; et eiusdem numeri filiis suis accepit uxores forinsecus. Qui septem annis iudicavit Israel;
JUDG|12|10|mortuusque est ac sepultus in Bethlehem.
JUDG|12|11|Cui successit Ahialon Zabulonites et iudicavit Israel decem annis;
JUDG|12|12|mortuusque est ac sepultus in Ahialon terrae Zabulon.
JUDG|12|13|Post hunc iudicavit Israel Abdon filius Illel Pharathonites.
JUDG|12|14|Qui habuit quadraginta filios et triginta ex eis nepotes ascendentes super septuaginta pullos asinarum. Et iudicavit Israel octo annis;
JUDG|12|15|mortuusque est ac sepultus in Pharathon terrae Ephraim in monte Amalecite.
JUDG|13|1|Rursumque filii Israel fece runt malum in conspectu Do mini, qui tradidit eos in manus Philisthinorum quadraginta annis.
JUDG|13|2|Erat autem vir quidam de Saraa et de stirpe Dan nomine Manue habens uxorem sterilem.
JUDG|13|3|Cui apparuit angelus Domini et dixit ad eam: " Ecce sterilis es et absque liberis, sed concipies et paries filium.
JUDG|13|4|Cave ergo, ne vinum bibas ac siceram nec immundum quidquam comedas,
JUDG|13|5|quia ecce concipies et paries filium, cuius non tanget caput novacula: erit enim puer nazaraeus Dei ex matris utero et ipse incipiet liberare Israel de manu Philisthinorum ".
JUDG|13|6|Quae cum venisset ad maritum, dixit ei: " Vir Dei venit ad me habens aspectum sicut angelus Domini, terribilis nimis. Non interrogavi eum, unde esset, nec ipse nomen suum mihi indicavit.
JUDG|13|7|Et dixit mihi: "Ecce concipies et paries filium; cave, ne vinum bibas et siceram et ne aliquo vescaris immundo: erit enim puer nazaraeus Dei ex utero matris usque ad diem mortis suae" ".
JUDG|13|8|Oravit itaque Manue Dominum et ait: " Obsecro, Domine, ut vir Dei, quem misisti, veniat iterum et doceat nos, quid debeamus facere de puero, qui nasciturus est ".
JUDG|13|9|Exaudivitque Deus precantem Manue, et venit rursum angelus Dei ad mulierem sedentem in agro. Manue autem maritus eius non erat cum ea.
JUDG|13|10|Festinavit ergo et cucurrit ad virum suum nuntiavitque ei dicens: " Ecce apparuit mihi vir, qui illo die venerat ad me ".
JUDG|13|11|Qui surrexit et secutus est uxorem suam veniensque ad virum dixit ei: " Tu es, qui locutus es mulieri? ". Et ille respondit: " Ego sum ".
JUDG|13|12|Cui Manue: " Quando, inquit, sermo tuus fuerit expletus, quid circa puerum observare et facere debemus? ".
JUDG|13|13|Dixitque angelus Domini ad Manue: " Ab omnibus, quae locutus sum uxori tuae, abstineat se;
JUDG|13|14|et, quidquid ex vinea nascitur, non comedat, vinum et siceram non bibat, nullo vescatur immundo et, quod ei praecepi, custodiat ".
JUDG|13|15|Dixitque Manue ad angelum Domini: " Obsecro, ut retineamus te et faciamus tibi haedum de capris ".
JUDG|13|16|Cui respondit angelus Domini: " Si me retines, non comedam panes tuos; sin autem vis holocaustum facere, offer illud Domino ". Et nesciebat Manue quod angelus Domini esset.
JUDG|13|17|Dixitque ad eum: " Quod est tibi nomen, ut, si sermo tuus fuerit expletus, honoremus te? ".
JUDG|13|18|Cui ille respondit: " Cur quaeris nomen meum, quod est mirabile? ".
JUDG|13|19|Tulit itaque Manue haedum de capris et oblationem similae et posuit super petram offerens Domino, qui facit mirabilia; ipse autem et uxor eius intuebantur.
JUDG|13|20|Cumque ascenderet flamma de altari in caelum, angelus Domini in flamma pariter ascendit. Quod cum vidisset Manue et uxor eius, proni ceciderunt in terram;
JUDG|13|21|et ultra non eis apparuit angelus Domini. Statimque intellexit Manue angelum esse Domini
JUDG|13|22|et dixit ad uxorem suam: " Morte moriemur, quia vidimus Deum ".
JUDG|13|23|Cui respondit mulier: " Si Dominus nos vellet occidere, de manibus nostris holocaustum et oblationem non suscepisset nec ostendisset nobis haec omnia neque talia dixisset ".
JUDG|13|24|Peperit itaque filium et vocavit nomen eius Samson. Crevitque puer, et benedixit ei Dominus.
JUDG|13|25|Coepitque spiritus Domini impellere eum in Castris Dan inter Saraa et Esthaol.
JUDG|14|1|Descendit igitur Samson in Thamna vidensque ibi mulie rem de filiabus Philisthim
JUDG|14|2|ascendit et nuntiavit patri suo et matri dicens: " Vidi mulierem in Thamna de filiabus Philisthinorum, quam quaeso ut mihi accipiatis uxorem.
JUDG|14|3|Cui dixerunt pater et mater sua: " Numquid non est mulier in filiabus fratrum tuorum et in omni populo meo, quia vis accipere uxorem de Philisthim, qui incircumcisi sunt? ". Dixitque Samson ad patrem suum: " Hanc mihi accipe, quia placuit oculis meis ".
JUDG|14|4|Parentes autem eius nesciebant quod res a Domino fieret, et quaereret occasionem contra Philisthim. Eo enim tempore Philisthim dominabantur Israeli.
JUDG|14|5|Descendit itaque Samson cum patre suo et matre in Thamna. Cumque venissent ad vineas oppidi, apparuit catulus leonis rugiens et occurrit ei.
JUDG|14|6|Irruit autem spiritus Domini in Samson, et dilaceravit leonem, quasi haedum in frusta concerperet, nihil omnino habens in manu; et hoc patri et matri noluit indicare.
JUDG|14|7|Descenditque et locutus est mulieri, quae placuerat oculis eius.
JUDG|14|8|Et post aliquot dies revertens, ut acciperet eam, declinavit, ut videret cadaver leonis; et ecce examen apum in corpore leonis erat ac favus mellis.
JUDG|14|9|Quem, cum sumpsisset in manibus, comedebat in via; veniensque ad patrem suum et matrem dedit eis partem, qui et ipsi comederunt. Nec tamen eis voluit indicare quod mel de corpore leonis assumpserat.
JUDG|14|10|Descendit itaque pater eius ad mulierem, et fecit ibi Samson convivium; sic enim iuvenes facere consuerant.
JUDG|14|11|Cum ergo cives loci illius vidissent eum, dederunt ei sodales triginta, qui essent cum eo.
JUDG|14|12|Quibus locutus est Samson: " Proponam vobis problema, quod si solveritis mihi intra septem dies convivii, dabo vobis triginta tunicas et totidem vestes mutatorias;
JUDG|14|13|sin autem non potueritis solvere, vos dabitis mihi triginta tunicas et eiusdem numeri vestes mutatorias ". Qui responderunt ei: " Propone problema, ut audiamus ".
JUDG|14|14|Dixitque eis: De comedente exivit cibus,et de forti est egressa dulcedo ".Nec potuerunt per tres dies propositionem solvere.
JUDG|14|15|Cumque adesset dies quartus, dixerunt ad uxorem Samson: " Blandire viro tuo et suade ei, ut indicet tibi quid significet problema. Quod si facere nolueris, incendemus et te et domum patris tui. An idcirco nos vocastis ad nuptias, ut spoliaretis? ".
JUDG|14|16|Quae fundebat apud Samson lacrimas et querebatur dicens: " Odisti me et non diligis; idcirco problema, quod proposuisti filiis populi mei, non vis mihi exponere ". At ille respondit: " Patri meo et matri nolui dicere et tibi indicare potero? ".
JUDG|14|17|Septem igitur diebus convivii flebat apud eum; tandemque die septimo, cum ei molesta esset, exposuit. Quae statim indicavit civibus suis,
JUDG|14|18|et illi dixerunt ei die septimo ante solis occubitum: Quid dulcius melle,et quid leone fortius? ".Qui ait ad eos: Si non arassetis in vitula mea,non invenissetis propositionem meam ".
JUDG|14|19|Irruit itaque in eo spiritus Domini, descenditque Ascalonem et percussit ibi triginta viros, quorum ablatas vestes dedit iis, qui problema solverant; iratusque nimis ascendit in domum patris sui.
JUDG|14|20|Uxor autem eius accepit maritum unum de amicis eius, qui erat pronubus.
JUDG|15|1|Post aliquantum autem tem poris, cum dies triticeae mes sis instarent, venit Samson invisere volens uxorem suam et attulit ei haedum de capris. Cumque ad eam vellet intrare, prohibuit eum pater illius
JUDG|15|2|dicens: " Putavi quod odisses eam et ideo tradidi illam amico tuo; sed habet sororem iuniorem, quae pulchrior illa est; sit tibi pro ea uxor ".
JUDG|15|3|Dixitque eis Samson: " Hac vice non erit culpa in me contra Philisthaeos, cum faciam eis mala ".
JUDG|15|4|Perrexitque et cepit trecentas vulpes caudasque earum iunxit ad caudas sumensque faces ligavit singulas in medio binarum caudarum;
JUDG|15|5|facibusque igne succensis, dimisit vulpes in segetes Philisthinorum. Et comportatae iam fruges et adhuc stantes in stipula concrematae sunt in tantum, ut vineas quoque et oliveta flamma consumeret.
JUDG|15|6|Dixeruntque Philisthim: " Quis fecit hanc rem? ". Quibus dictum est: " Samson gener Thamnathaei, quia tulit uxorem eius et alteri tradidit, haec operatus est ". Ascenderuntque Philisthim et combusserunt tam mulierem quam patrem eius.
JUDG|15|7|Quibus ait Samson: " Si talia facitis, utique ex vobis expetam ultionem et tunc quiescam ".
JUDG|15|8|Percussitque eos ingenti plaga, suram ad femur. Et descendens habitavit in spelunca petrae Etam.
JUDG|15|9|Igitur ascendentes Philisthim in terra Iudae castrametati sunt, et in Lehi (id est Maxilla) eorum est fusus exercitus.
JUDG|15|10|Dixeruntque ad eos viri de tribu Iudae: " Cur ascendistis adversum nos?. Qui responderunt: " Ut ligemus Samson venimus et reddamus ei, quae in nos operatus est ".
JUDG|15|11|Descenderunt ergo tria milia virorum de Iuda ad specum petrae Etam dixeruntque ad Samson: " Nescis quod Philisthim imperent nobis? Quare hoc nobis facere voluisti? ". Quibus ille ait: " Sicut fecerunt mihi, feci eis.
JUDG|15|12|" Ligare, inquiunt, te venimus et tradere in manus Philisthinorum ". " Iurate, respondit, mihi quod non me occidatis ".
JUDG|15|13|Dixerunt: " Non te occidemus, sed vinctum trademus ". Ligaveruntque eum duobus novis funibus et tulerunt de petra Etam.
JUDG|15|14|Qui cum venisset in Lehi, et Philisthim vociferantes occurrissent ei, irruit spiritus Domini in eum, et, sicut solent ad odorem ignis lina consumi, ita vincula, quibus brachia eius ligata erant, dissipata sunt et soluta.
JUDG|15|15|Inventamque maxillam asini recentem arripiens percussit in ea mille viros
JUDG|15|16|et ait: In maxilla asiniacervum feci ex eis!In mandibula asinipercussi mille viros! ".
JUDG|15|17|Cumque haec canens verba complesset, proiecit mandibulam de manu et vocavit nomen loci illius Ramathlehi (quod interpretatur Elevatio maxillae).
JUDG|15|18|Sitiensque valde clamavit ad Dominum et ait: " Tu dedisti in manu servi tui salutem hanc maximam atque victoriam; et en siti morior incidamque in manus incircumcisorum ".
JUDG|15|19|Aperuit itaque Deus fossam in Lehi, et egressae sunt inde aquae; quibus haustis, refocillavit spiritum et vires recepit. Idcirco appellatum est nomen fontis illius fons Invocantis, qui est in Lehi usque in praesentem diem.
JUDG|15|20|Iudicavitque Israel in diebus Philisthim viginti annis.
JUDG|16|1|Abiit Samson in Gazam et vidit ibi meretricem mulie rem ingressusque est ad eam.
JUDG|16|2|Cum nuntiatum esset Gazaeis intrasse urbem Samson, circuierunt et insidiabantur ei in porta civitatis; tota autem nocte quieverunt praestolantes, ut, facto mane, exeuntem occiderent.
JUDG|16|3|Dormivit autem Samson usque ad noctis medium et inde consurgens apprehendit ambas portae fores cum postibus suis et evellit eas cum sera, impositasque umeris portavit ad verticem montis, qui respicit Hebron.
JUDG|16|4|Post haec amavit mulierem, quae habitabat in valle Sorec et vocabatur Dalila.
JUDG|16|5|Veneruntque ad eam principes Philisthinorum atque dixerunt: " Decipe eum et disce ab illo in quo tantam habeat fortitudinem, et quomodo eum superare valeamus et vinctum humiliare; quod si feceris, dabimus tibi singuli mille centum argenteos ".
JUDG|16|6|Locuta est ergo Dalila ad Samson: " Dic mihi, obsecro, in quo sit tua maxima fortitudo, et quid sit, quo ligatus humilieris ".
JUDG|16|7|Cui respondit Samson: " Si septem nerviceis funibus necdum siccis et adhuc humentibus ligatus fuero, deficiam eroque ut ceteri homines ".
JUDG|16|8|Attuleruntque ad eam satrapae Philisthinorum septem funes, ut dixerat; quibus vinxit eum,
JUDG|16|9|latentibus apud se insidiis in cubiculo. Clamavitque ad eum: " Philisthim super te, Samson! ". Qui rupit vincula, quomodo si rumpat quis filum de stuppa tortum, cum odorem ignis acceperit; et non est cognitum in quo esset fortitudo eius.
JUDG|16|10|Dixitque ad eum Dalila: " Ecce illusisti mihi et falsum locutus es; saltem nunc indica mihi quo ligari debeas ".
JUDG|16|11|Cui ille respondit: " Si ligatus fuero novis funibus, qui numquam fuerunt in opere, infirmus ero et aliorum hominum similis ".
JUDG|16|12|Quibus rursum Dalila vinxit eum et clamavit: " Philisthim super te, Samson! ", in cubiculo insidiis praeparatis. Qui ita rupit vincula brachiorum quasi fila telarum.
JUDG|16|13|Dixitque Dalila rursum ad eum: " Usquequo decipis me et falsum loqueris? Ostende quo vinciri debeas ". Cui respondit Samson: " Si septem crines nexos capitis mei cum licio plexueris et paxillo fixeris, deficiam eroque ut ceteri homines ".
JUDG|16|14|Quae cum dormire eum fecisset et septem crines nexos capitis eius cum licio plexisset et paxillo fixisset, dixit ad eum: " Philisthim super te, Samson! ". Qui consurgens de somno extraxit paxillum cum navicula et licio.
JUDG|16|15|Dixitque ad eum Dalila: " Quomodo dicis quod ames me, cum animus tuus non sit mecum? Per tres vices mentitus es mihi et noluisti dicere in quo sit tua maxima fortitudo ".
JUDG|16|16|Cumque molesta ei esset et per multos dies iugiter eum urgeret, defecit anima eius et ad mortem usque lassata est.
JUDG|16|17|Tunc aperiens ei totum cor suum dixit ad eam: " Novacula numquam ascendit super caput meum, quia nazaraeus consecratus Deo sum de utero matris meae; si rasum fuerit caput meum, recedet a me fortitudo mea, et deficiam eroque ut ceteri homines ".
JUDG|16|18|Videns illa quod confessus ei esset omnem animum suum, misit ad principes Philisthinorum atque mandavit: " Ascendite adhuc semel, quia nunc mihi aperuit totum cor suum ". Qui ascenderunt, assumpta pecunia, quam promiserant.
JUDG|16|19|At illa dormire eum fecit super genua sua vocavitque tonsorem et fecit radere septem crines eius et coepit humiliare eum; statim enim ab eo fortitudo discessit.
JUDG|16|20|Dixitque: " Philisthim super te, Samson! ". Qui de somno consurgens dixit in animo suo: " Egrediar, sicut ante feci, et me excutiam ", nesciens quod Dominus recessisset ab eo.
JUDG|16|21|Quem cum apprehendissent Philisthim, statim eruerunt oculos eius et duxerunt Gazam vinctum duabus catenis aeneis et clausum in carcere molere fecerunt.
JUDG|16|22|Iamque capilli eius renasci coeperant, postquam rasi sunt.
JUDG|16|23|Principes autem Philisthinorum convenerunt in unum, ut immolarent hostias magnificas Dagon deo suo et epularentur dicentes: Tradidit deus nosterin manus nostrasinimicum nostrum Samson ".
JUDG|16|24|Quem etiam populus videns laudabat deum suum eademque dicebat: Tradidit deus noster in manus nostrasadversarium nostrum,qui vastavit terram nostramet occidit plurimos nostrum ".
JUDG|16|25|Cum enim iam hilariores essent, postulaverunt, ut vocaretur Samson et ante eos luderet. Qui adductus de carcere ludebat ante eos; feceruntque eum stare inter duas columnas.
JUDG|16|26|Qui dixit puero tenenti manum suam: " Dimitte me, ut tangam columnas, quibus imminet domus, et recliner super eas et paululum requiescam ".
JUDG|16|27|Domus autem plena erat virorum ac mulierum; et erant ibi omnes principes Philisthinorum, ac de tecto circiter tria milia utriusque sexus spectabant ludentem Samson.
JUDG|16|28|At ille invocavit Dominum dicens: " Domine Deus, memento mei! Et redde mihi tantum hac vice fortitudinem pristinam, Deus, ut ulciscar me de Philisthim saltem pro uno duorum luminum meorum! ".
JUDG|16|29|Et tangens ambas columnas medias, quibus innitebatur domus, obnixusque contra alteram earum dextera et contra alteram laeva
JUDG|16|30|ait: " Moriatur anima mea cum Philisthim! ". Concussisque fortiter columnis, cecidit domus super omnes principes et ceteram multitudinem, quae ibi erat; multoque plures interfecit moriens, quam ante vivus occiderat.
JUDG|16|31|Descendentes autem fratres eius et universa cognatio tulerunt corpus eius et sepelierunt inter Saraa et Esthaol in sepulcro patris sui Manue; iudicavitque Israel viginti annis.
JUDG|17|1|Fuit vir quidam de monte Ephraim nomine Michas,
JUDG|17|2|qui dixit matri suae: " Mille centum argenteos, qui ablati sunt a te et super quibus, me audiente, maledicens iuraveras, ecce ego habeo; ego abstuli ". Cui illa respondit: " Benedictus filius meus Domino! ".
JUDG|17|3|Reddidit ergo eos matri suae, quae dixit ei: " Consecravi et vovi argentum hoc Domino: de manu mea suscipiat pro filio meo, ut faciat sculptile atque conflatile. Et nunc trado illud tibi ".
JUDG|17|4|Reddiditque eos matri suae, quae tulit ducentos argenteos et dedit eos argentario, ut faceret ex eis sculptile atque conflatile, quod fuit in domo Michae,
JUDG|17|5|qui aediculam Dei habens fecit ephod ac theraphim implevitque unius filiorum suorum manum, et factus est ei sacerdos.
JUDG|17|6|In diebus illis non erat rex in Israel, sed unusquisque, quod sibi rectum videbatur, hoc faciebat.
JUDG|17|7|Fuit quoque adulescens de Bethlehem Iudae ex cognatione Iudae; eratque ipse Levites et habitabat ibi ut advena.
JUDG|17|8|Egressusque de civitate Bethlehem peregrinari voluit ubicumque sibi commodum repperisset. Cumque iter faciens venisset in monte Ephraim usque ad domum Michae,
JUDG|17|9|interrogatus est ab eo unde venisset. Qui respondit: " Levita sum de Bethlehem Iudae et vado, ut habitem, ubi potuero et utile mihi esse perspexero ".
JUDG|17|10|Dixitque Michas: " Mane apud me et esto mihi parens ac sacerdos; daboque tibi per annos singulos decem argenteos ac vestium apparatum et quae ad victum sunt necessaria ".
JUDG|17|11|Acquievit et mansit apud hominem fuitque illi quasi unus de filiis.
JUDG|17|12|Implevitque Michas manum eius et habuit puerum sacerdotem apud se,
JUDG|17|13|" nunc scio, dicens, quod benefaciet mihi Dominus habenti levitici generis sacerdotem ".
JUDG|18|1|In diebus illis non erat rex in Israel, et tribus Dan quaere bat possessionem sibi, ut habitaret in ea; usque ad illum enim diem inter ceteras tribus sortem non acceperat.
JUDG|18|2|Miserunt igitur filii Dan stirpis et familiae suae quinque viros fortissimos de Saraa et Esthaol, ut explorarent terram et diligenter inspicerent, dixeruntque eis: " Ite et considerate terram ". Qui cum venissent in montem Ephraim usque ad domum Michae, pernoctaverunt ibi.
JUDG|18|3|Cum essent prope domum Michae, agnoscentes vocem adulescentis Levitae declinaverant illuc dicentes ad eum: " Quis te huc adduxit? Quid hic agis? Quam ob causam huc venire voluisti? ".
JUDG|18|4|Qui respondit eis: " Haec et haec praestitit mihi Michas et me mercede conduxit, ut sim ei sacerdos ".
JUDG|18|5|Rogaveruntque eum, ut consuleret Deum, ut scire possent an prospero itinere pergerent, et res haberet effectum.
JUDG|18|6|Qui respondit eis: " Ite cum pace; Dominus respicit viam vestram et iter, quo pergitis ".
JUDG|18|7|Euntes itaque quinque viri venerunt Lais videruntque populum habitantem in ea absque ullo timore iuxta Sidoniorum consuetudinem, securum et quietum, nullo eis penitus resistente, magnarumque opum et procul a Sidoniis neque in societate cum Syria.
JUDG|18|8|Reversique ad fratres suos in Saraa et Esthaol et quid egissent sciscitantibus, responderunt:
JUDG|18|9|" Surgite, et ascendamus adversus eos. Vidimus enim terram valde opulentam et uberem, et vos neglegetis? Nolite cessare; eamus et possideamus eam.
JUDG|18|10|Intrabimus ad securos in regionem latissimam; tradetque nobis Deus locum, in quo nullius rei est penuria eorum, quae sunt in terra ".
JUDG|18|11|Profecti igitur sunt de cognatione Dan, de Saraa et Esthaol, sescenti viri accincti armis bellicis.
JUDG|18|12|Ascendentesque castrametati sunt in Cariathiarim Iudae, qui locus ex eo tempore Castrorum Dan nomen accepit et est post tergum Cariathiarim.
JUDG|18|13|Inde transierunt in montem Ephraim.Cumque venissent usque ad domum Michae,
JUDG|18|14|dixerunt quinque viri, qui prius missi fuerant ad considerandam terram Lais, fratribus suis: " Nostis quod in domibus istis sit ephod et theraphim et sculptile atque conflatile? Videte quid vobis placeat, ut faciatis ".
JUDG|18|15|Et, cum paululum declinassent, ingressi sunt domum adulescentis Levitae, domum Michae, salutaveruntque eum verbis pacificis.
JUDG|18|16|Sescenti autem viri, ita ut erant armati, stabant ante ostium.
JUDG|18|17|At illi, qui ingressi fuerant domum iuvenis, sculptile et ephod et theraphim atque conflatile tulerunt; et sacerdos stabat ante ostium et sescenti viri armati.
JUDG|18|18|Tulerunt igitur, qui intraverant domum, sculptile, ephod et theraphim atque conflatile. Quibus dixit sacerdos: " Quid facitis? ".
JUDG|18|19|Cui responderunt: " Tace et pone digitum super os tuum venique nobiscum, ut habeamus te patrem et sacerdotem. Quid tibi melius est, ut sis sacerdos in domo unius viri, an in una tribu et familia in Israel? ".
JUDG|18|20|Et gavisus est sacerdos tulitque ephod et theraphim ac sculptile et profectus est in medio populi.
JUDG|18|21|Qui cum pergerent et ante se ire fecissent parvulos et iumenta et omne, quod erat pretiosum,
JUDG|18|22|iamque a domo Michae essent procul, viri, qui habitabant in aedibus prope domum Michae, convocati secuti sunt filios Dan
JUDG|18|23|et post tergum clamare coeperunt. Qui cum respexissent, dixerunt ad Micham: " Quid tibi vis? Cur concurritis? ".
JUDG|18|24|Qui respondit: " Deos meos, quos mihi feci, tulistis, et sacerdotem et omnia, quae habeo, et dicitis: "Quid tibi est?" ".
JUDG|18|25|Dixeruntque ei filii Dan: " Cave, ne ultra loquaris ad nos, et irruant in te viri animo concitati, et ipse cum omni domo tua pereas ".
JUDG|18|26|Et sic, coepto itinere, perrexerunt. Videns autem Michas quod fortiores se essent, reversus est in domum suam.
JUDG|18|27|Sescenti autem viri tulerunt, quod Michas fecerat, et sacerdotem eius veneruntque in Lais ad populum quiescentem atque securum et percusserunt eos in ore gladii urbemque incendio tradiderunt,
JUDG|18|28|nullo penitus ferente praesidium, eo quod procul habitarent a Sidone neque cum Syria haberent quidquam societatis ac negotii.Erat autem civitas sita in regione Rohob; quam rursum exstruentes habitaverunt in ea,
JUDG|18|29|vocato nomine civitatis Dan iuxta vocabulum patris sui, quem genuerat Israel, quae prius Lais dicebatur.
JUDG|18|30|Posueruntque sibi sculptile; et Ionathan filius Gersam filii Moysi ac filii eius sacerdotes erant in tribu Dan usque ad diem captivitatis terrae;
JUDG|18|31|mansitque apud eos idolum Michae omni tempore, quo fuit domus Dei in Silo.
JUDG|18|32|In diebus illis non erat rex in Israel.
JUDG|19|1|Fuit quidam vir Levi tes habitans ut advena in extrema parte montis Ephraim, qui accepit concubinam de Bethlehem Iudae.
JUDG|19|2|Quae irritata reversa est in domum patris sui in Bethlehem mansitque apud eum quattuor mensibus.
JUDG|19|3|Secutusque est eam vir suus volens loqui ad cor eius et secum reducere habens in comitatu puerum et duos asinos. Quae suscepit eum et introduxit in domum patris sui. Quem cum socer eius vidisset, occurrit ei laetus
JUDG|19|4|et retinuit hominem. Mansitque gener in domo soceri tribus diebus comedens cum eo et bibens familiariter.
JUDG|19|5|Die autem quarto, cum de nocte consurrexissent, et ille proficisci vellet, socer ait ad eum: " Gusta prius pauxillum panis et conforta cor tuum et sic proficisceris ".
JUDG|19|6|Sederuntque ambo simul et comederunt ac biberunt. Dixitque pater puellae ad generum suum: " Quaeso te, ut hodie hic maneas, pariterque laetemur ".
JUDG|19|7|At ille consurgens coepit velle proficisci. Et nihilominus obnixe eum socer tenuit et apud se fecit manere.
JUDG|19|8|Mane autem facto, quinta die parabat Levites iter; cui socer rursum: " Oro te, inquit, ut confortes cor tuum". Et tardabant, donec declinaret dies; et ambo comederunt simul.
JUDG|19|9|Surrexitque adulescens, ut pergeret cum uxore sua et puero. Cui rursum locutus est socer eius pater puellae: " Considera quod dies ad occasum declivior sit et propinquet ad vesperum; manete apud me etiam hodie, pernocta hic et esto laeto animo, et cras mane proficiscemini, ut vadas in domum tuam ".
JUDG|19|10|Noluit gener acquiescere sermonibus eius, sed statim perrexit et venit contra Iebus, id est Ierusalem, ducens secum duos asinos onustos et concubinam.
JUDG|19|11|Iamque aderant iuxta Iebus, et dies mutabatur in noctem; dixitque puer ad dominum suum: " Veni, obsecro, declinemus ad urbem Iebusaeorum et maneamus in ea ".
JUDG|19|12|Cui respondit dominus: " Non ingrediamur oppidum gentis alienae, quae non est de filiis Israel, sed transibimus usque Gabaa ".
JUDG|19|13|Dixitque puero suo: "Veni, accedamus ad unum de locis et manebimus in Gabaa aut Rama ".
JUDG|19|14|Transierunt igitur Iebus et coeptum carpebant iter; occubuitque eis sol iuxta Gabaa, quae est in tribu Beniamin.
JUDG|19|15|Diverteruntque ad eam, ut manerent ibi; quo cum intrassent, sedebant in platea civitatis, et nullus eos recipere volebat hospitio.
JUDG|19|16|Et ecce apparuit homo senex revertens de agro et de opere suo vespere, qui et ipse erat de monte Ephraim et peregrinus habitabat in Gabaa; homines autem loci illius erant de tribu Beniamin.
JUDG|19|17|Elevatisque oculis, vidit senex sedentem hominem viatorem in platea civitatis et dixit ad eum: " Unde venis et quo vadis? ".
JUDG|19|18|Qui respondit ei: " Profecti sumus de Bethlehem Iudae et pergimus ad locum meum, qui est in extrema parte montis Ephraim, unde profectus sum in Bethlehem. Et nunc vado ad domum meam, nullusque sub tectum suum me vult recipere
JUDG|19|19|habentem paleas et pabulum pro asinis nostris et panem ac vinum in meos et ancillae tuae usus et pueri, qui cum servo tuo sunt; nulla re indigemus nisi hospitio ".
JUDG|19|20|Cui respondit senex: " Pax tecum sit! Ego praebebo omnia, quae necessaria sunt; tantum, quaeso, ne in platea maneas ".
JUDG|19|21|Introduxitque eum in domum suam et commixtum migma asinis praebuit; ac, postquam laverunt pedes suos, recepit eos in convivium.
JUDG|19|22|Illis laeto corde epulantibus, venerunt viri civitatis illius filii Belial et circumdantes domum senis fores pulsare coeperunt clamantes ad dominum domus atque dicentes: " Educ virum, qui ingressus est domum tuam, ut abutamur eo ".
JUDG|19|23|Egressusque est ad eos senex et ait: " Nolite, fratres, nolite facere malum hoc, quia ingressus est homo hospitium meum, et cessate ab hac stultitia.
JUDG|19|24|Habeo filiam virginem, et hic homo habet concubinam; educam eas ad vos, ut humilietis eas et faciatis eis, quod vobis placuerit; tantum, obsecro, ne scelus hoc operemini in virum ".
JUDG|19|25|Nolebant acquiescere sermonibus eius; quod cernens homo apprehendit et eduxit ad eos concubinam suam. Qua cum abusi essent et tota nocte ei illusissent, dimiserunt eam mane.
JUDG|19|26|At mulier, recedentibus tenebris, venit ad ostium domus, ubi manebat dominus suus, et ibi corruit.
JUDG|19|27|Mane facto surrexit homo et aperuit ostium, ut coeptam expleret viam; et ecce concubina eius iacebat ante ostium, sparsis in limine manibus.
JUDG|19|28|Cui ille loquebatur: " Surge, ut ambulemus ". Qua nihil respondente, intellegens quod erat mortua, tulit eam et imposuit asino; reversusque est in domum suam.
JUDG|19|29|Quam cum esset ingressus, arripuit gladium et cadaver uxoris secundum ossa sua in duodecim partes ac frusta concidens misit in omnes terminos Israel.
JUDG|19|30|Quod cum vidissent singuli, conclamabant: " Numquam res talis facta et visa est in Israel ex eo die, quo ascenderunt patres nostri de Aegypto, usque in praesens tempus! ". Praeceperat enim viris, quos miserat, dicens: Haec dicite omni viro Israel: Si factum est quidquam tale ex die, quo ascenderunt filii Israel de terra Aegypti, usque ad praesentem diem? Attendite ad hoc, consiliamini et decernite quid facto opus sit!".
JUDG|20|1|Egressi sunt itaque omnes fi lii Israel et pariter congrega ti, quasi vir unus, de Dan usque Bersabee et terra Galaad ad Dominum in Maspha.
JUDG|20|2|Omnisque populi anguli et cunctae tribus Israel in ecclesiam populi Dei convenerunt: quadringenta milia peditum pugnatorum.
JUDG|20|3|Nec latuit filios Beniamin, quod ascendissent filii Israel in Maspha. Interrogatusque Levita maritus mulieris interfectae quo modo tantum scelus perpetratum esset,
JUDG|20|4|respondit: " Veni in Gabaa Beniamin cum uxore mea illucque diverti.
JUDG|20|5|Et ecce homines civitatis illius circumdederunt nocte domum, in qua manebam, volentes me occidere et uxorem meam incredibili libidinis furore vexantes; denique mortua est.
JUDG|20|6|Quam arreptam in frusta concidi misique partes in omnes terminos possessionis Israel, quia fecerunt nefas et piaculum in Israel.
JUDG|20|7|Adestis omnes, filii Israel: decernite quid facere debeatis ".
JUDG|20|8|Stansque omnis populus quasi unius hominis sermone respondit: " Non recedemus in tabernacula nostra, nec suam quisquam intrabit domum,
JUDG|20|9|sed hoc contra Gabaa in commune faciemus secundum sortem:
JUDG|20|10|decem viri eligantur e centum ex omnibus tribubus Israel et centum de mille et mille de decem milibus, ut comportent exercitui cibaria illis, qui venerunt, ut reddant Gabaa Beniamin pro scelere, quod meretur ".
JUDG|20|11|Convenitque universus Israel ad civitatem quasi unus homo, eadem mente unoque consilio,
JUDG|20|12|et miserunt nuntios ad omnem tribum Beniamin, qui dicerent: " Quale nefas in vobis repertum est!
JUDG|20|13|Tradite homines filios Belial in Gabaa, qui hoc flagitium perpetrarunt, ut moriantur, et auferatur malum de Israel ".Qui noluerunt fratrum suorum filiorum Israel audire mandatum,
JUDG|20|14|sed ex cunctis urbibus, quae suae sortis erant, convenerunt in Gabaa, ut illis ferrent auxilium et contra universum Israel populum dimicarent.
JUDG|20|15|Recensitique sunt in die illa viginti sex milia de civitatibus Beniamin educentium gladium, praeter habitatores Gabaa, qui septingenti erant viri fortissimi.
JUDG|20|16|In universo hoc populo erant septingenti viri electi, qui sinistra pro dextra utebantur et sic fundis lapides ad certum iaciebant, ut capillum quoque possent percutere, et nequaquam in alteram partem ictus lapidis deferretur.
JUDG|20|17|Virorum quoque Israel, absque filiis Beniamin, recensita sunt quadringenta milia educentium gladios et paratorum ad pugnam.
JUDG|20|18|Qui surgentes venerunt in Bethel consulueruntque Deum atque dixerunt: " Quis erit in exercitu nostro princeps certaminis contra filios Beniamin?. Quibus respondit Dominus: " Iuda ascendet primus ".
JUDG|20|19|Statimque filii Israel surgentes mane castrametati sunt contra Gabaa;
JUDG|20|20|et inde procedentes ad pugnam contra Beniamin, contra urbem aciem direxerunt.
JUDG|20|21|Egressique filii Beniamin de Gabaa occiderunt de filiis Israel die illo viginti duo milia viros.
JUDG|20|22|Rursum filii Israel confortati in eodem loco, in quo prius certaverant, aciem direxerunt,
JUDG|20|23|ita tamen ut prius ascenderent et flerent coram Domino usque ad noctem consulerentque eum et dicerent: " Debeo ultra procedere ad dimicandum contra filios Beniamin fratres meos, an non? ". Quibus ille respondit: " Ascendite ad eos ".
JUDG|20|24|Cumque filii Israel altero die contra filios Beniamin ad proelium processissent,
JUDG|20|25|eruperunt filii Beniamin de Gabaa et occurrentes eis iterum decem et octo milia virorum educentium gladium prostraverunt.
JUDG|20|26|Quam ob rem omnes filii Israel, universus populus, venerunt in Bethel et sedentes flebant coram Domino ieiunaveruntque die illo usque ad vesperam et obtulerunt ei holocausta et pacificas victimas
JUDG|20|27|et super statu suo interrogaverunt. Eo tempore ibi erat arca foederis Dei,
JUDG|20|28|et Phinees filius Eleazari filii Aaron stabat coram eo. Consuluerunt igitur Dominum atque dixerunt: " Exire ultra debemus ad pugnam contra filios Beniamin fratres nostros, an quiescere? ". Quibus ait Dominus: " Ascendite, cras enim tradam eos in manus vestras ".
JUDG|20|29|Posueruntque filii Israel insidias per circuitum urbis Gabaa
JUDG|20|30|et tertia vice sicut semel et bis contra Beniamin et Gabaa exercitum produxerunt.
JUDG|20|31|Sed et filii Beniamin eruperunt in occursum populi et abstracti de civitate coeperunt caedere ex eis sicut primo et secundo die, per duas semitas terga vertentes, quarum una ferebat in Bethel, altera in Gabaa, atque prosternere in campo triginta circiter viros.
JUDG|20|32|Putaverunt enim solito eos more percussos cedere; qui fugam simulaverunt, ut abstraherent eos de civitate et quasi fugientes ad supradictas semitas perducerent.
JUDG|20|33|Omnes itaque viri Israel surgentes de sedibus suis tetenderunt aciem in loco, qui vocatur Baalthamar. Insidiae quoque eruperunt de loco suo, de regione in occidente Gabaa.
JUDG|20|34|Venerunt ergo adversus Gabaa decem milia virorum electorum de universo Israel. Ingravatumque est bellum contra filios Beniamin, et non intellexerunt quod ex omni parte illis instaret interitus.
JUDG|20|35|Percussitque eos Dominus in conspectu filiorum Israel, et interfecerunt ex eis in illo die viginti quinque milia et centum viros, omnes bellatores et educentes gladium.
JUDG|20|36|Filii autem Beniamin, cum se inferiores esse vidissent, coeperunt fugere. Quod cernentes filii Israel, dederunt eis ad fugiendum locum, quia confidebant in insidiis, quas iuxta urbem posuerant.
JUDG|20|37|Qui cum repente de latibulis surrexissent, irruerunt super Gabaa et ingressi celeriter percusserunt totam civitatem in ore gladii.
JUDG|20|38|Signum autem dederant filii Israel his, quos in insidiis collocaverant, ut ignem accenderent et, ascendente in altum fumo, captam urbem demonstrarent.
JUDG|20|39|Verterant ergo terga filii Israel in ipso certamine positi, et filii Beniamin putantes quod percussissent eos sicut in priore pugna, coeperant de exercitu eorum caedere triginta fere viros.
JUDG|20|40|Cum autem columna fumi de civitate conscendere coepisset, et Beniamin quoque retro aspiciens cerneret de civitate flammas in sublime ferri,
JUDG|20|41|cumque vir Israel versa facie aggrederetur, vir Beniamin conturbatus est, quia vidit se apprehensum a malo.
JUDG|20|42|Et ad viam deserti ire coeperunt, illuc quoque eos adversariis persequentibus. Sed et hi, qui urbem succenderant, occurrerunt eis,
JUDG|20|43|atque ita factum est ut ex utraque parte ab hostibus caederentur, nec erat eis ulla requies. Prostrati sunt usque ad orientalem plagam urbis Gabaa.
JUDG|20|44|Fuerunt autem, qui interfecti sunt de Beniamin, decem et octo milia virorum omnes robustissimi pugnatores.
JUDG|20|45|Qui remanserant, fugerunt in solitudinem et pergebant ad petram, cuius vocabulum est Remmon. Quasi racemos colligentes occiderunt in viis quinque milia viros. Et cum instantius eos persequerentur usque Gadaam, interfecerunt etiam alios duo milia.
JUDG|20|46|Et sic factum est ut omnes, qui ceciderant de Beniamin in die illa, essent viginti quinque milia pugnatores ad bella promptissimi.
JUDG|20|47|Remanserunt itaque, qui evadere potuerant et fugere in solitudinem, sescenti viri; sederuntque in petra Remmon mensibus quattuor.
JUDG|20|48|Regressi autem filii Israel ex civitatibus a viris usque ad iumenta, usque ad omne, quod inveniri poterat, gladio percusserunt, cunctasque urbes et viculos Beniamin vorax flamma consumpsit.
JUDG|21|1|Iuraverunt autem filii Israel in Maspha et dixerunt: " Nullus nostrum dabit filiis Beniamin de filiabus suis uxorem ".
JUDG|21|2|Venitque populus in Bethel, et in conspectu Dei sedentes usque ad vesperam levaverunt vocem et magno ululatu coeperunt flere dicentes:
JUDG|21|3|" Quare, Domine, Deus Israel, factum est hoc in populo tuo, ut hodie una tribus auferretur de Israel? ".
JUDG|21|4|Altera autem die diluculo consurgentes exstruxerunt altare obtuleruntque ibi holocausta et pacificas victimas
JUDG|21|5|et dixerunt: " Quis non ascendit in congregationem ad Dominum de universis tribubus Israel? ". Grandi enim se iuramento constrinxerant interfici eos, qui non ascendissent ad Dominum in Maspha.
JUDG|21|6|Ductique paenitentia filii Israel super fratre suo Beniamin coeperunt dicere: " Ablata est hodie una tribus de Israel.
JUDG|21|7|Quid faciemus, ut, qui remanserunt, uxores accipiant? Omnes enim in commune iuravimus per Dominum non daturos nos his filias nostras ".
JUDG|21|8|Idcirco dixerunt: " Quis est de universis tribubus Israel, qui non ascendit ad Dominum in Maspha? ". Et ecce nemo de Iabes Galaad in castra venerat ad congregationem,
JUDG|21|9|et, cum populus recenseretur, nullus ex eis repertus est.
JUDG|21|10|Misit itaque coetus decem milia viros robustissimos et praeceperunt eis: " Ite et percutite habitatores Iabes Galaad in ore gladii tam uxores quam parvulos eorum.
JUDG|21|11|Et hoc erit, quod observare debetis: Omne generis masculini et mulieres, quae cognoverunt viros, interficite; virgines autem reservate ".
JUDG|21|12|Inventaeque sunt de Iabes Galaad quadringentae virgines, quae nescierunt viri torum, et adduxerunt eas in castra in Silo in terra Chanaan.
JUDG|21|13|Misitque coetus nuntios ad filios Beniamin, qui erant in petra Remmon, et dederunt eis pacem.
JUDG|21|14|Veneruntque filii Beniamin in illo tempore, et datae sunt eis uxores de filiabus Iabes Galaad; alias autem non reppererunt, quas simili modo traderent.
JUDG|21|15|Populusque valde doluit de Beniamin, quia fecerat Dominus confractionem in tribubus Israel.
JUDG|21|16|Dixeruntque seniores coetus: " Quid faciemus reliquis, qui non acceperunt uxores? Omnes in Beniamin feminae conciderunt ".
JUDG|21|17|Et dixerunt: " Possessio eorum, qui effugerunt, erit Beniamin, ne una tribus deleatur ex Israel.
JUDG|21|18|Filias autem nostras eis dare non possumus, constricti hoc iuramento: Maledictus, qui dederit de filiabus suis uxorem Beniamin!" ".
JUDG|21|19|Ceperuntque consilium atque dixerunt: " Ecce sollemnitas Domini est in Silo anniversaria, quae sita est ad septentrionem urbis Bethel et ad orientalem plagam viae, quae de Bethel tendit ad Sichimam et ad meridiem oppidi Lebona ".
JUDG|21|20|Praeceperuntque filiis Beniamin atque dixerunt: "Ite et latitate in vineis;
JUDG|21|21|cumque videritis filias Silo ad ducendos choros ex more procedere, exite repente de vineis et rapite ex eis singuli uxores singulas et pergite in terram Beniamin ".
JUDG|21|22|Cumque venerint patres earum ac fratres et apud nos queri coeperint, dicemus eis: " Miseremini nostri et eorum; non enim acceperunt unusquisque uxorem in bello, et vos, si dedissetis eis, deliquissetis ".
JUDG|21|23|Feceruntque filii Beniamin, ut sibi fuerat imperatum, et iuxta numerum suum rapuerunt sibi de his, quae ducebant choros, uxores singulas; abieruntque in possessionem suam aedificantes urbes et habitantes in eis.
JUDG|21|24|Filii quoque Israel reversi sunt inde illo tempore unusquisque ad tribum et familiam suam in possessionem suam.
JUDG|21|25|In diebus illis non erat rex in Israel, sed unusquisque, quod sibi rectum videbatur, hoc faciebat.
