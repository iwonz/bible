2KGS|1|1|Praevaricatus est autem Moab in Israel, postquam mortuus est Achab.
2KGS|1|2|Ceciditque Ochozias per cancellos cenaculi sui, quod habebat in Samaria, et aegrotavit; misitque nuntios dicens ad eos: " Ite, consulite Beelzebub deum Accaron, utrum vivere queam de infirmitate mea hac ".
2KGS|1|3|Angelus autem Domini locutus est ad Eliam Thesbiten: " Surge, ascende in occursum nuntiorum regis Samariae et dices ad eos: Numquid non est Deus in Israel, ut eatis ad consulendum Beelzebub deum Accaron?
2KGS|1|4|Quam ob rem haec dicit Dominus: De lectulo, super quem ascendisti, non descendes, sed morte morieris ". Et abiit Elias.
2KGS|1|5|Reversique sunt nuntii ad Ochoziam, qui dixit eis: " Quare reversi estis? ".
2KGS|1|6|At illi responderunt ei: " Vir occurrit nobis et dixit ad nos: "Ite, revertimini ad regem, qui misit vos, et dicetis ei: Haec dicit Dominus: Numquid, quia non est Deus in Israel, mittis, ut consulatur Beelzebub deus Accaron? Idcirco de lectulo, super quem ascendisti, non descendes, sed morte morieris" ".
2KGS|1|7|Qui dixit eis: " Cuius figurae et habitus vir erat, qui occurrit vobis et locutus est verba haec? ".
2KGS|1|8|At illi dixerunt: " Vir in veste pilosa et zona pellicea accinctis renibus ". Qui ait: " Elias Thesbites est ".
2KGS|1|9|Misitque ad eum quinquagenarium principem et quinquaginta, qui erant sub eo; qui ascendit ad eum sedentique in vertice montis ait: " Homo Dei, rex praecepit, ut descendas ".
2KGS|1|10|Respondensque Elias dixit quinquagenario: " Si homo Dei sum, descendat ignis e caelo et devoret te et quinquaginta tuos ". Descendit itaque ignis e caelo et devoravit eum et quinquaginta, qui erant cum eo.
2KGS|1|11|Rursum misit ad eum principem quinquagenarium alterum et quinquaginta cum eo; qui locutus est illi: " Homo Dei, haec dicit rex: "Festina, descende!" ".
2KGS|1|12|Respondens Elias ait illis: " Si homo Dei ego sum, descendat ignis e caelo et devoret te et quinquaginta tuos ". Descendit ergo ignis Dei e caelo et devoravit illum et quinquaginta eius.
2KGS|1|13|Iterum misit principem quinquagenarium tertium et quinquaginta, qui erant cum eo; qui cum venisset, curvavit genua contra Eliam et precatus est eum et ait: " Homo Dei, noli despicere animam meam et animam servorum tuorum, qui mecum sunt.
2KGS|1|14|Ecce descendit ignis de caelo et devoravit duos principes quinquagenarios primos et quinquagenos, qui cum eis erant; sed nunc obsecro, ut miserearis animae meae ".
2KGS|1|15|Locutus est autem angelus Domini ad Eliam dicens: " Descende cum eo, ne timeas ". Surrexit igitur et descendit cum eo ad regem
2KGS|1|16|et locutus est ei: " Haec dicit Dominus: Quia misisti nuntios ad consulendum Beelzebub deum Accaron, quasi non esset Deus in Israel, a quo posses interrogare sermonem, ideo de lectulo, super quem ascendisti, non descendes, sed morte morieris ".
2KGS|1|17|Mortuus est ergo iuxta sermonem Domini, quem locutus est Elias. Et regnavit Ioram frater eius pro eo anno secundo Ioram filii Iosaphat regis Iudae; non enim habebat filium.
2KGS|1|18|Reliqua autem gestorum Ochoziae, quae operatus est, nonne haec scripta sunt in libro annalium regum Israel?
2KGS|2|1|Factum est autem cum levare vellet Dominus Eliam per turbi nem in caelum, ibant Elias et Eliseus de Galgalis;
2KGS|2|2|dixitque Elias ad Eliseum: " Sede hic, quia Dominus misit me usque Bethel ". Cui ait Eliseus: " Vivit Dominus, et vivit anima tua, quia non derelinquam te ". Cumque descendissent Bethel,
2KGS|2|3|egressi sunt filii prophetarum, qui erant in Bethel, ad Eliseum et dixerunt ei: "Numquid nosti quia hodie Dominus tollat dominum tuum desuper capite tuo? ". Qui respondit: " Et ego novi, silete ".
2KGS|2|4|Dixit autem ei Elias: " Elisee, sede hic, quia Dominus misit me in Iericho ". Et ille ait: " Vivit Dominus, et vivit anima tua, quia non derelinquam te ". Cumque venissent Ierichum,
2KGS|2|5|accesserunt filii prophetarum, qui erant in Iericho, ad Eliseum et dixerunt ei: " Numquid nosti quia hodie Dominus tollet dominum tuum desuper capite tuo? ". Et ait: " Et ego novi, silete ".
2KGS|2|6|Dixit autem ei Elias: " Sede hic, quia Dominus misit me ad Iordanem ". Qui ait: " Vivit Dominus, et vivit anima tua, quia non derelinquam te ". Ierunt igitur ambo pariter,
2KGS|2|7|et quinquaginta viri de filiis prophetarum secuti sunt, qui et steterunt e contra longe. Illi autem ambo stabant super Iordanem.
2KGS|2|8|Tulitque Elias pallium suum et involvit illud et percussit aquas, quae divisae sunt in utramque partem, et transierunt ambo per siccum.
2KGS|2|9|Cumque transissent, Elias dixit ad Eliseum: " Postula, quod vis, ut faciam tibi, antequam tollar a te ". Dixitque Eliseus: " Obsecro, ut fiant duae partes spiritus tui in me ".
2KGS|2|10|Qui respondit: " Rem difficilem postulasti. Attamen si videris me, quando tollor a te, erit tibi, quod petisti; si autem non videris, non erit ".
2KGS|2|11|Cumque pergerent et incedentes sermocinarentur, ecce currus igneus et equi ignei diviserunt utrumque; et ascendit Elias per turbinem in caelum.
2KGS|2|12|Eliseus autem videbat et clamabat: " Pater mi, pater mi, currus Israel et auriga eius! ". Et non vidit eum amplius; apprehenditque vestimenta sua et scidit illa in duas partes.
2KGS|2|13|Et levavit pallium Eliae, quod ceciderat ei, reversusque stetit super ripam Iordanis.
2KGS|2|14|Et pallio Eliae, quod ceciderat ei, percussit aquas et dixit: " Ubi est Deus Eliae etiam nunc? ". Percussitque aquas, et divisae sunt huc atque illuc, et transiit Eliseus.
2KGS|2|15|Videntes autem filii prophetarum, qui erant in Iericho de contra, dixerunt: " Requievit spiritus Eliae super Eliseum ". Et venientes in occursum eius adoraverunt eum proni in terram
2KGS|2|16|dixeruntque illi: " Ecce cum servis tuis sunt quinquaginta viri fortes, qui possunt ire et quaerere dominum tuum, ne forte tulerit eum spiritus Domini et proiecerit in uno montium aut in una vallium ". Qui ait: " Nolite mittere! ".
2KGS|2|17|Coegeruntque eum, donec acquiesceret et diceret: " Mittite ". Et miserunt quinquaginta viros. Qui cum quaesissent tribus diebus, non invenerunt
2KGS|2|18|et reversi sunt ad eum. At ille habitabat in Iericho dixitque eis: " Numquid non dixi vobis: Nolite ire?".
2KGS|2|19|Dixerunt quoque viri civitatis ad Eliseum: " Ecce habitatio civitatis huius optima est, sicut tu ipse, domine, perspicis; sed aquae pessimae sunt, et terra faciens abortium ".
2KGS|2|20|At ille ait: "Afferte mihi vas novum et mittite in illud sal ". Qui cum attulissent,
2KGS|2|21|egressus ad fontem aquarum misit in eum sal et ait: " Haec dicit Dominus: Sanavi aquas has, et non erit ultra in eis mors neque abortium ".
2KGS|2|22|Sanatae sunt ergo aquae usque ad diem hanc iuxta verbum Elisei, quod locutus est.
2KGS|2|23|Ascendit autem inde Bethel. Cumque ascenderet per viam, pueri parvi egressi sunt de civitate et illudebant ei dicentes: "Ascende, calve; ascende, calve! ".
2KGS|2|24|Qui cum respexisset, vidit eos et maledixit eis in nomine Domini; egressique sunt duo ursi de saltu et laceraverunt ex eis quadraginta duos pueros.
2KGS|2|25|Abiit autem inde in montem Carmeli et inde reversus est Samariam.
2KGS|3|1|Ioram vero filius Achab regnavit super Israel in Samaria anno decimo octavo Iosaphat regis Iudae regnavitque duodecim annis.
2KGS|3|2|Et fecit malum coram Domino, sed non sicut pater suus et mater; tulit enim lapidem Baal, quem fecerat pater eius.
2KGS|3|3|Verumtamen in peccatis Ieroboam filii Nabat, qui peccare fecit Israel, adhaesit nec recessit ab eis.
2KGS|3|4|Porro Mesa rex Moab nutriebat pecora multa et solvebat regi Israel centum milia agnorum et lanam centum milium arietum.
2KGS|3|5|Cumque mortuus fuisset Achab, praevaricatus est foedus, quod habebat cum rege Israel.
2KGS|3|6|Egressus est igitur rex Ioram in die illa de Samaria et recensuit universum Israel;
2KGS|3|7|profectusque misit ad Iosaphat regem Iudae dicens: " Rex Moab recessit a me. Vis venire mecum contra Moab ad proelium? ". Qui respondit: " Ascendam. Qui meus est tuus est, populus meus populus tuus, equi mei equi tui ".
2KGS|3|8|Dixitque: " Per quam viam ascendemus? ". At ille respondit: " Per desertum Idumaeae ".
2KGS|3|9|Perrexerunt igitur rex Israel et rex Iudae et rex Edom et circuierunt per viam septem dierum; nec erat aqua exercitui et iumentis, quae sequebantur eos.
2KGS|3|10|Dixitque rex Israel: " Heu! Congregavit nos Dominus tres reges, ut traderet in manu Moab ".
2KGS|3|11|Et ait Iosaphat: " Estne hic propheta Domini, ut interrogemus Dominum per eum? ". Et respondit unus de servis regis Israel: " Est hic Eliseus filius Saphat, qui fundebat aquam super manus Eliae ".
2KGS|3|12|Et ait Iosaphat: " Est apud eum sermo Domini ". Descenditque ad eum rex Israel et Iosaphat et rex Edom.
2KGS|3|13|Dixit autem Eliseus ad regem Israel: " Quid mihi et tibi est? Vade ad prophetas patris tui et ad prophetas matris tuae ". Et ait illi rex Israel: "Non, congregavit enim Dominus tres reges hos, ut traderet eos in manu Moab? ".
2KGS|3|14|Dixit autem Eliseus: " Vivit Dominus exercituum, in cuius conspectu sto, quod si non vultum Iosaphat regis Iudae revererer, ne attendissem quidem te nec respexissem;
2KGS|3|15|nunc autem adducite mihi psaltem ". Cumque caneret psaltes, facta est super eum manus Domini,
2KGS|3|16|et ait: " Haec dicit Dominus: Facite in torrente hoc fossas et fossas.
2KGS|3|17|Haec enim dicit Dominus: Non videbitis ventum neque pluviam, et torrens replebitur aquis; et bibetis vos et pecora et iumenta vestra.
2KGS|3|18|Parumque hoc est in conspectu Domini; insuper tradet etiam Moab in manu vestra,
2KGS|3|19|et percutietis omnem civitatem munitam et omnem urbem electam et universum lignum fructiferum succidetis cunctosque fontes aquarum obturabitis et omnem agrum egregium operietis lapidibus ".
2KGS|3|20|Factum est igitur mane, quando sacrificium offerri solet, et ecce aquae veniebant per viam Edom. Et repleta est terra aquis.
2KGS|3|21|Universi autem Moabitae audientes quod ascendissent reges, ut pugnarent adversum eos, convocaverunt omnes, qui accingi poterant balteo et desuper, et steterunt in terminis.
2KGS|3|22|Primoque mane surgentes et, orto iam sole super aquis, viderunt Moabitae e contra aquas rubras quasi sanguinem
2KGS|3|23|dixeruntque: "Sanguis est gladii! Pugnaverunt reges contra se et caesi sunt mutuo. Nunc perge ad praedam, Moab! ".
2KGS|3|24|Perrexeruntque in castra Israel. Porro consurgens Israel percussit Moab, at illi fugerunt coram eis. Venerunt igitur subsequentes et percutientes Moab.
2KGS|3|25|Et civitates destruxerunt et omnem agrum optimum mittentes singuli lapides repleverunt; et universos fontes aquarum obturaverunt et omnia ligna fructifera succiderunt, ita ut muri tantum Cirhareseth remanerent; et circumdederunt civitatem fundibularii et aggressi sunt.
2KGS|3|26|Quod cum vidisset rex Moab, praevaluisse scilicet hostes, tulit secum septingentos viros educentes gladium, ut irrumperet ad regem Edom; et non potuerunt.
2KGS|3|27|Arripiensque filium suum primogenitum, qui regnaturus erat pro eo, obtulit holocaustum super murum. Et facta est indignatio magna super Israel; statimque recesserunt ab eo et reversi sunt in terram suam.
2KGS|4|1|Mulier autem quaedam de uxoribus filiorum prophetarum clamabat ad Eliseum dicens: " Servus tuus vir meus mortuus est, et tu nosti quia servus tuus fuit timens Dominum; et ecce creditor venit, ut tollat duos filios meos ad serviendum sibi ".
2KGS|4|2|Cui dixit Eliseus: " Quid vis, ut faciam tibi? Dic mihi: Quid habes in domo tua? ". At illa respondit: " Non habeo ancilla tua quidquam in domo mea, nisi vasculum olei ".
2KGS|4|3|Cui ait: " Vade, pete mutuo ab omnibus vicinis tuis vasa vacua non pauca;
2KGS|4|4|et ingredere et claude ostium, cum intrinsecus fueris tu et filii tui, et mitte inde in omnia vasa haec et, cum plena fuerint, tolles ".
2KGS|4|5|Ivit itaque mulier et clausit ostium super se et super filios suos; illi offerebant vasa, et illa infundebat.
2KGS|4|6|Cumque plena fuissent vasa, dixit ad filium suum: " Affer mihi adhuc vas. Et ille respondit: " Non habeo ". Stetitque oleum.
2KGS|4|7|Venit autem illa et indicavit homini Dei. Et ille: " Vade, inquit, vende oleum et redde creditori tuo; tu autem et filii tui vivite de reliquo ".
2KGS|4|8|Facta est autem quaedam dies, et transibat Eliseus per Sunam. Erat autem ibi mulier magna, quae tenuit eum, ut comederet panem. Quotiescumque inde transibat, divertebat ad eam, ut comederet panem.
2KGS|4|9|Quae dixit ad virum suum: " Animadverto quod vir Dei sanctus est iste, qui transit per nos frequenter.
2KGS|4|10|Faciamus ergo cenaculum muratum parvum et ponamus ei in eo lectulum et mensam et sellam et candelabrum, ut, cum venerit ad nos, maneat ibi ".
2KGS|4|11|Facta est ergo dies quaedam, et veniens divertit in cenaculum et requievit ibi.
2KGS|4|12|Dixitque ad Giezi puerum suum: " Voca Sunamitin istam ". Qui cum vocasset eam, et illa stetisset coram eo,
2KGS|4|13|dixit ad puerum: " Loquere ad eam: Ecce sedule in omnibus ministrasti nobis; quid vis, ut faciam tibi? Numquid habes negotium et vis, ut loquar regi sive principi militiae? ". Quae respondit: " In medio populi mei habito ".
2KGS|4|14|Et ait: " Quid ergo vult, ut faciam ei? ". Dixitque Giezi: "Ne quaeras; filium enim non habet, et vir eius senex est ".
2KGS|4|15|Praecepit itaque, ut vocaret eam; quae cum vocata fuisset et stetisset ad ostium,
2KGS|4|16|dixit ad eam: " In tempore isto, in anno altero, amplexaberis filium ". At illa respondit: " Noli, quaeso, domine mi, vir Dei, noli mentiri ancillae tuae ".
2KGS|4|17|Et concepit mulier et peperit filium in tempore isto anni alterius, quo dixerat Eliseus.
2KGS|4|18|Crevit autem puer et, cum esset quaedam dies, et egressus isset ad patrem suum, ad messores,
2KGS|4|19|ait patri suo: " Caput meum, caput meum! ". At ille dixit servo: " Tolle et duc eum ad matrem suam ".
2KGS|4|20|Qui cum tulisset et adduxisset eum ad matrem suam, posuit eum illa super genua sua usque ad meridiem, et mortuus est.
2KGS|4|21|Ascendit autem et collocavit eum super lectulum hominis Dei et clausit ostium; et egressa
2KGS|4|22|vocavit virum suum et ait: "Mitte mecum, obsecro, unum de pueris et asinam, ut excurram usque ad hominem Dei et revertar ".
2KGS|4|23|Qui ait illi: " Quam ob causam vadis ad eum hodie? Non sunt calendae neque sabbatum ". Quae respondit: " Vale ".
2KGS|4|24|Stravitque asinam et praecepit puero: " Mina et propera, ne mihi moram facias in eundo, nisi praecepero tibi ".
2KGS|4|25|Profecta est igitur et venit ad virum Dei in montem Carmeli. Cumque vidisset eam vir Dei de contra, ait ad Giezi puerum suum: " Ecce Sunamitis illa.
2KGS|4|26|Vade cito in occursum eius et dic ei: Rectene agitur circa te et circa virum tuum et circa filium tuum? ". Quae respondit: " Recte ".
2KGS|4|27|Cumque venisset ad virum Dei in monte, apprehendit pedes eius; et accessit Giezi, ut amoveret eam, et ait homo Dei: " Dimitte illam; anima enim eius in amaritudine est, et Dominus celavit me et non indicavit mihi.
2KGS|4|28|Quae dixit illi: " Numquid petivi filium a domino meo? Numquid non dixi tibi: Ne illudas me? ".
2KGS|4|29|Et ille ait ad Giezi: " Accinge lumbos tuos et tolle baculum meum in manu tua et vade. Si occurrerit tibi homo, non salutes eum et, si salutaverit te quispiam, non respondeas illi. Et pones baculum meum super faciem pueri ".
2KGS|4|30|Porro mater pueri ait: " Vivit Dominus, et vivit anima tua, non dimittam te ". Surrexit ergo et secutus est eam.
2KGS|4|31|Giezi autem praecesserat eos et posuerat baculum super faciem pueri, et non erat vox neque sensus reversusque est in occursum eius et nuntiavit ei dicens: " Non evigilavit puer ".
2KGS|4|32|Ingressus est ergo Eliseus domum, et ecce puer mortuus iacebat in lectulo eius;
2KGS|4|33|ingressusque clausit ostium super se et puerum et oravit ad Dominum.
2KGS|4|34|Et ascendit et incubuit super puerum posuitque os suum super os eius et oculos suos super oculos eius et manus suas super manus eius et incurvavit se super eum, et calefacta est caro pueri.
2KGS|4|35|At ille reversus deambulavit in domo semel huc et illuc et ascendit et incubuit super eum, et sternutavit puer septies aperuitque oculos.
2KGS|4|36|Et ille vocavit Giezi et dixit ei: " Voca Sunamitin hanc ". Quae vocata ingressa est ad eum. Qui ait: " Tolle filium tuum ".
2KGS|4|37|Venit illa et corruit ad pedes eius et adoravit super terram; tulitque filium suum et egressa est.
2KGS|4|38|Et Eliseus reversus est in Galgala. Erat autem fames in terra, et filii prophetarum habitabant coram eo. Dixitque puero suo: " Pone ollam grandem et coque pulmentum filiis prophetarum ".
2KGS|4|39|Et egressus est unus in agrum, ut colligeret herbas agrestes; invenitque quasi vitem silvestrem et collegit ex ea colocynthidas agri. Et implevit pallium suum et reversus concidit in ollam pulmenti; nesciebat enim quid esset.
2KGS|4|40|Infuderunt ergo sociis, ut comederent. Cumque gustassent de coctione, exclamaverunt dicentes: " Mors in olla, vir Dei! ". Et non potuerunt comedere.
2KGS|4|41|At ille: " Afferte, inquit, farinam ". Cumque tulissent, misit in ollam et ait: " Infunde turbae, et comedat ". Et non fuit amplius quidquam amaritudinis in olla.
2KGS|4|42|Vir autem quidam venit de Baalsalisa deferens viro Dei panes primitiarum, viginti panes hordeaceos et frumentum novum in pera sua. At ille dixit: " Da populo, ut comedat ".
2KGS|4|43|Responditque ei minister eius: " Quantum est hoc, ut apponam coram centum viris? ". Rursum ille dixit: " Da populo, ut comedat. Haec enim dicit Dominus: "Comedent, et supererit" ".
2KGS|4|44|Posuit itaque coram eis, qui comederunt, et superfuit iuxta verbum Domini.
2KGS|5|1|Naaman princeps militiae regis Syriae erat vir magnus apud dominum suum et honoratus; per illum enim dedit Dominus salutem Syriae. Erat autem vir fortis leprosus.
2KGS|5|2|Porro de Syria egressa fuerat turma et captivam duxerat de terra Israel puellam parvulam, quae erat in obsequio uxoris Naaman.
2KGS|5|3|Quae ait ad dominam suam: " Utinam esset dominus meus ad prophetam, qui est in Samaria! Profecto curaret eum a lepra, quam habet ".
2KGS|5|4|Ingressus est itaque Naaman ad dominum suum et nuntiavit ei dicens: " Sic et sic locuta est puella de terra Israel ".
2KGS|5|5|Dixitque ei rex Syriae: " Vade, et mittam litteras ad regem Israel ". Qui cum profectus esset et tulisset secum decem talenta argenti et sex milia siclorum auri et decem mutatoria vestimentorum,
2KGS|5|6|detulit litteras ad regem Israel in haec verba: " Cum acceperis epistulam hanc, scito quod miserim ad te Naaman servum meum, ut cures eum a lepra sua ".
2KGS|5|7|Cumque legisset rex Israel litteras, scidit vestimenta sua et ait: " Numquid Deus sum, ut occidere possim et vivificare, quia iste mittit ad me, ut curem hominem a lepra sua? Animadvertite et videte quod occasiones quaerat adversum me ".
2KGS|5|8|Quod cum audisset Eliseus vir Dei, scidisse videlicet regem Israel vestimenta sua, misit ad eum dicens: " Quare scidisti vestimenta tua? Veniat ad me et sciat esse prophetam in Israel ".
2KGS|5|9|Venit ergo Naaman cum equis et curribus et stetit ad ostium domus Elisei.
2KGS|5|10|Misitque ad eum Eliseus nuntium dicens: " Vade et lavare septies in Iordane; et recipiet sanitatem caro tua, atque mundaberis ".
2KGS|5|11|Iratus Naaman recedebat dicens: " Putabam quod egrederetur ad me et stans invocaret nomen Domini Dei sui et tangeret manu sua locum leprae et curaret me.
2KGS|5|12|Numquid non meliores sunt Abana et Pharphar, fluvii Damasci, omnibus aquis Israel, ut laver in eis et munder? ". Cum ergo vertisset se et abiret indignans,
2KGS|5|13|accesserunt ad eum servi sui et locuti sunt ei: " Si rem grandem dixisset tibi propheta, certe faceres; quanto magis quia nunc dixit tibi: Lavare et mundaberis!" ".
2KGS|5|14|Descendit et intinxit se in Iordane septies iuxta sermonem viri Dei, et restituta est caro eius sicut caro pueri parvuli, et mundatus est.
2KGS|5|15|Reversusque ad virum Dei cum universo comitatu suo venit et stetit coram eo et ait: " Vere scio quod non sit Deus in universa terra, nisi tantum in Israel! Obsecro itaque, ut accipias benedictionem a servo tuo ".
2KGS|5|16|At ille respondit: " Vivit Dominus, ante quem sto, non accipiam ". Cumque vim faceret, penitus non acquievit.
2KGS|5|17|Dixitque Naaman: " Ut vis. Sed, obsecro, concedatur mihi servo tuo tantum terrae quantum onus duorum burdonum; non enim faciet ultra servus tuus holocaustum aut victimam diis alienis, nisi Domino.
2KGS|5|18|Hoc autem solum ignoscat Dominus servo tuo, quando ingreditur dominus meus templum Remmon, ut adoret ibi, et illo innitente super manum meam, si adoravero in templo Remmon, adorante eo in eodem loco, ut ignoscat mihi Dominus servo tuo pro hac re ".
2KGS|5|19|Qui dixit ei: " Vade in pace ". Abiit ergo ab eo viam modicam.
2KGS|5|20|Dixitque Giezi puer viri Dei: " Pepercit dominus meus Naaman Syro isti, ut non acciperet ab eo, quae attulit; vivit Dominus, curram post eum et accipiam ab eo aliquid ".
2KGS|5|21|Et secutus est Giezi post tergum Naaman. Quem cum vidisset ille currentem ad se, desiluit de curru in occursum eius et ait: " Rectene sunt omnia? ".
2KGS|5|22|Et ille ait: " Recte. Dominus meus misit me dicens: "Modo venerunt ad me duo adulescentes de monte Ephraim ex filiis prophetarum. Da eis talentum argenti et vestes mutatorias duplices" ".
2KGS|5|23|Dixitque Naaman: " Melius est, ut accipias duo talenta ". Et coegit eum ligavitque duo talenta argenti in duobus saccis et duplicia vestimenta et imposuit duobus pueris suis, qui et portaverunt coram eo.
2KGS|5|24|Cumque venisset ad collem, tulit de manu eorum et reposuit in domo; dimisitque viros et abierunt.
2KGS|5|25|Ipse autem ingressus stetit coram domino suo. Et dixit Eliseus: " Unde venis, Giezi? ". Qui respondit: " Non ivit servus tuus quoquam ".
2KGS|5|26|At ille: " Nonne, ait, cor meum in praesenti erat, quando reversus est homo de curru suo in occursum tui? Estne tempus accipere argentum et accipere vestes et oliveta et vineta et oves et boves et servos et ancillas?
2KGS|5|27|Sed et lepra Naaman adhaerebit tibi et semini tuo in sempiternum ". Et egressus est ab eo leprosus quasi nix.
2KGS|6|1|Dixerunt autem filii prophetarum ad Eliseum: " Ecce locus, in quo habitamus coram te, angustus est nobis.
2KGS|6|2|Eamus usque ad Iordanem, et tollant singuli de silva materias singulas, ut aedificemus nobis ibi locum ad habitandum ". Qui dixit: " Ite ".
2KGS|6|3|Et ait unus ex illis: " Veni ergo et tu cum servis tuis ". Respondit: " Ego veniam ".
2KGS|6|4|Et abiit cum eis. Cumque venissent ad Iordanem, caedebant ligna.
2KGS|6|5|Accidit autem, ut, cum unus materiam succidisset, caderet ferrum securis in aquam; exclamavitque ille et ait: " Heu, domine mi! Et hoc ipsum mutuo acceperam! ".
2KGS|6|6|Dixit autem homo Dei: " Ubi cecidit? ". At ille monstravit ei locum. Praecidit ergo lignum et misit illuc, natavitque ferrum.
2KGS|6|7|Et ait: " Tolle!". Qui extendit manum et tulit illud.
2KGS|6|8|Rex autem Syriae pugnabat contra Israel; consiliumque iniit cum servis suis dicens: " In loco illo et illo ponamus insidias ".
2KGS|6|9|Misit itaque vir Dei ad regem Israel dicens: " Cave, ne transeas in loco illo, quia ibi Syri in insidiis sunt ".
2KGS|6|10|Misit rex Israel ad locum, quem dixerat ei vir Dei et de quo praemonuerat eum, et observavit se ibi non semel neque bis.
2KGS|6|11|Conturbatumque est cor regis Syriae pro hac re et, convocatis servis suis, ait: " Quare non indicatis mihi quis proditor mei sit apud regem Israel? ".
2KGS|6|12|Dixitque unus servorum eius: " Nequaquam, domine mi rex. Sed Eliseus propheta, qui est in Israel, indicat regi Israel omnia verba, quaecumque locutus fueris in conclavi tuo ".
2KGS|6|13|Dixit eis: " Ite et videte ubi sit, ut mittam et capiam eum ". Annuntiaveruntque ei dicentes: " Ecce in Dothain ".
2KGS|6|14|Misit ergo illuc equos et currus et robur exercitus; qui cum venissent nocte, circumdederunt civitatem.
2KGS|6|15|Consurgens autem diluculo minister viri Dei egressus est viditque exercitum in circuitu civitatis et equos et currus nuntiavitque ei dicens: Heu, domine mi, quid faciemus? ".
2KGS|6|16|At ille respondit: "Noli timere; plures enim nobiscum sunt quam cum illis".
2KGS|6|17|Oravitque Eliseus dicens: " Domine, aperi oculos huius, ut videat ". Et aperuit Dominus oculos pueri, et vidit, et ecce mons plenus equorum et curruum igneorum in circuitu Elisei.
2KGS|6|18|Hostes vero descenderunt ad eum. Porro Eliseus oravit Dominum dicens: " Percute, obsecro, gentem hanc caecitate! ". Percussitque eos Dominus, ne viderent iuxta verbum Elisei.
2KGS|6|19|Dixit autem ad eos Eliseus: " Non est haec via, nec ista est civitas; sequimini me, et ostendam vobis virum, quem quaeritis ". Duxit ergo eos in Samariam.
2KGS|6|20|Cumque ingressi fuissent in Samaria, dixit Eliseus: " Domine, aperi oculos istorum, ut videant ". Aperuitque Dominus oculos eorum, et viderunt esse se in medio Samariae.
2KGS|6|21|Dixitque rex Israel ad Eliseum, cum vidisset eos: " Numquid percutiam eos, pater mi? ".
2KGS|6|22|At ille ait: " Non percuties; neque enim, quos cepisti gladio et arcu tuo, percutis. Pone panem et aquam coram eis, ut comedant et bibant et vadant ad dominum suum ".
2KGS|6|23|Appositaque est eis ciborum magna praeparatio, et comederunt et biberunt, et dimisit eos; abieruntque ad dominum suum, et ultra non venerunt turmae Syriae in terram Israel.
2KGS|6|24|Factum est autem post haec, congregavit Benadad rex Syriae universum exercitum suum et ascendit et obsidebat Samariam.
2KGS|6|25|Factaque est fames magna in Samaria et tamdiu obsessa est, donec venumdaretur caput asini octoginta argenteis et quarta pars cabi stercoris columbarum quinque argenteis.
2KGS|6|26|Cumque rex Israel transiret per murum, mulier exclamavit ad eum dicens: Salva me, domine mi rex! ".
2KGS|6|27|Qui ait: " Non, salvet te te Dominus. Unde salvare te possum? De area an de torculari? ". Dixitque ad eam rex: " Quid tibi vis? ". Quae respondit:
2KGS|6|28|" Mulier ista dixit mihi: "Da filium tuum, ut comedamus eum hodie, et filium meum comedemus cras".
2KGS|6|29|Coximus ergo filium meum et comedimus. Dixique ei die altera: Da filium tuum, ut comedamus eum; quae abscondit filium suum ".
2KGS|6|30|Quod cum audisset rex, scidit vestimenta sua. Et transibat super murum, viditque omnis populus cilicium, quo vestitus erat ad carnem intrinsecus.
2KGS|6|31|Et ait: " Haec mihi faciat Deus et haec addat, si steterit caput Elisei filii Saphat super eum hodie ".
2KGS|6|32|Eliseus autem sedebat in domo sua, et senes sedebant cum eo. Praemisit itaque rex virum. Sed antequam veniret nuntius, Eliseus dixit ad senes: " Numquid scitis quod miserit filius homicidae hic, ut praecidatur caput meum? Videte ergo, cum venerit nuntius, claudite ostium et non sinatis eum introire; ecce enim sonitus pedum domini eius post eum est ".
2KGS|6|33|Et adhuc illo loquente eis, apparuit rex, qui veniebat ad eum, et ait: Ecce, tantum malum a Domino est; quid amplius exspectabo a Domino? ".
2KGS|7|1|Dixit autem Eliseus: " Audite verbum Domini. Haec dicit Dominus: In tempore hoc cras modius similae uno statere erit, et duo modii hordei statere uno in porta Samariae ".
2KGS|7|2|Respondens dux, super cuius manum rex incumbebat, homini Dei ait: " Si Dominus fecerit etiam cataractas in caelo, numquid poterit esse, quod loqueris? ". Qui ait: " Videbis oculis tuis et inde non comedes ".
2KGS|7|3|Quattuor ergo viri erant leprosi iuxta introitum portae; qui dixerunt ad invicem: " Quid hic esse volumus, donec moriamur?
2KGS|7|4|Sive ingredi voluerimus civitatem, fame moriemur; sive manserimus hic, moriendum nobis est. Venite igitur, et transfugiamus ad castra Syriae. Si pepercerint nobis, vivemus; si autem occidere voluerint, nihilominus moriemur ".
2KGS|7|5|Surrexerunt igitur vesperi, ut venirent ad castra Syriae. Cumque venissent ad principium castrorum Syriae, nullum ibidem reppererunt.
2KGS|7|6|Siquidem Dominus sonitum audiri fecerat in castris Syriae curruum et equorum et exercitus plurimi; dixeruntque ad invicem: " Ecce mercede conduxit adversum nos rex Israel reges Hetthaeorum et Aegyptiorum, ut venirent contra nos ".
2KGS|7|7|Surrexerunt ergo et fugerunt in tenebris et dereliquerunt tentoria sua et equos et asinos, castra, sicut erant; fugeruntque animas tantum suas salvare cupientes.
2KGS|7|8|Igitur cum venissent leprosi illi ad principium castrorum, ingressi sunt unum tabernaculum et comederunt et biberunt; tuleruntque inde argentum et aurum et vestes et abierunt et absconderunt. Et rursum reversi sunt ad aliud tabernaculum, et inde similiter auferentes absconderunt.
2KGS|7|9|Dixeruntque ad invicem: " Non recte facimus; haec enim dies boni nuntii est, et nos tacemus. Si noluerimus nuntiare usque mane, sceleris arguemur; venite, eamus et nuntiemus in aula regis ".
2KGS|7|10|Cumque venissent, vocaverunt portarios civitatis et narraverunt eis dicentes: " Ivimus ad castra Syriae et nullum ibidem repperimus hominum nisi equos et asinos alligatos et tentoria, sicut erant ".
2KGS|7|11|Clamaverunt ergo portarii et nuntiaverunt in palatio regis intrinsecus.
2KGS|7|12|Qui surrexit nocte et ait ad servos suos: " Dico vobis quid fecerint nobis Syri. Sciunt quia fame laboramus, et idcirco egressi sunt de castris et latitant in agris dicentes: "Cum egressi fuerint de civitate, capiemus eos viventes, et tunc civitatem ingredi poterimus" ".
2KGS|7|13|Respondit autem unus servorum eius: " Tollamus quinque equos, qui remanserunt in urbe; fiant sicut universa multitudo Israel, quae consumpta est; mittamus ergo et videamus ".
2KGS|7|14|Adduxerunt ergo duos currus cum equis, misitque rex post exercitum Syrorum dicens: " Ite et videte ".
2KGS|7|15|Qui abierunt post eos usque ad Iordanem; ecce autem omnis via plena erat vestibus et vasis, quae proiecerant Syri, cum turbarentur. Reversique nuntii indicaverunt regi.
2KGS|7|16|Et egressus populus diripuit castra Syriae; factusque est modius similae statere uno, et duo modii hordei statere uno iuxta verbum Domini.
2KGS|7|17|Porro rex ducem illum, in cuius manu incumbebat, constituit ad portam; quem conculcavit turba in introitu, et mortuus est iuxta quod locutus fuerat vir Dei, quando descenderat rex ad eum.
2KGS|7|18|Factumque est secundum sermonem viri Dei, quem dixerat regi, quando ait: " Duo modii hordei statere uno erunt, et modius similae statere uno hoc eodem tempore cras in porta Samariae ";
2KGS|7|19|quando responderat dux ille viro Dei et dixerat: " Etiamsi Dominus fecerit cataractas in caelo, numquid fieri poterit, quod loqueris? ", et dixerat ei: " Videbis oculis tuis et inde non comedes ".
2KGS|7|20|Evenit ergo ei, sicut praedictum erat, et conculcavit eum populus in porta, et mortuus est.
2KGS|8|1|Eliseus autem locutus est ad mulierem, cuius vivere fecerat fi lium, dicens: " Surge, vade tu et domus tua et peregrinare ubicumque reppereris; vocavit enim Dominus famem, et veniet super terram septem annis ".
2KGS|8|2|Quae surrexit et fecit iuxta verbum hominis Dei et vadens cum domo sua peregrinata est in terra Philisthim septem annis.
2KGS|8|3|Cumque finiti essent anni septem, reversa est mulier de terra Philisthim; et egressa est, ut interpellaret regem pro domo sua et agris suis.
2KGS|8|4|Rex autem loquebatur cum Giezi puero viri Dei dicens: " Narra mihi omnia magnalia, quae fecit Eliseus ".
2KGS|8|5|Cumque ille narraret regi quomodo mortuum suscitasset, apparuit mulier, cuius vivificaverat filium, clamans ad regem pro domo sua et pro agris suis. Dixitque Giezi: " Domine mi rex, haec est mulier, et hic filius eius, quem suscitavit Eliseus ".
2KGS|8|6|Et interrogavit rex mulierem, quae narravit ei. Deditque ei rex eunuchum unum dicens: " Restitue ei omnia, quae sua sunt, et universos reditus agrorum a die, qua reliquit terram usque ad praesens ".
2KGS|8|7|Venit quoque Eliseus Damascum, et Benadad rex Syriae aegrotabat. Nuntiaveruntque ei dicentes: " Venit vir Dei huc ".
2KGS|8|8|Et ait rex ad Hazael: " Tolle tecum munera et vade in occursum viri Dei et consule Dominum per eum dicens: Si evadere potero de infirmitate mea hac? ".
2KGS|8|9|Ivit igitur Hazael in occursum eius habens secum munera et omnia bona Damasci, onera quadraginta camelorum. Cumque stetisset coram eo, ait: " Filius tuus Benadad rex Syriae misit me ad te dicens: "Si sanari potero de infirmitate mea hac?" ".
2KGS|8|10|Dixitque ei Eliseus: " Vade, dic ei: Sanaberis. Porro ostendit mihi Dominus quia morte morietur ".
2KGS|8|11|Stetitque facies eius, et conturbatus est usque ad suffusionem vultus flevitque vir Dei.
2KGS|8|12|Cui Hazael ait: " Quare dominus meus flet? ". At ille respondit: " Quia scio, quae facturus sis filiis Israel mala: civitates eorum munitas igne succendes et iuvenes eorum interficies gladio et parvulos eorum elides et praegnantes discindes ".
2KGS|8|13|Dixitque Hazael: " Quid enim sum servus tuus canis, ut faciam rem istam magnam? ". Et ait Eliseus: " Ostendit mihi Dominus te regem Syriae fore ".
2KGS|8|14|Qui cum recessisset ab Eliseo, venit ad dominum suum. Qui ait ei: " Quid tibi dixit Eliseus? ". At ille respondit: " Dixit mihi: Recipies sanitatem ".
2KGS|8|15|Cumque venisset dies altera, tulit stragulum et intinxit aqua et expandit super faciem eius, et mortuus est; regnavitque Hazael pro eo.
2KGS|8|16|Anno quinto Ioram filii Achab regis Israel - Iosaphat autem erat rex Iudae - regnavit Ioram filius Iosaphat regis Iudae.
2KGS|8|17|Triginta duorum erat annorum, cum regnare coepisset, et octo annis regnavit in Ierusalem.
2KGS|8|18|Ambulavitque in viis regum Israel, sicut ambulaverat domus Achab; filia enim Achab erat uxor eius. Et fecit, quod malum est coram Domino.
2KGS|8|19|Noluit autem Dominus disperdere Iudam propter David servum suum, sicut promiserat ei, ut daret illi lucernam et filiis eius cunctis diebus.
2KGS|8|20|In diebus eius recessit Edom, ne esset sub Iuda, et constituit sibi regem.
2KGS|8|21|Venitque Ioram Seira et omnis currus cum eo; et surrexit nocte percussitque Idumaeos, qui eum circumdederant, et principes curruum; et populus fugit in tabernacula sua.
2KGS|8|22|Recessit ergo Edom, ne esset sub Iuda, usque ad diem hanc. Tunc recessit et Lobna in tempore illo.
2KGS|8|23|Reliqua autem gestorum Ioram et universa, quae fecit, nonne haec scripta sunt in libro annalium regum Iudae?
2KGS|8|24|Et dormivit Ioram cum patribus suis sepultusque est cum eis in civitate David; et regnavit Ochozias filius eius pro eo.
2KGS|8|25|Anno duodecimo Ioram filii Achab regis Israel regnavit Ochozias filius Ioram regis Iudae.
2KGS|8|26|Viginti duorum annorum erat Ochozias, cum regnare coepisset, et uno anno regnavit in Ierusalem. Nomen matris eius Athalia filia Amri regis Israel.
2KGS|8|27|Et ambulavit in viis domus Achab et fecit, quod malum est coram Domino, sicut domus Achab; gener enim domus Achab fuit.
2KGS|8|28|Abiit quoque cum Ioram filio Achab ad proeliandum contra Hazael regem Syriae in Ramoth Galaad; et vulneraverunt Syri Ioram.
2KGS|8|29|Qui reversus est, ut curaretur in Iezrahel de vulneribus, quibus vulneraverant eum Syri in Rama proeliantem contra Hazael regem Syriae. Porro Ochozias filius Ioram rex Iudae descendit invisere Ioram filium Achab in Iezrahel, quia aegrotabat.
2KGS|9|1|Eliseus autem prophetes vocavit unum de filiis prophetarum et ait illi: Accinge lumbos tuos et tolle lenticulam olei hanc in manu tua et vade in Ramoth Galaad.
2KGS|9|2|Cumque veneris illuc, videbis Iehu filium Iosaphat filii Namsi et ingressus suscitabis eum de medio fratrum suorum et introduces interius cubiculum.
2KGS|9|3|Tenensque lenticulam olei fundes super caput eius et dices: " Haec dicit Dominus: Unxi te regem super Israel ". Aperiesque ostium et fugies et non ibi subsistes ".
2KGS|9|4|Abiit ergo adulescens puer prophetae Ramoth Galaad
2KGS|9|5|et ingressus est. Ecce autem principes exercitus sedebant, et ait: " Verbum mihi ad te, princeps ". Dixitque Iehu: " Ad quem ex omnibus nobis?. At ille dixit: " Ad te, o princeps ".
2KGS|9|6|Et surrexit et ingressus est cubiculum. At ille fudit oleum super caput eius et ait: " Haec dicit Dominus, Deus Israel: Unxi te regem super populum Domini, super Israel.
2KGS|9|7|Percuties domum Achab domini tui, ut ulciscar sanguinem servorum meorum prophetarum et sanguinem omnium servorum Domini de manu Iezabel.
2KGS|9|8|Perdamque omnem domum Achab et interficiam de Achab quidquid masculini sexus et impuberem et puberem in Israel.
2KGS|9|9|Et dabo domum Achab sicut domum Ieroboam filii Nabat et sicut domum Baasa filii Ahiae.
2KGS|9|10|Iezabel quoque comedent canes in agro Iezrahel, nec erit qui sepeliat eam ". Aperuitque ostium et fugit.
2KGS|9|11|Iehu autem egressus est ad servos domini sui, qui dixerunt ei: " Rectene sunt omnia? Quid venit insanus iste ad te? ". Qui ait eis: " Nostis hominem et loquelam eius ".
2KGS|9|12|At illi responderunt: " Mendacium! Narra nobis! ". Qui ait eis: " Haec et haec locutus est mihi dicens: "Haec dicit Dominus: Unxi te regem super Israel" ".
2KGS|9|13|Festinaverunt itaque et unusquisque tollens pallium suum posuerunt sub pedibus eius super structuram graduum et cecinerunt tuba atque dixerunt: " Regnavit Iehu! ".
2KGS|9|14|Coniuravit ergo Iehu filius Iosaphat filii Namsi contra Ioram. Porro Ioram defenderat Ramoth Galaad ipse et omnis Israel contra Hazael regem Syriae
2KGS|9|15|et reversus fuerat, ut curaretur in Iezrahel propter vulnera, quia percusserant eum Syri proeliantem contra Hazael regem Syriae. Dixitque Iehu: " Si placet vobis, nemo egrediatur profugus de civitate, ne vadat et nuntiet in Iezrahel ".
2KGS|9|16|Et ascendit et profectus est in Iezrahel; Ioram enim aegrotabat ibi, et Ochozias rex Iudae descenderat ad visitandum Ioram.
2KGS|9|17|Igitur speculator, qui stabat super turrim Iezrahel, vidit globum Iehu venientis et ait: " Video ego globum ". Dixitque Ioram: " Tolle equitem et mitte in occursum eorum, et dicat vadens: "Rectene sunt omnia?" ".
2KGS|9|18|Abiit igitur, qui ascenderat equum in occursum eius, et ait: " Haec dicit rex: Pacatane sunt omnia? ". Dixitque ei Iehu: " Quid tibi et paci? Transi et sequere me ". Nuntiavit quoque speculator dicens: " Venit nuntius ad eos et non revertitur ".
2KGS|9|19|Misit etiam equitem secundum; venitque ad eos et ait: " Haec dicit rex: Num pax est? ". Et ait Iehu: " Quid tibi et paci? Transi et sequere me ".
2KGS|9|20|Nuntiavit autem speculator dicens: " Venit usque ad eos et non revertitur. Est autem incessus quasi incessus Iehu filii Namsi; praeceps enim graditur ".
2KGS|9|21|Et ait Ioram: " Iunge currum! ". Iunxeruntque currum eius, et egressus est Ioram rex Israel et Ochozias rex Iudae singuli in curribus suis. Egressique sunt in occursum Iehu et invenerunt eum in agro Naboth Iezrahelitis.
2KGS|9|22|Cumque vidisset Ioram Iehu, dixit: " Estne pax, Iehu? ". At ille respondit: " Quae pax? Adhuc fornicationes Iezabel matris tuae et veneficia eius multa vigent! ".
2KGS|9|23|Convertit autem Ioram manum suam et fugiens ait ad Ochoziam: " Insidiae, Ochozia! ".
2KGS|9|24|Porro Iehu tetendit arcum manu et percussit Ioram inter scapulas. Et egressa est sagitta per cor eius; statimque corruit in curru suo.
2KGS|9|25|Dixitque Iehu ad Badacer ducem: " Tolle, proice eum in agro Naboth Iezrahelitae! Memento enim: ego et tu eramus cum his, qui vectabantur gemini post Achab patrem huius, quando Dominus onus hoc levavit super eum dicens:
2KGS|9|26|"Pro sanguine Naboth et pro sanguine filiorum eius, quem vidi heri, ait Dominus, reddam tibi in agro isto, dicit Dominus". Nunc igitur tolle, proice eum in agro iuxta verbum Domini ".
2KGS|9|27|Ochozias autem rex Iudae videns hoc fugit per viam Bethgan; persecutusque est eum Iehu et ait: " Etiam hunc percutite! ". Et percusserunt eum in curru suo in ascensu Gaver, qui est iuxta Ieblaam. Qui fugit in Mageddo et mortuus est ibi.
2KGS|9|28|Et imposuerunt eum servi eius super currum suum et tulerunt Ierusalem sepelieruntque in sepulcro cum patribus suis in civitate David.
2KGS|9|29|Anno undecimo Ioram filii Achab regnavit Ochozias super Iudam.
2KGS|9|30|Venit Iehu Iezrahel. Porro Iezabel, introitu eius audito, depinxit oculos suos stibio et ornavit caput suum et respexit per fenestram
2KGS|9|31|ingredientem Iehu per portam et ait: " Numquid pax esse potest Zamri, qui interfecit dominum suum? ".
2KGS|9|32|Levavitque Iehu faciem suam ad fenestram et ait: " Quis est mecum, quisnam? ". Et inclinaverunt se ad eum duo vel tres eunuchi.
2KGS|9|33|At ille dixit eis: " Praecipitate eam deorsum! ". Et praecipitaverunt eam; aspersusque est sanguine paries et equi, qui conculcaverunt eam.
2KGS|9|34|Cumque ingressus esset, ut comederet biberetque, ait: " Ite, videte maledictam illam et sepelite eam, quia filia regis est ".
2KGS|9|35|Cumque issent, ut sepelirent eam, non invenerunt nisi calvariam et pedes et summas manus.
2KGS|9|36|Reversique nuntiaverunt ei. Et ait Iehu: " Sermo Domini est, quem locutus est per servum suum Eliam Thesbiten dicens: In agro Iezrahel comedent canes carnes Iezabel;
2KGS|9|37|et erit cadaver Iezabel sicut stercus super faciem terrae in agro Iezrahel, ita ut non dicatur: "Haeccine est illa Iezabel" ".
2KGS|10|1|Erant autem Achab septuaginta filii in Samaria. Scripsit ergo Iehu litteras et misit in Samariam ad optimates civitatis et ad maiores natu et ad nutricios filiorum Achab dicens:
2KGS|10|2|" Statim ut acceperitis litteras has, qui habetis filios domini vestri et currus et equos et civitatem firmam et arma,
2KGS|10|3|eligite meliorem et iustiorem de filiis domini vestri et ponite eum super solium patris sui et pugnate pro domo domini vestri ".
2KGS|10|4|Timuerunt illi vehementer et dixerunt: " Ecce duo reges non potuerunt stare coram eo, et quomodo nos valebimus resistere? ".
2KGS|10|5|Miserunt ergo praepositus domus et praefectus civitatis et maiores natu et nutricii ad Iehu dicentes: " Servi tui sumus: quaecumque iusseris, faciemus nec constituemus regem; quodcumque tibi placet, fac ".
2KGS|10|6|Rescripsit autem eis litteras secundo dicens: " Si mei estis et oboeditis mihi, tollite capita virorum filiorum domini vestri et venite ad me hac eadem hora cras in Iezrahel ". Porro filii regis, septuaginta viri, apud optimates civitatis nutriebantur.
2KGS|10|7|Cumque venissent litterae ad eos, tulerunt filios regis et occiderunt septuaginta viros et posuerunt capita eorum in cophinis et miserunt ad eum in Iezrahel.
2KGS|10|8|Venit autem nuntius et indicavit ei dicens: " Attulerunt capita filiorum regis". Qui respondit: " Ponite ea duos acervos iuxta introitum portae usque mane ".
2KGS|10|9|Cumque diluxisset, egressus est et stans dixit ad omnem populum: " Vos iusti estis; ecce ego coniuravi contra dominum meum et interfeci eum, sed quis percussit omnes hos?
2KGS|10|10|Videte ergo nunc quoniam non cecidit de sermonibus Domini in terram, quos locutus est Dominus super domum Achab, et Dominus fecit, quod locutus est in manu servi sui Eliae ".
2KGS|10|11|Percussit igitur Iehu omnes, qui reliqui erant de domo Achab in Iezrahel, et universos optimates eius et notos et sacerdotes, donec non remanerent ex eo reliquiae.
2KGS|10|12|Et surrexit et intravit. Deinde profectus est in Samariam; cumque esset ad Betheced Pastorum in via,
2KGS|10|13|invenit fratres Ochoziae regis Iudae dixitque ad eos: " Quinam estis vos? ". At illi responderunt: " Fratres Ochoziae sumus et descendimus ad salutandos filios regis et filios dominae reginae ".
2KGS|10|14|Qui ait: " Comprehendite eos vivos ". Quos cum comprehendissent vivos, iugulaverunt eos iuxta cisternam Betheced, quadraginta duos viros, et non reliquit ex eis quemquam.
2KGS|10|15|Cumque abisset inde, invenit Ionadab filium Rechab in occursum sibi et benedixit ei. Et ait ad eum: " Numquid est cor tuum rectum sicut cor meum cum corde tuo? ". Et ait Ionadab: " Est ". " Si est, inquit, da manum tuam. Qui dedit manum suam. At ille levavit eum ad se in curru
2KGS|10|16|dixitque ad eum: " Veni mecum et vide zelum meum pro Domino ". Et impositum currui suo
2KGS|10|17|duxit in Samariam. Et percussit omnes, qui reliqui fuerant de Achab in Samaria usque ad unum, iuxta verbum Domini, quod locutus est per Eliam.
2KGS|10|18|Congregavit ergo Iehu omnem populum et dixit ad eos: " Achab coluit Baal parum, ego autem colam eum amplius.
2KGS|10|19|Nunc igitur omnes prophetas Baal et universos servos eius et cunctos sacerdotes ipsius vocate ad me; nullus sit qui non veniat. Sacrificium enim grande est mihi Baal; quicumque defuerit, non vivet ". Porro Iehu faciebat hoc insidiose, ut disperderet cultores Baal.
2KGS|10|20|Dixitque: " Sanctificate diem sollemnem Baal ". Vocaveruntque.
2KGS|10|21|Et misit Iehu in universos terminos Israel, et venerunt cuncti servi Baal; non fuit residuus, ne unus quidem qui non veniret. Et ingressi sunt templum Baal, et repleta est domus Baal a summo usque ad summum.
2KGS|10|22|Dixitque ei, qui erat super vestes: " Profer vestimenta universis servis Baal ". Et protulit eis vestes.
2KGS|10|23|Ingressusque Iehu et Ionadab filius Rechab templum Baal ait cultoribus Baal: " Perquirite et videte, ne quis forte vobiscum sit de servis Domini, sed ut sint soli servi Baal ".
2KGS|10|24|Ingressi sunt igitur, ut facerent victimas et holocausta; Iehu autem praeparaverat sibi foris octoginta viros et dixerat eis: " Quicumque permiserit fugere de hominibus his, quos ego adduxero in manus vestras, anima eius erit pro anima illius ".
2KGS|10|25|Factum est ergo cum completum esset holocaustum, praecepit Iehu cursoribus et ducibus suis: " Ingredimini et percutite eos; nullus evadat!. Percusseruntque eos cursores et duces ore gladii et proiecerunt. Tunc ierunt usque in dabir templi Baal.
2KGS|10|26|Et protulerunt lapidem Baal et combusserunt
2KGS|10|27|et comminuerunt eum. Destruxerunt quoque aedem Baal et fecerunt pro ea latrinas usque diem hanc.
2KGS|10|28|Delevit itaque Iehu Baal de Israel.
2KGS|10|29|Verumtamen a peccatis Ieroboam filii Nabat, qui peccare fecerat Israel, non recessit; nec dereliquit vitulos aureos, qui erant in Bethel et in Dan.
2KGS|10|30|Dixit autem Dominus ad Iehu: " Quia studiose fecisti, quod rectum erat in oculis meis et omnia quae erant in corde meo fecisti contra domum Achab, filii tui usque ad quartam generationem sedebunt super thronum Israel ".
2KGS|10|31|Porro Iehu non custodivit, ut ambularet in lege Domini, Dei Israel, in toto corde suo; non enim recessit a peccatis Ieroboam, qui peccare fecerat Israel.
2KGS|10|32|In diebus illis coepit Dominus discindere in Israel; percussitque eos Hazael in universis finibus Israel
2KGS|10|33|a Iordane contra orientalem plagam omnem terram Galaad et Gad et Ruben et Manasse, ab Aroer, quae est super torrentem Arnon, et Galaad et Basan.
2KGS|10|34|Reliqua autem gestorum Iehu et universa, quae fecit, et fortitudo eius, nonne haec scripta sunt in libro annalium regum Israel?
2KGS|10|35|Et dormivit Iehu cum patribus suis, sepelieruntque eum in Samaria; et regnavit Ioachaz filius eius pro eo.
2KGS|10|36|Dies autem, quos regnavit Iehu super Israel, viginti et octo anni sunt, in Samaria.
2KGS|11|1|Athalia vero mater Ochoziae videns mortuum filium suum surrexit et interfecit omne semen regium.
2KGS|11|2|Tollens autem Iosaba filia regis Ioram soror Ochoziae Ioas filium Ochoziae furata est eum de medio filiorum regis, qui interficiebantur, et nutricem eius in cubiculo lectulorum, et absconderunt eum a facie Athaliae, ut non interficeretur.
2KGS|11|3|Eratque cum ea in domo Domini clam sex annis; porro Athalia regnavit super terram.
2KGS|11|4|Anno autem septimo misit Ioiada et assumens centuriones Carum et cursorum introduxit ad se in templum Domini pepigitque cum eis foedus; et adiurans eos in domo Domini ostendit eis filium regis
2KGS|11|5|et praecepit illis dicens: " Hoc est, quod facere debetis: tertia pars vestrum introeat sabbato et observet excubitum domus regis;
2KGS|11|6|tertia autem pars ad portam Sur, et tertia pars sit ad portam, quae est post habitaculum cursorum, et custodietis excubitum domus per vices.
2KGS|11|7|Duae vero partes e vobis omnes egredientes sabbato custodiant excubias domus Domini circum regem.
2KGS|11|8|Et vallabitis eum habentes arma in manibus vestris; si quis autem ingressus fuerit saeptum templi, interficiatur; eritisque cum rege introeunte et egrediente.
2KGS|11|9|Et fecerunt centuriones iuxta omnia, quae praeceperat eis Ioiada sacerdos, et assumentes singuli viros suos, qui ingrediebantur sabbato, cum his, qui egrediebantur sabbato, venerunt ad Ioiada sacerdotem.
2KGS|11|10|Qui dedit centurionibus hastas et peltas regis David, quae erant in domo Domini.
2KGS|11|11|Et steterunt cursores singuli habentes arma in manu sua a parte templi dextera usque ad partem templi sinistram contra altare et aedem circum regem.
2KGS|11|12|Produxitque filium regis et dedit ei diadema et testimonium; feceruntque eum regem et unxerunt et plaudentes manu dixerunt: " Vivat rex! ".
2KGS|11|13|Audivit autem Athalia vocem populi et ingressa ad turbas in templum Domini
2KGS|11|14|vidit regem stantem super tribunal iuxta morem et principes et tubas prope eum omnemque populum terrae laetantem et canentem tubis; et scidit vestimenta sua clamavitque: " Coniuratio, coniuratio! ".
2KGS|11|15|Praecepit autem Ioiada sacerdos centurionibus, qui erant super exercitum, et ait eis: " Educite eam extra consaepta templi, et, quicumque secutus eam fuerit, feriatur gladio ". Dixerat enim sacerdos: " Non occidatur in templo Domini ".
2KGS|11|16|Imposueruntque ei manus et impegerunt eam per viam introitus Equorum in palatium, et interfecta est ibi.
2KGS|11|17|Pepigit igitur Ioiada foedus inter Dominum et inter regem et inter populum, ut esset populus Domini, et inter regem et populum.
2KGS|11|18|Ingressusque est omnis populus terrae templum Baal, et destruxerunt illud et aras eius et imagines contriverunt valide; Matthan quoque sacerdotem Baal occiderunt coram altaribus.Et posuit sacerdos custodias in domo Domini
2KGS|11|19|tulitque centuriones et Cares et cursores et omnem populum terrae; deduxeruntque regem de domo Domini. Et venerunt per viam portae Cursorum in palatium, et sedit super thronum regum.
2KGS|11|20|Laetatusque est omnis populus terrae, et civitas conquievit; Athalia autem occisa est gladio in domo regis.
2KGS|12|1|Septemque annorum erat Ioas, cum regnare coepisset.
2KGS|12|2|Anno septimo Iehu regnavit Ioas; quadraginta annis regnavit in Ierusalem. Nomen matris eius Sebia de Bersabee.
2KGS|12|3|Fecitque Ioas rectum coram Domino cunctis diebus, quibus docuit eum Ioiada sacerdos.
2KGS|12|4|Verumtamen excelsa non abstulit; adhuc populus immolabat et adolebat in excelsis.
2KGS|12|5|Dixitque Ioas ad sacerdotes: " Omnem pecuniam sanctorum, quae illata fuerit in templum Domini a praetereuntibus, quae offertur pro pretio animae, et quam sponte et arbitrio cordis sui inferunt in templum Domini,
2KGS|12|6|accipiant illam singuli sacerdotes a notis suis et instaurent sartatecta domus, si quid necessarium viderint instauratione ".
2KGS|12|7|Igitur usque ad vicesimum tertium annum regis Ioas non instauraverunt sacerdotes sartatecta templi.
2KGS|12|8|Vocavitque rex Ioas Ioiada pontificem et sacerdotes dicens eis: " Quare sartatecta non instauratis templi? Nolite ergo amplius accipere pecuniam a notis vestris, sed ad instaurationem templi reddite eam ".
2KGS|12|9|Acquieveruntque sacerdotes ultra non accipere pecuniam a populo nec instaurare sartatecta domus.
2KGS|12|10|Et tulit Ioiada pontifex gazophylacium unum aperuitque foramen desuper et posuit illud iuxta altare ad dexteram ingredientium domum Domini; mittebantque in eo sacerdotes, qui custodiebant ostia, omnem pecuniam, quae deferebatur ad templum Domini.
2KGS|12|11|Cumque viderent multam pecuniam esse in gazophylacio, ascendebat scriba regis et pontifex, colligebantque et numerabant pecuniam, quae inveniebatur in domo Domini,
2KGS|12|12|et dabant eam iuxta numerum atque mensuram in manu opificum, qui operibus praepositi erant in domo Domini; ipsique impendebant eam in fabris lignorum et in structoribus, qui operabantur in domo Domini,
2KGS|12|13|et in caementariis et in his, qui caedebant saxa, et ut emerent ligna et lapides de lapicidinis, ut instaurarentur sartatecta domus Domini, et pro universis, quae indigebant expensa ad muniendam domum.
2KGS|12|14|Verumtamen non fiebant pelves argenteae templi Domini et cultri et paterae et tubae, omne vas aureum et argenteum, de pecunia, quae inferebatur in templum Domini;
2KGS|12|15|opificibus enim dabatur, ut instauraretur templum Domini.
2KGS|12|16|Et non fiebat ratio his hominibus, qui accipiebant pecuniam, ut distribuerent eam operariis; illi enim in fide agebant.
2KGS|12|17|Pecuniam vero pro delicto et pecuniam pro peccatis non inferebatur in templum Domini, quia sacerdotum erat.
2KGS|12|18|Tunc ascendit Hazael rex Syriae et pugnabat contra Geth; cepitque eam et direxit faciem suam, ut ascenderet in Ierusalem.
2KGS|12|19|Quam ob rem tulit Ioas rex Iudae omnia sanctificata, quae consecraverant Iosaphat et Ioram et Ochozias patres eius reges Iudae, et quae ipse obtulerat, et universum aurum, quod inveniri potuit in thesauris templi Domini et in palatio regis, misitque Hazaeli regi Syriae; et recessit ab Ierusalem.
2KGS|12|20|Reliqua autem gestorum Ioas et universa, quae fecit, nonne haec scripta sunt in libro annalium regum Iudae?
2KGS|12|21|Surrexerunt autem servi eius et coniuraverunt inter se percusseruntque Ioas in domo Mello in descensu Sella.
2KGS|12|22|Iozachar namque filius Semath et Iozabad filius Somer servi eius percusserunt eum, et mortuus est; et sepelierunt eum cum patribus suis in civitate David. Regnavitque Amasias filius eius pro eo.
2KGS|13|1|Anno vicesimo tertio Ioas fi lii Ochoziae regis Iudae re gnavit Ioachaz filius Iehu super Israel in Samaria decem et septem annis.
2KGS|13|2|Et fecit malum coram Domino secutusque est peccatum Ieroboam filii Nabat, qui peccare fecit Israel; non declinavit ab eo.
2KGS|13|3|Iratusque est furor Domini contra Israel et tradidit eos in manu Hazael regis Syriae et in manu Benadad filii Hazael cunctis diebus.
2KGS|13|4|Deprecatus est autem Ioachaz faciem Domini, et audivit eum Dominus; vidit enim angustiam Israel, qua attriverat eos rex Syriae.
2KGS|13|5|Et dedit Dominus Israeli salvatorem, et liberatus est de manu Syriae; habitaveruntque filii Israel in tabernaculis suis sicut heri et nudiustertius.
2KGS|13|6|Verumtamen non recesserunt a peccatis domus Ieroboam, qui peccare fecit Israel; in ipsis ambulaverunt. Siquidem et palus permansit in Samaria.
2KGS|13|7|Et non reliquit Dominus Ioachaz de populo nisi quinquaginta equites et decem currus et decem milia peditum; interfecerat enim eos rex Syriae et redegerat quasi pulverem in tritura areae.
2KGS|13|8|Reliqua autem gestorum Ioachaz et universa, quae fecit, sed et fortitudo eius, nonne haec scripta sunt in libro annalium regum Israel?
2KGS|13|9|Dormivitque Ioachaz cum patribus suis, et sepelierunt eum in Samaria. Regnavitque Ioas filius eius pro eo.
2KGS|13|10|Anno tricesimo septimo Ioas regis Iudae regnavit Ioas filius Ioachaz super Israel in Samaria sedecim annis.
2KGS|13|11|Et fecit, quod malum est in conspectu Domini; non declinavit ab omnibus peccatis Ieroboam filii Nabat, qui peccare fecit Israel; in ipsis ambulavit.
2KGS|13|12|Reliqua autem gestorum Ioas et universa, quae fecit, sed et fortitudo eius, quomodo pugnaverit contra Amasiam regem Iudae, nonne haec scripta sunt in libro annalium regum Israel?
2KGS|13|13|Et dormivit Ioas cum patribus suis; Ieroboam autem sedit super solium eius. Porro Ioas sepultus est in Samaria cum regibus Israel.
2KGS|13|14|Eliseus autem aegrotabat infirmitate, qua et mortuus est; descenditque ad eum Ioas rex Israel et flebat coram eo dicebatque: " Pater mi, pater mi, currus Israel et auriga eius! ".
2KGS|13|15|Et ait illi Eliseus: "Affer arcum et sagittas". Cumque attulisset ad eum arcum et sagittas,
2KGS|13|16|dixit ad regem Israel: " Pone manum tuam super arcum ". Et, cum posuisset ille manum suam, superposuit Eliseus manus suas manibus regis
2KGS|13|17|et ait: " Aperi fenestram orientalem ". Cumque aperuisset, dixit Eliseus: "Iace sagittam!". Et iecit. Et ait Eliseus: " Sagitta salutis Domini, et sagitta salutis contra Syriam. Percutiesque Syriam in Aphec, donec consumas eam ".
2KGS|13|18|Et ait: " Tolle sagittas ". Qui cum tulisset, rursum dixit ei: " Percute iaculo terram!". Et, cum percussisset tribus vicibus et stetisset,
2KGS|13|19|iratus est contra eum vir Dei et ait: " Si percussisses quinquies aut sexies, percussisses Syriam usque ad consummationem; nunc autem tribus vicibus percuties eam ".
2KGS|13|20|Mortuus est ergo Eliseus, et sepelierunt eum. Latrunculi autem de Moab venerunt in terra in ipso anno.
2KGS|13|21|Quidam autem sepelientes hominem viderunt latrunculos et proiecerunt cadaver in sepulcro Elisei et abierunt. Quod cum tetigisset ossa Elisei, revixit homo et stetit super pedes suos.
2KGS|13|22|Igitur Hazael rex Syriae afflixit Israel cunctis diebus Ioachaz.
2KGS|13|23|Et misertus est Dominus eorum et reversus est ad eos propter pactum suum, quod habebat cum Abraham, Isaac et Iacob, et noluit disperdere eos neque proicere penitus usque in praesens tempus.
2KGS|13|24|Mortuus est autem Hazael rex Syriae; et regnavit Benadad filius eius pro eo.
2KGS|13|25|Porro Ioas filius Ioachaz tulit urbes de manu Benadad filii Hazael, quas tulerat de manu Ioachaz patris sui iure proelii; tribus vicibus percussit eum Ioas et reddidit civitates Israeli.
2KGS|14|1|Anno secundo Ioas filii Ioachaz regis Israel regnavit Amasias filius Ioas regis Iudae.
2KGS|14|2|Viginti quinque annorum erat, cum regnare coepisset, viginti autem et novem annis regnavit in Ierusalem. Nomen matris eius Ioaden de Ierusalem.
2KGS|14|3|Et fecit rectum coram Domino, verumtamen non ut David pater eius. Iuxta omnia, quae fecit Ioas pater suus, fecit,
2KGS|14|4|nisi hoc quod excelsa non abstulit; adhuc enim populus immolabat et adolebat in excelsis.
2KGS|14|5|Cumque obtinuisset regnum, percussit servos suos, qui interfecerant regem patrem suum;
2KGS|14|6|filios autem eorum, qui occiderant, non occidit, iuxta quod scriptum est in libro legis Moysi, sicut praecepit Dominus dicens: " Non morientur patres pro filiis, neque filii morientur pro patribus, sed unusquisque in peccato suo morietur ".
2KGS|14|7|Ipse percussit Edom in valle Salinarum decem milia et apprehendit Petram in proelio vocavitque nomen eius Iecethel usque in praesentem diem.
2KGS|14|8|Tunc misit Amasias nuntios ad Ioas filium Ioachaz filii Iehu regem Israel dicens: " Veni, et videamus nos ".
2KGS|14|9|Remisitque Ioas rex Israel ad Amasiam regem Iudae dicens: " Carduus Libani misit ad cedrum, quae est in Libano, dicens: "Da filiam tuam filio meo uxorem". Transieruntque bestiae agri, quae sunt in Libano, et conculcaverunt carduum.
2KGS|14|10|Percutiens invaluisti super Edom, et sublevavit te cor tuum; contentus esto gloria et sede in domo tua. Quare provocas malum, ut cadas tu et Iuda tecum? ".
2KGS|14|11|Et non acquievit Amasias.Ascenditque Ioas rex Israel, et viderunt se ipse et Amasias rex Iudae in Bethsames oppido Iudae.
2KGS|14|12|Percussusque est Iuda coram Israel, et fugerunt unusquisque in tabernacula sua.
2KGS|14|13|Amasiam vero regem Iudae filium Ioas filii Ochoziae cepit Ioas rex Israel in Bethsames et adduxit eum in Ierusalem. Et interrupit murum Ierusalem a porta Ephraim usque ad portam Anguli quadringentis cubitis.
2KGS|14|14|Tulitque omne aurum et argentum et universa vasa, quae inventa sunt in domo Domini et in thesauris regis, et obsides; et reversus est Samariam.
2KGS|14|15|Reliqua autem gestorum Ioas, quae fecit, et fortitudo eius, qua pugnavit contra Amasiam regem Iudae, nonne haec scripta sunt in libro annalium regum Israel?
2KGS|14|16|Dormivitque Ioas cum patribus suis et sepultus est in Samaria cum regibus Israel; et regnavit Ieroboam filius eius pro eo.
2KGS|14|17|Vixit autem Amasias filius Ioas rex Iudae, postquam mortuus est Ioas filius Ioachaz rex Israel, quindecim annis.
2KGS|14|18|Reliqua autem gestorum Amasiae, nonne haec scripta sunt in libro annalium regum Iudae?
2KGS|14|19|Factaque est contra eum coniuratio in Ierusalem, at ille fugit in Lachis; miseruntque post eum in Lachis et interfecerunt eum ibi.
2KGS|14|20|Et asportaverunt eum in equis; sepultusque est in Ierusalem cum patribus suis in civitate David.
2KGS|14|21|Tulit autem universus populus Iudae Azariam annos natum sedecim, et constituerunt eum regem pro patre eius Amasia.
2KGS|14|22|Ipse aedificavit Ailath et restituit eam Iudae, postquam dormivit rex cum patribus suis.
2KGS|14|23|Anno quinto decimo Amasiae filii Ioas regis Iudae regnavit Ieroboam filius Ioas regis Israel in Samaria quadraginta et uno anno.
2KGS|14|24|Et fecit, quod malum est coram Domino; non recessit ab omnibus peccatis Ieroboam filii Nabat, qui peccare fecit Israel.
2KGS|14|25|Ipse restituit terminos Israel ab introitu Emath usque ad mare Arabae iuxta sermonem Domini, Dei Israel, quem locutus est per servum suum Ionam filium Amathi prophetam, qui erat de Gethhepher.
2KGS|14|26|Vidit enim Dominus afflictionem Israel amaram nimis, et quod consumpti essent impuber et puber, et non esset qui auxiliaretur Israel.
2KGS|14|27|Nec locutus est Dominus, ut deleret nomen Israel de sub caelo, sed salvavit eos in manu Ieroboam filii Ioas.
2KGS|14|28|Reliqua autem gestorum Ieroboam et universa, quae fecit, et fortitudo eius, qua proeliatus est, et quomodo restituit, quod de finibus Damasci et Emath fuerat Iudae, Israeli, nonne haec scripta sunt in libro annalium regum Israel?
2KGS|14|29|Dormivitque Ieroboam cum patribus suis regibus Israel; et regnavit Zacharias filius eius pro eo.
2KGS|15|1|Anno vicesimo septimo Ieroboam regis Israel regnavit Azarias filius Amasiae regis Iudae.
2KGS|15|2|Sedecim annorum erat, cum regnare coepisset, et quinquaginta duobus annis regnavit in Ierusalem. Nomen matris eius Iechelia de Ierusalem.
2KGS|15|3|Fecitque, quod erat placitum coram Domino, iuxta omnia, quae fecit Amasias pater eius.
2KGS|15|4|Verumtamen excelsa non est demolitus; adhuc populus sacrificabat et adolebat in excelsis.
2KGS|15|5|Percussit autem Dominus regem, et fuit leprosus usque in diem mortis suae et habitabat in domo separata seorsum; Ioatham vero filius regis gubernabat palatium et iudicabat populum terrae.
2KGS|15|6|Reliqua autem gestorum Azariae et universa, quae fecit, nonne haec scripta sunt in libro annalium regum Iudae?
2KGS|15|7|Et dormivit Azarias cum patribus suis, sepelieruntque eum cum maioribus suis in civitate David; et regnavit Ioatham filius eius pro eo.
2KGS|15|8|Anno tricesimo octavo Azariae regis Iudae regnavit Zacharias filius Ieroboam super Israel in Samaria sex mensibus.
2KGS|15|9|Et fecit, quod malum est coram Domino, sicut fecerant patres eius; non recessit a peccatis Ieroboam filii Nabat, qui peccare fecit Israel.
2KGS|15|10|Coniuravit autem contra eum Sellum filius Iabes percussitque eum in Ieblaam et interfecit; regnavitque pro eo.
2KGS|15|11|Reliqua autem gestorum Zachariae, nonne haec scripta sunt in libro annalium regum Israel?
2KGS|15|12|Iste est sermo Domini, quem locutus est ad Iehu dicens: " Filii usque ad quartam generationem sedebunt de te super thronum Israel ". Factumque est ita.
2KGS|15|13|Sellum filius Iabes regnavit tricesimo nono anno Azariae regis Iudae; regnavit autem uno mense in Samaria.
2KGS|15|14|Et ascendit Manahem filius Gadi de Thersa venitque Samariam et percussit Sellum filium Iabes in Samaria et interfecit eum; regnavitque pro eo.
2KGS|15|15|Reliqua autem gestorum Sellum et coniuratio eius, per quam tetendit insidias, nonne haec scripta sunt in libro annalium regum Israel?
2KGS|15|16|Tunc percussit Manahem Thapsam et omnes, qui erant in ea, et terminos eius de Thersa; noluerant enim aperire ei. Et interfecit omnes praegnantes eius et scidit eas.
2KGS|15|17|Anno tricesimo nono Azariae regis Iudae regnavit Manahem filius Gadi super Israel decem annis in Samaria.
2KGS|15|18|Fecitque, quod erat malum coram Domino; non recessit a peccatis Ieroboam filii Nabat, qui peccare fecit Israel. In diebus eius
2KGS|15|19|venit Phul rex Assyriorum in terram, et dedit Manahem Phul mille talenta argenti, ut esset ei in auxilio et firmaret regnum eius.
2KGS|15|20|Indixitque Manahem argentum super Israel cunctis potentibus, ut daret regi Assyriorum, quinquaginta siclos argenti per singulos. Reversusque est rex Assyriorum et non est moratus in terra.
2KGS|15|21|Reliqua autem gestorum Manahem et universa, quae fecit, nonne haec scripta sunt in libro annalium regum Israel?
2KGS|15|22|Et dormivit Manahem cum patribus suis; regnavitque Phaceia filius eius pro eo.
2KGS|15|23|Anno quinquagesimo Azariae regis Iudae regnavit Phaceia filius Manahem super Israel in Samaria biennio.
2KGS|15|24|Et fecit, quod erat malum coram Domino; non recessit a peccatis Ieroboam filii Nabat, qui peccare fecit Israel.
2KGS|15|25|Coniuravit autem adversus eum Phacee filius Romeliae dux eius et percussit eum in Samaria in turre domus regiae, et cum eo erant quinquaginta viri de filiis Galaaditarum. Et interfecit eum regnavitque pro eo.
2KGS|15|26|Reliqua autem gestorum Phaceia et universa, quae fecit, nonne haec scripta sunt in libro annalium regum Israel?
2KGS|15|27|Anno quinquagesimo secundo Azariae regis Iudae regnavit Phacee filius Romeliae super Israel in Samaria viginti annis.
2KGS|15|28|Et fecit, quod malum erat coram Domino; non recessit a peccatis Ieroboam filii Nabat, qui peccare fecit Israel.
2KGS|15|29|In diebus Phacee regis Israel venit Theglathphalasar rex Assur et cepit Ahion et Abelbethmaacha et Ianoe et Cedes et Asor et Galaad et Galilaeam, universam terram Nephthali, et transtulit eos in Assur.
2KGS|15|30|Coniuravit autem et tetendit insidias Osee filius Ela contra Phacee filium Romeliae; et percussit eum et interfecit regnavitque pro eo vicesimo anno Ioatham filii Oziae.
2KGS|15|31|Reliqua autem gestorum Phacee et universa, quae fecit, nonne haec scripta sunt in libro annalium regum Israel?
2KGS|15|32|Anno secundo Phacee filii Romeliae regis Israel regnavit Ioatham filius Oziae regis Iudae.
2KGS|15|33|Viginti quinque annorum erat, cum regnare coepisset, et sedecim annis regnavit in Ierusalem. Nomen matris eius Ierusa filia Sadoc.
2KGS|15|34|Fecitque, quod erat placitum coram Domino; iuxta omnia, quae fecerat Ozias pater suus, operatus est.
2KGS|15|35|Verumtamen excelsa non abstulit; adhuc populus immolabat et adolebat in excelsis. Ipse aedificavit portam domus Domini superiorem.
2KGS|15|36|Reliqua autem gestorum Ioatham et universa, quae fecit, nonne haec scripta sunt in libro annalium regum Iudae?
2KGS|15|37|In diebus illis coepit Dominus mittere in Iudam Rasin regem Syriae et Phacee filium Romeliae.
2KGS|15|38|Et dormivit Ioatham cum patribus suis sepultusque est cum eis in civitate David patris sui; et regnavit Achaz filius eius pro eo.
2KGS|16|1|Anno septimo decimo Phacee filii Romeliae regnavit Achaz filius Ioatham regis Iudae.
2KGS|16|2|Viginti annorum erat Achaz, cum regnare coepisset, et sedecim annis regnavit in Ierusalem; non fecit, quod erat placitum in conspectu Domini Dei sui, sicut David pater eius,
2KGS|16|3|sed ambulavit in via regum Israel. Insuper et filium suum consecravit transferens per ignem secundum abominationes gentium, quas dissipavit Dominus coram filiis Israel;
2KGS|16|4|immolabat quoque et adolebat in excelsis et in collibus et sub omni ligno frondoso.
2KGS|16|5|Tunc ascendit Rasin rex Syriae et Phacee filius Romeliae rex Israel in Ierusalem ad proeliandum; cumque obsiderent Achaz, non valuerunt superare eum.
2KGS|16|6|In tempore illo restituit Rasin rex Syriae Ailath ad Edom et eiecit Iudaeos de Ailath; et Idumaei venerunt in Ailath et habitaverunt ibi usque in diem hanc.
2KGS|16|7|Misit autem Achaz nuntios ad Theglathphalasar regem Assyriorum dicens: " Servus tuus et filius tuus ego sum. Ascende et salvum me fac de manu regis Syriae et de manu regis Israel, qui consurrexerunt adversum me ".
2KGS|16|8|Et cum collegisset argentum et aurum, quod invenire potuit in domo Domini et in thesauris regis, misit regi Assyriorum munera.
2KGS|16|9|Qui et acquievit voluntati eius. Ascendit enim rex Assyriorum in Damascum et vastavit eam et transtulit habitatores eius in Cir; Rasin autem interfecit.
2KGS|16|10|Perrexitque rex Achaz in occursum Theglathphalasar regis Assyriorum in Damascum. Cumque vidisset altare Damasci, misit rex Achaz ad Uriam sacerdotem exemplar eius et descriptionem omnis operis eius.
2KGS|16|11|Exstruxitque Urias sacerdos altare; iuxta omnia, quae miserat rex Achaz de Damasco, ita fecit Urias sacerdos, donec veniret rex Achaz de Damasco.
2KGS|16|12|Cumque venisset rex de Damasco, vidit altare et accessit ad illud ascenditque
2KGS|16|13|et adolevit holocausta sua et oblationes et libavit libamina et fudit sanguinem pacificorum suorum super altare.
2KGS|16|14|Porro altare aeneum, quod erat coram Domino, transtulit de facie templi et de loco inter altare et templum Domini posuitque illud ex latere altaris ad aquilonem.
2KGS|16|15|Praecepit quoque rex Achaz Uriae sacerdoti dicens: " Super altare maius offer holocaustum matutinum et oblationem vespertinam et holocaustum regis et oblationem eius et holocaustum universi populi terrae et oblationem eorum et libamina eorum; et omnem sanguinem holocausti et universum sanguinem sacrificii super illud effundes. De altari vero aeneo erit mihi deliberandum ".
2KGS|16|16|Fecit igitur Urias sacerdos iuxta omnia, quae praeceperat rex Achaz.
2KGS|16|17|Excidit autem rex Achaz limbos basium et removit luterem, qui erat desuper, et mare deposuit de bobus aeneis, qui sustentabant illud, et posuit super pavimentum stratum lapide.
2KGS|16|18|Musach (id est Porticum) quoque sabbati, quod aedificatum erat in templo, et ingressum regis exterius convertit in templo Domini propter regem Assyriorum.
2KGS|16|19|Reliqua autem gestorum Achaz, quae fecit, nonne haec scripta sunt in libro annalium regum Iudae?
2KGS|16|20|Dormivitque Achaz cum patribus suis et sepultus est cum eis in civitate David; et regnavit Ezechias filius eius pro eo.
2KGS|17|1|Anno duodecimo Achaz regis Iudae regnavit Osee filius Ela in Samaria super Israel novem annis.
2KGS|17|2|Fecitque malum coram Domino, sed non sicut reges Israel, qui ante eum fuerant.
2KGS|17|3|Contra hunc ascendit Salmanasar rex Assyriorum; et factus est ei Osee servus reddebatque illi tributa.
2KGS|17|4|Cumque deprehendisset rex Assyriorum Osee quod rebellare nitens misisset nuntios ad Sua regem Aegypti nec praestaret tributa regi Assyriorum, sicut singulis annis solitus erat, apprehendit eum et vinctum misit in carcerem.
2KGS|17|5|Pervagatusque est omnem terram et ascendens Samariam obsedit eam tribus annis.
2KGS|17|6|Anno autem nono Osee cepit rex Assyriorum Samariam et transtulit Israel in Assur posuitque eos in Hala et iuxta Habor fluvium Gozan et in civitatibus Medorum.
2KGS|17|7|Factum est enim hoc, cum peccassent filii Israel Domino Deo suo, qui eduxerat eos de terra Aegypti, de manu pharaonis regis Aegypti: coluerunt deos alienos.
2KGS|17|8|Et ambulaverunt iuxta ritus gentium, quas consumpserat Dominus in conspectu filiorum Israel et regum Israel, qui similiter fecerant.
2KGS|17|9|Et offenderunt filii Israel operibus non rectis Dominum Deum suum et aedificaverunt sibi excelsa in cunctis urbibus suis a turre custodum usque ad civitatem munitam.
2KGS|17|10|Feceruntque sibi lapides et palos in omni colle sublimi et subter omne lignum nemorosum
2KGS|17|11|et adolebant ibi in omnibus excelsis sicut gentes, quas transtulerat Dominus a facie eorum; feceruntque pessima irritantes Dominum
2KGS|17|12|et coluerunt idola immunda, de quibus praecepit Dominus eis, ne facerent hoc.
2KGS|17|13|Et testificatus est Dominus in Israel et in Iuda per manum omnium prophetarum et videntium dicens: " Revertimini a viis vestris pessimis et custodite mandata mea et praecepta iuxta omnem legem, quam praecepi patribus vestris, et sicut misi ad vos in manu servorum meorum prophetarum.
2KGS|17|14|Qui non audierunt, sed induraverunt cervicem suam iuxta cervicem patrum suorum, qui noluerunt credere in Dominum Deum suum.
2KGS|17|15|Et abiecerunt legitima eius et pactum, quod pepigit cum patribus eorum, et testificationes, quibus contestatus est eos; secutique sunt vanitates et vani facti sunt et secuti sunt gentes, quae erant per circuitum eorum, super quibus praeceperat Dominus eis ut non facerent, sicut et illae faciebant.
2KGS|17|16|Et dereliquerunt omnia praecepta Domini Dei sui feceruntque sibi conflatiles duos vitulos et palum et adoraverunt universam militiam caeli servieruntque Baal
2KGS|17|17|et consecrabant filios suos et filias suas per ignem; et divinationibus inserviebant et auguriis et tradiderunt se, ut facerent malum coram Domino et irritarent eum.
2KGS|17|18|Iratusque est Dominus vehementer Israel et abstulit eos de conspectu suo, et non remansit nisi tribus Iudae tantummodo.
2KGS|17|19|Sed nec ipse Iuda custodivit mandata Domini Dei sui; verum ambulavit in erroribus Israel, quos operatus fuerat.
2KGS|17|20|Proiecitque Dominus omne semen Israel et afflixit eos et tradidit in manu diripientium, donec proiceret eos a facie sua,
2KGS|17|21|ex eo iam tempore, quo scissus est Israel a domo David, et constituerunt sibi regem Ieroboam filium Nabat; separavit enim Ieroboam Israel a Domino et peccare eos fecit peccatum magnum.
2KGS|17|22|Et ambulaverunt filii Israel in universis peccatis Ieroboam, quae fecerat; non recesserunt ab eis,
2KGS|17|23|usquequo auferret Dominus Israel a facie sua, sicut locutus fuerat in manu omnium servorum suorum prophetarum. Translatusque est Israel de terra sua in Assur usque in diem hanc.
2KGS|17|24|Adduxit autem rex Assyriorum de Babylone et de Chutha et de Ava et de Emath et de Sepharvaim et collocavit eos in civitatibus Samariae pro filiis Israel, qui possederunt Samariam et habitaverunt in urbibus eius.
2KGS|17|25|Cumque ibi habitare coepissent, non timebant Dominum. Et immisit eis Dominus leones, qui interficiebant inter eos.
2KGS|17|26|Nuntiatumque est regi Assyriorum et dictum: " Gentes, quas transtulisti et habitare fecisti in civitatibus Samariae, ignorant legitima Dei terrae; et immisit eis leones, et ecce interficiunt eos, eo quod ignorent ritum Dei terrae ".
2KGS|17|27|Praecepit autem rex Assyriorum dicens: " Ducite illuc unum de sacerdotibus, quos inde captivos adduxistis, et vadat et habitet cum eis et doceat eos legitima Dei terrae ".
2KGS|17|28|Igitur cum venisset unus de sacerdotibus his, qui captivi ducti fuerant de Samaria, habitavit in Bethel et docebat eos quomodo colerent Dominum.
2KGS|17|29|Et unaquaeque gens fabricata est deum suum; posueruntque eos in fanis excelsis, quae fecerant Samaritae, gens et gens in urbibus suis, in quibus habitabant.
2KGS|17|30|Viri enim Babylonii fecerunt Socchothbenoth, viri autem Chutheni fecerunt Nergel, et viri de Emath fecerunt Asima;
2KGS|17|31|porro Hevaei fecerunt Nebahaz et Tharthac, hi autem, qui erant de Sepharvaim, comburebant filios suos igne Adramelech et Anamelech diis Sepharvaim.
2KGS|17|32|Et nihilominus colebant Dominum. Fecerunt autem sibi de medio ipsorum sacerdotes excelsorum et ponebant eos in fanis excelsorum;
2KGS|17|33|et, cum Dominum colerent, diis quoque suis serviebant iuxta consuetudinem gentium, de quibus translati fuerant Samariam.
2KGS|17|34|Usque in praesentem diem morem sequuntur antiquum: non timent Dominum neque custodiunt instituta et iudicium ipsorum et legem et mandatum, quod praeceperat Dominus filiis Iacob, quem cognominavit Israel,
2KGS|17|35|et percusserat cum eis pactum et mandaverat eis dicens: " Nolite timere deos alienos et non adoretis eos neque colatis et non immoletis eis,
2KGS|17|36|sed Dominum, qui eduxit vos de terra Aegypti in fortitudine magna et in brachio extento, ipsum timete, illum adorate et ipsi immolate.
2KGS|17|37|Instituta quoque et iudicia et legem et mandatum, quod scripsit vobis, custodite, ut faciatis cunctis diebus; et non timeatis deos alienos.
2KGS|17|38|Et pactum, quod percussi vobiscum, nolite oblivisci nec timeatis deos alienos,
2KGS|17|39|sed Dominum Deum vestrum timete, et ipse eruet vos de manu omnium inimicorum vestrorum ".
2KGS|17|40|Illi vero non audierunt, sed iuxta consuetudinem suam pristinam perpetrabant.
2KGS|17|41|Fuerunt igitur gentes istae timentes quidem Dominum, sed nihilominus et idolis suis servientes; nam et filii eorum et nepotes, sicut fecerunt parentes sui, ita faciunt usque in praesentem diem.
2KGS|18|1|Anno tertio Osee filii Ela regis Israel regnavit Ezechias filius Achaz regis Iudae.
2KGS|18|2|Viginti quinque annorum erat, cum regnare coepisset, et viginti et novem annis regnavit in Ierusalem. Nomen matris eius Abi filia Zachariae.
2KGS|18|3|Fecitque, quod erat bonum coram Domino, iuxta omnia, quae fecerat David pater suus.
2KGS|18|4|Ipse dissipavit excelsa et contrivit lapides et succidit palum confregitque serpentem aeneum, quem fecerat Moyses; siquidem usque ad illud tempus filii Israel adolebant ei; vocabatur Nohestan.
2KGS|18|5|In Domino, Deo Israel, speravit. Itaque post eum non fuit similis ei de cunctis regibus Iudae sed neque in his, qui ante eum fuerunt.
2KGS|18|6|Et adhaesit Domino et non recessit a vestigiis eius fecitque mandata eius, quae praeceperat Dominus Moysi,
2KGS|18|7|unde et erat Dominus cum eo, et in cunctis, ad quae procedebat, prospere agebat.Rebellavit quoque contra regem Assyriorum et non servivit ei.
2KGS|18|8|Ipse percussit Philisthaeos usque Gazam et terminos eius, a turre custodum usque ad civitatem munitam.
2KGS|18|9|Anno quarto regis Ezechiae, qui erat annus septimus Osee filii Ela regis Israel, ascendit Salmanasar rex Assvriorum Samariam et oppugnavit eam
2KGS|18|10|et cepit. Post annos tres, anno sexto Ezechiae, id est nono anno Osee regis Israel, capta est Samaria.
2KGS|18|11|Et transtulit rex Assyriorum Israel in Assur collocavitque eos in Hala et Habor iuxta fluvium Gozan et in civitatibus Medorum,
2KGS|18|12|quia non audierunt vocem Domini Dei sui, sed praetergressi sunt pactum eius; omnia, quae praeceperat Moyses servus Domini, non audierunt neque fecerunt.
2KGS|18|13|Anno quarto decimo regis Ezechiae ascendit Sennacherib rex Assyriorum ad universas civitates Iudae munitas et cepit eas.
2KGS|18|14|Tunc misit Ezechias rex Iudae nuntios ad regem Assyriorum Lachis dicens: " Peccavi. Recede a me, et omne, quod imposueris mihi, feram ". Indixit itaque rex Assyriorum Ezechiae regi Iudae trecenta talenta argenti et triginta talenta auri;
2KGS|18|15|deditque Ezechias omne argentum, quod repertum fuerat in domo Domini et in thesauris regis.
2KGS|18|16|In tempore illo confregit Ezechias valvas templi Domini et postes, quos ipse inauraverat, et dedit aurum regi Assyriorum.
2KGS|18|17|Misit autem rex Assyriorum Tharthan et Rabsaris et Rabsacen de Lachis ad regem Ezechiam cum manu valida Ierusalem. Qui cum ascendissent, venerunt in Ierusalem et steterunt iuxta aquae ductum piscinae superioris, quae est in via agri fullonis,
2KGS|18|18|vocaveruntque regem. Egressus est autem ad eos Eliachim filius Helciae praepositus domus et Sobna scriba et Ioah filius Asaph a commentariis.
2KGS|18|19|Dixitque ad eos Rabsaces: " Loquimini Ezechiae: Haec dicit rex magnus, rex Assyriorum: Quae est ista fiducia, qua niteris?
2KGS|18|20|Forsitan putas verbum labiorum esse consilium et fortitudinem ad proelium? In quo confidis, ut audeas rebellare contra me?
2KGS|18|21|An speras in baculo arundineo atque confracto, Aegypto, super quem, si incubuerit homo, comminutus ingreditur manum eius et perforabit eam? Sic est pharao rex Aegypti omnibus, qui confidunt in eo.
2KGS|18|22|Quod si dixeritis mihi: "In Domino Deo nostro habemus fiduciam", nonne iste est, cuius abstulit Ezechias excelsa et altaria et praecepit Iudae et Ierusalem: "Ante altare hoc adorabitis in Ierusalem?".
2KGS|18|23|Nunc igitur spondete cum domino meo rege Assyriorum; dabo tibi duo milia equorum; et vide an habere valeas ascensores eorum.
2KGS|18|24|Et quomodo potes in fugam vertere unum satrapam de servis domini mei minimis? An fiduciam habes in Aegypto propter currus et equites?
2KGS|18|25|Numquid sine Domini voluntate ascendi ad locum istum, ut demolirer eum? Dominus dixit mihi: "Ascende ad terram hanc et demolire eam" ".
2KGS|18|26|Dixerunt autem Eliachim filius Helciae et Sobna et Ioah Rabsaci: " Precamur, ut loquaris nobis servis tuis Aramaice, siquidem intellegimus hanc linguam, et non loquaris nobis Iudaice, audiente populo, qui est super murum ".
2KGS|18|27|Responditque eis Rabsaces: " Numquid ad dominum tuum et ad te misit me dominus meus, ut loquerer sermones hos, et non ad viros, qui sedent super murum, ut comedant stercora sua et bibant urinam suam vobiscum? ".
2KGS|18|28|Stetit itaque Rabsaces et clamavit voce magna Iudaice et ait: " Audite verba regis magni, regis Assyriorum:
2KGS|18|29|Haec dicit rex: Non vos seducat Ezechias; non enim poterit eruere vos de manu mea!
2KGS|18|30|Neque fiduciam vobis tribuat super Domino dicens: "Eruens liberabit nos Dominus, et non tradetur civitas haec in manu regis Assyriorum".
2KGS|18|31|Nolite audire Ezechiam! Haec enim dicit rex Assyriorum: Facite mecum benedictionem et egredimini ad me, et comedet unusquisque de vinea sua et de ficu sua, et bibetis aquas de cisternis vestris,
2KGS|18|32|donec veniam et transferam vos in terram, quae similis terrae vestrae est, in terram fructiferam et fertilem vini, terram panis et vinearum, terram olivarum olei ac mellis; et vivetis et non moriemini. Nolite audire Ezechiam, qui vos decipit dicens: "Dominus liberabit nos!".
2KGS|18|33|Numquid liberaverunt dii gentium unusquisque terram suam de manu regis Assyriorum?
2KGS|18|34|Ubi sunt dii Emath et Arphad? Ubi sunt dii Sepharvaim, Ana et Ava? Numquid liberaverunt Samariam de manu mea?
2KGS|18|35|Quinam illi sunt in universis diis terrarum, qui eruerunt regionem suam de manu mea, ut possit eruere Dominus Ierusalem de manu mea? ".
2KGS|18|36|Tacuit itaque populus et non respondit ei quidquam; siquidem praeceptum regis acceperant, ut non responderent ei.
2KGS|18|37|Venitque Eliachim filius Helciae praepositus domus et Sobna scriba et Ioah filius Asaph a commentariis ad Ezechiam, scissis vestibus, et nuntiaverunt ei verba Rabsacis.
2KGS|19|1|Quae cum audisset rex Ezechias, scidit vestimenta sua et opertus est sacco ingressusque est domum Domini.
2KGS|19|2|Et misit Eliachim praepositum domus et Sobnam scribam et senes de sacerdotibus opertos saccis ad Isaiam prophetam filium Amos.
2KGS|19|3|Qui dixerunt: " Haec dicit Ezechias: Dies tribulationis et increpationis et blasphemiae dies iste; venerunt filii usque ad partum, et vires non habet parturiens.
2KGS|19|4|Forte audiet Dominus Deus tuus universa verba Rabsacis, quem misit rex Assyriorum dominus suus, ut exprobraret Deum viventem, et puniet verba, quae audivit Dominus Deus tuus; et fac orationem pro reliquiis, quae remanent ".
2KGS|19|5|Venerunt ergo servi regis Ezechiae ad Isaiam.
2KGS|19|6|Dixitque eis Isaias: " Haec dicetis domino vestro: Haec dicit Dominus: Noli timere a facie sermonum, quos audisti, quibus blasphemaverunt pueri regis Assyriorum me;
2KGS|19|7|ecce ego immittam ei spiritum, et audiet nuntium et revertetur in terram suam; et deiciam eum gladio in terra sua ".
2KGS|19|8|Reversus est igitur Rabsaces et invenit regem Assyriorum oppugnantem Lobnam; audierat enim quod recessisset de Lachis.
2KGS|19|9|Cumque audisset de Tharaca rege Aethiopiae dicentes: " Ecce egressus est, ut pugnet adversum te ", iterum misit nuntios ad Ezechiam dicens:
2KGS|19|10|" Haec dicite Ezechiae regi Iudae: Non te seducat Deus tuus, in quo habes fiduciam, neque dicas: "Non tradetur Ierusalem in manu regis Assyriorum".
2KGS|19|11|Tu enim ipse audisti, quae fecerint reges Assyriorum universis terris, quomodo vastaverint eas. Num ergo solus poteris liberari?
2KGS|19|12|Numquid liberaverunt dii gentium singulos, quos vastaverunt patres mei, Gozan videlicet et Charran et Reseph et filios Eden, qui erant in Thelassar?
2KGS|19|13|Ubi est rex Emath et rex Arphad et rex civitatis Sepharvaim, Ana et Ava? ".
2KGS|19|14|Itaque cum accepisset Ezechias litteras de manu nuntiorum et legisset eas, ascendit in domum Domini et expandit eas coram Domino
2KGS|19|15|et oravit in conspectu eius dicens: " Domine, Deus Israel, qui sedes super cherubim! Tu es Deus solus regnorum omnium terrae, tu fecisti caelum et terram.
2KGS|19|16|Inclina aurem tuam et audi; aperi, Domine, oculos tuos et vide et audi omnia verba Sennacherib, qui misit, ut exprobraret Deum viventem.
2KGS|19|17|Vere, Domine, dissipaverunt reges Assyriorum gentes et terras earum
2KGS|19|18|et miserunt deos eorum in ignem; non enim erant dii, sed opera manuum hominum ex ligno et lapide, et perdiderunt eos.
2KGS|19|19|Nunc igitur, Domine Deus noster, salvos nos fac de manu eius, ut sciant omnia regna terrae quia tu, Domine, es Deus solus ".
2KGS|19|20|Misit autem Isaias filius Amos ad Ezechiam dicens: " Haec dicit Dominus, Deus Israel: Quae deprecatus es me super Sennacherib rege Assyriorum, audivi.
2KGS|19|21|Iste est sermo, quem locutus est Dominus de eo:Sprevit te et subsannavit virgo filia Sion;post tergum tuum caputmovit filia Ierusalem.
2KGS|19|22|Cui exprobrasti et quem blasphemasti?Contra quem exaltasti vocemet elevasti in excelsum oculos tuos? Contra Sanctum Israel!
2KGS|19|23|Per manum servorum tuorumexprobrasti Dominoet dixisti: "In multitudine curruum meorumascendi excelsa montium in summitate Libaniet succidi sublimes cedros eius,electas abietes eius,et ingressus sum usque ad terminos eius,silvam condensam.
2KGS|19|24|Ego fodi et bibi aquas alienaset siccavi vestigiis pedum meorum omnes aquas Aegypti".
2KGS|19|25|Numquid non audisti,ab initio quid fecerim?Ex diebus antiquis plasmavi illudet nunc adduxi;eruntque in eradicationem,in acervos ruinarum civitates munitae.
2KGS|19|26|Et, qui sedent in eis breviata manu,contremuerunt et confusi sunt;facti sunt quasi fenum agriet gramen virens, herba tectorum, quae arefacta est, antequam veniret ad maturitatem.
2KGS|19|27|Sessionem tuamet egressum tuum et introitum tuum ego praesciviet furorem tuum contra me;
2KGS|19|28|insanisti in me,et superbia tua ascendit in aures meas.Ponam itaque circulum in naribus tuiset frenum in labris tuiset reducam te in viam,per quam venisti.
2KGS|19|29|Tibi autem, Ezechia, hoc erit signum:Comede hoc anno, quod reppereris, in secundo autem anno, quae sponte nascuntur;porro in anno tertio seminate et metite,plantate vineas et comedite fructum earum.
2KGS|19|30|Et, quodcumque reliquum fuerit de domo Iudae,mittet radicem deorsumet faciet fructum sursum;
2KGS|19|31|de Ierusalem quippe egredientur reliquiae,et, quod relinquetur, de monte Sion.Zelus Domini exercituum faciet hoc.
2KGS|19|32|Quam ob rem haec dicit Dominus de rege Assyriorum:Non ingredietur urbem hancnec mittet in eam sagittamnec occurret ei clipeonec fundet aggerem circa eam.
2KGS|19|33|Per viam, qua venit, reverteturet civitatem hanc non ingredietur, dicit Dominus.
2KGS|19|34|Protegamque urbem hanc et salvabo eampropter me et propter David servum meum ".
2KGS|19|35|Factum est igitur in nocte illa: egressus est angelus Domini et percussit in castris Assyriorum centum octoginta quinque milia. Cumque diluculo surrexissent, viderunt omnia corpora mortuorum.
2KGS|19|36|Et recedens abiit et reversus est Sennacherib rex Assyriorum et mansit in Nineve.
2KGS|19|37|Cumque adoraret in templo Nesroch dei sui, Adramelech et Sarasar filii eius percusserunt eum gladio fugeruntque in terram Armeniorum. Et regnavit Asarhaddon filius eius pro eo.
2KGS|20|1|In diebus illis aegrotavit Ezechias usque ad mortem. Et venit ad eum Isaias filius Amos prophetes dixitque ei: " Haec dicit Dominus: Dispone domui tuae, morieris enim et non vives ".
2KGS|20|2|Qui convertit faciem suam ad parietem et oravit Dominum dicens:
2KGS|20|3|" Obsecro, Domine, memento quomodo ambulaverim coram te in veritate et in corde perfecto et, quod placitum est coram te, fecerim ". Flevit itaque Ezechias fletu magno.
2KGS|20|4|Et antequam egrederetur Isaias mediam partem atrii, factus est sermo Domini ad eum dicens:
2KGS|20|5|" Revertere et dic Ezechiae duci populi mei: Haec dicit Dominus, Deus David patris tui: Audivi orationem tuam, vidi lacrimam tuam, et ecce sano te; die tertio ascendes templum Domini.
2KGS|20|6|Et addam diebus tuis quindecim annos; sed et de manu regis Assyriorum liberabo te et civitatem hanc et protegam urbem istam propter me et propter David servum meum ".
2KGS|20|7|Dixitque Isaias: " Afferte massam ficorum ". Quam cum attulissent et posuissent super ulcus eius, curatus est.
2KGS|20|8|Dixit autem Ezechias ad Isaiam: " Quod erit signum quia Dominus me sanabit et quia ascensurus sum die tertio templum Domini? ".
2KGS|20|9|Cui ait Isaias: " Hoc erit tibi signum a Domino quod facturus sit Dominus sermonem, quem locutus est: Vis ut accedat umbra decem gradibus, an ut revertatur totidem gradibus? ".
2KGS|20|10|Et ait Ezechias: " Facile est umbram descendere decem gradibus, nec hoc volo ut fiat, sed ut revertatur retrorsum decem gradibus ".
2KGS|20|11|Invocavit itaque Isaias propheta Dominum; et reduxit umbram per gradus, quibus iam descenderat in gradibus Achaz, retrorsum decem gradibus.
2KGS|20|12|In tempore illo misit Merodachbaladan filius Baladan rex Babyloniorum litteras et munera ad Ezechiam; audierat enim quod aegrotasset Ezechias.
2KGS|20|13|Laetatus est autem in adventu eorum Ezechias et ostendit eis totam domum thesauri sui, argentum et aurum et aromata et oleum optimum et domum vasorum suorum et omnia, quae inventa sunt in thesauris suis: non fuit, quod non monstraret eis Ezechias in domo sua et in omni potestate sua.
2KGS|20|14|Venit autem Isaias propheta ad regem Ezechiam dixitque ei: " Quid dixerunt viri isti et unde venerunt ad te? ". Cui ait Ezechias: " De terra longinqua venerunt, de Babylone ".
2KGS|20|15|At ille respondit: " Quid viderunt in domo tua? ". Ait Ezechias: " Omnia, quae sunt in domo mea viderunt; nihil est, quod non monstraverim eis in thesauris meis ".
2KGS|20|16|Dixit itaque Isaias Ezechiae: " Audi sermonem Domini:
2KGS|20|17|Ecce dies venient, et auferentur omnia, quae sunt in domo tua, et quae condiderunt patres tui usque in diem hanc, in Babylone; non remanebit quidquam, ait Dominus.
2KGS|20|18|Sed et de filiis tuis, qui egredientur ex te, quos generabis, tollentur et erunt eunuchi in palatio regis Babylonis ".
2KGS|20|19|Dixit Ezechias ad Isaiam: " Bonus sermo Domini, quem locutus es ". Et ait: " Nonne erit pax et securitas in diebus meis? ".
2KGS|20|20|Reliqua autem gestorum Ezechiae et omnis fortitudo eius, et quomodo fecerit piscinam et aquae ductum et introduxerit aquas in civitatem, nonne haec scripta sunt in libro annalium regum Iudae?
2KGS|20|21|Dormivitque Ezechias cum patribus suis; et regnavit Manasses filius eius pro eo.
2KGS|21|1|Duodecim annorum erat Manasses, cum regnare coe pisset, et quinquaginta quinque annis regnavit in Ierusalem. Nomen matris eius Haphsiba.
2KGS|21|2|Fecitque malum in conspectu Domini iuxta abominationes gentium, quas delevit Dominus a facie filiorum Israel.
2KGS|21|3|Conversusque est et aedificavit excelsa, quae dissipaverat Ezechias pater eius, et erexit aras Baal et fecit palum, sicut fecerat Achab rex Israel, et adoravit omnem militiam caeli et coluit eam.
2KGS|21|4|Exstruxitque aras in domo Domini, de qua dixit Dominus: " In Ierusalem ponam nomen meum ".
2KGS|21|5|Et exstruxit altaria universae militiae caeli in duobus atriis templi Domini
2KGS|21|6|et traduxit filium suum per ignem et hariolatus est et observavit auguria et constituit pythones et haruspices multiplicavit, ut faceret malum coram Domino et irritaret eum.
2KGS|21|7|Posuit quoque palum Aserae, quem fecerat, in templo, super quo locutus est Dominus ad David et ad Salomonem filium eius: " In templo hoc et in Ierusalem, quam elegi de cunctis tribubus Israel, ponam nomen meum in sempiternum;
2KGS|21|8|et ultra non faciam commoveri pedem Israel de terra, quam dedi patribus eorum, sic tamen si custodierint opere omnia, quae praecepi eis, et universam legem, quam mandavit eis servus meus Moyses ".
2KGS|21|9|Illi vero non audierunt, sed seducti sunt a Manasse, ut facerent malum plus quam gentes, quas contrivit Dominus a facie filiorum Israel.
2KGS|21|10|Locutusque est Dominus in manu servorum suorum prophetarum dicens:
2KGS|21|11|" Quia fecit Manasses rex Iudae abominationes istas pessimas super omnia, quae fecerunt Amorraei ante eum, et peccare fecit etiam Iudam in idolis suis,
2KGS|21|12|propterea haec dicit Dominus, Deus Israel: Ecce ego inducam mala super Ierusalem et Iudam, ut quicumque audierit, tinniant ambae aures eius.
2KGS|21|13|Et extendam super Ierusalem funiculum Samariae et pondus domus Achab et extergam Ierusalem sicut qui extergit vas, extergit et convertit super faciem eius.
2KGS|21|14|Et proiciam reliquias hereditatis meae et tradam eas in manu inimicorum eius; eruntque in vastitate et rapina cunctis adversariis suis,
2KGS|21|15|eo quod fecerint malum coram me et perseveraverint irritantes me ex die, qua egressi sunt patres eorum ex Aegypto, usque ad diem hanc ".
2KGS|21|16|Insuper et sanguinem innoxium fudit Manasses multum nimis, donec impleret Ierusalem usque ad summum, absque peccatis suis, quibus peccare fecit Iudam, ut faceret malum coram Domino.
2KGS|21|17|Reliqua autem gestorum Manasse et universa, quae fecit, et peccatum eius, quod peccavit, nonne haec scripta sunt in libro annalium regum Iudae?
2KGS|21|18|Dormivitque Manasses cum patribus suis et sepultus est in horto domus suae, in horto Oza; et regnavit Amon filius eius pro eo.
2KGS|21|19|Viginti et duo annorum erat Amon, cum regnare coepisset, duobusque annis regnavit in Ierusalem. Nomen matris eius Mesallemeth filia Harus de Ieteba.
2KGS|21|20|Fecitque malum in conspectu Domini, sicut fecerat Manasses pater eius,
2KGS|21|21|et ambulavit in omni via, per quam ambulaverat pater eius; servivitque idolis, quibus servierat pater suus, et adoravit ea.
2KGS|21|22|Et dereliquit Dominum, Deum patrum suorum et non ambulavit in via Domini.
2KGS|21|23|Tetenderuntque ei insidias servi sui et interfecerunt regem in domo sua;
2KGS|21|24|percussit autem populus terrae omnes, qui coniuraverant contra regem Amon, et constituerunt sibi regem Iosiam filium eius pro eo.
2KGS|21|25|Reliqua autem gestorum Amon, quae fecit, nonne haec scripta sunt in libro annalium regum Iudae?
2KGS|21|26|Sepelieruntque eum in sepulcro suo in horto Oza; et regnavit Iosias filius eius pro eo.
2KGS|22|1|Octo annorum erat Iosias, cum regnare coepisset, et tri ginta et uno anno regnavit in Ierusalem. Nomen matris eius Idida filia Adaia de Bascath.
2KGS|22|2|Fecitque, quod placitum erat coram Domino, et ambulavit per omnes vias David patris sui; non declinavit ad dexteram sive ad sinistram.
2KGS|22|3|Anno autem octavo decimo regis Iosiae misit rex Saphan filium Eseliae filii Mesullam scribam ad templum Domini dicens ei:
2KGS|22|4|" Vade ad Helciam sacerdotem magnum, ut effundatur pecunia, quae illata est in templum Domini, quam collegerunt ianitores a populo,
2KGS|22|5|deturque opificibus praepositis in domo Domini, qui et distribuent eam his, qui operantur in templo Domini ad instauranda sartatecta templi,
2KGS|22|6|tignariis videlicet et caementariis et his, qui interrupta componunt, et ut emantur ligna et lapides de lapicidinis ad instaurandum templum.
2KGS|22|7|Verumtamen non supputetur eis argentum, quod accipiunt, quia in potestate habent et in fide ".
2KGS|22|8|Dixit autem Helcias pontifex ad Saphan scribam: " Librum legis repperi in domo Domini! ". Deditque Helcias volumen Saphan, qui et legit illud.
2KGS|22|9|Venit quoque Saphan scriba ad regem et renuntiavit ei, quod praeceperat, et ait: " Effuderunt servi tui pecuniam, quae reperta est in domo, et dederunt opificibus praefectis operum templi Domini ".
2KGS|22|10|Narravitque Saphan scriba regi dicens: " Librum dedit mihi Helcias sacerdos ".Quem cum legisset Saphan coram rege,
2KGS|22|11|et audisset rex verba libri legis, scidit vestimenta sua
2KGS|22|12|et praecepit Helciae sacerdoti et Ahicam filio Saphan et Achobor filio Micha et Saphan scribae et Asaiae servo regis dicens:
2KGS|22|13|" Ite et consulite Dominum super me et super populo et super omni Iuda de verbis voluminis istius, quod inventum est; magna enim ira Domini succensa est contra nos, quia non audierunt patres nostri verba libri huius, ut facerent omne, quod scriptum est nobis ".
2KGS|22|14|Ierunt itaque Helcias sacerdos et Ahicam et Achobor et Saphan et Asaia ad Holdam propheten uxorem Sellum filii Thecuae filii Haraas custodis vestium, quae habitabat in Ierusalem in secunda, locutique sunt ad eam,
2KGS|22|15|et illa respondit eis: " Haec dicit Dominus, Deus Israel: Dicite viro, qui misit vos ad me:
2KGS|22|16|Haec dicit Dominus: Ecce ego adducam mala super locum hunc et super habitatores eius omnia verba libri, quae legit rex Iudae,
2KGS|22|17|quia dereliquerunt me et sacrificaverunt diis alienis irritantes me in cunctis operibus manuum suarum; et succendetur indignatio mea in loco hoc et non exstinguetur.
2KGS|22|18|Regi autem Iudae, qui misit vos, ut consuleretis Dominum, sic dicetis: Haec dicit Dominus, Deus Israel: Pro eo quod audisti verba voluminis,
2KGS|22|19|et perterritum est cor tuum, et humiliatus es coram Domino, auditis sermonibus contra locum istum et habitatores eius, quo videlicet fierent in stuporem et in maledictum, et scidisti vestimenta tua et flevisti coram me, et ego audivi, ait Dominus;
2KGS|22|20|idcirco colligam te ad patres tuos, et colligeris ad sepulcrum tuum in pace, ut non videant oculi tui omnia mala, quae inducturus sum super locum istum ". Et renuntiaverunt regi, quod dixerat.
2KGS|23|1|Qui misit, et congregati sunt ad eum omnes senes Iudae et Ierusalem;
2KGS|23|2|ascenditque rex templum Domini et omnes viri Iudae universique, qui habitabant in Ierusalem cum eo, sacerdotes et prophetae et omnis populus a parvo usque ad magnum. Legitque, cunctis audientibus, omnia verba libri foederis, qui inventus est in domo Domini.
2KGS|23|3|Stetitque rex super gradum suum et percussit foedus coram Domino, ut ambularent post Dominum et custodirent praecepta eius et testimonia et legitima in omni corde et in tota anima et suscitarent verba foederis huius, quae scripta erant in libro illo. Acquievitque universus populus pacto.
2KGS|23|4|Et praecepit rex Helciae pontifici et sacerdotibus secundi ordinis et ianitoribus, ut proicerent de templo Domini omnia vasa, quae facta fuerant Baal et Aserae et universae militiae caeli; et combussit ea foris Ierusalem in convalle Cedron et tulit pulverem eorum in Bethel.
2KGS|23|5|Et delevit aedituos, quos posuerant reges Iudae ad sacrificandum in excelsis per civitates Iudae et in circuitu Ierusalem, et eos, qui adolebant Baal et soli et lunae et duodecim signis et omni militiae caeli.
2KGS|23|6|Et efferri fecit palum de domo Domini foras Ierusalem in convalle Cedron et combussit eum ibi et redegit in pulverem et proiecit super sepulcrum vulgi.
2KGS|23|7|Destruxit quoque aediculas prostibulorum, quae erant in domo Domini, in quibus mulieres texebant vestes pro Asera.
2KGS|23|8|Congregavitque omnes sacerdotes de civitatibus Iudae et contaminavit excelsa, ubi sacrificabant sacerdotes, de Gabaa usque Bersabee; et destruxit excelsa pilosorum in introitu portae Iosue principis civitatis, ad sinistram ingredientis portam civitatis.
2KGS|23|9|Verumtamen non ascendebant sacerdotes excelsorum ad altare Domini in Ierusalem, sed tantum comedebant azyma in medio fratrum suorum.
2KGS|23|10|Contaminavit quoque Topheth, quod est in convalle Benennom, ut nemo consecraret filium suum aut filiam per ignem Moloch.
2KGS|23|11|Abstulit quoque equos, quos dederant reges Iudae soli in introitu templi Domini iuxta cubiculum Nathanmelech eunuchi, quod erat in Pharurim; currus autem solis combussit igne.
2KGS|23|12|Altaria quoque, quae erant super tectum cenaculi Achaz, quae fecerant reges Iudae, et altaria, quae fecerat Manasses in duobus atriis templi Domini, destruxit rex et contrivit ea ibi et dispersit cinerem eorum in torrentem Cedron.
2KGS|23|13|Excelsa quoque, quae erant ex adverso Ierusalem ad dexteram partem montis Perditionis, quae aedificaverat Salomon rex Israel Astharoth idolo Sidoniorum et Chamos idolo Moab et Melchom idolo filiorum Ammon, polluit rex;
2KGS|23|14|et contrivit lapides et succidit palos replevitque loca eorum ossibus mortuorum.
2KGS|23|15|Insuper et altare, quod erat in Bethel, excelsum, quod fecerat Ieroboam filius Nabat, qui peccare fecit Israel, etiam altare illud et excelsum destruxit atque combussit et comminuit in pulverem succenditque palum.
2KGS|23|16|Et conversus Iosias vidit ibi sepulcra, quae erant in monte, misitque et tulit ossa de sepulcris et combussit ea super altare et polluit illud iuxta verbum Domini, quod clamaverat vir Dei, cum staret Ieroboam in die festo ad altare. Et conversus elevavit oculos in sepulcrum viri Dei, qui clamaverat verba haec,
2KGS|23|17|et ait: " Quis est titulus ille, quem video? ". Responderuntque ei cives illius urbis: " Sepulcrum est hominis Dei, qui venit de Iuda et clamavit verba haec, quae fecisti super altare Bethel ".
2KGS|23|18|Et ait: " Dimittite eum; nemo commoveat ossa eius ". Et intacta manserunt ossa illius cum ossibus prophetae, qui venerat de Samaria.
2KGS|23|19|Insuper et omnia fana excelsorum, quae erant in civitatibus Samariae, quae fecerant reges Israel ad irritandum Dominum, abstulit Iosias et fecit eis secundum omnia opera, quae fecerat in Bethel.
2KGS|23|20|Et immolavit universos sacerdotes excelsorum, qui erant ibi super altaria, et combussit ossa humana super ea; reversusque est Ierusalem.
2KGS|23|21|Et praecepit omni populo dicens: " Facite Pascha Domino Deo vestro secundum quod scriptum est in libro foederis huius ".
2KGS|23|22|Nec enim factum est Pascha tale a diebus iudicum, qui iudicaverunt Israel, et omnibus diebus regum Israel et regum Iudae,
2KGS|23|23|sicut in octavo decimo anno regis Iosiae factum est Pascha istud Domino in Ierusalem.
2KGS|23|24|Sed et pythones et hariolos et theraphim et idola abominationesque omnes, quae erant in terra Iudae et in Ierusalem, abstulit Iosias, ut statueret verba legis, quae scripta sunt in libro, quem invenit Helcias sacerdos in templo Domini.
2KGS|23|25|Similis illi non fuit ante eum rex, qui reverteretur ad Dominum in omni corde suo et in tota anima sua et in universa virtute sua iuxta omnem legem Moysi, neque post eum surrexit similis illi.
2KGS|23|26|Verumtamen non est aversus Dominus ab ira furoris sui magni, quo iratus est furor eius contra Iudam propter omnes irritationes, quibus provocaverat eum Manasses.
2KGS|23|27|Dixit itaque Dominus: " Etiam Iudam auferam a facie mea, sicut abstuli Israel, et proiciam civitatem hanc, quam elegi, Ierusalem et domum, de qua dixi: Erit nomen meum ibi ".
2KGS|23|28|Reliqua autem gestorum Iosiae et universa, quae fecit, nonne haec scripta sunt in libro annalium regum Iudae?
2KGS|23|29|In diebus eius ascendit pharao Nechao rex Aegypti contra regem Assyriorum ad flumen Euphraten. Et abiit Iosias rex in occursum eius, qui occidit eum in Mageddo, cum vidisset eum.
2KGS|23|30|Et portaverunt eum in curru servi sui mortuum de Mageddo et pertulerunt in Ierusalem et sepelierunt eum in sepulcro suo. Tulitque populus terrae Ioachaz filium Iosiae et unxerunt eum et constituerunt eum regem pro patre suo.
2KGS|23|31|Viginti trium annorum erat Ioachaz, cum regnare coepisset, et tribus mensibus regnavit in Ierusalem. Nomen matris eius Amital filia Ieremiae de Lobna.
2KGS|23|32|Et fecit malum coram Domino iuxta omnia, quae fecerant patres eius.
2KGS|23|33|Vinxitque eum pharao Nechao in Rebla, quae est in terra Emath, ne regnaret in Ierusalem; et imposuit multam terrae centum talentis argenti et talento auri;
2KGS|23|34|regemque constituit pharao Nechao Eliachim filium Iosiae pro Iosia patre eius vertitque nomen eius Ioachim. Porro Ioachaz tulit, et venit in Aegyptum et mortuus est ibi.
2KGS|23|35|Argentum autem et aurum dedit Ioachim pharaoni, cum indixisset terrae, ut conferretur argentum iuxta praeceptum pharaonis; et secundum uniuscuiusque aestimationem exegit tam argentum quam aurum de populo terrae, ut daret pharaoni Nechao.
2KGS|23|36|Viginti quinque annorum erat Ioachim, cum regnare coepisset, et undecim annis regnavit in Ierusalem. Nomen matris eius Zebida filia Phadaia de Ruma.
2KGS|23|37|Et fecit malum coram Domino iuxta omnia, quae fecerant patres eius.
2KGS|24|1|In diebus eius ascendit Nabuchodonosor rex Babylonis, et factus est ei Ioachim servus tribus annis et rursum rebellavit contra eum.
2KGS|24|2|Immisitque ei Dominus turmas Chaldaeorum et turmas Syriae, turmas Moab et turmas filiorum Ammon; et immisit eas in Iudam, ut disperderent eum iuxta verbum Domini, quod locutus erat per servos suos prophetas.
2KGS|24|3|Factum est autem hoc propter iram Domini contra Iudam, ut auferret eum de conspectu suo propter peccata Manasse universa, quae fecit,
2KGS|24|4|et propter sanguinem innoxium, quem effudit et implevit Ierusalem cruore innocentium; et ob hanc rem noluit Dominus propitiari.
2KGS|24|5|Reliqua autem gestorum Ioachim et universa, quae fecit, nonne haec scripta sunt in libro annalium regum Iudae? Et dormivit Ioachim cum patribus suis;
2KGS|24|6|regnavitque Ioachin filius eius pro eo.
2KGS|24|7|Et ultra non addidit rex Aegypti ut egrederetur de terra sua; tulerat enim rex Babylonis a rivo Aegypti usque ad fluvium Euphraten omnia, quae fuerant regis Aegypti.
2KGS|24|8|Decem et octo annorum erat Ioachin, cum regnare coepisset, et tribus mensibus regnavit in Ierusalem. Nomen matris eius Naestha filia Elnathan de Ierusalem.
2KGS|24|9|Et fecit malum coram Domino iuxta omnia, quae fecerat pater eius.
2KGS|24|10|In tempore illo ascenderunt servi Nabuchodonosor regis Babylonis in Ierusalem, et venit urbs in obsidione.
2KGS|24|11|Venitque Nabuchodonosor rex Babylonis ad civitatem, cum servi eius oppugnarent eam;
2KGS|24|12|egressusque est Ioachin rex Iudae ad regem Babylonis ipse et mater eius et servi eius et principes eius et eunuchi eius; et cepit eum rex Babylonis anno octavo regni sui.
2KGS|24|13|Et protulit inde omnes thesauros domus Domini et thesauros domus regiae et concidit universa vasa aurea, quae fecerat Salomon rex Israel in templo Domini, iuxta verbum Domini.
2KGS|24|14|Et transtulit omnem Ierusalem et universos principes et omnes fortes exercitus decem milia in captivitatem et omnem artificem et clusorem; nihilque relictum est, exceptis pauperibus populi terrae.
2KGS|24|15|Transtulit quoque Ioachin in Babylonem; et matrem regis et uxores regis et eunuchos eius et cives validos terrae duxit in captivitatem de Ierusalem in Babylonem
2KGS|24|16|et omnes viros robustos septem milia et artifices et clusores mille, omnes viros fortes bellatores; duxitque eos rex Babylonis captivos in Babylonem.
2KGS|24|17|Et constituit Matthaniam patruum eius pro eo; imposuitque nomen ei Sedeciam.
2KGS|24|18|Vicesimum et primum annum aetatis habebat Sedecias, cum regnare coepisset, et undecim annis regnavit in Ierusalem. Nomen matris eius erat Amital filia Ieremiae de Lobna.
2KGS|24|19|Et fecit malum coram Domino iuxta omnia, quae fecerat Ioachim;
2KGS|24|20|irascebatur enim Dominus contra Ierusalem et contra Iudam, donec proiceret eos a facie sua.Recessitque Sedecias a rege Babylonis.
2KGS|25|1|Factum est autem anno nono regni eius, mense decimo, decima die mensis venit Nabuchodonosor rex Babylonis ipse et omnis exercitus eius in Ierusalem; et circumdederunt eam et exstruxerunt in circuitu eius munitiones.
2KGS|25|2|Et clausa est civitas atque vallata usque ad undecimum annum regis Sedeciae.
2KGS|25|3|Nona die mensis quarti praevaluit fames in civitate, nec erat panis populo terrae.
2KGS|25|4|Et interrupta est civitas, et omnes viri bellatores fugerunt exieruntque de civitate nocte per viam portae, quae est inter duplicem murum ad hortum regis, obsidentibus Chaldaeis in circuitu civitatem. Abierunt itaque per viam, quae ducit ad Arabam.
2KGS|25|5|Et persecutus est exercitus Chaldaeorum regem comprehenditque eum in planitie Iericho, et omnis exercitus eius dispersus est et reliquit eum.
2KGS|25|6|Apprehensum ergo regem duxerunt ad regem Babylonis in Rebla, qui locutus est cum eo iudicium.
2KGS|25|7|Filios autem Sedeciae occidit coram eo et oculos eius effodit vinxitque eum catenis aereis et adduxit in Babylonem.
2KGS|25|8|Mense quinto septima die mensis, ipse est annus nonus decimus regis Babylonis, venit Nabuzardan princeps satellitum servus regis Babylonis Ierusalem
2KGS|25|9|et succendit domum Domini et domum regis et omnes domos Ierusalem; omnemque domum combussit igne.
2KGS|25|10|Et muros Ierusalem in circuitu destruxit omnis exercitus Chaldaeorum, qui erat cum principe satellitum.
2KGS|25|11|Reliquam autem populi partem, qui remanserat in civitate, et perfugas, qui transfugerant ad regem Babylonis, et reliquum vulgus transtulit Nabuzardan princeps satellitum;
2KGS|25|12|et de pauperibus terrae reliquit in vinitores et agricolas.
2KGS|25|13|Columnas autem aereas, quae erant in templo Domini, et bases et mare aereum, quod erat in domo Domini, confregerunt Chaldaei et transtulerunt aes omnium in Babylonem.
2KGS|25|14|Ollas quoque et trullas et cultros et phialas et omnia vasa aerea, in quibus ministrabant, tulerunt;
2KGS|25|15|necnon thymiamateria et phialas, quae aurea aurea et quae argentea argentea, tulit princeps satellitum;
2KGS|25|16|columnas duas, mare unum et bases, quas fecerat Salomon templo Domini; non erat pondus aeris omnium horum vasorum.
2KGS|25|17|Decem et octo cubitos altitudinis habebat columna una et capitellum aereum super se altitudinis quinque cubitorum; et reticulum et malogranata super capitellum in circuitu omnia aerea; similem et columna secunda habebat ornatum.
2KGS|25|18|Tulit quoque princeps satellitum Saraiam sacerdotem primum et Sophoniam sacerdotem secundum et tres ianitores
2KGS|25|19|et de civitate eunuchum unum, qui erat praefectus super viros bellatores, et quinque viros de his, qui steterant coram rege, quos repperit in civitate, et scribam principis exercitus, qui probabat tirones de populo terrae, et sexaginta viros e populo terrae, qui inventi fuerant in civitate;
2KGS|25|20|quos tollens Nabuzardan princeps satellitum duxit ad regem Babylonis in Rebla,
2KGS|25|21|percussitque eos rex Babylonis et interfecit in Rebla in terra Emath.Et translatus est Iuda de terra sua.
2KGS|25|22|Populo autem, qui relictus erat in terra Iudae, quem dimiserat Nabuchodonosor rex Babylonis, praefecit Godoliam filium Ahicam filii Saphan.
2KGS|25|23|Quod cum audissent omnes duces militum, videlicet quod constituisset rex Babylonis Godoliam, ipsi et viri, qui erant cum eis, venerunt ad Godoliam in Maspha: Ismael filius Nathaniae et Iohanan filius Caree et Saraia filius Thanehumeth Netophathites et Iezonias filius Maachathitis, ipsi et socii eorum.
2KGS|25|24|Iuravitque eis Godolias et sociis eorum dicens: " Nolite timere a servis Chaldaeorum; manete in terra et servite regi Babylonis, et bene erit vobis ".
2KGS|25|25|Factum est autem in mense septimo venit Ismael filius Nathaniae filii Elisama de semine regio et decem viri cum eo; percusseruntque Godoliam, qui mortuus est, sed et Iudaeos et Chaldaeos, qui erant cum eo in Maspha.
2KGS|25|26|Consurgens autem populus a parvo usque ad magnum et principes militum venerunt in Aegyptum timentes Chaldaeos.
2KGS|25|27|Factum est vero anno tricesimo septimo transmigrationis Ioachin regis Iudae, mense duodecimo vicesima septima die mensis sublevavit Evilmerodach rex Babylonis anno, quo regnare coeperat, caput Ioachin regis Iudae de carcere.
2KGS|25|28|Et locutus est ei benigna et posuit thronum eius super thronos regum, qui erant cum eo in Babylone,
2KGS|25|29|et mutavit vestes eius, quas habuerat in carcere; et comedebat panem semper in conspectu eius cunctis diebus vitae suae.
2KGS|25|30|Annonam quoque constituit ei absque intermissione, quae et dabatur ei a rege per singulos dies omnibus diebus vitae suae.
