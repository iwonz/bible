HAG|1|1|In the second year of Darius the king, in the sixth month, on the first day of the month, the word of the LORD came by the hand of Haggai the prophet to Zerubbabel the son of Shealtiel, governor of Judah, and to Joshua the son of Jehozadak, the high priest:
HAG|1|2|"Thus says the LORD of hosts: These people say the time has not yet come to rebuild the house of the LORD."
HAG|1|3|Then the word of the LORD came by the hand of Haggai the prophet,
HAG|1|4|"Is it a time for you yourselves to dwell in your paneled houses, while this house lies in ruins?
HAG|1|5|Now, therefore, thus says the LORD of hosts: Consider your ways.
HAG|1|6|You have sown much, and harvested little. You eat, but you never have enough; you drink, but you never have your fill. You clothe yourselves, but no one is warm. And he who earns wages does so to put them into a bag with holes.
HAG|1|7|"Thus says the LORD of hosts: Consider your ways.
HAG|1|8|Go up to the hills and bring wood and build the house, that I may take pleasure in it and that I may be glorified, says the LORD.
HAG|1|9|You looked for much, and behold, it came to little. And when you brought it home, I blew it away. Why? declares the LORD of hosts. Because of my house that lies in ruins, while each of you busies himself with his own house.
HAG|1|10|Therefore the heavens above you have withheld the dew, and the earth has withheld its produce.
HAG|1|11|And I have called for a drought on the land and the hills, on the grain, the new wine, the oil, on what the ground brings forth, on man and beast, and on all their labors."
HAG|1|12|Then Zerubbabel the son of Shealtiel, and Joshua the son of Jehozadak, the high priest, with all the remnant of the people, obeyed the voice of the LORD their God, and the words of Haggai the prophet, as the LORD their God had sent him. And the people feared the LORD.
HAG|1|13|Then Haggai, the messenger of the LORD, spoke to the people with the LORD's message, "I am with you, declares the LORD."
HAG|1|14|And the LORD stirred up the spirit of Zerubbabel the son of Shealtiel, governor of Judah, and the spirit of Joshua the son of Jehozadak, the high priest, and the spirit of all the remnant of the people. And they came and worked on the house of the LORD of hosts, their God,
HAG|1|15|on the twenty-fourth day of the month, in the sixth month, in the second year of Darius the king.
HAG|2|1|In the seventh month, on the twenty-first day of the month, the word of the LORD came by the hand of Haggai the prophet,
HAG|2|2|"Speak now to Zerubbabel the son of Shealtiel, governor of Judah, and to Joshua the son of Jehozadak, the high priest, and to all the remnant of the people, and say,
HAG|2|3|'Who is left among you who saw this house in its former glory? How do you see it now? Is it not as nothing in your eyes?
HAG|2|4|Yet now be strong, O Zerubbabel, declares the LORD. Be strong, O Joshua, son of Jehozadak, the high priest. Be strong, all you people of the land, declares the LORD. Work, for I am with you, declares the LORD of hosts,
HAG|2|5|according to the covenant that I made with you when you came out of Egypt. My Spirit remains in your midst. Fear not.
HAG|2|6|For thus says the LORD of hosts: Yet once more, in a little while, I will shake the heavens and the earth and the sea and the dry land.
HAG|2|7|And I will shake all nations, so that the treasures of all nations shall come in, and I will fill this house with glory, says the LORD of hosts.
HAG|2|8|The silver is mine, and the gold is mine, declares the LORD of hosts.
HAG|2|9|The latter glory of this house shall be greater than the former, says the LORD of hosts. And in this place I will give peace, declares the LORD of hosts.'"
HAG|2|10|On the twenty-fourth day of the ninth month, in the second year of Darius, the word of the LORD came by Haggai the prophet,
HAG|2|11|"Thus says the LORD of hosts: Ask the priests about the law:
HAG|2|12|'If someone carries holy meat in the fold of his garment and touches with his fold bread or stew or wine or oil or any kind of food, does it become holy?'" The priests answered and said, "No."
HAG|2|13|Then Haggai said, "If someone who is unclean by contact with a dead body touches any of these, does it become unclean?" The priests answered and said, "It does become unclean."
HAG|2|14|Then Haggai answered and said, "So is it with this people, and with this nation before me, declares the LORD, and so with every work of their hands. And what they offer there is unclean.
HAG|2|15|Now then, consider from this day onward. Before stone was placed upon stone in the temple of the LORD,
HAG|2|16|how did you fare? When one came to a heap of twenty measures, there were but ten. When one came to the wine vat to draw fifty measures, there were but twenty.
HAG|2|17|I struck you and all the products of your toil with blight and with mildew and with hail, yet you did not turn to me, declares the LORD.
HAG|2|18|Consider from this day onward, from the twenty-fourth day of the ninth month. Since the day that the foundation of the LORD's temple was laid, consider:
HAG|2|19|Is the seed yet in the barn? Indeed, the vine, the fig tree, the pomegranate, and the olive tree have yielded nothing. But from this day on I will bless you."
HAG|2|20|The word of the LORD came a second time to Haggai on the twenty-fourth day of the month,
HAG|2|21|"Speak to Zerubbabel, governor of Judah, saying, I am about to shake the heavens and the earth,
HAG|2|22|and to overthrow the throne of kingdoms. I am about to destroy the strength of the kingdoms of the nations, and overthrow the chariots and their riders. And the horses and their riders shall go down, every one by the sword of his brother.
HAG|2|23|On that day, declares the LORD of hosts, I will take you, O Zerubbabel my servant, the son of Shealtiel, declares the LORD, and make you like a signet ring, for I have chosen you, declares the LORD of hosts."
