HAB|1|1|onus quod vidit Abacuc propheta
HAB|1|2|usquequo Domine clamabo et non exaudies vociferabor ad te vim patiens et non salvabis
HAB|1|3|quare ostendisti mihi iniquitatem et laborem videre praeda et iniustitia contra me et factum est iudicium et contradictio potentior
HAB|1|4|propter hoc lacerata est lex et non pervenit usque ad finem iudicium quia impius praevalet adversus iustum propterea egreditur iudicium perversum
HAB|1|5|aspicite in gentibus et videte et admiramini et obstupescite quia opus factum est in diebus vestris quod nemo credet cum narrabitur
HAB|1|6|quia ecce ego suscitabo Chaldeos gentem amaram et velocem ambulantem super latitudinem terrae ut possideat tabernacula non sua
HAB|1|7|horribilis et terribilis est ex semet ipsa iudicium et onus eius egredietur
HAB|1|8|leviores pardis equi eius et velociores lupis vespertinis et diffundentur equites eius equites namque eius de longe venient volabunt quasi aquila festinans ad comedendum
HAB|1|9|omnes ad praedam venient facies eorum ventus urens et congregabit quasi harenam captivitatem
HAB|1|10|et ipse de regibus triumphabit et tyranni ridiculi eius erunt ipse super omnem munitionem ridebit et conportabit aggerem et capiet eam
HAB|1|11|tunc mutabitur spiritus et pertransibit et corruet haec est fortitudo eius dei sui
HAB|1|12|numquid non tu a principio Domine Deus meus Sancte meus et non moriemur Domine in iudicium posuisti eum et fortem ut corriperes fundasti eum
HAB|1|13|mundi sunt oculi tui ne videas malum et respicere ad iniquitatem non poteris quare non respicis super inique agentes et taces devorante impio iustiorem se
HAB|1|14|et facies homines quasi pisces maris et quasi reptile non habens principem
HAB|1|15|totum in hamo sublevavit traxit illud in sagena sua et congregavit in rete suo super hoc laetabitur et exultabit
HAB|1|16|propterea immolabit sagenae suae et sacrificabit reti suo quia in ipsis incrassata est pars eius et cibus eius electus
HAB|1|17|propter hoc ergo expandit sagenam suam et semper interficere gentes non parcet
HAB|2|1|super custodiam meam stabo et figam gradum super munitionem et contemplabor ut videam quid dicatur mihi et quid respondeam ad arguentem me
HAB|2|2|et respondit mihi Dominus et dixit scribe visum et explana eum super tabulas ut percurrat qui legerit eum
HAB|2|3|quia adhuc visus procul et apparebit in finem et non mentietur si moram fecerit expecta illum quia veniens veniet et non tardabit
HAB|2|4|ecce qui incredulus est non erit recta anima eius in semet ipso iustus autem in fide sua vivet
HAB|2|5|et quomodo vinum potantem decipit sic erit vir superbus et non decorabitur qui dilatavit quasi infernus animam suam et ipse quasi mors et non adimpletur et congregabit ad se omnes gentes et coacervabit ad se omnes populos
HAB|2|6|numquid non omnes isti super eum parabolam sument et loquellam enigmatum eius et dicetur vae ei qui multiplicat non sua usquequo et adgravat contra se densum lutum
HAB|2|7|numquid non repente consurgent qui mordeant te et suscitabuntur lacerantes te et eris in rapinam eis
HAB|2|8|quia tu spoliasti gentes multas spoliabunt te omnes qui reliqui fuerint de populis propter sanguinem hominis et iniquitatem terrae civitatis et omnium habitantium in ea
HAB|2|9|vae qui congregat avaritiam malam domui suae ut sit in excelso nidus eius et liberari se putat de manu mali
HAB|2|10|cogitasti confusionem domui tuae concidisti populos multos et peccavit anima tua
HAB|2|11|quia lapis de pariete clamabit et lignum quod inter iuncturas aedificiorum est respondebit
HAB|2|12|vae qui aedificat civitatem in sanguinibus et praeparat urbem in iniquitate
HAB|2|13|numquid non haec a Domino sunt exercituum laborabunt enim populi in multo igni et gentes in vacuum et deficient
HAB|2|14|quia replebitur terra ut cognoscat gloriam Domini quasi aquae operientes mare
HAB|2|15|vae qui potum dat amico suo mittens fel suum et inebrians ut aspiciat nuditatem eius
HAB|2|16|repletus est ignominia pro gloria bibe tu quoque et consopire circumdabit te calix dexterae Domini et vomitus ignominiae super gloriam tuam
HAB|2|17|quia iniquitas Libani operiet te et vastitas animalium deterrebit eos de sanguinibus hominis et iniquitate terrae et civitatis et omnium habitantium in ea
HAB|2|18|quid prodest sculptile quia sculpsit illud fictor suus conflatile et imaginem falsam quia speravit in figmento fictor eius ut faceret simulacra muta
HAB|2|19|vae qui dicit ligno expergiscere surge lapidi tacenti numquid ipse docere poterit ecce iste coopertus est auro et argento et omnis spiritus non est in visceribus eius
HAB|2|20|Dominus autem in templo sancto suo sileat a facie eius omnis terra
HAB|3|1|oratio Abacuc prophetae pro ignorationibus
HAB|3|2|Domine audivi auditionem tuam et timui Domine opus tuum in medio annorum vivifica illud in medio annorum notum facies cum iratus fueris misericordiae recordaberis
HAB|3|3|Deus ab austro veniet et Sanctus de monte Pharan semper operuit caelos gloria eius et laudis eius plena est terra
HAB|3|4|splendor eius ut lux erit cornua in manibus eius ibi abscondita est fortitudo eius
HAB|3|5|ante faciem eius ibit mors et egredietur diabolus ante pedes eius
HAB|3|6|stetit et mensus est terram aspexit et dissolvit gentes et contriti sunt montes saeculi incurvati sunt colles mundi ab itineribus aeternitatis eius
HAB|3|7|pro iniquitate vidi tentoria Aethiopiae turbabuntur pelles terrae Madian
HAB|3|8|numquid in fluminibus iratus es Domine aut in fluminibus furor tuus vel in mari indignatio tua quia ascendes super equos tuos et quadrigae tuae salvatio
HAB|3|9|suscitans suscitabis arcum tuum iuramenta tribubus quae locutus es semper fluvios scindes terrae
HAB|3|10|viderunt te et doluerunt montes gurges aquarum transiit dedit abyssus vocem suam altitudo manus suas levavit
HAB|3|11|sol et luna steterunt in habitaculo suo in luce sagittarum tuarum ibunt in splendore fulgurantis hastae tuae
HAB|3|12|in fremitu conculcabis terram in furore obstupefacies gentes
HAB|3|13|egressus es in salutem populi tui in salutem cum christo tuo percussisti caput de domo impii denudasti fundamentum usque ad collum semper
HAB|3|14|maledixisti sceptris eius capiti bellatorum eius venientibus ut turbo ad dispergendum me exultatio eorum sicut eius qui devorat pauperem in abscondito
HAB|3|15|viam fecisti in mari equis tuis in luto aquarum multarum
HAB|3|16|audivi et conturbatus est venter meus ad vocem contremuerunt labia mea ingrediatur putredo in ossibus meis et subter me scateat ut requiescam in die tribulationis ut ascendam ad populum accinctum nostrum
HAB|3|17|ficus enim non florebit et non erit germen in vineis mentietur opus olivae et arva non adferent cibum abscidetur de ovili pecus et non erit armentum in praesepibus
HAB|3|18|ego autem in Domino gaudebo exultabo in Deo Iesu meo
HAB|3|19|Dominus Deus fortitudo mea et ponet pedes meos quasi cervorum et super excelsa mea deducet me victori in psalmis canentem
