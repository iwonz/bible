JOSH|1|1|耶和華的僕人 摩西 死了以後，耶和華對 摩西 的助手 嫩 的兒子 約書亞 說：
JOSH|1|2|「我的僕人 摩西 死了。現在你要起來，和眾百姓過這 約旦河 ，往我所要賜給 以色列 人的地去。
JOSH|1|3|凡你們腳掌所踏之地，我都照我所應許 摩西 的話賜給你們了。
JOSH|1|4|從曠野和這 黎巴嫩 ，直到 大河 ，就是 幼發拉底河 ， 赫 人的全地，又到 大海 日落的方向，都要作你們的疆土。
JOSH|1|5|你一生的日子，必無人能在你面前站立得住。我怎樣與 摩西 同在，也必照樣與你同在；我必不撇下你，也不丟棄你。
JOSH|1|6|你當剛強壯膽，因為你必使這百姓承受那地為業，就是我向他們列祖起誓要給他們的地。
JOSH|1|7|只要剛強，大大壯膽，謹守遵行我僕人 摩西 所吩咐你的一切律法，不可偏離左右，使你無論往哪裏去， 都可以順利。
JOSH|1|8|這律法書不可離開你的口，總要晝夜思想 ，好使你謹守遵行這書上所寫的一切話。如此，你的道路就可以亨通，凡事順利。
JOSH|1|9|我豈沒有吩咐你嗎？你當剛強壯膽，不要懼怕，也不要驚惶，因為你無論往哪裏去，耶和華你的上帝必與你同在。」
JOSH|1|10|於是， 約書亞 吩咐百姓的官長說：
JOSH|1|11|「你們要走遍營中，吩咐百姓說：『當預備食物， 因為三日之內你們要過這 約旦河 ，進去得耶和華－你們上帝賜給你們為業之地。』」
JOSH|1|12|約書亞 對 呂便 人、 迦得 人和 瑪拿西 半支派的人說：
JOSH|1|13|「你們要記得耶和華的僕人 摩西 所吩咐你們的話說：『耶和華－你們的上帝使你們得享安寧，必將這地賜給你們。』
JOSH|1|14|你們的妻子、孩子和牲畜可以留在 約旦河 東、 摩西 所給你們的地。但你們中間所有大能的勇士都要帶著兵器，在你們的弟兄前面過去，你們要幫助他們。
JOSH|1|15|等到耶和華使你們的弟兄和你們一樣得享平靜，並且得著耶和華－你們上帝所賜他們為業之地的時候，你們才可以回到你們所得之地，承受為業，就是耶和華的僕人 摩西 在 約旦河 東、向日出的方向所給你們的地。」
JOSH|1|16|他們回答 約書亞 說：「凡你吩咐我們的，我們都必做；凡你差我們去的地方，我們都必去。
JOSH|1|17|我們在一切事上怎樣聽從 摩西 ，也必照樣聽從你。惟願耶和華－你的上帝與你同在，像與 摩西 同在一樣。
JOSH|1|18|無論甚麼人違背你的命令，不聽從你所吩咐他的一切話，就必處死。你只要剛強壯膽！」
JOSH|2|1|嫩 的兒子 約書亞 從 什亭 暗中派兩個人作探子，說：「你們去窺探那地和 耶利哥 。」於是二人去了，來到一個名叫 喇合 的妓女家裏，在那裏睡覺。
JOSH|2|2|有人告訴 耶利哥 王說：「看哪，今夜有 以色列 人到這裏來窺探此地。」
JOSH|2|3|耶利哥 王派人到 喇合 那裏， 說：「你要交出那來到你這裏、進了你家的人，因為他們來是要窺探全地。」
JOSH|2|4|但女人已把二人藏起來，卻說：「那兩個人確實到我這裏來過，他們從哪裏來，我卻不知道。
JOSH|2|5|天黑、要關城門的時候，他們就出去了。他們往哪裏去我也不知道。你們趕快去追他們，就必追上。」
JOSH|2|6|其實，這女人已經領二人上了屋頂，把他們藏在她擺列在屋頂的的亞麻梗中。
JOSH|2|7|那些人就往 約旦河 的路上追趕他們，直到渡口。追趕他們的人一出去，城門就關了。
JOSH|2|8|二人還沒有睡之前，女人就上屋頂，到他們那裏，
JOSH|2|9|對他們說：「我知道耶和華已經把這地賜給你們了，並且我們也都懼怕你們。這地所有的居民在你們面前都融化了。
JOSH|2|10|因為我們聽見你們出 埃及 的時候，耶和華怎樣在你們前面使 紅海 的水乾了，並且你們怎樣處置 約旦河 東的兩個 亞摩利 王， 西宏 和 噩 ，把他們完全消滅。
JOSH|2|11|我們一聽見就膽戰心驚 ，人人因你們的緣故勇氣全失。耶和華－你們的上帝是天上地下的上帝。
JOSH|2|12|現在我既然恩待你們，求你們指著耶和華向我起誓，你們也要恩待我的父家。請你們給我一個確實的憑據，
JOSH|2|13|要救活我的父母、兄弟、姊妹，和所有屬他們的，拯救我們的性命脫離死亡。」
JOSH|2|14|那二人對她說：「我們願意以性命來替你們死。你們若不洩漏我們這件事，當耶和華將這地賜給我們的時候，我們必以慈愛和誠信待你。」
JOSH|2|15|於是女人用繩子把二人從窗戶縋下去，因為她的屋子是在城牆邊上，她也住在城牆上。
JOSH|2|16|她對他們說：「你們暫且往山上去，免得追趕的人遇見你們。要在那裏躲藏三天，等追趕的人回來，你們才可以走自己的路。」
JOSH|2|17|二人對她說：「你叫我們所起的誓與我們無關，
JOSH|2|18|除非，看哪，當我們來到這地的時候，你把這條朱紅線繩子繫在縋我們下去的窗戶上，並要叫你的父母、兄弟和你父的全家都聚集在你家中。
JOSH|2|19|凡離開你家門往街上去的，他的血必歸到自己頭上，與我們無關；凡在你家裏的，若有人下手害他，他的血就歸到我們頭上。
JOSH|2|20|你若洩漏我們這件事，你叫我們所起的誓 就與我們無關了。」
JOSH|2|21|女人說：「就照你們的話吧！」於是她送他們走了，就把朱紅繩子繫在窗戶上。
JOSH|2|22|二人離開，到山上去，在那裏停留三天，直等到追趕的人回去。追趕的人一路尋找，卻找不著。
JOSH|2|23|二人回來，下了山，過了河，來到 嫩 的兒子 約書亞 那裏，向他報告他們所遭遇的一切事。
JOSH|2|24|他們對 約書亞 說：「耶和華果然將那全地交在我們手中了，並且那地所有的居民在我們面前都融化了。」
JOSH|3|1|約書亞 清早起來，和 以色列 眾人起行，離開 什亭 ，來到 約旦河 ，過河以前住在那裏。
JOSH|3|2|過了三天，官長走遍營中，
JOSH|3|3|吩咐百姓說：「當你們看見 利未 家的祭司抬著耶和華－你們上帝的約櫃的時候，你們就要起行離開所住的地方，跟著約櫃走，
JOSH|3|4|使你們知道所當走的路，因為這條路是你們從來沒有走過的。只是你們要與約櫃相隔約二千肘，不可太靠近約櫃。」
JOSH|3|5|約書亞 吩咐百姓說：「你們要使自己分別為聖，因為明天耶和華必在你們中間行奇事。」
JOSH|3|6|約書亞 對祭司說：「你們抬起約櫃，在百姓的前面過去。」於是他們抬起約櫃，走在百姓前面。
JOSH|3|7|耶和華對 約書亞 說：「從今日起，我必使你在 以色列 眾人眼前被尊為大，使他們知道我怎樣與 摩西 同在，也必照樣與你同在。
JOSH|3|8|你要吩咐抬約櫃的祭司說：『你們到了 約旦河 的水邊，要在 約旦河 中站著。』」
JOSH|3|9|約書亞 對 以色列 人說：「你們近前，到這裏來，聽耶和華－你們上帝的話。」
JOSH|3|10|約書亞 說：「你們因這事會知道永生的上帝在你們中間，他必從你們面前趕出 迦南 人、 赫 人、 希未 人、 比利洗 人、 革迦撒 人、 亞摩利 人、 耶布斯 人。
JOSH|3|11|看哪！全地之主的約櫃必在你們的前面過去，到 約旦河 裏。
JOSH|3|12|現在， 你們要從 以色列 支派中選出十二個人，每支派一人。
JOSH|3|13|當抬耶和華全地之主約櫃的祭司，腳掌踏入 約旦河 水裏的時候， 約旦河 的水，就是從上往下流的水，必然中斷，豎立成壘。」
JOSH|3|14|百姓起行離開帳棚過 約旦河 的時候，抬約櫃的祭司在百姓的前面。
JOSH|3|15|那時正是收割的日子， 約旦河 的水漲滿兩岸。抬約櫃的人到了 約旦河 ，抬約櫃的祭司腳一入水邊，
JOSH|3|16|那從上往下流的水就在很遠的地方，在 撒拉但 旁邊的 亞當城 那裏停住，豎立成壘；那往 亞拉巴海 ，就是 鹽海 下流的水全然中斷。於是，百姓在 耶利哥 的對面過了河。
JOSH|3|17|抬耶和華約櫃的祭司在 約旦河 中的乾地上穩穩站著， 以色列 眾人都從乾地上過去，直到全國都過了 約旦河 。
JOSH|4|1|當全國都過了 約旦河 ，耶和華對 約書亞 說：
JOSH|4|2|「你要從百姓中選出十二個人，每支派一人，
JOSH|4|3|吩咐他們說：『你們從這裏，從 約旦河 中祭司的腳穩穩站立的地方，取十二塊石頭 ，一起帶過去，放在你們今夜住宿的地方。』」
JOSH|4|4|於是 約書亞 召集了他從 以色列 人中所選的十二個人，每支派一人。
JOSH|4|5|約書亞 對他們說：「你們要過去，到 約旦河 中，耶和華－你們上帝的約櫃前面，按 以色列 人支派的數目，每人各取一塊石頭扛在肩上。
JOSH|4|6|這些石頭在你們中間將成為記號。日後，你們的子孫問你們說：『這些石頭對你們有甚麼意思呢？』
JOSH|4|7|你們就對他們說：『這是因為 約旦河 的水在耶和華的約櫃前中斷；約櫃過 約旦河 的時候， 約旦河 的水就中斷了。這些石頭要作 以色列 人永遠的紀念。』」
JOSH|4|8|以色列 人就照 約書亞 所吩咐的做了。他們按 以色列 人支派的數目，從 約旦河 中取了十二塊石頭，正如耶和華所吩咐 約書亞 的。他們把石頭帶過去，到他們所住宿的地方，就放在那裏。
JOSH|4|9|約書亞 另外把十二塊石頭立在 約旦河 的中間，在抬約櫃祭司的腳站立的地方；直到今日，石頭還在那裏。
JOSH|4|10|抬約櫃的祭司站在 約旦河 的中間，直到耶和華命令 約書亞 告訴百姓的一切事辦完為止，正如 摩西 所吩咐 約書亞 的一切話。 於是，百姓急速過了河。
JOSH|4|11|全體百姓都過了河之後，耶和華的約櫃和祭司才過去，到百姓的前面。
JOSH|4|12|呂便 人、 迦得 人、 瑪拿西 半支派的人都照 摩西 所吩咐他們的，帶著兵器在 以色列 人的前面過去。
JOSH|4|13|約有四萬帶兵器的軍隊在耶和華面前過去，到 耶利哥 的平原，準備上陣。
JOSH|4|14|在那日，耶和華使 約書亞 在 以色列 眾人眼前被尊為大。在他一生的年日中，百姓敬服他，像從前敬服 摩西 一樣。
JOSH|4|15|耶和華對 約書亞 說：
JOSH|4|16|「你吩咐抬法櫃的祭司從 約旦河 上來。」
JOSH|4|17|約書亞 就吩咐祭司說：「你們從 約旦河 上來。」
JOSH|4|18|抬耶和華約櫃的祭司從 約旦河 中上來，腳掌一落乾地， 約旦河 的水就流回原處，仍舊漲滿兩岸。
JOSH|4|19|正月初十，百姓從 約旦河 上來，就在 耶利哥 東邊的 吉甲 安營。
JOSH|4|20|約書亞 把他們從 約旦河 取來的那十二塊石頭立在 吉甲 ，
JOSH|4|21|對 以色列 人說：「日後，你們的子孫問他們的父親說：『這些石頭是甚麼意思呢？』
JOSH|4|22|你們就讓你們的子孫知道，說：『 以色列 人曾走乾地過這 約旦河 。』
JOSH|4|23|因為耶和華－你們的上帝在你們前面使 約旦河 的水乾了，直到你們過來，就如耶和華－你們的上帝從前在我們前面使 紅海 乾了，直到我們過來一樣，
JOSH|4|24|要使地上萬民都知道，耶和華的手大有能力，也要使你們天天敬畏耶和華－你們的上帝。」
JOSH|5|1|約旦河 西 亞摩利 人的眾王和靠海 迦南 人的眾王，聽見耶和華在 以色列 人前面使 約旦河 的水乾了，直到他們過了河 ，眾王因 以色列 人的緣故都膽戰心驚，勇氣全失。
JOSH|5|2|那時，耶和華對 約書亞 說：「你要造火石刀，第二次為 以色列 人行割禮。」
JOSH|5|3|約書亞 就造了火石刀，在 哈爾拉勒山 為 以色列 人行割禮。
JOSH|5|4|約書亞 行割禮的原因是這樣：從 埃及 出來的眾百姓，所有能打仗的男丁，出了 埃及 以後，都死在曠野的路上。
JOSH|5|5|這些從 埃及 出來的眾百姓都受過割禮；但是那些出 埃及 以後，在曠野的路上所生的眾百姓卻沒有受過割禮。
JOSH|5|6|以色列 人在曠野走了四十年，直到那從 埃及 出來，全國能打仗的人都消滅了，因為他們沒有聽從耶和華的話。耶和華曾向他們起誓，必不容許他們看見耶和華向他們列祖起誓要給我們的地，就是流奶與蜜之地。
JOSH|5|7|他們的子孫，就是耶和華興起接續他們的，都沒有受過割禮；因為在路上他們沒有受割禮， 約書亞 就為他們行割禮。
JOSH|5|8|全國的人都受了割禮，留在營中自己的地方，直到痊癒。
JOSH|5|9|耶和華對 約書亞 說：「我今日將 埃及 的羞辱從你們身上除掉了。」因此，那地方名叫 吉甲 ，直到今日。
JOSH|5|10|以色列 人在 吉甲 安營。正月十四日晚上，他們在 耶利哥 的平原守逾越節。
JOSH|5|11|逾越節的第二日，他們吃了當地的出產，就在那一天，吃了無酵餅和烘過的穀物。
JOSH|5|12|他們吃了當地出產的第二日，嗎哪就停止了。 以色列 人不再有嗎哪了。那一年，他們就吃 迦南 地的出產。
JOSH|5|13|約書亞 靠近 耶利哥 的時候，舉目觀看，看哪，有一個人站在他對面，手裏拿著拔出來的刀。 約書亞 到他那裏，對他說：「你是屬我們的，還是屬我們敵人的呢？」
JOSH|5|14|他說：「不，我現在來是要作耶和華軍隊的元帥。」 約書亞 就臉伏於地下拜，說：「我主有甚麼話，請吩咐僕人吧！」
JOSH|5|15|耶和華軍隊的元帥對 約書亞 說：「把你腳上的鞋脫下來，因為你所站的地方是聖的。」 約書亞 就照著做了。
JOSH|6|1|耶利哥 的城門因 以色列 人的緣故，關得嚴緊，無人出入。
JOSH|6|2|耶和華對 約書亞 說：「看，我已經把 耶利哥城 和 耶利哥 王，以及大能的勇士，都交在你手中。
JOSH|6|3|你們要圍繞這城，所有的士兵繞城一次，六日你都要這樣做。
JOSH|6|4|七個祭司要拿七個羊角走在約櫃前。到了第七日，你們要圍繞這城七次，祭司也要吹角。
JOSH|6|5|羊角聲拖長的時候，你們一聽見角聲，眾百姓要大聲呼喊，城牆就必倒塌，各人要往前直上。」
JOSH|6|6|嫩 的兒子 約書亞 召了祭司來，對他們說：「你們抬起約櫃來，要有七個祭司拿七個羊角在耶和華的約櫃前。」
JOSH|6|7|他又對百姓說：「你們向前去圍繞那城，帶兵器的要在耶和華的約櫃前過去。」
JOSH|6|8|按照 約書亞 對百姓所說的，七個祭司拿了七個羊角在耶和華面前過去，他們吹著角，耶和華的約櫃在他們後面跟著。
JOSH|6|9|帶兵器的走在吹角的祭司前面，後隊跟著約櫃走，號角繼續在吹。
JOSH|6|10|約書亞 吩咐百姓說：「你們不可呼喊，不可讓人聽見你們的聲音，連一句話也不可出你們的口，直到我對你們說『呼喊』的那日，你們才呼喊。」
JOSH|6|11|這樣， 約書亞 使耶和華的約櫃圍繞那城，把城繞了一次。然後，眾人回到營裏，就在營裏住宿。
JOSH|6|12|約書亞 清早起來，祭司又抬起耶和華的約櫃。
JOSH|6|13|七個祭司拿七個羊角，走在耶和華的約櫃前，他們吹著角；帶兵器的走在他們前面，後隊跟著耶和華的約櫃走，號角繼續在吹。
JOSH|6|14|第二日，他們再把城圍繞一次，就回營裏去。六日都是這樣做。
JOSH|6|15|第七日清早黎明時，他們起來，以同樣的方式圍繞城七次；惟獨這一日他們圍繞城七次。
JOSH|6|16|到了第七次，祭司吹角的時候， 約書亞 對百姓說：「呼喊吧，因為耶和華已經把城交給你們了！
JOSH|6|17|這城和其中所有的都要永獻給耶和華作當毀滅的，只有妓女 喇合 與她家中所有的可以存活，因為她隱藏了我們所派的使者。
JOSH|6|18|但你們務必謹慎，不可取那當滅的物，免得你們受詛咒，取了那當滅的物，使 以色列 全營成為詛咒而遭受災禍。
JOSH|6|19|只有金子、銀子和銅鐵的器皿都要歸耶和華為聖，放入耶和華的庫房中。」
JOSH|6|20|於是百姓呼喊，祭司吹角。百姓一聽見角聲就大聲呼喊，城牆隨著倒塌。百姓上去進城，各人往前直上，把城奪取。
JOSH|6|21|他們把城中所有的，無論男女老少，牛羊和驢，都用刀殺盡。
JOSH|6|22|約書亞 對窺探這地的兩個人說：「你們進那妓女的家，照你們向她所起的誓，將那女人和她所有的都從那裏帶出來。」
JOSH|6|23|兩個作過探子的青年進去，把 喇合 與她的父母、兄弟，和她所有的帶出來，他們把她所有的親屬都帶出來，安置在 以色列 的營外。
JOSH|6|24|他們用火焚燒了那城和其中所有的，只有金子、銀子和銅鐵的器皿都放在耶和華殿的庫房中。
JOSH|6|25|至於妓女 喇合 和她父家，以及她所有的， 約書亞 保存了他們的性命。她就住在 以色列 中，直到今日，因為她隱藏了 約書亞 派來窺探 耶利哥 的使者。
JOSH|6|26|當時， 約書亞 叫眾人起誓說：「凡興起重修這 耶利哥城 的，當在耶和華面前受詛咒。 他立根基的時候，必喪長子， 安城門的時候，必喪幼子。」
JOSH|6|27|耶和華與 約書亞 同在， 約書亞 的名聲傳遍全地。
JOSH|7|1|以色列 人在當滅之物上犯了罪。 猶大 支派中， 謝拉 的曾孫， 撒底 的孫子， 迦米 的兒子 亞干 取了當滅之物，耶和華的怒氣就向 以色列 人發作。
JOSH|7|2|約書亞 從 耶利哥 派人往 伯特利 東邊，靠近 伯‧亞文 的 艾城 去，對他們說：「你們上去窺探那地。」那些人就上去窺探 艾城 。
JOSH|7|3|他們回到 約書亞 那裏，對他說：「眾百姓不必都上去，只要二、三千人上去就能攻取 艾城 ；不必勞動眾百姓都上去，因為他們人少。」
JOSH|7|4|於是百姓中約有三千人上那裏去，但他們竟在 艾城 的人面前逃跑。
JOSH|7|5|艾城 的人擊殺他們約三十六人，從城門前追趕他們，直到 示巴琳 ，在下坡的地方擊敗他們。他們都膽戰心驚，融化如水。
JOSH|7|6|約書亞 和 以色列 的長老就撕裂衣服，在耶和華的約櫃前臉伏於地，直到晚上。他們把灰撒在頭上。
JOSH|7|7|約書亞 說：「唉！主耶和華啊，你為甚麼領這百姓過 約旦河 ，把我們交在 亞摩利 人手中，使我們滅亡呢？我們不如住在 約旦河 的那邊！
JOSH|7|8|主啊，求求你， 以色列 人既在仇敵面前轉身逃跑，我還有甚麼可說的呢？
JOSH|7|9|迦南 人和這地所有的居民聽見了就必圍困我們，把我們的名從地上除去。那時，你為你至大的名要怎樣做呢？」
JOSH|7|10|耶和華對 約書亞 說：「起來！你的臉為何這樣俯伏呢？
JOSH|7|11|以色列 犯了罪，又違背了我所吩咐他們的約，又取了當滅之物。他們又偷竊，又行詭詐，又把那當滅的物與自己的器皿放在一起。
JOSH|7|12|因此， 以色列 人在仇敵面前站立不住。他們在仇敵面前轉身逃跑，因為他們成了當滅的物。你們若不把當滅的物從你們中間除掉，我就不再與你們同在了。
JOSH|7|13|你起來，去叫百姓分別為聖，說：『你們要為了明天使自己分別為聖，因為耶和華－ 以色列 的上帝這樣說： 以色列 啊，在你中間有當滅的物；你們若不把你們中間當滅之物除掉，你在仇敵面前必站立不住！』
JOSH|7|14|到了早晨，你們要按著支派近前來。耶和華所選的支派，要按著宗族近前來；耶和華所選的宗族，要按著家族近前來；耶和華所選的家族，要按著男丁，一個一個近前來。
JOSH|7|15|被選的人有當滅之物在他那裏，他和他所有的必被火焚燒，因為他違背了耶和華的約，又因他在 以色列 中做了愚妄的事。」
JOSH|7|16|於是， 約書亞 清早起來，召 以色列 按著支派近前來。選出來的是 猶大 支派。
JOSH|7|17|他召 猶大 的宗族近前來，選出來的是 謝拉 宗族。他召 謝拉 宗族，按著男丁 ，一個一個近前來，選出來的是 撒底 。
JOSH|7|18|他召 撒底 的家族，按著男丁，一個一個近前來，就選出 猶大 支派， 謝拉 的曾孫， 撒底 的孫子， 迦米 的兒子 亞干 。
JOSH|7|19|約書亞 對 亞干 說：「我兒，我勸你將榮耀歸給耶和華－ 以色列 的上帝，在他面前認罪，把你所做的事告訴我，不可向我隱瞞。」
JOSH|7|20|亞干 回答 約書亞 說：「我實在得罪了耶和華－ 以色列 的上帝。這是我所做的：
JOSH|7|21|我在所奪取的財物中看見一件美好的 示拿 外袍，二百舍客勒銀子，一條重五十舍客勒的金子。我貪愛這些物件，就拿去了。看哪，這些東西都埋在我帳棚內的地裏，銀子在外袍底下。」
JOSH|7|22|約書亞 就派使者跑到 亞干 的帳棚裏。看哪，那件外袍藏在他的帳棚裏，銀子在外袍底下。
JOSH|7|23|他們從帳棚裏把這些東西取出來，拿到 約書亞 和 以色列 眾人 那裏，倒在耶和華面前。
JOSH|7|24|約書亞 和 以色列 眾人把 謝拉 的曾孫 亞干 和那銀子、那件外袍、那條金子，以及 亞干 的兒女、牛、驢、羊、帳棚，和他所有的，都帶著上到 亞割谷 去。
JOSH|7|25|約書亞 說：「你為甚麼給我們招惹災禍呢？今日耶和華必使你遭受災禍。」於是 以色列 眾人用石頭打死他，用火焚燒他們，把石頭扔在其上。
JOSH|7|26|眾人在 亞干 身上堆了一大堆石頭，直存到今日。於是耶和華轉意，不發他的烈怒。因此，那地方名叫 亞割谷 ，直到今日。
JOSH|8|1|耶和華對 約書亞 說：「不要懼怕，也不要驚惶。你起來，率領所有作戰的士兵上 艾城 去。看，我已經把 艾城 的王和他的百姓、他的城，以及他的地，都交在你手裏。
JOSH|8|2|你怎樣處置 耶利哥 和 耶利哥 的王，也當照樣處置 艾城 和 艾城 的王。只是城內所奪的財物和牲畜，你們可以取為自己的掠物。你要在城的後面設下伏兵。
JOSH|8|3|於是， 約書亞 和所有作戰的士兵都起來，上 艾城 去。 約書亞 選了三萬大能的勇士，夜間派遣他們前去，
JOSH|8|4|吩咐他們說：「看，你們要在城的後面埋伏，不可離城太遠，各人都要準備。
JOSH|8|5|我與我所帶領的眾士兵要向城前進。城裏的人像上一次那樣出來迎擊我們的時候，我們就在他們面前逃跑。
JOSH|8|6|他們會出來追趕我們，直到我們引誘他們遠離那城。因為他們必說：『這些人像上次那樣在我們面前逃跑。』所以我們要在他們面前逃跑 。
JOSH|8|7|那時，你們就從埋伏的地方起來，奪取那城，因為耶和華－你們的上帝必把城交在你們的手裏。
JOSH|8|8|你們奪了城以後，要放火燒城，照耶和華的話去做。看，這是我吩咐你們的。」
JOSH|8|9|於是， 約書亞 派遣他們前去。他們行軍到埋伏的地方，伏在 伯特利 和 艾城 的中間，就是 艾城 的西邊。這夜， 約書亞 在士兵中間過夜。
JOSH|8|10|約書亞 清早起來，點齊士兵。他和 以色列 的長老在百姓前面上 艾城 去。
JOSH|8|11|所有跟他一起作戰的士兵都上去，向前逼近，來到城前，就在 艾城 北邊安營。 約書亞 與 艾城 之間隔著一個山谷。
JOSH|8|12|他選了約五千人，安排他們埋伏在 伯特利 和 艾城 的中間，就是 艾城 的西邊。
JOSH|8|13|於是，他們佈署軍隊，就是城北的全軍和城西的伏兵。當夜 約書亞 進入山谷之中。
JOSH|8|14|艾城 的王看見了，就和城裏的人清早起來，急忙出去，他和所有的士兵到了所定的地點，在 亞拉巴 前，迎擊 以色列 ，與之交戰；王並不知道城的後面有伏兵。
JOSH|8|15|約書亞 和 以色列 眾人在他們面前裝敗，往曠野的路逃跑。
JOSH|8|16|城內所有的百姓都被召來追趕他們。 艾城 的人追趕 約書亞 的時候，就被引誘遠離了城。
JOSH|8|17|艾城 和 伯特利 沒有一人不出來追趕 以色列 人的。他們撇下敞開的城門，去追趕 以色列 人。
JOSH|8|18|耶和華對 約書亞 說：「你向 艾城 伸出手裏的標槍，因為我要把那城交在你手裏。」 約書亞 就向那城伸出手裏的標槍。
JOSH|8|19|他一伸手，伏兵立刻從埋伏的地方衝出來，直攻入城，奪了它，立刻放火燒城。
JOSH|8|20|艾城 的人回頭，往後一看，看哪，城中煙氣沖天，他們向這邊或那邊都無處可逃。往曠野逃跑的百姓就轉身攻擊那些追趕他們的人。
JOSH|8|21|約書亞 和 以色列 眾人見伏兵已經奪了城，城中煙氣上騰，就轉身擊殺 艾城 的人。
JOSH|8|22|伏兵也出城追擊他們，他們就被 以色列 人前後夾攻，四面受敵。於是 以色列 人擊殺他們，沒有留下一個倖存者，也沒有一個逃脫。
JOSH|8|23|以色列 人生擒了 艾城 的王，把他解到 約書亞 那裏。
JOSH|8|24|以色列 人在田間和曠野殺盡了追趕他們的 艾城 所有的居民。他們全倒在刀下，直到滅盡。 以色列 眾人就回到 艾城 ，用刀殺了城中的人。
JOSH|8|25|當日殺死的人，連男帶女共有一萬二千，這也是 艾城 所有的人。
JOSH|8|26|約書亞 沒有收回手裏所伸出來的標槍，直到他滅絕 艾城 所有的居民。
JOSH|8|27|只是牲畜和城內所奪的財物， 以色列 人都照耶和華所吩咐 約書亞 的話，取為自己的掠物。
JOSH|8|28|約書亞 焚燒 艾城 ，使城成為永遠的廢墟，直到今日還是荒涼。
JOSH|8|29|他把 艾城 的王掛在樹上，直到晚上。日落的時候， 約書亞 吩咐人把屍首從樹上取下來，丟在城門口，並在屍首上堆了一大堆石頭，直存到今日。
JOSH|8|30|那時， 約書亞 在 以巴路山 上為耶和華－ 以色列 的上帝築一座壇。
JOSH|8|31|這壇是照耶和華的僕人 摩西 吩咐 以色列 人，用沒有動過鐵器的整塊石頭所築的，正如 摩西 律法書上所寫的。他們在這壇上給耶和華奉獻燔祭，又宰牲作為平安祭。
JOSH|8|32|約書亞 在那裏，當著 以色列 人面前，將 摩西 所寫的律法抄寫在石頭上。
JOSH|8|33|以色列 眾人，無論是本地人或寄居的，都和他們的長老、官長和審判官，站在約櫃兩旁，在抬耶和華約櫃的 利未 家的祭司面前，一半對著 基利心山 ，一半對著 以巴路山 ，照耶和華的僕人 摩西 先前所吩咐的，為 以色列 百姓祝福。
JOSH|8|34|隨後， 約書亞 將律法上祝福和詛咒的話，照著律法書上一切所寫的，宣讀一遍。
JOSH|8|35|摩西 所吩咐的一切話， 約書亞 在 以色列 全會眾和婦女、孩童，以及住在他們中間的外人面前，沒有一句不宣讀的。
JOSH|9|1|約旦河 西，住山區、低地和沿 大海 一帶直到 黎巴嫩 的諸王，就是 赫 人、 亞摩利 人、 迦南 人、 比利洗 人、 希未 人、 耶布斯 人的諸王，聽見這事，
JOSH|9|2|就都聚集，同心合意要與 約書亞 和 以色列 人作戰。
JOSH|9|3|基遍 的居民聽見 約書亞 向 耶利哥 和 艾城 所做的事，
JOSH|9|4|就設詭計，假扮使者 出去。他們拿舊布袋和破裂補過的舊皮酒袋馱在驢上，
JOSH|9|5|將補過的舊鞋穿在腳上，把舊衣服穿在身上，作食物的餅都又乾又長了霉 。
JOSH|9|6|他們到 吉甲 營中 約書亞 那裏，對他和 以色列 人說：「我們是從遠地來的，現在求你與我們立約。」
JOSH|9|7|以色列 人對 希未 人說：「或許你是住在我附近的。若是這樣，我怎能和你立約呢？」
JOSH|9|8|他們對 約書亞 說：「我們是你的僕人。」 約書亞 對他們說：「你們是甚麼人？是從哪裏來的？」
JOSH|9|9|他們對他說：「你的僕人是因耶和華－你上帝的名從極遠之地來的。我們聽見他的名聲，他在 埃及 所做的一切，
JOSH|9|10|以及他向 約旦河 東的兩個 亞摩利 王， 希實本 王 西宏 和在 亞斯她錄 的 巴珊 王 噩 所做的一切。
JOSH|9|11|我們的長老和我們當地所有的居民對我們說：『你們手裏要帶著路上用的乾糧去迎接 以色列 人，對他們說：我們是你們的僕人。現在求你們與我們立約。』
JOSH|9|12|我們出來要往你們這裏來的那日，這從我們家裏帶出來的餅是熱的；看哪，現在這餅又乾又長了霉。
JOSH|9|13|這些皮酒袋，我們盛酒的時候還是新的；看哪，現在已經破裂了。我們這些衣服和鞋，因為路途非常遙遠，也都穿舊了。」
JOSH|9|14|以色列 人收下他們的一些食物，但是沒有求問耶和華的指示。
JOSH|9|15|於是 約書亞 與他們建立和好關係，與他們立約，讓他們存活；會眾的領袖也向他們起誓。
JOSH|9|16|以色列 人與他們立約之後，過了三天才聽說他們是近鄰，住在附近。
JOSH|9|17|以色列 人起行，第三天就到了他們的城鎮，他們的城鎮是 基遍 、 基非拉 、 比錄 和 基列‧耶琳 。
JOSH|9|18|因為會眾的領袖已經指著耶和華－ 以色列 的上帝向他們起誓，所以 以色列 人不擊殺他們。全會眾就向領袖發怨言。
JOSH|9|19|眾領袖對全會眾說：「我們已經指著耶和華－ 以色列 的上帝向他們起誓，現在我們不能碰他們。
JOSH|9|20|我們要這樣對待他們，讓他們存活，免得因我們向他們所起的誓而憤怒臨到我們。」
JOSH|9|21|領袖對會眾說：「讓他們活著吧。」於是他們照領袖所說的，為全會眾作劈柴挑水的人。
JOSH|9|22|約書亞 召了他們來，對他們說：「你們為甚麼欺騙我們說：『我們離你們很遠』呢？其實你們就住在我們附近。
JOSH|9|23|現在你們當受詛咒！你們中間必不斷有人作奴僕，為我上帝的殿作劈柴挑水的人。」
JOSH|9|24|他們回答 約書亞 說：「因為確實有人告訴你的僕人，耶和華－你的上帝曾吩咐他的僕人 摩西 ，把這全地賜給你們，並要在你們面前除滅這地所有的居民。我們因你們的緣故很怕自己喪命，就做了這事。
JOSH|9|25|現在，看哪，我們在你手中，你看怎樣待我們是好的，是對的，就這樣做吧！」
JOSH|9|26|於是 約書亞 就這樣對待他們，他救了他們脫離 以色列 人的手， 以色列 人沒有殺他們。
JOSH|9|27|那日， 約書亞 分派他們到耶和華選擇的地方，為會眾和耶和華的壇劈柴挑水，直到今日。
JOSH|10|1|耶路撒冷 王 亞多尼‧洗德 聽見 約書亞 奪了 艾城 ，徹底毀滅，處置 艾城 和 艾城 的王像處置 耶利哥 和 耶利哥 的王一樣，又聽見 基遍 的居民與 以色列 人立了和約，住在他們中間，
JOSH|10|2|耶路撒冷 人就很懼怕，因為 基遍 是一座大城，如京城一樣，比 艾城 更大，並且城內的人都是勇士。
JOSH|10|3|耶路撒冷 王 亞多尼‧洗德 派人去見 希伯崙 王 何咸 、 耶末 王 毗蘭 、 拉吉 王 雅非亞 和 伊磯倫 王 底璧 ，說：
JOSH|10|4|「求你們上來幫助我，我們好攻打 基遍 ，因為它與 約書亞 和 以色列 人立了和約。」
JOSH|10|5|於是五個 亞摩利 王，就是 耶路撒冷 王、 希伯崙 王、 耶末 王、 拉吉 王和 伊磯倫 王，聯合上去，率領他們所有的軍隊，對著 基遍 安營，要攻打 基遍 。
JOSH|10|6|基遍 人就派人到 吉甲 的營中 約書亞 那裏，說：「不要袖手不顧你的僕人，求你趕快上來拯救我們，幫助我們，因為住山區 亞摩利 人的諸王已經聯合來攻擊我們。」
JOSH|10|7|於是 約書亞 和所有跟他一起作戰的士兵，以及大能的勇士，從 吉甲 上去。
JOSH|10|8|耶和華對 約書亞 說：「不要怕他們， 因為我已將他們交在你手裏，他們沒有一人能在你面前站立得住。」
JOSH|10|9|約書亞 就連夜從 吉甲 上去，猛然襲擊他們。
JOSH|10|10|耶和華使他們在 以色列 人面前潰亂。 約書亞 在 基遍 大大擊殺他們，在 伯‧和崙 的上坡路上追趕他們，擊殺他們，直到 亞西加 和 瑪基大 。
JOSH|10|11|他們在 以色列 人面前逃跑。正在 伯‧和崙 下坡的時候，耶和華從天上降下大冰雹 在他們身上，直降到 亞西加 ，打死他們。被冰雹打死的，比 以色列 人用刀殺死的還多。
JOSH|10|12|當耶和華將 亞摩利 人交給 以色列 人的那一日， 約書亞 向耶和華說話，在 以色列 人眼前說： 「太陽啊，停在 基遍 ； 月亮啊，停在 亞雅崙谷 。」
JOSH|10|13|太陽就停住，月亮就止住， 直到國民向敵人報仇。 這事豈不是寫在《雅煞珥書》上嗎？太陽停在天空當中，沒有急速下落，約有一整天。
JOSH|10|14|在這日以前，這日以後，耶和華聽人的聲音，沒有像這日的，這是因為耶和華為 以色列 作戰。
JOSH|10|15|約書亞 和跟他一起的 以色列 眾人回到 吉甲 的營中。
JOSH|10|16|那五個王逃跑，躲在 瑪基大 洞裏。
JOSH|10|17|有人告訴 約書亞 說：「那五個王已經找到了，都躲在 瑪基大 洞裏。」
JOSH|10|18|約書亞 說：「你們把幾塊大石頭滾到洞口，派人在那裏看守他們。
JOSH|10|19|你們卻不可停留，要追趕你們的仇敵，從後面攻擊他們，不讓他們進到自己的城鎮，因為耶和華－你們的上帝已經把他們交在你們手裏。」
JOSH|10|20|約書亞 和 以色列 人徹底擊敗他們，直到把他們滅盡，只剩下少許的人逃進堅固的城。
JOSH|10|21|眾百姓就安然回到 瑪基大 營中 ，到 約書亞 那裏。沒有人敢向 以色列 人饒舌。
JOSH|10|22|約書亞 說：「打開洞口，把那五個王從洞裏帶出來，到我這裏。」
JOSH|10|23|眾人就這樣做，把那五個王，就是 耶路撒冷 王、 希伯崙 王、 耶末 王、 拉吉 王和 伊磯倫 王，從洞裏帶出來，到 約書亞 那裏。
JOSH|10|24|他們帶出那五個王到 約書亞 那裏的時候， 約書亞 就召了 以色列 眾人來，對和他同去的軍官說：「你們近前來，把腳踏在這些王的頸項上。」他們就近前來，把腳踏在這些王的頸項上。
JOSH|10|25|約書亞 對他們說：「你們不要懼怕，也不要驚惶。當剛強壯膽，因為耶和華必這樣處置你們要攻打的所有仇敵。」
JOSH|10|26|隨後， 約書亞 把這五個王殺死，掛在五棵樹上。他們就被掛在樹上，直到晚上。
JOSH|10|27|日落的時候， 約書亞 吩咐人把屍首從樹上取下來，丟在他們躲過的洞裏，把幾塊大石頭放在洞口，直存到今日。
JOSH|10|28|當日， 約書亞 奪了 瑪基大 ，用刀擊殺城中的人和王，把城中所有人完全滅盡，沒有留下一個倖存者。他處置 瑪基大 王，像從前處置 耶利哥 王一樣。
JOSH|10|29|約書亞 和跟他一起的 以色列 眾人從 瑪基大 往 立拿 去，攻打 立拿 。
JOSH|10|30|耶和華將 立拿 和 立拿 的王也交在 以色列 人手裏。 約書亞 攻打這城，用刀擊殺了城中所有的人，沒有留下一個倖存者。他處置 立拿 王，像從前處置 耶利哥 王一樣。
JOSH|10|31|約書亞 和跟他一起的 以色列 眾人從 立拿 往 拉吉 去，對著 拉吉 安營，攻打這城。
JOSH|10|32|耶和華將 拉吉 交在 以色列 人的手裏。第二日 約書亞 就奪了 拉吉 ，用刀擊殺了城中所有的人，正如他向 立拿 一切所做的。
JOSH|10|33|那時 基色 王 何蘭 上來幫助 拉吉 ， 約書亞 就把他和他的百姓都擊殺了，沒有留下一個倖存者。
JOSH|10|34|約書亞 和跟他一起的 以色列 眾人從 拉吉 往 伊磯倫 去，對著 伊磯倫 安營，攻打這城。
JOSH|10|35|當日 約書亞 就奪了城，用刀擊殺了城中的人。那日， 約書亞 把城中所有的人完全滅盡，正如他向 拉吉 一切所做的。
JOSH|10|36|約書亞 和跟他一起的 以色列 眾人從 伊磯倫 上 希伯崙 去，攻打這城，
JOSH|10|37|奪了 希伯崙 ，用刀擊敗 希伯崙 、它的王和屬它的一切城鎮，以及城中所有的人；他沒有留下一個倖存者，正如他向 伊磯倫 所做的，把城中所有的人完全滅盡。
JOSH|10|38|約書亞 和跟他一起的 以色列 眾人回到 底璧 ，攻打這城，
JOSH|10|39|奪了 底璧 和屬它的一切城鎮，又擒獲它的王，用刀把城中所有的人完全滅盡，沒有留下一個倖存者。他處置 底璧 和它的王，像從前處置 希伯崙 ，處置 立拿 和它的王一樣。
JOSH|10|40|這樣， 約書亞 擊敗全地的人，就是山區、 尼革夫 、低地、山坡的人，和那裏的眾王，沒有留下一個倖存者。他把凡有氣息的完全滅盡，正如耶和華－ 以色列 的上帝所吩咐的。
JOSH|10|41|約書亞 從 加低斯‧巴尼亞 攻到 迦薩 ，又攻打 歌珊 全地，直到 基遍 。
JOSH|10|42|約書亞 一舉擊敗了這些王，奪了他們的地，因為耶和華－ 以色列 的上帝為 以色列 作戰。
JOSH|10|43|於是 約書亞 和跟他一起的 以色列 眾人回到 吉甲 的營中。
JOSH|11|1|夏瑣 王 耶賓 聽見了，就派人到 瑪頓 王 約巴 、 伸崙 王、 押煞 王，
JOSH|11|2|和北方山區、 基尼烈 南邊的 亞拉巴 、低地、西邊 多珥 山岡 的諸王，
JOSH|11|3|以及東方和西方的 迦南 人、山區的 亞摩利 人、 赫 人、 比利洗 人、 耶布斯 人，和 黑門山 下 米斯巴 地的 希未 人那裏。
JOSH|11|4|他們和他們的眾軍都出來，一大隊人馬，多如海邊的沙，並有極多的戰車戰馬。
JOSH|11|5|眾王組成聯軍，來到 米倫 水邊一同安營，要與 以色列 作戰。
JOSH|11|6|耶和華對 約書亞 說：「你不要怕他們。明日這時，我必把他們全部交給 以色列 人殺滅。你要砍斷他們馬的蹄筋，用火焚燒他們的戰車。」
JOSH|11|7|於是 約書亞 和所有跟他一起作戰的士兵，來到 米倫 水邊，突然攻擊他們。
JOSH|11|8|耶和華將他們交在 以色列 人手裏， 以色列 人就擊殺他們，追趕他們到 西頓 大城，到 米斯利弗‧瑪音 ，直到東邊 米斯巴 的山谷。 以色列 人擊殺他們，沒有留下一個倖存者。
JOSH|11|9|約書亞 照耶和華所吩咐他的去做，砍斷他們馬的蹄筋，用火焚燒他們的戰車。
JOSH|11|10|那時， 約書亞 轉回，奪了 夏瑣 ，用刀殺了 夏瑣 王。先前 夏瑣 在這些王國中是為首的。
JOSH|11|11|以色列 人用刀擊殺城中所有的人，把他們完全滅盡；凡有氣息的，沒有留下一個。 約書亞 又用火焚燒 夏瑣 。
JOSH|11|12|約書亞 奪了這些王的一切城鎮，擒獲了這些王，用刀殺了他們，把他們完全滅盡，正如耶和華的僕人 摩西 所吩咐的。
JOSH|11|13|至於造在山岡上的城鎮，除了 夏瑣 以外， 以色列 人都沒有焚燒。 約書亞 只焚燒了 夏瑣 。
JOSH|11|14|從那些城鎮所奪的財物和牲畜， 以色列 人都取為自己的掠物。至於所有的人，他們都用刀殺了，直到滅盡；凡有氣息的，沒有留下一個。
JOSH|11|15|耶和華怎樣吩咐他的僕人 摩西 ， 摩西 就這樣吩咐 約書亞 ， 約書亞 也照樣做了。凡耶和華所吩咐 摩西 的， 約書亞 沒有一件偏離不做的。
JOSH|11|16|約書亞 奪了那全地，就是山區、整個 尼革夫 、 歌珊 全地、低地、 亞拉巴 、 以色列 的山區和山下的低地，
JOSH|11|17|從上 西珥 的 哈拉山 ，直到 黑門山 下面 黎巴嫩 平原的 巴力‧迦得 。他擒獲了那裏的眾王，把他們殺死。
JOSH|11|18|約書亞 和這些王作戰了很長的一段日子。
JOSH|11|19|除了 希未 人 基遍 的居民之外，沒有一城與 以色列 人講和，都是 以色列 人作戰奪來的。
JOSH|11|20|因為耶和華的意思是要使他們的心剛硬，來與 以色列 人作戰，好使他們全被殺滅，不蒙憐憫，反被除滅，正如耶和華所吩咐 摩西 的。
JOSH|11|21|那時 約書亞 來到，剪除了住山區、 希伯崙 、 底璧 、 亞拿伯 、整個 猶大 山區和 以色列 山區的 亞衲 族人。 約書亞 把他們和他們的城鎮盡都毀滅。
JOSH|11|22|以色列 人的地中沒有留下一個 亞衲 族人，只有一些還留在 迦薩 、 迦特 和 亞實突 。
JOSH|11|23|這樣， 約書亞 照著耶和華所吩咐 摩西 的一切話奪了那全地，就按著 以色列 支派所得的份把地分給他們為業。於是國中太平，沒有戰爭了。
JOSH|12|1|這些是 以色列 人在 約旦河 東，向日出的方向，從 亞嫩谷 直到 黑門山 ，以及東邊 亞拉巴 的整個地區所擊殺的王和所得的地：
JOSH|12|2|有住 希實本 的 亞摩利 王 西宏 ，他統治的地從 亞嫩谷 邊的 亞羅珥 起，包括谷中之城和 基列 的一半，直到 亞捫 人邊界的 雅博河 ，
JOSH|12|3|以及從東邊的 亞拉巴 ，直到 基尼烈海 ，又向東通過 伯‧耶施末 的路，直到 亞拉巴 的海，就是 鹽海 ，再往南直到 毗斯迦山 斜坡的山腳。
JOSH|12|4|又有 巴珊 王 噩 ，他是 利乏音 人所剩下的，住在 亞斯她錄 和 以得來 。
JOSH|12|5|他統治的地是 黑門山 、 撒迦 、 巴珊 全地，直到 基述 人和 瑪迦 人的邊界，以及 基列 的一半，直到 希實本 王 西宏 的邊界。
JOSH|12|6|這兩個王是耶和華的僕人 摩西 和 以色列 人所擊殺的。耶和華的僕人 摩西 把他們的地賜給 呂便 人、 迦得 人和 瑪拿西 半支派的人為業。
JOSH|12|7|這些是 約書亞 和 以色列 人在 約旦河 西所擊殺的諸王，他們的地從 黎巴嫩 平原的 巴力‧迦得 ，直上到 西珥 的 哈拉山 。 約書亞 按著 以色列 支派所得的份把這地分給他們為業，
JOSH|12|8|就是 赫 人、 亞摩利 人、 迦南 人、 比利洗 人、 希未 人、 耶布斯 人的地，包括山區、低地、 亞拉巴 、山坡、曠野和 尼革夫 。
JOSH|12|9|這些王是： 耶利哥 王一人， 靠近 伯特利 的 艾城 王一人，
JOSH|12|10|耶路撒冷 王一人， 希伯崙 王一人，
JOSH|12|11|耶末 王一人， 拉吉 王一人，
JOSH|12|12|伊磯倫 王一人， 基色 王一人，
JOSH|12|13|底璧 王一人， 基德 王一人，
JOSH|12|14|何珥瑪 王一人， 亞拉得 王一人，
JOSH|12|15|立拿 王一人， 亞杜蘭 王一人，
JOSH|12|16|瑪基大 王一人， 伯特利 王一人，
JOSH|12|17|他普亞 王一人， 希弗 王一人，
JOSH|12|18|亞弗 王一人， 拉沙崙 王一人，
JOSH|12|19|瑪頓 王一人， 夏瑣 王一人，
JOSH|12|20|伸崙‧米崙 王一人 ， 押煞 王一人，
JOSH|12|21|他納 王一人， 米吉多 王一人，
JOSH|12|22|基低斯 王一人， 靠近 迦密 的 約念 王一人，
JOSH|12|23|多珥 山岡 的 多珥 王一人， 吉甲 的 戈印 王一人，
JOSH|12|24|得撒 王一人， 共三十一個王。
JOSH|13|1|約書亞 年紀老邁，耶和華對他說：「你年紀老邁了，還有極多剩下的未得之地。
JOSH|13|2|這是剩下的地： 非利士 人的全境和一切屬於 基述 人的，
JOSH|13|3|是從 埃及 東邊的 西曷河 往北，直到 以革倫 的邊界，算是屬 迦南 人的地，那裏有 非利士 人五個領袖統治 迦薩 人、 亞實突 人、 亞實基倫 人、 迦特 人、 以革倫 人；還有屬於 亞衛 人的，
JOSH|13|4|在南邊；還有 迦南 人的全地，以及 西頓 人的 米亞拉 到 亞弗 ，直到 亞摩利 人的邊界；
JOSH|13|5|還有 迦巴勒 人的地，以及向日出方向的 黎巴嫩 全地，從 黑門山 下的 巴力‧迦得 ，直到 哈馬口 ；
JOSH|13|6|從 黎巴嫩 直到 米斯利弗‧瑪音 ，一切山區的居民，就是所有的 西頓 人，我必在 以色列 人面前趕走他們。你只管照我所吩咐的，抽籤將這地分給 以色列 人為業。
JOSH|13|7|現在你要把這地分給九個支派和 瑪拿西 半個支派為業。
JOSH|13|8|呂便 、 迦得 二支派已經和 瑪拿西 另外半個支派得了產業，就是耶和華的僕人 摩西 在 約旦河 東所賜給他們的：
JOSH|13|9|從 亞嫩谷 邊的 亞羅珥 和谷中之城， 米底巴 的整個平原，直到 底本 ；
JOSH|13|10|還有在 希實本 作王的 亞摩利 王 西宏 的諸城，直到 亞捫 人的邊界；
JOSH|13|11|還有 基列 ， 基述 人和 瑪迦 人的邊界，整個 黑門山 、整個 巴珊 ，直到 撒迦 ；
JOSH|13|12|還有在 亞斯她錄 和 以得來 作王的 巴珊 王 噩 的整個國土， 噩 是 利乏音 人惟一存留的。 摩西 擊敗了這些人，把他們趕走。
JOSH|13|13|以色列 人卻沒有趕走 基述 人和 瑪迦 人； 基述 人和 瑪迦 人仍住在 以色列 中，直到今日。
JOSH|13|14|只是 利未 支派， 摩西 沒有分產業給他們。他們的產業是獻給耶和華－ 以色列 上帝的火祭，正如耶和華對他們說的。
JOSH|13|15|摩西 按著 呂便 支派的宗族分產業給他們。
JOSH|13|16|他們的地界是 亞嫩谷 邊的 亞羅珥 和谷中之城，靠近 米底巴 的整個平原；
JOSH|13|17|還有 希實本 和屬 希實本 平原的各城， 底本 、 巴末‧巴力 、 伯‧巴力‧勉 、
JOSH|13|18|雅雜 、 基底莫 、 米法押 、
JOSH|13|19|基列亭 、 西比瑪 、谷中山岡上的 細列‧沙轄 、
JOSH|13|20|伯‧毗珥 、 毗斯迦山 斜坡、 伯‧耶施末 ；
JOSH|13|21|還有平原的各城，和 亞摩利 王 西宏 的整個國土。這 西宏 曾在 希實本 作王， 摩西 把他和 米甸 的族長 以未 、 利金 、 蘇珥 、 戶珥 、 利巴 擊殺了；他們都是屬 西宏 的領袖，曾住在這地。
JOSH|13|22|以色列 人殺了這些人時，也用刀殺了 比珥 的兒子占卜的 巴蘭 。
JOSH|13|23|呂便 人的地界就是 約旦河 和靠近 約旦河 的地。以上是 呂便 人按著宗族所得為業的城鎮和所屬的村莊。
JOSH|13|24|摩西 按著 迦得 支派的宗族分產業給他們。
JOSH|13|25|他們的地界是 雅謝 和 基列 的各城，以及 亞捫 人之地的一半，直到 拉巴 前面的 亞羅珥 ；
JOSH|13|26|還有從 希實本 到 拉抹‧米斯巴 和 比多寧 ，又從 瑪哈念 到 底璧 的邊界，
JOSH|13|27|和谷中的 伯‧亞蘭 、 伯‧寧拉 、 疏割 、 撒分 ，就是 希實本 王 西宏 國土中其餘的地，以及 約旦河 與靠近 約旦河 的地，直到 基尼烈海 的邊緣，都在 約旦河 東。
JOSH|13|28|以上是 迦得 人按著宗族所得為業的城鎮和所屬的村莊。
JOSH|13|29|摩西 分產業給 瑪拿西 半支派，這是按著 瑪拿西 半支派的宗族分的。
JOSH|13|30|他們的地界是從 瑪哈念 起，包括整個 巴珊 全地，就是 巴珊 王 噩 的整個國土，以及在 巴珊 、 睚珥 的一切城鎮，共六十個；
JOSH|13|31|還有 基列 的一半，以及 巴珊 國的王 噩 的 亞斯她錄 和 以得來 兩座城。這些地是按著宗族分給 瑪拿西 兒子 瑪吉 子孫的，就是給 瑪吉 一半子孫的。
JOSH|13|32|以上是 摩西 在 約旦河 東， 耶利哥 對面的 摩押 平原所分配的產業。
JOSH|13|33|只是 利未 支派， 摩西 沒有把產業分給他們。耶和華－ 以色列 的上帝是他們的產業，正如耶和華對他們說的。
JOSH|14|1|這是 以色列 人在 迦南 地所得的產業，就是祭司 以利亞撒 和 嫩 的兒子 約書亞 ，以及 以色列 人各支派父系的領袖所分給他們的。
JOSH|14|2|他們照耶和華藉 摩西 所吩咐的，抽籤分產業給九個半支派。
JOSH|14|3|摩西 在 約旦河 東已經分了產業給另外兩個半支派。但是，他在他們中間沒有分產業給 利未 人。
JOSH|14|4|因 約瑟 的子孫成了兩個支派，就是 瑪拿西 和 以法蓮 。雖然他們沒有分地給 利未 人，卻給 利未 人城鎮居住，以及城鎮的郊外供他們牧養牲畜，安置財物。
JOSH|14|5|耶和華怎樣吩咐 摩西 ， 以色列 人就照樣做，把地分了。
JOSH|14|6|猶大 人來到 吉甲 ， 約書亞 那裏， 基尼洗 族 耶孚尼 的兒子 迦勒 對 約書亞 說：「耶和華在 加低斯‧巴尼亞 指著我和你對神人 摩西 所說的話，你都知道。
JOSH|14|7|耶和華的僕人 摩西 從 加低斯‧巴尼亞 差派我窺探這地的時候，我剛四十歲。我把心裏的話向他報告。
JOSH|14|8|雖然同我上去的眾弟兄使百姓膽戰心驚，我仍然專心跟從耶和華－我的上帝。
JOSH|14|9|那日， 摩西 起誓說：『你腳所踏之地必要歸你和你的子孫永遠為業，因為你專心跟從耶和華－我的上帝。』
JOSH|14|10|現在，看哪，耶和華照他所說的使我活了這四十五年。當 以色列 人在曠野飄流的時候，耶和華曾對 摩西 說了這話。現在，看哪，我已經八十五歲了。
JOSH|14|11|現今我還很健壯，像 摩西 差派我去的那天一樣；無論是戰爭，是出入，我現在的力量和那時的力量一樣。
JOSH|14|12|請你將耶和華那日所說的這山區給我。那日你也曾聽說，這裏有 亞衲 族人，以及寬大堅固的城，或許耶和華會照他所說的與我同在，我就把他們趕出去。」
JOSH|14|13|於是 約書亞 為 耶孚尼 的兒子 迦勒 祝福，把 希伯崙 給他為業。
JOSH|14|14|所以 希伯崙 成了 基尼洗 族 耶孚尼 的兒子 迦勒 的產業，直到今日，因為他專心跟從耶和華－ 以色列 的上帝。
JOSH|14|15|希伯崙 從前名叫 基列‧亞巴 ； 亞巴 是 亞衲 族最尊貴的人。於是國中太平，沒有戰爭了。
JOSH|15|1|猶大 支派按著宗族抽籤所得之地是在最南端，到 以東 的邊界，往南直到 尋 的曠野。
JOSH|15|2|他們南邊的地界是從 鹽海 的頂端，就是朝南的海灣開始，
JOSH|15|3|通到 亞克拉濱 斜坡的南邊，經過 尋 ，上到 加低斯‧巴尼亞 的南邊，又經過 希斯崙 ，上到 亞達珥 ，轉到 甲加 ，
JOSH|15|4|再經過 押們 ，順著 埃及 溪谷，這地界直通到海為止。這就是你們 南邊的地界。
JOSH|15|5|東邊的地界是從 鹽海 到 約旦河 口。北邊的地界是從 約旦河 口的海灣開始，
JOSH|15|6|這地界上到 伯‧曷拉 ，經過 伯‧亞拉巴 的北邊，這地界上到 呂便 之子 波罕 的磐石。
JOSH|15|7|這地界是從 亞割谷 往北上到 底璧 ，直向 亞都冥 斜坡對面的 吉甲 ，就是河的南邊，這地界再經過 隱‧示麥 泉，直通到 隱‧羅結 。
JOSH|15|8|這地界又上到 欣嫩子谷 ， 耶布斯 斜坡的南方， 耶布斯 就是 耶路撒冷 ，這地界又上到 欣嫩谷 西邊對面的山頂，就是在 利乏音谷 的最北端。
JOSH|15|9|這地界又從山頂延伸到 尼弗多亞 水泉，通到 以弗崙山 的城鎮，這地界又延伸到 巴拉 ， 巴拉 就是 基列‧耶琳 。
JOSH|15|10|這地界又從 巴拉 往西繞到 西珥山 ，經過 耶琳山 斜坡的北邊， 耶琳 就是 基撒崙 ，從那裏又下到 伯‧示麥 ，經過 亭拿 ，
JOSH|15|11|這地界通到 以革倫 斜坡的北邊。這地界又延伸到 施基崙 ，經過 巴拉山 到 雅比聶 ，這地界直通到海為止。
JOSH|15|12|西邊的地界就是 大海 和沿海一帶之地。這是 猶大 人按著宗族所得之地四圍的邊界。
JOSH|15|13|約書亞 照耶和華所指示的，把 猶大 人中的一份土地，就是 基列‧亞巴 ，分給 耶孚尼 的兒子 迦勒 。 亞巴 是 亞衲 族的祖先， 基列‧亞巴 就是 希伯崙 。
JOSH|15|14|迦勒 從那裏趕出 亞衲 的三族，就是 亞衲 族的 示篩 人、 亞希幔 人和 撻買 人。
JOSH|15|15|他又從那裏上去，攻擊 底璧 的居民，這 底璧 從前名叫 基列‧西弗 。
JOSH|15|16|迦勒 說：「誰能攻打 基列‧西弗 ，奪取那城，我就把我女兒 押撒 嫁給他。」
JOSH|15|17|迦勒 兄弟 基納斯 的兒子 俄陀聶 奪取了那城， 迦勒 就把女兒 押撒 嫁給他。
JOSH|15|18|押撒 來的時候，催促丈夫向她父親要一塊田。 押撒 一下驢， 迦勒 就對她說：「你要甚麼？」
JOSH|15|19|她說：「求你給我福分；你既然把我安置在 尼革夫 地，求你也給我水泉。」她父親就把上泉和下泉都賜給她。
JOSH|15|20|這是 猶大 支派按著宗族所得的產業。
JOSH|15|21|猶大 支派最南端，靠近 以東 邊界的城鎮，是 甲薛 、 以得 、 雅姑珥 、
JOSH|15|22|基拿 、 底摩拿 、 亞大達 、
JOSH|15|23|基低斯 、 夏瑣 、 以提楠 、
JOSH|15|24|西弗 、 提鍊 、 比亞綠 、
JOSH|15|25|夏瑣‧哈大他 、 加略‧希斯崙 ， 加略‧希斯崙 就是 夏瑣 ，
JOSH|15|26|亞曼 、 示瑪 、 摩拉大 、
JOSH|15|27|哈薩‧迦大 、 黑實門 、 伯‧帕列 、
JOSH|15|28|哈薩‧書亞 、 別是巴 、 比斯約他 、
JOSH|15|29|巴拉 、 以因 、 以森 、
JOSH|15|30|伊勒多臘 、 基失 、 何珥瑪 、
JOSH|15|31|洗革拉 、 麥瑪拿 、 三撒拿 、
JOSH|15|32|利巴勿 、 實忻 、 亞因 、 臨門 ，共二十九座城，還有所屬的村莊。
JOSH|15|33|在低地有 以實陶 、 瑣拉 、 亞實拿 、
JOSH|15|34|撒挪亞 、 隱‧干寧 、 他普亞 、 以楠 、
JOSH|15|35|耶末 、 亞杜蘭 、 梭哥 、 亞西加 、
JOSH|15|36|沙拉音 、 亞底他音 、 基底拉 、 基底羅他音 ，共十四座城，還有所屬的村莊。
JOSH|15|37|又有 洗楠 、 哈大沙 、 麥大‧迦得 、
JOSH|15|38|底連 、 米斯巴 、 約帖 、
JOSH|15|39|拉吉 、 波斯加 、 伊磯倫 、
JOSH|15|40|迦本 、 拉幔 、 基提利 、
JOSH|15|41|基低羅 、 伯‧大袞 、 拿瑪 、 瑪基大 ，共十六座城，還有所屬的村莊。
JOSH|15|42|又有 立拿 、 以帖 、 亞珊 、
JOSH|15|43|益弗他 、 亞實拿 、 尼悉 、
JOSH|15|44|基伊拉 、 亞革悉 、 瑪利沙 ，共九座城，還有所屬的村莊。
JOSH|15|45|又有 以革倫 和所屬的鄉鎮 與村莊，
JOSH|15|46|從 以革倫 直到海，一切靠近 亞實突 之地，以及所屬的村莊、
JOSH|15|47|亞實突 和所屬的鄉鎮與村莊， 迦薩 和所屬的鄉鎮與村莊，到 埃及 溪谷，直到 大海 以及沿海一帶之地。
JOSH|15|48|在山區有 沙密 、 雅提珥 、 梭哥 、
JOSH|15|49|大拿 、 基列‧薩拿 ， 基列‧薩拿 就是 底璧 ，
JOSH|15|50|亞拿伯 、 以實提莫 、 亞念 、
JOSH|15|51|歌珊 、 何崙 、 基羅 ，共十一座城，還有所屬的村莊。
JOSH|15|52|又有 亞拉 、 度瑪 、 以珊 、
JOSH|15|53|雅農 、 伯‧他普亞 、 亞非加 、
JOSH|15|54|宏他 、 基列‧亞巴 ， 基列‧亞巴 就是 希伯崙 ， 洗珥 ，共九座城，還有所屬的村莊。
JOSH|15|55|又有 瑪雲 、 迦密 、 西弗 、 淤他 、
JOSH|15|56|耶斯列 、 約甸 、 撒挪亞 、
JOSH|15|57|該隱 、 基比亞 、 亭拿 ，共十座城，還有所屬的村莊。
JOSH|15|58|又有 哈忽 、 伯‧夙 、 基突 、
JOSH|15|59|瑪臘 、 伯‧亞諾 、 伊勒提君 ，共六座城，還有所屬的村莊。
JOSH|15|60|又有 基列‧巴力 ， 基列‧巴力 就是 基列‧耶琳 ， 拉巴 ，共兩座城，還有所屬的村莊。
JOSH|15|61|在曠野有 伯‧亞拉巴 、 密丁 、 西迦迦 、
JOSH|15|62|匿珊 、 鹽城 、 隱‧基底 ，共六座城，還有所屬的村莊。
JOSH|15|63|至於住 耶路撒冷 的 耶布斯 人， 猶大 人不能把他們趕出去。於是， 耶布斯 人與 猶大 人同住在 耶路撒冷 ，直到今日。
JOSH|16|1|約瑟 的子孫抽籤所得之地是從靠近 耶利哥 的 約旦河 起，以 耶利哥 東邊的河水為邊界，經過曠野，從 耶利哥 上去，直到 伯特利 的山區；
JOSH|16|2|從 伯特利 又到 路斯 ，經過 亞基 人的邊界，直到 亞大錄 ；
JOSH|16|3|又往西，下到 押利提 人的邊界，到 下伯‧和崙 的邊界，到 基色 ，直通到海為止。
JOSH|16|4|約瑟 的兒子 瑪拿西 、 以法蓮 得了地業。
JOSH|16|5|以法蓮 子孫的地界，按著宗族所得的如下：他們地業的東界，是從 亞大錄‧亞達 到 上伯‧和崙 ，
JOSH|16|6|這地界直通到海。在北邊，這地界是從 密米他 ，向東繞到 他納‧示羅 ，又經過 雅挪哈 的東邊，
JOSH|16|7|從 雅挪哈 下到 亞大錄 和 拿拉 ，再到 耶利哥 ，直到 約旦河 為止。
JOSH|16|8|這地界又從 他普亞 ，順著 加拿河 往西延伸，直通到海為止。這就是 以法蓮 支派按著宗族所得的地業。
JOSH|16|9|在 瑪拿西 人地業的一切城鎮和所屬的村莊中，也保留一些城鎮給 以法蓮 的子孫。
JOSH|16|10|他們卻沒有趕出住在 基色 的 迦南 人。 迦南 人就住在 以法蓮 人中，成為服勞役的僕人，直到今日。
JOSH|17|1|瑪拿西 是 約瑟 的長子，這是他的支派抽籤所得之地。 瑪拿西 的長子， 基列 的父親 瑪吉 ，因為是勇士，就得了 基列 和 巴珊 。
JOSH|17|2|瑪拿西 其餘的子孫，就是 亞比以謝 的子孫， 希勒 的子孫， 亞斯烈 的子孫， 示劍 的子孫， 希弗 的子孫， 示米大 的子孫，都按著宗族抽籤得了地。這都是 約瑟 的兒子 瑪拿西 子孫中各宗族的男丁。
JOSH|17|3|瑪拿西 的玄孫， 瑪吉 的曾孫， 基列 的孫子， 希弗 的兒子 西羅非哈 沒有兒子，只有女兒。他的女兒名叫 瑪拉 、 挪阿 、 曷拉 、 密迦 、 得撒 。
JOSH|17|4|她們來到 以利亞撒 祭司和 嫩 的兒子 約書亞 以及眾領袖面前，說：「耶和華曾吩咐 摩西 在我們兄弟中分產業給我們。」於是 約書亞 照耶和華的指示，在她們叔伯中，把產業分給她們。
JOSH|17|5|除了 約旦河 東的 基列 和 巴珊 地之外，還有十份的地業是屬於 瑪拿西 的，
JOSH|17|6|因為 瑪拿西 支派的女子也在男子中分得產業。 基列 地屬於 瑪拿西 其餘的子孫。
JOSH|17|7|瑪拿西 的地界是從 亞設 起，到 示劍 前面的 密米他 ，往右 到 隱‧他普亞 居民之地。
JOSH|17|8|他普亞 地歸於 瑪拿西 ，只是 瑪拿西 邊界的 他普亞城 卻歸於 以法蓮 子孫。
JOSH|17|9|這地界從那裏下到 加拿河 。河南邊的城鎮雖然在 瑪拿西 境內，卻是屬於 以法蓮 的。 瑪拿西 的地界是在河的北邊直通到海為止。
JOSH|17|10|南邊屬於 以法蓮 ，北邊屬於 瑪拿西 ，以海為界；北邊達到 亞設 ，東邊達到 以薩迦 。
JOSH|17|11|瑪拿西 在 以薩迦 和 亞設 境內，有 伯‧善 和所屬的鄉鎮， 以伯蓮 和所屬的鄉鎮， 多珥 和所屬鄉鎮的居民；還有 隱‧多珥 和所屬鄉鎮的居民， 他納 和所屬鄉鎮的居民， 米吉多 和所屬鄉鎮的居民，共三個山岡 。
JOSH|17|12|只是 瑪拿西 的子孫不能趕出這些城鎮的居民， 迦南 人仍堅持住在那地。
JOSH|17|13|以色列 人強盛的時候，就叫 迦南 人做苦工，沒有把他們全然趕走。
JOSH|17|14|約瑟 的子孫對 約書亞 說：「耶和華到如今這樣賜福給我，我百姓眾多，你為甚麼只給我抽一籤，分一份的土地為業呢？」
JOSH|17|15|約書亞 對他們說：「如果你百姓眾多，而 以法蓮 山區太窄小，那麼你可以上 比利洗 人和 利乏音 人之地的樹林中，在那裏開墾。」
JOSH|17|16|約瑟 的子孫說：「那山區容不下我們，而且住平原的 迦南 人，就是住 伯‧善 和所屬的鄉鎮，以及住在 耶斯列 平原的人，都有鐵的戰車。」
JOSH|17|17|約書亞 對 約瑟 家，就是 以法蓮 和 瑪拿西 人，說：「你百姓眾多，並且強大，不可只有一籤而已。
JOSH|17|18|那山區也要歸你，雖然是樹林，你可以去開墾，邊緣之地也必歸你。 迦南 人縱然強盛，有鐵的戰車，你也能把他們趕出去。」
JOSH|18|1|以色列 全會眾都聚集在 示羅 ，把會幕設立在那裏。那地已經被他們征服了。
JOSH|18|2|以色列 人中剩下七個支派還沒有分得他們的地業。
JOSH|18|3|約書亞 對 以色列 人說：「耶和華－你們列祖的上帝所賜給你們的地，你們耽延不去得，要到幾時呢？
JOSH|18|4|你們每支派要選三個人，我好派他們去，他們要起身走遍那地，按照各支派應得的地業寫明，然後回到我這裏來。
JOSH|18|5|他們要把地分成七份。 猶大 在南方，住在他的境內。 約瑟 家在北方，住在他們的境內。
JOSH|18|6|你們把地劃成七份之後，就要把所寫的帶到我這裏來。我要在耶和華－我們的上帝面前，為你們抽籤。
JOSH|18|7|利未 人在你們中間沒有分得地業，因為耶和華祭司的職分就是他們的產業。 迦得 支派、 呂便 支派和 瑪拿西 半支派已經在 約旦河 東得了地業，是耶和華的僕人 摩西 給他們的。」
JOSH|18|8|那些去劃地的人起來正要去的時候， 約書亞 吩咐他們說：「你們去走遍那地，把地劃分以後，就回到我這裏來。我要在 示羅 這裏，在耶和華面前為你們抽籤。」
JOSH|18|9|那些人就去了，走遍那地，按照城鎮把地劃成七份，寫在冊上，回到 示羅 營中 約書亞 那裏。
JOSH|18|10|約書亞 就在 示羅 ，在耶和華面前為他們抽籤。 約書亞 按照 以色列 人的支派，在那裏把地分給他們。
JOSH|18|11|便雅憫 支派，按著宗族抽籤所得之地，是在 猶大 子孫和 約瑟 子孫之間。
JOSH|18|12|他們北邊的地界是從 約旦河 起，上到 耶利哥 斜坡的北邊，再往西上到山區，直到 伯‧亞文 的曠野。
JOSH|18|13|這地界從那裏往南經過 路斯 ，直到 路斯 的斜坡， 路斯 就是 伯特利 ，又下到 亞他錄‧亞達 ，直到 下伯‧和崙 南邊的山。
JOSH|18|14|這地界往西延伸，又轉向南，從 伯‧和崙 南邊對面的山，直通到 猶大 人的城 基列‧巴力 ， 基列‧巴力 就是 基列‧耶琳 。這就是西邊的地界。
JOSH|18|15|南邊是從 基列‧耶琳 的頂端為起點，這地界往西 通到 尼弗多亞 水泉，
JOSH|18|16|這地界又下到 欣嫩子谷 對面山的邊緣，就是 利乏音谷 的北邊；又下到 欣嫩谷 ，沿著 耶布斯 斜坡的南邊，下到 隱‧羅結 ；
JOSH|18|17|又往北轉彎，通到 隱‧示麥 ，直到 亞都冥 斜坡對面的 基利綠 ，又下到 呂便 之子 波罕 的磐石，
JOSH|18|18|又往北經過 亞拉巴 對面的斜坡 ，下到 亞拉巴 。
JOSH|18|19|這地界又經過 伯‧曷拉 斜坡的北邊，直通到 鹽海 的北灣，就是 約旦河 的南端為止。這就是南邊的地界。
JOSH|18|20|東邊的地界是 約旦河 。這是 便雅憫 人按著宗族，照著他們四圍的邊界所得的地業。
JOSH|18|21|便雅憫 支派按著宗族所得的城鎮就是： 耶利哥 、 伯‧曷拉 、 伊麥‧基悉 、
JOSH|18|22|伯‧亞拉巴 、 洗瑪臉 、 伯特利 、
JOSH|18|23|亞文 、 巴拉 、 俄弗拉 、
JOSH|18|24|基法‧阿摩尼 、 俄弗尼 和 迦巴 ，共十二座城，以及所屬的村莊；
JOSH|18|25|又有 基遍 、 拉瑪 、 比錄 、
JOSH|18|26|米斯巴 、 基非拉 、 摩撒 、
JOSH|18|27|利堅 、 伊利毗勒 、 他拉拉 、
JOSH|18|28|洗拉 、 以利弗 、 耶布斯 ， 耶布斯 就是 耶路撒冷 ， 基比亞 、 基列 ，共十四座城，以及所屬的村莊。這是 便雅憫 人按著宗族所得的地業。
JOSH|19|1|第二籤是 西緬 ，是 西緬 支派的人按著宗族抽出的，他們所得的地業是在 猶大 人地業的中間。
JOSH|19|2|他們所得為業之地是： 別是巴 ，或名 示巴 ， 摩拉大 、
JOSH|19|3|哈薩‧書亞 、 巴拉 、 以森 、
JOSH|19|4|伊勒多臘 、 比土力 、 何珥瑪 、
JOSH|19|5|洗革拉 、 伯‧瑪加博 、 哈薩‧蘇撒 、
JOSH|19|6|伯‧利巴勿 、 沙魯險 ，共十三座城，還有所屬的村莊；
JOSH|19|7|又有 亞因 、 利門 、 以帖 、 亞珊 ，共四座城，還有所屬的村莊；
JOSH|19|8|以及這些城鎮周圍一切的村莊，直到 巴拉‧比珥 ，就是 尼革夫 的 拉瑪 。這是 西緬 支派的人按著宗族所得的地業。
JOSH|19|9|西緬 人的地業取自 猶大 人的土地，因為 猶大 人所得的份過多，所以 西緬 人從 猶大 人的地業中取了地業。
JOSH|19|10|第三籤是 西布倫 人按著宗族抽到的。他們地業的邊界延伸到 撒立 。
JOSH|19|11|他們的地界往西，上到 瑪拉拉 ，達到 大巴設 ，又達到 約念 前面的河。
JOSH|19|12|又從 撒立 往東轉到向日出的方向，經過 吉斯綠‧他泊 的邊界，到 大比拉 ，又上到 雅非亞 。
JOSH|19|13|又從那裏往東，經過 迦特‧希弗 ，到 以特‧加汛 ，通到 臨門 ，延伸到 尼亞 。
JOSH|19|14|這地界在北邊繞過 尼亞 ，到 哈拿頓 ，直通到 伊弗他‧伊勒谷 ，
JOSH|19|15|包括 加他 、 拿哈拉 、 伸崙 、 以大拉 、 伯利恆 ，共十二座城，還有所屬的村莊。
JOSH|19|16|這些城鎮和所屬的村莊是 西布倫 人按著宗族所得的地業。
JOSH|19|17|第四籤是 以薩迦 ，是 以薩迦 人按著宗族抽出的。
JOSH|19|18|他們的地界是到 耶斯列 、 基蘇律 、 書念 、
JOSH|19|19|哈弗連 、 示按 、 亞拿哈拉 、
JOSH|19|20|拉璧 、 基善 、 亞別 、
JOSH|19|21|利篾 、 隱‧干寧 、 隱‧哈大 、 伯‧帕薛 。
JOSH|19|22|這地界達到 他泊 、 沙哈洗瑪 、 伯‧示麥 ，他們的地界直通到 約旦河 為止，共十六座城，還有所屬的村莊。
JOSH|19|23|這些城鎮和所屬的村莊是 以薩迦 支派的人按著宗族所得的地業。
JOSH|19|24|第五籤是 亞設 支派的人按著宗族抽出的。
JOSH|19|25|他們的地界是 黑甲 、 哈利 、 比田 、 押煞 、
JOSH|19|26|亞拉米勒 、 亞末 、 米沙勒 ，往西達到 迦密 ，又到 希曷‧立納 ，
JOSH|19|27|又轉到向日出方向的 伯‧大袞 ，達到 細步綸 ；又往北到 伊弗他‧伊勒谷 ，到 伯‧以墨 和 尼業 ，也通到 迦步勒 的左邊 ，
JOSH|19|28|又到 義伯崙 、 利合 、 哈們 、 加拿 ，直到 西頓 大城。
JOSH|19|29|這地界轉到 拉瑪 ，直到堅固的 推羅城 。這地界又轉到 何薩 ，靠近 亞革悉 一帶的地方 ，直通到海為止。
JOSH|19|30|又有 烏瑪 、 亞弗 、 利合 ，共二十二座城，還有所屬的村莊。
JOSH|19|31|這些城鎮和所屬的村莊是 亞設 支派的人按著宗族所得的地業。
JOSH|19|32|第六籤是 拿弗他利 人，是 拿弗他利 人按著宗族抽出的。
JOSH|19|33|他們的地界是從 希利弗 ，從 撒拿音 的橡樹、 亞大米‧尼吉 和 雅比聶 ，直到 拉共 ，直通到 約旦河 為止。
JOSH|19|34|這地界往西轉到 亞斯納‧他泊 ，從那裏通到 戶割 ，南邊達到 西布倫 ，西邊達到 亞設 ，向日出的方向達到 約旦河 的 猶大 。
JOSH|19|35|堅固的城有 西丁 、 側耳 、 哈末 、 拉甲 、 基尼烈 、
JOSH|19|36|亞大瑪 、 拉瑪 、 夏瑣 、
JOSH|19|37|基低斯 、 以得來 、 隱‧夏瑣 、
JOSH|19|38|以利穩 、 密大‧伊勒 、 和璉 、 伯‧亞納 、 伯‧示麥 ，共十九座城，還有所屬的村莊。
JOSH|19|39|這些城鎮和所屬的村莊是 拿弗他利 支派的人按著宗族所得的地業。
JOSH|19|40|但 支派，按著宗族，抽到第七籤。
JOSH|19|41|他們地業的邊界是 瑣拉 、 以實陶 、 伊珥‧示麥 、
JOSH|19|42|沙拉賓 、 亞雅崙 、 伊提拉 、
JOSH|19|43|以倫 、 亭拿 、 以革倫 、
JOSH|19|44|伊利提基 、 基比頓 、 巴拉 、
JOSH|19|45|伊胡得 、 比尼‧比拉 、 迦特‧臨門 、
JOSH|19|46|美‧耶昆 、 拉昆 ，以及 約帕 對面的地界。
JOSH|19|47|當 但 的子孫失去他們疆土的時候，就上去攻取 利善 ，用刀擊殺城中的人，得了那城，住在城中，以他們祖先 但 的名字將 利善 改名為 但 。
JOSH|19|48|這些城鎮和所屬的村莊是 但 支派的人按著宗族所得的地業。
JOSH|19|49|以色列 人按著疆土完成了地業的分配，就在他們中間把地給 嫩 的兒子 約書亞 為業。
JOSH|19|50|他們照著耶和華的指示，把 約書亞 所要的城，就是 以法蓮 山區的 亭拿‧西拉 給了他。 約書亞 修建那城，住在城中。
JOSH|19|51|這就是 以利亞撒 祭司和 嫩 的兒子 約書亞 ，以及 以色列 人各支派父系的領袖，在 示羅 會幕的門口，耶和華面前抽籤所分的地業。這樣， 他們就完成了分地的事。
JOSH|20|1|耶和華吩咐 約書亞 說：
JOSH|20|2|「你吩咐 以色列 人說：『你們要照我藉 摩西 所吩咐你們的，為自己設立逃城，
JOSH|20|3|使那無意中誤殺人的，可以逃到那裏。這些要作為你們逃避報血仇者的城。
JOSH|20|4|殺人者要逃到這些城中的一座，站在城門口，把他的事情陳訴給那城的長老聽。他們就要接他入城，給他地方，讓他住在他們中間。
JOSH|20|5|若是報血仇者追上了他，長老不可把他交在報血仇者的手裏，因為他是無意中殺了鄰舍的，並非過去彼此之間有仇恨。
JOSH|20|6|他要住在那城裏，直到他站在會眾面前受審判；等到當時的大祭司死後，殺人者才可以回到本城本家，就是他所逃出來的那城。』」
JOSH|20|7|於是， 以色列 人劃分 拿弗他利 山區 加利利 的 基低斯 、 以法蓮 山區的 示劍 和 猶大 山區的 基列‧亞巴 ， 基列‧亞巴 就是 希伯崙 。
JOSH|20|8|他們在 約旦河 的另一邊，就是 耶利哥 的東邊，從 呂便 支派中，在曠野的平原設立 比悉 ，從 迦得 支派中設立 基列 的 拉末 ，從 瑪拿西 支派中設立 巴珊 的 哥蘭 。
JOSH|20|9|這都是為 以色列 眾人和在他們中間寄居的外人所指定的城鎮，使凡誤殺人者可以逃到那裏，不至於死在報血仇者的手中，直到他站在會眾面前受審判 。
JOSH|21|1|利未 人的眾族長近前來到 以利亞撒 祭司和 嫩 的兒子 約書亞 ，以及 以色列 人各支派父系的領袖那裏，
JOSH|21|2|在 迦南 地的 示羅 對他們說：「從前耶和華曾藉著 摩西 吩咐給我們城鎮居住，以及城鎮的郊外供我們牧養牲畜。」
JOSH|21|3|於是 以色列 人照耶和華的指示，從自己的地業中，把這些城鎮和城鎮的郊外給了 利未 人。
JOSH|21|4|哥轄 族抽了籤。 利未 人中 亞倫 祭司的子孫，從 猶大 支派、 西緬 支派、 便雅憫 支派的地業中，抽籤得了十三座城。
JOSH|21|5|哥轄 其餘的子孫，從 以法蓮 支派、 但 支派、 瑪拿西 半支派宗族的地業中，抽籤得了十座城。
JOSH|21|6|革順 的子孫，從 以薩迦 支派、 亞設 支派、 拿弗他利 支派、住 巴珊 的 瑪拿西 半支派宗族的地業中，抽籤得了十三座城。
JOSH|21|7|米拉利 的子孫，按著宗族，從 呂便 支派、 迦得 支派、 西布倫 支派的地業中，得了十二座城。
JOSH|21|8|以色列 人照耶和華藉 摩西 所吩咐的，把這些城鎮和城鎮的郊外，抽籤給 利未 人。
JOSH|21|9|他們從 猶大 支派和 西緬 支派的地業中，給了以下所記名字的各城，
JOSH|21|10|就是給 利未 人 哥轄 宗族的 亞倫 子孫，因為他們抽到第一籤：
JOSH|21|11|把 猶大 山區的 基列‧亞巴 ，就是 希伯崙 ，和四圍的郊野給了他們。 亞巴 是 亞衲 族的祖先。
JOSH|21|12|但是，這城的田地和所屬的村莊卻給了 耶孚尼 的兒子 迦勒 為業。
JOSH|21|13|他們把 希伯崙 ，就是誤殺人的逃城和城的郊外，給了 亞倫 祭司的子孫；又給了 立拿 和城的郊外、
JOSH|21|14|雅提珥 和城的郊外、 以實提莫 和城的郊外、
JOSH|21|15|何崙 和城的郊外、 底璧 和城的郊外、
JOSH|21|16|亞因 和城的郊外、 淤他 和城的郊外，以及 伯‧示麥 和城的郊外，共九座城，都是從這二支派中分出來的。
JOSH|21|17|又從 便雅憫 支派的地業中給了 基遍 和城的郊外、 迦巴 和城的郊外、
JOSH|21|18|亞拿突 和城的郊外，以及 亞勒們 和城的郊外，共四座城。
JOSH|21|19|亞倫 子孫作祭司的共有十三座城，以及城的郊外。
JOSH|21|20|利未 人 哥轄 的宗族，就是 哥轄 其餘的子孫，抽籤所得的城是從 以法蓮 支派來的。
JOSH|21|21|他們把 以法蓮 山區的 示劍 ，就是誤殺人的逃城和城的郊外給了 哥轄 其餘的子孫；又給了 基色 和城的郊外、
JOSH|21|22|基伯先 和城的郊外，以及 伯‧和崙 和城的郊外，共四座城。
JOSH|21|23|又從 但 支派的地業中給了 伊利提基 和城的郊外、 基比頓 和城的郊外、
JOSH|21|24|亞雅崙 和城的郊外，以及 迦特‧臨門 和城的郊外，共四座城。
JOSH|21|25|又從 瑪拿西 半支派的地業中給了 他納 和城的郊外，以及 迦特‧臨門 和城的郊外，共兩座城。
JOSH|21|26|哥轄 其餘的子孫共有十座城，以及城的郊外。
JOSH|21|27|利未 人宗族中 革順 的子孫，從 瑪拿西 半支派的地業中所得的是 巴珊 的 哥蘭 ，就是誤殺人的逃城和城的郊外，以及 比‧施提拉 和城的郊外，共兩座城。
JOSH|21|28|從 以薩迦 支派的地業中所得的是 基善 和城的郊外、 大比拉 和城的郊外、
JOSH|21|29|耶末 和城的郊外，以及 隱‧干寧 和城的郊外，共四座城。
JOSH|21|30|從 亞設 支派的地業中所得的是 米沙勒 和城的郊外、 押頓 和城的郊外、
JOSH|21|31|黑甲 和城的郊外，以及 利合 和城的郊外，共四座城。
JOSH|21|32|從 拿弗他利 支派的地業中所得的是 加利利 的 基低斯 ，就是誤殺人的逃城和城的郊外、 哈末‧多珥 和城的郊外，以及 加珥坦 和城的郊外，共三座城。
JOSH|21|33|革順 人按著宗族共有十三個城，以及城的郊外。
JOSH|21|34|其餘的 利未 人，就是 米拉利 的子孫，按著宗族從 西布倫 支派的地業中所得的是 約念 和城的郊外、 加珥他 和城的郊外、
JOSH|21|35|丁拿 和城的郊外，以及 拿哈拉 和城的郊外，共四座城。
JOSH|21|36|從 呂便 支派的地業中所得的是 比悉 和城的郊外、 雅雜 和城的郊外、
JOSH|21|37|基底莫 和城的郊外，以及 米法押 和城的郊外，共四座城。
JOSH|21|38|從 迦得 支派的地業中所得的是 基列 的 拉末 ，就是誤殺人的逃城和城的郊外、 瑪哈念 和城的郊外、
JOSH|21|39|希實本 和城的郊外，以及 雅謝 和城的郊外，共四座城。
JOSH|21|40|利未 宗族其餘的人，就是 米拉利 的子孫，按著宗族抽籤所得的，共十二座城。
JOSH|21|41|利未 人在 以色列 人的地業中所得的城，共四十八個，還有城的郊外。
JOSH|21|42|這些城的四圍都有郊野，每個城都是如此。
JOSH|21|43|這樣，耶和華將從前向他們列祖起誓要給他們的全地賜給 以色列 人，他們就得了為業，住在其中。
JOSH|21|44|耶和華照著向他們列祖起誓所應許的一切，賜給他們全境安寧。他們所有的仇敵，沒有一個能在他們面前站立得住。耶和華把所有仇敵都交在他們手中。
JOSH|21|45|耶和華應許賜福給 以色列 家的話，一句都沒有落空，全都應驗了。
JOSH|22|1|此後， 約書亞 召了 呂便 人、 迦得 人和 瑪拿西 半支派的人來，
JOSH|22|2|對他們說：「耶和華的僕人 摩西 所吩咐你們的，你們都遵守了；我吩咐你們的話，你們也都聽從了。
JOSH|22|3|你們這許多日子，都沒有撇棄你們的弟兄，直到今日，並且遵守了耶和華你們上帝所吩咐的命令。
JOSH|22|4|如今耶和華－你們的上帝已經照著他所應許的，使你們的弟兄得享安寧。你們現在可以返回自己的帳棚，回到耶和華的僕人 摩西 在 約旦河 東所賜給你們為業之地。
JOSH|22|5|只是務要謹守遵行耶和華的僕人 摩西 所吩咐你們的誡命和律法，愛耶和華－你們的上帝，行他一切的道，守他的誡命，緊緊跟隨他，盡心盡性事奉他。」
JOSH|22|6|於是 約書亞 為他們祝福，送他們回去，他們就回到自己的帳棚去了。
JOSH|22|7|摩西 在 巴珊 曾把地業分給 瑪拿西 的半支派；然後 約書亞 在 約旦河 的西岸，在他們弟兄中，又把地業分給 瑪拿西 的另外半支派。 約書亞 送他們回帳棚的時候，為他們祝福，
JOSH|22|8|對他們說：「你們要把許多財物，許多牲畜，和金、銀、銅、鐵，以及許多衣服，帶回你們的帳棚去，要把你們從仇敵奪來的東西分給你們的眾弟兄。」
JOSH|22|9|於是 呂便 人、 迦得 人、 瑪拿西 半支派的人從 迦南 地的 示羅 起行，離開 以色列 人，回到他們已得為業的 基列 地，就是他們照耶和華藉 摩西 所吩咐而得的。
JOSH|22|10|呂便 人、 迦得 人和 瑪拿西 半支派的人到了 迦南 地的 約旦河 一帶地方，就在 約旦河 那裏築了一座壇，一座高大壯觀的壇。
JOSH|22|11|以色列 人聽見了，說：「看哪， 呂便 人、 迦得 人、 瑪拿西 半支派的人在 迦南 地對面， 約旦河 一帶地方， 以色列 人的境內，築了一座壇。」
JOSH|22|12|以色列 人一聽見，全會眾的 以色列 人就聚集在 示羅 ，要上去攻打他們。
JOSH|22|13|以色列 人派 以利亞撒 祭司的兒子 非尼哈 ，往 基列 地，到 呂便 人、 迦得 人和 瑪拿西 半支派的人那裏。
JOSH|22|14|和他同去的還有十個領袖， 以色列 每個支派在父家中各派一個領袖，這些人每一個在 以色列 族系中都是父家的領袖。
JOSH|22|15|他們來到 基列 地，到 呂便 人、 迦得 人和 瑪拿西 半支派的人那裏，對他們說：
JOSH|22|16|「耶和華全會眾這樣說：『你們今日離棄耶和華不跟從他，干犯 以色列 的上帝，悖逆耶和華，為自己築了一座壇，你們所犯的是何等的罪！
JOSH|22|17|從前我們在 毗珥 犯的罪孽，導致瘟疫臨到耶和華的會眾，甚至到今日都還沒有洗淨，這還算小事嗎？
JOSH|22|18|你們今日竟然離棄耶和華不跟從他！你們今日既然悖逆耶和華，明日他必向 以色列 全會眾發怒。
JOSH|22|19|若你們認為所得為業之地不潔淨，可以過來，到耶和華之地，就是耶和華的帳幕所居住之地，在我們中間得地業。你們卻不可悖逆耶和華，也不可背叛我們，在耶和華－我們上帝的壇以外為自己築壇。
JOSH|22|20|從前 謝拉 的曾孫 亞干 豈不是在那當滅的物上犯了罪，導致憤怒臨到 以色列 全會眾嗎？死在他所犯的罪中的，不只是他一個人而已！』」
JOSH|22|21|於是 呂便 人、 迦得 人、 瑪拿西 半支派的人回答 以色列 族系的領袖，說：
JOSH|22|22|「大能者上帝耶和華！大能者上帝耶和華！他已知道，願 以色列 人也知道，我們若有悖逆的行為，或是干犯耶和華，你今日就不要讓我們活著！
JOSH|22|23|若我們為自己築壇，離棄耶和華不跟從他，或將燔祭、素祭、平安祭獻在壇上，願耶和華親自追究。
JOSH|22|24|不是這樣！我們做這事的原因是懼怕將來你們的子孫對我們的子孫說：『你們與耶和華－ 以色列 的上帝有甚麼關係呢？
JOSH|22|25|因為耶和華以 約旦河 作我們和你們 呂便 人、 迦得 人的交界，所以你們在耶和華裏無份。』這樣，你們的子孫就使我們的子孫不再敬畏耶和華了。
JOSH|22|26|因此我們說：『不如為自己築一座壇，不是為獻燔祭，也不是為獻別樣的祭，
JOSH|22|27|而是為你我之間和後代子孫之間作證據，好使我們也在耶和華面前獻我們的燔祭、平安祭和別樣的祭來事奉他，免得你們的子孫將來對我們的子孫說，你們在耶和華裏無份。』
JOSH|22|28|所以我們說：『將來他們若對我們，或對我們的子孫這樣說，我們就可以回答說：你們看，我們列祖所築的壇是耶和華壇的樣式，這並不是為獻燔祭，也不是為獻別樣的祭，而是作為你們和我們之間的證據。』
JOSH|22|29|除了耶和華－我們上帝帳幕前的壇以外，我們絕沒有意思要為著獻燔祭、素祭和別樣的祭而另外築一座壇，悖逆耶和華，今日離棄不跟從他。」
JOSH|22|30|非尼哈 祭司與會眾中的領袖，就是與他同來那些 以色列 族系的領袖，聽見 呂便 人、 迦得 人、 瑪拿西 人所說的話，就都看為美。
JOSH|22|31|以利亞撒 祭司的兒子 非尼哈 對 呂便 人、 迦得 人、 瑪拿西 人說：「今日我們知道耶和華在我們中間，因為你們沒有向他犯悖逆的罪。現在你們把 以色列 人從耶和華的手中救出來了。」
JOSH|22|32|以利亞撒 祭司的兒子 非尼哈 與眾領袖離開了 呂便 人和 迦得 人，從 基列 地回 迦南 地，到了 以色列 人那裏，就把這事向他們回報。
JOSH|22|33|以色列 人看這事為美； 以色列 人就稱頌上帝，不再說要上去攻打 呂便 人和 迦得 人，毀壞他們所住的地了。
JOSH|22|34|呂便 人和 迦得 人給這壇起了名，因為這壇在我們之間見證耶和華是上帝。
JOSH|23|1|耶和華使 以色列 人從四圍所有的仇敵中得享安寧，已經有很多日子了。 約書亞 年紀老邁，
JOSH|23|2|就召了全 以色列 的眾長老、領袖、審判官和官長來，對他們說：「我年紀已經老邁。
JOSH|23|3|耶和華－你們的上帝因你們的緣故向這些國家所做的一切，你們都親眼看見了，那為你們作戰的是耶和華－你們的上帝。
JOSH|23|4|看，我已經把所剩下的列國，連同從 約旦河 起到 大海 日落的方向，我所剪除的列國，都抽籤分給你們各支派為業了。
JOSH|23|5|耶和華－你們的上帝必將他們從你們面前趕出去，使他們離開你們，你們就必得他們的地為業，正如耶和華－你們的上帝向你們所應許的。
JOSH|23|6|你們要大大壯膽，謹守遵行寫在 摩西 律法書上的一切話，不可偏離左右。
JOSH|23|7|不可與你們中間所剩下的這些國家往來。你們不可提他們神明的名，不可指著它們起誓，不可事奉它們，也不可敬拜它們。
JOSH|23|8|只要緊緊跟隨耶和華－你們的上帝，就像你們直到今日所做的。
JOSH|23|9|因為耶和華已經把又大又強的列國從你們面前趕出；直到今日，沒有一人能在你們面前站立得住。
JOSH|23|10|你們一人必追趕千人，因為耶和華－你們的上帝照他向你們所應許的，為你們作戰。
JOSH|23|11|你們要分外謹慎，愛耶和華－你們的上帝。
JOSH|23|12|你們若斷然轉離，緊緊跟隨你們中間所剩下的這些國家，彼此結親，互相往來，
JOSH|23|13|就要確實知道，耶和華－你們的上帝必不再將他們從你們面前趕出；他們卻要成為你們的羅網、圈套、肋上的鞭、眼中的刺，直到你們在耶和華－你們上帝所賜的這美地上滅亡。
JOSH|23|14|「看哪，我今日要走世人必走的路了。你們要一心一意知道，耶和華－你們上帝所應許要賜給你們的一切福氣，沒有一件落空，都應驗在你們身上了。
JOSH|23|15|耶和華－你們的上帝所應許的一切福氣怎樣臨到你們身上，耶和華也必照樣使各樣災禍臨到你們身上，直到他把你們從耶和華－你們上帝所賜給你們的這美地上除滅。
JOSH|23|16|你們若違背耶和華－你們上帝吩咐你們所守的約，去事奉別神，敬拜它們，耶和華的怒氣必向你們發作，使你們在他所賜給你們的美地上迅速滅亡。」
JOSH|24|1|約書亞 召集 以色列 的眾支派到 示劍 ，他召了 以色列 的長老、領袖、審判官和官長來；他們都站在上帝面前。
JOSH|24|2|約書亞 對眾百姓說：「耶和華－ 以色列 的上帝如此說：『古時你們的列祖，就是 亞伯拉罕 和 拿鶴 的父親 他拉 ，住在 大河 那邊事奉別神。
JOSH|24|3|我將你們的祖宗 亞伯拉罕 從 大河 那邊帶出來，領他走遍 迦南 全地，又使他的子孫眾多。我把 以撒 賜給他，
JOSH|24|4|我又把 雅各 和 以掃 賜給 以撒 ，將 西珥山 賜給 以掃 為業。但 雅各 和他的子孫下到 埃及 去了。
JOSH|24|5|我差遣 摩西 和 亞倫 ，照我在 埃及 中間所做的，降災與 埃及 ，然後把你們領出來。
JOSH|24|6|我領你們的祖宗出 埃及 ，你們就到了 紅海 。 埃及 人帶領戰車騎兵，追趕你們的祖宗到 紅海 。
JOSH|24|7|你們的祖宗哀求耶和華，他就用黑暗把你們和 埃及 人隔開了，又使海水衝向 埃及 人，淹沒他們。我在 埃及 所做的，你們都親眼見過。你們在曠野住了很多日子。
JOSH|24|8|我領你們到 約旦河 東 亞摩利 人所住之地。他們與你們爭戰，我把他們交在你們手中，你們就得了他們的地為業。我也在你們面前滅絕他們。
JOSH|24|9|那時， 摩押 王 西撥 的兒子 巴勒 起來攻擊 以色列 人，派人去召 比珥 的兒子 巴蘭 來詛咒你們。
JOSH|24|10|但我不願聽 巴蘭 ，所以他反而為你們連連祝福。這樣，我救了你們脫離他的手。
JOSH|24|11|你們過了 約旦河 ，來到 耶利哥 。 耶利哥 人、 亞摩利 人、 比利洗 人、 迦南 人、 赫 人、 革迦撒 人、 希未 人、 耶布斯 人都與你們爭戰，我卻把他們交在你們手裏。
JOSH|24|12|我派遣瘟疫 在你們前面，將 亞摩利 人的兩個王從你們面前趕出，並不是用你的刀，也不是用你的弓。
JOSH|24|13|我賜給你們的地，不是你們開墾的；我賜給你們的城鎮，不是你們建造的。你們卻住在其中，又得吃那不是你們栽植的葡萄園和橄欖園的果子。』
JOSH|24|14|「現在你們要敬畏耶和華，誠心誠意事奉他，除掉你們列祖在 大河 那邊和在 埃及 事奉的神明，事奉耶和華。
JOSH|24|15|若你們認為事奉耶和華不好，今日就可以選擇所要事奉的：是你們列祖在 大河 那邊所事奉的神明，或是你們所住這地 亞摩利 人的神明呢？至於我和我家，我們必定事奉耶和華。」
JOSH|24|16|百姓回答說：「我們絕不離棄耶和華去事奉別神。
JOSH|24|17|因為耶和華－我們的上帝曾領我們和我們的祖宗從 埃及 地為奴之家出來，在我們眼前行了那些大神蹟，並在我們所行的一切路上，和所經過的各民族中保護了我們。
JOSH|24|18|耶和華又把各民族和住此地的 亞摩利 人都從我們面前趕出去。所以，我們也必事奉耶和華，因為他是我們的上帝。」
JOSH|24|19|約書亞 對百姓說：「你們不能事奉耶和華，因為他是神聖的上帝，是忌邪 的上帝，必不赦免你們的過犯罪惡。
JOSH|24|20|你們若離棄耶和華去事奉外邦的神明，耶和華在降福之後，必轉而降禍給你們，把你們滅絕。」
JOSH|24|21|百姓對 約書亞 說：「不，我們要事奉耶和華。」
JOSH|24|22|約書亞 對百姓說：「你們選擇耶和華，要事奉他，你們自己作證吧！」他們說：「我們願意作證。」
JOSH|24|23|「現在，你們要除掉你們中間外邦的神明，專心歸向耶和華－ 以色列 的上帝。」
JOSH|24|24|百姓對 約書亞 說：「我們必事奉耶和華－我們的上帝，聽從他的話。」
JOSH|24|25|那日， 約書亞 就與百姓立約，在 示劍 為他們制定律例典章。
JOSH|24|26|約書亞 把這些話寫在上帝的律法書上，又拿一塊大石頭立在橡樹下耶和華聖所的旁邊。
JOSH|24|27|約書亞 對眾百姓說：「看哪，這石頭可以向我們作見證，因為它聽見了耶和華所吩咐我們的一切話；這石頭將向你們作見證，免得你們背叛你們的上帝。」
JOSH|24|28|於是 約書亞 解散百姓，各自回到自己的地業去了。
JOSH|24|29|這些事以後，耶和華的僕人， 嫩 的兒子 約書亞 死了，那時他一百一十歲。
JOSH|24|30|以色列 人把他葬在他自己地業的境內， 以法蓮 山區的 亭拿‧西拉 ，在 迦實山 的北邊。
JOSH|24|31|約書亞 在世的日子和他死了以後，那些知道耶和華為 以色列 所做一切事的長老還在世的時候， 以色列 人事奉耶和華。
JOSH|24|32|以色列 人把從 埃及 所帶來 約瑟 的骸骨安葬在 示劍 ，就是 雅各 從前用一百可錫塔 向 示劍 的父親 哈抹 的眾子所買的那塊地；這塊地就成了 約瑟 子孫的產業。
JOSH|24|33|亞倫 的兒子 以利亞撒 也死了，他們把他葬在他兒子 非尼哈 所得 以法蓮 山區的小山上 。
