OBAD|1|1|Visio Abdiae.Haec dicit Dominus Deus ad Edom.Auditum audivimus a Domino,et legatus ad gentes missus est: Surgite, et consurgamusadversus eum in proelium! ".
OBAD|1|2|" Ecce parvulum te dabo in gentibus,contemptibilis tu es valde.
OBAD|1|3|Superbia cordis tui decepit tehabitantem in scissuris petrae,exaltantem solium suum;qui dicit in corde suo:Quis detrahet me in terram?".
OBAD|1|4|Si exaltatus fueris ut aquilaet si inter sidera posueris nidum tuum,inde detraham te ",dicit Dominus.
OBAD|1|5|Si fures introissent ad te,si latrones per noctem,quomodo periisses!Nonne furati essent sufficientia sibi?Si vindemiatores introissent ad te,nonne racemos tantum reliquissent?
OBAD|1|6|Quomodo scrutati sunt Esau?Investigaverunt abscondita eius.
OBAD|1|7|Usque ad terminum eiecerunt te,omnes viri foederis tui deceperunt te,invaluerunt adversum te viri pacis tuae;qui comedunt tecum, ponent insidias subter te.Non est prudentia in eo.
OBAD|1|8|" Numquid non in die illa,dicit Dominus,perdam sapientes de Edomet prudentiam de monte Esau?
OBAD|1|9|Et timebunt fortes tui Theman,ut intereat omnis vir de monte Esau.
OBAD|1|10|Propter interfectionemet propter iniquitatemin fratrem tuum Iacoboperiet te confusio,et peribis in aeternum.
OBAD|1|11|In die cum stares ex adverso,quando capiebant alieni exercitum eius,et extranei ingrediebantur portas eiuset super Ierusalem mittebant sortem,tu quoque eras quasi unus ex eis ".
OBAD|1|12|Et non respicies diem fratris tui,diem calamitatis eius;et non laetaberis super filios Iudaein die perditionis eorum;et non magnificabis os tuumin die angustiae.
OBAD|1|13|Neque ingredieris portam populi meiin die ruinae eorum;neque respicies et tu malum eiusin die vastitatis illiuset non mittes manum in opes eiusin die vastitatis illius;
OBAD|1|14|neque stabis in exitibus,ut interficias eos, qui fugerint,et non trades reliquos eiusin die tribulationis.
OBAD|1|15|Quoniam iuxta est dies Dominisuper omnes gentes:sicut fecisti, fiet tibi,retributio tua convertetur in caput tuum.
OBAD|1|16|Quomodo enim bibistis super montem sanctum meum,bibent omnes gentes iugiter;et bibent et absorbebuntet erunt quasi non fuerint.
OBAD|1|17|Et in monte Sion erit salvatio,et erit sanctum;et possidebit domus Iacobeos, qui se possederant.
OBAD|1|18|Et erit domus Iacob ignis,et domus Ioseph flamma,et domus Esau stipula;et succendentur in eis, et devorabunt eos,et non erunt reliquiae domus Esau,quia Dominus locutus est.
OBAD|1|19|Et hereditabunt austrum,montem Esau,et Sephelam Philisthim;et possidebunt regionem Ephraimet regionem Samariae,et Beniamin possidebit Galaad;
OBAD|1|20|et transmigratio prima filiorum Israelpossidebit terram Chananaeorum usque ad Sareptam;et transmigratio Ierusalem, quae in Sapharad est,possidebit civitates austri.
OBAD|1|21|Et ascendent salvatores in montem Sioniudicare montem Esau,et erit Domino regnum.
