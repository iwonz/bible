EZEK|1|1|et factum est in tricesimo anno in quarto mense in quinta mensis cum essem in medio captivorum iuxta fluvium Chobar aperti sunt caeli et vidi visiones Dei
EZEK|1|2|in quinta mensis ipse est annus quintus transmigrationis regis Ioachin
EZEK|1|3|factum est verbum Domini ad Hiezecihel filium Buzi sacerdotem in terra Chaldeorum secus flumen Chobar et facta est super eum ibi manus Domini
EZEK|1|4|et vidi et ecce ventus turbinis veniebat ab aquilone et nubes magna et ignis involvens et splendor in circuitu eius et de medio eius quasi species electri id est de medio ignis
EZEK|1|5|et ex medio eorum similitudo quattuor animalium et hic aspectus eorum similitudo hominis in eis
EZEK|1|6|et quattuor facies uni et quattuor pinnae uni
EZEK|1|7|et pedes eorum pedes recti et planta pedis eorum quasi planta pedis vituli et scintillae quasi aspectus aeris candentis
EZEK|1|8|et manus hominis sub pinnis eorum in quattuor partibus et facies et pinnas per quattuor partes habebant
EZEK|1|9|iunctaeque erant pinnae eorum alterius ad alterum non revertebantur cum incederent sed unumquodque ante faciem suam gradiebatur
EZEK|1|10|similitudo autem vultus eorum facies hominis et facies leonis a dextris ipsorum quattuor facies autem bovis a sinistris ipsorum quattuor et facies aquilae ipsorum quattuor
EZEK|1|11|et facies eorum et pinnae eorum extentae desuper duae pinnae singulorum iungebantur et duae tegebant corpora eorum
EZEK|1|12|et unumquodque coram facie sua ambulabat ubi erat impetus spiritus illuc gradiebantur nec revertebantur cum ambularent
EZEK|1|13|et similitudo animalium aspectus eorum quasi carbonum ignis ardentium et quasi aspectus lampadarum haec erat visio discurrens in medio animalium splendor ignis et de igne fulgor egrediens
EZEK|1|14|et animalia ibant et revertebantur in similitudinem fulguris coruscantis
EZEK|1|15|cumque aspicerem animalia apparuit rota una super terram iuxta animalia habens quattuor facies
EZEK|1|16|et aspectus rotarum et opus earum quasi visio maris et una similitudo ipsarum quattuor et aspectus earum et opera quasi sit rota in medio rotae
EZEK|1|17|per quattuor partes earum euntes ibant et non revertebantur cum ambularent
EZEK|1|18|statura quoque erat rotis et altitudo et horribilis aspectus et totum corpus plenum oculis in circuitu ipsarum quattuor
EZEK|1|19|cumque ambularent animalia ambulabant pariter et rotae iuxta ea et cum elevarentur animalia de terra elevabantur simul et rotae
EZEK|1|20|quocumque ibat spiritus illuc eunte spiritu et rotae pariter levabantur sequentes eum spiritus enim vitae erat in rotis
EZEK|1|21|cum euntibus ibant et cum stantibus stabant et cum elevatis a terra pariter elevabantur et rotae sequentes ea quia spiritus vitae erat in rotis
EZEK|1|22|et similitudo super caput animalium firmamenti quasi aspectus cristalli horribilis et extenti super capita eorum desuper
EZEK|1|23|sub firmamento autem pinnae eorum rectae alterius ad alterum unumquodque duabus alis velabat corpus suum et alterum similiter velabatur
EZEK|1|24|et audiebam sonum alarum quasi sonum aquarum multarum quasi sonum sublimis Dei cum ambularent quasi sonus erat multitudinis ut sonus castrorum cumque starent dimittebantur pinnae eorum
EZEK|1|25|nam cum fieret vox supra firmamentum quod erat super caput eorum stabant et submittebant alas suas
EZEK|1|26|et super firmamentum quod erat inminens capiti eorum quasi aspectus lapidis sapphyri similitudo throni et super similitudinem throni similitudo quasi aspectus hominis desuper
EZEK|1|27|et vidi quasi speciem electri velut aspectum ignis intrinsecus eius per circuitum a lumbis eius et desuper et a lumbis eius usque deorsum vidi quasi speciem ignis splendentis in circuitu
EZEK|1|28|velut aspectum arcus cum fuerit in nube in die pluviae hic erat aspectus splendoris per gyrum
EZEK|2|1|haec visio similitudinis gloriae Domini et vidi et cecidi in faciem meam et audivi vocem loquentis et dixit ad me fili hominis sta supra pedes tuos et loquar tecum
EZEK|2|2|et ingressus est in me spiritus postquam locutus est mihi et statuit me supra pedes meos et audivi loquentem ad me
EZEK|2|3|et dicentem fili hominis mitto ego te ad filios Israhel ad gentes apostatrices quae recesserunt a me patres eorum praevaricati sunt pactum meum usque ad diem hanc
EZEK|2|4|et filii dura facie et indomabili corde sunt ad quos ego mitto te et dices ad eos haec dicit Dominus Deus
EZEK|2|5|si forte vel ipsi audiant et si forte quiescant quoniam domus exasperans est et scient quia propheta fuerit in medio eorum
EZEK|2|6|tu ergo fili hominis ne timeas eos neque sermones eorum metuas quoniam increduli et subversores sunt tecum et cum scorpionibus habitas verba eorum ne timeas et vultus eorum ne formides quia domus exasperans est
EZEK|2|7|loqueris ergo verba mea ad eos si forte audiant et quiescant quoniam inritatores sunt
EZEK|2|8|tu autem fili hominis audi quaecumque loquor ad te et noli esse exasperans sicut domus exasperatrix est aperi os tuum et comede quaecumque ego do tibi
EZEK|2|9|et vidi et ecce manus missa ad me in qua erat involutus liber et expandit illum coram me qui erat scriptus intus et foris et scriptae erant in eo lamentationes et carmen et vae
EZEK|3|1|et dixit ad me fili hominis quodcumque inveneris comede comede volumen istud et vadens loquere ad filios Israhel
EZEK|3|2|et aperui os meum et cibavit me volumine illo
EZEK|3|3|et dixit ad me fili hominis venter tuus comedet et viscera tua conplebuntur volumine isto quod ego do tibi et comedi illud et factum est in ore meo sicut mel dulce
EZEK|3|4|et dixit ad me fili hominis vade ad domum Israhel et loqueris verba mea ad eos
EZEK|3|5|non enim ad populum profundi sermonis et ignotae linguae tu mitteris ad domum Israhel
EZEK|3|6|neque ad populos multos profundi sermonis et ignotae linguae quorum non possis audire sermones et si ad illos mittereris ipsi audirent te
EZEK|3|7|domus autem Israhel nolent audire te quia nolunt audire me omnis quippe domus Israhel adtrita fronte est et duro corde
EZEK|3|8|ecce dedi faciem tuam valentiorem faciebus eorum et frontem tuam duriorem frontibus eorum
EZEK|3|9|ut adamantem et ut silicem dedi faciem tuam ne timeas eos neque metuas a facie eorum quia domus exasperans est
EZEK|3|10|et dixit ad me fili hominis omnes sermones meos quos loquor ad te adsume in corde tuo et auribus tuis audi
EZEK|3|11|et vade ingredere ad transmigrationem ad filios populi tui et loqueris ad eos et dices eis haec dicit Dominus Deus si forte audiant et quiescant
EZEK|3|12|et adsumpsit me spiritus et audivi post me vocem commotionis magnae benedicta gloria Domini de loco suo
EZEK|3|13|et vocem alarum animalium percutientium alteram ad alteram et vocem rotarum sequentium animalia et vocem commotionis magnae
EZEK|3|14|spiritus quoque levavit me et adsumpsit me et abii amarus in indignatione spiritus mei manus enim Domini erat mecum confortans me
EZEK|3|15|et veni ad transmigrationem acervum novarum frugum ad eos qui habitabant iuxta flumen Chobar et sedi ubi illi sedebant et mansi ibi septem diebus maerens in medio eorum
EZEK|3|16|cum autem pertransissent septem dies factum est verbum Domini ad me dicens
EZEK|3|17|fili hominis speculatorem dedi te domui Israhel et audies de ore meo verbum et adnuntiabis eis ex me
EZEK|3|18|si dicente me ad impium morte morieris non adnuntiaveris ei neque locutus fueris ut avertatur a via sua impia et vivat ipse impius in iniquitate sua morietur sanguinem autem eius de manu tua requiram
EZEK|3|19|si autem tu adnuntiaveris impio et ille non fuerit conversus ab impietate sua et via sua impia ipse quidem in iniquitate sua morietur tu autem animam tuam liberasti
EZEK|3|20|sed et si conversus iustus a iustitia sua fecerit iniquitatem ponam offendiculum coram eo ipse morietur quia non adnuntiasti ei in peccato suo morietur et non erunt in memoria iustitiae eius quas fecit sanguinem vero eius de manu tua requiram
EZEK|3|21|si autem tu adnuntiaveris iusto ut non peccet iustus et ille non peccaverit vivens vivet quia adnuntiasti ei et tu animam tuam liberasti
EZEK|3|22|et facta est super me manus Domini et dixit ad me surgens egredere in campum et ibi loquar tecum
EZEK|3|23|et surgens egressus sum in campum et ecce ibi gloria Domini stabat quasi gloria quam vidi iuxta fluvium Chobar et cecidi in faciem meam
EZEK|3|24|et ingressus est in me spiritus et statuit me super pedes meos et locutus est mihi et dixit ad me ingredere et includere in medio domus tuae
EZEK|3|25|et tu fili hominis ecce data sunt super te vincula et ligabunt te in eis et non egredieris in medio eorum
EZEK|3|26|et linguam tuam adherescere faciam palato tuo et eris mutus nec quasi vir obiurgans quia domus exasperans est
EZEK|3|27|cum autem locutus fuero tibi aperiam os tuum et dices ad eos haec dicit Dominus Deus qui audit audiat et qui quiescit quiescat quia domus exasperans est
EZEK|4|1|et tu fili hominis sume tibi laterem et pones eum coram te et describes in eo civitatem Hierusalem
EZEK|4|2|et ordinabis adversus eam obsidionem et aedificabis munitiones et conportabis aggerem et dabis contra eam castra et pones arietes in gyro
EZEK|4|3|et tu sume tibi sartaginem ferream et pones eam murum ferreum inter te et inter civitatem et obfirmabis faciem tuam ad eam et erit in obsidionem et circumdabis eam signum est domui Israhel
EZEK|4|4|et tu dormies super latus tuum sinistrum et pones iniquitates domus Israhel super eo numero dierum quibus dormies super illud et adsumes iniquitatem eorum
EZEK|4|5|ego autem dedi tibi annos iniquitatis eorum numero dierum trecentos et nonaginta dies et portabis iniquitatem domus Israhel
EZEK|4|6|et cum conpleveris haec dormies super latus tuum dextrum secundo et adsumes iniquitatem domus Iuda quadraginta diebus diem pro anno diem inquam pro anno dedi tibi
EZEK|4|7|et ad obsidionem Hierusalem convertes faciem tuam et brachium tuum erit exertum et prophetabis adversus eam
EZEK|4|8|ecce circumdedi te vinculis et non te convertes a latere tuo in latus aliud donec conpleas dies obsidionis tuae
EZEK|4|9|et tu sume tibi frumentum et hordeum et fabam et lentem et milium et viciam et mittes ea in vas unum et facies tibi panes numero dierum quibus dormies super latus tuum trecentis et nonaginta diebus comedes illud
EZEK|4|10|cibus autem tuus quo vesceris erit in pondere viginti stateres in die a tempore usque ad tempus comedes illud
EZEK|4|11|et aquam in mensura bibes sextam partem hin a tempore usque ad tempus bibes illud
EZEK|4|12|et quasi subcinericium hordiacium comedes illud et stercore quod egredietur de homine operies illud in oculis eorum
EZEK|4|13|et dixit Dominus sic comedent filii Israhel panem suum pollutum inter gentes ad quas eiciam eos
EZEK|4|14|et dixi ha ha ha Domine Deus ecce anima mea non est polluta et morticinum et laceratum a bestiis non comedi ab infantia mea usque nunc et non est ingressa os meum omnis caro inmunda
EZEK|4|15|et dixit ad me ecce dedi tibi fimum boum pro stercoribus humanis et facies panem tuum in eo
EZEK|4|16|et dixit ad me fili hominis ecce ego conteram baculum panis in Hierusalem et comedent panem in pondere et in sollicitudine et aquam in mensura et in angustia bibent
EZEK|4|17|ut deficientibus pane et aqua corruat unusquisque ad fratrem suum et contabescant in iniquitatibus suis
EZEK|5|1|et tu fili hominis sume tibi gladium acutum radentem pilos adsumes eum et duces per caput tuum et per barbam tuam et adsumes tibi stateram ponderis et divides eos
EZEK|5|2|tertiam partem igni conbures in medio civitatis iuxta conpletionem dierum obsidionis et adsumens tertiam partem concides gladio in circuitu eius tertiam vero aliam disperges in ventum et gladium nudabo post eos
EZEK|5|3|et sumes inde parvum numerum et ligabis eos in summitate pallii tui
EZEK|5|4|et ex eis rursum tolles et proicies in medio ignis et conbures eos igni ex eo egredietur ignis in omnem domum Israhel
EZEK|5|5|haec dicit Dominus Deus ista est Hierusalem in medio gentium posui eam et in circuitu eius terras
EZEK|5|6|et contempsit iudicia mea ut plus esset impia quam gentes et praecepta mea ultra quam terrae quae in circuitu eius sunt iudicia enim mea proiecerunt et in praeceptis meis non ambulaverunt
EZEK|5|7|idcirco haec dicit Dominus Deus quia superastis gentes quae in circuitu vestro sunt in praeceptis meis non ambulastis et iudicia mea non fecistis et iuxta iudicia gentium quae in circuitu vestro sunt non estis operati
EZEK|5|8|ideo haec dicit Dominus Deus ecce ego ad te et ipse ego faciam in medio tui iudicia in oculis gentium
EZEK|5|9|et faciam in te quae non feci et quibus similia ultra non faciam propter omnes abominationes tuas
EZEK|5|10|ideo patres comedent filios in medio tui et filii comedent patres suos et faciam in te iudicia et ventilabo universas reliquias tuas in omnem ventum
EZEK|5|11|idcirco vivo ego dicit Dominus Deus nisi pro eo quod sanctum meum violasti in omnibus offensionibus tuis et in omnibus abominationibus tuis ego quoque confringam et non parcet oculus meus et non miserebor
EZEK|5|12|tertia tui pars peste morietur et fame consumetur in medio tui et tertia tui pars gladio cadet in circuitu tuo tertiam vero partem tuam in omnem ventum dispergam et gladium evaginabo post eos
EZEK|5|13|et conpleam furorem meum et requiescere faciam indignationem meam in eis et consolabor et scient quia ego Dominus locutus sum in zelo meo cum implevero indignationem meam in eis
EZEK|5|14|et dabo te in desertum et in obprobrium in gentibus quae in circuitu tuo sunt in conspectu omnis praetereuntis
EZEK|5|15|et eris obprobrium et blasphemia exemplum et stupor in gentibus quae in circuitu tuo sunt cum fecero in te iudicia in furore et in indignatione et in increpationibus irae
EZEK|5|16|ego Dominus locutus sum quando misero sagittas famis pessimas in eos quae erunt mortiferae et quas mittam ut disperdam vos et famem congregabo super vos et conteram vobis baculum panis
EZEK|5|17|et inmittam in vos famem et bestias pessimas usque ad internicionem et pestilentia et sanguis transibunt per te et gladium inducam super te ego Dominus locutus sum
EZEK|6|1|et factus est sermo Domini ad me dicens
EZEK|6|2|fili hominis pone faciem tuam ad montes Israhel et prophetabis ad eos
EZEK|6|3|et dices montes Israhel audite verbum Domini Dei haec dicit Dominus Deus montibus et collibus rupibus et vallibus ecce ego inducam super vos gladium et disperdam excelsa vestra
EZEK|6|4|et demoliar aras vestras et confringentur simulacra vestra et deiciam interfectos vestros ante idola vestra
EZEK|6|5|et dabo cadavera filiorum Israhel ante faciem simulacrorum vestrorum et dispergam ossa vestra circum aras vestras
EZEK|6|6|in omnibus habitationibus vestris urbes desertae erunt et excelsa demolientur et dissipabuntur et interibunt arae vestrae et confringentur et cessabunt idola vestra et conterentur delubra vestra et delebuntur opera vestra
EZEK|6|7|et cadet interfectus in medio vestri et scietis quoniam ego Dominus
EZEK|6|8|et relinquam in vobis eos qui fugerint gladium in gentibus cum dispersero vos in terris
EZEK|6|9|et recordabuntur mei liberati vestri in gentibus ad quas captivi ducti sunt quia contrivi cor eorum fornicans et recedens a me et oculos eorum fornicantes post idola sua et displicebunt sibimet super malis quae fecerunt in universis abominationibus suis
EZEK|6|10|et scient quia ego Dominus non frustra locutus sum ut facerem eis malum hoc
EZEK|6|11|haec dicit Dominus Deus percute manu tua et adlide pedem tuum et dic eheu ad omnes abominationes malorum domus Israhel qui gladio fame peste ruituri sunt
EZEK|6|12|qui longe est peste morietur qui autem prope gladio corruet et qui relictus fuerit et obsessus fame morietur et conpleam indignationem meam in eis
EZEK|6|13|et scietis quia ego Dominus cum fuerint interfecti vestri in medio idolorum vestrorum in circuitu ararum vestrarum in omni colle excelso in cunctis summitatibus montium et subtus omne lignum nemorosum et subtus universam quercum frondosam locum ubi accenderunt tura redolentia universis idolis suis
EZEK|6|14|et extendam manum meam super eos et faciam terram desolatam et destitutam a deserto Deblatha in omnibus habitationibus eorum et scient quia ego Dominus
EZEK|7|1|et factus est sermo Domini ad me dicens
EZEK|7|2|et tu fili hominis haec dicit Dominus Deus terrae Israhel finis venit finis super quattuor plagas terrae
EZEK|7|3|nunc finis super te et emittam furorem meum in te et iudicabo te iuxta vias tuas et ponam contra te omnes abominationes tuas
EZEK|7|4|et non parcet oculus meus super te et non miserebor sed vias tuas ponam super te et abominationes tuae in medio tui erunt et scietis quia ego Dominus
EZEK|7|5|haec dicit Dominus Deus adflictio una adflictio ecce venit
EZEK|7|6|finis venit venit finis evigilavit adversum te ecce venit
EZEK|7|7|venit contractio super te qui habitas in terra venit tempus prope est dies occisionis et non gloriae montium
EZEK|7|8|nunc de propinquo effundam iram meam super te et conpleam furorem meum in te et iudicabo te iuxta vias tuas et inponam tibi omnia scelera tua
EZEK|7|9|et non parcet oculus meus neque miserebor sed vias tuas inponam tibi et abominationes tuae in medio tui erunt et scietis quia ego sum Dominus percutiens
EZEK|7|10|ecce dies ecce venit egressa est contractio floruit virga germinavit superbia
EZEK|7|11|iniquitas surrexit in virga impietatis non ex eis et non ex populo neque ex sonitu eorum et non erit requies in eis
EZEK|7|12|venit tempus adpropinquavit dies qui emit non laetetur et qui vendit non lugeat quia ira super omnem populum eius
EZEK|7|13|quia qui vendit ad id quod vendidit non revertetur et adhuc in viventibus vita eorum visio enim ad omnem multitudinem eius non regredietur et vir in iniquitate vitae suae non confortabitur
EZEK|7|14|canite tuba praeparentur omnes et non est qui vadat ad proelium ira enim mea super universum populum eius
EZEK|7|15|gladius foris pestis et fames intrinsecus qui in agro est gladio morietur et qui in civitate pestilentia et fame devorabuntur
EZEK|7|16|et salvabuntur qui fugerint ex eis et erunt in montibus quasi columbae convallium omnes trepidi unusquisque in iniquitate sua
EZEK|7|17|omnes manus dissolventur et omnia genua fluent aquis
EZEK|7|18|et accingent se ciliciis et operiet eos formido et in omni facie confusio et in universis capitibus eorum calvitium
EZEK|7|19|argentum eorum foris proicietur et aurum eorum in sterquilinium erit argentum eorum et aurum eorum non valebit liberare eos in die furoris Domini animam suam non saturabunt et ventres eorum non implebuntur quia scandalum iniquitatis eorum factum est
EZEK|7|20|et ornamentum monilium suorum in superbiam posuerunt et imagines abominationum suarum et simulacrorum fecerunt ex eo propter hoc dedi eis illud in inmunditiam
EZEK|7|21|et dabo illud in manus alienorum ad diripiendum et impiis terrae in praedam et contaminabunt illud
EZEK|7|22|et avertam faciem meam ab eis et violabunt arcanum meum et introibunt in illud emissarii et contaminabunt illud
EZEK|7|23|fac conclusionem quoniam terra plena est iudicio sanguinum et civitas plena iniquitate
EZEK|7|24|et adducam pessimos de gentibus et possidebunt domos eorum et quiescere faciam superbiam potentium et possidebunt sanctuaria eorum
EZEK|7|25|angustia superveniente requirent pacem et non erit
EZEK|7|26|conturbatio super conturbationem veniet et auditus super auditum et quaerent visionem de propheta et lex peribit a sacerdote et consilium a senioribus
EZEK|7|27|rex lugebit et princeps induetur maerore et manus populi terrae conturbabuntur secundum viam eorum faciam eis et secundum iudicia eorum iudicabo eos et scient quia ego Dominus
EZEK|8|1|et factum est in anno sexto in sexto mense in quinta mensis ego sedebam in domo mea et senes Iuda sedebant coram me et cecidit super me ibi manus Domini Dei
EZEK|8|2|et vidi et ecce similitudo quasi aspectus ignis ab aspectu lumborum eius et deorsum ignis et a lumbis eius et sursum quasi aspectus splendoris ut visio electri
EZEK|8|3|et emissa similitudo manus adprehendit me in cincinno capitis mei et elevavit me spiritus inter terram et caelum et adduxit in Hierusalem in visione Dei iuxta ostium interius quod respiciebat aquilonem ubi erat statutum idolum zeli ad provocandam aemulationem
EZEK|8|4|et ecce ibi gloria Dei Israhel secundum visionem quam videram in campo
EZEK|8|5|et dixit ad me fili hominis leva oculos tuos ad viam aquilonis et levavi oculos meos ad viam aquilonis et ecce ab aquilone portae altaris idolum zeli in ipso introitu
EZEK|8|6|et dixit ad me fili hominis putasne vides tu quid isti faciant abominationes magnas quas domus Israhel facit hic ut procul recedam a sanctuario meo et adhuc conversus videbis abominationes maiores
EZEK|8|7|et introduxit me ad ostium atrii et vidi et ecce foramen unum in pariete
EZEK|8|8|et dixit ad me fili hominis fode parietem et cum perfodissem parietem apparuit ostium unum
EZEK|8|9|et dixit ad me ingredere et vide abominationes pessimas quas isti faciunt hic
EZEK|8|10|et ingressus vidi et ecce omnis similitudo reptilium et animalium abominatio et universa idola domus Israhel depicta erant in pariete in circuitu per totum
EZEK|8|11|et septuaginta viri de senioribus domus Israhel et Hiezonias filius Saphan stabat in medio eorum stantium ante picturas et unusquisque habebat turibulum in manu sua et vapor nebulae de ture consurgebat
EZEK|8|12|et dixit ad me certe vides fili hominis quae seniores domus Israhel faciunt in tenebris unusquisque in abscondito cubiculi sui dicunt enim non videt Dominus nos dereliquit Dominus terram
EZEK|8|13|et dixit ad me adhuc conversus videbis abominationes maiores quas isti faciunt
EZEK|8|14|et introduxit me per ostium portae domus Domini quod respiciebat ad aquilonem et ecce ibi mulieres sedebant plangentes Adonidem
EZEK|8|15|et dixit ad me certe vidisti fili hominis adhuc conversus videbis abominationes maiores his
EZEK|8|16|et introduxit me in atrium domus Domini interius et ecce in ostio templi Domini inter vestibulum et altare quasi viginti quinque viri dorsa habentes contra templum Domini et facies ad orientem et adorabant ad ortum solis
EZEK|8|17|et dixit ad me certe vidisti fili hominis numquid leve est hoc domui Iuda ut facerent abominationes istas quas fecerunt hic quia replentes terram iniquitate conversi sunt ad inritandum me et ecce adplicant ramum ad nares suas
EZEK|8|18|ergo et ego faciam in furore non parcet oculus meus nec miserebor et cum clamaverint ad aures meas voce magna non exaudiam eos
EZEK|9|1|et clamavit in auribus meis voce magna dicens adpropinquaverunt visitationes urbis et unusquisque vas interfectionis habet in manu sua
EZEK|9|2|et ecce sex viri veniebant de via portae superioris quae respicit ad aquilonem et uniuscuiusque vas interitus in manu eius vir quoque unus in medio eorum vestitus lineis et atramentarium scriptoris ad renes eius et ingressi sunt et steterunt iuxta altare aereum
EZEK|9|3|et gloria Domini Israhel adsumpta est de cherub quae erat super eum ad limen domus et vocavit virum qui indutus erat lineis et atramentarium scriptoris habebat in lumbis suis
EZEK|9|4|et dixit Dominus ad eum transi per mediam civitatem in medio Hierusalem et signa thau super frontes virorum gementium et dolentium super cunctis abominationibus quae fiunt in medio eius
EZEK|9|5|et illis dixit audiente me transite per civitatem sequentes eum et percutite non parcat oculus vester neque misereamini
EZEK|9|6|senem adulescentulum et virginem parvulum et mulieres interficite usque ad internicionem omnem autem super quem videritis thau ne occidatis et a sanctuario meo incipite coeperunt ergo a viris senioribus qui erant ante faciem domus
EZEK|9|7|et dixit ad eos contaminate domum et implete atria interfectis egredimini et egressi sunt et percutiebant eos qui erant in civitate
EZEK|9|8|et caede conpleta remansi ego ruique super faciem meam et clamans aio heu heu heu Domine Deus ergone disperdes omnes reliquias Israhel effundens furorem tuum super Hierusalem
EZEK|9|9|et dixit ad me iniquitas domus Israhel et Iuda magna est nimis valde et repleta est terra sanguinibus et civitas repleta est aversione dixerunt enim dereliquit Dominus terram et Dominus non videt
EZEK|9|10|igitur et meus non parcet oculus neque miserebor viam eorum super caput eorum reddam
EZEK|9|11|et ecce vir qui indutus erat lineis qui habebat atramentarium in dorso suo respondit verbum dicens feci sicut praecepisti mihi
EZEK|10|1|et vidi et ecce in firmamento quod erat super caput cherubin quasi lapis sapphyrus quasi species similitudinis solii apparuit super ea
EZEK|10|2|et dixit ad virum qui indutus erat lineis et ait ingredere in medio rotarum quae sunt subtus cherub et imple manum tuam prunis ignis quae sunt inter cherubin et effunde super civitatem ingressusque est in conspectu meo
EZEK|10|3|cherubin autem stabant a dextris domus cum ingrederetur vir et nubes implevit atrium interius
EZEK|10|4|et elevata est gloria Domini desuper cherub ad limen domus et repleta est domus nube et atrium repletum est splendore gloriae Domini
EZEK|10|5|et sonitus alarum cherubin audiebatur usque ad atrium exterius quasi vox Dei omnipotentis loquentis
EZEK|10|6|cumque praecepisset viro qui indutus erat lineis dicens sume ignem de medio rotarum quae sunt inter cherubin ingressus ille stetit iuxta rotam
EZEK|10|7|et extendit cherub manum de medio cherubin ad ignem qui erat inter cherubin et sumpsit et dedit in manus eius qui indutus erat lineis qui accipiens egressus est
EZEK|10|8|et apparuit in cherubin similitudo manus hominis subtus pinnas eorum
EZEK|10|9|et vidi et ecce quattuor rotae iuxta cherubin rota una iuxta cherub unum et rota alia iuxta cherub unum species autem erat rotarum quasi visio lapidis chrysoliti
EZEK|10|10|et aspectus earum similitudo una quattuor quasi sit rota in medio rotae
EZEK|10|11|cumque ambularent in quattuor partes gradiebantur non revertebantur ambulantes sed ad locum ad quem ire declinabat quae prima erat sequebantur et ceterae nec convertebantur
EZEK|10|12|et omne corpus earum et colla et manus et pinnae et circuli plena erant oculis in circuitu quattuor rotarum
EZEK|10|13|et rotas istas vocavit volubiles audiente me
EZEK|10|14|quattuor autem facies habebat unum facies una facies cherub et facies secunda facies hominis et in tertio facies leonis et in quarto facies aquilae
EZEK|10|15|et elevata sunt cherubin ipsum est animal quod videram iuxta flumen Chobar
EZEK|10|16|cumque ambularent cherubin ibant pariter et rotae iuxta ea et cum levarent cherubin alas suas ut exaltarentur de terra non residebant rotae sed et ipsae iuxta erant
EZEK|10|17|stantibus illis stabant et cum elevatis elevabantur spiritus enim vitae erat in eis
EZEK|10|18|et egressa est gloria Domini a limine templi et stetit super cherubin
EZEK|10|19|et elevantia cherubin alas suas exaltata sunt a terra coram me et illis egredientibus rotae quoque subsecutae sunt et stetit in introitu portae domus Domini orientalis et gloria Dei Israhel erat super ea
EZEK|10|20|ipsum est animal quod vidi subter Deum Israhel iuxta fluvium Chobar et intellexi quia cherubin essent
EZEK|10|21|quattuor per quattuor vultus uni et quattuor alae uni et similitudo manus hominis sub alis eorum
EZEK|10|22|et similitudo vultuum eorum ipsi vultus quos videram iuxta fluvium Chobar et intuitus eorum et impetus singulorum ante faciem suam ingredi
EZEK|11|1|et elevavit me spiritus et introduxit me ad portam domus Domini orientalem quae respicit solis ortum et ecce in introitu portae viginti quinque viri et vidi in medio eorum Hiezoniam filium Azur et Pheltiam filium Banaiae principes populi
EZEK|11|2|dixitque ad me fili hominis hii viri qui cogitant iniquitatem et tractant consilium pessimum in urbe ista
EZEK|11|3|dicentes nonne dudum aedificatae sunt domus haec est lebes nos autem carnes
EZEK|11|4|idcirco vaticinare de eis vaticinare fili hominis
EZEK|11|5|et inruit in me spiritus Domini et dixit ad me loquere haec dicit Dominus sic locuti estis domus Israhel et cogitationes cordis vestri ego novi
EZEK|11|6|plurimos occidistis in urbe hac et implestis vias eius interfectis
EZEK|11|7|propterea haec dicit Dominus Deus interfecti vestri quos posuistis in medio eius hii sunt carnes et haec est lebes et educam vos de medio eius
EZEK|11|8|gladium metuistis et gladium inducam super vos ait Dominus Deus
EZEK|11|9|et eiciam vos de medio eius daboque vos in manu hostium et faciam in vobis iudicia
EZEK|11|10|gladio cadetis in finibus Israhel iudicabo vos et scietis quia ego Dominus
EZEK|11|11|haec non erit vobis in lebetem et vos non eritis in medio eius in carnes in finibus Israhel iudicabo vos
EZEK|11|12|et scietis quia ego Dominus qui in praeceptis meis non ambulastis et iudicia mea non fecistis sed iuxta iudicia gentium quae in circuitu vestro sunt estis operati
EZEK|11|13|et factum est cum prophetarem Pheltias filius Banaiae mortuus est et cecidi in faciem meam clamans voce magna et dixi heu heu heu Domine Deus consummationem tu facis reliquiarum Israhel
EZEK|11|14|et factum est verbum Domini ad me dicens
EZEK|11|15|fili hominis fratres tui fratres tui viri propinqui tui et omnis domus Israhel universi quibus dixerunt habitatores Hierusalem longe recedite a Domino nobis data est terra in possessionem
EZEK|11|16|propterea haec dicit Dominus Deus quia longe feci eos in gentibus et quia dispersi eos in terris ero eis in sanctificationem modicam in terris ad quas venerunt
EZEK|11|17|propterea loquere haec dicit Dominus Deus congregabo vos de populis et adunabo de terris in quibus dispersi estis daboque vobis humum Israhel
EZEK|11|18|et ingredientur illuc et auferent omnes offensiones cunctasque abominationes eius de illa
EZEK|11|19|et dabo eis cor unum et spiritum novum tribuam in visceribus eorum et auferam cor lapideum de carne eorum et dabo eis cor carneum
EZEK|11|20|ut in praeceptis meis ambulent et iudicia mea custodiant faciantque ea et sint mihi in populum et ego sim eis in Deum
EZEK|11|21|quorum cor post offendicula et abominationes suas ambulat horum viam in capite suo ponam dicit Dominus Deus
EZEK|11|22|et elevaverunt cherubin alas suas et rotae cum eis et gloria Dei Israhel erat super ea
EZEK|11|23|et ascendit gloria Domini de medio civitatis stetitque super montem qui est ad orientem urbis
EZEK|11|24|et spiritus levavit me adduxitque in Chaldeam ad transmigrationem in visione in spiritu Dei et sublata est a me visio quam videram
EZEK|11|25|et locutus sum ad transmigrationem omnia verba Domini quae ostenderat mihi
EZEK|12|1|et factus est sermo Domini ad me dicens
EZEK|12|2|fili hominis in medio domus exasperantis tu habitas qui oculos habent ad videndum et non vident et aures ad audiendum et non audiunt quia domus exasperans est
EZEK|12|3|tu ergo fili hominis fac tibi vasa transmigrationis et transmigrabis per diem coram eis transmigrabis autem de loco tuo ad locum alterum in conspectu eorum si forte aspiciant quia domus exasperans est
EZEK|12|4|et efferes foras vasa tua quasi vasa transmigrantis per diem in conspectu eorum tu autem egredieris vespere coram eis sicut egreditur migrans
EZEK|12|5|ante oculos eorum perfodi tibi parietem et egredieris per eum
EZEK|12|6|in conspectu eorum in umeris portaberis in caligine effereris faciem tuam velabis et non videbis terram quia portentum dedi te domui Israhel
EZEK|12|7|feci ergo sicut praeceperat mihi vasa mea protuli quasi vasa transmigrantis per diem et vespere perfodi mihi parietem manu in caligine egressus sum et in umeris portatus in conspectu eorum
EZEK|12|8|et factus est sermo Domini ad me mane dicens
EZEK|12|9|fili hominis numquid non dixerunt ad te domus Israhel domus exasperans quid tu facis
EZEK|12|10|dic ad eos haec dicit Dominus Deus super ducem onus istud qui est in Hierusalem et super omnem domum Israhel quae est in medio eorum
EZEK|12|11|dic ego portentum vestrum quomodo feci sic fiet illis in transmigrationem et captivitatem ibunt
EZEK|12|12|et dux qui est in medio eorum in umeris portabitur in caligine egredietur parietem perfodient ut educant eum facies eius operietur ut non videat oculo terram
EZEK|12|13|et extendam rete meum super illum et capietur in sagena mea et adducam eum in Babylonem in terram Chaldeorum et ipsam non videbit ibique morietur
EZEK|12|14|et omnes qui circa eum sunt praesidium eius et agmina eius dispergam in omnem ventum et gladium evaginabo post eos
EZEK|12|15|et scient quia ego Dominus quando dispersero illos in gentibus et disseminavero eos in terris
EZEK|12|16|et relinquam ex eis viros paucos a gladio et fame et pestilentia ut narrent omnia scelera eorum in gentibus ad quas ingredientur et scient quia ego Dominus
EZEK|12|17|et factus est sermo Domini ad me dicens
EZEK|12|18|fili hominis panem tuum in conturbatione comede sed et aquam tuam in festinatione et maerore bibe
EZEK|12|19|et dices ad populum terrae haec dicit Dominus Deus ad eos qui habitant in Hierusalem in terra Israhel panem suum in sollicitudine comedent et aquam suam in desolatione bibent ut desoletur terra a multitudine sua propter iniquitatem omnium qui habitant in ea
EZEK|12|20|et civitates quae nunc habitantur desolatae erunt terraque deserta et scietis quia ego Dominus
EZEK|12|21|et factus est sermo Domini ad me dicens
EZEK|12|22|fili hominis quod est proverbium istud vobis in terra Israhel dicentium in longum differentur dies et peribit omnis visio
EZEK|12|23|ideo dic ad eos haec dicit Dominus Deus quiescere faciam proverbium istud neque vulgo dicetur ultra in Israhel et loquere ad eos quod adpropinquaverint dies et sermo omnis visionis
EZEK|12|24|non enim erit ultra omnis visio cassa neque divinatio ambigua in medio filiorum Israhel
EZEK|12|25|quia ego Dominus loquar quodcumque locutus fuero verbum et fiet non prolongabitur amplius sed in diebus vestris domus exasperans loquar verbum et faciam illud dicit Dominus Deus
EZEK|12|26|et factus est sermo Domini ad me dicens
EZEK|12|27|fili hominis ecce domus Israhel dicentium visio quam hic videt in dies multos et in tempora longa iste prophetat
EZEK|12|28|propterea dic ad eos haec dicit Dominus Deus non prolongabitur ultra omnis sermo meus verbum quod locutus fuero conplebitur dicit Dominus Deus
EZEK|13|1|et factus est sermo Domini ad me dicens
EZEK|13|2|fili hominis vaticinare ad prophetas Israhel qui prophetant et dices prophetantibus de corde suo audite verbum Domini
EZEK|13|3|haec dicit Dominus Deus vae prophetis insipientibus qui sequuntur spiritum suum et nihil vident
EZEK|13|4|quasi vulpes in desertis prophetae tui Israhel erant
EZEK|13|5|non ascendistis ex adverso neque opposuistis murum pro domo Israhel ut staretis in proelio in die Domini
EZEK|13|6|vident vana et divinant mendacium dicentes ait Dominus cum Dominus non miserit eos et perseveraverunt confirmare sermonem
EZEK|13|7|numquid non visionem cassam vidistis et divinationem mendacem locuti estis et dicitis ait Dominus cum ego non sim locutus
EZEK|13|8|propterea haec dicit Dominus Deus quia locuti estis vana et vidistis mendacium ideo ecce ego ad vos ait Dominus Deus
EZEK|13|9|et erit manus mea super prophetas qui vident vana et divinant mendacium in concilio populi mei non erunt et in scriptura domus Israhel non scribentur nec in terra Israhel ingredientur et scietis quia ego Dominus Deus
EZEK|13|10|eo quod deceperint populum meum dicentes pax et non est pax et ipse aedificabat parietem illi autem liniebant eum luto absque paleis
EZEK|13|11|dic ad eos qui liniunt absque temperatura quod casurus sit erit enim imber inundans et dabo lapides praegrandes desuper inruentes et ventum procellae dissipantem
EZEK|13|12|siquidem ecce cecidit paries numquid non dicetur vobis ubi est litura quam levistis
EZEK|13|13|propterea haec dicit Dominus Deus et erumpere faciam spiritum tempestatum in indignatione mea et imber inundans in furore meo erit et lapides grandes in ira in consummationem
EZEK|13|14|et destruam parietem quem levistis absque temperamento et adaequabo eum terrae et revelabitur fundamentum eius et cadet et consumetur in medio eius et scietis quia ego sum Dominus
EZEK|13|15|et conplebo indignationem meam in parietem et in his qui linunt eum absque temperamento dicamque vobis non est paries et non sunt qui linunt eum
EZEK|13|16|prophetae Israhel qui prophetant ad Hierusalem et vident ei visionem pacis et non est pax ait Dominus Deus
EZEK|13|17|et tu fili hominis pone faciem tuam contra filias populi tui quae prophetant de corde suo et vaticinare super eas
EZEK|13|18|et dic haec ait Dominus Deus vae quae consuunt pulvillos sub omni cubito manus et faciunt cervicalia sub capite universae aetatis ad capiendas animas cum caperent animas populi mei vivificabant animas eorum
EZEK|13|19|et violabant me ad populum meum propter pugillum hordei et fragmen panis ut interficerent animas quae non moriuntur et vivificarent animas quae non vivunt mentientes populo meo credenti mendaciis
EZEK|13|20|propter hoc haec dicit Dominus Deus ecce ego ad pulvillos vestros quibus vos capitis animas volantes et disrumpam eos de brachiis vestris et dimittam animas quas vos capitis animas ad volandum
EZEK|13|21|et disrumpam cervicalia vestra et liberabo populum meum de manu vestra neque erunt ultra in manibus vestris ad praedandum et scietis quia ego Dominus
EZEK|13|22|pro eo quod maerere fecistis cor iusti mendaciter quem ego non contristavi et confortastis manus impii ut non reverteretur a via sua mala et viveret
EZEK|13|23|propterea vana non videbitis et divinationes non divinabitis amplius et eruam populum meum de manu vestra et scietis quoniam ego Dominus
EZEK|14|1|et venerunt ad me viri seniorum Israhel et sederunt coram me
EZEK|14|2|et factus est sermo Domini ad me dicens
EZEK|14|3|fili hominis viri isti posuerunt inmunditias suas in cordibus suis et scandalum iniquitatis suae statuerunt contra faciem suam numquid interrogatus respondebo eis
EZEK|14|4|propter hoc loquere eis et dices ad eos haec dicit Dominus Deus homo homo de domo Israhel qui posuerit inmunditias suas in corde suo et scandalum iniquitatis suae statuerit contra faciem suam et venerit ad prophetam interrogans per eum me ego Dominus respondebo ei in multitudine inmunditiarum suarum
EZEK|14|5|ut capiatur domus Israhel in corde suo quo recesserunt a me in cunctis idolis suis
EZEK|14|6|propterea dic ad domum Israhel haec dicit Dominus Deus convertimini et recedite ab idolis vestris et ab universis contaminationibus vestris avertite facies vestras
EZEK|14|7|quia homo homo de domo Israhel et de proselytis quicumque advena fuerit in Israhel si alienatus fuerit a me et posuerit idola sua in corde suo et scandalum iniquitatis suae statuerit contra faciem suam et venerit ad prophetam ut interroget per eum me ego Dominus respondebo ei per me
EZEK|14|8|et ponam faciem meam super hominem illum et faciam eum in exemplum et in proverbium et disperdam eum de medio populi mei et scietis quia ego Dominus
EZEK|14|9|et propheta cum erraverit et locutus fuerit verbum ego Dominus decepi prophetam illum et extendam manum meam super eum et delebo eum de medio populi mei Israhel
EZEK|14|10|et portabunt iniquitatem suam iuxta iniquitatem interrogantis sic iniquitas prophetae erit
EZEK|14|11|ut non erret ultra domus Israhel a me neque polluatur in universis praevaricationibus suis sed sit mihi in populum et ego sim eis in Deum ait Dominus exercituum
EZEK|14|12|et factus est sermo Domini ad me dicens
EZEK|14|13|fili hominis terra cum peccaverit mihi ut praevaricetur praevaricans extendam manum meam super eam et conteram virgam panis eius et inmittam in eam famem et interficiam de ea hominem et iumentum
EZEK|14|14|et si fuerint tres viri isti in medio eius Noe Danihel et Iob ipsi iustitia sua liberabunt animas suas ait Dominus exercituum
EZEK|14|15|quod si et bestias pessimas induxero super terram ut vastem eam et fuerit invia eo quod non sit pertransiens propter bestias
EZEK|14|16|tres viri isti qui fuerint in ea vivo ego dicit Dominus Deus quia nec filios nec filias liberabunt sed ipsi soli liberabuntur terra autem desolabitur
EZEK|14|17|vel si gladium induxero super terram illam et dixero gladio transi per terram et interfecero de ea hominem et iumentum
EZEK|14|18|et tres viri isti fuerint in medio eius vivo ego dicit Dominus Deus non liberabunt filios neque filias sed ipsi soli liberabuntur
EZEK|14|19|si autem et pestilentiam inmisero super terram illam et effudero indignationem meam super eam in sanguine ut auferam ex ea hominem et iumentum
EZEK|14|20|et Noe et Danihel et Iob fuerint in medio eius vivo ego dicit Dominus Deus quia filium et filiam non liberabunt sed ipsi iustitia sua liberabunt animas suas
EZEK|14|21|quoniam haec dicit Dominus Deus quod si et quattuor iudicia mea pessima gladium et famem et bestias malas et pestilentiam misero in Hierusalem ut interficiam de ea hominem et pecus
EZEK|14|22|tamen relinquetur in ea salvatio educentium filios et filias ecce ipsi egredientur ad vos et videbitis viam eorum et adinventiones eorum et consolabimini super malo quod induxi in Hierusalem in omnibus quae inportavi super eam
EZEK|14|23|et consolabuntur vos cum videritis viam eorum et adinventiones eorum et cognoscetis quod non frustra fecerim omnia quae feci in ea ait Dominus Deus
EZEK|15|1|et factus est sermo Domini ad me dicens
EZEK|15|2|fili hominis quid fiet ligno vitis ex omnibus lignis nemorum quae sunt inter ligna silvarum
EZEK|15|3|numquid tolletur de ea lignum ut fiat opus aut fabricabitur de ea paxillus ut dependeat in eo quodcumque vas
EZEK|15|4|ecce igni datum est in escam utramque partem eius consumpsit ignis et medietas eius redacta est in favillam numquid utile erit ad opus
EZEK|15|5|etiam cum esset integrum non erat aptum ad opus quanto magis cum ignis illud devoraverit et conbuserit nihil ex eo fiet operis
EZEK|15|6|propterea haec dicit Dominus Deus quomodo lignum vitis inter ligna silvarum quod dedi igni ad devorandum sic tradidi habitatores Hierusalem
EZEK|15|7|et ponam faciem meam in eos de igne egredientur et ignis consumet eos et scietis quia ego Dominus cum posuero faciem meam in eos
EZEK|15|8|et dedero terram inviam et desolatam eo quod praevaricatores extiterint dicit Dominus Deus
EZEK|16|1|et factus est sermo Domini ad me dicens
EZEK|16|2|fili hominis notas fac Hierusalem abominationes suas
EZEK|16|3|et dices haec dicit Dominus Deus Hierusalem radix tua et generatio tua de terra chananea pater tuus Amorreus et mater tua Cetthea
EZEK|16|4|et quando nata es in die ortus tui non est praecisus umbilicus tuus et in aqua non es lota in salutem nec sale salita nec involuta pannis
EZEK|16|5|non pepercit super te oculus ut facerem tibi unum de his miseratus tui sed proiecta es super faciem terrae in abiectione animae tuae in die qua nata es
EZEK|16|6|transiens autem per te vidi te conculcari in sanguine tuo et dixi tibi cum esses in sanguine tuo vive dixi inquam tibi in sanguine tuo vive
EZEK|16|7|multiplicatam quasi germen agri dedi te et multiplicata es et grandis effecta et ingressa es et pervenisti ad mundum muliebrem ubera tua intumuerunt et pilus tuus germinavit et eras nuda et confusionis plena
EZEK|16|8|et transivi per te et vidi te et ecce tempus tuum tempus amantium et expandi amictum meum super te et operui ignominiam tuam et iuravi tibi et ingressus sum pactum tecum ait Dominus Deus et facta es mihi
EZEK|16|9|et lavi te aqua et emundavi sanguinem tuum ex te et unxi te oleo
EZEK|16|10|et vestivi te discoloribus et calciavi te ianthino et cinxi te bysso et indui te subtilibus
EZEK|16|11|et ornavi te ornamento et dedi armillas in manibus tuis et torquem circa collum tuum
EZEK|16|12|et dedi inaurem super os tuum et circulos auribus tuis et coronam decoris in capite tuo
EZEK|16|13|et ornata es auro et argento et vestita es bysso et polymito et multicoloribus similam et mel et oleum comedisti et decora facta es vehementer nimis et profecisti in regnum
EZEK|16|14|et egressum est nomen tuum in gentes propter speciem tuam quia perfecta eras in decore meo quem posueram super te dicit Dominus Deus
EZEK|16|15|et habens fiduciam in pulchritudine tua fornicata es in nomine tuo et exposuisti fornicationem tuam omni transeunti ut eius fieres
EZEK|16|16|et sumens de vestimentis meis fecisti tibi excelsa hinc inde consuta et fornicata es super eis sicut non est factum neque futurum est
EZEK|16|17|et tulisti vasa decoris tui de auro meo et argento meo quae dedi tibi et fecisti tibi imagines masculinas et fornicata es in eis
EZEK|16|18|et sumpsisti vestimenta tua multicoloria et vestita es eis et oleum meum et thymiama meum posuisti coram eis
EZEK|16|19|et panem meum quem dedi tibi similam et oleum et mel quibus enutrivi te posuisti in conspectu eorum in odorem suavitatis et factum est ait Dominus Deus
EZEK|16|20|et tulisti filios tuos et filias tuas quas generasti mihi et immolasti eis ad devorandum numquid parva est fornicatio tua
EZEK|16|21|immolantis filios meos et dedisti illos consecrans eis
EZEK|16|22|et post omnes abominationes tuas et fornicationes non es recordata dierum adulescentiae tuae quando eras nuda et confusione plena conculcata in sanguine tuo
EZEK|16|23|et accidit post omnem malitiam tuam vae vae tibi ait Dominus Deus
EZEK|16|24|et aedificasti tibi lupanar et fecisti tibi prostibulum in cunctis plateis
EZEK|16|25|ad omne caput viae aedificasti signum prostitutionis tuae et abominabilem fecisti decorem tuum et divisisti pedes tuos omni transeunti et multiplicasti fornicationes tuas
EZEK|16|26|et fornicata es cum filiis Aegypti vicinis tuis magnarum carnium et multiplicasti fornicationem tuam ad inritandum me
EZEK|16|27|ecce ego extendi manum meam super te et auferam ius tuum et dabo te in animam odientium te filiarum Palestinarum quae erubescunt in via tua scelerata
EZEK|16|28|et fornicata es in filiis Assyriorum eo quod necdum fueris expleta et postquam fornicata es nec sic es satiata
EZEK|16|29|et multiplicasti fornicationem tuam in terra Chanaan cum Chaldeis et nec sic satiata es
EZEK|16|30|in quo mundabo cor tuum ait Dominus Deus cum facias omnia haec opera mulieris meretricis et procacis
EZEK|16|31|quia fabricasti lupanar tuum in capite omnis viae et excelsum tuum fecisti in omni platea nec facta es quasi meretrix fastidio augens pretium
EZEK|16|32|sed quasi mulier adultera quae super virum suum inducit alienos
EZEK|16|33|omnibus meretricibus dantur mercedes tu autem dedisti mercedes cunctis amatoribus tuis et donabas eis ut intrarent ad te undique ad fornicandum tecum
EZEK|16|34|factumque in te est contra consuetudinem mulierum in fornicationibus tuis et post te non erit fornicatio in eo enim quod dedisti mercedes et mercedes non accepisti factum est in te contrarium
EZEK|16|35|propterea meretrix audi verbum Domini
EZEK|16|36|haec dicit Dominus Deus quia effusum est aes tuum et revelata est ignominia tua in fornicationibus tuis super amatores tuos et super idola abominationum tuarum in sanguine filiorum tuorum quos dedisti eis
EZEK|16|37|ecce ego congregabo omnes amatores tuos quibus commixta es et omnes quos dilexisti cum universis quos oderas et congregabo eos super te undique et nudabo ignominiam tuam coram eis et videbunt omnem turpitudinem tuam
EZEK|16|38|et iudicabo te iudiciis adulterarum et effundentium sanguinem et dabo te in sanguinem furoris et zeli
EZEK|16|39|et dabo te in manus eorum et destruent lupanar tuum et demolientur prostibulum tuum et denudabunt te vestimentis tuis et auferent vasa decoris tui et derelinquent te nudam plenamque ignominia
EZEK|16|40|et adducent super te multitudinem et lapidabunt te lapidibus et trucidabunt te gladiis suis
EZEK|16|41|et conburent domos tuas igni et facient in te iudicia in oculis mulierum plurimarum et desines fornicari et mercedes ultra non dabis
EZEK|16|42|et requiescet indignatio mea in te et auferetur zelus meus a te et quiescam nec irascar amplius
EZEK|16|43|eo quod non fueris recordata dierum adulescentiae tuae et provocasti me in omnibus his quapropter et ego vias tuas in capite tuo dedi ait Dominus Deus et non feci iuxta scelera tua in omnibus abominationibus tuis
EZEK|16|44|ecce omnis qui dicit vulgo proverbium in te adsumet illud dicens sicut mater ita et filia eius
EZEK|16|45|filia matris tuae es tu quae proiecit virum suum et filios suos et soror sororum tuarum tu quae proiecerunt viros suos et filios suos mater vestra Cetthea et pater vester Amorreus
EZEK|16|46|et soror tua maior Samaria ipsa et filiae eius quae habitat ad sinistram tuam soror autem tua minor te quae habitat a dextris tuis Sodoma et filiae eius
EZEK|16|47|sed nec in viis earum ambulasti neque secundum scelera earum fecisti pauxillum minus paene sceleratiora fecisti illis in omnibus viis tuis
EZEK|16|48|vivo ego dicit Dominus Deus quia non fecit Sodoma soror tua ipsa et filiae eius sicut fecisti tu et filiae tuae
EZEK|16|49|ecce haec fuit iniquitas Sodomae sororis tuae superbia saturitas panis et abundantia et otium ipsius et filiarum eius et manum egeno et pauperi non porrigebant
EZEK|16|50|et elevatae sunt et fecerunt abominationes coram me et abstuli eas sicut vidisti
EZEK|16|51|et Samaria dimidium peccatorum tuorum non peccavit sed vicisti eas sceleribus tuis et iustificasti sorores tuas in omnibus abominationibus tuis quas operata es
EZEK|16|52|ergo et tu porta confusionem tuam quae vicisti sorores tuas peccatis tuis sceleratius agens ab eis iustificatae sunt enim a te ergo et tu confundere et porta ignominiam tuam quae iustificasti sorores tuas
EZEK|16|53|et convertam restituens eas conversione Sodomorum cum filiabus suis et conversione Samariae et filiarum eius et convertam reversionem tuam in medio earum
EZEK|16|54|ut portes ignominiam tuam et confundaris in omnibus quae fecisti consolans eas
EZEK|16|55|et soror tua Sodoma et filiae eius revertentur ad antiquitatem suam et Samaria et filiae eius revertentur ad antiquitatem suam et tu et filiae tuae revertimini ad antiquitatem vestram
EZEK|16|56|non fuit autem Sodoma soror tua audita in ore tuo in die superbiae tuae
EZEK|16|57|antequam revelaretur malitia tua sicut hoc tempore in obprobrium filiarum Syriae et cunctarum in circuitu tuo filiarum Palestinarum quae ambiunt te per gyrum
EZEK|16|58|scelus tuum et ignominiam tuam tu portasti ait Dominus Deus
EZEK|16|59|quia haec dicit Dominus Deus et faciam tibi sicut dispexisti iuramentum ut irritum faceres pactum
EZEK|16|60|et recordabor ego pacti mei tecum in diebus adulescentiae tuae et suscitabo tibi pactum sempiternum
EZEK|16|61|et recordaberis viarum tuarum et confunderis cum receperis sorores tuas te maiores cum minoribus tuis et dabo eas tibi in filias sed non ex pacto tuo
EZEK|16|62|et suscitabo ego pactum meum tecum et scies quia ego Dominus
EZEK|16|63|ut recorderis et confundaris et non sit tibi ultra aperire os prae confusione tua cum placatus fuero tibi in omnibus quae fecisti ait Dominus Deus
EZEK|17|1|et factum est verbum Domini ad me dicens
EZEK|17|2|fili hominis propone enigma et narra parabolam ad domum Israhel
EZEK|17|3|et dices haec dicit Dominus Deus aquila grandis magnarum alarum longo membrorum ductu plena plumis et varietate venit ad Libanum et tulit medullam cedri
EZEK|17|4|summitatem frondium eius avellit et transportavit eam in terram Chanaan in urbem negotiatorum posuit illam
EZEK|17|5|et tulit de semente terrae et posuit illud in terra pro semine ut firmaret radicem super aquas multas in superficie posuit illud
EZEK|17|6|cumque germinasset crevit in vineam latiorem humili statura respicientibus ramis eius ad eam et radices eius sub illa erunt facta est ergo vinea et fructificavit in palmites et emisit propagines
EZEK|17|7|et facta est aquila altera grandis magnis alis multisque plumis et ecce vinea ista quasi mittens radices suas ad eam palmites suos extendit ad illam ut inrigaret eam de areolis germinis sui
EZEK|17|8|in terra bona super aquas multas plantata est ut faciat frondes et portet fructum et sit in vineam grandem
EZEK|17|9|dic haec dicit Dominus Deus ergone prosperabitur nonne radices eius evellet et fructum eius distringet et siccabit omnes palmites germinis eius et arescet et non in brachio grandi neque in populo multo ut evelleret eam radicitus
EZEK|17|10|ecce plantata est ergone prosperabitur nonne cum tetigerit eam ventus urens siccabitur et in areis germinis sui arescet
EZEK|17|11|et factum est verbum Domini ad me dicens
EZEK|17|12|dic ad domum exasperantem nescitis quid ista significent dic ecce venit rex Babylonis Hierusalem et adsumet regem et principes eius et adducet eos ad semet ipsum in Babylonem
EZEK|17|13|et tollet de semine regni ferietque cum eo foedus et accipiet ab eo iusiurandum sed et fortes terrae tollet
EZEK|17|14|ut sit regnum humile et non elevetur sed custodiat pactum eius et servet illud
EZEK|17|15|qui recedens ab eo misit nuntios ad Aegyptum ut daret sibi equos et populum multum numquid prosperabitur vel consequetur salutem qui fecit haec et qui dissolvit pactum numquid effugiet
EZEK|17|16|vivo ego dicit Dominus Deus quoniam in loco regis qui constituit eum regem cuius fecit irritum iuramentum et solvit pactum quod habebat cum eo in medio Babylonis morietur
EZEK|17|17|et non in exercitu grandi neque in populo multo faciet contra eum Pharao proelium in iactu aggeris et in extructione vallorum ut interficiat animas multas
EZEK|17|18|spreverat enim iuramentum ut solveret foedus et ecce dedit manum suam et cum omnia haec fecerit non effugiet
EZEK|17|19|propterea haec dicit Dominus Deus vivo ego quoniam iuramentum quod sprevit et foedus quod praevaricatus est ponam in caput eius
EZEK|17|20|et expandam super eum rete meum et conprehendetur sagena mea et adducam eum in Babylonem et iudicabo illum ibi in praevaricatione qua despexit me
EZEK|17|21|et omnes profugi eius cum universo agmine gladio cadent residui autem in omnem ventum dispergentur et scietis quia ego Dominus locutus sum
EZEK|17|22|haec dicit Dominus Deus et sumam ego de medulla cedri sublimis et ponam de vertice ramorum eius tenerum distringam et plantabo super montem excelsum et eminentem
EZEK|17|23|in monte sublimi Israhel plantabo illud et erumpet in germen et faciet fructum et erit in cedrum magnam et habitabunt sub eo omnes volucres universum volatile sub umbra frondium eius nidificabit
EZEK|17|24|et scient omnia ligna regionis quia ego Dominus humiliavi lignum sublime et exaltavi lignum humile et siccavi lignum viride et frondere feci lignum aridum ego Dominus locutus sum et feci
EZEK|18|1|et factus est sermo Domini ad me dicens
EZEK|18|2|quid est quod inter vos parabolam vertitis in proverbium istud in terra Israhel dicentes patres comederunt uvam acerbam et dentes filiorum obstupescunt
EZEK|18|3|vivo ego dicit Dominus Deus si erit vobis ultra parabola haec in proverbium in Israhel
EZEK|18|4|ecce omnes animae meae sunt ut anima patris ita et anima filii mea est anima quae peccaverit ipsa morietur
EZEK|18|5|et vir si fuerit iustus et fecerit iudicium et iustitiam
EZEK|18|6|in montibus non comederit et oculos suos non levaverit ad idola domus Israhel et uxorem proximi sui non violaverit et ad mulierem menstruatam non accesserit
EZEK|18|7|et hominem non contristaverit pignus debitori reddiderit per vim nihil rapuerit panem suum esurienti dederit et nudum operuerit vestimento
EZEK|18|8|ad usuram non commodaverit et amplius non acceperit ab iniquitate averterit manum suam iudicium verum fecerit inter virum et virum
EZEK|18|9|in praeceptis meis ambulaverit et iudicia mea custodierit ut faciat veritatem hic iustus est vita vivet ait Dominus Deus
EZEK|18|10|quod si genuerit filium latronem effundentem sanguinem et fecerit unum de istis
EZEK|18|11|et haec quidem omnia non facientem sed in montibus comedentem et uxorem proximi sui polluentem
EZEK|18|12|egenum et pauperem contristantem rapientem rapinas pignus non reddentem et ad idola levantem oculos suos abominationem facientem
EZEK|18|13|ad usuram dantem et amplius accipientem numquid vivet non vivet cum universa detestanda haec fecerit morte morietur sanguis eius in ipso erit
EZEK|18|14|quod si genuerit filium qui videns omnia peccata patris sui quae fecit timuerit et non fecerit simile eis
EZEK|18|15|super montes non comederit et oculos suos non levaverit ad idola domus Israhel et uxorem proximi sui non violaverit
EZEK|18|16|et virum non contristaverit pignus non retinuerit et rapinam non rapuerit panem suum esurienti dederit et nudum operuerit vestimento
EZEK|18|17|a pauperis iniuria averterit manum suam usuram et superabundantiam non acceperit iudicia mea fecerit in praeceptis meis ambulaverit hic non morietur in iniquitate patris sui sed vita vivet
EZEK|18|18|pater eius quia calumniatus est et vim fecit fratri et malum operatus est in medio populi sui ecce mortuus est in iniquitate sua
EZEK|18|19|et dicitis quare non portavit filius iniquitatem patris videlicet quia filius iudicium et iustitiam operatus est omnia praecepta mea custodivit et fecit illa vita vivet
EZEK|18|20|anima quae peccaverit ipsa morietur filius non portabit iniquitatem patris et pater non portabit iniquitatem filii iustitia iusti super eum erit et impietas impii erit super eum
EZEK|18|21|si autem impius egerit paenitentiam ab omnibus peccatis suis quae operatus est et custodierit universa praecepta mea et fecerit iudicium et iustitiam vita vivet non morietur
EZEK|18|22|omnium iniquitatum eius quas operatus est non recordabor in iustitia sua quam operatus est vivet
EZEK|18|23|numquid voluntatis meae est mors impii dicit Dominus Deus et non ut convertatur a viis suis et vivat
EZEK|18|24|si autem averterit se iustus a iustitia sua et fecerit iniquitatem secundum omnes abominationes quas operari solet impius numquid vivet omnes iustitiae eius quas fecerat non recordabuntur in praevaricatione qua praevaricatus est et in peccato suo quod peccavit in ipsis morietur
EZEK|18|25|et dixistis non est aequa via Domini audite domus Israhel numquid via mea non est aequa et non magis viae vestrae pravae sunt
EZEK|18|26|cum enim averterit se iustus a iustitia sua et fecerit iniquitatem morietur in eis in iniustitia quam operatus est morietur
EZEK|18|27|et cum averterit se impius ab impietate sua quam operatus est et fecerit iudicium et iustitiam ipse animam suam vivificabit
EZEK|18|28|considerans enim et avertens se ab omnibus iniquitatibus suis quas operatus est vita vivet et non morietur
EZEK|18|29|et dicunt filii Israhel non est aequa via Domini numquid viae meae non sunt aequae domus Israhel et non magis viae vestrae pravae
EZEK|18|30|idcirco unumquemque iuxta vias suas iudicabo domus Israhel ait Dominus Deus convertimini et agite paenitentiam ab omnibus iniquitatibus vestris et non erit vobis in ruinam iniquitas
EZEK|18|31|proicite a vobis omnes praevaricationes vestras in quibus praevaricati estis et facite vobis cor novum et spiritum novum et quare moriemini domus Israhel
EZEK|18|32|quia nolo mortem morientis dicit Dominus Deus revertimini et vivite
EZEK|19|1|et tu adsume planctum super principes Israhel
EZEK|19|2|et dices quare mater tua leaena inter leones cubavit in medio leunculorum enutrivit catulos suos
EZEK|19|3|et eduxit unum de leunculis suis leo factus est et didicit capere praedam hominemque comedere
EZEK|19|4|et audierunt de eo gentes et non absque vulneribus suis ceperunt eum et adduxerunt eum in catenis in terram Aegypti
EZEK|19|5|quae cum vidisset quoniam infirmata est et periit expectatio eius tulit unum de leunculis suis leonem constituit eum
EZEK|19|6|qui incedebat inter leones et factus est leo didicit praedam capere et homines devorare
EZEK|19|7|didicit viduas facere et civitates eorum in desertum adducere et desolata est terra et plenitudo eius a voce rugitus illius
EZEK|19|8|et convenerunt adversum eum gentes undique de provinciis et expanderunt super eum rete suum in vulneribus earum captus est
EZEK|19|9|et miserunt eum in caveam in catenis adduxerunt eum ad regem Babylonis miseruntque eum in carcerem ne audiretur vox eius ultra super montes Israhel
EZEK|19|10|mater tua quasi vinea in sanguine tuo super aquam plantata fructus eius et frondes eius creverunt ex aquis multis
EZEK|19|11|et factae sunt ei virgae solidae in sceptra dominantium et exaltata est statura eius inter frondes et vidit altitudinem suam in multitudine palmitum suorum
EZEK|19|12|et evulsa est in ira in terramque proiecta et ventus urens siccavit fructum eius marcuerunt et arefactae sunt virgae roboris eius ignis comedit eam
EZEK|19|13|et nunc transplantata est in desertum in terra invia et sitienti
EZEK|19|14|et egressus est ignis de virga ramorum eius qui fructum eius comedit et non fuit in ea virga fortis sceptrum dominantium planctus est et erit in planctum
EZEK|20|1|et factum est in anno septimo in quinto mense in decima mensis venerunt viri de senioribus Israhel ut interrogarent Dominum et sederunt coram me
EZEK|20|2|et factus est sermo Domini ad me dicens
EZEK|20|3|fili hominis loquere senioribus Israhel et dices ad eos haec dicit Dominus Deus num ad interrogandum me vos venistis vivo ego quia non respondebo vobis ait Dominus Deus
EZEK|20|4|si iudicas eos si iudicas fili hominis abominationes patrum eorum ostende eis
EZEK|20|5|et dices ad eos haec dicit Dominus Deus in die qua elegi Israhel et levavi manum meam pro stirpe domus Iacob et apparui eis in terra Aegypti et levavi manum meam pro eis dicens ego Dominus Deus vester
EZEK|20|6|in die illa levavi manum meam pro eis ut educerem eos de terra Aegypti in terram quam provideram eis fluentem lacte et melle quae est egregia inter omnes terras
EZEK|20|7|et dixi ad eos unusquisque offensiones oculorum suorum abiciat et in idolis Aegypti nolite pollui ego Dominus Deus vester
EZEK|20|8|et inritaverunt me nolueruntque audire unusquisque abominationes oculorum suorum non proiecit nec idola Aegypti reliquerunt et dixi ut effunderem indignationem meam super eos et implerem iram meam in eis in medio terrae Aegypti
EZEK|20|9|et feci propter nomen meum ut non violaretur coram gentibus in quarum medio erant et inter quas apparui eis ut educerem eos de terra Aegypti
EZEK|20|10|eieci ergo eos de terra Aegypti et eduxi in desertum
EZEK|20|11|et dedi eis praecepta mea et iudicia mea ostendi eis quae faciat homo et vivat in eis
EZEK|20|12|insuper et sabbata mea dedi eis ut esset signum inter me et eos et scirent quia ego Dominus sanctificans eos
EZEK|20|13|et inritaverunt me domus Israhel in deserto in praeceptis meis non ambulaverunt et iudicia mea proiecerunt quae faciens homo vivet in eis et sabbata mea violaverunt vehementer dixi ergo ut effunderem furorem meum super eos in deserto et consumerem eos
EZEK|20|14|et feci propter nomen meum ne violaretur coram gentibus de quibus eieci eos in conspectu earum
EZEK|20|15|ego igitur levavi manum meam super eos in deserto ne inducerem eos in terram quam dedi eis fluentem lacte et melle praecipuam terrarum omnium
EZEK|20|16|quia iudicia mea proiecerunt et in praeceptis meis non ambulaverunt et sabbata mea violaverunt post idola enim cor eorum gradiebatur
EZEK|20|17|et pepercit oculus meus super eos ut non interficerem eos nec consumpsi eos in deserto
EZEK|20|18|dixi autem ad filios eorum in solitudine in praeceptis patrum vestrorum nolite incedere nec iudicia eorum custodiatis nec in idolis eorum polluamini
EZEK|20|19|ego Dominus Deus vester in praeceptis meis ambulate et iudicia mea custodite et facite ea
EZEK|20|20|et sabbata mea sanctificate ut sit signum inter me et vos et sciatur quia ego Dominus Deus vester
EZEK|20|21|et exacerbaverunt me filii in praeceptis meis non ambulaverunt et iudicia mea non custodierunt ut facerent ea quae cum fecerit homo vivet in eis et sabbata mea violaverunt et comminatus sum ut effunderem furorem meum super eos et implerem iram meam in eis in deserto
EZEK|20|22|averti autem manum meam et feci propter nomen meum ut non violaretur coram gentibus de quibus eieci eos in oculis earum
EZEK|20|23|iterum levavi manum meam in eos in solitudine ut dispergerem illos in nationes et ventilarem in terras
EZEK|20|24|eo quod iudicia mea non fecissent et praecepta mea reprobassent et sabbata mea violassent et post idola patrum suorum fuissent oculi eorum
EZEK|20|25|ergo et ego dedi eis praecepta non bona et iudicia in quibus non vivent
EZEK|20|26|et pollui eos in muneribus suis cum offerrent omne quod aperit vulvam propter delicta sua et scient quia ego Dominus
EZEK|20|27|quam ob rem loquere ad domum Israhel fili hominis et dices ad eos haec dicit Dominus Deus adhuc et in hoc blasphemaverunt me patres vestri cum sprevissent me contemnentes
EZEK|20|28|et induxissem eos in terram super quam levavi manum meam ut darem eis viderunt omnem collem excelsum et omne lignum nemorosum et immolaverunt ibi victimas suas et dederunt ibi inritationem oblationis suae et posuerunt ibi odorem suavitatis suae et libaverunt libationes suas
EZEK|20|29|et dixi ad eos quid est excelsum ad quod vos ingredimini et vocatum est nomen eius Excelsum usque ad hanc diem
EZEK|20|30|propterea dic ad domum Israhel haec dicit Dominus Deus certe in via patrum vestrorum vos polluimini et post offendicula eorum vos fornicamini
EZEK|20|31|et in oblatione donorum vestrorum cum transducitis filios vestros per ignem vos polluimini in omnibus idolis vestris usque hodie et ego respondebo vobis domus Israhel vivo ego dicit Dominus Deus quia non respondebo vobis
EZEK|20|32|neque cogitatio mentis vestrae fiet dicentium erimus sicut gentes et sicut cognationes terrae ut colamus ligna et lapides
EZEK|20|33|vivo ego dicit Dominus Deus quoniam in manu forti et brachio extento et in furore effuso regnabo super vos
EZEK|20|34|et educam vos de populis et congregabo vos de terris in quibus dispersi estis in manu valida et brachio extento et in furore effuso regnabo super vos
EZEK|20|35|et adducam vos in desertum populorum et iudicabor vobiscum ibi facie ad faciem
EZEK|20|36|sicut iudicio contendi adversum patres vestros in deserto terrae Aegypti sic iudicabo vos dicit Dominus Deus
EZEK|20|37|et subiciam vos sceptro meo et inducam vos in vinculis foederis
EZEK|20|38|et eligam de vobis transgressores et impios et de terra incolatus eorum educam eos et terram Israhel non ingredientur et scietis quia ego Dominus
EZEK|20|39|et vos domus Israhel haec dicit Dominus Deus singuli post idola vestra ambulate et servite eis quod si et in hoc non audieritis me et nomen meum sanctum pollueritis ultra in muneribus vestris et in idolis vestris
EZEK|20|40|in monte sancto meo in monte excelso Israhel ait Dominus Deus ibi serviet mihi omnis domus Israhel omnes inquam in terra in qua placebunt mihi et ibi quaeram primitias vestras et initium decimarum vestrarum in omnibus sanctificationibus vestris
EZEK|20|41|in odorem suavitatis suscipiam vos cum eduxero vos de populis et congregavero vos de terris in quas dispersi estis et sanctificabor in vobis in oculis nationum
EZEK|20|42|et scietis quia ego Dominus cum induxero vos ad terram Israhel in terram pro qua levavi manum meam ut darem eam patribus vestris
EZEK|20|43|et recordabimini ibi viarum vestrarum et omnium scelerum vestrorum quibus polluti estis in eis et displicebitis vobis in conspectu vestro in omnibus malitiis vestris quas fecistis
EZEK|20|44|et scietis quia ego Dominus cum benefecero vobis propter nomen meum non secundum vias vestras malas neque secundum scelera vestra pessima domus Israhel ait Dominus Deus
EZEK|20|45|et factus est sermo Domini ad me dicens
EZEK|20|46|fili hominis pone faciem tuam contra viam austri et stilla ad africum et propheta ad saltum agri meridiani
EZEK|20|47|et dices saltui meridiano audi verbum Domini haec dicit Dominus Deus ecce ego succendam in te ignem et conburam in te omne lignum viride et omne lignum aridum non extinguetur flamma succensionis et conburetur in ea omnis facies ab austro usque ad aquilonem
EZEK|20|48|et videbit universa caro quia ego Dominus succendi eam nec extinguetur
EZEK|20|49|et dixi ha ha ha Domine Deus ipsi dicunt de me numquid non per parabolas loquitur iste
EZEK|21|1|et factus est sermo Domini ad me dicens
EZEK|21|2|fili hominis pone faciem tuam ad Hierusalem et stilla ad sanctuaria et propheta contra humum Israhel
EZEK|21|3|et dices terrae Israhel haec dicit Dominus Deus ecce ego ad te et eiciam gladium meum de vagina sua et occidam in te iustum et impium
EZEK|21|4|pro eo autem quod occidi in te iustum et impium idcirco egredietur gladius meus de vagina sua ad omnem carnem ab austro ad aquilonem
EZEK|21|5|ut sciat omnis caro quia ego Dominus eduxi gladium meum de vagina sua inrevocabilem
EZEK|21|6|et tu fili hominis ingemesce in contritione lumborum et in amaritudinibus ingemesce coram eis
EZEK|21|7|cumque dixerint ad te quare tu gemis dices pro auditu quia venit et tabescet omne cor et dissolventur universae manus et infirmabitur omnis spiritus et per cuncta genua fluent aquae ecce venit et fiet ait Dominus Deus
EZEK|21|8|et factus est sermo Domini ad me dicens
EZEK|21|9|fili hominis propheta et dices haec dicit Dominus Deus loquere gladius gladius exacutus est et limatus
EZEK|21|10|ut caedat victimas exacutus est ut splendeat limatus est qui moves sceptrum filii mei succidisti omne lignum
EZEK|21|11|et dedi eum ad levigandum ut teneatur manu iste exacutus est gladius et iste limatus ut sit in manu interficientis
EZEK|21|12|clama et ulula fili hominis quia hic factus est in populo meo hic in cunctis ducibus Israhel qui fugerant gladio traditi sunt cum populo meo idcirco plaude super femur
EZEK|21|13|quia probatus est et hoc cum sceptrum subverterit et non erit dicit Dominus Deus
EZEK|21|14|tu ergo fili hominis propheta et percute manu ad manum et duplicetur gladius ac triplicetur gladius interfectorum hic est gladius occisionis magnae qui obstupescere eos facit
EZEK|21|15|et corde tabescere et multiplicat ruinas in omnibus portis eorum dedi conturbationem gladii acuti et limati ad fulgendum amicti ad caedem
EZEK|21|16|exacuere vade ad dextram sive ad sinistram quocumque faciei tuae est appetitus
EZEK|21|17|quin et ego plaudam manu ad manum et implebo indignationem meam ego Dominus locutus sum
EZEK|21|18|et factus est sermo Domini ad me dicens
EZEK|21|19|et tu fili hominis pone tibi duas vias ut veniat gladius regis Babylonis de terra una egredientur ambo et manu capiet coniecturam in capite viae civitatis coniciet
EZEK|21|20|viam pones ut veniat gladius ad Rabbath filiorum Ammon et ad Iudam in Hierusalem munitissimam
EZEK|21|21|stetit enim rex Babylonis in bivio in capite duarum viarum divinationem quaerens commiscens sagittas interrogavit idola exta consuluit
EZEK|21|22|ad dextram eius facta est divinatio super Hierusalem ut ponat arietes ut aperiat os in caede ut elevet vocem in ululatu ut ponat arietes contra portas ut conportet aggerem ut aedificet munitiones
EZEK|21|23|eritque quasi consulens frustra oraculum in oculis eorum et sabbatorum otium imitans ipse autem recordabitur iniquitatis ad capiendum
EZEK|21|24|idcirco haec dicit Dominus Deus pro eo quod recordati estis iniquitatis vestrae et revelastis praevaricationes vestras et apparuerunt peccata vestra in omnibus cogitationibus vestris pro eo inquam quod recordati estis manu capiemini
EZEK|21|25|tu autem profane impie dux Israhel cuius venit dies in tempore iniquitatis praefinita
EZEK|21|26|haec dicit Dominus Deus aufer cidarim tolle coronam nonne haec est quae humilem sublevavit et sublimem humiliavit
EZEK|21|27|iniquitatem iniquitatem iniquitatem ponam eam et hoc nunc factum est donec veniret cuius est iudicium et tradam ei
EZEK|21|28|et tu fili hominis propheta et dic haec dicit Dominus Deus ad filios Ammon et ad obprobrium eorum et dices mucro mucro evaginate ad occidendum limate ut interficias et fulgeas
EZEK|21|29|cum tibi viderentur vana et divinarentur mendacia ut dareris super colla vulneratorum impiorum quorum venit dies in tempore iniquitatis praefinita
EZEK|21|30|revertere ad vaginam tuam in loco in quo creatus es in terra nativitatis tuae iudicabo te
EZEK|21|31|et effundam super te indignationem meam in igne furoris mei sufflabo in te daboque te in manus hominum insipientium et fabricantium interitum
EZEK|21|32|igni eris cibus sanguis tuus erit in medio terrae oblivioni traderis quia ego Dominus locutus sum
EZEK|22|1|et factum est verbum Domini ad me dicens
EZEK|22|2|et tu fili hominis num iudicas num iudicas civitatem sanguinum
EZEK|22|3|et ostendes ei omnes abominationes suas et dices haec dicit Dominus Deus civitas effundens sanguinem in medio sui ut veniat tempus eius et quae fecit idola contra semet ipsam ut pollueretur
EZEK|22|4|in sanguine tuo qui a te effusus est deliquisti et in idolis tuis quae fecisti polluta es et adpropinquare fecisti dies tuos et adduxisti tempus annorum tuorum propterea dedi te obprobrium gentibus et inrisionem universis terris
EZEK|22|5|quae iuxta sunt et quae procul a te triumphabunt de te sordida nobilis grandis interitu
EZEK|22|6|ecce principes Israhel singuli in brachio suo fuerunt in te ad effundendum sanguinem
EZEK|22|7|patrem et matrem contumeliis adfecerunt in te advenam calumniati sunt in medio tui pupillum et viduam contristaverunt apud te
EZEK|22|8|sanctuaria mea sprevistis et sabbata mea polluistis
EZEK|22|9|viri detractores fuerunt in te ad effundendum sanguinem et super montes comederunt in te scelus operati sunt in medio tui
EZEK|22|10|verecundiora patris discoperuerunt in te inmunditiam menstruatae humiliaverunt in te
EZEK|22|11|et unusquisque in uxorem proximi sui operatus est abominationem et socer nurum suam polluit nefarie frater sororem suam filiam patris sui oppressit in te
EZEK|22|12|munera acceperunt apud te ad effundendum sanguinem usuram et superabundantiam accepisti et avare proximos tuos calumniabaris meique oblita es ait Dominus Deus
EZEK|22|13|ecce conplosi manus meas super avaritiam tuam quam fecisti et super sanguinem qui effusus est in medio tui
EZEK|22|14|numquid sustinebit cor tuum aut praevalebunt manus tuae in diebus quos ego faciam tibi ego Dominus locutus sum et faciam
EZEK|22|15|et dispergam te in nationes et ventilabo te in terras et deficere faciam inmunditiam tuam a te
EZEK|22|16|et possidebo te in conspectu gentium et scies quia ego Dominus
EZEK|22|17|et factum est verbum Domini ad me dicens
EZEK|22|18|fili hominis versa est mihi domus Israhel in scoriam omnes isti aes et stagnum et ferrum et plumbum in medio fornacis scoria argenti facti sunt
EZEK|22|19|propterea haec dicit Dominus Deus eo quod versi estis omnes in scoriam propterea ecce ego congregabo vos in medium Hierusalem
EZEK|22|20|congregatione argenti et aeris et ferri et stagni et plumbi in medium fornacis ut succendam in eam ignem ad conflandum sic congregabo in furore meo et in ira mea et requiescam et conflabo vos
EZEK|22|21|et congregabo vos et succendam vos in igne furoris mei et conflabimini in medio eius
EZEK|22|22|ut conflatur argentum in medio fornacis sic eritis in medio eius et scietis quia ego Dominus effuderim indignationem meam super vos
EZEK|22|23|et factum est verbum Domini ad me dicens
EZEK|22|24|fili hominis dic ei tu es terra inmunda et non conpluta in die furoris
EZEK|22|25|coniuratio prophetarum in medio eius sicut leo rugiens capiensque praedam animam devoraverunt opes et pretium acceperunt viduas eius multiplicaverunt in medio illius
EZEK|22|26|sacerdotes eius contempserunt legem meam et polluerunt sanctuaria mea inter sanctum et profanum non habuere distantiam et inter pollutum et mundum non intellexerunt et a sabbatis meis averterunt oculos suos et coinquinabar in medio eorum
EZEK|22|27|principes eius in medio illius quasi lupi rapientes praedam ad effundendum sanguinem et perdendas animas et avare sectanda lucra
EZEK|22|28|prophetae autem eius liniebant eos absque temperamento videntes vana et divinantes eis mendacium dicentes haec dicit Dominus Deus cum Dominus non sit locutus
EZEK|22|29|populi terrae calumniabantur calumniam et rapiebant violenter egenum et pauperem adfligebant et advenam opprimebant calumnia absque iudicio
EZEK|22|30|et quaesivi de eis virum qui interponeret sepem et staret oppositus contra me pro terra ne dissiparem eam et non inveni
EZEK|22|31|et effudi super eos indignationem meam in igne irae meae consumpsi eos viam eorum in caput eorum reddidi ait Dominus Deus
EZEK|23|1|et factus est sermo Domini ad me dicens
EZEK|23|2|fili hominis duae mulieres filiae matris unius fuerunt
EZEK|23|3|et fornicatae sunt in Aegypto in adulescentia sua fornicatae sunt ibi subacta sunt ubera earum et fractae sunt mammae pubertatis earum
EZEK|23|4|nomina autem earum Oolla maior et Ooliba soror eius et habui eas et pepererunt filios et filias porro earum nomina Samaria Oolla et Hierusalem Ooliba
EZEK|23|5|fornicata est igitur Oolla super me et insanivit in amatores suos in Assyrios propinquantes
EZEK|23|6|vestitos hyacintho principes et magistratus iuvenes cupidinis universos equites ascensores equorum
EZEK|23|7|et dedit fornicationes suas super eos electos filios Assyriorum universos et in omnibus in quos insanivit in inmunditiis eorum polluta est
EZEK|23|8|insuper et fornicationes suas quas habuerat in Aegypto non reliquit nam et illi dormierant cum ea in adulescentia eius et illi confregerant ubera pubertatis eius et effuderant fornicationem suam super eam
EZEK|23|9|propterea tradidi eam in manu amatorum suorum in manus filiorum Assur super quorum insanivit libidinem
EZEK|23|10|ipsi discoperuerunt ignominiam eius filios et filias illius tulerunt et ipsam occiderunt gladio et factae sunt famosae mulieres et iudicia perpetrarunt in ea
EZEK|23|11|quod cum vidisset soror eius Ooliba plus quam illa insanivit libidine et fornicationem suam super fornicationem sororis suae
EZEK|23|12|ad filios Assyriorum praebuit inpudenter ducibus et magistratibus ad se venientibus indutis veste varia equitibus qui vectabantur equis et adulescentibus forma cunctis egregia
EZEK|23|13|et vidi quod polluta esset via una ambarum
EZEK|23|14|et auxit fornicationes suas cumque vidisset viros depictos in pariete imagines Chaldeorum expressas coloribus
EZEK|23|15|et accinctos balteis renes et tiaras tinctas in capitibus eorum formam ducum omnium similitudinem filiorum Babylonis terraeque Chaldeorum in qua orti sunt
EZEK|23|16|et insanivit super eos concupiscentia oculorum suorum et misit nuntios ad eos in Chaldeam
EZEK|23|17|cumque venissent ad eam filii Babylonis ad cubile mammarum polluerunt eam stupris suis et polluta est ab eis et saturata est anima eius ab illis
EZEK|23|18|denudavit quoque fornicationes suas et discoperuit ignominiam suam et recessit anima mea ab ea sicut recesserat anima mea a sorore eius
EZEK|23|19|multiplicavit enim fornicationes suas recordans dies adulescentiae suae quibus fornicata est in terra Aegypti
EZEK|23|20|et insanivit libidine super concubitu eorum quorum carnes sunt ut carnes asinorum et sicut fluxus equorum fluxus eorum
EZEK|23|21|et visitasti scelus adulescentiae tuae quando subacta sunt in Aegypto ubera tua et confractae mammae pubertatis tuae
EZEK|23|22|propterea Ooliba haec dicit Dominus Deus ecce ego suscitabo omnes amatores tuos contra te de quibus satiata est anima tua et congregabo eos adversum te in circuitu
EZEK|23|23|filios Babylonis et universos Chaldeos nobiles tyrannosque et principes omnes filios Assyriorum iuvenes forma egregia duces et magistratus universos principes principum et nominatos ascensores equorum
EZEK|23|24|et venient super te instructi curru et rota multitudo populorum lorica et clypeo et galea armabuntur contra te undique et dabo coram eis iudicium et iudicabunt te iudiciis suis
EZEK|23|25|et ponam zelum meum in te quem exercent tecum in furore nasum tuum et aures tuas praecident et quae remanserint gladio concident ipsi filios tuos et filias tuas capient et novissimum tuum devorabitur igni
EZEK|23|26|et denudabunt te vestimentis tuis et tollent vasa gloriae tuae
EZEK|23|27|et requiescere faciam scelus tuum de te et fornicationem tuam de terra Aegypti nec levabis oculos tuos ad eos et Aegypti non recordaberis amplius
EZEK|23|28|quia haec dicit Dominus Deus ecce ego tradam te in manu eorum quos odisti in manu de quibus satiata est anima tua
EZEK|23|29|et agent tecum in odio et tollent omnes labores tuos et dimittent te nudam et ignominia plenam revelabitur ignominia fornicationum tuarum scelus tuum et fornicationes tuae
EZEK|23|30|fecerunt haec tibi quia fornicata es post gentes inter quas polluta es in idolis eorum
EZEK|23|31|in via sororis tuae ambulasti et dabo calicem eius in manu tua
EZEK|23|32|haec dicit Dominus Deus calicem sororis tuae bibes profundum et latum eris in derisum et in subsannationem quae es capacissima
EZEK|23|33|ebrietate et dolore repleberis calice maeroris et tristitiae calice sororis tuae Samariae
EZEK|23|34|et bibes illum et epotabis usque ad feces et fragmenta eius devorabis et ubera tua lacerabis quia ego locutus sum ait Dominus Deus
EZEK|23|35|propterea haec dicit Dominus Deus quia oblita es mei et proiecisti me post corpus tuum tu quoque porta scelus tuum et fornicationes tuas
EZEK|23|36|et ait Dominus ad me dicens fili hominis numquid iudicas Oollam et Oolibam et adnuntias eis scelera earum
EZEK|23|37|quia adulterae sunt et sanguis in manibus earum et cum idolis suis fornicatae sunt insuper et filios suos quos genuerunt mihi obtulerunt eis ad devorandum
EZEK|23|38|sed et hoc fecerunt mihi polluerunt sanctuarium meum in die illa et sabbata mea profanaverunt
EZEK|23|39|cumque immolarent filios suos idolis suis et ingrederentur sanctuarium meum in die illa ut polluerent illud etiam haec fecerunt in medio domus meae
EZEK|23|40|miserunt ad viros venientes de longe ad quos nuntium miserant itaque ecce venerunt quibus te lavisti et circumlevisti stibio oculos tuos et ornata es mundo muliebri
EZEK|23|41|sedisti in lecto pulcherrimo et mensa ordinata est ante te thymiama meum et unguentum meum posuisti super eam
EZEK|23|42|et vox multitudinis exultantis erat in ea et in viris qui de multitudine hominum adducebantur et veniebant de deserto posuerunt armillas in manibus eorum et coronas speciosas in capitibus eorum
EZEK|23|43|et dixi ei quae adtrita est in adulteriis nunc fornicabitur in fornicatione sua etiam haec
EZEK|23|44|et ingressi sunt ad eam quasi ad mulierem meretricem sic ingrediebantur ad Oollam et ad Oolibam mulieres nefarias
EZEK|23|45|viri ergo iusti sunt hii iudicabunt eas iudicio adulterarum et iudicio effundentium sanguinem quia adulterae sunt et sanguis in manibus earum
EZEK|23|46|haec enim dicit Dominus Deus adduc ad eas multitudinem et trade eas in tumultum et in rapinam
EZEK|23|47|et lapidentur lapidibus populorum et confodiantur gladiis eorum filios et filias earum interficient et domos earum igne succendent
EZEK|23|48|et auferam scelus de terra et discent omnes mulieres ne faciant secundum scelus earum
EZEK|23|49|et dabunt scelus vestrum super vos et peccata idolorum vestrorum portabitis et scietis quia ego Dominus Deus
EZEK|24|1|et factum est verbum Domini ad me in anno nono in mense decimo decima mensis dicens
EZEK|24|2|fili hominis scribe tibi nomen diei huius in qua confirmatus est rex Babylonis adversum Hierusalem hodie
EZEK|24|3|et dices per proverbium ad domum inritatricem parabolam et loqueris ad eos haec dicit Dominus Deus pone ollam pone inquam et mitte in ea aquam
EZEK|24|4|congere frusta eius in ea omnem partem bonam femur et armum electa et ossibus plena
EZEK|24|5|pinguissimum pecus adsume conpone quoque struices ossuum sub ea efferbuit coctio eius et discocta sunt ossa illius in medio eius
EZEK|24|6|propterea haec dicit Dominus Deus vae civitati sanguinum ollae cuius rubigo in ea est et rubigo eius non exivit de ea per partes et per partes suas eice eam non cecidit super eam sors
EZEK|24|7|sanguis enim eius in medio eius est super limpidissimam petram effudit illum non effudit illum super terram ut possit operiri pulvere
EZEK|24|8|ut superducerem indignationem meam et vindicta ulciscerer dedi sanguinem eius super petram limpidissimam ne operiretur
EZEK|24|9|propterea haec dicit Dominus Deus vae civitati sanguinum cuius ego grandem faciam pyram
EZEK|24|10|congere ossa quae igne succendam consumentur carnes et concoquetur universa conpositio et ossa tabescent
EZEK|24|11|pone quoque eam super prunas vacuam ut incalescat et liquefiat aes eius et confletur in medio eius inquinamentum eius et consumatur rubigo eius
EZEK|24|12|multo labore sudatum est et non exibit de ea nimia rubigo eius neque per ignem
EZEK|24|13|inmunditia tua execrabilis quia mundare te volui et non es mundata a sordibus tuis sed nec mundaberis prius donec quiescere faciam indignationem meam in te
EZEK|24|14|ego Dominus locutus sum venit et faciam non transeam nec parcam nec placabor iuxta vias tuas et iuxta adinventiones tuas iudicavi te dicit Dominus
EZEK|24|15|et factum est verbum Domini ad me dicens
EZEK|24|16|fili hominis ecce ego tollo a te desiderabile oculorum tuorum in plaga et non planges neque plorabis neque fluent lacrimae tuae
EZEK|24|17|ingemesce tacens mortuorum luctum non facies corona tua circumligata sit tibi et calciamenta tua erunt in pedibus tuis nec amictu ora velabis nec cibos lugentium comedes
EZEK|24|18|locutus sum ergo ad populum mane et mortua est uxor mea vesperi fecique mane sicut praeceperat mihi
EZEK|24|19|et dixit ad me populus quare non indicas nobis quid ista significent quae tu facis
EZEK|24|20|et dixi ad eos sermo Domini factus est ad me dicens
EZEK|24|21|loquere domui Israhel haec dicit Dominus Deus ecce ego polluam sanctuarium meum superbiam imperii vestri et desiderabile oculorum vestrorum et super quo pavet anima vestra et filii vestri et filiae quas reliquistis gladio cadent
EZEK|24|22|et facietis sicut feci ora amictu non velabitis et cibos lugentium non comedetis
EZEK|24|23|coronas habebitis in capitibus vestris et calciamenta in pedibus non plangetis neque flebitis sed tabescetis in iniquitatibus vestris et unusquisque gemet ad fratrem suum
EZEK|24|24|eritque Hiezecihel vobis in portentum iuxta omnia quae fecit facietis cum venerit istud et scietis quia ego Dominus Deus
EZEK|24|25|et tu fili hominis ecce in die quo tollam ab eis fortitudinem eorum et gaudium dignitatis et desiderium oculorum eorum super quo requiescunt animae eorum filios et filias eorum
EZEK|24|26|in die illa cum venerit fugiens ad te ut adnuntiet tibi
EZEK|24|27|in die inquam illa aperietur os tuum cum eo qui fugit et loqueris et non silebis ultra erisque eis in portentum et scietis quia ego Dominus
EZEK|25|1|et factus est sermo Domini ad me dicens
EZEK|25|2|fili hominis pone faciem tuam contra filios Ammon et prophetabis de eis
EZEK|25|3|et dices filiis Ammon audite verbum Domini Dei haec dicit Dominus Deus pro eo quod dixisti euge euge super sanctuarium meum quia pollutum est et super terram Israhel quoniam desolata est et super domum Iuda quoniam ducti sunt in captivitatem
EZEK|25|4|idcirco ego tradam te filiis orientalibus in hereditatem et conlocabunt caulas suas in te et ponent in te tentoria sua ipsi comedent fruges tuas et ipsi bibent lac tuum
EZEK|25|5|daboque Rabbath in habitaculum camelorum et filios Ammon in cubile pecorum et scietis quia ego Dominus
EZEK|25|6|quia haec dicit Dominus Deus pro eo quod plausisti manu et percussisti pede et gavisa es ex toto affectu super terram Israhel
EZEK|25|7|idcirco ecce ego extendam manum meam super te et tradam te in direptionem gentium et interficiam te de populis et perdam de terris et conteram et scies quia ego Dominus
EZEK|25|8|haec dicit Dominus Deus pro eo quod dixerunt Moab et Seir ecce sicut omnes gentes domus Iuda
EZEK|25|9|idcirco ecce ego aperiam umerum Moab de civitatibus de civitatibus inquam eius et de finibus eius inclitas terrae Bethiesimoth et Beelmeon et Cariathaim
EZEK|25|10|filiis orientis cum filiis Ammon et dabo eam in hereditatem ut non sit memoria ultra filiorum Ammon in gentibus
EZEK|25|11|et in Moab faciam iudicia et scient quia ego Dominus
EZEK|25|12|haec dicit Dominus Deus pro eo quod fecit Idumea ultionem ut se vindicaret de filiis Iuda peccavitque delinquens et vindictam expetivit de eis
EZEK|25|13|idcirco haec dicit Dominus Deus extendam manum meam super Idumeam et auferam de ea hominem et iumentum et faciam eam desertum ab austro et qui sunt in Daedan gladio cadent
EZEK|25|14|et dabo ultionem meam super Idumeam per manum populi mei Israhel et facient in Edom iuxta iram meam et furorem meum et scient vindictam meam dicit Dominus Deus
EZEK|25|15|haec dicit Dominus Deus pro eo quod fecerunt Palestini in vindictam et ulti se sunt toto animo interficientes et implentes inimicitias veteres
EZEK|25|16|propterea haec dicit Dominus Deus ecce ego extendam manum meam super Palestinos et interficiam interfectores et perdam reliquias maritimae regionis
EZEK|25|17|faciamque in eis ultiones magnas arguens in furore et scient quia ego Dominus cum dedero vindictam meam super eos
EZEK|26|1|et factum est in undecimo anno prima mensis factus est sermo Domini ad me dicens
EZEK|26|2|fili hominis pro eo quod dixit Tyrus de Hierusalem euge confractae sunt portae populorum conversa est ad me implebor deserta est
EZEK|26|3|propterea haec dicit Dominus Deus ecce ego super te Tyre et ascendere faciam ad te gentes multas sicut ascendit mare fluctuans
EZEK|26|4|et dissipabunt muros Tyri et destruent turres eius et radam pulverem eius de ea et dabo eam in limpidissimam petram
EZEK|26|5|siccatio sagenarum erit in medio maris quia ego locutus sum ait Dominus Deus et erit in direptionem gentibus
EZEK|26|6|filiae quoque eius quae sunt in agro gladio interficientur et scient quia ego Dominus
EZEK|26|7|quia haec dicit Dominus Deus ecce ego adducam ad Tyrum Nabuchodonosor regem Babylonis ab aquilone regem regum cum equis et curribus et equitibus et coetu populoque magno
EZEK|26|8|filias tuas quae sunt in agro gladio interficiet et circumdabit te munitionibus et conportabit aggerem in gyro et levabit contra te clypeum
EZEK|26|9|et vineas et arietes temperabit in muros tuos et turres tuas destruet in armatura sua
EZEK|26|10|inundatione equorum eius operiet te pulvis eorum a sonitu equitum et rotarum et curruum movebuntur muri tui dum ingressus fuerit portas tuas quasi per introitus urbis dissipatae
EZEK|26|11|ungulis equorum suorum conculcabit omnes plateas tuas populum tuum gladio caedet et statuae tuae nobiles in terram corruent
EZEK|26|12|vastabunt opes tuas diripient negotiationes tuas et destruent muros tuos et domos tuas praeclaras subvertent et lapides tuos et ligna tua et pulverem tuum in medio aquarum ponent
EZEK|26|13|et quiescere faciam multitudinem canticorum tuorum et sonitus cithararum tuarum non audietur amplius
EZEK|26|14|et dabo te in limpidissimam petram siccatio sagenarum eris nec aedificaberis ultra quia ego locutus sum dicit Dominus Deus
EZEK|26|15|haec dicit Dominus Deus Tyro numquid non a sonitu ruinae tuae et gemitu interfectorum tuorum cum occisi fuerint in medio tui commovebuntur insulae
EZEK|26|16|et descendent de sedibus suis omnes principes maris et auferent exuvias suas et vestimenta sua varia abicient et induentur stupore in terra sedebunt et adtoniti super repentino casu tuo admirabuntur
EZEK|26|17|et adsumentes super te lamentum dicent tibi quomodo peristi quae habitas in mari urbs inclita quae fuisti fortis in mari cum habitatoribus tuis quos formidabant universi
EZEK|26|18|nunc stupebunt naves in die pavoris tui et turbabuntur insulae in mari eo quod nullus egrediatur ex te
EZEK|26|19|quia haec dicit Dominus Deus cum dedero te urbem desolatam sicut civitates quae non habitantur et adduxero super te abyssum et operuerint te aquae multae
EZEK|26|20|et detraxero te cum his qui descendunt in lacum ad populum sempiternum et conlocavero te in terra novissima sicut solitudines veteres cum his qui deducuntur in lacum ut non habiteris porro dedero gloriam in terra viventium
EZEK|26|21|in nihilum redigam te et non eris et requisita non invenieris ultra in sempiternum dicit Dominus Deus
EZEK|27|1|et factum est verbum Domini ad me dicens
EZEK|27|2|tu ergo fili hominis adsume super Tyrum lamentum
EZEK|27|3|et dices Tyro quae habitat in introitu maris negotiationi populorum ad insulas multas haec dicit Dominus Deus o Tyre tu dixisti perfecti decoris ego sum
EZEK|27|4|et in corde maris sita finitimi tui qui te aedificaverunt impleverunt decorem tuum
EZEK|27|5|abietibus de Sanir extruxerunt te cum omnibus tabulatis maris cedrum de Libano tulerunt ut facerent tibi malum
EZEK|27|6|quercus de Basan dolaverunt in remos tuos transtra tua fecerunt tibi ex ebore indico et praetoriola de insulis Italiae
EZEK|27|7|byssus varia de Aegypto texta est tibi in velum ut poneretur in malo hyacinthus et purpura de insulis Elisa facta sunt operimentum tuum
EZEK|27|8|habitatores Sidonis et Aradii fuerunt remiges tui sapientes tui Tyre facti sunt gubernatores tui
EZEK|27|9|senes Bibli et prudentes eius habuerunt nautas ad ministerium variae supellectilis tuae omnes naves maris et nautae earum fuerunt in populo negotiationis tuae
EZEK|27|10|Persae et Lydi et Lybies erant in exercitu tuo viri bellatores tui clypeum et galeam suspenderunt in te pro ornatu tuo
EZEK|27|11|filii Aradii cum exercitu tuo erant super muros tuos in circuitu sed et Pigmei qui erant in turribus tuis faretras suas suspenderunt in muris tuis per gyrum ipsi conpleverunt pulchritudinem tuam
EZEK|27|12|Carthaginienses negotiatores tui a multitudine cunctarum divitiarum argento ferro stagno plumboque repleverunt nundinas tuas
EZEK|27|13|Graecia Thubal et Mosoch ipsi institores tui mancipia et vasa aerea adduxerunt populo tuo
EZEK|27|14|de domo Thogorma equos et equites et mulos adduxerunt ad forum tuum
EZEK|27|15|filii Dadan negotiatores tui insulae multae negotiatio manus tuae dentes eburneos et hebeninos commutaverunt in pretio tuo
EZEK|27|16|Syrus negotiator tuus propter multitudinem operum tuorum gemmam purpuram et scutulata et byssum et sericum et chodchod proposuerunt in mercatu tuo
EZEK|27|17|Iuda et terra Israhel ipsi institores tui in frumento primo balsamum et mel et oleum et resinam proposuerunt in nundinis tuis
EZEK|27|18|Damascenus negotiator tuus in multitudine operum tuorum in multitudine diversarum opum in vino pingui in lanis coloris optimi
EZEK|27|19|Dan et Graecia et Mozel in nundinis tuis proposuerunt ferrum fabrefactum stacte et calamus in negotiatione tua
EZEK|27|20|Dadan institores tui in tapetibus ad sedendum
EZEK|27|21|Arabia et universi principes Cedar ipsi negotiatores manus tuae cum agnis et arietibus et hedis venerunt ad te negotiatores tui
EZEK|27|22|venditores Saba et Reema ipsi negotiatores tui cum universis primis aromatibus et lapide pretioso et auro quod proposuerunt in mercatu tuo
EZEK|27|23|Aran et Chenne et Eden negotiatores Saba Assur Chelmad venditores tui
EZEK|27|24|ipsi negotiatores tui multifariam involucris hyacinthi et polymitorum gazarumque pretiosarum quae obvolutae et adstrictae erant funibus cedros quoque habebant in negotiationibus tuis
EZEK|27|25|naves maris principes tuae in negotiatione tua et repleta es et glorificata nimis in corde maris
EZEK|27|26|in aquis multis adduxerunt te remiges tui ventus auster contrivit te in corde maris
EZEK|27|27|divitiae tuae et thesauri tui et multiplex instrumentum tuum nautae tui et gubernatores tui qui tenebant supellectilem tuam et populo tuo praeerant viri quoque bellatores tui qui erant in te cum universa multitudine tua quae est in medio tui cadent in corde maris in die ruinae tuae
EZEK|27|28|a sonitu clamoris gubernatorum tuorum conturbabuntur classes
EZEK|27|29|et descendent de navibus suis omnes qui tenebant remum nautae et universi gubernatores maris in terra stabunt
EZEK|27|30|et heiulabunt super te voce magna et clamabunt amare et superiacient pulverem capitibus suis et cinere conspergentur
EZEK|27|31|et radent super te calvitium et accingentur ciliciis et plorabunt te in amaritudine animae ploratu amarissimo
EZEK|27|32|et adsument super te carmen lugubre et plangent te quae est ut Tyrus quae obmutuit in medio maris
EZEK|27|33|quae in exitu negotiationum tuarum de mari implesti populos multos in multitudine divitiarum tuarum et populorum tuorum ditasti reges terrae
EZEK|27|34|nunc contrita es a mari in profundis aquarum opes tuae et omnis multitudo tua quae erat in medio tui ceciderunt
EZEK|27|35|universi habitatores insularum obstipuerunt super te et reges earum omnes tempestate perculsi mutaverunt vultus
EZEK|27|36|negotiatores populorum sibilaverunt super te ad nihilum deducta es et non eris usque in perpetuum
EZEK|28|1|et factus est sermo Domini ad me dicens
EZEK|28|2|fili hominis dic principi Tyri haec dicit Dominus Deus eo quod elevatum est cor tuum et dixisti Deus ego sum et in cathedra Dei sedi in corde maris cum sis homo et non Deus et dedisti cor tuum quasi cor Dei
EZEK|28|3|ecce sapientior es tu Danihele omne secretum non est absconditum a te
EZEK|28|4|in sapientia et prudentia tua fecisti tibi fortitudinem et adquisisti aurum et argentum in thesauris tuis
EZEK|28|5|in multitudine sapientiae tuae et in negotiatione tua multiplicasti tibi fortitudinem et elevatum est cor tuum in robore tuo
EZEK|28|6|propterea haec dicit Dominus Deus eo quod elevatum est cor tuum quasi cor Dei
EZEK|28|7|idcirco ecce ego adducam super te alienos robustissimos gentium et nudabunt gladios suos super pulchritudinem sapientiae tuae et polluent decorem tuum
EZEK|28|8|interficient et detrahent te et morieris interitu occisorum in corde maris
EZEK|28|9|numquid dicens loqueris Deus ego sum coram interficientibus te cum sis homo et non Deus in manu occidentium te
EZEK|28|10|morte incircumcisorum morieris in manu alienorum quia ego locutus sum ait Dominus Deus
EZEK|28|11|et factus est sermo Domini ad me dicens fili hominis leva planctum super regem Tyri
EZEK|28|12|et dices ei haec dicit Dominus Deus tu signaculum similitudinis plenus sapientia et perfectus decore
EZEK|28|13|in deliciis paradisi Dei fuisti omnis lapis pretiosus operimentum tuum sardius topazius et iaspis chrysolitus et onyx et berillus sapphyrus et carbunculus et zmaragdus aurum opus decoris tui et foramina tua in die qua conditus es praeparata sunt
EZEK|28|14|tu cherub extentus et protegens et posui te in monte sancto Dei in medio lapidum ignitorum ambulasti
EZEK|28|15|perfectus in viis tuis a die conditionis tuae donec inventa est iniquitas in te
EZEK|28|16|in multitudine negotiationis tuae repleta sunt interiora tua iniquitate et peccasti et eieci te de monte Dei et perdidi te o cherub protegens de medio lapidum ignitorum
EZEK|28|17|elevatum est cor tuum in decore tuo perdidisti sapientiam tuam in decore tuo in terram proieci te ante faciem regum dedi te ut cernerent te
EZEK|28|18|in multitudine iniquitatum tuarum et iniquitate negotiationis tuae polluisti sanctificationem tuam producam ergo ignem de medio tui qui comedat te et dabo te in cinerem super terram in conspectu omnium videntium te
EZEK|28|19|omnes qui viderint te in gentibus obstupescent super te nihili factus es et non eris in perpetuum
EZEK|28|20|et factus est sermo Domini ad me dicens
EZEK|28|21|fili hominis pone faciem tuam contra Sidonem et prophetabis de ea
EZEK|28|22|et dices haec dicit Dominus Deus ecce ego ad te Sidon et glorificabor in medio tui et scient quia ego Dominus cum fecero in ea iudicia et sanctificatus fuero in ea
EZEK|28|23|et inmittam ei pestilentiam et sanguinem in plateis eius et corruent interfecti in medio eius gladio per circuitum et scient quia ego Dominus
EZEK|28|24|et non erit ultra domui Israhel offendiculum amaritudinis et spina dolorem inferens undique per circuitum eorum qui adversantur eis et scient quia ego Dominus Deus
EZEK|28|25|haec dicit Dominus Deus quando congregavero domum Israhel de populis in quibus dispersi sunt sanctificabor in eis coram gentibus et habitabunt in terra sua quam dedi servo meo Iacob
EZEK|28|26|et habitabunt in ea securi et aedificabunt domos plantabuntque vineas et habitabunt confidenter cum fecero iudicia in omnibus qui adversantur eis per circuitum et scient quia ego Dominus Deus eorum
EZEK|29|1|in anno decimo in decimo mense undecima mensis factum est verbum Domini ad me dicens
EZEK|29|2|fili hominis pone faciem tuam contra Pharaonem regem Aegypti et prophetabis de eo et de Aegypto universa
EZEK|29|3|loquere et dices haec dicit Dominus Deus ecce ego ad te Pharao rex Aegypti draco magne qui cubas in medio fluminum tuorum et dicis meus est fluvius et ego feci memet ipsum
EZEK|29|4|et ponam frenum in maxillis tuis et adglutinabo pisces fluminum tuorum squamis tuis et extraham te de medio fluminum tuorum et universi pisces tui squamis tuis adherebunt
EZEK|29|5|et proiciam te in desertum et omnes pisces fluminis tui super faciem terrae cades non colligeris neque congregaberis bestiis terrae et volatilibus caeli dedi te ad devorandum
EZEK|29|6|et scient omnes habitatores Aegypti quia ego Dominus pro eo quod fuisti baculus harundineus domui Israhel
EZEK|29|7|quando adprehenderunt te manu et confractus es et lacerasti omnem umerum eorum et innitentibus eis super te comminutus es et dissolvisti omnes renes eorum
EZEK|29|8|propterea haec dicit Dominus Deus ecce ego adducam super te gladium et interficiam de te hominem et iumentum
EZEK|29|9|et erit terra Aegypti in desertum et solitudinem et scient quia ego Dominus eo quod dixerit fluvius meus est et ego feci
EZEK|29|10|idcirco ecce ego ad te et ad flumina tua daboque terram Aegypti in solitudines gladio dissipatam a turre Syenes usque ad terminos Aethiopiae
EZEK|29|11|non pertransibit eam pes hominis neque pes iumenti gradietur in ea et non habitabitur quadraginta annis
EZEK|29|12|daboque terram Aegypti desertam in medio terrarum desertarum et civitates eius in medio urbium subversarum erunt desolatae quadraginta annis et dispergam Aegyptios in nationes et ventilabo eos in terras
EZEK|29|13|quia haec dicit Dominus Deus post finem quadraginta annorum congregabo Aegyptum de populis in quibus dispersi fuerunt
EZEK|29|14|et reducam captivitatem Aegypti et conlocabo eos in terra Fatures in terra nativitatis suae et erunt ibi in regnum humile
EZEK|29|15|inter regna cetera erit humillima et non elevabitur ultra super nationes et inminuam eos ne imperent gentibus
EZEK|29|16|neque erunt ultra domui Israhel in confidentia docentes iniquitatem ut fugiant et sequantur eos et scient quia ego Dominus Deus
EZEK|29|17|et factum est in vicesimo et septimo anno in primo in una mensis factum est verbum Domini ad me dicens
EZEK|29|18|fili hominis Nabuchodonosor rex Babylonis servire fecit exercitum suum servitute magna adversum Tyrum omne caput decalvatum et omnis umerus depilatus est et merces non est reddita ei neque exercitui eius de Tyro pro servitute qua servivit mihi adversum eam
EZEK|29|19|propterea haec dicit Dominus Deus ecce ego dabo Nabuchodonosor regem Babylonis in terra Aegypti et accipiet multitudinem eius et depraedabitur manubias eius et diripiet spolia eius et erit merces exercitui illius
EZEK|29|20|et operi pro quo servivit adversum eam dedi ei terram Aegypti pro eo quod laboraverunt mihi ait Dominus Deus
EZEK|29|21|in die illo pullulabit cornu domui Israhel et tibi dabo apertum os in medio eorum et scient quoniam ego Dominus
EZEK|30|1|et factum est verbum Domini ad me dicens
EZEK|30|2|fili hominis propheta et dic haec dicit Dominus Deus ululate vae vae diei
EZEK|30|3|quia iuxta est dies et adpropinquavit dies Domini dies nubis tempus gentium erit
EZEK|30|4|et veniet gladius in Aegyptum et erit pavor in Aethiopia cum ceciderint vulnerati in Aegypto et ablata fuerit multitudo illius et destructa fundamenta eius
EZEK|30|5|Aethiopia et Lybia et Lydii et omne reliquum vulgus et Chub et filii terrae foederis cum eis gladio cadent
EZEK|30|6|haec dicit Dominus Deus et corruent fulcientes Aegyptum et destruetur superbia imperii eius a turre Syenes gladio cadent in ea ait Dominus exercituum
EZEK|30|7|et dissipabuntur in medio terrarum desolatarum et urbes eius in medio civitatum desertarum erunt
EZEK|30|8|et scient quoniam ego Dominus cum dedero ignem in Aegyptum et adtriti fuerint omnes auxiliatores eius
EZEK|30|9|in die illa egredientur nuntii a facie mea in trieribus ad conterendam Aethiopiae confidentiam et erit pavor in eis in die Aegypti quia absque dubio veniet
EZEK|30|10|haec dicit Dominus Deus et cessare faciam multitudinem Aegypti in manu Nabuchodonosor regis Babylonis
EZEK|30|11|ipse et populus eius cum eo fortissimi gentium adducentur ad disperdendam terram et evaginabunt gladios suos super Aegyptum et implebunt terram interfectis
EZEK|30|12|et faciam alveos fluminum aridos et tradam terram in manu pessimorum et dissipabo terram et plenitudinem eius in manu alienorum ego Dominus locutus sum
EZEK|30|13|haec dicit Dominus Deus et disperdam simulacra et cessare faciam idola de Memphis et dux de terra Aegypti non erit amplius et dabo terrorem in terra Aegypti
EZEK|30|14|et disperdam terram Fatures et dabo ignem in Tafnis et faciam iudicia in Alexandriam
EZEK|30|15|et effundam indignationem meam super Pelusium robur Aegypti et interficiam multitudinem Alexandriae
EZEK|30|16|et dabo ignem in Aegypto quasi parturiens dolebit Pelusium et Alexandria erit dissipata et in Memphis angustiae cotidianae
EZEK|30|17|iuvenes Eliupoleos et Bubasti gladio cadent et ipsae captivae ducentur
EZEK|30|18|et in Tafnis nigrescet dies cum contrivero ibi sceptra Aegypti et defecerit in ea superbia potentiae eius ipsam nubes operiet filiae autem eius in captivitatem ducentur
EZEK|30|19|et faciam iudicia in Aegypto et scient quia ego Dominus
EZEK|30|20|et factum est in undecimo anno in primo in septima mensis factum est verbum Domini ad me dicens
EZEK|30|21|fili hominis brachium Pharao regis Aegypti confregi et ecce non est obvolutum ut restitueretur ei sanitas ut ligaretur pannis et farciretur linteolis et recepto robore posset tenere gladium
EZEK|30|22|propterea haec dicit Dominus Deus ecce ego ad Pharao regem Aegypti et comminuam brachium eius forte sed confractum et deiciam gladium de manu eius
EZEK|30|23|et dispergam Aegyptum in gentibus et ventilabo eos in terris
EZEK|30|24|et confortabo brachia regis Babylonis daboque gladium meum in manu eius et confringam brachia Pharaonis et gement gemitibus interfecti coram facie eius
EZEK|30|25|et confortabo brachia regis Babylonis et brachia Pharaonis concident et scient quia ego Dominus cum dedero gladium meum in manu regis Babylonis et extenderit eum super terram Aegypti
EZEK|30|26|et dispergam Aegyptum in nationes et ventilabo eos in terris et scient quia ego Dominus
EZEK|31|1|et factum est in undecimo anno tertio una mensis factum est verbum Domini ad me dicens
EZEK|31|2|fili hominis dic Pharaoni regi Aegypti et populo eius cui similis factus es in magnitudine tua
EZEK|31|3|ecce Assur quasi cedrus in Libano pulcher ramis et frondibus nemorosus excelsusque altitudine et inter condensas frondes elevatum est cacumen eius
EZEK|31|4|aquae nutrierunt illum abyssus exaltavit eum flumina eius manabant in circuitu radicum eius et rivos suos emisit ad universa ligna regionis
EZEK|31|5|propterea elevata est altitudo eius super omnia ligna regionis et multiplicata sunt arbusta eius et elevati sunt rami eius prae aquis multis
EZEK|31|6|cumque extendisset umbram suam in ramis eius fecerunt nidos omnia volatilia caeli et sub frondibus eius genuerunt omnes bestiae saltuum et sub umbraculo illius habitabat coetus gentium plurimarum
EZEK|31|7|eratque pulcherrimus in magnitudine sua et in dilatatione arbustorum suorum erat enim radix illius iuxta aquas multas
EZEK|31|8|cedri non fuerunt altiores illo in paradiso Dei abietes non adaequaverunt summitatem eius et platani non fuerunt aequae frondibus illius omne lignum paradisi Dei non est adsimilatum illi et pulchritudini eius
EZEK|31|9|quoniam speciosum feci eum et multis condensisque frondibus et aemulata sunt eum omnia ligna voluptatis quae erant in paradiso Dei
EZEK|31|10|propterea haec dicit Dominus Deus pro eo quod sublimatus est in altitudine et dedit summitatem suam virentem atque condensam et elevatum est cor eius in altitudine sua
EZEK|31|11|tradidi eum in manu fortissimi gentium faciens faciet ei iuxta impietatem eius eieci eum
EZEK|31|12|et succident illum alieni et crudelissimi nationum et proicient eum super montes et in cunctis convallibus corruent rami eius et confringentur arbusta eius in universis rupibus terrae et recedent de umbraculo eius omnes populi terrae et relinquent eum
EZEK|31|13|in ruina eius habitaverunt omnia volatilia caeli et in ramis eius fuerunt universae bestiae regionis
EZEK|31|14|quam ob rem non elevabuntur in altitudine sua omnia ligna aquarum neque ponent sublimitatem suam inter nemorosa atque frondosa nec stabunt in sublimitate eorum omnia quae inrigantur aquis quia omnes traditi sunt in mortem ad terram ultimam in medio filiorum hominum ad eos qui descendunt in lacum
EZEK|31|15|haec dicit Dominus Deus in die quando descendit ad inferos indixi luctum operui eum abysso et prohibui flumina eius et coercui aquas multas contristatus est super eum Libanus et omnia ligna agri concussa sunt
EZEK|31|16|a sonitu ruinae eius commovi gentes cum deducerem eum ad infernum cum his qui descendebant in lacum et consolata sunt in terra infima omnia ligna voluptatis egregia atque praeclara in Libano universa quae inrigabantur aquis
EZEK|31|17|nam et ipsi cum ea descendent ad infernum ad interfectos gladio et brachium uniuscuiusque sedebit sub umbraculo eius in medio nationum
EZEK|31|18|cui adsimilatus es o inclite atque sublimis inter ligna voluptatis ecce deductus es cum lignis voluptatis ad terram ultimam in medio incircumcisorum dormies cum his qui interfecti sunt gladio ipse est Pharao et omnis multitudo eius dicit Dominus Deus
EZEK|32|1|et factum est duodecimo anno in mense duodecimo in una mensis factum est verbum Domini ad me dicens
EZEK|32|2|fili hominis adsume lamentum super Pharao regem Aegypti et dices ad eum leoni gentium adsimilatus es et draconi qui est in mari et ventilabas cornu in fluminibus tuis et conturbabas aquas pedibus tuis et conculcabas flumina eorum
EZEK|32|3|propterea haec dicit Dominus Deus expandam super te rete meum in multitudine populorum multorum et extrahent te in sagena mea
EZEK|32|4|et proiciam te in terram super faciem agri abiciam te et habitare faciam super te omnia volatilia caeli et saturabo de te bestias universae terrae
EZEK|32|5|et dabo carnes tuas super montes et implebo colles tuos sanie tua
EZEK|32|6|et inrigabo terram pedore sanguinis tui super montes et valles implebuntur ex te
EZEK|32|7|et operiam cum extinctus fueris caelos et nigrescere faciam stellas eius solem nube tegam et luna non dabit lumen suum
EZEK|32|8|omnia luminaria caeli maerere faciam super te et dabo tenebras super terram tuam dicit Dominus Deus
EZEK|32|9|et inritabo cor populorum multorum cum induxero contritionem tuam in gentibus super terras quas nescis
EZEK|32|10|et stupescere faciam super te populos multos et reges eorum horrore nimio formidabunt super te cum volare coeperit gladius meus super facies eorum et obstupescent repente singuli pro anima sua in die ruinae suae
EZEK|32|11|quia haec dicit Dominus Deus gladius regis Babylonis veniet tibi
EZEK|32|12|in gladiis fortium deiciam multitudinem tuam inexpugnabiles gentes omnes heae et vastabunt superbiam Aegypti et dissipabitur multitudo eius
EZEK|32|13|et perdam omnia iumenta eius quae erant super aquas plurimas et non conturbabit eas pes hominis ultra neque ungula iumentorum turbabit eas
EZEK|32|14|tunc purissimas reddam aquas eorum et flumina eorum quasi oleum adducam ait Dominus Deus
EZEK|32|15|cum dedero terram Aegypti desolatam deseretur autem terra a plenitudine sua quando percussero omnes habitatores eius et scient quia ego Dominus
EZEK|32|16|planctus est et plangent eum filiae gentium plangent eum super Aegypto et super multitudine eius plangent eum ait Dominus Deus
EZEK|32|17|et factum est in duodecimo anno in quintadecima mensis factum est verbum Domini ad me dicens
EZEK|32|18|fili hominis cane lugubre super multitudine Aegypti et detrahe eam ipsam et filias gentium robustarum ad terram ultimam cum his qui descendunt in lacum
EZEK|32|19|quo pulchrior es descende et dormi cum incircumcisis
EZEK|32|20|in medio interfectorum gladio cadent gladius datus est adtraxerunt eam et omnes populos eius
EZEK|32|21|loquentur ei potentissimi robustorum de medio inferni qui cum auxiliatoribus eius descenderunt et dormierunt incircumcisi interfecti gladio
EZEK|32|22|ibi Assur et omnis multitudo eius in circuitu illius sepulchra eius omnes interfecti et qui ceciderunt gladio
EZEK|32|23|quorum data sunt sepulchra in novissimis laci et facta est multitudo eius per gyrum sepulchri eius universi interfecti cadentesque gladio qui dederant quondam formidinem in terra viventium
EZEK|32|24|ibi Aelam et omnis multitudo eius per gyrum sepulchri sui omnes hii interfecti ruentesque gladio qui descenderunt incircumcisi ad terram ultimam qui posuerunt terrorem suum in terra viventium et portaverunt ignominiam suam cum his qui descendunt in lacum
EZEK|32|25|in medio interfectorum posuerunt cubile eius in universis populis eius in circuitu eius sepulchrum illius omnes hii incircumcisi interfectique gladio dederant enim terrorem in terra viventium et portaverunt ignominiam suam cum his qui descendunt in lacum in medio interfectorum positi sunt
EZEK|32|26|ibi Mosoch et Thubal et omnis multitudo eius in circuitu illius sepulchra eius omnes hii incircumcisi interfectique et cadentes gladio quia dederunt formidinem suam in terra viventium
EZEK|32|27|et non dormient cum fortibus cadentibusque et incircumcisis qui descenderunt ad infernum cum armis suis et posuerunt gladios suos sub capitibus suis et fuerunt iniquitates eorum in ossibus eorum quia terror fortium facti sunt in terra viventium
EZEK|32|28|et tu ergo in medio incircumcisorum contereris et dormies cum interfectis gladio
EZEK|32|29|ibi Idumea et reges eius omnes duces eius qui dati sunt cum exercitu suo cum interfectis gladio et qui cum incircumcisis dormierunt et cum his qui descenderunt in lacum
EZEK|32|30|ibi principes aquilonis omnes et universi venatores qui deducti sunt cum interfectis paventes et in sua fortitudine confusi qui dormierunt incircumcisi cum interfectis gladio et portaverunt confusionem suam cum his qui descendunt in lacum
EZEK|32|31|vidit eos Pharao et consolatus est super universa multitudine sua quae interfecta est gladio Pharao et omnis exercitus eius ait Dominus Deus
EZEK|32|32|quia dedi terrorem meum in terra viventium et dormivit in medio incircumcisorum cum interfectis gladio Pharao et omnis multitudo eius ait Dominus Deus
EZEK|33|1|et factum est verbum Domini ad me dicens
EZEK|33|2|fili hominis loquere ad filios populi tui et dices ad eos terra cum induxero super eam gladium et tulerit populus terrae virum unum de novissimis suis et constituerit eum super se speculatorem
EZEK|33|3|et ille viderit gladium venientem super terram et cecinerit bucina et adnuntiaverit populo
EZEK|33|4|audiens autem quisquis ille est sonum bucinae non se observaverit veneritque gladius et tulerit eum sanguis ipsius super caput eius erit
EZEK|33|5|sonum bucinae audivit et non se observavit sanguis eius in ipso erit si autem custodierit animam suam salvavit
EZEK|33|6|quod si speculator viderit gladium venientem et non insonuerit bucina et populus non se custodierit veneritque gladius et tulerit de eis animam ille quidem in iniquitate sua captus est sanguinem autem eius de manu speculatoris requiram
EZEK|33|7|et tu fili hominis speculatorem dedi te domui Israhel audiens ergo ex ore meo sermonem adnuntiabis eis ex me
EZEK|33|8|si me dicente ad impium impie morte morieris non fueris locutus ut se custodiat impius a via sua ipse impius in iniquitate sua morietur sanguinem autem eius de manu tua requiram
EZEK|33|9|si autem adnuntiante te ad impium ut a viis suis convertatur non fuerit conversus a via sua ipse in iniquitate sua morietur porro tu animam tuam liberasti
EZEK|33|10|tu ergo fili hominis dic ad domum Israhel sic locuti estis dicentes iniquitates nostrae et peccata nostra super nos sunt et in ipsis nos tabescimus quomodo ergo vivere poterimus
EZEK|33|11|dic ad eos vivo ego dicit Dominus Deus nolo mortem impii sed ut revertatur impius a via sua et vivat convertimini a viis vestris pessimis et quare moriemini domus Israhel
EZEK|33|12|tu itaque fili hominis dic ad filios populi tui iustitia iusti non liberabit eum in quacumque die peccaverit et impietas impii non nocebit ei in quacumque die conversus fuerit ab impietate sua et iustus non poterit vivere in iustitia sua in quacumque die peccaverit
EZEK|33|13|etiam si dixero iusto quod vita vivat et confisus in iustitia sua fecerit iniquitatem omnes iustitiae eius oblivioni tradentur et in iniquitate sua quam operatus est in ipsa morietur
EZEK|33|14|sin autem dixero impio morte morieris et egerit paenitentiam a peccato suo feceritque iudicium et iustitiam
EZEK|33|15|pignus restituerit ille impius rapinamque reddiderit in mandatis vitae ambulaverit nec fecerit quicquam iniustum vita vivet et non morietur
EZEK|33|16|omnia peccata eius quae peccavit non inputabuntur ei iudicium et iustitiam fecit vita vivet
EZEK|33|17|et dixerunt filii populi tui non est aequi ponderis via Domini et ipsorum via iniusta est
EZEK|33|18|cum enim recesserit iustus a iustitia sua feceritque iniquitatem morietur in eis
EZEK|33|19|et cum recesserit impius ab impietate sua feceritque iudicium et iustitiam vivet in eis
EZEK|33|20|et dicitis non est recta via Domini unumquemque iuxta vias suas iudicabo de vobis domus Israhel
EZEK|33|21|et factum est in duodecimo anno in duodecimo mense in quinta mensis transmigrationis nostrae venit ad me qui fugerat de Hierusalem dicens vastata est civitas
EZEK|33|22|manus autem Domini facta fuerat ad me vespere antequam veniret qui fugerat aperuitque os meum donec veniret ad me mane et aperto ore meo non silui amplius
EZEK|33|23|et factum est verbum Domini ad me dicens
EZEK|33|24|fili hominis qui habitant in ruinosis his super humum Israhel loquentes aiunt unus erat Abraham et hereditate possedit terram nos autem multi nobis data est terra in possessionem
EZEK|33|25|idcirco dices ad eos haec dicit Dominus Deus qui in sanguine comeditis et oculos vestros levatis ad inmunditias vestras et sanguinem funditis numquid terram hereditate possidebitis
EZEK|33|26|stetistis in gladiis vestris fecistis abominationes et unusquisque uxorem proximi sui polluit et terram hereditate possidebitis
EZEK|33|27|haec dices ad eos sic dicit Dominus Deus vivo ego quia qui in ruinosis habitant gladio cadent et qui in agro est bestiis tradetur ad devorandum qui autem in praesidiis et in speluncis sunt peste morientur
EZEK|33|28|et dabo terram in solitudinem et desertum et deficiet superba fortitudo eius et desolabuntur montes Israhel eo quod nullus sit qui per eos transeat
EZEK|33|29|et scient quia ego Dominus cum dedero terram desolatam et desertam propter universas abominationes suas quas operati sunt
EZEK|33|30|et tu fili hominis filii populi tui qui loquuntur de te iuxta muros et in ostiis domorum et dicunt unus ad alterum vir ad proximum suum loquentes venite et audiamus qui sit sermo egrediens a Domino
EZEK|33|31|et veniunt ad te quasi si ingrediatur populus et sedent coram te populus meus et audiunt sermones tuos et non faciunt eos quia in canticum oris sui vertunt illos et avaritiam suam sequitur cor eorum
EZEK|33|32|et es eis quasi carmen musicum quod suavi dulcique sono canitur et audient verba tua et non facient ea
EZEK|33|33|et cum venerit quod praedictum est ecce enim venit tunc scient quod prophetes fuerit inter eos
EZEK|34|1|et factum est verbum Domini ad me dicens
EZEK|34|2|fili hominis propheta de pastoribus Israhel propheta et dices pastoribus haec dicit Dominus Deus vae pastoribus Israhel qui pascebant semet ipsos nonne greges pascuntur a pastoribus
EZEK|34|3|lac comedebatis et lanis operiebamini et quod crassum erat occidebatis gregem autem meum non pascebatis
EZEK|34|4|quod infirmum fuit non consolidastis et quod aegrotum non sanastis quod fractum est non alligastis et quod abiectum est non reduxistis quod perierat non quaesistis sed cum austeritate imperabatis eis et cum potentia
EZEK|34|5|et dispersae sunt oves meae eo quod non esset pastor et factae sunt in devorationem omnium bestiarum agri et dispersae sunt
EZEK|34|6|erraverunt greges mei in cunctis montibus et in universo colle excelso et super omnem faciem terrae dispersi sunt greges mei et non erat qui requireret non erat inquam qui requireret
EZEK|34|7|propterea pastores audite verbum Domini
EZEK|34|8|vivo ego dicit Dominus Deus quia pro eo quod facti sunt greges mei in rapinam et oves meae in devorationem omnium bestiarum agri eo quod non esset pastor neque enim quaesierunt pastores gregem meum sed pascebant pastores semet ipsos et greges meos non pascebant
EZEK|34|9|propterea pastores audite verbum Domini
EZEK|34|10|haec dicit Dominus Deus ecce ego ipse super pastores requiram gregem meum de manu eorum et cessare eos faciam ut ultra non pascant gregem nec pascant amplius pastores semet ipsos et liberabo gregem meum de ore eorum et non erunt ultra eis in escam
EZEK|34|11|quia haec dicit Dominus Deus ecce ego ipse requiram oves meas et visitabo eas
EZEK|34|12|sicut visitat pastor gregem suum in die quando fuerit in medio ovium suarum dissipatarum sic visitabo oves meas et liberabo eas de omnibus locis quo dispersae fuerant in die nubis et caliginis
EZEK|34|13|et educam eas de populis et congregabo eas de terris et inducam eas in terram suam et pascam eas in montibus Israhel in rivis et in cunctis sedibus terrae
EZEK|34|14|in pascuis uberrimis pascam eas et in montibus excelsis Israhel erunt pascuae eorum ibi requiescent in herbis virentibus et in pascuis pinguibus pascentur super montes Israhel
EZEK|34|15|ego pascam oves meas et ego eas accubare faciam dicit Dominus Deus
EZEK|34|16|quod perierat requiram et quod abiectum erat reducam et quod confractum fuerat alligabo et quod infirmum erat consolidabo et quod pingue et forte custodiam et pascam illas in iudicio
EZEK|34|17|vos autem greges mei haec dicit Dominus Deus ecce ego iudico inter pecus et pecus arietum et hircorum
EZEK|34|18|nonne satis vobis erat pascuam bonam depasci insuper et reliquias pascuarum vestrarum conculcastis pedibus vestris et cum purissimam aquam biberetis reliquam pedibus vestris turbabatis
EZEK|34|19|et oves meae his quae conculcata pedibus vestris fuerant pascebantur et quae pedes vestri turbaverant haec bibebant
EZEK|34|20|propterea haec dicit Dominus Deus ad eos ecce ego ipse iudico inter pecus pingue et macilentum
EZEK|34|21|pro eo quod lateribus et umeris inpingebatis et cornibus vestris ventilabatis omnia infirma pecora donec dispergerentur foras
EZEK|34|22|salvabo gregem meum et non erit ultra in rapinam et iudicabo inter pecus et pecus
EZEK|34|23|et suscitabo super ea pastorem unum qui pascat ea servum meum David ipse pascet ea et ipse erit eis in pastorem
EZEK|34|24|ego autem Dominus ero eis in Deum et servus meus David princeps in medio eorum ego Dominus locutus sum
EZEK|34|25|et faciam cum eis pactum pacis et cessare faciam bestias pessimas de terra et qui habitant in deserto securi dormient in saltibus
EZEK|34|26|et ponam eos in circuitu collis mei benedictionem et deducam imbrem in tempore suo pluviae benedictionis erunt
EZEK|34|27|et dabit lignum agri fructum suum et terra dabit germen suum et erunt in terra sua absque timore et scient quia ego Dominus cum contrivero catenas iugi eorum et eruero eos de manu imperantium sibi
EZEK|34|28|et non erunt ultra in rapinam gentibus neque bestiae terrae devorabunt eos sed habitabunt confidenter absque ullo terrore
EZEK|34|29|et suscitabo eis germen nominatum et non erunt ultra inminuti fame in terra neque portabunt amplius obprobria gentium
EZEK|34|30|et scient quia ego Dominus Deus eorum cum eis et ipsi populus meus domus Israhel ait Dominus Deus
EZEK|34|31|vos autem greges mei greges pascuae meae homines estis et ego Dominus Deus vester dicit Dominus Deus
EZEK|35|1|et factus est sermo Domini ad me dicens
EZEK|35|2|fili hominis pone faciem tuam adversum montem Seir et prophetabis de eo et dices illi
EZEK|35|3|haec dicit Dominus Deus ecce ego ad te mons Seir et extendam manum meam super te et dabo te desolatum atque desertum
EZEK|35|4|urbes tuas demoliar et tu desertus eris et scies quia ego Dominus
EZEK|35|5|eo quod fueris inimicus sempiternus et concluseris filios Israhel in manus gladii in tempore adflictionis eorum in tempore iniquitatis extremae
EZEK|35|6|propterea vivo ego dicit Dominus Deus quoniam sanguini tradam te et sanguis te persequetur et cum sanguinem oderis sanguis persequetur te
EZEK|35|7|et dabo montem Seir desolatum et desertum et auferam de eo euntem et redeuntem
EZEK|35|8|et implebo montes eius occisorum suorum in collibus tuis et in vallibus tuis atque in torrentibus interfecti gladio cadent
EZEK|35|9|in solitudines sempiternas tradam te et civitates tuae non habitabuntur et scietis quoniam ego Dominus
EZEK|35|10|eo quod dixeris duae gentes et duae terrae meae erunt et hereditate possidebo eas cum Dominus esset ibi
EZEK|35|11|propterea vivo ego dicit Dominus Deus quia faciam iuxta iram tuam et secundum zelum tuum quem fecisti odio habens eos et notus efficiar per eos cum te iudicavero
EZEK|35|12|et scies quia ego Dominus audivi universa obprobria tua quae locutus es de montibus Israhel dicens deserti nobis dati sunt ad devorandum
EZEK|35|13|et insurrexistis super me ore vestro et rogastis adversum me verba vestra ego audivi
EZEK|35|14|haec dicit Dominus Deus laetante universa terra in solitudinem te redigam
EZEK|35|15|sicuti gavisus es super hereditatem domus Israhel eo quod fuerit dissipata sic faciam tibi dissipatus eris mons Seir et Idumea omnis et scient quia ego Dominus
EZEK|36|1|tu autem fili hominis propheta super montes Israhel et dices montes Israhel audite verbum Domini
EZEK|36|2|haec dicit Dominus Deus eo quod dixerit inimicus de vobis euge altitudines sempiternae in hereditatem datae sunt nobis
EZEK|36|3|propterea vaticinare et dic haec dicit Dominus Deus pro eo quod desolati estis et conculcati per circuitum et facti in hereditatem reliquis gentibus et ascendistis super labium linguae et obprobrium populi
EZEK|36|4|propterea montes Israhel audite verbum Domini Dei haec dicit Dominus Deus montibus et collibus torrentibus vallibusque et desertis parietinis et urbibus derelictis quae depopulatae sunt et subsannatae a reliquis gentibus per circuitum
EZEK|36|5|propterea haec dicit Dominus Deus quoniam in igne zeli mei locutus sum de reliquis gentibus et de Idumea universa qui dederunt terram meam sibi in hereditatem cum gaudio et toto corde ex animo et eiecerunt eam ut vastarent
EZEK|36|6|idcirco vaticinare super humum Israhel et dices montibus et collibus iugis et vallibus haec dicit Dominus Deus ecce ego in zelo meo et in furore meo locutus sum eo quod confusionem gentium sustinueritis
EZEK|36|7|idcirco haec dicit Dominus Deus ego levavi manum meam ut gentes quae in circuitu vestro sunt ipsae confusionem suam portent
EZEK|36|8|vos autem montes Israhel ramos vestros germinetis et fructum vestrum adferatis populo meo Israhel prope est enim ut veniat
EZEK|36|9|quia ecce ego ad vos et convertar ad vos et arabimini et accipietis sementem
EZEK|36|10|et multiplicabo in vobis homines omnemque domum Israhel et habitabuntur civitates et ruinosa instaurabuntur
EZEK|36|11|et replebo vos hominibus et iumentis et multiplicabuntur et crescent et habitari vos faciam sicut a principio bonisque donabo maioribus quam habuistis ab initio et scietis quia ego Dominus
EZEK|36|12|et adducam super vos homines populum meum Israhel et hereditate possidebunt te et eris eis in hereditatem et non addes ultra ut absque eis sis
EZEK|36|13|haec dicit Dominus Deus pro eo quod dicunt de vobis devoratrix hominum es et suffocans gentem tuam
EZEK|36|14|propterea homines non comedes amplius et gentem tuam non necabis ultra ait Dominus Deus
EZEK|36|15|nec auditam faciam in te amplius confusionem gentium et obprobrium populorum nequaquam portabis et gentem tuam non amittes amplius ait Dominus Deus
EZEK|36|16|et factum est verbum Domini ad me dicens
EZEK|36|17|fili hominis domus Israhel habitaverunt in humo sua et polluerunt eam in viis suis et in studiis suis iuxta inmunditiam menstruatae facta est via eorum coram me
EZEK|36|18|et effudi indignationem meam super eos pro sanguine quem fuderunt super terram et in idolis suis polluerunt eam
EZEK|36|19|et dispersi eos in gentes et ventilati sunt in terris iuxta vias eorum et adinventiones iudicavi eos
EZEK|36|20|et ingressi sunt ad gentes ad quas introierunt et polluerunt nomen sanctum meum cum diceretur de eis populus Domini iste est et de terra eius egressi sunt
EZEK|36|21|et peperci nomini meo sancto quod polluerat domus Israhel in gentibus ad quas ingressi sunt
EZEK|36|22|idcirco dices domui Israhel haec dicit Dominus Deus non propter vos ego faciam domus Israhel sed propter nomen sanctum meum quod polluistis in gentibus ad quas intrastis
EZEK|36|23|et sanctificabo nomen meum magnum quod pollutum est inter gentes quod polluistis in medio earum ut sciant gentes quia ego Dominus ait Dominus exercituum cum sanctificatus fuero in vobis coram eis
EZEK|36|24|tollam quippe vos de gentibus et congregabo de universis terris et adducam vos in terram vestram
EZEK|36|25|et effundam super vos aquam mundam et mundabimini ab omnibus inquinamentis vestris et ab universis idolis vestris mundabo vos
EZEK|36|26|et dabo vobis cor novum et spiritum novum ponam in medio vestri et auferam cor lapideum de carne vestra et dabo vobis cor carneum
EZEK|36|27|et spiritum meum ponam in medio vestri et faciam ut in praeceptis meis ambuletis et iudicia mea custodiatis et operemini
EZEK|36|28|et habitabitis in terra quam dedi patribus vestris et eritis mihi in populum et ego ero vobis in Deum
EZEK|36|29|et salvabo vos ex universis inquinamentis vestris et vocabo frumentum et multiplicabo illud et non inponam in vobis famem
EZEK|36|30|et multiplicabo fructum ligni et genimina agri ut non portetis ultra obprobrium famis in gentibus
EZEK|36|31|et recordabimini viarum vestrarum pessimarum studiorumque non bonorum et displicebunt vobis iniquitates vestrae et scelera vestra
EZEK|36|32|non propter vos ego faciam ait Dominus Deus notum sit vobis confundimini et erubescite super viis vestris domus Israhel
EZEK|36|33|haec dicit Dominus Deus in die qua mundavero vos ex omnibus iniquitatibus vestris et habitari fecero urbes et instauravero ruinosa
EZEK|36|34|et terra deserta fuerit exculta quae quondam erat desolata in oculis omnis viatoris
EZEK|36|35|dicent terra illa inculta facta est ut hortus voluptatis et civitates desertae et destitutae atque suffossae munitae sederunt
EZEK|36|36|et scient gentes quaecumque derelictae fuerint in circuitu vestro quia ego Dominus aedificavi dissipata plantavique inculta ego Dominus locutus sum et fecerim
EZEK|36|37|haec dicit Dominus Deus adhuc in hoc invenient me domus Israhel ut faciam eis multiplicabo eos sicut gregem hominum
EZEK|36|38|ut gregem sanctum ut gregem Hierusalem in sollemnitatibus eius sic erunt civitates desertae plenaeque gregibus hominum et scient quia ego Dominus
EZEK|37|1|facta est super me manus Domini et eduxit me in spiritu Domini et dimisit me in medio campi qui erat plenus ossibus
EZEK|37|2|et circumduxit me per ea in gyro erant autem multa valde super faciem campi siccaque vehementer
EZEK|37|3|et dixit ad me fili hominis putasne vivent ossa ista et dixi Domine Deus tu nosti
EZEK|37|4|et dixit ad me vaticinare de ossibus istis et dices eis ossa arida audite verbum Domini
EZEK|37|5|haec dicit Dominus Deus ossibus his ecce ego intromittam in vos spiritum et vivetis
EZEK|37|6|et dabo super vos nervos et succrescere faciam super vos carnes et superextendam in vobis cutem et dabo vobis spiritum et vivetis et scietis quia ego Dominus
EZEK|37|7|et prophetavi sicut praeceperat mihi factus est autem sonitus prophetante me et ecce commotio et accesserunt ossa ad ossa unumquodque ad iuncturam suam
EZEK|37|8|et vidi et ecce super ea nervi et carnes ascenderunt et extenta est in eis cutis desuper et spiritum non habebant
EZEK|37|9|et dixit ad me vaticinare ad spiritum vaticinare fili hominis et dices ad spiritum haec dicit Dominus Deus a quattuor ventis veni spiritus et insufla super interfectos istos et revivescant
EZEK|37|10|et prophetavi sicut praeceperat mihi et ingressus est in ea spiritus et vixerunt steteruntque super pedes suos exercitus grandis nimis valde
EZEK|37|11|et dixit ad me fili hominis ossa haec universa domus Israhel est ipsi dicunt aruerunt ossa nostra et periit spes nostra et abscisi sumus
EZEK|37|12|propterea vaticinare et dices ad eos haec dicit Dominus Deus ecce ego aperiam tumulos vestros et educam vos de sepulchris vestris populus meus et inducam vos in terram Israhel
EZEK|37|13|et scietis quia ego Dominus cum aperuero sepulchra vestra et eduxero vos de tumulis vestris populus meus
EZEK|37|14|et dedero spiritum meum in vobis et vixeritis et requiescere vos faciam super humum vestram et scietis quia ego Dominus locutus sum et feci ait Dominus Deus
EZEK|37|15|et factus est sermo Domini ad me dicens
EZEK|37|16|et tu fili hominis sume tibi lignum unum et scribe super illud Iudae et filiorum Israhel sociis eius et tolle lignum alterum et scribe super eum Ioseph lignum Ephraim et cunctae domui Israhel sociorumque eius
EZEK|37|17|et adiunge illa unum ad alterum tibi in lignum unum et erunt in unionem in manu tua
EZEK|37|18|cum autem dixerint ad te filii populi tui loquentes nonne indicas nobis quid in his tibi velis
EZEK|37|19|loqueris ad eos haec dicit Dominus Deus ecce ego adsumam lignum Ioseph quod est in manu Ephraim et tribus Israhel quae iunctae sunt ei et dabo eas pariter cum ligno Iuda et faciam eas in lignum unum et erunt unum in manu eius
EZEK|37|20|erunt autem ligna super quae scripseris in manu tua in oculis eorum
EZEK|37|21|et dices ad eos haec dicit Dominus Deus ecce ego adsumam filios Israhel de medio nationum ad quas abierunt et congregabo eos undique et adducam eos ad humum suam
EZEK|37|22|et faciam eos gentem unam in terra in montibus Israhel et rex unus erit omnibus imperans et non erunt ultra duae gentes nec dividentur amplius in duo regna
EZEK|37|23|neque polluentur ultra in idolis suis et abominationibus suis et in cunctis iniquitatibus suis et salvos eos faciam de universis sedibus suis in quibus peccaverunt et mundabo eos et erunt mihi populus et ego ero eis Deus
EZEK|37|24|et servus meus David rex super eos et pastor unus erit omnium eorum in iudiciis meis ambulabunt et mandata mea custodient et facient ea
EZEK|37|25|et habitabunt super terram quam dedi servo meo Iacob in qua habitaverunt patres vestri et habitabunt super eam ipsi et filii eorum et filii filiorum eorum usque in sempiternum et David servus meus princeps eorum in perpetuum
EZEK|37|26|et percutiam illis foedus pacis pactum sempiternum erit eis et fundabo eos et multiplicabo et dabo sanctificationem meam in medio eorum in perpetuum
EZEK|37|27|et erit tabernaculum meum in eis et ero eis Deus et ipsi erunt mihi populus
EZEK|37|28|et scient gentes quia ego Dominus sanctificator Israhel cum fuerit sanctificatio mea in medio eorum in perpetuum
EZEK|38|1|et factus est sermo Domini ad me dicens
EZEK|38|2|fili hominis pone faciem tuam contra Gog terram Magog principem capitis Mosoch et Thubal et vaticinare de eo
EZEK|38|3|et dices ad eum haec dicit Dominus Deus ecce ego ad te Gog principem capitis Mosoch et Thubal
EZEK|38|4|et circumagam te et ponam frenum in maxillis tuis et educam te et omnem exercitum tuum equos et equites vestitos loricis universos multitudinem magnam hastam et clypeum arripientium et gladium
EZEK|38|5|Persae Aethiopes et Lybies cum eis omnes scutati et galeati
EZEK|38|6|Gomer et universa agmina eius domus Thogorma latera aquilonis et totum robur eius populique multi tecum
EZEK|38|7|praepara et instrue te et omnem multitudinem tuam quae coacervata est ad te et esto eis in praeceptum
EZEK|38|8|post dies multos visitaberis in novissimo annorum venies ad terram quae reversa est a gladio congregata est de populis multis ad montes Israhel qui fuerunt deserti iugiter haec de populis educta est et habitaverunt in ea confidenter universi
EZEK|38|9|ascendens autem quasi tempestas venies et quasi nubes ut operias terram tu et omnia agmina tua et populi multi tecum
EZEK|38|10|haec dicit Dominus Deus in die illa ascendent sermones super cor tuum et cogitabis cogitationem pessimam
EZEK|38|11|et dices ascendam ad terram absque muro veniam ad quiescentes habitantesque secure omnes habitant sine muro vectes et portae non sunt eis
EZEK|38|12|ut diripias spolia et invadas praedam ut inferas manum tuam super eos qui deserti fuerant et postea restituti et super populum qui est congregatus ex gentibus qui possidere coepit et esse habitator umbilici terrae
EZEK|38|13|Seba et Dedan et negotiatores Tharsis et omnes leones eius dicent tibi numquid ad sumenda spolia tu venis ecce ad diripiendam praedam congregasti multitudinem tuam ut tollas argentum et aurum auferas supellectilem atque substantiam et diripias manubias infinitas
EZEK|38|14|propterea vaticinare fili hominis et dices ad Gog haec dicit Dominus Deus numquid non in die illo cum habitaverit populus meus Israhel confidenter scies
EZEK|38|15|et venies de loco tuo a lateribus aquilonis tu et populi multi tecum ascensores equorum universi coetus magnus et exercitus vehemens
EZEK|38|16|et ascendes super populum meum Israhel quasi nubes ut operias terram in novissimis diebus eris et adducam te super terram meam ut sciant gentes me cum sanctificatus fuero in te in oculis eorum o Gog
EZEK|38|17|haec dicit Dominus Deus tu ergo ille es de quo locutus sum in diebus antiquis in manu servorum meorum prophetarum Israhel qui prophetaverunt in diebus illorum temporum ut adducerem te super eos
EZEK|38|18|et erit in die illa in die adventus Gog super terram Israhel ait Dominus Deus ascendet indignatio mea in furore meo
EZEK|38|19|et in zelo meo in igne irae meae locutus sum quia in die illa erit commotio magna super terram Israhel
EZEK|38|20|et commovebuntur a facie mea pisces maris et volucres caeli et bestiae agri et omne reptile quod movetur super humum cunctique homines qui sunt super faciem terrae et subvertentur montes et cadent sepes et omnis murus in terra corruet
EZEK|38|21|et convocabo adversum eum in cunctis montibus meis gladium ait Dominus Deus gladius uniuscuiusque in fratrem suum dirigetur
EZEK|38|22|et iudicabo eum peste et sanguine et imbre vehementi et lapidibus inmensis ignem et sulphur pluam super eum et super exercitum eius et super populos multos qui sunt cum eo
EZEK|38|23|et magnificabor et sanctificabor et notus ero in oculis gentium multarum et scient quia ego Dominus
EZEK|39|1|tu autem fili hominis vaticinare adversum Gog et dices haec dicit Dominus Deus ecce ego super te Gog principem capitis Mosoch et Thubal
EZEK|39|2|et circumagam te et seducam te et ascendere faciam de lateribus aquilonis et adducam te super montes Israhel
EZEK|39|3|et percutiam arcum tuum in manu sinistra tua et sagittas tuas de manu dextera tua deiciam
EZEK|39|4|super montes Israhel cades tu et omnia agmina tua et populi qui sunt tecum feris avibus omnique volatili et bestiis terrae dedi te devorandum
EZEK|39|5|super faciem agri cades quia ego locutus sum ait Dominus Deus
EZEK|39|6|et emittam ignem in Magog et in his qui habitant in insulis confidenter et scient quia ego Dominus
EZEK|39|7|et nomen sanctum meum notum faciam in medio populi mei Israhel et non polluam nomen sanctum meum amplius et scient gentes quia ego Dominus Sanctus Israhel
EZEK|39|8|ecce venit et factum est ait Dominus Deus haec est dies de qua locutus sum
EZEK|39|9|et egredientur habitatores de civitatibus Israhel et succendent et conburent arma clypeum et hastas arcum et sagittas et baculos manus et contos et succendent ea igne septem annis
EZEK|39|10|et non portabunt ligna de regionibus neque succident de saltibus quoniam arma succendent igne et depraedabuntur eos quibus praedae fuerant et diripient vastatores suos ait Dominus Deus
EZEK|39|11|et erit in die illa dabo Gog locum nominatum sepulchrum in Israhel vallem Viatorum ad orientem maris quae obstupescere facit praetereuntes et sepelient ibi Gog et omnem multitudinem eius et vocabitur vallis Multitudinis Gog
EZEK|39|12|et sepelient eos domus Israhel ut mundent terram septem mensibus
EZEK|39|13|sepeliet autem omnis populus terrae et erit eis nominata dies in qua glorificatus sum ait Dominus Deus
EZEK|39|14|et viros iugiter constituent lustrantes terram qui sepeliant et requirant eos qui remanserant super faciem terrae ut emundent eam post menses autem septem quaerere incipient
EZEK|39|15|et circumibunt peragrantes terram cumque viderint os hominis statuent iuxta illud titulum donec sepeliant illud pollinctores in valle Multitudinis Gog
EZEK|39|16|nomen autem civitatis Amona et mundabunt terram
EZEK|39|17|tu ergo fili hominis haec dicit Dominus Deus dic omni volucri et universis avibus cunctisque bestiis agri convenite properate concurrite undique ad victimam meam quam ego immolo vobis victimam grandem super montes Israhel ut comedatis carnes et bibatis sanguinem
EZEK|39|18|carnes fortium comedetis et sanguinem principum terrae bibetis arietum agnorum et hircorum taurorumque altilium et pinguium omnium
EZEK|39|19|et comedetis adipem in saturitate et bibetis sanguinem in ebrietate de victima quam ego immolabo vobis
EZEK|39|20|et saturabimini super mensam meam de equo et de equite forti et de universis viris bellatoribus ait Dominus Deus
EZEK|39|21|et ponam gloriam meam in gentibus et videbunt omnes gentes iudicium meum quod fecerim et manum meam quam posuerim super eos
EZEK|39|22|et scient domus Israhel quia ego Dominus Deus eorum a die illa et deinceps
EZEK|39|23|et scient gentes quoniam in iniquitate sua capta sit domus Israhel eo quod reliquerint me et absconderim faciem meam ab eis et tradiderim eos in manu hostium et ceciderint in gladio universi
EZEK|39|24|iuxta inmunditiam eorum et scelus feci eis et abscondi faciem meam ab illis
EZEK|39|25|propterea haec dicit Dominus Deus nunc reducam captivitatem Iacob et miserebor omnis domus Israhel et adsumam zelum pro nomine sancto meo
EZEK|39|26|et portabunt confusionem suam et omnem praevaricationem quam praevaricati sunt in me cum habitaverint in terra sua confidenter neminem formidantes
EZEK|39|27|et reduxero eos de populis et congregavero de terris inimicorum suorum et sanctificatus fuero in eis in oculis gentium plurimarum
EZEK|39|28|et scient quia ego Dominus Deus eorum eo quod transtulerim eos in nationes et congregavero eos super terram suam et non dereliquerim quemquam ex eis ibi
EZEK|39|29|et non abscondam ultra faciem meam ab eis eo quod effuderim spiritum meum super omnem domum Israhel ait Dominus Deus
EZEK|40|1|in vicesimo et quinto anno transmigrationis nostrae in exordio anni decima mensis quartodecimo anno postquam percussa est civitas in ipsa hac die facta est super me manus Domini et adduxit me illuc
EZEK|40|2|in visionibus Dei adduxit me in terram Israhel et dimisit me super montem excelsum nimis super quem erat quasi aedificium civitatis vergentis ad austrum
EZEK|40|3|et introduxit me illuc et ecce vir cuius erat species quasi species aeris et funiculus lineus in manu eius et calamus mensurae in manu eius stabat autem in porta
EZEK|40|4|et locutus est ad me idem vir fili hominis vide oculis tuis et auribus tuis audi et pone cor tuum in omnia quae ego ostendam tibi quia ut ostendantur tibi adductus es huc adnuntia omnia quae tu vides domui Israhel
EZEK|40|5|et ecce murus forinsecus in circuitu domus undique et in manu viri calamus mensurae sex cubitorum et palmo et mensus est latitudinem aedificii calamo uno altitudinem quoque calamo uno
EZEK|40|6|et venit ad portam quae respiciebat viam orientalem et ascendit per gradus eius et mensus est limen portae calamo uno latitudinem id est limen unum calamo uno in latitudine
EZEK|40|7|et thalamum uno calamo in longum et uno calamo in latum et inter thalamos quinque cubitos
EZEK|40|8|et limen portae iuxta vestibulum portae intrinsecus calamo uno
EZEK|40|9|et mensus est vestibulum portae octo cubitorum et frontem eius duobus cubitis vestibulum autem portae erat intrinsecus
EZEK|40|10|porro thalami portae ad viam orientalem tres hinc et tres inde mensura una trium et mensura una frontium ex utraque parte
EZEK|40|11|et mensus est latitudinem liminis portae decem cubitorum et longitudinem portae tredecim cubitorum
EZEK|40|12|et marginem ante thalamos cubiti unius et cubitus unus finis utrimque thalami autem sex cubitorum erant hinc et inde
EZEK|40|13|et mensus est portam a tecto thalami usque ad tectum eius latitudinem viginti et quinque cubitorum ostium contra ostium
EZEK|40|14|et fecit frontes per sexaginta cubitos et ad frontem atrium portae undique per circuitum
EZEK|40|15|et ante faciem portae quae pertingebat usque ad faciem vestibuli portae interioris quinquaginta cubitos
EZEK|40|16|et fenestras obliquas in thalamis et in frontibus eorum quae erant intra portam undique per circuitum similiter autem erant et in vestibulis fenestrae per gyrum intrinsecus et ante frontes pictura palmarum
EZEK|40|17|et eduxit me ad atrium exterius et ecce gazofilacia et pavimentum stratum lapide in atrio per circuitum triginta gazofilacia in circuitu pavimenti
EZEK|40|18|et pavimentum in fronte portarum secundum longitudinem portarum erat inferius
EZEK|40|19|et mensus est latitudinem a facie portae inferioris usque ad frontem atrii interioris extrinsecus centum cubitos ad orientem et ad aquilonem
EZEK|40|20|portam quoque quae respiciebat viam aquilonis atrii exterioris mensus est tam in longitudine quam in latitudine
EZEK|40|21|et thalamos eius tres hinc et tres inde et frontem eius et vestibulum eius secundum mensuram portae prioris quinquaginta cubitorum longitudinem eius et latitudinem viginti quinque cubitorum
EZEK|40|22|fenestrae autem eius et vestibulum et scalpturae secundum mensuram portae quae respiciebat ad orientem et septem graduum erat ascensus eius et vestibulum ante eam
EZEK|40|23|et porta atrii interioris contra portam aquilonis et orientalem et mensus est a porta usque ad portam centum cubitos
EZEK|40|24|et duxit me ad viam australem et ecce porta quae respiciebat ad austrum et mensus est frontem eius et vestibulum eius iuxta mensuras superiores
EZEK|40|25|et fenestras eius et vestibula in circuitu sicut fenestras ceteras quinquaginta cubitorum longitudine et latitudine viginti quinque cubitorum
EZEK|40|26|et in gradibus septem ascendebatur ad eam et vestibulum ante fores eius et celatae palmae erant una hinc et altera inde in fronte eius
EZEK|40|27|et porta atrii interioris in via australi et mensus est a porta usque ad portam in via australi centum cubitos
EZEK|40|28|et introduxit me in atrium interius ad portam australem et mensus est portam iuxta mensuras superiores
EZEK|40|29|thalamum eius et frontem eius et vestibulum eius hisdem mensuris et fenestras eius et vestibulorum eius in circuitu quinquaginta cubitos longitudinis et latitudinis viginti quinque cubitos
EZEK|40|30|et vestibulum per gyrum longitudine viginti quinque cubitorum et latitudine quinque cubitorum
EZEK|40|31|et vestibulum eius ad atrium exterius et palmas eius in fronte et octo gradus erant quibus ascendebatur per eam
EZEK|40|32|et introduxit me in atrium interius per viam orientalem et mensus est portam secundum mensuras superiores
EZEK|40|33|thalamum eius et frontem eius et vestibula eius sicut supra et fenestras eius et vestibuli eius in circuitu longitudine quinquaginta cubitorum et latitudine viginti quinque cubitorum
EZEK|40|34|et vestibulum eius id est atrii exterioris et palmae celatae in fronte eius hinc et inde et in octo gradibus ascensus eius
EZEK|40|35|et introduxit me ad portam quae respiciebat ad aquilonem et mensus est secundum mensuras superiores
EZEK|40|36|thalamum eius frontem eius vestibulum eius et fenestras eius per circuitum longitudine quinquaginta cubitorum et latitudine viginti quinque cubitorum
EZEK|40|37|vestibulum eius in atrium exterius et celatura palmarum in fronte illius hinc et inde et in octo gradibus ascensus eius
EZEK|40|38|et per singula gazofilacia ostium in frontibus portarum ibi lavabunt holocaustum
EZEK|40|39|et in vestibulo portae duae mensae hinc et duae mensae inde ut immoletur super eas holocaustum et pro peccato et pro delicto
EZEK|40|40|et ad latus exterius quod ascendit ad ostium portae quae pergit ad aquilonem duae mensae et ad latus alterum ante vestibulum portae duae mensae
EZEK|40|41|quattuor mensae hinc et quattuor mensae inde per latera portae octo mensae erunt super quas immolabunt
EZEK|40|42|quattuor autem mensae ad holocaustum de lapidibus quadris extructae longitudine cubiti unius et dimidii et latitudine cubiti unius et dimidii et altitudine cubiti unius super quas ponant vasa in quibus immolatur holocaustum et victima
EZEK|40|43|et labia earum palmi unius reflexa intrinsecus per circuitum super mensas autem carnes oblationis
EZEK|40|44|et extra portam interiorem gazofilacia cantorum in atrio interiori quod erat in latere portae respicientis ad aquilonem et facies eorum contra viam australem una ex latere portae orientalis quae respiciebat ad viam aquilonis
EZEK|40|45|et dixit ad me hoc est gazofilacium quod respicit viam meridianam sacerdotum qui excubant in custodiis templi
EZEK|40|46|porro gazofilacium quod respicit ad viam aquilonis sacerdotum erit qui excubant ad ministerium altaris isti sunt filii Sadoc qui accedunt de filiis Levi ad Dominum ut ministrent ei
EZEK|40|47|et mensus est atrium longitudine centum cubitorum et latitudine centum cubitorum per quadrum et altare ante faciem templi
EZEK|40|48|et introduxit me in vestibulum templi et mensus est vestibulum quinque cubitis hinc et quinque cubitis inde et latitudinem portae trium cubitorum hinc et trium cubitorum inde
EZEK|40|49|longitudinem autem vestibuli viginti cubitorum et latitudinem undecim cubitorum et octo gradibus ascendebatur ad eam et columnae erant in frontibus una hinc et altera inde
EZEK|41|1|et introduxit me in templum et mensus est frontes sex cubitos latitudinis hinc et sex cubitos latitudinis inde latitudinem tabernaculi
EZEK|41|2|et latitudo portae decem cubitorum erat et latera portae quinque cubitis hinc et quinque cubitis inde et mensus est longitudinem eius quadraginta cubitorum et latitudinem viginti cubitorum
EZEK|41|3|et introgressus intrinsecus mensus est in fronte portae duos cubitos et portam sex cubitorum et latitudinem portae septem cubitorum
EZEK|41|4|et mensus est longitudinem eius viginti cubitorum et latitudinem viginti cubitorum ante faciem templi et dixit ad me hoc est sanctum sanctorum
EZEK|41|5|et mensus est parietem domus sex cubitorum et latitudinem lateris quattuor cubitorum undique per circuitum domus
EZEK|41|6|latera autem latus ad latus bis triginta tria et erant eminentia quae ingrederentur per parietem domus in lateribus per circuitum ut continerent et non adtingerent parietem templi
EZEK|41|7|et platea erat in rotundum ascendens sursum per cocleam et in cenaculum templi deferebat per gyrum idcirco latius erat templum in superioribus et sic de inferioribus ascendebatur ad superiora in medium
EZEK|41|8|et vidi in domo altitudinem per circuitum fundata latera ad mensuram calami sex cubitorum spatio
EZEK|41|9|et latitudinem per parietem lateris forinsecus quinque cubitorum et interior domus in lateribus domus
EZEK|41|10|et inter gazofilacia latitudinem viginti cubitorum in circuitu domus undique
EZEK|41|11|et ostium lateris ad orationem ostium unum ad viam aquilonis et ostium unum ad viam australem et latitudinem loci ad orationem quinque cubitorum in circuitu
EZEK|41|12|et aedificium quod erat separatum versumque ad viam respicientem ad mare latitudinis septuaginta cubitorum paries autem aedificii quinque cubitorum latitudinis per circuitum et longitudo eius nonaginta cubitorum
EZEK|41|13|et mensus est domus longitudinem centum cubitorum et quod separatum erat aedificium et parietes eius longitudinis centum cubitorum
EZEK|41|14|latitudo autem ante faciem domus et eius quod erat separatum contra orientem centum cubitorum
EZEK|41|15|et mensus est longitudinem aedificii contra faciem eius quod erat separatum ad dorsum ekthetas ex utraque parte centum cubitorum et templum interius et vestibula atrii
EZEK|41|16|limina et fenestras obliquas et ekthetas in circuitu per tres partes contra uniuscuiusque limen stratumque ligno per gyrum in circuitu terra autem usque ad fenestras et fenestrae clausae super ostia
EZEK|41|17|et usque ad domum interiorem et forinsecus per omnem parietem in circuitu intrinsecus et forinsecus ad mensuram
EZEK|41|18|et fabrefacta cherubin et palmae et palma inter cherub et cherub duasque facies habebat cherub
EZEK|41|19|faciem hominis iuxta palmam ex hac parte et faciem leonis iuxta palmam ex alia parte expressam per omnem domum in circuitu
EZEK|41|20|de terra usque ad superiora portae cherubin et palmae celatae erant in pariete templi
EZEK|41|21|limen quadrangulum et facies sanctuarii aspectus contra aspectum
EZEK|41|22|altaris lignei trium cubitorum altitudo et longitudo eius duo cubitorum et anguli eius et longitudo eius et parietes eius lignei et locutus est ad me haec est mensa coram Domino
EZEK|41|23|et duo ostia erant in templo et in sanctuario
EZEK|41|24|et in duobus ostiis ex utraque parte bina erant ostiola quae in se invicem plicabantur bina enim ostia erant ex utraque parte ostiorum
EZEK|41|25|et celata erant in ipsis ostiis templi cherubin et scalptura palmarum sicut in parietibus quoque expressa erat quam ob rem erant et grossiora ligna in vestibuli fronte forinsecus
EZEK|41|26|super quae fenestrae obliquae et similitudo palmarum hinc atque inde in umerulis vestibuli secundum latera domus latitudinemque parietum
EZEK|42|1|et eduxit me in atrium exterius per viam ducentem ad aquilonem et eduxit me in gazofilacium quod erat contra separatum aedificium et contra aedem vergentem ad aquilonem
EZEK|42|2|in facie longitudinis centum cubitos ostii aquilonis et latitudinis quinquaginta cubitos
EZEK|42|3|contra viginti cubitos atrii interioris et contra pavimentum stratum lapide atrii exterioris ubi erat porticus iuncta porticui triplici
EZEK|42|4|et ante gazofilacia deambulatio decem cubitorum latitudinis ad interiora respiciens viae cubiti unius et ostia earum ad aquilonem
EZEK|42|5|ubi erant gazofilacia in superioribus humiliora quia subportabant porticus quae ex illis eminebant de inferioribus et de mediis aedificii
EZEK|42|6|tristega enim erant et non habebant columnas sicut erant columnae atriorum propterea eminebant de inferioribus et de mediis a terra
EZEK|42|7|et peribolus exterior secundum gazofilacia quae erant in via atrii exterioris ante gazofilacia longitudo eius quinquaginta cubitorum
EZEK|42|8|quia longitudo erat gazofilaciorum atrii exterioris quinquaginta cubitorum et longitudo ante faciem templi centum cubitorum
EZEK|42|9|et erat subter gazofilacia haec introitus ab oriente ingredientium in ea de atrio exteriori
EZEK|42|10|in latitudine periboli atrii quod erat contra viam orientalem in facie aedificii separati et erant ante aedificium gazofilacia
EZEK|42|11|et via ante faciem eorum iuxta similitudinem gazofilaciorum quae erant in via aquilonis secundum longitudinem eorum sic et latitudo eorum et omnis introitus eorum et similitudines et ostia eorum
EZEK|42|12|secundum ostia gazofilaciorum quae erant in via respiciente ad notum ostium in capite viae quae via erat ante vestibulum separatum per viam orientalem ingredientibus
EZEK|42|13|et dixit ad me gazofilacia aquilonis et gazofilacia austri quae sunt ante aedificium separatum haec sunt gazofilacia sancta in quibus vescuntur sacerdotes qui adpropinquant ad Dominum in sancta sanctorum ibi ponent sancta sanctorum et oblationem pro peccato et pro delicto locus enim sanctus est
EZEK|42|14|cum autem ingressi fuerint sacerdotes non egredientur de sanctis in atrium exterius et ibi reponent vestimenta sua in quibus ministrant quia sancta sunt vestienturque vestimentis aliis et sic procedent ad populum
EZEK|42|15|cumque conplesset mensuras domus interioris eduxit me per viam portae quae respiciebat ad viam orientalem et mensus est eam undique per circuitum
EZEK|42|16|mensus autem est contra ventum orientalem calamo mensurae quingentos calamos in calamo mensurae per circuitum
EZEK|42|17|et mensus est contra ventum aquilonem quingentos calamos in calamo mensurae per gyrum
EZEK|42|18|et ad ventum australem mensus est quingentos calamos in calamo mensurae per circuitum
EZEK|42|19|et ad ventum occidentalem mensus est quingentos calamos in calamo mensurae
EZEK|42|20|per quattuor ventos mensus est illud murum eius undique per circuitum longitudine quingentorum cubitorum et latitudine quingentorum cubitorum dividentem inter sanctuarium et vulgi locum
EZEK|43|1|et duxit me ad portam quae respiciebat ad viam orientalem
EZEK|43|2|et ecce gloria Dei Israhel ingrediebatur per viam orientalem et vox erat ei quasi vox aquarum multarum et terra splendebat a maiestate eius
EZEK|43|3|et vidi visionem secundum speciem quam videram quando venit ut disperderet civitatem et species secundum aspectum quem videram iuxta fluvium Chobar et cecidi super faciem meam
EZEK|43|4|et maiestas Domini ingressa est templum per viam portae quae respiciebat ad orientem
EZEK|43|5|et levavit me spiritus et introduxit me in atrium interius et ecce repleta erat gloria Domini domus
EZEK|43|6|et audivi loquentem ad me de domo et vir qui stabat iuxta me
EZEK|43|7|dixit ad me fili hominis locus solii mei et locus vestigiorum pedum meorum ubi habito in medio filiorum Israhel in aeternum et non polluent ultra domus Israhel nomen sanctum meum ipsi et reges eorum in fornicationibus suis et in ruinis regum suorum et in excelsis
EZEK|43|8|qui fabricati sunt limen suum iuxta limen meum et postes suos iuxta postes meos et murus erat inter me et eos et polluerunt nomen sanctum meum in abominationibus quas fecerunt propter quod consumpsi eos in ira mea
EZEK|43|9|nunc ergo repellant procul fornicationem suam et ruinas regum suorum a me et habitabo in medio eorum semper
EZEK|43|10|tu autem fili hominis ostende domui Israhel templum et confundantur ab iniquitatibus suis et metiantur fabricam
EZEK|43|11|et erubescant ex omnibus quae fecerunt figuram domus et fabricae eius exitus et introitus et omnem descriptionem eius et universa praecepta eius cunctumque ordinem eius et omnes leges eius ostende eis et scribes in oculis eorum et custodiant omnes descriptiones eius et praecepta illius et faciant ea
EZEK|43|12|ista est lex domus in summitate montis omnes fines eius in circuitu sanctum sanctorum est haec ergo est lex domus
EZEK|43|13|istae autem mensurae altaris in cubito verissimo qui habebat cubitum et palmum in sinu eius erat cubitus et cubitus in latitudine et definitio usque ad labium eius in circuitu palmus unus haec quoque erat fossa altaris
EZEK|43|14|et de sinu terrae usque ad crepidinem novissimam duo cubiti et latitudo cubiti unius et a crepidine maiori usque ad crepidinem minorem quattuor cubiti et latitudo unius cubiti
EZEK|43|15|ipse autem arihel quattuor cubitorum et ab arihel usque sursum cornua quattuor
EZEK|43|16|et arihel duodecim cubitorum in longitudine per duodecim cubitos latitudinis quadrangulatum aequis lateribus
EZEK|43|17|et crepido quattuordecim cubitorum longitudinis per quattuordecim latitudinis in quattuor angulis eius et corona in circuitu eius dimidii cubitus et sinus eius unius cubiti per circuitum gradus autem eius versi ad orientem
EZEK|43|18|et dixit ad me fili hominis haec dicit Dominus Deus hii sunt ritus altaris in quacumque die fuerit fabricatum ut offeratur super illud holocaustum et effundatur sanguis
EZEK|43|19|et dabis sacerdotibus Levitis qui sunt de semine Sadoc qui accedunt ad me ait Dominus Deus ut offerant mihi vitulum de armento pro peccato
EZEK|43|20|et adsumens de sanguine eius pones super quattuor cornua eius et super quattuor angulos crepidinis et super coronam in circuitu et mundabis illud et expiabis
EZEK|43|21|et tolles vitulum qui oblatus fuerit pro peccato et conbures illum in separato loco domus extra sanctuarium
EZEK|43|22|et in die secunda offeres hircum caprarum inmaculatum pro peccato et expiabunt altare sicut expiaverunt in vitulo
EZEK|43|23|cumque conpleveris expians illud offeres vitulum de armento inmaculatum et arietem de grege inmaculatum
EZEK|43|24|et offeres eos in conspectu Domini et mittent sacerdotes super eos sal et offerent eos holocaustum Domino
EZEK|43|25|septem diebus facies hircum pro peccato cotidie et vitulum de armento et arietem de pecoribus inmaculatos offerent
EZEK|43|26|septem diebus expiabunt altare et mundabunt illud et implebunt manum eius
EZEK|43|27|expletis autem diebus in die octava et ultra facient sacerdotes super altare holocausta vestra et quae pro pace offerunt et placatus ero vobis ait Dominus Deus
EZEK|44|1|et convertit me ad viam portae sanctuarii exterioris quae respiciebat ad orientem et erat clausa
EZEK|44|2|et dixit Dominus ad me porta haec clausa erit non aperietur et vir non transiet per eam quoniam Dominus Deus Israhel ingressus est per eam eritque clausa
EZEK|44|3|principi princeps ipse sedebit in ea ut comedat panem coram Domino per viam vestibuli portae ingredietur et per viam eius egredietur
EZEK|44|4|et adduxit me per viam portae aquilonis in conspectu domus et vidi et ecce implevit gloria Domini domum Domini et cecidi in faciem meam
EZEK|44|5|et dixit ad me Dominus fili hominis pone cor tuum et vide oculis tuis et auribus tuis audi omnia quae ego loquor ad te de universis caerimoniis domus Domini et de cunctis legibus eius et pones cor tuum in viis templi per omnes exitus sanctuarii
EZEK|44|6|et dices ad exasperantem me domum Israhel haec dicit Dominus Deus sufficiant vobis omnia scelera vestra domus Israhel
EZEK|44|7|eo quod inducitis filios alienos incircumcisos corde et incircumcisos carne ut sint in sanctuario meo et polluant domum meam et offertis panes meos adipem et sanguinem et dissolvitis pactum meum in omnibus sceleribus vestris
EZEK|44|8|et non servastis praecepta sanctuarii mei et posuistis custodes observationum mearum in sanctuario meo vobismet ipsis
EZEK|44|9|haec dicit Dominus Deus omnis alienigena incircumcisus corde et incircumcisus carne non ingredietur sanctuarium meum omnis filius alienus qui est in medio filiorum Israhel
EZEK|44|10|sed et Levitae qui longe recesserunt a me in errore filiorum Israhel et erraverunt a me post idola sua et portaverunt iniquitatem suam
EZEK|44|11|erunt in sanctuario meo aeditui et ianitores portarum domus et ministri domus ipsi mactabunt holocaustosin et victimas populi et ipsi stabunt in conspectu eorum ut ministrent eis
EZEK|44|12|pro eo quod ministraverunt illis in conspectu idolorum suorum et facti sunt domui Israhel in offendiculum iniquitatis idcirco levavi manum meam super eos dicit Dominus Deus et portaverunt iniquitatem suam
EZEK|44|13|et non adpropinquabunt ad me ut sacerdotio fungantur mihi neque accedent ad omne sanctuarium meum iuxta sancta sanctorum sed portabunt confusionem suam et scelera sua quae fecerunt
EZEK|44|14|et dabo eos ianitores domus in omni ministerio eius et universis quae fiunt in ea
EZEK|44|15|sacerdotes autem Levitae filii Sadoc qui custodierunt caerimonias sanctuarii mei cum errarent filii Israhel a me ipsi accedent ad me ut ministrent mihi et stabunt in conspectu meo ut offerant mihi adipem et sanguinem ait Dominus Deus
EZEK|44|16|ipsi ingredientur sanctuarium meum et ipsi accedent ad mensam meam ut ministrent mihi et custodiant caerimonias meas
EZEK|44|17|cumque ingredientur portas atrii interioris vestibus lineis induentur nec ascendet super eos quicquam laneum quando ministrant in portis atrii interioris et intrinsecus
EZEK|44|18|vittae lineae erunt in capitibus eorum et feminalia linea erunt in lumbis eorum et non accingentur in sudore
EZEK|44|19|cumque egredientur atrium exterius ad populum exuent se vestimenta sua in quibus ministraverunt et reponent ea in gazofilacio sanctuarii et vestient se vestimentis aliis et non sanctificabunt populum in vestibus suis
EZEK|44|20|caput autem suum non radent neque comam nutrient sed tondentes adtondent capita sua
EZEK|44|21|et vinum non bibet omnis sacerdos quando ingressurus est atrium interius
EZEK|44|22|et viduam et repudiatam non accipient uxores sed virgines de semine domus Israhel sed et viduam quae fuerit vidua a sacerdote accipient
EZEK|44|23|et populum meum docebunt quid sit inter sanctum et pollutum et inter mundum et inmundum ostendent eis
EZEK|44|24|et cum fuerit controversia stabunt in iudiciis meis et iudicabunt leges meas et praecepta mea in omnibus sollemnitatibus meis custodient et sabbata mea sanctificabunt
EZEK|44|25|et ad mortuum hominem non ingredientur ne polluantur nisi ad patrem et matrem et filium et filiam et fratrem et sororem quae alterum virum non habuit in quibus contaminabuntur
EZEK|44|26|et postquam fuerit emundatus septem dies numerabuntur ei
EZEK|44|27|et in die introitus sui in sanctuarium ad atrium interius ut ministret mihi in sanctuario offeret pro peccato suo ait Dominus Deus
EZEK|44|28|erit autem eis hereditas ego hereditas eorum et possessionem non dabitis eis in Israhel ego enim possessio eorum
EZEK|44|29|victimam et pro peccato et pro delicto ipsi comedent et omne votum in Israhel ipsorum erit
EZEK|44|30|et primitiva omnium primogenitorum et omnia libamenta ex omnibus quae offeruntur sacerdotum erunt et primitiva ciborum vestrorum dabitis sacerdoti ut reponat benedictionem domui suae
EZEK|44|31|omne morticinum et captum a bestia de avibus et de pecoribus non comedent sacerdotes
EZEK|45|1|cumque coeperitis terram dividere sortito separate primitias Domino sanctificatum de terra longitudine viginti quinque milia et latitudine decem milia sanctificatum erit in omni termino eius per circuitum
EZEK|45|2|et erit ex omni parte sanctificatum quingentos per quingentos quadrifariam per circuitum et quinquaginta cubitis in suburbana eius per gyrum
EZEK|45|3|et a mensura ista mensurabis longitudinem viginti quinque milium et latitudinem decem milium et in ipso erit templum sanctumque sanctorum
EZEK|45|4|sanctificatum de terra erit sacerdotibus ministris sanctuarii qui accedunt ad ministerium Domini et erit eis locus in domos et in sanctuarium sanctitatis
EZEK|45|5|viginti quinque autem milia longitudinis et decem milia latitudinis erunt Levitis qui ministrant domui ipsi possidebunt viginti gazofilacia
EZEK|45|6|et possessionem civitatis dabitis quinque milia latitudinis et longitudinis viginti quinque milia secundum separationem sanctuarii omni domui Israhel
EZEK|45|7|principi quoque hinc et inde in separationem sanctuarii et in possessionem civitatis contra faciem separationis sanctuarii et contra faciem possessionis urbis a latere maris usque ad mare et a latere orientis usque ad orientem longitudinem autem iuxta unamquamque partium a termino occidentali usque ad terminum orientalem
EZEK|45|8|de terra erit ei possessio in Israhel et non depopulabuntur ultra principes populum meum sed terram dabunt domui Israhel secundum tribus eorum
EZEK|45|9|haec dicit Dominus Deus sufficiat vobis principes Israhel iniquitatem et rapinas intermittite et iudicium et iustitiam facite separate confinia vestra a populo meo ait Dominus Deus
EZEK|45|10|statera iusta et oephi iustum et batus iustus erit vobis
EZEK|45|11|oephi et batus aequalia et unius mensurae erunt ut capiat decimam partem chori batus et decimam partem chori oephi iuxta mensuram chori erit aequa libratio eorum
EZEK|45|12|siclus autem viginti obolos habeat porro viginti sicli et viginti quinque sicli et quindecim sicli minam facient
EZEK|45|13|et haec sunt primitiae quas tolletis sextam partem oephi de choro frumenti et sextam partem oephi de choro hordei
EZEK|45|14|mensura quoque olei batus olei decima pars chori est et decem bati chorum faciunt quia decem bati implent chorum
EZEK|45|15|et arietem unum de grege ducentorum de his quae nutriunt Israhel in sacrificium et in holocaustum et in pacifica ad expiandum pro eis ait Dominus Deus
EZEK|45|16|omnis populus terrae tenebitur primitiis his principi in Israhel
EZEK|45|17|et super principem erunt holocausta et sacrificium et libamina in sollemnitatibus et in kalendis et in sabbatis in universis sollemnitatibus domus Israhel ipse faciat pro peccato sacrificium et holocaustum et pacifica ad expiandum pro domo Israhel
EZEK|45|18|haec dicit Dominus Deus in primo mense una mensis sumes vitulum de armento inmaculatum et expiabis sanctuarium
EZEK|45|19|et tollet sacerdos de sanguine quod erit pro peccato et ponet in postibus domus et in quattuor angulis crepidinis altaris et in postibus portae atrii interioris
EZEK|45|20|et sic facies in septima mensis pro unoquoque qui ignoravit et errore deceptus est et expiabitis pro domo
EZEK|45|21|in primo mense quartadecima die mensis erit vobis paschae sollemnitas septem diebus azyma comedentur
EZEK|45|22|et faciet princeps in die illa pro se et pro universo populo terrae vitulum pro peccato
EZEK|45|23|et in septem dierum sollemnitate faciet holocaustum Domino septem vitulos et septem arietes inmaculatos cotidie septem diebus et pro peccato hircum caprarum cotidie
EZEK|45|24|et sacrificium oephi per vitulum et oephi per arietem faciet et olei hin per singula oephi
EZEK|45|25|septimo mense quintadecima die mensis in sollemnitate faciet sicut supra dicta sunt per septem dies tam pro peccato quam pro holocausto et in sacrificio et in oleo
EZEK|46|1|haec dicit Dominus Deus porta atrii interioris quae respicit ad orientem erit clausa sex diebus in quibus opus fit die autem sabbati aperietur sed et in die kalendarum aperietur
EZEK|46|2|et intrabit princeps per viam vestibuli portae de foris et stabit in limine portae et facient sacerdotes holocaustum eius et pacifica eius et adorabit super limen portae et egredietur porta autem non claudetur usque ad vesperam
EZEK|46|3|et adorabit populus terrae ad ostium portae illius in sabbatis et in kalendis coram Domino
EZEK|46|4|holocaustum autem hoc offeret princeps Domino in die sabbati sex agnos inmaculatos et arietem inmaculatum
EZEK|46|5|et sacrificium oephi per arietem agnis autem sacrificium quod dederit manus eius et olei hin per singula oephi
EZEK|46|6|in die autem kalendarum vitulum de armento inmaculatum et sex agni et arietes inmaculati erunt
EZEK|46|7|et oephi per vitulum oephi quoque per arietem faciet sacrificium agnis autem sicut invenerit manus eius et olei hin per singula oephi
EZEK|46|8|cumque ingressurus est princeps per viam vestibuli portae ingrediatur et per eandem viam exeat
EZEK|46|9|et cum intrabit populus terrae in conspectu Domini in sollemnitatibus qui ingreditur per portam aquilonis ut adoret egrediatur per viam portae meridianae porro qui ingreditur per viam portae meridianae egrediatur per viam portae aquilonis non revertetur per viam portae per quam ingressus est sed e regione illius egredietur
EZEK|46|10|princeps autem in medio eorum cum ingredientibus ingredietur et cum egredientibus egredietur
EZEK|46|11|et in nundinis et in sollemnitatibus erit sacrificium oephi per vitulum et oephi per arietem agnis autem erit sacrificium sicut invenerit manus eius et olei hin per singula oephi
EZEK|46|12|cum autem fecerit princeps spontaneum holocaustum aut pacifica voluntaria Domino aperietur ei porta quae respicit ad orientem et faciet holocaustum suum et pacifica sua sicut fieri solet in die sabbati et egredietur claudeturque porta postquam exierit
EZEK|46|13|et agnum eiusdem anni inmaculatum faciet holocaustum cotidie Domino semper mane faciet illud
EZEK|46|14|et sacrificium faciet super eo cata mane mane sextam partem oephi et de oleo tertiam partem hin ut misceatur similae sacrificium Domino legitimum iuge atque perpetuum
EZEK|46|15|faciet agnum et sacrificium et oleum cata mane mane holocaustum sempiternum
EZEK|46|16|haec dicit Dominus Deus si dederit princeps donum alicui de filiis suis hereditas eius filiorum suorum erit possidebunt ea hereditarie
EZEK|46|17|si autem dederit legatum de hereditate sua uni servorum suorum erit illius usque ad annum remissionis et revertetur ad principem hereditas autem eius filiis eius erit
EZEK|46|18|et non accipiet princeps de hereditate populi per violentiam et de possessione eorum sed de possessione sua hereditatem dabit filiis suis ut non dispergatur populus meus unusquisque a possessione sua
EZEK|46|19|et introduxit me per ingressum qui erat ex latere portae in gazofilacia sanctuarii ad sacerdotes quae respiciebant ad aquilonem et erat ibi locus vergens ad occidentem
EZEK|46|20|et dixit ad me iste est locus ubi coquent sacerdotes pro delicto et pro peccato ubi coquent sacrificium ut non efferant in atrio exteriori et sanctificetur populus
EZEK|46|21|et eduxit me in atrium exterius et circumduxit me per quattuor angulos atrii et ecce atriolum erat in angulo atrii atriola singula per angulos atrii
EZEK|46|22|in quattuor angulos atrii atriola disposita quadraginta cubitorum per longum et triginta per latum mensurae unius quattuor erant
EZEK|46|23|et paries per circuitum ambiens quattuor atriola et culinae fabricatae erant subter porticus per gyrum
EZEK|46|24|et dixit ad me haec est domus culinarum in qua coquent ministri domus Domini victimas populi
EZEK|47|1|et convertit me ad portam domus et ecce aquae egrediebantur subter limen domus ad orientem facies enim domus respiciebat ad orientem aquae autem descendebant in latus templi dextrum ad meridiem altaris
EZEK|47|2|et eduxit me per viam portae aquilonis et convertit me ad viam foras portam exteriorem viam quae respiciebat ad orientem et ecce aquae redundantes a latere dextro
EZEK|47|3|cum egrederetur vir ad orientem qui habebat funiculum in manu sua et mensus est mille cubitos et transduxit me per aquam usque ad talos
EZEK|47|4|rursumque mensus est mille et transduxit me per aquam usque ad genua
EZEK|47|5|et mensus est mille et transduxit me per aquam usque ad renes et mensus est mille torrentem quem non potui pertransire quoniam intumuerant aquae profundae torrentis qui non potest transvadari
EZEK|47|6|et dixit ad me certe vidisti fili hominis et duxit me et convertit ad ripam torrentis
EZEK|47|7|cumque me convertissem ecce in ripa torrentis ligna multa nimis ex utraque parte
EZEK|47|8|et ait ad me aquae istae quae egrediuntur ad tumulos sabuli orientalis et descendunt ad plana deserti intrabunt mare et exibunt et sanabuntur aquae
EZEK|47|9|et omnis anima vivens quae serpit quocumque venerit torrens vivet et erunt pisces multi satis postquam venerint illuc aquae istae et sanabuntur et vivent omnia ad quae venerit torrens
EZEK|47|10|vivent et stabunt super illa piscatores ab Engaddi usque ad Engallim siccatio sagenarum erunt plurimae species erunt piscium eius sicut pisces maris magni multitudinis nimiae
EZEK|47|11|in litoribus autem eius et in palustribus non sanabuntur quia in salinas dabuntur
EZEK|47|12|et super torrentem orietur in ripis eius ex utraque parte omne lignum pomiferum non defluet folium ex eo et non deficiet fructus eius per singulos menses adferet primitiva quia aquae eius de sanctuario egredientur et erunt fructus eius in cibum et folia eius ad medicinam
EZEK|47|13|haec dicit Dominus Deus hic est terminus in quo possidebitis terram in duodecim tribubus Israhel quia Ioseph duplicem funiculum habet
EZEK|47|14|possidebitis autem eam singuli aeque ut frater suus quam levavi manum meam ut darem patribus vestris et cadet terra haec vobis in possessionem
EZEK|47|15|hic est autem terminus terrae ad plagam septentrionalem a mari magno via Bethalon venientibus Sadada
EZEK|47|16|Emath Berotha Sabarim quae est inter terminum Damasci et confinium Emath domus Atticon quae est iuxta terminos Auran
EZEK|47|17|et erit terminus a mari usque ad atrium Aenon terminus Damasci et ab aquilone ad aquilonem et terminus Emath plaga autem septentrionalis
EZEK|47|18|porro plaga orientalis de medio Auran et de medio Damasci et de medio Galaad et de medio terrae Israhel Iordanis disterminans ad mare orientale metiemini etiam plagam orientalem
EZEK|47|19|plaga autem australis meridiana a Thamar usque ad aquas Contradictionis Cades et torrens usque ad mare magnum et plaga ad meridiem australis
EZEK|47|20|et plaga maris mare magnum a confinio per directum donec venias Emath haec est plaga maris
EZEK|47|21|et dividetis terram istam vobis per tribus Israhel
EZEK|47|22|et mittetis eam in hereditatem vobis et advenis qui accesserint ad vos qui genuerint filios in medio vestrum et erunt vobis sicut indigenae inter filios Israhel vobiscum divident possessionem in medio tribuum Israhel
EZEK|47|23|in tribu autem quacumque fuerit advena ibi dabitis possessionem illi ait Dominus Deus
EZEK|48|1|et haec nomina tribuum a finibus aquilonis iuxta viam Aethlon pergentibus Emath atrium Aenon terminus Damasci ad aquilonem iuxta Emath et erit ei plaga orientalis mare Dan una
EZEK|48|2|et ad terminum Dan a plaga orientali usque ad plagam maris Aser una
EZEK|48|3|et super terminum Aser a plaga orientali usque ad plagam maris Nepthalim una
EZEK|48|4|et super terminum Nepthalim a plaga orientali usque ad plagam maris Manasse una
EZEK|48|5|et super terminum Manasse a plaga orientali usque ad plagam maris Ephraim una
EZEK|48|6|et super terminum Ephraim a plaga orientali usque ad plagam maris Ruben una
EZEK|48|7|et super terminum Ruben a plaga orientali usque ad plagam maris Iuda una
EZEK|48|8|et super terminum Iuda a plaga orientali usque ad plagam maris erunt primitiae quas separabitis viginti quinque milibus latitudinis et longitudinis sicuti singulae partes a plaga orientali usque ad plagam maris et erit sanctuarium in medio eius
EZEK|48|9|primitiae quas separastis Domino longitudo viginti quinque milibus et latitudo decem milibus
EZEK|48|10|hae autem erunt primitiae sanctuarii sacerdotum ad aquilonem viginti quinque milia et ad mare latitudinis decem milia sed et ad orientem latitudinis decem milia et ad meridiem longitudinis viginti quinque milia et erit sanctuarium Domini in medio eius
EZEK|48|11|sacerdotibus sanctuarium erit de filiis Sadoc qui custodierunt caerimonias meas et non erraverunt cum errarent filii Israhel sicut erraverunt et Levitae
EZEK|48|12|et erunt eis primitiae de primitiis terrae sanctum sanctorum iuxta terminum Levitarum
EZEK|48|13|sed et Levitis similiter iuxta fines sacerdotum viginti quinque milia longitudinis et latitudinis decem milia omnis longitudo viginti et quinque milium et latitudo decem milium
EZEK|48|14|et non venundabunt ex eo neque mutabunt nec transferentur primitiae terrae quia sanctificatae sunt Domino
EZEK|48|15|quinque milia autem quae supersunt in latitudine per viginti quinque milia profana erunt urbis in habitaculum et in suburbana et erit civitas in medio eius
EZEK|48|16|et heae mensurae eius ad plagam septentrionalem quingenti et quattuor milia et ad plagam meridianam quingenti et quattuor milia et ad plagam orientalem quingenti et quattuor milia et ad plagam occidentalem quingenti et quattuor milia
EZEK|48|17|erunt autem suburbana civitatis ad aquilonem ducenti quinquaginta et in meridie ducenti quinquaginta et ad orientem ducenti quinquaginta et ad mare ducenti quinquaginta
EZEK|48|18|quod autem reliquum fuerit in longitudine secundum primitias sanctuarii decem milia in orientem et decem milia ad occidentem erunt sicut primitiae sanctuarii et erunt fruges eius in panes his qui serviunt civitati
EZEK|48|19|servientes autem civitati operabuntur ex omnibus tribubus Israhel
EZEK|48|20|omnes primitiae viginti quinque milium per viginti quinque milia in quadrum separabuntur in primitias sanctuarii et possessionem civitatis
EZEK|48|21|quod autem reliquum fuerit principis erit ex omni parte primitiarum sanctuarii et possessionis civitatis e regione viginti quinque milium primitiarum usque ad terminum orientalem sed et ad mare e regione viginti quinque milium usque ad terminum maris similiter in partibus principis erit et erunt primitiae sanctuarii et sanctuarium templi in medio eius
EZEK|48|22|de possessione autem Levitarum et de possessione civitatis in medio partium principis erit inter terminum Iuda et inter terminum Beniamin et ad principem pertinebit
EZEK|48|23|et reliquis tribubus a plaga orientali usque ad plagam occidentalem Beniamin una
EZEK|48|24|et contra terminum Beniamin a plaga orientali usque ad plagam occidentalem Symeon una
EZEK|48|25|et super terminum Symeonis a plaga orientali usque ad plagam occidentis Isachar una
EZEK|48|26|et super terminum Isachar a plaga orientali usque ad plagam occidentalem Zabulon una
EZEK|48|27|et super terminum Zabulon a plaga orientali usque ad plagam maris Gad una
EZEK|48|28|et super terminum Gad ad plagam austri in meridiem et erit finis de Thamar usque ad aquas Contradictionis Cades hereditas contra mare magnum
EZEK|48|29|haec est terra quam mittetis in sortem tribubus Israhel et hae partitiones earum ait Dominus Deus
EZEK|48|30|et hii egressus civitatis a plaga septentrionali quingentos et quattuor milia mensurabis
EZEK|48|31|et portae civitatis in nominibus tribuum Israhel portae tres a septentrione porta Ruben una porta Iudae una porta Levi una
EZEK|48|32|et ad plagam orientalem quingentos et quattuor milia et portae tres porta Ioseph una porta Beniamin una porta Dan una
EZEK|48|33|et ad plagam meridianam quingentos et quattuor milia metieris portam Symeonis unam portam Isachar unam portam Zabulon unam
EZEK|48|34|et ad plagam occidentalem quingenti et quattuor milia portae eorum tres porta Gad una porta Aser una porta Nepthalim una
EZEK|48|35|per circuitum decem et octo milia et nomen civitatis ex illa die Dominus ibidem
