EPH|1|1|Paulus apostolus Christi Iesu per voluntatem Dei sanctis omnibus qui sunt Ephesi et fidelibus in Christo Iesu
EPH|1|2|gratia vobis et pax a Deo Patre nostro et Domino Iesu Christo
EPH|1|3|benedictus Deus et Pater Domini nostri Iesu Christi qui benedixit nos in omni benedictione spiritali in caelestibus in Christo
EPH|1|4|sicut elegit nos in ipso ante mundi constitutionem ut essemus sancti et inmaculati in conspectu eius in caritate
EPH|1|5|qui praedestinavit nos in adoptionem filiorum per Iesum Christum in ipsum secundum propositum voluntatis suae
EPH|1|6|in laudem gloriae gratiae suae in qua gratificavit nos in dilecto
EPH|1|7|in quo habemus redemptionem per sanguinem eius remissionem peccatorum secundum divitias gratiae eius
EPH|1|8|quae superabundavit in nobis in omni sapientia et prudentia
EPH|1|9|ut notum faceret nobis sacramentum voluntatis suae secundum bonum placitum eius quod proposuit in eo
EPH|1|10|in dispensationem plenitudinis temporum instaurare omnia in Christo quae in caelis et quae in terra sunt in ipso
EPH|1|11|in quo etiam sorte vocati sumus praedestinati secundum propositum eius qui omnia operatur secundum consilium voluntatis suae
EPH|1|12|ut simus in laudem gloriae eius qui ante speravimus in Christo
EPH|1|13|in quo et vos cum audissetis verbum veritatis evangelium salutis vestrae in quo et credentes signati estis Spiritu promissionis Sancto
EPH|1|14|qui est pignus hereditatis nostrae in redemptionem adquisitionis in laudem gloriae ipsius
EPH|1|15|propterea et ego audiens fidem vestram quae est in Domino Iesu et dilectionem in omnes sanctos
EPH|1|16|non cesso gratias agens pro vobis memoriam vestri faciens in orationibus meis
EPH|1|17|ut Deus Domini nostri Iesu Christi Pater gloriae det vobis spiritum sapientiae et revelationis in agnitione eius
EPH|1|18|inluminatos oculos cordis vestri ut sciatis quae sit spes vocationis eius quae divitiae gloriae hereditatis eius in sanctis
EPH|1|19|et quae sit supereminens magnitudo virtutis eius in nos qui credidimus secundum operationem potentiae virtutis eius
EPH|1|20|quam operatus est in Christo suscitans illum a mortuis et constituens ad dexteram suam in caelestibus
EPH|1|21|supra omnem principatum et potestatem et virtutem et dominationem et omne nomen quod nominatur non solum in hoc saeculo sed et in futuro
EPH|1|22|et omnia subiecit sub pedibus eius et ipsum dedit caput supra omnia ecclesiae
EPH|1|23|quae est corpus ipsius plenitudo eius qui omnia in omnibus adimpletur
EPH|2|1|et vos cum essetis mortui delictis et peccatis vestris
EPH|2|2|in quibus aliquando ambulastis secundum saeculum mundi huius secundum principem potestatis aeris huius spiritus qui nunc operatur in filios diffidentiae
EPH|2|3|in quibus et nos omnes aliquando conversati sumus in desideriis carnis nostrae facientes voluntates carnis et cogitationum et eramus natura filii irae sicut et ceteri
EPH|2|4|Deus autem qui dives est in misericordia propter nimiam caritatem suam qua dilexit nos
EPH|2|5|et cum essemus mortui peccatis convivificavit nos Christo gratia estis salvati
EPH|2|6|et conresuscitavit et consedere fecit in caelestibus in Christo Iesu
EPH|2|7|ut ostenderet in saeculis supervenientibus abundantes divitias gratiae suae in bonitate super nos in Christo Iesu
EPH|2|8|gratia enim estis salvati per fidem et hoc non ex vobis Dei enim donum est
EPH|2|9|non ex operibus ut ne quis glorietur
EPH|2|10|ipsius enim sumus factura creati in Christo Iesu in operibus bonis quae praeparavit Deus ut in illis ambulemus
EPH|2|11|propter quod memores estote quod aliquando vos gentes in carne qui dicimini praeputium ab ea quae dicitur circumcisio in carne manufacta
EPH|2|12|quia eratis illo in tempore sine Christo alienati a conversatione Israhel et hospites testamentorum promissionis spem non habentes et sine Deo in mundo
EPH|2|13|nunc autem in Christo Iesu vos qui aliquando eratis longe facti estis prope in sanguine Christi
EPH|2|14|ipse est enim pax nostra qui fecit utraque unum et medium parietem maceriae solvens inimicitiam in carne sua
EPH|2|15|legem mandatorum decretis evacuans ut duos condat in semet ipsum in unum novum hominem faciens pacem
EPH|2|16|et reconciliet ambos in uno corpore Deo per crucem interficiens inimicitiam in semet ipso
EPH|2|17|et veniens evangelizavit pacem vobis qui longe fuistis et pacem his qui prope
EPH|2|18|quoniam per ipsum habemus accessum ambo in uno Spiritu ad Patrem
EPH|2|19|ergo iam non estis hospites et advenae sed estis cives sanctorum et domestici Dei
EPH|2|20|superaedificati super fundamentum apostolorum et prophetarum ipso summo angulari lapide Christo Iesu
EPH|2|21|in quo omnis aedificatio constructa crescit in templum sanctum in Domino
EPH|2|22|in quo et vos coaedificamini in habitaculum Dei in Spiritu
EPH|3|1|huius rei gratia ego Paulus vinctus Christi Iesu pro vobis gentibus
EPH|3|2|si tamen audistis dispensationem gratiae Dei quae data est mihi in vobis
EPH|3|3|quoniam secundum revelationem notum mihi factum est sacramentum sicut supra scripsi in brevi
EPH|3|4|prout potestis legentes intellegere prudentiam meam in mysterio Christi
EPH|3|5|quod aliis generationibus non est agnitum filiis hominum sicuti nunc revelatum est sanctis apostolis eius et prophetis in Spiritu
EPH|3|6|esse gentes coheredes et concorporales et conparticipes promissionis in Christo Iesu per evangelium
EPH|3|7|cuius factus sum minister secundum donum gratiae Dei quae data est mihi secundum operationem virtutis eius
EPH|3|8|mihi omnium sanctorum minimo data est gratia haec in gentibus evangelizare ininvestigabiles divitias Christi
EPH|3|9|et inluminare omnes quae sit dispensatio sacramenti absconditi a saeculis in Deo qui omnia creavit
EPH|3|10|ut innotescat principibus et potestatibus in caelestibus per ecclesiam multiformis sapientia Dei
EPH|3|11|secundum praefinitionem saeculorum quam fecit in Christo Iesu Domino nostro
EPH|3|12|in quo habemus fiduciam et accessum in confidentia per fidem eius
EPH|3|13|propter quod peto ne deficiatis in tribulationibus meis pro vobis quae est gloria vestra
EPH|3|14|huius rei gratia flecto genua mea ad Patrem Domini nostri Iesu Christi
EPH|3|15|ex quo omnis paternitas in caelis et in terra nominatur
EPH|3|16|ut det vobis secundum divitias gloriae suae virtute corroborari per Spiritum eius in interiore homine
EPH|3|17|habitare Christum per fidem in cordibus vestris in caritate radicati et fundati
EPH|3|18|ut possitis conprehendere cum omnibus sanctis quae sit latitudo et longitudo et sublimitas et profundum
EPH|3|19|scire etiam supereminentem scientiae caritatem Christi ut impleamini in omnem plenitudinem Dei
EPH|3|20|ei autem qui potens est omnia facere superabundanter quam petimus aut intellegimus secundum virtutem quae operatur in nobis
EPH|3|21|ipsi gloria in ecclesia et in Christo Iesu in omnes generationes saeculi saeculorum amen
EPH|4|1|obsecro itaque vos ego vinctus in Domino ut digne ambuletis vocatione qua vocati estis
EPH|4|2|cum omni humilitate et mansuetudine cum patientia subportantes invicem in caritate
EPH|4|3|solliciti servare unitatem spiritus in vinculo pacis
EPH|4|4|unum corpus et unus spiritus sicut vocati estis in una spe vocationis vestrae
EPH|4|5|unus Dominus una fides unum baptisma
EPH|4|6|unus Deus et Pater omnium qui super omnes et per omnia et in omnibus nobis
EPH|4|7|unicuique autem nostrum data est gratia secundum mensuram donationis Christi
EPH|4|8|propter quod dicit ascendens in altum captivam duxit captivitatem dedit dona hominibus
EPH|4|9|quod autem ascendit quid est nisi quia et descendit primum in inferiores partes terrae
EPH|4|10|qui descendit ipse est et qui ascendit super omnes caelos ut impleret omnia
EPH|4|11|et ipse dedit quosdam quidem apostolos quosdam autem prophetas alios vero evangelistas alios autem pastores et doctores
EPH|4|12|ad consummationem sanctorum in opus ministerii in aedificationem corporis Christi
EPH|4|13|donec occurramus omnes in unitatem fidei et agnitionis Filii Dei in virum perfectum in mensuram aetatis plenitudinis Christi
EPH|4|14|ut iam non simus parvuli fluctuantes et circumferamur omni vento doctrinae in nequitia hominum in astutia ad circumventionem erroris
EPH|4|15|veritatem autem facientes in caritate crescamus in illo per omnia qui est caput Christus
EPH|4|16|ex quo totum corpus conpactum et conexum per omnem iuncturam subministrationis secundum operationem in mensuram uniuscuiusque membri augmentum corporis facit in aedificationem sui in caritate
EPH|4|17|hoc igitur dico et testificor in Domino ut iam non ambuletis sicut gentes ambulant in vanitate sensus sui
EPH|4|18|tenebris obscuratum habentes intellectum alienati a vita Dei per ignorantiam quae est in illis propter caecitatem cordis ipsorum
EPH|4|19|qui desperantes semet ipsos tradiderunt inpudicitiae in operationem inmunditiae omnis in avaritia
EPH|4|20|vos autem non ita didicistis Christum
EPH|4|21|si tamen illum audistis et in ipso edocti estis sicut est veritas in Iesu
EPH|4|22|deponere vos secundum pristinam conversationem veterem hominem qui corrumpitur secundum desideria erroris
EPH|4|23|renovamini autem spiritu mentis vestrae
EPH|4|24|et induite novum hominem qui secundum Deum creatus est in iustitia et sanctitate veritatis
EPH|4|25|propter quod deponentes mendacium loquimini veritatem unusquisque cum proximo suo quoniam sumus invicem membra
EPH|4|26|irascimini et nolite peccare sol non occidat super iracundiam vestram
EPH|4|27|nolite locum dare diabolo
EPH|4|28|qui furabatur iam non furetur magis autem laboret operando manibus quod bonum est ut habeat unde tribuat necessitatem patienti
EPH|4|29|omnis sermo malus ex ore vestro non procedat sed si quis bonus ad aedificationem oportunitatis ut det gratiam audientibus
EPH|4|30|et nolite contristare Spiritum Sanctum Dei in quo signati estis in die redemptionis
EPH|4|31|omnis amaritudo et ira et indignatio et clamor et blasphemia tollatur a vobis cum omni malitia
EPH|4|32|estote autem invicem benigni misericordes donantes invicem sicut et Deus in Christo donavit nobis
EPH|5|1|estote ergo imitatores Dei sicut filii carissimi
EPH|5|2|et ambulate in dilectione sicut et Christus dilexit nos et tradidit se ipsum pro nobis oblationem et hostiam Deo in odorem suavitatis
EPH|5|3|fornicatio autem et omnis inmunditia aut avaritia nec nominetur in vobis sicut decet sanctos
EPH|5|4|aut turpitudo aut stultiloquium aut scurrilitas quae ad rem non pertinent sed magis gratiarum actio
EPH|5|5|hoc enim scitote intellegentes quod omnis fornicator aut inmundus aut avarus quod est idolorum servitus non habet hereditatem in regno Christi et Dei
EPH|5|6|nemo vos seducat inanibus verbis propter haec enim venit ira Dei in filios diffidentiae
EPH|5|7|nolite ergo effici participes eorum
EPH|5|8|eratis enim aliquando tenebrae nunc autem lux in Domino ut filii lucis ambulate
EPH|5|9|fructus enim lucis est in omni bonitate et iustitia et veritate
EPH|5|10|probantes quid sit beneplacitum Deo
EPH|5|11|et nolite communicare operibus infructuosis tenebrarum magis autem et redarguite
EPH|5|12|quae enim in occulto fiunt ab ipsis turpe est et dicere
EPH|5|13|omnia autem quae arguuntur a lumine manifestantur omne enim quod manifestatur lumen est
EPH|5|14|propter quod dicit surge qui dormis et exsurge a mortuis et inluminabit tibi Christus
EPH|5|15|videte itaque fratres quomodo caute ambuletis non quasi insipientes sed ut sapientes
EPH|5|16|redimentes tempus quoniam dies mali sunt
EPH|5|17|propterea nolite fieri inprudentes sed intellegentes quae sit voluntas Domini
EPH|5|18|et nolite inebriari vino in quo est luxuria sed implemini Spiritu
EPH|5|19|loquentes vobismet ipsis in psalmis et hymnis et canticis spiritalibus cantantes et psallentes in cordibus vestris Domino
EPH|5|20|gratias agentes semper pro omnibus in nomine Domini nostri Iesu Christi Deo et Patri
EPH|5|21|subiecti invicem in timore Christi
EPH|5|22|mulieres viris suis subditae sint sicut Domino
EPH|5|23|quoniam vir caput est mulieris sicut Christus caput est ecclesiae ipse salvator corporis
EPH|5|24|sed ut ecclesia subiecta est Christo ita et mulieres viris suis in omnibus
EPH|5|25|viri diligite uxores sicut et Christus dilexit ecclesiam et se ipsum tradidit pro ea
EPH|5|26|ut illam sanctificaret mundans lavacro aquae in verbo
EPH|5|27|ut exhiberet ipse sibi gloriosam ecclesiam non habentem maculam aut rugam aut aliquid eiusmodi sed ut sit sancta et inmaculata
EPH|5|28|ita et viri debent diligere uxores suas ut corpora sua qui suam uxorem diligit se ipsum diligit
EPH|5|29|nemo enim umquam carnem suam odio habuit sed nutrit et fovet eam sicut et Christus ecclesiam
EPH|5|30|quia membra sumus corporis eius de carne eius et de ossibus eius
EPH|5|31|propter hoc relinquet homo patrem et matrem suam et adherebit uxori suae et erunt duo in carne una
EPH|5|32|sacramentum hoc magnum est ego autem dico in Christo et in ecclesia
EPH|5|33|verumtamen et vos singuli unusquisque suam uxorem sicut se ipsum diligat uxor autem ut timeat virum
EPH|6|1|filii oboedite parentibus vestris in Domino hoc enim est iustum
EPH|6|2|honora patrem tuum et matrem quod est mandatum primum in promissione
EPH|6|3|ut bene sit tibi et sis longevus super terram
EPH|6|4|et patres nolite ad iracundiam provocare filios vestros sed educate illos in disciplina et correptione Domini
EPH|6|5|servi oboedite dominis carnalibus cum timore et tremore in simplicitate cordis vestri sicut Christo
EPH|6|6|non ad oculum servientes quasi hominibus placentes sed ut servi Christi facientes voluntatem Dei ex animo
EPH|6|7|cum bona voluntate servientes sicut Domino et non hominibus
EPH|6|8|scientes quoniam unusquisque quodcumque fecerit bonum hoc percipiet a Domino sive servus sive liber
EPH|6|9|et domini eadem facite illis remittentes minas scientes quia et illorum et vester Dominus est in caelis et personarum acceptio non est apud eum
EPH|6|10|de cetero fratres confortamini in Domino et in potentia virtutis eius
EPH|6|11|induite vos arma Dei ut possitis stare adversus insidias diaboli
EPH|6|12|quia non est nobis conluctatio adversus carnem et sanguinem sed adversus principes et potestates adversus mundi rectores tenebrarum harum contra spiritalia nequitiae in caelestibus
EPH|6|13|propterea accipite armaturam Dei ut possitis resistere in die malo et omnibus perfectis stare
EPH|6|14|state ergo succincti lumbos vestros in veritate et induti loricam iustitiae
EPH|6|15|et calciati pedes in praeparatione evangelii pacis
EPH|6|16|in omnibus sumentes scutum fidei in quo possitis omnia tela nequissimi ignea extinguere
EPH|6|17|et galeam salutis adsumite et gladium Spiritus quod est verbum Dei
EPH|6|18|per omnem orationem et obsecrationem orantes omni tempore in Spiritu et in ipso vigilantes in omni instantia et obsecratione pro omnibus sanctis
EPH|6|19|et pro me ut detur mihi sermo in apertione oris mei cum fiducia notum facere mysterium evangelii
EPH|6|20|pro quo legatione fungor in catena ita ut in ipso audeam prout oportet me loqui
EPH|6|21|ut autem et vos sciatis quae circa me sunt quid agam omnia nota vobis faciet Tychicus carissimus frater et fidelis minister in Domino
EPH|6|22|quem misi ad vos in hoc ipsum ut cognoscatis quae circa nos sunt et consoletur corda vestra
EPH|6|23|pax fratribus et caritas cum fide a Deo Patre et Domino Iesu Christo
EPH|6|24|gratia cum omnibus qui diligunt Dominum nostrum Iesum Christum in incorruptione
