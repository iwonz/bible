2THESS|1|1|Paul, Silas and Timothy, To the church of the Thessalonians in God our Father and the Lord Jesus Christ:
2THESS|1|2|Grace and peace to you from God the Father and the Lord Jesus Christ.
2THESS|1|3|We ought always to thank God for you, brothers, and rightly so, because your faith is growing more and more, and the love every one of you has for each other is increasing.
2THESS|1|4|Therefore, among God's churches we boast about your perseverance and faith in all the persecutions and trials you are enduring.
2THESS|1|5|All this is evidence that God's judgment is right, and as a result you will be counted worthy of the kingdom of God, for which you are suffering.
2THESS|1|6|God is just: He will pay back trouble to those who trouble you
2THESS|1|7|and give relief to you who are troubled, and to us as well. This will happen when the Lord Jesus is revealed from heaven in blazing fire with his powerful angels.
2THESS|1|8|He will punish those who do not know God and do not obey the gospel of our Lord Jesus.
2THESS|1|9|They will be punished with everlasting destruction and shut out from the presence of the Lord and from the majesty of his power
2THESS|1|10|on the day he comes to be glorified in his holy people and to be marveled at among all those who have believed. This includes you, because you believed our testimony to you.
2THESS|1|11|With this in mind, we constantly pray for you, that our God may count you worthy of his calling, and that by his power he may fulfill every good purpose of yours and every act prompted by your faith.
2THESS|1|12|We pray this so that the name of our Lord Jesus may be glorified in you, and you in him, according to the grace of our God and the Lord Jesus Christ.
2THESS|2|1|Concerning the coming of our Lord Jesus Christ and our being gathered to him, we ask you, brothers,
2THESS|2|2|not to become easily unsettled or alarmed by some prophecy, report or letter supposed to have come from us, saying that the day of the Lord has already come.
2THESS|2|3|Don't let anyone deceive you in any way, for that day will not come until the rebellion occurs and the man of lawlessness is revealed, the man doomed to destruction.
2THESS|2|4|He will oppose and will exalt himself over everything that is called God or is worshiped, so that he sets himself up in God's temple, proclaiming himself to be God.
2THESS|2|5|Don't you remember that when I was with you I used to tell you these things?
2THESS|2|6|And now you know what is holding him back, so that he may be revealed at the proper time.
2THESS|2|7|For the secret power of lawlessness is already at work; but the one who now holds it back will continue to do so till he is taken out of the way.
2THESS|2|8|And then the lawless one will be revealed, whom the Lord Jesus will overthrow with the breath of his mouth and destroy by the splendor of his coming.
2THESS|2|9|The coming of the lawless one will be in accordance with the work of Satan displayed in all kinds of counterfeit miracles, signs and wonders,
2THESS|2|10|and in every sort of evil that deceives those who are perishing. They perish because they refused to love the truth and so be saved.
2THESS|2|11|For this reason God sends them a powerful delusion so that they will believe the lie
2THESS|2|12|and so that all will be condemned who have not believed the truth but have delighted in wickedness.
2THESS|2|13|But we ought always to thank God for you, brothers loved by the Lord, because from the beginning God chose you to be saved through the sanctifying work of the Spirit and through belief in the truth.
2THESS|2|14|He called you to this through our gospel, that you might share in the glory of our Lord Jesus Christ.
2THESS|2|15|So then, brothers, stand firm and hold to the teachings we passed on to you, whether by word of mouth or by letter.
2THESS|2|16|May our Lord Jesus Christ himself and God our Father, who loved us and by his grace gave us eternal encouragement and good hope,
2THESS|2|17|encourage your hearts and strengthen you in every good deed and word.
2THESS|3|1|Finally, brothers, pray for us that the message of the Lord may spread rapidly and be honored, just as it was with you.
2THESS|3|2|And pray that we may be delivered from wicked and evil men, for not everyone has faith.
2THESS|3|3|But the Lord is faithful, and he will strengthen and protect you from the evil one.
2THESS|3|4|We have confidence in the Lord that you are doing and will continue to do the things we command.
2THESS|3|5|May the Lord direct your hearts into God's love and Christ's perseverance.
2THESS|3|6|In the name of the Lord Jesus Christ, we command you, brothers, to keep away from every brother who is idle and does not live according to the teaching you received from us.
2THESS|3|7|For you yourselves know how you ought to follow our example. We were not idle when we were with you,
2THESS|3|8|nor did we eat anyone's food without paying for it. On the contrary, we worked night and day, laboring and toiling so that we would not be a burden to any of you.
2THESS|3|9|We did this, not because we do not have the right to such help, but in order to make ourselves a model for you to follow.
2THESS|3|10|For even when we were with you, we gave you this rule: "If a man will not work, he shall not eat."
2THESS|3|11|We hear that some among you are idle. They are not busy; they are busybodies.
2THESS|3|12|Such people we command and urge in the Lord Jesus Christ to settle down and earn the bread they eat.
2THESS|3|13|And as for you, brothers, never tire of doing what is right.
2THESS|3|14|If anyone does not obey our instruction in this letter, take special note of him. Do not associate with him, in order that he may feel ashamed.
2THESS|3|15|Yet do not regard him as an enemy, but warn him as a brother.
2THESS|3|16|Now may the Lord of peace himself give you peace at all times and in every way. The Lord be with all of you.
2THESS|3|17|I, Paul, write this greeting in my own hand, which is the distinguishing mark in all my letters. This is how I write.
2THESS|3|18|The grace of our Lord Jesus Christ be with you all.
