2CHR|1|1|Solomon the son of David established himself in his kingdom, and the LORD his God was with him and made him exceedingly great.
2CHR|1|2|Solomon spoke to all Israel, to the commanders of thousands and of hundreds, to the judges, and to all the leaders in all Israel, the heads of fathers' houses.
2CHR|1|3|And Solomon, and all the assembly with him, went to the high place that was at Gibeon, for the tent of meeting of God, which Moses the servant of the LORD had made in the wilderness, was there.
2CHR|1|4|(But David had brought up the ark of God from Kiriath-jearim to the place that David had prepared for it, for he had pitched a tent for it in Jerusalem.)
2CHR|1|5|Moreover, the bronze altar that Bezalel the son of Uri, son of Hur, had made, was there before the tabernacle of the LORD. And Solomon and the assembly resorted to it.
2CHR|1|6|And Solomon went up there to the bronze altar before the LORD, which was at the tent of meeting, and offered a thousand burnt offerings on it.
2CHR|1|7|In that night God appeared to Solomon, and said to him, "Ask what I shall give you."
2CHR|1|8|And Solomon said to God, "You have shown great and steadfast love to David my father, and have made me king in his place.
2CHR|1|9|O LORD God, let your word to David my father be now fulfilled, for you have made me king over a people as numerous as the dust of the earth.
2CHR|1|10|Give me now wisdom and knowledge to go out and come in before this people, for who can govern this people of yours, which is so great?"
2CHR|1|11|God answered Solomon, "Because this was in your heart, and you have not asked possessions, wealth, honor, or the life of those who hate you, and have not even asked long life, but have asked wisdom and knowledge for yourself that you may govern my people over whom I have made you king,
2CHR|1|12|wisdom and knowledge are granted to you. I will also give you riches, possessions, and honor, such as none of the kings had who were before you, and none after you shall have the like."
2CHR|1|13|So Solomon came from the high place at Gibeon, from before the tent of meeting, to Jerusalem. And he reigned over Israel.
2CHR|1|14|Solomon gathered together chariots and horsemen. He had 1,400 chariots and 12,000 horsemen, whom he stationed in the chariot cities and with the king in Jerusalem.
2CHR|1|15|And the king made silver and gold as common in Jerusalem as stone, and he made cedar as plentiful as the sycamore of the Shephelah.
2CHR|1|16|And Solomon's import of horses was from Egypt and Kue, and the king's traders would buy them from Kue for a price.
2CHR|1|17|They imported a chariot from Egypt for 600 shekels of silver, and a horse for 150. Likewise through them these were exported to all the kings of the Hittites and the kings of Syria.
2CHR|2|1|Now Solomon purposed to build a temple for the name of the LORD, and a royal palace for himself.
2CHR|2|2|And Solomon assigned 70,000 men to bear burdens and 80,000 to quarry in the hill country, and 3,600 to oversee them.
2CHR|2|3|And Solomon sent word to Hiram the king of Tyre: "As you dealt with David my father and sent him cedar to build himself a house to dwell in, so deal with me.
2CHR|2|4|Behold, I am about to build a house for the name of the LORD my God and dedicate it to him for the burning of incense of sweet spices before him, and for the regular arrangement of the showbread, and for burnt offerings morning and evening, on the Sabbaths and the new moons and the appointed feasts of the LORD our God, as ordained forever for Israel.
2CHR|2|5|The house that I am to build will be great, for our God is greater than all gods.
2CHR|2|6|But who is able to build him a house, since heaven, even highest heaven, cannot contain him? Who am I to build a house for him, except as a place to make offerings before him?
2CHR|2|7|So now send me a man skilled to work in gold, silver, bronze, and iron, and in purple, crimson, and blue fabrics, trained also in engraving, to be with the skilled workers who are with me in Judah and Jerusalem, whom David my father provided.
2CHR|2|8|Send me also cedar, cypress, and algum timber from Lebanon, for I know that your servants know how to cut timber in Lebanon. And my servants will be with your servants,
2CHR|2|9|to prepare timber for me in abundance, for the house I am to build will be great and wonderful.
2CHR|2|10|I will give for your servants, the woodsmen who cut timber, 20,000 cors of crushed wheat, 20,000 cors of barley, 20,000 baths of wine, and 20,000 baths of oil."
2CHR|2|11|Then Hiram the king of Tyre answered in a letter that he sent to Solomon, "Because the LORD loves his people, he has made you king over them."
2CHR|2|12|Hiram also said, "Blessed be the LORD God of Israel, who made heaven and earth, who has given King David a wise son, who has discretion and understanding, who will build a temple for the LORD and a royal palace for himself.
2CHR|2|13|"Now I have sent a skilled man, who has understanding, Huram-abi,
2CHR|2|14|the son of a woman of the daughters of Dan, and his father was a man of Tyre. He is trained to work in gold, silver, bronze, iron, stone, and wood, and in purple, blue, and crimson fabrics and fine linen, and to do all sorts of engraving and execute any design that may be assigned him, with your craftsmen, the craftsmen of my lord, David your father.
2CHR|2|15|Now therefore the wheat and barley, oil and wine, of which my lord has spoken, let him send to his servants.
2CHR|2|16|And we will cut whatever timber you need from Lebanon and bring it to you in rafts by sea to Joppa, so that you may take it up to Jerusalem."
2CHR|2|17|Then Solomon counted all the resident aliens who were in the land of Israel, after the census of them that David his father had taken, and there were found 153,600.
2CHR|2|18|Seventy thousand of them he assigned to bear burdens, 80,000 to quarry in the hill country, and 3,600 as overseers to make the people work.
2CHR|3|1|Then Solomon began to build the house of the LORD in Jerusalem on Mount Moriah, where the LORD had appeared to David his father, at the place that David had appointed, on the threshing floor of Ornan the Jebusite.
2CHR|3|2|He began to build in the second month of the fourth year of his reign.
2CHR|3|3|These are Solomon's measurements for building the house of God: the length, in cubits of the old standard, was sixty cubits, and the breadth twenty cubits.
2CHR|3|4|The vestibule in front of the nave of the house was twenty cubits long, equal to the width of the house, and its height was 120 cubits. He overlaid it on the inside with pure gold.
2CHR|3|5|The nave he lined with cypress and covered it with fine gold and made palms and chains on it.
2CHR|3|6|He adorned the house with settings of precious stones. The gold was gold of Parvaim.
2CHR|3|7|So he lined the house with gold- its beams, its thresholds, its walls, and its doors- and he carved cherubim on the walls.
2CHR|3|8|And he made the Most Holy Place. Its length, corresponding to the breadth of the house, was twenty cubits, and its breadth was twenty cubits. He overlaid it with 600 talents of fine gold.
2CHR|3|9|The weight of gold for the nails was fifty shekels. And he overlaid the upper chambers with gold.
2CHR|3|10|In the Most Holy Place he made two cherubim of wood and overlaid them with gold.
2CHR|3|11|The wings of the cherubim together extended twenty cubits: one wing of the one, of five cubits, touched the wall of the house, and its other wing, of five cubits, touched the wing of the other cherub;
2CHR|3|12|and of this cherub, one wing, of five cubits, touched the wall of the house, and the other wing, also of five cubits, was joined to the wing of the first cherub.
2CHR|3|13|The wings of these cherubim extended twenty cubits. The cherubim stood on their feet, facing the nave.
2CHR|3|14|And he made the veil of blue and purple and crimson fabrics and fine linen, and he worked cherubim on it.
2CHR|3|15|In front of the house he made two pillars thirty-five cubits high, with a capital of five cubits on the top of each.
2CHR|3|16|He made chains like a necklace and put them on the tops of the pillars, and he made a hundred pomegranates and put them on the chains.
2CHR|3|17|He set up the pillars in front of the temple, one on the south, the other on the north; that on the south he called Jachin, and that on the north Boaz.
2CHR|4|1|He made an altar of bronze, twenty cubits long and twenty cubits wide and ten cubits high.
2CHR|4|2|Then he made the sea of cast metal. It was round, ten cubits from brim to brim, and five cubits high, and a line of thirty cubits measured its circumference.
2CHR|4|3|Under it were figures of gourds, for ten cubits, compassing the sea all around. The gourds were in two rows, cast with it when it was cast.
2CHR|4|4|It stood on twelve oxen, three facing north, three facing west, three facing south, and three facing east. The sea was set on them, and all their rear parts were inward.
2CHR|4|5|Its thickness was a handbreadth. And its brim was made like the brim of a cup, like the flower of a lily. It held 3,000 baths.
2CHR|4|6|He also made ten basins in which to wash, and set five on the south side, and five on the north side. In these they were to rinse off what was used for the burnt offering, and the sea was for the priests to wash in.
2CHR|4|7|And he made ten golden lampstands as prescribed, and set them in the temple, five on the south side and five on the north.
2CHR|4|8|He also made ten tables and placed them in the temple, five on the south side and five on the north. And he made a hundred basins of gold.
2CHR|4|9|He made the court of the priests and the great court and doors for the court and overlaid their doors with bronze.
2CHR|4|10|And he set the sea at the southeast corner of the house.
2CHR|4|11|Hiram also made the pots, the shovels, and the basins. So Hiram finished the work that he did for King Solomon on the house of God:
2CHR|4|12|the two pillars, the bowls, and the two capitals on the top of the pillars; and the two latticeworks to cover the two bowls of the capitals that were on the top of the pillars;
2CHR|4|13|and the 400 pomegranates for the two latticeworks, two rows of pomegranates for each latticework, to cover the two bowls of the capitals that were on the pillars.
2CHR|4|14|He made the stands also, and the basins on the stands,
2CHR|4|15|and the one sea, and the twelve oxen underneath it.
2CHR|4|16|The pots, the shovels, the forks, and all the equipment for these, Huram-abi made of burnished bronze for King Solomon for the house of the LORD.
2CHR|4|17|In the plain of the Jordan the king cast them, in the clay ground between Succoth and Zeredah.
2CHR|4|18|Solomon made all these things in great quantities, for the weight of the bronze was not sought.
2CHR|4|19|So Solomon made all the vessels that were in the house of God: the golden altar, the tables for the bread of the Presence,
2CHR|4|20|the lampstands and their lamps of pure gold to burn before the inner sanctuary, as prescribed;
2CHR|4|21|the flowers, the lamps, and the tongs, of purest gold;
2CHR|4|22|the snuffers, basins, dishes for incense, and fire pans, of pure gold, and the sockets of the temple, for the inner doors to the Most Holy Place and for the doors of the nave of the temple were of gold.
2CHR|5|1|Thus all the work that Solomon did for the house of the LORD was finished. And Solomon brought in the things that David his father had dedicated, and stored the silver, the gold, and all the vessels in the treasuries of the house of God.
2CHR|5|2|Then Solomon assembled the elders of Israel and all the heads of the tribes, the leaders of the fathers' houses of the people of Israel, in Jerusalem, to bring up the ark of the covenant of the LORD out of the city of David, which is Zion.
2CHR|5|3|And all the men of Israel assembled before the king at the feast that is in the seventh month.
2CHR|5|4|And all the elders of Israel came, and the Levites took up the ark.
2CHR|5|5|And they brought up the ark, the tent of meeting, and all the holy vessels that were in the tent; the Levitical priests brought them up.
2CHR|5|6|And King Solomon and all the congregation of Israel, who had assembled before him, were before the ark, sacrificing so many sheep and oxen that they could not be counted or numbered.
2CHR|5|7|Then the priests brought the ark of the covenant of the LORD to its place, in the inner sanctuary of the house, in the Most Holy Place, underneath the wings of the cherubim.
2CHR|5|8|The cherubim spread out their wings over the place of the ark, so that the cherubim made a covering above the ark and its poles.
2CHR|5|9|And the poles were so long that the ends of the poles were seen from the Holy Place before the inner sanctuary, but they could not be seen from outside. And they are there to this day.
2CHR|5|10|There was nothing in the ark except the two tablets that Moses put there at Horeb, where the LORD made a covenant with the people of Israel, when they came out of Egypt.
2CHR|5|11|And when the priests came out of the Holy Place (for all the priests who were present had consecrated themselves, without regard to their divisions,
2CHR|5|12|and all the Levitical singers, Asaph, Heman, and Jeduthun, their sons and kinsmen, arrayed in fine linen, with cymbals, harps, and lyres, stood east of the altar with 120 priests who were trumpeters;
2CHR|5|13|and it was the duty of the trumpeters and singers to make themselves heard in unison in praise and thanksgiving to the LORD), and when the song was raised, with trumpets and cymbals and other musical instruments, in praise to the LORD, "For he is good, for his steadfast love endures forever," the house, the house of the LORD, was filled with a cloud,
2CHR|5|14|so that the priests could not stand to minister because of the cloud, for the glory of the LORD filled the house of God.
2CHR|6|1|Then Solomon said, "The LORD has said that he would dwell in thick darkness.
2CHR|6|2|But I have built you an exalted house, a place for you to dwell in forever."
2CHR|6|3|Then the king turned around and blessed all the assembly of Israel, while all the assembly of Israel stood.
2CHR|6|4|And he said, "Blessed be the LORD, the God of Israel, who with his hand has fulfilled what he promised with his mouth to David my father, saying,
2CHR|6|5|'Since the day that I brought my people out of the land of Egypt, I chose no city out of all the tribes of Israel in which to build a house, that my name might be there, and I chose no man as prince over my people Israel;
2CHR|6|6|but I have chosen Jerusalem that my name may be there, and I have chosen David to be over my people Israel.'
2CHR|6|7|Now it was in the heart of David my father to build a house for the name of the LORD, the God of Israel.
2CHR|6|8|But the LORD said to David my father, 'Whereas it was in your heart to build a house for my name, you did well that it was in your heart.
2CHR|6|9|Nevertheless, it is not you who shall build the house, but your son who shall be born to you shall build the house for my name.'
2CHR|6|10|Now the LORD has fulfilled his promise that he made. For I have risen in the place of David my father and sit on the throne of Israel, as the LORD promised, and I have built the house for the name of the LORD, the God of Israel.
2CHR|6|11|And there I have set the ark, in which is the covenant of the LORD that he made with the people of Israel."
2CHR|6|12|Then Solomon stood before the altar of the LORD in the presence of all the assembly of Israel and spread out his hands.
2CHR|6|13|Solomon had made a bronze platform five cubits long, five cubits wide, and three cubits high, and had set it in the court, and he stood on it. Then he knelt on his knees in the presence of all the assembly of Israel, and spread out his hands toward heaven,
2CHR|6|14|and said, "O LORD, God of Israel, there is no God like you, in heaven or on earth, keeping covenant and showing steadfast love to your servants who walk before you with all their heart,
2CHR|6|15|who have kept with your servant David my father what you declared to him. You spoke with your mouth, and with your hand have fulfilled it this day.
2CHR|6|16|Now therefore, O LORD, God of Israel, keep for your servant David my father what you have promised him, saying, 'You shall not lack a man to sit before me on the throne of Israel, if only your sons pay close attention to their way, to walk in my law as you have walked before me.'
2CHR|6|17|Now therefore, O LORD, God of Israel, let your word be confirmed, which you have spoken to your servant David.
2CHR|6|18|"But will God indeed dwell with man on the earth? Behold, heaven and the highest heaven cannot contain you, how much less this house that I have built!
2CHR|6|19|Yet have regard to the prayer of your servant and to his plea, O LORD my God, listening to the cry and to the prayer that your servant prays before you,
2CHR|6|20|that your eyes may be open day and night toward this house, the place where you have promised to set your name, that you may listen to the prayer that your servant offers toward this place.
2CHR|6|21|And listen to the pleas of your servant and of your people Israel, when they pray toward this place. And listen from heaven your dwelling place, and when you hear, forgive.
2CHR|6|22|"If a man sins against his neighbor and is made to take an oath and comes and swears his oath before your altar in this house,
2CHR|6|23|then hear from heaven and act and judge your servants, repaying the guilty by bringing his conduct on his own head, and vindicating the righteous by rewarding him according to his righteousness.
2CHR|6|24|"If your people Israel are defeated before the enemy because they have sinned against you, and they turn again and acknowledge your name and pray and plead with you in this house,
2CHR|6|25|then hear from heaven and forgive the sin of your people Israel and bring them again to the land that you gave to them and to their fathers.
2CHR|6|26|"When heaven is shut up and there is no rain because they have sinned against you, if they pray toward this place and acknowledge your name and turn from their sin, when you afflict them,
2CHR|6|27|then hear in heaven and forgive the sin of your servants, your people Israel, when you teach them the good way in which they should walk, and grant rain upon your land, which you have given to your people as an inheritance.
2CHR|6|28|"If there is famine in the land, if there is pestilence or blight or mildew or locust or caterpillar, if their enemies besiege them in the land at their gates, whatever plague, whatever sickness there is,
2CHR|6|29|whatever prayer, whatever plea is made by any man or by all your people Israel, each knowing his own affliction and his own sorrow and stretching out his hands toward this house,
2CHR|6|30|then hear from heaven your dwelling place and forgive and render to each whose heart you know, according to all his ways, for you, you only, know the hearts of the children of mankind,
2CHR|6|31|that they may fear you and walk in your ways all the days that they live in the land that you gave to our fathers.
2CHR|6|32|"Likewise, when a foreigner, who is not of your people Israel, comes from a far country for the sake of your great name and your mighty hand and your outstretched arm, when he comes and prays toward this house,
2CHR|6|33|hear from heaven your dwelling place and do according to all for which the foreigner calls to you, in order that all the peoples of the earth may know your name and fear you, as do your people Israel, and that they may know that this house that I have built is called by your name.
2CHR|6|34|"If your people go out to battle against their enemies, by whatever way you shall send them, and they pray to you toward this city that you have chosen and the house that I have built for your name,
2CHR|6|35|then hear from heaven their prayer and their plea, and maintain their cause.
2CHR|6|36|"If they sin against you- for there is no one who does not sin- and you are angry with them and give them to an enemy, so that they are carried away captive to a land far or near,
2CHR|6|37|yet if they turn their heart in the land to which they have been carried captive, and repent and plead with you in the land of their captivity, saying, 'We have sinned and have acted perversely and wickedly,'
2CHR|6|38|if they repent with all their mind and with all their heart in the land of their captivity to which they were carried captive, and pray toward their land, which you gave to their fathers, the city that you have chosen and the house that I have built for your name,
2CHR|6|39|then hear from heaven your dwelling place their prayer and their pleas, and maintain their cause and forgive your people who have sinned against you.
2CHR|6|40|Now, O my God, let your eyes be open and your ears attentive to the prayer of this place.
2CHR|6|41|"And now arise, O LORD God, and go to your resting place, you and the ark of your might. Let your priests, O LORD God, be clothed with salvation, and let your saints rejoice in your goodness.
2CHR|6|42|O LORD God, do not turn away the face of your anointed one! Remember your steadfast love for David your servant."
2CHR|7|1|As soon as Solomon finished his prayer, fire came down from heaven and consumed the burnt offering and the sacrifices, and the glory of the LORD filled the temple.
2CHR|7|2|And the priests could not enter the house of the LORD, because the glory of the LORD filled the LORD's house.
2CHR|7|3|When all the people of Israel saw the fire come down and the glory of the LORD on the temple, they bowed down with their faces to the ground on the pavement and worshiped and gave thanks to the LORD, saying, "For he is good, for his steadfast love endures forever."
2CHR|7|4|Then the king and all the people offered sacrifice before the LORD.
2CHR|7|5|King Solomon offered as a sacrifice 22,000 oxen and 120,000 sheep. So the king and all the people dedicated the house of God.
2CHR|7|6|The priests stood at their posts; the Levites also, with the instruments for music to the LORD that King David had made for giving thanks to the LORD- for his steadfast love endures forever- whenever David offered praises by their ministry; opposite them the priests sounded trumpets, and all Israel stood.
2CHR|7|7|And Solomon consecrated the middle of the court that was before the house of the LORD, for there he offered the burnt offering and the fat of the peace offerings, because the bronze altar Solomon had made could not hold the burnt offering and the grain offering and the fat.
2CHR|7|8|At that time Solomon held the feast for seven days, and all Israel with him, a very great assembly, from Lebo-hamath to the Brook of Egypt.
2CHR|7|9|And on the eighth day they held a solemn assembly, for they had kept the dedication of the altar seven days and the feast seven days.
2CHR|7|10|On the twenty-third day of the seventh month he sent the people away to their homes, joyful and glad of heart for the prosperity that the LORD had granted to David and to Solomon and to Israel his people.
2CHR|7|11|Thus Solomon finished the house of the LORD and the king's house. All that Solomon had planned to do in the house of the LORD and in his own house he successfully accomplished.
2CHR|7|12|Then the LORD appeared to Solomon in the night and said to him: "I have heard your prayer and have chosen this place for myself as a house of sacrifice.
2CHR|7|13|When I shut up the heavens so that there is no rain, or command the locust to devour the land, or send pestilence among my people,
2CHR|7|14|if my people who are called by my name humble themselves, and pray and seek my face and turn from their wicked ways, then I will hear from heaven and will forgive their sin and heal their land.
2CHR|7|15|Now my eyes will be open and my ears attentive to the prayer that is made in this place.
2CHR|7|16|For now I have chosen and consecrated this house that my name may be there forever. My eyes and my heart will be there for all time.
2CHR|7|17|And as for you, if you will walk before me as David your father walked, doing according to all that I have commanded you and keeping my statutes and my rules,
2CHR|7|18|then I will establish your royal throne, as I covenanted with David your father, saying, 'You shall not lack a man to rule Israel.'
2CHR|7|19|"But if you turn aside and forsake my statutes and my commandments that I have set before you, and go and serve other gods and worship them,
2CHR|7|20|then I will pluck you up from my land that I have given you, and this house that I have consecrated for my name, I will cast out of my sight, and I will make it a proverb and a byword among all peoples.
2CHR|7|21|And at this house, which was exalted, everyone passing by will be astonished and say, 'Why has the LORD done thus to this land and to this house?'
2CHR|7|22|Then they will say, 'Because they abandoned the LORD, the God of their fathers who brought them out of the land of Egypt and laid hold on other gods and worshiped them and served them. Therefore he has brought all this disaster on them.'"
2CHR|8|1|At the end of twenty years, in which Solomon had built the house of the LORD and his own house,
2CHR|8|2|Solomon rebuilt the cities that Hiram had given to him, and settled the people of Israel in them.
2CHR|8|3|And Solomon went to Hamath-zobah and took it.
2CHR|8|4|He built Tadmor in the wilderness and all the store cities that he built in Hamath.
2CHR|8|5|He also built Upper Beth-horon and Lower Beth-horon, fortified cities with walls, gates, and bars,
2CHR|8|6|and Baalath, and all the store cities that Solomon had and all the cities for his chariots and the cities for his horsemen, and whatever Solomon desired to build in Jerusalem, in Lebanon, and in all the land of his dominion.
2CHR|8|7|All the people who were left of the Hittites, the Amorites, the Perizzites, the Hivites, and the Jebusites, who were not of Israel,
2CHR|8|8|from their descendants who were left after them in the land, whom the people of Israel had not destroyed- these Solomon drafted as forced labor, and so they are to this day.
2CHR|8|9|But of the people of Israel Solomon made no slaves for his work; they were soldiers, and his officers, the commanders of his chariots, and his horsemen.
2CHR|8|10|And these were the chief officers of King Solomon, 250, who exercised authority over the people.
2CHR|8|11|Solomon brought Pharaoh's daughter up from the city of David to the house that he had built for her, for he said, "My wife shall not live in the house of David king of Israel, for the places to which the ark of the LORD has come are holy."
2CHR|8|12|Then Solomon offered up burnt offerings to the LORD on the altar of the LORD that he had built before the vestibule,
2CHR|8|13|as the duty of each day required, offering according to the commandment of Moses for the Sabbaths, the new moons, and the three annual feasts- the Feast of Unleavened Bread, the Feast of Weeks, and the Feast of Booths.
2CHR|8|14|According to the ruling of David his father, he appointed the divisions of the priests for their service, and the Levites for their offices of praise and ministry before the priests as the duty of each day required, and the gatekeepers in their divisions at each gate, for so David the man of God had commanded.
2CHR|8|15|And they did not turn aside from what the king had commanded the priests and Levites concerning any matter and concerning the treasuries.
2CHR|8|16|Thus was accomplished all the work of Solomon from the day the foundation of the house of the LORD was laid until it was finished. So the house of the LORD was completed.
2CHR|8|17|Then Solomon went to Ezion-geber and Eloth on the shore of the sea, in the land of Edom.
2CHR|8|18|And Hiram sent to him by the hand of his servants ships and servants familiar with the sea, and they went to Ophir together with the servants of Solomon and brought from there 450 talents of gold and brought it to King Solomon.
2CHR|9|1|Now when the queen of Sheba heard of the fame of Solomon, she came to Jerusalem to test him with hard questions, having a very great retinue and camels bearing spices and very much gold and precious stones. And when she came to Solomon, she told him all that was on her mind.
2CHR|9|2|And Solomon answered all her questions. There was nothing hidden from Solomon that he could not explain to her.
2CHR|9|3|And when the queen of Sheba had seen the wisdom of Solomon, the house that he had built,
2CHR|9|4|the food of his table, the seating of his officials, and the attendance of his servants, and their clothing, his cupbearers, and their clothing, and his burnt offerings that he offered at the house of the LORD, there was no more breath in her.
2CHR|9|5|And she said to the king, "The report was true that I heard in my own land of your words and of your wisdom,
2CHR|9|6|but I did not believe the reports until I came and my own eyes had seen it. And behold, half the greatness of your wisdom was not told me; you surpass the report that I heard.
2CHR|9|7|Happy are your wives! Happy are these your servants, who continually stand before you and hear your wisdom!
2CHR|9|8|Blessed be the LORD your God, who has delighted in you and set you on his throne as king for the LORD your God! Because your God loved Israel and would establish them forever, he has made you king over them, that you may execute justice and righteousness."
2CHR|9|9|Then she gave the king 120 talents of gold, and a very great quantity of spices, and precious stones. There were no spices such as those that the queen of Sheba gave to King Solomon.
2CHR|9|10|Moreover, the servants of Hiram and the servants of Solomon, who brought gold from Ophir, brought algum wood and precious stones.
2CHR|9|11|And the king made from the algum wood supports for the house of the LORD and for the king's house, lyres also and harps for the singers. There never was seen the like of them before in the land of Judah.
2CHR|9|12|And King Solomon gave to the queen of Sheba all that she desired, whatever she asked besides what she had brought to the king. So she turned and went back to her own land with her servants.
2CHR|9|13|Now the weight of gold that came to Solomon in one year was 666 talents of gold,
2CHR|9|14|besides that which the explorers and merchants brought. And all the kings of Arabia and the governors of the land brought gold and silver to Solomon.
2CHR|9|15|King Solomon made 200 large shields of beaten gold; 600 shekels of beaten gold went into each shield.
2CHR|9|16|And he made 300 shields of beaten gold; 300 shekels of gold went into each shield; and the king put them in the House of the Forest of Lebanon.
2CHR|9|17|The king also made a great ivory throne and overlaid it with pure gold.
2CHR|9|18|The throne had six steps and a footstool of gold, which were attached to the throne, and on each side of the seat were arm rests and two lions standing beside the arm rests,
2CHR|9|19|while twelve lions stood there, one on each end of a step on the six steps. Nothing like it was ever made for any kingdom.
2CHR|9|20|All King Solomon's drinking vessels were of gold, and all the vessels of the House of the Forest of Lebanon were of pure gold. Silver was not considered as anything in the days of Solomon.
2CHR|9|21|For the king's ships went to Tarshish with the servants of Hiram. Once every three years the ships of Tarshish used to come bringing gold, silver, ivory, apes, and peacocks.
2CHR|9|22|Thus King Solomon excelled all the kings of the earth in riches and in wisdom.
2CHR|9|23|And all the kings of the earth sought the presence of Solomon to hear his wisdom, which God had put into his mind.
2CHR|9|24|Every one of them brought his present, articles of silver and of gold, garments, myrrh, spices, horses, and mules, so much year by year.
2CHR|9|25|And Solomon had 4,000 stalls for horses and chariots, and 12,000 horsemen, whom he stationed in the chariot cities and with the king in Jerusalem.
2CHR|9|26|And he ruled over all the kings from the Euphrates to the land of the Philistines and to the border of Egypt.
2CHR|9|27|And the king made silver as common in Jerusalem as stone, and he made cedar as plentiful as the sycamore of the Shephelah.
2CHR|9|28|And horses were imported for Solomon from Egypt and from all lands.
2CHR|9|29|Now the rest of the acts of Solomon, from first to last, are they not written in the history of Nathan the prophet, and in the prophecy of Ahijah the Shilonite, and in the visions of Iddo the seer concerning Jeroboam the son of Nebat?
2CHR|9|30|Solomon reigned in Jerusalem over all Israel forty years.
2CHR|9|31|And Solomon slept with his fathers and was buried in the city of David his father, and Rehoboam his son reigned in his place.
2CHR|10|1|Rehoboam went to Shechem, for all Israel had come to Shechem to make him king.
2CHR|10|2|And as soon as Jeroboam the son of Nebat heard of it (for he was in Egypt, where he had fled from King Solomon), then Jeroboam returned from Egypt.
2CHR|10|3|And they sent and called him. And Jeroboam and all Israel came and said to Rehoboam,
2CHR|10|4|"Your father made our yoke heavy. Now therefore lighten the hard service of your father and his heavy yoke on us, and we will serve you."
2CHR|10|5|He said to them, "Come to me again in three days." So the people went away.
2CHR|10|6|Then King Rehoboam took counsel with the old men, who had stood before Solomon his father while he was yet alive, saying, "How do you advise me to answer this people?"
2CHR|10|7|And they said to him, "If you will be good to this people and please them and speak good words to them, then they will be your servants forever."
2CHR|10|8|But he abandoned the counsel that the old men gave him, and took counsel with the young men who had grown up with him and stood before him.
2CHR|10|9|And he said to them, "What do you advise that we answer this people who have said to me, 'Lighten the yoke that your father put on us'?"
2CHR|10|10|And the young men who had grown up with him said to him, "Thus shall you speak to the people who said to you, 'Your father made our yoke heavy, but you lighten it for us'; thus shall you say to them, 'My little finger is thicker than my father's thighs.
2CHR|10|11|And now, whereas my father laid on you a heavy yoke, I will add to your yoke. My father disciplined you with whips, but I will discipline you with scorpions.'"
2CHR|10|12|So Jeroboam and all the people came to Rehoboam the third day, as the king said, "Come to me again the third day."
2CHR|10|13|And the king answered them harshly; and forsaking the counsel of the old men,
2CHR|10|14|King Rehoboam spoke to them according to the counsel of the young men, saying, "My father made your yoke heavy, but I will add to it. My father disciplined you with whips, but I will discipline you with scorpions."
2CHR|10|15|So the king did not listen to the people, for it was a turn of affairs brought about by God that the LORD might fulfill his word, which he spoke by Ahijah the Shilonite to Jeroboam the son of Nebat.
2CHR|10|16|And when all Israel saw that the king did not listen to them, the people answered the king, "What portion have we in David? We have no inheritance in the son of Jesse. Each of you to your tents, O Israel! Look now to your own house, David." So all Israel went to their tents.
2CHR|10|17|But Rehoboam reigned over the people of Israel who lived in the cities of Judah.
2CHR|10|18|Then King Rehoboam sent Hadoram, who was taskmaster over the forced labor, and the people of Israel stoned him to death with stones. And King Rehoboam quickly mounted his chariot to flee to Jerusalem.
2CHR|10|19|So Israel has been in rebellion against the house of David to this day.
2CHR|11|1|When Rehoboam came to Jerusalem, he assembled the house of Judah and Benjamin, 180,000 chosen warriors, to fight against Israel, to restore the kingdom to Rehoboam.
2CHR|11|2|But the word of the LORD came to Shemaiah the man of God:
2CHR|11|3|"Say to Rehoboam the son of Solomon, king of Judah, and to all Israel in Judah and Benjamin,
2CHR|11|4|'Thus says the LORD, You shall not go up or fight against your relatives. Return every man to his home, for this thing is from me.'"So they listened to the word of the LORD and returned and did not go against Jeroboam.
2CHR|11|5|Rehoboam lived in Jerusalem, and he built cities for defense in Judah.
2CHR|11|6|He built Bethlehem, Etam, Tekoa,
2CHR|11|7|Beth-zur, Soco, Adullam,
2CHR|11|8|Gath, Mareshah, Ziph,
2CHR|11|9|Adoraim, Lachish, Azekah,
2CHR|11|10|Zorah, Aijalon, and Hebron, fortified cities that are in Judah and in Benjamin.
2CHR|11|11|He made the fortresses strong, and put commanders in them, and stores of food, oil, and wine.
2CHR|11|12|And he put shields and spears in all the cities and made them very strong. So he held Judah and Benjamin.
2CHR|11|13|And the priests and the Levites who were in all Israel presented themselves to him from all places where they lived.
2CHR|11|14|For the Levites left their common lands and their holdings and came to Judah and Jerusalem, because Jeroboam and his sons cast them out from serving as priests of the LORD,
2CHR|11|15|and he appointed his own priests for the high places and for the goat idols and for the calves that he had made.
2CHR|11|16|And those who had set their hearts to seek the LORD God of Israel came after them from all the tribes of Israel to Jerusalem to sacrifice to the LORD, the God of their fathers.
2CHR|11|17|They strengthened the kingdom of Judah, and for three years they made Rehoboam the son of Solomon secure, for they walked for three years in the way of David and Solomon.
2CHR|11|18|Rehoboam took as wife Mahalath the daughter of Jerimoth the son of David, and of Abihail the daughter of Eliab the son of Jesse,
2CHR|11|19|and she bore him sons, Jeush, Shemariah, and Zaham.
2CHR|11|20|After her he took Maacah the daughter of Absalom, who bore him Abijah, Attai, Ziza, and Shelomith.
2CHR|11|21|Rehoboam loved Maacah the daughter of Absalom above all his wives and concubines (he took eighteen wives and sixty concubines, and fathered twenty-eight sons and sixty daughters).
2CHR|11|22|And Rehoboam appointed Abijah the son of Maacah as chief prince among his brothers, for he intended to make him king.
2CHR|11|23|And he dealt wisely and distributed some of his sons through all the districts of Judah and Benjamin, in all the fortified cities, and he gave them abundant provisions and procured wives for them.
2CHR|12|1|When the rule of Rehoboam was established and he was strong, he abandoned the law of the LORD, and all Israel with him.
2CHR|12|2|In the fifth year of King Rehoboam, because they had been unfaithful to the LORD, Shishak king of Egypt came up against Jerusalem
2CHR|12|3|with 1,200 chariots and 60,000 horsemen. And the people were without number who came with him from Egypt- Libyans, Sukkiim, and Ethiopians.
2CHR|12|4|And he took the fortified cities of Judah and came as far as Jerusalem.
2CHR|12|5|Then Shemaiah the prophet came to Rehoboam and to the princes of Judah, who had gathered at Jerusalem because of Shishak, and said to them, "Thus says the LORD, 'You abandoned me, so I have abandoned you to the hand of Shishak.'"
2CHR|12|6|Then the princes of Israel and the king humbled themselves and said, "The LORD is righteous."
2CHR|12|7|When the LORD saw that they humbled themselves, the word of the LORD came to Shemaiah: "They have humbled themselves. I will not destroy them, but I will grant them some deliverance, and my wrath shall not be poured out on Jerusalem by the hand of Shishak.
2CHR|12|8|Nevertheless, they shall be servants to him, that they may know my service and the service of the kingdoms of the countries."
2CHR|12|9|So Shishak king of Egypt came up against Jerusalem. He took away the treasures of the house of the LORD and the treasures of the king's house. He took away everything. He also took away the shields of gold that Solomon had made,
2CHR|12|10|and King Rehoboam made in their place shields of bronze and committed them to the hands of the officers of the guard, who kept the door of the king's house.
2CHR|12|11|And as often as the king went into the house of the LORD, the guard came and carried them and brought them back to the guardroom.
2CHR|12|12|And when he humbled himself the wrath of the LORD turned from him, so as not to make a complete destruction. Moreover, conditions were good in Judah.
2CHR|12|13|So King Rehoboam grew strong in Jerusalem and reigned. Rehoboam was forty-one years old when he began to reign, and he reigned seventeen years in Jerusalem, the city that the LORD had chosen out of all the tribes of Israel to put his name there. His mother's name was Naamah the Ammonite.
2CHR|12|14|And he did evil, for he did not set his heart to seek the LORD.
2CHR|12|15|Now the acts of Rehoboam, from first to last, are they not written in the chronicles of Shemaiah the prophet and of Iddo the seer? There were continual wars between Rehoboam and Jeroboam.
2CHR|12|16|And Rehoboam slept with his fathers and was buried in the city of David, and Abijah his son reigned in his place.
2CHR|13|1|In the eighteenth year of King Jeroboam, Abijah began to reign over Judah.
2CHR|13|2|He reigned for three years in Jerusalem. His mother's name was Micaiah the daughter of Uriel of Gibeah. Now there was war between Abijah and Jeroboam.
2CHR|13|3|Abijah went out to battle, having an army of valiant men of war, 400,000 chosen men. And Jeroboam drew up his line of battle against him with 800,000 chosen mighty warriors.
2CHR|13|4|Then Abijah stood up on Mount Zemaraim that is in the hill country of Ephraim and said, "Hear me, O Jeroboam and all Israel!
2CHR|13|5|Ought you not to know that the LORD God of Israel gave the kingship over Israel forever to David and his sons by a covenant of salt?
2CHR|13|6|Yet Jeroboam the son of Nebat, a servant of Solomon the son of David, rose up and rebelled against his lord,
2CHR|13|7|and certain worthless scoundrels gathered about him and defied Rehoboam the son of Solomon, when Rehoboam was young and irresolute and could not withstand them.
2CHR|13|8|"And now you think to withstand the kingdom of the LORD in the hand of the sons of David, because you are a great multitude and have with you the golden calves that Jeroboam made you for gods.
2CHR|13|9|Have you not driven out the priests of the LORD, the sons of Aaron, and the Levites, and made priests for yourselves like the peoples of other lands? Whoever comes for ordination with a young bull or seven rams becomes a priest of what are no gods.
2CHR|13|10|But as for us, the LORD is our God, and we have not forsaken him. We have priests ministering to the LORD who are sons of Aaron, and Levites for their service.
2CHR|13|11|They offer to the LORD every morning and every evening burnt offerings and incense of sweet spices, set out the showbread on the table of pure gold, and care for the golden lampstand that its lamps may burn every evening. For we keep the charge of the LORD our God, but you have forsaken him.
2CHR|13|12|Behold, God is with us at our head, and his priests with their battle trumpets to sound the call to battle against you. O sons of Israel, do not fight against the LORD, the God of your fathers, for you cannot succeed."
2CHR|13|13|Jeroboam had sent an ambush around to come upon them from behind. Thus his troops were in front of Judah, and the ambush was behind them.
2CHR|13|14|And when Judah looked, behold, the battle was in front of and behind them. And they cried to the LORD, and the priests blew the trumpets.
2CHR|13|15|Then the men of Judah raised the battle shout. And when the men of Judah shouted, God defeated Jeroboam and all Israel before Abijah and Judah.
2CHR|13|16|The men of Israel fled before Judah, and God gave them into their hand.
2CHR|13|17|Abijah and his people struck them with great force, so there fell slain of Israel 500,000 chosen men.
2CHR|13|18|Thus the men of Israel were subdued at that time, and the men of Judah prevailed, because they relied on the LORD, the God of their fathers.
2CHR|13|19|And Abijah pursued Jeroboam and took cities from him, Bethel with its villages and Jeshanah with its villages and Ephron with its villages.
2CHR|13|20|Jeroboam did not recover his power in the days of Abijah. And the LORD struck him down, and he died.
2CHR|13|21|But Abijah grew mighty. And he took fourteen wives and had twenty-two sons and sixteen daughters.
2CHR|13|22|The rest of the acts of Abijah, his ways and his sayings, are written in the story of the prophet Iddo.
2CHR|14|1|Abijah slept with his fathers, and they buried him in the city of David. And Asa his son reigned in his place. In his days the land had rest for ten years.
2CHR|14|2|And Asa did what was good and right in the eyes of the LORD his God.
2CHR|14|3|He took away the foreign altars and the high places and broke down the pillars and cut down the Asherim
2CHR|14|4|and commanded Judah to seek the LORD, the God of their fathers, and to keep the law and the commandment.
2CHR|14|5|He also took out of all the cities of Judah the high places and the incense altars. And the kingdom had rest under him.
2CHR|14|6|He built fortified cities in Judah, for the land had rest. He had no war in those years, for the LORD gave him peace.
2CHR|14|7|And he said to Judah, "Let us build these cities and surround them with walls and towers, gates and bars. The land is still ours, because we have sought the LORD our God. We have sought him, and he has given us peace on every side." So they built and prospered.
2CHR|14|8|And Asa had an army of 300,000 from Judah, armed with large shields and spears, and 280,000 men from Benjamin that carried shields and drew bows. All these were mighty men of valor.
2CHR|14|9|Zerah the Ethiopian came out against them with an army of a million men and 300 chariots, and came as far as Mareshah.
2CHR|14|10|And Asa went out to meet him, and they drew up their lines of battle in the Valley of Zephathah at Mareshah.
2CHR|14|11|And Asa cried to the LORD his God, "O LORD, there is none like you to help, between the mighty and the weak. Help us, O LORD our God, for we rely on you, and in your name we have come against this multitude. O LORD, you are our God; let not man prevail against you."
2CHR|14|12|So the LORD defeated the Ethiopians before Asa and before Judah, and the Ethiopians fled.
2CHR|14|13|Asa and the people who were with him pursued them as far as Gerar, and the Ethiopians fell until none remained alive, for they were broken before the LORD and his army. The men of Judah carried away very much spoil.
2CHR|14|14|And they attacked all the cities around Gerar, for the fear of the LORD was upon them. They plundered all the cities, for there was much plunder in them.
2CHR|14|15|And they struck down the tents of those who had livestock and carried away sheep in abundance and camels. Then they returned to Jerusalem.
2CHR|15|1|The Spirit of God came upon Azariah the son of Oded,
2CHR|15|2|and he went out to meet Asa and said to him, "Hear me, Asa, and all Judah and Benjamin: The LORD is with you while you are with him. If you seek him, he will be found by you, but if you forsake him, he will forsake you.
2CHR|15|3|For a long time Israel was without the true God, and without a teaching priest and without law,
2CHR|15|4|but when in their distress they turned to the LORD, the God of Israel, and sought him, he was found by them.
2CHR|15|5|In those times there was no peace to him who went out or to him who came in, for great disturbances afflicted all the inhabitants of the lands.
2CHR|15|6|They were broken in pieces. Nation was crushed by nation and city by city, for God troubled them with every sort of distress.
2CHR|15|7|But you, take courage! Do not let you hands be weak, for your work shall be rewarded."
2CHR|15|8|As soon as Asa heard these words, the prophecy of Azariah the son of Oded, he took courage and put away the detestable idols from all the land of Judah and Benjamin and from the cities that he had taken in the hill country of Ephraim, and he repaired the altar of the LORD that was in front of the vestibule of the house of the LORD.
2CHR|15|9|And he gathered all Judah and Benjamin, and those from Ephraim, Manasseh, and Simeon who were residing with them, for great numbers had deserted to him from Israel when they saw that the LORD his God was with him.
2CHR|15|10|They were gathered at Jerusalem in the third month of the fifteenth year of the reign of Asa.
2CHR|15|11|They sacrificed to the LORD on that day from the spoil that they had brought 700 oxen and 7,000 sheep.
2CHR|15|12|And they entered into a covenant to seek the LORD, the God of their fathers, with all their heart and with all their soul,
2CHR|15|13|but that whoever would not seek the LORD, the God of Israel, should be put to death, whether young or old, man or woman.
2CHR|15|14|They swore an oath to the LORD with a loud voice and with shouting and with trumpets and with horns.
2CHR|15|15|And all Judah rejoiced over the oath, for they had sworn with all their heart and had sought him with their whole desire, and he was found by them, and the LORD gave them rest all around.
2CHR|15|16|Even Maacah, his mother, King Asa removed from being queen mother because she had made a detestable image for Asherah. Asa cut down her image, crushed it, and burned it at the brook Kidron.
2CHR|15|17|But the high places were not taken out of Israel. Nevertheless, the heart of Asa was wholly true all his days.
2CHR|15|18|And he brought into the house of God the sacred gifts of his father and his own sacred gifts, silver, and gold, and vessels.
2CHR|15|19|And there was no more war until the thirty-fifth year of the reign of Asa.
2CHR|16|1|In the thirty-sixth year of the reign of Asa, Baasha king of Israel went up against Judah and built Ramah, that he might permit no one to go out or come in to Asa king of Judah.
2CHR|16|2|Then Asa took silver and gold from the treasures of the house of the LORD and the king's house and sent them to Ben-hadad king of Syria, who lived in Damascus, saying,
2CHR|16|3|"There is a covenant between me and you, as there was between my father and your father. Behold, I am sending to you silver and gold. Go, break your covenant with Baasha king of Israel, that he may withdraw from me."
2CHR|16|4|And Ben-hadad listened to King Asa and sent the commanders of his armies against the cities of Israel, and they conquered Ijon, Dan, Abel-maim, and all the store cities of Naphtali.
2CHR|16|5|And when Baasha heard of it, he stopped building Ramah and let his work cease.
2CHR|16|6|Then King Asa took all Judah, and they carried away the stones of Ramah and its timber, with which Baasha had been building, and with them he built Geba and Mizpah.
2CHR|16|7|At that time Hanani the seer came to Asa king of Judah and said to him, "Because you relied on the king of Syria, and did not rely on the LORD your God, the army of the king of Syria has escaped you.
2CHR|16|8|Were not the Ethiopians and the Libyans a huge army with very many chariots and horsemen? Yet because you relied on the LORD, he gave them into your hand.
2CHR|16|9|For the eyes of the LORD run to and fro throughout the whole earth, to give strong support to those whose heart is blameless toward him. You have done foolishly in this, for from now on you will have wars."
2CHR|16|10|Then Asa was angry with the seer and put him in the stocks in prison, for he was in a rage with him because of this. And Asa inflicted cruelties upon some of the people at the same time.
2CHR|16|11|The acts of Asa, from first to last, are written in the Book of the Kings of Judah and Israel.
2CHR|16|12|In the thirty-ninth year of his reign Asa was diseased in his feet, and his disease became severe. Yet even in his disease he did not seek the LORD, but sought help from physicians.
2CHR|16|13|And Asa slept with his fathers, dying in the forty-first year of his reign.
2CHR|16|14|They buried him in the tomb that he had cut for himself in the city of David. They laid him on a bier that had been filled with various kinds of spices prepared by the perfumer's art, and they made a very great fire in his honor.
2CHR|17|1|Jehoshaphat his son reigned in his place and strengthened himself against Israel.
2CHR|17|2|He placed forces in all the fortified cities of Judah and set garrisons in the land of Judah, and in the cities of Ephraim that Asa his father had captured.
2CHR|17|3|The LORD was with Jehoshaphat, because he walked in the earlier ways of his father David. He did not seek the Baals,
2CHR|17|4|but sought the God of his father and walked in his commandments, and not according to the practices of Israel.
2CHR|17|5|Therefore the LORD established the kingdom in his hand. And all Judah brought tribute to Jehoshaphat, and he had great riches and honor.
2CHR|17|6|His heart was courageous in the ways of the LORD. And furthermore, he took the high places and the Asherim out of Judah.
2CHR|17|7|In the third year of his reign he sent his officials, Ben-hail, Obadiah, Zechariah, Nethanel, and Micaiah, to teach in the cities of Judah;
2CHR|17|8|and with them the Levites, Shemaiah, Nethaniah, Zebadiah, Asahel, Shemiramoth, Jehonathan, Adonijah, Tobijah, and Tobadonijah; and with these Levites, the priests Elishama and Jehoram.
2CHR|17|9|And they taught in Judah, having the Book of the Law of the LORD with them. They went about through all the cities of Judah and taught among the people.
2CHR|17|10|And the fear of the LORD fell upon all the kingdoms of the lands that were around Judah, and they made no war against Jehoshaphat.
2CHR|17|11|Some of the Philistines brought Jehoshaphat presents and silver for tribute, and the Arabians also brought him 7,700 rams and 7,700 goats.
2CHR|17|12|And Jehoshaphat grew steadily greater. He built in Judah fortresses and store cities,
2CHR|17|13|and he had large supplies in the cities of Judah. He had soldiers, mighty men of valor, in Jerusalem.
2CHR|17|14|This was the muster of them by fathers' houses: Of Judah, the commanders of thousands: Adnah the commander, with 300,000 mighty men of valor;
2CHR|17|15|and next to him Jehohanan the commander, with 280,000;
2CHR|17|16|and next to him Amasiah the son of Zichri, a volunteer for the service of the LORD, with 200,000 mighty men of valor.
2CHR|17|17|Of Benjamin: Eliada, a mighty man of valor, with 200,000 men armed with bow and shield;
2CHR|17|18|and next to him Jehozabad with 180,000 armed for war.
2CHR|17|19|These were in the service of the king, besides those whom the king had placed in the fortified cities throughout all Judah.
2CHR|18|1|Now Jehoshaphat had great riches and honor, and he made a marriage alliance with Ahab.
2CHR|18|2|After some years he went down to Ahab in Samaria. And Ahab killed an abundance of sheep and oxen for him and for the people who were with him, and induced him to go up against Ramoth-gilead.
2CHR|18|3|Ahab king of Israel said to Jehoshaphat king of Judah, "Will you go with me to Ramoth-gilead?" He answered him, "I am as you are, my people as your people. We will be with you in the war."
2CHR|18|4|And Jehoshaphat said to the king of Israel, "Inquire first for the word of the LORD."
2CHR|18|5|Then the king of Israel gathered the prophets together, four hundred men, and said to them, "Shall we go to battle against Ramoth-gilead, or shall I refrain?" And they said, "Go up, for God will give it into the hand of the king."
2CHR|18|6|But Jehoshaphat said, "Is there not here another prophet of the LORD of whom we may inquire?"
2CHR|18|7|And the king of Israel said to Jehoshaphat, "There is yet one man by whom we may inquire of the LORD, Micaiah the son of Imlah; but I hate him, for he never prophesies good concerning me, but always evil." And Jehoshaphat said, "Let not the king say so."
2CHR|18|8|Then the king of Israel summoned an officer and said, "Bring quickly Micaiah the son of Imlah."
2CHR|18|9|Now the king of Israel and Jehoshaphat the king of Judah were sitting on their thrones, arrayed in their robes. And they were sitting at the threshing floor at the entrance of the gate of Samaria, and all the prophets were prophesying before them.
2CHR|18|10|And Zedekiah the son of Chenaanah made for himself horns of iron and said, "Thus says the LORD, 'With these you shall push the Syrians until they are destroyed.'"
2CHR|18|11|And all the prophets prophesied so and said, "Go up to Ramoth-gilead and triumph. The LORD will give it into the hand of the king."
2CHR|18|12|And the messenger who went to summon Micaiah said to him, "Behold, the words of the prophets with one accord are favorable to the king. Let your word be like the word of one of them, and speak favorably."
2CHR|18|13|But Micaiah said, "As the LORD lives, what my God says, that I will speak."
2CHR|18|14|And when he had come to the king, the king said to him, "Micaiah, shall we go to Ramoth-gilead to battle, or shall I refrain?" And he answered, "Go up and triumph; they will be given into your hand."
2CHR|18|15|But the king said to him, "How many times shall I make you swear that you speak to me nothing but the truth in the name of the LORD?"
2CHR|18|16|And he said, "I saw all Israel scattered on the mountains, as sheep that have no shepherd. And the LORD said, 'These have no master; let each return to his home in peace.'"
2CHR|18|17|And the king of Israel said to Jehoshaphat, "Did I not tell you that he would not prophesy good concerning me, but evil?"
2CHR|18|18|And Micaiah said, "Therefore hear the word of the LORD: I saw the LORD sitting on his throne, and all the host of heaven standing on his right hand and on his left.
2CHR|18|19|And the LORD said, 'Who will entice Ahab the king of Israel, that he may go up and fall at Ramoth-gilead?' And one said one thing, and another said another.
2CHR|18|20|Then a spirit came forward and stood before the LORD, saying, 'I will entice him.' And the LORD said to him, 'By what means?'
2CHR|18|21|And he said, 'I will go out, and will be a lying spirit in the mouth of all his prophets.' And he said, 'You are to entice him, and you shall succeed; go out and do so.'
2CHR|18|22|Now therefore behold, the LORD has put a lying spirit in the mouth of these your prophets. The LORD has declared disaster concerning you."
2CHR|18|23|Then Zedekiah the son of Chenaanah came near and struck Micaiah on the cheek and said, "Which way did the Spirit of the LORD go from me to speak to you?"
2CHR|18|24|And Micaiah said, "Behold, you shall see on that day when you go into an inner chamber to hide yourself."
2CHR|18|25|And the king of Israel said, "Seize Micaiah and take him back to Amon the governor of the city and to Joash the king's son,
2CHR|18|26|and say, 'Thus says the king, Put this fellow in prison and feed him with meager rations of bread and water until I return in peace.'"
2CHR|18|27|And Micaiah said, "If you return in peace, the LORD has not spoken by me." And he said, "Hear, all you peoples!"
2CHR|18|28|So the king of Israel and Jehoshaphat the king of Judah went up to Ramoth-gilead.
2CHR|18|29|And the king of Israel said to Jehoshaphat, "I will disguise myself and go into battle, but you wear your robes." And the king of Israel disguised himself, and they went into battle.
2CHR|18|30|Now the king of Syria had commanded the captains of his chariots, "Fight with neither small nor great, but only with the king of Israel."
2CHR|18|31|As soon as the captains of the chariots saw Jehoshaphat, they said, "It is the king of Israel." So they turned to fight against him. And Jehoshaphat cried out, and the LORD helped him; God drew them away from him.
2CHR|18|32|For as soon as the captains of the chariots saw that it was not the king of Israel, they turned back from pursuing him.
2CHR|18|33|But a certain man drew his bow at random and struck the king of Israel between the scale armor and the breastplate. Therefore he said to the driver of his chariot, "Turn around and carry me out of the battle, for I am wounded."
2CHR|18|34|And the battle continued that day, and the king of Israel was propped up in his chariot facing the Syrians until evening. Then at sunset he died.
2CHR|19|1|Jehoshaphat the king of Judah returned in safety to his house in Jerusalem.
2CHR|19|2|But Jehu the son of Hanani the seer went out to meet him and said to King Jehoshaphat, "Should you help the wicked and love those who hate the LORD? Because of this, wrath has gone out against you from the LORD.
2CHR|19|3|Nevertheless, some good is found in you, for you destroyed the Asherahs out of the land, and have set your heart to seek God."
2CHR|19|4|Jehoshaphat lived at Jerusalem. And he went out again among the people, from Beersheba to the hill country of Ephraim, and brought them back to the LORD, the God of their fathers.
2CHR|19|5|He appointed judges in the land in all the fortified cities of Judah, city by city,
2CHR|19|6|and said to the judges, "Consider what you do, for you judge not for man but for the LORD. He is with you in giving judgment.
2CHR|19|7|Now then, let the fear of the LORD be upon you. Be careful what you do, for there is no injustice with the LORD our God, or partiality or taking bribes."
2CHR|19|8|Moreover, in Jerusalem Jehoshaphat appointed certain Levites and priests and heads of families of Israel, to give judgment for the LORD and to decide disputed cases. They had their seat at Jerusalem.
2CHR|19|9|And he charged them: "Thus you shall do in the fear of the LORD, in faithfulness, and with your whole heart:
2CHR|19|10|whenever a case comes to you from your brothers who live in their cities, concerning bloodshed, law or commandment, statutes or rules, then you shall warn them, that they may not incur guilt before the LORD and wrath may not come upon you and your brothers. Thus you shall do, and you will not incur guilt.
2CHR|19|11|And behold, Amariah the chief priest is over you in all matters of the LORD; and Zebadiah the son of Ishmael, the governor of the house of Judah, in all the king's matters, and the Levites will serve you as officers. Deal courageously, and may the LORD be with the upright!"
2CHR|20|1|After this the Moabites and Ammonites, and with them some of the Meunites, came against Jehoshaphat for battle.
2CHR|20|2|Some men came and told Jehoshaphat, "A great multitude is coming against you from Edom, from beyond the sea; and, behold, they are in Hazazon-tamar" (that is, Engedi).
2CHR|20|3|Then Jehoshaphat was afraid and set his face to seek the LORD, and proclaimed a fast throughout all Judah.
2CHR|20|4|And Judah assembled to seek help from the LORD; from all the cities of Judah they came to seek the LORD.
2CHR|20|5|And Jehoshaphat stood in the assembly of Judah and Jerusalem, in the house of the LORD, before the new court,
2CHR|20|6|and said, "O LORD, God of our fathers, are you not God in heaven? You rule over all the kingdoms of the nations. In your hand are power and might, so that none is able to withstand you.
2CHR|20|7|Did you not, our God, drive out the inhabitants of this land before your people Israel, and give it forever to the descendants of Abraham your friend?
2CHR|20|8|And they have lived in it and have built for you in it a sanctuary for your name, saying,
2CHR|20|9|'If disaster comes upon us, the sword, judgment, or pestilence, or famine, we will stand before this house and before you- for your name is in this house- and cry out to you in our affliction, and you will hear and save.'
2CHR|20|10|And now behold, the men of Ammon and Moab and Mount Seir, whom you would not let Israel invade when they came from the land of Egypt, and whom they avoided and did not destroy-
2CHR|20|11|behold, they reward us by coming to drive us out of your possession, which you have given us to inherit.
2CHR|20|12|O our God, will you not execute judgment on them? For we are powerless against this great horde that is coming against us. We do not know what to do, but our eyes are on you."
2CHR|20|13|Meanwhile all Judah stood before the LORD, with their little ones, their wives, and their children.
2CHR|20|14|And the Spirit of the LORD came upon Jahaziel the son of Zechariah, son of Benaiah, son of Jeiel, son of Mattaniah, a Levite of the sons of Asaph, in the midst of the assembly.
2CHR|20|15|And he said, "Listen, all Judah and inhabitants of Jerusalem and King Jehoshaphat: Thus says the LORD to you, 'Do not be afraid and do not be dismayed at this great horde, for the battle is not yours but God's.
2CHR|20|16|Tomorrow go down against them. Behold, they will come up by the ascent of Ziz. You will find them at the end of the valley, east of the wilderness of Jeruel.
2CHR|20|17|You will not need to fight in this battle. Stand firm, hold your position, and see the salvation of the LORD on your behalf, O Judah and Jerusalem.' Do not be afraid and do not be dismayed. Tomorrow go out against them, and the LORD will be with you."
2CHR|20|18|Then Jehoshaphat bowed his head with his face to the ground, and all Judah and the inhabitants of Jerusalem fell down before the LORD, worshiping the LORD.
2CHR|20|19|And the Levites, of the Kohathites and the Korahites, stood up to praise the LORD, the God of Israel, with a very loud voice.
2CHR|20|20|And they rose early in the morning and went out into the wilderness of Tekoa. And when they went out, Jehoshaphat stood and said, "Hear me, Judah and inhabitants of Jerusalem! Believe in the LORD your God, and you will be established; believe his prophets, and you will succeed."
2CHR|20|21|And when he had taken counsel with the people, he appointed those who were to sing to the LORD and praise him in holy attire, as they went before the army, and say, "Give thanks to the LORD, for his steadfast love endures forever."
2CHR|20|22|And when they began to sing and praise, the LORD set an ambush against the men of Ammon, Moab, and Mount Seir, who had come against Judah, so that they were routed.
2CHR|20|23|For the men of Ammon and Moab rose against the inhabitants of Mount Seir, devoting them to destruction, and when they had made an end of the inhabitants of Seir, they all helped to destroy one another.
2CHR|20|24|When Judah came to the watchtower of the wilderness, they looked toward the horde, and behold, there were dead bodies lying on the ground; none had escaped.
2CHR|20|25|When Jehoshaphat and his people came to take their spoil, they found among them, in great numbers, goods, clothing, and precious things, which they took for themselves until they could carry no more. They were three days in taking the spoil, it was so much.
2CHR|20|26|On the fourth day they assembled in the Valley of Beracah, for there they blessed the LORD. Therefore the name of that place has been called the Valley of Beracah to this day.
2CHR|20|27|Then they returned, every man of Judah and Jerusalem, and Jehoshaphat at their head, returning to Jerusalem with joy, for the LORD had made them rejoice over their enemies.
2CHR|20|28|They came to Jerusalem with harps and lyres and trumpets, to the house of the LORD.
2CHR|20|29|And the fear of God came on all the kingdoms of the countries when they heard that the LORD had fought against the enemies of Israel.
2CHR|20|30|So the realm of Jehoshaphat was quiet, for his God gave him rest all around.
2CHR|20|31|Thus Jehoshaphat reigned over Judah. He was thirty-five years old when he began to reign, and he reigned twenty-five years in Jerusalem. His mother's name was Azubah the daughter of Shilhi.
2CHR|20|32|He walked in the way of Asa his father and did not turn aside from it, doing what was right in the sight of the LORD.
2CHR|20|33|The high places, however, were not taken away; the people had not yet set their hearts upon the God of their fathers.
2CHR|20|34|Now the rest of the acts of Jehoshaphat, from first to last, are written in the chronicles of Jehu the son of Hanani, which are recorded in the Book of the Kings of Israel.
2CHR|20|35|After this Jehoshaphat king of Judah joined with Ahaziah king of Israel, who acted wickedly.
2CHR|20|36|He joined him in building ships to go to Tarshish, and they built the ships in Ezion-geber.
2CHR|20|37|Then Eliezer the son of Dodavahu of Mareshah prophesied against Jehoshaphat, saying, "Because you have joined with Ahaziah, the LORD will destroy what you have made." And the ships were wrecked and were not able to go to Tarshish.
2CHR|21|1|Jehoshaphat slept with his fathers and was buried with his fathers in the city of David, and Jehoram his son reigned in his place.
2CHR|21|2|He had brothers, the sons of Jehoshaphat: Azariah, Jehiel, Zechariah, Azariah, Michael, and Shephatiah; all these were the sons of Jehoshaphat king of Judah.
2CHR|21|3|Their father gave them great gifts of silver, gold, and valuable possessions, together with fortified cities in Judah, but he gave the kingdom to Jehoram, because he was the firstborn.
2CHR|21|4|When Jehoram had ascended the throne of his father and was established, he killed all his brothers with the sword, and also some of the princes of Israel.
2CHR|21|5|Jehoram was thirty-two years old when he became king, and he reigned eight years in Jerusalem.
2CHR|21|6|And he walked in the way of the kings of Israel, as the house of Ahab had done, for the daughter of Ahab was his wife. And he did what was evil in the sight of the LORD.
2CHR|21|7|Yet the LORD was not willing to destroy the house of David, because of the covenant that he had made with David, and since he had promised to give a lamp to him and to his sons forever.
2CHR|21|8|In his days Edom revolted from the rule of Judah and set up a king of their own.
2CHR|21|9|Then Jehoram passed over with his commanders and all his chariots, and he rose by night and struck the Edomites who had surrounded him and his chariot commanders.
2CHR|21|10|So Edom revolted from the rule of Judah to this day. At that time Libnah also revolted from his rule, because he had forsaken the LORD, the God of his fathers.
2CHR|21|11|Moreover, he made high places in the hill country of Judah and led the inhabitants of Jerusalem into whoredom and made Judah go astray.
2CHR|21|12|And a letter came to him from Elijah the prophet, saying, "Thus says the LORD, the God of David your father, 'Because you have not walked in the ways of Jehoshaphat your father, or in the ways of Asa king of Judah,
2CHR|21|13|but have walked in the way of the kings of Israel and have enticed Judah and the inhabitants of Jerusalem into whoredom, as the house of Ahab led Israel into whoredom, and also you have killed your brothers, of your father's house, who were better than yourself,
2CHR|21|14|behold, the LORD will bring a great plague on your people, your children, your wives, and all your possessions,
2CHR|21|15|and you yourself will have a severe sickness with a disease of your bowels, until your bowels come out because of the disease, day by day.'"
2CHR|21|16|And the LORD stirred up against Jehoram the anger of the Philistines and of the Arabians who are near the Ethiopians.
2CHR|21|17|And they came up against Judah and invaded it and carried away all the possessions they found that belonged to the king's house, and also his sons and his wives, so that no son was left to him except Jehoahaz, his youngest son.
2CHR|21|18|And after all this the LORD struck him in his bowels with an incurable disease.
2CHR|21|19|In course of time, at the end of two years, his bowels came out because of the disease, and he died in great agony. His people made no fire in his honor, like the fires made for his fathers.
2CHR|21|20|He was thirty-two years old when he began to reign, and he reigned eight years in Jerusalem. And he departed with no one's regret. They buried him in the city of David, but not in the tombs of the kings.
2CHR|22|1|And the inhabitants of Jerusalem made Ahaziah his youngest son king in his place, for the band of men that came with the Arabians to the camp had killed all the older sons. So Ahaziah the son of Jehoram king of Judah reigned.
2CHR|22|2|Ahaziah was twenty-two years old when he began to reign, and he reigned one year in Jerusalem. His mother's name was Athaliah, the granddaughter of Omri.
2CHR|22|3|He also walked in the ways of the house of Ahab, for his mother was his counselor in doing wickedly.
2CHR|22|4|He did what was evil in the sight of the LORD, as the house of Ahab had done. For after the death of his father they were his counselors, to his undoing.
2CHR|22|5|He even followed their counsel and went with Jehoram the son of Ahab king of Israel to make war against Hazael king of Syria at Ramoth-gilead. And the Syrians wounded Joram,
2CHR|22|6|and he returned to be healed in Jezreel of the wounds that he had received at Ramah, when he fought against Hazael king of Syria. And Ahaziah the son of Jehoram king of Judah went down to see Joram the son of Ahab in Jezreel, because he was wounded.
2CHR|22|7|But it was ordained by God that the downfall of Ahaziah should come about through his going to visit Joram. For when he came there, he went out with Jehoram to meet Jehu the son of Nimshi, whom the LORD had anointed to destroy the house of Ahab.
2CHR|22|8|And when Jehu was executing judgment on the house of Ahab, he met the princes of Judah and the sons of Ahaziah's brothers, who attended Ahaziah, and he killed them.
2CHR|22|9|He searched for Ahaziah, and he was captured while hiding in Samaria, and he was brought to Jehu and put to death. They buried him, for they said, "He is the grandson of Jehoshaphat, who sought the LORD with all his heart." And the house of Ahaziah had no one able to rule the kingdom.
2CHR|22|10|Now when Athaliah the mother of Ahaziah saw that her son was dead, she arose and destroyed all the royal family of the house of Judah.
2CHR|22|11|But Jehoshabeath, the daughter of the king, took Joash the son of Ahaziah and stole him away from among the king's sons who were about to be put to death, and she put him and his nurse in a bedroom. Thus Jehoshabeath, the daughter of King Jehoram and wife of Jehoiada the priest, because she was a sister of Ahaziah, hid him from Athaliah, so that she did not put him to death.
2CHR|22|12|And he remained with them six years, hidden in the house of God, while Athaliah reigned over the land.
2CHR|23|1|But in the seventh year Jehoiada took courage and entered into a covenant with the commanders of hundreds, Azariah the son of Jeroham, Ishmael the son of Jehohanan, Azariah the son of Obed, Maaseiah the son of Adaiah, and Elishaphat the son of Zichri.
2CHR|23|2|And they went about through Judah and gathered the Levites from all the cities of Judah, and the heads of fathers' houses of Israel, and they came to Jerusalem.
2CHR|23|3|And all the assembly made a covenant with the king in the house of God. And Jehoiada said to them, "Behold, the king's son! Let him reign, as the LORD spoke concerning the sons of David.
2CHR|23|4|This is the thing that you shall do: of you priests and Levites who come off duty on the Sabbath, one third shall be gatekeepers,
2CHR|23|5|and one third shall be at the king's house and one third at the Gate of the Foundation. And all the people shall be in the courts of the house of the LORD.
2CHR|23|6|Let no one enter the house of the LORD except the priests and ministering Levites. They may enter, for they are holy, but all the people shall keep the charge of the LORD.
2CHR|23|7|The Levites shall surround the king, each with his weapons in his hand. And whoever enters the house shall be put to death. Be with the king when he comes in and when he goes out."
2CHR|23|8|The Levites and all Judah did according to all that Jehoiada the priest commanded, and they each brought his men, who were to go off duty on the Sabbath, with those who were to come on duty on the Sabbath, for Jehoiada the priest did not dismiss the divisions.
2CHR|23|9|And Jehoiada the priest gave to the captains the spears and the large and small shields that had been King David's, which were in the house of God.
2CHR|23|10|And he set all the people as a guard for the king, every man with his weapon in his hand, from the south side of the house to the north side of the house, around the altar and the house.
2CHR|23|11|Then they brought out the king's son and put the crown on him and gave him the testimony. And they proclaimed him king, and Jehoiada and his sons anointed him, and they said, "Long live the king."
2CHR|23|12|When Athaliah heard the noise of the people running and praising the king, she went into the house of the LORD to the people.
2CHR|23|13|And when she looked, there was the king standing by his pillar at the entrance, and the captains and the trumpeters beside the king, and all the people of the land rejoicing and blowing trumpets, and the singers with their musical instruments leading in the celebration. And Athaliah tore her clothes and cried, "Treason! Treason!"
2CHR|23|14|Then Jehoiada the priest brought out the captains who were set over the army, saying to them, "Bring her out between the ranks, and anyone who follows her is to be put to death with the sword." For the priest said, "Do not put her to death in the house of the LORD."
2CHR|23|15|So they laid hands on her, and she went into the entrance of the horse gate of the king's house, and they put her to death there.
2CHR|23|16|And Jehoiada made a covenant between himself and all the people and the king that they should be the LORD's people.
2CHR|23|17|Then all the people went to the house of Baal and tore it down; his altars and his images they broke in pieces, and they killed Mattan the priest of Baal before the altars.
2CHR|23|18|And Jehoiada posted watchmen for the house of the LORD under the direction of the Levitical priests and the Levites whom David had organized to be in charge of the house of the LORD, to offer burnt offerings to the LORD, as it is written in the Law of Moses, with rejoicing and with singing, according to the order of David.
2CHR|23|19|He stationed the gatekeepers at the gates of the house of the LORD so that no one should enter who was in any way unclean.
2CHR|23|20|And he took the captains, the nobles, the governors of the people, and all the people of the land, and they brought the king down from the house of the LORD, marching through the upper gate to the king's house. And they set the king on the royal throne.
2CHR|23|21|So all the people of the land rejoiced, and the city was quiet after Athaliah had been put to death with the sword.
2CHR|24|1|Joash was seven years old when he began to reign, and he reigned forty years in Jerusalem. His mother's name was Zibiah of Beersheba.
2CHR|24|2|And Joash did what was right in the eyes of the LORD all the days of Jehoiada the priest.
2CHR|24|3|Jehoiada got for him two wives, and he had sons and daughters.
2CHR|24|4|After this Joash decided to restore the house of the LORD.
2CHR|24|5|And he gathered the priests and the Levites and said to them, "Go out to the cities of Judah and gather from all Israel money to repair the house of your God from year to year, and see that you act quickly." But the Levites did not act quickly.
2CHR|24|6|So the king summoned Jehoiada the chief and said to him, "Why have you not required the Levites to bring in from Judah and Jerusalem the tax levied by Moses, the servant of the LORD, and the congregation of Israel for the tent of testimony?"
2CHR|24|7|For the sons of Athaliah, that wicked woman, had broken into the house of God, and had also used all the dedicated things of the house of the LORD for the Baals.
2CHR|24|8|So the king commanded, and they made a chest and set it outside the gate of the house of the LORD.
2CHR|24|9|And proclamation was made throughout Judah and Jerusalem to bring in for the LORD the tax that Moses the servant of God laid on Israel in the wilderness.
2CHR|24|10|And all the princes and all the people rejoiced and brought their tax and dropped it into the chest until they had finished.
2CHR|24|11|And whenever the chest was brought to the king's officers by the Levites, when they saw that there was much money in it, the king's secretary and the officer of the chief priest would come and empty the chest and take it and return it to its place. Thus they did day after day, and collected money in abundance.
2CHR|24|12|And the king and Jehoiada gave it to those who had charge of the work of the house of the LORD, and they hired masons and carpenters to restore the house of the LORD, and also workers in iron and bronze to repair the house of the LORD.
2CHR|24|13|So those who were engaged in the work labored, and the repairing went forward in their hands, and they restored the house of God to its proper condition and strengthened it.
2CHR|24|14|And when they had finished, they brought the rest of the money before the king and Jehoiada, and with it were made utensils for the house of the LORD, both for the service and for the burnt offerings, and dishes for incense and vessels of gold and silver. And they offered burnt offerings in the house of the LORD regularly all the days of Jehoiada.
2CHR|24|15|But Jehoiada grew old and full of days, and died. He was 130 years old at his death.
2CHR|24|16|And they buried him in the city of David among the kings, because he had done good in Israel, and toward God and his house.
2CHR|24|17|Now after the death of Jehoiada the princes of Judah came and paid homage to the king. Then the king listened to them.
2CHR|24|18|And they abandoned the house of the LORD, the God of their fathers, and served the Asherim and the idols. And wrath came upon Judah and Jerusalem for this guilt of theirs.
2CHR|24|19|Yet he sent prophets among them to bring them back to the LORD. These testified against them, but they would not pay attention.
2CHR|24|20|Then the Spirit of God clothed Zechariah the son of Jehoiada the priest, and he stood above the people, and said to them, "Thus says God, 'Why do you break the commandments of the LORD, so that you cannot prosper? Because you have forsaken the LORD, he has forsaken you.'"
2CHR|24|21|But they conspired against him, and by command of the king they stoned him with stones in the court of the house of the LORD.
2CHR|24|22|Thus Joash the king did not remember the kindness that Jehoiada, Zechariah's father, had shown him, but killed his son. And when he was dying, he said, "May the LORD see and avenge!"
2CHR|24|23|At the end of the year the army of the Syrians came up against Joash. They came to Judah and Jerusalem and destroyed all the princes of the people from among the people and sent all their spoil to the king of Damascus.
2CHR|24|24|Though the army of the Syrians had come with few men, the LORD delivered into their hand a very great army, because Judah had forsaken the LORD, the God of their fathers. Thus they executed judgment on Joash.
2CHR|24|25|When they had departed from him, leaving him severely wounded, his servants conspired against him because of the blood of the son of Jehoiada the priest, and killed him on his bed. So he died, and they buried him in the city of David, but they did not bury him in the tombs of the kings.
2CHR|24|26|Those who conspired against him were Zabad the son of Shimeath the Ammonite, and Jehozabad the son of Shimrith the Moabite.
2CHR|24|27|Accounts of his sons and of the many oracles against him and of the rebuilding of the house of God are written in the Story of the Book of the Kings. And Amaziah his son reigned in his place.
2CHR|25|1|Amaziah was twenty-five years old when he began to reign, and he reigned twenty-nine years in Jerusalem. His mother's name was Jehoaddan of Jerusalem.
2CHR|25|2|And he did what was right in the eyes of the LORD, yet not with a whole heart.
2CHR|25|3|And as soon as the royal power was firmly his, he killed his servants who had struck down the king his father.
2CHR|25|4|But he did not put their children to death, according to what is written in the Law, in the Book of Moses, where the LORD commanded, "Fathers shall not die because of their children, nor children die because of their fathers, but each one shall die for his own sin."
2CHR|25|5|Then Amaziah assembled the men of Judah and set them by fathers' houses under commanders of thousands and of hundreds for all Judah and Benjamin. He mustered those twenty years old and upward, and found that they were 300,000 choice men, fit for war, able to handle spear and shield.
2CHR|25|6|He hired also 100,000 mighty men of valor from Israel for 100 talents of silver.
2CHR|25|7|But a man of God came to him and said, "O king, do not let the army of Israel go with you, for the LORD is not with Israel, with all these Ephraimites.
2CHR|25|8|But go, act, be strong for the battle. Why should you suppose that God will cast you down before the enemy? For God has power to help or to cast down."
2CHR|25|9|And Amaziah said to the man of God, "But what shall we do about the hundred talents that I have given to the army of Israel?" The man of God answered, "The LORD is able to give you much more than this."
2CHR|25|10|Then Amaziah discharged the army that had come to him from Ephraim to go home again. And they became very angry with Judah and returned home in fierce anger.
2CHR|25|11|But Amaziah took courage and led out his people and went to the Valley of Salt and struck down 10,000 men of Seir.
2CHR|25|12|The men of Judah captured another 10,000 alive and took them to the top of a rock and threw them down from the top of the rock, and they were all dashed to pieces.
2CHR|25|13|But the men of the army whom Amaziah sent back, not letting them go with him to battle, raided the cities of Judah, from Samaria to Beth-horon, and struck down 3,000 people in them and took much spoil.
2CHR|25|14|After Amaziah came from striking down the Edomites, he brought the gods of the men of Seir and set them up as his gods and worshiped them, making offerings to them.
2CHR|25|15|Therefore the LORD was angry with Amaziah and sent to him a prophet, who said to him, "Why have you sought the gods of a people who did not deliver their own people from your hand?"
2CHR|25|16|But as he was speaking, the king said to him, "Have we made you a royal counselor? Stop! Why should you be struck down?" So the prophet stopped, but said, "I know that God has determined to destroy you, because you have done this and have not listened to my counsel."
2CHR|25|17|Then Amaziah king of Judah took counsel and sent to Joash the son of Jehoahaz, son of Jehu, king of Israel, saying, "Come, let us look one another in the face."
2CHR|25|18|And Joash the king of Israel sent word to Amaziah king of Judah, "A thistle on Lebanon sent to a cedar on Lebanon, saying, 'Give your daughter to my son for a wife,' and a wild beast of Lebanon passed by and trampled down the thistle.
2CHR|25|19|You say, 'See, I have struck down Edom,' and your heart has lifted you up in boastfulness. But now stay at home. Why should you provoke trouble so that you fall, you and Judah with you?"
2CHR|25|20|But Amaziah would not listen, for it was of God, in order that he might give them into the hand of their enemies, because they had sought the gods of Edom.
2CHR|25|21|So Joash king of Israel went up, and he and Amaziah king of Judah faced one another in battle at Beth-shemesh, which belongs to Judah.
2CHR|25|22|And Judah was defeated by Israel, and every man fled to his home.
2CHR|25|23|And Joash king of Israel captured Amaziah king of Judah, the son of Joash, son of Ahaziah, at Beth-shemesh, and brought him to Jerusalem and broke down the wall of Jerusalem for 400 cubits, from the Ephraim Gate to the Corner Gate.
2CHR|25|24|And he seized all the gold and silver, and all the vessels that were found in the house of God, in the care of Obed-edom. He seized also the treasuries of the king's house, also hostages, and he returned to Samaria.
2CHR|25|25|Amaziah the son of Joash, king of Judah, lived fifteen years after the death of Joash the son of Jehoahaz, king of Israel.
2CHR|25|26|Now the rest of the deeds of Amaziah, from first to last, are they not written in the Book of the Kings of Judah and Israel?
2CHR|25|27|From the time when he turned away from the LORD they made a conspiracy against him in Jerusalem, and he fled to Lachish. But they sent after him to Lachish and put him to death there.
2CHR|25|28|And they brought him upon horses, and he was buried with his fathers in the city of David.
2CHR|26|1|And all the people of Judah took Uzziah, who was sixteen years old, and made him king instead of his father Amaziah.
2CHR|26|2|He built Eloth and restored it to Judah, after the king slept with his fathers.
2CHR|26|3|Uzziah was sixteen years old when he began to reign, and he reigned fifty-two years in Jerusalem. His mother's name was Jecoliah of Jerusalem.
2CHR|26|4|And he did what was right in the eyes of the LORD, according to all that his father Amaziah had done.
2CHR|26|5|He set himself to seek God in the days of Zechariah, who instructed him in the fear of God, and as long as he sought the LORD, God made him prosper.
2CHR|26|6|He went out and made war against the Philistines and broke through the wall of Gath and the wall of Jabneh and the wall of Ashdod, and he built cities in the territory of Ashdod and elsewhere among the Philistines.
2CHR|26|7|God helped him against the Philistines and against the Arabians who lived in Gurbaal and against the Meunites.
2CHR|26|8|The Ammonites paid tribute to Uzziah, and his fame spread even to the border of Egypt, for he became very strong.
2CHR|26|9|Moreover, Uzziah built towers in Jerusalem at the Corner Gate and at the Valley Gate and at the Angle, and fortified them.
2CHR|26|10|And he built towers in the wilderness and cut out many cisterns, for he had large herds, both in the Shephelah and in the plain, and he had farmers and vinedressers in the hills and in the fertile lands, for he loved the soil.
2CHR|26|11|Moreover, Uzziah had an army of soldiers, fit for war, in divisions according to the numbers in the muster made by Jeiel the secretary and Maaseiah the officer, under the direction of Hananiah, one of the king's commanders.
2CHR|26|12|The whole number of the heads of fathers' houses of mighty men of valor was 2,600.
2CHR|26|13|Under their command was an army of 307,500, who could make war with mighty power, to help the king against the enemy.
2CHR|26|14|And Uzziah prepared for all the army shields, spears, helmets, coats of mail, bows, and stones for slinging.
2CHR|26|15|In Jerusalem he made engines, invented by skillful men, to be on the towers and the corners, to shoot arrows and great stones. And his fame spread far, for he was marvelously helped, till he was strong.
2CHR|26|16|But when he was strong, he grew proud, to his destruction. For he was unfaithful to the LORD his God and entered the temple of the LORD to burn incense on the altar of incense.
2CHR|26|17|But Azariah the priest went in after him, with eighty priests of the LORD who were men of valor,
2CHR|26|18|and they withstood King Uzziah and said to him, "It is not for you, Uzziah, to burn incense to the LORD, but for the priests the sons of Aaron, who are consecrated to burn incense. Go out of the sanctuary, for you have done wrong, and it will bring you no honor from the LORD God."
2CHR|26|19|Then Uzziah was angry. Now he had a censer in his hand to burn incense, and when he became angry with the priests, leprosy broke out on his forehead in the presence of the priests in the house of the LORD, by the altar of incense.
2CHR|26|20|And Azariah the chief priest and all the priests looked at him, and behold, he was leprous in his forehead! And they rushed him out quickly, and he himself hurried to go out, because the LORD had struck him.
2CHR|26|21|And King Uzziah was a leper to the day of his death, and being a leper lived in a separate house, for he was excluded from the house of the LORD. And Jotham his son was over the king's household, governing the people of the land.
2CHR|26|22|Now the rest of the acts of Uzziah, from first to last, Isaiah the prophet the son of Amoz wrote.
2CHR|26|23|And Uzziah slept with his fathers, and they buried him with his fathers in the burial field that belonged to the kings, for they said, "He is a leper." And Jotham his son reigned in his place.
2CHR|27|1|Jotham was twenty-five years old when he began to reign, and he reigned sixteen years in Jerusalem. His mother's name was Jerushah the daughter of Zadok.
2CHR|27|2|And he did what was right in the eyes of the LORD according to all that his father Uzziah had done, except he did not enter the temple of the LORD. But the people still followed corrupt practices.
2CHR|27|3|He built the upper gate of the house of the LORD and did much building on the wall of Ophel.
2CHR|27|4|Moreover, he built cities in the hill country of Judah, and forts and towers on the wooded hills.
2CHR|27|5|He fought with the king of the Ammonites and prevailed against them. And the Ammonites gave him that year 100 talents of silver, and 10,000 cors of wheat and 10,000 of barley. The Ammonites paid him the same amount in the second and the third years.
2CHR|27|6|So Jotham became mighty, because he ordered his ways before the LORD his God.
2CHR|27|7|Now the rest of the acts of Jotham, and all his wars and his ways, behold, they are written in the Book of the Kings of Israel and Judah.
2CHR|27|8|He was twenty-five years old when he began to reign, and he reigned sixteen years in Jerusalem.
2CHR|27|9|And Jotham slept with his fathers, and they buried him in the city of David, and Ahaz his son reigned in his place.
2CHR|28|1|Ahaz was twenty years old when he began to reign, and he reigned sixteen years in Jerusalem. And he did not do what was right in the eyes of the LORD, as his father David had done,
2CHR|28|2|but he walked in the ways of the kings of Israel. He even made metal images for the Baals,
2CHR|28|3|and he made offerings in the Valley of the Son of Hinnom and burned his sons as an offering, according to the abominations of the nations whom the LORD drove out before the people of Israel.
2CHR|28|4|And he sacrificed and made offerings on the high places and on the hills and under every green tree.
2CHR|28|5|Therefore the LORD his God gave him into the hand of the king of Syria, who defeated him and took captive a great number of his people and brought them to Damascus. He was also given into the hand of the king of Israel, who struck him with great force.
2CHR|28|6|For Pekah the son of Remaliah killed 120,000 from Judah in one day, all of them men of valor, because they had forsaken the LORD, the God of their fathers.
2CHR|28|7|And Zichri, a mighty man of Ephraim, killed Maaseiah the king's son and Azrikam the commander of the palace and Elkanah the next in authority to the king.
2CHR|28|8|The men of Israel took captive 200,000 of their relatives, women, sons, and daughters. They also took much spoil from them and brought the spoil to Samaria.
2CHR|28|9|But a prophet of the LORD was there, whose name was Oded, and he went out to meet the army that came to Samaria and said to them, "Behold, because the LORD, the God of your fathers, was angry with Judah, he gave them into your hand, but you have killed them in a rage that has reached up to heaven.
2CHR|28|10|And now you intend to subjugate the people of Judah and Jerusalem, male and female, as your slaves. Have you not sins of your own against the LORD your God?
2CHR|28|11|Now hear me, and send back the captives from your relatives whom you have taken, for the fierce wrath of the LORD is upon you."
2CHR|28|12|Certain chiefs also of the men of Ephraim, Azariah the son of Johanan, Berechiah the son of Meshillemoth, Jehizkiah the son of Shallum, and Amasa the son of Hadlai, stood up against those who were coming from the war
2CHR|28|13|and said to them, "You shall not bring the captives in here, for you propose to bring upon us guilt against the LORD in addition to our present sins and guilt. For our guilt is already great, and there is fierce wrath against Israel."
2CHR|28|14|So the armed men left the captives and the spoil before the princes and all the assembly.
2CHR|28|15|And the men who have been mentioned by name rose and took the captives, and with the spoil they clothed all who were naked among them. They clothed them, gave them sandals, provided them with food and drink, and anointed them, and carrying all the feeble among them on donkeys, they brought them to their kinsfolk at Jericho, the city of palm trees. Then they returned to Samaria.
2CHR|28|16|At that time King Ahaz sent to the king of Assyria for help.
2CHR|28|17|For the Edomites had again invaded and defeated Judah and carried away captives.
2CHR|28|18|And the Philistines had made raids on the cities in the Shephelah and the Negeb of Judah, and had taken Beth-shemesh, Aijalon, Gederoth, Soco with its villages, Timnah with its villages, and Gimzo with its villages. And they settled there.
2CHR|28|19|For the LORD humbled Judah because of Ahaz king of Israel, for he had made Judah act sinfully and had been very unfaithful to the LORD.
2CHR|28|20|So Tiglath-pileser king of Assyria came against him and afflicted him instead of strengthening him.
2CHR|28|21|For Ahaz took a portion from the house of the LORD and the house of the king and of the princes, and gave tribute to the king of Assyria, but it did not help him.
2CHR|28|22|In the time of his distress he became yet more faithless to the LORD- this same King Ahaz.
2CHR|28|23|For he sacrificed to the gods of Damascus that had defeated him and said, "Because the gods of the kings of Syria helped them, I will sacrifice to them that they may help me." But they were the ruin of him and of all Israel.
2CHR|28|24|And Ahaz gathered together the vessels of the house of God and cut in pieces the vessels of the house of God, and he shut up the doors of the house of the LORD, and he made himself altars in every corner of Jerusalem.
2CHR|28|25|In every city of Judah he made high places to make offerings to other gods, provoking to anger the LORD, the God of his fathers.
2CHR|28|26|Now the rest of his acts and all his ways, from first to last, behold, they are written in the Book of the Kings of Judah and Israel.
2CHR|28|27|And Ahaz slept with his fathers, and they buried him in the city, in Jerusalem, for they did not bring him into the tombs of the kings of Israel. And Hezekiah his son reigned in his place.
2CHR|29|1|Hezekiah began to reign when he was twenty-five years old, and he reigned twenty-nine years in Jerusalem. His mother's name was Abijah the daughter of Zechariah.
2CHR|29|2|And he did what was right in the eyes of the LORD, according to all that David his father had done.
2CHR|29|3|In the first year of his reign, in the first month, he opened the doors of the house of the LORD and repaired them.
2CHR|29|4|He brought in the priests and the Levites and assembled them in the square on the east
2CHR|29|5|and said to them, "Hear me, Levites! Now consecrate yourselves, and consecrate the house of the LORD, the God of your fathers, and carry out the filth from the Holy Place.
2CHR|29|6|For our fathers have been unfaithful and have done what was evil in the sight of the LORD our God. They have forsaken him and have turned away their faces from the habitation of the LORD and turned their backs.
2CHR|29|7|They also shut the doors of the vestibule and put out the lamps and have not burned incense or offered burnt offerings in the Holy Place to the God of Israel.
2CHR|29|8|Therefore the wrath of the LORD came on Judah and Jerusalem, and he has made them an object of horror, of astonishment, and of hissing, as you see with your own eyes.
2CHR|29|9|For behold, our fathers have fallen by the sword, and our sons and our daughters and our wives are in captivity for this.
2CHR|29|10|Now it is in my heart to make a covenant with the LORD, the God of Israel, in order that his fierce anger may turn away from us.
2CHR|29|11|My sons, do not now be negligent, for the LORD has chosen you to stand in his presence, to minister to him and to be his ministers and make offerings to him."
2CHR|29|12|Then the Levites arose, Mahath the son of Amasai, and Joel the son of Azariah, of the sons of the Kohathites; and of the sons of Merari, Kish the son of Abdi, and Azariah the son of Jehallelel; and of the Gershonites, Joah the son of Zimmah, and Eden the son of Joah;
2CHR|29|13|and of the sons of Elizaphan, Shimri and Jeuel; and of the sons of Asaph, Zechariah and Mattaniah;
2CHR|29|14|and of the sons of Heman, Jehuel and Shimei; and of the sons of Jeduthun, Shemaiah and Uzziel.
2CHR|29|15|They gathered their brothers and consecrated themselves and went in as the king had commanded, by the words of the LORD, to cleanse the house of the LORD.
2CHR|29|16|The priests went into the inner part of the house of the LORD to cleanse it, and they brought out all the uncleanness that they found in the temple of the LORD into the court of the house of the LORD. And the Levites took it and carried it out to the brook Kidron.
2CHR|29|17|They began to consecrate on the first day of the first month, and on the eighth day of the month they came to the vestibule of the LORD. Then for eight days they consecrated the house of the LORD, and on the sixteenth day of the first month they finished.
2CHR|29|18|Then they went in to Hezekiah the king and said, "We have cleansed all the house of the LORD, the altar of burnt offering and all its utensils, and the table for the showbread and all its utensils.
2CHR|29|19|All the utensils that King Ahaz discarded in his reign when he was faithless, we have made ready and consecrated, and behold, they are before the altar of the LORD."
2CHR|29|20|Then Hezekiah the king rose early and gathered the officials of the city and went up to the house of the LORD.
2CHR|29|21|And they brought seven bulls, seven rams, seven lambs, and seven male goats for a sin offering for the kingdom and for the sanctuary and for Judah. And he commanded the priests the sons of Aaron to offer them on the altar of the LORD.
2CHR|29|22|So they slaughtered the bulls, and the priests received the blood and threw it against the altar. And they slaughtered the rams and their blood was thrown against the altar. And they slaughtered the lambs and their blood was thrown against the altar.
2CHR|29|23|Then the goats for the sin offering were brought to the king and the assembly, and they laid their hands on them,
2CHR|29|24|and the priests slaughtered them and made a sin offering with their blood on the altar, to make atonement for all Israel. For the king commanded that the burnt offering and the sin offering should be made for all Israel.
2CHR|29|25|And he stationed the Levites in the house of the LORD with cymbals, harps, and lyres, according to the commandment of David and of Gad the king's seer and of Nathan the prophet, for the commandment was from the LORD through his prophets.
2CHR|29|26|The Levites stood with the instruments of David, and the priests with the trumpets.
2CHR|29|27|Then Hezekiah commanded that the burnt offering be offered on the altar. And when the burnt offering began, the song to the LORD began also, and the trumpets, accompanied by the instruments of David king of Israel.
2CHR|29|28|The whole assembly worshiped, and the singers sang and the trumpeters sounded. All this continued until the burnt offering was finished.
2CHR|29|29|When the offering was finished, the king and all who were present with him bowed themselves and worshiped.
2CHR|29|30|And Hezekiah the king and the officials commanded the Levites to sing praises to the LORD with the words of David and of Asaph the seer. And they sang praises with gladness, and they bowed down and worshiped.
2CHR|29|31|Then Hezekiah said, "You have now consecrated yourselves to the LORD. Come near; bring sacrifices and thank offerings to the house of the LORD." And the assembly brought sacrifices and thank offerings, and all who were of a willing heart brought burnt offerings.
2CHR|29|32|The number of the burnt offerings that the assembly brought was 70 bulls, 100 rams, and 200 lambs; all these were for a burnt offering to the LORD.
2CHR|29|33|And the consecrated offerings were 600 bulls and 3,000 sheep.
2CHR|29|34|But the priests were too few and could not flay all the burnt offerings, so until other priests had consecrated themselves, their brothers the Levites helped them, until the work was finished- for the Levites were more upright in heart than the priests in consecrating themselves.
2CHR|29|35|Besides the great number of burnt offerings, there was the fat of the peace offerings, and there were the drink offerings for the burnt offerings. Thus the service of the house of the LORD was restored.
2CHR|29|36|And Hezekiah and all the people rejoiced because God had prepared for the people, for the thing came about suddenly.
2CHR|30|1|Hezekiah sent to all Israel and Judah, and wrote letters also to Ephraim and Manasseh, that they should come to the house of the LORD at Jerusalem to keep the Passover to the LORD, the God of Israel.
2CHR|30|2|For the king and his princes and all the assembly in Jerusalem had taken counsel to keep the Passover in the second month-
2CHR|30|3|for they could not keep it at that time because the priests had not consecrated themselves in sufficient number, nor had the people assembled in Jerusalem-
2CHR|30|4|and the plan seemed right to the king and all the assembly.
2CHR|30|5|So they decreed to make a proclamation throughout all Israel, from Beersheba to Dan, that the people should come and keep the Passover to the LORD, the God of Israel, at Jerusalem, for they had not kept it as often as prescribed.
2CHR|30|6|So couriers went throughout all Israel and Judah with letters from the king and his princes, as the king had commanded, saying, "O people of Israel, return to the LORD, the God of Abraham, Isaac, and Israel, that he may turn again to the remnant of you who have escaped from the hand of the kings of Assyria.
2CHR|30|7|Do not be like your fathers and your brothers, who were faithless to the LORD God of their fathers, so that he made them a desolation, as you see.
2CHR|30|8|Do not now be stiff-necked as your fathers were, but yield yourselves to the LORD and come to his sanctuary, which he has consecrated forever, and serve the LORD your God, that his fierce anger may turn away from you.
2CHR|30|9|For if you return to the LORD, your brothers and your children will find compassion with their captors and return to this land. For the LORD your God is gracious and merciful and will not turn away his face from you, if you return to him."
2CHR|30|10|So the couriers went from city to city through the country of Ephraim and Manasseh, and as far as Zebulun, but they laughed them to scorn and mocked them.
2CHR|30|11|However, some men of Asher, of Manasseh, and of Zebulun humbled themselves and came to Jerusalem.
2CHR|30|12|The hand of God was also on Judah to give them one heart to do what the king and the princes commanded by the word of the LORD.
2CHR|30|13|And many people came together in Jerusalem to keep the Feast of Unleavened Bread in the second month, a very great assembly.
2CHR|30|14|They set to work and removed the altars that were in Jerusalem, and all the altars for burning incense they took away and threw into the Kidron valley.
2CHR|30|15|And they slaughtered the Passover lamb on the fourteenth day of the second month. And the priests and the Levites were ashamed, so that they consecrated themselves and brought burnt offerings into the house of the LORD.
2CHR|30|16|They took their accustomed posts according to the Law of Moses the man of God. The priests threw the blood that they received from the hand of the Levites.
2CHR|30|17|For there were many in the assembly who had not consecrated themselves. Therefore the Levites had to slaughter the Passover lamb for everyone who was not clean, to consecrate it to the LORD.
2CHR|30|18|For a majority of the people, many of them from Ephraim, Manasseh, Issachar, and Zebulun, had not cleansed themselves, yet they ate the Passover otherwise than as prescribed. For Hezekiah had prayed for them, saying, "May the good LORD pardon everyone
2CHR|30|19|who sets his heart to seek God, the LORD, the God of his fathers, even though not according to the sanctuary's rules of cleanness."
2CHR|30|20|And the LORD heard Hezekiah and healed the people.
2CHR|30|21|And the people of Israel who were present at Jerusalem kept the Feast of Unleavened Bread seven days with great gladness, and the Levites and the priests praised the LORD day by day, singing with all their might to the LORD.
2CHR|30|22|And Hezekiah spoke encouragingly to all the Levites who showed good skill in the service of the LORD. So they ate the food of the festival for seven days, sacrificing peace offerings and giving thanks to the LORD, the God of their fathers.
2CHR|30|23|Then the whole assembly agreed together to keep the feast for another seven days. So they kept it for another seven days with gladness.
2CHR|30|24|For Hezekiah king of Judah gave the assembly 1,000 bulls and 7,000 sheep for offerings, and the princes gave the assembly 1,000 bulls and 10,000 sheep. And the priests consecrated themselves in great numbers.
2CHR|30|25|The whole assembly of Judah, and the priests and the Levites, and the whole assembly that came out of Israel, and the sojourners who came out of the land of Israel, and the sojourners who lived in Judah, rejoiced.
2CHR|30|26|So there was great joy in Jerusalem, for since the time of Solomon the son of David king of Israel there had been nothing like this in Jerusalem.
2CHR|30|27|Then the priests and the Levites arose and blessed the people, and their voice was heard, and their prayer came to his holy habitation in heaven.
2CHR|31|1|Now when all this was finished, all Israel who were present went out to the cities of Judah and broke in pieces the pillars and cut down the Asherim and broke down the high places and the altars throughout all Judah and Benjamin, and in Ephraim and Manasseh, until they had destroyed them all. Then all the people of Israel returned to their cities, every man to his possession.
2CHR|31|2|And Hezekiah appointed the divisions of the priests and of the Levites, division by division, each according to his service, the priests and the Levites, for burnt offerings and peace offerings, to minister in the gates of the camp of the LORD and to give thanks and praise.
2CHR|31|3|The contribution of the king from his own possessions was for the burnt offerings: the burnt offerings of morning and evening, and the burnt offerings for the Sabbaths, the new moons, and the appointed feasts, as it is written in the Law of the LORD.
2CHR|31|4|And he commanded the people who lived in Jerusalem to give the portion due to the priests and the Levites, that they might give themselves to the Law of the LORD.
2CHR|31|5|As soon as the command was spread abroad, the people of Israel gave in abundance the firstfruits of grain, wine, oil, honey, and of all the produce of the field. And they brought in abundantly the tithe of everything.
2CHR|31|6|And the people of Israel and Judah who lived in the cities of Judah also brought in the tithe of cattle and sheep, and the tithe of the dedicated things that had been dedicated to the LORD their God, and laid them in heaps.
2CHR|31|7|In the third month they began to pile up the heaps, and finished them in the seventh month.
2CHR|31|8|When Hezekiah and the princes came and saw the heaps, they blessed the LORD and his people Israel.
2CHR|31|9|And Hezekiah questioned the priests and the Levites about the heaps.
2CHR|31|10|Azariah the chief priest, who was of the house of Zadok, answered him, "Since they began to bring the contributions into the house of the LORD, we have eaten and had enough and have plenty left, for the LORD has blessed his people, so that we have this large amount left."
2CHR|31|11|Then Hezekiah commanded them to prepare chambers in the house of the LORD, and they prepared them.
2CHR|31|12|And they faithfully brought in the contributions, the tithes, and the dedicated things. The chief officer in charge of them was Conaniah the Levite, with Shimei his brother as second,
2CHR|31|13|while Jehiel, Azaziah, Nahath, Asahel, Jerimoth, Jozabad, Eliel, Ismachiah, Mahath, and Benaiah were overseers assisting Conaniah and Shimei his brother, by the appointment of Hezekiah the king and Azariah the chief officer of the house of God.
2CHR|31|14|And Kore the son of Imnah the Levite, keeper of the east gate, was over the freewill offerings to God, to apportion the contribution reserved for the LORD and the most holy offerings.
2CHR|31|15|Eden, Miniamin, Jeshua, Shemaiah, Amariah, and Shecaniah were faithfully assisting him in the cities of the priests, to distribute the portions to their brothers, old and young alike, by divisions,
2CHR|31|16|except those enrolled by genealogy, males from three years old and upwards- all who entered the house of the LORD as the duty of each day required- for their service according to their offices, by their divisions.
2CHR|31|17|The enrollment of the priests was according to their fathers' houses; that of the Levites from twenty years old and upwards was according to their offices, by their divisions.
2CHR|31|18|They were enrolled with all their little children, their wives, their sons, and their daughters, the whole assembly, for they were faithful in keeping themselves holy.
2CHR|31|19|And for the sons of Aaron, the priests, who were in the fields of common land belonging to their cities, there were men in the several cities who were designated by name to distribute portions to every male among the priests and to everyone among the Levites who was enrolled.
2CHR|31|20|Thus Hezekiah did throughout all Judah, and he did what was good and right and faithful before the LORD his God.
2CHR|31|21|And every work that he undertook in the service of the house of God and in accordance with the law and the commandments, seeking his God, he did with all his heart, and prospered.
2CHR|32|1|After these things and these acts of faithfulness, Sennacherib king of Assyria came and invaded Judah and encamped against the fortified cities, thinking to win them for himself.
2CHR|32|2|And when Hezekiah saw that Sennacherib had come and intended to fight against Jerusalem,
2CHR|32|3|he planned with his officers and his mighty men to stop the water of the springs that were outside the city; and they helped him.
2CHR|32|4|A great many people were gathered, and they stopped all the springs and the brook that flowed through the land, saying, "Why should the kings of Assyria come and find much water?"
2CHR|32|5|He set to work resolutely and built up all the wall that was broken down and raised towers upon it, and outside it he built another wall, and he strengthened the Millo in the city of David. He also made weapons and shields in abundance.
2CHR|32|6|And he set combat commanders over the people and gathered them together to him in the square at the gate of the city and spoke encouragingly to them, saying,
2CHR|32|7|"Be strong and courageous. Do not be afraid or dismayed before the king of Assyria and all the horde that is with him, for there are more with us than with him.
2CHR|32|8|With him is an arm of flesh, but with us is the LORD our God, to help us and to fight our battles." And the people took confidence from the words of Hezekiah king of Judah.
2CHR|32|9|After this, Sennacherib, king of Assyria, who was besieging Lachish with all his forces, sent his servants to Jerusalem to Hezekiah king of Judah and to all the people of Judah who were in Jerusalem, saying,
2CHR|32|10|"Thus says Sennacherib king of Assyria, 'On what are you trusting, that you endure the siege in Jerusalem?
2CHR|32|11|Is not Hezekiah misleading you, that he may give you over to die by famine and by thirst, when he tells you, "The LORD our God will deliver us from the hand of the king of Assyria"?
2CHR|32|12|Has not this same Hezekiah taken away his high places and his altars and commanded Judah and Jerusalem, "Before one altar you shall worship, and on it you shall burn your sacrifices"?
2CHR|32|13|Do you not know what I and my fathers have done to all the peoples of other lands? Were the gods of the nations of those lands at all able to deliver their lands out of my hand?
2CHR|32|14|Who among all the gods of those nations that my fathers devoted to destruction was able to deliver his people from my hand, that your God should be able to deliver you from my hand?
2CHR|32|15|Now, therefore, do not let Hezekiah deceive you or mislead you in this fashion, and do not believe him, for no god of any nation or kingdom has been able to deliver his people from my hand or from the hand of my fathers. How much less will your God deliver you out of my hand!'"
2CHR|32|16|And his servants said still more against the Lord GOD and against his servant Hezekiah.
2CHR|32|17|And he wrote letters to cast contempt on the LORD, the God of Israel and to speak against him, saying, "Like the gods of the nations of the lands who have not delivered their people from my hands, so the God of Hezekiah will not deliver his people from my hand."
2CHR|32|18|And they shouted it with a loud voice in the language of Judah to the people of Jerusalem who were on the wall, to frighten and terrify them, in order that they might take the city.
2CHR|32|19|And they spoke of the God of Jerusalem as they spoke of the gods of the peoples of the earth, which are the work of men's hands.
2CHR|32|20|Then Hezekiah the king and Isaiah the prophet, the son of Amoz, prayed because of this and cried to heaven.
2CHR|32|21|And the LORD sent an angel, who cut off all the mighty warriors and commanders and officers in the camp of the king of Assyria. So he returned with shame of face to his own land. And when he came into the house of his god, some of his own sons struck him down there with the sword.
2CHR|32|22|So the LORD saved Hezekiah and the inhabitants of Jerusalem from the hand of Sennacherib king of Assyria and from the hand of all his enemies, and he provided for them on every side.
2CHR|32|23|And many brought gifts to the LORD to Jerusalem and precious things to Hezekiah king of Judah, so that he was exalted in the sight of all nations from that time onward.
2CHR|32|24|In those days Hezekiah became sick and was at the point of death, and he prayed to the LORD, and he answered him and gave him a sign.
2CHR|32|25|But Hezekiah did not make return according to the benefit done to him, for his heart was proud. Therefore wrath came upon him and Judah and Jerusalem.
2CHR|32|26|But Hezekiah humbled himself for the pride of his heart, both he and the inhabitants of Jerusalem, so that the wrath of the LORD did not come upon them in the days of Hezekiah.
2CHR|32|27|And Hezekiah had very great riches and honor, and he made for himself treasuries for silver, for gold, for precious stones, for spices, for shields, and for all kinds of costly vessels;
2CHR|32|28|storehouses also for the yield of grain, wine, and oil; and stalls for all kinds of cattle, and sheepfolds.
2CHR|32|29|He likewise provided cities for himself, and flocks and herds in abundance, for God had given him very great possessions.
2CHR|32|30|This same Hezekiah closed the upper outlet of the waters of Gihon and directed them down to the west side of the city of David. And Hezekiah prospered in all his works.
2CHR|32|31|And so in the matter of the envoys of the princes of Babylon, who had been sent to him to inquire about the sign that had been done in the land, God left him to himself, in order to test him and to know all that was in his heart.
2CHR|32|32|Now the rest of the acts of Hezekiah and his good deeds, behold, they are written in the vision of Isaiah the prophet the son of Amoz, in the Book of the Kings of Judah and Israel.
2CHR|32|33|And Hezekiah slept with his fathers, and they buried him in the upper part of the tombs of the sons of David, and all Judah and the inhabitants of Jerusalem did him honor at his death. And Manasseh his son reigned in his place.
2CHR|33|1|Manasseh was twelve years old when he began to reign, and he reigned fifty-five years in Jerusalem.
2CHR|33|2|And he did what was evil in the sight of the LORD, according to the abominations of the nations whom the LORD drove out before the people of Israel.
2CHR|33|3|For he rebuilt the high places that his father Hezekiah had broken down, and he erected altars to the Baals, and made Asherahs, and worshiped all the host of heaven and served them.
2CHR|33|4|And he built altars in the house of the LORD, of which the LORD had said, "In Jerusalem shall my name be forever."
2CHR|33|5|And he built altars for all the host of heaven in the two courts of the house of the LORD.
2CHR|33|6|And he burned his sons as an offering in the Valley of the Son of Hinnom, and used fortune-telling and omens and sorcery, and dealt with mediums and with wizards. He did much evil in the sight of the LORD, provoking him to anger.
2CHR|33|7|And the carved image of the idol that he had made he set in the house of God, of which God said to David and to Solomon his son, "In this house, and in Jerusalem, which I have chosen out of all the tribes of Israel, I will put my name forever,
2CHR|33|8|and I will no more remove the foot of Israel from the land that I appointed for your fathers, if only they will be careful to do all that I have commanded them, all the law, the statutes, and the rules given through Moses."
2CHR|33|9|Manasseh led Judah and the inhabitants of Jerusalem astray, to do more evil than the nations whom the LORD destroyed before the people of Israel.
2CHR|33|10|The LORD spoke to Manasseh and to his people, but they paid no attention.
2CHR|33|11|Therefore the LORD brought upon them the commanders of the army of the king of Assyria, who captured Manasseh with hooks and bound him with chains of bronze and brought him to Babylon.
2CHR|33|12|And when he was in distress, he entreated the favor of the LORD his God and humbled himself greatly before the God of his fathers.
2CHR|33|13|He prayed to him, and God was moved by his entreaty and heard his plea and brought him again to Jerusalem into his kingdom. Then Manasseh knew that the LORD was God.
2CHR|33|14|Afterward he built an outer wall for the city of David west of Gihon, in the valley, and for the entrance into the Fish Gate, and carried it around Ophel, and raised it to a very great height. He also put commanders of the army in all the fortified cities in Judah.
2CHR|33|15|And he took away the foreign gods and the idol from the house of the LORD, and all the altars that he had built on the mountain of the house of the LORD and in Jerusalem, and he threw them outside of the city.
2CHR|33|16|He also restored the altar of the LORD and offered on it sacrifices of peace offerings and of thanksgiving, and he commanded Judah to serve the LORD, the God of Israel.
2CHR|33|17|Nevertheless, the people still sacrificed at the high places, but only to the LORD their God.
2CHR|33|18|Now the rest of the acts of Manasseh, and his prayer to his God, and the words of the seers who spoke to him in the name of the LORD, the God of Israel, behold, they are in the Chronicles of the Kings of Israel.
2CHR|33|19|And his prayer, and how God was moved by his entreaty, and all his sin and his faithlessness, and the sites on which he built high places and set up the Asherim and the images, before he humbled himself, behold, they are written in the Chronicles of the Seers.
2CHR|33|20|So Manasseh slept with his fathers, and they buried him in his house, and Amon his son reigned in his place.
2CHR|33|21|Amon was twenty-two years old when he began to reign, and he reigned two years in Jerusalem.
2CHR|33|22|And he did what was evil in the sight of the LORD, as Manasseh his father had done. Amon sacrificed to all the images that Manasseh his father had made, and served them.
2CHR|33|23|And he did not humble himself before the LORD, as Manasseh his father had humbled himself, but this Amon incurred guilt more and more.
2CHR|33|24|And his servants conspired against him and put him to death in his house.
2CHR|33|25|But the people of the land struck down all those who had conspired against King Amon. And the people of the land made Josiah his son king in his place.
2CHR|34|1|Josiah was eight years old when he began to reign, and he reigned thirty-one years in Jerusalem.
2CHR|34|2|And he did what was right in the eyes of the LORD, and walked in the ways of David his father; and he did not turn aside to the right hand or to the left.
2CHR|34|3|For in the eighth year of his reign, while he was yet a boy, he began to seek the God of David his father, and in the twelfth year he began to purge Judah and Jerusalem of the high places, the Asherim, and the carved and the metal images.
2CHR|34|4|And they chopped down the altars of the Baals in his presence, and he cut down the incense altars that stood above them. And he broke in pieces the Asherim and the carved and the metal images, and he made dust of them and scattered it over the graves of those who had sacrificed to them.
2CHR|34|5|He also burned the bones of the priests on their altars and cleansed Judah and Jerusalem.
2CHR|34|6|And in the cities of Manasseh, Ephraim, and Simeon, and as far as Naphtali, in their ruins all around,
2CHR|34|7|he broke down the altars and beat the Asherim and the images into powder and cut down all the incense altars throughout all the land of Israel. Then he returned to Jerusalem.
2CHR|34|8|Now in the eighteenth year of his reign, when he had cleansed the land and the house, he sent Shaphan the son of Azaliah, and Maaseiah the governor of the city, and Joah the son of Joahaz, the recorder, to repair the house of the LORD his God.
2CHR|34|9|They came to Hilkiah the high priest and gave him the money that had been brought into the house of God, which the Levites, the keepers of the threshold, had collected from Manasseh and Ephraim and from all the remnant of Israel and from all Judah and Benjamin and from the inhabitants of Jerusalem.
2CHR|34|10|And they gave it to the workmen who were working in the house of the LORD. And the workmen who were working in the house of the LORD gave it for repairing and restoring the house.
2CHR|34|11|They gave it to the carpenters and the builders to buy quarried stone, and timber for binders and beams for the buildings that the kings of Judah had let go to ruin.
2CHR|34|12|And the men did the work faithfully. Over them were set Jahath and Obadiah the Levites, of the sons of Merari, and Zechariah and Meshullam, of the sons of the Kohathites, to have oversight. The Levites, all who were skillful with instruments of music,
2CHR|34|13|were over the burden bearers and directed all who did work in every kind of service, and some of the Levites were scribes and officials and gatekeepers.
2CHR|34|14|While they were bringing out the money that had been brought into the house of the LORD, Hilkiah the priest found the Book of the Law of the LORD given through Moses.
2CHR|34|15|Then Hilkiah answered and said to Shaphan the secretary, "I have found the Book of the Law in the house of the LORD." And Hilkiah gave the book to Shaphan.
2CHR|34|16|Shaphan brought the book to the king, and further reported to the king, "All that was committed to your servants they are doing.
2CHR|34|17|They have emptied out the money that was found in the house of the LORD and have given it into the hand of the overseers and the workmen."
2CHR|34|18|Then Shaphan the secretary told the king, "Hilkiah the priest has given me a book." And Shaphan read from it before the king.
2CHR|34|19|And when the king heard the words of the Law, he tore his clothes.
2CHR|34|20|And the king commanded Hilkiah, Ahikam the son of Shaphan, Abdon the son of Micah, Shaphan the secretary, and Asaiah the king's servant, saying,
2CHR|34|21|"Go, inquire of the LORD for me and for those who are left in Israel and in Judah, concerning the words of the book that has been found. For great is the wrath of the LORD that is poured out on us, because our fathers have not kept the word of the LORD, to do according to all that is written in this book."
2CHR|34|22|So Hilkiah and those whom the king had sent went to Huldah the prophetess, the wife of Shallum the son of Tokhath, son of Hasrah, keeper of the wardrobe (now she lived in Jerusalem in the Second Quarter) and spoke to her to that effect.
2CHR|34|23|And she said to them, "Thus says the LORD, the God of Israel: 'Tell the man who sent you to me,
2CHR|34|24|Thus says the LORD, behold, I will bring disaster upon this place and upon its inhabitants, all the curses that are written in the book that was read before the king of Judah.
2CHR|34|25|Because they have forsaken me and have made offerings to other gods, that they might provoke me to anger with all the works of their hands, therefore my wrath will be poured out on this place and will not be quenched.
2CHR|34|26|But to the king of Judah, who sent you to inquire of the LORD, thus shall you say to him, Thus says the LORD, the God of Israel: Regarding the words that you have heard,
2CHR|34|27|because your heart was tender and you humbled yourself before God when you heard his words against this place and its inhabitants, and you have humbled yourself before me and have torn your clothes and wept before me, I also have heard you, declares the LORD.
2CHR|34|28|Behold, I will gather you to your fathers, and you shall be gathered to your grave in peace, and your eyes shall not see all the disaster that I will bring upon this place and its inhabitants.'"And they brought back word to the king.
2CHR|34|29|Then the king sent and gathered together all the elders of Judah and Jerusalem.
2CHR|34|30|And the king went up to the house of the LORD, with all the men of Judah and the inhabitants of Jerusalem and the priests and the Levites, all the people both great and small. And he read in their hearing all the words of the Book of the Covenant that had been found in the house of the LORD.
2CHR|34|31|And the king stood in his place and made a covenant before the LORD, to walk after the LORD and to keep his commandments and his testimonies and his statutes, with all his heart and all his soul, to perform the words of the covenant that were written in this book.
2CHR|34|32|Then he made all who were present in Jerusalem and in Benjamin stand to it. And the inhabitants of Jerusalem did according to the covenant of God, the God of their fathers.
2CHR|34|33|And Josiah took away all the abominations from all the territory that belonged to the people of Israel and made all who were present in Israel serve the LORD their God. All his days they did not turn away from following the LORD, the God of their fathers.
2CHR|35|1|Josiah kept a Passover to the LORD in Jerusalem. And they slaughtered the Passover lamb on the fourteenth day of the first month.
2CHR|35|2|He appointed the priests to their offices and encouraged them in the service of the house of the LORD.
2CHR|35|3|And he said to the Levites who taught all Israel and who were holy to the LORD, "Put the holy ark in the house that Solomon the son of David, king of Israel, built. You need not carry it on your shoulders. Now serve the LORD your God and his people Israel.
2CHR|35|4|Prepare yourselves according to your fathers' houses by your divisions, as prescribed in the writing of David king of Israel and the document of Solomon his son.
2CHR|35|5|And stand in the Holy Place according to the groupings of the fathers' houses of your brothers the lay people, and according to the division of the Levites by fathers' household.
2CHR|35|6|And slaughter the Passover lamb, and consecrate yourselves, and prepare for your brothers, to do according to the word of the LORD by Moses."
2CHR|35|7|Then Josiah contributed to the lay people, as Passover offerings for all who were present, lambs and young goats from the flock to the number of 30,000, and 3,000 bulls; these were from the king's possessions.
2CHR|35|8|And his officials contributed willingly to the people, to the priests, and to the Levites. Hilkiah, Zechariah, and Jehiel, the chief officers of the house of God, gave to the priests for the Passover offerings 2,600 Passover lambs and 300 bulls.
2CHR|35|9|Conaniah also, and Shemaiah and Nethanel his brothers, and Hashabiah and Jeiel and Jozabad, the chiefs of the Levites, gave to the Levites for the Passover offerings 5,000 lambs and young goats and 500 bulls.
2CHR|35|10|When the service had been prepared for, the priests stood in their place, and the Levites in their divisions according to the king's command.
2CHR|35|11|And they slaughtered the Passover lamb, and the priests threw the blood that they received from them while the Levites flayed the sacrifices.
2CHR|35|12|And they set aside the burnt offerings that they might distribute them according to the groupings of the fathers' houses of the lay people, to offer to the LORD, as it is written in the Book of Moses. And so they did with the bulls.
2CHR|35|13|And they roasted the Passover lamb with fire according to the rule; and they boiled the holy offerings in pots, in cauldrons, and in pans, and carried them quickly to all the lay people.
2CHR|35|14|And afterward they prepared for themselves and for the priests, because the priests the sons of Aaron were offering the burnt offerings and the fat parts until night; so the Levites prepared for themselves and for the priests the sons of Aaron.
2CHR|35|15|The singers, the sons of Asaph, were in their place according to the command of David, and Asaph, and Heman, and Jeduthun the king's seer; and the gatekeepers were at each gate. They did not need to depart from their service, for their brothers the Levites prepared for them.
2CHR|35|16|So all the service of the LORD was prepared that day, to keep the Passover and to offer burnt offerings on the altar of the LORD, according to the command of King Josiah.
2CHR|35|17|And the people of Israel who were present kept the Passover at that time, and the Feast of Unleavened Bread seven days.
2CHR|35|18|No Passover like it had been kept in Israel since the days of Samuel the prophet. None of the kings of Israel had kept such a Passover as was kept by Josiah, and the priests and the Levites, and all Judah and Israel who were present, and the inhabitants of Jerusalem.
2CHR|35|19|In the eighteenth year of the reign of Josiah this Passover was kept.
2CHR|35|20|After all this, when Josiah had prepared the temple, Neco king of Egypt went up to fight at Carchemish on the Euphrates and Josiah went out to meet him.
2CHR|35|21|But he sent envoys to him, saying, "What have we to do with each other, king of Judah? I am not coming against you this day, but against the house with which I am at war. And God has commanded me to hurry. Cease opposing God, who is with me, lest he destroy you."
2CHR|35|22|Nevertheless, Josiah did not turn away from him, but disguised himself in order to fight with him. He did not listen to the words of Neco from the mouth of God, but came to fight in the plain of Megiddo.
2CHR|35|23|And the archers shot King Josiah. And the king said to his servants, "Take me away, for I am badly wounded."
2CHR|35|24|So his servants took him out of the chariot and carried him in his second chariot and brought him to Jerusalem. And he died and was buried in the tombs of his fathers. All Judah and Jerusalem mourned for Josiah.
2CHR|35|25|Jeremiah also uttered a lament for Josiah; and all the singing men and singing women have spoken of Josiah in their laments to this day. They made these a rule in Israel; behold, they are written in the Laments.
2CHR|35|26|Now the rest of the acts of Josiah, and his good deeds according to what is written in the Law of the LORD,
2CHR|35|27|and his acts, first and last, behold, they are written in the Book of the Kings of Israel and Judah.
2CHR|36|1|The people of the land took Jehoahaz the son of Josiah and made him king in his father's place in Jerusalem.
2CHR|36|2|Jehoahaz was twenty-three years old when he began to reign, and he reigned three months in Jerusalem.
2CHR|36|3|Then the king of Egypt deposed him in Jerusalem and laid on the land a tribute of a hundred talents of silver and a talent of gold.
2CHR|36|4|And the king of Egypt made Eliakim his brother king over Judah and Jerusalem, and changed his name to Jehoiakim. But Neco took Jehoahaz his brother and carried him to Egypt.
2CHR|36|5|Jehoiakim was twenty-five years old when he began to reign, and he reigned eleven years in Jerusalem. He did what was evil in the sight of the LORD his God.
2CHR|36|6|Against him came up Nebuchadnezzar king of Babylon and bound him in chains to take him to Babylon.
2CHR|36|7|Nebuchadnezzar also carried part of the vessels of the house of the LORD to Babylon and put them in his palace in Babylon.
2CHR|36|8|Now the rest of the acts of Jehoiakim, and the abominations that he did, and what was found against him, behold, they are written in the Book of the Kings of Israel and Judah. And Jehoiachin his son reigned in his place.
2CHR|36|9|Jehoiachin was eight years old when he became king, and he reigned three months and ten days in Jerusalem. He did what was evil in the sight of the LORD.
2CHR|36|10|In the spring of the year King Nebuchadnezzar sent and brought him to Babylon, with the precious vessels of the house of the LORD, and made his brother Zedekiah king over Judah and Jerusalem.
2CHR|36|11|Zedekiah was twenty-one years old when he began to reign, and he reigned eleven years in Jerusalem.
2CHR|36|12|He did what was evil in the sight of the LORD his God. He did not humble himself before Jeremiah the prophet, who spoke from the mouth of the LORD.
2CHR|36|13|He also rebelled against King Nebuchadnezzar, who had made him swear by God. He stiffened his neck and hardened his heart against turning to the LORD, the God of Israel.
2CHR|36|14|All the officers of the priests and the people likewise were exceedingly unfaithful, following all the abominations of the nations. And they polluted the house of the LORD that he had made holy in Jerusalem.
2CHR|36|15|The LORD, the God of their fathers, sent persistently to them by his messengers, because he had compassion on his people and on his dwelling place.
2CHR|36|16|But they kept mocking the messengers of God, despising his words and scoffing at his prophets, until the wrath of the LORD rose against his people, until there was no remedy.
2CHR|36|17|Therefore he brought up against them the king of the Chaldeans, who killed their young men with the sword in the house of their sanctuary and had no compassion on young man or virgin, old man or aged. He gave them all into his hand.
2CHR|36|18|And all the vessels of the house of God, great and small, and the treasures of the house of the LORD, and the treasures of the king and of his princes, all these he brought to Babylon.
2CHR|36|19|And they burned the house of God and broke down the wall of Jerusalem and burned all its palaces with fire and destroyed all its precious vessels.
2CHR|36|20|He took into exile in Babylon those who had escaped from the sword, and they became servants to him and to his sons until the establishment of the kingdom of Persia,
2CHR|36|21|to fulfill the word of the LORD by the mouth of Jeremiah, until the land had enjoyed its Sabbaths. All the days that it lay desolate it kept Sabbath, to fulfill seventy years.
2CHR|36|22|Now in the first year of Cyrus king of Persia, that the word of the LORD by the mouth of Jeremiah might be fulfilled, the LORD stirred up the spirit of Cyrus king of Persia, so that he made a proclamation throughout all his kingdom and also put it in writing:
2CHR|36|23|"Thus says Cyrus king of Persia, 'The LORD, the God of heaven, has given me all the kingdoms of the earth, and he has charged me to build him a house at Jerusalem, which is in Judah. Whoever is among you of all his people, may the LORD his God be with him. Let him go up.'"
