GAL|1|1|我使徒 保羅 和所有跟我一起的弟兄，寫信給 加拉太 的眾教會。我作使徒不是由於人，也不是藉著人，而是藉著耶穌基督與使他從死人中復活的父上帝。
GAL|1|2|
GAL|1|3|願恩惠、平安 從我們的父上帝和主耶穌基督歸給你們！
GAL|1|4|基督照我們父上帝的旨意，為我們的罪捨己，要救我們脫離現今這罪惡的世代。
GAL|1|5|願榮耀歸給上帝，直到永永遠遠。阿們！
GAL|1|6|我很驚訝你們這麼快就離開那位藉著基督之 恩呼召你們的上帝，而去隨從別的福音；
GAL|1|7|其實並沒有另一個福音，不過有些人騷擾你們，要把基督的福音更改了。
GAL|1|8|但無論是我們或是天上來的使者，若傳福音給你們 ，與我們所傳給你們的不同，他該受詛咒！
GAL|1|9|我們已經說了，現在我再說，若有人傳福音給你們，與你們以往所領受的不同，他該受詛咒！
GAL|1|10|我現在是要得人的心，還是要得上帝的心呢？難道我在討人的喜歡嗎？我若仍舊想討人的喜歡，我就不是基督的僕人了。
GAL|1|11|弟兄們，我要你們知道，我所傳的福音不是按照人的意思；
GAL|1|12|因為我不是從人領受的，也不是人教導我的，而是藉著耶穌基督的啟示而來。
GAL|1|13|你們聽說過從前我在 猶太 教中的行徑，我怎樣竭力壓迫殘害上帝的教會。
GAL|1|14|在 猶太 教中，我比本國許多同輩的人更激進，為我祖宗的傳統更熱心。
GAL|1|15|然而，那位把我從母腹裏分別出來、又施恩呼召我的上帝 ，既然樂意
GAL|1|16|把他兒子啟示在我心裏，讓我在外邦人中傳揚他，我就沒有跟有血有肉的人商量，
GAL|1|17|也沒有上 耶路撒冷 去見那些比我先作使徒的，惟獨到 阿拉伯 去，後來又回到 大馬士革 。
GAL|1|18|過了三年，我才上 耶路撒冷 去見 磯法 ，和他同住了十五天。
GAL|1|19|至於別的使徒，除了主的兄弟 雅各 ，我都沒有見過。
GAL|1|20|我現在寫給你們的是在上帝面前說的，不說謊話。
GAL|1|21|以後我到了 敘利亞 和 基利家 一帶；
GAL|1|22|那時，在基督裏的 猶太 各教會都沒有見過我的面。
GAL|1|23|不過他們聽說「那從前壓迫我們的，現在竟傳揚他原先所殘害的信仰」。
GAL|1|24|他們就為我的緣故歸榮耀給上帝。
GAL|2|1|過了十四年，我再上 耶路撒冷 去， 巴拿巴 同行，也帶了 提多 一起去。
GAL|2|2|我是奉了啟示上去的；我把在外邦人中所傳的福音對弟兄們說明，我是私下對那些有名望的人說的，免得我現在或是從前都徒然奔跑了。
GAL|2|3|但跟我同去的 提多 ，雖是 希臘 人，也沒有勉強他受割禮；
GAL|2|4|因為有偷著混進來的假弟兄，暗中窺探我們在基督耶穌裏擁有的自由，要使我們作奴隸，
GAL|2|5|可是，為要使福音的真理仍存在你們中間，我們一點也沒有讓步順服他們。
GAL|2|6|至於那些有名望的，不論他們是何等人，都與我無關；上帝不以外貌取人。那些有名望的，並沒有加增我甚麼。
GAL|2|7|相反地，他們看見了主託付我傳福音給未受割禮的人，正如主託付 彼得 傳福音給受割禮的人；
GAL|2|8|那感動 彼得 、叫他為受割禮的人作使徒的，也感動我，叫我為外邦人作使徒。
GAL|2|9|那些被認為是教會柱石的 雅各 、 磯法 、 約翰 知道上帝所賜給我的恩典，就跟我和 巴拿巴 握右手以示合作，同意我們往外邦人那裏去，他們往受割禮的人那裏去。
GAL|2|10|他們只要求我們記念窮人，這也是我一向熱心在做的。
GAL|2|11|後來， 磯法 到了 安提阿 ，因為他有可責之處，我就當面反對他。
GAL|2|12|從 雅各 那裏來的人未到以前，他和外邦人一同吃飯，及至他們來到，他因怕奉割禮的人就退出，跟外邦人疏遠了。
GAL|2|13|其餘的 猶太 人也都隨著他裝假，甚至連 巴拿巴 也隨夥裝假。
GAL|2|14|但我一看見他們做得不對，與福音的真理不合，就在眾人面前對 磯法 說：「你既是 猶太 人，卻按照外邦人的樣子，不按照 猶太 人的樣子生活，怎麼能勉強外邦人按照 猶太 人的樣子生活呢？」
GAL|2|15|我們生來就是 猶太 人，不是外邦罪人；
GAL|2|16|可是我們知道，人稱義不是因律法的行為，而是因信耶穌基督 ，我們也信了基督耶穌，為要使我們因信基督稱義，不因律法的行為稱義，因為，凡血肉之軀沒有一個能因律法的行為稱義。
GAL|2|17|我們若求在基督裏稱義，自己卻還被視為罪人，那麼，基督是罪的用人嗎？絕對不是！
GAL|2|18|如果我重新建造我所拆毀的，這就證明自己是違犯律法的人。
GAL|2|19|我因律法而向律法死了，使我可以向上帝活著。我已經與基督同釘十字架，
GAL|2|20|現在活著的不再是我，乃是基督在我裏面活著；並且我如今在肉身活著，是因信上帝的兒子而活；他是愛我，為我捨己。
GAL|2|21|我不廢掉上帝的恩；如果義是藉著律法而獲得，那麼基督就白白死了。
GAL|3|1|無知的 加拉太 人哪，耶穌基督釘十字架，已經活現在你們眼前，誰又迷惑了你們呢？
GAL|3|2|這是我惟一要問你們的：你們領受了聖靈，是因律法的行為或是因聽信福音呢？
GAL|3|3|你們既然以聖靈開始，如今竟要以肉身終結嗎？你們是這樣的無知嗎？
GAL|3|4|你們受這麼多的苦都是徒然的嗎？如果真是徒然的，
GAL|3|5|那麼，上帝賜給你們聖靈，又在你們中間行異能，是因律法的行為或是因聽信福音呢？
GAL|3|6|正如 亞伯拉罕 「信了上帝，這就算他為義」。
GAL|3|7|所以，你們知道：有信心的人才是 亞伯拉罕 的子孫。
GAL|3|8|聖經既然預先看見上帝要使外邦人因信稱義，預先傳福音給 亞伯拉罕 ，說：「萬國都必因你得福。」
GAL|3|9|可見，那有信心的人和有信心的 亞伯拉罕 一同得福。
GAL|3|10|凡出於律法的行為都是受詛咒的，因為經上記著：「凡不持守律法書上所記的一切而去行的，都是受詛咒的。」
GAL|3|11|沒有一個人靠著律法在上帝面前稱義，這是明顯的，因為經上說：「義人必因信得生。」
GAL|3|12|律法並不出於信，而是說：「行這些事的就必因此得生。」
GAL|3|13|既然基督為我們成了詛咒，就把我們從律法的詛咒中贖出來。因為經上記著：「凡掛在木頭上的都是受詛咒的。」
GAL|3|14|這是要使 亞伯拉罕 的福，因著基督耶穌臨到外邦人，使我們能因信得著所應許的聖靈。
GAL|3|15|弟兄們，我照著人的觀點說，人的遺囑一經確定，沒有人能廢棄或加增。
GAL|3|16|那些應許原是向 亞伯拉罕 和他後裔說的，並不是說「和眾後裔」，指許多人，而是說「和你那個後裔」，指一個人，就是基督。
GAL|3|17|我是這麼說，上帝預先所立的約不能被四百三十年以後的律法廢掉，使應許失效。
GAL|3|18|因為承受產業若是出於律法，就不再是出於應許；但上帝是憑著應許把產業賜給 亞伯拉罕 。
GAL|3|19|這樣說來，為甚麼要有律法呢？律法是為過犯的緣故而加上去的，等候那蒙應許的子孫來到才結束，是藉著天使經中保之手而設立的。
GAL|3|20|但中保本不是為單方設立的；上帝卻是一位。
GAL|3|21|這樣，律法是與上帝的 應許對立嗎？絕對不是！如果律法的頒佈能使人得生命，義就誠然出於律法了。
GAL|3|22|但聖經把萬物都圈在罪裏，為要使因信耶穌基督 而來的應許歸給信的人。
GAL|3|23|但這「信」還未來以前，我們被看守在律法之下，像被圈住，直到那將來的「信」顯明出來。
GAL|3|24|這樣，律法是我們的啟蒙教師，直到基督來了 ，好使我們因信稱義。
GAL|3|25|但這「信」既然來到，我們從此就不在啟蒙教師的手下了。
GAL|3|26|其實，你們藉著信，在基督耶穌裏都成為上帝的兒女。
GAL|3|27|你們凡受洗歸入基督的都披戴基督了：
GAL|3|28|不再分 猶太 人或 希臘 人，不再分為奴的自主的，不再分男的女的，因為你們在基督耶穌裏都成為一了。
GAL|3|29|既然你們屬於基督，你們就是 亞伯拉罕 的子孫，是照著應許承受產業的了。
GAL|4|1|我說，雖然那承受產業的是整個產業的主人，但在未成年的時候卻與奴隸毫無分別，
GAL|4|2|仍是在監護人和管家的手下，直等他父親預定的時候來到。
GAL|4|3|我們也是一樣，在未成年的時候，被世上粗淺的學說 所奴役，也是如此。
GAL|4|4|等到時候成熟，上帝就差遣他的兒子，為女子所生，且生在律法之下，
GAL|4|5|為要把律法之下的人贖出來，使我們獲得兒子的名分。
GAL|4|6|因為你們是兒子，上帝就差他兒子的靈進入我們 的心，呼叫：「阿爸，父！」
GAL|4|7|可見，你不再是奴隸，而是兒子了，既然是兒子，就靠著上帝也成為後嗣了。
GAL|4|8|但從前不認識上帝的時候，你們是給那些本來不是上帝的神明作奴隸；
GAL|4|9|現在你們既然認識上帝，更可說是被上帝所認識的，怎麼還要轉回那懦弱無用的粗淺學說 ，情願再給它們作奴隸呢？
GAL|4|10|你們竟又謹守日子、月份、節期、年份，
GAL|4|11|我為你們擔心，惟恐我在你們身上是枉費工夫了。
GAL|4|12|弟兄們，我勸你們，要像我一樣，因為我也像你們一樣。你們一點沒有虧負我。
GAL|4|13|你們知道，我因為身體有疾病才有第一次傳福音給你們的機會。
GAL|4|14|雖然你們為我身體的緣故受試煉，卻沒有輕看我，也沒有厭棄我，反倒接待我如同上帝的使者，如同基督耶穌。
GAL|4|15|你們當日的好意哪裏去了呢？那時若辦得到，你們就是把自己的眼睛挖出來給我，也都情願。這是我可以給你們作證的。
GAL|4|16|如今我把真理告訴你們，倒成了你們的仇敵嗎？
GAL|4|17|那些熱心待你們的人，不懷好意，是要隔絕你們，好使你們熱心待他們。
GAL|4|18|在善事上，時刻熱心待別人原是好的，卻不只是我與你們同在的時候才這樣。
GAL|4|19|我的孩子們哪，我為你們再受生產之苦，直等到基督成形在你們心裏 。
GAL|4|20|我期望現今就在你們那裏，可以改變我的口氣，因為我為你們心裏難過。
GAL|4|21|你們這願意在律法之下的人，請告訴我，你們沒有聽見律法嗎？
GAL|4|22|因為律法上記著， 亞伯拉罕 有兩個兒子，一個是使女生的，一個是自由的婦人生的。
GAL|4|23|那使女所生的是按著肉體生的；那自由的婦人所生的是憑著應許生的。
GAL|4|24|這是比方：那兩個婦人就是兩個約；一個婦人是出於 西奈山 ，生子為奴，就是 夏甲 。
GAL|4|25|這 夏甲 是指著 阿拉伯 的 西奈山 ，與現在的 耶路撒冷 同類，因為 耶路撒冷 和她的兒女都是為奴的。
GAL|4|26|但另一婦人就是在上的 耶路撒冷 ，是自由的，她是我們的母親。
GAL|4|27|因為經上記著： 不懷孕、不生養的，你要歡樂； 未曾經過產難的，你要高聲歡呼； 因為沒有丈夫的，比有丈夫的有更多的兒女。
GAL|4|28|弟兄們，你們是憑著應許作兒女的，如同 以撒 一樣。
GAL|4|29|當時，那按著肉體生的迫害了那按著聖靈生的，現在也是這樣。
GAL|4|30|然而經上是怎麼說的呢？是說：「把使女和她兒子趕出去！因為使女的兒子絕不能與自由婦人的兒子一同承受產業。」
GAL|4|31|弟兄們，這樣看來，我們不是使女的兒女，而是自由婦人的兒女了。
GAL|5|1|基督釋放了我們，為使我們得自由。所以要站穩了，不要再被奴隸的軛挾制。
GAL|5|2|我— 保羅 告訴你們，你們若受割禮，基督就對你們無益了。
GAL|5|3|我再指著凡受割禮的人確實地說，他有義務遵行全部的律法。
GAL|5|4|你們這要靠律法稱義的是與基督隔絕，從恩典中墜落了。
GAL|5|5|至於我們，我們是靠著聖靈，憑著信心，等候所盼望的義。
GAL|5|6|因為在基督耶穌裏，受割禮不受割禮都沒有功效，惟獨使人發出仁愛的信心才有功效。
GAL|5|7|你們向來跑得好，誰攔阻了你們，使你們不順從真理呢？
GAL|5|8|這樣的勸導不是出於那召你們的。
GAL|5|9|一點麵酵能使全團都發起來。
GAL|5|10|我在主裏深信你們必不懷別樣的心；但騷擾你們的，無論是誰，必須承受懲罰。
GAL|5|11|弟兄們，我若仍舊傳割禮，為甚麼還受迫害呢？若是這樣，十字架絆倒人的地方就沒有了。
GAL|5|12|恨不得那騷擾你們的人把自己閹割了。
GAL|5|13|弟兄們，你們蒙召是要得自由；只是不可把這自由當作放縱情慾的機會，總要用愛心互相服侍。
GAL|5|14|因為全部律法都包括在「愛鄰 如己」這一句話之內了。
GAL|5|15|你們要謹慎，你們若相咬相吞，恐怕要彼此消滅了。
GAL|5|16|我說，你們要順著聖靈而行，絕不可滿足肉體的情慾。
GAL|5|17|因為肉體的情慾和聖靈相爭，聖靈和肉體相爭，這兩個彼此敵對，使你們不能做所願意做的。
GAL|5|18|但你們若被聖靈引導，就不在律法之下。
GAL|5|19|情慾的事都是顯而易見的；就如淫亂、污穢、放蕩、
GAL|5|20|拜偶像、行邪術、仇恨、紛爭、忌恨、憤怒、自私、分派、結黨、
GAL|5|21|嫉妒 、醉酒、荒宴等類。我從前告訴過你們，現在又告訴你們，做這樣事的人必不能承受上帝的國。
GAL|5|22|聖靈的果子就是仁愛、喜樂、和平、忍耐、恩慈、良善、信實、
GAL|5|23|溫柔、節制。這樣的事沒有律法禁止。
GAL|5|24|凡屬基督耶穌 的人，是已經把肉體與肉體的邪情私慾同釘在十字架上了。
GAL|5|25|我們若靠著聖靈而活，也要靠著聖靈行事。
GAL|5|26|不要貪圖虛名，彼此惹氣，互相嫉妒。
GAL|6|1|弟兄們，若有人偶然被過犯所勝，你們屬靈的人就要用溫柔的心把他挽回過來；自己也要留意，免得也被引誘。
GAL|6|2|你們各人的重擔要互相擔當，這樣就會成全 基督的律法。
GAL|6|3|人若沒有甚麼了不起，還自以為了不起的，就是自欺。
GAL|6|4|各人要省察自己的行為；這樣，他所誇口的只在自己，而不在別人。
GAL|6|5|因為人人必須擔當自己的擔子。
GAL|6|6|在真道上受教的，要把一切美好的東西與施教的人分享。
GAL|6|7|不要自欺；上帝是輕慢不得的，因為人種的是甚麼，收的也是甚麼。
GAL|6|8|順著肉體撒種的，必從肉體收敗壞；順著聖靈撒種的，必從聖靈收永生。
GAL|6|9|我們行善不可喪志，因為若不灰心，到了適當的時候就有收成。
GAL|6|10|所以，一有機會就要向眾人行善，向信徒一家的人更要這樣。
GAL|6|11|你們看我親手寫給你們的字是何等的大！
GAL|6|12|那些想要炫耀外表的人才勉強你們受割禮，無非是怕自己為基督的十字架受迫害。
GAL|6|13|他們那些受割禮的，連自己也不守律法；他們要你們受割禮，不過是要拿你們的肉體誇口。
GAL|6|14|但我絕不以別的誇口，只誇我們主耶穌基督的十字架；因這十字架 ，就我而論，世界已經釘在十字架上；就世界而論，我已經釘在十字架上。
GAL|6|15|受割禮或不受割禮都無關緊要，要緊的就是作新造的人。
GAL|6|16|凡照這準則行的人，願平安 憐憫，加給他們，和上帝的 以色列 民。
GAL|6|17|從今以後，不要有人再攪擾我，因為我身上帶著耶穌的印記。
GAL|6|18|弟兄們，願我們主耶穌基督的恩與你們的靈同在。阿們！
