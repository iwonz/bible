HAB|1|1|Пророческое видение, которое видел пророк Аввакум.
HAB|1|2|Доколе, Господи, я буду взывать, и Ты не слышишь, буду вопиять к Тебе о насилии, и Ты не спасаешь?
HAB|1|3|Для чего даешь мне видеть злодейство и смотреть на бедствия? Грабительство и насилие предо мною, и восстает вражда и поднимается раздор.
HAB|1|4|От этого закон потерял силу, и суда правильного нет: так как нечестивый одолевает праведного, то и суд происходит превратный.
HAB|1|5|Посмотрите между народами и внимательно вглядитесь, и вы сильно изумитесь; ибо Я сделаю во дни ваши такое дело, которому вы не поверили бы, если бы вам рассказывали.
HAB|1|6|Ибо вот, Я подниму Халдеев, народ жестокий и необузданный, который ходит по широтам земли, чтобы завладеть не принадлежащими ему селениями.
HAB|1|7|Страшен и грозен он; от него самого происходит суд его и власть его.
HAB|1|8|Быстрее барсов кони его и прытче вечерних волков; скачет в разные стороны конница его; издалека приходят всадники его, прилетают как орел, бросающийся на добычу.
HAB|1|9|Весь он идет для грабежа; устремив лице свое вперед, он забирает пленников, как песок.
HAB|1|10|И над царями он издевается, и князья служат ему посмешищем; над всякою крепостью он смеется: насыплет осадный вал и берет ее.
HAB|1|11|Тогда надмевается дух его, и он ходит и буйствует; сила его – бог его.
HAB|1|12|Но не Ты ли издревле Господь Бог мой, Святый мой? мы не умрем! Ты, Господи, только для суда попустил его. Скала моя! для наказания Ты назначил его.
HAB|1|13|Чистым очам Твоим не свойственно глядеть на злодеяния, и смотреть на притеснение Ты не можешь; для чего же Ты смотришь на злодеев и безмолвствуешь, когда нечестивец поглощает того, кто праведнее его,
HAB|1|14|и оставляешь людей как рыбу в море, как пресмыкающихся, у которых нет властителя?
HAB|1|15|Всех их таскает удою, захватывает в сеть свою и забирает их в неводы свои, и от того радуется и торжествует.
HAB|1|16|За то приносит жертвы сети своей и кадит неводу своему, потому что от них тучна часть его и роскошна пища его.
HAB|1|17|Неужели для этого он должен опорожнять свою сеть и непрестанно избивать народы без пощады?
HAB|2|1|На стражу мою стал я и, стоя на башне, наблюдал, чтобы узнать, что скажет Он во мне, и что мне отвечать по жалобе моей?
HAB|2|2|И отвечал мне Господь и сказал: запиши видение и начертай ясно на скрижалях, чтобы читающий легко мог прочитать,
HAB|2|3|ибо видение относится еще к определенному времени и говорит о конце и не обманет; и хотя бы и замедлило, жди его, ибо непременно сбудется, не отменится.
HAB|2|4|Вот, душа надменная не успокоится, а праведный своею верою жив будет.
HAB|2|5|Надменный человек, как бродящее вино, не успокаивается, так что расширяет душу свою как ад, и как смерть он ненасытен, и собирает к себе все народы, и захватывает себе все племена.
HAB|2|6|Но не все ли они будут произносить о нем притчу и насмешливую песнь: "горе тому, кто без меры обогащает себя не своим, – на долго ли? – и обременяет себя залогами!"
HAB|2|7|Не восстанут ли внезапно те, которые будут терзать тебя, и не поднимутся ли против тебя грабители, и ты достанешься им на расхищение?
HAB|2|8|Так как ты ограбил многие народы, то и тебя ограбят все остальные народы за пролитие крови человеческой, за разорение страны, города и всех живущих в нем.
HAB|2|9|Горе тому, кто жаждет неправедных приобретений для дома своего, чтобы устроить гнездо свое на высоте и тем обезопасить себя от руки несчастья!
HAB|2|10|Бесславие измыслил ты для твоего дома, истребляя многие народы, и согрешил против души твоей.
HAB|2|11|Камни из стен возопиют и перекладины из дерева будут отвечать им:
HAB|2|12|"горе строящему город на крови и созидающему крепости неправдою!"
HAB|2|13|Вот, не от Господа ли Саваофа это, что народы трудятся для огня и племена мучат себя напрасно?
HAB|2|14|Ибо земля наполнится познанием славы Господа, как воды наполняют море.
HAB|2|15|Горе тебе, который подаешь ближнему твоему питье с примесью злобы твоей и делаешь его пьяным, чтобы видеть срамоту его!
HAB|2|16|Ты пресытился стыдом вместо славы; пей же и ты и показывай срамоту, – обратится и к тебе чаша десницы Господней и посрамление на славу твою.
HAB|2|17|Ибо злодейство твое на Ливане обрушится на тебя за истребление устрашенных животных, за пролитие крови человеческой, за опустошение страны, города и всех живущих в нем.
HAB|2|18|Что за польза от истукана, сделанного художником, этого литаго лжеучителя, хотя ваятель, делая немые кумиры, полагается на свое произведение?
HAB|2|19|Горе тому, кто говорит дереву: "встань!" и бессловесному камню: "пробудись!" Научит ли он чему–нибудь? Вот, он обложен золотом и серебром, но дыхания в нем нет.
HAB|2|20|А Господь – во святом храме Своем: да молчит вся земля пред лицем Его!
HAB|3|1|Молитва Аввакума пророка, для пения.
HAB|3|2|Господи! услышал я слух Твой и убоялся. Господи! соверши дело Твое среди лет, среди лет яви его; во гневе вспомни о милости.
HAB|3|3|Бог от Фемана грядет и Святый – от горы Фаран. Покрыло небеса величие Его, и славою Его наполнилась земля.
HAB|3|4|Блеск ее – как солнечный свет; от руки Его лучи, и здесь тайник Его силы!
HAB|3|5|Пред лицем Его идет язва, а по стопам Его – жгучий ветер.
HAB|3|6|Он стал и поколебал землю; воззрел, и в трепет привел народы; вековые горы распались, первобытные холмы опали; пути Его вечные.
HAB|3|7|Грустными видел я шатры Ефиопские; сотряслись палатки земли Мадиамской.
HAB|3|8|Разве на реки воспылал, Господи, гнев Твой? разве на реки – негодование Твое, или на море – ярость Твоя, что Ты восшел на коней Твоих, на колесницы Твои спасительные?
HAB|3|9|Ты обнажил лук Твой по клятвенному обетованию, данному коленам. Ты потоками рассек землю.
HAB|3|10|Увидев Тебя, вострепетали горы, ринулись воды; бездна дала голос свой, высоко подняла руки свои;
HAB|3|11|солнце и луна остановились на месте своем пред светом летающих стрел Твоих, пред сиянием сверкающих копьев Твоих.
HAB|3|12|Во гневе шествуешь Ты по земле и в негодовании попираешь народы.
HAB|3|13|Ты выступаешь для спасения народа Твоего, для спасения помазанного Твоего. Ты сокрушаешь главу нечестивого дома, обнажая его от основания до верха.
HAB|3|14|Ты пронзаешь копьями его главу вождей его, когда они как вихрь ринулись разбить меня, в радости, как бы думая поглотить бедного скрытно.
HAB|3|15|Ты с конями Твоими проложил путь по морю, через пучину великих вод.
HAB|3|16|Я услышал, и вострепетала внутренность моя; при вести о сем задрожали губы мои, боль проникла в кости мои, и колеблется место подо мною; а я должен быть спокоен в день бедствия, когда придет на народ мой грабитель его.
HAB|3|17|Хотя бы не расцвела смоковница и не было плода на виноградных лозах, и маслина изменила, и нива не дала пищи, хотя бы не стало овец в загоне и рогатого скота в стойлах, –
HAB|3|18|но и тогда я буду радоваться о Господе и веселиться о Боге спасения моего.
HAB|3|19|Господь Бог – сила моя: Он сделает ноги мои как у оленя и на высоты мои возведет меня! (Начальнику хора).
