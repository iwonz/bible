PS|1|1|Blessed is the man who does not walk in the counsel of the wicked or stand in the way of sinners or sit in the seat of mockers.
PS|1|2|But his delight is in the law of the LORD, and on his law he meditates day and night.
PS|1|3|He is like a tree planted by streams of water, which yields its fruit in season and whose leaf does not wither. Whatever he does prospers.
PS|1|4|Not so the wicked! They are like chaff that the wind blows away.
PS|1|5|Therefore the wicked will not stand in the judgment, nor sinners in the assembly of the righteous.
PS|1|6|For the LORD watches over the way of the righteous, but the way of the wicked will perish.
PS|2|1|Why do the nations conspire and the peoples plot in vain?
PS|2|2|The kings of the earth take their stand and the rulers gather together against the LORD and against his Anointed One.
PS|2|3|"Let us break their chains," they say, "and throw off their fetters."
PS|2|4|The One enthroned in heaven laughs; the Lord scoffs at them.
PS|2|5|Then he rebukes them in his anger and terrifies them in his wrath, saying,
PS|2|6|"I have installed my King on Zion, my holy hill."
PS|2|7|I will proclaim the decree of the LORD: He said to me, "You are my Son; today I have become your Father.
PS|2|8|Ask of me, and I will make the nations your inheritance, the ends of the earth your possession.
PS|2|9|You will rule them with an iron scepter; you will dash them to pieces like pottery."
PS|2|10|Therefore, you kings, be wise; be warned, you rulers of the earth.
PS|2|11|Serve the LORD with fear and rejoice with trembling.
PS|2|12|Kiss the Son, lest he be angry and you be destroyed in your way, for his wrath can flare up in a moment. Blessed are all who take refuge in him.
PS|3|1|O LORD, how many are my foes! How many rise up against me!
PS|3|2|Many are saying of me, "God will not deliver him." Selah
PS|3|3|But you are a shield around me, O LORD; you bestow glory on me and lift up my head.
PS|3|4|To the LORD I cry aloud, and he answers me from his holy hill. Selah
PS|3|5|I lie down and sleep; I wake again, because the LORD sustains me.
PS|3|6|I will not fear the tens of thousands drawn up against me on every side.
PS|3|7|Arise, O LORD! Deliver me, O my God! Strike all my enemies on the jaw; break the teeth of the wicked.
PS|3|8|From the LORD comes deliverance. May your blessing be on your people. Selah
PS|4|1|Answer me when I call to you, O my righteous God. Give me relief from my distress; be merciful to me and hear my prayer.
PS|4|2|How long, O men, will you turn my glory into shame? How long will you love delusions and seek false gods? Selah
PS|4|3|Know that the LORD has set apart the godly for himself; the LORD will hear when I call to him.
PS|4|4|In your anger do not sin; when you are on your beds, search your hearts and be silent. Selah
PS|4|5|Offer right sacrifices and trust in the LORD.
PS|4|6|Many are asking, "Who can show us any good?" Let the light of your face shine upon us, O LORD.
PS|4|7|You have filled my heart with greater joy than when their grain and new wine abound.
PS|4|8|I will lie down and sleep in peace, for you alone, O LORD, make me dwell in safety.
PS|5|1|Give ear to my words, O LORD, consider my sighing.
PS|5|2|Listen to my cry for help, my King and my God, for to you I pray.
PS|5|3|In the morning, O LORD, you hear my voice; in the morning I lay my requests before you and wait in expectation.
PS|5|4|You are not a God who takes pleasure in evil; with you the wicked cannot dwell.
PS|5|5|The arrogant cannot stand in your presence; you hate all who do wrong.
PS|5|6|You destroy those who tell lies; bloodthirsty and deceitful men the LORD abhors.
PS|5|7|But I, by your great mercy, will come into your house; in reverence will I bow down toward your holy temple.
PS|5|8|Lead me, O LORD, in your righteousness because of my enemies- make straight your way before me.
PS|5|9|Not a word from their mouth can be trusted; their heart is filled with destruction. Their throat is an open grave; with their tongue they speak deceit.
PS|5|10|Declare them guilty, O God! Let their intrigues be their downfall. Banish them for their many sins, for they have rebelled against you.
PS|5|11|But let all who take refuge in you be glad; let them ever sing for joy. Spread your protection over them, that those who love your name may rejoice in you.
PS|5|12|For surely, O LORD, you bless the righteous; you surround them with your favor as with a shield.
PS|6|1|O LORD, do not rebuke me in your anger or discipline me in your wrath.
PS|6|2|Be merciful to me, LORD, for I am faint; O LORD, heal me, for my bones are in agony.
PS|6|3|My soul is in anguish. How long, O LORD, how long?
PS|6|4|Turn, O LORD, and deliver me; save me because of your unfailing love.
PS|6|5|No one remembers you when he is dead. Who praises you from the grave?
PS|6|6|I am worn out from groaning; all night long I flood my bed with weeping and drench my couch with tears.
PS|6|7|My eyes grow weak with sorrow; they fail because of all my foes.
PS|6|8|Away from me, all you who do evil, for the LORD has heard my weeping.
PS|6|9|The LORD has heard my cry for mercy; the LORD accepts my prayer.
PS|6|10|All my enemies will be ashamed and dismayed; they will turn back in sudden disgrace.
PS|7|1|O LORD my God, I take refuge in you; save and deliver me from all who pursue me,
PS|7|2|or they will tear me like a lion and rip me to pieces with no one to rescue me.
PS|7|3|O LORD my God, if I have done this and there is guilt on my hands-
PS|7|4|if I have done evil to him who is at peace with me or without cause have robbed my foe-
PS|7|5|then let my enemy pursue and overtake me; let him trample my life to the ground and make me sleep in the dust. Selah
PS|7|6|Arise, O LORD, in your anger; rise up against the rage of my enemies. Awake, my God; decree justice.
PS|7|7|Let the assembled peoples gather around you. Rule over them from on high;
PS|7|8|let the LORD judge the peoples. Judge me, O LORD, according to my righteousness, according to my integrity, O Most High.
PS|7|9|O righteous God, who searches minds and hearts, bring to an end the violence of the wicked and make the righteous secure.
PS|7|10|My shield is God Most High, who saves the upright in heart.
PS|7|11|God is a righteous judge, a God who expresses his wrath every day.
PS|7|12|If he does not relent, he will sharpen his sword; he will bend and string his bow.
PS|7|13|He has prepared his deadly weapons; he makes ready his flaming arrows.
PS|7|14|He who is pregnant with evil and conceives trouble gives birth to disillusionment.
PS|7|15|He who digs a hole and scoops it out falls into the pit he has made.
PS|7|16|The trouble he causes recoils on himself; his violence comes down on his own head.
PS|7|17|I will give thanks to the LORD because of his righteousness and will sing praise to the name of the LORD Most High.
PS|8|1|O LORD, our Lord, how majestic is your name in all the earth! You have set your glory above the heavens.
PS|8|2|From the lips of children and infants you have ordained praise because of your enemies, to silence the foe and the avenger.
PS|8|3|When I consider your heavens, the work of your fingers, the moon and the stars, which you have set in place,
PS|8|4|what is man that you are mindful of him, the son of man that you care for him?
PS|8|5|You made him a little lower than the heavenly beings and crowned him with glory and honor.
PS|8|6|You made him ruler over the works of your hands; you put everything under his feet:
PS|8|7|all flocks and herds, and the beasts of the field,
PS|8|8|the birds of the air, and the fish of the sea, all that swim the paths of the seas.
PS|8|9|O LORD, our Lord, how majestic is your name in all the earth!
PS|9|1|I will praise you, O LORD, with all my heart; I will tell of all your wonders.
PS|9|2|I will be glad and rejoice in you; I will sing praise to your name, O Most High.
PS|9|3|My enemies turn back; they stumble and perish before you.
PS|9|4|For you have upheld my right and my cause; you have sat on your throne, judging righteously.
PS|9|5|You have rebuked the nations and destroyed the wicked; you have blotted out their name for ever and ever.
PS|9|6|Endless ruin has overtaken the enemy, you have uprooted their cities; even the memory of them has perished.
PS|9|7|The LORD reigns forever; he has established his throne for judgment.
PS|9|8|He will judge the world in righteousness; he will govern the peoples with justice.
PS|9|9|The LORD is a refuge for the oppressed, a stronghold in times of trouble.
PS|9|10|Those who know your name will trust in you, for you, LORD, have never forsaken those who seek you.
PS|9|11|Sing praises to the LORD, enthroned in Zion; proclaim among the nations what he has done.
PS|9|12|For he who avenges blood remembers; he does not ignore the cry of the afflicted.
PS|9|13|O LORD, see how my enemies persecute me! Have mercy and lift me up from the gates of death,
PS|9|14|that I may declare your praises in the gates of the Daughter of Zion and there rejoice in your salvation.
PS|9|15|The nations have fallen into the pit they have dug; their feet are caught in the net they have hidden.
PS|9|16|The LORD is known by his justice; the wicked are ensnared by the work of their hands. Higgaion. Selah
PS|9|17|The wicked return to the grave, all the nations that forget God.
PS|9|18|But the needy will not always be forgotten, nor the hope of the afflicted ever perish.
PS|9|19|Arise, O LORD, let not man triumph; let the nations be judged in your presence.
PS|9|20|Strike them with terror, O LORD; let the nations know they are but men. Selah
PS|10|1|Why, O LORD, do you stand far off? Why do you hide yourself in times of trouble?
PS|10|2|In his arrogance the wicked man hunts down the weak, who are caught in the schemes he devises.
PS|10|3|He boasts of the cravings of his heart; he blesses the greedy and reviles the LORD.
PS|10|4|In his pride the wicked does not seek him; in all his thoughts there is no room for God.
PS|10|5|His ways are always prosperous; he is haughty and your laws are far from him; he sneers at all his enemies.
PS|10|6|He says to himself, "Nothing will shake me; I'll always be happy and never have trouble."
PS|10|7|His mouth is full of curses and lies and threats; trouble and evil are under his tongue.
PS|10|8|He lies in wait near the villages; from ambush he murders the innocent, watching in secret for his victims.
PS|10|9|He lies in wait like a lion in cover; he lies in wait to catch the helpless; he catches the helpless and drags them off in his net.
PS|10|10|His victims are crushed, they collapse; they fall under his strength.
PS|10|11|He says to himself, "God has forgotten; he covers his face and never sees."
PS|10|12|Arise, LORD! Lift up your hand, O God. Do not forget the helpless.
PS|10|13|Why does the wicked man revile God? Why does he say to himself, "He won't call me to account"?
PS|10|14|But you, O God, do see trouble and grief; you consider it to take it in hand. The victim commits himself to you; you are the helper of the fatherless.
PS|10|15|Break the arm of the wicked and evil man; call him to account for his wickedness that would not be found out.
PS|10|16|The LORD is King for ever and ever; the nations will perish from his land.
PS|10|17|You hear, O LORD, the desire of the afflicted; you encourage them, and you listen to their cry,
PS|10|18|defending the fatherless and the oppressed, in order that man, who is of the earth, may terrify no more.
PS|11|1|In the LORD I take refuge. How then can you say to me: "Flee like a bird to your mountain.
PS|11|2|For look, the wicked bend their bows; they set their arrows against the strings to shoot from the shadows at the upright in heart.
PS|11|3|When the foundations are being destroyed, what can the righteous do?"
PS|11|4|The LORD is in his holy temple; the LORD is on his heavenly throne. He observes the sons of men; his eyes examine them.
PS|11|5|The LORD examines the righteous, but the wicked and those who love violence his soul hates.
PS|11|6|On the wicked he will rain fiery coals and burning sulfur; a scorching wind will be their lot.
PS|11|7|For the LORD is righteous, he loves justice; upright men will see his face.
PS|12|1|Help, LORD, for the godly are no more; the faithful have vanished from among men.
PS|12|2|Everyone lies to his neighbor; their flattering lips speak with deception.
PS|12|3|May the LORD cut off all flattering lips and every boastful tongue
PS|12|4|that says, "We will triumph with our tongues; we own our lips -who is our master?"
PS|12|5|"Because of the oppression of the weak and the groaning of the needy, I will now arise," says the LORD. "I will protect them from those who malign them."
PS|12|6|And the words of the LORD are flawless, like silver refined in a furnace of clay, purified seven times.
PS|12|7|O LORD, you will keep us safe and protect us from such people forever.
PS|12|8|The wicked freely strut about when what is vile is honored among men.
PS|13|1|How long, O LORD? Will you forget me forever? How long will you hide your face from me?
PS|13|2|How long must I wrestle with my thoughts and every day have sorrow in my heart? How long will my enemy triumph over me?
PS|13|3|Look on me and answer, O LORD my God. Give light to my eyes, or I will sleep in death;
PS|13|4|my enemy will say, "I have overcome him," and my foes will rejoice when I fall.
PS|13|5|But I trust in your unfailing love; my heart rejoices in your salvation.
PS|13|6|I will sing to the LORD, for he has been good to me.
PS|14|1|The fool says in his heart, "There is no God." They are corrupt, their deeds are vile; there is no one who does good.
PS|14|2|The LORD looks down from heaven on the sons of men to see if there are any who understand, any who seek God.
PS|14|3|All have turned aside, they have together become corrupt; there is no one who does good, not even one.
PS|14|4|Will evildoers never learn- those who devour my people as men eat bread and who do not call on the LORD?
PS|14|5|There they are, overwhelmed with dread, for God is present in the company of the righteous.
PS|14|6|You evildoers frustrate the plans of the poor, but the LORD is their refuge.
PS|14|7|Oh, that salvation for Israel would come out of Zion! When the LORD restores the fortunes of his people, let Jacob rejoice and Israel be glad!
PS|15|1|LORD, who may dwell in your sanctuary? Who may live on your holy hill?
PS|15|2|He whose walk is blameless and who does what is righteous, who speaks the truth from his heart
PS|15|3|and has no slander on his tongue, who does his neighbor no wrong and casts no slur on his fellowman,
PS|15|4|who despises a vile man but honors those who fear the LORD, who keeps his oath even when it hurts,
PS|15|5|who lends his money without usury and does not accept a bribe against the innocent. He who does these things will never be shaken.
PS|16|1|Keep me safe, O God, for in you I take refuge.
PS|16|2|I said to the LORD, "You are my Lord; apart from you I have no good thing."
PS|16|3|As for the saints who are in the land, they are the glorious ones in whom is all my delight.
PS|16|4|The sorrows of those will increase who run after other gods. I will not pour out their libations of blood or take up their names on my lips.
PS|16|5|LORD, you have assigned me my portion and my cup; you have made my lot secure.
PS|16|6|The boundary lines have fallen for me in pleasant places; surely I have a delightful inheritance.
PS|16|7|I will praise the LORD, who counsels me; even at night my heart instructs me.
PS|16|8|I have set the LORD always before me. Because he is at my right hand, I will not be shaken.
PS|16|9|Therefore my heart is glad and my tongue rejoices; my body also will rest secure,
PS|16|10|because you will not abandon me to the grave, nor will you let your Holy One see decay.
PS|16|11|You have made known to me the path of life; you will fill me with joy in your presence, with eternal pleasures at your right hand.
PS|17|1|Hear, O LORD, my righteous plea; listen to my cry. Give ear to my prayer- it does not rise from deceitful lips.
PS|17|2|May my vindication come from you; may your eyes see what is right.
PS|17|3|Though you probe my heart and examine me at night, though you test me, you will find nothing; I have resolved that my mouth will not sin.
PS|17|4|As for the deeds of men- by the word of your lips I have kept myself from the ways of the violent.
PS|17|5|My steps have held to your paths; my feet have not slipped.
PS|17|6|I call on you, O God, for you will answer me; give ear to me and hear my prayer.
PS|17|7|Show the wonder of your great love, you who save by your right hand those who take refuge in you from their foes.
PS|17|8|Keep me as the apple of your eye; hide me in the shadow of your wings
PS|17|9|from the wicked who assail me, from my mortal enemies who surround me.
PS|17|10|They close up their callous hearts, and their mouths speak with arrogance.
PS|17|11|They have tracked me down, they now surround me, with eyes alert, to throw me to the ground.
PS|17|12|They are like a lion hungry for prey, like a great lion crouching in cover.
PS|17|13|Rise up, O LORD, confront them, bring them down; rescue me from the wicked by your sword.
PS|17|14|O LORD, by your hand save me from such men, from men of this world whose reward is in this life. You still the hunger of those you cherish; their sons have plenty, and they store up wealth for their children.
PS|17|15|And I-in righteousness I will see your face; when I awake, I will be satisfied with seeing your likeness.
PS|18|1|I love you, O LORD, my strength.
PS|18|2|The LORD is my rock, my fortress and my deliverer; my God is my rock, in whom I take refuge. He is my shield and the horn of my salvation, my stronghold.
PS|18|3|I call to the LORD, who is worthy of praise, and I am saved from my enemies.
PS|18|4|The cords of death entangled me; the torrents of destruction overwhelmed me.
PS|18|5|The cords of the grave coiled around me; the snares of death confronted me.
PS|18|6|In my distress I called to the LORD; I cried to my God for help. From his temple he heard my voice; my cry came before him, into his ears.
PS|18|7|The earth trembled and quaked, and the foundations of the mountains shook; they trembled because he was angry.
PS|18|8|Smoke rose from his nostrils; consuming fire came from his mouth, burning coals blazed out of it.
PS|18|9|He parted the heavens and came down; dark clouds were under his feet.
PS|18|10|He mounted the cherubim and flew; he soared on the wings of the wind.
PS|18|11|He made darkness his covering, his canopy around him- the dark rain clouds of the sky.
PS|18|12|Out of the brightness of his presence clouds advanced, with hailstones and bolts of lightning.
PS|18|13|The LORD thundered from heaven; the voice of the Most High resounded.
PS|18|14|He shot his arrows and scattered the enemies, great bolts of lightning and routed them.
PS|18|15|The valleys of the sea were exposed and the foundations of the earth laid bare at your rebuke, O LORD, at the blast of breath from your nostrils.
PS|18|16|He reached down from on high and took hold of me; he drew me out of deep waters.
PS|18|17|He rescued me from my powerful enemy, from my foes, who were too strong for me.
PS|18|18|They confronted me in the day of my disaster, but the LORD was my support.
PS|18|19|He brought me out into a spacious place; he rescued me because he delighted in me.
PS|18|20|The LORD has dealt with me according to my righteousness; according to the cleanness of my hands he has rewarded me.
PS|18|21|For I have kept the ways of the LORD; I have not done evil by turning from my God.
PS|18|22|All his laws are before me; I have not turned away from his decrees.
PS|18|23|I have been blameless before him and have kept myself from sin.
PS|18|24|The LORD has rewarded me according to my righteousness, according to the cleanness of my hands in his sight.
PS|18|25|To the faithful you show yourself faithful, to the blameless you show yourself blameless,
PS|18|26|to the pure you show yourself pure, but to the crooked you show yourself shrewd.
PS|18|27|You save the humble but bring low those whose eyes are haughty.
PS|18|28|You, O LORD, keep my lamp burning; my God turns my darkness into light.
PS|18|29|With your help I can advance against a troop; with my God I can scale a wall.
PS|18|30|As for God, his way is perfect; the word of the LORD is flawless. He is a shield for all who take refuge in him.
PS|18|31|For who is God besides the LORD? And who is the Rock except our God?
PS|18|32|It is God who arms me with strength and makes my way perfect.
PS|18|33|He makes my feet like the feet of a deer; he enables me to stand on the heights.
PS|18|34|He trains my hands for battle; my arms can bend a bow of bronze.
PS|18|35|You give me your shield of victory, and your right hand sustains me; you stoop down to make me great.
PS|18|36|You broaden the path beneath me, so that my ankles do not turn.
PS|18|37|I pursued my enemies and overtook them; I did not turn back till they were destroyed.
PS|18|38|I crushed them so that they could not rise; they fell beneath my feet.
PS|18|39|You armed me with strength for battle; you made my adversaries bow at my feet.
PS|18|40|You made my enemies turn their backs in flight, and I destroyed my foes.
PS|18|41|They cried for help, but there was no one to save them- to the LORD, but he did not answer.
PS|18|42|I beat them as fine as dust borne on the wind; I poured them out like mud in the streets.
PS|18|43|You have delivered me from the attacks of the people; you have made me the head of nations; people I did not know are subject to me.
PS|18|44|As soon as they hear me, they obey me; foreigners cringe before me.
PS|18|45|They all lose heart; they come trembling from their strongholds.
PS|18|46|The LORD lives! Praise be to my Rock! Exalted be God my Savior!
PS|18|47|He is the God who avenges me, who subdues nations under me,
PS|18|48|who saves me from my enemies. You exalted me above my foes; from violent men you rescued me.
PS|18|49|Therefore I will praise you among the nations, O LORD; I will sing praises to your name.
PS|18|50|He gives his king great victories; he shows unfailing kindness to his anointed, to David and his descendants forever.
PS|19|1|The heavens declare the glory of God; the skies proclaim the work of his hands.
PS|19|2|Day after day they pour forth speech; night after night they display knowledge.
PS|19|3|There is no speech or language where their voice is not heard.
PS|19|4|Their voice goes out into all the earth, their words to the ends of the world. In the heavens he has pitched a tent for the sun,
PS|19|5|which is like a bridegroom coming forth from his pavilion, like a champion rejoicing to run his course.
PS|19|6|It rises at one end of the heavens and makes its circuit to the other; nothing is hidden from its heat.
PS|19|7|The law of the LORD is perfect, reviving the soul. The statutes of the LORD are trustworthy, making wise the simple.
PS|19|8|The precepts of the LORD are right, giving joy to the heart. The commands of the LORD are radiant, giving light to the eyes.
PS|19|9|The fear of the LORD is pure, enduring forever. The ordinances of the LORD are sure and altogether righteous.
PS|19|10|They are more precious than gold, than much pure gold; they are sweeter than honey, than honey from the comb.
PS|19|11|By them is your servant warned; in keeping them there is great reward.
PS|19|12|Who can discern his errors? Forgive my hidden faults.
PS|19|13|Keep your servant also from willful sins; may they not rule over me. Then will I be blameless, innocent of great transgression.
PS|19|14|May the words of my mouth and the meditation of my heart be pleasing in your sight, O Lord, my Rock and my Redeemer.
PS|20|1|May the LORD answer you when you are in distress; may the name of the God of Jacob protect you.
PS|20|2|May he send you help from the sanctuary and grant you support from Zion.
PS|20|3|May he remember all your sacrifices and accept your burnt offerings. Selah
PS|20|4|May he give you the desire of your heart and make all your plans succeed.
PS|20|5|We will shout for joy when you are victorious and will lift up our banners in the name of our God. May the LORD grant all your requests.
PS|20|6|Now I know that the LORD saves his anointed; he answers him from his holy heaven with the saving power of his right hand.
PS|20|7|Some trust in chariots and some in horses, but we trust in the name of the LORD our God.
PS|20|8|They are brought to their knees and fall, but we rise up and stand firm.
PS|20|9|O LORD, save the king! Answer us when we call!
PS|21|1|O LORD, the king rejoices in your strength. How great is his joy in the victories you give!
PS|21|2|You have granted him the desire of his heart and have not withheld the request of his lips. Selah
PS|21|3|You welcomed him with rich blessings and placed a crown of pure gold on his head.
PS|21|4|He asked you for life, and you gave it to him- length of days, for ever and ever.
PS|21|5|Through the victories you gave, his glory is great; you have bestowed on him splendor and majesty.
PS|21|6|Surely you have granted him eternal blessings and made him glad with the joy of your presence.
PS|21|7|For the king trusts in the LORD; through the unfailing love of the Most High he will not be shaken.
PS|21|8|Your hand will lay hold on all your enemies; your right hand will seize your foes.
PS|21|9|At the time of your appearing you will make them like a fiery furnace. In his wrath the LORD will swallow them up, and his fire will consume them.
PS|21|10|You will destroy their descendants from the earth, their posterity from mankind.
PS|21|11|Though they plot evil against you and devise wicked schemes, they cannot succeed;
PS|21|12|for you will make them turn their backs when you aim at them with drawn bow.
PS|21|13|Be exalted, O LORD, in your strength; we will sing and praise your might.
PS|22|1|My God, my God, why have you forsaken me? Why are you so far from saving me, so far from the words of my groaning?
PS|22|2|O my God, I cry out by day, but you do not answer, by night, and am not silent.
PS|22|3|Yet you are enthroned as the Holy One; you are the praise of Israel.
PS|22|4|In you our fathers put their trust; they trusted and you delivered them.
PS|22|5|They cried to you and were saved; in you they trusted and were not disappointed.
PS|22|6|But I am a worm and not a man, scorned by men and despised by the people.
PS|22|7|All who see me mock me; they hurl insults, shaking their heads:
PS|22|8|"He trusts in the LORD; let the LORD rescue him. Let him deliver him, since he delights in him."
PS|22|9|Yet you brought me out of the womb; you made me trust in you even at my mother's breast.
PS|22|10|From birth I was cast upon you; from my mother's womb you have been my God.
PS|22|11|Do not be far from me, for trouble is near and there is no one to help.
PS|22|12|Many bulls surround me; strong bulls of Bashan encircle me.
PS|22|13|Roaring lions tearing their prey open their mouths wide against me.
PS|22|14|I am poured out like water, and all my bones are out of joint. My heart has turned to wax; it has melted away within me.
PS|22|15|My strength is dried up like a potsherd, and my tongue sticks to the roof of my mouth; you lay me in the dust of death.
PS|22|16|Dogs have surrounded me; a band of evil men has encircled me, they have pierced my hands and my feet.
PS|22|17|I can count all my bones; people stare and gloat over me.
PS|22|18|They divide my garments among them and cast lots for my clothing.
PS|22|19|But you, O LORD, be not far off; O my Strength, come quickly to help me.
PS|22|20|Deliver my life from the sword, my precious life from the power of the dogs.
PS|22|21|Rescue me from the mouth of the lions; save me from the horns of the wild oxen.
PS|22|22|I will declare your name to my brothers; in the congregation I will praise you.
PS|22|23|You who fear the LORD, praise him! All you descendants of Jacob, honor him! Revere him, all you descendants of Israel!
PS|22|24|For he has not despised or disdained the suffering of the afflicted one; he has not hidden his face from him but has listened to his cry for help.
PS|22|25|From you comes the theme of my praise in the great assembly; before those who fear you will I fulfill my vows.
PS|22|26|The poor will eat and be satisfied; they who seek the LORD will praise him- may your hearts live forever!
PS|22|27|All the ends of the earth will remember and turn to the LORD, and all the families of the nations will bow down before him,
PS|22|28|for dominion belongs to the LORD and he rules over the nations.
PS|22|29|All the rich of the earth will feast and worship; all who go down to the dust will kneel before him- those who cannot keep themselves alive.
PS|22|30|Posterity will serve him; future generations will be told about the Lord.
PS|22|31|They will proclaim his righteousness to a people yet unborn- for he has done it.
PS|23|1|The LORD is my shepherd, I shall not be in want.
PS|23|2|He makes me lie down in green pastures, he leads me beside quiet waters,
PS|23|3|he restores my soul. He guides me in paths of righteousness for his name's sake.
PS|23|4|Even though I walk through the valley of the shadow of death, I will fear no evil, for you are with me; your rod and your staff, they comfort me.
PS|23|5|You prepare a table before me in the presence of my enemies. You anoint my head with oil; my cup overflows.
PS|23|6|Surely goodness and love will follow me all the days of my life, and I will dwell in the house of the LORD forever.
PS|24|1|The earth is the LORD's, and everything in it, the world, and all who live in it;
PS|24|2|for he founded it upon the seas and established it upon the waters.
PS|24|3|Who may ascend the hill of the LORD? Who may stand in his holy place?
PS|24|4|He who has clean hands and a pure heart, who does not lift up his soul to an idol or swear by what is false.
PS|24|5|He will receive blessing from the LORD and vindication from God his Savior.
PS|24|6|Such is the generation of those who seek him, who seek your face, O God of Jacob. Selah
PS|24|7|Lift up your heads, O you gates; be lifted up, you ancient doors, that the King of glory may come in.
PS|24|8|Who is this King of glory? The LORD strong and mighty, the LORD mighty in battle.
PS|24|9|Lift up your heads, O you gates; lift them up, you ancient doors, that the King of glory may come in.
PS|24|10|Who is he, this King of glory? The LORD Almighty- he is the King of glory. Selah
PS|25|1|To you, O LORD, I lift up my soul;
PS|25|2|in you I trust, O my God. Do not let me be put to shame, nor let my enemies triumph over me.
PS|25|3|No one whose hope is in you will ever be put to shame, but they will be put to shame who are treacherous without excuse.
PS|25|4|Show me your ways, O LORD, teach me your paths;
PS|25|5|guide me in your truth and teach me, for you are God my Savior, and my hope is in you all day long.
PS|25|6|Remember, O LORD, your great mercy and love, for they are from of old.
PS|25|7|Remember not the sins of my youth and my rebellious ways; according to your love remember me, for you are good, O LORD.
PS|25|8|Good and upright is the LORD; therefore he instructs sinners in his ways.
PS|25|9|He guides the humble in what is right and teaches them his way.
PS|25|10|All the ways of the LORD are loving and faithful for those who keep the demands of his covenant.
PS|25|11|For the sake of your name, O LORD, forgive my iniquity, though it is great.
PS|25|12|Who, then, is the man that fears the LORD? He will instruct him in the way chosen for him.
PS|25|13|He will spend his days in prosperity, and his descendants will inherit the land.
PS|25|14|The LORD confides in those who fear him; he makes his covenant known to them.
PS|25|15|My eyes are ever on the LORD, for only he will release my feet from the snare.
PS|25|16|Turn to me and be gracious to me, for I am lonely and afflicted.
PS|25|17|The troubles of my heart have multiplied; free me from my anguish.
PS|25|18|Look upon my affliction and my distress and take away all my sins.
PS|25|19|See how my enemies have increased and how fiercely they hate me!
PS|25|20|Guard my life and rescue me; let me not be put to shame, for I take refuge in you.
PS|25|21|May integrity and uprightness protect me, because my hope is in you.
PS|25|22|Redeem Israel, O God, from all their troubles!
PS|26|1|Vindicate me, O LORD, for I have led a blameless life; I have trusted in the LORD without wavering.
PS|26|2|Test me, O LORD, and try me, examine my heart and my mind;
PS|26|3|for your love is ever before me, and I walk continually in your truth.
PS|26|4|I do not sit with deceitful men, nor do I consort with hypocrites;
PS|26|5|I abhor the assembly of evildoers and refuse to sit with the wicked.
PS|26|6|I wash my hands in innocence, and go about your altar, O LORD,
PS|26|7|proclaiming aloud your praise and telling of all your wonderful deeds.
PS|26|8|I love the house where you live, O LORD, the place where your glory dwells.
PS|26|9|Do not take away my soul along with sinners, my life with bloodthirsty men,
PS|26|10|in whose hands are wicked schemes, whose right hands are full of bribes.
PS|26|11|But I lead a blameless life; redeem me and be merciful to me.
PS|26|12|My feet stand on level ground; in the great assembly I will praise the LORD.
PS|27|1|The LORD is my light and my salvation- whom shall I fear? The LORD is the stronghold of my life- of whom shall I be afraid?
PS|27|2|When evil men advance against me to devour my flesh, when my enemies and my foes attack me, they will stumble and fall.
PS|27|3|Though an army besiege me, my heart will not fear; though war break out against me, even then will I be confident.
PS|27|4|One thing I ask of the LORD, this is what I seek: that I may dwell in the house of the LORD all the days of my life, to gaze upon the beauty of the LORD and to seek him in his temple.
PS|27|5|For in the day of trouble he will keep me safe in his dwelling; he will hide me in the shelter of his tabernacle and set me high upon a rock.
PS|27|6|Then my head will be exalted above the enemies who surround me; at his tabernacle will I sacrifice with shouts of joy; I will sing and make music to the LORD.
PS|27|7|Hear my voice when I call, O LORD; be merciful to me and answer me.
PS|27|8|My heart says of you, "Seek his face!" Your face, LORD, I will seek.
PS|27|9|Do not hide your face from me, do not turn your servant away in anger; you have been my helper. Do not reject me or forsake me, O God my Savior.
PS|27|10|Though my father and mother forsake me, the LORD will receive me.
PS|27|11|Teach me your way, O LORD; lead me in a straight path because of my oppressors.
PS|27|12|Do not turn me over to the desire of my foes, for false witnesses rise up against me, breathing out violence.
PS|27|13|I am still confident of this: I will see the goodness of the LORD in the land of the living.
PS|27|14|Wait for the LORD; be strong and take heart and wait for the LORD.
PS|28|1|To you I call, O LORD my Rock; do not turn a deaf ear to me. For if you remain silent, I will be like those who have gone down to the pit.
PS|28|2|Hear my cry for mercy as I call to you for help, as I lift up my hands toward your Most Holy Place.
PS|28|3|Do not drag me away with the wicked, with those who do evil, who speak cordially with their neighbors but harbor malice in their hearts.
PS|28|4|Repay them for their deeds and for their evil work; repay them for what their hands have done and bring back upon them what they deserve.
PS|28|5|Since they show no regard for the works of the LORD and what his hands have done, he will tear them down and never build them up again.
PS|28|6|Praise be to the LORD, for he has heard my cry for mercy.
PS|28|7|The LORD is my strength and my shield; my heart trusts in him, and I am helped. My heart leaps for joy and I will give thanks to him in song.
PS|28|8|The LORD is the strength of his people, a fortress of salvation for his anointed one.
PS|28|9|Save your people and bless your inheritance; be their shepherd and carry them forever.
PS|29|1|Ascribe to the LORD, O mighty ones, ascribe to the LORD glory and strength.
PS|29|2|Ascribe to the LORD the glory due his name; worship the LORD in the splendor of his holiness.
PS|29|3|The voice of the LORD is over the waters; the God of glory thunders, the LORD thunders over the mighty waters.
PS|29|4|The voice of the LORD is powerful; the voice of the LORD is majestic.
PS|29|5|The voice of the LORD breaks the cedars; the LORD breaks in pieces the cedars of Lebanon.
PS|29|6|He makes Lebanon skip like a calf, Sirion like a young wild ox.
PS|29|7|The voice of the LORD strikes with flashes of lightning.
PS|29|8|The voice of the LORD shakes the desert; the LORD shakes the Desert of Kadesh.
PS|29|9|The voice of the LORD twists the oaks and strips the forests bare. And in his temple all cry, "Glory!"
PS|29|10|The LORD sits enthroned over the flood; the LORD is enthroned as King forever.
PS|29|11|The LORD gives strength to his people; the LORD blesses his people with peace.
PS|30|1|I will exalt you, O LORD, for you lifted me out of the depths and did not let my enemies gloat over me.
PS|30|2|O LORD my God, I called to you for help and you healed me.
PS|30|3|O LORD, you brought me up from the grave; you spared me from going down into the pit.
PS|30|4|Sing to the LORD, you saints of his; praise his holy name.
PS|30|5|For his anger lasts only a moment, but his favor lasts a lifetime; weeping may remain for a night, but rejoicing comes in the morning.
PS|30|6|When I felt secure, I said, "I will never be shaken."
PS|30|7|O LORD, when you favored me, you made my mountain stand firm; but when you hid your face, I was dismayed.
PS|30|8|To you, O LORD, I called; to the Lord I cried for mercy:
PS|30|9|"What gain is there in my destruction, in my going down into the pit? Will the dust praise you? Will it proclaim your faithfulness?
PS|30|10|Hear, O LORD, and be merciful to me; O LORD, be my help."
PS|30|11|You turned my wailing into dancing; you removed my sackcloth and clothed me with joy,
PS|30|12|that my heart may sing to you and not be silent. O LORD my God, I will give you thanks forever.
PS|31|1|In you, O LORD, I have taken refuge; let me never be put to shame; deliver me in your righteousness.
PS|31|2|Turn your ear to me, come quickly to my rescue; be my rock of refuge, a strong fortress to save me.
PS|31|3|Since you are my rock and my fortress, for the sake of your name lead and guide me.
PS|31|4|Free me from the trap that is set for me, for you are my refuge.
PS|31|5|Into your hands I commit my spirit; redeem me, O LORD, the God of truth.
PS|31|6|I hate those who cling to worthless idols; I trust in the LORD.
PS|31|7|I will be glad and rejoice in your love, for you saw my affliction and knew the anguish of my soul.
PS|31|8|You have not handed me over to the enemy but have set my feet in a spacious place.
PS|31|9|Be merciful to me, O LORD, for I am in distress; my eyes grow weak with sorrow, my soul and my body with grief.
PS|31|10|My life is consumed by anguish and my years by groaning; my strength fails because of my affliction, and my bones grow weak.
PS|31|11|Because of all my enemies, I am the utter contempt of my neighbors; I am a dread to my friends- those who see me on the street flee from me.
PS|31|12|I am forgotten by them as though I were dead; I have become like broken pottery.
PS|31|13|For I hear the slander of many; there is terror on every side; they conspire against me and plot to take my life.
PS|31|14|But I trust in you, O LORD; I say, "You are my God."
PS|31|15|My times are in your hands; deliver me from my enemies and from those who pursue me.
PS|31|16|Let your face shine on your servant; save me in your unfailing love.
PS|31|17|Let me not be put to shame, O LORD, for I have cried out to you; but let the wicked be put to shame and lie silent in the grave.
PS|31|18|Let their lying lips be silenced, for with pride and contempt they speak arrogantly against the righteous.
PS|31|19|How great is your goodness, which you have stored up for those who fear you, which you bestow in the sight of men on those who take refuge in you.
PS|31|20|In the shelter of your presence you hide them from the intrigues of men; in your dwelling you keep them safe from accusing tongues.
PS|31|21|Praise be to the LORD, for he showed his wonderful love to me when I was in a besieged city.
PS|31|22|In my alarm I said, "I am cut off from your sight!" Yet you heard my cry for mercy when I called to you for help.
PS|31|23|Love the LORD, all his saints! The LORD preserves the faithful, but the proud he pays back in full.
PS|31|24|Be strong and take heart, all you who hope in the LORD.
PS|32|1|Blessed is he whose transgressions are forgiven, whose sins are covered.
PS|32|2|Blessed is the man whose sin the LORD does not count against him and in whose spirit is no deceit.
PS|32|3|When I kept silent, my bones wasted away through my groaning all day long.
PS|32|4|For day and night your hand was heavy upon me; my strength was sapped as in the heat of summer. Selah
PS|32|5|Then I acknowledged my sin to you and did not cover up my iniquity. I said, "I will confess my transgressions to the LORD "- and you forgave the guilt of my sin. Selah
PS|32|6|Therefore let everyone who is godly pray to you while you may be found; surely when the mighty waters rise, they will not reach him.
PS|32|7|You are my hiding place; you will protect me from trouble and surround me with songs of deliverance. Selah
PS|32|8|I will instruct you and teach you in the way you should go; I will counsel you and watch over you.
PS|32|9|Do not be like the horse or the mule, which have no understanding but must be controlled by bit and bridle or they will not come to you.
PS|32|10|Many are the woes of the wicked, but the LORD's unfailing love surrounds the man who trusts in him.
PS|32|11|Rejoice in the LORD and be glad, you righteous; sing, all you who are upright in heart!
PS|33|1|Sing joyfully to the LORD, you righteous; it is fitting for the upright to praise him.
PS|33|2|Praise the LORD with the harp; make music to him on the ten-stringed lyre.
PS|33|3|Sing to him a new song; play skillfully, and shout for joy.
PS|33|4|For the word of the LORD is right and true; he is faithful in all he does.
PS|33|5|The LORD loves righteousness and justice; the earth is full of his unfailing love.
PS|33|6|By the word of the LORD were the heavens made, their starry host by the breath of his mouth.
PS|33|7|He gathers the waters of the sea into jars; he puts the deep into storehouses.
PS|33|8|Let all the earth fear the LORD; let all the people of the world revere him.
PS|33|9|For he spoke, and it came to be; he commanded, and it stood firm.
PS|33|10|The LORD foils the plans of the nations; he thwarts the purposes of the peoples.
PS|33|11|But the plans of the LORD stand firm forever, the purposes of his heart through all generations.
PS|33|12|Blessed is the nation whose God is the LORD, the people he chose for his inheritance.
PS|33|13|From heaven the LORD looks down and sees all mankind;
PS|33|14|from his dwelling place he watches all who live on earth-
PS|33|15|he who forms the hearts of all, who considers everything they do.
PS|33|16|No king is saved by the size of his army; no warrior escapes by his great strength.
PS|33|17|A horse is a vain hope for deliverance; despite all its great strength it cannot save.
PS|33|18|But the eyes of the LORD are on those who fear him, on those whose hope is in his unfailing love,
PS|33|19|to deliver them from death and keep them alive in famine.
PS|33|20|We wait in hope for the LORD; he is our help and our shield.
PS|33|21|In him our hearts rejoice, for we trust in his holy name.
PS|33|22|May your unfailing love rest upon us, O LORD, even as we put our hope in you.
PS|34|1|I will extol the LORD at all times; his praise will always be on my lips.
PS|34|2|My soul will boast in the LORD; let the afflicted hear and rejoice.
PS|34|3|Glorify the LORD with me; let us exalt his name together.
PS|34|4|I sought the LORD, and he answered me; he delivered me from all my fears.
PS|34|5|Those who look to him are radiant; their faces are never covered with shame.
PS|34|6|This poor man called, and the LORD heard him; he saved him out of all his troubles.
PS|34|7|The angel of the LORD encamps around those who fear him, and he delivers them.
PS|34|8|Taste and see that the LORD is good; blessed is the man who takes refuge in him.
PS|34|9|Fear the LORD, you his saints, for those who fear him lack nothing.
PS|34|10|The lions may grow weak and hungry, but those who seek the LORD lack no good thing.
PS|34|11|Come, my children, listen to me; I will teach you the fear of the LORD.
PS|34|12|Whoever of you loves life and desires to see many good days,
PS|34|13|keep your tongue from evil and your lips from speaking lies.
PS|34|14|Turn from evil and do good; seek peace and pursue it.
PS|34|15|The eyes of the LORD are on the righteous and his ears are attentive to their cry;
PS|34|16|the face of the LORD is against those who do evil, to cut off the memory of them from the earth.
PS|34|17|The righteous cry out, and the LORD hears them; he delivers them from all their troubles.
PS|34|18|The LORD is close to the brokenhearted and saves those who are crushed in spirit.
PS|34|19|A righteous man may have many troubles, but the LORD delivers him from them all;
PS|34|20|he protects all his bones, not one of them will be broken.
PS|34|21|Evil will slay the wicked; the foes of the righteous will be condemned.
PS|34|22|The LORD redeems his servants; no one will be condemned who takes refuge in him.
PS|35|1|Contend, O LORD, with those who contend with me; fight against those who fight against me.
PS|35|2|Take up shield and buckler; arise and come to my aid.
PS|35|3|Brandish spear and javelin against those who pursue me. Say to my soul, "I am your salvation."
PS|35|4|May those who seek my life be disgraced and put to shame; may those who plot my ruin be turned back in dismay.
PS|35|5|May they be like chaff before the wind, with the angel of the LORD driving them away;
PS|35|6|may their path be dark and slippery, with the angel of the LORD pursuing them.
PS|35|7|Since they hid their net for me without cause and without cause dug a pit for me,
PS|35|8|may ruin overtake them by surprise- may the net they hid entangle them, may they fall into the pit, to their ruin.
PS|35|9|Then my soul will rejoice in the LORD and delight in his salvation.
PS|35|10|My whole being will exclaim, "Who is like you, O LORD? You rescue the poor from those too strong for them, the poor and needy from those who rob them."
PS|35|11|Ruthless witnesses come forward; they question me on things I know nothing about.
PS|35|12|They repay me evil for good and leave my soul forlorn.
PS|35|13|Yet when they were ill, I put on sackcloth and humbled myself with fasting. When my prayers returned to me unanswered,
PS|35|14|I went about mourning as though for my friend or brother. I bowed my head in grief as though weeping for my mother.
PS|35|15|But when I stumbled, they gathered in glee; attackers gathered against me when I was unaware. They slandered me without ceasing.
PS|35|16|Like the ungodly they maliciously mocked; they gnashed their teeth at me.
PS|35|17|O Lord, how long will you look on? Rescue my life from their ravages, my precious life from these lions.
PS|35|18|I will give you thanks in the great assembly; among throngs of people I will praise you.
PS|35|19|Let not those gloat over me who are my enemies without cause; let not those who hate me without reason maliciously wink the eye.
PS|35|20|They do not speak peaceably, but devise false accusations against those who live quietly in the land.
PS|35|21|They gape at me and say, "Aha! Aha! With our own eyes we have seen it."
PS|35|22|O LORD, you have seen this; be not silent. Do not be far from me, O Lord.
PS|35|23|Awake, and rise to my defense! Contend for me, my God and Lord.
PS|35|24|Vindicate me in your righteousness, O LORD my God; do not let them gloat over me.
PS|35|25|Do not let them think, "Aha, just what we wanted!" or say, "We have swallowed him up."
PS|35|26|May all who gloat over my distress be put to shame and confusion; may all who exalt themselves over me be clothed with shame and disgrace.
PS|35|27|May those who delight in my vindication shout for joy and gladness; may they always say, "The LORD be exalted, who delights in the well-being of his servant."
PS|35|28|My tongue will speak of your righteousness and of your praises all day long.
PS|36|1|An oracle is within my heart concerning the sinfulness of the wicked: There is no fear of God before his eyes.
PS|36|2|For in his own eyes he flatters himself too much to detect or hate his sin.
PS|36|3|The words of his mouth are wicked and deceitful; he has ceased to be wise and to do good.
PS|36|4|Even on his bed he plots evil; he commits himself to a sinful course and does not reject what is wrong.
PS|36|5|Your love, O LORD, reaches to the heavens, your faithfulness to the skies.
PS|36|6|Your righteousness is like the mighty mountains, your justice like the great deep. O LORD, you preserve both man and beast.
PS|36|7|How priceless is your unfailing love! Both high and low among men find refuge in the shadow of your wings.
PS|36|8|They feast on the abundance of your house; you give them drink from your river of delights.
PS|36|9|For with you is the fountain of life; in your light we see light.
PS|36|10|Continue your love to those who know you, your righteousness to the upright in heart.
PS|36|11|May the foot of the proud not come against me, nor the hand of the wicked drive me away.
PS|36|12|See how the evildoers lie fallen- thrown down, not able to rise!
PS|37|1|Do not fret because of evil men or be envious of those who do wrong;
PS|37|2|for like the grass they will soon wither, like green plants they will soon die away.
PS|37|3|Trust in the LORD and do good; dwell in the land and enjoy safe pasture.
PS|37|4|Delight yourself in the LORD and he will give you the desires of your heart.
PS|37|5|Commit your way to the LORD; trust in him and he will do this:
PS|37|6|He will make your righteousness shine like the dawn, the justice of your cause like the noonday sun.
PS|37|7|Be still before the LORD and wait patiently for him; do not fret when men succeed in their ways, when they carry out their wicked schemes.
PS|37|8|Refrain from anger and turn from wrath; do not fret-it leads only to evil.
PS|37|9|For evil men will be cut off, but those who hope in the LORD will inherit the land.
PS|37|10|A little while, and the wicked will be no more; though you look for them, they will not be found.
PS|37|11|But the meek will inherit the land and enjoy great peace.
PS|37|12|The wicked plot against the righteous and gnash their teeth at them;
PS|37|13|but the Lord laughs at the wicked, for he knows their day is coming.
PS|37|14|The wicked draw the sword and bend the bow to bring down the poor and needy, to slay those whose ways are upright.
PS|37|15|But their swords will pierce their own hearts, and their bows will be broken.
PS|37|16|Better the little that the righteous have than the wealth of many wicked;
PS|37|17|for the power of the wicked will be broken, but the LORD upholds the righteous.
PS|37|18|The days of the blameless are known to the LORD, and their inheritance will endure forever.
PS|37|19|In times of disaster they will not wither; in days of famine they will enjoy plenty.
PS|37|20|But the wicked will perish: The LORD's enemies will be like the beauty of the fields, they will vanish-vanish like smoke.
PS|37|21|The wicked borrow and do not repay, but the righteous give generously;
PS|37|22|those the LORD blesses will inherit the land, but those he curses will be cut off.
PS|37|23|If the LORD delights in a man's way, he makes his steps firm;
PS|37|24|though he stumble, he will not fall, for the LORD upholds him with his hand.
PS|37|25|I was young and now I am old, yet I have never seen the righteous forsaken or their children begging bread.
PS|37|26|They are always generous and lend freely; their children will be blessed.
PS|37|27|Turn from evil and do good; then you will dwell in the land forever.
PS|37|28|For the LORD loves the just and will not forsake his faithful ones. They will be protected forever, but the offspring of the wicked will be cut off;
PS|37|29|the righteous will inherit the land and dwell in it forever.
PS|37|30|The mouth of the righteous man utters wisdom, and his tongue speaks what is just.
PS|37|31|The law of his God is in his heart; his feet do not slip.
PS|37|32|The wicked lie in wait for the righteous, seeking their very lives;
PS|37|33|but the LORD will not leave them in their power or let them be condemned when brought to trial.
PS|37|34|Wait for the LORD and keep his way. He will exalt you to inherit the land; when the wicked are cut off, you will see it.
PS|37|35|I have seen a wicked and ruthless man flourishing like a green tree in its native soil,
PS|37|36|but he soon passed away and was no more; though I looked for him, he could not be found.
PS|37|37|Consider the blameless, observe the upright; there is a future for the man of peace.
PS|37|38|But all sinners will be destroyed; the future of the wicked will be cut off.
PS|37|39|The salvation of the righteous comes from the LORD; he is their stronghold in time of trouble.
PS|37|40|The LORD helps them and delivers them; he delivers them from the wicked and saves them, because they take refuge in him.
PS|38|1|O LORD, do not rebuke me in your anger or discipline me in your wrath.
PS|38|2|For your arrows have pierced me, and your hand has come down upon me.
PS|38|3|Because of your wrath there is no health in my body; my bones have no soundness because of my sin.
PS|38|4|My guilt has overwhelmed me like a burden too heavy to bear.
PS|38|5|My wounds fester and are loathsome because of my sinful folly.
PS|38|6|I am bowed down and brought very low; all day long I go about mourning.
PS|38|7|My back is filled with searing pain; there is no health in my body.
PS|38|8|I am feeble and utterly crushed; I groan in anguish of heart.
PS|38|9|All my longings lie open before you, O Lord; my sighing is not hidden from you.
PS|38|10|My heart pounds, my strength fails me; even the light has gone from my eyes.
PS|38|11|My friends and companions avoid me because of my wounds; my neighbors stay far away.
PS|38|12|Those who seek my life set their traps, those who would harm me talk of my ruin; all day long they plot deception.
PS|38|13|I am like a deaf man, who cannot hear, like a mute, who cannot open his mouth;
PS|38|14|I have become like a man who does not hear, whose mouth can offer no reply.
PS|38|15|I wait for you, O LORD; you will answer, O Lord my God.
PS|38|16|For I said, "Do not let them gloat or exalt themselves over me when my foot slips."
PS|38|17|For I am about to fall, and my pain is ever with me.
PS|38|18|I confess my iniquity; I am troubled by my sin.
PS|38|19|Many are those who are my vigorous enemies; those who hate me without reason are numerous.
PS|38|20|Those who repay my good with evil slander me when I pursue what is good.
PS|38|21|O LORD, do not forsake me; be not far from me, O my God.
PS|38|22|Come quickly to help me, O Lord my Savior.
PS|39|1|I said, "I will watch my ways and keep my tongue from sin; I will put a muzzle on my mouth as long as the wicked are in my presence."
PS|39|2|But when I was silent and still, not even saying anything good, my anguish increased.
PS|39|3|My heart grew hot within me, and as I meditated, the fire burned; then I spoke with my tongue:
PS|39|4|"Show me, O LORD, my life's end and the number of my days; let me know how fleeting is my life.
PS|39|5|You have made my days a mere handbreadth; the span of my years is as nothing before you. Each man's life is but a breath. Selah
PS|39|6|Man is a mere phantom as he goes to and fro: He bustles about, but only in vain; he heaps up wealth, not knowing who will get it.
PS|39|7|"But now, Lord, what do I look for? My hope is in you.
PS|39|8|Save me from all my transgressions; do not make me the scorn of fools.
PS|39|9|I was silent; I would not open my mouth, for you are the one who has done this.
PS|39|10|Remove your scourge from me; I am overcome by the blow of your hand.
PS|39|11|You rebuke and discipline men for their sin; you consume their wealth like a moth- each man is but a breath. Selah
PS|39|12|"Hear my prayer, O LORD, listen to my cry for help; be not deaf to my weeping. For I dwell with you as an alien, a stranger, as all my fathers were.
PS|39|13|Look away from me, that I may rejoice again before I depart and am no more."
PS|40|1|I waited patiently for the LORD; he turned to me and heard my cry.
PS|40|2|He lifted me out of the slimy pit, out of the mud and mire; he set my feet on a rock and gave me a firm place to stand.
PS|40|3|He put a new song in my mouth, a hymn of praise to our God. Many will see and fear and put their trust in the LORD.
PS|40|4|Blessed is the man who makes the LORD his trust, who does not look to the proud, to those who turn aside to false gods.
PS|40|5|Many, O LORD my God, are the wonders you have done. The things you planned for us no one can recount to you; were I to speak and tell of them, they would be too many to declare.
PS|40|6|Sacrifice and offering you did not desire, but my ears you have pierced,; burnt offerings and sin offerings you did not require.
PS|40|7|Then I said, "Here I am, I have come- it is written about me in the scroll.
PS|40|8|I desire to do your will, O my God; your law is within my heart."
PS|40|9|I proclaim righteousness in the great assembly; I do not seal my lips, as you know, O LORD.
PS|40|10|I do not hide your righteousness in my heart; I speak of your faithfulness and salvation. I do not conceal your love and your truth from the great assembly.
PS|40|11|Do not withhold your mercy from me, O LORD; may your love and your truth always protect me.
PS|40|12|For troubles without number surround me; my sins have overtaken me, and I cannot see. They are more than the hairs of my head, and my heart fails within me.
PS|40|13|Be pleased, O LORD, to save me; O LORD, come quickly to help me.
PS|40|14|May all who seek to take my life be put to shame and confusion; may all who desire my ruin be turned back in disgrace.
PS|40|15|May those who say to me, "Aha! Aha!" be appalled at their own shame.
PS|40|16|But may all who seek you rejoice and be glad in you; may those who love your salvation always say, "The LORD be exalted!"
PS|40|17|Yet I am poor and needy; may the Lord think of me. You are my help and my deliverer; O my God, do not delay.
PS|41|1|Blessed is he who has regard for the weak; the LORD delivers him in times of trouble.
PS|41|2|The LORD will protect him and preserve his life; he will bless him in the land and not surrender him to the desire of his foes.
PS|41|3|The LORD will sustain him on his sickbed and restore him from his bed of illness.
PS|41|4|I said, "O LORD, have mercy on me; heal me, for I have sinned against you."
PS|41|5|My enemies say of me in malice, "When will he die and his name perish?"
PS|41|6|Whenever one comes to see me, he speaks falsely, while his heart gathers slander; then he goes out and spreads it abroad.
PS|41|7|All my enemies whisper together against me; they imagine the worst for me, saying,
PS|41|8|"A vile disease has beset him; he will never get up from the place where he lies."
PS|41|9|Even my close friend, whom I trusted, he who shared my bread, has lifted up his heel against me.
PS|41|10|But you, O LORD, have mercy on me; raise me up, that I may repay them.
PS|41|11|I know that you are pleased with me, for my enemy does not triumph over me.
PS|41|12|In my integrity you uphold me and set me in your presence forever.
PS|41|13|Praise be to the LORD, the God of Israel, from everlasting to everlasting. Amen and Amen.
PS|42|1|As the deer pants for streams of water, so my soul pants for you, O God.
PS|42|2|My soul thirsts for God, for the living God. When can I go and meet with God?
PS|42|3|My tears have been my food day and night, while men say to me all day long, "Where is your God?"
PS|42|4|These things I remember as I pour out my soul: how I used to go with the multitude, leading the procession to the house of God, with shouts of joy and thanksgiving among the festive throng.
PS|42|5|Why are you downcast, O my soul? Why so disturbed within me? Put your hope in God, for I will yet praise him, my Savior and
PS|42|6|my God. My soul is downcast within me; therefore I will remember you from the land of the Jordan, the heights of Hermon-from Mount Mizar.
PS|42|7|Deep calls to deep in the roar of your waterfalls; all your waves and breakers have swept over me.
PS|42|8|By day the LORD directs his love, at night his song is with me- a prayer to the God of my life.
PS|42|9|I say to God my Rock, "Why have you forgotten me? Why must I go about mourning, oppressed by the enemy?"
PS|42|10|My bones suffer mortal agony as my foes taunt me, saying to me all day long, "Where is your God?"
PS|42|11|Why are you downcast, O my soul? Why so disturbed within me? Put your hope in God, for I will yet praise him, my Savior and my God.
PS|43|1|Vindicate me, O God, and plead my cause against an ungodly nation; rescue me from deceitful and wicked men.
PS|43|2|You are God my stronghold. Why have you rejected me? Why must I go about mourning, oppressed by the enemy?
PS|43|3|Send forth your light and your truth, let them guide me; let them bring me to your holy mountain, to the place where you dwell.
PS|43|4|Then will I go to the altar of God, to God, my joy and my delight. I will praise you with the harp, O God, my God.
PS|43|5|Why are you downcast, O my soul? Why so disturbed within me? Put your hope in God, for I will yet praise him, my Savior and my God.
PS|44|1|We have heard with our ears, O God; our fathers have told us what you did in their days, in days long ago.
PS|44|2|With your hand you drove out the nations and planted our fathers; you crushed the peoples and made our fathers flourish.
PS|44|3|It was not by their sword that they won the land, nor did their arm bring them victory; it was your right hand, your arm, and the light of your face, for you loved them.
PS|44|4|You are my King and my God, who decrees victories for Jacob.
PS|44|5|Through you we push back our enemies; through your name we trample our foes.
PS|44|6|I do not trust in my bow, my sword does not bring me victory;
PS|44|7|but you give us victory over our enemies, you put our adversaries to shame.
PS|44|8|In God we make our boast all day long, and we will praise your name forever. Selah
PS|44|9|But now you have rejected and humbled us; you no longer go out with our armies.
PS|44|10|You made us retreat before the enemy, and our adversaries have plundered us.
PS|44|11|You gave us up to be devoured like sheep and have scattered us among the nations.
PS|44|12|You sold your people for a pittance, gaining nothing from their sale.
PS|44|13|You have made us a reproach to our neighbors, the scorn and derision of those around us.
PS|44|14|You have made us a byword among the nations; the peoples shake their heads at us.
PS|44|15|My disgrace is before me all day long, and my face is covered with shame
PS|44|16|at the taunts of those who reproach and revile me, because of the enemy, who is bent on revenge.
PS|44|17|All this happened to us, though we had not forgotten you or been false to your covenant.
PS|44|18|Our hearts had not turned back; our feet had not strayed from your path.
PS|44|19|But you crushed us and made us a haunt for jackals and covered us over with deep darkness.
PS|44|20|If we had forgotten the name of our God or spread out our hands to a foreign god,
PS|44|21|would not God have discovered it, since he knows the secrets of the heart?
PS|44|22|Yet for your sake we face death all day long; we are considered as sheep to be slaughtered.
PS|44|23|Awake, O Lord! Why do you sleep? Rouse yourself! Do not reject us forever.
PS|44|24|Why do you hide your face and forget our misery and oppression?
PS|44|25|We are brought down to the dust; our bodies cling to the ground.
PS|44|26|Rise up and help us; redeem us because of your unfailing love.
PS|45|1|My heart is stirred by a noble theme as I recite my verses for the king; my tongue is the pen of a skillful writer.
PS|45|2|You are the most excellent of men and your lips have been anointed with grace, since God has blessed you forever.
PS|45|3|Gird your sword upon your side, O mighty one; clothe yourself with splendor and majesty.
PS|45|4|In your majesty ride forth victoriously in behalf of truth, humility and righteousness; let your right hand display awesome deeds.
PS|45|5|Let your sharp arrows pierce the hearts of the king's enemies; let the nations fall beneath your feet.
PS|45|6|Your throne, O God, will last for ever and ever; a scepter of justice will be the scepter of your kingdom.
PS|45|7|You love righteousness and hate wickedness; therefore God, your God, has set you above your companions by anointing you with the oil of joy.
PS|45|8|All your robes are fragrant with myrrh and aloes and cassia; from palaces adorned with ivory the music of the strings makes you glad.
PS|45|9|Daughters of kings are among your honored women; at your right hand is the royal bride in gold of Ophir.
PS|45|10|Listen, O daughter, consider and give ear: Forget your people and your father's house.
PS|45|11|The king is enthralled by your beauty; honor him, for he is your lord.
PS|45|12|The Daughter of Tyre will come with a gift, men of wealth will seek your favor.
PS|45|13|All glorious is the princess within her chamber; her gown is interwoven with gold.
PS|45|14|In embroidered garments she is led to the king; her virgin companions follow her and are brought to you.
PS|45|15|They are led in with joy and gladness; they enter the palace of the king.
PS|45|16|Your sons will take the place of your fathers; you will make them princes throughout the land.
PS|45|17|I will perpetuate your memory through all generations; therefore the nations will praise you for ever and ever.
PS|46|1|God is our refuge and strength, an ever-present help in trouble.
PS|46|2|Therefore we will not fear, though the earth give way and the mountains fall into the heart of the sea,
PS|46|3|though its waters roar and foam and the mountains quake with their surging. Selah
PS|46|4|There is a river whose streams make glad the city of God, the holy place where the Most High dwells.
PS|46|5|God is within her, she will not fall; God will help her at break of day.
PS|46|6|Nations are in uproar, kingdoms fall; he lifts his voice, the earth melts.
PS|46|7|The LORD Almighty is with us; the God of Jacob is our fortress. Selah
PS|46|8|Come and see the works of the LORD, the desolations he has brought on the earth.
PS|46|9|He makes wars cease to the ends of the earth; he breaks the bow and shatters the spear, he burns the shields with fire.
PS|46|10|"Be still, and know that I am God; I will be exalted among the nations, I will be exalted in the earth."
PS|46|11|The LORD Almighty is with us; the God of Jacob is our fortress. Selah
PS|47|1|Clap your hands, all you nations; shout to God with cries of joy.
PS|47|2|How awesome is the LORD Most High, the great King over all the earth!
PS|47|3|He subdued nations under us, peoples under our feet.
PS|47|4|He chose our inheritance for us, the pride of Jacob, whom he loved. Selah
PS|47|5|God has ascended amid shouts of joy, the LORD amid the sounding of trumpets.
PS|47|6|Sing praises to God, sing praises; sing praises to our King, sing praises.
PS|47|7|For God is the King of all the earth; sing to him a psalm of praise.
PS|47|8|God reigns over the nations; God is seated on his holy throne.
PS|47|9|The nobles of the nations assemble as the people of the God of Abraham, for the kings of the earth belong to God; he is greatly exalted.
PS|48|1|Great is the LORD, and most worthy of praise, in the city of our God, his holy mountain.
PS|48|2|It is beautiful in its loftiness, the joy of the whole earth. Like the utmost heights of Zaphon is Mount Zion, the city of the Great King.
PS|48|3|God is in her citadels; he has shown himself to be her fortress.
PS|48|4|When the kings joined forces, when they advanced together,
PS|48|5|they saw her and were astounded; they fled in terror.
PS|48|6|Trembling seized them there, pain like that of a woman in labor.
PS|48|7|You destroyed them like ships of Tarshish shattered by an east wind.
PS|48|8|As we have heard, so have we seen in the city of the LORD Almighty, in the city of our God: God makes her secure forever. Selah
PS|48|9|Within your temple, O God, we meditate on your unfailing love.
PS|48|10|Like your name, O God, your praise reaches to the ends of the earth; your right hand is filled with righteousness.
PS|48|11|Mount Zion rejoices, the villages of Judah are glad because of your judgments.
PS|48|12|Walk about Zion, go around her, count her towers,
PS|48|13|consider well her ramparts, view her citadels, that you may tell of them to the next generation.
PS|48|14|For this God is our God for ever and ever; he will be our guide even to the end.
PS|49|1|Hear this, all you peoples; listen, all who live in this world,
PS|49|2|both low and high, rich and poor alike:
PS|49|3|My mouth will speak words of wisdom; the utterance from my heart will give understanding.
PS|49|4|I will turn my ear to a proverb; with the harp I will expound my riddle:
PS|49|5|Why should I fear when evil days come, when wicked deceivers surround me-
PS|49|6|those who trust in their wealth and boast of their great riches?
PS|49|7|No man can redeem the life of another or give to God a ransom for him-
PS|49|8|the ransom for a life is costly, no payment is ever enough-
PS|49|9|that he should live on forever and not see decay.
PS|49|10|For all can see that wise men die; the foolish and the senseless alike perish and leave their wealth to others.
PS|49|11|Their tombs will remain their houses forever, their dwellings for endless generations, though they had named lands after themselves.
PS|49|12|But man, despite his riches, does not endure; he is like the beasts that perish.
PS|49|13|This is the fate of those who trust in themselves, and of their followers, who approve their sayings. Selah
PS|49|14|Like sheep they are destined for the grave, and death will feed on them. The upright will rule over them in the morning; their forms will decay in the grave, far from their princely mansions.
PS|49|15|But God will redeem my life from the grave; he will surely take me to himself. Selah
PS|49|16|Do not be overawed when a man grows rich, when the splendor of his house increases;
PS|49|17|for he will take nothing with him when he dies, his splendor will not descend with him.
PS|49|18|Though while he lived he counted himself blessed- and men praise you when you prosper-
PS|49|19|he will join the generation of his fathers, who will never see the light of life.
PS|49|20|A man who has riches without understanding is like the beasts that perish.
PS|50|1|The Mighty One, God, the LORD, speaks and summons the earth from the rising of the sun to the place where it sets.
PS|50|2|From Zion, perfect in beauty, God shines forth.
PS|50|3|Our God comes and will not be silent; a fire devours before him, and around him a tempest rages.
PS|50|4|He summons the heavens above, and the earth, that he may judge his people:
PS|50|5|"Gather to me my consecrated ones, who made a covenant with me by sacrifice."
PS|50|6|And the heavens proclaim his righteousness, for God himself is judge. Selah
PS|50|7|"Hear, O my people, and I will speak, O Israel, and I will testify against you: I am God, your God.
PS|50|8|I do not rebuke you for your sacrifices or your burnt offerings, which are ever before me.
PS|50|9|I have no need of a bull from your stall or of goats from your pens,
PS|50|10|for every animal of the forest is mine, and the cattle on a thousand hills.
PS|50|11|I know every bird in the mountains, and the creatures of the field are mine.
PS|50|12|If I were hungry I would not tell you, for the world is mine, and all that is in it.
PS|50|13|Do I eat the flesh of bulls or drink the blood of goats?
PS|50|14|Sacrifice thank offerings to God, fulfill your vows to the Most High,
PS|50|15|and call upon me in the day of trouble; I will deliver you, and you will honor me."
PS|50|16|But to the wicked, God says: "What right have you to recite my laws or take my covenant on your lips?
PS|50|17|You hate my instruction and cast my words behind you.
PS|50|18|When you see a thief, you join with him; you throw in your lot with adulterers.
PS|50|19|You use your mouth for evil and harness your tongue to deceit.
PS|50|20|You speak continually against your brother and slander your own mother's son.
PS|50|21|These things you have done and I kept silent; you thought I was altogether like you. But I will rebuke you and accuse you to your face.
PS|50|22|"Consider this, you who forget God, or I will tear you to pieces, with none to rescue:
PS|50|23|He who sacrifices thank offerings honors me, and he prepares the way so that I may show him the salvation of God."
PS|51|1|Have mercy on me, O God, according to your unfailing love; according to your great compassion blot out my transgressions.
PS|51|2|Wash away all my iniquity and cleanse me from my sin.
PS|51|3|For I know my transgressions, and my sin is always before me.
PS|51|4|Against you, you only, have I sinned and done what is evil in your sight, so that you are proved right when you speak and justified when you judge.
PS|51|5|Surely I was sinful at birth, sinful from the time my mother conceived me.
PS|51|6|Surely you desire truth in the inner parts; you teach me wisdom in the inmost place.
PS|51|7|Cleanse me with hyssop, and I will be clean; wash me, and I will be whiter than snow.
PS|51|8|Let me hear joy and gladness; let the bones you have crushed rejoice.
PS|51|9|Hide your face from my sins and blot out all my iniquity.
PS|51|10|Create in me a pure heart, O God, and renew a steadfast spirit within me.
PS|51|11|Do not cast me from your presence or take your Holy Spirit from me.
PS|51|12|Restore to me the joy of your salvation and grant me a willing spirit, to sustain me.
PS|51|13|Then I will teach transgressors your ways, and sinners will turn back to you.
PS|51|14|Save me from bloodguilt, O God, the God who saves me, and my tongue will sing of your righteousness.
PS|51|15|O Lord, open my lips, and my mouth will declare your praise.
PS|51|16|You do not delight in sacrifice, or I would bring it; you do not take pleasure in burnt offerings.
PS|51|17|The sacrifices of God are a broken spirit; a broken and contrite heart, O God, you will not despise.
PS|51|18|In your good pleasure make Zion prosper; build up the walls of Jerusalem.
PS|51|19|Then there will be righteous sacrifices, whole burnt offerings to delight you; then bulls will be offered on your altar.
PS|52|1|Why do you boast of evil, you mighty man? Why do you boast all day long, you who are a disgrace in the eyes of God?
PS|52|2|Your tongue plots destruction; it is like a sharpened razor, you who practice deceit.
PS|52|3|You love evil rather than good, falsehood rather than speaking the truth. Selah
PS|52|4|You love every harmful word, O you deceitful tongue!
PS|52|5|Surely God will bring you down to everlasting ruin: He will snatch you up and tear you from your tent; he will uproot you from the land of the living. Selah
PS|52|6|The righteous will see and fear; they will laugh at him, saying,
PS|52|7|"Here now is the man who did not make God his stronghold but trusted in his great wealth and grew strong by destroying others!"
PS|52|8|But I am like an olive tree flourishing in the house of God; I trust in God's unfailing love for ever and ever.
PS|52|9|I will praise you forever for what you have done; in your name I will hope, for your name is good. I will praise you in the presence of your saints.
PS|53|1|The fool says in his heart, "There is no God." They are corrupt, and their ways are vile; there is no one who does good.
PS|53|2|God looks down from heaven on the sons of men to see if there are any who understand, any who seek God.
PS|53|3|Everyone has turned away, they have together become corrupt; there is no one who does good, not even one.
PS|53|4|Will the evildoers never learn- those who devour my people as men eat bread and who do not call on God?
PS|53|5|There they were, overwhelmed with dread, where there was nothing to dread. God scattered the bones of those who attacked you; you put them to shame, for God despised them.
PS|53|6|Oh, that salvation for Israel would come out of Zion! When God restores the fortunes of his people, let Jacob rejoice and Israel be glad!
PS|54|1|Save me, O God, by your name; vindicate me by your might.
PS|54|2|Hear my prayer, O God; listen to the words of my mouth.
PS|54|3|Strangers are attacking me; ruthless men seek my life- men without regard for God. Selah
PS|54|4|Surely God is my help; the Lord is the one who sustains me.
PS|54|5|Let evil recoil on those who slander me; in your faithfulness destroy them.
PS|54|6|I will sacrifice a freewill offering to you; I will praise your name, O LORD, for it is good.
PS|54|7|For he has delivered me from all my troubles, and my eyes have looked in triumph on my foes.
PS|55|1|Listen to my prayer, O God, do not ignore my plea;
PS|55|2|hear me and answer me. My thoughts trouble me and I am distraught
PS|55|3|at the voice of the enemy, at the stares of the wicked; for they bring down suffering upon me and revile me in their anger.
PS|55|4|My heart is in anguish within me; the terrors of death assail me.
PS|55|5|Fear and trembling have beset me; horror has overwhelmed me.
PS|55|6|I said, "Oh, that I had the wings of a dove! I would fly away and be at rest-
PS|55|7|I would flee far away and stay in the desert; Selah
PS|55|8|I would hurry to my place of shelter, far from the tempest and storm."
PS|55|9|Confuse the wicked, O Lord, confound their speech, for I see violence and strife in the city.
PS|55|10|Day and night they prowl about on its walls; malice and abuse are within it.
PS|55|11|Destructive forces are at work in the city; threats and lies never leave its streets.
PS|55|12|If an enemy were insulting me, I could endure it; if a foe were raising himself against me, I could hide from him.
PS|55|13|But it is you, a man like myself, my companion, my close friend,
PS|55|14|with whom I once enjoyed sweet fellowship as we walked with the throng at the house of God.
PS|55|15|Let death take my enemies by surprise; let them go down alive to the grave, for evil finds lodging among them.
PS|55|16|But I call to God, and the LORD saves me.
PS|55|17|Evening, morning and noon I cry out in distress, and he hears my voice.
PS|55|18|He ransoms me unharmed from the battle waged against me, even though many oppose me.
PS|55|19|God, who is enthroned forever, will hear them and afflict them- Selah men who never change their ways and have no fear of God.
PS|55|20|My companion attacks his friends; he violates his covenant.
PS|55|21|His speech is smooth as butter, yet war is in his heart; his words are more soothing than oil, yet they are drawn swords.
PS|55|22|Cast your cares on the LORD and he will sustain you; he will never let the righteous fall.
PS|55|23|But you, O God, will bring down the wicked into the pit of corruption; bloodthirsty and deceitful men will not live out half their days. But as for me, I trust in you.
PS|56|1|Be merciful to me, O God, for men hotly pursue me; all day long they press their attack.
PS|56|2|My slanderers pursue me all day long; many are attacking me in their pride.
PS|56|3|When I am afraid, I will trust in you.
PS|56|4|In God, whose word I praise, in God I trust; I will not be afraid. What can mortal man do to me?
PS|56|5|All day long they twist my words; they are always plotting to harm me.
PS|56|6|They conspire, they lurk, they watch my steps, eager to take my life.
PS|56|7|On no account let them escape; in your anger, O God, bring down the nations.
PS|56|8|Record my lament; list my tears on your scroll - are they not in your record?
PS|56|9|Then my enemies will turn back when I call for help. By this I will know that God is for me.
PS|56|10|In God, whose word I praise, in the LORD, whose word I praise-
PS|56|11|in God I trust; I will not be afraid. What can man do to me?
PS|56|12|I am under vows to you, O God; I will present my thank offerings to you.
PS|56|13|For you have delivered me from death and my feet from stumbling, that I may walk before God in the light of life.
PS|57|1|Have mercy on me, O God, have mercy on me, for in you my soul takes refuge. I will take refuge in the shadow of your wings until the disaster has passed.
PS|57|2|I cry out to God Most High, to God, who fulfills {his purpose} for me.
PS|57|3|He sends from heaven and saves me, rebuking those who hotly pursue me; Selah God sends his love and his faithfulness.
PS|57|4|I am in the midst of lions; I lie among ravenous beasts- men whose teeth are spears and arrows, whose tongues are sharp swords.
PS|57|5|Be exalted, O God, above the heavens; let your glory be over all the earth.
PS|57|6|They spread a net for my feet- I was bowed down in distress. They dug a pit in my path- but they have fallen into it themselves. Selah
PS|57|7|My heart is steadfast, O God, my heart is steadfast; I will sing and make music.
PS|57|8|Awake, my soul! Awake, harp and lyre! I will awaken the dawn.
PS|57|9|I will praise you, O Lord, among the nations; I will sing of you among the peoples.
PS|57|10|For great is your love, reaching to the heavens; your faithfulness reaches to the skies.
PS|57|11|Be exalted, O God, above the heavens; let your glory be over all the earth.
PS|58|1|Do you rulers indeed speak justly? Do you judge uprightly among men?
PS|58|2|No, in your heart you devise injustice, and your hands mete out violence on the earth.
PS|58|3|Even from birth the wicked go astray; from the womb they are wayward and speak lies.
PS|58|4|Their venom is like the venom of a snake, like that of a cobra that has stopped its ears,
PS|58|5|that will not heed the tune of the charmer, however skillful the enchanter may be.
PS|58|6|Break the teeth in their mouths, O God; tear out, O LORD, the fangs of the lions!
PS|58|7|Let them vanish like water that flows away; when they draw the bow, let their arrows be blunted.
PS|58|8|Like a slug melting away as it moves along, like a stillborn child, may they not see the sun.
PS|58|9|Before your pots can feel the heat of the thorns- whether they be green or dry-the wicked will be swept away.
PS|58|10|The righteous will be glad when they are avenged, when they bathe their feet in the blood of the wicked.
PS|58|11|Then men will say, "Surely the righteous still are rewarded; surely there is a God who judges the earth."
PS|59|1|Deliver me from my enemies, O God; protect me from those who rise up against me.
PS|59|2|Deliver me from evildoers and save me from bloodthirsty men.
PS|59|3|See how they lie in wait for me! Fierce men conspire against me for no offense or sin of mine, O LORD.
PS|59|4|I have done no wrong, yet they are ready to attack me. Arise to help me; look on my plight!
PS|59|5|O LORD God Almighty, the God of Israel, rouse yourself to punish all the nations; show no mercy to wicked traitors. Selah
PS|59|6|They return at evening, snarling like dogs, and prowl about the city.
PS|59|7|See what they spew from their mouths- they spew out swords from their lips, and they say, "Who can hear us?"
PS|59|8|But you, O LORD, laugh at them; you scoff at all those nations.
PS|59|9|O my Strength, I watch for you; you, O God, are my fortress,
PS|59|10|my loving God. God will go before me and will let me gloat over those who slander me.
PS|59|11|But do not kill them, O Lord our shield, or my people will forget. In your might make them wander about, and bring them down.
PS|59|12|For the sins of their mouths, for the words of their lips, let them be caught in their pride. For the curses and lies they utter,
PS|59|13|consume them in wrath, consume them till they are no more. Then it will be known to the ends of the earth that God rules over Jacob. Selah
PS|59|14|They return at evening, snarling like dogs, and prowl about the city.
PS|59|15|They wander about for food and howl if not satisfied.
PS|59|16|But I will sing of your strength, in the morning I will sing of your love; for you are my fortress, my refuge in times of trouble.
PS|59|17|O my Strength, I sing praise to you; you, O God, are my fortress, my loving God.
PS|60|1|You have rejected us, O God, and burst forth upon us; you have been angry-now restore us!
PS|60|2|You have shaken the land and torn it open; mend its fractures, for it is quaking.
PS|60|3|You have shown your people desperate times; you have given us wine that makes us stagger.
PS|60|4|But for those who fear you, you have raised a banner to be unfurled against the bow. Selah
PS|60|5|Save us and help us with your right hand, that those you love may be delivered.
PS|60|6|God has spoken from his sanctuary: "In triumph I will parcel out Shechem and measure off the Valley of Succoth.
PS|60|7|Gilead is mine, and Manasseh is mine; Ephraim is my helmet, Judah my scepter.
PS|60|8|Moab is my washbasin, upon Edom I toss my sandal; over Philistia I shout in triumph."
PS|60|9|Who will bring me to the fortified city? Who will lead me to Edom?
PS|60|10|Is it not you, O God, you who have rejected us and no longer go out with our armies?
PS|60|11|Give us aid against the enemy, for the help of man is worthless.
PS|60|12|With God we will gain the victory, and he will trample down our enemies.
PS|61|1|Hear my cry, O God; listen to my prayer.
PS|61|2|From the ends of the earth I call to you, I call as my heart grows faint; lead me to the rock that is higher than I.
PS|61|3|For you have been my refuge, a strong tower against the foe.
PS|61|4|I long to dwell in your tent forever and take refuge in the shelter of your wings. Selah
PS|61|5|For you have heard my vows, O God; you have given me the heritage of those who fear your name.
PS|61|6|Increase the days of the king's life, his years for many generations.
PS|61|7|May he be enthroned in God's presence forever; appoint your love and faithfulness to protect him.
PS|61|8|Then will I ever sing praise to your name and fulfill my vows day after day.
PS|62|1|My soul finds rest in God alone; my salvation comes from him.
PS|62|2|He alone is my rock and my salvation; he is my fortress, I will never be shaken.
PS|62|3|How long will you assault a man? Would all of you throw him down- this leaning wall, this tottering fence?
PS|62|4|They fully intend to topple him from his lofty place; they take delight in lies. With their mouths they bless, but in their hearts they curse. Selah
PS|62|5|Find rest, O my soul, in God alone; my hope comes from him.
PS|62|6|He alone is my rock and my salvation; he is my fortress, I will not be shaken.
PS|62|7|My salvation and my honor depend on God; he is my mighty rock, my refuge.
PS|62|8|Trust in him at all times, O people; pour out your hearts to him, for God is our refuge. Selah
PS|62|9|Lowborn men are but a breath, the highborn are but a lie; if weighed on a balance, they are nothing; together they are only a breath.
PS|62|10|Do not trust in extortion or take pride in stolen goods; though your riches increase, do not set your heart on them.
PS|62|11|One thing God has spoken, two things have I heard: that you, O God, are strong,
PS|62|12|and that you, O Lord, are loving. Surely you will reward each person according to what he has done.
PS|63|1|O God, you are my God, earnestly I seek you; my soul thirsts for you, my body longs for you, in a dry and weary land where there is no water.
PS|63|2|I have seen you in the sanctuary and beheld your power and your glory.
PS|63|3|Because your love is better than life, my lips will glorify you.
PS|63|4|I will praise you as long as I live, and in your name I will lift up my hands.
PS|63|5|My soul will be satisfied as with the richest of foods; with singing lips my mouth will praise you.
PS|63|6|On my bed I remember you; I think of you through the watches of the night.
PS|63|7|Because you are my help, I sing in the shadow of your wings.
PS|63|8|My soul clings to you; your right hand upholds me.
PS|63|9|They who seek my life will be destroyed; they will go down to the depths of the earth.
PS|63|10|They will be given over to the sword and become food for jackals.
PS|63|11|But the king will rejoice in God; all who swear by God's name will praise him, while the mouths of liars will be silenced.
PS|64|1|Hear me, O God, as I voice my complaint; protect my life from the threat of the enemy.
PS|64|2|Hide me from the conspiracy of the wicked, from that noisy crowd of evildoers.
PS|64|3|They sharpen their tongues like swords and aim their words like deadly arrows.
PS|64|4|They shoot from ambush at the innocent man; they shoot at him suddenly, without fear.
PS|64|5|They encourage each other in evil plans, they talk about hiding their snares; they say, "Who will see them?"
PS|64|6|They plot injustice and say, "We have devised a perfect plan!" Surely the mind and heart of man are cunning.
PS|64|7|But God will shoot them with arrows; suddenly they will be struck down.
PS|64|8|He will turn their own tongues against them and bring them to ruin; all who see them will shake their heads in scorn.
PS|64|9|All mankind will fear; they will proclaim the works of God and ponder what he has done.
PS|64|10|Let the righteous rejoice in the LORD and take refuge in him; let all the upright in heart praise him!
PS|65|1|Praise awaits you, O God, in Zion; to you our vows will be fulfilled.
PS|65|2|O you who hear prayer, to you all men will come.
PS|65|3|When we were overwhelmed by sins, you forgave our transgressions.
PS|65|4|Blessed are those you choose and bring near to live in your courts! We are filled with the good things of your house, of your holy temple.
PS|65|5|You answer us with awesome deeds of righteousness, O God our Savior, the hope of all the ends of the earth and of the farthest seas,
PS|65|6|who formed the mountains by your power, having armed yourself with strength,
PS|65|7|who stilled the roaring of the seas, the roaring of their waves, and the turmoil of the nations.
PS|65|8|Those living far away fear your wonders; where morning dawns and evening fades you call forth songs of joy.
PS|65|9|You care for the land and water it; you enrich it abundantly. The streams of God are filled with water to provide the people with grain, for so you have ordained it.
PS|65|10|You drench its furrows and level its ridges; you soften it with showers and bless its crops.
PS|65|11|You crown the year with your bounty, and your carts overflow with abundance.
PS|65|12|The grasslands of the desert overflow; the hills are clothed with gladness.
PS|65|13|The meadows are covered with flocks and the valleys are mantled with grain; they shout for joy and sing.
PS|66|1|Shout with joy to God, all the earth!
PS|66|2|Sing the glory of his name; make his praise glorious!
PS|66|3|Say to God, "How awesome are your deeds! So great is your power that your enemies cringe before you.
PS|66|4|All the earth bows down to you; they sing praise to you, they sing praise to your name." Selah
PS|66|5|Come and see what God has done, how awesome his works in man's behalf!
PS|66|6|He turned the sea into dry land, they passed through the waters on foot- come, let us rejoice in him.
PS|66|7|He rules forever by his power, his eyes watch the nations- let not the rebellious rise up against him. Selah
PS|66|8|Praise our God, O peoples, let the sound of his praise be heard;
PS|66|9|he has preserved our lives and kept our feet from slipping.
PS|66|10|For you, O God, tested us; you refined us like silver.
PS|66|11|You brought us into prison and laid burdens on our backs.
PS|66|12|You let men ride over our heads; we went through fire and water, but you brought us to a place of abundance.
PS|66|13|I will come to your temple with burnt offerings and fulfill my vows to you-
PS|66|14|vows my lips promised and my mouth spoke when I was in trouble.
PS|66|15|I will sacrifice fat animals to you and an offering of rams; I will offer bulls and goats. Selah
PS|66|16|Come and listen, all you who fear God; let me tell you what he has done for me.
PS|66|17|I cried out to him with my mouth; his praise was on my tongue.
PS|66|18|If I had cherished sin in my heart, the Lord would not have listened;
PS|66|19|but God has surely listened and heard my voice in prayer.
PS|66|20|Praise be to God, who has not rejected my prayer or withheld his love from me!
PS|67|1|May God be gracious to us and bless us and make his face shine upon us, Selah
PS|67|2|that your ways may be known on earth, your salvation among all nations.
PS|67|3|May the peoples praise you, O God; may all the peoples praise you.
PS|67|4|May the nations be glad and sing for joy, for you rule the peoples justly and guide the nations of the earth. Selah
PS|67|5|May the peoples praise you, O God; may all the peoples praise you.
PS|67|6|Then the land will yield its harvest, and God, our God, will bless us.
PS|67|7|God will bless us, and all the ends of the earth will fear him.
PS|68|1|May God arise, may his enemies be scattered; may his foes flee before him.
PS|68|2|As smoke is blown away by the wind, may you blow them away; as wax melts before the fire, may the wicked perish before God.
PS|68|3|But may the righteous be glad and rejoice before God; may they be happy and joyful.
PS|68|4|Sing to God, sing praise to his name, extol him who rides on the clouds - his name is the LORD - and rejoice before him.
PS|68|5|A father to the fatherless, a defender of widows, is God in his holy dwelling.
PS|68|6|God sets the lonely in families, he leads forth the prisoners with singing; but the rebellious live in a sun-scorched land.
PS|68|7|When you went out before your people, O God, when you marched through the wasteland, Selah
PS|68|8|the earth shook, the heavens poured down rain, before God, the One of Sinai, before God, the God of Israel.
PS|68|9|You gave abundant showers, O God; you refreshed your weary inheritance.
PS|68|10|Your people settled in it, and from your bounty, O God, you provided for the poor.
PS|68|11|The Lord announced the word, and great was the company of those who proclaimed it:
PS|68|12|"Kings and armies flee in haste; in the camps men divide the plunder.
PS|68|13|Even while you sleep among the campfires, the wings of my dove are sheathed with silver, its feathers with shining gold."
PS|68|14|When the Almighty scattered the kings in the land, it was like snow fallen on Zalmon.
PS|68|15|The mountains of Bashan are majestic mountains; rugged are the mountains of Bashan.
PS|68|16|Why gaze in envy, O rugged mountains, at the mountain where God chooses to reign, where the LORD himself will dwell forever?
PS|68|17|The chariots of God are tens of thousands and thousands of thousands; the Lord has come from Sinai into his sanctuary.
PS|68|18|When you ascended on high, you led captives in your train; you received gifts from men, even from the rebellious- that you, O LORD God, might dwell there.
PS|68|19|Praise be to the Lord, to God our Savior, who daily bears our burdens. Selah
PS|68|20|Our God is a God who saves; from the Sovereign LORD comes escape from death.
PS|68|21|Surely God will crush the heads of his enemies, the hairy crowns of those who go on in their sins.
PS|68|22|The Lord says, "I will bring them from Bashan; I will bring them from the depths of the sea,
PS|68|23|that you may plunge your feet in the blood of your foes, while the tongues of your dogs have their share."
PS|68|24|Your procession has come into view, O God, the procession of my God and King into the sanctuary.
PS|68|25|In front are the singers, after them the musicians; with them are the maidens playing tambourines.
PS|68|26|Praise God in the great congregation; praise the LORD in the assembly of Israel.
PS|68|27|There is the little tribe of Benjamin, leading them, there the great throng of Judah's princes, and there the princes of Zebulun and of Naphtali.
PS|68|28|Summon your power, O God; show us your strength, O God, as you have done before.
PS|68|29|Because of your temple at Jerusalem kings will bring you gifts.
PS|68|30|Rebuke the beast among the reeds, the herd of bulls among the calves of the nations. Humbled, may it bring bars of silver. Scatter the nations who delight in war.
PS|68|31|Envoys will come from Egypt; Cush will submit herself to God.
PS|68|32|Sing to God, O kingdoms of the earth, sing praise to the Lord, Selah
PS|68|33|to him who rides the ancient skies above, who thunders with mighty voice.
PS|68|34|Proclaim the power of God, whose majesty is over Israel, whose power is in the skies.
PS|68|35|You are awesome, O God, in your sanctuary; the God of Israel gives power and strength to his people. Praise be to God!
PS|69|1|Save me, O God, for the waters have come up to my neck.
PS|69|2|I sink in the miry depths, where there is no foothold. I have come into the deep waters; the floods engulf me.
PS|69|3|I am worn out calling for help; my throat is parched. My eyes fail, looking for my God.
PS|69|4|Those who hate me without reason outnumber the hairs of my head; many are my enemies without cause, those who seek to destroy me. I am forced to restore what I did not steal.
PS|69|5|You know my folly, O God; my guilt is not hidden from you.
PS|69|6|May those who hope in you not be disgraced because of me, O Lord, the LORD Almighty; may those who seek you not be put to shame because of me, O God of Israel.
PS|69|7|For I endure scorn for your sake, and shame covers my face.
PS|69|8|I am a stranger to my brothers, an alien to my own mother's sons;
PS|69|9|for zeal for your house consumes me, and the insults of those who insult you fall on me.
PS|69|10|When I weep and fast, I must endure scorn;
PS|69|11|when I put on sackcloth, people make sport of me.
PS|69|12|Those who sit at the gate mock me, and I am the song of the drunkards.
PS|69|13|But I pray to you, O LORD, in the time of your favor; in your great love, O God, answer me with your sure salvation.
PS|69|14|Rescue me from the mire, do not let me sink; deliver me from those who hate me, from the deep waters.
PS|69|15|Do not let the floodwaters engulf me or the depths swallow me up or the pit close its mouth over me.
PS|69|16|Answer me, O LORD, out of the goodness of your love; in your great mercy turn to me.
PS|69|17|Do not hide your face from your servant; answer me quickly, for I am in trouble.
PS|69|18|Come near and rescue me; redeem me because of my foes.
PS|69|19|You know how I am scorned, disgraced and shamed; all my enemies are before you.
PS|69|20|Scorn has broken my heart and has left me helpless; I looked for sympathy, but there was none, for comforters, but I found none.
PS|69|21|They put gall in my food and gave me vinegar for my thirst.
PS|69|22|May the table set before them become a snare; may it become retribution and a trap.
PS|69|23|May their eyes be darkened so they cannot see, and their backs be bent forever.
PS|69|24|Pour out your wrath on them; let your fierce anger overtake them.
PS|69|25|May their place be deserted; let there be no one to dwell in their tents.
PS|69|26|For they persecute those you wound and talk about the pain of those you hurt.
PS|69|27|Charge them with crime upon crime; do not let them share in your salvation.
PS|69|28|May they be blotted out of the book of life and not be listed with the righteous.
PS|69|29|I am in pain and distress; may your salvation, O God, protect me.
PS|69|30|I will praise God's name in song and glorify him with thanksgiving.
PS|69|31|This will please the LORD more than an ox, more than a bull with its horns and hoofs.
PS|69|32|The poor will see and be glad- you who seek God, may your hearts live!
PS|69|33|The LORD hears the needy and does not despise his captive people.
PS|69|34|Let heaven and earth praise him, the seas and all that move in them,
PS|69|35|for God will save Zion and rebuild the cities of Judah. Then people will settle there and possess it;
PS|69|36|the children of his servants will inherit it, and those who love his name will dwell there.
PS|70|1|Hasten, O God, to save me; O LORD, come quickly to help me.
PS|70|2|May those who seek my life be put to shame and confusion; may all who desire my ruin be turned back in disgrace.
PS|70|3|May those who say to me, "Aha! Aha!" turn back because of their shame.
PS|70|4|But may all who seek you rejoice and be glad in you; may those who love your salvation always say, "Let God be exalted!"
PS|70|5|Yet I am poor and needy; come quickly to me, O God. You are my help and my deliverer; O LORD, do not delay.
PS|71|1|In you, O LORD, I have taken refuge; let me never be put to shame.
PS|71|2|Rescue me and deliver me in your righteousness; turn your ear to me and save me.
PS|71|3|Be my rock of refuge, to which I can always go; give the command to save me, for you are my rock and my fortress.
PS|71|4|Deliver me, O my God, from the hand of the wicked, from the grasp of evil and cruel men.
PS|71|5|For you have been my hope, O Sovereign LORD, my confidence since my youth.
PS|71|6|From birth I have relied on you; you brought me forth from my mother's womb. I will ever praise you.
PS|71|7|I have become like a portent to many, but you are my strong refuge.
PS|71|8|My mouth is filled with your praise, declaring your splendor all day long.
PS|71|9|Do not cast me away when I am old; do not forsake me when my strength is gone.
PS|71|10|For my enemies speak against me; those who wait to kill me conspire together.
PS|71|11|They say, "God has forsaken him; pursue him and seize him, for no one will rescue him."
PS|71|12|Be not far from me, O God; come quickly, O my God, to help me.
PS|71|13|May my accusers perish in shame; may those who want to harm me be covered with scorn and disgrace.
PS|71|14|But as for me, I will always have hope; I will praise you more and more.
PS|71|15|My mouth will tell of your righteousness, of your salvation all day long, though I know not its measure.
PS|71|16|I will come and proclaim your mighty acts, O Sovereign LORD; I will proclaim your righteousness, yours alone.
PS|71|17|Since my youth, O God, you have taught me, and to this day I declare your marvelous deeds.
PS|71|18|Even when I am old and gray, do not forsake me, O God, till I declare your power to the next generation, your might to all who are to come.
PS|71|19|Your righteousness reaches to the skies, O God, you who have done great things. Who, O God, is like you?
PS|71|20|Though you have made me see troubles, many and bitter, you will restore my life again; from the depths of the earth you will again bring me up.
PS|71|21|You will increase my honor and comfort me once again.
PS|71|22|I will praise you with the harp for your faithfulness, O my God; I will sing praise to you with the lyre, O Holy One of Israel.
PS|71|23|My lips will shout for joy when I sing praise to you- I, whom you have redeemed.
PS|71|24|My tongue will tell of your righteous acts all day long, for those who wanted to harm me have been put to shame and confusion.
PS|72|1|Endow the king with your justice, O God, the royal son with your righteousness.
PS|72|2|He will judge your people in righteousness, your afflicted ones with justice.
PS|72|3|The mountains will bring prosperity to the people, the hills the fruit of righteousness.
PS|72|4|He will defend the afflicted among the people and save the children of the needy; he will crush the oppressor.
PS|72|5|He will endure as long as the sun, as long as the moon, through all generations.
PS|72|6|He will be like rain falling on a mown field, like showers watering the earth.
PS|72|7|In his days the righteous will flourish; prosperity will abound till the moon is no more.
PS|72|8|He will rule from sea to sea and from the River to the ends of the earth.
PS|72|9|The desert tribes will bow before him and his enemies will lick the dust.
PS|72|10|The kings of Tarshish and of distant shores will bring tribute to him; the kings of Sheba and Seba will present him gifts.
PS|72|11|All kings will bow down to him and all nations will serve him.
PS|72|12|For he will deliver the needy who cry out, the afflicted who have no one to help.
PS|72|13|He will take pity on the weak and the needy and save the needy from death.
PS|72|14|He will rescue them from oppression and violence, for precious is their blood in his sight.
PS|72|15|Long may he live! May gold from Sheba be given him. May people ever pray for him and bless him all day long.
PS|72|16|Let grain abound throughout the land; on the tops of the hills may it sway. Let its fruit flourish like Lebanon; let it thrive like the grass of the field.
PS|72|17|May his name endure forever; may it continue as long as the sun. All nations will be blessed through him, and they will call him blessed.
PS|72|18|Praise be to the LORD God, the God of Israel, who alone does marvelous deeds.
PS|72|19|Praise be to his glorious name forever; may the whole earth be filled with his glory. Amen and Amen.
PS|72|20|This concludes the prayers of David son of Jesse.
PS|73|1|A psalm of Asaph. Surely God is good to Israel, to those who are pure in heart.
PS|73|2|But as for me, my feet had almost slipped; I had nearly lost my foothold.
PS|73|3|For I envied the arrogant when I saw the prosperity of the wicked.
PS|73|4|They have no struggles; their bodies are healthy and strong.
PS|73|5|They are free from the burdens common to man; they are not plagued by human ills.
PS|73|6|Therefore pride is their necklace; they clothe themselves with violence.
PS|73|7|From their callous hearts comes iniquity; the evil conceits of their minds know no limits.
PS|73|8|They scoff, and speak with malice; in their arrogance they threaten oppression.
PS|73|9|Their mouths lay claim to heaven, and their tongues take possession of the earth.
PS|73|10|Therefore their people turn to them and drink up waters in abundance.
PS|73|11|They say, "How can God know? Does the Most High have knowledge?"
PS|73|12|This is what the wicked are like- always carefree, they increase in wealth.
PS|73|13|Surely in vain have I kept my heart pure; in vain have I washed my hands in innocence.
PS|73|14|All day long I have been plagued; I have been punished every morning.
PS|73|15|If I had said, "I will speak thus," I would have betrayed your children.
PS|73|16|When I tried to understand all this, it was oppressive to me
PS|73|17|till I entered the sanctuary of God; then I understood their final destiny.
PS|73|18|Surely you place them on slippery ground; you cast them down to ruin.
PS|73|19|How suddenly are they destroyed, completely swept away by terrors!
PS|73|20|As a dream when one awakes, so when you arise, O Lord, you will despise them as fantasies.
PS|73|21|When my heart was grieved and my spirit embittered,
PS|73|22|I was senseless and ignorant; I was a brute beast before you.
PS|73|23|Yet I am always with you; you hold me by my right hand.
PS|73|24|You guide me with your counsel, and afterward you will take me into glory.
PS|73|25|Whom have I in heaven but you? And earth has nothing I desire besides you.
PS|73|26|My flesh and my heart may fail, but God is the strength of my heart and my portion forever.
PS|73|27|Those who are far from you will perish; you destroy all who are unfaithful to you.
PS|73|28|But as for me, it is good to be near God. I have made the Sovereign LORD my refuge; I will tell of all your deeds.
PS|74|1|Why have you rejected us forever, O God? Why does your anger smolder against the sheep of your pasture?
PS|74|2|Remember the people you purchased of old, the tribe of your inheritance, whom you redeemed- Mount Zion, where you dwelt.
PS|74|3|Turn your steps toward these everlasting ruins, all this destruction the enemy has brought on the sanctuary.
PS|74|4|Your foes roared in the place where you met with us; they set up their standards as signs.
PS|74|5|They behaved like men wielding axes to cut through a thicket of trees.
PS|74|6|They smashed all the carved paneling with their axes and hatchets.
PS|74|7|They burned your sanctuary to the ground; they defiled the dwelling place of your Name.
PS|74|8|They said in their hearts, "We will crush them completely!" They burned every place where God was worshiped in the land.
PS|74|9|We are given no miraculous signs; no prophets are left, and none of us knows how long this will be.
PS|74|10|How long will the enemy mock you, O God? Will the foe revile your name forever?
PS|74|11|Why do you hold back your hand, your right hand? Take it from the folds of your garment and destroy them!
PS|74|12|But you, O God, are my king from of old; you bring salvation upon the earth.
PS|74|13|It was you who split open the sea by your power; you broke the heads of the monster in the waters.
PS|74|14|It was you who crushed the heads of Leviathan and gave him as food to the creatures of the desert.
PS|74|15|It was you who opened up springs and streams; you dried up the ever flowing rivers.
PS|74|16|The day is yours, and yours also the night; you established the sun and moon.
PS|74|17|It was you who set all the boundaries of the earth; you made both summer and winter.
PS|74|18|Remember how the enemy has mocked you, O LORD, how foolish people have reviled your name.
PS|74|19|Do not hand over the life of your dove to wild beasts; do not forget the lives of your afflicted people forever.
PS|74|20|Have regard for your covenant, because haunts of violence fill the dark places of the land.
PS|74|21|Do not let the oppressed retreat in disgrace; may the poor and needy praise your name.
PS|74|22|Rise up, O God, and defend your cause; remember how fools mock you all day long.
PS|74|23|Do not ignore the clamor of your adversaries, the uproar of your enemies, which rises continually.
PS|75|1|We give thanks to you, O God, we give thanks, for your Name is near; men tell of your wonderful deeds.
PS|75|2|You say, "I choose the appointed time; it is I who judge uprightly.
PS|75|3|When the earth and all its people quake, it is I who hold its pillars firm. Selah
PS|75|4|To the arrogant I say, 'Boast no more,' and to the wicked, 'Do not lift up your horns.
PS|75|5|Do not lift your horns against heaven; do not speak with outstretched neck.'"
PS|75|6|No one from the east or the west or from the desert can exalt a man.
PS|75|7|But it is God who judges: He brings one down, he exalts another.
PS|75|8|In the hand of the LORD is a cup full of foaming wine mixed with spices; he pours it out, and all the wicked of the earth drink it down to its very dregs.
PS|75|9|As for me, I will declare this forever; I will sing praise to the God of Jacob.
PS|75|10|I will cut off the horns of all the wicked, but the horns of the righteous will be lifted up.
PS|76|1|In Judah God is known; his name is great in Israel.
PS|76|2|His tent is in Salem, his dwelling place in Zion.
PS|76|3|There he broke the flashing arrows, the shields and the swords, the weapons of war. Selah
PS|76|4|You are resplendent with light, more majestic than mountains rich with game.
PS|76|5|Valiant men lie plundered, they sleep their last sleep; not one of the warriors can lift his hands.
PS|76|6|At your rebuke, O God of Jacob, both horse and chariot lie still.
PS|76|7|You alone are to be feared. Who can stand before you when you are angry?
PS|76|8|From heaven you pronounced judgment, and the land feared and was quiet-
PS|76|9|when you, O God, rose up to judge, to save all the afflicted of the land. Selah
PS|76|10|Surely your wrath against men brings you praise, and the survivors of your wrath are restrained.
PS|76|11|Make vows to the LORD your God and fulfill them; let all the neighboring lands bring gifts to the One to be feared.
PS|76|12|He breaks the spirit of rulers; he is feared by the kings of the earth.
PS|77|1|I cried out to God for help; I cried out to God to hear me.
PS|77|2|When I was in distress, I sought the Lord; at night I stretched out untiring hands and my soul refused to be comforted.
PS|77|3|I remembered you, O God, and I groaned; I mused, and my spirit grew faint. Selah
PS|77|4|You kept my eyes from closing; I was too troubled to speak.
PS|77|5|I thought about the former days, the years of long ago;
PS|77|6|I remembered my songs in the night. My heart mused and my spirit inquired:
PS|77|7|"Will the Lord reject forever? Will he never show his favor again?
PS|77|8|Has his unfailing love vanished forever? Has his promise failed for all time?
PS|77|9|Has God forgotten to be merciful? Has he in anger withheld his compassion?" Selah
PS|77|10|Then I thought, "To this I will appeal: the years of the right hand of the Most High."
PS|77|11|I will remember the deeds of the LORD; yes, I will remember your miracles of long ago.
PS|77|12|I will meditate on all your works and consider all your mighty deeds.
PS|77|13|Your ways, O God, are holy. What god is so great as our God?
PS|77|14|You are the God who performs miracles; you display your power among the peoples.
PS|77|15|With your mighty arm you redeemed your people, the descendants of Jacob and Joseph. Selah
PS|77|16|The waters saw you, O God, the waters saw you and writhed; the very depths were convulsed.
PS|77|17|The clouds poured down water, the skies resounded with thunder; your arrows flashed back and forth.
PS|77|18|Your thunder was heard in the whirlwind, your lightning lit up the world; the earth trembled and quaked.
PS|77|19|Your path led through the sea, your way through the mighty waters, though your footprints were not seen.
PS|77|20|You led your people like a flock by the hand of Moses and Aaron.
PS|78|1|O my people, hear my teaching; listen to the words of my mouth.
PS|78|2|I will open my mouth in parables, I will utter hidden things, things from of old-
PS|78|3|what we have heard and known, what our fathers have told us.
PS|78|4|We will not hide them from their children; we will tell the next generation the praiseworthy deeds of the LORD, his power, and the wonders he has done.
PS|78|5|He decreed statutes for Jacob and established the law in Israel, which he commanded our forefathers to teach their children,
PS|78|6|so the next generation would know them, even the children yet to be born, and they in turn would tell their children.
PS|78|7|Then they would put their trust in God and would not forget his deeds but would keep his commands.
PS|78|8|They would not be like their forefathers- a stubborn and rebellious generation, whose hearts were not loyal to God, whose spirits were not faithful to him.
PS|78|9|The men of Ephraim, though armed with bows, turned back on the day of battle;
PS|78|10|they did not keep God's covenant and refused to live by his law.
PS|78|11|They forgot what he had done, the wonders he had shown them.
PS|78|12|He did miracles in the sight of their fathers in the land of Egypt, in the region of Zoan.
PS|78|13|He divided the sea and led them through; he made the water stand firm like a wall.
PS|78|14|He guided them with the cloud by day and with light from the fire all night.
PS|78|15|He split the rocks in the desert and gave them water as abundant as the seas;
PS|78|16|he brought streams out of a rocky crag and made water flow down like rivers.
PS|78|17|But they continued to sin against him, rebelling in the desert against the Most High.
PS|78|18|They willfully put God to the test by demanding the food they craved.
PS|78|19|They spoke against God, saying, "Can God spread a table in the desert?
PS|78|20|When he struck the rock, water gushed out, and streams flowed abundantly. But can he also give us food? Can he supply meat for his people?"
PS|78|21|When the LORD heard them, he was very angry; his fire broke out against Jacob, and his wrath rose against Israel,
PS|78|22|for they did not believe in God or trust in his deliverance.
PS|78|23|Yet he gave a command to the skies above and opened the doors of the heavens;
PS|78|24|he rained down manna for the people to eat, he gave them the grain of heaven.
PS|78|25|Men ate the bread of angels; he sent them all the food they could eat.
PS|78|26|He let loose the east wind from the heavens and led forth the south wind by his power.
PS|78|27|He rained meat down on them like dust, flying birds like sand on the seashore.
PS|78|28|He made them come down inside their camp, all around their tents.
PS|78|29|They ate till they had more than enough, for he had given them what they craved.
PS|78|30|But before they turned from the food they craved, even while it was still in their mouths,
PS|78|31|God's anger rose against them; he put to death the sturdiest among them, cutting down the young men of Israel.
PS|78|32|In spite of all this, they kept on sinning; in spite of his wonders, they did not believe.
PS|78|33|So he ended their days in futility and their years in terror.
PS|78|34|Whenever God slew them, they would seek him; they eagerly turned to him again.
PS|78|35|They remembered that God was their Rock, that God Most High was their Redeemer.
PS|78|36|But then they would flatter him with their mouths, lying to him with their tongues;
PS|78|37|their hearts were not loyal to him, they were not faithful to his covenant.
PS|78|38|Yet he was merciful; he forgave their iniquities and did not destroy them. Time after time he restrained his anger and did not stir up his full wrath.
PS|78|39|He remembered that they were but flesh, a passing breeze that does not return.
PS|78|40|How often they rebelled against him in the desert and grieved him in the wasteland!
PS|78|41|Again and again they put God to the test; they vexed the Holy One of Israel.
PS|78|42|They did not remember his power- the day he redeemed them from the oppressor,
PS|78|43|the day he displayed his miraculous signs in Egypt, his wonders in the region of Zoan.
PS|78|44|He turned their rivers to blood; they could not drink from their streams.
PS|78|45|He sent swarms of flies that devoured them, and frogs that devastated them.
PS|78|46|He gave their crops to the grasshopper, their produce to the locust.
PS|78|47|He destroyed their vines with hail and their sycamore-figs with sleet.
PS|78|48|He gave over their cattle to the hail, their livestock to bolts of lightning.
PS|78|49|He unleashed against them his hot anger, his wrath, indignation and hostility- a band of destroying angels.
PS|78|50|He prepared a path for his anger; he did not spare them from death but gave them over to the plague.
PS|78|51|He struck down all the firstborn of Egypt, the firstfruits of manhood in the tents of Ham.
PS|78|52|But he brought his people out like a flock; he led them like sheep through the desert.
PS|78|53|He guided them safely, so they were unafraid; but the sea engulfed their enemies.
PS|78|54|Thus he brought them to the border of his holy land, to the hill country his right hand had taken.
PS|78|55|He drove out nations before them and allotted their lands to them as an inheritance; he settled the tribes of Israel in their homes.
PS|78|56|But they put God to the test and rebelled against the Most High; they did not keep his statutes.
PS|78|57|Like their fathers they were disloyal and faithless, as unreliable as a faulty bow.
PS|78|58|They angered him with their high places; they aroused his jealousy with their idols.
PS|78|59|When God heard them, he was very angry; he rejected Israel completely.
PS|78|60|He abandoned the tabernacle of Shiloh, the tent he had set up among men.
PS|78|61|He sent the ark of his might into captivity, his splendor into the hands of the enemy.
PS|78|62|He gave his people over to the sword; he was very angry with his inheritance.
PS|78|63|Fire consumed their young men, and their maidens had no wedding songs;
PS|78|64|their priests were put to the sword, and their widows could not weep.
PS|78|65|Then the Lord awoke as from sleep, as a man wakes from the stupor of wine.
PS|78|66|He beat back his enemies; he put them to everlasting shame.
PS|78|67|Then he rejected the tents of Joseph, he did not choose the tribe of Ephraim;
PS|78|68|but he chose the tribe of Judah, Mount Zion, which he loved.
PS|78|69|He built his sanctuary like the heights, like the earth that he established forever.
PS|78|70|He chose David his servant and took him from the sheep pens;
PS|78|71|from tending the sheep he brought him to be the shepherd of his people Jacob, of Israel his inheritance.
PS|78|72|And David shepherded them with integrity of heart; with skillful hands he led them.
PS|79|1|O God, the nations have invaded your inheritance; they have defiled your holy temple, they have reduced Jerusalem to rubble.
PS|79|2|They have given the dead bodies of your servants as food to the birds of the air, the flesh of your saints to the beasts of the earth.
PS|79|3|They have poured out blood like water all around Jerusalem, and there is no one to bury the dead.
PS|79|4|We are objects of reproach to our neighbors, of scorn and derision to those around us.
PS|79|5|How long, O LORD? Will you be angry forever? How long will your jealousy burn like fire?
PS|79|6|Pour out your wrath on the nations that do not acknowledge you, on the kingdoms that do not call on your name;
PS|79|7|for they have devoured Jacob and destroyed his homeland.
PS|79|8|Do not hold against us the sins of the fathers; may your mercy come quickly to meet us, for we are in desperate need.
PS|79|9|Help us, O God our Savior, for the glory of your name; deliver us and forgive our sins for your name's sake.
PS|79|10|Why should the nations say, "Where is their God?" Before our eyes, make known among the nations that you avenge the outpoured blood of your servants.
PS|79|11|May the groans of the prisoners come before you; by the strength of your arm preserve those condemned to die.
PS|79|12|Pay back into the laps of our neighbors seven times the reproach they have hurled at you, O Lord.
PS|79|13|Then we your people, the sheep of your pasture, will praise you forever; from generation to generation we will recount your praise.
PS|80|1|Hear us, O Shepherd of Israel, you who lead Joseph like a flock; you who sit enthroned between the cherubim, shine forth
PS|80|2|before Ephraim, Benjamin and Manasseh. Awaken your might; come and save us.
PS|80|3|Restore us, O God; make your face shine upon us, that we may be saved.
PS|80|4|O LORD God Almighty, how long will your anger smolder against the prayers of your people?
PS|80|5|You have fed them with the bread of tears; you have made them drink tears by the bowlful.
PS|80|6|You have made us a source of contention to our neighbors, and our enemies mock us.
PS|80|7|Restore us, O God Almighty; make your face shine upon us, that we may be saved.
PS|80|8|You brought a vine out of Egypt; you drove out the nations and planted it.
PS|80|9|You cleared the ground for it, and it took root and filled the land.
PS|80|10|The mountains were covered with its shade, the mighty cedars with its branches.
PS|80|11|It sent out its boughs to the Sea, its shoots as far as the River.
PS|80|12|Why have you broken down its walls so that all who pass by pick its grapes?
PS|80|13|Boars from the forest ravage it and the creatures of the field feed on it.
PS|80|14|Return to us, O God Almighty! Look down from heaven and see! Watch over this vine,
PS|80|15|the root your right hand has planted, the son you have raised up for yourself.
PS|80|16|Your vine is cut down, it is burned with fire; at your rebuke your people perish.
PS|80|17|Let your hand rest on the man at your right hand, the son of man you have raised up for yourself.
PS|80|18|Then we will not turn away from you; revive us, and we will call on your name.
PS|80|19|Restore us, O LORD God Almighty; make your face shine upon us, that we may be saved.
PS|81|1|Sing for joy to God our strength; shout aloud to the God of Jacob!
PS|81|2|Begin the music, strike the tambourine, play the melodious harp and lyre.
PS|81|3|Sound the ram's horn at the New Moon, and when the moon is full, on the day of our Feast;
PS|81|4|this is a decree for Israel, an ordinance of the God of Jacob.
PS|81|5|He established it as a statute for Joseph when he went out against Egypt, where we heard a language we did not understand.
PS|81|6|He says, "I removed the burden from their shoulders; their hands were set free from the basket.
PS|81|7|In your distress you called and I rescued you, I answered you out of a thundercloud; I tested you at the waters of Meribah. Selah
PS|81|8|"Hear, O my people, and I will warn you- if you would but listen to me, O Israel!
PS|81|9|You shall have no foreign god among you; you shall not bow down to an alien god.
PS|81|10|I am the LORD your God, who brought you up out of Egypt. Open wide your mouth and I will fill it.
PS|81|11|"But my people would not listen to me; Israel would not submit to me.
PS|81|12|So I gave them over to their stubborn hearts to follow their own devices.
PS|81|13|"If my people would but listen to me, if Israel would follow my ways,
PS|81|14|how quickly would I subdue their enemies and turn my hand against their foes!
PS|81|15|Those who hate the LORD would cringe before him, and their punishment would last forever.
PS|81|16|But you would be fed with the finest of wheat; with honey from the rock I would satisfy you."
PS|82|1|God presides in the great assembly; he gives judgment among the "gods":
PS|82|2|"How long will you defend the unjust and show partiality to the wicked? Selah
PS|82|3|Defend the cause of the weak and fatherless; maintain the rights of the poor and oppressed.
PS|82|4|Rescue the weak and needy; deliver them from the hand of the wicked.
PS|82|5|"They know nothing, they understand nothing. They walk about in darkness; all the foundations of the earth are shaken.
PS|82|6|"I said, 'You are "gods"; you are all sons of the Most High.'
PS|82|7|But you will die like mere men; you will fall like every other ruler."
PS|82|8|Rise up, O God, judge the earth, for all the nations are your inheritance.
PS|83|1|O God, do not keep silent; be not quiet, O God, be not still.
PS|83|2|See how your enemies are astir, how your foes rear their heads.
PS|83|3|With cunning they conspire against your people; they plot against those you cherish.
PS|83|4|"Come," they say, "let us destroy them as a nation, that the name of Israel be remembered no more."
PS|83|5|With one mind they plot together; they form an alliance against you-
PS|83|6|the tents of Edom and the Ishmaelites, of Moab and the Hagrites,
PS|83|7|Gebal, Ammon and Amalek, Philistia, with the people of Tyre.
PS|83|8|Even Assyria has joined them to lend strength to the descendants of Lot. Selah
PS|83|9|Do to them as you did to Midian, as you did to Sisera and Jabin at the river Kishon,
PS|83|10|who perished at Endor and became like refuse on the ground.
PS|83|11|Make their nobles like Oreb and Zeeb, all their princes like Zebah and Zalmunna,
PS|83|12|who said, "Let us take possession of the pasturelands of God."
PS|83|13|Make them like tumbleweed, O my God, like chaff before the wind.
PS|83|14|As fire consumes the forest or a flame sets the mountains ablaze,
PS|83|15|so pursue them with your tempest and terrify them with your storm.
PS|83|16|Cover their faces with shame so that men will seek your name, O LORD.
PS|83|17|May they ever be ashamed and dismayed; may they perish in disgrace.
PS|83|18|Let them know that you, whose name is the LORD - that you alone are the Most High over all the earth.
PS|84|1|How lovely is your dwelling place, O LORD Almighty!
PS|84|2|My soul yearns, even faints, for the courts of the LORD; my heart and my flesh cry out for the living God.
PS|84|3|Even the sparrow has found a home, and the swallow a nest for herself, where she may have her young- a place near your altar, O LORD Almighty, my King and my God.
PS|84|4|Blessed are those who dwell in your house; they are ever praising you. Selah
PS|84|5|Blessed are those whose strength is in you, who have set their hearts on pilgrimage.
PS|84|6|As they pass through the Valley of Baca, they make it a place of springs; the autumn rains also cover it with pools.
PS|84|7|They go from strength to strength, till each appears before God in Zion.
PS|84|8|Hear my prayer, O LORD God Almighty; listen to me, O God of Jacob. Selah
PS|84|9|Look upon our shield, O God; look with favor on your anointed one.
PS|84|10|Better is one day in your courts than a thousand elsewhere; I would rather be a doorkeeper in the house of my God than dwell in the tents of the wicked.
PS|84|11|For the LORD God is a sun and shield; the LORD bestows favor and honor; no good thing does he withhold from those whose walk is blameless.
PS|84|12|O LORD Almighty, blessed is the man who trusts in you.
PS|85|1|You showed favor to your land, O LORD; you restored the fortunes of Jacob.
PS|85|2|You forgave the iniquity of your people and covered all their sins. Selah
PS|85|3|You set aside all your wrath and turned from your fierce anger.
PS|85|4|Restore us again, O God our Savior, and put away your displeasure toward us.
PS|85|5|Will you be angry with us forever? Will you prolong your anger through all generations?
PS|85|6|Will you not revive us again, that your people may rejoice in you?
PS|85|7|Show us your unfailing love, O LORD, and grant us your salvation.
PS|85|8|I will listen to what God the LORD will say; he promises peace to his people, his saints- but let them not return to folly.
PS|85|9|Surely his salvation is near those who fear him, that his glory may dwell in our land.
PS|85|10|Love and faithfulness meet together; righteousness and peace kiss each other.
PS|85|11|Faithfulness springs forth from the earth, and righteousness looks down from heaven.
PS|85|12|The LORD will indeed give what is good, and our land will yield its harvest.
PS|85|13|Righteousness goes before him and prepares the way for his steps.
PS|86|1|Hear, O LORD, and answer me, for I am poor and needy.
PS|86|2|Guard my life, for I am devoted to you. You are my God; save your servant who trusts in you.
PS|86|3|Have mercy on me, O Lord, for I call to you all day long.
PS|86|4|Bring joy to your servant, for to you, O Lord, I lift up my soul.
PS|86|5|You are forgiving and good, O Lord, abounding in love to all who call to you.
PS|86|6|Hear my prayer, O LORD; listen to my cry for mercy.
PS|86|7|In the day of my trouble I will call to you, for you will answer me.
PS|86|8|Among the gods there is none like you, O Lord; no deeds can compare with yours.
PS|86|9|All the nations you have made will come and worship before you, O Lord; they will bring glory to your name.
PS|86|10|For you are great and do marvelous deeds; you alone are God.
PS|86|11|Teach me your way, O LORD, and I will walk in your truth; give me an undivided heart, that I may fear your name.
PS|86|12|I will praise you, O Lord my God, with all my heart; I will glorify your name forever.
PS|86|13|For great is your love toward me; you have delivered me from the depths of the grave.
PS|86|14|The arrogant are attacking me, O God; a band of ruthless men seeks my life- men without regard for you.
PS|86|15|But you, O Lord, are a compassionate and gracious God, slow to anger, abounding in love and faithfulness.
PS|86|16|Turn to me and have mercy on me; grant your strength to your servant and save the son of your maidservant.
PS|86|17|Give me a sign of your goodness, that my enemies may see it and be put to shame, for you, O LORD, have helped me and comforted me.
PS|87|1|He has set his foundation on the holy mountain;
PS|87|2|the LORD loves the gates of Zion more than all the dwellings of Jacob.
PS|87|3|Glorious things are said of you, O city of God: Selah
PS|87|4|"I will record Rahab and Babylon among those who acknowledge me- Philistia too, and Tyre, along with Cush - and will say, 'This one was born in Zion.'"
PS|87|5|Indeed, of Zion it will be said, "This one and that one were born in her, and the Most High himself will establish her."
PS|87|6|The LORD will write in the register of the peoples: "This one was born in Zion." Selah
PS|87|7|As they make music they will sing, "All my fountains are in you."
PS|88|1|O LORD, the God who saves me, day and night I cry out before you.
PS|88|2|May my prayer come before you; turn your ear to my cry.
PS|88|3|For my soul is full of trouble and my life draws near the grave.
PS|88|4|I am counted among those who go down to the pit; I am like a man without strength.
PS|88|5|I am set apart with the dead, like the slain who lie in the grave, whom you remember no more, who are cut off from your care.
PS|88|6|You have put me in the lowest pit, in the darkest depths.
PS|88|7|Your wrath lies heavily upon me; you have overwhelmed me with all your waves. Selah
PS|88|8|You have taken from me my closest friends and have made me repulsive to them. I am confined and cannot escape;
PS|88|9|my eyes are dim with grief. I call to you, O LORD, every day; I spread out my hands to you.
PS|88|10|Do you show your wonders to the dead? Do those who are dead rise up and praise you? Selah
PS|88|11|Is your love declared in the grave, your faithfulness in Destruction?
PS|88|12|Are your wonders known in the place of darkness, or your righteous deeds in the land of oblivion?
PS|88|13|But I cry to you for help, O LORD; in the morning my prayer comes before you.
PS|88|14|Why, O LORD, do you reject me and hide your face from me?
PS|88|15|From my youth I have been afflicted and close to death; I have suffered your terrors and am in despair.
PS|88|16|Your wrath has swept over me; your terrors have destroyed me.
PS|88|17|All day long they surround me like a flood; they have completely engulfed me.
PS|88|18|You have taken my companions and loved ones from me; the darkness is my closest friend.
PS|89|1|I will sing of the LORD's great love forever; with my mouth I will make your faithfulness known through all generations.
PS|89|2|I will declare that your love stands firm forever, that you established your faithfulness in heaven itself.
PS|89|3|You said, "I have made a covenant with my chosen one, I have sworn to David my servant,
PS|89|4|'I will establish your line forever and make your throne firm through all generations.'" Selah
PS|89|5|The heavens praise your wonders, O LORD, your faithfulness too, in the assembly of the holy ones.
PS|89|6|For who in the skies above can compare with the LORD? Who is like the LORD among the heavenly beings?
PS|89|7|In the council of the holy ones God is greatly feared; he is more awesome than all who surround him.
PS|89|8|O LORD God Almighty, who is like you? You are mighty, O LORD, and your faithfulness surrounds you.
PS|89|9|You rule over the surging sea; when its waves mount up, you still them.
PS|89|10|You crushed Rahab like one of the slain; with your strong arm you scattered your enemies.
PS|89|11|The heavens are yours, and yours also the earth; you founded the world and all that is in it.
PS|89|12|You created the north and the south; Tabor and Hermon sing for joy at your name.
PS|89|13|Your arm is endued with power; your hand is strong, your right hand exalted.
PS|89|14|Righteousness and justice are the foundation of your throne; love and faithfulness go before you.
PS|89|15|Blessed are those who have learned to acclaim you, who walk in the light of your presence, O LORD.
PS|89|16|They rejoice in your name all day long; they exult in your righteousness.
PS|89|17|For you are their glory and strength, and by your favor you exalt our horn.
PS|89|18|Indeed, our shield belongs to the LORD, our king to the Holy One of Israel.
PS|89|19|Once you spoke in a vision, to your faithful people you said: "I have bestowed strength on a warrior; I have exalted a young man from among the people.
PS|89|20|I have found David my servant; with my sacred oil I have anointed him.
PS|89|21|My hand will sustain him; surely my arm will strengthen him.
PS|89|22|No enemy will subject him to tribute; no wicked man will oppress him.
PS|89|23|I will crush his foes before him and strike down his adversaries.
PS|89|24|My faithful love will be with him, and through my name his horn will be exalted.
PS|89|25|I will set his hand over the sea, his right hand over the rivers.
PS|89|26|He will call out to me, 'You are my Father, my God, the Rock my Savior.'
PS|89|27|I will also appoint him my firstborn, the most exalted of the kings of the earth.
PS|89|28|I will maintain my love to him forever, and my covenant with him will never fail.
PS|89|29|I will establish his line forever, his throne as long as the heavens endure.
PS|89|30|"If his sons forsake my law and do not follow my statutes,
PS|89|31|if they violate my decrees and fail to keep my commands,
PS|89|32|I will punish their sin with the rod, their iniquity with flogging;
PS|89|33|but I will not take my love from him, nor will I ever betray my faithfulness.
PS|89|34|I will not violate my covenant or alter what my lips have uttered.
PS|89|35|Once for all, I have sworn by my holiness- and I will not lie to David-
PS|89|36|that his line will continue forever and his throne endure before me like the sun;
PS|89|37|it will be established forever like the moon, the faithful witness in the sky." Selah
PS|89|38|But you have rejected, you have spurned, you have been very angry with your anointed one.
PS|89|39|You have renounced the covenant with your servant and have defiled his crown in the dust.
PS|89|40|You have broken through all his walls and reduced his strongholds to ruins.
PS|89|41|All who pass by have plundered him; he has become the scorn of his neighbors.
PS|89|42|You have exalted the right hand of his foes; you have made all his enemies rejoice.
PS|89|43|You have turned back the edge of his sword and have not supported him in battle.
PS|89|44|You have put an end to his splendor and cast his throne to the ground.
PS|89|45|You have cut short the days of his youth; you have covered him with a mantle of shame. Selah
PS|89|46|How long, O LORD? Will you hide yourself forever? How long will your wrath burn like fire?
PS|89|47|Remember how fleeting is my life. For what futility you have created all men!
PS|89|48|What man can live and not see death, or save himself from the power of the grave? Selah
PS|89|49|O Lord, where is your former great love, which in your faithfulness you swore to David?
PS|89|50|Remember, Lord, how your servant has been mocked, how I bear in my heart the taunts of all the nations,
PS|89|51|the taunts with which your enemies have mocked, O LORD, with which they have mocked every step of your anointed one.
PS|89|52|Praise be to the LORD forever! Amen and Amen. BOOK IV Psalms 90-106
PS|90|1|Lord, you have been our dwelling place throughout all generations.
PS|90|2|Before the mountains were born or you brought forth the earth and the world, from everlasting to everlasting you are God.
PS|90|3|You turn men back to dust, saying, "Return to dust, O sons of men."
PS|90|4|For a thousand years in your sight are like a day that has just gone by, or like a watch in the night.
PS|90|5|You sweep men away in the sleep of death; they are like the new grass of the morning-
PS|90|6|though in the morning it springs up new, by evening it is dry and withered.
PS|90|7|We are consumed by your anger and terrified by your indignation.
PS|90|8|You have set our iniquities before you, our secret sins in the light of your presence.
PS|90|9|All our days pass away under your wrath; we finish our years with a moan.
PS|90|10|The length of our days is seventy years- or eighty, if we have the strength; yet their span is but trouble and sorrow, for they quickly pass, and we fly away.
PS|90|11|Who knows the power of your anger? For your wrath is as great as the fear that is due you.
PS|90|12|Teach us to number our days aright, that we may gain a heart of wisdom.
PS|90|13|Relent, O LORD! How long will it be? Have compassion on your servants.
PS|90|14|Satisfy us in the morning with your unfailing love, that we may sing for joy and be glad all our days.
PS|90|15|Make us glad for as many days as you have afflicted us, for as many years as we have seen trouble.
PS|90|16|May your deeds be shown to your servants, your splendor to their children.
PS|90|17|May the favor of the Lord our God rest upon us; establish the work of our hands for us- yes, establish the work of our hands.
PS|91|1|He who dwells in the shelter of the Most High will rest in the shadow of the Almighty.
PS|91|2|I will say of the LORD, "He is my refuge and my fortress, my God, in whom I trust."
PS|91|3|Surely he will save you from the fowler's snare and from the deadly pestilence.
PS|91|4|He will cover you with his feathers, and under his wings you will find refuge; his faithfulness will be your shield and rampart.
PS|91|5|You will not fear the terror of night, nor the arrow that flies by day,
PS|91|6|nor the pestilence that stalks in the darkness, nor the plague that destroys at midday.
PS|91|7|A thousand may fall at your side, ten thousand at your right hand, but it will not come near you.
PS|91|8|You will only observe with your eyes and see the punishment of the wicked.
PS|91|9|If you make the Most High your dwelling- even the LORD, who is my refuge-
PS|91|10|then no harm will befall you, no disaster will come near your tent.
PS|91|11|For he will command his angels concerning you to guard you in all your ways;
PS|91|12|they will lift you up in their hands, so that you will not strike your foot against a stone.
PS|91|13|You will tread upon the lion and the cobra; you will trample the great lion and the serpent.
PS|91|14|"Because he loves me," says the LORD, "I will rescue him; I will protect him, for he acknowledges my name.
PS|91|15|He will call upon me, and I will answer him; I will be with him in trouble, I will deliver him and honor him.
PS|91|16|With long life will I satisfy him and show him my salvation."
PS|92|1|It is good to praise the LORD and make music to your name, O Most High,
PS|92|2|to proclaim your love in the morning and your faithfulness at night,
PS|92|3|to the music of the ten-stringed lyre and the melody of the harp.
PS|92|4|For you make me glad by your deeds, O LORD; I sing for joy at the works of your hands.
PS|92|5|How great are your works, O LORD, how profound your thoughts!
PS|92|6|The senseless man does not know, fools do not understand,
PS|92|7|that though the wicked spring up like grass and all evildoers flourish, they will be forever destroyed.
PS|92|8|But you, O LORD, are exalted forever.
PS|92|9|For surely your enemies, O LORD, surely your enemies will perish; all evildoers will be scattered.
PS|92|10|You have exalted my horn like that of a wild ox; fine oils have been poured upon me.
PS|92|11|My eyes have seen the defeat of my adversaries; my ears have heard the rout of my wicked foes.
PS|92|12|The righteous will flourish like a palm tree, they will grow like a cedar of Lebanon;
PS|92|13|planted in the house of the LORD, they will flourish in the courts of our God.
PS|92|14|They will still bear fruit in old age, they will stay fresh and green,
PS|92|15|proclaiming, "The LORD is upright; he is my Rock, and there is no wickedness in him."
PS|93|1|The LORD reigns, he is robed in majesty; the LORD is robed in majesty and is armed with strength. The world is firmly established; it cannot be moved.
PS|93|2|Your throne was established long ago; you are from all eternity.
PS|93|3|The seas have lifted up, O LORD, the seas have lifted up their voice; the seas have lifted up their pounding waves.
PS|93|4|Mightier than the thunder of the great waters, mightier than the breakers of the sea- the LORD on high is mighty.
PS|93|5|Your statutes stand firm; holiness adorns your house for endless days, O LORD.
PS|94|1|O LORD, the God who avenges, O God who avenges, shine forth.
PS|94|2|Rise up, O Judge of the earth; pay back to the proud what they deserve.
PS|94|3|How long will the wicked, O LORD, how long will the wicked be jubilant?
PS|94|4|They pour out arrogant words; all the evildoers are full of boasting.
PS|94|5|They crush your people, O LORD; they oppress your inheritance.
PS|94|6|They slay the widow and the alien; they murder the fatherless.
PS|94|7|They say, "The LORD does not see; the God of Jacob pays no heed."
PS|94|8|Take heed, you senseless ones among the people; you fools, when will you become wise?
PS|94|9|Does he who implanted the ear not hear? Does he who formed the eye not see?
PS|94|10|Does he who disciplines nations not punish? Does he who teaches man lack knowledge?
PS|94|11|The LORD knows the thoughts of man; he knows that they are futile.
PS|94|12|Blessed is the man you discipline, O LORD, the man you teach from your law;
PS|94|13|you grant him relief from days of trouble, till a pit is dug for the wicked.
PS|94|14|For the LORD will not reject his people; he will never forsake his inheritance.
PS|94|15|Judgment will again be founded on righteousness, and all the upright in heart will follow it.
PS|94|16|Who will rise up for me against the wicked? Who will take a stand for me against evildoers?
PS|94|17|Unless the LORD had given me help, I would soon have dwelt in the silence of death.
PS|94|18|When I said, "My foot is slipping," your love, O LORD, supported me.
PS|94|19|When anxiety was great within me, your consolation brought joy to my soul.
PS|94|20|Can a corrupt throne be allied with you- one that brings on misery by its decrees?
PS|94|21|They band together against the righteous and condemn the innocent to death.
PS|94|22|But the LORD has become my fortress, and my God the rock in whom I take refuge.
PS|94|23|He will repay them for their sins and destroy them for their wickedness; the LORD our God will destroy them.
PS|95|1|Come, let us sing for joy to the LORD; let us shout aloud to the Rock of our salvation.
PS|95|2|Let us come before him with thanksgiving and extol him with music and song.
PS|95|3|For the LORD is the great God, the great King above all gods.
PS|95|4|In his hand are the depths of the earth, and the mountain peaks belong to him.
PS|95|5|The sea is his, for he made it, and his hands formed the dry land.
PS|95|6|Come, let us bow down in worship, let us kneel before the LORD our Maker;
PS|95|7|for he is our God and we are the people of his pasture, the flock under his care. Today, if you hear his voice,
PS|95|8|do not harden your hearts as you did at Meribah, as you did that day at Massah in the desert,
PS|95|9|where your fathers tested and tried me, though they had seen what I did.
PS|95|10|For forty years I was angry with that generation; I said, "They are a people whose hearts go astray, and they have not known my ways."
PS|95|11|So I declared on oath in my anger, "They shall never enter my rest."
PS|96|1|Sing to the LORD a new song; sing to the LORD, all the earth.
PS|96|2|Sing to the LORD, praise his name; proclaim his salvation day after day.
PS|96|3|Declare his glory among the nations, his marvelous deeds among all peoples.
PS|96|4|For great is the LORD and most worthy of praise; he is to be feared above all gods.
PS|96|5|For all the gods of the nations are idols, but the LORD made the heavens.
PS|96|6|Splendor and majesty are before him; strength and glory are in his sanctuary.
PS|96|7|Ascribe to the LORD, O families of nations, ascribe to the LORD glory and strength.
PS|96|8|Ascribe to the LORD the glory due his name; bring an offering and come into his courts.
PS|96|9|Worship the LORD in the splendor of his holiness; tremble before him, all the earth.
PS|96|10|Say among the nations, "The LORD reigns." The world is firmly established, it cannot be moved; he will judge the peoples with equity.
PS|96|11|Let the heavens rejoice, let the earth be glad; let the sea resound, and all that is in it;
PS|96|12|let the fields be jubilant, and everything in them. Then all the trees of the forest will sing for joy;
PS|96|13|they will sing before the LORD, for he comes, he comes to judge the earth. He will judge the world in righteousness and the peoples in his truth.
PS|97|1|The LORD reigns, let the earth be glad; let the distant shores rejoice.
PS|97|2|Clouds and thick darkness surround him; righteousness and justice are the foundation of his throne.
PS|97|3|Fire goes before him and consumes his foes on every side.
PS|97|4|His lightning lights up the world; the earth sees and trembles.
PS|97|5|The mountains melt like wax before the LORD, before the Lord of all the earth.
PS|97|6|The heavens proclaim his righteousness, and all the peoples see his glory.
PS|97|7|All who worship images are put to shame, those who boast in idols- worship him, all you gods!
PS|97|8|Zion hears and rejoices and the villages of Judah are glad because of your judgments, O LORD.
PS|97|9|For you, O LORD, are the Most High over all the earth; you are exalted far above all gods.
PS|97|10|Let those who love the LORD hate evil, for he guards the lives of his faithful ones and delivers them from the hand of the wicked.
PS|97|11|Light is shed upon the righteous and joy on the upright in heart.
PS|97|12|Rejoice in the LORD, you who are righteous, and praise his holy name.
PS|98|1|Sing to the LORD a new song, for he has done marvelous things; his right hand and his holy arm have worked salvation for him.
PS|98|2|The LORD has made his salvation known and revealed his righteousness to the nations.
PS|98|3|He has remembered his love and his faithfulness to the house of Israel; all the ends of the earth have seen the salvation of our God.
PS|98|4|Shout for joy to the LORD, all the earth, burst into jubilant song with music;
PS|98|5|make music to the LORD with the harp, with the harp and the sound of singing,
PS|98|6|with trumpets and the blast of the ram's horn- shout for joy before the LORD, the King.
PS|98|7|Let the sea resound, and everything in it, the world, and all who live in it.
PS|98|8|Let the rivers clap their hands, Let the mountains sing together for joy;
PS|98|9|let them sing before the LORD, for he comes to judge the earth. He will judge the world in righteousness and the peoples with equity.
PS|99|1|The LORD reigns, let the nations tremble; he sits enthroned between the cherubim, let the earth shake.
PS|99|2|Great is the LORD in Zion; he is exalted over all the nations.
PS|99|3|Let them praise your great and awesome name- he is holy.
PS|99|4|The King is mighty, he loves justice- you have established equity; in Jacob you have done what is just and right.
PS|99|5|Exalt the LORD our God and worship at his footstool; he is holy.
PS|99|6|Moses and Aaron were among his priests, Samuel was among those who called on his name; they called on the LORD and he answered them.
PS|99|7|He spoke to them from the pillar of cloud; they kept his statutes and the decrees he gave them.
PS|99|8|O LORD our God, you answered them; you were to Israel a forgiving God, though you punished their misdeeds.
PS|99|9|Exalt the LORD our God and worship at his holy mountain, for the LORD our God is holy.
PS|100|1|Shout for joy to the LORD, all the earth.
PS|100|2|Worship the LORD with gladness; come before him with joyful songs.
PS|100|3|Know that the LORD is God. It is he who made us, and we are his; we are his people, the sheep of his pasture.
PS|100|4|Enter his gates with thanksgiving and his courts with praise; give thanks to him and praise his name.
PS|100|5|For the LORD is good and his love endures forever; his faithfulness continues through all generations.
PS|101|1|I will sing of your love and justice; to you, O LORD, I will sing praise.
PS|101|2|I will be careful to lead a blameless life- when will you come to me? I will walk in my house with blameless heart.
PS|101|3|I will set before my eyes no vile thing. The deeds of faithless men I hate; they will not cling to me.
PS|101|4|Men of perverse heart shall be far from me; I will have nothing to do with evil.
PS|101|5|Whoever slanders his neighbor in secret, him will I put to silence; whoever has haughty eyes and a proud heart, him will I not endure.
PS|101|6|My eyes will be on the faithful in the land, that they may dwell with me; he whose walk is blameless will minister to me.
PS|101|7|No one who practices deceit will dwell in my house; no one who speaks falsely will stand in my presence.
PS|101|8|Every morning I will put to silence all the wicked in the land; I will cut off every evildoer from the city of the LORD.
PS|102|1|Hear my prayer, O LORD; let my cry for help come to you.
PS|102|2|Do not hide your face from me when I am in distress. Turn your ear to me; when I call, answer me quickly.
PS|102|3|For my days vanish like smoke; my bones burn like glowing embers.
PS|102|4|My heart is blighted and withered like grass; I forget to eat my food.
PS|102|5|Because of my loud groaning I am reduced to skin and bones.
PS|102|6|I am like a desert owl, like an owl among the ruins.
PS|102|7|I lie awake; I have become like a bird alone on a roof.
PS|102|8|All day long my enemies taunt me; those who rail against me use my name as a curse.
PS|102|9|For I eat ashes as my food and mingle my drink with tears
PS|102|10|because of your great wrath, for you have taken me up and thrown me aside.
PS|102|11|My days are like the evening shadow; I wither away like grass.
PS|102|12|But you, O LORD, sit enthroned forever; your renown endures through all generations.
PS|102|13|You will arise and have compassion on Zion, for it is time to show favor to her; the appointed time has come.
PS|102|14|For her stones are dear to your servants; her very dust moves them to pity.
PS|102|15|The nations will fear the name of the LORD, all the kings of the earth will revere your glory.
PS|102|16|For the LORD will rebuild Zion and appear in his glory.
PS|102|17|He will respond to the prayer of the destitute; he will not despise their plea.
PS|102|18|Let this be written for a future generation, that a people not yet created may praise the LORD:
PS|102|19|"The LORD looked down from his sanctuary on high, from heaven he viewed the earth,
PS|102|20|to hear the groans of the prisoners and release those condemned to death."
PS|102|21|So the name of the LORD will be declared in Zion and his praise in Jerusalem
PS|102|22|when the peoples and the kingdoms assemble to worship the LORD.
PS|102|23|In the course of my life he broke my strength; he cut short my days.
PS|102|24|So I said: "Do not take me away, O my God, in the midst of my days; your years go on through all generations.
PS|102|25|In the beginning you laid the foundations of the earth, and the heavens are the work of your hands.
PS|102|26|They will perish, but you remain; they will all wear out like a garment. Like clothing you will change them and they will be discarded.
PS|102|27|But you remain the same, and your years will never end.
PS|102|28|The children of your servants will live in your presence; their descendants will be established before you."
PS|103|1|Praise the LORD, O my soul; all my inmost being, praise his holy name.
PS|103|2|Praise the LORD, O my soul, and forget not all his benefits-
PS|103|3|who forgives all your sins and heals all your diseases,
PS|103|4|who redeems your life from the pit and crowns you with love and compassion,
PS|103|5|who satisfies your desires with good things so that your youth is renewed like the eagle's.
PS|103|6|The LORD works righteousness and justice for all the oppressed.
PS|103|7|He made known his ways to Moses, his deeds to the people of Israel:
PS|103|8|The LORD is compassionate and gracious, slow to anger, abounding in love.
PS|103|9|He will not always accuse, nor will he harbor his anger forever;
PS|103|10|he does not treat us as our sins deserve or repay us according to our iniquities.
PS|103|11|For as high as the heavens are above the earth, so great is his love for those who fear him;
PS|103|12|as far as the east is from the west, so far has he removed our transgressions from us.
PS|103|13|As a father has compassion on his children, so the LORD has compassion on those who fear him;
PS|103|14|for he knows how we are formed, he remembers that we are dust.
PS|103|15|As for man, his days are like grass, he flourishes like a flower of the field;
PS|103|16|the wind blows over it and it is gone, and its place remembers it no more.
PS|103|17|But from everlasting to everlasting the LORD's love is with those who fear him, and his righteousness with their children's children-
PS|103|18|with those who keep his covenant and remember to obey his precepts.
PS|103|19|The LORD has established his throne in heaven, and his kingdom rules over all.
PS|103|20|Praise the LORD, you his angels, you mighty ones who do his bidding, who obey his word.
PS|103|21|Praise the LORD, all his heavenly hosts, you his servants who do his will.
PS|103|22|Praise the LORD, all his works everywhere in his dominion. Praise the LORD, O my soul.
PS|104|1|Praise the LORD, O my soul. O LORD my God, you are very great; you are clothed with splendor and majesty.
PS|104|2|He wraps himself in light as with a garment; he stretches out the heavens like a tent
PS|104|3|and lays the beams of his upper chambers on their waters. He makes the clouds his chariot and rides on the wings of the wind.
PS|104|4|He makes winds his messengers, flames of fire his servants.
PS|104|5|He set the earth on its foundations; it can never be moved.
PS|104|6|You covered it with the deep as with a garment; the waters stood above the mountains.
PS|104|7|But at your rebuke the waters fled, at the sound of your thunder they took to flight;
PS|104|8|they flowed over the mountains, they went down into the valleys, to the place you assigned for them.
PS|104|9|You set a boundary they cannot cross; never again will they cover the earth.
PS|104|10|He makes springs pour water into the ravines; it flows between the mountains.
PS|104|11|They give water to all the beasts of the field; the wild donkeys quench their thirst.
PS|104|12|The birds of the air nest by the waters; they sing among the branches.
PS|104|13|He waters the mountains from his upper chambers; the earth is satisfied by the fruit of his work.
PS|104|14|He makes grass grow for the cattle, and plants for man to cultivate- bringing forth food from the earth:
PS|104|15|wine that gladdens the heart of man, oil to make his face shine, and bread that sustains his heart.
PS|104|16|The trees of the LORD are well watered, the cedars of Lebanon that he planted.
PS|104|17|There the birds make their nests; the stork has its home in the pine trees.
PS|104|18|The high mountains belong to the wild goats; the crags are a refuge for the coneys.
PS|104|19|The moon marks off the seasons, and the sun knows when to go down.
PS|104|20|You bring darkness, it becomes night, and all the beasts of the forest prowl.
PS|104|21|The lions roar for their prey and seek their food from God.
PS|104|22|The sun rises, and they steal away; they return and lie down in their dens.
PS|104|23|Then man goes out to his work, to his labor until evening.
PS|104|24|How many are your works, O LORD! In wisdom you made them all; the earth is full of your creatures.
PS|104|25|There is the sea, vast and spacious, teeming with creatures beyond number- living things both large and small.
PS|104|26|There the ships go to and fro, and the leviathan, which you formed to frolic there.
PS|104|27|These all look to you to give them their food at the proper time.
PS|104|28|When you give it to them, they gather it up; when you open your hand, they are satisfied with good things.
PS|104|29|When you hide your face, they are terrified; when you take away their breath, they die and return to the dust.
PS|104|30|When you send your Spirit, they are created, and you renew the face of the earth.
PS|104|31|May the glory of the LORD endure forever; may the LORD rejoice in his works-
PS|104|32|he who looks at the earth, and it trembles, who touches the mountains, and they smoke.
PS|104|33|I will sing to the LORD all my life; I will sing praise to my God as long as I live.
PS|104|34|May my meditation be pleasing to him, as I rejoice in the LORD.
PS|104|35|But may sinners vanish from the earth and the wicked be no more. Praise the LORD, O my soul. Praise the LORD.
PS|105|1|Give thanks to the LORD, call on his name; make known among the nations what he has done.
PS|105|2|Sing to him, sing praise to him; tell of all his wonderful acts.
PS|105|3|Glory in his holy name; let the hearts of those who seek the LORD rejoice.
PS|105|4|Look to the LORD and his strength; seek his face always.
PS|105|5|Remember the wonders he has done, his miracles, and the judgments he pronounced,
PS|105|6|O descendants of Abraham his servant, O sons of Jacob, his chosen ones.
PS|105|7|He is the LORD our God; his judgments are in all the earth.
PS|105|8|He remembers his covenant forever, the word he commanded, for a thousand generations,
PS|105|9|the covenant he made with Abraham, the oath he swore to Isaac.
PS|105|10|He confirmed it to Jacob as a decree, to Israel as an everlasting covenant:
PS|105|11|"To you I will give the land of Canaan as the portion you will inherit."
PS|105|12|When they were but few in number, few indeed, and strangers in it,
PS|105|13|they wandered from nation to nation, from one kingdom to another.
PS|105|14|He allowed no one to oppress them; for their sake he rebuked kings:
PS|105|15|"Do not touch my anointed ones; do my prophets no harm."
PS|105|16|He called down famine on the land and destroyed all their supplies of food;
PS|105|17|and he sent a man before them- Joseph, sold as a slave.
PS|105|18|They bruised his feet with shackles, his neck was put in irons,
PS|105|19|till what he foretold came to pass, till the word of the LORD proved him true.
PS|105|20|The king sent and released him, the ruler of peoples set him free.
PS|105|21|He made him master of his household, ruler over all he possessed,
PS|105|22|to instruct his princes as he pleased and teach his elders wisdom.
PS|105|23|Then Israel entered Egypt; Jacob lived as an alien in the land of Ham.
PS|105|24|The LORD made his people very fruitful; he made them too numerous for their foes,
PS|105|25|whose hearts he turned to hate his people, to conspire against his servants.
PS|105|26|He sent Moses his servant, and Aaron, whom he had chosen.
PS|105|27|They performed his miraculous signs among them, his wonders in the land of Ham.
PS|105|28|He sent darkness and made the land dark- for had they not rebelled against his words?
PS|105|29|He turned their waters into blood, causing their fish to die.
PS|105|30|Their land teemed with frogs, which went up into the bedrooms of their rulers.
PS|105|31|He spoke, and there came swarms of flies, and gnats throughout their country.
PS|105|32|He turned their rain into hail, with lightning throughout their land;
PS|105|33|he struck down their vines and fig trees and shattered the trees of their country.
PS|105|34|He spoke, and the locusts came, grasshoppers without number;
PS|105|35|they ate up every green thing in their land, ate up the produce of their soil.
PS|105|36|Then he struck down all the firstborn in their land, the firstfruits of all their manhood.
PS|105|37|He brought out Israel, laden with silver and gold, and from among their tribes no one faltered.
PS|105|38|Egypt was glad when they left, because dread of Israel had fallen on them.
PS|105|39|He spread out a cloud as a covering, and a fire to give light at night.
PS|105|40|They asked, and he brought them quail and satisfied them with the bread of heaven.
PS|105|41|He opened the rock, and water gushed out; like a river it flowed in the desert.
PS|105|42|For he remembered his holy promise given to his servant Abraham.
PS|105|43|He brought out his people with rejoicing, his chosen ones with shouts of joy;
PS|105|44|he gave them the lands of the nations, and they fell heir to what others had toiled for-
PS|105|45|that they might keep his precepts and observe his laws. Praise the LORD.
PS|106|1|Praise the LORD. Give thanks to the LORD, for he is good; his love endures forever.
PS|106|2|Who can proclaim the mighty acts of the LORD or fully declare his praise?
PS|106|3|Blessed are they who maintain justice, who constantly do what is right.
PS|106|4|Remember me, O LORD, when you show favor to your people, come to my aid when you save them,
PS|106|5|that I may enjoy the prosperity of your chosen ones, that I may share in the joy of your nation and join your inheritance in giving praise.
PS|106|6|We have sinned, even as our fathers did; we have done wrong and acted wickedly.
PS|106|7|When our fathers were in Egypt, they gave no thought to your miracles; they did not remember your many kindnesses, and they rebelled by the sea, the Red Sea.
PS|106|8|Yet he saved them for his name's sake, to make his mighty power known.
PS|106|9|He rebuked the Red Sea, and it dried up; he led them through the depths as through a desert.
PS|106|10|He saved them from the hand of the foe; from the hand of the enemy he redeemed them.
PS|106|11|The waters covered their adversaries; not one of them survived.
PS|106|12|Then they believed his promises and sang his praise.
PS|106|13|But they soon forgot what he had done and did not wait for his counsel.
PS|106|14|In the desert they gave in to their craving; in the wasteland they put God to the test.
PS|106|15|So he gave them what they asked for, but sent a wasting disease upon them.
PS|106|16|In the camp they grew envious of Moses and of Aaron, who was consecrated to the LORD.
PS|106|17|The earth opened up and swallowed Dathan; it buried the company of Abiram.
PS|106|18|Fire blazed among their followers; a flame consumed the wicked.
PS|106|19|At Horeb they made a calf and worshiped an idol cast from metal.
PS|106|20|They exchanged their Glory for an image of a bull, which eats grass.
PS|106|21|They forgot the God who saved them, who had done great things in Egypt,
PS|106|22|miracles in the land of Ham and awesome deeds by the Red Sea.
PS|106|23|So he said he would destroy them- had not Moses, his chosen one, stood in the breach before him to keep his wrath from destroying them.
PS|106|24|Then they despised the pleasant land; they did not believe his promise.
PS|106|25|They grumbled in their tents and did not obey the LORD.
PS|106|26|So he swore to them with uplifted hand that he would make them fall in the desert,
PS|106|27|make their descendants fall among the nations and scatter them throughout the lands.
PS|106|28|They yoked themselves to the Baal of Peor and ate sacrifices offered to lifeless gods;
PS|106|29|they provoked the LORD to anger by their wicked deeds, and a plague broke out among them.
PS|106|30|But Phinehas stood up and intervened, and the plague was checked.
PS|106|31|This was credited to him as righteousness for endless generations to come.
PS|106|32|By the waters of Meribah they angered the LORD, and trouble came to Moses because of them;
PS|106|33|for they rebelled against the Spirit of God, and rash words came from Moses' lips.
PS|106|34|They did not destroy the peoples as the LORD had commanded them,
PS|106|35|but they mingled with the nations and adopted their customs.
PS|106|36|They worshiped their idols, which became a snare to them.
PS|106|37|They sacrificed their sons and their daughters to demons.
PS|106|38|They shed innocent blood, the blood of their sons and daughters, whom they sacrificed to the idols of Canaan, and the land was desecrated by their blood.
PS|106|39|They defiled themselves by what they did; by their deeds they prostituted themselves.
PS|106|40|Therefore the LORD was angry with his people and abhorred his inheritance.
PS|106|41|He handed them over to the nations, and their foes ruled over them.
PS|106|42|Their enemies oppressed them and subjected them to their power.
PS|106|43|Many times he delivered them, but they were bent on rebellion and they wasted away in their sin.
PS|106|44|But he took note of their distress when he heard their cry;
PS|106|45|for their sake he remembered his covenant and out of his great love he relented.
PS|106|46|He caused them to be pitied by all who held them captive.
PS|106|47|Save us, O LORD our God, and gather us from the nations, that we may give thanks to your holy name and glory in your praise.
PS|106|48|Praise be to the LORD, the God of Israel, from everlasting to everlasting. Let all the people say, "Amen!" Praise the LORD.
PS|107|1|Give thanks to the LORD, for he is good; his love endures forever.
PS|107|2|Let the redeemed of the LORD say this- those he redeemed from the hand of the foe,
PS|107|3|those he gathered from the lands, from east and west, from north and south.
PS|107|4|Some wandered in desert wastelands, finding no way to a city where they could settle.
PS|107|5|They were hungry and thirsty, and their lives ebbed away.
PS|107|6|Then they cried out to the LORD in their trouble, and he delivered them from their distress.
PS|107|7|He led them by a straight way to a city where they could settle.
PS|107|8|Let them give thanks to the LORD for his unfailing love and his wonderful deeds for men,
PS|107|9|for he satisfies the thirsty and fills the hungry with good things.
PS|107|10|Some sat in darkness and the deepest gloom, prisoners suffering in iron chains,
PS|107|11|for they had rebelled against the words of God and despised the counsel of the Most High.
PS|107|12|So he subjected them to bitter labor; they stumbled, and there was no one to help.
PS|107|13|Then they cried to the LORD in their trouble, and he saved them from their distress.
PS|107|14|He brought them out of darkness and the deepest gloom and broke away their chains.
PS|107|15|Let them give thanks to the LORD for his unfailing love and his wonderful deeds for men,
PS|107|16|for he breaks down gates of bronze and cuts through bars of iron.
PS|107|17|Some became fools through their rebellious ways and suffered affliction because of their iniquities.
PS|107|18|They loathed all food and drew near the gates of death.
PS|107|19|Then they cried to the LORD in their trouble, and he saved them from their distress.
PS|107|20|He sent forth his word and healed them; he rescued them from the grave.
PS|107|21|Let them give thanks to the LORD for his unfailing love and his wonderful deeds for men.
PS|107|22|Let them sacrifice thank offerings and tell of his works with songs of joy.
PS|107|23|Others went out on the sea in ships; they were merchants on the mighty waters.
PS|107|24|They saw the works of the LORD, his wonderful deeds in the deep.
PS|107|25|For he spoke and stirred up a tempest that lifted high the waves.
PS|107|26|They mounted up to the heavens and went down to the depths; in their peril their courage melted away.
PS|107|27|They reeled and staggered like drunken men; they were at their wits' end.
PS|107|28|Then they cried out to the LORD in their trouble, and he brought them out of their distress.
PS|107|29|He stilled the storm to a whisper; the waves of the sea were hushed.
PS|107|30|They were glad when it grew calm, and he guided them to their desired haven.
PS|107|31|Let them give thanks to the LORD for his unfailing love and his wonderful deeds for men.
PS|107|32|Let them exalt him in the assembly of the people and praise him in the council of the elders.
PS|107|33|He turned rivers into a desert, flowing springs into thirsty ground,
PS|107|34|and fruitful land into a salt waste, because of the wickedness of those who lived there.
PS|107|35|He turned the desert into pools of water and the parched ground into flowing springs;
PS|107|36|there he brought the hungry to live, and they founded a city where they could settle.
PS|107|37|They sowed fields and planted vineyards that yielded a fruitful harvest;
PS|107|38|he blessed them, and their numbers greatly increased, and he did not let their herds diminish.
PS|107|39|Then their numbers decreased, and they were humbled by oppression, calamity and sorrow;
PS|107|40|he who pours contempt on nobles made them wander in a trackless waste.
PS|107|41|But he lifted the needy out of their affliction and increased their families like flocks.
PS|107|42|The upright see and rejoice, but all the wicked shut their mouths.
PS|107|43|Whoever is wise, let him heed these things and consider the great love of the LORD.
PS|108|1|My heart is steadfast, O God; I will sing and make music with all my soul.
PS|108|2|Awake, harp and lyre! I will awaken the dawn.
PS|108|3|I will praise you, O LORD, among the nations; I will sing of you among the peoples.
PS|108|4|For great is your love, higher than the heavens; your faithfulness reaches to the skies.
PS|108|5|Be exalted, O God, above the heavens, and let your glory be over all the earth.
PS|108|6|Save us and help us with your right hand, that those you love may be delivered.
PS|108|7|God has spoken from his sanctuary: "In triumph I will parcel out Shechem and measure off the Valley of Succoth.
PS|108|8|Gilead is mine, Manasseh is mine; Ephraim is my helmet, Judah my scepter.
PS|108|9|Moab is my washbasin, upon Edom I toss my sandal; over Philistia I shout in triumph."
PS|108|10|Who will bring me to the fortified city? Who will lead me to Edom?
PS|108|11|Is it not you, O God, you who have rejected us and no longer go out with our armies?
PS|108|12|Give us aid against the enemy, for the help of man is worthless.
PS|108|13|With God we will gain the victory, and he will trample down our enemies.
PS|109|1|O God, whom I praise, do not remain silent,
PS|109|2|for wicked and deceitful men have opened their mouths against me; they have spoken against me with lying tongues.
PS|109|3|With words of hatred they surround me; they attack me without cause.
PS|109|4|In return for my friendship they accuse me, but I am a man of prayer.
PS|109|5|They repay me evil for good, and hatred for my friendship.
PS|109|6|Appoint an evil man to oppose him; let an accuser stand at his right hand.
PS|109|7|When he is tried, let him be found guilty, and may his prayers condemn him.
PS|109|8|May his days be few; may another take his place of leadership.
PS|109|9|May his children be fatherless and his wife a widow.
PS|109|10|May his children be wandering beggars; may they be driven from their ruined homes.
PS|109|11|May a creditor seize all he has; may strangers plunder the fruits of his labor.
PS|109|12|May no one extend kindness to him or take pity on his fatherless children.
PS|109|13|May his descendants be cut off, their names blotted out from the next generation.
PS|109|14|May the iniquity of his fathers be remembered before the LORD; may the sin of his mother never be blotted out.
PS|109|15|May their sins always remain before the LORD, that he may cut off the memory of them from the earth.
PS|109|16|For he never thought of doing a kindness, but hounded to death the poor and the needy and the brokenhearted.
PS|109|17|He loved to pronounce a curse- may it come on him; he found no pleasure in blessing- may it be far from him.
PS|109|18|He wore cursing as his garment; it entered into his body like water, into his bones like oil.
PS|109|19|May it be like a cloak wrapped about him, like a belt tied forever around him.
PS|109|20|May this be the LORD's payment to my accusers, to those who speak evil of me.
PS|109|21|But you, O Sovereign LORD, deal well with me for your name's sake; out of the goodness of your love, deliver me.
PS|109|22|For I am poor and needy, and my heart is wounded within me.
PS|109|23|I fade away like an evening shadow; I am shaken off like a locust.
PS|109|24|My knees give way from fasting; my body is thin and gaunt.
PS|109|25|I am an object of scorn to my accusers; when they see me, they shake their heads.
PS|109|26|Help me, O LORD my God; save me in accordance with your love.
PS|109|27|Let them know that it is your hand, that you, O LORD, have done it.
PS|109|28|They may curse, but you will bless; when they attack they will be put to shame, but your servant will rejoice.
PS|109|29|My accusers will be clothed with disgrace and wrapped in shame as in a cloak.
PS|109|30|With my mouth I will greatly extol the LORD; in the great throng I will praise him.
PS|109|31|For he stands at the right hand of the needy one, to save his life from those who condemn him.
PS|110|1|The LORD says to my Lord: "Sit at my right hand until I make your enemies a footstool for your feet."
PS|110|2|The LORD will extend your mighty scepter from Zion; you will rule in the midst of your enemies.
PS|110|3|Your troops will be willing on your day of battle. Arrayed in holy majesty, from the womb of the dawn you will receive the dew of your youth.
PS|110|4|The LORD has sworn and will not change his mind: "You are a priest forever, in the order of Melchizedek."
PS|110|5|The Lord is at your right hand; he will crush kings on the day of his wrath.
PS|110|6|He will judge the nations, heaping up the dead and crushing the rulers of the whole earth.
PS|110|7|He will drink from a brook beside the way; therefore he will lift up his head.
PS|111|1|Praise the LORD. I will extol the LORD with all my heart in the council of the upright and in the assembly.
PS|111|2|Great are the works of the LORD; they are pondered by all who delight in them.
PS|111|3|Glorious and majestic are his deeds, and his righteousness endures forever.
PS|111|4|He has caused his wonders to be remembered; the LORD is gracious and compassionate.
PS|111|5|He provides food for those who fear him; he remembers his covenant forever.
PS|111|6|He has shown his people the power of his works, giving them the lands of other nations.
PS|111|7|The works of his hands are faithful and just; all his precepts are trustworthy.
PS|111|8|They are steadfast for ever and ever, done in faithfulness and uprightness.
PS|111|9|He provided redemption for his people; he ordained his covenant forever- holy and awesome is his name.
PS|111|10|The fear of the LORD is the beginning of wisdom; all who follow his precepts have good understanding. To him belongs eternal praise.
PS|112|1|Praise the LORD. Blessed is the man who fears the LORD, who finds great delight in his commands.
PS|112|2|His children will be mighty in the land; the generation of the upright will be blessed.
PS|112|3|Wealth and riches are in his house, and his righteousness endures forever.
PS|112|4|Even in darkness light dawns for the upright, for the gracious and compassionate and righteous man.
PS|112|5|Good will come to him who is generous and lends freely, who conducts his affairs with justice.
PS|112|6|Surely he will never be shaken; a righteous man will be remembered forever.
PS|112|7|He will have no fear of bad news; his heart is steadfast, trusting in the LORD.
PS|112|8|His heart is secure, he will have no fear; in the end he will look in triumph on his foes.
PS|112|9|He has scattered abroad his gifts to the poor, his righteousness endures forever; his horn will be lifted high in honor.
PS|112|10|The wicked man will see and be vexed, he will gnash his teeth and waste away; the longings of the wicked will come to nothing.
PS|113|1|Praise the LORD. Praise, O servants of the LORD, praise the name of the LORD.
PS|113|2|Let the name of the LORD be praised, both now and forevermore.
PS|113|3|From the rising of the sun to the place where it sets, the name of the LORD is to be praised.
PS|113|4|The LORD is exalted over all the nations, his glory above the heavens.
PS|113|5|Who is like the LORD our God, the One who sits enthroned on high,
PS|113|6|who stoops down to look on the heavens and the earth?
PS|113|7|He raises the poor from the dust and lifts the needy from the ash heap;
PS|113|8|he seats them with princes, with the princes of their people.
PS|113|9|He settles the barren woman in her home as a happy mother of children. Praise the LORD.
PS|114|1|When Israel came out of Egypt, the house of Jacob from a people of foreign tongue,
PS|114|2|Judah became God's sanctuary, Israel his dominion.
PS|114|3|The sea looked and fled, the Jordan turned back;
PS|114|4|the mountains skipped like rams, the hills like lambs.
PS|114|5|Why was it, O sea, that you fled, O Jordan, that you turned back,
PS|114|6|you mountains, that you skipped like rams, you hills, like lambs?
PS|114|7|Tremble, O earth, at the presence of the Lord, at the presence of the God of Jacob,
PS|114|8|who turned the rock into a pool, the hard rock into springs of water.
PS|115|1|Not to us, O LORD, not to us but to your name be the glory, because of your love and faithfulness.
PS|115|2|Why do the nations say, "Where is their God?"
PS|115|3|Our God is in heaven; he does whatever pleases him.
PS|115|4|But their idols are silver and gold, made by the hands of men.
PS|115|5|They have mouths, but cannot speak, eyes, but they cannot see;
PS|115|6|they have ears, but cannot hear, noses, but they cannot smell;
PS|115|7|they have hands, but cannot feel, feet, but they cannot walk; nor can they utter a sound with their throats.
PS|115|8|Those who make them will be like them, and so will all who trust in them.
PS|115|9|O house of Israel, trust in the LORD - he is their help and shield.
PS|115|10|O house of Aaron, trust in the LORD - he is their help and shield.
PS|115|11|You who fear him, trust in the LORD - he is their help and shield.
PS|115|12|The LORD remembers us and will bless us: He will bless the house of Israel, he will bless the house of Aaron,
PS|115|13|he will bless those who fear the LORD - small and great alike.
PS|115|14|May the LORD make you increase, both you and your children.
PS|115|15|May you be blessed by the LORD, the Maker of heaven and earth.
PS|115|16|The highest heavens belong to the LORD, but the earth he has given to man.
PS|115|17|It is not the dead who praise the LORD, those who go down to silence;
PS|115|18|it is we who extol the LORD, both now and forevermore. Praise the LORD.
PS|116|1|I love the LORD, for he heard my voice; he heard my cry for mercy.
PS|116|2|Because he turned his ear to me, I will call on him as long as I live.
PS|116|3|The cords of death entangled me, the anguish of the grave came upon me; I was overcome by trouble and sorrow.
PS|116|4|Then I called on the name of the LORD: "O LORD, save me!"
PS|116|5|The LORD is gracious and righteous; our God is full of compassion.
PS|116|6|The LORD protects the simplehearted; when I was in great need, he saved me.
PS|116|7|Be at rest once more, O my soul, for the LORD has been good to you.
PS|116|8|For you, O LORD, have delivered my soul from death, my eyes from tears, my feet from stumbling,
PS|116|9|that I may walk before the LORD in the land of the living.
PS|116|10|I believed; therefore I said, "I am greatly afflicted."
PS|116|11|And in my dismay I said, "All men are liars."
PS|116|12|How can I repay the LORD for all his goodness to me?
PS|116|13|I will lift up the cup of salvation and call on the name of the LORD.
PS|116|14|I will fulfill my vows to the LORD in the presence of all his people.
PS|116|15|Precious in the sight of the LORD is the death of his saints.
PS|116|16|O LORD, truly I am your servant; I am your servant, the son of your maidservant; you have freed me from my chains.
PS|116|17|I will sacrifice a thank offering to you and call on the name of the LORD.
PS|116|18|I will fulfill my vows to the LORD in the presence of all his people,
PS|116|19|in the courts of the house of the LORD - in your midst, O Jerusalem. Praise the LORD.
PS|117|1|Praise the LORD, all you nations; extol him, all you peoples.
PS|117|2|For great is his love toward us, and the faithfulness of the LORD endures forever. Praise the LORD.
PS|118|1|Give thanks to the LORD, for he is good; his love endures forever.
PS|118|2|Let Israel say: "His love endures forever."
PS|118|3|Let the house of Aaron say: "His love endures forever."
PS|118|4|Let those who fear the LORD say: "His love endures forever."
PS|118|5|In my anguish I cried to the LORD, and he answered by setting me free.
PS|118|6|The LORD is with me; I will not be afraid. What can man do to me?
PS|118|7|The LORD is with me; he is my helper. I will look in triumph on my enemies.
PS|118|8|It is better to take refuge in the LORD than to trust in man.
PS|118|9|It is better to take refuge in the LORD than to trust in princes.
PS|118|10|All the nations surrounded me, but in the name of the LORD I cut them off.
PS|118|11|They surrounded me on every side, but in the name of the LORD I cut them off.
PS|118|12|They swarmed around me like bees, but they died out as quickly as burning thorns; in the name of the LORD I cut them off.
PS|118|13|I was pushed back and about to fall, but the LORD helped me.
PS|118|14|The LORD is my strength and my song; he has become my salvation.
PS|118|15|Shouts of joy and victory resound in the tents of the righteous: "The LORD's right hand has done mighty things!
PS|118|16|The LORD's right hand is lifted high; the LORD's right hand has done mighty things!"
PS|118|17|I will not die but live, and will proclaim what the LORD has done.
PS|118|18|The LORD has chastened me severely, but he has not given me over to death.
PS|118|19|Open for me the gates of righteousness; I will enter and give thanks to the LORD.
PS|118|20|This is the gate of the LORD through which the righteous may enter.
PS|118|21|I will give you thanks, for you answered me; you have become my salvation.
PS|118|22|The stone the builders rejected has become the capstone;
PS|118|23|the LORD has done this, and it is marvelous in our eyes.
PS|118|24|This is the day the LORD has made; let us rejoice and be glad in it.
PS|118|25|O LORD, save us; O LORD, grant us success.
PS|118|26|Blessed is he who comes in the name of the LORD. From the house of the LORD we bless you.
PS|118|27|The LORD is God, and he has made his light shine upon us. With boughs in hand, join in the festal procession up to the horns of the altar.
PS|118|28|You are my God, and I will give you thanks; you are my God, and I will exalt you.
PS|118|29|Give thanks to the LORD, for he is good; his love endures forever.
PS|119|1|Blessed are they whose ways are blameless, who walk according to the law of the LORD.
PS|119|2|Blessed are they who keep his statutes and seek him with all their heart.
PS|119|3|They do nothing wrong; they walk in his ways.
PS|119|4|You have laid down precepts that are to be fully obeyed.
PS|119|5|Oh, that my ways were steadfast in obeying your decrees!
PS|119|6|Then I would not be put to shame when I consider all your commands.
PS|119|7|I will praise you with an upright heart as I learn your righteous laws.
PS|119|8|I will obey your decrees; do not utterly forsake me.
PS|119|9|How can a young man keep his way pure? By living according to your word.
PS|119|10|I seek you with all my heart; do not let me stray from your commands.
PS|119|11|I have hidden your word in my heart that I might not sin against you.
PS|119|12|Praise be to you, O LORD; teach me your decrees.
PS|119|13|With my lips I recount all the laws that come from your mouth.
PS|119|14|I rejoice in following your statutes as one rejoices in great riches.
PS|119|15|I meditate on your precepts and consider your ways.
PS|119|16|I delight in your decrees; I will not neglect your word.
PS|119|17|Do good to your servant, and I will live; I will obey your word.
PS|119|18|Open my eyes that I may see wonderful things in your law.
PS|119|19|I am a stranger on earth; do not hide your commands from me.
PS|119|20|My soul is consumed with longing for your laws at all times.
PS|119|21|You rebuke the arrogant, who are cursed and who stray from your commands.
PS|119|22|Remove from me scorn and contempt, for I keep your statutes.
PS|119|23|Though rulers sit together and slander me, your servant will meditate on your decrees.
PS|119|24|Your statutes are my delight; they are my counselors.
PS|119|25|I am laid low in the dust; preserve my life according to your word.
PS|119|26|I recounted my ways and you answered me; teach me your decrees.
PS|119|27|Let me understand the teaching of your precepts; then I will meditate on your wonders.
PS|119|28|My soul is weary with sorrow; strengthen me according to your word.
PS|119|29|Keep me from deceitful ways; be gracious to me through your law.
PS|119|30|I have chosen the way of truth; I have set my heart on your laws.
PS|119|31|I hold fast to your statutes, O LORD; do not let me be put to shame.
PS|119|32|I run in the path of your commands, for you have set my heart free.
PS|119|33|Teach me, O LORD, to follow your decrees; then I will keep them to the end.
PS|119|34|Give me understanding, and I will keep your law and obey it with all my heart.
PS|119|35|Direct me in the path of your commands, for there I find delight.
PS|119|36|Turn my heart toward your statutes and not toward selfish gain.
PS|119|37|Turn my eyes away from worthless things; preserve my life according to your word.
PS|119|38|Fulfill your promise to your servant, so that you may be feared.
PS|119|39|Take away the disgrace I dread, for your laws are good.
PS|119|40|How I long for your precepts! Preserve my life in your righteousness.
PS|119|41|May your unfailing love come to me, O LORD, your salvation according to your promise;
PS|119|42|then I will answer the one who taunts me, for I trust in your word.
PS|119|43|Do not snatch the word of truth from my mouth, for I have put my hope in your laws.
PS|119|44|I will always obey your law, for ever and ever.
PS|119|45|I will walk about in freedom, for I have sought out your precepts.
PS|119|46|I will speak of your statutes before kings and will not be put to shame,
PS|119|47|for I delight in your commands because I love them.
PS|119|48|I lift up my hands to your commands, which I love, and I meditate on your decrees.
PS|119|49|Remember your word to your servant, for you have given me hope.
PS|119|50|My comfort in my suffering is this: Your promise preserves my life.
PS|119|51|The arrogant mock me without restraint, but I do not turn from your law.
PS|119|52|I remember your ancient laws, O LORD, and I find comfort in them.
PS|119|53|Indignation grips me because of the wicked, who have forsaken your law.
PS|119|54|Your decrees are the theme of my song wherever I lodge.
PS|119|55|In the night I remember your name, O LORD, and I will keep your law.
PS|119|56|This has been my practice: I obey your precepts.
PS|119|57|You are my portion, O LORD; I have promised to obey your words.
PS|119|58|I have sought your face with all my heart; be gracious to me according to your promise.
PS|119|59|I have considered my ways and have turned my steps to your statutes.
PS|119|60|I will hasten and not delay to obey your commands.
PS|119|61|Though the wicked bind me with ropes, I will not forget your law.
PS|119|62|At midnight I rise to give you thanks for your righteous laws.
PS|119|63|I am a friend to all who fear you, to all who follow your precepts.
PS|119|64|The earth is filled with your love, O LORD; teach me your decrees.
PS|119|65|Do good to your servant according to your word, O LORD.
PS|119|66|Teach me knowledge and good judgment, for I believe in your commands.
PS|119|67|Before I was afflicted I went astray, but now I obey your word.
PS|119|68|You are good, and what you do is good; teach me your decrees.
PS|119|69|Though the arrogant have smeared me with lies, I keep your precepts with all my heart.
PS|119|70|Their hearts are callous and unfeeling, but I delight in your law.
PS|119|71|It was good for me to be afflicted so that I might learn your decrees.
PS|119|72|The law from your mouth is more precious to me than thousands of pieces of silver and gold.
PS|119|73|Your hands made me and formed me; give me understanding to learn your commands.
PS|119|74|May those who fear you rejoice when they see me, for I have put my hope in your word.
PS|119|75|I know, O LORD, that your laws are righteous, and in faithfulness you have afflicted me.
PS|119|76|May your unfailing love be my comfort, according to your promise to your servant.
PS|119|77|Let your compassion come to me that I may live, for your law is my delight.
PS|119|78|May the arrogant be put to shame for wronging me without cause; but I will meditate on your precepts.
PS|119|79|May those who fear you turn to me, those who understand your statutes.
PS|119|80|May my heart be blameless toward your decrees, that I may not be put to shame.
PS|119|81|My soul faints with longing for your salvation, but I have put my hope in your word.
PS|119|82|My eyes fail, looking for your promise; I say, "When will you comfort me?"
PS|119|83|Though I am like a wineskin in the smoke, I do not forget your decrees.
PS|119|84|How long must your servant wait? When will you punish my persecutors?
PS|119|85|The arrogant dig pitfalls for me, contrary to your law.
PS|119|86|All your commands are trustworthy; help me, for men persecute me without cause.
PS|119|87|They almost wiped me from the earth, but I have not forsaken your precepts.
PS|119|88|Preserve my life according to your love, and I will obey the statutes of your mouth.
PS|119|89|Your word, O LORD, is eternal; it stands firm in the heavens.
PS|119|90|Your faithfulness continues through all generations; you established the earth, and it endures.
PS|119|91|Your laws endure to this day, for all things serve you.
PS|119|92|If your law had not been my delight, I would have perished in my affliction.
PS|119|93|I will never forget your precepts, for by them you have preserved my life.
PS|119|94|Save me, for I am yours; I have sought out your precepts.
PS|119|95|The wicked are waiting to destroy me, but I will ponder your statutes.
PS|119|96|To all perfection I see a limit; but your commands are boundless.
PS|119|97|Oh, how I love your law! I meditate on it all day long.
PS|119|98|Your commands make me wiser than my enemies, for they are ever with me.
PS|119|99|I have more insight than all my teachers, for I meditate on your statutes.
PS|119|100|I have more understanding than the elders, for I obey your precepts.
PS|119|101|I have kept my feet from every evil path so that I might obey your word.
PS|119|102|I have not departed from your laws, for you yourself have taught me.
PS|119|103|How sweet are your words to my taste, sweeter than honey to my mouth!
PS|119|104|I gain understanding from your precepts; therefore I hate every wrong path.
PS|119|105|Your word is a lamp to my feet and a light for my path.
PS|119|106|I have taken an oath and confirmed it, that I will follow your righteous laws.
PS|119|107|I have suffered much; preserve my life, O LORD, according to your word.
PS|119|108|Accept, O LORD, the willing praise of my mouth, and teach me your laws.
PS|119|109|Though I constantly take my life in my hands, I will not forget your law.
PS|119|110|The wicked have set a snare for me, but I have not strayed from your precepts.
PS|119|111|Your statutes are my heritage forever; they are the joy of my heart.
PS|119|112|My heart is set on keeping your decrees to the very end.
PS|119|113|I hate double-minded men, but I love your law.
PS|119|114|You are my refuge and my shield; I have put my hope in your word.
PS|119|115|Away from me, you evildoers, that I may keep the commands of my God!
PS|119|116|Sustain me according to your promise, and I will live; do not let my hopes be dashed.
PS|119|117|Uphold me, and I will be delivered; I will always have regard for your decrees.
PS|119|118|You reject all who stray from your decrees, for their deceitfulness is in vain.
PS|119|119|All the wicked of the earth you discard like dross; therefore I love your statutes.
PS|119|120|My flesh trembles in fear of you; I stand in awe of your laws.
PS|119|121|I have done what is righteous and just; do not leave me to my oppressors.
PS|119|122|Ensure your servant's well-being; let not the arrogant oppress me.
PS|119|123|My eyes fail, looking for your salvation, looking for your righteous promise.
PS|119|124|Deal with your servant according to your love and teach me your decrees.
PS|119|125|I am your servant; give me discernment that I may understand your statutes.
PS|119|126|It is time for you to act, O LORD; your law is being broken.
PS|119|127|Because I love your commands more than gold, more than pure gold,
PS|119|128|and because I consider all your precepts right, I hate every wrong path.
PS|119|129|Your statutes are wonderful; therefore I obey them.
PS|119|130|The unfolding of your words gives light; it gives understanding to the simple.
PS|119|131|I open my mouth and pant, longing for your commands.
PS|119|132|Turn to me and have mercy on me, as you always do to those who love your name.
PS|119|133|Direct my footsteps according to your word; let no sin rule over me.
PS|119|134|Redeem me from the oppression of men, that I may obey your precepts.
PS|119|135|Make your face shine upon your servant and teach me your decrees.
PS|119|136|Streams of tears flow from my eyes, for your law is not obeyed.
PS|119|137|Righteous are you, O LORD, and your laws are right.
PS|119|138|The statutes you have laid down are righteous; they are fully trustworthy.
PS|119|139|My zeal wears me out, for my enemies ignore your words.
PS|119|140|Your promises have been thoroughly tested, and your servant loves them.
PS|119|141|Though I am lowly and despised, I do not forget your precepts.
PS|119|142|Your righteousness is everlasting and your law is true.
PS|119|143|Trouble and distress have come upon me, but your commands are my delight.
PS|119|144|Your statutes are forever right; give me understanding that I may live.
PS|119|145|I call with all my heart; answer me, O LORD, and I will obey your decrees.
PS|119|146|I call out to you; save me and I will keep your statutes.
PS|119|147|I rise before dawn and cry for help; I have put my hope in your word.
PS|119|148|My eyes stay open through the watches of the night, that I may meditate on your promises.
PS|119|149|Hear my voice in accordance with your love; preserve my life, O LORD, according to your laws.
PS|119|150|Those who devise wicked schemes are near, but they are far from your law.
PS|119|151|Yet you are near, O LORD, and all your commands are true.
PS|119|152|Long ago I learned from your statutes that you established them to last forever.
PS|119|153|Look upon my suffering and deliver me, for I have not forgotten your law.
PS|119|154|Defend my cause and redeem me; preserve my life according to your promise.
PS|119|155|Salvation is far from the wicked, for they do not seek out your decrees.
PS|119|156|Your compassion is great, O LORD; preserve my life according to your laws.
PS|119|157|Many are the foes who persecute me, but I have not turned from your statutes.
PS|119|158|I look on the faithless with loathing, for they do not obey your word.
PS|119|159|See how I love your precepts; preserve my life, O LORD, according to your love.
PS|119|160|All your words are true; all your righteous laws are eternal.
PS|119|161|Rulers persecute me without cause, but my heart trembles at your word.
PS|119|162|I rejoice in your promise like one who finds great spoil.
PS|119|163|I hate and abhor falsehood but I love your law.
PS|119|164|Seven times a day I praise you for your righteous laws.
PS|119|165|Great peace have they who love your law, and nothing can make them stumble.
PS|119|166|I wait for your salvation, O LORD, and I follow your commands.
PS|119|167|I obey your statutes, for I love them greatly.
PS|119|168|I obey your precepts and your statutes, for all my ways are known to you.
PS|119|169|May my cry come before you, O LORD; give me understanding according to your word.
PS|119|170|May my supplication come before you; deliver me according to your promise.
PS|119|171|May my lips overflow with praise, for you teach me your decrees.
PS|119|172|May my tongue sing of your word, for all your commands are righteous.
PS|119|173|May your hand be ready to help me, for I have chosen your precepts.
PS|119|174|I long for your salvation, O LORD, and your law is my delight.
PS|119|175|Let me live that I may praise you, and may your laws sustain me.
PS|119|176|I have strayed like a lost sheep. Seek your servant, for I have not forgotten your commands.
PS|120|1|I call on the LORD in my distress, and he answers me.
PS|120|2|Save me, O LORD, from lying lips and from deceitful tongues.
PS|120|3|What will he do to you, and what more besides, O deceitful tongue?
PS|120|4|He will punish you with a warrior's sharp arrows, with burning coals of the broom tree.
PS|120|5|Woe to me that I dwell in Meshech, that I live among the tents of Kedar!
PS|120|6|Too long have I lived among those who hate peace.
PS|120|7|I am a man of peace; but when I speak, they are for war.
PS|121|1|I lift up my eyes to the hills- where does my help come from?
PS|121|2|My help comes from the LORD, the Maker of heaven and earth.
PS|121|3|He will not let your foot slip- he who watches over you will not slumber;
PS|121|4|indeed, he who watches over Israel will neither slumber nor sleep.
PS|121|5|The LORD watches over you- the LORD is your shade at your right hand;
PS|121|6|the sun will not harm you by day, nor the moon by night.
PS|121|7|The LORD will keep you from all harm- he will watch over your life;
PS|121|8|the LORD will watch over your coming and going both now and forevermore.
PS|122|1|I rejoiced with those who said to me, "Let us go to the house of the LORD."
PS|122|2|Our feet are standing in your gates, O Jerusalem.
PS|122|3|Jerusalem is built like a city that is closely compacted together.
PS|122|4|That is where the tribes go up, the tribes of the LORD, to praise the name of the LORD according to the statute given to Israel.
PS|122|5|There the thrones for judgment stand, the thrones of the house of David.
PS|122|6|Pray for the peace of Jerusalem: "May those who love you be secure.
PS|122|7|May there be peace within your walls and security within your citadels."
PS|122|8|For the sake of my brothers and friends, I will say, "Peace be within you."
PS|122|9|For the sake of the house of the LORD our God, I will seek your prosperity.
PS|123|1|I lift up my eyes to you, to you whose throne is in heaven.
PS|123|2|As the eyes of slaves look to the hand of their master, as the eyes of a maid look to the hand of her mistress, so our eyes look to the LORD our God, till he shows us his mercy.
PS|123|3|Have mercy on us, O LORD, have mercy on us, for we have endured much contempt.
PS|123|4|We have endured much ridicule from the proud, much contempt from the arrogant.
PS|124|1|If the LORD had not been on our side- let Israel say-
PS|124|2|if the LORD had not been on our side when men attacked us,
PS|124|3|when their anger flared against us, they would have swallowed us alive;
PS|124|4|the flood would have engulfed us, the torrent would have swept over us,
PS|124|5|the raging waters would have swept us away.
PS|124|6|Praise be to the LORD, who has not let us be torn by their teeth.
PS|124|7|We have escaped like a bird out of the fowler's snare; the snare has been broken, and we have escaped.
PS|124|8|Our help is in the name of the LORD, the Maker of heaven and earth.
PS|125|1|Those who trust in the LORD are like Mount Zion, which cannot be shaken but endures forever.
PS|125|2|As the mountains surround Jerusalem, so the LORD surrounds his people both now and forevermore.
PS|125|3|The scepter of the wicked will not remain over the land allotted to the righteous, for then the righteous might use their hands to do evil.
PS|125|4|Do good, O LORD, to those who are good, to those who are upright in heart.
PS|125|5|But those who turn to crooked ways the LORD will banish with the evildoers. Peace be upon Israel.
PS|126|1|When the LORD brought back the captives to Zion, we were like men who dreamed.
PS|126|2|Our mouths were filled with laughter, our tongues with songs of joy. Then it was said among the nations, "The LORD has done great things for them."
PS|126|3|The LORD has done great things for us, and we are filled with joy.
PS|126|4|Restore our fortunes, O LORD, like streams in the Negev.
PS|126|5|Those who sow in tears will reap with songs of joy.
PS|126|6|He who goes out weeping, carrying seed to sow, will return with songs of joy, carrying sheaves with him.
PS|127|1|Unless the LORD builds the house, its builders labor in vain. Unless the LORD watches over the city, the watchmen stand guard in vain.
PS|127|2|In vain you rise early and stay up late, toiling for food to eat- for he grants sleep to those he loves.
PS|127|3|Sons are a heritage from the LORD, children a reward from him.
PS|127|4|Like arrows in the hands of a warrior are sons born in one's youth.
PS|127|5|Blessed is the man whose quiver is full of them. They will not be put to shame when they contend with their enemies in the gate.
PS|128|1|Blessed are all who fear the LORD, who walk in his ways.
PS|128|2|You will eat the fruit of your labor; blessings and prosperity will be yours.
PS|128|3|Your wife will be like a fruitful vine within your house; your sons will be like olive shoots around your table.
PS|128|4|Thus is the man blessed who fears the LORD.
PS|128|5|May the LORD bless you from Zion all the days of your life; may you see the prosperity of Jerusalem,
PS|128|6|and may you live to see your children's children. Peace be upon Israel.
PS|129|1|They have greatly oppressed me from my youth- let Israel say-
PS|129|2|they have greatly oppressed me from my youth, but they have not gained the victory over me.
PS|129|3|Plowmen have plowed my back and made their furrows long.
PS|129|4|But the LORD is righteous; he has cut me free from the cords of the wicked.
PS|129|5|May all who hate Zion be turned back in shame.
PS|129|6|May they be like grass on the roof, which withers before it can grow;
PS|129|7|with it the reaper cannot fill his hands, nor the one who gathers fill his arms.
PS|129|8|May those who pass by not say, "The blessing of the LORD be upon you; we bless you in the name of the LORD."
PS|130|1|Out of the depths I cry to you, O LORD;
PS|130|2|O Lord, hear my voice. Let your ears be attentive to my cry for mercy.
PS|130|3|If you, O LORD, kept a record of sins, O Lord, who could stand?
PS|130|4|But with you there is forgiveness; therefore you are feared.
PS|130|5|I wait for the LORD, my soul waits, and in his word I put my hope.
PS|130|6|My soul waits for the Lord more than watchmen wait for the morning, more than watchmen wait for the morning.
PS|130|7|O Israel, put your hope in the LORD, for with the LORD is unfailing love and with him is full redemption.
PS|130|8|He himself will redeem Israel from all their sins.
PS|131|1|My heart is not proud, O LORD, my eyes are not haughty; I do not concern myself with great matters or things too wonderful for me.
PS|131|2|But I have stilled and quieted my soul; like a weaned child with its mother, like a weaned child is my soul within me.
PS|131|3|O Israel, put your hope in the LORD both now and forevermore.
PS|132|1|O LORD, remember David and all the hardships he endured.
PS|132|2|He swore an oath to the LORD and made a vow to the Mighty One of Jacob:
PS|132|3|"I will not enter my house or go to my bed-
PS|132|4|I will allow no sleep to my eyes, no slumber to my eyelids,
PS|132|5|till I find a place for the LORD, a dwelling for the Mighty One of Jacob."
PS|132|6|We heard it in Ephrathah, we came upon it in the fields of Jaar:
PS|132|7|"Let us go to his dwelling place; let us worship at his footstool-
PS|132|8|arise, O LORD, and come to your resting place, you and the ark of your might.
PS|132|9|May your priests be clothed with righteousness; may your saints sing for joy."
PS|132|10|For the sake of David your servant, do not reject your anointed one.
PS|132|11|The LORD swore an oath to David, a sure oath that he will not revoke: "One of your own descendants I will place on your throne-
PS|132|12|if your sons keep my covenant and the statutes I teach them, then their sons will sit on your throne for ever and ever."
PS|132|13|For the LORD has chosen Zion, he has desired it for his dwelling:
PS|132|14|"This is my resting place for ever and ever; here I will sit enthroned, for I have desired it-
PS|132|15|I will bless her with abundant provisions; her poor will I satisfy with food.
PS|132|16|I will clothe her priests with salvation, and her saints will ever sing for joy.
PS|132|17|"Here I will make a horn grow for David and set up a lamp for my anointed one.
PS|132|18|I will clothe his enemies with shame, but the crown on his head will be resplendent."
PS|133|1|How good and pleasant it is when brothers live together in unity!
PS|133|2|It is like precious oil poured on the head, running down on the beard, running down on Aaron's beard, down upon the collar of his robes.
PS|133|3|It is as if the dew of Hermon were falling on Mount Zion. For there the LORD bestows his blessing, even life forevermore.
PS|134|1|Praise the LORD, all you servants of the LORD who minister by night in the house of the LORD.
PS|134|2|Lift up your hands in the sanctuary and praise the LORD.
PS|134|3|May the LORD, the Maker of heaven and earth, bless you from Zion.
PS|135|1|Praise the LORD. Praise the name of the LORD; praise him, you servants of the LORD,
PS|135|2|you who minister in the house of the LORD, in the courts of the house of our God.
PS|135|3|Praise the LORD, for the LORD is good; sing praise to his name, for that is pleasant.
PS|135|4|For the LORD has chosen Jacob to be his own, Israel to be his treasured possession.
PS|135|5|I know that the LORD is great, that our Lord is greater than all gods.
PS|135|6|The LORD does whatever pleases him, in the heavens and on the earth, in the seas and all their depths.
PS|135|7|He makes clouds rise from the ends of the earth; he sends lightning with the rain and brings out the wind from his storehouses.
PS|135|8|He struck down the firstborn of Egypt, the firstborn of men and animals.
PS|135|9|He sent his signs and wonders into your midst, O Egypt, against Pharaoh and all his servants.
PS|135|10|He struck down many nations and killed mighty kings-
PS|135|11|Sihon king of the Amorites, Og king of Bashan and all the kings of Canaan-
PS|135|12|and he gave their land as an inheritance, an inheritance to his people Israel.
PS|135|13|Your name, O LORD, endures forever, your renown, O LORD, through all generations.
PS|135|14|For the LORD will vindicate his people and have compassion on his servants.
PS|135|15|The idols of the nations are silver and gold, made by the hands of men.
PS|135|16|They have mouths, but cannot speak, eyes, but they cannot see;
PS|135|17|they have ears, but cannot hear, nor is there breath in their mouths.
PS|135|18|Those who make them will be like them, and so will all who trust in them.
PS|135|19|O house of Israel, praise the LORD; O house of Aaron, praise the LORD;
PS|135|20|O house of Levi, praise the LORD; you who fear him, praise the LORD.
PS|135|21|Praise be to the LORD from Zion, to him who dwells in Jerusalem. Praise the LORD.
PS|136|1|Give thanks to the LORD, for he is good. His love endures forever.
PS|136|2|Give thanks to the God of gods. His love endures forever.
PS|136|3|Give thanks to the Lord of lords: His love endures forever.
PS|136|4|to him who alone does great wonders, His love endures forever.
PS|136|5|who by his understanding made the heavens, His love endures forever.
PS|136|6|who spread out the earth upon the waters, His love endures forever.
PS|136|7|who made the great lights- His love endures forever.
PS|136|8|the sun to govern the day, His love endures forever.
PS|136|9|the moon and stars to govern the night; His love endures forever.
PS|136|10|to him who struck down the firstborn of Egypt His love endures forever.
PS|136|11|and brought Israel out from among them His love endures forever.
PS|136|12|with a mighty hand and outstretched arm; His love endures forever.
PS|136|13|to him who divided the Red Sea asunder His love endures forever.
PS|136|14|and brought Israel through the midst of it, His love endures forever.
PS|136|15|but swept Pharaoh and his army into the Red Sea; His love endures forever.
PS|136|16|to him who led his people through the desert, His love endures forever.
PS|136|17|who struck down great kings, His love endures forever.
PS|136|18|and killed mighty kings- His love endures forever.
PS|136|19|Sihon king of the Amorites His love endures forever.
PS|136|20|and Og king of Bashan- His love endures forever.
PS|136|21|and gave their land as an inheritance, His love endures forever.
PS|136|22|an inheritance to his servant Israel; His love endures forever.
PS|136|23|to the One who remembered us in our low estate His love endures forever.
PS|136|24|and freed us from our enemies, His love endures forever.
PS|136|25|and who gives food to every creature. His love endures forever.
PS|136|26|Give thanks to the God of heaven. His love endures forever.
PS|137|1|By the rivers of Babylon we sat and wept when we remembered Zion.
PS|137|2|There on the poplars we hung our harps,
PS|137|3|for there our captors asked us for songs, our tormentors demanded songs of joy; they said, "Sing us one of the songs of Zion!"
PS|137|4|How can we sing the songs of the LORD while in a foreign land?
PS|137|5|If I forget you, O Jerusalem, may my right hand forget its skill.
PS|137|6|May my tongue cling to the roof of my mouth if I do not remember you, if I do not consider Jerusalem my highest joy.
PS|137|7|Remember, O LORD, what the Edomites did on the day Jerusalem fell. "Tear it down," they cried, "tear it down to its foundations!"
PS|137|8|O Daughter of Babylon, doomed to destruction, happy is he who repays you for what you have done to us-
PS|137|9|he who seizes your infants and dashes them against the rocks.
PS|138|1|I will praise you, O LORD, with all my heart; before the "gods" I will sing your praise.
PS|138|2|I will bow down toward your holy temple and will praise your name for your love and your faithfulness, for you have exalted above all things your name and your word.
PS|138|3|When I called, you answered me; you made me bold and stouthearted.
PS|138|4|May all the kings of the earth praise you, O LORD, when they hear the words of your mouth.
PS|138|5|May they sing of the ways of the LORD, for the glory of the LORD is great.
PS|138|6|Though the LORD is on high, he looks upon the lowly, but the proud he knows from afar.
PS|138|7|Though I walk in the midst of trouble, you preserve my life; you stretch out your hand against the anger of my foes, with your right hand you save me.
PS|138|8|The LORD will fulfill his purpose for me; your love, O LORD, endures forever- do not abandon the works of your hands.
PS|139|1|O LORD, you have searched me and you know me.
PS|139|2|You know when I sit and when I rise; you perceive my thoughts from afar.
PS|139|3|You discern my going out and my lying down; you are familiar with all my ways.
PS|139|4|Before a word is on my tongue you know it completely, O LORD.
PS|139|5|You hem me in-behind and before; you have laid your hand upon me.
PS|139|6|Such knowledge is too wonderful for me, too lofty for me to attain.
PS|139|7|Where can I go from your Spirit? Where can I flee from your presence?
PS|139|8|If I go up to the heavens, you are there; if I make my bed in the depths, you are there.
PS|139|9|If I rise on the wings of the dawn, if I settle on the far side of the sea,
PS|139|10|even there your hand will guide me, your right hand will hold me fast.
PS|139|11|If I say, "Surely the darkness will hide me and the light become night around me,"
PS|139|12|even the darkness will not be dark to you; the night will shine like the day, for darkness is as light to you.
PS|139|13|For you created my inmost being; you knit me together in my mother's womb.
PS|139|14|I praise you because I am fearfully and wonderfully made; your works are wonderful, I know that full well.
PS|139|15|My frame was not hidden from you when I was made in the secret place. When I was woven together in the depths of the earth,
PS|139|16|your eyes saw my unformed body. All the days ordained for me were written in your book before one of them came to be.
PS|139|17|How precious to me are your thoughts, O God! How vast is the sum of them!
PS|139|18|Were I to count them, they would outnumber the grains of sand. When I awake, I am still with you.
PS|139|19|If only you would slay the wicked, O God! Away from me, you bloodthirsty men!
PS|139|20|They speak of you with evil intent; your adversaries misuse your name.
PS|139|21|Do I not hate those who hate you, O LORD, and abhor those who rise up against you?
PS|139|22|I have nothing but hatred for them; I count them my enemies.
PS|139|23|Search me, O God, and know my heart; test me and know my anxious thoughts.
PS|139|24|See if there is any offensive way in me, and lead me in the way everlasting.
PS|140|1|Rescue me, O LORD, from evil men; protect me from men of violence,
PS|140|2|who devise evil plans in their hearts and stir up war every day.
PS|140|3|They make their tongues as sharp as a serpent's; the poison of vipers is on their lips. Selah
PS|140|4|Keep me, O LORD, from the hands of the wicked; protect me from men of violence who plan to trip my feet.
PS|140|5|Proud men have hidden a snare for me; they have spread out the cords of their net and have set traps for me along my path. Selah
PS|140|6|O LORD, I say to you, "You are my God." Hear, O LORD, my cry for mercy.
PS|140|7|O Sovereign LORD, my strong deliverer, who shields my head in the day of battle-
PS|140|8|do not grant the wicked their desires, O LORD; do not let their plans succeed, or they will become proud. Selah
PS|140|9|Let the heads of those who surround me be covered with the trouble their lips have caused.
PS|140|10|Let burning coals fall upon them; may they be thrown into the fire, into miry pits, never to rise.
PS|140|11|Let slanderers not be established in the land; may disaster hunt down men of violence.
PS|140|12|I know that the LORD secures justice for the poor and upholds the cause of the needy.
PS|140|13|Surely the righteous will praise your name and the upright will live before you.
PS|141|1|O LORD, I call to you; come quickly to me. Hear my voice when I call to you.
PS|141|2|May my prayer be set before you like incense; may the lifting up of my hands be like the evening sacrifice.
PS|141|3|Set a guard over my mouth, O LORD; keep watch over the door of my lips.
PS|141|4|Let not my heart be drawn to what is evil, to take part in wicked deeds with men who are evildoers; let me not eat of their delicacies.
PS|141|5|Let a righteous man strike me-it is a kindness; let him rebuke me-it is oil on my head. My head will not refuse it. Yet my prayer is ever against the deeds of evildoers;
PS|141|6|their rulers will be thrown down from the cliffs, and the wicked will learn that my words were well spoken.
PS|141|7|They will say, "As one plows and breaks up the earth, so our bones have been scattered at the mouth of the grave. "
PS|141|8|But my eyes are fixed on you, O Sovereign LORD; in you I take refuge-do not give me over to death.
PS|141|9|Keep me from the snares they have laid for me, from the traps set by evildoers.
PS|141|10|Let the wicked fall into their own nets, while I pass by in safety.
PS|142|1|I cry aloud to the LORD; I lift up my voice to the LORD for mercy.
PS|142|2|I pour out my complaint before him; before him I tell my trouble.
PS|142|3|When my spirit grows faint within me, it is you who know my way. In the path where I walk men have hidden a snare for me.
PS|142|4|Look to my right and see; no one is concerned for me. I have no refuge; no one cares for my life.
PS|142|5|I cry to you, O LORD; I say, "You are my refuge, my portion in the land of the living."
PS|142|6|Listen to my cry, for I am in desperate need; rescue me from those who pursue me, for they are too strong for me.
PS|142|7|Set me free from my prison, that I may praise your name. Then the righteous will gather about me because of your goodness to me.
PS|143|1|O LORD, hear my prayer, listen to my cry for mercy; in your faithfulness and righteousness come to my relief.
PS|143|2|Do not bring your servant into judgment, for no one living is righteous before you.
PS|143|3|The enemy pursues me, he crushes me to the ground; he makes me dwell in darkness like those long dead.
PS|143|4|So my spirit grows faint within me; my heart within me is dismayed.
PS|143|5|I remember the days of long ago; I meditate on all your works and consider what your hands have done.
PS|143|6|I spread out my hands to you; my soul thirsts for you like a parched land. Selah
PS|143|7|Answer me quickly, O LORD; my spirit fails. Do not hide your face from me or I will be like those who go down to the pit.
PS|143|8|Let the morning bring me word of your unfailing love, for I have put my trust in you. Show me the way I should go, for to you I lift up my soul.
PS|143|9|Rescue me from my enemies, O LORD, for I hide myself in you.
PS|143|10|Teach me to do your will, for you are my God; may your good Spirit lead me on level ground.
PS|143|11|For your name's sake, O LORD, preserve my life; in your righteousness, bring me out of trouble.
PS|143|12|In your unfailing love, silence my enemies; destroy all my foes, for I am your servant.
PS|144|1|Praise be to the LORD my Rock, who trains my hands for war, my fingers for battle.
PS|144|2|He is my loving God and my fortress, my stronghold and my deliverer, my shield, in whom I take refuge, who subdues peoples under me.
PS|144|3|O LORD, what is man that you care for him, the son of man that you think of him?
PS|144|4|Man is like a breath; his days are like a fleeting shadow.
PS|144|5|Part your heavens, O LORD, and come down; touch the mountains, so that they smoke.
PS|144|6|Send forth lightning and scatter {the enemies}; shoot your arrows and rout them.
PS|144|7|Reach down your hand from on high; deliver me and rescue me from the mighty waters, from the hands of foreigners
PS|144|8|whose mouths are full of lies, whose right hands are deceitful.
PS|144|9|I will sing a new song to you, O God; on the ten-stringed lyre I will make music to you,
PS|144|10|to the One who gives victory to kings, who delivers his servant David from the deadly sword.
PS|144|11|Deliver me and rescue me from the hands of foreigners whose mouths are full of lies, whose right hands are deceitful.
PS|144|12|Then our sons in their youth will be like well-nurtured plants, and our daughters will be like pillars carved to adorn a palace.
PS|144|13|Our barns will be filled with every kind of provision. Our sheep will increase by thousands, by tens of thousands in our fields;
PS|144|14|our oxen will draw heavy loads. There will be no breaching of walls, no going into captivity, no cry of distress in our streets.
PS|144|15|Blessed are the people of whom this is true; blessed are the people whose God is the LORD.
PS|145|1|I will exalt you, my God the King; I will praise your name for ever and ever.
PS|145|2|Every day I will praise you and extol your name for ever and ever.
PS|145|3|Great is the LORD and most worthy of praise; his greatness no one can fathom.
PS|145|4|One generation will commend your works to another; they will tell of your mighty acts.
PS|145|5|They will speak of the glorious splendor of your majesty, and I will meditate on your wonderful works.
PS|145|6|They will tell of the power of your awesome works, and I will proclaim your great deeds.
PS|145|7|They will celebrate your abundant goodness and joyfully sing of your righteousness.
PS|145|8|The LORD is gracious and compassionate, slow to anger and rich in love.
PS|145|9|The LORD is good to all; he has compassion on all he has made.
PS|145|10|All you have made will praise you, O LORD; your saints will extol you.
PS|145|11|They will tell of the glory of your kingdom and speak of your might,
PS|145|12|so that all men may know of your mighty acts and the glorious splendor of your kingdom.
PS|145|13|Your kingdom is an everlasting kingdom, and your dominion endures through all generations. The LORD is faithful to all his promises and loving toward all he has made.
PS|145|14|The LORD upholds all those who fall and lifts up all who are bowed down.
PS|145|15|The eyes of all look to you, and you give them their food at the proper time.
PS|145|16|You open your hand and satisfy the desires of every living thing.
PS|145|17|The LORD is righteous in all his ways and loving toward all he has made.
PS|145|18|The LORD is near to all who call on him, to all who call on him in truth.
PS|145|19|He fulfills the desires of those who fear him; he hears their cry and saves them.
PS|145|20|The LORD watches over all who love him, but all the wicked he will destroy.
PS|145|21|My mouth will speak in praise of the LORD. Let every creature praise his holy name for ever and ever.
PS|146|1|Praise the LORD. Praise the LORD, O my soul.
PS|146|2|I will praise the LORD all my life; I will sing praise to my God as long as I live.
PS|146|3|Do not put your trust in princes, in mortal men, who cannot save.
PS|146|4|When their spirit departs, they return to the ground; on that very day their plans come to nothing.
PS|146|5|Blessed is he whose help is the God of Jacob, whose hope is in the LORD his God,
PS|146|6|the Maker of heaven and earth, the sea, and everything in them- the LORD, who remains faithful forever.
PS|146|7|He upholds the cause of the oppressed and gives food to the hungry. The LORD sets prisoners free,
PS|146|8|the LORD gives sight to the blind, the LORD lifts up those who are bowed down, the LORD loves the righteous.
PS|146|9|The LORD watches over the alien and sustains the fatherless and the widow, but he frustrates the ways of the wicked.
PS|146|10|The LORD reigns forever, your God, O Zion, for all generations. Praise the LORD.
PS|147|1|Praise the LORD. How good it is to sing praises to our God, how pleasant and fitting to praise him!
PS|147|2|The LORD builds up Jerusalem; he gathers the exiles of Israel.
PS|147|3|He heals the brokenhearted and binds up their wounds.
PS|147|4|He determines the number of the stars and calls them each by name.
PS|147|5|Great is our Lord and mighty in power; his understanding has no limit.
PS|147|6|The LORD sustains the humble but casts the wicked to the ground.
PS|147|7|Sing to the LORD with thanksgiving; make music to our God on the harp.
PS|147|8|He covers the sky with clouds; he supplies the earth with rain and makes grass grow on the hills.
PS|147|9|He provides food for the cattle and for the young ravens when they call.
PS|147|10|His pleasure is not in the strength of the horse, nor his delight in the legs of a man;
PS|147|11|the LORD delights in those who fear him, who put their hope in his unfailing love.
PS|147|12|Extol the LORD, O Jerusalem; praise your God, O Zion,
PS|147|13|for he strengthens the bars of your gates and blesses your people within you.
PS|147|14|He grants peace to your borders and satisfies you with the finest of wheat.
PS|147|15|He sends his command to the earth; his word runs swiftly.
PS|147|16|He spreads the snow like wool and scatters the frost like ashes.
PS|147|17|He hurls down his hail like pebbles. Who can withstand his icy blast?
PS|147|18|He sends his word and melts them; he stirs up his breezes, and the waters flow.
PS|147|19|He has revealed his word to Jacob, his laws and decrees to Israel.
PS|147|20|He has done this for no other nation; they do not know his laws. Praise the LORD.
PS|148|1|Praise the LORD. Praise the LORD from the heavens, praise him in the heights above.
PS|148|2|Praise him, all his angels, praise him, all his heavenly hosts.
PS|148|3|Praise him, sun and moon, praise him, all you shining stars.
PS|148|4|Praise him, you highest heavens and you waters above the skies.
PS|148|5|Let them praise the name of the LORD, for he commanded and they were created.
PS|148|6|He set them in place for ever and ever; he gave a decree that will never pass away.
PS|148|7|Praise the LORD from the earth, you great sea creatures and all ocean depths,
PS|148|8|lightning and hail, snow and clouds, stormy winds that do his bidding,
PS|148|9|you mountains and all hills, fruit trees and all cedars,
PS|148|10|wild animals and all cattle, small creatures and flying birds,
PS|148|11|kings of the earth and all nations, you princes and all rulers on earth,
PS|148|12|young men and maidens, old men and children.
PS|148|13|Let them praise the name of the LORD, for his name alone is exalted; his splendor is above the earth and the heavens.
PS|148|14|He has raised up for his people a horn, the praise of all his saints, of Israel, the people close to his heart. Praise the LORD.
PS|149|1|Praise the LORD. Sing to the LORD a new song, his praise in the assembly of the saints.
PS|149|2|Let Israel rejoice in their Maker; let the people of Zion be glad in their King.
PS|149|3|Let them praise his name with dancing and make music to him with tambourine and harp.
PS|149|4|For the LORD takes delight in his people; he crowns the humble with salvation.
PS|149|5|Let the saints rejoice in this honor and sing for joy on their beds.
PS|149|6|May the praise of God be in their mouths and a double-edged sword in their hands,
PS|149|7|to inflict vengeance on the nations and punishment on the peoples,
PS|149|8|to bind their kings with fetters, their nobles with shackles of iron,
PS|149|9|to carry out the sentence written against them. This is the glory of all his saints. Praise the LORD.
PS|150|1|Praise the LORD. Praise God in his sanctuary; praise him in his mighty heavens.
PS|150|2|Praise him for his acts of power; praise him for his surpassing greatness.
PS|150|3|Praise him with the sounding of the trumpet, praise him with the harp and lyre,
PS|150|4|praise him with tambourine and dancing, praise him with the strings and flute,
PS|150|5|praise him with the clash of cymbals, praise him with resounding cymbals.
PS|150|6|Let everything that has breath praise the LORD. Praise the LORD.
