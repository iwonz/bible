2COR|1|1|Paulus apostolus Iesu Christi per voluntatem Dei et Timotheus frater ecclesiae Dei quae est Corinthi cum sanctis omnibus qui sunt in universa Achaia
2COR|1|2|gratia vobis et pax a Deo Patre nostro et Domino Iesu Christo
2COR|1|3|benedictus Deus et Pater Domini nostri Iesu Christi Pater misericordiarum et Deus totius consolationis
2COR|1|4|qui consolatur nos in omni tribulatione nostra ut possimus et ipsi consolari eos qui in omni pressura sunt per exhortationem qua exhortamur et ipsi a Deo
2COR|1|5|quoniam sicut abundant passiones Christi in nobis ita et per Christum abundat consolatio nostra
2COR|1|6|sive autem tribulamur pro vestra exhortatione et salute sive exhortamur pro vestra exhortatione quae operatur in tolerantia earundem passionum quas et nos patimur
2COR|1|7|et spes nostra firma pro vobis scientes quoniam sicut socii passionum estis sic eritis et consolationis
2COR|1|8|non enim volumus ignorare vos fratres de tribulatione nostra quae facta est in Asia quoniam supra modum gravati sumus supra virtutem ita ut taederet nos etiam vivere
2COR|1|9|sed ipsi in nobis ipsis responsum mortis habuimus ut non simus fidentes in nobis sed in Deo qui suscitat mortuos
2COR|1|10|qui de tantis periculis eripuit nos et eruet in quem speramus quoniam et adhuc eripiet
2COR|1|11|adiuvantibus et vobis in oratione pro nobis ut ex multis personis eius quae in nobis est donationis per multos gratiae agantur pro nobis
2COR|1|12|nam gloria nostra haec est testimonium conscientiae nostrae quod in simplicitate et sinceritate Dei et non in sapientia carnali sed in gratia Dei conversati sumus in mundo abundantius autem ad vos
2COR|1|13|non enim alia scribimus vobis quam quae legistis et cognoscitis spero autem quod usque in finem cognoscetis
2COR|1|14|sicut et cognovistis nos ex parte quia gloria vestra sumus sicut et vos nostra in die Domini nostri Iesu Christi
2COR|1|15|et hac confidentia volui prius venire ad vos ut secundam gratiam haberetis
2COR|1|16|et per vos transire in Macedoniam et iterum a Macedonia venire ad vos et a vobis deduci in Iudaeam
2COR|1|17|cum hoc ergo voluissem numquid levitate usus sum aut quae cogito secundum carnem cogito ut sit apud me est et non
2COR|1|18|fidelis autem Deus quia sermo noster qui fit apud vos non est in illo est et non
2COR|1|19|Dei enim Filius Iesus Christus qui in vobis per nos praedicatus est per me et Silvanum et Timotheum non fuit est et non sed est in illo fuit
2COR|1|20|quotquot enim promissiones Dei sunt in illo est ideo et per ipsum amen Deo ad gloriam nostram
2COR|1|21|qui autem confirmat nos vobiscum in Christum et qui unxit nos Deus
2COR|1|22|et qui signavit nos et dedit pignus Spiritus in cordibus nostris
2COR|1|23|ego autem testem Deum invoco in animam meam quod parcens vobis non veni ultra Corinthum
2COR|1|24|non quia dominamur fidei vestrae sed adiutores sumus gaudii vestri nam fide stetistis
2COR|2|1|statui autem hoc ipse apud me ne iterum in tristitia venirem ad vos
2COR|2|2|si enim ego contristo vos et quis est qui me laetificet nisi qui contristatur ex me
2COR|2|3|et hoc ipsum scripsi ut non cum venero tristitiam super tristitiam habeam de quibus oportuerat me gaudere confidens in omnibus vobis quia meum gaudium omnium vestrum est
2COR|2|4|nam ex multa tribulatione et angustia cordis scripsi vobis per multas lacrimas non ut contristemini sed ut sciatis quam caritatem habeo abundantius in vobis
2COR|2|5|si quis autem contristavit non me contristavit sed ex parte ut non onerem omnes vos
2COR|2|6|sufficit illi qui eiusmodi est obiurgatio haec quae fit a pluribus
2COR|2|7|ita ut e contra magis donetis et consolemini ne forte abundantiori tristitia absorbeatur qui eiusmodi est
2COR|2|8|propter quod obsecro vos ut confirmetis in illum caritatem
2COR|2|9|ideo enim et scripsi ut cognoscam experimentum vestrum an in omnibus oboedientes sitis
2COR|2|10|cui autem aliquid donatis et ego nam et ego quod donavi si quid donavi propter vos in persona Christi
2COR|2|11|ut non circumveniamur a Satana non enim ignoramus cogitationes eius
2COR|2|12|cum venissem autem Troadem propter evangelium Christi et ostium mihi apertum esset in Domino
2COR|2|13|non habui requiem spiritui meo eo quod non invenerim Titum fratrem meum sed valefaciens eis profectus sum in Macedoniam
2COR|2|14|Deo autem gratias qui semper triumphat nos in Christo Iesu et odorem notitiae suae manifestat per nos in omni loco
2COR|2|15|quia Christi bonus odor sumus Deo in his qui salvi fiunt et in his qui pereunt
2COR|2|16|aliis quidem odor mortis in mortem aliis autem odor vitae in vitam et ad haec quis tam idoneus
2COR|2|17|non enim sumus sicut plurimi adulterantes verbum Dei sed ex sinceritate sed sicut ex Deo coram Deo in Christo loquimur
2COR|3|1|incipimus iterum nosmet ipsos commendare aut numquid egemus sicut quidam commendaticiis epistulis ad vos aut ex vobis
2COR|3|2|epistula nostra vos estis scripta in cordibus nostris quae scitur et legitur ab omnibus hominibus
2COR|3|3|manifestati quoniam epistula estis Christi ministrata a nobis et scripta non atramento sed Spiritu Dei vivi non in tabulis lapideis sed in tabulis cordis carnalibus
2COR|3|4|fiduciam autem talem habemus per Christum ad Deum
2COR|3|5|non quod sufficientes simus cogitare aliquid a nobis quasi ex nobis sed sufficientia nostra ex Deo est
2COR|3|6|qui et idoneos nos fecit ministros novi testamenti non litterae sed Spiritus littera enim occidit Spiritus autem vivificat
2COR|3|7|quod si ministratio mortis litteris deformata in lapidibus fuit in gloria ita ut non possent intendere filii Israhel in faciem Mosi propter gloriam vultus eius quae evacuatur
2COR|3|8|quomodo non magis ministratio Spiritus erit in gloria
2COR|3|9|nam si ministratio damnationis gloria est multo magis abundat ministerium iustitiae in gloria
2COR|3|10|nam nec glorificatum est quod claruit in hac parte propter excellentem gloriam
2COR|3|11|si enim quod evacuatur per gloriam est multo magis quod manet in gloria est
2COR|3|12|habentes igitur talem spem multa fiducia utimur
2COR|3|13|et non sicut Moses ponebat velamen super faciem suam ut non intenderent filii Israhel in faciem eius quod evacuatur
2COR|3|14|sed obtusi sunt sensus eorum usque in hodiernum enim diem id ipsum velamen in lectione veteris testamenti manet non revelatum quoniam in Christo evacuatur
2COR|3|15|sed usque in hodiernum diem cum legitur Moses velamen est positum super cor eorum
2COR|3|16|cum autem conversus fuerit ad Deum aufertur velamen
2COR|3|17|Dominus autem Spiritus est ubi autem Spiritus Domini ibi libertas
2COR|3|18|nos vero omnes revelata facie gloriam Domini speculantes in eandem imaginem transformamur a claritate in claritatem tamquam a Domini Spiritu
2COR|4|1|ideo habentes hanc ministrationem iuxta quod misericordiam consecuti sumus non deficimus
2COR|4|2|sed abdicamus occulta dedecoris non ambulantes in astutia neque adulterantes verbum Dei sed in manifestatione veritatis commendantes nosmet ipsos ad omnem conscientiam hominum coram Deo
2COR|4|3|quod si etiam opertum est evangelium nostrum in his qui pereunt est opertum
2COR|4|4|in quibus deus huius saeculi excaecavit mentes infidelium ut non fulgeat inluminatio evangelii gloriae Christi qui est imago Dei
2COR|4|5|non enim nosmet ipsos praedicamus sed Iesum Christum Dominum nos autem servos vestros per Iesum
2COR|4|6|quoniam Deus qui dixit de tenebris lucem splendescere qui inluxit in cordibus nostris ad inluminationem scientiae claritatis Dei in facie Christi Iesu
2COR|4|7|habemus autem thesaurum istum in vasis fictilibus ut sublimitas sit virtutis Dei et non ex nobis
2COR|4|8|in omnibus tribulationem patimur sed non angustiamur aporiamur sed non destituimur
2COR|4|9|persecutionem patimur sed non derelinquimur deicimur sed non perimus
2COR|4|10|semper mortificationem Iesu in corpore nostro circumferentes ut et vita Iesu in corporibus nostris manifestetur
2COR|4|11|semper enim nos qui vivimus in mortem tradimur propter Iesum ut et vita Iesu manifestetur in carne nostra mortali
2COR|4|12|ergo mors in nobis operatur vita autem in vobis
2COR|4|13|habentes autem eundem spiritum fidei sicut scriptum est credidi propter quod locutus sum et nos credimus propter quod et loquimur
2COR|4|14|scientes quoniam qui suscitavit Iesum et nos cum Iesu suscitabit et constituet vobiscum
2COR|4|15|omnia enim propter vos ut gratia abundans per multos gratiarum actione abundet in gloriam Dei
2COR|4|16|propter quod non deficimus sed licet is qui foris est noster homo corrumpitur tamen is qui intus est renovatur de die in diem
2COR|4|17|id enim quod in praesenti est momentaneum et leve tribulationis nostrae supra modum in sublimitatem aeternum gloriae pondus operatur nobis
2COR|4|18|non contemplantibus nobis quae videntur sed quae non videntur quae enim videntur temporalia sunt quae autem non videntur aeterna sunt
2COR|5|1|scimus enim quoniam si terrestris domus nostra huius habitationis dissolvatur quod aedificationem ex Deo habeamus domum non manufactam aeternam in caelis
2COR|5|2|nam et in hoc ingemescimus habitationem nostram quae de caelo est superindui cupientes
2COR|5|3|si tamen vestiti non nudi inveniamur
2COR|5|4|nam et qui sumus in tabernaculo ingemescimus gravati eo quod nolumus expoliari sed supervestiri ut absorbeatur quod mortale est a vita
2COR|5|5|qui autem efficit nos in hoc ipsum Deus qui dedit nobis pignus Spiritus
2COR|5|6|audentes igitur semper et scientes quoniam dum sumus in corpore peregrinamur a Domino
2COR|5|7|per fidem enim ambulamus et non per speciem
2COR|5|8|audemus autem et bonam voluntatem habemus magis peregrinari a corpore et praesentes esse ad Deum
2COR|5|9|et ideo contendimus sive absentes sive praesentes placere illi
2COR|5|10|omnes enim nos manifestari oportet ante tribunal Christi ut referat unusquisque propria corporis prout gessit sive bonum sive malum
2COR|5|11|scientes ergo timorem Domini hominibus suademus Deo autem manifesti sumus spero autem et in conscientiis vestris manifestos nos esse
2COR|5|12|non iterum nos commendamus vobis sed occasionem damus vobis gloriandi pro nobis ut habeatis ad eos qui in facie gloriantur et non in corde
2COR|5|13|sive enim mente excedimus Deo sive sobrii sumus vobis
2COR|5|14|caritas enim Christi urget nos aestimantes hoc quoniam si unus pro omnibus mortuus est ergo omnes mortui sunt
2COR|5|15|et pro omnibus mortuus est ut et qui vivunt iam non sibi vivant sed ei qui pro ipsis mortuus est et resurrexit
2COR|5|16|itaque nos ex hoc neminem novimus secundum carnem et si cognovimus secundum carnem Christum sed nunc iam non novimus
2COR|5|17|si qua ergo in Christo nova creatura vetera transierunt ecce facta sunt nova
2COR|5|18|omnia autem ex Deo qui reconciliavit nos sibi per Christum et dedit nobis ministerium reconciliationis
2COR|5|19|quoniam quidem Deus erat in Christo mundum reconcilians sibi non reputans illis delicta ipsorum et posuit in nobis verbum reconciliationis
2COR|5|20|pro Christo ergo legationem fungimur tamquam Deo exhortante per nos obsecramus pro Christo reconciliamini Deo
2COR|5|21|eum qui non noverat peccatum pro nobis peccatum fecit ut nos efficeremur iustitia Dei in ipso
2COR|6|1|adiuvantes autem et exhortamur ne in vacuum gratiam Dei recipiatis
2COR|6|2|ait enim tempore accepto exaudivi te et in die salutis adiuvavi te ecce nunc tempus acceptabile ecce nunc dies salutis
2COR|6|3|nemini dantes ullam offensionem ut non vituperetur ministerium
2COR|6|4|sed in omnibus exhibeamus nosmet ipsos sicut Dei ministros in multa patientia in tribulationibus in necessitatibus in angustiis
2COR|6|5|in plagis in carceribus in seditionibus in laboribus in vigiliis in ieiuniis
2COR|6|6|in castitate in scientia in longanimitate in suavitate in Spiritu Sancto in caritate non ficta
2COR|6|7|in verbo veritatis in virtute Dei per arma iustitiae a dextris et sinistris
2COR|6|8|per gloriam et ignobilitatem per infamiam et bonam famam ut seductores et veraces sicut qui ignoti et cogniti
2COR|6|9|quasi morientes et ecce vivimus ut castigati et non mortificati
2COR|6|10|quasi tristes semper autem gaudentes sicut egentes multos autem locupletantes tamquam nihil habentes et omnia possidentes
2COR|6|11|os nostrum patet ad vos o Corinthii cor nostrum dilatatum est
2COR|6|12|non angustiamini in nobis angustiamini autem in visceribus vestris
2COR|6|13|eandem autem habentes remunerationem tamquam filiis dico dilatamini et vos
2COR|6|14|nolite iugum ducere cum infidelibus quae enim participatio iustitiae cum iniquitate aut quae societas luci ad tenebras
2COR|6|15|quae autem conventio Christi ad Belial aut quae pars fideli cum infidele
2COR|6|16|qui autem consensus templo Dei cum idolis vos enim estis templum Dei vivi sicut dicit Deus quoniam inhabitabo in illis et inambulabo et ero illorum Deus et ipsi erunt mihi populus
2COR|6|17|propter quod exite de medio eorum et separamini dicit Dominus et inmundum ne tetigeritis
2COR|6|18|et ego recipiam vos et ero vobis in patrem et vos eritis mihi in filios et filias dicit Dominus omnipotens
2COR|7|1|has igitur habentes promissiones carissimi mundemus nos ab omni inquinamento carnis et spiritus perficientes sanctificationem in timore Dei
2COR|7|2|capite nos neminem laesimus neminem corrupimus neminem circumvenimus
2COR|7|3|non ad condemnationem dico praedixi enim quod in cordibus nostris estis ad conmoriendum et ad convivendum
2COR|7|4|multa mihi fiducia est apud vos multa mihi gloriatio pro vobis repletus sum consolatione superabundo gaudio in omni tribulatione nostra
2COR|7|5|nam et cum venissemus Macedoniam nullam requiem habuit caro nostra sed omnem tribulationem passi foris pugnae intus timores
2COR|7|6|sed qui consolatur humiles consolatus est nos Deus in adventu Titi
2COR|7|7|non solum autem in adventu eius sed etiam in solacio quo consolatus est in vobis referens nobis vestrum desiderium vestrum fletum vestram aemulationem pro me ita ut magis gauderem
2COR|7|8|quoniam et si contristavi vos in epistula non me paenitet et si paeniteret videns quod epistula illa et si ad horam vos contristavit
2COR|7|9|nunc gaudeo non quia contristati estis sed quia contristati estis ad paenitentiam contristati enim estis secundum Deum ut in nullo detrimentum patiamini ex nobis
2COR|7|10|quae enim secundum Deum tristitia est paenitentiam in salutem stabilem operatur saeculi autem tristitia mortem operatur
2COR|7|11|ecce enim hoc ipsum secundum Deum contristari vos quantam in vobis operatur sollicitudinem sed defensionem sed indignationem sed timorem sed desiderium sed aemulationem sed vindictam in omnibus exhibuistis vos incontaminatos esse negotio
2COR|7|12|igitur et si scripsi vobis non propter eum qui fecit iniuriam nec propter eum qui passus est sed ad manifestandam sollicitudinem nostram quam pro vobis habemus ad vos coram Deo
2COR|7|13|ideo consolati sumus in consolatione autem nostra abundantius magis gavisi sumus super gaudium Titi quia refectus est spiritus eius ab omnibus vobis
2COR|7|14|et si quid apud illum de vobis gloriatus sum non sum confusus sed sicut omnia vobis in veritate locuti sumus ita et gloriatio nostra quae fuit ad Titum veritas facta est
2COR|7|15|et viscera eius abundantius in vos sunt reminiscentis omnium vestrum oboedientiam quomodo cum timore et tremore excepistis eum
2COR|7|16|gaudeo quod in omnibus confido in vobis
2COR|8|1|notam autem facimus vobis fratres gratiam Dei quae data est in ecclesiis Macedoniae
2COR|8|2|quod in multo experimento tribulationis abundantia gaudii ipsorum et altissima paupertas eorum abundavit in divitias simplicitatis eorum
2COR|8|3|quia secundum virtutem testimonium illis reddo et supra virtutem voluntarii fuerunt
2COR|8|4|cum multa exhortatione obsecrantes nos gratiam et communicationem ministerii quod fit in sanctos
2COR|8|5|et non sicut speravimus sed semet ipsos dederunt primum Domino deinde nobis per voluntatem Dei
2COR|8|6|ita ut rogaremus Titum ut quemadmodum coepit ita et perficiat in vos etiam gratiam istam
2COR|8|7|sed sicut in omnibus abundatis fide et sermone et scientia et omni sollicitudine et caritate vestra in nos ut et in hac gratia abundetis
2COR|8|8|non quasi imperans dico sed per aliorum sollicitudinem etiam vestrae caritatis ingenitum bonum conprobans
2COR|8|9|scitis enim gratiam Domini nostri Iesu Christi quoniam propter vos egenus factus est cum esset dives ut illius inopia vos divites essetis
2COR|8|10|et consilium in hoc do hoc enim vobis utile est qui non solum facere sed et velle coepistis ab anno priore
2COR|8|11|nunc vero et facto perficite ut quemadmodum promptus est animus voluntatis ita sit et perficiendi ex eo quod habetis
2COR|8|12|si enim voluntas prompta est secundum id quod habet accepta est non secundum quod non habet
2COR|8|13|non enim ut aliis sit remissio vobis autem tribulatio sed ex aequalitate
2COR|8|14|in praesenti tempore vestra abundantia illorum inopiam suppleat ut et illorum abundantia vestrae inopiae sit supplementum ut fiat aequalitas sicut scriptum est
2COR|8|15|qui multum non abundavit et qui modicum non minoravit
2COR|8|16|gratias autem Deo qui dedit eandem sollicitudinem pro vobis in corde Titi
2COR|8|17|quoniam exhortationem quidem suscepit sed cum sollicitior esset sua voluntate profectus est ad vos
2COR|8|18|misimus etiam cum illo fratrem cuius laus est in evangelio per omnes ecclesias
2COR|8|19|non solum autem sed et ordinatus ab ecclesiis comes peregrinationis nostrae in hac gratia quae ministratur a nobis ad Domini gloriam et destinatam voluntatem nostram
2COR|8|20|devitantes hoc ne quis nos vituperet in hac plenitudine quae ministratur a nobis
2COR|8|21|providemus enim bona non solum coram Deo sed etiam coram hominibus
2COR|8|22|misimus autem cum illis et fratrem nostrum quem probavimus in multis saepe sollicitum esse nunc autem multo sollicitiorem confidentia multa in vos
2COR|8|23|sive pro Tito qui est socius meus et in vos adiutor sive fratres nostri apostoli ecclesiarum gloriae Christi
2COR|8|24|ostensionem ergo quae est caritatis vestrae et nostrae gloriae pro vobis in illos ostendite in faciem ecclesiarum
2COR|9|1|nam de ministerio quod fit in sanctos ex abundanti est mihi scribere vobis
2COR|9|2|scio enim promptum animum vestrum pro quo de vobis glorior apud Macedonas quoniam Achaia parata est ab anno praeterito et vestra aemulatio provocavit plurimos
2COR|9|3|misi autem fratres ut ne quod gloriamur de vobis evacuetur in hac parte ut quemadmodum dixi parati sitis
2COR|9|4|ne cum venerint mecum Macedones et invenerint vos inparatos erubescamus nos ut non dicamus vos in hac substantia
2COR|9|5|necessarium ergo existimavi rogare fratres ut praeveniant ad vos et praeparent repromissam benedictionem hanc paratam esse sic quasi benedictionem non quasi avaritiam
2COR|9|6|hoc autem qui parce seminat parce et metet et qui seminat in benedictionibus de benedictionibus et metet
2COR|9|7|unusquisque prout destinavit corde suo non ex tristitia aut ex necessitate hilarem enim datorem diligit Deus
2COR|9|8|potens est autem Deus omnem gratiam abundare facere in vobis ut in omnibus semper omnem sufficientiam habentes abundetis in omne opus bonum
2COR|9|9|sicut scriptum est dispersit dedit pauperibus iustitia eius manet in aeternum
2COR|9|10|qui autem administrat semen seminanti et panem ad manducandum praestabit et multiplicabit semen vestrum et augebit incrementa frugum iustitiae vestrae
2COR|9|11|ut in omnibus locupletati abundetis in omnem simplicitatem quae operatur per nos gratiarum actionem Deo
2COR|9|12|quoniam ministerium huius officii non solum supplet ea quae desunt sanctis sed etiam abundat per multas gratiarum actiones in Domino
2COR|9|13|per probationem ministerii huius glorificantes Deum in oboedientia confessionis vestrae in evangelium Christi et simplicitate communicationis in illos et in omnes
2COR|9|14|et ipsorum obsecratione pro vobis desiderantium vos propter eminentem gratiam Dei in vobis
2COR|9|15|gratias Deo super inenarrabili dono eius
2COR|10|1|ipse autem ego Paulus obsecro vos per mansuetudinem et modestiam Christi qui in facie quidem humilis inter vos absens autem confido in vobis
2COR|10|2|rogo autem ne praesens audeam per eam confidentiam qua existimo audere in quosdam qui arbitrantur nos tamquam secundum carnem ambulemus
2COR|10|3|in carne enim ambulantes non secundum carnem militamus
2COR|10|4|nam arma militiae nostrae non carnalia sed potentia Deo ad destructionem munitionum consilia destruentes
2COR|10|5|et omnem altitudinem extollentem se adversus scientiam Dei et in captivitatem redigentes omnem intellectum in obsequium Christi
2COR|10|6|et in promptu habentes ulcisci omnem inoboedientiam cum impleta fuerit vestra oboedientia
2COR|10|7|quae secundum faciem sunt videte si quis confidit sibi Christi se esse hoc cogitet iterum apud se quia sicut ipse Christi est ita et nos
2COR|10|8|nam et si amplius aliquid gloriatus fuero de potestate nostra quam dedit Dominus in aedificationem et non in destructionem vestram non erubescam
2COR|10|9|ut autem non existimer tamquam terrere vos per epistulas
2COR|10|10|quoniam quidem epistulae inquiunt graves sunt et fortes praesentia autem corporis infirma et sermo contemptibilis
2COR|10|11|hoc cogitet qui eiusmodi est quia quales sumus verbo per epistulas absentes tales et praesentes in facto
2COR|10|12|non enim audemus inserere aut conparare nos quibusdam qui se ipsos commendant sed ipsi in nobis nosmet ipsos metientes et conparantes nosmet ipsos nobis
2COR|10|13|nos autem non in inmensum gloriabimur sed secundum mensuram regulae quam mensus est nobis Deus mensuram pertingendi usque ad vos
2COR|10|14|non enim quasi non pertingentes ad vos superextendimus nos usque ad vos enim pervenimus in evangelio Christi
2COR|10|15|non in inmensum gloriantes in alienis laboribus spem autem habentes crescentis fidei vestrae in vobis magnificari secundum regulam nostram in abundantiam
2COR|10|16|etiam in illa quae ultra vos sunt evangelizare non in aliena regula in his quae praeparata sunt gloriari
2COR|10|17|qui autem gloriatur in Domino glorietur
2COR|10|18|non enim qui se ipsum commendat ille probatus est sed quem Dominus commendat
2COR|11|1|utinam sustineretis modicum quid insipientiae meae sed et subportate me
2COR|11|2|aemulor enim vos Dei aemulatione despondi enim vos uni viro virginem castam exhibere Christo
2COR|11|3|timeo autem ne sicut serpens Evam seduxit astutia sua ita corrumpantur sensus vestri et excidant a simplicitate quae est in Christo
2COR|11|4|nam si is qui venit alium Christum praedicat quem non praedicavimus aut alium spiritum accipitis quem non accepistis aut aliud evangelium quod non recepistis recte pateremini
2COR|11|5|existimo enim nihil me minus fecisse magnis apostolis
2COR|11|6|et si inperitus sermone sed non scientia in omnibus autem manifestatus sum vobis
2COR|11|7|aut numquid peccatum feci me ipsum humilians ut vos exaltemini quoniam gratis evangelium Dei evangelizavi vobis
2COR|11|8|alias ecclesias expoliavi accipiens stipendium ad ministerium vestrum
2COR|11|9|et cum essem apud vos et egerem nulli onerosus fui nam quod mihi deerat suppleverunt fratres qui venerunt a Macedonia et in omnibus sine onere me vobis servavi et servabo
2COR|11|10|est veritas Christi in me quoniam haec gloria non infringetur in me in regionibus Achaiae
2COR|11|11|quare quia non diligo vos Deus scit
2COR|11|12|quod autem facio et faciam ut amputem occasionem eorum qui volunt occasionem ut in quo gloriantur inveniantur sicut et nos
2COR|11|13|nam eiusmodi pseudoapostoli operarii subdoli transfigurantes se in apostolos Christi
2COR|11|14|et non mirum ipse enim Satanas transfigurat se in angelum lucis
2COR|11|15|non est ergo magnum si ministri eius transfigurentur velut ministri iustitiae quorum finis erit secundum opera ipsorum
2COR|11|16|iterum dico ne quis me putet insipientem alioquin velut insipientem accipite me ut et ego modicum quid glorier
2COR|11|17|quod loquor non loquor secundum Dominum sed quasi in insipientia in hac substantia gloriae
2COR|11|18|quoniam multi gloriantur secundum carnem et ego gloriabor
2COR|11|19|libenter enim suffertis insipientes cum sitis ipsi sapientes
2COR|11|20|sustinetis enim si quis vos in servitutem redigit si quis devorat si quis accipit si quis extollitur si quis in faciem vos caedit
2COR|11|21|secundum ignobilitatem dico quasi nos infirmi fuerimus in quo quis audet in insipientia dico audeo et ego
2COR|11|22|Hebraei sunt et ego Israhelitae sunt et ego semen Abrahae sunt et ego
2COR|11|23|ministri Christi sunt minus sapiens dico plus ego in laboribus plurimis in carceribus abundantius in plagis supra modum in mortibus frequenter
2COR|11|24|a Iudaeis quinquies quadragenas una minus accepi
2COR|11|25|ter virgis caesus sum semel lapidatus sum ter naufragium feci nocte et die in profundo maris fui
2COR|11|26|in itineribus saepe periculis fluminum periculis latronum periculis ex genere periculis ex gentibus periculis in civitate periculis in solitudine periculis in mari periculis in falsis fratribus
2COR|11|27|in labore et aerumna in vigiliis multis in fame et siti in ieiuniis multis in frigore et nuditate
2COR|11|28|praeter illa quae extrinsecus sunt instantia mea cotidiana sollicitudo omnium ecclesiarum
2COR|11|29|quis infirmatur et non infirmor quis scandalizatur et ego non uror
2COR|11|30|si gloriari oportet quae infirmitatis meae sunt gloriabor
2COR|11|31|Deus et Pater Domini Iesu scit qui est benedictus in saecula quod non mentior
2COR|11|32|Damasci praepositus gentis Aretae regis custodiebat civitatem Damascenorum ut me conprehenderet
2COR|11|33|et per fenestram in sporta dimissus sum per murum et effugi manus eius
2COR|12|1|si gloriari oportet non expedit quidem veniam autem ad visiones et revelationes Domini
2COR|12|2|scio hominem in Christo ante annos quattuordecim sive in corpore nescio sive extra corpus nescio Deus scit raptum eiusmodi usque ad tertium caelum
2COR|12|3|et scio huiusmodi hominem sive in corpore sive extra corpus nescio Deus scit
2COR|12|4|quoniam raptus est in paradisum et audivit arcana verba quae non licet homini loqui
2COR|12|5|pro eiusmodi gloriabor pro me autem nihil gloriabor nisi in infirmitatibus meis
2COR|12|6|nam et si voluero gloriari non ero insipiens veritatem enim dicam parco autem ne quis in me existimet supra id quod videt me aut audit ex me
2COR|12|7|et ne magnitudo revelationum extollat me datus est mihi stimulus carnis meae angelus Satanae ut me colaphizet
2COR|12|8|propter quod ter Dominum rogavi ut discederet a me
2COR|12|9|et dixit mihi sufficit tibi gratia mea nam virtus in infirmitate perficitur libenter igitur gloriabor in infirmitatibus meis ut inhabitet in me virtus Christi
2COR|12|10|propter quod placeo mihi in infirmitatibus in contumeliis in necessitatibus in persecutionibus in angustiis pro Christo cum enim infirmor tunc potens sum
2COR|12|11|factus sum insipiens vos me coegistis ego enim debui a vobis commendari nihil enim minus fui ab his qui sunt supra modum apostoli tametsi nihil sum
2COR|12|12|signa tamen apostoli facta sunt super vos in omni patientia signis et prodigiis et virtutibus
2COR|12|13|quid est enim quod minus habuistis prae ceteris ecclesiis nisi quod ego ipse non gravavi vos donate mihi hanc iniuriam
2COR|12|14|ecce tertio hoc paratus sum venire ad vos et non ero gravis vobis non enim quaero quae vestra sunt sed vos nec enim debent filii parentibus thesaurizare sed parentes filiis
2COR|12|15|ego autem libentissime inpendam et superinpendar ipse pro animabus vestris licet plus vos diligens minus diligar
2COR|12|16|sed esto ego vos non gravavi sed cum essem astutus dolo vos cepi
2COR|12|17|numquid per aliquem eorum quos misi ad vos circumveni vos
2COR|12|18|rogavi Titum et misi cum illo fratrem numquid Titus vos circumvenit nonne eodem spiritu ambulavimus nonne hisdem vestigiis
2COR|12|19|olim putatis quod excusemus nos apud vos coram Deo in Christo loquimur omnia autem carissimi propter vestram aedificationem
2COR|12|20|timeo enim ne forte cum venero non quales volo inveniam vos et ego inveniar a vobis qualem non vultis ne forte contentiones aemulationes animositates dissensiones detractiones susurrationes inflationes seditiones sint inter vos
2COR|12|21|ne iterum cum venero humiliet me Deus apud vos et lugeam multos ex his qui ante peccaverunt et non egerunt paenitentiam super inmunditia et fornicatione et inpudicitia quam gesserunt
2COR|13|1|ecce tertio hoc venio ad vos in ore duorum vel trium testium stabit omne verbum
2COR|13|2|praedixi et praedico ut praesens bis et nunc absens his qui ante peccaverunt et ceteris omnibus quoniam si venero iterum non parcam
2COR|13|3|an experimentum quaeritis eius qui in me loquitur Christi qui in vos non infirmatur sed potens est in vobis
2COR|13|4|nam et si crucifixus est ex infirmitate sed vivit ex virtute Dei nam et nos infirmi sumus in illo sed vivemus cum eo ex virtute Dei in vobis
2COR|13|5|vosmet ipsos temptate si estis in fide ipsi vos probate an non cognoscitis vos ipsos quia Christus Iesus in vobis est nisi forte reprobi estis
2COR|13|6|spero autem quod cognoscetis quia nos non sumus reprobi
2COR|13|7|oramus autem Deum ut nihil mali faciatis non ut nos probati pareamus sed ut vos quod bonum est faciatis nos autem ut reprobi simus
2COR|13|8|non enim possumus aliquid adversus veritatem sed pro veritate
2COR|13|9|gaudemus enim quando nos infirmi sumus vos autem potentes estis hoc et oramus vestram consummationem
2COR|13|10|ideo haec absens scribo ut non praesens durius agam secundum potestatem quam Dominus dedit mihi in aedificationem et non in destructionem
2COR|13|11|de cetero fratres gaudete perfecti estote exhortamini idem sapite pacem habete et Deus dilectionis et pacis erit vobiscum
2COR|13|12|salutate invicem in osculo sancto salutant vos sancti omnes
2COR|13|13|gratia Domini nostri Iesu Christi et caritas Dei et communicatio Sancti Spiritus cum omnibus vobis amen
