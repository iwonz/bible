MIC|1|1|Verbum Domini, quod factum est ad Michaeam Morasthiten in diebus Ioatham, Achaz, Ezechiae regum Iudae, quod vidit super Samariam et Ierusalem.
MIC|1|2|Audite, populi omnes,et attendat terra et plenitudo eius;et sit Dominus Deus vobis in testem,Dominus de templo sancto suo.
MIC|1|3|Quia ecce Dominus egreditur de loco suoet descendet et calcabitsuper excelsa terrae;
MIC|1|4|et liquescent montes subtus eum,et valles scindentursicut cera a facie ignis,sicut aquae, quae decurrunt in praeceps.
MIC|1|5|In scelere Iacob omne istudet in peccatis domus Israel.Quod scelus Iacob?Nonne Samaria?Et quae excelsa Iudae?Nonne Ierusalem?
MIC|1|6|Et ponam Samariam in acervum lapidum,in agrum, ubi plantatur vinea;et detraham in vallem lapides eiuset fundamenta eius revelabo.
MIC|1|7|Et omnia sculptilia eius concidentur,et omnes mercedes eius comburentur igne,et omnia idola eius ponam in perditionem,quia de mercedibus meretricis congregata suntet usque ad mercedem meretricis revertentur.
MIC|1|8|Super hoc plangam et ululabo;vadam spoliatus et nudus,faciam planctum velut thoumet luctum quasi struthionum,
MIC|1|9|quia desperata est plaga eius,quia venit usque ad Iudam,tetigit portam populi meiusque ad Ierusalem.
MIC|1|10|In Geth nolite annuntiare,lacrimis ne ploretis,in Bethleaphra in pulvere volutamini.
MIC|1|11|Et transite vobis, habitatores Saphir,confusi ignominia;non sunt egressi habitatores Saanan.Planctus Betheselauferet a vobis mansionem suam.
MIC|1|12|Profecto trement de bonohabitatores Maroth,quia descendit malum a Dominoin portam Ierusalem.
MIC|1|13|Iungite quadrigae equos, habitatores Lachis;principium peccati est filiae Sion,quia in te inventa sunt scelera Israel.
MIC|1|14|Propterea dabis dimissionemsuper Moresethgeth.Domus Achzib in deceptionemregibus Israel.
MIC|1|15|Adhuc expugnatorem adducam tibi,quae habitas in Maresa;usque Odollam venietgloria Israel.
MIC|1|16|Decalvare et tonderesuper filios deliciarum tuarum;dilata calvitium tuum sicut aquila, quoniam captivi ducti sunt ex te.
MIC|2|1|Vae, qui cogitant iniquitatemet operantur malum in cubilibus suis!In luce matutina faciunt illud,quoniam est in potestate manus eorum.
MIC|2|2|Concupiscunt agros, et violenter tollunt,domos, et rapiunt.Et opprimunt virum et domum eius,hominem et hereditatem eius.
MIC|2|3|Idcirco haec dicit Dominus: Ecce ego cogitosuper familiam istam malum,unde non auferetiscolla vestra;et non ambulabitis erecti,quoniam tempus pessimum est.
MIC|2|4|In die illasumetur super vos parabola,et assumetur lamentum dicentium: "Depopulatione vastati sumus;pars populi mei commutatur,quam nemo ei restituet;infideli regiones nostrae dividuntur".
MIC|2|5|Propter hoc non erit tibimittens funiculum sortisin coetu Domini ".
MIC|2|6|" Ne vaticinemini! ". " Vaticinentur,non vaticinentur de his,non cedet confusio! ".
MIC|2|7|Numquid maledicta est domus Iacob?Numquid abbreviatus est spiritus Domini,aut tales sunt actiones eius?Nonne verba eius bona suntcum eo, qui recte graditur?
MIC|2|8|Vos autem contra populum meumut adversarium consurgitis.Desuper tunica pallium tollitis ei;qui transibant fiducialiter,fiunt quasi bello capti.
MIC|2|9|Mulieres populi mei eicitisde domo deliciarum suarum;a parvulis earum aufertisdecorem meum in perpetuum.
MIC|2|10|" Surgite et ite,quia non habetis hic requiem! ".Propter immunditiam peribitisperditione pessima.
MIC|2|11|Si esset vir vento excitatuset mendacium loqueretur: Vaticinabor tibi de vino et sicera ",hic esset vates populi istius.
MIC|2|12|Congregatione congregabo, Iacob, totum te;in unum conducam reliquias Israel,pariter ponam illum quasi gregem in ovili,quasi pecus in medio pascuae;et tumultuabuntur a multitudine hominum.
MIC|2|13|Ascendet enim pandens iter ante eos;erumpent et transibunt portam, egredientur per eam.Et transibit rex eorum coram eis,et Dominus in capite eorum.
MIC|3|1|Et dixi: Audite, principes Iacobet duces domus Israel:Numquid non vestrum est scire iudicium? ".
MIC|3|2|Sed odio habetis bonum et diligitis malum.Violenter tollitis pelles eorum desuper eoset carnem eorum desuper ossibus eorum.
MIC|3|3|Qui comedunt carnem populi meiet pellem eorum desuper excoriant; et ossa eorum confringuntet secant sicut carnem assam in lebeteet quasi carnem in medio ollae.
MIC|3|4|Tunc clamabunt ad Dominum,et non exaudiet eoset abscondet faciem suam ab eisin tempore illo,sicut pessima fecerunt opera sua.
MIC|3|5|Haec dicit Dominus super prophetas,qui seducunt populum meum,qui cum habent, quid mordeant dentibus suis,praedicant pacem;et, si quis non dederit in ore eorum quippiam,sanctificant super eum proelium.
MIC|3|6|Propterea nox vobis sine visione erit,et tenebrae vobis sine divinatione; et occumbet sol super prophetas,et obtenebrabitur super eos dies.
MIC|3|7|Et confundentur videntes,et confundentur divini,et operient labia sua omnes,quia non est responsum Dei.
MIC|3|8|Verumtamen ego repletus sumfortitudine spiritus Domini,iudicio et virtute,ut annuntiem Iacob scelus suumet Israel peccatum suum.
MIC|3|9|Audite hoc, principes domus Iacobet iudices domus Israel,qui abominamini iudiciumet omnia recta pervertitis,
MIC|3|10|qui aedificatis Sion in sanguinibuset Ierusalem in iniquitate.
MIC|3|11|Principes eius in muneribus iudicant,et sacerdotes eius in mercede docent,et prophetae eius in pecunia divinant;et super Dominum requiescunt dicentes: Numquid non Dominus in medio nostrum?Non venient super nos mala ".
MIC|3|12|Propter hoc causa vestriSion quasi ager arabitur,et Ierusalem quasi acervus lapidum erit,et mons templi in excelsa silvarum.
MIC|4|1|Et erit in novissimis diebus:Erit mons domus Dominipraeparatus in vertice montiumet sublimis super colles;et fluent ad eum populi.
MIC|4|2|Et properabunt gentes multae et dicent: Venite, ascendamus ad montem Dominiet ad domum Dei Iacob,et docebit nos de viis suis,et ibimus in semitis eius ";quia de Sion egredietur lex,et verbum Domini de Ierusalem.
MIC|4|3|Et iudicabit inter populos multoset decernet gentibus fortibus usque in longinquum;et concident gladios suos in vomereset hastas suas in falces;non sumet gens adversus gentem gladium,et non discent ultra belligerare.
MIC|4|4|Et sedebit unusquisque subtus vitem suamet subtus ficum suam,et non erit qui deterreat;quia os Domini exercituum locutum est.
MIC|4|5|Quia omnes populi ambulabuntunusquisque in nomine dei sui;nos autem ambulabimus in nomine DominiDei nostri in aeternum et ultra.
MIC|4|6|" In die illa, dicit Dominus,congregabo claudicantem,et eam, quam eieceram, colligamet quam afflixeram;
MIC|4|7|et ponam claudicantem in reliquiaset eam, quae laboraverat, in gentem robustam ".Et regnabit Dominus super eos in monte Sionex hoc nunc et usque in aeternum.
MIC|4|8|Et tu, turris gregis,collis filiae Sion,usque ad te veniet et pervenietpotestas prima,regnum filiae Ierusalem.
MIC|4|9|Nunc quare clamas clamore magno?Numquid rex non est in te,aut consiliarius tuus periit,quia comprehendit te dolor sicut parturientem?
MIC|4|10|Dole et satage,filia Sion, quasi parturiens;quia nunc egredieris de civitateet habitabis in campoet venies usque ad Babylonem;ibi liberaberis,ibi redimet te Dominusde manu inimicorum tuorum.
MIC|4|11|Nunc autem congregatae sunt super tegentes multae,quae dicunt: "Profanetur,et aspiciat in Sion oculus noster ".
MIC|4|12|Ipsi autem non cognoveruntcogitationes Dominiet non intellexerunt consilium eius,quia congregavit eos quasi manipulos in area.
MIC|4|13|Surge et tritura, filia Sion,quia cornu tuum ponam ferreumet ungulas tuas ponam aereas,et comminues populos multoset vovebis Domino rapinas eorumet divitias eorum Domino universae terrae.
MIC|4|14|Nunc incide te, filia incisionis!Obsidionem posuerunt super nos;in virga percutiuntmaxillam iudicis Israel.
MIC|5|1|Sed tu, Bethlehem Ephratha,parvulus in milibus Iudae,ex te mihi egredietur,qui sit dominator in Israel;et egressus eius a temporibus antiquis,a diebus aeternitatis.
MIC|5|2|Propter hoc dabit eosusque ad tempus, in quo parturiens pariet;et reliquiae fratrum eiusconvertentur ad filios Israel.
MIC|5|3|Et stabit et pascet in fortitudine Domini,in sublimitate nominis Domini Dei sui;et habitabunt secure, quia nunc magnus eritusque ad terminos terrae,
MIC|5|4|et erit iste pax.Assyrius cum venerit in terram nostramet quando calcaverit in domibus nostris,suscitabimus super eum septem pastoreset octo primates hominum.
MIC|5|5|Et pascent terram Assyriae in gladio et terram Nemrod in lanceis;et liberabit ab Assyrio,cum venerit in terram nostramet cum calcaverit in finibus nostris.
MIC|5|6|Et erunt reliquiae Iacobin medio populorum multorumquasi ros a Dominoet quasi imbres super herbam,quae non exspectat virumet non praestolatur filios homi num.
MIC|5|7|Et erunt reliquiae Iacob in gentibus,in medio populorum multorum,quasi leo in iumentis silvarumet quasi catulus leonis in gregibus pecorum;qui cum transierit et conculcaverit et ceperit,non est qui eruat.
MIC|5|8|Exaltabitur manus tua super hostes tuos,et omnes inimici tui interibunt.
MIC|5|9|"Et erit in die illa,dicit Dominus,auferam equos tuos de medio tuiet disperdam quadrigas tuas
MIC|5|10|et perdam civitates terrae tuaeet destruam omnes munitiones tuas.
MIC|5|11|Et auferam veneficia de manu tua,et divini non erunt in te.
MIC|5|12|Et perire faciam sculptilia tuaet lapides tuos de medio tui,et non adorabis ultraopera manuum tuarum;
MIC|5|13|et evellam palos tuos de medio tuiet conteram idola tua.
MIC|5|14|Et faciam in furoreet in indignatione ultionemin omnibus gentibus,quae non audierunt ".
MIC|6|1|Audite, quae Dominus loqui tur: Surge, contende iudicio coram montibus,et audiant colles vocem tuam ".
MIC|6|2|Audite, montes, iudicium Domini,et auscultate, fundamenta terrae;quia iudicium Domini cum populo suo,et cum Israel iudicio contendit.
MIC|6|3|" Popule meus, quid feci tibiet quid molestus fui tibi?Responde mihi.
MIC|6|4|Ego eduxi te de terra Aegyptiet de domo servientium liberavi teet misi ante faciem tuam Moysenet Aaron et Mariam.
MIC|6|5|Popule meus, memento, quaeso,quid cogitaverit Balac rex Moab,et quid responderit ei Balaam filius Beor,de Settim usque ad Galgalam,ut cognoscas iustitias Domini ".
MIC|6|6|" Quid dignum offeram Domino,dum curvo genu Deo excelso?Numquid offeram ei holocautomataet vitulos anniculos?
MIC|6|7|Numquid placebunt Domino milia arietum,multa milia torrentium olei?Numquid dabo primogenitum meum pro scelere meo,fructum ventris mei pro peccato animae meae?".
MIC|6|8|Indicatum est tibi, o homo, quid sit bonum,et quid Dominus quaerat a te:utique facere iudicium et diligere caritatemet sollicitum ambulare cum Deo tuo.
MIC|6|9|Vox Domini ad civitatem clamat et sapientia est timere nomen tuum -: Audite, tribus et coetus civitatis!
MIC|6|10|Numquid tolerabo batum iniquumet ephi minus maledictum?
MIC|6|11|Numquid iustificabo stateram impiamet saccelli pondera dolosa?
MIC|6|12|Quia divites eius repleti sunt iniquitate,et habitantes in ea loquebantur mendacium,et lingua eorum fraudulenta in ore eorum.
MIC|6|13|Ego ergo coepi percutere teperditione super peccatis tuis.
MIC|6|14|Tu comedes et non saturaberis,et sordes tuae in medio tui.Tu removebis et non salvabis;et, quos salvaveris, in gladium dabo.
MIC|6|15|Tu seminabis et non metes,tu calcabis olivam et non ungeris oleo,mustum et non bibes vinum.
MIC|6|16|Custodisti praecepta Amriet omne opus domus Achab;et ambulasti in voluntatibus eorum,ut darem te in perditionemet habitantes tuos in sibilum:et opprobrium populorum portabitis ".
MIC|7|1|Vae mihi, quia factum est mihisicut congregata messe,sicut collecta vindemia!Non est botrus ad comedendum,nec praecoqua ficus, quam desideravit anima mea.
MIC|7|2|Periit pius de terra,et rectus in hominibus non est;omnes in sanguine insidiantur,vir fratrem suum rete venatur.
MIC|7|3|Ad malum manus eorum paratae sunt;princeps postulat,et iudex est pro mercede,et magnus manifestat desiderium animae suae;vae eis, qui pervertunt illud!
MIC|7|4|Qui optimus in eis, est quasi paliurus,et, qui rectus, quasi spina de saepe; dies speculatorum tuorum, visitatio tua venit:nunc erit confusio eorum.
MIC|7|5|Nolite credere amico,nolite confidere in proximo;ab ea, quae dormit in sinu tuo,custodi claustra oris tui;
MIC|7|6|quia filius contumeliam facit patri,filia consurgit adversus matrem suam,nurus adversus socrum suam:inimici hominis domestici eius.
MIC|7|7|Ego autem ad Dominum aspiciam,exspectabo Deum salvatorem meum; audiet me Deus meus.
MIC|7|8|Ne laeteris, inimica mea, super mequia cecidi: consurgam;cum sedeo in tenebris,Dominus lux mea est.
MIC|7|9|Iram Domini porto,quoniam peccavi ei,donec iudicet causam meamet faciat iudicium meum;educet me in lucem,videbo iustitiam eius.
MIC|7|10|Et aspiciet inimica meaet operietur confusione,quae dicit ad me: Ubi est Dominus Deus tuus? ".Oculi mei videbunt in eam;nunc erit in conculcationemut lutum platearum.
MIC|7|11|Dies veniet ut aedificentur maceriae tuae;in die illa dilatabuntur fines tui.
MIC|7|12|In die illa usque ad te venienthabitantes ab Assyria usque ad Aegyptumet ab Aegypto usque ad flumenet a mari usque ad mareet a monte usque ad montem.
MIC|7|13|Terra autem erit in desolationempropter habitatores suoset propter fructum operum eorum.
MIC|7|14|Pasce populum tuum in virga tua,gregem hereditatis tuae,habitantes solos in saltu,in medio hortorum;pascantur Basan et Galaadiuxta dies antiquos.
MIC|7|15|Secundum dies egressionis tuae de terra Aegyptiostende nobis mirabilia.
MIC|7|16|Videbunt gentes et confundentursuper omni fortitudine sua,ponent manum super os,aures eorum surdae erunt;
MIC|7|17|lingent pulverem sicut serpens,velut reptilia terrae.Trementes exibunt de aedibus suis " ad Dominum Deum nostrum "formidabunt et timebunt te.
MIC|7|18|Quis Deus similis tui,qui aufers iniquitatemet transis peccatumreliquiarum hereditatis tuae?Non servat in aeternum furorem suum,quoniam volens misericordiam est.
MIC|7|19|Revertetur et miserebitur nostri,calcabit iniquitates nostraset proiciet in profundum marisomnia peccata nostra.
MIC|7|20|Dabis veritatem Iacob,misericordiam Abraham,quae iurasti patribus nostrisa diebus antiquis.
