2SAM|1|1|factum est autem postquam mortuus est Saul ut David reverteretur a caede Amalech et maneret in Siceleg dies duos
2SAM|1|2|in die autem tertia apparuit homo veniens de castris Saul veste conscissa et pulvere aspersus caput et ut venit ad David cecidit super faciem suam et adoravit
2SAM|1|3|dixitque ad eum David unde venis qui ait ad eum de castris Israhel fugi
2SAM|1|4|et dixit ad eum David quod est verbum quod factum est indica mihi qui ait fugit populus e proelio et multi corruentes e populo mortui sunt sed et Saul et Ionathan filius eius interierunt
2SAM|1|5|dixitque David ad adulescentem qui nuntiabat unde scis quia mortuus est Saul et Ionathan filius eius
2SAM|1|6|ait adulescens qui narrabat ei casu veni in montem Gelboe et Saul incumbebat super hastam suam porro currus et equites adpropinquabant ei
2SAM|1|7|et conversus post tergum suum vidensque me vocavit cui cum respondissem adsum
2SAM|1|8|dixit mihi quisnam es tu et aio ad eum Amalechites sum
2SAM|1|9|et locutus est mihi sta super me et interfice me quoniam tenent me angustiae et adhuc tota anima in me est
2SAM|1|10|stansque super eum occidi illum sciebam enim quod vivere non poterat post ruinam et tuli diadema quod erat in capite eius et armillam de brachio illius et adtuli ad te dominum meum huc
2SAM|1|11|adprehendens autem David vestimenta sua scidit omnesque viri qui erant cum eo
2SAM|1|12|et planxerunt et fleverunt et ieiunaverunt usque ad vesperam super Saul et super Ionathan filium eius et super populum Domini et super domum Israhel quod corruissent gladio
2SAM|1|13|dixitque David ad iuvenem qui nuntiaverat ei unde es qui respondit filius hominis advenae amalechitae ego sum
2SAM|1|14|et ait ad eum David quare non timuisti mittere manum tuam ut occideres christum Domini
2SAM|1|15|vocansque David unum de pueris ait accedens inrue in eum qui percussit illum et mortuus est
2SAM|1|16|et ait ad eum David sanguis tuus super caput tuum os enim tuum locutum est adversum te dicens ego interfeci christum Domini
2SAM|1|17|planxit autem David planctum huiuscemodi super Saul et super Ionathan filium eius
2SAM|1|18|et praecepit ut docerent filios Iuda arcum sicut scriptum est in libro Iustorum
2SAM|1|19|incliti Israhel super montes tuos interfecti sunt quomodo ceciderunt fortes
2SAM|1|20|nolite adnuntiare in Geth neque adnuntietis in conpetis Ascalonis ne forte laetentur filiae Philisthim ne exultent filiae incircumcisorum
2SAM|1|21|montes Gelboe nec ros nec pluviae veniant super vos neque sint agri primitiarum quia ibi abiectus est clypeus fortium clypeus Saul quasi non esset unctus oleo
2SAM|1|22|a sanguine interfectorum ab adipe fortium sagitta Ionathan numquam rediit retrorsum et gladius Saul non est reversus inanis
2SAM|1|23|Saul et Ionathan amabiles et decori in vita sua in morte quoque non sunt divisi aquilis velociores leonibus fortiores
2SAM|1|24|filiae Israhel super Saul flete qui vestiebat vos coccino in deliciis qui praebebat ornamenta aurea cultui vestro
2SAM|1|25|quomodo ceciderunt fortes in proelio Ionathan in excelsis tuis occisus est
2SAM|1|26|doleo super te frater mi Ionathan decore nimis et amabilis super amorem mulierum
2SAM|1|27|quomodo ceciderunt robusti et perierunt arma bellica
2SAM|2|1|igitur post haec consuluit David Dominum dicens num ascendam in unam de civitatibus Iuda et ait Dominus ad eum ascende dixitque David quo ascendam et respondit ei in Hebron
2SAM|2|2|ascendit ergo David et duae uxores eius Ahinoem Iezrahelites et Abigail uxor Nabal Carmeli
2SAM|2|3|sed et viros qui erant cum eo duxit David singulos cum domo sua et manserunt in oppidis Hebron
2SAM|2|4|veneruntque viri Iuda et unxerunt ibi David ut regnaret super domum Iuda et nuntiatum est David quod viri Iabesgalaad sepelissent Saul
2SAM|2|5|misit ergo David nuntios ad viros Iabesgalaad dixitque ad eos benedicti vos Domino qui fecistis misericordiam hanc cum domino vestro Saul et sepelistis eum
2SAM|2|6|et nunc retribuet quidem vobis Dominus misericordiam et veritatem sed et ego reddam gratiam eo quod feceritis verbum istud
2SAM|2|7|confortentur manus vestrae et estote filii fortitudinis licet enim mortuus sit dominus vester Saul tamen me unxit domus Iuda regem sibi
2SAM|2|8|Abner autem filius Ner princeps exercitus Saul tulit Hisboseth filium Saul et circumduxit eum per Castra
2SAM|2|9|regemque constituit super Galaad et super Gesuri et super Iezrahel et super Ephraim et super Beniamin et super Israhel universum
2SAM|2|10|quadraginta annorum erat Hisboseth filius Saul cum regnare coepisset super Israhel et duobus annis regnavit sola autem domus Iuda sequebatur David
2SAM|2|11|et fuit numerus dierum quos commoratus est David imperans in Hebron super domum Iuda septem annorum et sex mensuum
2SAM|2|12|egressusque Abner filius Ner et pueri Hisboseth filii Saul de Castris in Gabaon
2SAM|2|13|porro Ioab filius Sarviae et pueri David egressi sunt et occurrerunt eis iuxta piscinam Gabaon et cum in unum convenissent e regione sederunt hii ex una parte piscinae et illi ex altera
2SAM|2|14|dixitque Abner ad Ioab surgant pueri et ludant coram nobis et respondit Ioab surgant
2SAM|2|15|surrexerunt ergo et transierunt numero duodecim de Beniamin ex parte Hisboseth filii Saul et duodecim de pueris David
2SAM|2|16|adprehensoque unusquisque capite conparis sui defixit gladium in latus contrarii et ceciderunt simul vocatumque est nomen loci illius ager Robustorum in Gabaon
2SAM|2|17|et ortum est bellum durum satis in die illa fugatusque est Abner et viri Israhel a pueris David
2SAM|2|18|erant autem ibi tres filii Sarviae Ioab et Abisai et Asahel porro Asahel cursor velocissimus fuit quasi unus ex capreis quae morantur in silvis
2SAM|2|19|persequebatur autem Asahel Abner et non declinavit ad dexteram sive ad sinistram omittens persequi Abner
2SAM|2|20|respexit itaque Abner post tergum suum et ait tune es Asahel qui respondit ego sum
2SAM|2|21|dixitque ei Abner vade ad dextram sive ad sinistram et adprehende unum de adulescentibus et tolle tibi spolia eius noluit autem Asahel omittere quin urgueret eum
2SAM|2|22|rursumque locutus est Abner ad Asahel recede noli me sequi ne conpellar confodere te in terra et levare non potero faciem meam ad Ioab fratrem tuum
2SAM|2|23|qui audire contempsit et noluit declinare percussit ergo eum Abner aversa hasta in inguine et transfodit et mortuus est in eodem loco omnesque qui transiebant per locum in quo ceciderat Asahel et mortuus erat subsistebant
2SAM|2|24|persequentibus autem Ioab et Abisai fugientem Abner sol occubuit et venerunt usque ad collem Aquaeductus qui est ex adverso vallis et itineris deserti in Gabaon
2SAM|2|25|congregatique sunt filii Beniamin ad Abner et conglobati in unum cuneum steterunt in summitate tumuli unius
2SAM|2|26|et exclamavit Abner ad Ioab et ait num usque ad internicionem tuus mucro desaeviet an ignoras quod periculosa sit desperatio usquequo non dicis populo ut omittat persequi fratres suos
2SAM|2|27|et ait Ioab vivit Dominus si locutus fuisses mane recessisset populus persequens fratrem suum
2SAM|2|28|insonuit ergo Ioab bucina et stetit omnis exercitus nec persecuti sunt ultra Israhel neque iniere certamen
2SAM|2|29|Abner autem et viri eius abierunt per campestria tota nocte illa et transierunt Iordanem et lustrata omni Bethoron venerunt ad Castra
2SAM|2|30|porro Ioab reversus omisso Abner congregavit omnem populum et defuerunt de pueris David decem et novem viri excepto Asahele
2SAM|2|31|servi autem David percusserunt de Beniamin et de viris qui erant cum Abner trecentos sexaginta qui et mortui sunt
2SAM|2|32|tuleruntque Asahel et sepelierunt eum in sepulchro patris sui in Bethleem et ambulaverunt tota nocte Ioab et viri qui erant cum eo et in ipso crepusculo pervenerunt in Hebron
2SAM|3|1|facta est ergo longa concertatio inter domum Saul et inter domum David David proficiens et semper se ipso robustior domus autem Saul decrescens cotidie
2SAM|3|2|nati quoque sunt filii David in Hebron fuitque primogenitus eius Amnon de Ahinoem Iezrahelitide
2SAM|3|3|et post eum Chelaab de Abigail uxore Nabal Carmeli porro tertius Absalom filius Maacha filiae Tholomai regis Gessur
2SAM|3|4|quartus autem Adonias filius Aggith et quintus Safathia filius Abital
2SAM|3|5|sextus quoque Iethraam de Agla uxore David hii nati sunt David in Hebron
2SAM|3|6|cum ergo esset proelium inter domum Saul et domum David Abner filius Ner regebat domum Saul
2SAM|3|7|fuerat autem Sauli concubina nomine Respha filia Ahia dixitque Hisboseth ad Abner
2SAM|3|8|quare ingressus es ad concubinam patris mei qui iratus nimis propter verba Hisboseth ait numquid caput canis ego sum adversum Iuda hodie qui fecerim misericordiam super domum Saul patris tui et super fratres et proximos eius et non tradidi te in manu David et tu requisisti in me quod argueres pro muliere hodie
2SAM|3|9|haec faciat Deus Abner et haec addat ei nisi quomodo iuravit Dominus David sic faciam cum eo
2SAM|3|10|ut transferatur regnum de domo Saul et elevetur thronus David super Israhel et super Iudam a Dan usque Bersabee
2SAM|3|11|et non potuit respondere ei quicquam quia metuebat illum
2SAM|3|12|misit ergo Abner nuntios ad David pro se dicentes cuius est terra et loquerentur fac mecum amicitias et erit manus mea tecum et reducam ad te universum Israhel
2SAM|3|13|qui ait optime ego faciam tecum amicitias sed unam rem peto a te dicens non videbis faciem meam antequam adduxeris Michol filiam Saul et sic venies et videbis me
2SAM|3|14|misit autem David nuntios ad Hisboseth filium Saul dicens redde uxorem meam Michol quam despondi mihi centum praeputiis Philisthim
2SAM|3|15|misit ergo Hisboseth et tulit eam a viro suo Faltihel filio Lais
2SAM|3|16|sequebaturque eam vir suus plorans usque Baurim et dixit ad eum Abner vade revertere qui reversus est
2SAM|3|17|sermonem quoque intulit Abner ad seniores Israhel dicens tam heri quam nudius tertius quaerebatis David ut regnaret super vos
2SAM|3|18|nunc ergo facite quoniam Dominus locutus est ad David dicens in manu servi mei David salvabo populum meum Israhel de manu Philisthim et omnium inimicorum eius
2SAM|3|19|locutus est autem Abner etiam ad Beniamin et abiit ut loqueretur ad David in Hebron omnia quae placuerant Israhel et universo Beniamin
2SAM|3|20|venitque ad David in Hebron cum viginti viris et fecit David Abner et viris eius qui venerant cum eo convivium
2SAM|3|21|et dixit Abner ad David surgam ut congregem ad te dominum meum regem omnem Israhel et ineam tecum foedus et imperes omnibus sicut desiderat anima tua cum ergo deduxisset David Abner et ille isset in pace
2SAM|3|22|statim pueri David et Ioab venerunt caesis latronibus cum praeda magna nimis Abner autem non erat cum David in Hebron quia iam dimiserat eum et profectus fuerat in pace
2SAM|3|23|et Ioab et omnis exercitus qui erat cum eo postea venerant nuntiatum est itaque Ioab a narrantibus venit Abner filius Ner ad regem et dimisit eum et abiit in pace
2SAM|3|24|et ingressus est Ioab ad regem et ait quid fecisti ecce venit Abner ad te quare dimisisti eum et abiit et recessit
2SAM|3|25|ignoras Abner filium Ner quoniam ad hoc venit ut deciperet te et sciret exitum tuum et introitum tuum et nosset omnia quae agis
2SAM|3|26|egressus itaque Ioab a David misit nuntios post Abner et reduxit eum a cisterna Sira ignorante David
2SAM|3|27|cumque redisset Abner in Hebron seorsum abduxit eum Ioab ad medium portae ut loqueretur ei in dolo et percussit illum ibi in inguine et mortuus est in ultionem sanguinis Asahel fratris eius
2SAM|3|28|quod cum audisset David rem iam gestam ait mundus ego sum et regnum meum apud Dominum usque in sempiternum a sanguine Abner filii Ner
2SAM|3|29|et veniat super caput Ioab et super omnem domum patris eius nec deficiat de domo Ioab fluxum seminis sustinens et leprosus tenens fusum et cadens gladio et indigens pane
2SAM|3|30|igitur Ioab et Abisai frater eius interfecerunt Abner eo quod occidisset Asahel fratrem eorum in Gabaon in proelio
2SAM|3|31|dixit autem David ad Ioab et ad omnem populum qui erat cum eo scindite vestimenta vestra et accingimini saccis et plangite ante exequias Abner porro rex David sequebatur feretrum
2SAM|3|32|cumque sepelissent Abner in Hebron levavit rex vocem suam et flevit super tumulum Abner flevit autem et omnis populus
2SAM|3|33|plangensque rex Abner ait nequaquam ut mori solent ignavi mortuus est Abner
2SAM|3|34|manus tuae non sunt ligatae et pedes tui non sunt conpedibus adgravati sed sicut solent cadere coram filiis iniquitatis corruisti congeminansque omnis populus flevit super eum
2SAM|3|35|cumque venisset universa multitudo cibum capere cum David clara adhuc die iuravit David dicens haec faciat mihi Deus et haec addat si ante occasum solis gustavero panem vel aliud quicquam
2SAM|3|36|omnisque populus audivit et placuerunt eis cuncta quae fecit rex in conspectu totius populi
2SAM|3|37|et cognovit omne vulgus et universus Israhel in die illa quoniam non actum fuisset a rege ut occideretur Abner filius Ner
2SAM|3|38|dixit quoque rex ad servos suos num ignoratis quoniam princeps et maximus cecidit hodie in Israhel
2SAM|3|39|ego autem adhuc delicatus et unctus rex porro viri isti filii Sarviae duri mihi sunt retribuat Dominus facienti malum iuxta malitiam suam
2SAM|4|1|audivit autem filius Saul quod cecidisset Abner in Hebron et dissolutae sunt manus eius omnisque Israhel perturbatus est
2SAM|4|2|duo autem viri principes latronum erant filio Saul nomen uni Baana et nomen alteri Rechab filii Remmon Berothitae de filiis Beniamin siquidem et Beroth reputata est in Beniamin
2SAM|4|3|et fugerunt Berothitae in Getthaim fueruntque ibi advenae usque in tempus illud
2SAM|4|4|erat autem Ionathan filio Saul filius debilis pedibus quinquennis enim fuit quando venit nuntius de Saul et Ionathan ex Iezrahel tollens itaque eum nutrix sua fugit cumque festinaret ut fugeret cecidit et claudus effectus est habuitque vocabulum Mifiboseth
2SAM|4|5|venientes igitur filii Remmon Berothitae Rechab et Baana ingressi sunt fervente die domum Hisboseth qui dormiebat super stratum suum meridie
2SAM|4|6|ingressi sunt autem domum adsumentes spicas tritici et percusserunt eum in inguine Rechab et Baana frater eius et fugerunt
2SAM|4|7|cum autem ingressi fuissent domum ille dormiebat super lectulum suum in conclavi et percutientes interfecerunt eum sublatoque capite eius abierunt per viam deserti tota nocte
2SAM|4|8|et adtulerunt caput Hisboseth ad David in Hebron dixeruntque ad regem ecce caput Hisboseth filii Saul inimici tui qui quaerebat animam tuam et dedit Dominus domino meo regi ultiones hodie de Saul et de semine eius
2SAM|4|9|respondens autem David Rechab et Baana fratri eius filiis Remmon Berothei dixit ad eos vivit Dominus qui eruit animam meam de omni angustia
2SAM|4|10|quoniam eum qui adnuntiaverat mihi et dixerat mortuus est Saul qui putabat se prospera nuntiare tenui et occidi in Siceleg cui oportebat me dare mercedem pro nuntio
2SAM|4|11|quanto magis nunc cum homines impii interfecerint virum innoxium in domo sua super lectulum suum non quaeram sanguinem eius de manu vestra et auferam vos de terra
2SAM|4|12|praecepit itaque David pueris et interfecerunt eos praecidentesque manus et pedes eorum suspenderunt eos super piscinam in Hebron caput autem Hisboseth tulerunt et sepelierunt in sepulchro Abner in Hebron
2SAM|5|1|et venerunt universae tribus Israhel ad David in Hebron dicentes ecce nos os tuum et caro tua sumus
2SAM|5|2|sed et heri et nudius tertius cum esset Saul rex super nos tu eras educens et reducens Israhel dixit autem Dominus ad te tu pasces populum meum Israhel et tu eris dux super Israhel
2SAM|5|3|venerunt quoque et senes de Israhel ad regem in Hebron et percussit cum eis rex David foedus in Hebron coram Domino unxeruntque David in regem super Israhel
2SAM|5|4|filius triginta annorum erat David cum regnare coepisset et quadraginta annis regnavit
2SAM|5|5|in Hebron regnavit super Iudam septem annis et sex mensibus in Hierusalem autem regnavit triginta tribus annis super omnem Israhel et Iudam
2SAM|5|6|et abiit rex et omnes viri qui erant cum eo in Hierusalem ad Iebuseum habitatorem terrae dictumque est ad David ab eis non ingredieris huc nisi abstuleris caecos et claudos dicentes non ingredietur David huc
2SAM|5|7|cepit autem David arcem Sion haec est civitas David
2SAM|5|8|proposuerat enim in die illa praemium qui percussisset Iebuseum et tetigisset domatum fistulas et claudos et caecos odientes animam David idcirco dicitur in proverbio caecus et claudus non intrabunt templum
2SAM|5|9|habitavit autem David in arce et vocavit eam civitatem David et aedificavit per gyrum a Mello et intrinsecus
2SAM|5|10|et ingrediebatur proficiens atque succrescens et Dominus Deus exercituum erat cum eo
2SAM|5|11|misit quoque Hiram rex Tyri nuntios ad David et ligna cedrina et artifices lignorum artificesque lapidum ad parietes et aedificaverunt domum David
2SAM|5|12|et cognovit David quoniam confirmasset eum Dominus regem super Israhel et quoniam exaltasset regnum eius super populum suum Israhel
2SAM|5|13|accepit ergo adhuc concubinas et uxores de Hierusalem postquam venerat de Hebron natique sunt David et alii filii et filiae
2SAM|5|14|et haec nomina eorum qui nati sunt ei in Hierusalem Samua et Sobab et Nathan et Salomon
2SAM|5|15|et Ibaar et Helisua et Nepheg
2SAM|5|16|et Iafia et Helisama et Helida et Helifeleth
2SAM|5|17|audierunt vero Philisthim quod unxissent David regem super Israhel et ascenderunt universi ut quaererent David quod cum audisset David descendit in praesidium
2SAM|5|18|Philisthim autem venientes diffusi sunt in valle Raphaim
2SAM|5|19|et consuluit David Dominum dicens si ascendam ad Philisthim et si dabis eos in manu mea et dixit Dominus ad David ascende quia tradens dabo Philisthim in manu tua
2SAM|5|20|venit ergo David in Baalpharasim et percussit eos ibi et dixit divisit Dominus inimicos meos coram me sicut dividuntur aquae propterea vocatum est nomen loci illius Baalpharasim
2SAM|5|21|et reliquerunt ibi sculptilia sua quae tulit David et viri eius
2SAM|5|22|et addiderunt adhuc Philisthim ut ascenderent et diffusi sunt in valle Raphaim
2SAM|5|23|consuluit autem David Dominum qui respondit non ascendas sed gyra post tergum eorum et venies ad eos ex adverso pirorum
2SAM|5|24|et cum audieris sonitum gradientis in cacumine pirorum tunc inibis proelium quia tunc egredietur Dominus ante faciem tuam ut percutiat castra Philisthim
2SAM|5|25|fecit itaque David sicut ei praeceperat Dominus et percussit Philisthim de Gabee usque dum venias Gezer
2SAM|6|1|congregavit autem rursum David omnes electos ex Israhel triginta milia
2SAM|6|2|surrexitque et abiit et universus populus qui erat cum eo de viris Iuda ut adducerent arcam Dei super quam invocatum est nomen Domini exercituum sedentis in cherubin super eam
2SAM|6|3|et inposuerunt arcam Domini super plaustrum novum tuleruntque eam de domo Abinadab qui erat in Gabaa Oza autem et Haio filii Abinadab minabant plaustrum novum
2SAM|6|4|cumque tulissent eam de domo Abinadab qui erat in Gabaa custodiens arcam Dei Haio praecedebat arcam
2SAM|6|5|David autem et omnis Israhel ludebant coram Domino in omnibus lignis fabrefactis et citharis et lyris et tympanis et sistris et cymbalis
2SAM|6|6|postquam autem venerunt ad aream Nachon extendit manum Oza ad arcam Dei et tenuit eam quoniam calcitrabant boves
2SAM|6|7|iratusque est indignatione Dominus contra Ozam et percussit eum super temeritate qui mortuus est ibi iuxta arcam Dei
2SAM|6|8|contristatus autem est David eo quod percussisset Dominus Ozam et vocatum est nomen loci illius Percussio Oza usque in diem hanc
2SAM|6|9|et extimuit David Dominum in die illa dicens quomodo ingredietur ad me arca Domini
2SAM|6|10|et noluit devertere ad se arcam Domini in civitate David sed devertit eam in domo Obededom Getthei
2SAM|6|11|et habitavit arca Domini in domo Obededom Getthei tribus mensibus et benedixit Dominus Obededom et omnem domum eius
2SAM|6|12|nuntiatumque est regi David benedixit Dominus Obededom et omnia eius propter arcam Dei abiit ergo David et adduxit arcam Dei de domo Obededom in civitatem David cum gaudio
2SAM|6|13|cumque transcendissent qui portabant arcam Domini sex passus immolabat bovem et arietem
2SAM|6|14|et David saltabat totis viribus ante Dominum porro David erat accinctus ephod lineo
2SAM|6|15|et David et omnis domus Israhel ducebant arcam testamenti Domini in iubilo et in clangore bucinae
2SAM|6|16|cumque intrasset arca Domini civitatem David Michol filia Saul prospiciens per fenestram vidit regem David subsilientem atque saltantem coram Domino et despexit eum in corde suo
2SAM|6|17|et introduxerunt arcam Domini et posuerunt eam in loco suo in medio tabernaculi quod tetenderat ei David et obtulit David holocausta coram Domino et pacifica
2SAM|6|18|cumque conplesset offerens holocaustum et pacifica benedixit populo in nomine Domini exercituum
2SAM|6|19|et partitus est multitudini universae Israhel tam viro quam mulieri singulis collyridam panis unam et assaturam bubulae carnis unam et similam frixam oleo et abiit omnis populus unusquisque in domum suam
2SAM|6|20|reversusque est et David ut benediceret domui suae et egressa Michol filia Saul in occursum David ait quam gloriosus fuit hodie rex Israhel discoperiens se ante ancillas servorum suorum et nudatus est quasi si nudetur unus de scurris
2SAM|6|21|dixitque David ad Michol ante Dominum qui elegit me potius quam patrem tuum et quam omnem domum eius et praecepit mihi ut essem dux super populum Domini Israhel
2SAM|6|22|et ludam et vilior fiam plus quam factus sum et ero humilis in oculis meis et cum ancillis de quibus locuta es gloriosior apparebo
2SAM|6|23|igitur Michol filiae Saul non est natus filius usque ad diem mortis suae
2SAM|7|1|factum est autem cum sedisset rex in domo sua et Dominus dedisset ei requiem undique ab universis inimicis suis
2SAM|7|2|dixit ad Nathan prophetam videsne quod ego habitem in domo cedrina et arca Dei posita sit in medio pellium
2SAM|7|3|dixitque Nathan ad regem omne quod est in corde tuo vade fac quia Dominus tecum est
2SAM|7|4|factum est autem in nocte illa et ecce sermo Domini ad Nathan dicens
2SAM|7|5|vade et loquere ad servum meum David haec dicit Dominus numquid tu aedificabis mihi domum ad habitandum
2SAM|7|6|neque enim habitavi in domo ex die qua eduxi filios Israhel de terra Aegypti usque in diem hanc sed ambulans ambulabam in tabernaculo et in tentorio
2SAM|7|7|per cuncta loca quae transivi cum omnibus filiis Israhel numquid loquens locutus sum ad unam de tribubus Israhel cui praecepi ut pasceret populum meum Israhel dicens quare non aedificastis mihi domum cedrinam
2SAM|7|8|et nunc haec dices servo meo David haec dicit Dominus exercituum ego tuli te de pascuis sequentem greges ut esses dux super populum meum Israhel
2SAM|7|9|et fui tecum in omnibus ubicumque ambulasti et interfeci universos inimicos tuos a facie tua fecique tibi nomen grande iuxta nomen magnorum qui sunt in terra
2SAM|7|10|et ponam locum populo meo Israhel et plantabo eum et habitabit sub eo et non turbabitur amplius nec addent filii iniquitatis ut adfligant eum sicut prius
2SAM|7|11|ex die qua constitui iudices super populum meum Israhel et requiem dabo tibi ab omnibus inimicis tuis praedicitque tibi Dominus quod domum faciat tibi Dominus
2SAM|7|12|cumque conpleti fuerint dies tui et dormieris cum patribus tuis suscitabo semen tuum post te quod egredietur de utero tuo et firmabo regnum eius
2SAM|7|13|ipse aedificabit domum nomini meo et stabiliam thronum regni eius usque in sempiternum
2SAM|7|14|ego ero ei in patrem et ipse erit mihi in filium qui si inique aliquid gesserit arguam eum in virga virorum et in plagis filiorum hominum
2SAM|7|15|misericordiam autem meam non auferam ab eo sicut abstuli a Saul quem amovi a facie tua
2SAM|7|16|et fidelis erit domus tua et regnum tuum usque in aeternum ante faciem tuam et thronus tuus erit firmus iugiter
2SAM|7|17|secundum omnia verba haec et iuxta universam visionem istam sic locutus est Nathan ad David
2SAM|7|18|ingressus est autem rex David et sedit coram Domino et dixit quis ego sum Domine Deus et quae domus mea quia adduxisti me hucusque
2SAM|7|19|sed et hoc parum visum est in conspectu tuo Domine Deus nisi loquereris etiam de domo servi tui in longinquum ista est enim lex Adam Domine Deus
2SAM|7|20|quid ergo addere poterit adhuc David ut loquatur ad te tu enim scis servum tuum Domine Deus
2SAM|7|21|propter verbum tuum et secundum cor tuum fecisti omnia magnalia haec ita ut notum faceres servo tuo
2SAM|7|22|idcirco magnificatus es Domine Deus quia non est similis tui neque est deus extra te in omnibus quae audivimus auribus nostris
2SAM|7|23|quae est autem ut populus tuus Israhel gens in terra propter quam ivit Deus ut redimeret eam sibi in populum et poneret sibi nomen faceretque eis magnalia et horribilia super terram a facie populi tui quem redemisti tibi ex Aegypto gentem et deum eius
2SAM|7|24|et firmasti tibi populum tuum Israhel in populum sempiternum et tu Domine factus es eis in Deum
2SAM|7|25|nunc ergo Domine Deus verbum quod locutus es super servum tuum et super domum eius suscita in sempiternum et fac sicut locutus es
2SAM|7|26|et magnificetur nomen tuum usque in sempiternum atque dicatur Dominus exercituum Deus super Israhel et domus servi tui David erit stabilita coram Domino
2SAM|7|27|quia tu Domine exercituum Deus Israhel revelasti aurem servi tui dicens domum aedificabo tibi propterea invenit servus tuus cor suum ut oraret te oratione hac
2SAM|7|28|nunc ergo Domine Deus tu es Deus et verba tua erunt vera locutus es enim ad servum tuum bona haec
2SAM|7|29|incipe igitur et benedic domui servi tui ut sit in sempiternum coram te quia tu Domine Deus locutus es et benedictione tua benedicetur domus servi tui in sempiternum
2SAM|8|1|factum est autem post haec percussit David Philisthim et humiliavit eos et tulit David frenum tributi de manu Philisthim
2SAM|8|2|et percussit Moab et mensus est eos funiculo coaequans terrae mensus est autem duos funiculos unum ad occidendum et unum ad vivificandum factusque est Moab David serviens sub tributo
2SAM|8|3|et percussit David Adadezer filium Roob regem Soba quando profectus est ut dominaretur super flumen Eufraten
2SAM|8|4|et captis David ex parte eius mille septingentis equitibus et viginti milibus peditum subnervavit omnes iugales curruum dereliquit autem ex eis centum currus
2SAM|8|5|venit quoque Syria Damasci ut praesidium ferret Adadezer regi Soba et percussit David de Syria viginti duo milia virorum
2SAM|8|6|et posuit David praesidium in Syria Damasci factaque est Syria David serviens sub tributo servavit Dominus David in omnibus ad quaecumque profectus est
2SAM|8|7|et tulit David arma aurea quae habebant servi Adadezer et detulit ea in Hierusalem
2SAM|8|8|et de Bete et de Beroth civitatibus Adadezer tulit rex David aes multum nimis
2SAM|8|9|audivit autem Thou rex Emath quod percussisset David omne robur Adadezer
2SAM|8|10|et misit Thou Ioram filium suum ad regem David ut salutaret eum congratulans et gratias ageret eo quod expugnasset Adadezer et percussisset eum hostis quippe erat Thou Adadezer et in manu eius erant vasa argentea et vasa aurea et vasa aerea
2SAM|8|11|quae et ipsa sanctificavit rex David Domino cum argento et auro quae sanctificaverat de universis gentibus quas subegerat
2SAM|8|12|de Syria et Moab et filiis Ammon et Philisthim et Amalech et de manubiis Adadezer filii Roob regis Soba
2SAM|8|13|fecit quoque sibi David nomen cum reverteretur capta Syria in valle Salinarum caesis duodecim milibus
2SAM|8|14|et posuit in Idumea custodes statuitque praesidium et facta est universa Idumea serviens David et servavit Dominus David in omnibus ad quaecumque profectus est
2SAM|8|15|et regnavit David super omnem Israhel faciebat quoque David iudicium et iustitiam omni populo suo
2SAM|8|16|Ioab autem filius Sarviae erat super exercitum porro Iosaphat filius Ahilud erat a commentariis
2SAM|8|17|et Sadoc filius Achitob et Ahimelech filius Abiathar sacerdotes et Saraias scriba
2SAM|8|18|Banaias autem filius Ioiada super Cherethi et Felethi filii autem David sacerdotes erant
2SAM|9|1|et dixit David putasne est aliquis qui remanserit de domo Saul ut faciam cum eo misericordiam propter Ionathan
2SAM|9|2|erat autem de domo Saul servus nomine Siba quem cum vocasset rex ad se dixit ei tune es Siba et ille respondit ego sum servus tuus
2SAM|9|3|et ait rex num superest aliquis de domo Saul ut faciam cum eo misericordiam Dei dixitque Siba regi superest filius Ionathan debilis pedibus
2SAM|9|4|ubi inquit est et Siba ad regem ecce ait in domo est Machir filii Amihel in Lodabar
2SAM|9|5|misit ergo rex David et tulit eum de domo Machir filii Amihel de Lodabar
2SAM|9|6|cum autem venisset Mifiboseth filius Ionathan filii Saul ad David corruit in faciem suam et adoravit dixitque David Mifiboseth qui respondit adsum servus tuus
2SAM|9|7|et ait ei David ne timeas quia faciens faciam in te misericordiam propter Ionathan patrem tuum et restituam tibi omnes agros Saul patris tui et tu comedes panem in mensa mea semper
2SAM|9|8|qui adorans eum dixit quis ego sum servus tuus quoniam respexisti super canem mortuum similem mei
2SAM|9|9|vocavit itaque rex Sibam puerum Saul et dixit ei omnia quaecumque fuerunt Saul et universam domum eius dedi filio domini tui
2SAM|9|10|operare igitur ei terram tu et filii tui et servi tui et inferes filio domini tui cibos ut alatur Mifiboseth autem filius domini tui comedet semper panem super mensam meam erant autem Sibae quindecim filii et viginti servi
2SAM|9|11|dixitque Siba ad regem sicut iussisti domine mi rex servo tuo sic faciet servus tuus et Mifiboseth comedet super mensam tuam quasi unus de filiis regis
2SAM|9|12|habebat autem Mifiboseth filium parvulum nomine Micha omnis vero cognatio domus Siba serviebat Mifiboseth
2SAM|9|13|porro Mifiboseth habitabat in Hierusalem quia de mensa regis iugiter vescebatur et erat claudus utroque pede
2SAM|10|1|factum est autem post haec ut moreretur rex filiorum Ammon et regnaret Anon filius eius pro eo
2SAM|10|2|dixitque David faciam misericordiam cum Anon filio Naas sicut fecit pater eius mecum misericordiam misit ergo David consolans eum per servos suos super patris interitu cum autem venissent servi David in terram filiorum Ammon
2SAM|10|3|dixerunt principes filiorum Ammon ad Anon dominum suum putas quod propter honorem patris tui David miserit ad te consolatores et non ideo ut investigaret et exploraret civitatem et everteret eam misit David servos suos ad te
2SAM|10|4|tulit itaque Anon servos David rasitque dimidiam partem barbae eorum et praecidit vestes eorum medias usque ad nates et dimisit eos
2SAM|10|5|quod cum nuntiatum esset David misit in occursum eorum erant enim viri confusi turpiter valde et mandavit eis David manete Hiericho donec crescat barba vestra et tunc revertimini
2SAM|10|6|videntes autem filii Ammon quod iniuriam fecissent David miserunt et conduxerunt mercede Syrum Roob et Syrum Soba viginti milia peditum et a rege Maacha mille viros et ab Histob duodecim milia virorum
2SAM|10|7|quod cum audisset David misit Ioab et omnem exercitum bellatorum
2SAM|10|8|egressi sunt ergo filii Ammon et direxerunt aciem ante ipsum introitum portae Syrus autem Soba et Roob et Histob et Maacha seorsum erant in campo
2SAM|10|9|videns igitur Ioab quod praeparatum esset adversum se proelium et ex adverso et post tergum elegit ex omnibus electis Israhel et instruxit aciem contra Syrum
2SAM|10|10|reliquam autem partem populi tradidit Abisai fratri suo qui direxit aciem adversum filios Ammon
2SAM|10|11|et ait Ioab si praevaluerint adversum me Syri eris mihi in adiutorium si autem filii Ammon praevaluerint adversum te auxiliabor tibi
2SAM|10|12|esto vir fortis et pugnemus pro populo nostro et civitate Dei nostri Dominus autem faciet quod bonum est in conspectu suo
2SAM|10|13|iniit itaque Ioab et populus qui erat cum eo certamen contra Syros qui statim fugerunt a facie eius
2SAM|10|14|filii autem Ammon videntes quod fugissent Syri fugerunt et ipsi a facie Abisai et ingressi sunt civitatem reversusque est Ioab a filiis Ammon et venit Hierusalem
2SAM|10|15|videntes igitur Syri quoniam corruissent coram Israhel congregati sunt pariter
2SAM|10|16|misitque Adadezer et eduxit Syros qui erant trans Fluvium et adduxit exercitum eorum Sobach autem magister militiae Adadezer erat princeps eorum
2SAM|10|17|quod cum nuntiatum esset David contraxit omnem Israhelem et transivit Iordanem venitque in Helema et direxerunt aciem Syri ex adverso David et pugnaverunt contra eum
2SAM|10|18|fugeruntque Syri a facie Israhel et occidit David de Syris septingentos currus et quadraginta milia equitum et Sobach principem militiae percussit qui statim mortuus est
2SAM|10|19|videntes autem universi reges qui erant in praesidio Adadezer victos se ab Israhel fecerunt pacem cum Israhel et servierunt eis timueruntque Syri auxilium praebere filiis Ammon
2SAM|11|1|factum est ergo vertente anno eo tempore quo solent reges ad bella procedere misit David Ioab et servos suos cum eo et universum Israhel et vastaverunt filios Ammon et obsederunt Rabba David autem remansit in Hierusalem
2SAM|11|2|dum haec agerentur accidit ut surgeret David de stratu suo post meridiem et deambularet in solario domus regiae viditque mulierem se lavantem ex adverso super solarium suum erat autem mulier pulchra valde
2SAM|11|3|misit ergo rex et requisivit quae esset mulier nuntiatumque ei est quod ipsa esset Bethsabee filia Heliam uxor Uriae Hetthei
2SAM|11|4|missis itaque David nuntiis tulit eam quae cum ingressa esset ad illum dormivit cum ea statimque sanctificata est ab inmunditia sua
2SAM|11|5|et reversa est domum suam concepto fetu mittensque nuntiavit David et ait concepi
2SAM|11|6|misit autem David ad Ioab dicens mitte ad me Uriam Hettheum misitque Ioab Uriam ad David
2SAM|11|7|et venit Urias ad David quaesivitque David quam recte ageret Ioab et populus et quomodo administraretur bellum
2SAM|11|8|et dixit David ad Uriam vade in domum tuam et lava pedes tuos egressus est Urias de domo regis secutusque est eum cibus regius
2SAM|11|9|dormivit autem Urias ante portam domus regiae cum aliis servis domini sui et non descendit ad domum suam
2SAM|11|10|nuntiatumque est David a dicentibus non ivit Urias ad domum suam et ait David ad Uriam numquid non de via venisti quare non descendisti ad domum tuam
2SAM|11|11|et ait Urias ad David arca et Israhel et Iuda habitant in papilionibus et dominus meus Ioab et servi domini mei super faciem terrae manent et ego ingrediar domum meam ut comedam et bibam et dormiam cum uxore mea per salutem tuam et per salutem animae tuae quod non faciam rem hanc
2SAM|11|12|ait ergo David ad Uriam mane hic etiam hodie et cras dimittam te mansit Urias in Hierusalem die illa et altera
2SAM|11|13|et vocavit eum David ut comederet coram se et biberet et inebriavit eum qui egressus vespere dormivit in stratu suo cum servis domini sui et in domum suam non descendit
2SAM|11|14|factum est ergo mane et scripsit David epistulam ad Ioab misitque per manum Uriae
2SAM|11|15|scribens in epistula ponite Uriam ex adverso belli ubi fortissimum proelium est et derelinquite eum ut percussus intereat
2SAM|11|16|igitur cum Ioab obsideret urbem posuit Uriam in loco quo sciebat viros esse fortissimos
2SAM|11|17|egressique viri de civitate bellabant adversum Ioab et ceciderunt de populo servorum David et mortuus est etiam Urias Hettheus
2SAM|11|18|misit itaque Ioab et nuntiavit David omnia verba proelii
2SAM|11|19|praecepitque nuntio dicens cum conpleveris universos sermones belli ad regem
2SAM|11|20|si eum videris indignari et dixerit quare accessistis ad murum ut proeliaremini an ignorabatis quod multa desuper ex muro tela mittantur
2SAM|11|21|quis percussit Abimelech filium Hieroboseth nonne mulier misit super eum fragmen molae de muro et interfecit eum in Thebes quare iuxta murum accessistis dices etiam servus tuus Urias Hettheus occubuit
2SAM|11|22|abiit ergo nuntius et venit et narravit David omnia quae ei praeceperat Ioab
2SAM|11|23|et dixit nuntius ad David praevaluerunt adversum nos viri et egressi sunt ad nos in agrum nos autem facto impetu persecuti eos sumus usque ad portam civitatis
2SAM|11|24|et direxerunt iacula sagittarii ad servos tuos ex muro desuper mortuique sunt de servis regis quin etiam servus tuus Urias Hettheus mortuus est
2SAM|11|25|et dixit David ad nuntium haec dices Ioab non te frangat ista res varius enim eventus est proelii et nunc hunc nunc illum consumit gladius conforta bellatores tuos adversum urbem ut destruas eam et exhortare eos
2SAM|11|26|audivit autem uxor Uriae quod mortuus esset Urias vir suus et planxit eum
2SAM|11|27|transactoque luctu misit David et introduxit eam domum suam et facta est ei uxor peperitque ei filium et displicuit verbum hoc quod fecerat David coram Domino
2SAM|12|1|misit ergo Dominus Nathan ad David qui cum venisset ad eum dixit ei duo viri erant in civitate una unus dives et alter pauper
2SAM|12|2|dives habebat oves et boves plurimos valde
2SAM|12|3|pauper autem nihil habebat omnino praeter ovem unam parvulam quam emerat et nutrierat et quae creverat apud eum cum filiis eius simul de pane illius comedens et de calice eius bibens et in sinu illius dormiens eratque illi sicut filia
2SAM|12|4|cum autem peregrinus quidam venisset ad divitem parcens ille sumere de ovibus et de bubus suis ut exhiberet convivium peregrino illi qui venerat ad se tulit ovem viri pauperis et praeparavit cibos homini qui venerat ad se
2SAM|12|5|iratus autem indignatione David adversus hominem illum nimis dixit ad Nathan vivit Dominus quoniam filius mortis est vir qui fecit hoc
2SAM|12|6|ovem reddet in quadruplum eo quod fecerit verbum istud et non pepercerit
2SAM|12|7|dixit autem Nathan ad David tu es ille vir haec dicit Dominus Deus Israhel ego unxi te in regem super Israhel et ego erui te de manu Saul
2SAM|12|8|et dedi tibi domum domini tui et uxores domini tui in sinu tuo dedique tibi domum Israhel et Iuda et si parva sunt ista adiciam tibi multo maiora
2SAM|12|9|quare ergo contempsisti verbum Domini ut faceres malum in conspectu meo Uriam Hettheum percussisti gladio et uxorem illius accepisti uxorem et interfecisti eum gladio filiorum Ammon
2SAM|12|10|quam ob rem non recedet gladius de domo tua usque in sempiternum eo quod despexeris me et tuleris uxorem Uriae Hetthei ut esset uxor tua
2SAM|12|11|itaque haec dicit Dominus ecce ego suscitabo super te malum de domo tua et tollam uxores tuas in oculis tuis et dabo proximo tuo et dormiet cum uxoribus tuis in oculis solis huius
2SAM|12|12|tu enim fecisti abscondite ego vero faciam verbum istud in conspectu omnis Israhel et in conspectu solis
2SAM|12|13|et dixit David ad Nathan peccavi Domino dixitque Nathan ad David Dominus quoque transtulit peccatum tuum non morieris
2SAM|12|14|verumtamen quoniam blasphemare fecisti inimicos Domini propter verbum hoc filius qui natus est tibi morte morietur
2SAM|12|15|et reversus est Nathan domum suam percussitque Dominus parvulum quem pepererat uxor Uriae David et desperatus est
2SAM|12|16|deprecatusque est David Dominum pro parvulo et ieiunavit David ieiunio et ingressus seorsum iacuit super terram
2SAM|12|17|venerunt autem seniores domus eius cogentes eum ut surgeret de terra qui noluit neque comedit cum eis cibum
2SAM|12|18|accidit autem die septima ut moreretur infans timueruntque servi David nuntiare ei quod mortuus esset parvulus dixerunt enim ecce cum parvulus adhuc viveret loquebamur ad eum et non audiebat vocem nostram quanto magis si dixerimus mortuus est puer se adfliget
2SAM|12|19|cum ergo vidisset David servos suos musitantes intellexit quod mortuus esset infantulus dixitque ad servos suos num mortuus est puer qui responderunt ei mortuus est
2SAM|12|20|surrexit igitur David de terra et lotus unctusque est cumque mutasset vestem ingressus est domum Domini et adoravit et venit in domum suam petivitque ut ponerent ei panem et comedit
2SAM|12|21|dixerunt autem ei servi sui quis est sermo quem fecisti propter infantem cum adhuc viveret ieiunasti et flebas mortuo autem puero surrexisti et comedisti panem
2SAM|12|22|qui ait propter infantem dum adhuc viveret ieiunavi et flevi dicebam enim quis scit si forte donet eum mihi Dominus et vivet infans
2SAM|12|23|nunc autem quia mortuus est quare ieiuno numquid potero revocare eum amplius ego vadam magis ad eum ille vero non revertetur ad me
2SAM|12|24|et consolatus est David Bethsabee uxorem suam ingressusque ad eam dormivit cum ea quae genuit filium et vocavit nomen eius Salomon et Dominus dilexit eum
2SAM|12|25|misitque in manu Nathan prophetae et vocavit nomen eius Amabilis Domino eo quod diligeret eum Dominus
2SAM|12|26|igitur pugnabat Ioab contra Rabbath filiorum Ammon et expugnabat urbem regiam
2SAM|12|27|misitque Ioab nuntios ad David dicens dimicavi adversum Rabbath et capienda est urbs Aquarum
2SAM|12|28|nunc igitur congrega reliquam partem populi et obside civitatem et cape eam ne cum a me vastata fuerit urbs nomini meo adscribatur victoria
2SAM|12|29|congregavit itaque David omnem populum et profectus est adversum Rabbath cumque dimicasset cepit eam
2SAM|12|30|et tulit diadema regis eorum de capite eius pondo auri talentum habens gemmas pretiosissimas et inpositum est super caput David sed et praedam civitatis asportavit multam valde
2SAM|12|31|populum quoque eius adducens serravit et circumegit super eos ferrata carpenta divisitque cultris et transduxit in typo laterum sic fecit universis civitatibus filiorum Ammon et reversus est David et omnis exercitus Hierusalem
2SAM|13|1|factum est autem post haec ut Absalom filii David sororem speciosissimam vocabulo Thamar adamaret Amnon filius David
2SAM|13|2|et deperiret eam valde ita ut aegrotaret propter amorem eius quia cum esset virgo difficile ei videbatur ut quippiam inhoneste ageret cum ea
2SAM|13|3|erat autem Amnonis amicus nomine Ionadab filius Semaa fratris David vir prudens valde
2SAM|13|4|qui dixit ad eum quare sic adtenuaris macie fili regis per singulos dies cur non indicas mihi dixitque ei Amnon Thamar sororem Absalom fratris mei amo
2SAM|13|5|cui respondit Ionadab cuba super lectulum tuum et languorem simula cumque venerit pater tuus ut visitet te dic ei veniat oro Thamar soror mea ut det mihi cibum et faciat pulmentum ut comedam de manu eius
2SAM|13|6|accubuit itaque Amnon et quasi aegrotare coepit cumque venisset rex ad visitandum eum ait Amnon ad regem veniat obsecro Thamar soror mea ut faciat in oculis meis duas sorbitiunculas et cibum capiam de manu eius
2SAM|13|7|misit ergo David ad Thamar domum dicens veni in domum Amnon fratris tui et fac ei pulmentum
2SAM|13|8|venitque Thamar in domum Amnon fratris sui ille autem iacebat quae tollens farinam commiscuit et liquefaciens in oculis eius coxit sorbitiunculas
2SAM|13|9|tollensque quod coxerat effudit et posuit coram eo et noluit comedere dixitque Amnon eicite universos a me cumque eiecissent omnes
2SAM|13|10|dixit Amnon ad Thamar infer cibum in conclave ut vescar de manu tua tulit ergo Thamar sorbitiunculas quas fecerat et intulit ad Amnon fratrem suum in conclave
2SAM|13|11|cumque obtulisset ei cibum adprehendit eam et ait veni cuba mecum soror mea
2SAM|13|12|quae respondit ei noli frater mi noli opprimere me neque enim hoc fas est in Israhel noli facere stultitiam hanc
2SAM|13|13|et ego enim ferre non potero obprobrium meum et tu eris quasi unus de insipientibus in Israhel quin potius loquere ad regem et non negabit me tibi
2SAM|13|14|noluit autem adquiescere precibus eius sed praevalens viribus oppressit eam et cubavit cum illa
2SAM|13|15|et exosam eam habuit Amnon magno odio nimis ita ut maius esset odium quo oderat eam amore quo ante dilexerat dixitque ei Amnon surge vade
2SAM|13|16|quae respondit ei maius est hoc malum quod nunc agis adversum me quam quod ante fecisti expellens me et noluit audire eam
2SAM|13|17|sed vocato puero qui ministrabat ei dixit eice hanc a me foras et claude ostium post eam
2SAM|13|18|quae induta erat talari tunica huiuscemodi enim filiae regis virgines vestibus utebantur eiecit itaque eam minister illius foras clausitque fores post eam
2SAM|13|19|quae aspergens cinerem capiti suo scissa talari tunica inpositisque manibus super caput suum ibat ingrediens et clamans
2SAM|13|20|dixit autem ei Absalom frater suus num Amnon frater tuus concubuit tecum sed nunc soror tace frater tuus est neque adfligas cor tuum pro re hac mansit itaque Thamar contabescens in domo Absalom fratris sui
2SAM|13|21|cum autem audisset rex David verba haec contristatus est valde
2SAM|13|22|porro non est locutus Absalom ad Amnon nec malum nec bonum oderat enim Absalom Amnon eo quod violasset Thamar sororem suam
2SAM|13|23|factum est autem post tempus biennii ut tonderentur oves Absalom in Baalasor quae est iuxta Ephraim et vocavit Absalom omnes filios regis
2SAM|13|24|venitque ad regem et ait ad eum ecce tondentur oves servi tui veniat oro rex cum servis suis ad servum suum
2SAM|13|25|dixitque rex ad Absalom noli fili mi noli rogare ut veniamus omnes et gravemus te cum autem cogeret eum et noluisset ire benedixit ei
2SAM|13|26|et ait Absalom si non vis venire veniat obsecro nobiscum saltem Amnon frater meus dixitque ad eum rex non est necesse ut vadat tecum
2SAM|13|27|coegit itaque eum Absalom et dimisit cum eo Amnon et universos filios regis
2SAM|13|28|praeceperat autem Absalom pueris suis dicens observate cum temulentus fuerit Amnon vino et dixero vobis percutite eum et interficite nolite timere ego enim sum qui praecepi vobis roboramini et estote viri fortes
2SAM|13|29|fecerunt ergo pueri Absalom adversum Amnon sicut praeceperat eis Absalom surgentesque omnes filii regis ascenderunt singuli mulas suas et fugerunt
2SAM|13|30|cumque adhuc pergerent in itinere fama praevenit ad David dicens percussit Absalom omnes filios regis et non remansit ex eis saltem unus
2SAM|13|31|surrexit itaque rex et scidit vestimenta sua et cecidit super terram et omnes servi ipsius qui adsistebant ei sciderunt vestimenta sua
2SAM|13|32|respondens autem Ionadab filius Samaa fratris David dixit ne aestimet dominus meus quod omnes pueri filii regis occisi sint Amnon solus mortuus est quoniam in ore Absalom erat positus ex die qua oppressit Thamar sororem eius
2SAM|13|33|nunc ergo ne ponat dominus meus rex super cor suum verbum istud dicens omnes filii regis occisi sunt quoniam Amnon solus mortuus est
2SAM|13|34|fugit autem Absalom et levavit puer speculator oculos suos et aspexit et ecce populus multus veniebat per iter devium ex latere montis
2SAM|13|35|dixit autem Ionadab ad regem ecce filii regis adsunt iuxta verbum servi tui sic factum est
2SAM|13|36|cumque cessasset loqui apparuerunt et filii regis et intrantes levaverunt vocem suam et fleverunt sed et rex et omnes servi eius fleverunt ploratu magno nimis
2SAM|13|37|porro Absalom fugiens abiit ad Tholomai filium Amiur regem Gessur luxit ergo David filium suum cunctis diebus
2SAM|13|38|Absalom autem cum fugisset et venisset in Gessur fuit ibi tribus annis
2SAM|13|39|cessavitque David rex persequi Absalom eo quod consolatus esset super Amnon interitu
2SAM|14|1|intellegens autem Ioab filius Sarviae quod cor regis versum esset ad Absalom
2SAM|14|2|misit Thecuam et tulit inde mulierem sapientem dixitque ad eam lugere te simula et induere veste lugubri et ne unguaris oleo ut sis quasi mulier plurimo iam tempore lugens mortuum
2SAM|14|3|et ingredieris ad regem et loqueris ad eum sermones huiuscemodi posuit autem Ioab verba in ore eius
2SAM|14|4|itaque cum ingressa fuisset mulier thecuites ad regem cecidit coram eo super terram et adoravit et dixit serva me rex
2SAM|14|5|et ait ad eam rex quid causae habes quae respondit heu mulier vidua ego sum mortuus est enim vir meus
2SAM|14|6|et ancillae tuae erant duo filii qui rixati sunt adversum se in agro nullusque erat qui eos prohibere posset et percussit alter alterum et interfecit eum
2SAM|14|7|et ecce consurgens universa cognatio adversum ancillam tuam dicit trade eum qui percussit fratrem suum ut occidamus eum pro anima fratris sui quem interfecit et deleamus heredem et quaerunt extinguere scintillam meam quae relicta est ut non supersit viro meo nomen et reliquiae super terram
2SAM|14|8|et ait rex ad mulierem vade in domum tuam et ego iubebo pro te
2SAM|14|9|dixitque mulier thecuites ad regem in me domine mi rex iniquitas et in domum patris mei rex autem et thronus eius sit innocens
2SAM|14|10|et ait rex qui contradixerit tibi adduc eum ad me et ultra non addet ut tangat te
2SAM|14|11|quae ait recordetur rex Domini Dei sui ut non multiplicentur proximi sanguinis ad ulciscendum et nequaquam interficient filium meum qui ait vivit Dominus quia non cadet de capillis filii tui super terram
2SAM|14|12|dixit ergo mulier loquatur ancilla tua ad dominum meum regem verbum et ait loquere
2SAM|14|13|dixitque mulier quare cogitasti istiusmodi rem contra populum Dei et locutus est rex verbum istud ut peccet et non reducat eiectum suum
2SAM|14|14|omnes morimur et quasi aquae delabimur in terram quae non revertuntur nec vult perire Deus animam sed retractat cogitans ne penitus pereat qui abiectus est
2SAM|14|15|nunc igitur veni ut loquar ad regem dominum meum verbum hoc praesente populo et dixit ancilla tua loquar ad regem si quo modo faciat rex verbum ancillae suae
2SAM|14|16|et audivit rex ut liberaret ancillam suam de manu omnium qui volebant delere me et filium meum simul de hereditate Dei
2SAM|14|17|dicat ergo ancilla tua ut fiat verbum domini mei regis quasi sacrificium sicut enim angelus Dei sic est dominus meus rex ut nec benedictione nec maledictione moveatur unde et Dominus Deus tuus est tecum
2SAM|14|18|et respondens rex dixit ad mulierem ne abscondas a me verbum quod te interrogo dixitque mulier loquere domine mi rex
2SAM|14|19|et ait rex numquid manus Ioab tecum est in omnibus istis respondit mulier et ait per salutem animae tuae domine mi rex nec ad dextram nec ad sinistram est ex omnibus his quae locutus est dominus meus rex servus enim tuus Ioab ipse praecepit mihi et ipse posuit in os ancillae tuae omnia verba haec
2SAM|14|20|ut verterem figuram sermonis huius servus tuus Ioab praecepit istud tu autem domine mi sapiens es sicut habet sapientiam angelus Dei ut intellegas omnia super terram
2SAM|14|21|et ait rex ad Ioab ecce placatus feci verbum tuum vade igitur et revoca puerum Absalom
2SAM|14|22|cadensque Ioab super faciem suam in terram adoravit et benedixit regi et dixit Ioab hodie intellexit servus tuus quia inveni gratiam in oculis tuis domine mi rex fecisti enim sermonem servi tui
2SAM|14|23|surrexit ergo Ioab et abiit in Gessur et adduxit Absalom in Hierusalem
2SAM|14|24|dixit autem rex revertatur in domum suam et faciem meam non videat reversus est itaque Absalom in domum suam et faciem regis non vidit
2SAM|14|25|porro sicut Absalom vir non erat pulcher in omni Israhel et decorus nimis a vestigio pedis usque ad verticem non erat in eo ulla macula
2SAM|14|26|et quando tondebatur capillum semel autem in anno tondebatur quia gravabat eum caesaries ponderabat capillos capitis sui ducentis siclis pondere publico
2SAM|14|27|nati sunt autem Absalom filii tres et filia una nomine Thamar eleganti forma
2SAM|14|28|mansitque Absalom Hierusalem duobus annis et faciem regis non vidit
2SAM|14|29|misit itaque ad Ioab ut mitteret eum ad regem qui noluit venire ad eum cumque secundo misisset et ille noluisset venire
2SAM|14|30|dixit servis suis scitis agrum Ioab iuxta agrum meum habentem messem hordei ite igitur et succendite eum igni succenderunt ergo servi Absalom segetem igni
2SAM|14|31|surrexitque Ioab et venit ad Absalom in domum eius et dixit quare succenderunt servi tui segetem meam igni
2SAM|14|32|et respondit Absalom ad Ioab misi ad te obsecrans ut venires ad me et mitterem te ad regem ut diceres ei quare veni de Gessur melius mihi erat ibi esse obsecro ergo ut videam faciem regis quod si memor est iniquitatis meae interficiat me
2SAM|14|33|ingressus Ioab ad regem nuntiavit ei vocatusque Absalom intravit ad regem et adoravit super faciem terrae coram eo osculatusque est rex Absalom
2SAM|15|1|igitur post haec fecit sibi Absalom currum et equites et quinquaginta viros qui praecederent eum
2SAM|15|2|et mane consurgens Absalom stabat iuxta introitum portae et omnem virum qui habebat negotium ut veniret ad regis iudicium vocabat Absalom ad se et dicebat de qua civitate es tu qui respondens aiebat ex una tribu Israhel ego sum servus tuus
2SAM|15|3|respondebatque ei Absalom videntur mihi sermones tui boni et iusti sed non est qui te audiat constitutus a rege dicebatque Absalom
2SAM|15|4|quis me constituat iudicem super terram ut ad me veniant omnes qui habent negotium et iuste iudicem
2SAM|15|5|sed et cum accederet ad eum homo ut salutaret illum extendebat manum suam et adprehendens osculabatur eum
2SAM|15|6|faciebatque hoc omni Israhel qui veniebat ad iudicium ut audiretur a rege et sollicitabat corda virorum Israhel
2SAM|15|7|post quattuor autem annos dixit Absalom ad regem vadam et reddam vota mea quae vovi Domino in Hebron
2SAM|15|8|vovens enim vovit servus tuus cum esset in Gessur Syriae dicens si reduxerit me Dominus in Hierusalem sacrificabo Domino
2SAM|15|9|dixitque ei rex vade in pace et surrexit et abiit in Hebron
2SAM|15|10|misit autem Absalom exploratores in universas tribus Israhel dicens statim ut audieritis clangorem bucinae dicite regnavit Absalom in Hebron
2SAM|15|11|porro cum Absalom ierunt ducenti viri de Hierusalem vocati euntes simplici corde et causam penitus ignorantes
2SAM|15|12|accersivit quoque Absalom Ahitofel Gilonitem consiliarium David de civitate sua Gilo cum immolaret victimas et facta est coniuratio valida populusque concurrens augebatur cum Absalom
2SAM|15|13|venit igitur nuntius ad David dicens toto corde universus Israhel sequitur Absalom
2SAM|15|14|et ait David servis suis qui erant cum eo in Hierusalem surgite fugiamus neque enim erit nobis effugium a facie Absalom festinate egredi ne forte veniens occupet nos et inpellat super nos ruinam et percutiat civitatem in ore gladii
2SAM|15|15|dixeruntque servi regis ad eum omnia quaecumque praeceperit dominus noster rex libenter exsequimur servi tui
2SAM|15|16|egressus est ergo rex et universa domus eius pedibus suis et dereliquit rex decem mulieres concubinas ad custodiendam domum
2SAM|15|17|egressusque rex et omnis Israhel pedibus suis stetit procul a domo
2SAM|15|18|et universi servi eius ambulabant iuxta eum et legiones Cherethi et Felethi et omnes Getthei sescenti viri qui secuti eum fuerant de Geth praecedebant regem
2SAM|15|19|dixit autem rex ad Ethai Gettheum cur venis nobiscum revertere et habita cum rege quia peregrinus es et egressus de loco tuo
2SAM|15|20|heri venisti et hodie inpelleris nobiscum egredi ego autem vadam quo iturus sum revertere et reduc tecum fratres tuos ostendisti gratiam et fidem
2SAM|15|21|et respondit Ethai regi dicens vivit Dominus et vivit dominus meus rex quoniam in quocumque loco fueris domine mi rex sive in morte sive in vita ibi erit servus tuus
2SAM|15|22|et ait David Ethai veni et transi et transivit Ethai Gettheus et omnes viri qui cum eo erant et reliqua multitudo
2SAM|15|23|omnesque flebant voce magna et universus populus transiebat rex quoque transgrediebatur torrentem Cedron et cunctus populus incedebat contra viam quae respicit ad desertum
2SAM|15|24|venit autem et Sadoc et universi Levitae cum eo portantes arcam foederis Dei et deposuerunt arcam Dei et ascendit Abiathar donec expletus est omnis populus qui egressus fuerat de civitate
2SAM|15|25|et dixit rex ad Sadoc reporta arcam Dei in urbem si invenero gratiam in oculis Domini reducet me et ostendet mihi eam et tabernaculum suum
2SAM|15|26|si autem dixerit non places praesto sum faciat quod bonum est coram se
2SAM|15|27|et dixit rex ad Sadoc sacerdotem o videns revertere in civitatem in pace et Achimaas filius tuus et Ionathan filius Abiathar duo filii vestri sint vobiscum
2SAM|15|28|ecce ego abscondar in campestribus deserti donec veniat sermo a vobis indicans mihi
2SAM|15|29|reportaverunt igitur Sadoc et Abiathar arcam Dei Hierusalem et manserunt ibi
2SAM|15|30|porro David ascendebat clivum Olivarum scandens et flens operto capite et nudis pedibus incedens sed et omnis populus qui erat cum eo operto capite ascendebat plorans
2SAM|15|31|nuntiatum est autem David quod et Ahitofel esset in coniuratione cum Absalom dixitque David infatua quaeso consilium Ahitofel Domine
2SAM|15|32|cumque ascenderet David summitatem montis in quo adoraturus erat Dominum ecce occurrit ei Husai Arachites scissa veste et terra pleno capite
2SAM|15|33|et dixit ei David si veneris mecum eris mihi oneri
2SAM|15|34|si autem in civitatem revertaris et dixeris Absalom servus tuus sum rex sicut fui servus patris tui sic ero servus tuus dissipabis consilium Ahitofel
2SAM|15|35|habes autem tecum Sadoc et Abiathar sacerdotes et omne verbum quodcumque audieris de domo regis indicabis Sadoc et Abiathar sacerdotibus
2SAM|15|36|sunt autem cum eis duo filii eorum Achimaas Sadoc et Ionathan Abiathar et mittetis per eos ad me omne verbum quod audieritis
2SAM|15|37|veniente ergo Husai amico David in civitatem Absalom quoque ingressus est Hierusalem
2SAM|16|1|cumque David transisset paululum montis verticem apparuit Siba puer Mifiboseth in occursum eius cum duobus asinis qui onerati erant ducentis panibus et centum alligaturis uvae passae et centum massis palatarum et utribus vini
2SAM|16|2|et dixit rex Sibae quid sibi volunt haec responditque Siba asini domestici regis ut sedeant et panes et palatae ad vescendum pueris tuis vinum autem ut bibat si quis defecerit in deserto
2SAM|16|3|et ait rex ubi est filius domini tui responditque Siba regi remansit in Hierusalem dicens hodie restituet mihi domus Israhel regnum patris mei
2SAM|16|4|et ait rex Sibae tua sint omnia quae fuerunt Mifiboseth dixitque Siba adoro inveniam gratiam coram te domine mi rex
2SAM|16|5|venit ergo rex David usque Baurim et ecce egrediebatur inde vir de cognatione domus Saul nomine Semei filius Gera procedebat egrediens et maledicebat
2SAM|16|6|mittebatque lapides contra David et contra universos servos regis David omnis autem populus et universi bellatores a dextro et sinistro latere regis incedebant
2SAM|16|7|ita autem loquebatur Semei cum malediceret regi egredere egredere vir sanguinum et vir Belial
2SAM|16|8|reddidit tibi Dominus universum sanguinem domus Saul quoniam invasisti regnum pro eo et dedit Dominus regnum in manu Absalom filii tui et ecce premunt te mala tua quoniam vir sanguinum es
2SAM|16|9|dixit autem Abisai filius Sarviae regi quare maledicit canis hic moriturus domino meo regi vadam et amputabo caput eius
2SAM|16|10|et ait rex quid mihi et vobis filii Sarviae dimittite eum maledicat Dominus enim praecepit ei ut malediceret David et quis est qui audeat dicere quare sic fecerit
2SAM|16|11|et ait rex Abisai et universis servis suis ecce filius meus qui egressus est de utero meo quaerit animam meam quanto magis nunc filius Iemini dimittite eum ut maledicat iuxta praeceptum Domini
2SAM|16|12|si forte respiciat Dominus adflictionem meam et reddat mihi bonum pro maledictione hac hodierna
2SAM|16|13|ambulabat itaque David et socii eius per viam cum eo Semei autem per iugum montis ex latere contra illum gradiebatur maledicens et mittens lapides adversum eum terramque spargens
2SAM|16|14|venit itaque rex et universus populus cum eo lassus et refocilati sunt ibi
2SAM|16|15|Absalom autem et omnis populus Israhel ingressi sunt Hierusalem sed et Ahitofel cum eo
2SAM|16|16|cum autem venisset Husai Arachites amicus David ad Absalom locutus est ad eum salve rex salve rex
2SAM|16|17|ad quem Absalom haec est inquit gratia tua ad amicum tuum quare non isti cum amico tuo
2SAM|16|18|responditque Husai ad Absalom nequaquam quia illius ero quem elegit Dominus et omnis hic populus et universus Israhel et cum eo manebo
2SAM|16|19|sed ut et hoc inferam cui ego serviturus sum nonne filio regis sicut parui patri tuo sic parebo et tibi
2SAM|16|20|dixit autem Absalom ad Ahitofel inite consilium quid agere debeamus
2SAM|16|21|et ait Ahitofel ad Absalom ingredere ad concubinas patris tui quas dimisit ad custodiendam domum ut cum audierit omnis Israhel quod foedaveris patrem tuum roborentur manus eorum tecum
2SAM|16|22|tetenderunt igitur Absalom tabernaculum in solario ingressusque est ad concubinas patris sui coram universo Israhel
2SAM|16|23|consilium autem Ahitofel quod dabat in diebus illis quasi si quis consuleret Deum sic erat omne consilium Ahitofel et cum esset cum David et cum esset cum Absalom
2SAM|17|1|dixit igitur Ahitofel ad Absalom eligam mihi duodecim milia virorum et consurgens persequar David hac nocte
2SAM|17|2|et inruens super eum quippe qui lassus est et solutis manibus percutiam eum cumque fugerit omnis populus qui cum eo est percutiam regem desolatum
2SAM|17|3|et reducam universum populum quomodo omnis reverti solet unum enim virum tu quaeris et omnis populus erit in pace
2SAM|17|4|placuitque sermo eius Absalom et cunctis maioribus natu Israhel
2SAM|17|5|ait autem Absalom vocate et Husai Arachiten et audiamus quid etiam ipse dicat
2SAM|17|6|cumque venisset Husai ad Absalom ait Absalom ad eum huiuscemodi sermonem locutus est Ahitofel facere debemus an non quod das consilium
2SAM|17|7|et dixit Husai ad Absalom non bonum consilium quod dedit Ahitofel hac vice
2SAM|17|8|et rursum intulit Husai tu nosti patrem tuum et viros qui cum eo sunt esse fortissimos et amaro animo veluti si ursa raptis catulis in saltu saeviat sed et pater tuus vir bellator est nec morabitur cum populo
2SAM|17|9|forsitan nunc latitat in foveis aut in uno quo voluerit loco et cum ceciderit unus quilibet in principio audiet quicumque audierit et dicet facta est plaga in populo qui sequebatur Absalom
2SAM|17|10|et fortissimus quoque cuius cor est quasi leonis pavore solvetur scit enim omnis populus Israhel fortem esse patrem tuum et robustos omnes qui cum eo sunt
2SAM|17|11|sed hoc mihi videtur rectum esse consilium congregetur ad te universus Israhel a Dan usque Bersabee quasi harena maris innumerabilis et tu eris in medio eorum
2SAM|17|12|et inruemus super eum in quocumque loco fuerit inventus et operiemus eum sicut cadere solet ros super terram et non relinquemus de viris qui cum eo sunt ne unum quidem
2SAM|17|13|quod si urbem aliquam fuerit ingressus circumdabit omnis Israhel civitati illi funes et trahemus eam in torrentem ut non repperiatur nec calculus quidem ex ea
2SAM|17|14|dixitque Absalom et omnis vir Israhel melius consilium Husai Arachitae consilio Ahitofel Domini autem nutu dissipatum est consilium Ahitofel utile ut induceret Dominus super Absalom malum
2SAM|17|15|et ait Husai Sadoc et Abiathar sacerdotibus hoc et hoc modo consilium dedit Ahitofel Absalom et senibus Israhel et ego tale et tale dedi consilium
2SAM|17|16|nunc ergo mittite cito et nuntiate David dicentes ne moremini nocte hac in campestribus deserti sed absque dilatione transgredere ne forte absorbeatur rex et omnis populus qui cum eo est
2SAM|17|17|Ionathan autem et Achimaas stabant iuxta fontem Rogel abiit ancilla et nuntiavit eis et illi profecti sunt ut referrent ad regem David nuntium non enim poterant videri aut introire civitatem
2SAM|17|18|vidit autem eos quidam puer et indicavit Absalom illi vero concito gradu ingressi sunt domum cuiusdam viri in Baurim qui habebat puteum in vestibulo suo et descenderunt in eum
2SAM|17|19|tulit autem mulier et expandit velamen super os putei quasi siccans ptisanas et sic res latuit
2SAM|17|20|cumque venissent servi Absalom ad mulierem in domum dixerunt ubi est Achimaas et Ionathan et respondit eis mulier transierunt gustata paululum aqua at hii qui quaerebant cum non repperissent reversi sunt Hierusalem
2SAM|17|21|cumque abissent ascenderunt illi de puteo et pergentes nuntiaverunt regi David atque dixerunt surgite transite cito fluvium quoniam huiuscemodi dedit consilium contra vos Ahitofel
2SAM|17|22|surrexit ergo David et omnis populus qui erat cum eo et transierunt Iordanem donec dilucesceret et ne unus quidem residuus fuit qui non transisset fluvium
2SAM|17|23|porro Ahitofel videns quod non fuisset factum consilium suum stravit asinum suum et surrexit et abiit in domum suam et in civitatem suam et disposita domo sua suspendio interiit et sepultus est in sepulchro patris sui
2SAM|17|24|David autem venit in Castra et Absalom transivit Iordanem ipse et omnis vir Israhel cum eo
2SAM|17|25|Amasam vero constituit Absalom pro Ioab super exercitum Amasa autem erat filius viri qui vocabatur Iethra de Hiesreli qui ingressus est ad Abigail filiam Naas sororem Sarviae quae fuit mater Ioab
2SAM|17|26|et castrametatus est Israhel cum Absalom in terra Galaad
2SAM|17|27|cumque venisset David in Castra Sobi filius Naas de Rabbath filiorum Ammon et Machir filius Ammihel de Lodabar et Berzellai Galaadites de Rogelim
2SAM|17|28|obtulerunt ei stratoria et tappetia et vasa fictilia frumentum et hordeum et farinam pulentam et fabam et lentem frixum cicer
2SAM|17|29|et mel et butyrum oves et pingues vitulos dederuntque David et populo qui cum eo erat ad vescendum suspicati enim sunt populum fame et siti fatigari in deserto
2SAM|18|1|igitur considerato David populo suo constituit super eum tribunos et centuriones
2SAM|18|2|et dedit populi tertiam partem sub manu Ioab et tertiam in manu Abisai filii Sarviae fratris Ioab et tertiam sub manu Ethai qui erat de Geth dixitque rex ad populum egrediar et ego vobiscum
2SAM|18|3|et respondit populus non exibis sive enim fugerimus non magnopere ad eos de nobis pertinebit sive media pars ceciderit e nobis non satis curabunt quia tu unus pro decem milibus conputaris melius est igitur ut sis nobis in urbe praesidio
2SAM|18|4|ad quos rex ait quod vobis rectum videtur hoc faciam stetit ergo rex iuxta portam egrediebaturque populus per turmas suas centeni et milleni
2SAM|18|5|et praecepit rex Ioab et Abisai et Ethai dicens servate mihi puerum Absalom et omnis populus audiebat praecipientem regem cunctis principibus pro Absalom
2SAM|18|6|itaque egressus est populus in campum contra Israhel et factum est proelium in saltu Ephraim
2SAM|18|7|et caesus est ibi populus Israhel ab exercitu David factaque est ibi plaga magna in die illa viginti milium
2SAM|18|8|fuit autem ibi proelium dispersum super faciem omnis terrae et multo plures erant quos saltus consumpserat de populo quam hii quos voraverat gladius in die illa
2SAM|18|9|accidit autem ut occurreret Absalom servis David sedens mulo cumque ingressus fuisset mulus subter condensam quercum et magnam adhesit caput eius quercui et illo suspenso inter caelum et terram mulus cui sederat pertransivit
2SAM|18|10|vidit autem hoc quispiam et nuntiavit Ioab dicens vidi Absalom pendere de quercu
2SAM|18|11|et ait Ioab viro qui nuntiaverat ei si vidisti quare non confodisti eum cum terra et ego dedissem tibi decem argenti siclos et unum balteum
2SAM|18|12|qui dixit ad Ioab si adpenderes in manibus meis mille argenteos nequaquam mitterem manum meam in filium regis audientibus enim nobis praecepit rex tibi et Abisai et Ethai dicens custodite mihi puerum Absalom
2SAM|18|13|sed et si fecissem contra animam meam audacter nequaquam hoc regem latere potuisset et tu stares ex adverso
2SAM|18|14|et ait Ioab non sicut tu vis sed adgrediar eum coram te tulit ergo tres lanceas in manu sua et infixit eas in corde Absalom cumque adhuc palpitaret herens in quercu
2SAM|18|15|cucurrerunt decem iuvenes armigeri Ioab et percutientes interfecerunt eum
2SAM|18|16|cecinit autem Ioab bucina et retinuit populum ne persequeretur fugientem Israhel volens parcere multitudini
2SAM|18|17|et tulerunt Absalom et proiecerunt eum in saltu in foveam grandem et conportaverunt super eum acervum lapidum magnum nimis omnis autem Israhel fugit in tabernacula sua
2SAM|18|18|porro Absalom erexerat sibi cum adhuc viveret titulum qui est in valle Regis dixerat enim non habeo filium et hoc erit monumentum nominis mei vocavitque titulum nomine suo et appellatur manus Absalom usque ad hanc diem
2SAM|18|19|Achimaas autem filius Sadoc ait curram et nuntiabo regi quia iudicium fecerit ei Dominus de manu inimicorum eius
2SAM|18|20|ad quem Ioab dixit non eris nuntius in hac die sed nuntiabis in alia hodie nolo te nuntiare filius enim regis est mortuus
2SAM|18|21|et ait Ioab Chusi vade et nuntia regi quae vidisti adoravit Chusi Ioab et cucurrit
2SAM|18|22|rursum autem Achimaas filius Sadoc dixit ad Ioab quid inpedit si etiam ego curram post Chusi dixitque Ioab quid vis currere fili mi non eris boni nuntii baiulus
2SAM|18|23|qui respondit quid enim si cucurrero et ait ei curre currens ergo Achimaas per viam conpendii transivit Chusi
2SAM|18|24|David autem sedebat inter duas portas speculator vero qui erat in fastigio portae super murum elevans oculos vidit hominem currentem solum
2SAM|18|25|et exclamans indicavit regi dixitque rex si solus est bonus est nuntius in ore eius properante autem illo et accedente propius
2SAM|18|26|vidit speculator hominem alterum currentem et vociferans in culmine ait apparet mihi homo currens solus dixitque rex et iste bonus est nuntius
2SAM|18|27|speculator autem contemplor ait cursum prioris quasi cursum Achimaas filii Sadoc et ait rex vir bonus est et nuntium portans bonum venit
2SAM|18|28|clamans autem Achimaas dixit ad regem salve et adorans regem coram eo pronus in terram ait benedictus Dominus Deus tuus qui conclusit homines qui levaverunt manus suas contra dominum meum regem
2SAM|18|29|et ait rex estne pax puero Absalom dixitque Achimaas vidi tumultum magnum cum mitteret Ioab servus tuus o rex me servum tuum nescio aliud
2SAM|18|30|ad quem rex transi ait et sta hic cumque ille transisset et staret
2SAM|18|31|apparuit Chusi et veniens ait bonum adporto nuntium domine mi rex iudicavit enim pro te Dominus hodie de manu omnium qui surrexerunt contra te
2SAM|18|32|dixit autem rex ad Chusi estne pax puero Absalom cui respondens Chusi fiant inquit sicut puer inimici domini mei regis et universi qui consurgunt adversum eum in malum
2SAM|18|33|contristatus itaque rex ascendit cenaculum portae et flevit et sic loquebatur vadens fili mi Absalom fili mi Absalom quis mihi tribuat ut ego moriar pro te Absalom fili mi fili mi
2SAM|19|1|nuntiatum est autem Ioab quod rex fleret et lugeret filium suum
2SAM|19|2|et versa est victoria in die illa in luctum omni populo audivit enim populus in die illa dici dolet rex super filio suo
2SAM|19|3|et declinabat populus in die illa ingredi civitatem quomodo declinare solet populus versus et fugiens de proelio
2SAM|19|4|porro rex operuit caput suum et clamabat voce magna fili mi Absalom Absalom fili mi fili mi
2SAM|19|5|ingressus ergo Ioab ad regem in domo dixit confudisti hodie vultus omnium servorum tuorum qui salvam fecerunt animam tuam et animam filiorum tuorum et filiarum tuarum et animam uxorum tuarum et animam concubinarum tuarum
2SAM|19|6|diligis odientes te et odio habes diligentes te et ostendisti hodie quia non curas de ducibus tuis et de servis tuis et vere cognovi modo quia si Absalom viveret et nos omnes occubuissemus tunc placeret tibi
2SAM|19|7|nunc igitur surge et procede et adloquens satisfac servis tuis iuro enim tibi per Dominum quod si non exieris ne unus quidem remansurus sit tecum nocte hac et peius erit hoc tibi quam omnia mala quae venerunt super te ab adulescentia tua usque in praesens
2SAM|19|8|surrexit ergo rex et sedit in porta et omni populo nuntiatum est quod rex sederet in porta venitque universa multitudo coram rege Israhel autem fugit in tabernacula sua
2SAM|19|9|omnis quoque populus certabat in cunctis tribubus Israhel dicens rex liberavit nos de manu inimicorum nostrorum ipse salvavit nos de manu Philisthinorum et nunc fugit de terra propter Absalom
2SAM|19|10|Absalom autem quem unximus super nos mortuus est in bello usquequo siletis et non reducitis regem
2SAM|19|11|rex vero David misit ad Sadoc et ad Abiathar sacerdotes dicens loquimini ad maiores natu Iuda dicentes cur venitis novissimi ad reducendum regem in domum suam sermo autem omnis Israhel pervenerat ad regem in domo eius
2SAM|19|12|fratres mei vos os meum et caro mea vos quare novissimi reducitis regem
2SAM|19|13|et Amasae dicite nonne os meum es et caro mea haec faciat mihi Deus et haec addat si non magister militiae fueris coram me omni tempore pro Ioab
2SAM|19|14|et inclinavit cor omnium virorum Iuda quasi viri unius miseruntque ad regem dicentes revertere tu et omnes servi tui
2SAM|19|15|et reversus est rex et venit usque ad Iordanem et Iuda venit in Galgala ut occurreret regi et transduceret eum Iordanem
2SAM|19|16|festinavit autem Semei filius Gera filii Iemini de Baurim et descendit cum viris Iuda in occursum regis David
2SAM|19|17|cum mille viris de Beniamin et Siba puer de domo Saul et quindecim filii eius ac viginti servi erant cum eo et inrumpentes Iordanem ante regem
2SAM|19|18|transierunt vada ut transducerent domum regis et facerent iuxta iussionem eius Semei autem filius Gera prostratus coram rege cum iam transisset Iordanem
2SAM|19|19|dixit ad eum ne reputes mihi domine mi iniquitatem neque memineris iniuriam servi tui in die qua egressus es domine mi rex de Hierusalem neque ponas rex in corde tuo
2SAM|19|20|agnosco enim servus tuus peccatum meum et idcirco hodie primus veni de omni domo Ioseph descendique in occursum domini mei regis
2SAM|19|21|respondens vero Abisai filius Sarviae dixit numquid pro his verbis non occidetur Semei quia maledixit christo Domini
2SAM|19|22|et ait David quid mihi et vobis filii Sarviae cur efficimini mihi hodie in Satan ergone hodie interficietur vir in Israhel an ignoro hodie me factum regem super Israhel
2SAM|19|23|et ait rex Semei non morieris iuravitque ei
2SAM|19|24|Mifiboseth quoque filius Saul descendit in occursum regis inlotis pedibus et intonsa barba vestesque suas non laverat a die qua egressus fuerat rex usque ad diem reversionis eius in pace
2SAM|19|25|cumque Hierusalem occurrisset regi dixit ei rex quare non venisti mecum Mifiboseth
2SAM|19|26|qui respondens ait domine mi rex servus meus contempsit me dixi ei ego famulus tuus ut sterneret mihi asinum et ascendens abirem cum rege claudus enim sum servus tuus
2SAM|19|27|insuper et accusavit me servum tuum ad te dominum meum regem tu autem domine mi rex sicut angelus Dei fac quod placitum est tibi
2SAM|19|28|neque enim fuit domus patris mei nisi morti obnoxia domino meo regi tu autem posuisti me servum tuum inter convivas mensae tuae quid igitur habeo iustae querellae aut quid possum ultra vociferari ad regem
2SAM|19|29|ait ergo ei rex quid ultra loqueris fixum est quod locutus sum tu et Siba dividite possessiones
2SAM|19|30|responditque Mifiboseth regi etiam cuncta accipiat postquam reversus est dominus meus rex pacifice in domum suam
2SAM|19|31|Berzellai quoque Galaadites descendens de Rogelim transduxit regem Iordanem paratus etiam ultra fluvium prosequi eum
2SAM|19|32|erat autem Berzellai Galaadites senex valde id est octogenarius et ipse praebuit alimenta regi cum moraretur in Castris fuit quippe vir dives nimis
2SAM|19|33|dixit itaque rex ad Berzellai veni mecum ut requiescas secure mecum in Hierusalem
2SAM|19|34|et ait Berzellai ad regem quot sunt dies annorum vitae meae ut ascendam cum rege Hierusalem
2SAM|19|35|octogenarius sum hodie numquid vigent sensus mei ad discernendum suave aut amarum aut delectare potest servum tuum cibus et potus vel audire ultra possum vocem cantorum atque cantricum quare servus tuus fit oneri domino meo regi
2SAM|19|36|paululum procedam famulus tuus ab Iordane tecum nec indigeo hac vicissitudine
2SAM|19|37|sed obsecro ut revertar servus tuus et moriar in civitate mea iuxta sepulchrum patris mei et matris meae est autem servus tuus Chamaam ipse vadat tecum domine mi rex et fac ei quod tibi bonum videtur
2SAM|19|38|dixitque rex mecum transeat Chamaam et ego faciam ei quicquid tibi placuerit et omne quod petieris a me inpetrabis
2SAM|19|39|cumque transisset universus populus et rex Iordanem osculatus est rex Berzellai et benedixit ei et ille reversus est in locum suum
2SAM|19|40|transivit ergo rex in Galgalam et Chamaam cum eo omnis autem populus Iuda transduxerat regem et media tantum pars adfuerat de populo Israhel
2SAM|19|41|itaque omnes viri Israhel concurrentes ad regem dixerunt ei quare te furati sunt fratres nostri viri Iuda et transduxerunt regem et domum eius Iordanem omnesque viros David cum eo
2SAM|19|42|et respondit omnis vir Iuda ad viros Israhel quia propior mihi est rex cur irasceris super hac re numquid comedimus aliquid ex rege aut munera nobis data sunt
2SAM|19|43|et respondit vir Israhel ad viros Iuda et ait decem partibus maior ego sum apud regem magisque ad me pertinet David quam ad te cur mihi fecisti iniuriam et non mihi nuntiatum est priori ut reducerem regem meum durius autem responderunt viri Iuda viris Israhel
2SAM|20|1|accidit quoque ut ibi esset vir Belial nomine Seba filius Bochri vir iemineus et cecinit bucina et ait non est nobis pars in David neque hereditas in filio Isai vir in tabernacula tua Israhel
2SAM|20|2|et separatus est omnis Israhel a David secutusque est Seba filium Bochri viri autem Iuda adheserunt regi suo a Iordane usque Hierusalem
2SAM|20|3|cumque venisset rex in domum suam Hierusalem tulit decem mulieres concubinas quas dereliquerat ad custodiendam domum et tradidit eas in custodiam alimenta eis praebens et non est ingressus ad eas sed erant clausae usque ad diem mortis suae in viduitate viventes
2SAM|20|4|dixit autem rex Amasae convoca mihi omnes viros Iuda in diem tertium et tu adesto praesens
2SAM|20|5|abiit ergo Amasa ut convocaret Iudam et moratus est extra placitum quod ei constituerat
2SAM|20|6|ait autem David ad Abisai nunc magis adflicturus est nos Seba filius Bochri quam Absalom tolle igitur servos domini tui et persequere eum ne forte inveniat civitates munitas et effugiat nos
2SAM|20|7|egressi sunt ergo cum eo viri Ioab Cherethi quoque et Felethi et omnes robusti exierunt de Hierusalem ad persequendum Seba filium Bochri
2SAM|20|8|cumque illi essent iuxta lapidem grandem qui est in Gabaon Amasa veniens occurrit eis porro Ioab vestitus erat tunica stricta ad mensuram habitus sui et desuper accinctus gladio dependente usque ad ilia in vagina qui fabrefactus levi motu egredi poterat et percutere
2SAM|20|9|dixit itaque Ioab ad Amasa salve mi frater et tenuit manu dextra mentum Amasae quasi osculans eum
2SAM|20|10|porro Amasa non observavit gladium quem habebat Ioab qui percussit eum in latere et effudit intestina eius in terram nec secundum vulnus adposuit Ioab autem et Abisai frater eius persecuti sunt Seba filium Bochri
2SAM|20|11|interea quidam viri cum stetissent iuxta cadaver Amasae de sociis Ioab dixerunt ecce qui esse voluit pro Ioab comes David pro Ioab
2SAM|20|12|Amasa autem conspersus sanguine iacebat in media via vidit hoc quidam vir quod subsisteret omnis populus ad videndum eum et amovit Amasam de via in agrum operuitque eum vestimento ne subsisterent transeuntes propter eum
2SAM|20|13|amoto igitur illo de via transiebat omnis vir sequens Ioab ad persequendum Seba filium Bochri
2SAM|20|14|porro ille transierat per omnes tribus Israhel in Abelam et in Bethmacha omnesque electi congregati fuerant ad eum
2SAM|20|15|venerunt itaque et obpugnabant eum in Abela et in Bethmacha et circumdederunt munitionibus civitatem et obsessa est urbs omnis autem turba quae erat cum Ioab moliebatur destruere muros
2SAM|20|16|et exclamavit mulier sapiens de civitate audite audite dicite Ioab adpropinqua huc et loquar tecum
2SAM|20|17|qui cum accessisset ad eam ait illi tu es Ioab et ille respondit ego ad quem sic locuta est audi sermones ancillae tuae qui respondit audio
2SAM|20|18|rursumque illa sermo inquit dicebatur in veteri proverbio qui interrogant interrogent in Abela et sic perficiebant
2SAM|20|19|nonne ego sum quae respondeo veritatem Israhel et tu quaeris subruere civitatem et evertere matrem in Israhel quare praecipitas hereditatem Domini
2SAM|20|20|respondensque Ioab ait absit absit hoc a me non praecipito neque demolior
2SAM|20|21|non se sic habet res sed homo de monte Ephraim Seba filius Bochri cognomine levavit manum contra regem David tradite illum solum et recedemus a civitate et ait mulier ad Ioab ecce caput eius mittetur ad te per murum
2SAM|20|22|ingressa est ergo ad omnem populum et locuta est eis sapienter qui abscisum caput Seba filii Bochri proiecerunt ad Ioab et ille cecinit tuba et recesserunt ab urbe unusquisque in tabernacula sua Ioab autem reversus est Hierusalem ad regem
2SAM|20|23|fuit ergo Ioab super omnem exercitum Israhel Banaias autem filius Ioiadae super Cheretheos et Feletheos
2SAM|20|24|Aduram vero super tributa porro Iosaphat filius Ahilud a commentariis
2SAM|20|25|Sia autem scriba Sadoc vero et Abiathar sacerdotes
2SAM|20|26|Hira autem Hiaiarites erat sacerdos David
2SAM|21|1|facta est quoque fames in diebus David tribus annis iugiter et consuluit David oraculum Domini dixitque Dominus propter Saul et domum eius et sanguinem quia occidit Gabaonitas
2SAM|21|2|vocatis ergo Gabaonitis rex dixit ad eos porro Gabaonitae non sunt de filiis Israhel sed reliquiae Amorreorum filii quippe Israhel iuraverant eis et voluit Saul percutere eos zelo quasi pro filiis Israhel et Iuda
2SAM|21|3|dixit ergo David ad Gabaonitas quid faciam vobis et quod erit vestri piaculum ut benedicatis hereditati Domini
2SAM|21|4|dixeruntque ei Gabaonitae non est nobis super argento et auro quaestio contra Saul et contra domum eius neque volumus ut interficiatur homo de Israhel ad quos ait quid ergo vultis ut faciam vobis
2SAM|21|5|qui dixerunt regi virum qui adtrivit nos et oppressit inique ita delere debemus ut ne unus quidem residuus sit de stirpe eius in cunctis finibus Israhel
2SAM|21|6|dentur nobis septem viri de filiis eius et crucifigamus eos Domino in Gabaath Saul quondam electi Domini et ait rex ego dabo
2SAM|21|7|pepercitque rex Mifiboseth filio Ionathan filii Saul propter iusiurandum Domini quod fuerat inter David et inter Ionathan filium Saul
2SAM|21|8|tulit itaque rex duos filios Respha filiae Ahia quos peperit Saul Armoni et Mifiboseth et quinque filios Michol filiae Saul quos genuerat Hadriheli filio Berzellai qui fuit de Molathi
2SAM|21|9|et dedit eos in manu Gabaonitarum qui crucifixerunt illos in monte coram Domino et ceciderunt hii septem simul occisi in diebus messis primis incipiente messione hordei
2SAM|21|10|tollens autem Respha filia Ahia cilicium substravit sibi super petram ab initio messis donec stillaret aqua super eos de caelo et non dimisit aves lacerare eos per diem neque bestias per noctem
2SAM|21|11|et nuntiata sunt David quae fecerat Respha filia Ahia concubina Saul
2SAM|21|12|et abiit David et tulit ossa Saul et ossa Ionathan filii eius a viris Iabesgalaad qui furati fuerant ea de platea Bethsan in qua suspenderant eos Philisthim cum interfecissent Saul in Gelboe
2SAM|21|13|et asportavit inde ossa Saul et ossa Ionathan filii eius et colligentes ossa eorum qui adfixi fuerant
2SAM|21|14|sepelierunt ea cum ossibus Saul et Ionathan filii eius in terra Beniamin in latere in sepulchro Cis patris eius feceruntque omnia quae praeceperat rex et repropitiatus est Deus terrae post haec
2SAM|21|15|factum est autem rursum proelium Philisthinorum adversum Israhel et descendit David et servi eius cum eo et pugnabant contra Philisthim deficiente autem David
2SAM|21|16|Iesbidenob qui fuit de genere Arafa cuius ferrum hastae trecentas uncias adpendebat et accinctus erat ense novo nisus est percutere David
2SAM|21|17|praesidioque ei fuit Abisai filius Sarviae et percussum Philistheum interfecit tunc iuraverunt viri David dicentes non egredieris nobiscum in bellum ne extinguas lucernam Israhel
2SAM|21|18|secundum quoque fuit bellum in Gob contra Philistheos tunc percussit Sobbochai de Usathi Seph de stirpe Arafa
2SAM|21|19|tertium quoque fuit bellum in Gob contra Philistheos in quo percussit Adeodatus filius Saltus polymitarius bethleemites Goliath Gettheum cuius hastile hastae erat quasi liciatorium texentium
2SAM|21|20|quartum bellum fuit in Geth in quo vir excelsus qui senos in manibus pedibusque habebat digitos id est viginti et quattuor et erat de origine Arafa
2SAM|21|21|blasphemavit Israhel percussit autem eum Ionathan filius Sammaa fratris David
2SAM|21|22|hii quattuor nati sunt de Arafa in Geth et ceciderunt in manu David et servorum eius
2SAM|22|1|locutus est autem David Domino verba carminis huius in die qua liberavit eum Dominus de manu omnium inimicorum suorum et de manu Saul
2SAM|22|2|et ait Dominus petra mea et robur meum et salvator meus
2SAM|22|3|Deus meus fortis meus sperabo in eum scutum meum et cornu salutis meae elevator meus et refugium meum salvator meus de iniquitate liberabis me
2SAM|22|4|laudabilem invocabo Dominum et ab inimicis meis salvus ero
2SAM|22|5|quia circumdederunt me contritiones mortis torrentes Belial terruerunt me
2SAM|22|6|funes inferi circumdederunt me praevenerunt me laquei mortis
2SAM|22|7|in tribulatione mea invocabo Dominum et ad Deum meum clamabo et exaudiet de templo suo vocem meam et clamor meus veniet ad aures eius
2SAM|22|8|commota est et contremuit terra fundamenta montium concussa sunt et conquassata quoniam iratus est
2SAM|22|9|ascendit fumus de naribus eius et ignis de ore eius voravit carbones incensi sunt ab eo
2SAM|22|10|et inclinavit caelos et descendit et caligo sub pedibus eius
2SAM|22|11|et ascendit super cherubin et volavit et lapsus est super pinnas venti
2SAM|22|12|posuit tenebras in circuitu suo latibulum cribrans aquas de nubibus caelorum
2SAM|22|13|prae fulgore in conspectu eius succensi sunt carbones ignis
2SAM|22|14|tonabit de caelis Dominus et Excelsus dabit vocem suam
2SAM|22|15|misit sagittas et dissipavit eos fulgur et consumpsit eos
2SAM|22|16|et apparuerunt effusiones maris et revelata sunt fundamenta orbis ab increpatione Domini ab inspiratione spiritus furoris eius
2SAM|22|17|misit de excelso et adsumpsit me extraxit me de aquis multis
2SAM|22|18|liberavit me ab inimico meo potentissimo ab his qui oderant me quoniam robustiores me erant
2SAM|22|19|praevenit me in die adflictionis meae et factus est Dominus firmamentum meum
2SAM|22|20|et eduxit me in latitudinem liberavit me quia placuit ei
2SAM|22|21|retribuet mihi Dominus secundum iustitiam meam et secundum munditiam manuum mearum reddet mihi
2SAM|22|22|quia custodivi vias Domini et non egi impie a Deo meo
2SAM|22|23|omnia enim iudicia eius in conspectu meo et praecepta eius non amovi a me
2SAM|22|24|et ero perfectus cum eo et custodiam me ab iniquitate mea
2SAM|22|25|et restituet Dominus mihi secundum iustitiam meam et secundum munditiam manuum mearum in conspectu oculorum suorum
2SAM|22|26|cum sancto sanctus eris et cum robusto perfectus
2SAM|22|27|cum electo electus eris et cum perverso perverteris
2SAM|22|28|et populum pauperem salvum facies oculisque tuis excelsos humiliabis
2SAM|22|29|quia tu lucerna mea Domine et Domine inluminabis tenebras meas
2SAM|22|30|in te enim curram accinctus in Deo meo transiliam murum
2SAM|22|31|Deus inmaculata via eius eloquium Domini igne examinatum scutum est omnium sperantium in se
2SAM|22|32|quis est deus praeter Dominum et quis fortis praeter Deum nostrum
2SAM|22|33|Deus qui accingit me fortitudine et conplanavit perfectam viam meam
2SAM|22|34|coaequans pedes meos cervis et super excelsa mea statuens me
2SAM|22|35|docens manus meas ad proelium et conponens quasi arcum aereum brachia mea
2SAM|22|36|dedisti mihi clypeum salutis tuae et mansuetudo mea multiplicavit me
2SAM|22|37|dilatabis gressus meos subtus me et non deficient tali mei
2SAM|22|38|persequar inimicos meos et conteram et non revertar donec consumam eos
2SAM|22|39|consumam eos et confringam ut non consurgant cadent sub pedibus meis
2SAM|22|40|accinxisti me fortitudine ad proelium incurvabis resistentes mihi sub me
2SAM|22|41|inimicos meos dedisti mihi dorsum odientes me et disperdam eos
2SAM|22|42|clamabunt et non erit qui salvet ad Dominum et non exaudiet eos
2SAM|22|43|delebo eos ut pulverem terrae quasi lutum platearum comminuam eos atque conpingam
2SAM|22|44|salvabis me a contradictionibus populi mei custodies in caput gentium populus quem ignoro serviet mihi
2SAM|22|45|filii alieni resistent mihi auditu auris oboedient mihi
2SAM|22|46|filii alieni defluxerunt et contrahentur in angustiis suis
2SAM|22|47|vivit Dominus et benedictus Deus meus et exaltabitur Deus fortis salutis meae
2SAM|22|48|Deus qui das vindictas mihi et deicis populos sub me
2SAM|22|49|qui educis me ab inimicis meis et a resistentibus mihi elevas me a viro iniquo liberabis me
2SAM|22|50|propterea confitebor tibi Domine in gentibus et nomini tuo cantabo
2SAM|22|51|magnificanti salutes regis sui et facienti misericordiam christo suo David et semini eius in sempiternum
2SAM|23|1|haec autem sunt verba novissima quae dixit David filius Isai dixit vir cui constitutum est de christo Dei Iacob egregius psalta Israhel
2SAM|23|2|spiritus Domini locutus est per me et sermo eius per linguam meam
2SAM|23|3|dixit Deus Israhel mihi locutus est Fortis Israhel dominator hominum iustus dominator in timore Dei
2SAM|23|4|sicut lux aurorae oriente sole mane absque nubibus rutilat et sicut pluviis germinat herba de terra
2SAM|23|5|nec tanta est domus mea apud Deum ut pactum aeternum iniret mecum firmum in omnibus atque munitum cuncta enim salus mea et omnis voluntas nec est quicquam ex ea quod non germinet
2SAM|23|6|praevaricatores autem quasi spinae evellentur universi quae non tolluntur manibus
2SAM|23|7|et si quis tangere voluerit eas armabitur ferro et ligno lanceato igneque succensae conburentur usque ad nihilum
2SAM|23|8|haec nomina fortium David Sedens in cathedra sapientissimus princeps inter tres ipse est quasi tenerrimus ligni vermiculus qui octingentos interfecit impetu uno
2SAM|23|9|post hunc Eleazar filius patrui eius Ahoi inter tres fortes qui erant cum David quando exprobraverunt Philisthim et congregati sunt illuc in proelium
2SAM|23|10|cumque ascendissent viri Israhel ipse stetit et percussit Philistheos donec deficeret manus eius et obrigesceret cum gladio fecitque Dominus salutem magnam in die illa et populus qui fugerat reversus est ad caesorum spolia detrahenda
2SAM|23|11|et post hunc Semma filius Age de Arari et congregati sunt Philisthim in statione erat quippe ibi ager plenus lente cumque fugisset populus a facie Philisthim
2SAM|23|12|stetit ille in medio agri et tuitus est eum percussitque Philistheos et fecit Dominus salutem magnam
2SAM|23|13|necnon ante descenderant tres qui erant principes inter triginta et venerant tempore messis ad David in speluncam Odollam castra autem Philisthim erant posita in valle Gigantum
2SAM|23|14|et David erat in praesidio porro statio Philisthinorum tunc erat in Bethleem
2SAM|23|15|desideravit igitur David et ait si quis mihi daret potum aquae de cisterna quae est in Bethleem iuxta portam
2SAM|23|16|inruperunt ergo tres fortes castra Philisthinorum et hauserunt aquam de cisterna Bethleem quae erat iuxta portam et adtulerunt ad David at ille noluit bibere sed libavit illam Domino
2SAM|23|17|dicens propitius mihi sit Dominus ne faciam hoc num sanguinem hominum istorum qui profecti sunt et animarum periculum bibam noluit ergo bibere haec fecerunt tres robustissimi
2SAM|23|18|Abisai quoque frater Ioab filius Sarviae princeps erat de tribus ipse est qui elevavit hastam suam contra trecentos quos interfecit nominatus in tribus
2SAM|23|19|et inter tres nobilior eratque eorum princeps sed usque ad tres primos non pervenerat
2SAM|23|20|et Banaias filius Ioiada viri fortissimi magnorum operum de Capsehel ipse percussit duos leones Moab et ipse descendit et percussit leonem in media cisterna diebus nivis
2SAM|23|21|ipse quoque interfecit virum aegyptium virum dignum spectaculo habentem in manu hastam itaque cum descendisset ad eum in virga vi extorsit hastam de manu Aegyptii et interfecit eum hasta sua
2SAM|23|22|haec fecit Banaias filius Ioiadae
2SAM|23|23|et ipse nominatus inter tres robustos qui erant inter triginta nobiliores verumtamen usque ad tres non pervenerat fecitque eum David sibi auricularium a secreto
2SAM|23|24|Asahel frater Ioab inter triginta Eleanan filius patrui eius de Bethleem
2SAM|23|25|Semma de Arari Helica de Arodi
2SAM|23|26|Helas de Felthi Hira filius Aces de Thecua
2SAM|23|27|Abiezer de Anathoth Mobonnai de Usathi
2SAM|23|28|Selmon Aohites Maharai Netophathites
2SAM|23|29|Heled filius Banaa et ipse Netophathites Hithai filius Ribai de Gebeeth filiorum Beniamin
2SAM|23|30|Banahi Aufrathonites Heddai de torrente Gaas
2SAM|23|31|Abialbon Arbathites Azmaveth de Beromi
2SAM|23|32|Eliaba de Salboni filii Iasen Ionathan
2SAM|23|33|Semma de Horodi Haiam filius Sarar Arorites
2SAM|23|34|Elifeleth filius Aasbai filii Maachathi Heliam filius Ahitofel Gelonites
2SAM|23|35|Esrai de Carmelo Farai de Arbi
2SAM|23|36|Igaal filius Nathan de Soba Bonni de Gaddi
2SAM|23|37|Selech de Ammoni Naharai Berothites armiger Ioab filii Sarviae
2SAM|23|38|Hira Hiethrites Gareb et ipse Hiethrites
2SAM|23|39|Urias Hettheus omnes triginta septem
2SAM|24|1|et addidit furor Domini irasci contra Israhel commovitque David in eis dicentem vade numera Israhel et Iudam
2SAM|24|2|dixitque rex ad Ioab principem exercitus sui perambula omnes tribus Israhel a Dan usque Bersabee et numerate populum ut sciam numerum eius
2SAM|24|3|dixitque Ioab regi adaugeat Dominus Deus tuus ad populum quantus nunc est iterumque centuplicet in conspectu domini mei regis sed quid sibi dominus meus rex vult in re huiuscemodi
2SAM|24|4|obtinuit autem sermo regis verba Ioab et principum exercitus egressusque est Ioab et principes militum a facie regis ut numerarent populum Israhel
2SAM|24|5|cumque pertransissent Iordanem venerunt in Aroer ad dextram urbis quae est in valle Gad
2SAM|24|6|et per Iazer transierunt in Galaad et in terram inferiorem Hodsi et venerunt in Dan silvestria circumeuntesque iuxta Sidonem
2SAM|24|7|transierunt propter moenia Tyri et omnem terram Hevei et Chananei veneruntque ad meridiem Iuda in Bersabee
2SAM|24|8|et lustrata universa terra adfuerunt post novem menses et viginti dies in Hierusalem
2SAM|24|9|dedit ergo Ioab numerum descriptionis populi regi et inventa sunt de Israhel octingenta milia virorum fortium qui educerent gladium et de Iuda quingenta milia pugnatorum
2SAM|24|10|percussit autem cor David eum postquam numeratus est populus et dixit David ad Dominum peccavi valde in hoc facto sed precor Domine ut transferas iniquitatem servi tui quia stulte egi nimis
2SAM|24|11|surrexit itaque David mane et sermo Domini factus est ad Gad propheten et videntem David dicens
2SAM|24|12|vade et loquere ad David haec dicit Dominus trium tibi datur optio elige unum quod volueris ex his ut faciam tibi
2SAM|24|13|cumque venisset Gad ad David nuntiavit ei dicens aut septem annis veniet tibi fames in terra tua aut tribus mensibus fugies adversarios tuos et illi persequentur aut certe tribus diebus erit pestilentia in terra tua nunc ergo delibera et vide quem respondeam ei qui me misit sermonem
2SAM|24|14|dixit autem David ad Gad artor nimis sed melius est ut incidam in manu Domini multae enim misericordiae eius sunt quam in manu hominis
2SAM|24|15|inmisitque Dominus pestilentiam in Israhel de mane usque ad tempus constitutum et mortui sunt ex populo a Dan usque Bersabee septuaginta milia virorum
2SAM|24|16|cumque extendisset manum angelus Dei super Hierusalem ut disperderet eam misertus est Dominus super adflictione et ait angelo percutienti populum sufficit nunc contine manum tuam erat autem angelus Domini iuxta aream Areuna Iebusei
2SAM|24|17|dixitque David ad Dominum cum vidisset angelum caedentem populum ego sum qui peccavi ego inique egi isti qui oves sunt quid fecerunt vertatur obsecro manus tua contra me et contra domum patris mei
2SAM|24|18|venit autem Gad ad David in die illa et dixit ei ascende constitue Domino altare in area Areuna Iebusei
2SAM|24|19|et ascendit David iuxta sermonem Gad quem praeceperat ei Dominus
2SAM|24|20|conspiciensque Areuna animadvertit regem et servos eius transire ad se
2SAM|24|21|et egressus adoravit regem prono vultu in terra et ait quid causae est ut veniat dominus meus rex ad servum suum cui David ait ut emam a te aream et aedificem altare Domino et cesset interfectio quae grassatur in populo
2SAM|24|22|et ait Areuna ad David accipiat et offerat dominus meus rex sicut ei placet habes boves in holocaustum et plaustrum et iuga boum in usum lignorum
2SAM|24|23|omnia dedit Areuna rex regi dixitque Areuna ad regem Dominus Deus tuus suscipiat votum tuum
2SAM|24|24|cui respondens rex ait nequaquam ut vis sed emam pretio a te et non offeram Domino Deo meo holocausta gratuita emit ergo David aream et boves argenti siclis quinquaginta
2SAM|24|25|et aedificavit ibi David altare Domino et obtulit holocausta et pacifica et repropitiatus est Dominus terrae et cohibita est plaga ab Israhel
