2COR|1|1|Paul, an apostle of Christ Jesus by the will of God, and Timothy our brother, To the church of God that is at Corinth, with all the saints who are in the whole of Achaia:
2COR|1|2|Grace to you and peace from God our Father and the Lord Jesus Christ.
2COR|1|3|Blessed be the God and Father of our Lord Jesus Christ, the Father of mercies and God of all comfort,
2COR|1|4|who comforts us in all our affliction, so that we may be able to comfort those who are in any affliction, with the comfort with which we ourselves are comforted by God.
2COR|1|5|For as we share abundantly in Christ's sufferings, so through Christ we share abundantly in comfort too.
2COR|1|6|If we are afflicted, it is for your comfort and salvation; and if we are comforted, it is for your comfort, which you experience when you patiently endure the same sufferings that we suffer.
2COR|1|7|Our hope for you is unshaken, for we know that as you share in our sufferings, you will also share in our comfort.
2COR|1|8|For we do not want you to be ignorant, brothers, of the affliction we experienced in Asia. For we were so utterly burdened beyond our strength that we despaired of life itself.
2COR|1|9|Indeed, we felt that we had received the sentence of death. But that was to make us rely not on ourselves but on God who raises the dead.
2COR|1|10|He delivered us from such a deadly peril, and he will deliver us. On him we have set our hope that he will deliver us again.
2COR|1|11|You also must help us by prayer, so that many will give thanks on our behalf for the blessing granted us through the prayers of many.
2COR|1|12|For our boast is this: the testimony of our conscience that we behaved in the world with simplicity and godly sincerity, not by earthly wisdom but by the grace of God, and supremely so toward you.
2COR|1|13|For we are not writing to you anything other than what you read and acknowledge and I hope you will fully acknowledge-
2COR|1|14|just as you did partially acknowledge us, that on the day of our Lord Jesus you will boast of us as we will boast of you.
2COR|1|15|Because I was sure of this, I wanted to come to you first, so that you might have a second experience of grace.
2COR|1|16|I wanted to visit you on my way to Macedonia, and to come back to you from Macedonia and have you send me on my way to Judea.
2COR|1|17|Was I vacillating when I wanted to do this? Do I make my plans according to the flesh, ready to say "Yes, yes" and "No, no" at the same time?
2COR|1|18|As surely as God is faithful, our word to you has not been Yes and No.
2COR|1|19|For the Son of God, Jesus Christ, whom we proclaimed among you, Silvanus and Timothy and I, was not Yes and No, but in him it is always Yes.
2COR|1|20|For all the promises of God find their Yes in him. That is why it is through him that we utter our Amen to God for his glory.
2COR|1|21|And it is God who establishes us with you in Christ, and has anointed us,
2COR|1|22|and who has also put his seal on us and given us his Spirit in our hearts as a guarantee.
2COR|1|23|But I call God to witness against me- it was to spare you that I refrained from coming again to Corinth.
2COR|1|24|Not that we lord it over your faith, but we work with you for your joy, for you stand firm in your faith.
2COR|2|1|For I made up my mind not to make another painful visit to you.
2COR|2|2|For if I cause you pain, who is there to make me glad but the one whom I have pained?
2COR|2|3|And I wrote as I did, so that when I came I might not suffer pain from those who should have made me rejoice, for I felt sure of all of you, that my joy would be the joy of you all.
2COR|2|4|For I wrote to you out of much affliction and anguish of heart and with many tears, not to cause you pain but to let you know the abundant love that I have for you.
2COR|2|5|Now if anyone has caused pain, he has caused it not to me, but in some measure- not to put it too severely- to all of you.
2COR|2|6|For such a one, this punishment by the majority is enough,
2COR|2|7|so you should rather turn to forgive and comfort him, or he may be overwhelmed by excessive sorrow.
2COR|2|8|So I beg you to reaffirm your love for him.
2COR|2|9|For this is why I wrote, that I might test you and know whether you are obedient in everything.
2COR|2|10|Anyone whom you forgive, I also forgive. What I have forgiven, if I have forgiven anything, has been for your sake in the presence of Christ,
2COR|2|11|so that we would not be outwitted by Satan; for we are not ignorant of his designs.
2COR|2|12|When I came to Troas to preach the gospel of Christ, even though a door was opened for me in the Lord,
2COR|2|13|my spirit was not at rest because I did not find my brother Titus there. So I took leave of them and went on to Macedonia.
2COR|2|14|But thanks be to God, who in Christ always leads us in triumphal procession, and through us spreads the fragrance of the knowledge of him everywhere.
2COR|2|15|For we are the aroma of Christ to God among those who are being saved and among those who are perishing,
2COR|2|16|to one a fragrance from death to death, to the other a fragrance from life to life. Who is sufficient for these things?
2COR|2|17|For we are not, like so many, peddlers of God's word, but as men of sincerity, as commissioned by God, in the sight of God we speak in Christ.
2COR|3|1|Are we beginning to commend ourselves again? Or do we need, as some do, letters of recommendation to you, or from you?
2COR|3|2|You yourselves are our letter of recommendation, written on our hearts, to be known and read by all.
2COR|3|3|And you show that you are a letter from Christ delivered by us, written not with ink but with the Spirit of the living God, not on tablets of stone but on tablets of human hearts.
2COR|3|4|Such is the confidence that we have through Christ toward God.
2COR|3|5|Not that we are sufficient in ourselves to claim anything as coming from us, but our sufficiency is from God,
2COR|3|6|who has made us competent to be ministers of a new covenant, not of the letter but of the Spirit. For the letter kills, but the Spirit gives life.
2COR|3|7|Now if the ministry of death, carved in letters on stone, came with such glory that the Israelites could not gaze at Moses' face because of its glory, which was being brought to an end,
2COR|3|8|will not the ministry of the Spirit have even more glory?
2COR|3|9|For if there was glory in the ministry of condemnation, the ministry of righteousness must far exceed it in glory.
2COR|3|10|Indeed, in this case, what once had glory has come to have no glory at all, because of the glory that surpasses it.
2COR|3|11|For if what was being brought to an end came with glory, much more will what is permanent have glory.
2COR|3|12|Since we have such a hope, we are very bold,
2COR|3|13|not like Moses, who would put a veil over his face so that the Israelites might not gaze at the outcome of what was being brought to an end.
2COR|3|14|But their minds were hardened. For to this day, when they read the old covenant, that same veil remains unlifted, because only through Christ is it taken away.
2COR|3|15|Yes, to this day whenever Moses is read a veil lies over their hearts.
2COR|3|16|But when one turns to the Lord, the veil is removed.
2COR|3|17|Now the Lord is the Spirit, and where the Spirit of the Lord is, there is freedom.
2COR|3|18|And we all, with unveiled face, beholding the glory of the Lord, are being transformed into the same image from one degree of glory to another. For this comes from the Lord who is the Spirit.
2COR|4|1|Therefore, having this ministry by the mercy of God, we do not lose heart.
2COR|4|2|But we have renounced disgraceful, underhanded ways. We refuse to practice cunning or to tamper with God's word, but by the open statement of the truth we would commend ourselves to everyone's conscience in the sight of God.
2COR|4|3|And even if our gospel is veiled, it is veiled only to those who are perishing.
2COR|4|4|In their case the god of this world has blinded the minds of the unbelievers, to keep them from seeing the light of the gospel of the glory of Christ, who is the image of God.
2COR|4|5|For what we proclaim is not ourselves, but Jesus Christ as Lord, with ourselves as your servants for Jesus' sake.
2COR|4|6|For God, who said, "Let light shine out of darkness," has shone in our hearts to give the light of the knowledge of the glory of God in the face of Jesus Christ.
2COR|4|7|But we have this treasure in jars of clay, to show that the surpassing power belongs to God and not to us.
2COR|4|8|We are afflicted in every way, but not crushed; perplexed, but not driven to despair;
2COR|4|9|persecuted, but not forsaken; struck down, but not destroyed;
2COR|4|10|always carrying in the body the death of Jesus, so that the life of Jesus may also be manifested in our bodies.
2COR|4|11|For we who live are always being given over to death for Jesus' sake, so that the life of Jesus also may be manifested in our mortal flesh.
2COR|4|12|So death is at work in us, but life in you.
2COR|4|13|Since we have the same spirit of faith according to what has been written, "I believed, and so I spoke," we also believe, and so we also speak,
2COR|4|14|knowing that he who raised the Lord Jesus will raise us also with Jesus and bring us with you into his presence.
2COR|4|15|For it is all for your sake, so that as grace extends to more and more people it may increase thanksgiving, to the glory of God.
2COR|4|16|So we do not lose heart. Though our outer nature is wasting away, our inner nature is being renewed day by day.
2COR|4|17|For this slight momentary affliction is preparing for us an eternal weight of glory beyond all comparison,
2COR|4|18|as we look not to the things that are seen but to the things that are unseen. For the things that are seen are transient, but the things that are unseen are eternal.
2COR|5|1|For we know that if the tent, which is our earthly home, is destroyed, we have a building from God, a house not made with hands, eternal in the heavens.
2COR|5|2|For in this tent we groan, longing to put on our heavenly dwelling,
2COR|5|3|if indeed by putting it on we may not be found naked.
2COR|5|4|For while we are still in this tent, we groan, being burdened--not that we would be unclothed, but that we would be further clothed, so that what is mortal may be swallowed up by life.
2COR|5|5|He who has prepared us for this very thing is God, who has given us the Spirit as a guarantee.
2COR|5|6|So we are always of good courage. We know that while we are at home in the body we are away from the Lord,
2COR|5|7|for we walk by faith, not by sight.
2COR|5|8|Yes, we are of good courage, and we would rather be away from the body and at home with the Lord.
2COR|5|9|So whether we are at home or away, we make it our aim to please him.
2COR|5|10|For we must all appear before the judgment seat of Christ, so that each one may receive what is due for what he has done in the body, whether good or evil.
2COR|5|11|Therefore, knowing the fear of the Lord, we persuade others. But what we are is known to God, and I hope it is known also to your conscience.
2COR|5|12|We are not commending ourselves to you again but giving you cause to boast about us, so that you may be able to answer those who boast about outward appearance and not about what is in the heart.
2COR|5|13|For if we are beside ourselves, it is for God; if we are in our right mind, it is for you.
2COR|5|14|For the love of Christ controls us, because we have concluded this: that one has died for all, therefore all have died;
2COR|5|15|and he died for all, that those who live might no longer live for themselves but for him who for their sake died and was raised.
2COR|5|16|From now on, therefore, we regard no one according to the flesh. Even though we once regarded Christ according to the flesh, we regard him thus no longer.
2COR|5|17|Therefore, if anyone is in Christ, he is a new creation. The old has passed away; behold, the new has come.
2COR|5|18|All this is from God, who through Christ reconciled us to himself and gave us the ministry of reconciliation;
2COR|5|19|that is, in Christ God was reconciling the world to himself, not counting their trespasses against them, and entrusting to us the message of reconciliation.
2COR|5|20|Therefore, we are ambassadors for Christ, God making his appeal through us. We implore you on behalf of Christ, be reconciled to God.
2COR|5|21|For our sake he made him to be sin who knew no sin, so that in him we might become the righteousness of God.
2COR|6|1|Working together with him, then, we appeal to you not to receive the grace of God in vain.
2COR|6|2|For he says, "In a favorable time I listened to you, and in a day of salvation I have helped you." Behold, now is the favorable time; behold, now is the day of salvation.
2COR|6|3|We put no obstacle in anyone's way, so that no fault may be found with our ministry,
2COR|6|4|but as servants of God we commend ourselves in every way: by great endurance, in afflictions, hardships, calamities,
2COR|6|5|beatings, imprisonments, riots, labors, sleepless nights, hunger;
2COR|6|6|by purity, knowledge, patience, kindness, the Holy Spirit, genuine love,
2COR|6|7|by truthful speech, and the power of God; with the weapons of righteousness for the right hand and for the left;
2COR|6|8|through honor and dishonor, through slander and praise. We are treated as impostors, and yet are true;
2COR|6|9|as unknown, and yet well known; as dying, and behold, we live; as punished, and yet not killed;
2COR|6|10|as sorrowful, yet always rejoicing; as poor, yet making many rich; as having nothing, yet possessing everything.
2COR|6|11|We have spoken freely to you, Corinthians; our heart is wide open.
2COR|6|12|You are not restricted by us, but you are restricted in your own affections.
2COR|6|13|In return (I speak as to children) widen your hearts also.
2COR|6|14|Do not be unequally yoked with unbelievers. For what partnership has righteousness with lawlessness? Or what fellowship has light with darkness?
2COR|6|15|What accord has Christ with Belial? Or what portion does a believer share with an unbeliever?
2COR|6|16|What agreement has the temple of God with idols? For we are the temple of the living God; as God said, "I will make my dwelling among them and walk among them, and I will be their God, and they shall be my people.
2COR|6|17|Therefore go out from their midst, and be separate from them, says the Lord, and touch no unclean thing; then I will welcome you,
2COR|6|18|and I will be a father to you, and you shall be sons and daughters to me, says the Lord Almighty."
2COR|7|1|Since we have these promises, beloved, let us cleanse ourselves from every defilement of body and spirit, bringing holiness to completion in the fear of God.
2COR|7|2|Make room in your hearts for us. We have wronged no one, we have corrupted no one, we have taken advantage of no one.
2COR|7|3|I do not say this to condemn you, for I said before that you are in our hearts, to die together and to live together.
2COR|7|4|I am acting with great boldness toward you; I have great pride in you; I am filled with comfort. In all our affliction, I am overflowing with joy.
2COR|7|5|For even when we came into Macedonia, our bodies had no rest, but we were afflicted at every turn- fighting without and fear within.
2COR|7|6|But God, who comforts the downcast, comforted us by the coming of Titus,
2COR|7|7|and not only by his coming but also by the comfort with which he was comforted by you, as he told us of your longing, your mourning, your zeal for me, so that I rejoiced still more.
2COR|7|8|For even if I made you grieve with my letter, I do not regret it- though I did regret it, for I see that that letter grieved you, though only for a while.
2COR|7|9|As it is, I rejoice, not because you were grieved, but because you were grieved into repenting. For you felt a godly grief, so that you suffered no loss through us.
2COR|7|10|For godly grief produces a repentance that leads to salvation without regret, whereas worldly grief produces death.
2COR|7|11|For see what earnestness this godly grief has produced in you, but also what eagerness to clear yourselves, what indignation, what fear, what longing, what zeal, what punishment! At every point you have proved yourselves innocent in the matter.
2COR|7|12|So although I wrote to you, it was not for the sake of the one who did the wrong, nor for the sake of the one who suffered the wrong, but in order that your earnestness for us might be revealed to you in the sight of God.
2COR|7|13|Therefore we are comforted. And besides our own comfort, we rejoiced still more at the joy of Titus, because his spirit has been refreshed by you all.
2COR|7|14|For whatever boasts I made to him about you, I was not put to shame. But just as everything we said to you was true, so also our boasting before Titus has proved true.
2COR|7|15|And his affection for you is even greater, as he remembers the obedience of you all, how you received him with fear and trembling.
2COR|7|16|I rejoice, because I have perfect confidence in you.
2COR|8|1|We want you to know, brothers, about the grace of God that has been given among the churches of Macedonia,
2COR|8|2|for in a severe test of affliction, their abundance of joy and their extreme poverty have overflowed in a wealth of generosity on their part.
2COR|8|3|For they gave according to their means, as I can testify, and beyond their means, of their own free will,
2COR|8|4|begging us earnestly for the favor of taking part in the relief of the saints-
2COR|8|5|and this, not as we expected, but they gave themselves first to the Lord and then by the will of God to us.
2COR|8|6|Accordingly, we urged Titus that as he had started, so he should complete among you this act of grace.
2COR|8|7|But as you excel in everything- in faith, in speech, in knowledge, in all earnestness, and in our love for you- see that you excel in this act of grace also.
2COR|8|8|I say this not as a command, but to prove by the earnestness of others that your love also is genuine.
2COR|8|9|For you know the grace of our Lord Jesus Christ, that though he was rich, yet for your sake he became poor, so that you by his poverty might become rich.
2COR|8|10|And in this matter I give my judgment: this benefits you, who a year ago started not only to do this work but also to desire to do it.
2COR|8|11|So now finish doing it as well, so that your readiness in desiring it may be matched by your completing it out of what you have.
2COR|8|12|For if the readiness is there, it is acceptable according to what a person has, not according to what he does not have.
2COR|8|13|I do not mean that others should be eased and you burdened, but that as a matter of fairness
2COR|8|14|your abundance at the present time should supply their need, so that their abundance may supply your need, that there may be fairness.
2COR|8|15|As it is written, "Whoever gathered much had nothing left over, and whoever gathered little had no lack."
2COR|8|16|But thanks be to God, who put into the heart of Titus the same earnest care I have for you.
2COR|8|17|For he not only accepted our appeal, but being himself very earnest he is going to you of his own accord.
2COR|8|18|With him we are sending the brother who is famous among all the churches for his preaching of the gospel.
2COR|8|19|And not only that, but he has been appointed by the churches to travel with us as we carry out this act of grace that is being ministered by us, for the glory of the Lord himself and to show our good will.
2COR|8|20|We take this course so that no one should blame us about this generous gift that is being administered by us,
2COR|8|21|for we aim at what is honorable not only in the Lord's sight but also in the sight of man.
2COR|8|22|And with them we are sending our brother whom we have often tested and found earnest in many matters, but who is now more earnest than ever because of his great confidence in you.
2COR|8|23|As for Titus, he is my partner and fellow worker for your benefit. And as for our brothers, they are messengers of the churches, the glory of Christ.
2COR|8|24|So give proof before the churches of your love and of our boasting about you to these men.
2COR|9|1|Now it is superfluous for me to write to you about the ministry for the saints,
2COR|9|2|for I know your readiness, of which I boast about you to the people of Macedonia, saying that Achaia has been ready since last year. And your zeal has stirred up most of them.
2COR|9|3|But I am sending the brothers so that our boasting about you may not prove vain in this matter, so that you may be ready, as I said you would be.
2COR|9|4|Otherwise, if some Macedonians come with me and find that you are not ready, we would be humiliated- to say nothing of you- for being so confident.
2COR|9|5|So I thought it necessary to urge the brothers to go on ahead to you and arrange in advance for the gift you have promised, so that it may be ready as a willing gift, not as an exaction.
2COR|9|6|The point is this: whoever sows sparingly will also reap sparingly, and whoever sows bountifully will also reap bountifully.
2COR|9|7|Each one must give as he has made up his mind, not reluctantly or under compulsion, for God loves a cheerful giver.
2COR|9|8|And God is able to make all grace abound to you, so that having all sufficiency in all things at all times, you may abound in every good work.
2COR|9|9|As it is written, "He has distributed freely, he has given to the poor; his righteousness endures forever."
2COR|9|10|He who supplies seed to the sower and bread for food will supply and multiply your seed for sowing and increase the harvest of your righteousness.
2COR|9|11|You will be enriched in every way for all your generosity, which through us will produce thanksgiving to God.
2COR|9|12|For the ministry of this service is not only supplying the needs of the saints, but is also overflowing in many thanksgivings to God.
2COR|9|13|By their approval of this service, they will glorify God because of your submission flowing from your confession of the gospel of Christ, and the generosity of your contribution for them and for all others,
2COR|9|14|while they long for you and pray for you, because of the surpassing grace of God upon you.
2COR|9|15|Thanks be to God for his inexpressible gift!
2COR|10|1|I, Paul, myself entreat you, by the meekness and gentleness of Christ- I who am humble when face to face with you, but bold toward you when I am away!-
2COR|10|2|I beg of you that when I am present I may not have to show boldness with such confidence as I count on showing against some who suspect us of walking according to the flesh.
2COR|10|3|For though we walk in the flesh, we are not waging war according to the flesh.
2COR|10|4|For the weapons of our warfare are not of the flesh but have divine power to destroy strongholds. We destroy arguments
2COR|10|5|and every lofty opinion raised against the knowledge of God, and take every thought captive to obey Christ,
2COR|10|6|being ready to punish every disobedience, when your obedience is complete.
2COR|10|7|Look at what is before your eyes. If anyone is confident that he is Christ's, let him remind himself that just as he is Christ's, so also are we.
2COR|10|8|For even if I boast a little too much of our authority, which the Lord gave for building you up and not for destroying you, I will not be ashamed.
2COR|10|9|I do not want to appear to be frightening you with my letters.
2COR|10|10|For they say, "His letters are weighty and strong, but his bodily presence is weak, and his speech of no account."
2COR|10|11|Let such a person understand that what we say by letter when absent, we do when present.
2COR|10|12|Not that we dare to classify or compare ourselves with some of those who are commending themselves. But when they measure themselves by one another and compare themselves with one another, they are without understanding.
2COR|10|13|But we will not boast beyond limits, but will boast only with regard to the area of influence God assigned to us, to reach even to you.
2COR|10|14|For we are not overextending ourselves, as though we did not reach you. We were the first to come all the way to you with the gospel of Christ.
2COR|10|15|We do not boast beyond limit in the labors of others. But our hope is that as your faith increases, our area of influence among you may be greatly enlarged,
2COR|10|16|so that we may preach the gospel in lands beyond you, without boasting of work already done in another's area of influence.
2COR|10|17|"Let the one who boasts, boast in the Lord."
2COR|10|18|For it is not the one who commends himself who is approved, but the one whom the Lord commends.
2COR|11|1|I wish you would bear with me in a little foolishness. Do bear with me!
2COR|11|2|I feel a divine jealousy for you, for I betrothed you to one husband, to present you as a pure virgin to Christ.
2COR|11|3|But I am afraid that as the serpent deceived Eve by his cunning, your thoughts will be led astray from a sincere and pure devotion to Christ.
2COR|11|4|For if someone comes and proclaims another Jesus than the one we proclaimed, or if you receive a different spirit from the one you received, or if you accept a different gospel from the one you accepted, you put up with it readily enough.
2COR|11|5|I consider that I am not in the least inferior to these super-apostles.
2COR|11|6|Even if I am unskilled in speaking, I am not so in knowledge; indeed, in every way we have made this plain to you in all things.
2COR|11|7|Or did I commit a sin in humbling myself so that you might be exalted, because I preached God's gospel to you free of charge?
2COR|11|8|I robbed other churches by accepting support from them in order to serve you.
2COR|11|9|And when I was with you and was in need, I did not burden anyone, for the brothers who came from Macedonia supplied my need. So I refrained and will refrain from burdening you in any way.
2COR|11|10|As the truth of Christ is in me, this boasting of mine will not be silenced in the regions of Achaia.
2COR|11|11|And why? Because I do not love you? God knows I do!
2COR|11|12|And what I do I will continue to do, in order to undermine the claim of those who would like to claim that in their boasted mission they work on the same terms as we do.
2COR|11|13|For such men are false apostles, deceitful workmen, disguising themselves as apostles of Christ.
2COR|11|14|And no wonder, for even Satan disguises himself as an angel of light.
2COR|11|15|So it is no surprise if his servants, also, disguise themselves as servants of righteousness. Their end will correspond to their deeds.
2COR|11|16|I repeat, let no one think me foolish. But even if you do, accept me as a fool, so that I too may boast a little.
2COR|11|17|What I am saying with this boastful confidence, I say not with the Lord's authority but as a fool.
2COR|11|18|Since many boast according to the flesh, I too will boast.
2COR|11|19|For you gladly bear with fools, being wise yourselves!
2COR|11|20|For you bear it if someone makes slaves of you, or devours you, or takes advantage of you, or puts on airs, or strikes you in the face.
2COR|11|21|To my shame, I must say, we were too weak for that! But whatever anyone else dares to boast of- I am speaking as a fool- I also dare to boast of that.
2COR|11|22|Are they Hebrews? So am I. Are they Israelites? So am I. Are they offspring of Abraham? So am I.
2COR|11|23|Are they servants of Christ? I am a better one- I am talking like a madman- with far greater labors, far more imprisonments, with countless beatings, and often near death.
2COR|11|24|Five times I received at the hands of the Jews the forty lashes less one.
2COR|11|25|Three times I was beaten with rods. Once I was stoned. Three times I was shipwrecked; a night and a day I was adrift at sea;
2COR|11|26|on frequent journeys, in danger from rivers, danger from robbers, danger from my own people, danger from Gentiles, danger in the city, danger in the wilderness, danger at sea, danger from false brothers;
2COR|11|27|in toil and hardship, through many a sleepless night, in hunger and thirst, often without food, in cold and exposure.
2COR|11|28|And, apart from other things, there is the daily pressure on me of my anxiety for all the churches.
2COR|11|29|Who is weak, and I am not weak? Who is made to fall, and I am not indignant?
2COR|11|30|If I must boast, I will boast of the things that show my weakness.
2COR|11|31|The God and Father of the Lord Jesus, he who is blessed forever, knows that I am not lying.
2COR|11|32|At Damascus, the governor under King Aretas was guarding the city of Damascus in order to seize me,
2COR|11|33|but I was let down in a basket through a window in the wall and escaped his hands.
2COR|12|1|I must go on boasting. Though there is nothing to be gained by it, I will go on to visions and revelations of the Lord.
2COR|12|2|I know a man in Christ who fourteen years ago was caught up to the third heaven- whether in the body or out of the body I do not know, God knows.
2COR|12|3|And I know that this man was caught up into paradise- whether in the body or out of the body I do not know, God knows-
2COR|12|4|and he heard things that cannot be told, which man may not utter.
2COR|12|5|On behalf of this man I will boast, but on my own behalf I will not boast, except of my weaknesses.
2COR|12|6|Though if I should wish to boast, I would not be a fool, for I would be speaking the truth. But I refrain from it, so that no one may think more of me than he sees in me or hears from me.
2COR|12|7|So to keep me from being too elated by the surpassing greatness of the revelations, a thorn was given me in the flesh, a messenger of Satan to harass me, to keep me from being too elated.
2COR|12|8|Three times I pleaded with the Lord about this, that it should leave me.
2COR|12|9|But he said to me, "My grace is sufficient for you, for my power is made perfect in weakness." Therefore I will boast all the more gladly of my weaknesses, so that the power of Christ may rest upon me.
2COR|12|10|For the sake of Christ, then, I am content with weaknesses, insults, hardships, persecutions, and calamities. For when I am weak, then I am strong.
2COR|12|11|I have been a fool! You forced me to it, for I ought to have been commended by you. For I was not at all inferior to these super-apostles, even though I am nothing.
2COR|12|12|The signs of a true apostle were performed among you with utmost patience, with signs and wonders and mighty works.
2COR|12|13|For in what were you less favored than the rest of the churches, except that I myself did not burden you? Forgive me this wrong!
2COR|12|14|Here for the third time I am ready to come to you. And I will not be a burden, for I seek not what is yours but you. For children are not obligated to save up for their parents, but parents for their children.
2COR|12|15|I will most gladly spend and be spent for your souls. If I love you more, am I to be loved less?
2COR|12|16|But granting that I myself did not burden you, I was crafty, you say, and got the better of you by deceit.
2COR|12|17|Did I take advantage of you through any of those whom I sent to you?
2COR|12|18|I urged Titus to go, and sent the brother with him. Did Titus take advantage of you? Did we not act in the same spirit? Did we not take the same steps?
2COR|12|19|Have you been thinking all along that we have been defending ourselves to you? It is in the sight of God that we have been speaking in Christ, and all for your upbuilding, beloved.
2COR|12|20|For I fear that perhaps when I come I may find you not as I wish, and that you may find me not as you wish- that perhaps there may be quarreling, jealousy, anger, hostility, slander, gossip, conceit, and disorder.
2COR|12|21|I fear that when I come again my God may humble me before you, and I may have to mourn over many of those who sinned earlier and have not repented of the impurity, sexual immorality, and sensuality that they have practiced.
2COR|13|1|This is the third time I am coming to you. Every charge must be established by the evidence of two or three witnesses.
2COR|13|2|I warned those who sinned before and all the others, and I warn them now while absent, as I did when present on my second visit, that if I come again I will not spare them-
2COR|13|3|since you seek proof that Christ is speaking in me. He is not weak in dealing with you, but is powerful among you.
2COR|13|4|For he was crucified in weakness, but lives by the power of God. For we also are weak in him, but in dealing with you we will live with him by the power of God.
2COR|13|5|Examine yourselves, to see whether you are in the faith. Test yourselves. Or do you not realize this about yourselves, that Jesus Christ is in you?- unless indeed you fail to meet the test!
2COR|13|6|I hope you will find out that we have not failed the test.
2COR|13|7|But we pray to God that you may not do wrong- not that we may appear to have met the test, but that you may do what is right, though we may seem to have failed.
2COR|13|8|For we cannot do anything against the truth, but only for the truth.
2COR|13|9|For we are glad when we are weak and you are strong. Your restoration is what we pray for.
2COR|13|10|For this reason I write these things while I am away from you, that when I come I may not have to be severe in my use of the authority that the Lord has given me for building up and not for tearing down.
2COR|13|11|Finally, brothers, rejoice. Aim for restoration, comfort one another, agree with one another, live in peace; and the God of love and peace will be with you.
2COR|13|12|Greet one another with a holy kiss.
2COR|13|13|All the saints greet you.
2COR|13|14|The grace of the Lord Jesus Christ and the love of God and the fellowship of the Holy Spirit be with you all.
