EZEK|1|1|И было в тридцатый год, в четвертый [месяц], в пятый [день] месяца, когда я находился среди переселенцев при реке Ховаре, отверзлись небеса, и я видел видения Божии.
EZEK|1|2|В пятый [день] месяца (это был пятый год от пленения царя Иоакима),
EZEK|1|3|было слово Господне к Иезекиилю, сыну Вузия, священнику, в земле Халдейской, при реке Ховаре; и была на нем там рука Господня.
EZEK|1|4|И я видел, и вот, бурный ветер шел от севера, великое облако и клубящийся огонь, и сияние вокруг него,
EZEK|1|5|а из средины его как бы свет пламени из средины огня; и из средины его видно было подобие четырех животных, – и таков был вид их: облик их был, как у человека;
EZEK|1|6|и у каждого четыре лица, и у каждого из них четыре крыла;
EZEK|1|7|а ноги их – ноги прямые, и ступни ног их – как ступня ноги у тельца, и сверкали, как блестящая медь.
EZEK|1|8|И руки человеческие были под крыльями их, на четырех сторонах их;
EZEK|1|9|и лица у них и крылья у них – у всех четырех; крылья их соприкасались одно к другому; во время шествия своего они не оборачивались, а шли каждое по направлению лица своего.
EZEK|1|10|Подобие лиц их – лице человека и лице льва с правой стороны у всех их четырех; а с левой стороны лице тельца у всех четырех и лице орла у всех четырех.
EZEK|1|11|И лица их и крылья их сверху были разделены, но у каждого два крыла соприкасались одно к другому, а два покрывали тела их.
EZEK|1|12|И шли они, каждое в ту сторону, которая пред лицем его; куда дух хотел идти, туда и шли; во время шествия своего не оборачивались.
EZEK|1|13|И вид этих животных был как вид горящих углей, как вид лампад; [огонь] ходил между животными, и сияние от огня и молния исходила из огня.
EZEK|1|14|И животные быстро двигались туда и сюда, как сверкает молния.
EZEK|1|15|И смотрел я на животных, и вот, на земле подле этих животных по одному колесу перед четырьмя лицами их.
EZEK|1|16|Вид колес и устроение их – как вид топаза, и подобие у всех четырех одно; и по виду их и по устроению их казалось, будто колесо находилось в колесе.
EZEK|1|17|Когда они шли, шли на четыре свои стороны; во время шествия не оборачивались.
EZEK|1|18|А ободья их – высоки и страшны были они; ободья их у всех четырех вокруг полны были глаз.
EZEK|1|19|И когда шли животные, шли и колеса подле [них]; а когда животные поднимались от земли, тогда поднимались и колеса.
EZEK|1|20|Куда дух хотел идти, туда шли и они; куда бы ни пошел дух, и колеса поднимались наравне с ними, ибо дух животных [был] в колесах.
EZEK|1|21|Когда шли те, шли и они; и когда те стояли, стояли и они; и когда те поднимались от земли, тогда наравне с ними поднимались и колеса, ибо дух животных [был] в колесах.
EZEK|1|22|Над головами животных было подобие свода, как вид изумительного кристалла, простертого сверху над головами их.
EZEK|1|23|А под сводом простирались крылья их прямо одно к другому, и у каждого были два крыла, которые покрывали их, у каждого два крыла покрывали тела их.
EZEK|1|24|И когда они шли, я слышал шум крыльев их, как бы шум многих вод, как бы глас Всемогущего, сильный шум, как бы шум в воинском стане; [а] когда они останавливались, опускали крылья свои.
EZEK|1|25|И голос был со свода, который над головами их; когда они останавливались, тогда опускали крылья свои.
EZEK|1|26|А над сводом, который над головами их, [было] подобие престола по виду как бы из камня сапфира; а над подобием престола было как бы подобие человека вверху на нем.
EZEK|1|27|И видел я как бы пылающий металл, как бы вид огня внутри него вокруг; от вида чресл его и выше и от вида чресл его и ниже я видел как бы некий огонь, и сияние [было] вокруг него.
EZEK|1|28|В каком виде бывает радуга на облаках во время дождя, такой вид имело это сияние кругом.
EZEK|2|1|Такое было видение подобия славы Господней. Увидев это, я пал на лице свое, и слышал глас Глаголющего, и Он сказал мне: сын человеческий! стань на ноги твои, и Я буду говорить с тобою.
EZEK|2|2|И когда Он говорил мне, вошел в меня дух и поставил меня на ноги мои, и я слышал Говорящего мне.
EZEK|2|3|И Он сказал мне: сын человеческий! Я посылаю тебя к сынам Израилевым, к людям непокорным, которые возмутились против Меня; они и отцы их изменники предо Мною до сего самого дня.
EZEK|2|4|И эти сыны с огрубелым лицем и с жестоким сердцем; к ним Я посылаю тебя, и ты скажешь им: "так говорит Господь Бог!"
EZEK|2|5|Будут ли они слушать, или не будут, ибо они мятежный дом; но пусть знают, что был пророк среди них.
EZEK|2|6|А ты, сын человеческий, не бойся их и не бойся речей их, если они волчцами и тернами будут для тебя, и ты будешь жить у скорпионов; не бойся речей их и не страшись лица их, ибо они мятежный дом;
EZEK|2|7|и говори им слова Мои, будут ли они слушать, или не будут, ибо они упрямы.
EZEK|2|8|Ты же, сын человеческий, слушай, что Я буду говорить тебе; не будь упрям, как этот мятежный дом; открой уста твои и съешь, что Я дам тебе.
EZEK|2|9|И увидел я, и вот, рука простерта ко мне, и вот, в ней книжный свиток.
EZEK|2|10|И Он развернул его передо мною, и вот, свиток исписан был внутри и снаружи, и написано на нем: "плач, и стон, и горе".
EZEK|3|1|И сказал мне: сын человеческий! съешь, что перед тобою, съешь этот свиток, и иди, говори дому Израилеву.
EZEK|3|2|Тогда я открыл уста мои, и Он дал мне съесть этот свиток;
EZEK|3|3|и сказал мне: сын человеческий! напитай чрево твое и наполни внутренность твою этим свитком, который Я даю тебе; и я съел, и было в устах моих сладко, как мед.
EZEK|3|4|И Он сказал мне: сын человеческий! встань и иди к дому Израилеву, и говори им Моими словами;
EZEK|3|5|ибо не к народу с речью невнятною и с непонятным языком ты посылаешься, но к дому Израилеву,
EZEK|3|6|не к народам многим с невнятною речью и с непонятным языком, которых слов ты не разумел бы; да если бы Я послал тебя и к ним, то они послушались бы тебя;
EZEK|3|7|а дом Израилев не захочет слушать тебя; ибо они не хотят слушать Меня, потому что весь дом Израилев с крепким лбом и жестоким сердцем.
EZEK|3|8|Вот, Я сделал и твое лице крепким против лиц их, и твое чело крепким против их лба.
EZEK|3|9|Как алмаз, который крепче камня, сделал Я чело твое; не бойся их и не страшись перед лицем их, ибо они мятежный дом.
EZEK|3|10|И сказал мне: сын человеческий! все слова Мои, которые буду говорить тебе, прими сердцем твоим и выслушай ушами твоими;
EZEK|3|11|встань и пойди к переселенным, к сынам народа твоего, и говори к ним, и скажи им: "так говорит Господь Бог!" будут ли они слушать, или не будут.
EZEK|3|12|И поднял меня дух; и я слышал позади себя великий громовой голос: "благословенна слава Господа от места своего!"
EZEK|3|13|и также шум крыльев животных, соприкасающихся одно к другому, и стук колес подле них, и звук сильного грома.
EZEK|3|14|И дух поднял меня, и взял меня. И шел я в огорчении, с встревоженным духом; и рука Господня была крепко на мне.
EZEK|3|15|И пришел я к переселенным в Тел–Авив, живущим при реке Ховаре, и остановился там, где они жили, и провел среди них семь дней в изумлении.
EZEK|3|16|По прошествии же семи дней было ко мне слово Господне:
EZEK|3|17|сын человеческий! Я поставил тебя стражем дому Израилеву, и ты будешь слушать слово из уст Моих, и будешь вразумлять их от Меня.
EZEK|3|18|Когда Я скажу беззаконнику: "смертью умрешь!", а ты не будешь вразумлять его и говорить, чтобы остеречь беззаконника от беззаконного пути его, чтобы он жив был, то беззаконник тот умрет в беззаконии своем, и Я взыщу кровь его от рук твоих.
EZEK|3|19|Но если ты вразумлял беззаконника, а он не обратился от беззакония своего и от беззаконного пути своего, то он умрет в беззаконии своем, а ты спас душу твою.
EZEK|3|20|И если праведник отступит от правды своей и поступит беззаконно, когда Я положу пред ним преткновение, и он умрет, то, если ты не вразумлял его, он умрет за грех свой, и не припомнятся ему праведные дела его, какие делал он; и Я взыщу кровь его от рук твоих.
EZEK|3|21|Если же ты будешь вразумлять праведника, чтобы праведник не согрешил, и он не согрешит, то и он жив будет, потому что был вразумлен, и ты спас душу твою.
EZEK|3|22|И была на мне там рука Господа, и Он сказал мне: встань и выйди в поле, и Я буду говорить там с тобою.
EZEK|3|23|И встал я, и вышел в поле; и вот, там стояла слава Господня, как слава, которую видел я при реке Ховаре; и пал я на лице свое.
EZEK|3|24|И вошел в меня дух, и поставил меня на ноги мои, и Он говорил со мною, и сказал мне: иди и запрись в доме твоем.
EZEK|3|25|И ты, сын человеческий, – вот, возложат на тебя узы, и свяжут тебя ими, и не будешь ходить среди них.
EZEK|3|26|И язык твой Я прилеплю к гортани твоей, и ты онемеешь, и не будешь обличителем их, ибо они мятежный дом.
EZEK|3|27|А когда Я буду говорить с тобою, тогда открою уста твои, и ты будешь говорить им: "так говорит Господь Бог!" кто хочет слушать, слушай; а кто не хочет слушать, не слушай: ибо они мятежный дом.
EZEK|4|1|И ты, сын человеческий, возьми себе кирпич и положи его перед собою, и начертай на нем город Иерусалим;
EZEK|4|2|и устрой осаду против него, и сделай укрепление против него, и насыпь вал вокруг него, и расположи стан против него, и расставь кругом против него стенобитные машины;
EZEK|4|3|и возьми себе железную доску, и поставь ее [как бы] железную стену между тобою и городом, и обрати на него лице твое, и он будет в осаде, и ты осаждай его. Это будет знамением дому Израилеву.
EZEK|4|4|Ты же ложись на левый бок твой и положи на него беззаконие дома Израилева: по числу дней, в которые будешь лежать на нем, ты будешь нести беззаконие их.
EZEK|4|5|И Я определил тебе годы беззакония их числом дней: триста девяносто дней ты будешь нести беззаконие дома Израилева.
EZEK|4|6|И когда исполнишь это, то вторично ложись уже на правый бок, и сорок дней неси на себе беззаконие дома Иудина, день за год, день за год Я определил тебе.
EZEK|4|7|И обрати лице твое и обнаженную правую руку твою на осаду Иерусалима, и пророчествуй против него.
EZEK|4|8|Вот, Я возложил на тебя узы, и ты не повернешься с одного бока на другой, доколе не исполнишь дней осады твоей.
EZEK|4|9|Возьми себе пшеницы и ячменя, и бобов, и чечевицы, и пшена, и полбы, и всыпь их в один сосуд, и сделай себе из них хлебы, по числу дней, в которые ты будешь лежать на боку твоем; триста девяносто дней ты будешь есть их.
EZEK|4|10|И пищу твою, которою будешь питаться, ешь весом по двадцати сиклей в день; от времени до времени ешь это.
EZEK|4|11|И воду пей мерою, по шестой части гина пей; от времени до времени пей так.
EZEK|4|12|И ешь, как ячменные лепешки, и пеки их при глазах их на человеческом кале.
EZEK|4|13|И сказал Господь: так сыны Израилевы будут есть нечистый хлеб свой среди тех народов, к которым Я изгоню их.
EZEK|4|14|Тогда сказал я: о, Господи Боже! душа моя никогда не осквернялась, и мертвечины и растерзанного зверем я не ел от юности моей доныне; и никакое нечистое мясо не входило в уста мои.
EZEK|4|15|И сказал Он мне: вот, Я дозволяю тебе, вместо человеческого кала, коровий помет, и на нем приготовляй хлеб твой.
EZEK|4|16|И сказал мне: сын человеческий! вот, Я сокрушу в Иерусалиме опору хлебную, и будут есть хлеб весом и в печали, и воду будут пить мерою и в унынии,
EZEK|4|17|потому что у них будет недостаток в хлебе и воде; и они с ужасом будут смотреть друг на друга, и исчахнут в беззаконии своем.
EZEK|5|1|А ты, сын человеческий, возьми себе острый нож, бритву брадобреев возьми себе, и води ею по голове твоей и по бороде твоей, и возьми себе весы, и раздели волосы на части.
EZEK|5|2|Третью часть сожги огнем посреди города, когда исполнятся дни осады; третью часть возьми и изруби ножом в окрестностях его; и третью часть развей по ветру; а Я обнажу меч вслед за ними.
EZEK|5|3|И возьми из этого небольшое число, и завяжи их у себя в полы.
EZEK|5|4|Но и из этого еще возьми, и брось в огонь, и сожги это в огне. Оттуда выйдет огонь на весь дом Израилев.
EZEK|5|5|Так говорит Господь Бог: это Иерусалим! Я поставил его среди народов, и вокруг него – земли.
EZEK|5|6|А он поступил против постановлений Моих нечестивее язычников, и против уставов Моих – хуже, нежели земли вокруг него; ибо они отвергли постановления Мои и по уставам Моим не поступают.
EZEK|5|7|Посему так говорит Господь Бог: за то, что вы умножили беззакония ваши более, нежели язычники, которые вокруг вас, по уставам Моим не поступаете и постановлений Моих не исполняете, и даже не поступаете и по постановлениям язычников, которые вокруг вас, –
EZEK|5|8|посему так говорит Господь Бог: вот и Я против тебя, Я Сам, и произведу среди тебя суд перед глазами язычников.
EZEK|5|9|И сделаю над тобою то, чего Я никогда не делал и чему подобного впредь не буду делать, за все твои мерзости.
EZEK|5|10|За то отцы будут есть сыновей среди тебя, и сыновья будут есть отцов своих; и произведу над тобою суд, и весь остаток твой развею по всем ветрам.
EZEK|5|11|Посему, – живу Я, говорит Господь Бог, – за то, что ты осквернил святилище Мое всеми мерзостями твоими и всеми гнусностями твоими, Я умалю тебя, и не пожалеет око Мое, и Я не помилую тебя.
EZEK|5|12|Третья часть у тебя умрет от язвы и погибнет от голода среди тебя; третья часть падет от меча в окрестностях твоих; а третью часть развею по всем ветрам, и обнажу меч вслед за ними.
EZEK|5|13|И совершится гнев Мой, и утолю ярость Мою над ними, и удовлетворюсь; и узнают, что Я, Господь, говорил в ревности Моей, когда совершится над ними ярость Моя.
EZEK|5|14|И сделаю тебя пустынею и поруганием среди народов, которые вокруг тебя, перед глазами всякого мимоходящего.
EZEK|5|15|И будешь посмеянием и поруганием, примером и ужасом у народов, которые вокруг тебя, когда Я произведу над тобою суд во гневе и ярости, и в яростных казнях; – Я, Господь, изрек сие; –
EZEK|5|16|и когда пошлю на них лютые стрелы голода, которые будут губить, когда пошлю их на погибель вашу, и усилю голод между вами, и сокрушу хлебную опору у вас,
EZEK|5|17|и пошлю на вас голод и лютых зверей, и обесчадят тебя; и язва и кровь пройдет по тебе, и меч наведу на тебя; Я, Господь, изрек сие.
EZEK|6|1|И было ко мне слово Господне:
EZEK|6|2|сын человеческий! обрати лице твое к горам Израилевым и прореки на них,
EZEK|6|3|и скажи: горы Израилевы! слушайте слово Господа Бога. Так говорит Господь Бог горам и холмам, долинам и лощинам: вот, Я наведу на вас меч, и разрушу высоты ваши;
EZEK|6|4|и жертвенники ваши будут опустошены, столбы ваши в честь солнца будут разбиты, и повергну убитых ваших перед идолами вашими;
EZEK|6|5|и положу трупы сынов Израилевых перед идолами их, и рассыплю кости ваши вокруг жертвенников ваших.
EZEK|6|6|Во всех местах вашего жительства города будут опустошены и высоты разрушены, для того, чтобы опустошены и разрушены были жертвенники ваши, чтобы сокрушены и уничтожены были идолы ваши, и разбиты солнечные столбы ваши, и изгладились произведения ваши.
EZEK|6|7|И будут падать среди вас убитые, и узнаете, что Я Господь.
EZEK|6|8|Но Я сберегу остаток, так что будут у вас среди народов уцелевшие от меча, когда вы будете рассеяны по землям.
EZEK|6|9|И вспомнят о Мне уцелевшие ваши среди народов, куда будут отведены в плен, когда Я приведу в сокрушение блудное сердце их, отпавшее от Меня, и глаза их, блудившие вслед идолов; и они к самим себе почувствуют отвращение за то зло, какое они делали во всех мерзостях своих;
EZEK|6|10|и узнают, что Я Господь; не напрасно говорил Я, что наведу на них такое бедствие.
EZEK|6|11|Так говорит Господь Бог: всплесни руками твоими и топни ногою твоею, и скажи: горе за все гнусные злодеяния дома Израилева! падут они от меча, голода и моровой язвы.
EZEK|6|12|Кто вдали, тот умрет от моровой язвы; а кто близко, тот падет от меча; а оставшийся и уцелевший умрет от голода; так совершу над ними гнев Мой.
EZEK|6|13|И узнаете, что Я Господь, когда пораженные будут [лежать] между идолами своими вокруг жертвенников их, на всяком высоком холме, на всех вершинах гор и под всяким зеленеющим деревом, и под всяким ветвистым дубом, на том месте, где они приносили благовонные курения всем идолам своим.
EZEK|6|14|И простру на них руку Мою, и сделаю землю пустынею и степью, от пустыни Дивлаф, во всех местах жительства их, и узнают, что Я Господь.
EZEK|7|1|И было ко мне слово Господне:
EZEK|7|2|и ты, сын человеческий, [скажи]: так говорит Господь Бог; земле Израилевой конец, – конец пришел на четыре края земли.
EZEK|7|3|Вот конец тебе; и пошлю на тебя гнев Мой, и буду судить тебя по путям твоим, и возложу на тебя все мерзости твои.
EZEK|7|4|И не пощадит тебя око Мое, и не помилую, и воздам тебе по путям твоим, и мерзости твои с тобою будут, и узнаете, что Я Господь.
EZEK|7|5|Так говорит Господь Бог: беда единственная, вот, идет беда.
EZEK|7|6|Конец пришел, пришел конец, встал на тебя; вот дошла,
EZEK|7|7|дошла напасть до тебя, житель земли! приходит время, приближается день смятения, а не веселых восклицаний на горах.
EZEK|7|8|Вот, скоро изолью на тебя ярость Мою и совершу над тобою гнев Мой, и буду судить тебя по путям твоим, и возложу на тебя все мерзости твои.
EZEK|7|9|И не пощадит тебя око Мое, и не помилую. По путям твоим воздам тебе, и мерзости твои с тобою будут; и узнаете, что Я Господь каратель.
EZEK|7|10|Вот день! вот пришла, наступила напасть! жезл вырос, гордость разрослась.
EZEK|7|11|Восстает сила на жезл нечестия; ничего [не останется] от них, и от богатства их, и от шума их, и от пышности их.
EZEK|7|12|Пришло время, наступил день; купивший не радуйся, и продавший не плачь; ибо гнев над всем множеством их.
EZEK|7|13|Ибо продавший не возвратится к проданному, хотя бы и остались они в живых; ибо пророческое видение о всем множестве их не отменится, и никто своим беззаконием не укрепит своей жизни.
EZEK|7|14|Затрубят в трубу, и все готовится, но никто не идет на войну: ибо гнев Мой над всем множеством их.
EZEK|7|15|Вне дома меч, а в доме мор и голод. Кто в поле, тот умрет от меча; а кто в городе, того пожрут голод и моровая язва.
EZEK|7|16|А уцелевшие из них убегут и будут на горах, как голуби долин; все они будут стонать, каждый за свое беззаконие.
EZEK|7|17|У всех руки опустятся, и у всех колени задрожат, [как] вода.
EZEK|7|18|Тогда они препояшутся вретищем, и обоймет их трепет; и у всех на лицах будет стыд, и у всех на головах плешь.
EZEK|7|19|Серебро свое они выбросят на улицы, и золото у них будет в пренебрежении. Серебро их и золото их не сильно будет спасти их в день ярости Господа. Они не насытят ими душ своих и не наполнят утроб своих; ибо оно было поводом к беззаконию их.
EZEK|7|20|И в красных нарядах своих они превращали его в гордость, и делали из него изображения гнусных своих истуканов; за то и сделаю его нечистым для них;
EZEK|7|21|и отдам его в руки чужим в добычу и беззаконникам земли на расхищение, и они осквернят его.
EZEK|7|22|И отвращу от них лице Мое, и осквернят сокровенное Мое; и придут туда грабители, и осквернят его.
EZEK|7|23|Сделай цепь, ибо земля эта наполнена кровавыми злодеяниями, и город полон насилий.
EZEK|7|24|Я приведу злейших из народов, и завладеют домами их. И положу конец надменности сильных, и будут осквернены святыни их.
EZEK|7|25|Идет пагуба; будут искать мира, и не найдут.
EZEK|7|26|Беда пойдет за бедою и весть за вестью; и будут просить у пророка видения, и не станет учения у священника и совета у старцев.
EZEK|7|27|Царь будет сетовать, и князь облечется в ужас, и у народа земли будут дрожать руки. Поступлю с ними по путям их, и по судам их буду судить их; и узнают, что Я Господь.
EZEK|8|1|И было в шестом году, в шестом [месяце], в пятый день месяца, сидел я в доме моем, и старейшины Иудейские сидели перед лицем моим, и низошла на меня там рука Господа Бога.
EZEK|8|2|И увидел я: и вот подобие [мужа], как бы огненное, и от чресл его и ниже – огонь, и от чресл его и выше – как бы сияние, как бы свет пламени.
EZEK|8|3|И простер Он как бы руку, и взял меня за волоса головы моей, и поднял меня дух между землею и небом, и принес меня в видениях Божиих в Иерусалим ко входу внутренних ворот, обращенных к северу, где поставлен был идол ревности, возбуждающий ревнование.
EZEK|8|4|И вот, там была слава Бога Израилева, подобная той, какую я видел на поле.
EZEK|8|5|И сказал мне: сын человеческий! подними глаза твои к северу. И я поднял глаза мои к северу, и вот, с северной стороны у ворот жертвенника – тот идол ревности при входе.
EZEK|8|6|И сказал Он мне: сын человеческий! видишь ли ты, что они делают? великие мерзости, какие делает дом Израилев здесь, чтобы Я удалился от святилища Моего? но обратись, и ты увидишь еще большие мерзости.
EZEK|8|7|И привел меня ко входу во двор, и я взглянул, и вот в стене скважина.
EZEK|8|8|И сказал мне: сын человеческий! прокопай стену; и я прокопал стену, и вот какая–то дверь.
EZEK|8|9|И сказал мне: войди и посмотри на отвратительные мерзости, какие они делают здесь.
EZEK|8|10|И вошел я, и вижу, и вот всякие изображения пресмыкающихся и нечистых животных и всякие идолы дома Израилева, написанные по стенам кругом.
EZEK|8|11|И семьдесят мужей из старейшин дома Израилева стоят перед ними, и Иезания, сын Сафанов, среди них; и у каждого в руке свое кадило, и густое облако курений возносится кверху.
EZEK|8|12|И сказал мне: видишь ли, сын человеческий, что делают старейшины дома Израилева в темноте, каждый в расписанной своей комнате? ибо говорят: "не видит нас Господь, оставил Господь землю сию".
EZEK|8|13|И сказал мне: обратись, и увидишь еще большие мерзости, какие они делают.
EZEK|8|14|И привел меня ко входу в ворота дома Господня, которые к северу, и вот, там сидят женщины, плачущие по Фаммузе,
EZEK|8|15|и сказал мне: видишь ли, сын человеческий? обратись, и еще увидишь большие мерзости.
EZEK|8|16|И ввел меня во внутренний двор дома Господня, и вот у дверей храма Господня, между притвором и жертвенником, около двадцати пяти мужей [стоят] спинами своими ко храму Господню, а лицами своими на восток, и кланяются на восток солнцу.
EZEK|8|17|И сказал мне: видишь ли, сын человеческий? мало ли дому Иудину, чтобы делать такие мерзости, какие они делают здесь? но они еще землю наполнили нечестием, и сугубо прогневляют Меня; и вот, они ветви подносят к носам своим.
EZEK|8|18|За то и Я стану действовать с яростью; не пожалеет око Мое, и не помилую; и хотя бы они взывали в уши Мои громким голосом, не услышу их.
EZEK|9|1|И возгласил в уши мои великим гласом, говоря: пусть приблизятся каратели города, каждый со своим губительным орудием в руке своей.
EZEK|9|2|И вот, шесть человек идут от верхних ворот, обращенных к северу, и у каждого в руке губительное орудие его, и между ними один, одетый в льняную одежду, у которого при поясе его прибор писца. И пришли и стали подле медного жертвенника.
EZEK|9|3|И слава Бога Израилева сошла с Херувима, на котором была, к порогу дома. И призвал Он человека, одетого в льняную одежду, у которого при поясе прибор писца.
EZEK|9|4|И сказал ему Господь: пройди посреди города, посреди Иерусалима, и на челах людей скорбящих, воздыхающих о всех мерзостях, совершающихся среди него, сделай знак.
EZEK|9|5|А тем сказал в слух мой: идите за ним по городу и поражайте; пусть не жалеет око ваше, и не щадите;
EZEK|9|6|старика, юношу и девицу, и младенца и жен бейте до смерти, но не троньте ни одного человека, на котором знак, и начните от святилища Моего. И начали они с тех старейшин, которые были перед домом.
EZEK|9|7|И сказал им: оскверните дом, и наполните дворы убитыми, и выйдите. И вышли, и стали убивать в городе.
EZEK|9|8|И когда они их убили, а я остался, тогда я пал на лице свое и возопил, и сказал: о, Господи Боже! неужели Ты погубишь весь остаток Израиля, изливая гнев Твой на Иерусалим?
EZEK|9|9|И сказал Он мне: нечестие дома Израилева и Иудина велико, весьма велико; и земля сия полна крови, и город исполнен неправды; ибо они говорят: "оставил Господь землю сию, и не видит Господь".
EZEK|9|10|За то и Мое око не пощадит, и не помилую; обращу поведение их на их голову.
EZEK|9|11|И вот человек, одетый в льняную одежду, у которого при поясе прибор писца, дал ответ и сказал: я сделал, как Ты повелел мне.
EZEK|10|1|И видел я, и вот на своде, который над главами Херувимов, как бы камень сапфир, как бы нечто, похожее на престол, видимо было над ними.
EZEK|10|2|И говорил Он человеку, одетому в льняную одежду, и сказал: войди между колесами под Херувимов и возьми полные пригоршни горящих угольев между Херувимами, и брось на город; и он вошел в моих глазах.
EZEK|10|3|Херувимы же стояли по правую сторону дома, когда вошел тот человек, и облако наполняло внутренний двор.
EZEK|10|4|И поднялась слава Господня с Херувима к порогу дома, и дом наполнился облаком, и двор наполнился сиянием славы Господа.
EZEK|10|5|И шум от крыльев Херувимов слышен был даже на внешнем дворе, как бы глас Бога Всемогущего, когда Он говорит.
EZEK|10|6|И когда Он дал повеление человеку, одетому в льняную одежду, сказав: "возьми огня между колесами, между Херувимами", и когда он вошел и стал у колеса, –
EZEK|10|7|тогда из среды Херувимов один Херувим простер руку свою к огню, который между Херувимами, и взял и дал в пригоршни одетому в льняную одежду. Он взял и вышел.
EZEK|10|8|И видно было у Херувимов подобие рук человеческих под крыльями их.
EZEK|10|9|И видел я: и вот четыре колеса подле Херувимов, по одному колесу подле каждого Херувима, и колеса по виду как бы из камня топаза.
EZEK|10|10|И по виду все четыре сходны, как будто бы колесо находилось в колесе.
EZEK|10|11|Когда шли они, то шли на четыре свои стороны; во время шествия своего не оборачивались, но к тому месту, куда обращена была голова, и они туда шли; во время шествия своего не оборачивались.
EZEK|10|12|И все тело их, и спина их, и руки их, и крылья их, и колеса кругом были полны очей, все четыре колеса их.
EZEK|10|13|К колесам сим, как я слышал, сказано было: "галгал".
EZEK|10|14|И у каждого [из] животных четыре лица: первое лице – лице херувимово, второе лице – лице человеческое, третье лице львиное и четвертое лице орлиное.
EZEK|10|15|Херувимы поднялись. Это были те же животные, которых видел я при реке Ховаре.
EZEK|10|16|И когда шли Херувимы, тогда шли подле них и колеса; и когда Херувимы поднимали крылья свои, чтобы подняться от земли, и колеса не отделялись, но были при них.
EZEK|10|17|Когда те стояли, стояли и они; когда те поднимались, поднимались и они; ибо в них [был] дух животных.
EZEK|10|18|И отошла слава Господня от порога дома и стала над Херувимами.
EZEK|10|19|И подняли Херувимы крылья свои, и поднялись в глазах моих от земли; когда они уходили, то и колеса подле них; и стали у входа в восточные врата Дома Господня, и слава Бога Израилева вверху над ними.
EZEK|10|20|Это были те же животные, которых видел я в подножии Бога Израилева при реке Ховаре. И я узнал, что это Херувимы.
EZEK|10|21|У каждого по четыре лица, и у каждого по четыре крыла, и под крыльями их подобие рук человеческих.
EZEK|10|22|А подобие лиц их то же, какие лица видел я при реке Ховаре, – и вид их, и сами они. Каждый шел прямо в ту сторону, которая была перед лицем его.
EZEK|11|1|И поднял меня дух, и привел меня к восточным воротам дома Господня, которые обращены к востоку. И вот, у входа в ворота двадцать пять человек; и между ними я видел Иазанию, сына Азурова, и Фалтию, сына Ванеева, князей народа.
EZEK|11|2|И Он сказал мне: сын человеческий! вот люди, у которых на уме беззаконие и которые дают худой совет в городе сем,
EZEK|11|3|говоря: "еще не близко; будем строить домы; он котел, а мы мясо".
EZEK|11|4|Посему изреки на них пророчество, пророчествуй, сын человеческий.
EZEK|11|5|И нисшел на меня Дух Господень и сказал мне: скажи, так говорит Господь: что говорите вы, дом Израилев, и что на ум вам приходит, это Я знаю.
EZEK|11|6|Много убитых ваших вы положили в сем городе и улицы его наполнили трупами.
EZEK|11|7|Посему так говорит Господь Бог: убитые ваши, которых вы положили среди него, суть мясо, а он – котел; но вас Я выведу из него.
EZEK|11|8|Вы боитесь меча, и Я наведу на вас меч, говорит Господь Бог.
EZEK|11|9|И выведу вас из него, и отдам вас в руку чужих, и произведу над вами суд.
EZEK|11|10|От меча падете; на пределах Израилевых будут судить вас, и узнаете, что Я Господь.
EZEK|11|11|Он не будет для вас котлом, и вы не будете мясом в нем; на пределах Израилевых буду судить вас.
EZEK|11|12|И узнаете, что Я Господь; ибо по заповедям Моим вы не ходили и уставов Моих не выполняли, а поступали по уставам народов, окружающих вас.
EZEK|11|13|И было, когда я пророчествовал, Фалтия, сын Ванеев, умер. И пал я на лице, и возопил громким голосом, и сказал: о, Господи Боже! неужели Ты хочешь до конца истребить остаток Израиля?
EZEK|11|14|И было ко мне слово Господне:
EZEK|11|15|сын человеческий! твоим братьям, твоим братьям, твоим единокровным и всему дому Израилеву, всем им говорят живущие в Иерусалиме: "живите вдали от Господа; нам во владение отдана эта земля".
EZEK|11|16|На это скажи: так говорит Господь Бог: хотя Я и удалил их к народам и хотя рассеял их по землям, но Я буду для них некоторым святилищем в тех землях, куда пошли они.
EZEK|11|17|Затем скажи: так говорит Господь Бог: Я соберу вас из народов, и возвращу вас из земель, в которые вы рассеяны; и дам вам землю Израилеву.
EZEK|11|18|И придут туда, и извергнут из нее все гнусности ее и все мерзости ее.
EZEK|11|19|И дам им сердце единое, и дух новый вложу в них, и возьму из плоти их сердце каменное, и дам им сердце плотяное,
EZEK|11|20|чтобы они ходили по заповедям Моим, и соблюдали уставы Мои, и выполняли их; и будут Моим народом, а Я буду их Богом.
EZEK|11|21|А чье сердце увлечется вслед гнусностей их и мерзостей их, поведение тех обращу на их голову, говорит Господь Бог.
EZEK|11|22|Тогда Херувимы подняли крылья свои, и колеса подле них; и слава Бога Израилева вверху над ними.
EZEK|11|23|И поднялась слава Господа из среды города и остановилась над горою, которая на восток от города.
EZEK|11|24|И дух поднял меня и перенес меня в Халдею, к переселенцам, в видении, Духом Божиим. И отошло от меня видение, которое я видел.
EZEK|11|25|И я пересказал переселенцам все слова Господа, которые Он открыл мне.
EZEK|12|1|И было ко мне слово Господне:
EZEK|12|2|сын человеческий! ты живешь среди дома мятежного; у них есть глаза, чтобы видеть, а не видят; у них есть уши, чтобы слышать, а не слышат; потому что они – мятежный дом.
EZEK|12|3|Ты же, сын человеческий, изготовь себе нужное для переселения, и среди дня переселяйся перед глазами их, и переселяйся с места твоего в другое место перед глазами их; может быть, они уразумеют, хотя они – дом мятежный;
EZEK|12|4|и вещи твои вынеси, как вещи нужные при переселении, днем, перед глазами их, и сам выйди вечером перед глазами их, как выходят для переселения.
EZEK|12|5|Перед глазами их проломай себе отверстие в стене, и вынеси через него.
EZEK|12|6|Перед глазами их возьми ношу на плечо, впотьмах вынеси ее, лице твое закрой, чтобы не видеть земли; ибо Я поставил тебя знамением дому Израилеву.
EZEK|12|7|И сделал я, как повелено было мне; вещи мои, как вещи нужные при переселении, вынес днем, а вечером проломал себе рукою отверстие в стене, впотьмах вынес ношу и поднял на плечо перед глазами их.
EZEK|12|8|И было ко мне слово Господне поутру:
EZEK|12|9|сын человеческий! не говорил ли тебе дом Израилев, дом мятежный: "что ты делаешь?"
EZEK|12|10|Скажи им: так говорит Господь Бог: это – предвещание для начальствующего в Иерусалиме и для всего дома Израилева, который находится там.
EZEK|12|11|Скажи: я знамение для вас; что делаю я, то будет с ними, – в переселение, в плен пойдут они.
EZEK|12|12|И начальствующий, который среди них, впотьмах поднимет [ношу] на плечо и выйдет. Стену проломают, чтобы отправить [его] через нее; он закроет лице свое, так что не увидит глазами земли сей.
EZEK|12|13|И раскину на него сеть Мою, и будет пойман в тенета Мои, и отведу его в Вавилон, в землю Халдейскую, но он не увидит ее, и там умрет.
EZEK|12|14|А всех, которые вокруг него, споборников его и все войско его развею по всем ветрам, и обнажу вслед их меч.
EZEK|12|15|И узнают, что Я Господь, когда рассею их по народам и развею их по землям.
EZEK|12|16|Но небольшое число их Я сохраню от меча, голода и язвы, чтобы они рассказали у народов, к которым пойдут, о всех своих мерзостях; и узнают, что Я Господь.
EZEK|12|17|И было ко мне слово Господне:
EZEK|12|18|сын человеческий! хлеб твой ешь с трепетом, и воду твою пей с дрожанием и печалью.
EZEK|12|19|И скажи народу земли: так говорит Господь Бог о жителях Иерусалима, о земле Израилевой: они хлеб свой будут есть с печалью и воду свою будут пить в унынии, потому что земля его будет лишена всего изобилия своего за неправды всех живущих на ней.
EZEK|12|20|И будут разорены населенные города, и земля сделается пустою, и узнаете, что Я Господь.
EZEK|12|21|И было ко мне слово Господне:
EZEK|12|22|сын человеческий! что за поговорка у вас, в земле Израилевой: "много дней пройдет, и всякое пророческое видение исчезнет"?
EZEK|12|23|Посему скажи им: так говорит Господь Бог: уничтожу эту поговорку, и не будут уже употреблять такой поговорки у Израиля; но скажи им: близки дни и исполнение всякого видения пророческого.
EZEK|12|24|Ибо уже не останется втуне никакое видение пророческое, и ни одно предвещание не будет ложным в доме Израилевом.
EZEK|12|25|Ибо Я Господь, Я говорю; и слово, которое Я говорю, исполнится, и не будет отложено; в ваши дни, мятежный дом, Я изрек слово, и исполню его, говорит Господь Бог.
EZEK|12|26|И было ко мне слово Господне:
EZEK|12|27|сын человеческий! вот, дом Израилев говорит: "пророческое видение, которое видел он, [сбудется] после многих дней, и он пророчествует об отдаленных временах".
EZEK|12|28|Посему скажи им: так говорит Господь Бог: ни одно из слов Моих уже не будет отсрочено, но слово, которое Я скажу, сбудется, говорит Господь Бог.
EZEK|13|1|И было ко мне слово Господне:
EZEK|13|2|сын человеческий! изреки пророчество на пророков Израилевых пророчествующих, и скажи пророкам от собственного сердца: слушайте слово Господне!
EZEK|13|3|Так говорит Господь Бог: горе безумным пророкам, которые водятся своим духом и ничего не видели!
EZEK|13|4|Пророки твои, Израиль, как лисицы в развалинах.
EZEK|13|5|В проломы вы не входите и не ограждаете стеною дома Израилева, чтобы твердо стоять в сражении в день Господа.
EZEK|13|6|Они видят пустое и предвещают ложь, говоря: "Господь сказал"; а Господь не посылал их; и обнадеживают, что слово сбудется.
EZEK|13|7|Не пустое ли видение видели вы? и не лживое ли предвещание изрекаете, говоря: "Господь сказал", а Я не говорил?
EZEK|13|8|Посему так говорит Господь Бог: так как вы говорите пустое и видите в видениях ложь, за то вот Я – на вас, говорит Господь Бог.
EZEK|13|9|И будет рука Моя против этих пророков, видящих пустое и предвещающих ложь; в совете народа Моего они не будут, и в список дома Израилева не впишутся, и в землю Израилеву не войдут; и узнаете, что Я Господь Бог.
EZEK|13|10|За то, что они вводят народ Мой в заблуждение, говоря: "мир", тогда как нет мира; и когда он строит стену, они обмазывают ее грязью,
EZEK|13|11|скажи обмазывающим стену грязью, что она упадет. Пойдет проливной дождь, и вы, каменные градины, падете, и бурный ветер разорвет ее.
EZEK|13|12|И вот, падет стена; тогда не скажут ли вам: "где та обмазка, которою вы обмазывали?"
EZEK|13|13|Посему так говорит Господь Бог: Я пущу бурный ветер во гневе Моем, и пойдет проливной дождь в ярости Моей, и камни града в негодовании Моем, для истребления.
EZEK|13|14|И разрушу стену, которую вы обмазывали грязью, и повергну ее на землю, и откроется основание ее, и падет, и вы вместе с нею погибнете; и узнаете, что Я Господь.
EZEK|13|15|И истощу ярость Мою на стене и на обмазывающих ее грязью, и скажу вам: нет стены, и нет обмазывавших ее,
EZEK|13|16|пророков Израилевых, которые пророчествовали Иерусалиму и возвещали ему видения мира, тогда как нет мира, говорит Господь Бог.
EZEK|13|17|Ты же, сын человеческий, обрати лице твое к дщерям народа твоего, пророчествующим от собственного своего сердца, и изреки на них пророчество,
EZEK|13|18|и скажи: так говорит Господь Бог: горе сшивающим чародейные мешочки под мышки и делающим покрывала для головы всякого роста, чтобы уловлять души! Неужели, уловляя души народа Моего, вы спасете ваши души?
EZEK|13|19|И бесславите Меня пред народом Моим за горсти ячменя и за куски хлеба, умерщвляя души, которые не должны умереть, и оставляя жизнь душам, которые не должны жить, обманывая народ, который слушает ложь.
EZEK|13|20|Посему так говорит Господь Бог: вот, Я – на ваши чародейные мешочки, которыми вы там уловляете души, чтобы они прилетали, и вырву их из–под мышц ваших, и пущу на свободу души, которые вы уловляете, чтобы прилетали к вам.
EZEK|13|21|И раздеру покрывала ваши, и избавлю народ Мой от рук ваших, и не будут уже в ваших руках добычею, и узнаете, что Я Господь.
EZEK|13|22|За то, что вы ложью опечаливаете сердце праведника, которое Я не хотел опечаливать, и поддерживаете руки беззаконника, чтобы он не обратился от порочного пути своего и не сохранил жизни своей, –
EZEK|13|23|за это уже не будете иметь пустых видений и впредь не будете предугадывать; и Я избавлю народ Мой от рук ваших, и узнаете, что Я Господь.
EZEK|14|1|И пришли ко мне несколько человек из старейшин Израилевых и сели перед лицем моим.
EZEK|14|2|И было ко мне слово Господне:
EZEK|14|3|сын человеческий! Сии люди допустили идолов своих в сердце свое и поставили соблазн нечестия своего перед лицем своим: могу ли Я отвечать им?
EZEK|14|4|Посему говори с ними и скажи им: так говорит Господь Бог: если кто из дома Израилева допустит идолов своих в сердце свое и поставит соблазн нечестия своего перед лицем своим, и придет к пророку, – то Я, Господь, могу ли, при множестве идолов его, дать ему ответ?
EZEK|14|5|Пусть дом Израилев поймет в сердце своем, что все они через своих идолов сделались чужими для Меня.
EZEK|14|6|Посему скажи дому Израилеву: так говорит Господь Бог: обратитесь и отвратитесь от идолов ваших, и от всех мерзостей ваших отвратите лице ваше.
EZEK|14|7|Ибо если кто из дома Израилева и из пришельцев, которые живут у Израиля, отложится от Меня и допустит идолов своих в сердце свое, и поставит соблазн нечестия своего перед лицем своим, и придет к пророку вопросить Меня через него, – то Я, Господь, дам ли ему ответ от Себя?
EZEK|14|8|Я обращу лице Мое против того человека и сокрушу его в знамение и притчу, и истреблю его из народа Моего, и узнаете, что Я Господь.
EZEK|14|9|А если пророк допустит обольстить себя и скажет слово так, как бы Я, Господь, научил этого пророка, то Я простру на него руку Мою и истреблю его из народа Моего, Израиля.
EZEK|14|10|И понесут вину беззакония своего: какова вина вопрошающего, такова будет вина и пророка,
EZEK|14|11|чтобы впредь дом Израилев не уклонялся от Меня и чтобы более не оскверняли себя всякими беззакониями своими, но чтобы были Моим народом, и Я был их Богом, говорит Господь Бог.
EZEK|14|12|И было ко мне слово Господне:
EZEK|14|13|сын человеческий! если бы какая земля согрешила предо Мною, вероломно отступив от Меня, и Я простер на нее руку Мою, и истребил в ней хлебную опору, и послал на нее голод, и стал губить на ней людей и скот;
EZEK|14|14|и если бы нашлись в ней сии три мужа: Ной, Даниил и Иов, – то они праведностью своею спасли бы только свои души, говорит Господь Бог.
EZEK|14|15|Или, если бы Я послал на эту землю лютых зверей, которые осиротили бы ее, и она по причине зверей сделалась пустою и непроходимою:
EZEK|14|16|то сии три мужа среди нее, – живу Я, говорит Господь Бог, – не спасли бы ни сыновей, ни дочерей, а они, только они спаслись бы, земля же сделалась бы пустынею.
EZEK|14|17|Или, если бы Я навел на ту землю меч и сказал: "меч, пройди по земле!", и стал истреблять на ней людей и скот,
EZEK|14|18|то сии три мужа среди нее, – живу Я, говорит Господь Бог, – не спасли бы ни сыновей, ни дочерей, а они только спаслись бы.
EZEK|14|19|Или, если бы Я послал на ту землю моровую язву и излил на нее ярость Мою в кровопролитии, чтобы истребить на ней людей и скот:
EZEK|14|20|то Ной, Даниил и Иов среди нее, – живу Я, говорит Господь Бог, – не спасли бы ни сыновей, ни дочерей; праведностью своею они спасли бы только свои души.
EZEK|14|21|Ибо так говорит Господь Бог: если и четыре тяжкие казни Мои: меч, и голод, и лютых зверей, и моровую язву пошлю на Иерусалим, чтобы истребить в нем людей и скот,
EZEK|14|22|и тогда останется в нем остаток, сыновья и дочери, которые будут выведены оттуда; вот, они выйдут к вам, и вы увидите поведение их и дела их, и утешитесь о том бедствии, которое Я навел на Иерусалим, о всем, что Я навел на него.
EZEK|14|23|Они утешат вас, когда вы увидите поведение их и дела их; и узнаете, что Я не напрасно сделал все то, что сделал в нем, говорит Господь Бог.
EZEK|15|1|И было ко мне слово Господне:
EZEK|15|2|сын человеческий! какое преимущество имеет дерево виноградной лозы перед всяким другим деревом и ветви виноградной лозы – между деревами в лесу?
EZEK|15|3|Берут ли от него кусок на какое–либо изделие? Берут ли от него хотя на гвоздь, чтобы вешать на нем какую–либо вещь?
EZEK|15|4|Вот, оно отдается огню на съедение; оба конца его огонь поел, и обгорела середина его: годится ли оно на какое–нибудь изделие?
EZEK|15|5|И тогда, как оно было цело, не годилось ни на какое изделие; тем паче, когда огонь поел его, и оно обгорело, годится ли оно на какое–нибудь изделие?
EZEK|15|6|Посему так говорит Господь Бог: как дерево виноградной лозы между деревами лесными Я отдал огню на съедение, так отдам ему и жителей Иерусалима.
EZEK|15|7|И обращу лице Мое против них; из одного огня выйдут, и другой огонь пожрет их, – и узнаете, что Я Господь, когда обращу против них лице Мое.
EZEK|15|8|И сделаю эту землю пустынею за то, что они вероломно поступали, говорит Господь Бог.
EZEK|16|1|И было ко мне слово Господне:
EZEK|16|2|сын человеческий! выскажи Иерусалиму мерзости его
EZEK|16|3|и скажи: так говорит Господь Бог [дщери] Иерусалима: твой корень и твоя родина в земле Ханаанской; отец твой Аморрей, и мать твоя Хеттеянка;
EZEK|16|4|при рождении твоем, в день, когда ты родилась, пупа твоего не отрезали, и водою ты не была омыта для очищения, и солью не была осолена, и пеленами не повита.
EZEK|16|5|Ничей глаз не сжалился над тобою, чтобы из милости к тебе сделать тебе что–нибудь из этого; но ты выброшена была на поле, по презрению к жизни твоей, в день рождения твоего.
EZEK|16|6|И проходил Я мимо тебя, и увидел тебя, брошенную на попрание в кровях твоих, и сказал тебе: "в кровях твоих живи!" Так, Я сказал тебе: "в кровях твоих живи!"
EZEK|16|7|Умножил тебя как полевые растения; ты выросла и стала большая, и достигла превосходной красоты: поднялись груди, и волоса у тебя выросли; но ты была нага и непокрыта.
EZEK|16|8|И проходил Я мимо тебя, и увидел тебя, и вот, это было время твое, время любви; и простер Я воскрилия [риз] Моих на тебя, и покрыл наготу твою; и поклялся тебе и вступил в союз с тобою, говорит Господь Бог, – и ты стала Моею.
EZEK|16|9|Омыл Я тебя водою и смыл с тебя кровь твою и помазал тебя елеем.
EZEK|16|10|И надел на тебя узорчатое платье, и обул тебя в сафьяные сандалии, и опоясал тебя виссоном, и покрыл тебя шелковым покрывалом.
EZEK|16|11|И нарядил тебя в наряды, и положил на руки твои запястья и на шею твою ожерелье.
EZEK|16|12|И дал тебе кольцо на твой нос и серьги к ушам твоим и на голову твою прекрасный венец.
EZEK|16|13|Так украшалась ты золотом и серебром, и одежда твоя [была] виссон и шелк и узорчатые ткани; питалась ты хлебом из лучшей пшеничной муки, медом и елеем, и была чрезвычайно красива, и достигла царственного величия.
EZEK|16|14|И пронеслась по народам слава твоя ради красоты твоей, потому что она была вполне совершенна при том великолепном наряде, который Я возложил на тебя, говорит Господь Бог.
EZEK|16|15|Но ты понадеялась на красоту твою, и, пользуясь славою твоею, стала блудить и расточала блудодейство твое на всякого мимоходящего, отдаваясь ему.
EZEK|16|16|И взяла из одежд твоих, и сделала себе разноцветные высоты, и блудодействовала на них, как никогда не случится и не будет.
EZEK|16|17|И взяла нарядные твои вещи из Моего золота и из Моего серебра, которые Я дал тебе, и сделала себе мужские изображения, и блудодействовала с ними.
EZEK|16|18|И взяла узорчатые платья твои, и одела их ими, и ставила перед ними елей Мой и фимиам Мой,
EZEK|16|19|и хлеб Мой, который Я давал тебе, пшеничную муку, и елей, и мед, которыми Я питал тебя, ты поставляла перед ними в приятное благовоние; и это было, говорит Господь Бог.
EZEK|16|20|И взяла сыновей твоих и дочерей твоих, которых ты родила Мне, и приносила в жертву на снедение им. Мало ли тебе было блудодействовать?
EZEK|16|21|Но ты и сыновей Моих заколала и отдавала им, проводя их [через] [огонь].
EZEK|16|22|И при всех твоих мерзостях и блудодеяниях твоих ты не вспомнила о днях юности твоей, когда ты была нага и непокрыта и брошена в крови твоей на попрание.
EZEK|16|23|И после всех злодеяний твоих, – горе, горе тебе! говорит Господь Бог, –
EZEK|16|24|ты построила себе блудилища и наделала себе возвышений на всякой площади;
EZEK|16|25|при начале всякой дороги устроила себе возвышения, позорила красоту твою и раскидывала ноги твои для всякого мимоходящего, и умножила блудодеяния твои.
EZEK|16|26|Блудила с сыновьями Египта, соседями твоими, людьми великорослыми, и умножала блудодеяния твои, прогневляя Меня.
EZEK|16|27|И вот, Я простер на тебя руку Мою, и уменьшил назначенное тебе, и отдал тебя на произвол ненавидящим тебя дочерям Филистимским, которые устыдились срамного поведения твоего.
EZEK|16|28|И блудила ты с сынами Ассура и не насытилась; блудила с ними, но тем не удовольствовалась;
EZEK|16|29|и умножила блудодеяния твои в земле Ханаанской до Халдеи, но и тем не удовольствовалась.
EZEK|16|30|Как истомлено должно быть сердце твое, говорит Господь Бог, когда ты все это делала, как необузданная блудница!
EZEK|16|31|Когда ты строила себе блудилища при начале всякой дороги и делала себе возвышения на всякой площади, ты была не как блудница, потому что отвергала подарки,
EZEK|16|32|но как прелюбодейная жена, принимающая вместо своего мужа чужих.
EZEK|16|33|Всем блудницам дают подарки, а ты сама давала подарки всем любовникам твоим и подкупала их, чтобы они со всех сторон приходили к тебе блудить с тобою.
EZEK|16|34|У тебя в блудодеяниях твоих было противное тому, что бывает с женщинами: не за тобою гонялись, но ты давала подарки, а тебе не давали подарков; и потому ты поступала в противность другим.
EZEK|16|35|Посему выслушай, блудница, слово Господне!
EZEK|16|36|Так говорит Господь Бог: за то, что ты так сыпала деньги твои, и в блудодеяниях твоих раскрываема была нагота твоя перед любовниками твоими и перед всеми мерзкими идолами твоими, и за кровь сыновей твоих, которых ты отдавала им, –
EZEK|16|37|за то вот, Я соберу всех любовников твоих, которыми ты услаждалась и которых ты любила, со всеми теми, которых ненавидела, и соберу их отовсюду против тебя, и раскрою перед ними наготу твою, и увидят весь срам твой.
EZEK|16|38|Я буду судить тебя судом прелюбодейц и проливающих кровь, – и предам тебя кровавой ярости и ревности;
EZEK|16|39|предам тебя в руки их и они разорят блудилища твои, и раскидают возвышения твои, и сорвут с тебя одежды твои, и возьмут наряды твои, и оставят тебя нагою и непокрытою.
EZEK|16|40|И созовут на тебя собрание, и побьют тебя камнями, и разрубят тебя мечами своими.
EZEK|16|41|Сожгут домы твои огнем и совершат над тобою суд перед глазами многих жен; и положу конец блуду твоему, и не будешь уже давать подарков.
EZEK|16|42|И утолю над тобою гнев Мой, и отступит от тебя негодование Мое, и успокоюсь, и уже не буду гневаться.
EZEK|16|43|За то, что ты не вспомнила о днях юности твоей и всем этим раздражала Меня, вот, и Я поведение твое обращу на [твою] голову, говорит Господь Бог, чтобы ты не предавалась более разврату после всех твоих мерзостей.
EZEK|16|44|Вот, всякий, кто говорит притчами, может сказать о тебе: "какова мать, такова и дочь".
EZEK|16|45|Ты дочь в мать твою, которая бросила мужа своего и детей своих, – и ты сестра в сестер твоих, которые бросили мужей своих и детей своих. Мать ваша Хеттеянка, и отец ваш Аморрей.
EZEK|16|46|Большая же сестра твоя – Самария, с дочерями своими живущая влево от тебя; а меньшая сестра твоя, живущая от тебя вправо, есть Содома с дочерями ее.
EZEK|16|47|Но ты и не их путями ходила и не по их мерзостям поступала; этого было мало: ты поступала развратнее их на всех путях твоих.
EZEK|16|48|Живу Я, говорит Господь Бог; Содома, сестра твоя, не делала того сама и ее дочери, что делала ты и дочери твои.
EZEK|16|49|Вот в чем было беззаконие Содомы, сестры твоей и дочерей ее: в гордости, пресыщении и праздности, и она руки бедного и нищего не поддерживала.
EZEK|16|50|И возгордились они, и делали мерзости пред лицем Моим, и, увидев это, Я отверг их.
EZEK|16|51|И Самария половины грехов твоих не нагрешила; ты превзошла их мерзостями твоими, и через твои мерзости, какие делала ты, сестры твои оказались правее тебя.
EZEK|16|52|Неси же посрамление твое и ты, которая осуждала сестер твоих; по грехам твоим, какими ты опозорила себя более их, они правее тебя. Красней же от стыда и ты, и неси посрамление твое, так оправдав сестер твоих.
EZEK|16|53|Но Я возвращу плен их, плен Содомы и дочерей ее, плен Самарии и дочерей ее, и между ними плен плененных твоих,
EZEK|16|54|дабы ты несла посрамление твое и стыдилась всего того, что делала, служа для них утешением.
EZEK|16|55|И сестры твои, Содома и дочери ее, возвратятся в прежнее состояние свое; и Самария и дочери ее возвратятся в прежнее состояние свое, и ты и дочери твои возвратитесь в прежнее состояние ваше.
EZEK|16|56|О сестре твоей Содоме и помина не было в устах твоих во дни гордыни твоей,
EZEK|16|57|доколе еще не открыто было нечестие твое, как во время посрамления от дочерей Сирии и всех окружавших ее, от дочерей Филистимы, смотревших на тебя с презрением со всех сторон.
EZEK|16|58|За разврат твой и за мерзости твои терпишь ты, говорит Господь.
EZEK|16|59|Ибо так говорит Господь Бог: Я поступлю с тобою, как поступила ты, презрев клятву нарушением союза.
EZEK|16|60|Но Я вспомню союз Мой с тобою во дни юности твоей, и восстановлю с тобою вечный союз.
EZEK|16|61|И ты вспомнишь о путях твоих, и будет стыдно тебе, когда станешь принимать к себе сестер твоих, больших тебя, как и меньших тебя, и когда Я буду давать тебе их в дочерей, но не от твоего союза.
EZEK|16|62|Я восстановлю союз Мой с тобою, и узнаешь, что Я Господь,
EZEK|16|63|для того, чтобы ты помнила и стыдилась, и чтобы вперед нельзя было тебе и рта открыть от стыда, когда Я прощу тебе все, что ты делала, говорит Господь Бог.
EZEK|17|1|И было ко мне слово Господне:
EZEK|17|2|сын человеческий! предложи загадку и скажи притчу к дому Израилеву.
EZEK|17|3|Скажи: так говорит Господь Бог: большой орел с большими крыльями, с длинными перьями, пушистый, пестрый, прилетел на Ливан и снял с кедра верхушку,
EZEK|17|4|сорвал верхний из молодых побегов его и принес его в землю Ханаанскую, в городе торговцев положил его;
EZEK|17|5|и взял от семени этой земли, и посадил на земле семени, поместил у больших вод, как сажают иву.
EZEK|17|6|И оно выросло, и сделалось виноградною лозою, широкою, низкою ростом, которой ветви клонились к ней, и корни ее были под нею же, и стало виноградною лозою, и дало отрасли, и пустило ветви.
EZEK|17|7|И еще был орел с большими крыльями и пушистый; и вот, эта виноградная лоза потянулась к нему своими корнями и простерла к нему ветви свои, чтобы он поливал ее из борозд рассадника своего.
EZEK|17|8|Она была посажена на хорошем поле, у больших вод, так что могла пускать ветви и приносить плод, сделаться лозою великолепною.
EZEK|17|9|Скажи: так говорит Господь Бог: будет ли ей успех? Не вырвут ли корней ее, и не оборвут ли плодов ее, так что она засохнет? все молодые ветви, отросшие от нее, засохнут. И не с большою силою и не со многими людьми сорвут ее с корней ее.
EZEK|17|10|И вот, хотя она посажена, но будет ли успех? Не иссохнет ли она, как скоро коснется ее восточный ветер? иссохнет на грядах, где выросла.
EZEK|17|11|И было ко мне слово Господне:
EZEK|17|12|скажи мятежному дому: разве не знаете, что это значит? – Скажи: вот, пришел царь Вавилонский в Иерусалим, и взял царя его и князей его, и привел их к себе в Вавилон.
EZEK|17|13|И взял [другого] из царского рода, и заключил с ним союз, и обязал его клятвою, и взял сильных земли той с собою,
EZEK|17|14|чтобы царство было покорное, чтобы не могло подняться, чтобы сохраняем был союз и стоял твердо.
EZEK|17|15|Но тот отложился от него, послав послов своих в Египет, чтобы дали ему коней и много людей. Будет ли ему успех? Уцелеет ли тот, кто это делает? Он нарушил союз и уцелеет ли?
EZEK|17|16|Живу Я, говорит Господь Бог: в местопребывании царя, который поставил его царем, и которому данную клятву он презрел, и нарушил союз свой с ним, он умрет у него в Вавилоне.
EZEK|17|17|С великою силою и с многочисленным народом фараон ничего не сделает для него в этой войне, когда будет насыпан вал и построены будут осадные башни на погибель многих душ.
EZEK|17|18|Он презрел клятву, чтобы нарушить союз, и вот, дал руку свою и сделал все это; он не уцелеет.
EZEK|17|19|Посему так говорит Господь Бог: живу Я! клятву Мою, которую он презрел, и союз Мой, который он нарушил, Я обращу на его голову.
EZEK|17|20|И закину на него сеть Мою, и пойман будет в тенета Мои; и приведу его в Вавилон, и там буду судиться с ним за вероломство его против Меня.
EZEK|17|21|А все беглецы его из всех полков его падут от меча, а оставшиеся развеяны будут по всем ветрам; и узнаете, что Я, Господь, сказал это.
EZEK|17|22|Так говорит Господь Бог: и возьму Я с вершины высокого кедра, и посажу; с верхних побегов его оторву нежную отрасль и посажу на высокой и величественной горе.
EZEK|17|23|На высокой горе Израилевой посажу его, и пустит ветви, и принесет плод, и сделается величественным кедром, и будут обитать под ним всякие птицы, всякие пернатые будут обитать в тени ветвей его.
EZEK|17|24|И узнают все дерева полевые, что Я, Господь, высокое дерево понижаю, низкое дерево повышаю, зеленеющее дерево иссушаю, а сухое дерево делаю цветущим: Я, Господь, сказал, и сделаю.
EZEK|18|1|И было ко мне слово Господне:
EZEK|18|2|зачем вы употребляете в земле Израилевой эту пословицу, говоря: "отцы ели кислый виноград, а у детей на зубах оскомина"?
EZEK|18|3|Живу Я! говорит Господь Бог, – не будут вперед говорить пословицу эту в Израиле.
EZEK|18|4|Ибо вот, все души – Мои: как душа отца, так и душа сына – Мои: душа согрешающая, та умрет.
EZEK|18|5|Если кто праведен и творит суд и правду,
EZEK|18|6|на горах жертвенного не ест и к идолам дома Израилева не обращает глаз своих, жены ближнего своего не оскверняет и к своей жене во время очищения нечистот ее не приближается,
EZEK|18|7|никого не притесняет, должнику возвращает залог его, хищения не производит, хлеб свой дает голодному и нагого покрывает одеждою,
EZEK|18|8|в рост не отдает и лихвы не берет, от неправды удерживает руку свою, суд человеку с человеком производит правильный,
EZEK|18|9|поступает по заповедям Моим и соблюдает постановления Мои искренно: то он праведник, он непременно будет жив, говорит Господь Бог.
EZEK|18|10|Но если у него родился сын разбойник, проливающий кровь, и делает что–нибудь из всего того,
EZEK|18|11|чего он сам не делал совсем, и на горах ест жертвенное, и жену ближнего своего оскверняет,
EZEK|18|12|бедного и нищего притесняет, насильно отнимает, залога не возвращает, и к идолам обращает глаза свои, делает мерзость,
EZEK|18|13|в рост дает, и берет лихву; то будет ли он жив? [Нет], он не будет жив. Кто делает все такие мерзости, тот непременно умрет, кровь его будет на нем.
EZEK|18|14|Но если у кого родился сын, который, видя все грехи отца своего, какие он делает, видит и не делает подобного им:
EZEK|18|15|на горах жертвенного не ест, к идолам дома Израилева не обращает глаз своих, жены ближнего своего не оскверняет,
EZEK|18|16|и человека не притесняет, залога не берет, и насильно не отнимает, хлеб свой дает голодному, и нагого покрывает одеждою,
EZEK|18|17|от [обиды] бедному удерживает руку свою, роста и лихвы не берет, исполняет Мои повеления и поступает по заповедям Моим, – то сей не умрет за беззаконие отца своего; он будет жив.
EZEK|18|18|А отец его, так как он жестоко притеснял, грабил брата и недоброе делал среди народа своего, вот, он умрет за свое беззаконие.
EZEK|18|19|Вы говорите: "почему же сын не несет вины отца своего?" Потому что сын поступает законно и праведно, все уставы Мои соблюдает и исполняет их; он будет жив.
EZEK|18|20|Душа согрешающая, она умрет; сын не понесет вины отца, и отец не понесет вины сына, правда праведного при нем и остается, и беззаконие беззаконного при нем и остается.
EZEK|18|21|И беззаконник, если обратится от всех грехов своих, какие делал, и будет соблюдать все уставы Мои и поступать законно и праведно, жив будет, не умрет.
EZEK|18|22|Все преступления его, какие делал он, не припомнятся ему: в правде своей, которую будет делать, он жив будет.
EZEK|18|23|Разве Я хочу смерти беззаконника? говорит Господь Бог. Не того ли, чтобы он обратился от путей своих и был жив?
EZEK|18|24|И праведник, если отступит от правды своей и будет поступать неправедно, будет делать все те мерзости, какие делает беззаконник, будет ли он жив? все добрые дела его, какие он делал, не припомнятся; за беззаконие свое, какое делает, и за грехи свои, в каких грешен, он умрет.
EZEK|18|25|Но вы говорите: "неправ путь Господа!" Послушайте, дом Израилев! Мой ли путь неправ? не ваши ли пути неправы?
EZEK|18|26|Если праведник отступает от правды своей и делает беззаконие и за то умирает, то он умирает за беззаконие свое, которое сделал.
EZEK|18|27|И беззаконник, если обращается от беззакония своего, какое делал, и творит суд и правду, – к жизни возвратит душу свою.
EZEK|18|28|Ибо он увидел и обратился от всех преступлений своих, какие делал; он будет жив, не умрет.
EZEK|18|29|А дом Израилев говорит: "неправ путь Господа!" Мои ли пути неправы, дом Израилев? не ваши ли пути неправы?
EZEK|18|30|Посему Я буду судить вас, дом Израилев, каждого по путям его, говорит Господь Бог; покайтесь и обратитесь от всех преступлений ваших, чтобы нечестие не было вам преткновением.
EZEK|18|31|Отвергните от себя все грехи ваши, которыми согрешали вы, и сотворите себе новое сердце и новый дух; и зачем вам умирать, дом Израилев?
EZEK|18|32|Ибо Я не хочу смерти умирающего, говорит Господь Бог; но обратитесь, и живите!
EZEK|19|1|А ты подними плач о князьях Израиля
EZEK|19|2|и скажи: что за львица мать твоя? расположилась среди львов, между молодыми львами растила львенков своих.
EZEK|19|3|И вскормила одного из львенков своих; он сделался молодым львом и научился ловить добычу, ел людей.
EZEK|19|4|И услышали о нем народы; он пойман был в яму их, и в цепях отвели его в землю Египетскую.
EZEK|19|5|И когда, пождав, увидела она, что надежда ее пропала, тогда взяла другого из львенков своих и сделала его молодым львом.
EZEK|19|6|И, сделавшись молодым львом, он стал ходить между львами и научился ловить добычу, ел людей
EZEK|19|7|и осквернял вдов их и города их опустошал; и опустела земля и все селения ее от рыкания его.
EZEK|19|8|Тогда восстали на него народы из окрестных областей и раскинули на него сеть свою; он пойман был в яму их.
EZEK|19|9|И посадили его в клетку на цепи и отвели его к царю Вавилонскому; отвели его в крепость, чтобы не слышен уже был голос его на горах Израилевых.
EZEK|19|10|Твоя мать была, как виноградная лоза, посаженная у воды; плодовита и ветвиста была она от обилия воды.
EZEK|19|11|И были у нее ветви крепкие для скипетров властителей, и высоко поднялся ствол ее между густыми ветвями; и выдавалась она высотою своею со множеством ветвей своих.
EZEK|19|12|Но во гневе вырвана, брошена на землю, и восточный ветер иссушил плод ее; отторжены и иссохли крепкие ветви ее, огонь пожрал их.
EZEK|19|13|А теперь она пересажена в пустыню, в землю сухую и жаждущую.
EZEK|19|14|И вышел огонь из ствола ветвей ее, пожрал плоды ее и не осталось на ней ветвей крепких для скипетра властителя. Это плачевная песнь, и останется для плача.
EZEK|20|1|В седьмом году, в пятом [месяце], в десятый день месяца, пришли мужи из старейшин Израилевых вопросить Господа и сели перед лицем моим.
EZEK|20|2|И было ко мне слово Господне:
EZEK|20|3|сын человеческий! говори со старейшинами Израилевыми и скажи им: так говорит Господь Бог: вы пришли вопросить Меня? Живу Я, не дам вам ответа, говорит Господь Бог.
EZEK|20|4|Хочешь ли судиться с ними, хочешь ли судиться, сын человеческий? выскажи им мерзости отцов их
EZEK|20|5|и скажи им: так говорит Господь Бог: в тот день, когда Я избрал Израиля и, подняв руку Мою, [поклялся] племени дома Иаковлева, и открыл Себя им в земле Египетской, и, подняв руку, сказал им: "Я Господь Бог ваш!" –
EZEK|20|6|в тот день, подняв руку Мою, Я поклялся им вывести их из земли Египетской в землю, которую Я усмотрел для них, текущую молоком и медом, красу всех земель,
EZEK|20|7|и сказал им: отвергните каждый мерзости от очей ваших и не оскверняйте себя идолами Египетскими: Я Господь Бог ваш.
EZEK|20|8|Но они возмутились против Меня и не хотели слушать Меня; никто не отверг мерзостей от очей своих и не оставил идолов Египетских. И Я сказал: изолью на них гнев Мой, истощу на них ярость Мою среди земли Египетской.
EZEK|20|9|Но Я поступил ради имени Моего, чтобы оно не хулилось перед народами, среди которых находились они и перед глазами которых Я открыл Себя им, чтобы вывести их из земли Египетской.
EZEK|20|10|И Я вывел их из земли Египетской и привел их в пустыню,
EZEK|20|11|и дал им заповеди Мои, и объявил им Мои постановления, исполняя которые человек жив был бы через них;
EZEK|20|12|дал им также субботы Мои, чтобы они были знамением между Мною и ими, чтобы знали, что Я Господь, освящающий их.
EZEK|20|13|Но дом Израилев возмутился против Меня в пустыне: по заповедям Моим не поступали и отвергли постановления Мои, исполняя которые человек жив был бы через них, и субботы Мои нарушали, и Я сказал: изолью на них ярость Мою в пустыне, чтобы истребить их.
EZEK|20|14|Но Я поступил ради имени Моего, чтобы оно не хулилось перед народами, в глазах которых Я вывел их.
EZEK|20|15|Даже Я, подняв руку Мою против них в пустыне, [поклялся], что не введу их в землю, которую Я назначил, – текущую молоком и медом, красу всех земель, –
EZEK|20|16|за то, что они отвергли постановления Мои, и не поступали по заповедям Моим, и нарушали субботы Мои; ибо сердце их стремилось к идолам их.
EZEK|20|17|Но око Мое пожалело погубить их; и Я не истребил их в пустыне.
EZEK|20|18|И говорил Я сыновьям их в пустыне: не ходите по правилам отцов ваших, и не соблюдайте установлений их, и не оскверняйте себя идолами их.
EZEK|20|19|Я Господь Бог ваш: по Моим заповедям поступайте, и Мои уставы соблюдайте, и исполняйте их.
EZEK|20|20|И святите субботы Мои, чтобы они были знамением между Мною и вами, дабы вы знали, что Я Господь Бог ваш.
EZEK|20|21|Но и сыновья возмутились против Меня: по заповедям Моим не поступали и уставов Моих не соблюдали, не исполняли того, что исполняя, человек был бы жив, нарушали субботы Мои, – и Я сказал: изолью на них гнев Мой, истощу над ними ярость Мою в пустыне;
EZEK|20|22|но Я отклонил руку Мою и поступил ради имени Моего, чтобы оно не хулилось перед народами, перед глазами которых Я вывел их.
EZEK|20|23|Также, подняв руку Мою в пустыне, Я [поклялся] рассеять их по народам и развеять их по землям
EZEK|20|24|за то, что они постановлений Моих не исполняли и заповеди Мои отвергли, и нарушали субботы мои, и глаза их обращались к идолам отцов их.
EZEK|20|25|И попустил им учреждения недобрые и постановления, от которых они не могли быть живы,
EZEK|20|26|и попустил им оскверниться жертвоприношениями их, когда они стали проводить через огонь всякий первый плод утробы, чтобы разорить их, дабы знали, что Я Господь.
EZEK|20|27|Посему говори дому Израилеву, сын человеческий, и скажи им: так говорит Господь Бог: вот чем еще хулили Меня отцы ваши, вероломно поступая против Меня:
EZEK|20|28|Я привел их в землю, которую клятвенно обещал дать им, подняв руку Мою, – а они, высмотрев себе всякий высокий холм и всякое ветвистое дерево, стали заколать там жертвы свои, и ставили там оскорбительные для Меня приношения свои и благовонные курения свои, и возливали там возлияния свои.
EZEK|20|29|И Я говорил им: что это за высота, куда ходите вы? поэтому именем Бама называется она и до сего дня.
EZEK|20|30|Посему скажи дому Израилеву: так говорит Господь Бог: не оскверняете ли вы себя по примеру отцов ваших и не блудодействуете ли вслед мерзостей их?
EZEK|20|31|Принося дары ваши и проводя сыновей ваших через огонь, вы оскверняете себя всеми идолами вашими до сего дня, и хотите вопросить Меня, дом Израилев? живу Я, говорит Господь Бог, не дам вам ответа.
EZEK|20|32|И что приходит вам на ум, совсем не сбудется. Вы говорите: "будем, как язычники, как племена иноземные, служить дереву и камню".
EZEK|20|33|Живу Я, говорит Господь Бог: рукою крепкою и мышцею простертою и излиянием ярости буду господствовать над вами.
EZEK|20|34|И выведу вас из народов и из стран, по которым вы рассеяны, и соберу вас рукою крепкою и мышцею простертою и излиянием ярости.
EZEK|20|35|И приведу вас в пустыню народов, и там буду судиться с вами лицом к лицу.
EZEK|20|36|Как Я судился с отцами вашими в пустыне земли Египетской, так буду судиться с вами, говорит Господь Бог.
EZEK|20|37|И проведу вас под жезлом и введу вас в узы завета.
EZEK|20|38|И выделю из вас мятежников и непокорных Мне. Из земли пребывания их выведу их, но в землю Израилеву они не войдут, и узнаете, что Я Господь.
EZEK|20|39|А вы, дом Израилев, – так говорит Господь Бог, – идите каждый к своим идолам и служите им, если Меня не слушаете, но не оскверняйте более святаго имени Моего дарами вашими и идолами вашими,
EZEK|20|40|потому что на Моей святой горе, на горе высокой Израилевой, – говорит Господь Бог, – там будет служить Мне весь дом Израилев, – весь, сколько ни есть его на земле; там Я с благоволением приму их, и там потребую приношений ваших и начатков ваших со всеми святынями вашими.
EZEK|20|41|Приму вас, как благовонное курение, когда выведу вас из народов и соберу вас из стран, по которым вы рассеяны, и буду святиться в вас перед глазами народов.
EZEK|20|42|И узнаете, что Я Господь, когда введу вас в землю Израилеву, – в землю, которую Я [клялся] дать отцам вашим, подняв руку Мою.
EZEK|20|43|И вспомните там о путях ваших и обо всех делах ваших, какими вы оскверняли себя, и возгнушаетесь самими собою за все злодеяния ваши, какие вы делали.
EZEK|20|44|И узнаете, что Я Господь, когда буду поступать с вами ради имени Моего, не по злым вашим путям и вашим делам развратным, дом Израилев, – говорит Господь Бог.
EZEK|21|1|И было ко мне слово Господне:
EZEK|21|2|сын человеческий! обрати лице твое на путь к полудню, и произнеси слово на полдень, и изреки пророчество на лес южного поля.
EZEK|21|3|И скажи южному лесу: слушай слово Господа; так говорит Господь Бог: вот, Я зажгу в тебе огонь, и он пожрет в тебе всякое дерево зеленеющее и всякое дерево сухое; не погаснет пылающий пламень, и все будет опалено им от юга до севера.
EZEK|21|4|И увидит всякая плоть, что Я, Господь, зажег его, и он не погаснет.
EZEK|21|5|И сказал я: о, Господи Боже! они говорят обо мне: "не говорит ли он притчи?"
EZEK|21|6|И было ко мне слово Господне:
EZEK|21|7|сын человеческий! обрати лице твое к Иерусалиму и произнеси слово на святилища, и изреки пророчество на землю Израилеву,
EZEK|21|8|и скажи земле Израилевой: так говорит Господь Бог: вот, Я – на тебя, и извлеку меч Мой из ножен его и истреблю у тебя праведного и нечестивого.
EZEK|21|9|А для того, чтобы истребить у тебя праведного и нечестивого, меч Мой из ножен своих пойдет на всякую плоть от юга до севера.
EZEK|21|10|И узнает всякая плоть, что Я, Господь, извлек меч Мой из ножен его, и он уже не возвратится.
EZEK|21|11|Ты же, сын человеческий, стенай, сокрушая бедра твои, и в горести стенай перед глазами их.
EZEK|21|12|И когда скажут тебе: "отчего ты стенаешь?", скажи: "от слуха, что идет", – и растает всякое сердце, и все руки опустятся, и всякий дух изнеможет, и все колени задрожат, как вода. Вот, это придет и сбудется, говорит Господь Бог.
EZEK|21|13|И было ко мне слово Господне:
EZEK|21|14|сын человеческий! изреки пророчество и скажи: так говорит Господь Бог: скажи: меч, меч наострен и вычищен;
EZEK|21|15|наострен для того, чтобы больше заколать; вычищен, чтобы сверкал, как молния. Радоваться ли нам, что жезл сына Моего презирает всякое дерево?
EZEK|21|16|Я дал его вычистить, чтобы взять в руку; уже наострен этот меч и вычищен, чтобы отдать его в руку убийцы.
EZEK|21|17|Стенай и рыдай, сын человеческий, ибо он – на народ Мой, на всех князей Израиля; они отданы будут под меч с народом Моим; посему ударяй себя по бедрам.
EZEK|21|18|Ибо он уже испытан. И что, если он презирает и жезл? сей не устоит, говорит Господь Бог.
EZEK|21|19|Ты же, сын человеческий, пророчествуй и ударяй рукою об руку; и удвоится меч и утроится, меч на поражаемых, меч на поражение великого, проникающий во внутренность жилищ их.
EZEK|21|20|Чтобы растаяли сердца и чтобы павших было более, Я у всех ворот их поставлю грозный меч, увы! сверкающий, как молния, наостренный для заклания.
EZEK|21|21|Соберись и иди направо или иди налево, куда бы ни обратилось лице твое.
EZEK|21|22|И Я буду рукоплескать и утолю гнев Мой; Я, Господь, сказал.
EZEK|21|23|И было ко мне слово Господне:
EZEK|21|24|и ты, сын человеческий, представь себе две дороги, по которым должно идти мечу царя Вавилонского, – обе они должны выходить из одной земли; и начертай руку, начертай при начале дорог в города.
EZEK|21|25|Представь дорогу, по которой меч шел бы в Равву сынов Аммоновых и в Иудею, в укрепленный Иерусалим;
EZEK|21|26|потому что царь Вавилонский остановился на распутье, при начале двух дорог, для гаданья: трясет стрелы, вопрошает терафимов, рассматривает печень.
EZEK|21|27|В правой руке у него гаданье: "в Иерусалим", где должно поставить тараны, открыть для побоища уста, возвысить голос для военного крика, подвести тараны к воротам, насыпать вал, построить осадные башни.
EZEK|21|28|Это гаданье показалось в глазах их лживым; но так как они клялись клятвою, то он, вспомнив о таком их вероломстве, положил взять его.
EZEK|21|29|Посему так говорит Господь Бог: так как вы сами приводите на память беззаконие ваше, делая явными преступления ваши, выставляя на вид грехи ваши во всех делах ваших, и сами приводите это на память, то вы будете взяты руками.
EZEK|21|30|И ты, недостойный, преступный вождь Израиля, которого день наступил ныне, когда нечестию его положен будет конец!
EZEK|21|31|так говорит Господь Бог: сними с себя диадему и сложи венец; этого уже не будет; униженное возвысится и высокое унизится.
EZEK|21|32|Низложу, низложу, низложу и его не будет, доколе не придет Тот, Кому [принадлежит] он, и Я дам Ему.
EZEK|21|33|И ты, сын человеческий, изреки пророчество и скажи: так говорит Господь Бог о сынах Аммона и о поношении их; и скажи: меч, меч обнажен для заклания, вычищен для истребления, чтобы сверкал, как молния,
EZEK|21|34|чтобы, тогда как представляют тебе пустые видения и ложно гадают тебе, и тебя приложил к обезглавленным нечестивцам, которых день наступил, когда нечестию их положен будет конец.
EZEK|21|35|Возвратить ли его в ножны его? – на месте, где ты сотворен, на земле происхождения твоего буду судить тебя:
EZEK|21|36|и изолью на тебя негодование Мое, дохну на тебя огнем ярости Моей и отдам тебя в руки людей свирепых, опытных в убийстве.
EZEK|21|37|Ты будешь пищею огню, кровь твоя останется на земле; не будут и вспоминать о тебе; ибо Я, Господь, сказал это.
EZEK|22|1|И было ко мне слово Господне:
EZEK|22|2|и ты, сын человеческий, хочешь ли судить, судить город кровей? выскажи ему все мерзости его.
EZEK|22|3|И скажи: так говорит Господь Бог: о, город, проливающий кровь среди себя, чтобы наступило время твое, и делающий у себя идолов, чтобы осквернять себя!
EZEK|22|4|Кровью, которую ты пролил, ты сделал себя виновным, и идолами, каких ты наделал, ты осквернил себя, и приблизил дни твои и достиг годины твоей. За это отдам тебя на посмеяние народам, на поругание всем землям.
EZEK|22|5|Близкие и далекие от тебя будут ругаться над тобою, осквернившим имя твое, прославившимся буйством.
EZEK|22|6|Вот, начальствующие у Израиля, каждый по мере сил своих, были у тебя, чтобы проливать кровь.
EZEK|22|7|У тебя отца и мать злословят, пришельцу делают обиду среди тебя, сироту и вдову притесняют у тебя.
EZEK|22|8|Святынь Моих ты не уважаешь и субботы Мои нарушаешь.
EZEK|22|9|Клеветники находятся в тебе, чтобы проливать кровь, и на горах едят у тебя [идоложертвенное], среди тебя производят гнусность.
EZEK|22|10|Наготу отца открывают у тебя, жену во время очищения нечистот ее насилуют у тебя.
EZEK|22|11|Иной делает мерзость с женою ближнего своего, иной оскверняет сноху свою, иной насилует сестру свою, дочь отца своего.
EZEK|22|12|Взятки берут у тебя, чтобы проливать кровь; ты берешь рост и лихву и насилием вымогаешь корысть у ближнего твоего, а Меня забыл, говорит Господь Бог.
EZEK|22|13|И вот, Я всплеснул руками Моими о корыстолюбии твоем, какое обнаруживается у тебя, и о кровопролитии, которое совершается среди тебя.
EZEK|22|14|Устоит ли сердце твое, будут ли тверды руки твои в те дни, в которые буду действовать против тебя? Я, Господь, сказал и сделаю.
EZEK|22|15|И рассею тебя по народам, и развею тебя по землям, и положу конец мерзостям твоим среди тебя.
EZEK|22|16|И сделаешь сам себя презренным перед глазами народов, и узнаешь, что Я Господь.
EZEK|22|17|И было ко мне слово Господне:
EZEK|22|18|сын человеческий! дом Израилев сделался у Меня изгарью; все они – олово, медь и железо и свинец в горниле, сделались, как изгарь серебра.
EZEK|22|19|Посему так говорит Господь Бог: так как все вы сделались изгарью, за то вот, Я соберу вас в Иерусалим.
EZEK|22|20|Как в горнило кладут вместе серебро, и медь, и железо, и свинец, и олово, чтобы раздуть на них огонь и расплавить; так Я во гневе Моем и в ярости Моей соберу, и положу, и расплавлю вас.
EZEK|22|21|Соберу вас и дохну на вас огнем негодования Моего, и расплавитесь среди него.
EZEK|22|22|Как серебро расплавляется в горниле, так расплавитесь и вы среди него, и узнаете, что Я, Господь, излил ярость Мою на вас.
EZEK|22|23|И было ко мне слово Господне:
EZEK|22|24|сын человеческий! скажи ему: ты – земля неочищенная, не орошаемая дождем в день гнева!
EZEK|22|25|Заговор пророков ее среди нее – как лев рыкающий, терзающий добычу; съедают души, обирают имущество и драгоценности, и умножают число вдов.
EZEK|22|26|Священники ее нарушают закон Мой и оскверняют святыни Мои, не отделяют святаго от несвятаго и не указывают различия между чистым и нечистым, и от суббот Моих они закрыли глаза свои, и Я уничижен у них.
EZEK|22|27|Князья у нее как волки, похищающие добычу; проливают кровь, губят души, чтобы приобрести корысть.
EZEK|22|28|А пророки ее все замазывают грязью, видят пустое и предсказывают им ложное, говоря: "так говорит Господь Бог", тогда как не говорил Господь.
EZEK|22|29|А в народе угнетают друг друга, грабят и притесняют бедного и нищего, и пришельца угнетают несправедливо.
EZEK|22|30|Искал Я у них человека, который поставил бы стену и стал бы предо Мною в проломе за сию землю, чтобы Я не погубил ее, но не нашел.
EZEK|22|31|Итак изолью на них негодование Мое, огнем ярости Моей истреблю их, поведение их обращу им на голову, говорит Господь Бог.
EZEK|23|1|И было ко мне слово Господне:
EZEK|23|2|сын человеческий! были две женщины, дочери одной матери,
EZEK|23|3|и блудили они в Египте, блудили в своей молодости; там измяты груди их, и там растлили девственные сосцы их.
EZEK|23|4|Имена им: большой – Огола, а сестре ее – Оголива. И были они Моими, и рождали сыновей и дочерей; и именовались – Огола Самариею, а Оголива Иерусалимом.
EZEK|23|5|И стала Огола блудить от Меня и пристрастилась к своим любовникам, к Ассириянам, к соседям своим,
EZEK|23|6|к одевавшимся в ткани яхонтового цвета, к областеначальникам и градоправителям, ко всем красивым юношам, всадникам, ездящим на конях;
EZEK|23|7|и расточала блудодеяния свои со всеми отборными из сынов Ассура, и оскверняла себя всеми идолами тех, к кому ни пристращалась;
EZEK|23|8|не переставала блудить и с Египтянами, потому что они с нею спали в молодости ее и растлевали девственные сосцы ее, и изливали на нее похоть свою.
EZEK|23|9|За то Я и отдал ее в руки любовников ее, в руки сынов Ассура, к которым она пристрастилась.
EZEK|23|10|Они открыли наготу ее, взяли сыновей ее и дочерей ее, а ее убили мечом. И она сделалась позором между женщинами, когда совершили над нею казнь.
EZEK|23|11|Сестра ее, Оголива, видела это, и еще развращеннее была в любви своей, и блужение ее превзошло блужение сестры ее.
EZEK|23|12|Она пристрастилась к сынам Ассуровым, к областеначальникам и градоправителям, соседям ее, пышно одетым, к всадникам, ездящим на конях, ко всем отборным юношам.
EZEK|23|13|И Я видел, что она осквернила себя, [и что] у обеих их одна дорога.
EZEK|23|14|Но эта еще умножила блудодеяния свои, потому что, увидев вырезанных на стене мужчин, красками нарисованные изображения Халдеев,
EZEK|23|15|опоясанных по чреслам своим поясом, с роскошными на голове их повязками, имеющих вид военачальников, похожих на сынов Вавилона, которых родина земля Халдейская,
EZEK|23|16|она влюбилась в них по одному взгляду очей своих и послала к ним в Халдею послов.
EZEK|23|17|И пришли к ней сыны Вавилона на любовное ложе, и осквернили ее блудодейством своим, и она осквернила себя ими; и отвратилась от них душа ее.
EZEK|23|18|Когда же она явно предалась блудодеяниям своим и открыла наготу свою, тогда и от нее отвратилась душа Моя, как отвратилась душа Моя от сестры ее.
EZEK|23|19|И она умножала блудодеяния свои, вспоминая дни молодости своей, когда блудила в земле Египетской;
EZEK|23|20|и пристрастилась к любовникам своим, у которых плоть – плоть ослиная, и похоть, как у жеребцов.
EZEK|23|21|Так ты вспомнила распутство молодости твоей, когда Египтяне жали сосцы твои из–за девственных грудей твоих.
EZEK|23|22|Посему, Оголива, так говорит Господь Бог: вот, Я возбужу против тебя любовников твоих, от которых отвратилась душа твоя, и приведу их против тебя со всех сторон:
EZEK|23|23|сынов Вавилона и всех Халдеев, из Пехода, из Шоа и Коа, и с ними всех сынов Ассура, красивых юношей, областеначальников и градоправителей, сановных и именитых, всех искусных наездников.
EZEK|23|24|И придут на тебя с оружием, с конями и колесницами и с множеством народа, и обступят тебя кругом в латах, со щитами и в шлемах, и отдам им тебя на суд, и будут судить тебя своим судом.
EZEK|23|25|И обращу ревность Мою против тебя, и поступят с тобою яростно: отрежут у тебя нос и уши, а остальное твое от меча падет; возьмут сыновей твоих и дочерей твоих, а остальное твое огнем будет пожрано;
EZEK|23|26|и снимут с тебя одежды твои, возьмут наряды твои.
EZEK|23|27|И положу конец распутству твоему и блужению твоему, принесенному из земли Египетской, и не будешь обращать к ним глаз твоих, и о Египте уже не вспомнишь.
EZEK|23|28|Ибо так говорит Господь Бог: вот, Я предаю тебя в руки тех, которых ты возненавидела, в руки тех, от которых отвратилась душа твоя.
EZEK|23|29|И поступят с тобою жестоко, и возьмут у тебя все, нажитое трудами, и оставят тебя нагою и непокрытою, и открыта будет срамная нагота твоя, и распутство твое, и блудодейство твое.
EZEK|23|30|Это будет сделано с тобою за блудодейство твое с народами, которых идолами ты осквернила себя.
EZEK|23|31|Ты ходила дорогою сестры твоей; за то и дам в руку тебе чашу ее.
EZEK|23|32|Так говорит Господь Бог: ты будешь пить чашу сестры твоей, глубокую и широкую, и подвергнешься посмеянию и позору, по огромной вместительности ее.
EZEK|23|33|Опьянения и горести будешь исполнена: чаша ужаса и опустошения – чаша сестры твоей, Самарии!
EZEK|23|34|И выпьешь ее, и осушишь, и черепки ее оближешь, и груди твои истерзаешь: ибо Я сказал это, говорит Господь Бог.
EZEK|23|35|Посему так говорит Господь Бог: так как ты забыла Меня и отвратилась от Меня, то и терпи за беззаконие твое и за блудодейство твое.
EZEK|23|36|И сказал мне Господь: сын человеческий! хочешь ли судить Оголу и Оголиву? выскажи им мерзости их;
EZEK|23|37|ибо они прелюбодействовали, и кровь на руках их, и с идолами своими прелюбодействовали, и сыновей своих, которых родили Мне, через огонь проводили в пищу им.
EZEK|23|38|Еще вот что они делали Мне: оскверняли святилище Мое в тот же день, и нарушали субботы Мои;
EZEK|23|39|потому что, когда они заколали детей своих для идолов своих, в тот же день приходили в святилище Мое, чтобы осквернять его: вот как поступали они в доме Моем!
EZEK|23|40|Кроме сего посылали за людьми, приходившими издалека; к ним отправляли послов, и вот, они приходили, и ты для них умывалась, сурьмила глаза твои и украшалась нарядами,
EZEK|23|41|и садились на великолепное ложе, перед которым приготовляем был стол и на котором предлагала ты благовонные курения Мои и елей Мой.
EZEK|23|42|И раздавался голос народа, ликовавшего у нее, и к людям из толпы народной вводимы были пьяницы из пустыни; и они возлагали на руки их запястья и на головы их красивые венки.
EZEK|23|43|Тогда сказал Я об одряхлевшей в прелюбодействе: теперь кончатся блудодеяния ее вместе с нею.
EZEK|23|44|Но приходили к ней, как приходят к жене блуднице, так приходили к Оголе и Оголиве, к распутным женам.
EZEK|23|45|Но мужи праведные будут судить их; они будут судить их судом прелюбодейц и судом проливающих кровь, потому что они прелюбодейки, и у них кровь на руках.
EZEK|23|46|Ибо так сказал Господь Бог: созвать на них собрание и предать их озлоблению и грабежу.
EZEK|23|47|И собрание побьет их камнями, и изрубит их мечами своими, и убьет сыновей их и дочерей их, и домы их сожжет огнем.
EZEK|23|48|Так положу конец распутству на сей земле, и все женщины примут урок, и не будут делать срамных дел подобно вам;
EZEK|23|49|и возложат на вас ваше распутство, и понесете наказание за грехи с идолами вашими, и узнаете, что Я Господь Бог.
EZEK|24|1|И было ко мне слово Господне в девятом году, в десятом месяце, в десятый день месяца:
EZEK|24|2|сын человеческий! запиши себе имя этого дня, этого самого дня: в этот самый день царь Вавилонский подступит к Иерусалиму.
EZEK|24|3|И произнеси на мятежный дом притчу, и скажи им: так говорит Господь Бог: поставь котел, поставь и налей в него воды;
EZEK|24|4|сложи в него куски мяса, все лучшие куски, бедра и плеча, и наполни отборными костями;
EZEK|24|5|отборных овец возьми, и [разожги] под ним кости, и кипяти до того, чтобы и кости разварились в нем.
EZEK|24|6|Посему так говорит Господь Бог: горе городу кровей! горе котлу, в котором есть накипь и с которого накипь его не сходит! кусок за куском его выбрасывайте из него, не выбирая по жребию.
EZEK|24|7|Ибо кровь его среди него; он оставил ее на голой скале; не на землю проливал ее, где она могла бы покрыться пылью.
EZEK|24|8|Чтобы возбудить гнев для совершения мщения, Я оставил кровь его на голой скале, чтобы она не скрылась.
EZEK|24|9|Посему так говорит Господь Бог: горе городу кровей! и Я разложу большой костер.
EZEK|24|10|Прибавь дров, разведи огонь, вывари мясо; пусть все сгустится, и кости перегорят.
EZEK|24|11|И когда котел будет пуст, поставь его на уголья, чтобы он разгорелся, и чтобы медь его раскалилась, и расплавилась в нем нечистота его, и вся накипь его исчезла.
EZEK|24|12|Труд будет тяжелый; но большая накипь его не сойдет с него; и в огне [останется] на нем накипь его.
EZEK|24|13|В нечистоте твоей такая мерзость, что, сколько Я ни чищу тебя, ты все нечист; от нечистоты твоей ты и впредь не очистишься, доколе ярости Моей Я не утолю над тобою.
EZEK|24|14|Я Господь, Я говорю: это придет и Я сделаю; не отменю и не пощажу, и не помилую. По путям твоим и по делам твоим будут судить тебя, говорит Господь Бог.
EZEK|24|15|И было ко мне слово Господне:
EZEK|24|16|сын человеческий! вот, Я возьму у тебя язвою утеху очей твоих; но ты не сетуй и не плачь, и слезы да не выступают у тебя;
EZEK|24|17|вздыхай в безмолвии, плача по умершим не совершай; но обвязывай себя повязкою и обувай ноги твои в обувь твою, и бороды не закрывай, и хлеба от чужих не ешь.
EZEK|24|18|И после того, как говорил я поутру слово к народу, вечером умерла жена моя, и на другой день я сделал так, как повелено было мне.
EZEK|24|19|И сказал мне народ: не скажешь ли нам, какое для нас значение в том, что ты делаешь?
EZEK|24|20|И сказал я им: ко мне было слово Господне:
EZEK|24|21|скажи дому Израилеву: так говорит Господь Бог: вот, Я отдам на поругание святилище Мое, опору силы вашей, утеху очей ваших и отраду души вашей, а сыновья ваши и дочери ваши, которых вы оставили, падут от меча.
EZEK|24|22|И вы будете делать то же, что делал я; бороды не будете закрывать, и хлеба от чужих не будете есть;
EZEK|24|23|и повязки ваши будут на головах ваших, и обувь ваша на ногах ваших; не будете сетовать и плакать, но будете истаявать от грехов ваших и воздыхать друг перед другом.
EZEK|24|24|И будет для вас Иезекииль знамением: все, что он делал, и вы будете делать; и когда это сбудется, узнаете, что Я Господь Бог.
EZEK|24|25|А что до тебя, сын человеческий, то в тот день, когда Я возьму у них украшение славы их, утеху очей их и отраду души их, сыновей их и дочерей их, –
EZEK|24|26|в тот день придет к тебе спасшийся [оттуда], чтобы подать весть в уши твои.
EZEK|24|27|В тот день при этом спасшемся откроются уста твои, и ты будешь говорить, и не останешься уже безмолвным, и будешь знамением для них, и узнают, что Я Господь.
EZEK|25|1|И было ко мне слово Господне:
EZEK|25|2|сын человеческий! обрати лице твое к сынам Аммоновым и изреки на них пророчество,
EZEK|25|3|и скажи сынам Аммоновым: слушайте слово Господа Бога: так говорит Господь Бог: за то, что ты о святилище Моем говоришь: "а! а!", потому что оно поругано, – и о земле Израилевой, потому что она опустошена, и о доме Иудином, потому что они пошли в плен, –
EZEK|25|4|за то вот, Я отдам тебя в наследие сынам востока, и построят у тебя овчарни свои, и поставят у тебя шатры свои, и будут есть плоды твои и пить молоко твое.
EZEK|25|5|Я сделаю Равву стойлом для верблюдов, и сынов Аммоновых – пастухами овец, и узнаете, что Я Господь.
EZEK|25|6|Ибо так говорит Господь Бог: за то, что ты рукоплескал и топал ногою, и со всем презрением к земле Израилевой душевно радовался, –
EZEK|25|7|за то вот, Я простру руку Мою на тебя и отдам тебя на расхищение народам, и истреблю тебя из числа народов, и изглажу тебя из числа земель; сокрушу тебя, и узнаешь, что Я Господь.
EZEK|25|8|Так говорит Господь Бог: за то, что Моав и Сеир говорят: "вот и дом Иудин, как все народы!",
EZEK|25|9|за то вот, Я, [начиная] от городов, от всех пограничных городов его, красы земли, от Беф–Иешимофа, Ваалмеона и Кириафаима, открою бок Моава
EZEK|25|10|для сынов востока и отдам его в наследие [им], вместе с сынами Аммоновыми, чтобы сыны Аммона не упоминались более среди народов.
EZEK|25|11|И над Моавом произведу суд, и узнают, что Я Господь.
EZEK|25|12|Так говорит Господь Бог: за то, что Едом жестоко мстил дому Иудину и тяжко согрешил, совершая над ним мщение,
EZEK|25|13|за то, так говорит Господь Бог: простру руку Мою на Едома и истреблю у него людей и скот, и сделаю его пустынею; от Фемана до Дедана все падут от меча.
EZEK|25|14|И совершу мщение Мое над Едомом рукою народа Моего, Израиля; и они будут действовать в Идумее по Моему гневу и Моему негодованию, и узнают мщение Мое, говорит Господь Бог.
EZEK|25|15|Так говорит Господь Бог: за то, что Филистимляне поступили мстительно и мстили с презрением в душе, на погибель, по вечной неприязни,
EZEK|25|16|за то, так говорит Господь Бог: вот, Я простру руку Мою на Филистимлян, и истреблю Критян, и уничтожу остаток их на берегу моря;
EZEK|25|17|и совершу над ними великое мщение наказаниями яростными; и узнают, что Я Господь, когда совершу над ними Мое мщение.
EZEK|26|1|В одиннадцатом году, в первый день первого месяца, было ко мне слово Господне:
EZEK|26|2|сын человеческий! за то, что Тир говорит о Иерусалиме: "а! а! он сокрушен – врата народов; он обращается ко мне; наполнюсь; он опустошен", –
EZEK|26|3|за то, так говорит Господь Бог: вот, Я – на тебя, Тир, и подниму на тебя многие народы, как море поднимает волны свои.
EZEK|26|4|И разобьют стены Тира и разрушат башни его; и вымету из него прах его и сделаю его голою скалою.
EZEK|26|5|Местом для расстилания сетей будет он среди моря; ибо Я сказал это, говорит Господь Бог: и будет он на расхищение народам.
EZEK|26|6|А дочери его, которые на земле, убиты будут мечом, и узнают, что Я Господь.
EZEK|26|7|Ибо так говорит Господь Бог: вот, Я приведу против Тира от севера Навуходоносора, царя Вавилонского, царя царей, с конями и с колесницами, и со всадниками, и с войском, и с многочисленным народом.
EZEK|26|8|Дочерей твоих на земле он побьет мечом и устроит против тебя осадные башни, и насыплет против тебя вал, и поставит против тебя щиты;
EZEK|26|9|и к стенам твоим придвинет стенобитные машины и башни твои разрушит секирами своими.
EZEK|26|10|От множества коней его покроет тебя пыль, от шума всадников и колес и колесниц потрясутся стены твои, когда он будет входить в ворота твои, как входят в разбитый город.
EZEK|26|11|Копытами коней своих он истопчет все улицы твои, народ твой побьет мечом и памятники могущества твоего повергнет на землю.
EZEK|26|12|И разграбят богатство твое, и расхитят товары твои, и разрушат стены твои, и разобьют красивые домы твои, и камни твои и дерева твои, и землю твою бросят в воду.
EZEK|26|13|И прекращу шум песней твоих, и звук цитр твоих уже не будет слышен.
EZEK|26|14|И сделаю тебя голою скалою, будешь местом для расстилания сетей; не будешь вновь построен: ибо Я, Господь, сказал это, говорит Господь Бог.
EZEK|26|15|Так говорит Господь Бог Тиру: от шума падения твоего, от стона раненых, когда будет производимо среди тебя избиение, не содрогнутся ли острова?
EZEK|26|16|И сойдут все князья моря с престолов своих, и сложат с себя мантии свои, и снимут с себя узорчатые одежды свои, облекутся в трепет, сядут на землю, и ежеминутно будут содрогаться и изумляться о тебе.
EZEK|26|17|И поднимут плач о тебе и скажут тебе: как погиб ты, населенный мореходцами, город знаменитый, который был силен на море, сам и жители его, наводившие страх на всех обитателей его!
EZEK|26|18|Ныне, в день падения твоего, содрогнулись острова; острова на море приведены в смятение погибелью твоею.
EZEK|26|19|Ибо так говорит Господь Бог: когда Я сделаю тебя городом опустелым, подобным городам необитаемым, когда подниму на тебя пучину, и покроют тебя большие воды;
EZEK|26|20|тогда низведу тебя с отходящими в могилу к народу давно бывшему, и помещу тебя в преисподних земли, в пустынях вечных, с отшедшими в могилу, чтобы ты не был более населен; и явлю Я славу на земле живых.
EZEK|26|21|Ужасом сделаю тебя, и не будет тебя, и будут искать тебя, но уже не найдут тебя во веки, говорит Господь Бог.
EZEK|27|1|И было ко мне слово Господне:
EZEK|27|2|и ты, сын человеческий, подними плач о Тире
EZEK|27|3|и скажи Тиру, поселившемуся на выступах в море, торгующему с народами на многих островах: так говорит Господь Бог: Тир! ты говоришь: "я совершенство красоты!"
EZEK|27|4|Пределы твои в сердце морей; строители твои усовершили красоту твою:
EZEK|27|5|из Сенирских кипарисов устроили все помосты твои; брали с Ливана кедр, чтобы сделать на тебе мачты;
EZEK|27|6|из дубов Васанских делали весла твои; скамьи твои делали из букового дерева, с оправою из слоновой кости с островов Киттимских;
EZEK|27|7|узорчатые полотна из Египта употреблялись на паруса твои и служили флагом; голубого и пурпурового цвета ткани с островов Елисы были покрывалом твоим.
EZEK|27|8|Жители Сидона и Арвада были у тебя гребцами; свои знатоки были у тебя, Тир; они были у тебя кормчими.
EZEK|27|9|Старшие из Гевала и знатоки его были у тебя, чтобы заделывать пробоины твои. Всякие морские корабли и корабельщики их находились у тебя для производства торговли твоей.
EZEK|27|10|Перс и Лидиянин и Ливиец находились в войске твоем и были у тебя ратниками, вешали на тебе щит и шлем; они придавали тебе величие.
EZEK|27|11|Сыны Арвада с собственным твоим войском стояли кругом на стенах твоих, и Гамадимы были на башнях твоих; кругом по стенам твоим они вешали колчаны свои; они довершали красу твою.
EZEK|27|12|Фарсис, торговец твой, по множеству всякого богатства, платил за товары твои серебром, железом, свинцом и оловом.
EZEK|27|13|Иаван, Фувал и Мешех торговали с тобою, выменивая товары твои на души человеческие и медную посуду.
EZEK|27|14|Из дома Фогарма за товары твои доставляли тебе лошадей и строевых коней и лошаков.
EZEK|27|15|Сыны Дедана торговали с тобою; многие острова производили с тобою мену, в уплату тебе доставляли слоновую кость и черное дерево.
EZEK|27|16|По причине большого торгового производства твоего торговали с тобою Арамеяне; за товары твои они платили карбункулами, тканями пурпуровыми, узорчатыми, и виссонами, и кораллами, и рубинами.
EZEK|27|17|Иудея и земля Израилева торговали с тобою; за товар твой платили пшеницею Миннифскою и сластями, и медом, и деревянным маслом, и бальзамом.
EZEK|27|18|Дамаск, по причине большого торгового производства твоего, по изобилию всякого богатства, торговал с тобою вином Хелбонским и белою шерстью.
EZEK|27|19|Дан и Иаван из Узала платили тебе за товары твои выделанным железом; кассия и благовонная трость шли на обмен тебе.
EZEK|27|20|Дедан торговал с тобою драгоценными попонами для верховой езды.
EZEK|27|21|Аравия и все князья Кидарские производили мену с тобою: ягнят и баранов и козлов променивали тебе.
EZEK|27|22|Купцы из Савы и Раемы торговали с тобою всякими лучшими благовониями и всякими дорогими камнями, и золотом платили за товары твои.
EZEK|27|23|Харан и Хане и Еден, купцы Савейские, Ассур и Хилмад торговали с тобою.
EZEK|27|24|Они торговали с тобою драгоценными одеждами, шелковыми и узорчатыми материями, которые они привозили на твои рынки в дорогих ящиках, сделанных из кедра и хорошо упакованных.
EZEK|27|25|Фарсисские корабли были твоими караванами в твоей торговле, и ты сделался богатым и весьма славным среди морей.
EZEK|27|26|Гребцы твои завели тебя в большие воды; восточный ветер разбил тебя среди морей.
EZEK|27|27|Богатство твое и товары твои, все склады твои, корабельщики твои и кормчие твои, заделывавшие пробоины твои и распоряжавшиеся торговлею твоею, и все ратники твои, какие у тебя были, и все множество народа в тебе, в день падения твоего упадет в сердце морей.
EZEK|27|28|От вопля кормчих твоих содрогнутся окрестности.
EZEK|27|29|И с кораблей своих сойдут все гребцы, корабельщики, все кормчие моря, и станут на землю;
EZEK|27|30|и зарыдают о тебе громким голосом, и горько застенают, посыпав пеплом головы свои и валяясь во прахе;
EZEK|27|31|и остригут по тебе волосы догола, и опояшутся вретищами, и заплачут о тебе от душевной скорби горьким плачем;
EZEK|27|32|и в сетовании своем поднимут плачевную песнь о тебе, и так зарыдают о тебе: "кто как Тир, так разрушенный посреди моря!
EZEK|27|33|Когда приходили с морей товары твои, ты насыщал многие народы; множеством богатства твоего и торговлею твоею обогащал царей земли.
EZEK|27|34|А когда ты разбит морями в пучине вод, товары твои и все толпившееся в тебе упало.
EZEK|27|35|Все обитатели островов ужаснулись о тебе, и цари их содрогнулись, изменились в лицах.
EZEK|27|36|Торговцы других народов свистнули о тебе; ты сделался ужасом, – и не будет тебя во веки".
EZEK|28|1|И было ко мне слово Господне:
EZEK|28|2|сын человеческий! скажи начальствующему в Тире: так говорит Господь Бог: за то, что вознеслось сердце твое и ты говоришь: "я бог, восседаю на седалище божием, в сердце морей", и будучи человеком, а не Богом, ставишь ум твой наравне с умом Божиим, –
EZEK|28|3|вот, ты премудрее Даниила, нет тайны, сокрытой от тебя;
EZEK|28|4|твоею мудростью и твоим разумом ты приобрел себе богатство и в сокровищницы твои собрал золота и серебра;
EZEK|28|5|большою мудростью твоею, посредством торговли твоей, ты умножил богатство твое, и ум твой возгордился богатством твоим, –
EZEK|28|6|за то так говорит Господь Бог: так как ты ум твой ставишь наравне с умом Божиим,
EZEK|28|7|вот, Я приведу на тебя иноземцев, лютейших из народов, и они обнажат мечи свои против красы твоей мудрости и помрачат блеск твой;
EZEK|28|8|низведут тебя в могилу, и умрешь в сердце морей смертью убитых.
EZEK|28|9|Скажешь ли тогда перед твоим убийцею: "я бог", тогда как в руке поражающего тебя ты будешь человек, а не бог?
EZEK|28|10|Ты умрешь от руки иноземцев смертью необрезанных; ибо Я сказал это, говорит Господь Бог.
EZEK|28|11|И было ко мне слово Господне:
EZEK|28|12|сын человеческий! плачь о царе Тирском и скажи ему: так говорит Господь Бог: ты печать совершенства, полнота мудрости и венец красоты.
EZEK|28|13|Ты находился в Едеме, в саду Божием; твои одежды были украшены всякими драгоценными камнями; рубин, топаз и алмаз, хризолит, оникс, яспис, сапфир, карбункул и изумруд и золото, все, искусно усаженное у тебя в гнездышках и нанизанное на тебе, приготовлено было в день сотворения твоего.
EZEK|28|14|Ты был помазанным херувимом, чтобы осенять, и Я поставил тебя на то; ты был на святой горе Божией, ходил среди огнистых камней.
EZEK|28|15|Ты совершен был в путях твоих со дня сотворения твоего, доколе не нашлось в тебе беззакония.
EZEK|28|16|От обширности торговли твоей внутреннее твое исполнилось неправды, и ты согрешил; и Я низвергнул тебя, как нечистого, с горы Божией, изгнал тебя, херувим осеняющий, из среды огнистых камней.
EZEK|28|17|От красоты твоей возгордилось сердце твое, от тщеславия твоего ты погубил мудрость твою; за то Я повергну тебя на землю, перед царями отдам тебя на позор.
EZEK|28|18|Множеством беззаконий твоих в неправедной торговле твоей ты осквернил святилища твои; и Я извлеку из среды тебя огонь, который и пожрет тебя: и Я превращу тебя в пепел на земле перед глазами всех, видящих тебя.
EZEK|28|19|Все, знавшие тебя среди народов, изумятся о тебе; ты сделаешься ужасом, и не будет тебя во веки.
EZEK|28|20|И было ко мне слово Господне:
EZEK|28|21|сын человеческий! обрати лице твое к Сидону и изреки на него пророчество,
EZEK|28|22|и скажи: вот, Я – на тебя, Сидон, и прославлюсь среди тебя, и узнают, что Я Господь, когда произведу суд над ним и явлю в нем святость Мою;
EZEK|28|23|и пошлю на него моровую язву и кровопролитие на улицы его, и падут среди него убитые мечом, пожирающим его отовсюду; и узнают, что Я Господь.
EZEK|28|24|И не будет он впредь для дома Израилева колючим терном и причиняющим боль волчцом, более всех соседей зложелательствующим ему, и узнают, что Я Господь Бог.
EZEK|28|25|Так говорит Господь Бог: когда Я соберу дом Израилев из народов, между которыми они рассеяны, и явлю в них святость Мою перед глазами племен, и они будут жить на земле своей, которую Я дал рабу Моему Иакову:
EZEK|28|26|тогда они будут жить на ней безопасно, и построят домы, и насадят виноградники, и будут жить в безопасности, потому что Я произведу суд над всеми зложелателями их вокруг них, и узнают, что Я Господь Бог их.
EZEK|29|1|В десятом году, в десятом [месяце], в двенадцатый [день] месяца, было ко мне слово Господне:
EZEK|29|2|сын человеческий! обрати лице твое к фараону, царю Египетскому, и изреки пророчество на него и на весь Египет.
EZEK|29|3|Говори и скажи: так говорит Господь Бог: вот, Я – на тебя, фараон, царь Египетский, большой крокодил, который, лежа среди рек своих, говоришь: "моя река, и я создал ее для себя".
EZEK|29|4|Но Я вложу крюк в челюсти твои и к чешуе твоей прилеплю рыб из рек твоих, и вытащу тебя из рек твоих со всею рыбою рек твоих, прилипшею к чешуе твоей;
EZEK|29|5|и брошу тебя в пустыне, тебя и всю рыбу из рек твоих, ты упадешь на открытое поле, не уберут и не подберут тебя; отдам тебя на съедение зверям земным и птицам небесным.
EZEK|29|6|И узнают все обитатели Египта, что Я Господь; потому что они дому Израилеву были подпорою тростниковою.
EZEK|29|7|Когда они ухватились за тебя рукою, ты расщепился и все плечо исколол им; и когда они оперлись о тебя, ты сломился и изранил все чресла им.
EZEK|29|8|Посему так говорит Господь Бог: вот, Я наведу на тебя меч, и истреблю у тебя людей и скот.
EZEK|29|9|И сделается земля Египетская пустынею и степью; и узнают, что Я Господь. Так как он говорит: "моя река, и я создал ее";
EZEK|29|10|то вот, Я – на реки твои, и сделаю землю Египетскую пустынею из пустынь от Мигдола до Сиены, до самого предела Ефиопии.
EZEK|29|11|Не будет проходить по ней нога человеческая, и нога скотов не будет проходить по ней, и не будут обитать на ней сорок лет.
EZEK|29|12|И сделаю землю Египетскую пустынею среди земель опустошенных; и города ее среди опустелых городов будут пустыми сорок лет, и рассею Египтян по народам, и развею их по землям.
EZEK|29|13|Ибо так говорит Господь Бог: по окончании сорока лет Я соберу Египтян из народов, между которыми они будут рассеяны;
EZEK|29|14|и возвращу плен Египта, и обратно приведу их в землю Пафрос, в землю происхождения их, и там они будут царством слабым.
EZEK|29|15|Оно будет слабее [других] царств, и не будет более возноситься над народами; Я умалю их, чтобы они не господствовали над народами.
EZEK|29|16|И не будут впредь дому Израилеву опорою, припоминающею беззаконие их, когда они обращались к нему; и узнают, что Я Господь Бог.
EZEK|29|17|В двадцать седьмом году, в первом [месяце], в первый [день] месяца, было ко мне слово Господне:
EZEK|29|18|сын человеческий! Навуходоносор, царь Вавилонский, утомил свое войско большими работами при Тире; все головы оплешивели и все плечи стерты; а ни ему, ни войску его нет вознаграждения от Тира за работы, которые он употребил против него.
EZEK|29|19|Посему так говорит Господь Бог: вот, Я Навуходоносору, царю Вавилонскому, даю землю Египетскую, чтобы он обобрал богатство ее и произвел грабеж в ней, и ограбил награбленное ею, и это будет вознаграждением войску его.
EZEK|29|20|В награду за дело, которое он произвел в нем, Я отдаю ему землю Египетскую, потому что они делали это для Меня, сказал Господь Бог.
EZEK|29|21|В тот день возвращу рог дому Израилеву, и тебе открою уста среди них, и узнают, что Я Господь.
EZEK|30|1|И было ко мне слово Господне:
EZEK|30|2|сын человеческий! изреки пророчество и скажи: так говорит Господь Бог: рыдайте! о, злосчастный день!
EZEK|30|3|Ибо близок день, так! близок день Господа, день мрачный; година народов наступает.
EZEK|30|4|И пойдет меч на Египет, и ужас распространится в Ефиопии, когда в Египте будут падать пораженные, когда возьмут богатство его, и основания его будут разрушены;
EZEK|30|5|Ефиопия и Ливия, и Лидия, и весь смешанный народ, и Хуб, и сыны земли завета вместе с ними падут от меча.
EZEK|30|6|Так говорит Господь: падут подпоры Египта, и упадет гордыня могущества его; от Мигдола до Сиены будут падать в нем от меча, сказал Господь Бог.
EZEK|30|7|И опустеет он среди опустошенных земель, и города его будут среди опустошенных городов.
EZEK|30|8|И узнают, что Я Господь, когда пошлю огонь на Египет, и все подпоры его будут сокрушены.
EZEK|30|9|В тот день пойдут от Меня вестники на кораблях, чтобы устрашить беспечных Ефиоплян, и распространится у них ужас, как в день Египта; ибо вот, он идет.
EZEK|30|10|Так говорит Господь Бог: положу конец многолюдству Египта рукою Навуходоносора, царя Вавилонского.
EZEK|30|11|Он и с ним народ его, лютейший из народов, приведены будут на погибель сей земли, и обнажат мечи свои на Египет, и наполнят землю пораженными.
EZEK|30|12|И реки сделаю сушею и предам землю в руки злым, и рукою иноземцев опустошу землю и все, наполняющее ее. Я, Господь, сказал это.
EZEK|30|13|Так говорит Господь Бог: истреблю идолов и уничтожу лжебогов в Мемфисе, и из земли Египетской не будет уже властителя, и наведу страх на землю Египетскую.
EZEK|30|14|И опустошу Пафрос и пошлю огонь на Цоан, и произведу суд над Но.
EZEK|30|15|И изолью ярость Мою на Син, крепость Египта, и истреблю многолюдие в Но.
EZEK|30|16|И пошлю огонь на Египет; вострепещет Син, и Но рушится, и на Мемфис нападут враги среди дня.
EZEK|30|17|Молодые люди Она и Бубаста падут от меча, а прочие пойдут в плен.
EZEK|30|18|И в Тафнисе померкнет день, когда Я сокрушу там ярмо Египта, и прекратится в нем гордое могущество его. Облако закроет его, и дочери его пойдут в плен.
EZEK|30|19|Так произведу Я суд над Египтом, и узнают, что Я Господь.
EZEK|30|20|В одиннадцатом году, в первом месяце, в седьмой [день] месяца, было ко мне слово Господне:
EZEK|30|21|сын человеческий! Я уже сокрушил мышцу фараону, царю Египетскому; и вот, она еще не обвязана для излечения ее и не обвита врачебными перевязками, от которых она получила бы силу держать меч.
EZEK|30|22|Посему так говорит Господь Бог: вот, Я – на фараона, царя Египетского, и сокрушу мышцы его, здоровую и переломленную, так что меч выпадет из руки его.
EZEK|30|23|И рассею Египтян по народам, и развею их по землям.
EZEK|30|24|А мышцы царя Вавилонского сделаю крепкими и дам ему меч Мой в руку, мышцы же фараона сокрушу, и он изъязвленный будет сильно стонать перед ним.
EZEK|30|25|Укреплю мышцы царя Вавилонского, а мышцы у фараона опустятся; и узнают, что Я Господь, когда меч Мой дам в руку царю Вавилонскому, и он прострет его на землю Египетскую.
EZEK|30|26|И рассею Египтян по народам, и развею их по землям, и узнают, что Я Господь.
EZEK|31|1|В одиннадцатом году, в третьем [месяце], в первый день месяца, было ко мне слово Господне:
EZEK|31|2|сын человеческий! скажи фараону, царю Египетскому, и народу его: кому ты равняешь себя в величии твоем?
EZEK|31|3|Вот, Ассур был кедр на Ливане, с красивыми ветвями и тенистою листвою, и высокий ростом; вершина его находилась среди толстых сучьев.
EZEK|31|4|Воды растили его, бездна поднимала его, реки ее окружали питомник его, и она протоки свои посылала ко всем деревам полевым.
EZEK|31|5|От того высота его перевысила все дерева полевые, и сучьев на нем было много, и ветви его умножались, и сучья его становились длинными от множества вод, когда он разрастался.
EZEK|31|6|На сучьях его вили гнезда всякие птицы небесные, под ветвями его выводили детей всякие звери полевые, и под тенью его жили всякие многочисленные народы.
EZEK|31|7|Он красовался высотою роста своего, длиною ветвей своих, ибо корень его был у великих вод.
EZEK|31|8|Кедры в саду Божием не затемняли его; кипарисы не равнялись сучьям его, и каштаны не были величиною с ветви его, ни одно дерево в саду Божием не равнялось с ним красотою своею.
EZEK|31|9|Я украсил его множеством ветвей его, так что все дерева Едемские в саду Божием завидовали ему.
EZEK|31|10|Посему так сказал Господь Бог: за то, что ты высок стал ростом и вершину твою выставил среди толстых сучьев, и сердце его возгордилось величием его, –
EZEK|31|11|за то Я отдал его в руки властителю народов; он поступил с ним, как надобно; за беззаконие его Я отверг его.
EZEK|31|12|И срубили его чужеземцы, лютейшие из народов, и повергли его на горы; и на все долины упали ветви его; и сучья его сокрушились на всех лощинах земли, и из–под тени его ушли все народы земли, и оставили его.
EZEK|31|13|На обломках его поместились всякие птицы небесные, и в сучьях были всякие полевые звери.
EZEK|31|14|Это для того, чтобы никакие дерева при водах не величались высоким ростом своим и не поднимали вершины своей из среды толстых сучьев, и чтобы не прилеплялись к ним из–за высоты их дерева, пьющие воду; ибо все они будут преданы смерти, в преисподнюю страну вместе с сынами человеческими, отшедшими в могилу.
EZEK|31|15|Так говорит Господь Бог: в тот день, когда он сошел в могилу, Я сделал сетование о нем, затворил ради него бездну и остановил реки ее, и задержал большие воды и омрачил по нем Ливан, и все дерева полевые были в унынии по нем.
EZEK|31|16|Шумом падения его Я привел в трепет народы, когда низвел его в преисподнюю, к отшедшим в могилу, и обрадовались в преисподней стране все дерева Едема, отличные и наилучшие Ливанские, все, пьющие воду;
EZEK|31|17|ибо и они с ним отошли в преисподнюю, к пораженным мечом, и союзники его, жившие под тенью его, среди народов.
EZEK|31|18|Итак которому из дерев Едемских равнялся ты в славе и величии? Но теперь наравне с деревами Едемскими ты будешь низведен в преисподнюю, будешь лежать среди необрезанных, с пораженными мечом. Это фараон и все множество народа его, говорит Господь Бог.
EZEK|32|1|В двенадцатом году, в двенадцатом месяце, в первый [день] месяца, было ко мне слово Господне:
EZEK|32|2|сын человеческий! подними плач о фараоне, царе Египетском, и скажи ему: ты как молодой лев между народами и как чудовище в морях, кидаешься в реках твоих, и мутишь ногами твоими воды, и попираешь потоки их.
EZEK|32|3|Так говорит Господь Бог: Я закину на тебя сеть Мою в собрании многих народов, и они вытащат тебя Моею мрежею.
EZEK|32|4|И выкину тебя на землю, на открытом поле брошу тебя, и будут садиться на тебя всякие небесные птицы, и насыщаться тобою звери всей земли.
EZEK|32|5|И раскидаю мясо твое по горам, и долины наполню твоими трупами.
EZEK|32|6|И землю плавания твоего напою кровью твоею до самых гор; и рытвины будут наполнены тобою.
EZEK|32|7|И когда ты угаснешь, закрою небеса и звезды их помрачу, солнце закрою облаком, и луна не будет светить светом своим.
EZEK|32|8|Все светила, светящиеся на небе, помрачу над тобою и на землю твою наведу тьму, говорит Господь Бог.
EZEK|32|9|Приведу в смущение сердце многих народов, когда разглашу о падении твоем между народами, по землям, которых ты не знал.
EZEK|32|10|И приведу тобою в ужас многие народы, и цари их содрогнутся о тебе в страхе, когда мечом Моим потрясу перед лицем их, и поминутно будут трепетать каждый за душу свою в день падения твоего.
EZEK|32|11|Ибо так говорит Господь Бог: меч царя Вавилонского придет на тебя.
EZEK|32|12|От мечей сильных падет народ твой; все они – лютейшие из народов, и уничтожат гордость Египта, и погибнет все множество его.
EZEK|32|13|И истреблю весь скот его при великих водах, и вперед не будет мутить их нога человеческая, и копыта скота не будут мутить их.
EZEK|32|14|Тогда дам покой водам их, и сделаю, что реки их потекут, как масло, говорит Господь Бог.
EZEK|32|15|Когда сделаю землю Египетскую пустынею, и когда лишится земля всего, наполняющего ее; когда поражу всех живущих на ней, тогда узнают, что Я Господь.
EZEK|32|16|Вот плачевная песнь, которую будут петь; дочери народов будут петь ее; о Египте и обо всем множестве его будут петь ее, говорит Господь Бог.
EZEK|32|17|В двенадцатом году, в пятнадцатый [день того же] месяца, было ко мне слово Господне:
EZEK|32|18|сын человеческий! оплачь народ Египетский, и низринь его, его и дочерей знаменитых народов в преисподнюю, с отходящими в могилу.
EZEK|32|19|Кого ты превосходишь? сойди, и лежи с необрезанными.
EZEK|32|20|Те падут среди убитых мечом, и он отдан мечу; влеките его и все множество его.
EZEK|32|21|Среди преисподней будут говорить о нем и о союзниках его первые из героев; они пали и лежат там между необрезанными, сраженные мечом.
EZEK|32|22|Там Ассур и все полчище его, вокруг него гробы их, все пораженные, павшие от меча.
EZEK|32|23|Гробы его поставлены в самой глубине преисподней, и полчище его вокруг гробницы его, все пораженные, павшие от меча, те, которые распространяли ужас на земле живых.
EZEK|32|24|Так Елам со всем множеством своим вокруг гробницы его, все они пораженные, павшие от меча, которые необрезанными сошли в преисподнюю, которые распространили собою ужас на земле живых и несут позор свой с отшедшими в могилу.
EZEK|32|25|Среди пораженных дали ложе ему со всем множеством его; вокруг него гробы их, все необрезанные, пораженные мечом; и как они распространяли ужас на земле живых, то и несут на себе позор наравне с отшедшими в могилу и положены среди пораженных.
EZEK|32|26|Там Мешех и Фувал со всем множеством своим; вокруг него гробы их, все необрезанные, пораженные мечом, потому что они распространяли ужас на земле живых.
EZEK|32|27|Не должны ли [и] они лежать с павшими героями необрезанными, которые с воинским оружием своим сошли в преисподнюю и мечи свои положили себе под головы, и осталось беззаконие их на костях их, потому что они, как сильные, были ужасом на земле живых.
EZEK|32|28|И ты будешь сокрушен среди необрезанных и лежать с пораженными мечом.
EZEK|32|29|Там Едом и цари его и все князья его, которые при всей своей храбрости положены среди пораженных мечом; они лежат с необрезанными и сошедшими в могилу.
EZEK|32|30|Там властелины севера, все они и все Сидоняне, которые сошли туда с пораженными, быв посрамлены в могуществе своем, наводившем ужас, и лежат они с необрезанными, пораженными мечом, и несут позор свой с отшедшими в могилу.
EZEK|32|31|Увидит их фараон и утешится о всем множестве своем, пораженном мечом, фараон и все войско его, говорит Господь Бог.
EZEK|32|32|Ибо Я распространю страх Мой на земле живых, и положен будет фараон и все множество его среди необрезанных с пораженными мечом, говорит Господь Бог.
EZEK|33|1|И было ко мне слово Господне:
EZEK|33|2|сын человеческий! изреки слово к сынам народа твоего и скажи им: если Я на какую–либо землю наведу меч, и народ той земли возьмет из среды себя человека и поставит его у себя стражем;
EZEK|33|3|и он, увидев меч, идущий на землю, затрубит в трубу и предостережет народ;
EZEK|33|4|и если кто будет слушать голос трубы, но не остережет себя, – то, когда меч придет и захватит его, кровь его будет на его голове.
EZEK|33|5|Голос трубы он слышал, но не остерег себя, кровь его на нем будет; а кто остерегся, тот спас жизнь свою.
EZEK|33|6|Если же страж видел идущий меч и не затрубил в трубу, и народ не был предостережен, – то, когда придет меч и отнимет у кого из них жизнь, сей схвачен будет за грех свой, но кровь его взыщу от руки стража.
EZEK|33|7|И тебя, сын человеческий, Я поставил стражем дому Израилеву, и ты будешь слышать из уст Моих слово и вразумлять их от Меня.
EZEK|33|8|Когда Я скажу беззаконнику: "беззаконник! ты смертью умрешь", а ты не будешь ничего говорить, чтобы предостеречь беззаконника от пути его, – то беззаконник тот умрет за грех свой, но кровь его взыщу от руки твоей.
EZEK|33|9|Если же ты остерегал беззаконника от пути его, чтобы он обратился от него, но он от пути своего не обратился, – то он умирает за грех свой, а ты спас душу твою.
EZEK|33|10|И ты, сын человеческий, скажи дому Израилеву: вы говорите так: "преступления наши и грехи наши на нас, и мы истаеваем в них: как же можем мы жить?"
EZEK|33|11|Скажи им: живу Я, говорит Господь Бог: не хочу смерти грешника, но чтобы грешник обратился от пути своего и жив был. Обратитесь, обратитесь от злых путей ваших; для чего умирать вам, дом Израилев?
EZEK|33|12|И ты, сын человеческий, скажи сынам народа твоего: праведность праведника не спасет в день преступления его, и беззаконник за беззаконие свое не падет в день обращения от беззакония своего, равно как и праведник в день согрешения своего не может остаться в живых за свою праведность.
EZEK|33|13|Когда Я скажу праведнику, что он будет жив, а он понадеется на свою праведность и сделает неправду, – то все праведные дела его не помянутся, и он умрет от неправды своей, какую сделал.
EZEK|33|14|А когда скажу беззаконнику: "ты смертью умрешь", и он обратится от грехов своих и будет творить суд и правду,
EZEK|33|15|[если] этот беззаконник возвратит залог, за похищенное заплатит, будет ходить по законам жизни, не делая ничего худого, – то он будет жив, не умрет.
EZEK|33|16|Ни один из грехов его, какие он сделал, не помянется ему; он стал творить суд и правду, он будет жив.
EZEK|33|17|А сыны народа твоего говорят: "неправ путь Господа", тогда как их путь неправ.
EZEK|33|18|Когда праведник отступил от праведности своей и начал делать беззаконие, – то он умрет за то.
EZEK|33|19|И когда беззаконник обратился от беззакония своего и стал творить суд и правду, он будет за то жив.
EZEK|33|20|А вы говорите: "неправ путь Господа!" Я буду судить вас, дом Израилев, каждого по путям его.
EZEK|33|21|В двенадцатом году нашего переселения, в десятом [месяце], в пятый [день] месяца, пришел ко мне один из спасшихся из Иерусалима и сказал: "разрушен город!"
EZEK|33|22|Но еще до прихода сего спасшегося вечером была на мне рука Господа, и Он открыл мне уста, прежде нежели тот пришел ко мне поутру. И открылись уста мои, и я уже не был безмолвен.
EZEK|33|23|И было ко мне слово Господне:
EZEK|33|24|сын человеческий! живущие на опустелых местах в земле Израилевой говорят: "Авраам был один, и получил во владение землю сию, а нас много; [итак] нам дана земля сия во владение".
EZEK|33|25|Посему скажи им: так говорит Господь Бог: вы едите с кровью и поднимаете глаза ваши к идолам вашим, и проливаете кровь; и хотите владеть землею?
EZEK|33|26|Вы опираетесь на меч ваш, делаете мерзости, оскверняете один жену другого, и хотите владеть землею?
EZEK|33|27|Вот что скажи им: так говорит Господь Бог: живу Я! те, которые на местах разоренных, падут от меча; а кто в поле, того отдам зверям на съедение; а которые в укреплениях и пещерах, те умрут от моровой язвы.
EZEK|33|28|И сделаю землю пустынею из пустынь, и гордое могущество ее престанет, и горы Израилевы опустеют, так что не будет проходящих.
EZEK|33|29|И узнают, что Я Господь, когда сделаю землю пустынею из пустынь за все мерзости их, какие они делали.
EZEK|33|30|А о тебе, сын человеческий, сыны народа твоего разговаривают у стен и в дверях домов и говорят один другому, брат брату: "пойдите и послушайте, какое слово вышло от Господа".
EZEK|33|31|И они приходят к тебе, как на народное сходбище, и садится перед лицем твоим народ Мой, и слушают слова твои, но не исполняют их; ибо они в устах своих делают из этого забаву, сердце их увлекается за корыстью их.
EZEK|33|32|И вот, ты для них – как забавный певец с приятным голосом и хорошо играющий; они слушают слова твои, но не исполняют их.
EZEK|33|33|Но когда сбудется, – вот, уже и сбывается, – тогда узнают, что среди них был пророк.
EZEK|34|1|И было ко мне слово Господне:
EZEK|34|2|сын человеческий! изреки пророчество на пастырей Израилевых, изреки пророчество и скажи им, пастырям: так говорит Господь Бог: горе пастырям Израилевым, которые пасли себя самих! не стадо ли должны пасти пастыри?
EZEK|34|3|Вы ели тук и волною одевались, откормленных овец заколали, [а] стада не пасли.
EZEK|34|4|Слабых не укрепляли, и больной овцы не врачевали, и пораненной не перевязывали, и угнанной не возвращали, и потерянной не искали, а правили ими с насилием и жестокостью.
EZEK|34|5|И рассеялись они без пастыря и, рассеявшись, сделались пищею всякому зверю полевому.
EZEK|34|6|Блуждают овцы Мои по всем горам и по всякому высокому холму, и по всему лицу земли рассеялись овцы Мои, и никто не разведывает о них, и никто не ищет их.
EZEK|34|7|Посему, пастыри, выслушайте слово Господне.
EZEK|34|8|Живу Я! говорит Господь Бог; за то, что овцы Мои оставлены были на расхищение и без пастыря сделались овцы Мои пищею всякого зверя полевого, и пастыри Мои не искали овец Моих, и пасли пастыри самих себя, а овец Моих не пасли, –
EZEK|34|9|за то, пастыри, выслушайте слово Господне.
EZEK|34|10|Так говорит Господь Бог: вот, Я – на пастырей, и взыщу овец Моих от руки их, и не дам им более пасти овец, и не будут более пастыри пасти самих себя, и исторгну овец Моих из челюстей их, и не будут они пищею их.
EZEK|34|11|Ибо так говорит Господь Бог: вот, Я Сам отыщу овец Моих и осмотрю их.
EZEK|34|12|Как пастух поверяет стадо свое в тот день, когда находится среди стада своего рассеянного, так Я пересмотрю овец Моих и высвобожу их из всех мест, в которые они были рассеяны в день облачный и мрачный.
EZEK|34|13|И выведу их из народов, и соберу их из стран, и приведу их в землю их, и буду пасти их на горах Израилевых, при потоках и на всех обитаемых местах земли сей.
EZEK|34|14|Буду пасти их на хорошей пажити, и загон их будет на высоких горах Израилевых; там они будут отдыхать в хорошем загоне и будут пастись на тучной пажити, на горах Израилевых.
EZEK|34|15|Я буду пасти овец Моих и Я буду покоить их, говорит Господь Бог.
EZEK|34|16|Потерявшуюся отыщу и угнанную возвращу, и пораненную перевяжу, и больную укреплю, а разжиревшую и буйную истреблю; буду пасти их по правде.
EZEK|34|17|Вас же, овцы Мои, – так говорит Господь Бог, – вот, Я буду судить между овцою и овцою, между бараном и козлом.
EZEK|34|18|Разве мало вам того, что пасетесь на хорошей пажити, а между тем остальное на пажити вашей топчете ногами вашими, пьете чистую воду, а оставшуюся мутите ногами вашими,
EZEK|34|19|так что овцы Мои должны питаться тем, что потоптано ногами вашими, и пить то, что возмущено ногами вашими?
EZEK|34|20|Посему так говорит им Господь Бог: вот, Я Сам буду судить между овцою тучною и овцою тощею.
EZEK|34|21|Так как вы толкаете боком и плечом, и рогами своими бодаете всех слабых, доколе не вытолкаете их вон, –
EZEK|34|22|то Я спасу овец Моих, и они не будут уже расхищаемы, и рассужу между овцою и овцою.
EZEK|34|23|И поставлю над ними одного пастыря, который будет пасти их, раба Моего Давида; он будет пасти их и он будет у них пастырем.
EZEK|34|24|И Я, Господь, буду их Богом, и раб Мой Давид будет князем среди них. Я, Господь, сказал это.
EZEK|34|25|И заключу с ними завет мира и удалю с земли лютых зверей, так что безопасно будут жить в степи и спать в лесах.
EZEK|34|26|Дарую им и окрестностям холма Моего благословение, и дождь буду ниспосылать в свое время; это будут дожди благословения.
EZEK|34|27|И полевое дерево будет давать плод свой, и земля будет давать произведения свои; и будут они безопасны на земле своей, и узнают, что Я Господь, когда сокрушу связи ярма их и освобожу их из руки поработителей их.
EZEK|34|28|Они не будут уже добычею для народов, и полевые звери не будут пожирать их; они будут жить безопасно, и никто не будет устрашать [их].
EZEK|34|29|И произведу у них насаждение славное, и не будут уже погибать от голода на земле и терпеть посрамления от народов.
EZEK|34|30|И узнают, что Я, Господь Бог их, с ними, и они, дом Израилев, Мой народ, говорит Господь Бог,
EZEK|34|31|и что вы – овцы Мои, овцы паствы Моей; вы – человеки, [а] Я Бог ваш, говорит Господь Бог.
EZEK|35|1|И было ко мне слово Господне:
EZEK|35|2|сын человеческий! обрати лице твое к горе Сеир и изреки на нее пророчество
EZEK|35|3|и скажи ей: так говорит Господь Бог: вот, Я – на тебя, гора Сеир! и простру на тебя руку Мою и сделаю тебя пустою и необитаемою.
EZEK|35|4|Города твои превращу в развалины, и ты сама опустеешь и узнаешь, что Я Господь.
EZEK|35|5|Так как у тебя вечная вражда, и ты предавала сынов Израилевых в руки мечу во время несчастья их, во время окончательной гибели:
EZEK|35|6|за это – живу Я! говорит Господь Бог – сделаю тебя кровью, и кровь будет преследовать тебя; так как ты не ненавидела крови, то кровь и будет преследовать тебя.
EZEK|35|7|И сделаю гору Сеир пустою и безлюдною степью и истреблю на ней приходящего и возвращающегося.
EZEK|35|8|И наполню высоты ее убитыми ее; на холмах твоих и в долинах твоих, и во всех рытвинах твоих будут падать сраженные мечом.
EZEK|35|9|Сделаю тебя пустынею вечною, и в городах твоих не будут жить, и узнаете, что Я Господь.
EZEK|35|10|Так как ты говорила: "эти два народа и эти две земли будут мои, и мы завладеем ими, хотя и Господь был там":
EZEK|35|11|за то, – живу Я! говорит Господь Бог, – поступлю с тобою по мере ненависти твоей и зависти твоей, какую ты выказала из ненависти твоей к ним, и явлю Себя им, когда буду судить тебя.
EZEK|35|12|И узнаешь, что Я, Господь, слышал все глумления твои, какие ты произносила на горы Израилевы, говоря: "опустели! нам отданы на съедение!"
EZEK|35|13|Вы величались предо Мною языком вашим и умножали речи ваши против Меня; Я слышал это.
EZEK|35|14|Так говорит Господь Бог: когда вся земля будет радоваться, Я сделаю тебя пустынею.
EZEK|35|15|Как ты радовалась тому, что удел дома Израилева опустел, так сделаю Я и с тобою: опустошена будешь, гора Сеир, и вся Идумея вместе, и узнают, что Я Господь.
EZEK|36|1|И ты, сын человеческий, изреки пророчество на горы Израилевы и скажи: горы Израилевы! слушайте слово Господне.
EZEK|36|2|Так говорит Господь Бог: так как враг говорит о вас: "а! а! и вечные высоты достались нам в удел",
EZEK|36|3|то изреки пророчество и скажи: так говорит Господь Бог: за то, именно за то, что опустошают вас и поглощают вас со всех сторон, чтобы вы сделались достоянием прочих народов и подверглись злоречию и пересудам людей, –
EZEK|36|4|за это, горы Израилевы, выслушайте слово Господа Бога: так говорит Господь Бог горам и холмам, лощинам и долинам, и опустелым развалинам, и оставленным городам, которые сделались добычею и посмеянием прочим окрестным народам;
EZEK|36|5|за это так говорит Господь Бог: в огне ревности Моей Я изрек слово на прочие народы и на всю Идумею, которые назначили землю Мою во владение себе, с сердечною радостью и с презрением в душе обрекая ее в добычу себе.
EZEK|36|6|Посему изреки пророчество о земле Израилевой и скажи горам и холмам, лощинам и долинам: так говорит Господь Бог: вот, Я изрек сие в ревности Моей и в ярости Моей, потому что вы несете на себе посмеяние от народов.
EZEK|36|7|Посему так говорит Господь Бог: Я поднял руку Мою с клятвою, что народы, которые вокруг вас, сами понесут срам свой.
EZEK|36|8|А вы, горы Израилевы, распустите ветви ваши и будете приносить плоды ваши народу Моему Израилю; ибо они скоро придут.
EZEK|36|9|Ибо вот, Я к вам обращусь, и вы будете возделываемы и засеваемы.
EZEK|36|10|И поселю на вас множество людей, весь дом Израилев, весь, и заселены будут города и застроены развалины.
EZEK|36|11|И умножу на вас людей и скот, и они будут плодиться и размножаться, и заселю вас, как было в прежние времена ваши, и буду благотворить вам больше, нежели в прежние времена ваши, и узнаете, что Я Господь.
EZEK|36|12|И приведу на вас людей, народ Мой, Израиля, и они будут владеть тобою, [земля]! и ты будешь наследием их и не будешь более делать их бездетными.
EZEK|36|13|Так говорит Господь Бог: за то, что говорят о вас: "ты – [земля], поедающая людей и делающая народ твой бездетным":
EZEK|36|14|за то уже не будешь поедать людей и народа твоего не будешь вперед делать бездетным, говорит Господь Бог.
EZEK|36|15|И не будешь более слышать посмеяния от народов, и поругания от племен не понесешь уже на себе, и народа твоего вперед не будешь делать бездетным, говорит Господь Бог.
EZEK|36|16|И было ко мне слово Господне:
EZEK|36|17|сын человеческий! когда дом Израилев жил на земле своей, он осквернял ее поведением своим и делами своими; путь их пред лицем Моим был как нечистота женщины во время очищения ее.
EZEK|36|18|И Я излил на них гнев Мой за кровь, которую они проливали на этой земле, и за то, что они оскверняли ее идолами своими.
EZEK|36|19|И Я рассеял их по народам, и они развеяны по землям; Я судил их по путям их и по делам их.
EZEK|36|20|И пришли они к народам, куда пошли, и обесславили святое имя Мое, потому что о них говорят: "они – народ Господа, и вышли из земли Его".
EZEK|36|21|И пожалел Я святое имя Мое, которое обесславил дом Израилев у народов, куда пришел.
EZEK|36|22|Посему скажи дому Израилеву: так говорит Господь Бог: не для вас Я сделаю это, дом Израилев, а ради святаго имени Моего, которое вы обесславили у народов, куда пришли.
EZEK|36|23|И освящу великое имя Мое, бесславимое у народов, среди которых вы обесславили его, и узнают народы, что Я Господь, говорит Господь Бог, когда явлю на вас святость Мою перед глазами их.
EZEK|36|24|И возьму вас из народов, и соберу вас из всех стран, и приведу вас в землю вашу.
EZEK|36|25|И окроплю вас чистою водою, и вы очиститесь от всех скверн ваших, и от всех идолов ваших очищу вас.
EZEK|36|26|И дам вам сердце новое, и дух новый дам вам; и возьму из плоти вашей сердце каменное, и дам вам сердце плотяное.
EZEK|36|27|Вложу внутрь вас дух Мой и сделаю то, что вы будете ходить в заповедях Моих и уставы Мои будете соблюдать и выполнять.
EZEK|36|28|И будете жить на земле, которую Я дал отцам вашим, и будете Моим народом, и Я буду вашим Богом.
EZEK|36|29|И освобожу вас от всех нечистот ваших, и призову хлеб, и умножу его, и не дам вам терпеть голода.
EZEK|36|30|И умножу плоды на деревах и произведения полей, чтобы вперед не терпеть вам поношения от народов из–за голода.
EZEK|36|31|Тогда вспомните о злых путях ваших и недобрых делах ваших и почувствуете отвращение к самим себе за беззакония ваши и за мерзости ваши.
EZEK|36|32|Не ради вас Я сделаю это, говорит Господь Бог, да будет вам известно. Краснейте и стыдитесь путей ваших, дом Израилев.
EZEK|36|33|Так говорит Господь Бог: в тот день, когда очищу вас от всех беззаконий ваших и населю города, и обстроены будут развалины,
EZEK|36|34|и опустошенная земля будет возделываема, быв пустынею в глазах всякого мимоходящего,
EZEK|36|35|тогда скажут: "эта опустелая земля сделалась, как сад Едемский; и эти развалившиеся и опустелые и разоренные города укреплены и населены".
EZEK|36|36|И узнают народы, которые останутся вокруг вас, что Я, Господь, вновь созидаю разрушенное, засаждаю опустелое. Я, Господь, сказал – и сделал.
EZEK|36|37|Так говорит Господь Бог: вот, еще и в том явлю милость Мою дому Израилеву, умножу их людьми как стадо.
EZEK|36|38|Как много бывает жертвенных овец в Иерусалиме во время праздников его, так полны будут людьми опустелые города, и узнают, что Я Господь.
EZEK|37|1|Была на мне рука Господа, и Господь вывел меня духом и поставил меня среди поля, и оно было полно костей,
EZEK|37|2|и обвел меня кругом около них, и вот весьма много их на поверхности поля, и вот они весьма сухи.
EZEK|37|3|И сказал мне: сын человеческий! оживут ли кости сии? Я сказал: Господи Боже! Ты знаешь это.
EZEK|37|4|И сказал мне: изреки пророчество на кости сии и скажи им: "кости сухие! слушайте слово Господне!"
EZEK|37|5|Так говорит Господь Бог костям сим: вот, Я введу дух в вас, и оживете.
EZEK|37|6|И обложу вас жилами, и выращу на вас плоть, и покрою вас кожею, и введу в вас дух, и оживете, и узнаете, что Я Господь.
EZEK|37|7|Я изрек пророчество, как повелено было мне; и когда я пророчествовал, произошел шум, и вот движение, и стали сближаться кости, кость с костью своею.
EZEK|37|8|И видел я: и вот, жилы были на них, и плоть выросла, и кожа покрыла их сверху, а духа не было в них.
EZEK|37|9|Тогда сказал Он мне: изреки пророчество духу, изреки пророчество, сын человеческий, и скажи духу: так говорит Господь Бог: от четырех ветров приди, дух, и дохни на этих убитых, и они оживут.
EZEK|37|10|И я изрек пророчество, как Он повелел мне, и вошел в них дух, и они ожили, и стали на ноги свои – весьма, весьма великое полчище.
EZEK|37|11|И сказал Он мне: сын человеческий! кости сии – весь дом Израилев. Вот, они говорят: "иссохли кости наши, и погибла надежда наша, мы оторваны от корня".
EZEK|37|12|Посему изреки пророчество и скажи им: так говорит Господь Бог: вот, Я открою гробы ваши и выведу вас, народ Мой, из гробов ваших и введу вас в землю Израилеву.
EZEK|37|13|И узнаете, что Я Господь, когда открою гробы ваши и выведу вас, народ Мой, из гробов ваших,
EZEK|37|14|и вложу в вас дух Мой, и оживете, и помещу вас на земле вашей, и узнаете, что Я, Господь, сказал это – и сделал, говорит Господь.
EZEK|37|15|И было ко мне слово Господне:
EZEK|37|16|ты же, сын человеческий, возьми себе один жезл и напиши на нем: "Иуде и сынам Израилевым, союзным с ним"; и еще возьми жезл и напиши на нем: "Иосифу"; это жезл Ефрема и всего дома Израилева, союзного с ним.
EZEK|37|17|И сложи их у себя один с другим в один жезл, чтобы они в руке твоей были одно.
EZEK|37|18|И когда спросят у тебя сыны народа твоего: "не объяснишь ли нам, что это у тебя?",
EZEK|37|19|тогда скажи им: так говорит Господь Бог: вот, Я возьму жезл Иосифов, который в руке Ефрема и союзных с ним колен Израилевых, и приложу их к нему, к жезлу Иуды, и сделаю их одним жезлом, и будут одно в руке Моей.
EZEK|37|20|Когда же оба жезла, на которых ты напишешь, будут в руке твоей перед глазами их,
EZEK|37|21|то скажи им: так говорит Господь Бог: вот, Я возьму сынов Израилевых из среды народов, между которыми они находятся, и соберу их отовсюду и приведу их в землю их.
EZEK|37|22|На этой земле, на горах Израиля Я сделаю их одним народом, и один Царь будет царем у всех их, и не будут более двумя народами, и уже не будут вперед разделяться на два царства.
EZEK|37|23|И не будут уже осквернять себя идолами своими и мерзостями своими и всякими пороками своими, и освобожу их из всех мест жительства их, где они грешили, и очищу их, и будут Моим народом, и Я буду их Богом.
EZEK|37|24|А раб Мой Давид будет Царем над ними и Пастырем всех их, и они будут ходить в заповедях Моих, и уставы Мои будут соблюдать и выполнять их.
EZEK|37|25|И будут жить на земле, которую Я дал рабу Моему Иакову, на которой жили отцы их; там будут жить они и дети их, и дети детей их во веки; и раб Мой Давид будет князем у них вечно.
EZEK|37|26|И заключу с ними завет мира, завет вечный будет с ними. И устрою их, и размножу их, и поставлю среди них святилище Мое на веки.
EZEK|37|27|И будет у них жилище Мое, и буду их Богом, а они будут Моим народом.
EZEK|37|28|И узнают народы, что Я Господь, освящающий Израиля, когда святилище Мое будет среди них во веки.
EZEK|38|1|И было ко мне слово Господне:
EZEK|38|2|сын человеческий! обрати лице твое к Гогу в земле Магог, князю Роша, Мешеха и Фувала, и изреки на него пророчество
EZEK|38|3|и скажи: так говорит Господь Бог: вот, Я – на тебя, Гог, князь Роша, Мешеха и Фувала!
EZEK|38|4|И поверну тебя, и вложу удила в челюсти твои, и выведу тебя и все войско твое, коней и всадников, всех в полном вооружении, большое полчище, в бронях и со щитами, всех вооруженных мечами,
EZEK|38|5|Персов, Ефиоплян и Ливийцев с ними, всех со щитами и в шлемах,
EZEK|38|6|Гомера со всеми отрядами его, дом Фогарма, от пределов севера, со всеми отрядами его, многие народы с тобою.
EZEK|38|7|Готовься и снаряжайся, ты и все полчища твои, собравшиеся к тебе, и будь им вождем.
EZEK|38|8|После многих дней ты понадобишься; в последние годы ты придешь в землю, избавленную от меча, собранную из многих народов, на горы Израилевы, которые были в постоянном запустении, но теперь жители ее будут возвращены из народов, и все они будут жить безопасно.
EZEK|38|9|И поднимешься, как буря, пойдешь, как туча, чтобы покрыть землю, ты и все полчища твои и многие народы с тобою.
EZEK|38|10|Так говорит Господь Бог: в тот день придут тебе на сердце мысли, и ты задумаешь злое предприятие
EZEK|38|11|и скажешь: "поднимусь я на землю неогражденную, пойду на беззаботных, живущих беспечно, – все они живут без стен, и нет у них ни запоров, ни дверей, –
EZEK|38|12|чтобы произвести грабеж и набрать добычи, наложить руку на вновь заселенные развалины и на народ, собранный из народов, занимающийся хозяйством и торговлею, живущий на вершине земли".
EZEK|38|13|Сава и Дедан и купцы Фарсисские со всеми молодыми львами их скажут тебе: "ты пришел, чтобы произвести грабеж, собрал полчище твое, чтобы набрать добычи, взять серебро и золото, отнять скот и имущество, захватить большую добычу?"
EZEK|38|14|Посему изреки пророчество, сын человеческий, и скажи Гогу: так говорит Господь Бог: не так ли? в тот день, когда народ Мой Израиль будет жить безопасно, ты узнаешь это;
EZEK|38|15|и пойдешь с места твоего, от пределов севера, ты и многие народы с тобою, все сидящие на конях, сборище великое и войско многочисленное.
EZEK|38|16|И поднимешься на народ Мой, на Израиля, как туча, чтобы покрыть землю: это будет в последние дни, и Я приведу тебя на землю Мою, чтобы народы узнали Меня, когда Я над тобою, Гог, явлю святость Мою пред глазами их.
EZEK|38|17|Так говорит Господь Бог: не ты ли тот самый, о котором Я говорил в древние дни чрез рабов Моих, пророков Израилевых, которые пророчествовали в те времена, что Я приведу тебя на них?
EZEK|38|18|И будет в тот день, когда Гог придет на землю Израилеву, говорит Господь Бог, гнев Мой воспылает в ярости Моей.
EZEK|38|19|И в ревности Моей, в огне негодования Моего Я сказал: истинно в тот день произойдет великое потрясение на земле Израилевой.
EZEK|38|20|И вострепещут от лица Моего рыбы морские и птицы небесные, и звери полевые и все пресмыкающееся, ползающее по земле, и все люди, которые на лице земли, и обрушатся горы, и упадут утесы, и все стены падут на землю.
EZEK|38|21|И по всем горам Моим призову меч против него, говорит Господь Бог; меч каждого человека будет против брата его.
EZEK|38|22|И буду судиться с ним моровою язвою и кровопролитием, и пролью на него и на полки его и на многие народы, которые с ним, всепотопляющий дождь и каменный град, огонь и серу;
EZEK|38|23|и покажу Мое величие и святость Мою, и явлю Себя пред глазами многих народов, и узнают, что Я Господь.
EZEK|39|1|Ты же, сын человеческий, изреки пророчество на Гога и скажи: так говорит Господь Бог: вот, Я – на тебя, Гог, князь Роша, Мешеха и Фувала!
EZEK|39|2|И поверну тебя, и поведу тебя, и выведу тебя от краев севера, и приведу тебя на горы Израилевы.
EZEK|39|3|И выбью лук твой из левой руки твоей, и выброшу стрелы твои из правой руки твоей.
EZEK|39|4|Падешь ты на горах Израилевых, ты и все полки твои, и народы, которые с тобою; отдам тебя на съедение всякого рода хищным птицам и зверям полевым.
EZEK|39|5|На открытом поле падешь; ибо Я сказал это, говорит Господь Бог.
EZEK|39|6|И пошлю огонь на землю Магог и на жителей островов, живущих беспечно, и узнают, что Я Господь.
EZEK|39|7|И явлю святое имя Мое среди народа Моего, Израиля, и не дам вперед бесславить святаго имени Моего, и узнают народы, что Я Господь, Святый в Израиле.
EZEK|39|8|Вот, это придет и сбудется, говорит Господь Бог, – это тот день, о котором Я сказал.
EZEK|39|9|Тогда жители городов Израилевых выйдут, и разведут огонь, и будут сожигать оружие, щиты и латы, луки и стрелы, и булавы и копья; семь лет буду жечь их.
EZEK|39|10|И не будут носить дров с поля, ни рубить из лесов, но будут жечь только оружие; и ограбят грабителей своих, и оберут обирателей своих, говорит Господь Бог.
EZEK|39|11|И будет в тот день: дам Гогу место для могилы в Израиле, долину прохожих на восток от моря, и она будет задерживать прохожих; и похоронят там Гога и все полчище его, и будут называть ее долиною полчища Гогова.
EZEK|39|12|И дом Израилев семь месяцев будет хоронить их, чтобы очистить землю.
EZEK|39|13|И весь народ земли будет хоронить [их], и знаменит будет у них день, в который Я прославлю Себя, говорит Господь Бог.
EZEK|39|14|И назначат людей, которые постоянно обходили бы землю и с помощью прохожих погребали бы оставшихся на поверхности земли, для очищения ее; по прошествии семи месяцев они начнут делать поиски;
EZEK|39|15|и когда кто из обходящих землю увидит кость человеческую, то поставит возле нее знак, доколе погребатели не похоронят ее в долине полчища Гогова.
EZEK|39|16|И будет имя городу: Гамона. И так очистят они землю.
EZEK|39|17|Ты же, сын человеческий, так говорит Господь Бог, скажи всякого рода птицам и всем зверям полевым: собирайтесь и идите, со всех сторон сходитесь к жертве Моей, которую Я заколю для вас, к великой жертве на горах Израилевых; и будете есть мясо и пить кровь.
EZEK|39|18|Мясо мужей сильных будете есть, и будете пить кровь князей земли, баранов, ягнят, козлов и тельцов, всех откормленных на Васане;
EZEK|39|19|и будете есть жир до сытости и пить кровь до опьянения от жертвы Моей, которую Я заколю для вас.
EZEK|39|20|И насытитесь за столом Моим конями и всадниками, мужами сильными и всякими людьми военными, говорит Господь Бог.
EZEK|39|21|И явлю славу Мою между народами, и все народы увидят суд Мой, который Я произведу, и руку Мою, которую Я наложу на них.
EZEK|39|22|И будет знать дом Израилев, что Я Господь Бог их, от сего дня и далее.
EZEK|39|23|И узнают народы, что дом Израилев был переселен за неправду свою; за то, что они поступали вероломно предо Мною, Я сокрыл от них лице Мое и отдал их в руки врагов их, и все они пали от меча.
EZEK|39|24|За нечистоты их и за их беззаконие Я сделал это с ними, и сокрыл от них лице Мое.
EZEK|39|25|Посему так говорит Господь Бог: ныне возвращу плен Иакова, и помилую весь дом Израиля, и возревную по святом имени Моем.
EZEK|39|26|И почувствуют они бесчестие свое и все беззакония свои, какие делали предо Мною, когда будут жить на земле своей безопасно, и никто не будет устрашать их,
EZEK|39|27|когда Я возвращу их из народов, и соберу их из земель врагов их, и явлю в них святость Мою пред глазами многих народов.
EZEK|39|28|И узнают, что Я Господь Бог их, когда, рассеяв их между народами, опять соберу их в землю их и не оставлю уже там ни одного из них;
EZEK|39|29|и не буду уже скрывать от них лица Моего, потому что Я изолью дух Мой на дом Израилев, говорит Господь Бог.
EZEK|40|1|В двадцать пятом году по переселении нашем, в начале года, в десятый [день] месяца, в четырнадцатом году по разрушении города, в тот самый день была на мне рука Господа, и Он повел меня туда.
EZEK|40|2|В видениях Божиих привел Он меня в землю Израилеву и поставил меня на весьма высокой горе, и на ней, с южной стороны, были как бы городские здания;
EZEK|40|3|и привел меня туда. И вот муж, которого вид как бы вид блестящей меди, и льняная вервь в руке его и трость измерения, и стоял он у ворот.
EZEK|40|4|И сказал мне этот муж: "сын человеческий! смотри глазами твоими и слушай ушами твоими, и прилагай сердце твое ко всему, что я буду показывать тебе, ибо ты для того и приведен сюда, чтоб я показал тебе [это]; все, что увидишь, возвести дому Израилеву".
EZEK|40|5|И вот, вне храма стена со всех сторон [его], и в руке того мужа трость измерения в шесть локтей, [считая каждый локоть] в локоть с ладонью; и намерил он в этом здании одну трость толщины и одну трость вышины.
EZEK|40|6|Потом пошел к воротам, обращенным лицом к востоку, и взошел по ступеням их, и нашел меры в одном пороге ворот одну трость ширины и в другом пороге одну трость ширины.
EZEK|40|7|И в каждой боковой комнате одна трость длины и одна трость ширины, а между комнатами пять локтей, и в пороге ворот у притвора ворот внутри одна же трость.
EZEK|40|8|И смерил он в притворе ворот внутри одну трость,
EZEK|40|9|а в притворе у ворот намерил восемь локтей и два локтя в столбах. Этот притвор у ворот со стороны храма.
EZEK|40|10|Боковых комнат у восточных ворот три – с одной стороны и три – с другой; одна мера во всех трех и одна мера в столбах с той и другой стороны.
EZEK|40|11|Ширины в отверстии ворот он намерил десять локтей, а длины ворот тринадцать локтей.
EZEK|40|12|А перед комнатами выступ в один локоть, и в один же локоть с другой стороны выступ; эти комнаты с одной стороны [имели] шесть локтей и шесть же локтей с другой стороны.
EZEK|40|13|Потом намерил он в воротах от крыши одной комнаты до крыши другой двадцать пять локтей ширины; дверь была против двери.
EZEK|40|14|А в столбах он насчитал шестьдесят локтей, в каждом столбе около двора и у ворот,
EZEK|40|15|и от передней стороны входа в ворота до передней стороны внутренних ворот пятьдесят локтей.
EZEK|40|16|Решетчатые окна были и в боковых комнатах и в столбах их, внутрь ворот кругом, также и в притворах окна были кругом на внутреннюю сторону, и на столбах – пальмы.
EZEK|40|17|И привел он меня на внешний двор, и вот там комнаты, и каменный помост кругом двора был сделан; тридцать комнат на том помосте.
EZEK|40|18|И помост этот был по бокам ворот, соответственно длине ворот; этот помост был ниже.
EZEK|40|19|И намерил он в ширину от нижних ворот до внешнего края внутреннего двора сто локтей, к востоку и к северу.
EZEK|40|20|Он измерил также длину и ширину ворот внешнего двора, обращенных лицом к северу,
EZEK|40|21|и боковые комнаты при них, три с одной стороны и три с другой; и столбы их, и выступы их были такой же меры, как у прежних ворот: длина их пятьдесят локтей, а ширина двадцать пять локтей.
EZEK|40|22|И окна их, и выступы их, и пальмы их – той же меры, как у ворот, обращенных лицом к востоку; и входят к ним семью ступенями, и перед ними выступы.
EZEK|40|23|И во внутренний двор есть ворота против ворот северных и восточных; и намерил он от ворот до ворот сто локтей.
EZEK|40|24|И повел меня на юг, и вот там ворота южные; и намерил он в столбах и выступах такую же меру.
EZEK|40|25|И окна в них и в преддвериях их такие же, как те окна: длина пятьдесят локтей, а ширины двадцать пять локтей.
EZEK|40|26|Подъем к ним – в семь ступеней, и преддверия перед ними; и пальмовые украшения – одно с той стороны и одно с другой на столбах их.
EZEK|40|27|И во внутренний двор были южные ворота; и намерил он от ворот до ворот южных сто локтей.
EZEK|40|28|И привел он меня через южные ворота во внутренний двор; и намерил в южных воротах ту же меру.
EZEK|40|29|И боковые комнаты их, и столбы их, и притворы их – той же меры, и окна в них в притворах их были кругом; всего в длину пятьдесят локтей, а в ширину двадцать пять локтей.
EZEK|40|30|Притворы были кругом длиною в двадцать пять локтей, а шириною в пять локтей.
EZEK|40|31|И притворы были у них на внешний двор, и пальмы были на столбах их; подъем к ним – в восемь ступеней.
EZEK|40|32|И повел меня восточными воротами на внутренний двор; и намерил в этих воротах ту же меру.
EZEK|40|33|И боковые комнаты их, и столбы их, и притворы их были той же меры; и окна в них и притворах их были кругом; длина пятьдесят локтей, а ширина двадцать пять локтей.
EZEK|40|34|Притворы у них были на внешний двор, и пальмы на столбах их с той и другой стороны; подъем к ним – в восемь ступеней.
EZEK|40|35|Потом привел меня к северным воротам, и намерил в них ту же меру.
EZEK|40|36|Боковые комнаты при них, столбы их и притворы их, и окна в них были кругом; всего в длину пятьдесят локтей, и в ширину двадцать пять локтей.
EZEK|40|37|Притворы у них были на внешний двор, и пальмы на столбах их с той и с другой стороны; подъем к ним – в восемь ступеней.
EZEK|40|38|Была также комната, со входом в нее, у столбов ворот: там омывают жертвы всесожжения.
EZEK|40|39|А в притворе у ворот два стола с одной стороны и два с другой стороны, чтобы заколать на них жертвы всесожжения и жертвы за грех и жертвы за преступление.
EZEK|40|40|И у наружного бока при входе в отверстие северных ворот были два стола, и у другого бока, подле притвора у ворот, два стола.
EZEK|40|41|Четыре стола с одной стороны и четыре стола с другой стороны, по бокам ворот: [всего] восемь столов, на которых заколают [жертвы].
EZEK|40|42|И четыре стола для приготовления всесожжения были из тесаных камней, длиною в полтора локтя, и шириною в полтора локтя, а вышиною в один локоть; на них кладут орудия для заклания жертвы всесожжения и [других] жертв.
EZEK|40|43|И крюки в одну ладонь приделаны были к стенам здания кругом, а на столах клали жертвенное мясо.
EZEK|40|44|Снаружи внутренних ворот были комнаты для певцов; на внутреннем дворе, сбоку северных ворот, одна обращена лицом к югу, а другая, сбоку южных ворот, обращена лицом к северу.
EZEK|40|45|И сказал он мне: "эта комната, которая лицом к югу, для священников, бодрствующих на страже храма;
EZEK|40|46|а комната, которая лицом к северу, для священников, бодрствующих на страже жертвенника: это сыны Садока, которые одни из сынов Левия приближаются к Господу, чтобы служить Ему".
EZEK|40|47|И намерил он во дворе сто локтей длины и сто локтей ширины: [он] был четыреугольный; а перед храмом стоял жертвенник.
EZEK|40|48|И привел он меня к притвору храма, и намерил в столбах притвора пять локтей с одной стороны и пять локтей с другой; а в воротах три локтя ширины с одной стороны и три локтя с другой.
EZEK|40|49|Длина притвора – в двадцать локтей, а ширина – в одиннадцать локтей, и всходят в него по десяти ступеням; и были подпоры у столбов, одна с одной стороны, а другая с другой.
EZEK|41|1|Потом ввел меня в храм и намерил в столбах шесть локтей ширины с одной стороны и шесть локтей ширины с другой стороны, в ширину скинии.
EZEK|41|2|В дверях десять локтей ширины, и по бокам дверей пять локтей с одной стороны и пять локтей с другой стороны; и намерил длины в храме сорок локтей, а ширины двадцать локтей.
EZEK|41|3|И пошел внутрь, и намерил в столбах у дверей два локтя и в дверях шесть локтей, а ширина двери – в семь локтей.
EZEK|41|4|И отмерил в нем двадцать локтей в длину и двадцать локтей в ширину храма, и сказал мне: "это – Святое Святых".
EZEK|41|5|И намерил в стене храма шесть локтей, а ширины в боковых комнатах, кругом храма, по четыре локтя.
EZEK|41|6|Боковых комнат было тридцать три, комната подле комнаты; они вдаются в стену, которая у храма для комнат кругом, так что они в связи с нею, но стены самого храма не касаются.
EZEK|41|7|И он более и более расширялся кругом вверх боковыми комнатами, потому что окружность храма восходила выше и выше вокруг храма, и потому храм имел большую ширину вверху, и из нижнего этажа восходили в верхний через средний.
EZEK|41|8|И я видел верх дома во всю окружность; боковые комнаты в основании имели там меры цельную трость, шесть полных локтей.
EZEK|41|9|Ширина стены боковых комнат, выходящих наружу, пять локтей, и открытое пространство есть подле боковых комнат храма.
EZEK|41|10|И между комнатами расстояние двадцать локтей кругом всего храма.
EZEK|41|11|Двери боковых комнат [ведут] на открытое пространство, одни двери – на северную сторону, а другие двери – на южную сторону; а ширина этого открытого пространства – пять локтей кругом.
EZEK|41|12|Здание перед площадью на западной стороне – шириною в семьдесят локтей; стена же этого здания – в пять локтей ширины кругом, а длина ее – девяносто локтей.
EZEK|41|13|И намерил он в храме сто локтей длины, и в площади и в пристройке, и в стенах его также сто локтей длины.
EZEK|41|14|И ширина храма по лицевой стороне и площади к востоку сто же локтей.
EZEK|41|15|И в длине здания перед площадью на задней стороне ее с боковыми комнатами его по ту и другую сторону он намерил сто локтей, со внутренностью храма и притворами двора.
EZEK|41|16|Дверные брусья и решетчатые окна, и боковые комнаты кругом, во всех трех [ярусах], против порогов обшиты деревом и от пола по окна; окна были закрыты.
EZEK|41|17|От верха дверей как внутри храма, так и снаружи, и по всей стене кругом, внутри и снаружи, были резные изображения,
EZEK|41|18|сделаны были херувимы и пальмы: пальма между двумя херувимами, и у каждого херувима два лица.
EZEK|41|19|С одной стороны к пальме обращено лицо человеческое, а с другой стороны к пальме – лице львиное; так сделано во всем храме кругом.
EZEK|41|20|От пола до верха дверей сделаны были херувимы и пальмы, также и по стене храма.
EZEK|41|21|В храме были четырехугольные дверные косяки, и святилище имело такой же вид, как я видел.
EZEK|41|22|Жертвенник был деревянный в три локтя вышины и в два локтя длины; и углы его, и подножие его, и стенки его – из дерева. И сказал он мне: "это трапеза, которая пред Господом".
EZEK|41|23|В храме и во святилище по две двери,
EZEK|41|24|и двери сии о двух досках, обе доски подвижные, две у одной двери и две доски у другой;
EZEK|41|25|и сделаны на них, на дверях храма, херувимы и пальмы такие же, какие сделаны по стенам; а перед притвором снаружи был деревянный помост.
EZEK|41|26|И решетчатые окна с пальмами, по ту и другую сторону, были по бокам притвора и в боковых комнатах храма и на деревянной обшивке.
EZEK|42|1|И вывел меня ко внешнему двору северною дорогою, и привел меня к комнатам, которые против площади и против здания на севере,
EZEK|42|2|к тому месту, которое у северных дверей имеет в длину сто локтей, а в ширину пятьдесят локтей.
EZEK|42|3|Напротив двадцати [локтей] внутреннего двора и напротив помоста, который на внешнем дворе, были галерея против галереи в три яруса.
EZEK|42|4|А перед комнатами ход в десять локтей ширины, а внутрь в один локоть; двери их лицом к северу.
EZEK|42|5|Верхние комнаты уже, потому что галереи отнимают у них несколько против нижних и средних [комнат] этого здания.
EZEK|42|6|Они в три яруса, и таких столбов, какие на дворах, нет у них; потому они и сделаны уже против нижних и средних комнат, начиная от пола.
EZEK|42|7|А наружная стена напротив этих комнат от внешнего двора, составляющая лицевую сторону комнат, имеет длины пятьдесят локтей;
EZEK|42|8|потому что [и] комнаты на внешнем дворе занимают длины только пятьдесят локтей, и вот перед храмом сто локтей.
EZEK|42|9|А снизу ход к этим комнатам с восточной стороны, когда подходят к ним со внешнего двора.
EZEK|42|10|В ширину стены двора к востоку перед площадью и перед зданием были комнаты.
EZEK|42|11|И ход перед ними такой же, как и у тех комнат, которые обращены к северу, такая же длина, как и у тех, и такая же ширина, и все выходы их, и устройство их, и двери их такие же, как и у тех.
EZEK|42|12|Такие же двери, как и у комнат, которые на юг, и для входа в них дверь у самой дороги, которая шла прямо вдоль стены на восток.
EZEK|42|13|И сказал он мне: "комнаты на север [и] комнаты на юг, которые перед площадью, суть комнаты священные, в которых священники, приближающиеся к Господу, съедают священнейшие жертвы; там же они кладут священнейшие жертвы, и хлебное приношение, и жертву за грех, и жертву за преступление, ибо это место святое.
EZEK|42|14|Когда войдут [туда] священники, то они не должны выходить из этого святаго места на внешний двор, доколе не оставят там одежд своих, в которых служили, ибо они священны; они должны надеть на себя другие одежды и тогда выходить к народу".
EZEK|42|15|Когда кончил он измерения внутреннего храма, то вывел меня воротами, обращенными лицом к востоку, и стал измерять его кругом.
EZEK|42|16|Он измерил восточную сторону тростью измерения и [намерил] тростью измерения всего пятьсот тростей;
EZEK|42|17|в северной стороне той же тростью измерения намерил всего пятьсот тростей;
EZEK|42|18|в южной стороне намерил тростью измерения также пятьсот тростей.
EZEK|42|19|Поворотив к западной стороне, намерил тростью измерения пятьсот тростей.
EZEK|42|20|Со всех четырех сторон он измерил его; кругом него была стена длиною в пятьсот [тростей] и в пятьсот [тростей] шириною, чтобы отделить святое место от несвятого.
EZEK|43|1|И привел меня к воротам, к тем воротам, которые обращены лицом к востоку.
EZEK|43|2|И вот, слава Бога Израилева шла от востока, и глас Его – как шум вод многих, и земля осветилась от славы Его.
EZEK|43|3|Это видение было такое же, какое я видел прежде, точно такое, какое я видел, когда приходил возвестить гибель городу, и видения, подобные видениям, какие видел я у реки Ховара. И я пал на лице мое.
EZEK|43|4|И слава Господа вошла в храм путем ворот, обращенных лицом к востоку.
EZEK|43|5|И поднял меня дух, и ввел меня во внутренний двор, и вот, слава Господа наполнила весь храм.
EZEK|43|6|И я слышал кого–то, говорящего мне из храма, а тот муж стоял подле меня,
EZEK|43|7|и сказал мне: сын человеческий! это место престола Моего и место стопам ног Моих, где Я буду жить среди сынов Израилевых во веки; и дом Израилев не будет более осквернять святаго имени Моего, ни они, ни цари их, блужением своим и трупами царей своих на высотах их.
EZEK|43|8|Они ставили порог свой у порога Моего и вереи дверей своих подле Моих верей, так что одна стена [была] между Мною и ими, и оскверняли святое имя Мое мерзостями своими, какие делали, и за то Я погубил их во гневе Моем.
EZEK|43|9|А теперь они удалят от Меня блужение свое и трупы царей своих, и Я буду жить среди них во веки.
EZEK|43|10|Ты, сын человеческий, возвести дому Израилеву о храме сем, чтобы они устыдились беззаконий своих и чтобы сняли с него меру.
EZEK|43|11|И если они устыдятся всего того, что делали, то покажи им вид храма и расположение его, и выходы его, и входы его, и все очертания его, и все уставы его, и все образы его, и все законы его, и напиши при глазах их, чтобы они сохраняли все очертания его и все уставы его и поступали по ним.
EZEK|43|12|Вот закон храма: на вершине горы все пространство его вокруг – Святое Святых; вот закон храма!
EZEK|43|13|И вот размеры жертвенника локтями, [считая] локоть в локоть с ладонью: основание в локоть, ширина в локоть же, и пояс по всем краям его в одну пядень; и вот задняя сторона жертвенника.
EZEK|43|14|От основания, что в земле, до нижнего выступа два локтя, а шириною он в один локоть; от малого выступа до большого выступа четыре локтя, а ширина его – в один локоть.
EZEK|43|15|Самый жертвенник вышиною в четыре локтя; и из жертвенника [поднимаются] вверх четыре рога.
EZEK|43|16|Жертвенник имеет двенадцать [локтей] длины [и] двенадцать ширины; он четырехугольный на все свои четыре стороны.
EZEK|43|17|А в площадке четырнадцать [локтей] длины и четырнадцать ширины на все четыре стороны ее, и вокруг нее пояс в пол–локтя, а основание ее в локоть вокруг, ступени же к нему – с востока.
EZEK|43|18|И сказал он мне: сын человеческий! так говорит Господь Бог: вот уставы жертвенника к тому дню, когда он будет сделан для приношения на нем всесожжений и для кропления на него кровью.
EZEK|43|19|Священникам от колена Левиина, которые из племени Садока, приближающимся ко Мне, чтобы служить Мне, говорит Господь Бог, дай тельца из стада волов, в жертву за грех.
EZEK|43|20|И возьми крови его, и покропи на четыре рога его, и на четыре угла площадки, и на пояс кругом, и так очисти его и освяти его.
EZEK|43|21|И возьми тельца, [в жертву] за грех, и сожги его на назначенном месте дома вне святилища.
EZEK|43|22|А на другой день в жертву за грех принеси из козьего стада козла без порока, и пусть очистят жертвенник так же, как очищали тельцом.
EZEK|43|23|Когда же кончишь очищение, приведи из стада волов тельца без порока и из стада овец овна без порока;
EZEK|43|24|и принеси их пред лице Господа; и священники бросят на них соли, и вознесут их во всесожжение Господу.
EZEK|43|25|Семь дней приноси в жертву за грех по козлу в день; также пусть приносят в жертву по тельцу из стада волов и по овну из стада овец без порока.
EZEK|43|26|Семь дней они должны очищать жертвенник и освящать его и наполнять руки свои.
EZEK|43|27|По окончании же сих дней, в восьмой день и далее, священники будут возносить на жертвеннике ваши всесожжения и благодарственные жертвы; и Я буду милостив к вам, говорит Господь Бог.
EZEK|44|1|И привел он меня обратно ко внешним воротам святилища, обращенным лицом на восток, и они были затворены.
EZEK|44|2|И сказал мне Господь: ворота сии будут затворены, не отворятся, и никакой человек не войдет ими, ибо Господь, Бог Израилев, вошел ими, и они будут затворены.
EZEK|44|3|Что до князя, он, [как] князь, сядет в них, чтобы есть хлеб пред Господом; войдет путем притвора этих ворот, и тем же путем выйдет.
EZEK|44|4|Потом привел меня путем ворот северных перед лице храма, и я видел, и вот, слава Господа наполняла дом Господа, и пал я на лице мое.
EZEK|44|5|И сказал мне Господь: сын человеческий! прилагай сердце твое [ко] [всему], и смотри глазами твоими, и слушай ушами твоими все, что Я говорю тебе о всех постановлениях дома Господа и всех законах его; и прилагай сердце твое ко входу в храм и ко всем выходам из святилища.
EZEK|44|6|И скажи мятежному дому Израилеву: так говорит Господь Бог: довольно вам, дом Израилев, делать все мерзости ваши,
EZEK|44|7|вводить сынов чужой, необрезанных сердцем и необрезанных плотью, чтобы они были в Моем святилище и оскверняли храм Мой, подносить хлеб Мой, тук и кровь, и разрушать завет Мой всякими мерзостями вашими.
EZEK|44|8|Вы не исполняли стражи у святынь Моих, а ставили вместо себя их для стражи в Моем святилище.
EZEK|44|9|Так говорит Господь Бог: никакой сын чужой, необрезанный сердцем и необрезанный плотью, не должен входить во святилище Мое, даже и тот сын чужой, который [живет] среди сынов Израиля.
EZEK|44|10|Равно и левиты, которые удалились от Меня во время отступничества Израилева, которые, оставив Меня, блуждали вслед идолов своих, понесут наказание за вину свою.
EZEK|44|11|Они будут служить во святилище Моем, как сторожа у ворот храма и прислужники у храма; они будут заколать для народа всесожжение и другие жертвы, и будут стоять пред ними для служения им.
EZEK|44|12|За то, что они служили им пред идолами их и были для дома Израилева соблазном к нечестию, Я поднял на них руку Мою, говорит Господь Бог, и они понесут наказание за вину свою;
EZEK|44|13|они не будут приближаться ко Мне, чтобы священнодействовать предо Мною и приступать ко всем святыням Моим, к Святому Святых, но будут нести на себе бесславие свое и мерзости свои, какие делали.
EZEK|44|14|Сделаю их стражами храма для всех служб его и для всего, что производится в нем.
EZEK|44|15|А священники из колена Левиина, сыны Садока, которые, во время отступления сынов Израилевых от Меня, постоянно стояли на страже святилища Моего, те будут приближаться ко Мне, чтобы служить Мне, и будут предстоять пред лицем Моим, чтобы приносить Мне тук и кровь, говорит Господь Бог.
EZEK|44|16|Они будут входить во святилище Мое и приближаться к трапезе Моей, чтобы служить Мне и соблюдать стражу Мою.
EZEK|44|17|Когда придут к воротам внутреннего двора, тогда оденутся в одежды льняные, а шерстяное не должно быть на них во время служения их в воротах внутреннего двора и внутри храма.
EZEK|44|18|Увясла на головах их должны быть также льняные; и исподняя одежда на чреслах их должна быть также льняная; в поту они не должны опоясываться.
EZEK|44|19|А когда надобно будет выйти на внешний двор, на внешний двор к народу, тогда они должны будут снять одежды свои, в которых они служили, и оставить их в священных комнатах, и одеться в другие одежды, чтобы священными одеждами своими не прикасаться к народу.
EZEK|44|20|И головы своей они не должны брить, и не должны отпускать волос, а пусть непременно стригут головы свои.
EZEK|44|21|И вина не должен пить ни один священник, когда идет во внутренний двор.
EZEK|44|22|Ни вдовы, ни разведенной с мужем они не должны брать себе в жены, а только могут брать себе девиц из племени дома Израилева и вдову, оставшуюся вдовою от священника.
EZEK|44|23|Они должны учить народ Мой отличать священное от несвященного и объяснять им, что нечисто и что чисто.
EZEK|44|24|При спорных делах они должны присутствовать в суде, и по уставам Моим судить их, и наблюдать законы Мои и постановления Мои о всех праздниках Моих, и свято хранить субботы Мои.
EZEK|44|25|К мертвому человеку никто из них не должен подходить, чтобы не сделаться нечистым; только ради отца и матери, ради сына и дочери, брата и сестры, которая не была замужем, можно им сделать себя нечистыми.
EZEK|44|26|По очищении же такого, еще семь дней надлежит отсчитать ему.
EZEK|44|27|И в тот день, когда ему надобно будет приступать ко святыне во внутреннем дворе, чтобы служить при святыне, он должен принести жертву за грех, говорит Господь Бог.
EZEK|44|28|А что до удела их, то Я их удел. И владения не давайте им в Израиле: Я их владение.
EZEK|44|29|Они будут есть от хлебного приношения, от жертвы за грех и жертвы за преступление; и все заклятое у Израиля им же принадлежит.
EZEK|44|30|И начатки из всех плодов ваших и всякого рода приношения, из чего ни состояли бы приношения ваши, принадлежат священникам; и начатки молотого вами отдавайте священнику, чтобы над домом твоим почивало благословение.
EZEK|44|31|Никакой мертвечины и ничего, растерзанного зверем, ни из птиц, ни из скота, не должны есть священники.
EZEK|45|1|Когда будете по жребию делить землю на уделы, тогда отделите священный участок Господу в двадцать пять тысяч [тростей] длины и десять тысяч ширины; да будет свято это место во всем объеме своем, кругом.
EZEK|45|2|От него к святилищу отойдет четырехугольник по пятисот [тростей] кругом, и кругом него площадь в пятьдесят локтей.
EZEK|45|3|Из этой меры отмерь двадцать пять тысяч [тростей] в длину и десять тысяч в ширину, где будет находиться святилище, Святое Святых.
EZEK|45|4|Эта священная часть земли принадлежать будет священникам, служителям святилища, приступающим к служению Господу: это будет для них местом для домов и святынею для святилища.
EZEK|45|5|Двадцать пять тысяч [тростей] длины и десять тысяч ширины будут принадлежать левитам, служителям храма, как их владение для обитания их.
EZEK|45|6|И во владение городу дайте пять тысяч ширины и двадцать пять тысяч длины, против священного места, отделенного Господу; это принадлежать должно всему дому Израилеву.
EZEK|45|7|И князю [дайте] долю по ту и другую сторону, как подле священного места, отделенного [Господу], так и подле городского владения, к западу с западной стороны и к востоку с восточной стороны, длиною наравне с одним из оных уделов от западного предела до восточного.
EZEK|45|8|Это его земля, его владение в Израиле, чтобы князья Мои вперед не теснили народа Моего и чтобы предоставили землю дому Израилеву по коленам его.
EZEK|45|9|Так говорит Господь Бог: довольно вам, князья Израилевы! отложите обиды и угнетения и творите суд и правду, перестаньте вытеснять народ Мой из владения его, говорит Господь Бог.
EZEK|45|10|Да будут у вас правильные весы и правильная ефа и правильный бат.
EZEK|45|11|Ефа и бат должны быть одинаковой меры, так чтобы бат вмещал в себе десятую часть хомера и ефа десятую часть хомера; мера их должна определяться по хомеру.
EZEK|45|12|В сикле двадцать гер; а двадцать сиклей, двадцать пять сиклей и пятнадцать сиклей составлять будут у вас мину.
EZEK|45|13|Вот дань, какую вы должны давать [князю]: шестую часть ефы от хомера пшеницы и шестую часть ефы от хомера ячменя;
EZEK|45|14|постановление об елее: от кора елея десятую часть бата; десять батов [составят] хомер, потому что в хомере десять батов;
EZEK|45|15|одну овцу от стада в двести овец с тучной пажити Израиля: все это для хлебного приношения и всесожжения, и благодарственной жертвы, в очищение их, говорит Господь Бог.
EZEK|45|16|Весь народ земли обязывается делать сие приношение князю в Израиле.
EZEK|45|17|А на обязанности князя будут лежать всесожжение и хлебное приношение, и возлияние в праздники и в новомесячия, и в субботы, во все торжества дома Израилева; он должен будет приносить жертву за грех и хлебное приношение, и всесожжение, и жертву благодарственную для очищения дома Израилева.
EZEK|45|18|Так говорит Господь Бог: в первом [месяце], в первый [день] месяца, возьми из стада волов тельца без порока, и очисти святилище.
EZEK|45|19|Священник пусть возьмет крови от этой жертвы за грех и покропит ею на вереи храма и на четыре угла площадки у жертвенника и на вереи ворот внутреннего двора.
EZEK|45|20|То же сделай и в седьмой [день] месяца за согрешающих умышленно и по простоте, и так очищайте храм.
EZEK|45|21|В первом [месяце], в четырнадцатый день месяца, должна быть у вас Пасха, праздник семидневный, когда должно есть опресноки.
EZEK|45|22|В этот день князь за себя и за весь народ земли принесет тельца в жертву за грех.
EZEK|45|23|И в эти семь дней праздника он должен приносить во всесожжение Господу каждый день по семи тельцов и по семи овнов без порока, и в жертву за грех каждый день по козлу из козьего стада.
EZEK|45|24|Хлебного приношения он должен приносить по ефе на тельца и по ефе на овна и по гину елея на ефу.
EZEK|45|25|В седьмом [месяце], в пятнадцатый день месяца, в праздник, в течение семи дней он должен приносить то же: такую же жертву за грех, такое же всесожжение, и столько же хлебного приношения и столько же елея.
EZEK|46|1|Так говорит Господь Бог: ворота внутреннего двора, обращенные лицом к востоку, должны быть заперты в продолжение шести рабочих дней, а в субботний день они должны быть отворены и в день новомесячия должны быть отворены.
EZEK|46|2|Князь пойдет через внешний притвор ворот и станет у вереи этих ворот; и священники совершат его всесожжение и его благодарственную жертву; и он у порога ворот поклонится [Господу], и выйдет, а ворота остаются незапертыми до вечера.
EZEK|46|3|И народ земли будет поклоняться пред Господом, при входе в ворота, в субботы и новомесячия.
EZEK|46|4|Всесожжение, которое князь принесет Господу в субботний день, должно быть из шести агнцев без порока и из овна без порока;
EZEK|46|5|хлебного приношения ефа на овна, а на агнцев хлебного приношения, сколько рука его подаст, а елея гин на ефу.
EZEK|46|6|В день новомесячия будут приносимы им из стада волов телец без порока, также шесть агнцев и овен без порока.
EZEK|46|7|Хлебного приношения он принесет ефу на тельца и ефу на овна, а на агнцев, сколько рука его подаст, и елея гин на ефу.
EZEK|46|8|И когда приходить будет князь, то должен входить через притвор ворот и тем же путем выходить.
EZEK|46|9|А когда народ земли будет приходить пред лице Господа в праздники, то вошедший северными воротами для поклонения должен выходить воротами южными, а вошедший южными воротами должен выходить воротами северными; он не должен выходить теми же воротами, которыми вошел, а должен выходить противоположными.
EZEK|46|10|И князь должен находиться среди них; когда они входят, входит и он; и когда они выходят, выходит и он.
EZEK|46|11|И в праздники и в торжественные дни хлебного приношения [от] [него] должно быть по ефе на тельца и по ефе на овна, а на агнцев, сколько подаст рука его, и елея по гину на ефу.
EZEK|46|12|А если князь, по усердию своему, захочет принести всесожжение или благодарственную жертву Господу, то должны отворить ему ворота, обращенные к востоку, и он совершит свое всесожжение и свою благодарственную жертву так же, как совершил в субботний день, и после сего он выйдет, и по выходе его ворота запрутся.
EZEK|46|13|Каждый день приноси Господу во всесожжение однолетнего агнца без порока; каждое утро приноси его.
EZEK|46|14|А хлебного приношения прилагай к нему каждое утро шестую часть ефы и елея третью часть гина, чтобы растворить муку; таково вечное постановление о хлебном приношении Господу, навсегда.
EZEK|46|15|Пусть приносят во всесожжение агнца и хлебное приношение и елей каждое утро постоянно.
EZEK|46|16|Так говорит Господь Бог: если князь дает кому из сыновей своих подарок, то это должно пойти в наследство и его сыновьям; это владение их должно быть наследственным.
EZEK|46|17|Если же он даст из наследия своего кому–либо из рабов своих подарок, то это будет принадлежать ему только до года освобождения, и тогда возвратится к князю. Только к сыновьям его должно переходить наследие его.
EZEK|46|18|Но князь не может брать из наследственного участка народа, вытесняя их из владения их; из своего только владения он может уделять детям своим, чтобы никто из народа Моего не был изгоняем из своего владения.
EZEK|46|19|И привел он меня тем ходом, который сбоку ворот, к священным комнатам для священников, обращенным к северу, и вот там одно место на краю к западу.
EZEK|46|20|И сказал мне: "это – место, где священники должны варить жертву за преступление и жертву за грех, где должны печь хлебное приношение, не вынося его на внешний двор, для освящения народа".
EZEK|46|21|И вывел меня на внешний двор, и провел меня по четырем углам двора, и вот, в каждом углу двора еще двор.
EZEK|46|22|Во всех четырех углах двора были покрытые дворы в сорок [локтей] длины и тридцать ширины, одной меры во всех четырех углах.
EZEK|46|23|И кругом всех их четырех – стены, а у стен сделаны очаги кругом.
EZEK|46|24|И сказал мне: "вот поварни, в которых служители храма варят жертвы народные".
EZEK|47|1|Потом привел он меня обратно к дверям храма, и вот, из–под порога храма течет вода на восток, ибо храм стоял лицом на восток, и вода текла из–под правого бока храма, по южную сторону жертвенника.
EZEK|47|2|И вывел меня северными воротами, и внешним путем обвел меня к внешним воротам, путем, обращенным к востоку; и вот, вода течет по правую сторону.
EZEK|47|3|Когда тот муж пошел на восток, то в руке держал шнур, и отмерил тысячу локтей, и повел меня по воде; воды было по лодыжку.
EZEK|47|4|И [еще] отмерил тысячу, и повел меня по воде; воды было по колено. И еще отмерил тысячу, и повел меня; воды было по поясницу.
EZEK|47|5|И еще отмерил тысячу, и уже тут был такой поток, через который я не мог идти, потому что вода была так высока, что надлежало плыть, а переходить нельзя было этот поток.
EZEK|47|6|И сказал мне: "видел, сын человеческий?" и повел меня обратно к берегу этого потока.
EZEK|47|7|И когда я пришел назад, и вот, на берегах потока много было дерев по ту и другую сторону.
EZEK|47|8|И сказал мне: эта вода течет в восточную сторону земли, сойдет на равнину и войдет в море; и воды его сделаются здоровыми.
EZEK|47|9|И всякое живущее существо, пресмыкающееся там, где войдут две струи, будет живо; и рыбы будет весьма много, потому что войдет туда эта вода, и воды [в море] сделаются здоровыми, и, куда войдет этот поток, все будет живо там.
EZEK|47|10|И будут стоять подле него рыболовы от Ен–Гадди до Эглаима, будут закидывать сети. Рыба будет в своем виде и, как в большом море, рыбы будет весьма много.
EZEK|47|11|Болота его и лужи его, которые не сделаются здоровыми, будут оставлены для соли.
EZEK|47|12|У потока по берегам его, с той и другой стороны, будут расти всякие дерева, доставляющие пищу: листья их не будут увядать, и плоды на них не будут истощаться; каждый месяц будут созревать новые, потому что вода для них течет из святилища; плоды их будут употребляемы в пищу, а листья на врачевание.
EZEK|47|13|Так говорит Господь Бог: вот распределение, по которому вы должны разделить землю в наследие двенадцати коленам Израилевым: Иосифу два удела.
EZEK|47|14|И наследуйте ее, как один, так и другой; так как Я, подняв руку Мою, клялся отдать ее отцам вашим, то и будет земля сия наследием вашим.
EZEK|47|15|И вот предел земли: на северном конце, начиная от великого моря, через Хетлон, по дороге в Цедад,
EZEK|47|16|Емаф, Берот, Сивраим, находящийся между Дамасскою и Емафскою областями Гацар–Тихон, который на границе Аврана.
EZEK|47|17|И будет граница от моря до Гацар–Енон, граница с Дамаском, и далее на севере область Емаф; и вот северный край.
EZEK|47|18|Черту восточного края ведите между Авраном и Дамаском, между Галаадом и землею Израильскою, по Иордану, от северного края до восточного моря; это восточный край.
EZEK|47|19|А южный край с полуденной стороны от Тамары до вод пререкания при Кадисе, и по течению потока до великого моря; это полуденный край на юге.
EZEK|47|20|Западный же предел – великое море, от южной границы до места против Емафа; это западный край.
EZEK|47|21|И разделите себе землю сию на уделы по коленам Израилевым.
EZEK|47|22|И разделите ее по жребию в наследие себе и иноземцам, живущим у вас, которые родили у вас детей; и они среди сынов Израилевых должны считаться наравне с природными жителями, и они с вами войдут в долю среди колен Израилевых.
EZEK|47|23|В котором колене живет иноземец, в том и дайте ему наследие его, говорит Господь Бог.
EZEK|48|1|Вот имена колен. На северном краю по дороге от Хетлона, ведущей в Емаф, Гацар–Енон, от северной границы Дамаска по пути к Емафу: все это от востока до моря один удел Дану.
EZEK|48|2|Подле границы Дана, от восточного края до западного, это один удел Асиру.
EZEK|48|3|Подле границы Асира, от восточного края до западного, это один удел Неффалиму.
EZEK|48|4|Подле границы Неффалима, от восточного края до западного, это один удел Манассии.
EZEK|48|5|Подле границы Манассии, от восточного края до западного, это один удел Ефрему.
EZEK|48|6|Подле границы Ефрема, от восточного края до западного, это один удел Рувиму.
EZEK|48|7|Подле границы Рувима, от восточного края до западного, это один удел Иуде.
EZEK|48|8|А подле границы Иуды, от восточного края до западного, священный участок, шириною в двадцать пять тысяч [тростей], а длиною наравне с другими уделами, от восточного края до западного; среди него будет святилище.
EZEK|48|9|Участок, который вы посвятите Господу, длиною будет в двадцать пять тысяч, а шириною в десять тысяч [тростей].
EZEK|48|10|И этот священный участок должен принадлежать священникам, к северу двадцать пять тысяч и к морю в ширину десять тысяч, и к востоку в ширину десять тысяч, а к югу в длину двадцать пять тысяч [тростей], и среди него будет святилище Господне.
EZEK|48|11|Это посвятите священникам из сынов Садока, которые стояли на страже Моей, которые во время отступничества сынов Израилевых не отступили от Меня, как отступили [другие] левиты.
EZEK|48|12|Им будет принадлежать эта часть земли из священного участка, святыня из святынь, у предела левитов.
EZEK|48|13|И левиты получат также у священнического предела двадцать пять тысяч в длину и десять тысяч [тростей] в ширину; вся длина двадцать пять тысяч, а ширина десять тысяч [тростей].
EZEK|48|14|И из этой части они не могут ни продать, ни променять; и начатки земли не могут переходить к другим, потому что это святыня Господня.
EZEK|48|15|А остальные пять тысяч в ширину с двадцатью пятью тысячами [в] [длину] назначаются для города в общее употребление, на заселение и на предместья; город будет в средине.
EZEK|48|16|И вот размеры его: северная сторона четыре тысячи пятьсот и южная сторона четыре тысячи пятьсот, восточная сторона четыре тысячи пятьсот и западная сторона четыре тысячи пятьсот [тростей].
EZEK|48|17|А предместья города к северу двести пятьдесят, и к востоку двести пятьдесят, и к югу двести пятьдесят, и к западу двести пятьдесят [тростей].
EZEK|48|18|А что остается из длины против священного участка, десять тысяч к востоку и десять тысяч к западу, против священного участка, произведения с этой земли должны быть для продовольствия работающих в городе.
EZEK|48|19|Работать же в городе могут работники из всех колен Израилевых.
EZEK|48|20|Весь отделенный участок в двадцать пять тысяч длины и в двадцать пять тысяч ширины, четырехугольный, выделите в священный удел, со включением владений города;
EZEK|48|21|а остальное князю. Как со стороны священного участка, так и со стороны владений города, против двадцати пяти тысяч [тростей] до восточной границы участка, и на запад против двадцати пяти тысяч у западной границы соразмерно с сими уделами, удел князю, так что священный участок и святилище будет в средине его.
EZEK|48|22|И то, что от владений левитских [и] от владений города остается в промежутке, принадлежит также князю; промежуток между границею Иуды и между границею Вениамина будет принадлежать князю.
EZEK|48|23|Остальное же от колен, от восточного края до западного – один удел Вениамину.
EZEK|48|24|Подле границы Вениамина, от восточного края до западного – один удел Симеону.
EZEK|48|25|Подле границы Симеона, от восточного края до западного – один удел Иссахару.
EZEK|48|26|Подле границы Иссахара, от восточного края до западного – один удел Завулону.
EZEK|48|27|Подле границы Завулона, от восточного края до западного – один удел Гаду.
EZEK|48|28|А подле границы Гада на южной стороне идет южный предел от Тамары к водам пререкания при Кадисе, вдоль потока до великого моря.
EZEK|48|29|Вот земля, которую вы по жребию разделите коленам Израилевым, и вот участки их, говорит Господь Бог.
EZEK|48|30|И вот выходы города: с северной стороны меры четыре тысячи пятьсот;
EZEK|48|31|и ворота города называются именами колен Израилевых; к северу трое ворот: ворота Рувимовы одни, ворота Иудины одни, ворота Левиины одни.
EZEK|48|32|И с восточной стороны [меры] четыре тысячи пятьсот, и трое ворот: ворота Иосифовы одни, ворота Вениаминовы одни, ворота Дановы одни;
EZEK|48|33|и с южной стороны меры четыре тысячи пятьсот, и трое ворот: ворота Симеоновы одни, ворота Иссахаровы одни, ворота Завулоновы одни.
EZEK|48|34|С морской стороны [меры] четыре тысячи пятьсот, ворот здесь трое же: ворота Гадовы одни, ворота Асировы одни, ворота Неффалимовы одни.
EZEK|48|35|Всего кругом восемнадцать тысяч. А имя городу с того дня будет: "Господь там".
