JAS|1|1|James, a servant of God and of the Lord Jesus Christ, to the twelve tribes which are scattered abroad, greeting.
JAS|1|2|My brethren, count it all joy when ye fall into divers temptations;
JAS|1|3|Knowing this, that the trying of your faith worketh patience.
JAS|1|4|But let patience have her perfect work, that ye may be perfect and entire, wanting nothing.
JAS|1|5|If any of you lack wisdom, let him ask of God, that giveth to all men liberally, and upbraideth not; and it shall be given him.
JAS|1|6|But let him ask in faith, nothing wavering. For he that wavereth is like a wave of the sea driven with the wind and tossed.
JAS|1|7|For let not that man think that he shall receive any thing of the Lord.
JAS|1|8|A double minded man is unstable in all his ways.
JAS|1|9|Let the brother of low degree rejoice in that he is exalted:
JAS|1|10|But the rich, in that he is made low: because as the flower of the grass he shall pass away.
JAS|1|11|For the sun is no sooner risen with a burning heat, but it withereth the grass, and the flower thereof falleth, and the grace of the fashion of it perisheth: so also shall the rich man fade away in his ways.
JAS|1|12|Blessed is the man that endureth temptation: for when he is tried, he shall receive the crown of life, which the Lord hath promised to them that love him.
JAS|1|13|Let no man say when he is tempted, I am tempted of God: for God cannot be tempted with evil, neither tempteth he any man:
JAS|1|14|But every man is tempted, when he is drawn away of his own lust, and enticed.
JAS|1|15|Then when lust hath conceived, it bringeth forth sin: and sin, when it is finished, bringeth forth death.
JAS|1|16|Do not err, my beloved brethren.
JAS|1|17|Every good gift and every perfect gift is from above, and cometh down from the Father of lights, with whom is no variableness, neither shadow of turning.
JAS|1|18|Of his own will begat he us with the word of truth, that we should be a kind of firstfruits of his creatures.
JAS|1|19|Wherefore, my beloved brethren, let every man be swift to hear, slow to speak, slow to wrath:
JAS|1|20|For the wrath of man worketh not the righteousness of God.
JAS|1|21|Wherefore lay apart all filthiness and superfluity of naughtiness, and receive with meekness the engrafted word, which is able to save your souls.
JAS|1|22|But be ye doers of the word, and not hearers only, deceiving your own selves.
JAS|1|23|For if any be a hearer of the word, and not a doer, he is like unto a man beholding his natural face in a glass:
JAS|1|24|For he beholdeth himself, and goeth his way, and straightway forgetteth what manner of man he was.
JAS|1|25|But whoso looketh into the perfect law of liberty, and continueth therein, he being not a forgetful hearer, but a doer of the work, this man shall be blessed in his deed.
JAS|1|26|If any man among you seem to be religious, and bridleth not his tongue, but deceiveth his own heart, this man's religion is vain.
JAS|1|27|Pure religion and undefiled before God and the Father is this, To visit the fatherless and widows in their affliction, and to keep himself unspotted from the world.
JAS|2|1|My brethren, have not the faith of our Lord Jesus Christ, the Lord of glory, with respect of persons.
JAS|2|2|For if there come unto your assembly a man with a gold ring, in goodly apparel, and there come in also a poor man in vile raiment;
JAS|2|3|And ye have respect to him that weareth the gay clothing, and say unto him, Sit thou here in a good place; and say to the poor, Stand thou there, or sit here under my footstool:
JAS|2|4|Are ye not then partial in yourselves, and are become judges of evil thoughts?
JAS|2|5|Hearken, my beloved brethren, Hath not God chosen the poor of this world rich in faith, and heirs of the kingdom which he hath promised to them that love him?
JAS|2|6|But ye have despised the poor. Do not rich men oppress you, and draw you before the judgment seats?
JAS|2|7|Do not they blaspheme that worthy name by the which ye are called?
JAS|2|8|If ye fulfil the royal law according to the scripture, Thou shalt love thy neighbour as thyself, ye do well:
JAS|2|9|But if ye have respect to persons, ye commit sin, and are convinced of the law as transgressors.
JAS|2|10|For whosoever shall keep the whole law, and yet offend in one point, he is guilty of all.
JAS|2|11|For he that said, Do not commit adultery, said also, Do not kill. Now if thou commit no adultery, yet if thou kill, thou art become a transgressor of the law.
JAS|2|12|So speak ye, and so do, as they that shall be judged by the law of liberty.
JAS|2|13|For he shall have judgment without mercy, that hath shewed no mercy; and mercy rejoiceth against judgment.
JAS|2|14|What doth it profit, my brethren, though a man say he hath faith, and have not works? can faith save him?
JAS|2|15|If a brother or sister be naked, and destitute of daily food,
JAS|2|16|And one of you say unto them, Depart in peace, be ye warmed and filled; notwithstanding ye give them not those things which are needful to the body; what doth it profit?
JAS|2|17|Even so faith, if it hath not works, is dead, being alone.
JAS|2|18|Yea, a man may say, Thou hast faith, and I have works: shew me thy faith without thy works, and I will shew thee my faith by my works.
JAS|2|19|Thou believest that there is one God; thou doest well: the devils also believe, and tremble.
JAS|2|20|But wilt thou know, O vain man, that faith without works is dead?
JAS|2|21|Was not Abraham our father justified by works, when he had offered Isaac his son upon the altar?
JAS|2|22|Seest thou how faith wrought with his works, and by works was faith made perfect?
JAS|2|23|And the scripture was fulfilled which saith, Abraham believed God, and it was imputed unto him for righteousness: and he was called the Friend of God.
JAS|2|24|Ye see then how that by works a man is justified, and not by faith only.
JAS|2|25|Likewise also was not Rahab the harlot justified by works, when she had received the messengers, and had sent them out another way?
JAS|2|26|For as the body without the spirit is dead, so faith without works is dead also.
JAS|3|1|My brethren, be not many masters, knowing that we shall receive the greater condemnation.
JAS|3|2|For in many things we offend all. If any man offend not in word, the same is a perfect man, and able also to bridle the whole body.
JAS|3|3|Behold, we put bits in the horses' mouths, that they may obey us; and we turn about their whole body.
JAS|3|4|Behold also the ships, which though they be so great, and are driven of fierce winds, yet are they turned about with a very small helm, whithersoever the governor listeth.
JAS|3|5|Even so the tongue is a little member, and boasteth great things. Behold, how great a matter a little fire kindleth!
JAS|3|6|And the tongue is a fire, a world of iniquity: so is the tongue among our members, that it defileth the whole body, and setteth on fire the course of nature; and it is set on fire of hell.
JAS|3|7|For every kind of beasts, and of birds, and of serpents, and of things in the sea, is tamed, and hath been tamed of mankind:
JAS|3|8|But the tongue can no man tame; it is an unruly evil, full of deadly poison.
JAS|3|9|Therewith bless we God, even the Father; and therewith curse we men, which are made after the similitude of God.
JAS|3|10|Out of the same mouth proceedeth blessing and cursing. My brethren, these things ought not so to be.
JAS|3|11|Doth a fountain send forth at the same place sweet water and bitter?
JAS|3|12|Can the fig tree, my brethren, bear olive berries? either a vine, figs? so can no fountain both yield salt water and fresh.
JAS|3|13|Who is a wise man and endued with knowledge among you? let him shew out of a good conversation his works with meekness of wisdom.
JAS|3|14|But if ye have bitter envying and strife in your hearts, glory not, and lie not against the truth.
JAS|3|15|This wisdom descendeth not from above, but is earthly, sensual, devilish.
JAS|3|16|For where envying and strife is, there is confusion and every evil work.
JAS|3|17|But the wisdom that is from above is first pure, then peaceable, gentle, and easy to be intreated, full of mercy and good fruits, without partiality, and without hypocrisy.
JAS|3|18|And the fruit of righteousness is sown in peace of them that make peace.
JAS|4|1|From whence come wars and fightings among you? come they not hence, even of your lusts that war in your members?
JAS|4|2|Ye lust, and have not: ye kill, and desire to have, and cannot obtain: ye fight and war, yet ye have not, because ye ask not.
JAS|4|3|Ye ask, and receive not, because ye ask amiss, that ye may consume it upon your lusts.
JAS|4|4|Ye adulterers and adulteresses, know ye not that the friendship of the world is enmity with God? whosoever therefore will be a friend of the world is the enemy of God.
JAS|4|5|Do ye think that the scripture saith in vain, The spirit that dwelleth in us lusteth to envy?
JAS|4|6|But he giveth more grace. Wherefore he saith, God resisteth the proud, but giveth grace unto the humble.
JAS|4|7|Submit yourselves therefore to God. Resist the devil, and he will flee from you.
JAS|4|8|Draw nigh to God, and he will draw nigh to you. Cleanse your hands, ye sinners; and purify your hearts, ye double minded.
JAS|4|9|Be afflicted, and mourn, and weep: let your laughter be turned to mourning, and your joy to heaviness.
JAS|4|10|Humble yourselves in the sight of the Lord, and he shall lift you up.
JAS|4|11|Speak not evil one of another, brethren. He that speaketh evil of his brother, and judgeth his brother, speaketh evil of the law, and judgeth the law: but if thou judge the law, thou art not a doer of the law, but a judge.
JAS|4|12|There is one lawgiver, who is able to save and to destroy: who art thou that judgest another?
JAS|4|13|Go to now, ye that say, To day or to morrow we will go into such a city, and continue there a year, and buy and sell, and get gain:
JAS|4|14|Whereas ye know not what shall be on the morrow. For what is your life? It is even a vapour, that appeareth for a little time, and then vanisheth away.
JAS|4|15|For that ye ought to say, If the Lord will, we shall live, and do this, or that.
JAS|4|16|But now ye rejoice in your boastings: all such rejoicing is evil.
JAS|4|17|Therefore to him that knoweth to do good, and doeth it not, to him it is sin.
JAS|5|1|Go to now, ye rich men, weep and howl for your miseries that shall come upon you.
JAS|5|2|Your riches are corrupted, and your garments are motheaten.
JAS|5|3|Your gold and silver is cankered; and the rust of them shall be a witness against you, and shall eat your flesh as it were fire. Ye have heaped treasure together for the last days.
JAS|5|4|Behold, the hire of the labourers who have reaped down your fields, which is of you kept back by fraud, crieth: and the cries of them which have reaped are entered into the ears of the Lord of sabaoth.
JAS|5|5|Ye have lived in pleasure on the earth, and been wanton; ye have nourished your hearts, as in a day of slaughter.
JAS|5|6|Ye have condemned and killed the just; and he doth not resist you.
JAS|5|7|Be patient therefore, brethren, unto the coming of the Lord. Behold, the husbandman waiteth for the precious fruit of the earth, and hath long patience for it, until he receive the early and latter rain.
JAS|5|8|Be ye also patient; stablish your hearts: for the coming of the Lord draweth nigh.
JAS|5|9|Grudge not one against another, brethren, lest ye be condemned: behold, the judge standeth before the door.
JAS|5|10|Take, my brethren, the prophets, who have spoken in the name of the Lord, for an example of suffering affliction, and of patience.
JAS|5|11|Behold, we count them happy which endure. Ye have heard of the patience of Job, and have seen the end of the Lord; that the Lord is very pitiful, and of tender mercy.
JAS|5|12|But above all things, my brethren, swear not, neither by heaven, neither by the earth, neither by any other oath: but let your yea be yea; and your nay, nay; lest ye fall into condemnation.
JAS|5|13|Is any among you afflicted? let him pray. Is any merry? let him sing psalms.
JAS|5|14|Is any sick among you? let him call for the elders of the church; and let them pray over him, anointing him with oil in the name of the Lord:
JAS|5|15|And the prayer of faith shall save the sick, and the Lord shall raise him up; and if he have committed sins, they shall be forgiven him.
JAS|5|16|Confess your faults one to another, and pray one for another, that ye may be healed. The effectual fervent prayer of a righteous man availeth much.
JAS|5|17|Elias was a man subject to like passions as we are, and he prayed earnestly that it might not rain: and it rained not on the earth by the space of three years and six months.
JAS|5|18|And he prayed again, and the heaven gave rain, and the earth brought forth her fruit.
JAS|5|19|Brethren, if any of you do err from the truth, and one convert him;
JAS|5|20|Let him know, that he which converteth the sinner from the error of his way shall save a soul from death, and shall hide a multitude of sins.
