JUDE|1|1|Jude, the servant of Jesus Christ, and brother of James, to them that are sanctified by God the Father, and preserved in Jesus Christ, and called:
JUDE|1|2|Mercy unto you, and peace, and love, be multiplied.
JUDE|1|3|Beloved, when I gave all diligence to write unto you of the common salvation, it was needful for me to write unto you, and exhort you that ye should earnestly contend for the faith which was once delivered unto the saints.
JUDE|1|4|For there are certain men crept in unawares, who were before of old ordained to this condemnation, ungodly men, turning the grace of our God into lasciviousness, and denying the only Lord God, and our Lord Jesus Christ.
JUDE|1|5|I will therefore put you in remembrance, though ye once knew this, how that the Lord, having saved the people out of the land of Egypt, afterward destroyed them that believed not.
JUDE|1|6|And the angels which kept not their first estate, but left their own habitation, he hath reserved in everlasting chains under darkness unto the judgment of the great day.
JUDE|1|7|Even as Sodom and Gomorrha, and the cities about them in like manner, giving themselves over to fornication, and going after strange flesh, are set forth for an example, suffering the vengeance of eternal fire.
JUDE|1|8|Likewise also these filthy dreamers defile the flesh, despise dominion, and speak evil of dignities.
JUDE|1|9|Yet Michael the archangel, when contending with the devil he disputed about the body of Moses, durst not bring against him a railing accusation, but said, The Lord rebuke thee.
JUDE|1|10|But these speak evil of those things which they know not: but what they know naturally, as brute beasts, in those things they corrupt themselves.
JUDE|1|11|Woe unto them! for they have gone in the way of Cain, and ran greedily after the error of Balaam for reward, and perished in the gainsaying of Core.
JUDE|1|12|These are spots in your feasts of charity, when they feast with you, feeding themselves without fear: clouds they are without water, carried about of winds; trees whose fruit withereth, without fruit, twice dead, plucked up by the roots;
JUDE|1|13|Raging waves of the sea, foaming out their own shame; wandering stars, to whom is reserved the blackness of darkness for ever.
JUDE|1|14|And Enoch also, the seventh from Adam, prophesied of these, saying, Behold, the Lord cometh with ten thousands of his saints,
JUDE|1|15|To execute judgment upon all, and to convince all that are ungodly among them of all their ungodly deeds which they have ungodly committed, and of all their hard speeches which ungodly sinners have spoken against him.
JUDE|1|16|These are murmurers, complainers, walking after their own lusts; and their mouth speaketh great swelling words, having men's persons in admiration because of advantage.
JUDE|1|17|But, beloved, remember ye the words which were spoken before of the apostles of our Lord Jesus Christ;
JUDE|1|18|How that they told you there should be mockers in the last time, who should walk after their own ungodly lusts.
JUDE|1|19|These be they who separate themselves, sensual, having not the Spirit.
JUDE|1|20|But ye, beloved, building up yourselves on your most holy faith, praying in the Holy Ghost,
JUDE|1|21|Keep yourselves in the love of God, looking for the mercy of our Lord Jesus Christ unto eternal life.
JUDE|1|22|And of some have compassion, making a difference:
JUDE|1|23|And others save with fear, pulling them out of the fire; hating even the garment spotted by the flesh.
JUDE|1|24|Now unto him that is able to keep you from falling, and to present you faultless before the presence of his glory with exceeding joy,
JUDE|1|25|To the only wise God our Saviour, be glory and majesty, dominion and power, both now and ever. Amen.
