ACTS|1|1|Первую книгу написал я [к тебе], Феофил, о всем, что Иисус делал и чему учил от начала
ACTS|1|2|до того дня, в который Он вознесся, дав Святым Духом повеления Апостолам, которых Он избрал,
ACTS|1|3|которым и явил Себя живым, по страдании Своем, со многими верными доказательствами, в продолжение сорока дней являясь им и говоря о Царствии Божием.
ACTS|1|4|И, собрав их, Он повелел им: не отлучайтесь из Иерусалима, но ждите обещанного от Отца, о чем вы слышали от Меня,
ACTS|1|5|ибо Иоанн крестил водою, а вы, через несколько дней после сего, будете крещены Духом Святым.
ACTS|1|6|Посему они, сойдясь, спрашивали Его, говоря: не в сие ли время, Господи, восстановляешь Ты царство Израилю?
ACTS|1|7|Он же сказал им: не ваше дело знать времена или сроки, которые Отец положил в Своей власти,
ACTS|1|8|но вы примете силу, когда сойдет на вас Дух Святый; и будете Мне свидетелями в Иерусалиме и во всей Иудее и Самарии и даже до края земли.
ACTS|1|9|Сказав сие, Он поднялся в глазах их, и облако взяло Его из вида их.
ACTS|1|10|И когда они смотрели на небо, во время восхождения Его, вдруг предстали им два мужа в белой одежде
ACTS|1|11|и сказали: мужи Галилейские! что вы стоите и смотрите на небо? Сей Иисус, вознесшийся от вас на небо, придет таким же образом, как вы видели Его восходящим на небо.
ACTS|1|12|Тогда они возвратились в Иерусалим с горы, называемой Елеон, которая находится близ Иерусалима, в расстоянии субботнего пути.
ACTS|1|13|И, придя, взошли в горницу, где и пребывали, Петр и Иаков, Иоанн и Андрей, Филипп и Фома, Варфоломей и Матфей, Иаков Алфеев и Симон Зилот, и Иуда, [брат] Иакова.
ACTS|1|14|Все они единодушно пребывали в молитве и молении, с [некоторыми] женами и Мариею, Материю Иисуса, и с братьями Его.
ACTS|1|15|И в те дни Петр, став посреди учеников, сказал
ACTS|1|16|было же собрание человек около ста двадцати: мужи братия! Надлежало исполниться тому, что в Писании предрек Дух Святый устами Давида об Иуде, бывшем вожде тех, которые взяли Иисуса;
ACTS|1|17|он был сопричислен к нам и получил жребий служения сего;
ACTS|1|18|но приобрел землю неправедною мздою, и когда низринулся, расселось чрево его, и выпали все внутренности его;
ACTS|1|19|и это сделалось известно всем жителям Иерусалима, так что земля та на отечественном их наречии названа Акелдама, то есть земля крови.
ACTS|1|20|В книге же Псалмов написано: да будет двор его пуст, и да не будет живущего в нем; и: достоинство его да приимет другой.
ACTS|1|21|Итак надобно, чтобы один из тех, которые находились с нами во все время, когда пребывал и обращался с нами Господь Иисус,
ACTS|1|22|начиная от крещения Иоаннова до того дня, в который Он вознесся от нас, был вместе с нами свидетелем воскресения Его.
ACTS|1|23|И поставили двоих: Иосифа, называемого Варсавою, который прозван Иустом, и Матфия;
ACTS|1|24|и помолились и сказали: Ты, Господи, Сердцеведец всех, покажи из сих двоих одного, которого Ты избрал
ACTS|1|25|принять жребий сего служения и Апостольства, от которого отпал Иуда, чтобы идти в свое место.
ACTS|1|26|И бросили о них жребий, и выпал жребий Матфию, и он сопричислен к одиннадцати Апостолам.
ACTS|2|1|При наступлении дня Пятидесятницы все они были единодушно вместе.
ACTS|2|2|И внезапно сделался шум с неба, как бы от несущегося сильного ветра, и наполнил весь дом, где они находились.
ACTS|2|3|И явились им разделяющиеся языки, как бы огненные, и почили по одному на каждом из них.
ACTS|2|4|И исполнились все Духа Святаго, и начали говорить на иных языках, как Дух давал им провещевать.
ACTS|2|5|В Иерусалиме же находились Иудеи, люди набожные, из всякого народа под небом.
ACTS|2|6|Когда сделался этот шум, собрался народ, и пришел в смятение, ибо каждый слышал их говорящих его наречием.
ACTS|2|7|И все изумлялись и дивились, говоря между собою: сии говорящие не все ли Галилеяне?
ACTS|2|8|Как же мы слышим каждый собственное наречие, в котором родились.
ACTS|2|9|Парфяне, и Мидяне, и Еламиты, и жители Месопотамии, Иудеи и Каппадокии, Понта и Асии,
ACTS|2|10|Фригии и Памфилии, Египта и частей Ливии, прилежащих к Киринее, и пришедшие из Рима, Иудеи и прозелиты,
ACTS|2|11|критяне и аравитяне, слышим их нашими языками говорящих о великих [делах] Божиих?
ACTS|2|12|И изумлялись все и, недоумевая, говорили друг другу: что это значит?
ACTS|2|13|А иные, насмехаясь, говорили: они напились сладкого вина.
ACTS|2|14|Петр же, став с одиннадцатью, возвысил голос свой и возгласил им: мужи Иудейские, и все живущие в Иерусалиме! сие да будет вам известно, и внимайте словам моим:
ACTS|2|15|они не пьяны, как вы думаете, ибо теперь третий час дня;
ACTS|2|16|но это есть предреченное пророком Иоилем:
ACTS|2|17|И будет в последние дни, говорит Бог, излию от Духа Моего на всякую плоть, и будут пророчествовать сыны ваши и дочери ваши; и юноши ваши будут видеть видения, и старцы ваши сновидениями вразумляемы будут.
ACTS|2|18|И на рабов Моих и на рабынь Моих в те дни излию от Духа Моего, и будут пророчествовать.
ACTS|2|19|И покажу чудеса на небе вверху и знамения на земле внизу, кровь и огонь и курение дыма.
ACTS|2|20|Солнце превратится во тьму, и луна – в кровь, прежде нежели наступит день Господень, великий и славный.
ACTS|2|21|И будет: всякий, кто призовет имя Господне, спасется.
ACTS|2|22|Мужи Израильские! выслушайте слова сии: Иисуса Назорея, Мужа, засвидетельствованного вам от Бога силами и чудесами и знамениями, которые Бог сотворил через Него среди вас, как и сами знаете,
ACTS|2|23|Сего, по определенному совету и предведению Божию преданного, вы взяли и, пригвоздив руками беззаконных, убили;
ACTS|2|24|но Бог воскресил Его, расторгнув узы смерти, потому что ей невозможно было удержать Его.
ACTS|2|25|Ибо Давид говорит о Нем: видел я пред собою Господа всегда, ибо Он одесную меня, дабы я не поколебался.
ACTS|2|26|От того возрадовалось сердце мое и возвеселился язык мой; даже и плоть моя упокоится в уповании,
ACTS|2|27|ибо Ты не оставишь души моей в аде и не дашь святому Твоему увидеть тления.
ACTS|2|28|Ты дал мне познать путь жизни, Ты исполнишь меня радостью пред лицем Твоим.
ACTS|2|29|Мужи братия! да будет позволено с дерзновением сказать вам о праотце Давиде, что он и умер и погребен, и гроб его у нас до сего дня.
ACTS|2|30|Будучи же пророком и зная, что Бог с клятвою обещал ему от плода чресл его воздвигнуть Христа во плоти и посадить на престоле его,
ACTS|2|31|Он прежде сказал о воскресении Христа, что не оставлена душа Его в аде, и плоть Его не видела тления.
ACTS|2|32|Сего Иисуса Бог воскресил, чему все мы свидетели.
ACTS|2|33|Итак Он, быв вознесен десницею Божиею и приняв от Отца обетование Святаго Духа, излил то, что вы ныне видите и слышите.
ACTS|2|34|Ибо Давид не восшел на небеса; но сам говорит: сказал Господь Господу моему: седи одесную Меня,
ACTS|2|35|доколе положу врагов Твоих в подножие ног Твоих.
ACTS|2|36|Итак твердо знай, весь дом Израилев, что Бог соделал Господом и Христом Сего Иисуса, Которого вы распяли.
ACTS|2|37|Услышав это, они умилились сердцем и сказали Петру и прочим Апостолам: что нам делать, мужи братия?
ACTS|2|38|Петр же сказал им: покайтесь, и да крестится каждый из вас во имя Иисуса Христа для прощения грехов; и получите дар Святаго Духа.
ACTS|2|39|Ибо вам принадлежит обетование и детям вашим и всем дальним, кого ни призовет Господь Бог наш.
ACTS|2|40|И другими многими словами он свидетельствовал и увещевал, говоря: спасайтесь от рода сего развращенного.
ACTS|2|41|Итак охотно принявшие слово его крестились, и присоединилось в тот день душ около трех тысяч.
ACTS|2|42|И они постоянно пребывали в учении Апостолов, в общении и преломлении хлеба и в молитвах.
ACTS|2|43|Был же страх на всякой душе; и много чудес и знамений совершилось через Апостолов в Иерусалиме.
ACTS|2|44|Все же верующие были вместе и имели все общее.
ACTS|2|45|И продавали имения и всякую собственность, и разделяли всем, смотря по нужде каждого.
ACTS|2|46|И каждый день единодушно пребывали в храме и, преломляя по домам хлеб, принимали пищу в веселии и простоте сердца,
ACTS|2|47|хваля Бога и находясь в любви у всего народа. Господь же ежедневно прилагал спасаемых к Церкви.
ACTS|3|1|Петр и Иоанн шли вместе в храм в час молитвы девятый.
ACTS|3|2|И был человек, хромой от чрева матери его, которого носили и сажали каждый день при дверях храма, называемых Красными, просить милостыни у входящих в храм.
ACTS|3|3|Он, увидев Петра и Иоанна перед входом в храм, просил у них милостыни.
ACTS|3|4|Петр с Иоанном, всмотревшись в него, сказали: взгляни на нас.
ACTS|3|5|И он пристально смотрел на них, надеясь получить от них что–нибудь.
ACTS|3|6|Но Петр сказал: серебра и золота нет у меня; а что имею, то даю тебе: во имя Иисуса Христа Назорея встань и ходи.
ACTS|3|7|И, взяв его за правую руку, поднял; и вдруг укрепились его ступни и колени,
ACTS|3|8|и вскочив, стал, и начал ходить, и вошел с ними в храм, ходя и скача, и хваля Бога.
ACTS|3|9|И весь народ видел его ходящим и хвалящим Бога;
ACTS|3|10|и узнали его, что это был тот, который сидел у Красных дверей храма для милостыни; и исполнились ужаса и изумления от случившегося с ним.
ACTS|3|11|И как исцеленный хромой не отходил от Петра и Иоанна, то весь народ в изумлении сбежался к ним в притвор, называемый Соломонов.
ACTS|3|12|Увидев это, Петр сказал народу: мужи Израильские! что дивитесь сему, или что смотрите на нас, как будто бы мы своею силою или благочестием сделали то, что он ходит?
ACTS|3|13|Бог Авраама и Исаака и Иакова, Бог отцов наших, прославил Сына Своего Иисуса, Которого вы предали и от Которого отреклись перед лицом Пилата, когда он полагал освободить Его.
ACTS|3|14|Но вы от Святого и Праведного отреклись, и просили даровать вам человека убийцу,
ACTS|3|15|а Начальника жизни убили. Сего Бог воскресил из мертвых, чему мы свидетели.
ACTS|3|16|И ради веры во имя Его, имя Его укрепило сего, которого вы видите и знаете, и вера, которая от Него, даровала ему исцеление сие перед всеми вами.
ACTS|3|17|Впрочем я знаю, братия, что вы, как и начальники ваши, сделали это по неведению;
ACTS|3|18|Бог же, как предвозвестил устами всех Своих пророков пострадать Христу, так и исполнил.
ACTS|3|19|Итак покайтесь и обратитесь, чтобы загладились грехи ваши,
ACTS|3|20|да придут времена отрады от лица Господа, и да пошлет Он предназначенного вам Иисуса Христа,
ACTS|3|21|Которого небо должно было принять до времен совершения всего, что говорил Бог устами всех святых Своих пророков от века.
ACTS|3|22|Моисей сказал отцам: Господь Бог ваш воздвигнет вам из братьев ваших Пророка, как меня, слушайтесь Его во всем, что Он ни будет говорить вам;
ACTS|3|23|и будет, что всякая душа, которая не послушает Пророка того, истребится из народа.
ACTS|3|24|И все пророки, от Самуила и после него, сколько их ни говорили, также предвозвестили дни сии.
ACTS|3|25|Вы сыны пророков и завета, который завещевал Бог отцам вашим, говоря Аврааму: и в семени твоем благословятся все племена земные.
ACTS|3|26|Бог, воскресив Сына Своего Иисуса, к вам первым послал Его благословить вас, отвращая каждого от злых дел ваших.
ACTS|4|1|Когда они говорили к народу, к ним приступили священники и начальники стражи при храме и саддукеи,
ACTS|4|2|досадуя на то, что они учат народ и проповедуют в Иисусе воскресение из мертвых;
ACTS|4|3|и наложили на них руки и отдали [их] под стражу до утра; ибо уже был вечер.
ACTS|4|4|Многие же из слушавших слово уверовали; и было число таковых людей около пяти тысяч.
ACTS|4|5|На другой день собрались в Иерусалим начальники их и старейшины, и книжники,
ACTS|4|6|и Анна первосвященник, и Каиафа, и Иоанн, и Александр, и прочие из рода первосвященнического;
ACTS|4|7|и, поставив их посреди, спрашивали: какою силою или каким именем вы сделали это?
ACTS|4|8|Тогда Петр, исполнившись Духа Святаго, сказал им: начальники народа и старейшины Израильские!
ACTS|4|9|Если от нас сегодня требуют ответа в благодеянии человеку немощному, как он исцелен,
ACTS|4|10|то да будет известно всем вам и всему народу Израильскому, что именем Иисуса Христа Назорея, Которого вы распяли, Которого Бог воскресил из мертвых, Им поставлен он перед вами здрав.
ACTS|4|11|Он есть камень, пренебреженный вами зиждущими, но сделавшийся главою угла, и нет ни в ком ином спасения,
ACTS|4|12|ибо нет другого имени под небом, данного человекам, которым надлежало бы нам спастись.
ACTS|4|13|Видя смелость Петра и Иоанна и приметив, что они люди некнижные и простые, они удивлялись, между тем узнавали их, что они были с Иисусом;
ACTS|4|14|видя же исцеленного человека, стоящего с ними, ничего не могли сказать вопреки.
ACTS|4|15|И, приказав им выйти вон из синедриона, рассуждали между собою,
ACTS|4|16|говоря: что нам делать с этими людьми? Ибо всем, живущим в Иерусалиме, известно, что ими сделано явное чудо, и мы не можем отвергнуть [сего];
ACTS|4|17|но, чтобы более не разгласилось это в народе, с угрозою запретим им, чтобы не говорили об имени сем никому из людей.
ACTS|4|18|И, призвав их, приказали им отнюдь не говорить и не учить о имени Иисуса.
ACTS|4|19|Но Петр и Иоанн сказали им в ответ: судите, справедливо ли пред Богом слушать вас более, нежели Бога?
ACTS|4|20|Мы не можем не говорить того, что видели и слышали.
ACTS|4|21|Они же, пригрозив, отпустили их, не находя возможности наказать их, по причине народа; потому что все прославляли Бога за происшедшее.
ACTS|4|22|Ибо лет более сорока было тому человеку, над которым сделалось сие чудо исцеления.
ACTS|4|23|Быв отпущены, они пришли к своим и пересказали, что говорили им первосвященники и старейшины.
ACTS|4|24|Они же, выслушав, единодушно возвысили голос к Богу и сказали: Владыко Боже, сотворивший небо и землю и море и все, что в них!
ACTS|4|25|Ты устами отца нашего Давида, раба Твоего, сказал Духом Святым: что мятутся язычники, и народы замышляют тщетное?
ACTS|4|26|Восстали цари земные, и князи собрались вместе на Господа и на Христа Его.
ACTS|4|27|Ибо поистине собрались в городе сем на Святаго Сына Твоего Иисуса, помазанного Тобою, Ирод и Понтий Пилат с язычниками и народом Израильским,
ACTS|4|28|чтобы сделать то, чему быть предопределила рука Твоя и совет Твой.
ACTS|4|29|И ныне, Господи, воззри на угрозы их, и дай рабам Твоим со всею смелостью говорить слово Твое,
ACTS|4|30|тогда как Ты простираешь руку Твою на исцеления и на соделание знамений и чудес именем Святаго Сына Твоего Иисуса.
ACTS|4|31|И, по молитве их, поколебалось место, где они были собраны, и исполнились все Духа Святаго, и говорили слово Божие с дерзновением.
ACTS|4|32|У множества же уверовавших было одно сердце и одна душа; и никто ничего из имения своего не называл своим, но все у них было общее.
ACTS|4|33|Апостолы же с великою силою свидетельствовали о воскресении Господа Иисуса Христа; и великая благодать была на всех их.
ACTS|4|34|Не было между ними никого нуждающегося; ибо все, которые владели землями или домами, продавая их, приносили цену проданного
ACTS|4|35|и полагали к ногам Апостолов; и каждому давалось, в чем кто имел нужду.
ACTS|4|36|Так Иосия, прозванный от Апостолов Варнавою, что значит – сын утешения, левит, родом Кипрянин,
ACTS|4|37|у которого была своя земля, продав ее, принес деньги и положил к ногам Апостолов.
ACTS|5|1|Некоторый же муж, именем Анания, с женою своею Сапфирою, продав имение,
ACTS|5|2|утаил из цены, с ведома и жены своей, а некоторую часть принес и положил к ногам Апостолов.
ACTS|5|3|Но Петр сказал: Анания! Для чего [ты допустил] сатане вложить в сердце твое [мысль] солгать Духу Святому и утаить из цены земли?
ACTS|5|4|Чем ты владел, не твое ли было, и приобретенное продажею не в твоей ли власти находилось? Для чего ты положил это в сердце твоем? Ты солгал не человекам, а Богу.
ACTS|5|5|Услышав сии слова, Анания пал бездыханен; и великий страх объял всех, слышавших это.
ACTS|5|6|И встав, юноши приготовили его к погребению и, вынеся, похоронили.
ACTS|5|7|Часа через три после сего пришла и жена его, не зная о случившемся.
ACTS|5|8|Петр же спросил ее: скажи мне, за столько ли продали вы землю? Она сказала: да, за столько.
ACTS|5|9|Но Петр сказал ей: что это согласились вы искусить Духа Господня? вот, входят в двери погребавшие мужа твоего; и тебя вынесут.
ACTS|5|10|Вдруг она упала у ног его и испустила дух. И юноши, войдя, нашли ее мертвою и, вынеся, похоронили подле мужа ее.
ACTS|5|11|И великий страх объял всю церковь и всех слышавших это.
ACTS|5|12|Руками же Апостолов совершались в народе многие знамения и чудеса; и все единодушно пребывали в притворе Соломоновом.
ACTS|5|13|Из посторонних же никто не смел пристать к ним, а народ прославлял их.
ACTS|5|14|Верующих же более и более присоединялось к Господу, множество мужчин и женщин,
ACTS|5|15|так что выносили больных на улицы и полагали на постелях и кроватях, дабы хотя тень проходящего Петра осенила кого из них.
ACTS|5|16|Сходились также в Иерусалим многие из окрестных городов, неся больных и нечистыми духами одержимых, которые и исцелялись все.
ACTS|5|17|Первосвященник же и с ним все, принадлежавшие к ереси саддукейской, исполнились зависти,
ACTS|5|18|и наложили руки свои на Апостолов, и заключили их в народную темницу.
ACTS|5|19|Но Ангел Господень ночью отворил двери темницы и, выведя их, сказал:
ACTS|5|20|идите и, став в храме, говорите народу все сии слова жизни.
ACTS|5|21|Они, выслушав, вошли утром в храм и учили. Между тем первосвященник и которые с ним, придя, созвали синедрион и всех старейшин из сынов Израилевых и послали в темницу привести [Апостолов].
ACTS|5|22|Но служители, придя, не нашли их в темнице и, возвратившись, донесли,
ACTS|5|23|говоря: темницу мы нашли запертою со всею предосторожностью и стражей стоящими перед дверями; но, отворив, не нашли в ней никого.
ACTS|5|24|Когда услышали эти слова первосвященник, начальник стражи и [прочие] первосвященники, недоумевали, что бы это значило.
ACTS|5|25|Пришел же некто и донес им, говоря: вот, мужи, которых вы заключили в темницу, стоят в храме и учат народ.
ACTS|5|26|Тогда начальник стражи пошел со служителями и привел их без принуждения, потому что боялись народа, чтобы не побили их камнями.
ACTS|5|27|Приведя же их, поставили в синедрионе; и спросил их первосвященник, говоря:
ACTS|5|28|не запретили ли мы вам накрепко учить о имени сем? и вот, вы наполнили Иерусалим учением вашим и хотите навести на нас кровь Того Человека.
ACTS|5|29|Петр же и Апостолы в ответ сказали: должно повиноваться больше Богу, нежели человекам.
ACTS|5|30|Бог отцов наших воскресил Иисуса, Которого вы умертвили, повесив на древе.
ACTS|5|31|Его возвысил Бог десницею Своею в Начальника и Спасителя, дабы дать Израилю покаяние и прощение грехов.
ACTS|5|32|Свидетели Ему в сем мы и Дух Святый, Которого Бог дал повинующимся Ему.
ACTS|5|33|Слышав это, они разрывались от гнева и умышляли умертвить их.
ACTS|5|34|Встав же в синедрионе, некто фарисей, именем Гамалиил, законоучитель, уважаемый всем народом, приказал вывести Апостолов на короткое время,
ACTS|5|35|а им сказал: мужи Израильские! подумайте сами с собою о людях сих, что вам с ними делать.
ACTS|5|36|Ибо незадолго перед сим явился Февда, выдавая себя за кого–то великого, и к нему пристало около четырехсот человек; но он был убит, и все, которые слушались его, рассеялись и исчезли.
ACTS|5|37|После него во время переписи явился Иуда Галилеянин и увлек за собою довольно народа; но он погиб, и все, которые слушались его, рассыпались.
ACTS|5|38|И ныне, говорю вам, отстаньте от людей сих и оставьте их; ибо если это предприятие и это дело – от человеков, то оно разрушится,
ACTS|5|39|а если от Бога, то вы не можете разрушить его; [берегитесь], чтобы вам не оказаться и богопротивниками.
ACTS|5|40|Они послушались его; и, призвав Апостолов, били [их] и, запретив им говорить о имени Иисуса, отпустили их.
ACTS|5|41|Они же пошли из синедриона, радуясь, что за имя Господа Иисуса удостоились принять бесчестие.
ACTS|5|42|И всякий день в храме и по домам не переставали учить и благовествовать об Иисусе Христе.
ACTS|6|1|В эти дни, когда умножились ученики, произошел у Еллинистов ропот на Евреев за то, что вдовицы их пренебрегаемы были в ежедневном раздаянии потребностей.
ACTS|6|2|Тогда двенадцать [Апостолов], созвав множество учеников, сказали: нехорошо нам, оставив слово Божие, пещись о столах.
ACTS|6|3|Итак, братия, выберите из среды себя семь человек изведанных, исполненных Святаго Духа и мудрости; их поставим на эту службу,
ACTS|6|4|а мы постоянно пребудем в молитве и служении слова.
ACTS|6|5|И угодно было это предложение всему собранию; и избрали Стефана, мужа, исполненного веры и Духа Святаго, и Филиппа, и Прохора, и Никанора, и Тимона, и Пармена, и Николая Антиохийца, обращенного из язычников;
ACTS|6|6|их поставили перед Апостолами, и [сии], помолившись, возложили на них руки.
ACTS|6|7|И слово Божие росло, и число учеников весьма умножалось в Иерусалиме; и из священников очень многие покорились вере.
ACTS|6|8|А Стефан, исполненный веры и силы, совершал великие чудеса и знамения в народе.
ACTS|6|9|Некоторые из так называемой синагоги Либертинцев и Киринейцев и Александрийцев и некоторые из Киликии и Асии вступили в спор со Стефаном;
ACTS|6|10|но не могли противостоять мудрости и Духу, Которым он говорил.
ACTS|6|11|Тогда научили они некоторых сказать: мы слышали, как он говорил хульные слова на Моисея и на Бога.
ACTS|6|12|И возбудили народ и старейшин и книжников и, напав, схватили его и повели в синедрион.
ACTS|6|13|И представили ложных свидетелей, которые говорили: этот человек не перестает говорить хульные слова на святое место сие и на закон.
ACTS|6|14|Ибо мы слышали, как он говорил, что Иисус Назорей разрушит место сие и переменит обычаи, которые передал нам Моисей.
ACTS|6|15|И все, сидящие в синедрионе, смотря на него, видели лице его, как лице Ангела.
ACTS|7|1|Тогда сказал первосвященник: так ли это?
ACTS|7|2|Но он сказал: мужи братия и отцы! послушайте. Бог славы явился отцу нашему Аврааму в Месопотамии, прежде переселения его в Харран,
ACTS|7|3|и сказал ему: выйди из земли твоей и из родства твоего и из дома отца твоего, и пойди в землю, которую покажу тебе.
ACTS|7|4|Тогда он вышел из земли Халдейской и поселился в Харране; а оттуда, по смерти отца его, переселил его [Бог] в сию землю, в которой вы ныне живете.
ACTS|7|5|И не дал ему на ней наследства ни на стопу ноги, а обещал дать ее во владение ему и потомству его по нем, когда еще был он бездетен.
ACTS|7|6|И сказал ему Бог, что потомки его будут переселенцами в чужой земле и будут в порабощении и притеснении лет четыреста.
ACTS|7|7|Но Я, сказал Бог, произведу суд над тем народом, у которого они будут в порабощении; и после того они выйдут и будут служить Мне на сем месте.
ACTS|7|8|И дал ему завет обрезания. По сем родил он Исаака и обрезал его в восьмой день; а Исаак [родил] Иакова, Иаков же двенадцать патриархов.
ACTS|7|9|Патриархи, по зависти, продали Иосифа в Египет; но Бог был с ним,
ACTS|7|10|и избавил его от всех скорбей его, и даровал мудрость ему и благоволение царя Египетского фараона, [который] и поставил его начальником над Египтом и над всем домом своим.
ACTS|7|11|И пришел голод и великая скорбь на всю землю Египетскую и Ханаанскую, и отцы наши не находили пропитания.
ACTS|7|12|Иаков же, услышав, что есть хлеб в Египте, послал [туда] отцов наших в первый раз.
ACTS|7|13|А когда они пришли во второй раз, Иосиф открылся братьям своим, и известен стал фараону род Иосифов.
ACTS|7|14|Иосиф, послав, призвал отца своего Иакова и все родство свое, душ семьдесят пять.
ACTS|7|15|Иаков перешел в Египет, и скончался сам и отцы наши;
ACTS|7|16|и перенесены были в Сихем и положены во гробе, который купил Авраам ценою серебра у сынов Еммора Сихемова.
ACTS|7|17|А по мере, как приближалось время [исполниться] обетованию, о котором клялся Бог Аврааму, народ возрастал и умножался в Египте,
ACTS|7|18|до тех пор, как восстал иной царь, который не знал Иосифа.
ACTS|7|19|Сей, ухищряясь против рода нашего, притеснял отцов наших, принуждая их бросать детей своих, чтобы не оставались в живых.
ACTS|7|20|В это время родился Моисей, и был прекрасен пред Богом. Три месяца он был питаем в доме отца своего.
ACTS|7|21|А когда был брошен, взяла его дочь фараонова и воспитала его у себя, как сына.
ACTS|7|22|И научен был Моисей всей мудрости Египетской, и был силен в словах и делах.
ACTS|7|23|Когда же исполнилось ему сорок лет, пришло ему на сердце посетить братьев своих, сынов Израилевых.
ACTS|7|24|И, увидев одного из них обижаемого, вступился и отмстил за оскорбленного, поразив Египтянина.
ACTS|7|25|Он думал, поймут братья его, что Бог рукою его дает им спасение; но они не поняли.
ACTS|7|26|На следующий день, когда некоторые из них дрались, он явился и склонял их к миру, говоря: вы братья; зачем обижаете друг друга?
ACTS|7|27|Но обижающий ближнего оттолкнул его, сказав: кто тебя поставил начальником и судьею над нами?
ACTS|7|28|Не хочешь ли ты убить и меня, как вчера убил Египтянина?
ACTS|7|29|От сих слов Моисей убежал и сделался пришельцем в земле Мадиамской, где родились от него два сына.
ACTS|7|30|По исполнении сорока лет явился ему в пустыне горы Синая Ангел Господень в пламени горящего тернового куста.
ACTS|7|31|Моисей, увидев, дивился видению; а когда подходил рассмотреть, был к нему глас Господень:
ACTS|7|32|Я Бог отцов твоих, Бог Авраама и Бог Исаака и Бог Иакова. Моисей, объятый трепетом, не смел смотреть.
ACTS|7|33|И сказал ему Господь: сними обувь с ног твоих, ибо место, на котором ты стоишь, есть земля святая.
ACTS|7|34|Я вижу притеснение народа Моего в Египте, и слышу стенание его, и нисшел избавить его: итак пойди, Я пошлю тебя в Египет.
ACTS|7|35|Сего Моисея, которого они отвергли, сказав: кто тебя поставил начальником и судьею? сего Бог чрез Ангела, явившегося ему в терновом кусте, послал начальником и избавителем.
ACTS|7|36|Сей вывел их, сотворив чудеса и знамения в земле Египетской, и в Чермном море, и в пустыне в продолжение сорока лет.
ACTS|7|37|Это тот Моисей, который сказал сынам Израилевым: Пророка воздвигнет вам Господь Бог ваш из братьев ваших, как меня; Его слушайте.
ACTS|7|38|Это тот, который был в собрании в пустыне с Ангелом, говорившим ему на горе Синае, и с отцами нашими, и который принял живые слова, чтобы передать нам,
ACTS|7|39|которому отцы наши не хотели быть послушными, но отринули его и обратились сердцами своими к Египту,
ACTS|7|40|сказав Аарону: сделай нам богов, которые предшествовали бы нам; ибо с Моисеем, который вывел нас из земли Египетской, не знаем, что случилось.
ACTS|7|41|И сделали в те дни тельца, и принесли жертву идолу, и веселились перед делом рук своих.
ACTS|7|42|Бог же отвратился и оставил их служить воинству небесному, как написано в книге пророков: дом Израилев! приносили ли вы Мне заколения и жертвы в продолжение сорока лет в пустыне?
ACTS|7|43|Вы приняли скинию Молохову и звезду бога вашего Ремфана, изображения, которые вы сделали, чтобы поклоняться им: и Я переселю вас далее Вавилона.
ACTS|7|44|Скиния свидетельства была у отцов наших в пустыне, как повелел Говоривший Моисею сделать ее по образцу, им виденному.
ACTS|7|45|Отцы наши с Иисусом, взяв ее, внесли во владения народов, изгнанных Богом от лица отцов наших. [Так было] до дней Давида.
ACTS|7|46|Сей обрел благодать пред Богом и молил, [чтобы] найти жилище Богу Иакова.
ACTS|7|47|Соломон же построил Ему дом.
ACTS|7|48|Но Всевышний не в рукотворенных храмах живет, как говорит пророк:
ACTS|7|49|Небо – престол Мой, и земля – подножие ног Моих. Какой дом созиждете Мне, говорит Господь, или какое место для покоя Моего?
ACTS|7|50|Не Моя ли рука сотворила все сие?
ACTS|7|51|Жестоковыйные! люди с необрезанным сердцем и ушами! вы всегда противитесь Духу Святому, как отцы ваши, так и вы.
ACTS|7|52|Кого из пророков не гнали отцы ваши? Они убили предвозвестивших пришествие Праведника, Которого предателями и убийцами сделались ныне вы, –
ACTS|7|53|вы, которые приняли закон при служении Ангелов и не сохранили.
ACTS|7|54|Слушая сие, они рвались сердцами своими и скрежетали на него зубами.
ACTS|7|55|Стефан же, будучи исполнен Духа Святаго, воззрев на небо, увидел славу Божию и Иисуса, стоящего одесную Бога,
ACTS|7|56|и сказал: вот, я вижу небеса отверстые и Сына Человеческого, стоящего одесную Бога.
ACTS|7|57|Но они, закричав громким голосом, затыкали уши свои, и единодушно устремились на него,
ACTS|7|58|и, выведя за город, стали побивать его камнями. Свидетели же положили свои одежды у ног юноши, именем Савла,
ACTS|7|59|и побивали камнями Стефана, который молился и говорил: Господи Иисусе! приими дух мой.
ACTS|7|60|И, преклонив колени, воскликнул громким голосом: Господи! не вмени им греха сего. И, сказав сие, почил.
ACTS|8|1|Савл же одобрял убиение его. В те дни произошло великое гонение на церковь в Иерусалиме; и все, кроме Апостолов, рассеялись по разным местам Иудеи и Самарии.
ACTS|8|2|Стефана же погребли мужи благоговейные, и сделали великий плач по нем.
ACTS|8|3|А Савл терзал церковь, входя в домы и влача мужчин и женщин, отдавал в темницу.
ACTS|8|4|Между тем рассеявшиеся ходили и благовествовали слово.
ACTS|8|5|Так Филипп пришел в город Самарийский и проповедывал им Христа.
ACTS|8|6|Народ единодушно внимал тому, что говорил Филипп, слыша и видя, какие он творил чудеса.
ACTS|8|7|Ибо нечистые духи из многих, одержимых ими, выходили с великим воплем, а многие расслабленные и хромые исцелялись.
ACTS|8|8|И была радость великая в том городе.
ACTS|8|9|Находился же в городе некоторый муж, именем Симон, который перед тем волхвовал и изумлял народ Самарийский, выдавая себя за кого–то великого.
ACTS|8|10|Ему внимали все, от малого до большого, говоря: сей есть великая сила Божия.
ACTS|8|11|А внимали ему потому, что он немалое время изумлял их волхвованиями.
ACTS|8|12|Но, когда поверили Филиппу, благовествующему о Царствии Божием и о имени Иисуса Христа, то крестились и мужчины и женщины.
ACTS|8|13|Уверовал и сам Симон и, крестившись, не отходил от Филиппа; и, видя совершающиеся великие силы и знамения, изумлялся.
ACTS|8|14|Находившиеся в Иерусалиме Апостолы, услышав, что Самаряне приняли слово Божие, послали к ним Петра и Иоанна,
ACTS|8|15|которые, придя, помолились о них, чтобы они приняли Духа Святаго.
ACTS|8|16|Ибо Он не сходил еще ни на одного из них, а только были они крещены во имя Господа Иисуса.
ACTS|8|17|Тогда возложили руки на них, и они приняли Духа Святаго.
ACTS|8|18|Симон же, увидев, что через возложение рук Апостольских подается Дух Святый, принес им деньги,
ACTS|8|19|говоря: дайте и мне власть сию, чтобы тот, на кого я возложу руки, получал Духа Святаго.
ACTS|8|20|Но Петр сказал ему: серебро твое да будет в погибель с тобою, потому что ты помыслил дар Божий получить за деньги.
ACTS|8|21|Нет тебе в сем части и жребия, ибо сердце твое неправо пред Богом.
ACTS|8|22|Итак покайся в сем грехе твоем, и молись Богу: может быть, опустится тебе помысел сердца твоего;
ACTS|8|23|ибо вижу тебя исполненного горькой желчи и в узах неправды.
ACTS|8|24|Симон же сказал в ответ: помолитесь вы за меня Господу, дабы не постигло меня ничто из сказанного вами.
ACTS|8|25|Они же, засвидетельствовав и проповедав слово Господне, обратно пошли в Иерусалим и во многих селениях Самарийских проповедали Евангелие.
ACTS|8|26|А Филиппу Ангел Господень сказал: встань и иди на полдень, на дорогу, идущую из Иерусалима в Газу, на ту, которая пуста.
ACTS|8|27|Он встал и пошел. И вот, муж Ефиоплянин, евнух, вельможа Кандакии, царицы Ефиопской, хранитель всех сокровищ ее, приезжавший в Иерусалим для поклонения,
ACTS|8|28|возвращался и, сидя на колеснице своей, читал пророка Исаию.
ACTS|8|29|Дух сказал Филиппу: подойди и пристань к сей колеснице.
ACTS|8|30|Филипп подошел и, услышав, что он читает пророка Исаию, сказал: разумеешь ли, что читаешь?
ACTS|8|31|Он сказал: как могу разуметь, если кто не наставит меня? и попросил Филиппа взойти и сесть с ним.
ACTS|8|32|А место из Писания, которое он читал, было сие: как овца, веден был Он на заклание, и, как агнец пред стригущим его безгласен, так Он не отверзает уст Своих.
ACTS|8|33|В уничижении Его суд Его совершился. Но род Его кто разъяснит? ибо вземлется от земли жизнь Его.
ACTS|8|34|Евнух же сказал Филиппу: прошу тебя [сказать]: о ком пророк говорит это? о себе ли, или о ком другом?
ACTS|8|35|Филипп отверз уста свои и, начав от сего Писания, благовествовал ему об Иисусе.
ACTS|8|36|Между тем, продолжая путь, они приехали к воде; и евнух сказал: вот вода; что препятствует мне креститься?
ACTS|8|37|Филипп же сказал ему: если веруешь от всего сердца, можно. Он сказал в ответ: верую, что Иисус Христос есть Сын Божий.
ACTS|8|38|И приказал остановить колесницу, и сошли оба в воду, Филипп и евнух; и крестил его.
ACTS|8|39|Когда же они вышли из воды, Дух Святый сошел на евнуха, а Филиппа восхитил Ангел Господень, и евнух уже не видел его, и продолжал путь, радуясь.
ACTS|8|40|А Филипп оказался в Азоте и, проходя, благовествовал всем городам, пока пришел в Кесарию.
ACTS|9|1|Савл же, еще дыша угрозами и убийством на учеников Господа, пришел к первосвященнику
ACTS|9|2|и выпросил у него письма в Дамаск к синагогам, чтобы, кого найдет последующих сему учению, и мужчин и женщин, связав, приводить в Иерусалим.
ACTS|9|3|Когда же он шел и приближался к Дамаску, внезапно осиял его свет с неба.
ACTS|9|4|Он упал на землю и услышал голос, говорящий ему: Савл, Савл! что ты гонишь Меня?
ACTS|9|5|Он сказал: кто Ты, Господи? Господь же сказал: Я Иисус, Которого ты гонишь. Трудно тебе идти против рожна.
ACTS|9|6|Он в трепете и ужасе сказал: Господи! что повелишь мне делать? и Господь [сказал] ему: встань и иди в город; и сказано будет тебе, что тебе надобно делать.
ACTS|9|7|Люди же, шедшие с ним, стояли в оцепенении, слыша голос, а никого не видя.
ACTS|9|8|Савл встал с земли, и с открытыми глазами никого не видел. И повели его за руки, и привели в Дамаск.
ACTS|9|9|И три дня он не видел, и не ел, и не пил.
ACTS|9|10|В Дамаске был один ученик, именем Анания; и Господь в видении сказал ему: Анания! Он сказал: я, Господи.
ACTS|9|11|Господь же [сказал] ему: встань и пойди на улицу, так называемую Прямую, и спроси в Иудином доме Тарсянина, по имени Савла; он теперь молится,
ACTS|9|12|и видел в видении мужа, именем Ананию, пришедшего к нему и возложившего на него руку, чтобы он прозрел.
ACTS|9|13|Анания отвечал: Господи! я слышал от многих о сем человеке, сколько зла сделал он святым Твоим в Иерусалиме;
ACTS|9|14|и здесь имеет от первосвященников власть вязать всех, призывающих имя Твое.
ACTS|9|15|Но Господь сказал ему: иди, ибо он есть Мой избранный сосуд, чтобы возвещать имя Мое перед народами и царями и сынами Израилевыми.
ACTS|9|16|И Я покажу ему, сколько он должен пострадать за имя Мое.
ACTS|9|17|Анания пошел и вошел в дом и, возложив на него руки, сказал: брат Савл! Господь Иисус, явившийся тебе на пути, которым ты шел, послал меня, чтобы ты прозрел и исполнился Святаго Духа.
ACTS|9|18|И тотчас как бы чешуя отпала от глаз его, и вдруг он прозрел; и, встав, крестился,
ACTS|9|19|и, приняв пищи, укрепился. И был Савл несколько дней с учениками в Дамаске.
ACTS|9|20|И тотчас стал проповедывать в синагогах об Иисусе, что Он есть Сын Божий.
ACTS|9|21|И все слышавшие дивились и говорили: не тот ли это самый, который гнал в Иерусалиме призывающих имя сие? да и сюда за тем пришел, чтобы вязать их и вести к первосвященникам.
ACTS|9|22|А Савл более и более укреплялся и приводил в замешательство Иудеев, живущих в Дамаске, доказывая, что Сей есть Христос.
ACTS|9|23|Когда же прошло довольно времени, Иудеи согласились убить его.
ACTS|9|24|Но Савл узнал об этом умысле их. А они день и ночь стерегли у ворот, чтобы убить его.
ACTS|9|25|Ученики же ночью, взяв его, спустили по стене в корзине.
ACTS|9|26|Савл прибыл в Иерусалим и старался пристать к ученикам; но все боялись его, не веря, что он ученик.
ACTS|9|27|Варнава же, взяв его, пришел к Апостолам и рассказал им, как на пути он видел Господа, и что говорил ему Господь, и как он в Дамаске смело проповедывал во имя Иисуса.
ACTS|9|28|И пребывал он с ними, входя и исходя, в Иерусалиме, и смело проповедывал во имя Господа Иисуса.
ACTS|9|29|Говорил также и состязался с Еллинистами; а они покушались убить его.
ACTS|9|30|Братия, узнав [о сем], отправили его в Кесарию и препроводили в Тарс.
ACTS|9|31|Церкви же по всей Иудее, Галилее и Самарии были в покое, назидаясь и ходя в страхе Господнем; и, при утешении от Святаго Духа, умножались.
ACTS|9|32|Случилось, что Петр, обходя всех, пришел и к святым, живущим в Лидде.
ACTS|9|33|Там нашел он одного человека, именем Энея, который восемь уже лет лежал в постели в расслаблении.
ACTS|9|34|Петр сказал ему: Эней! исцеляет тебя Иисус Христос; встань с постели твоей. И он тотчас встал.
ACTS|9|35|И видели его все, живущие в Лидде и в Сароне, которые и обратились к Господу.
ACTS|9|36|В Иоппии находилась одна ученица, именем Тавифа, что значит: "серна"; она была исполнена добрых дел и творила много милостынь.
ACTS|9|37|Случилось в те дни, что она занемогла и умерла. Ее омыли и положили в горнице.
ACTS|9|38|А как Лидда была близ Иоппии, то ученики, услышав, что Петр находится там, послали к нему двух человек просить, чтобы он не замедлил придти к ним.
ACTS|9|39|Петр, встав, пошел с ними; и когда он прибыл, ввели его в горницу, и все вдовицы со слезами предстали перед ним, показывая рубашки и платья, какие делала Серна, живя с ними.
ACTS|9|40|Петр выслал всех вон и, преклонив колени, помолился, и, обратившись к телу, сказал: Тавифа! встань. И она открыла глаза свои и, увидев Петра, села.
ACTS|9|41|Он, подав ей руку, поднял ее, и, призвав святых и вдовиц, поставил ее перед ними живою.
ACTS|9|42|Это сделалось известным по всей Иоппии, и многие уверовали в Господа.
ACTS|9|43|И довольно дней пробыл он в Иоппии у некоторого Симона кожевника.
ACTS|10|1|В Кесарии был некоторый муж, именем Корнилий, сотник из полка, называемого Италийским,
ACTS|10|2|благочестивый и боящийся Бога со всем домом своим, творивший много милостыни народу и всегда молившийся Богу.
ACTS|10|3|Он в видении ясно видел около девятого часа дня Ангела Божия, который вошел к нему и сказал ему: Корнилий!
ACTS|10|4|Он же, взглянув на него и испугавшись, сказал: что, Господи? [Ангел] отвечал ему: молитвы твои и милостыни твои пришли на память пред Богом.
ACTS|10|5|Итак пошли людей в Иоппию и призови Симона, называемого Петром.
ACTS|10|6|Он гостит у некоего Симона кожевника, которого дом находится при море; он скажет тебе слова, которыми спасешься ты и весь дом твой.
ACTS|10|7|Когда Ангел, говоривший с Корнилием, отошел, то он, призвав двоих из своих слуг и благочестивого воина из находившихся при нем
ACTS|10|8|и, рассказав им все, послал их в Иоппию.
ACTS|10|9|На другой день, когда они шли и приближались к городу, Петр около шестого часа взошел на верх дома помолиться.
ACTS|10|10|И почувствовал он голод, и хотел есть. Между тем, как приготовляли, он пришел в исступление
ACTS|10|11|и видит отверстое небо и сходящий к нему некоторый сосуд, как бы большое полотно, привязанное за четыре угла и опускаемое на землю;
ACTS|10|12|в нем находились всякие четвероногие земные, звери, пресмыкающиеся и птицы небесные.
ACTS|10|13|И был глас к нему: встань, Петр, заколи и ешь.
ACTS|10|14|Но Петр сказал: нет, Господи, я никогда не ел ничего скверного или нечистого.
ACTS|10|15|Тогда в другой раз [был] глас к нему: что Бог очистил, того ты не почитай нечистым.
ACTS|10|16|Это было трижды; и сосуд опять поднялся на небо.
ACTS|10|17|Когда же Петр недоумевал в себе, что бы значило видение, которое он видел, – вот, мужи, посланные Корнилием, расспросив о доме Симона, остановились у ворот,
ACTS|10|18|и, крикнув, спросили: здесь ли Симон, называемый Петром?
ACTS|10|19|Между тем, как Петр размышлял о видении, Дух сказал ему: вот, три человека ищут тебя;
ACTS|10|20|встань, сойди и иди с ними, нимало не сомневаясь; ибо Я послал их.
ACTS|10|21|Петр, сойдя к людям, присланным к нему от Корнилия, сказал: я тот, которого вы ищете; за каким делом пришли вы?
ACTS|10|22|Они же сказали: Корнилий сотник, муж добродетельный и боящийся Бога, одобряемый всем народом Иудейским, получил от святаго Ангела повеление призвать тебя в дом свой и послушать речей твоих.
ACTS|10|23|Тогда Петр, пригласив их, угостил. А на другой день, встав, пошел с ними, и некоторые из братий Иоппийских пошли с ним.
ACTS|10|24|В следующий день пришли они в Кесарию. Корнилий же ожидал их, созвав родственников своих и близких друзей.
ACTS|10|25|Когда Петр входил, Корнилий встретил его и поклонился, пав к ногам его.
ACTS|10|26|Петр же поднял его, говоря: встань; я тоже человек.
ACTS|10|27|И, беседуя с ним, вошел [в дом], и нашел многих собравшихся.
ACTS|10|28|И сказал им: вы знаете, что Иудею возбранено сообщаться или сближаться с иноплеменником; но мне Бог открыл, чтобы я не почитал ни одного человека скверным или нечистым.
ACTS|10|29|Посему я, будучи позван, и пришел беспрекословно. Итак спрашиваю: для какого дела вы призвали меня?
ACTS|10|30|Корнилий сказал: четвертого дня я постился до теперешнего часа, и в девятом часу молился в своем доме, и вот, стал предо мною муж в светлой одежде,
ACTS|10|31|и говорит: Корнилий! услышана молитва твоя, и милостыни твои воспомянулись пред Богом.
ACTS|10|32|Итак пошли в Иоппию и призови Симона, называемого Петром; он гостит в доме кожевника Симона при море; он придет и скажет тебе.
ACTS|10|33|Тотчас послал я к тебе, и ты хорошо сделал, что пришел. Теперь все мы предстоим пред Богом, чтобы выслушать все, что повелено тебе от Бога.
ACTS|10|34|Петр отверз уста и сказал: истинно познаю, что Бог нелицеприятен,
ACTS|10|35|но во всяком народе боящийся Его и поступающий по правде приятен Ему.
ACTS|10|36|Он послал сынам Израилевым слово, благовествуя мир чрез Иисуса Христа; Сей есть Господь всех.
ACTS|10|37|Вы знаете происходившее по всей Иудее, начиная от Галилеи, после крещения, проповеданного Иоанном:
ACTS|10|38|как Бог Духом Святым и силою помазал Иисуса из Назарета, и Он ходил, благотворя и исцеляя всех, обладаемых диаволом, потому что Бог был с Ним.
ACTS|10|39|И мы свидетели всего, что сделал Он в стране Иудейской и в Иерусалиме, и что наконец Его убили, повесив на древе.
ACTS|10|40|Сего Бог воскресил в третий день, и дал Ему являться
ACTS|10|41|не всему народу, но свидетелям, предъизбранным от Бога, нам, которые с Ним ели и пили, по воскресении Его из мертвых.
ACTS|10|42|И Он повелел нам проповедывать людям и свидетельствовать, что Он есть определенный от Бога Судия живых и мертвых.
ACTS|10|43|О Нем все пророки свидетельствуют, что всякий верующий в Него получит прощение грехов именем Его.
ACTS|10|44|Когда Петр еще продолжал эту речь, Дух Святый сошел на всех, слушавших слово.
ACTS|10|45|И верующие из обрезанных, пришедшие с Петром, изумились, что дар Святаго Духа излился и на язычников,
ACTS|10|46|ибо слышали их говорящих языками и величающих Бога. Тогда Петр сказал:
ACTS|10|47|кто может запретить креститься водою тем, которые, как и мы, получили Святаго Духа?
ACTS|10|48|И велел им креститься во имя Иисуса Христа. Потом они просили его пробыть у них несколько дней.
ACTS|11|1|Услышали Апостолы и братия, бывшие в Иудее, что и язычники приняли слово Божие.
ACTS|11|2|И когда Петр пришел в Иерусалим, обрезанные упрекали его,
ACTS|11|3|говоря: ты ходил к людям необрезанным и ел с ними.
ACTS|11|4|Петр же начал пересказывать им по порядку, говоря:
ACTS|11|5|в городе Иоппии я молился, и в исступлении видел видение: сходил некоторый сосуд, как бы большое полотно, за четыре угла спускаемое с неба, и спустилось ко мне.
ACTS|11|6|Я посмотрел в него и, рассматривая, увидел четвероногих земных, зверей, пресмыкающихся и птиц небесных.
ACTS|11|7|И услышал я голос, говорящий мне: встань, Петр, заколи и ешь.
ACTS|11|8|Я же сказал: нет, Господи, ничего скверного или нечистого никогда не входило в уста мои.
ACTS|11|9|И отвечал мне голос вторично с неба: что Бог очистил, того ты не почитай нечистым.
ACTS|11|10|Это было трижды, и опять поднялось все на небо.
ACTS|11|11|И вот, в тот самый час три человека стали перед домом, в котором я был, посланные из Кесарии ко мне.
ACTS|11|12|Дух сказал мне, чтобы я шел с ними, нимало не сомневаясь. Пошли со мною и сии шесть братьев, и мы пришли в дом [того] человека.
ACTS|11|13|Он рассказал нам, как он видел в доме своем Ангела святого, который стал и сказал ему: пошли в Иоппию людей и призови Симона, называемого Петром;
ACTS|11|14|он скажет тебе слова, которыми спасешься ты и весь дом твой.
ACTS|11|15|Когда же начал я говорить, сошел на них Дух Святый, как и на нас вначале.
ACTS|11|16|Тогда вспомнил я слово Господа, как Он говорил: "Иоанн крестил водою, а вы будете крещены Духом Святым".
ACTS|11|17|Итак, если Бог дал им такой же дар, как и нам, уверовавшим в Господа Иисуса Христа, то кто же я, чтобы мог воспрепятствовать Богу?
ACTS|11|18|Выслушав это, они успокоились и прославили Бога, говоря: видно, и язычникам дал Бог покаяние в жизнь.
ACTS|11|19|Между тем рассеявшиеся от гонения, бывшего после Стефана, прошли до Финикии и Кипра и Антиохии, никому не проповедуя слово, кроме Иудеев.
ACTS|11|20|Были же некоторые из них Кипряне и Киринейцы, которые, придя в Антиохию, говорили Еллинам, благовествуя Господа Иисуса.
ACTS|11|21|И была рука Господня с ними, и великое число, уверовав, обратилось к Господу.
ACTS|11|22|Дошел слух о сем до церкви Иерусалимской, и поручили Варнаве идти в Антиохию.
ACTS|11|23|Он, прибыв и увидев благодать Божию, возрадовался и убеждал всех держаться Господа искренним сердцем;
ACTS|11|24|ибо он был муж добрый и исполненный Духа Святаго и веры. И приложилось довольно народа к Господу.
ACTS|11|25|Потом Варнава пошел в Тарс искать Савла и, найдя его, привел в Антиохию.
ACTS|11|26|Целый год собирались они в церкви и учили немалое число людей, и ученики в Антиохии в первый раз стали называться Христианами.
ACTS|11|27|В те дни пришли из Иерусалима в Антиохию пророки.
ACTS|11|28|И один из них, по имени Агав, встав, предвозвестил Духом, что по всей вселенной будет великий голод, который и был при кесаре Клавдии.
ACTS|11|29|Тогда ученики положили, каждый по достатку своему, послать пособие братьям, живущим в Иудее,
ACTS|11|30|что и сделали, послав [собранное] к пресвитерам через Варнаву и Савла.
ACTS|12|1|В то время царь Ирод поднял руки на некоторых из принадлежащих к церкви, чтобы сделать им зло,
ACTS|12|2|и убил Иакова, брата Иоаннова, мечом.
ACTS|12|3|Видя же, что это приятно Иудеям, вслед за тем взял и Петра, – тогда были дни опресноков, –
ACTS|12|4|и, задержав его, посадил в темницу, и приказал четырем четверицам воинов стеречь его, намереваясь после Пасхи вывести его к народу.
ACTS|12|5|Итак Петра стерегли в темнице, между тем церковь прилежно молилась о нем Богу.
ACTS|12|6|Когда же Ирод хотел вывести его, в ту ночь Петр спал между двумя воинами, скованный двумя цепями, и стражи у дверей стерегли темницу.
ACTS|12|7|И вот, Ангел Господень предстал, и свет осиял темницу. [Ангел], толкнув Петра в бок, пробудил его и сказал: встань скорее. И цепи упали с рук его.
ACTS|12|8|И сказал ему Ангел: опояшься и обуйся. Он сделал так. Потом говорит ему: надень одежду твою и иди за мною.
ACTS|12|9|[Петр] вышел и следовал за ним, не зная, что делаемое Ангелом было действительно, а думая, что видит видение.
ACTS|12|10|Пройдя первую и вторую стражу, они пришли к железным воротам, ведущим в город, которые сами собою отворились им: они вышли, и прошли одну улицу, и вдруг Ангела не стало с ним.
ACTS|12|11|Тогда Петр, придя в себя, сказал: теперь я вижу воистину, что Господь послал Ангела Своего и избавил меня из руки Ирода и от всего, чего ждал народ Иудейский.
ACTS|12|12|И, осмотревшись, пришел к дому Марии, матери Иоанна, называемого Марком, где многие собрались и молились.
ACTS|12|13|Когда же Петр постучался у ворот, то вышла послушать служанка, именем Рода,
ACTS|12|14|и, узнав голос Петра, от радости не отворила ворот, но, вбежав, объявила, что Петр стоит у ворот.
ACTS|12|15|А те сказали ей: в своем ли ты уме? Но она утверждала свое. Они же говорили: это Ангел его.
ACTS|12|16|Между тем Петр продолжал стучать. Когда же отворили, то увидели его и изумились.
ACTS|12|17|Он же, дав знак рукою, чтобы молчали, рассказал им, как Господь вывел его из темницы, и сказал: уведомьте о сем Иакова и братьев. Потом, выйдя, пошел в другое место.
ACTS|12|18|По наступлении дня между воинами сделалась большая тревога о том, что сделалось с Петром.
ACTS|12|19|Ирод же, поискав его и не найдя, судил стражей и велел казнить их. Потом он отправился из Иудеи в Кесарию и [там] оставался.
ACTS|12|20|Ирод был раздражен на Тирян и Сидонян; они же, согласившись, пришли к нему и, склонив на свою сторону Власта, постельника царского, просили мира, потому что область их питалась от [области] царской.
ACTS|12|21|В назначенный день Ирод, одевшись в царскую одежду, сел на возвышенном месте и говорил к ним;
ACTS|12|22|а народ восклицал: [это] голос Бога, а не человека.
ACTS|12|23|Но вдруг Ангел Господень поразил его за то, что он не воздал славы Богу; и он, быв изъеден червями, умер.
ACTS|12|24|Слово же Божие росло и распространялось.
ACTS|12|25|А Варнава и Савл, по исполнении поручения, возвратились из Иерусалима в Антиохию, взяв с собою и Иоанна, прозванного Марком.
ACTS|13|1|В Антиохии, в тамошней церкви были некоторые пророки и учители: Варнава, и Симеон, называемый Нигер, и Луций Киринеянин, и Манаил, совоспитанник Ирода четвертовластника, и Савл.
ACTS|13|2|Когда они служили Господу и постились, Дух Святый сказал: отделите Мне Варнаву и Савла на дело, к которому Я призвал их.
ACTS|13|3|Тогда они, совершив пост и молитву и возложив на них руки, отпустили их.
ACTS|13|4|Сии, быв посланы Духом Святым, пришли в Селевкию, а оттуда отплыли в Кипр;
ACTS|13|5|и, быв в Саламине, проповедывали слово Божие в синагогах Иудейских; имели же при себе и Иоанна для служения.
ACTS|13|6|Пройдя весь остров до Пафа, нашли они некоторого волхва, лжепророка, Иудеянина, именем Вариисуса,
ACTS|13|7|который находился с проконсулом Сергием Павлом, мужем разумным. Сей, призвав Варнаву и Савла, пожелал услышать слово Божие.
ACTS|13|8|А Елима волхв ибо то значит имя его противился им, стараясь отвратить проконсула от веры.
ACTS|13|9|Но Савл, он же и Павел, исполнившись Духа Святаго и устремив на него взор,
ACTS|13|10|сказал: о, исполненный всякого коварства и всякого злодейства, сын диавола, враг всякой правды! перестанешь ли ты совращать с прямых путей Господних?
ACTS|13|11|И ныне вот, рука Господня на тебя: ты будешь слеп и не увидишь солнца до времени. И вдруг напал на него мрак и тьма, и он, обращаясь туда и сюда, искал вожатого.
ACTS|13|12|Тогда проконсул, увидев происшедшее, уверовал, дивясь учению Господню.
ACTS|13|13|Отплыв из Пафа, Павел и бывшие при нем прибыли в Пергию, в Памфилии. Но Иоанн, отделившись от них, возвратился в Иерусалим.
ACTS|13|14|Они же, проходя от Пергии, прибыли в Антиохию Писидийскую и, войдя в синагогу в день субботний, сели.
ACTS|13|15|После чтения закона и пророков, начальники синагоги послали сказать им: мужи братия! если у вас есть слово наставления к народу, говорите.
ACTS|13|16|Павел, встав и дав знак рукою, сказал: мужи Израильтяне и боящиеся Бога! послушайте.
ACTS|13|17|Бог народа сего избрал отцов наших и возвысил сей народ во время пребывания в земле Египетской, и мышцею вознесенною вывел их из нее,
ACTS|13|18|и около сорока лет времени питал их в пустыне.
ACTS|13|19|И, истребив семь народов в земле Ханаанской, разделил им в наследие землю их.
ACTS|13|20|И после сего, около четырехсот пятидесяти лет, давал им судей до пророка Самуила.
ACTS|13|21|Потом просили они царя, и Бог дал им Саула, сына Кисова, мужа из колена Вениаминова. [Так прошло] лет сорок.
ACTS|13|22|Отринув его, поставил им царем Давида, о котором и сказал, свидетельствуя: нашел Я мужа по сердцу Моему, Давида, сына Иессеева, который исполнит все хотения Мои.
ACTS|13|23|Из его–то потомства Бог по обетованию воздвиг Израилю Спасителя Иисуса.
ACTS|13|24|Перед самым явлением Его Иоанн проповедывал крещение покаяния всему народу Израильскому.
ACTS|13|25|При окончании же поприща своего, Иоанн говорил: за кого почитаете вы меня? я не тот; но вот, идет за мною, у Которого я недостоин развязать обувь на ногах.
ACTS|13|26|Мужи братия, дети рода Авраамова, и боящиеся Бога между вами! вам послано слово спасения сего.
ACTS|13|27|Ибо жители Иерусалима и начальники их, не узнав Его и осудив, исполнили слова пророческие, читаемые каждую субботу,
ACTS|13|28|и, не найдя в Нем никакой вины, достойной смерти, просили Пилата убить Его.
ACTS|13|29|Когда же исполнили все написанное о Нем, то, сняв с древа, положили Его во гроб.
ACTS|13|30|Но Бог воскресил Его из мертвых.
ACTS|13|31|Он в продолжение многих дней являлся тем, которые вышли с Ним из Галилеи в Иерусалим и которые ныне суть свидетели Его перед народом.
ACTS|13|32|И мы благовествуем вам, что обетование, данное отцам, Бог исполнил нам, детям их, воскресив Иисуса,
ACTS|13|33|как и во втором псалме написано: Ты Сын Мой: Я ныне родил Тебя.
ACTS|13|34|А что воскресил Его из мертвых, так что Он уже не обратится в тление, [о сем] сказал так: Я дам вам милости, [обещанные] Давиду, верно.
ACTS|13|35|Посему и в другом [месте] говорит: не дашь Святому Твоему увидеть тление.
ACTS|13|36|Давид, в свое время послужив изволению Божию, почил и приложился к отцам своим, и увидел тление;
ACTS|13|37|а Тот, Которого Бог воскресил, не увидел тления.
ACTS|13|38|Итак, да будет известно вам, мужи братия, что ради Него возвещается вам прощение грехов;
ACTS|13|39|и во всем, в чем вы не могли оправдаться законом Моисеевым, оправдывается Им всякий верующий.
ACTS|13|40|Берегитесь же, чтобы не пришло на вас сказанное у пророков:
ACTS|13|41|смотрите, презрители, подивитесь и исчезните; ибо Я делаю дело во дни ваши, дело, которому не поверили бы вы, если бы кто рассказывал вам.
ACTS|13|42|При выходе их из Иудейской синагоги язычники просили их говорить о том же в следующую субботу.
ACTS|13|43|Когда же собрание было распущено, то многие Иудеи и чтители [Бога], обращенные из язычников, последовали за Павлом и Варнавою, которые, беседуя с ними, убеждали их пребывать в благодати Божией.
ACTS|13|44|В следующую субботу почти весь город собрался слушать слово Божие.
ACTS|13|45|Но Иудеи, увидев народ, исполнились зависти и, противореча и злословя, сопротивлялись тому, что говорил Павел.
ACTS|13|46|Тогда Павел и Варнава с дерзновением сказали: вам первым надлежало быть проповедану слову Божию, но как вы отвергаете его и сами себя делаете недостойными вечной жизни, то вот, мы обращаемся к язычникам.
ACTS|13|47|Ибо так заповедал нам Господь: Я положил Тебя во свет язычникам, чтобы Ты был во спасение до края земли.
ACTS|13|48|Язычники, слыша это, радовались и прославляли слово Господне, и уверовали все, которые были предуставлены к вечной жизни.
ACTS|13|49|И слово Господне распространялось по всей стране.
ACTS|13|50|Но Иудеи, подстрекнув набожных и почетных женщин и первых в городе [людей], воздвигли гонение на Павла и Варнаву и изгнали их из своих пределов.
ACTS|13|51|Они же, отрясши на них прах от ног своих, пошли в Иконию.
ACTS|13|52|А ученики исполнялись радости и Духа Святаго.
ACTS|14|1|В Иконии они вошли вместе в Иудейскую синагогу и говорили так, что уверовало великое множество Иудеев и Еллинов.
ACTS|14|2|А неверующие Иудеи возбудили и раздражили против братьев сердца язычников.
ACTS|14|3|Впрочем они пробыли [здесь] довольно времени, смело действуя о Господе, Который, во свидетельство слову благодати Своей, творил руками их знамения и чудеса.
ACTS|14|4|Между тем народ в городе разделился: и одни были на стороне Иудеев, а другие на стороне Апостолов.
ACTS|14|5|Когда же язычники и Иудеи со своими начальниками устремились на них, чтобы посрамить и побить их камнями,
ACTS|14|6|они, узнав [о сем], удалились в Ликаонские города Листру и Дервию и в окрестности их,
ACTS|14|7|и там благовествовали.
ACTS|14|8|В Листре некоторый муж, не владевший ногами, сидел, будучи хром от чрева матери своей, и никогда не ходил.
ACTS|14|9|Он слушал говорившего Павла, который, взглянув на него и увидев, что он имеет веру для получения исцеления,
ACTS|14|10|сказал громким голосом: тебе говорю во имя Господа Иисуса Христа: стань на ноги твои прямо. И он тотчас вскочил и стал ходить.
ACTS|14|11|Народ же, увидев, что сделал Павел, возвысил свой голос, говоря по–ликаонски: боги в образе человеческом сошли к нам.
ACTS|14|12|И называли Варнаву Зевсом, а Павла Ермием, потому что он начальствовал в слове.
ACTS|14|13|Жрец же [идола] Зевса, находившегося перед их городом, приведя к воротам волов и [принеся] венки, хотел вместе с народом совершить жертвоприношение.
ACTS|14|14|Но Апостолы Варнава и Павел, услышав [о сем], разодрали свои одежды и, бросившись в народ, громогласно говорили:
ACTS|14|15|мужи! что вы это делаете? И мы – подобные вам человеки, и благовествуем вам, чтобы вы обратились от сих ложных к Богу Живому, Который сотворил небо и землю, и море, и все, что в них,
ACTS|14|16|Который в прошедших родах попустил всем народам ходить своими путями,
ACTS|14|17|хотя и не переставал свидетельствовать о Себе благодеяниями, подавая нам с неба дожди и времена плодоносные и исполняя пищею и веселием сердца наши.
ACTS|14|18|И, говоря сие, они едва убедили народ не приносить им жертвы и идти каждому домой. Между тем, как они, оставаясь там, учили,
ACTS|14|19|из Антиохии и Иконии пришли некоторые Иудеи и, когда [Апостолы] смело проповедывали, убедили народ отстать от них, говоря: они не говорят ничего истинного, а все лгут. И, возбудив народ, побили Павла камнями и вытащили за город, почитая его умершим.
ACTS|14|20|Когда же ученики собрались около него, он встал и пошел в город, а на другой день удалился с Варнавою в Дервию.
ACTS|14|21|Проповедав Евангелие сему городу и приобретя довольно учеников, они обратно проходили Листру, Иконию и Антиохию,
ACTS|14|22|утверждая души учеников, увещевая пребывать в вере и [поучая], что многими скорбями надлежит нам войти в Царствие Божие.
ACTS|14|23|Рукоположив же им пресвитеров к каждой церкви, они помолились с постом и предали их Господу, в Которого уверовали.
ACTS|14|24|Потом, пройдя через Писидию, пришли в Памфилию,
ACTS|14|25|и, проповедав слово Господне в Пергии, сошли в Атталию;
ACTS|14|26|а оттуда отплыли в Антиохию, откуда были преданы благодати Божией на дело, которое и исполнили.
ACTS|14|27|Прибыв туда и собрав церковь, они рассказали все, что сотворил Бог с ними и как Он отверз дверь веры язычникам.
ACTS|14|28|И пребывали там немалое время с учениками.
ACTS|15|1|Некоторые, пришедшие из Иудеи, учили братьев: если не обрежетесь по обряду Моисееву, не можете спастись.
ACTS|15|2|Когда же произошло разногласие и немалое состязание у Павла и Варнавы с ними, то положили Павлу и Варнаве и некоторым другим из них отправиться по сему делу к Апостолам и пресвитерам в Иерусалим.
ACTS|15|3|Итак, быв провожены церковью, они проходили Финикию и Самарию, рассказывая об обращении язычников, и производили радость великую во всех братиях.
ACTS|15|4|По прибытии же в Иерусалим они были приняты церковью, Апостолами и пресвитерами, и возвестили все, что Бог сотворил с ними и как отверз дверь веры язычникам.
ACTS|15|5|Тогда восстали некоторые из фарисейской ереси уверовавшие и говорили, что должно обрезывать [язычников] и заповедывать соблюдать закон Моисеев.
ACTS|15|6|Апостолы и пресвитеры собрались для рассмотрения сего дела.
ACTS|15|7|По долгом рассуждении Петр, встав, сказал им: мужи братия! вы знаете, что Бог от дней первых избрал из нас [меня], чтобы из уст моих язычники услышали слово Евангелия и уверовали;
ACTS|15|8|и Сердцеведец Бог дал им свидетельство, даровав им Духа Святаго, как и нам;
ACTS|15|9|и не положил никакого различия между нами и ими, верою очистив сердца их.
ACTS|15|10|Что же вы ныне искушаете Бога, [желая] возложить на выи учеников иго, которого не могли понести ни отцы наши, ни мы?
ACTS|15|11|Но мы веруем, что благодатию Господа Иисуса Христа спасемся, как и они.
ACTS|15|12|Тогда умолкло все собрание и слушало Варнаву и Павла, рассказывавших, какие знамения и чудеса сотворил Бог через них среди язычников.
ACTS|15|13|После же того, как они умолкли, начал речь Иаков и сказал: мужи братия! послушайте меня.
ACTS|15|14|Симон изъяснил, как Бог первоначально призрел на язычников, чтобы составить из них народ во имя Свое.
ACTS|15|15|И с сим согласны слова пророков, как написано:
ACTS|15|16|Потом обращусь и воссоздам скинию Давидову падшую, и то, что в ней разрушено, воссоздам, и исправлю ее,
ACTS|15|17|чтобы взыскали Господа прочие человеки и все народы, между которыми возвестится имя Мое, говорит Господь, творящий все сие.
ACTS|15|18|Ведомы Богу от вечности все дела Его.
ACTS|15|19|Посему я полагаю не затруднять обращающихся к Богу из язычников,
ACTS|15|20|а написать им, чтобы они воздерживались от оскверненного идолами, от блуда, удавленины и крови, и чтобы не делали другим того, чего не хотят себе.
ACTS|15|21|Ибо [закон] Моисеев от древних родов по всем городам имеет проповедующих его и читается в синагогах каждую субботу.
ACTS|15|22|Тогда Апостолы и пресвитеры со всею церковью рассудили, избрав из среды себя мужей, послать их в Антиохию с Павлом и Варнавою, [именно]: Иуду, прозываемого Варсавою, и Силу, мужей, начальствующих между братиями,
ACTS|15|23|написав и вручив им следующее: "Апостолы и пресвитеры и братия – находящимся в Антиохии, Сирии и Киликии братиям из язычников: радоваться.
ACTS|15|24|Поелику мы услышали, что некоторые, вышедшие от нас, смутили вас [своими] речами и поколебали ваши души, говоря, что должно обрезываться и соблюдать закон, чего мы им не поручали,
ACTS|15|25|то мы, собравшись, единодушно рассудили, избрав мужей, послать их к вам с возлюбленными нашими Варнавою и Павлом,
ACTS|15|26|человеками, предавшими души свои за имя Господа нашего Иисуса Христа.
ACTS|15|27|Итак мы послали Иуду и Силу, которые изъяснят вам то же и словесно.
ACTS|15|28|Ибо угодно Святому Духу и нам не возлагать на вас никакого бремени более, кроме сего необходимого:
ACTS|15|29|воздерживаться от идоложертвенного и крови, и удавленины, и блуда, и не делать другим того, чего себе не хотите. Соблюдая сие, хорошо сделаете. Будьте здравы".
ACTS|15|30|Итак, отправленные пришли в Антиохию и, собрав людей, вручили письмо.
ACTS|15|31|Они же, прочитав, возрадовались о сем наставлении.
ACTS|15|32|Иуда и Сила, будучи также пророками, обильным словом преподали наставление братиям и утвердили их.
ACTS|15|33|Пробыв там [некоторое] время, они с миром отпущены были братиями к Апостолам.
ACTS|15|34|Но Силе рассудилось остаться там. (А Иуда возвратился в Иерусалим.)
ACTS|15|35|Павел же и Варнава жили в Антиохии, уча и благовествуя, вместе с другими многими, слово Господне.
ACTS|15|36|По некотором времени Павел сказал Варнаве: пойдем опять, посетим братьев наших по всем городам, в которых мы проповедали слово Господне, как они живут.
ACTS|15|37|Варнава хотел взять с собою Иоанна, называемого Марком.
ACTS|15|38|Но Павел полагал не брать отставшего от них в Памфилии и не шедшего с ними на дело, на которое они были посланы.
ACTS|15|39|Отсюда произошло огорчение, так что они разлучились друг с другом; и Варнава, взяв Марка, отплыл в Кипр;
ACTS|15|40|а Павел, избрав себе Силу, отправился, быв поручен братиями благодати Божией,
ACTS|15|41|и проходил Сирию и Киликию, утверждая церкви.
ACTS|16|1|Дошел он до Дервии и Листры. И вот, там был некоторый ученик, именем Тимофей, которого мать была Иудеянка уверовавшая, а отец Еллин,
ACTS|16|2|и о котором свидетельствовали братия, находившиеся в Листре и Иконии.
ACTS|16|3|Его пожелал Павел взять с собою; и, взяв, обрезал его ради Иудеев, находившихся в тех местах; ибо все знали об отце его, что он был Еллин.
ACTS|16|4|Проходя же по городам, они предавали [верным] соблюдать определения, постановленные Апостолами и пресвитерами в Иерусалиме.
ACTS|16|5|И церкви утверждались верою и ежедневно увеличивались числом.
ACTS|16|6|Пройдя через Фригию и Галатийскую страну, они не были допущены Духом Святым проповедывать слово в Асии.
ACTS|16|7|Дойдя до Мисии, предпринимали идти в Вифинию; но Дух не допустил их.
ACTS|16|8|Миновав же Мисию, сошли они в Троаду.
ACTS|16|9|И было ночью видение Павлу: предстал некий муж, Македонянин, прося его и говоря: приди в Македонию и помоги нам.
ACTS|16|10|После сего видения, тотчас мы положили отправиться в Македонию, заключая, что призывал нас Господь благовествовать там.
ACTS|16|11|Итак, отправившись из Троады, мы прямо прибыли в Самофракию, а на другой день в Неаполь,
ACTS|16|12|оттуда же в Филиппы: это первый город в той части Македонии, колония. В этом городе мы пробыли несколько дней.
ACTS|16|13|В день же субботний мы вышли за город к реке, где, по обыкновению, был молитвенный дом, и, сев, разговаривали с собравшимися [там] женщинами.
ACTS|16|14|И одна женщина из города Фиатир, именем Лидия, торговавшая багряницею, чтущая Бога, слушала; и Господь отверз сердце ее внимать тому, что говорил Павел.
ACTS|16|15|Когда же крестилась она и домашние ее, то просила нас, говоря: если вы признали меня верною Господу, то войдите в дом мой и живите [у] [меня]. И убедила нас.
ACTS|16|16|Случилось, что, когда мы шли в молитвенный дом, встретилась нам одна служанка, одержимая духом прорицательным, которая через прорицание доставляла большой доход господам своим.
ACTS|16|17|Идя за Павлом и за нами, она кричала, говоря: сии человеки – рабы Бога Всевышнего, которые возвещают нам путь спасения.
ACTS|16|18|Это она делала много дней. Павел, вознегодовав, обратился и сказал духу: именем Иисуса Христа повелеваю тебе выйти из нее. И [дух] вышел в тот же час.
ACTS|16|19|Тогда господа ее, видя, что исчезла надежда дохода их, схватили Павла и Силу и повлекли на площадь к начальникам.
ACTS|16|20|И, приведя их к воеводам, сказали: сии люди, будучи Иудеями, возмущают наш город
ACTS|16|21|и проповедуют обычаи, которых нам, Римлянам, не следует ни принимать, ни исполнять.
ACTS|16|22|Народ также восстал на них, а воеводы, сорвав с них одежды, велели бить их палками
ACTS|16|23|и, дав им много ударов, ввергли в темницу, приказав темничному стражу крепко стеречь их.
ACTS|16|24|Получив такое приказание, он ввергнул их во внутреннюю темницу и ноги их забил в колоду.
ACTS|16|25|Около полуночи Павел и Сила, молясь, воспевали Бога; узники же слушали их.
ACTS|16|26|Вдруг сделалось великое землетрясение, так что поколебалось основание темницы; тотчас отворились все двери, и у всех узы ослабели.
ACTS|16|27|Темничный же страж, пробудившись и увидев, что двери темницы отворены, извлек меч и хотел умертвить себя, думая, что узники убежали.
ACTS|16|28|Но Павел возгласил громким голосом, говоря: не делай себе никакого зла, ибо все мы здесь.
ACTS|16|29|Он потребовал огня, вбежал [в темницу] и в трепете припал к Павлу и Силе,
ACTS|16|30|и, выведя их вон, сказал: государи [мои]! что мне делать, чтобы спастись?
ACTS|16|31|Они же сказали: веруй в Господа Иисуса Христа, и спасешься ты и весь дом твой.
ACTS|16|32|И проповедали слово Господне ему и всем, бывшим в доме его.
ACTS|16|33|И, взяв их в тот час ночи, он омыл раны их и немедленно крестился сам и все [домашние] его.
ACTS|16|34|И, приведя их в дом свой, предложил трапезу и возрадовался со всем домом своим, что уверовал в Бога.
ACTS|16|35|Когда же настал день, воеводы послали городских служителей сказать: отпусти тех людей.
ACTS|16|36|Темничный страж объявил о сем Павлу: воеводы прислали отпустить вас; итак выйдите теперь и идите с миром.
ACTS|16|37|Но Павел сказал к ним: нас, Римских граждан, без суда всенародно били и бросили в темницу, а теперь тайно выпускают? нет, пусть придут и сами выведут нас.
ACTS|16|38|Городские служители пересказали эти слова воеводам, и те испугались, услышав, что это Римские граждане.
ACTS|16|39|И, придя, извинились перед ними и, выведя, просили удалиться из города.
ACTS|16|40|Они же, выйдя из темницы, пришли к Лидии и, увидев братьев, поучали их, и отправились.
ACTS|17|1|Пройдя через Амфиполь и Аполлонию, они пришли в Фессалонику, где была Иудейская синагога.
ACTS|17|2|Павел, по своему обыкновению, вошел к ним и три субботы говорил с ними из Писаний,
ACTS|17|3|открывая и доказывая им, что Христу надлежало пострадать и воскреснуть из мертвых и что Сей Христос есть Иисус, Которого я проповедую вам.
ACTS|17|4|И некоторые из них уверовали и присоединились к Павлу и Силе, как из Еллинов, чтущих [Бога], великое множество, так и из знатных женщин немало.
ACTS|17|5|Но неуверовавшие Иудеи, возревновав и взяв с площади некоторых негодных людей, собрались толпою и возмущали город и, приступив к дому Иасона, домогались вывести их к народу.
ACTS|17|6|Не найдя же их, повлекли Иасона и некоторых братьев к городским начальникам, крича, что эти всесветные возмутители пришли и сюда,
ACTS|17|7|а Иасон принял их, и все они поступают против повелений кесаря, почитая другого царем, Иисуса.
ACTS|17|8|И встревожили народ и городских начальников, слушавших это.
ACTS|17|9|Но [сии], получив удостоверение от Иасона и прочих, отпустили их.
ACTS|17|10|Братия же немедленно ночью отправили Павла и Силу в Верию, куда они прибыв, пошли в синагогу Иудейскую.
ACTS|17|11|Здешние были благомысленнее Фессалоникских: они приняли слово со всем усердием, ежедневно разбирая Писания, точно ли это так.
ACTS|17|12|И многие из них уверовали, и из Еллинских почетных женщин и из мужчин немало.
ACTS|17|13|Но когда Фессалоникские Иудеи узнали, что и в Верии проповедано Павлом слово Божие, то пришли и туда, возбуждая и возмущая народ.
ACTS|17|14|Тогда братия тотчас отпустили Павла, как будто идущего к морю; а Сила и Тимофей остались там.
ACTS|17|15|Сопровождавшие Павла проводили его до Афин и, получив приказание к Силе и Тимофею, чтобы они скорее пришли к нему, отправились.
ACTS|17|16|В ожидании их в Афинах Павел возмутился духом при виде этого города, полного идолов.
ACTS|17|17|Итак он рассуждал в синагоге с Иудеями и с чтущими [Бога], и ежедневно на площади со встречающимися.
ACTS|17|18|Некоторые из эпикурейских и стоических философов стали спорить с ним; и одни говорили: "что хочет сказать этот суеслов?", а другие: "кажется, он проповедует о чужих божествах", потому что он благовествовал им Иисуса и воскресение.
ACTS|17|19|И, взяв его, привели в ареопаг и говорили: можем ли мы знать, что это за новое учение, проповедуемое тобою?
ACTS|17|20|Ибо что–то странное ты влагаешь в уши наши. Посему хотим знать, что это такое?
ACTS|17|21|Афиняне же все и живущие [у них] иностранцы ни в чем охотнее не проводили время, как в том, чтобы говорить или слушать что – нибудь новое.
ACTS|17|22|И, став Павел среди ареопага, сказал: Афиняне! по всему вижу я, что вы как бы особенно набожны.
ACTS|17|23|Ибо, проходя и осматривая ваши святыни, я нашел и жертвенник, на котором написано "неведомому Богу". Сего–то, Которого вы, не зная, чтите, я проповедую вам.
ACTS|17|24|Бог, сотворивший мир и все, что в нем, Он, будучи Господом неба и земли, не в рукотворенных храмах живет
ACTS|17|25|и не требует служения рук человеческих, [как бы] имеющий в чем–либо нужду, Сам дая всему жизнь и дыхание и все.
ACTS|17|26|От одной крови Он произвел весь род человеческий для обитания по всему лицу земли, назначив предопределенные времена и пределы их обитанию,
ACTS|17|27|дабы они искали Бога, не ощутят ли Его и не найдут ли, хотя Он и недалеко от каждого из нас:
ACTS|17|28|ибо мы Им живем и движемся и существуем, как и некоторые из ваших стихотворцев говорили: "мы Его и род".
ACTS|17|29|Итак мы, будучи родом Божиим, не должны думать, что Божество подобно золоту, или серебру, или камню, получившему образ от искусства и вымысла человеческого.
ACTS|17|30|Итак, оставляя времена неведения, Бог ныне повелевает людям всем повсюду покаяться,
ACTS|17|31|ибо Он назначил день, в который будет праведно судить вселенную, посредством предопределенного Им Мужа, подав удостоверение всем, воскресив Его из мертвых.
ACTS|17|32|Услышав о воскресении мертвых, одни насмехались, а другие говорили: об этом послушаем тебя в другое время.
ACTS|17|33|Итак Павел вышел из среды их.
ACTS|17|34|Некоторые же мужи, пристав к нему, уверовали; между ними был Дионисий Ареопагит и женщина, именем Дамарь, и другие с ними.
ACTS|18|1|После сего Павел, оставив Афины, пришел в Коринф;
ACTS|18|2|И, нашед некоторого Иудея, именем Акилу, родом Понтянина, недавно пришедшего из Италии, и Прискиллу, жену его, – потому что Клавдий повелел всем Иудеям удалиться из Рима, – пришел к ним,
ACTS|18|3|и, по одинаковости ремесла, остался у них и работал; ибо ремеслом их было делание палаток.
ACTS|18|4|Во всякую же субботу он говорил в синагоге и убеждал Иудеев и Еллинов.
ACTS|18|5|А когда пришли из Македонии Сила и Тимофей, то Павел понуждаем был духом свидетельствовать Иудеям, что Иисус есть Христос.
ACTS|18|6|Но как они противились и злословили, то он, отрясши одежды свои, сказал к ним: кровь ваша на главах ваших; я чист; отныне иду к язычникам.
ACTS|18|7|И пошел оттуда, и пришел к некоторому чтущему Бога, именем Иусту, которого дом был подле синагоги.
ACTS|18|8|Крисп же, начальник синагоги, уверовал в Господа со всем домом своим, и многие из Коринфян, слушая, уверовали и крестились.
ACTS|18|9|Господь же в видении ночью сказал Павлу: не бойся, но говори и не умолкай,
ACTS|18|10|ибо Я с тобою, и никто не сделает тебе зла, потому что у Меня много людей в этом городе.
ACTS|18|11|И он оставался там год и шесть месяцев, поучая их слову Божию.
ACTS|18|12|Между тем, во время проконсульства Галлиона в Ахаии, напали Иудеи единодушно на Павла и привели его пред судилище,
ACTS|18|13|говоря, что он учит людей чтить Бога не по закону.
ACTS|18|14|Когда же Павел хотел открыть уста, Галлион сказал Иудеям: Иудеи! если бы какая–нибудь была обида или злой умысел, то я имел бы причину выслушать вас,
ACTS|18|15|но когда идет спор об учении и об именах и о законе вашем, то разбирайте сами; я не хочу быть судьею в этом.
ACTS|18|16|И прогнал их от судилища.
ACTS|18|17|А все Еллины, схватив Сосфена, начальника синагоги, били его перед судилищем; и Галлион нимало не беспокоился о том.
ACTS|18|18|Павел, пробыв еще довольно дней, простился с братиями и отплыл в Сирию, – и с ним Акила и Прискилла, – остригши голову в Кенхреях, по обету.
ACTS|18|19|Достигнув Ефеса, оставил их там, а сам вошел в синагогу и рассуждал с Иудеями.
ACTS|18|20|Когда же они просили его побыть у них долее, он не согласился,
ACTS|18|21|а простился с ними, сказав: мне нужно непременно провести приближающийся праздник в Иерусалиме; к вам же возвращусь опять, если будет угодно Богу. И отправился из Ефеса. (Акила же и Прискилла остались в Ефесе).
ACTS|18|22|Побывав в Кесарии, он приходил [в Иерусалим], приветствовал церковь и отошел в Антиохию.
ACTS|18|23|И, проведя [там] несколько времени, вышел, и проходил по порядку страну Галатийскую и Фригию, утверждая всех учеников.
ACTS|18|24|Некто Иудей, именем Аполлос, родом из Александрии, муж красноречивый и сведущий в Писаниях, пришел в Ефес.
ACTS|18|25|Он был наставлен в начатках пути Господня и, горя духом, говорил и учил о Господе правильно, зная только крещение Иоанново.
ACTS|18|26|Он начал смело говорить в синагоге. Услышав его, Акила и Прискилла приняли его и точнее объяснили ему путь Господень.
ACTS|18|27|А когда он вознамерился идти в Ахаию, то братия послали к [тамошним] ученикам, располагая их принять его; и он, прибыв туда, много содействовал уверовавшим благодатью,
ACTS|18|28|ибо он сильно опровергал Иудеев всенародно, доказывая Писаниями, что Иисус есть Христос.
ACTS|19|1|Во время пребывания Аполлоса в Коринфе Павел, пройдя верхние страны, прибыл в Ефес и, найдя [там] некоторых учеников,
ACTS|19|2|сказал им: приняли ли вы Святаго Духа, уверовав? Они же сказали ему: мы даже и не слыхали, есть ли Дух Святый.
ACTS|19|3|Он сказал им: во что же вы крестились? Они отвечали: во Иоанново крещение.
ACTS|19|4|Павел сказал: Иоанн крестил крещением покаяния, говоря людям, чтобы веровали в Грядущего по нем, то есть во Христа Иисуса.
ACTS|19|5|Услышав это, они крестились во имя Господа Иисуса,
ACTS|19|6|и, когда Павел возложил на них руки, нисшел на них Дух Святый, и они стали говорить [иными] языками и пророчествовать.
ACTS|19|7|Всех их было человек около двенадцати.
ACTS|19|8|Придя в синагогу, он небоязненно проповедывал три месяца, беседуя и удостоверяя о Царствии Божием.
ACTS|19|9|Но как некоторые ожесточились и не верили, злословя путь Господень перед народом, то он, оставив их, отделил учеников, и ежедневно проповедывал в училище некоего Тиранна.
ACTS|19|10|Это продолжалось до двух лет, так что все жители Асии слышали проповедь о Господе Иисусе, как Иудеи, так и Еллины.
ACTS|19|11|Бог же творил немало чудес руками Павла,
ACTS|19|12|так что на больных возлагали платки и опоясания с тела его, и у них прекращались болезни, и злые духи выходили из них.
ACTS|19|13|Даже некоторые из скитающихся Иудейских заклинателей стали употреблять над имеющими злых духов имя Господа Иисуса, говоря: заклинаем вас Иисусом, Которого Павел проповедует.
ACTS|19|14|Это делали какие–то семь сынов Иудейского первосвященника Скевы.
ACTS|19|15|Но злой дух сказал в ответ: Иисуса знаю, и Павел мне известен, а вы кто?
ACTS|19|16|И бросился на них человек, в котором был злой дух, и, одолев их, взял над ними такую силу, что они, нагие и избитые, выбежали из того дома.
ACTS|19|17|Это сделалось известно всем живущим в Ефесе Иудеям и Еллинам, и напал страх на всех их, и величаемо было имя Господа Иисуса.
ACTS|19|18|Многие же из уверовавших приходили, исповедуя и открывая дела свои.
ACTS|19|19|А из занимавшихся чародейством довольно многие, собрав книги свои, сожгли перед всеми, и сложили цены их, и оказалось их на пятьдесят тысяч [драхм].
ACTS|19|20|С такою силою возрастало и возмогало слово Господне.
ACTS|19|21|Когда же это совершилось, Павел положил в духе, пройдя Македонию и Ахаию, идти в Иерусалим, сказав: побывав там, я должен видеть и Рим.
ACTS|19|22|И, послав в Македонию двоих из служивших ему, Тимофея и Ераста, сам остался на время в Асии.
ACTS|19|23|В то время произошел немалый мятеж против пути Господня,
ACTS|19|24|ибо некто серебряник, именем Димитрий, делавший серебряные храмы Артемиды и доставлявший художникам немалую прибыль,
ACTS|19|25|собрав их и других подобных ремесленников, сказал: друзья! вы знаете, что от этого ремесла зависит благосостояние наше;
ACTS|19|26|между тем вы видите и слышите, что не только в Ефесе, но почти во всей Асии этот Павел своими убеждениями совратил немалое число людей, говоря, что делаемые руками человеческими не суть боги.
ACTS|19|27|А это нам угрожает тем, что не только ремесло наше придет в презрение, но и храм великой богини Артемиды ничего не будет значить, и испровергнется величие той, которую почитает вся Асия и вселенная.
ACTS|19|28|Выслушав это, они исполнились ярости и стали кричать, говоря: велика Артемида Ефесская!
ACTS|19|29|И весь город наполнился смятением. Схватив Македонян Гаия и Аристарха, спутников Павловых, они единодушно устремились на зрелище.
ACTS|19|30|Когда же Павел хотел войти в народ, ученики не допустили его.
ACTS|19|31|Также и некоторые из Асийских начальников, будучи друзьями его, послав к нему, просили не показываться на зрелище.
ACTS|19|32|Между тем одни кричали одно, а другие другое, ибо собрание было беспорядочное, и большая часть [собравшихся] не знали, зачем собрались.
ACTS|19|33|По предложению Иудеев, из народа вызван был Александр. Дав знак рукою, Александр хотел говорить к народу.
ACTS|19|34|Когда же узнали, что он Иудей, то закричали все в один голос, и около двух часов кричали: велика Артемида Ефесская!
ACTS|19|35|Блюститель же порядка, утишив народ, сказал: мужи Ефесские! какой человек не знает, что город Ефес есть служитель великой богини Артемиды и Диопета?
ACTS|19|36|Если же в этом нет спора, то надобно вам быть спокойными и не поступать опрометчиво.
ACTS|19|37|А вы привели этих мужей, которые ни храма Артемидина не обокрали, ни богини вашей не хулили.
ACTS|19|38|Если же Димитрий и другие с ним художники имеют жалобу на кого–нибудь, то есть судебные собрания и есть проконсулы: пусть жалуются друг на друга.
ACTS|19|39|А если вы ищете чего–нибудь другого, то это будет решено в законном собрании.
ACTS|19|40|Ибо мы находимся в опасности – за происшедшее ныне быть обвиненными в возмущении, так как нет никакой причины, которою мы могли бы оправдать такое сборище. Сказав это, он распустил собрание.
ACTS|20|1|По прекращении мятежа Павел, призвав учеников и дав им наставления и простившись с ними, вышел и пошел в Македонию.
ACTS|20|2|Пройдя же те места и преподав [верующим] обильные наставления, пришел в Елладу.
ACTS|20|3|[Там] пробыл он три месяца. Когда же, по случаю возмущения, сделанного против него Иудеями, он хотел отправиться в Сирию, то пришло ему на мысль возвратиться через Македонию.
ACTS|20|4|Его сопровождали до Асии Сосипатр Пирров, Вериянин, и из Фессалоникийцев Аристарх и Секунд, и Гаий Дервянин и Тимофей, и Асийцы Тихик и Трофим.
ACTS|20|5|Они, пойдя вперед, ожидали нас в Троаде.
ACTS|20|6|А мы, после дней опресночных, отплыли из Филипп и дней в пять прибыли к ним в Троаду, где пробыли семь дней.
ACTS|20|7|В первый же день недели, когда ученики собрались для преломления хлеба, Павел, намереваясь отправиться в следующий день, беседовал с ними и продолжил слово до полуночи.
ACTS|20|8|В горнице, где мы собрались, было довольно светильников.
ACTS|20|9|Во время продолжительной беседы Павловой один юноша, именем Евтих, сидевший на окне, погрузился в глубокий сон и, пошатнувшись, сонный упал вниз с третьего жилья, и поднят мертвым.
ACTS|20|10|Павел, сойдя, пал на него и, обняв его, сказал: не тревожьтесь, ибо душа его в нем.
ACTS|20|11|Взойдя же и преломив хлеб и вкусив, беседовал довольно, даже до рассвета, и потом вышел.
ACTS|20|12|Между тем отрока привели живого, и немало утешились.
ACTS|20|13|Мы пошли вперед на корабль и поплыли в Асс, чтобы взять оттуда Павла; ибо он так приказал нам, намереваясь сам идти пешком.
ACTS|20|14|Когда же он сошелся с нами в Ассе, то, взяв его, мы прибыли в Митилину.
ACTS|20|15|И, отплыв оттуда, в следующий день мы остановились против Хиоса, а на другой пристали к Самосу и, побывав в Трогиллии, в следующий [день] прибыли в Милит,
ACTS|20|16|ибо Павлу рассудилось миновать Ефес, чтобы не замедлить ему в Асии; потому что он поспешал, если можно, в день Пятидесятницы быть в Иерусалиме.
ACTS|20|17|Из Милита же послав в Ефес, он призвал пресвитеров церкви,
ACTS|20|18|и, когда они пришли к нему, он сказал им: вы знаете, как я с первого дня, в который пришел в Асию, все время был с вами,
ACTS|20|19|работая Господу со всяким смиренномудрием и многими слезами, среди искушений, приключавшихся мне по злоумышлениям Иудеев;
ACTS|20|20|как я не пропустил ничего полезного, о чем вам не проповедывал бы и чему не учил бы вас всенародно и по домам,
ACTS|20|21|возвещая Иудеям и Еллинам покаяние пред Богом и веру в Господа нашего Иисуса Христа.
ACTS|20|22|И вот, ныне я, по влечению Духа, иду в Иерусалим, не зная, что там встретится со мною;
ACTS|20|23|только Дух Святый по всем городам свидетельствует, говоря, что узы и скорби ждут меня.
ACTS|20|24|Но я ни на что не взираю и не дорожу своею жизнью, только бы с радостью совершить поприще мое и служение, которое я принял от Господа Иисуса, проповедать Евангелие благодати Божией.
ACTS|20|25|И ныне, вот, я знаю, что уже не увидите лица моего все вы, между которыми ходил я, проповедуя Царствие Божие.
ACTS|20|26|Посему свидетельствую вам в нынешний день, что чист я от крови всех,
ACTS|20|27|ибо я не упускал возвещать вам всю волю Божию.
ACTS|20|28|Итак внимайте себе и всему стаду, в котором Дух Святый поставил вас блюстителями, пасти Церковь Господа и Бога, которую Он приобрел Себе Кровию Своею.
ACTS|20|29|Ибо я знаю, что, по отшествии моем, войдут к вам лютые волки, не щадящие стада;
ACTS|20|30|и из вас самих восстанут люди, которые будут говорить превратно, дабы увлечь учеников за собою.
ACTS|20|31|Посему бодрствуйте, памятуя, что я три года день и ночь непрестанно со слезами учил каждого из вас.
ACTS|20|32|И ныне предаю вас, братия, Богу и слову благодати Его, могущему назидать [вас] более и дать вам наследие со всеми освященными.
ACTS|20|33|Ни серебра, ни золота, ни одежды я ни от кого не пожелал:
ACTS|20|34|сами знаете, что нуждам моим и [нуждам] бывших при мне послужили руки мои сии.
ACTS|20|35|Во всем показал я вам, что, так трудясь, надобно поддерживать слабых и памятовать слова Господа Иисуса, ибо Он Сам сказал: "блаженнее давать, нежели принимать".
ACTS|20|36|Сказав это, он преклонил колени свои и со всеми ими помолился.
ACTS|20|37|Тогда немалый плач был у всех, и, падая на выю Павла, целовали его,
ACTS|20|38|скорбя особенно от сказанного им слова, что они уже не увидят лица его. И провожали его до корабля.
ACTS|21|1|Когда же мы, расставшись с ними, отплыли, то прямо пришли в Кос, на другой день в Родос и оттуда в Патару,
ACTS|21|2|и, найдя корабль, идущий в Финикию, взошли на него и отплыли.
ACTS|21|3|Быв в виду Кипра и оставив его слева, мы плыли в Сирию, и пристали в Тире, ибо тут надлежало сложить груз с корабля.
ACTS|21|4|И, найдя учеников, пробыли там семь дней. Они, по [внушению] Духа, говорили Павлу, чтобы он не ходил в Иерусалим.
ACTS|21|5|Проведя эти дни, мы вышли и пошли, и нас провожали все с женами и детьми даже за город; а на берегу, преклонив колени, помолились.
ACTS|21|6|И, простившись друг с другом, мы вошли в корабль, а они возвратились домой.
ACTS|21|7|Мы же, совершив плавание, прибыли из Тира в Птолемаиду, где, приветствовав братьев, пробыли у них один день.
ACTS|21|8|А на другой день Павел и мы, бывшие с ним, выйдя, пришли в Кесарию и, войдя в дом Филиппа благовестника, одного из семи [диаконов], остались у него.
ACTS|21|9|У него были четыре дочери девицы, пророчествующие.
ACTS|21|10|Между тем как мы пребывали у них многие дни, пришел из Иудеи некто пророк, именем Агав,
ACTS|21|11|и, войдя к нам, взял пояс Павлов и, связав себе руки и ноги, сказал: так говорит Дух Святый: мужа, чей этот пояс, так свяжут в Иерусалиме Иудеи и предадут в руки язычников.
ACTS|21|12|Когда же мы услышали это, то и мы и тамошние просили, чтобы он не ходил в Иерусалим.
ACTS|21|13|Но Павел в ответ сказал: что вы делаете? что плачете и сокрушаете сердце мое? я не только хочу быть узником, но готов умереть в Иерусалиме за имя Господа Иисуса.
ACTS|21|14|Когда же мы не могли уговорить его, то успокоились, сказав: да будет воля Господня!
ACTS|21|15|После сих дней, приготовившись, пошли мы в Иерусалим.
ACTS|21|16|С нами шли и некоторые ученики из Кесарии, провожая [нас] к некоему давнему ученику, Мнасону Кипрянину, у которого можно было бы нам жить.
ACTS|21|17|По прибытии нашем в Иерусалим братия радушно приняли нас.
ACTS|21|18|На другой день Павел пришел с нами к Иакову; пришли и все пресвитеры.
ACTS|21|19|Приветствовав их, [Павел] рассказывал подробно, что сотворил Бог у язычников служением его.
ACTS|21|20|Они же, выслушав, прославили Бога и сказали ему: видишь, брат, сколько тысяч уверовавших Иудеев, и все они ревнители закона.
ACTS|21|21|А о тебе наслышались они, что ты всех Иудеев, живущих между язычниками, учишь отступлению от Моисея, говоря, чтобы они не обрезывали детей своих и не поступали по обычаям.
ACTS|21|22|Итак что же? Верно соберется народ; ибо услышат, что ты пришел.
ACTS|21|23|Сделай же, что мы скажем тебе: есть у нас четыре человека, имеющие на себе обет.
ACTS|21|24|Взяв их, очистись с ними, и возьми на себя издержки на [жертву] за них, чтобы остригли себе голову, и узнают все, что слышанное ими о тебе несправедливо, но что и сам ты продолжаешь соблюдать закон.
ACTS|21|25|А об уверовавших язычниках мы писали, положив, чтобы они ничего такого не наблюдали, а только хранили себя от идоложертвенного, от крови, от удавленины и от блуда.
ACTS|21|26|Тогда Павел, взяв тех мужей и очистившись с ними, в следующий день вошел в храм и объявил окончание дней очищения, когда должно быть принесено за каждого из них приношение.
ACTS|21|27|Когда же семь дней оканчивались, тогда Асийские Иудеи, увидев его в храме, возмутили весь народ и наложили на него руки,
ACTS|21|28|крича: мужи Израильские, помогите! этот человек всех повсюду учит против народа и закона и места сего; притом и Еллинов ввел в храм и осквернил святое место сие.
ACTS|21|29|Ибо перед тем они видели с ним в городе Трофима Ефесянина и думали, что Павел его ввел в храм.
ACTS|21|30|Весь город пришел в движение, и сделалось стечение народа; и, схватив Павла, повлекли его вон из храма, и тотчас заперты были двери.
ACTS|21|31|Когда же они хотели убить его, до тысяченачальника полка дошла весть, что весь Иерусалим возмутился.
ACTS|21|32|Он, тотчас взяв воинов и сотников, устремился на них; они же, увидев тысяченачальника и воинов, перестали бить Павла.
ACTS|21|33|Тогда тысяченачальник, приблизившись, взял его и велел сковать двумя цепями, и спрашивал: кто он, и что сделал.
ACTS|21|34|В народе одни кричали одно, а другие другое. Он же, не могши по причине смятения узнать ничего верного, повелел вести его в крепость.
ACTS|21|35|Когда же он был на лестнице, то воинам пришлось нести его по причине стеснения от народа,
ACTS|21|36|ибо множество народа следовало и кричало: смерть ему!
ACTS|21|37|При входе в крепость Павел сказал тысяченачальнику: можно ли мне сказать тебе нечто? А тот сказал: ты знаешь по–гречески?
ACTS|21|38|Так не ты ли тот Египтянин, который перед сими днями произвел возмущение и вывел в пустыню четыре тысячи человек разбойников?
ACTS|21|39|Павел же сказал: я Иудеянин, Тарсянин, гражданин небезызвестного Киликийского города; прошу тебя, позволь мне говорить к народу.
ACTS|21|40|Когда же тот позволил, Павел, стоя на лестнице, дал знак рукою народу; и, когда сделалось глубокое молчание, начал говорить на еврейском языке так:
ACTS|22|1|Мужи братия и отцы! выслушайте теперь мое оправдание перед вами.
ACTS|22|2|Услышав же, что он заговорил с ними на еврейском языке, они еще более утихли. Он сказал:
ACTS|22|3|я Иудеянин, родившийся в Тарсе Киликийском, воспитанный в сем городе при ногах Гамалиила, тщательно наставленный в отеческом законе, ревнитель по Боге, как и все вы ныне.
ACTS|22|4|Я даже до смерти гнал [последователей] сего учения, связывая и предавая в темницу и мужчин и женщин,
ACTS|22|5|как засвидетельствует о мне первосвященник и все старейшины, от которых и письма взяв к братиям, живущим в Дамаске, я шел, чтобы тамошних привести в оковах в Иерусалим на истязание.
ACTS|22|6|Когда же я был в пути и приближался к Дамаску, около полудня вдруг осиял меня великий свет с неба.
ACTS|22|7|Я упал на землю и услышал голос, говоривший мне: Савл, Савл! что ты гонишь Меня?
ACTS|22|8|Я отвечал: кто Ты, Господи? Он сказал мне: Я Иисус Назорей, Которого ты гонишь.
ACTS|22|9|Бывшие же со мною свет видели, и пришли в страх; но голоса Говорившего мне не слыхали.
ACTS|22|10|Тогда я сказал: Господи! что мне делать? Господь же сказал мне: встань и иди в Дамаск, и там тебе сказано будет все, что назначено тебе делать.
ACTS|22|11|А как я от славы света того лишился зрения, то бывшие со мною за руку привели меня в Дамаск.
ACTS|22|12|Некто Анания, муж благочестивый по закону, одобряемый всеми Иудеями, живущими в Дамаске,
ACTS|22|13|пришел ко мне и, подойдя, сказал мне: брат Савл! прозри. И я тотчас увидел его.
ACTS|22|14|Он же сказал мне: Бог отцов наших предъизбрал тебя, чтобы ты познал волю Его, увидел Праведника и услышал глас из уст Его,
ACTS|22|15|потому что ты будешь Ему свидетелем пред всеми людьми о том, что ты видел и слышал.
ACTS|22|16|Итак, что ты медлишь? Встань, крестись и омой грехи твои, призвав имя Господа Иисуса,
ACTS|22|17|Когда же я возвратился в Иерусалим и молился в храме, пришел я в исступление,
ACTS|22|18|и увидел Его, и Он сказал мне: поспеши и выйди скорее из Иерусалима, потому что [здесь] не примут твоего свидетельства о Мне.
ACTS|22|19|Я сказал: Господи! им известно, что я верующих в Тебя заключал в темницы и бил в синагогах,
ACTS|22|20|и когда проливалась кровь Стефана, свидетеля Твоего, я там стоял, одобрял убиение его и стерег одежды побивавших его.
ACTS|22|21|И Он сказал мне: иди; Я пошлю тебя далеко к язычникам.
ACTS|22|22|До этого слова слушали его; а за сим подняли крик, говоря: истреби от земли такого! ибо ему не должно жить.
ACTS|22|23|Между тем как они кричали, метали одежды и бросали пыль на воздух,
ACTS|22|24|тысяченачальник повелел ввести его в крепость, приказав бичевать его, чтобы узнать, по какой причине так кричали против него.
ACTS|22|25|Но когда растянули его ремнями, Павел сказал стоявшему сотнику: разве вам позволено бичевать Римского гражданина, да и без суда?
ACTS|22|26|Услышав это, сотник подошел и донес тысяченачальнику, говоря: смотри, что ты хочешь делать? этот человек – Римский гражданин.
ACTS|22|27|Тогда тысяченачальник, подойдя к нему, сказал: скажи мне, ты Римский гражданин? Он сказал: да.
ACTS|22|28|Тысяченачальник отвечал: я за большие деньги приобрел это гражданство. Павел же сказал: а я и родился в нем.
ACTS|22|29|Тогда тотчас отступили от него хотевшие пытать его. А тысяченачальник, узнав, что он Римский гражданин, испугался, что связал его.
ACTS|22|30|На другой день, желая достоверно узнать, в чем обвиняют его Иудеи, освободил его от оков и повелел собраться первосвященникам и всему синедриону и, выведя Павла, поставил его перед ними.
ACTS|23|1|Павел, устремив взор на синедрион, сказал: мужи братия! я всею доброю совестью жил пред Богом до сего дня.
ACTS|23|2|Первосвященник же Анания стоявшим перед ним приказал бить его по устам.
ACTS|23|3|Тогда Павел сказал ему: Бог будет бить тебя, стена подбеленная! ты сидишь, чтобы судить по закону, и, вопреки закону, велишь бить меня.
ACTS|23|4|Предстоящие же сказали: первосвященника Божия поносишь?
ACTS|23|5|Павел сказал: я не знал, братия, что он первосвященник; ибо написано: начальствующего в народе твоем не злословь.
ACTS|23|6|Узнав же Павел, что [тут] одна часть саддукеев, а другая фарисеев, возгласил в синедрионе: мужи братия! я фарисей, сын фарисея; за чаяние воскресения мертвых меня судят.
ACTS|23|7|Когда же он сказал это, произошла распря между фарисеями и саддукеями, и собрание разделилось.
ACTS|23|8|Ибо саддукеи говорят, что нет воскресения, ни Ангела, ни духа; а фарисеи признают и то и другое.
ACTS|23|9|Сделался большой крик; и, встав, книжники фарисейской стороны спорили, говоря: ничего худого мы не находим в этом человеке; если же дух или Ангел говорил ему, не будем противиться Богу.
ACTS|23|10|Но как раздор увеличился, то тысяченачальник, опасаясь, чтобы они не растерзали Павла, повелел воинам сойти взять его из среды их и отвести в крепость.
ACTS|23|11|В следующую ночь Господь, явившись ему, сказал: дерзай, Павел; ибо, как ты свидетельствовал о Мне в Иерусалиме, так надлежит тебе свидетельствовать и в Риме.
ACTS|23|12|С наступлением дня некоторые Иудеи сделали умысел, и заклялись не есть и не пить, доколе не убьют Павла.
ACTS|23|13|Было же более сорока сделавших такое заклятие.
ACTS|23|14|Они, придя к первосвященникам и старейшинам, сказали: мы клятвою заклялись не есть ничего, пока не убьем Павла.
ACTS|23|15|Итак ныне же вы с синедрионом дайте знать тысяченачальнику, чтобы он завтра вывел его к вам, как будто вы хотите точнее рассмотреть дело о нем; мы же, прежде нежели он приблизится, готовы убить его.
ACTS|23|16|Услышав о сем умысле, сын сестры Павловой пришел и, войдя в крепость, уведомил Павла.
ACTS|23|17|Павел же, призвав одного из сотников, сказал: отведи этого юношу к тысяченачальнику, ибо он имеет нечто сказать ему.
ACTS|23|18|Тот, взяв его, привел к тысяченачальнику и сказал: узник Павел, призвав меня, просил отвести к тебе этого юношу, который имеет нечто сказать тебе.
ACTS|23|19|Тысяченачальник, взяв его за руку и отойдя с ним в сторону, спрашивал: что такое имеешь ты сказать мне?
ACTS|23|20|Он отвечал, что Иудеи согласились просить тебя, чтобы ты завтра вывел Павла пред синедрион, как будто они хотят точнее исследовать дело о нем.
ACTS|23|21|Но ты не слушай их; ибо его подстерегают более сорока человек из них, которые заклялись не есть и не пить, доколе не убьют его; и они теперь готовы, ожидая твоего распоряжения.
ACTS|23|22|Тогда тысяченачальник отпустил юношу, сказав: никому не говори, что ты объявил мне это.
ACTS|23|23|И, призвав двух сотников, сказал: приготовьте мне воинов [пеших] двести, конных семьдесят и стрелков двести, чтобы с третьего часа ночи шли в Кесарию.
ACTS|23|24|Приготовьте также ослов, чтобы, посадив Павла, препроводить его к правителю Феликсу.
ACTS|23|25|Написал и письмо следующего содержания:
ACTS|23|26|"Клавдий Лисий достопочтенному правителю Феликсу – радоваться.
ACTS|23|27|Сего человека Иудеи схватили и готовы были убить; я, придя с воинами, отнял его, узнав, что он Римский гражданин.
ACTS|23|28|Потом, желая узнать, в чем обвиняли его, привел его в синедрион их
ACTS|23|29|и нашел, что его обвиняют в спорных мнениях, касающихся закона их, но что нет в нем никакой вины, достойной смерти или оков.
ACTS|23|30|А как до меня дошло, что Иудеи злоумышляют на этого человека, то я немедленно послал его к тебе, приказав и обвинителям говорить на него перед тобою. Будь здоров".
ACTS|23|31|Итак воины, по [данному] им приказанию, взяв Павла, повели ночью в Антипатриду.
ACTS|23|32|А на другой день, предоставив конным идти с ним, возвратились в крепость.
ACTS|23|33|А те, придя в Кесарию и отдав письмо правителю, представили ему и Павла.
ACTS|23|34|Правитель, прочитав письмо, спросил, из какой он области, и, узнав, что из Киликии, сказал:
ACTS|23|35|я выслушаю тебя, когда явятся твои обвинители. И повелел ему быть под стражею в Иродовой претории.
ACTS|24|1|Через пять дней пришел первосвященник Анания со старейшинами и с некоторым ритором Тертуллом, которые жаловались правителю на Павла.
ACTS|24|2|Когда же он был призван, то Тертулл начал обвинять его, говоря:
ACTS|24|3|всегда и везде со всякою благодарностью признаем мы, что тебе, достопочтенный Феликс, обязаны мы многим миром, и твоему попечению благоустроением сего народа.
ACTS|24|4|Но, чтобы много не утруждать тебя, прошу тебя выслушать нас кратко, со свойственным тебе снисхождением.
ACTS|24|5|Найдя сего человека язвою [общества], возбудителем мятежа между иудеями, живущими по вселенной, и представителем Назорейской ереси,
ACTS|24|6|который отважился даже осквернить храм, мы взяли его и хотели судить его по нашему закону.
ACTS|24|7|Но тысяченачальник Лисий, придя, с великим насилием взял его из рук наших и послал к тебе,
ACTS|24|8|повелев и нам, обвинителям его, идти к тебе. Ты можешь сам, разобрав, узнать от него о всем том, в чем мы обвиняем его.
ACTS|24|9|И Иудеи подтвердили, сказав, что это так.
ACTS|24|10|Павел же, когда правитель дал ему знак говорить, отвечал: зная, что ты многие годы справедливо судишь народ сей, я тем свободнее буду защищать мое дело.
ACTS|24|11|Ты можешь узнать, что не более двенадцати дней тому, как я пришел в Иерусалим для поклонения.
ACTS|24|12|И ни в святилище, ни в синагогах, ни по городу они не находили меня с кем–либо спорящим или производящим народное возмущение,
ACTS|24|13|и не могут доказать того, в чем теперь обвиняют меня.
ACTS|24|14|Но в том признаюсь тебе, что по учению, которое они называют ересью, я действительно служу Богу отцов [моих], веруя всему, написанному в законе и пророках,
ACTS|24|15|имея надежду на Бога, что будет воскресение мертвых, праведных и неправедных, чего и сами они ожидают.
ACTS|24|16|Посему и сам подвизаюсь всегда иметь непорочную совесть пред Богом и людьми.
ACTS|24|17|После многих лет я пришел, чтобы доставить милостыню народу моему и приношения.
ACTS|24|18|При сем нашли меня, очистившегося в храме не с народом и не с шумом.
ACTS|24|19|[Это были] некоторые Асийские Иудеи, которым надлежало бы предстать пред тебя и обвинять меня, если что имеют против меня.
ACTS|24|20|Или пусть сии самые скажут, какую нашли они во мне неправду, когда я стоял перед синедрионом,
ACTS|24|21|разве только то одно слово, которое громко произнес я, стоя между ними, что за [учение о] воскресении мертвых я ныне судим вами.
ACTS|24|22|Выслушав это, Феликс отсрочил [дело] их, сказав: рассмотрю ваше дело, когда придет тысяченачальник Лисий, и я обстоятельно узнаю об этом учении.
ACTS|24|23|А Павла приказал сотнику стеречь, но не стеснять его и не запрещать никому из его близких служить ему или приходить к нему.
ACTS|24|24|Через несколько дней Феликс, придя с Друзиллою, женою своею, Иудеянкою, призвал Павла, и слушал его о вере во Христа Иисуса.
ACTS|24|25|И как он говорил о правде, о воздержании и о будущем суде, то Феликс пришел в страх и отвечал: теперь пойди, а когда найду время, позову тебя.
ACTS|24|26|Притом же надеялся он, что Павел даст ему денег, чтобы отпустил его: посему часто призывал его и беседовал с ним.
ACTS|24|27|Но по прошествии двух лет на место Феликса поступил Порций Фест. Желая доставить удовольствие Иудеям, Феликс оставил Павла в узах.
ACTS|25|1|Фест, прибыв в область, через три дня отправился из Кесарии в Иерусалим.
ACTS|25|2|Тогда первосвященник и знатнейшие из Иудеев явились к нему [с] [жалобою] на Павла и убеждали его,
ACTS|25|3|прося, чтобы он сделал милость, вызвал его в Иерусалим; и злоумышляли убить его на дороге.
ACTS|25|4|Но Фест отвечал, что Павел содержится в Кесарии под стражею и что он сам скоро отправится туда.
ACTS|25|5|Итак, сказал он, которые из вас могут, пусть пойдут со мною, и если есть что–нибудь за этим человеком, пусть обвиняют его.
ACTS|25|6|Пробыв же у них не больше восьми или десяти дней, возвратился в Кесарию, и на другой день, сев на судейское место, повелел привести Павла.
ACTS|25|7|Когда он явился, стали кругом пришедшие из Иерусалима Иудеи, принося на Павла многие и тяжкие обвинения, которых не могли доказать.
ACTS|25|8|Он же в оправдание свое сказал: я не сделал никакого преступления ни против закона Иудейского, ни против храма, ни против кесаря.
ACTS|25|9|Фест, желая сделать угождение Иудеям, сказал в ответ Павлу: хочешь ли идти в Иерусалим, чтобы я там судил тебя в этом?
ACTS|25|10|Павел сказал: я стою перед судом кесаревым, где мне и следует быть судиму. Иудеев я ничем не обидел, как и ты хорошо знаешь.
ACTS|25|11|Ибо, если я неправ и сделал что–нибудь, достойное смерти, то не отрекаюсь умереть; а если ничего того нет, в чем сии обвиняют меня, то никто не может выдать меня им. Требую суда кесарева.
ACTS|25|12|Тогда Фест, поговорив с советом, отвечал: ты потребовал суда кесарева, к кесарю и отправишься.
ACTS|25|13|Через несколько дней царь Агриппа и Вереника прибыли в Кесарию поздравить Феста.
ACTS|25|14|И как они провели там много дней, то Фест предложил царю дело Павлово, говоря: [здесь] есть человек, оставленный Феликсом в узах,
ACTS|25|15|на которого, в бытность мою в Иерусалиме, [с жалобою] явились первосвященники и старейшины Иудейские, требуя осуждения его.
ACTS|25|16|Я отвечал им, что у Римлян нет обыкновения выдавать какого–нибудь человека на смерть, прежде нежели обвиняемый будет иметь обвинителей налицо и получит свободу защищаться против обвинения.
ACTS|25|17|Когда же они пришли сюда, то, без всякого отлагательства, на другой же день сел я на судейское место и повелел привести того человека.
ACTS|25|18|Обступив его, обвинители не представили ни одного из обвинений, какие я предполагал;
ACTS|25|19|но они имели некоторые споры с ним об их Богопочитании и о каком–то Иисусе умершем, о Котором Павел утверждал, что Он жив.
ACTS|25|20|Затрудняясь в решении этого вопроса, я сказал: хочет ли он идти в Иерусалим и там быть судимым в этом?
ACTS|25|21|Но как Павел потребовал, чтобы он оставлен был на рассмотрение Августово, то я велел содержать его под стражею до тех пор, как пошлю его к кесарю.
ACTS|25|22|Агриппа же сказал Фесту: хотел бы и я послушать этого человека. Завтра же, отвечал тот, услышишь его.
ACTS|25|23|На другой день, когда Агриппа и Вереника пришли с великою пышностью и вошли в судебную палату с тысяченачальниками и знатнейшими гражданами, по приказанию Феста приведен был Павел.
ACTS|25|24|И сказал Фест: царь Агриппа и все присутствующие с нами мужи! вы видите того, против которого все множество Иудеев приступали ко мне в Иерусалиме и здесь и кричали, что ему не должно более жить.
ACTS|25|25|Но я нашел, что он не сделал ничего, достойного смерти; и как он сам потребовал суда у Августа, то я решился послать его [к нему].
ACTS|25|26|Я не имею ничего верного написать о нем государю; посему привел его пред вас, и особенно пред тебя, царь Агриппа, дабы, по рассмотрении, было мне что написать.
ACTS|25|27|Ибо, мне кажется, нерассудительно послать узника и не показать обвинений на него.
ACTS|26|1|Агриппа сказал Павлу: позволяется тебе говорить за себя. Тогда Павел, простерши руку, стал говорить в свою защиту:
ACTS|26|2|царь Агриппа! почитаю себя счастливым, что сегодня могу защищаться перед тобою во всем, в чем обвиняют меня Иудеи,
ACTS|26|3|тем более, что ты знаешь все обычаи и спорные мнения Иудеев. Посему прошу тебя выслушать меня великодушно.
ACTS|26|4|Жизнь мою от юности [моей], которую сначала проводил я среди народа моего в Иерусалиме, знают все Иудеи;
ACTS|26|5|они издавна знают обо мне, если захотят свидетельствовать, что я жил фарисеем по строжайшему в нашем вероисповедании учению.
ACTS|26|6|И ныне я стою перед судом за надежду на обетование, данное от Бога нашим отцам,
ACTS|26|7|которого исполнение надеются увидеть наши двенадцать колен, усердно служа [Богу] день и ночь. За сию–то надежду, царь Агриппа, обвиняют меня Иудеи.
ACTS|26|8|Что же? Неужели вы невероятным почитаете, что Бог воскрешает мертвых?
ACTS|26|9|Правда, и я думал, что мне должно много действовать против имени Иисуса Назорея.
ACTS|26|10|Это я и делал в Иерусалиме: получив власть от первосвященников, я многих святых заключал в темницы, и, когда убивали их, я подавал на то голос;
ACTS|26|11|и по всем синагогам я многократно мучил их и принуждал хулить [Иисуса] и, в чрезмерной против них ярости, преследовал даже и в чужих городах.
ACTS|26|12|Для сего, идя в Дамаск со властью и поручением от первосвященников,
ACTS|26|13|среди дня на дороге я увидел, государь, с неба свет, превосходящий солнечное сияние, осиявший меня и шедших со мною.
ACTS|26|14|Все мы упали на землю, и я услышал голос, говоривший мне на еврейском языке: Савл, Савл! что ты гонишь Меня? Трудно тебе идти против рожна.
ACTS|26|15|Я сказал: кто Ты, Господи? Он сказал: "Я Иисус, Которого ты гонишь.
ACTS|26|16|Но встань и стань на ноги твои; ибо Я для того и явился тебе, чтобы поставить тебя служителем и свидетелем того, что ты видел и что Я открою тебе,
ACTS|26|17|избавляя тебя от народа Иудейского и от язычников, к которым Я теперь посылаю тебя
ACTS|26|18|открыть глаза им, чтобы они обратились от тьмы к свету и от власти сатаны к Богу, и верою в Меня получили прощение грехов и жребий с освященными".
ACTS|26|19|Поэтому, царь Агриппа, я не воспротивился небесному видению,
ACTS|26|20|но сперва жителям Дамаска и Иерусалима, потом всей земле Иудейской и язычникам проповедывал, чтобы они покаялись и обратились к Богу, делая дела, достойные покаяния.
ACTS|26|21|За это схватили меня Иудеи в храме и покушались растерзать.
ACTS|26|22|Но, получив помощь от Бога, я до сего дня стою, свидетельствуя малому и великому, ничего не говоря, кроме того, о чем пророки и Моисей говорили, что это будет,
ACTS|26|23|[то есть] что Христос имел пострадать и, восстав первый из мертвых, возвестить свет народу (Иудейскому) и язычникам.
ACTS|26|24|Когда он так защищался, Фест громким голосом сказал: безумствуешь ты, Павел! большая ученость доводит тебя до сумасшествия.
ACTS|26|25|Нет, достопочтенный Фест, сказал он, я не безумствую, но говорю слова истины и здравого смысла.
ACTS|26|26|Ибо знает об этом царь, перед которым и говорю смело. Я отнюдь не верю, чтобы от него было что–нибудь из сего скрыто; ибо это не в углу происходило.
ACTS|26|27|Веришь ли, царь Агриппа, пророкам? Знаю, что веришь.
ACTS|26|28|Агриппа сказал Павлу: ты немного не убеждаешь меня сделаться Христианином.
ACTS|26|29|Павел сказал: молил бы я Бога, чтобы мало ли, много ли, не только ты, но и все, слушающие меня сегодня, сделались такими, как я, кроме этих уз.
ACTS|26|30|Когда он сказал это, царь и правитель, Вереника и сидевшие с ними встали;
ACTS|26|31|и, отойдя в сторону, говорили между собою, что этот человек ничего, достойного смерти или уз, не делает.
ACTS|26|32|И сказал Агриппа Фесту: можно было бы освободить этого человека, если бы он не потребовал суда у кесаря. Посему и решился правитель послать его к кесарю.
ACTS|27|1|Когда решено было плыть нам в Италию, то отдали Павла и некоторых других узников сотнику Августова полка, именем Юлию.
ACTS|27|2|Мы взошли на Адрамитский корабль и отправились, намереваясь плыть около Асийских мест. С нами был Аристарх, Македонянин из Фессалоники.
ACTS|27|3|На другой [день] пристали к Сидону. Юлий, поступая с Павлом человеколюбиво, позволил ему сходить к друзьям и воспользоваться их усердием.
ACTS|27|4|Отправившись оттуда, мы приплыли в Кипр, по причине противных ветров,
ACTS|27|5|и, переплыв море против Киликии и Памфилии, прибыли в Миры Ликийские.
ACTS|27|6|Там сотник нашел Александрийский корабль, плывущий в Италию, и посадил нас на него.
ACTS|27|7|Медленно плавая многие дни и едва поровнявшись с Книдом, по причине неблагоприятного нам ветра, мы подплыли к Криту при Салмоне.
ACTS|27|8|Пробравшись же с трудом мимо него, прибыли к одному месту, называемому Хорошие Пристани, близ которого был город Ласея.
ACTS|27|9|Но как прошло довольно времени, и плавание было уже опасно, потому что и пост уже прошел, то Павел советовал,
ACTS|27|10|говоря им: мужи! я вижу, что плавание будет с затруднениями и с большим вредом не только для груза и корабля, но и для нашей жизни.
ACTS|27|11|Но сотник более доверял кормчему и начальнику корабля, нежели словам Павла.
ACTS|27|12|А как пристань не была приспособлена к зимовке, то многие давали совет отправиться оттуда, чтобы, если можно, дойти до Финика, пристани Критской, лежащей против юго–западного и северо–западного ветра, и [там] перезимовать.
ACTS|27|13|Подул южный ветер, и они, подумав, что уже получили желаемое, отправились, и поплыли поблизости Крита.
ACTS|27|14|Но скоро поднялся против него ветер бурный, называемый эвроклидон.
ACTS|27|15|Корабль схватило так, что он не мог противиться ветру, и мы носились, отдавшись волнам.
ACTS|27|16|И, набежав на один островок, называемый Клавдой, мы едва могли удержать лодку.
ACTS|27|17|Подняв ее, стали употреблять пособия и обвязывать корабль; боясь же, чтобы не сесть на мель, спустили парус и таким образом носились.
ACTS|27|18|На другой день, по причине сильного обуревания, начали выбрасывать [груз],
ACTS|27|19|а на третий мы своими руками побросали с корабля вещи.
ACTS|27|20|Но как многие дни не видно было ни солнца, ни звезд и продолжалась немалая буря, то наконец исчезала всякая надежда к нашему спасению.
ACTS|27|21|И как долго не ели, то Павел, став посреди них, сказал: мужи! надлежало послушаться меня и не отходить от Крита, чем и избежали бы сих затруднений и вреда.
ACTS|27|22|Теперь же убеждаю вас ободриться, потому что ни одна душа из вас не погибнет, а только корабль.
ACTS|27|23|Ибо Ангел Бога, Которому принадлежу я и Которому служу, явился мне в эту ночь
ACTS|27|24|и сказал: "не бойся, Павел! тебе должно предстать пред кесаря, и вот, Бог даровал тебе всех плывущих с тобою".
ACTS|27|25|Посему ободритесь, мужи, ибо я верю Богу, что будет так, как мне сказано.
ACTS|27|26|Нам должно быть выброшенными на какой–нибудь остров.
ACTS|27|27|В четырнадцатую ночь, как мы носимы были в Адриатическом море, около полуночи корабельщики стали догадываться, что приближаются к какой–то земле,
ACTS|27|28|и, вымерив глубину, нашли двадцать сажен; потом на небольшом расстоянии, вымерив опять, нашли пятнадцать сажен.
ACTS|27|29|Опасаясь, чтобы не попасть на каменистые места, бросили с кормы четыре якоря, и ожидали дня.
ACTS|27|30|Когда же корабельщики хотели бежать с корабля и спускали на море лодку, делая вид, будто хотят бросить якоря с носа,
ACTS|27|31|Павел сказал сотнику и воинам: если они не останутся на корабле, то вы не можете спастись.
ACTS|27|32|Тогда воины отсекли веревки у лодки, и она упала.
ACTS|27|33|Перед наступлением дня Павел уговаривал всех принять пищу, говоря: сегодня четырнадцатый день, как вы, в ожидании, остаетесь без пищи, не вкушая ничего.
ACTS|27|34|Потому прошу вас принять пищу: это послужит к сохранению вашей жизни; ибо ни у кого из вас не пропадет волос с головы.
ACTS|27|35|Сказав это и взяв хлеб, он возблагодарил Бога перед всеми и, разломив, начал есть.
ACTS|27|36|Тогда все ободрились и также приняли пищу.
ACTS|27|37|Было же всех нас на корабле двести семьдесят шесть душ.
ACTS|27|38|Насытившись же пищею, стали облегчать корабль, выкидывая пшеницу в море.
ACTS|27|39|Когда настал день, земли не узнавали, а усмотрели только некоторый залив, имеющий [отлогий] берег, к которому и решились, если можно, пристать с кораблем.
ACTS|27|40|И, подняв якоря, пошли по морю и, развязав рули и подняв малый парус по ветру, держали к берегу.
ACTS|27|41|Попали на косу, и корабль сел на мель. Нос увяз и остался недвижим, а корма разбивалась силою волн.
ACTS|27|42|Воины согласились было умертвить узников, чтобы кто–нибудь, выплыв, не убежал.
ACTS|27|43|Но сотник, желая спасти Павла, удержал их от сего намерения, и велел умеющим плавать первым броситься и выйти на землю,
ACTS|27|44|прочим же [спасаться] кому на досках, а кому на чем–нибудь от корабля; и таким образом все спаслись на землю.
ACTS|28|1|Спасшись же, бывшие с Павлом узнали, что остров называется Мелит.
ACTS|28|2|Иноплеменники оказали нам немалое человеколюбие, ибо они, по причине бывшего дождя и холода, разложили огонь и приняли всех нас.
ACTS|28|3|Когда же Павел набрал множество хвороста и клал на огонь, тогда ехидна, выйдя от жара, повисла на руке его.
ACTS|28|4|Иноплеменники, когда увидели висящую на руке его змею, говорили друг другу: верно этот человек – убийца, когда его, спасшегося от моря, суд [Божий] не оставляет жить.
ACTS|28|5|Но он, стряхнув змею в огонь, не потерпел никакого вреда.
ACTS|28|6|Они ожидали было, что у него будет воспаление, или он внезапно упадет мертвым; но, ожидая долго и видя, что не случилось с ним никакой беды, переменили мысли и говорили, что он Бог.
ACTS|28|7|Около того места были поместья начальника острова, именем Публия; он принял нас и три дня дружелюбно угощал.
ACTS|28|8|Отец Публия лежал, страдая горячкою и болью в животе; Павел вошел к нему, помолился и, возложив на него руки свои, исцелил его.
ACTS|28|9|После сего события и прочие на острове, имевшие болезни, приходили и были исцеляемы,
ACTS|28|10|и оказывали нам много почести и при отъезде снабдили нужным.
ACTS|28|11|Через три месяца мы отплыли на Александрийском корабле, называемом Диоскуры, зимовавшем на том острове,
ACTS|28|12|и, приплыв в Сиракузы, пробыли там три дня.
ACTS|28|13|Оттуда отплыв, прибыли в Ригию; и как через день подул южный ветер, прибыли на второй день в Путеол,
ACTS|28|14|где нашли братьев, и были упрошены пробыть у них семь дней, а потом пошли в Рим.
ACTS|28|15|Тамошние братья, услышав о нас, вышли нам навстречу до Аппиевой площади и трех гостиниц. Увидев их, Павел возблагодарил Бога и ободрился.
ACTS|28|16|Когда же пришли мы в Рим, то сотник передал узников военачальнику, а Павлу позволено жить особо с воином, стерегущим его.
ACTS|28|17|Через три дня Павел созвал знатнейших из Иудеев и, когда они сошлись, говорил им: мужи братия! не сделав ничего против народа или отеческих обычаев, я в узах из Иерусалима предан в руки Римлян.
ACTS|28|18|Они, судив меня, хотели освободить, потому что нет во мне никакой вины, достойной смерти;
ACTS|28|19|но так как Иудеи противоречили, то я принужден был потребовать суда у кесаря, впрочем не с тем, чтобы обвинить в чем–либо мой народ.
ACTS|28|20|По этой причине я и призвал вас, чтобы увидеться и поговорить с вами, ибо за надежду Израилеву обложен я этими узами.
ACTS|28|21|Они же сказали ему: мы ни писем не получали о тебе из Иудеи, ни из приходящих братьев никто не известил о тебе и не сказал чего–либо худого.
ACTS|28|22|Впрочем желательно нам слышать от тебя, как ты мыслишь; ибо известно нам, что об этом учении везде спорят.
ACTS|28|23|И, назначив ему день, очень многие пришли к нему в гостиницу; и он от утра до вечера излагал им [учение] о Царствии Божием, приводя свидетельства и удостоверяя их о Иисусе из закона Моисеева и пророков.
ACTS|28|24|Одни убеждались словами его, а другие не верили.
ACTS|28|25|Будучи же не согласны между собою, они уходили, когда Павел сказал следующие слова: хорошо Дух Святый сказал отцам нашим через пророка Исаию:
ACTS|28|26|пойди к народу сему и скажи: слухом услышите, и не уразумеете, и очами смотреть будете, и не увидите.
ACTS|28|27|Ибо огрубело сердце людей сих, и ушами с трудом слышат, и очи свои сомкнули, да не узрят очами, и не услышат ушами, и не уразумеют сердцем, и не обратятся, чтобы Я исцелил их.
ACTS|28|28|Итак да будет вам известно, что спасение Божие послано язычникам: они и услышат.
ACTS|28|29|Когда он сказал это, Иудеи ушли, много споря между собою.
ACTS|28|30|И жил Павел целых два года на своем иждивении и принимал всех, приходивших к нему,
ACTS|28|31|проповедуя Царствие Божие и уча о Господе Иисусе Христе со всяким дерзновением невозбранно.
