2TIM|1|1|奉上帝旨意，按照基督耶穌裏所應許的生命，作基督耶穌使徒的 保羅 ，
2TIM|1|2|寫信給我親愛的兒子 提摩太 。願恩惠、憐憫、平安 從父上帝和我們的主基督耶穌歸給你！
2TIM|1|3|我感謝上帝，就是我接續祖先用純潔的良心所事奉的上帝，在祈禱中晝夜不停地想念你。
2TIM|1|4|我一想起你的眼淚，就急切想見你，好讓我滿心快樂。
2TIM|1|5|我記得你無偽的信心，這信心先存在你外祖母 羅以 和你母親 友妮基 的心裏，我深信也存在你的心裏。
2TIM|1|6|為這緣故，我提醒你要把上帝藉著我按手所給你的恩賜再如火挑旺起來。
2TIM|1|7|因為上帝賜給我們的不是膽怯的心，而是剛強、仁愛、自制的心。
2TIM|1|8|所以，不要以給我們的主作見證為恥，也不要以我這為主被囚的為恥；總要靠著上帝的大能，與我為福音同受苦難。
2TIM|1|9|上帝救了我們， 以聖召召我們， 不是按我們的行為， 而是按他的旨意和恩典； 這恩典是萬古之先 在基督耶穌裏賜給我們的，
2TIM|1|10|但如今 藉著我們的救主基督耶穌的顯現已經表明出來； 他把死廢去， 藉著福音，將不朽的生命彰顯出來。
2TIM|1|11|我為這福音奉派作傳道，作使徒，作教師。
2TIM|1|12|為這緣故，我也受這些苦難。然而，我不以為恥，因為我知道我所信的是誰，也深信他能保全他所交託我的 ，直到那日。
2TIM|1|13|你從我聽到那健全的言論，要用在基督耶穌裏的信心和愛心常常守著，作為規範。
2TIM|1|14|你要靠著那住在我們裏面的聖靈，牢牢守住所交託給你那美好的事。
2TIM|1|15|你知道，所有在 亞細亞 的人都離棄了我，其中有 腓吉路 和 黑摩其尼 。
2TIM|1|16|願主憐憫 阿尼色弗 一家的人，因為他屢次令我欣慰。他不以我的鐵鏈為恥，
2TIM|1|17|反而一到 羅馬 就急切尋找我，並且找到了。
2TIM|1|18|願主使他在那日能蒙主的憐憫。他在 以弗所 怎樣多服事我，你是清楚知道的。
2TIM|2|1|我兒啊，你要在基督耶穌的恩典上剛強起來。
2TIM|2|2|你在許多見證人面前聽見我所教導的，也要交託給那忠心而又能教導別人的人。
2TIM|2|3|你要和我同受苦難，作基督耶穌的精兵。
2TIM|2|4|凡當兵的，不讓世務纏身，好使那招他當兵的人喜悅。
2TIM|2|5|運動員在比賽的時候，不按規則就不能得冠冕。
2TIM|2|6|勤勞的農夫理當先得糧食。
2TIM|2|7|我所說的話，你要考慮，因為主必在凡事上給你聰明。
2TIM|2|8|要記得耶穌基督，他是 大衛 的後裔，從死人中復活；這就是我所傳的福音。
2TIM|2|9|我為這福音受苦難，甚至像犯人一樣被捆綁，然而上帝的話沒有被捆綁。
2TIM|2|10|所以，我為了選民事事忍耐，為使他們也能得到那在基督耶穌裏的救恩和永遠的榮耀。
2TIM|2|11|這話是可信的： 我們若與基督同死，也必與他同活；
2TIM|2|12|我們若忍耐到底，也必和他一同作王。 我們若不認他，他也必不認我們；
2TIM|2|13|我們縱然失信，他仍是可信的， 因為他不能否認自己。
2TIM|2|14|你要向眾人提醒這些事，在上帝 面前囑咐他們不可在言詞上爭辯；這是沒有益處的，只能傷害聽的人。
2TIM|2|15|你當竭力在上帝面前作一個經得起考驗、無愧的工人，按著正意講解真理的話。
2TIM|2|16|要遠避世俗的空談，因為這等空談會使人進到更不敬虔的地步。
2TIM|2|17|他們的話如同毒瘡越爛越大；其中有 許米乃 和 腓理徒 ，
2TIM|2|18|他們偏離了真理，說復活的事已過去，敗壞了好些人的信心。
2TIM|2|19|然而，上帝堅固的根基屹立不移；上面有這印記說：「主認得他自己的人」，又說：「凡稱呼主名的人總要離開不義。」
2TIM|2|20|大戶人家不但有金器銀器，也有木器瓦器；有作為貴重之用的，有作為卑賤之用的。
2TIM|2|21|人若自潔，脫離卑賤的事，必成為貴重的器皿，成為聖潔，合乎主用，預備行各樣的善事。
2TIM|2|22|你要逃避年輕人的私慾，同那以純潔的心求告主的人追求公義、信實、仁愛、和平。
2TIM|2|23|但要棄絕那愚拙無知的辯論，因為你知道這等事只會引起爭辯。
2TIM|2|24|主的僕人不可爭辯，只要溫和待人，善於教導，恆心忍耐，
2TIM|2|25|用溫柔勸導反對的人。也許上帝會給他們悔改的心能明白真理，
2TIM|2|26|讓他們這些已被魔鬼擄去順從他詭計的人能醒悟過來，脫離他的羅網。
2TIM|3|1|你該知道，末世必有艱難的日子來到。
2TIM|3|2|那時人會專愛自己，貪愛錢財，自誇，狂傲，毀謗，違背父母，忘恩負義，心不聖潔，
2TIM|3|3|沒有親情，抗拒和解，好說讒言，不能節制，性情兇暴，不愛良善，
2TIM|3|4|賣主賣友，任意妄為，自高自大，愛好宴樂，不愛上帝，
2TIM|3|5|有敬虔的外貌，卻背棄了敬虔的實質，這等人你要避開。
2TIM|3|6|他們當中有人潛入別人家裏，操縱無知的婦女；這些婦女被罪惡壓制，被各樣的私慾引誘，
2TIM|3|7|雖然常常學習，終久無法達到明白真理的地步。
2TIM|3|8|從前 雅尼 和 佯庇 怎樣反對 摩西 ，這等人也怎樣抵擋真理；他們的心地敗壞，信仰經不起考驗。
2TIM|3|9|然而，他們沒有進步，因為他們的愚昧必在眾人面前顯露出來，像那兩人一樣。
2TIM|3|10|但你已經追隨了我的教導、行為、志向、信心、寬容、愛心、忍耐，
2TIM|3|11|以及我在 安提阿 、 以哥念 、 路司得 所遭遇的迫害和苦難。我忍受了何等的迫害！但從這一切苦難中，主都把我救了出來。
2TIM|3|12|其實，凡立志在基督耶穌裏敬虔度日的，也都將受迫害。
2TIM|3|13|只是作惡的和騙人的將變本加厲，迷惑人也被人迷惑。
2TIM|3|14|至於你，你要持守所學習的和所確信的，因為你知道是跟誰學的，
2TIM|3|15|並且知道你從小明白聖經，這聖經能使你因在基督耶穌裏的信 有得救的智慧。
2TIM|3|16|聖經都是上帝所默示的 ，於教訓、督責、使人歸正、教導人學義都是有益的，
2TIM|3|17|叫屬上帝的人得以完全，預備行各樣的善事。
2TIM|4|1|我在上帝面前，並在將來審判活人死人的基督耶穌面前，憑著他的顯現和他的國度鄭重地勸戒你：
2TIM|4|2|務要傳道；無論得時不得時總要專心，並以百般的忍耐和各樣的教導責備人，警戒人，勸勉人。
2TIM|4|3|因為時候將到，那時人會厭煩健全的教導，耳朵發癢，就隨心所欲地增添好些教師，
2TIM|4|4|並且掩耳不聽真理，偏向無稽的傳說。
2TIM|4|5|至於你，凡事要謹慎，忍受苦難，做傳福音的工作，盡你的職分。
2TIM|4|6|至於我，我已經被澆獻，離世的時候到了。
2TIM|4|7|那美好的仗我已經打過了，當跑的路我已經跑盡了，該信的道我已經守住了。
2TIM|4|8|從此以後，有公義的冠冕為我存留，就是按著公義審判的主到了那日要賜給我的；不但賜給我，也賜給凡愛慕他顯現的人。
2TIM|4|9|你要趕緊到我這裏來。
2TIM|4|10|因為 底馬 貪愛現今的世界，已經離棄我，往 帖撒羅尼迦 去了； 革勒士 往 加拉太 去； 提多 往 撻馬太 去；
2TIM|4|11|只有 路加 在我這裏。你來的時候把 馬可 帶來，因為他在服事 上於我有益。
2TIM|4|12|我已經打發 推基古 往 以弗所 去。
2TIM|4|13|我在 特羅亞 留給 加布 的那件外衣，你來的時候要帶來，那些書也帶來，特別是那幾卷羊皮的書。
2TIM|4|14|銅匠 亞歷山大 多方害我；主必照他所行的報應他。
2TIM|4|15|你也要防備他，因為他極力抗拒我們的話。
2TIM|4|16|我初次上訴時，沒有人前來幫助，竟都離棄了我，但願這罪不歸在他們身上。
2TIM|4|17|惟有主站在我身邊，加給我力量，使我能把福音完整地傳開，讓所有的外邦人都聽見；我也從獅子口裏被救出來。
2TIM|4|18|主必救我脫離一切的兇惡，也必救我進他的天國。願榮耀歸給他，直到永永遠遠。阿們！
2TIM|4|19|請向 百基拉 、 亞居拉 和 阿尼色弗 一家的人問安。
2TIM|4|20|以拉都 在 哥林多 住下了。 特羅非摩 病了，我把他留在 米利都 。
2TIM|4|21|你要趕緊在冬天以前到我這裏來。 友布羅 、 布田 、 利奴 、 革老底亞 和眾弟兄都向你問安。
2TIM|4|22|願主與你的靈同在！願恩惠與你們同在！
