OBAD|1|1|Видіння Овдія. Так сказав Господь Бог на Едом: Почули ми вістку від Господа, і посланий був між народів посол, щоб сказати: Уставайте, і станьмо на нього до бою!
OBAD|1|2|Оце Я малим тебе дав між народи, ти дуже погорджений.
OBAD|1|3|Гордість серця твого обманила тебе, який перебуваєш по щілинах скельних, у високім сидінні своїм, що говориш у серці своєму: Хто скине на землю мене?
OBAD|1|4|Якщо б ти піднісся, немов той орел, і якщо б ти кубло своє склав поміж зорями, то й звідти Я скину тебе, промовляє Господь!
OBAD|1|5|Чи ж до тебе злодії приходили, чи нічні ті грабіжники, такий ти понищений! чи ж вони не накрали б собі скільки треба? Якщо б до тебе прийшли збирачі винограду, чи ж вони не лишили б хоч вибірків?
OBAD|1|6|Як Ісав перешуканий, як криївки його переглянені!
OBAD|1|7|Аж до границі прогнали тебе, обманять тебе твої всі союзники, переможуть тебе твої приятелі! Ті, що хліб твій їдять, пастку розставлять на тебе, нема в тому розуму!
OBAD|1|8|Чи ж не станеться це того дня, промовляє Господь, і вигублю Я мудреців із Едому, а розум з гори Ісавової?
OBAD|1|9|І настрашене буде лицарство твоє, о Темане, щоб був витятий кожен з Ісава убивством.
OBAD|1|10|Через насилля на Якова на брата твого сором покриє тебе, і ти витятий будеш навіки.
OBAD|1|11|Того дня, коли став ти навпроти, того дня, як чужі полонили були його військо, і коли чужинці в його брами ввійшли і жереба кидали про Єрусалим, то й ти був, як один з них!
OBAD|1|12|І тому не дивися на день свого брата, на день лиха його, і не тішся з Юдиних синів у день їхньої згуби, і не розкривай своїх уст у день утиску.
OBAD|1|13|І не входь ти до брами народу Мого у день лиха його, і не приглядайся до зла його й ти в день нещастя його, і не простягайте своєї руки до багатства його в день нещастя його!
OBAD|1|14|І на роздоріжжі не стій, щоб витинати його втікачів, і в день утиску не видавай його решток!
OBAD|1|15|Бо близький день Господній над усіма народами, як зробив ти, то так і тобі буде зроблено: вернеться на твою голову чин твій!
OBAD|1|16|Бо як ви пили на святій Моїй горі, так народи усі завжди питимуть! І будуть пити вони, і будуть хлептати, і стануть вони, немов їх не було.
OBAD|1|17|А на Сіонській горі буде спасіння, і буде святою вона, і спадки свої вже посяде дім Яковів.
OBAD|1|18|І дім Якова стане огнем, і дім Йосипа полум'ям, а дім Ісава соломою, і будуть палати вони проти них, і їх пожеруть, і останку не буде із дому Ісава, бо Господь це сказав.
OBAD|1|19|І посядуть південні Ісавову гору, а мешканці долин филистимлян, і посядуть Єфремове поле та поле самарійське, а Веніямин Ґілеад.
OBAD|1|20|А полонені війська Ізраїлевих синів заволодіють тим, що хананейське аж до Цорфату, а єрусалимські вигнанці в неволі, що в Сефараді, посядуть міста полудневі.
OBAD|1|21|І спасителі прийдуть на гору Сіон, щоб гору Ісава судити, і царство Господнє настане!
