HAB|1|1|哈巴谷 先知所看见的默示。
HAB|1|2|耶和华啊，我呼求， 你不应允，要到几时呢？ 我向你呼喊“暴力！” 你还不拯救？
HAB|1|3|你为何使我看见罪孽？ 你为何坐视奸恶呢？ 毁灭和凶暴在我面前， 争执与纷争不断发生。
HAB|1|4|因此律法无效， 公理从未彰显。 因恶人围困义人， 所以公理遭受扭曲。
HAB|1|5|你们要向列国观看 ，注意看， 要惊奇，再惊奇！ 因为在你们的日子，有一件事发生 ， 尽管有人说了，你们还是不信。
HAB|1|6|看哪，我必兴起 迦勒底 人， 就是那残忍暴躁之民，通行遍地， 霸占不属自己的住处。
HAB|1|7|他威武可畏， 审判与威权都由他而出。
HAB|1|8|他的马比豹更快， 比晚上 的野狼更猛。 他的战马跳跃， 他的战马从远方而来 ； 他们飞跑，如鹰急速抓食，
HAB|1|9|都为施行残暴而来， 他们的脸面向东 ， 聚集俘虏，多如尘沙。
HAB|1|10|他讥诮列王， 嘲讽领袖， 嗤笑一切堡垒， 堆土攻取它。
HAB|1|11|那时，他如风猛然扫过， 他背叛，显为有罪； 他以自己的力量为神明。
HAB|1|12|耶和华－我的上帝，我的圣者啊， 你不是从亘古就有吗？ 我们必不致死。 耶和华啊，你派他为要行审判； 磐石啊，你立他为要惩治人。
HAB|1|13|你的眼目清洁， 不看邪恶，也不看奸恶， 为何你却看着人行诡诈呢？ 恶人吞灭比自己公义的人， 为何你保持沉默呢？
HAB|1|14|你为何使人如海中的鱼， 又如无人管辖的爬行动物呢？
HAB|1|15|他用钩子把他们全拉上来， 用罗网捕获他们， 拉渔网聚集他们。 因此，他欢喜快乐，
HAB|1|16|向罗网献祭， 向渔网烧香； 因为他藉此得丰盛的收获 与肥美的食物。
HAB|1|17|但他岂可因此屡屡倒空罗网 ， 时常杀戮列国的人，毫不顾惜呢？
HAB|2|1|我要站在我的了望台， 立在城楼 上观看， 看耶和华要对我说什么， 我可用什么话向他诉冤。
HAB|2|2|耶和华回答我，说： 将这默示清楚地写在看板上， 使人容易朗读 。
HAB|2|3|因为这默示有一定日期， 论及终局，绝不落空。 它虽然耽延，你要等候； 因为它必临到，不再迟延。
HAB|2|4|看哪，恶人自高自大，心不正直； 惟义人必因他的信得生 。
HAB|2|5|他因酒诡诈、 狂傲、不安于位； 他张开喉咙 ，好像阴间， 如死亡不能知足， 他聚集万国， 招聚万民全归自己。
HAB|2|6|这些人岂不都要提起诗歌和俗语，嘲讽他说： 祸哉！你增添不属自己的财物， 靠押金发财，要到几时呢？
HAB|2|7|咬伤你的 岂不忽然兴起， 扰害你的岂不突然崛起， 你就成为他们的掳物吗？
HAB|2|8|因你抢夺许多国家， 流人的血，向土地、城镇和全城的居民施行残暴， 各国残存之民都必抢夺你。
HAB|2|9|祸哉！那为本家积蓄不义之财、 在高处搭窝、指望得免灾祸的人！
HAB|2|10|你图谋剪除许多民族，犯了罪， 使自己的家蒙羞，自害己命。
HAB|2|11|墙里的石头要呼叫， 屋内的栋梁必应声。
HAB|2|12|祸哉！那以鲜血建城、 以罪孽造镇的人！
HAB|2|13|看哪，这不都是 出于万军之耶和华吗？ 万民劳碌得来的被火焚烧， 万族辛苦建造的，归于虚空。
HAB|2|14|全地都必认识耶和华的荣耀， 好像水充满海洋一般。
HAB|2|15|祸哉！那给邻舍酒喝，加上毒物 ， 使人喝醉，为要看见他们下体的人！
HAB|2|16|你满受羞辱，不得荣耀； 你也喝吧，显明你是未受割礼的 ！ 耶和华右手的杯必传到你那里， 你的荣耀就变为羞辱。
HAB|2|17|黎巴嫩 所受的残暴必淹没你， 野兽所遭遇的毁灭使你惊吓 ； 因你流人的血， 向土地、城镇和全城的居民施行残暴。
HAB|2|18|偶像有什么益处呢？ 制造者雕刻它， 铸成偶像，作虚假的教师； 制造者倚靠的是自己所做的哑巴偶像。
HAB|2|19|祸哉！那对木头说“醒起”， 对哑巴石头说“起来”的人！ 偶像岂能教导人呢？ 看哪，它以金银包裹，其中并无气息。
HAB|2|20|惟耶和华在他的圣殿中， 全地都当在他面前肃静。
HAB|3|1|哈巴谷 先知的祷告，调用流离歌。
HAB|3|2|耶和华啊，我听见你的名声； 耶和华啊，我惧怕你的作为。 求你在这些年间 复兴你的作为， 在这些年间将它显明出来 ； 在发怒的时候以怜悯为念。
HAB|3|3|上帝从 提幔 而来， 圣者从 巴兰山 临到； 他的荣光遮蔽诸天， 颂赞遍满全地。
HAB|3|4|他的辉煌如同日光， 从他手里发出光芒， 那里 隐藏他的能力。
HAB|3|5|在他前面有瘟疫流行， 在他脚下有热症发出。
HAB|3|6|他站立，震动 大地， 他观看，震动列国。 永久的山崩裂， 长存的岭塌陷， 他的作为与古时一样。
HAB|3|7|我见 古珊 的帐棚遭难， 米甸 地的幔子动摇。
HAB|3|8|耶和华啊，你岂是向江河发怒， 向江河生气， 向海洋发烈怒吗？ 你骑在马上， 坐在得胜的战车上，
HAB|3|9|你的弓全然显露 ， 箭是发誓的言语 ； 你以江河分开大地。
HAB|3|10|山岭见你，无不战抖； 大水泛滥而过， 深渊发声， 汹涌翻腾 。
HAB|3|11|因你的箭射出光芒， 你的枪闪出光耀， 日月都停在原处。
HAB|3|12|你发怒遍行大地， 以怒气责打列国，如打谷一般。
HAB|3|13|你出来拯救你的百姓， 拯救你的受膏者； 你打破恶人之家的头， 暴露其根基，直到颈项 。
HAB|3|14|你以其戈矛刺透他战士的头； 他们如旋风将我 刮散， 他们喜爱暗中吞吃困苦的人。
HAB|3|15|你骑马践踏海， 践踏汹涌的大水。
HAB|3|16|我听见这声音，身体战兢， 嘴唇发颤， 骨中朽烂， 在所立之处战兢 ； 但我安静等候 灾难之日临到那上来侵犯我们的民 。
HAB|3|17|虽然无花果树不发旺， 葡萄树不结果， 橄榄树也不收成， 田地不出粮食， 圈中绝了羊， 棚内也没有牛；
HAB|3|18|然而，我要因耶和华欢欣， 因救我的上帝喜乐。
HAB|3|19|主耶和华是我的力量， 他使我的脚快如母鹿， 又使我稳行在高处。 这歌交给圣咏团长，用丝弦的乐器。
