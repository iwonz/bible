JOHN|1|1|В начале было Слово, и Слово было у Бога, и Слово было Бог.
JOHN|1|2|Оно было в начале у Бога.
JOHN|1|3|Все чрез Него начало быть, и без Него ничто не начало быть, что начало быть.
JOHN|1|4|В Нем была жизнь, и жизнь была свет человеков.
JOHN|1|5|И свет во тьме светит, и тьма не объяла его.
JOHN|1|6|Был человек, посланный от Бога; имя ему Иоанн.
JOHN|1|7|Он пришел для свидетельства, чтобы свидетельствовать о Свете, дабы все уверовали чрез него.
JOHN|1|8|Он не был свет, но [был послан], чтобы свидетельствовать о Свете.
JOHN|1|9|Был Свет истинный, Который просвещает всякого человека, приходящего в мир.
JOHN|1|10|В мире был, и мир чрез Него начал быть, и мир Его не познал.
JOHN|1|11|Пришел к своим, и свои Его не приняли.
JOHN|1|12|А тем, которые приняли Его, верующим во имя Его, дал власть быть чадами Божиими,
JOHN|1|13|которые ни от крови, ни от хотения плоти, ни от хотения мужа, но от Бога родились.
JOHN|1|14|И Слово стало плотию, и обитало с нами, полное благодати и истины; и мы видели славу Его, славу, как Единородного от Отца.
JOHN|1|15|Иоанн свидетельствует о Нем и, восклицая, говорит: Сей был Тот, о Котором я сказал, что Идущий за мною стал впереди меня, потому что был прежде меня.
JOHN|1|16|И от полноты Его все мы приняли и благодать на благодать,
JOHN|1|17|ибо закон дан чрез Моисея; благодать же и истина произошли чрез Иисуса Христа.
JOHN|1|18|Бога не видел никто никогда; Единородный Сын, сущий в недре Отчем, Он явил.
JOHN|1|19|И вот свидетельство Иоанна, когда Иудеи прислали из Иерусалима священников и левитов спросить его: кто ты?
JOHN|1|20|Он объявил, и не отрекся, и объявил, что я не Христос.
JOHN|1|21|И спросили его: что же? ты Илия? Он сказал: нет. Пророк? Он отвечал: нет.
JOHN|1|22|Сказали ему: кто же ты? чтобы нам дать ответ пославшим нас: что ты скажешь о себе самом?
JOHN|1|23|Он сказал: я глас вопиющего в пустыне: исправьте путь Господу, как сказал пророк Исаия.
JOHN|1|24|А посланные были из фарисеев;
JOHN|1|25|И они спросили его: что же ты крестишь, если ты ни Христос, ни Илия, ни пророк?
JOHN|1|26|Иоанн сказал им в ответ: я крещу в воде; но стоит среди вас [Некто], Которого вы не знаете.
JOHN|1|27|Он–то Идущий за мною, но Который стал впереди меня. Я недостоин развязать ремень у обуви Его.
JOHN|1|28|Это происходило в Вифаваре при Иордане, где крестил Иоанн.
JOHN|1|29|На другой день видит Иоанн идущего к нему Иисуса и говорит: вот Агнец Божий, Который берет [на Себя] грех мира.
JOHN|1|30|Сей есть, о Котором я сказал: за мною идет Муж, Который стал впереди меня, потому что Он был прежде меня.
JOHN|1|31|Я не знал Его; но для того пришел крестить в воде, чтобы Он явлен был Израилю.
JOHN|1|32|И свидетельствовал Иоанн, говоря: я видел Духа, сходящего с неба, как голубя, и пребывающего на Нем.
JOHN|1|33|Я не знал Его; но Пославший меня крестить в воде сказал мне: на Кого увидишь Духа сходящего и пребывающего на Нем, Тот есть крестящий Духом Святым.
JOHN|1|34|И я видел и засвидетельствовал, что Сей есть Сын Божий.
JOHN|1|35|На другой день опять стоял Иоанн и двое из учеников его.
JOHN|1|36|И, увидев идущего Иисуса, сказал: вот Агнец Божий.
JOHN|1|37|Услышав от него сии слова, оба ученика пошли за Иисусом.
JOHN|1|38|Иисус же, обратившись и увидев их идущих, говорит им: что вам надобно? Они сказали Ему: Равви, – что значит: учитель, – где живешь?
JOHN|1|39|Говорит им: пойдите и увидите. Они пошли и увидели, где Он живет; и пробыли у Него день тот. Было около десятого часа.
JOHN|1|40|Один из двух, слышавших от Иоанна [об Иисусе] и последовавших за Ним, был Андрей, брат Симона Петра.
JOHN|1|41|Он первый находит брата своего Симона и говорит ему: мы нашли Мессию, что значит: Христос;
JOHN|1|42|и привел его к Иисусу. Иисус же, взглянув на него, сказал: ты – Симон, сын Ионин; ты наречешься Кифа, что значит: камень Петр.
JOHN|1|43|На другой день [Иисус] восхотел идти в Галилею, и находит Филиппа и говорит ему: иди за Мною.
JOHN|1|44|Филипп же был из Вифсаиды, из [одного] города с Андреем и Петром.
JOHN|1|45|Филипп находит Нафанаила и говорит ему: мы нашли Того, о Котором писали Моисей в законе и пророки, Иисуса, сына Иосифова, из Назарета.
JOHN|1|46|Но Нафанаил сказал ему: из Назарета может ли быть что доброе? Филипп говорит ему: пойди и посмотри.
JOHN|1|47|Иисус, увидев идущего к Нему Нафанаила, говорит о нем: вот подлинно Израильтянин, в котором нет лукавства.
JOHN|1|48|Нафанаил говорит Ему: почему Ты знаешь меня? Иисус сказал ему в ответ: прежде нежели позвал тебя Филипп, когда ты был под смоковницею, Я видел тебя.
JOHN|1|49|Нафанаил отвечал Ему: Равви! Ты Сын Божий, Ты Царь Израилев.
JOHN|1|50|Иисус сказал ему в ответ: ты веришь, потому что Я тебе сказал: Я видел тебя под смоковницею; увидишь больше сего.
JOHN|1|51|И говорит ему: истинно, истинно говорю вам: отныне будете видеть небо отверстым и Ангелов Божиих восходящих и нисходящих к Сыну Человеческому.
JOHN|2|1|На третий день был брак в Кане Галилейской, и Матерь Иисуса была там.
JOHN|2|2|Был также зван Иисус и ученики Его на брак.
JOHN|2|3|И как недоставало вина, то Матерь Иисуса говорит Ему: вина нет у них.
JOHN|2|4|Иисус говорит Ей: что Мне и Тебе, Жено? еще не пришел час Мой.
JOHN|2|5|Матерь Его сказала служителям: что скажет Он вам, то сделайте.
JOHN|2|6|Было же тут шесть каменных водоносов, стоявших [по обычаю] очищения Иудейского, вмещавших по две или по три меры.
JOHN|2|7|Иисус говорит им: наполните сосуды водою. И наполнили их до верха.
JOHN|2|8|И говорит им: теперь почерпните и несите к распорядителю пира. И понесли.
JOHN|2|9|Когда же распорядитель отведал воды, сделавшейся вином, – а он не знал, откуда [это вино], знали только служители, почерпавшие воду, – тогда распорядитель зовет жениха
JOHN|2|10|и говорит ему: всякий человек подает сперва хорошее вино, а когда напьются, тогда худшее; а ты хорошее вино сберег доселе.
JOHN|2|11|Так положил Иисус начало чудесам в Кане Галилейской и явил славу Свою; и уверовали в Него ученики Его.
JOHN|2|12|После сего пришел Он в Капернаум, Сам и Матерь Его, и братья его, и ученики Его; и там пробыли немного дней.
JOHN|2|13|Приближалась Пасха Иудейская, и Иисус пришел в Иерусалим
JOHN|2|14|и нашел, что в храме продавали волов, овец и голубей, и сидели меновщики денег.
JOHN|2|15|И, сделав бич из веревок, выгнал из храма всех, [также] и овец и волов; и деньги у меновщиков рассыпал, а столы их опрокинул.
JOHN|2|16|И сказал продающим голубей: возьмите это отсюда и дома Отца Моего не делайте домом торговли.
JOHN|2|17|При сем ученики Его вспомнили, что написано: ревность по доме Твоем снедает Меня.
JOHN|2|18|На это Иудеи сказали: каким знамением докажешь Ты нам, что [имеешь] [власть] так поступать?
JOHN|2|19|Иисус сказал им в ответ: разрушьте храм сей, и Я в три дня воздвигну его.
JOHN|2|20|На это сказали Иудеи: сей храм строился сорок шесть лет, и Ты в три дня воздвигнешь его?
JOHN|2|21|А Он говорил о храме тела Своего.
JOHN|2|22|Когда же воскрес Он из мертвых, то ученики Его вспомнили, что Он говорил это, и поверили Писанию и слову, которое сказал Иисус.
JOHN|2|23|И когда Он был в Иерусалиме на празднике Пасхи, то многие, видя чудеса, которые Он творил, уверовали во имя Его.
JOHN|2|24|Но Сам Иисус не вверял Себя им, потому что знал всех
JOHN|2|25|и не имел нужды, чтобы кто засвидетельствовал о человеке, ибо Сам знал, что в человеке.
JOHN|3|1|Между фарисеями был некто, именем Никодим, [один] из начальников Иудейских.
JOHN|3|2|Он пришел к Иисусу ночью и сказал Ему: Равви! мы знаем, что Ты учитель, пришедший от Бога; ибо таких чудес, какие Ты творишь, никто не может творить, если не будет с ним Бог.
JOHN|3|3|Иисус сказал ему в ответ: истинно, истинно говорю тебе, если кто не родится свыше, не может увидеть Царствия Божия.
JOHN|3|4|Никодим говорит Ему: как может человек родиться, будучи стар? неужели может он в другой раз войти в утробу матери своей и родиться?
JOHN|3|5|Иисус отвечал: истинно, истинно говорю тебе, если кто не родится от воды и Духа, не может войти в Царствие Божие.
JOHN|3|6|Рожденное от плоти есть плоть, а рожденное от Духа есть дух.
JOHN|3|7|Не удивляйся тому, что Я сказал тебе: должно вам родиться свыше.
JOHN|3|8|Дух дышит, где хочет, и голос его слышишь, а не знаешь, откуда приходит и куда уходит: так бывает со всяким, рожденным от Духа.
JOHN|3|9|Никодим сказал Ему в ответ: как это может быть?
JOHN|3|10|Иисус отвечал и сказал ему: ты – учитель Израилев, и этого ли не знаешь?
JOHN|3|11|Истинно, истинно говорю тебе: мы говорим о том, что знаем, и свидетельствуем о том, что видели, а вы свидетельства Нашего не принимаете.
JOHN|3|12|Если Я сказал вам о земном, и вы не верите, – как поверите, если буду говорить вам о небесном?
JOHN|3|13|Никто не восходил на небо, как только сшедший с небес Сын Человеческий, сущий на небесах.
JOHN|3|14|И как Моисей вознес змию в пустыне, так должно вознесену быть Сыну Человеческому,
JOHN|3|15|дабы всякий, верующий в Него, не погиб, но имел жизнь вечную.
JOHN|3|16|Ибо так возлюбил Бог мир, что отдал Сына Своего Единородного, дабы всякий верующий в Него, не погиб, но имел жизнь вечную.
JOHN|3|17|Ибо не послал Бог Сына Своего в мир, чтобы судить мир, но чтобы мир спасен был чрез Него.
JOHN|3|18|Верующий в Него не судится, а неверующий уже осужден, потому что не уверовал во имя Единородного Сына Божия.
JOHN|3|19|Суд же состоит в том, что свет пришел в мир; но люди более возлюбили тьму, нежели свет, потому что дела их были злы;
JOHN|3|20|ибо всякий, делающий злое, ненавидит свет и не идет к свету, чтобы не обличились дела его, потому что они злы,
JOHN|3|21|а поступающий по правде идет к свету, дабы явны были дела его, потому что они в Боге соделаны.
JOHN|3|22|После сего пришел Иисус с учениками Своими в землю Иудейскую и там жил с ними и крестил.
JOHN|3|23|А Иоанн также крестил в Еноне, близ Салима, потому что там было много воды; и приходили [туда] и крестились,
JOHN|3|24|ибо Иоанн еще не был заключен в темницу.
JOHN|3|25|Тогда у Иоанновых учеников произошел спор с Иудеями об очищении.
JOHN|3|26|И пришли к Иоанну и сказали ему: равви! Тот, Который был с тобою при Иордане и о Котором ты свидетельствовал, вот Он крестит, и все идут к Нему.
JOHN|3|27|Иоанн сказал в ответ: не может человек ничего принимать [на] [себя], если не будет дано ему с неба.
JOHN|3|28|Вы сами мне свидетели в том, что я сказал: не я Христос, но я послан пред Ним.
JOHN|3|29|Имеющий невесту есть жених, а друг жениха, стоящий и внимающий ему, радостью радуется, слыша голос жениха. Сия–то радость моя исполнилась.
JOHN|3|30|Ему должно расти, а мне умаляться.
JOHN|3|31|Приходящий свыше и есть выше всех; а сущий от земли земной и есть и говорит, как сущий от земли; Приходящий с небес есть выше всех,
JOHN|3|32|и что Он видел и слышал, о том и свидетельствует; и никто не принимает свидетельства Его.
JOHN|3|33|Принявший Его свидетельство сим запечатлел, что Бог истинен,
JOHN|3|34|ибо Тот, Которого послал Бог, говорит слова Божии; ибо не мерою дает Бог Духа.
JOHN|3|35|Отец любит Сына и все дал в руку Его.
JOHN|3|36|Верующий в Сына имеет жизнь вечную, а не верующий в Сына не увидит жизни, но гнев Божий пребывает на нем.
JOHN|4|1|Когда же узнал Иисус о [дошедшем до] фарисеев слухе, что Он более приобретает учеников и крестит, нежели Иоанн, –
JOHN|4|2|хотя Сам Иисус не крестил, а ученики Его, –
JOHN|4|3|то оставил Иудею и пошел опять в Галилею.
JOHN|4|4|Надлежало же Ему проходить через Самарию.
JOHN|4|5|Итак приходит Он в город Самарийский, называемый Сихарь, близ участка земли, данного Иаковом сыну своему Иосифу.
JOHN|4|6|Там был колодезь Иаковлев. Иисус, утрудившись от пути, сел у колодезя. Было около шестого часа.
JOHN|4|7|Приходит женщина из Самарии почерпнуть воды. Иисус говорит ей: дай Мне пить.
JOHN|4|8|Ибо ученики Его отлучились в город купить пищи.
JOHN|4|9|Женщина Самарянская говорит Ему: как ты, будучи Иудей, просишь пить у меня, Самарянки? ибо Иудеи с Самарянами не сообщаются.
JOHN|4|10|Иисус сказал ей в ответ: если бы ты знала дар Божий и Кто говорит тебе: дай Мне пить, то ты сама просила бы у Него, и Он дал бы тебе воду живую.
JOHN|4|11|Женщина говорит Ему: господин! тебе и почерпнуть нечем, а колодезь глубок; откуда же у тебя вода живая?
JOHN|4|12|Неужели ты больше отца нашего Иакова, который дал нам этот колодезь и сам из него пил, и дети его, и скот его?
JOHN|4|13|Иисус сказал ей в ответ: всякий, пьющий воду сию, возжаждет опять,
JOHN|4|14|а кто будет пить воду, которую Я дам ему, тот не будет жаждать вовек; но вода, которую Я дам ему, сделается в нем источником воды, текущей в жизнь вечную.
JOHN|4|15|Женщина говорит Ему: господин! дай мне этой воды, чтобы мне не иметь жажды и не приходить сюда черпать.
JOHN|4|16|Иисус говорит ей: пойди, позови мужа твоего и приди сюда.
JOHN|4|17|Женщина сказала в ответ: у меня нет мужа. Иисус говорит ей: правду ты сказала, что у тебя нет мужа,
JOHN|4|18|ибо у тебя было пять мужей, и тот, которого ныне имеешь, не муж тебе; это справедливо ты сказала.
JOHN|4|19|Женщина говорит Ему: Господи! вижу, что Ты пророк.
JOHN|4|20|Отцы наши поклонялись на этой горе, а вы говорите, что место, где должно поклоняться, находится в Иерусалиме.
JOHN|4|21|Иисус говорит ей: поверь Мне, что наступает время, когда и не на горе сей, и не в Иерусалиме будете поклоняться Отцу.
JOHN|4|22|Вы не знаете, чему кланяетесь, а мы знаем, чему кланяемся, ибо спасение от Иудеев.
JOHN|4|23|Но настанет время и настало уже, когда истинные поклонники будут поклоняться Отцу в духе и истине, ибо таких поклонников Отец ищет Себе.
JOHN|4|24|Бог есть дух, и поклоняющиеся Ему должны поклоняться в духе и истине.
JOHN|4|25|Женщина говорит Ему: знаю, что придет Мессия, то есть Христос; когда Он придет, то возвестит нам все.
JOHN|4|26|Иисус говорит ей: это Я, Который говорю с тобою.
JOHN|4|27|В это время пришли ученики Его, и удивились, что Он разговаривал с женщиною; однакож ни один не сказал: чего Ты требуешь? или: о чем говоришь с нею?
JOHN|4|28|Тогда женщина оставила водонос свой и пошла в город, и говорит людям:
JOHN|4|29|пойдите, посмотрите Человека, Который сказал мне все, что я сделала: не Он ли Христос?
JOHN|4|30|Они вышли из города и пошли к Нему.
JOHN|4|31|Между тем ученики просили Его, говоря: Равви! ешь.
JOHN|4|32|Но Он сказал им: у Меня есть пища, которой вы не знаете.
JOHN|4|33|Посему ученики говорили между собою: разве кто принес Ему есть?
JOHN|4|34|Иисус говорит им: Моя пища есть творить волю Пославшего Меня и совершить дело Его.
JOHN|4|35|Не говорите ли вы, что еще четыре месяца, и наступит жатва? А Я говорю вам: возведите очи ваши и посмотрите на нивы, как они побелели и поспели к жатве.
JOHN|4|36|Жнущий получает награду и собирает плод в жизнь вечную, так что и сеющий и жнущий вместе радоваться будут,
JOHN|4|37|ибо в этом случае справедливо изречение: один сеет, а другой жнет.
JOHN|4|38|Я послал вас жать то, над чем вы не трудились: другие трудились, а вы вошли в труд их.
JOHN|4|39|И многие Самаряне из города того уверовали в Него по слову женщины, свидетельствовавшей, что Он сказал ей все, что она сделала.
JOHN|4|40|И потому, когда пришли к Нему Самаряне, то просили Его побыть у них; и Он пробыл там два дня.
JOHN|4|41|И еще большее число уверовали по Его слову.
JOHN|4|42|А женщине той говорили: уже не по твоим речам веруем, ибо сами слышали и узнали, что Он истинно Спаситель мира, Христос.
JOHN|4|43|По прошествии же двух дней Он вышел оттуда и пошел в Галилею,
JOHN|4|44|ибо Сам Иисус свидетельствовал, что пророк не имеет чести в своем отечестве.
JOHN|4|45|Когда пришел Он в Галилею, то Галилеяне приняли Его, видев все, что Он сделал в Иерусалиме в праздник, – ибо и они ходили на праздник.
JOHN|4|46|Итак Иисус опять пришел в Кану Галилейскую, где претворил воду в вино. В Капернауме был некоторый царедворец, у которого сын был болен.
JOHN|4|47|Он, услышав, что Иисус пришел из Иудеи в Галилею, пришел к Нему и просил Его придти и исцелить сына его, который был при смерти.
JOHN|4|48|Иисус сказал ему: вы не уверуете, если не увидите знамений и чудес.
JOHN|4|49|Царедворец говорит Ему: Господи! приди, пока не умер сын мой.
JOHN|4|50|Иисус говорит ему: пойди, сын твой здоров. Он поверил слову, которое сказал ему Иисус, и пошел.
JOHN|4|51|На дороге встретили его слуги его и сказали: сын твой здоров.
JOHN|4|52|Он спросил у них: в котором часу стало ему легче? Ему сказали: вчера в седьмом часу горячка оставила его.
JOHN|4|53|Из этого отец узнал, что это был тот час, в который Иисус сказал ему: сын твой здоров, и уверовал сам и весь дом его.
JOHN|4|54|Это второе чудо сотворил Иисус, возвратившись из Иудеи в Галилею.
JOHN|5|1|После сего был праздник Иудейский, и пришел Иисус в Иерусалим.
JOHN|5|2|Есть же в Иерусалиме у Овечьих [ворот] купальня, называемая по–еврейски Вифезда, при которой было пять крытых ходов.
JOHN|5|3|В них лежало великое множество больных, слепых, хромых, иссохших, ожидающих движения воды,
JOHN|5|4|ибо Ангел Господень по временам сходил в купальню и возмущал воду, и кто первый входил [в нее] по возмущении воды, тот выздоравливал, какою бы ни был одержим болезнью.
JOHN|5|5|Тут был человек, находившийся в болезни тридцать восемь лет.
JOHN|5|6|Иисус, увидев его лежащего и узнав, что он лежит уже долгое время, говорит ему: хочешь ли быть здоров?
JOHN|5|7|Больной отвечал Ему: так, Господи; но не имею человека, который опустил бы меня в купальню, когда возмутится вода; когда же я прихожу, другой уже сходит прежде меня.
JOHN|5|8|Иисус говорит ему: встань, возьми постель твою и ходи.
JOHN|5|9|И он тотчас выздоровел, и взял постель свою и пошел. Было же это в день субботний.
JOHN|5|10|Посему Иудеи говорили исцеленному: сегодня суббота; не должно тебе брать постели.
JOHN|5|11|Он отвечал им: Кто меня исцелил, Тот мне сказал: возьми постель твою и ходи.
JOHN|5|12|Его спросили: кто Тот Человек, Который сказал тебе: возьми постель твою и ходи?
JOHN|5|13|Исцеленный же не знал, кто Он, ибо Иисус скрылся в народе, бывшем на том месте.
JOHN|5|14|Потом Иисус встретил его в храме и сказал ему: вот, ты выздоровел; не греши больше, чтобы не случилось с тобою чего хуже.
JOHN|5|15|Человек сей пошел и объявил Иудеям, что исцеливший его есть Иисус.
JOHN|5|16|И стали Иудеи гнать Иисуса и искали убить Его за то, что Он делал такие [дела] в субботу.
JOHN|5|17|Иисус же говорил им: Отец Мой доныне делает, и Я делаю.
JOHN|5|18|И еще более искали убить Его Иудеи за то, что Он не только нарушал субботу, но и Отцем Своим называл Бога, делая Себя равным Богу.
JOHN|5|19|На это Иисус сказал: истинно, истинно говорю вам: Сын ничего не может творить Сам от Себя, если не увидит Отца творящего: ибо, что творит Он, то и Сын творит также.
JOHN|5|20|Ибо Отец любит Сына и показывает Ему все, что творит Сам; и покажет Ему дела больше сих, так что вы удивитесь.
JOHN|5|21|Ибо, как Отец воскрешает мертвых и оживляет, так и Сын оживляет, кого хочет.
JOHN|5|22|Ибо Отец и не судит никого, но весь суд отдал Сыну,
JOHN|5|23|дабы все чтили Сына, как чтут Отца. Кто не чтит Сына, тот не чтит и Отца, пославшего Его.
JOHN|5|24|Истинно, истинно говорю вам: слушающий слово Мое и верующий в Пославшего Меня имеет жизнь вечную, и на суд не приходит, но перешел от смерти в жизнь.
JOHN|5|25|Истинно, истинно говорю вам: наступает время, и настало уже, когда мертвые услышат глас Сына Божия и, услышав, оживут.
JOHN|5|26|Ибо, как Отец имеет жизнь в Самом Себе, так и Сыну дал иметь жизнь в Самом Себе.
JOHN|5|27|И дал Ему власть производить и суд, потому что Он есть Сын Человеческий.
JOHN|5|28|Не дивитесь сему; ибо наступает время, в которое все, находящиеся в гробах, услышат глас Сына Божия;
JOHN|5|29|и изыдут творившие добро в воскресение жизни, а делавшие зло – в воскресение осуждения.
JOHN|5|30|Я ничего не могу творить Сам от Себя. Как слышу, так и сужу, и суд Мой праведен; ибо не ищу Моей воли, но воли пославшего Меня Отца.
JOHN|5|31|Если Я свидетельствую Сам о Себе, то свидетельство Мое не есть истинно.
JOHN|5|32|Есть другой, свидетельствующий о Мне; и Я знаю, что истинно то свидетельство, которым он свидетельствует о Мне.
JOHN|5|33|Вы посылали к Иоанну, и он засвидетельствовал об истине.
JOHN|5|34|Впрочем Я не от человека принимаю свидетельство, но говорю это для того, чтобы вы спаслись.
JOHN|5|35|Он был светильник, горящий и светящий; а вы хотели малое время порадоваться при свете его.
JOHN|5|36|Я же имею свидетельство больше Иоаннова: ибо дела, которые Отец дал Мне совершить, самые дела сии, Мною творимые, свидетельствуют о Мне, что Отец послал Меня.
JOHN|5|37|И пославший Меня Отец Сам засвидетельствовал о Мне. А вы ни гласа Его никогда не слышали, ни лица Его не видели;
JOHN|5|38|и не имеете слова Его пребывающего в вас, потому что вы не веруете Тому, Которого Он послал.
JOHN|5|39|Исследуйте Писания, ибо вы думаете чрез них иметь жизнь вечную; а они свидетельствуют о Мне.
JOHN|5|40|Но вы не хотите придти ко Мне, чтобы иметь жизнь.
JOHN|5|41|Не принимаю славы от человеков,
JOHN|5|42|но знаю вас: вы не имеете в себе любви к Богу.
JOHN|5|43|Я пришел во имя Отца Моего, и не принимаете Меня; а если иной придет во имя свое, его примете.
JOHN|5|44|Как вы можете веровать, когда друг от друга принимаете славу, а славы, которая от Единого Бога, не ищете?
JOHN|5|45|Не думайте, что Я буду обвинять вас пред Отцем: есть на вас обвинитель Моисей, на которого вы уповаете.
JOHN|5|46|Ибо если бы вы верили Моисею, то поверили бы и Мне, потому что он писал о Мне.
JOHN|5|47|Если же его писаниям не верите, как поверите Моим словам?
JOHN|6|1|После сего пошел Иисус на ту сторону моря Галилейского, [в] [окрестности] Тивериады.
JOHN|6|2|За Ним последовало множество народа, потому что видели чудеса, которые Он творил над больными.
JOHN|6|3|Иисус взошел на гору и там сидел с учениками Своими.
JOHN|6|4|Приближалась же Пасха, праздник Иудейский.
JOHN|6|5|Иисус, возведя очи и увидев, что множество народа идет к Нему, говорит Филиппу: где нам купить хлебов, чтобы их накормить?
JOHN|6|6|Говорил же это, испытывая его; ибо Сам знал, что хотел сделать.
JOHN|6|7|Филипп отвечал Ему: им на двести динариев не довольно будет хлеба, чтобы каждому из них досталось хотя понемногу.
JOHN|6|8|Один из учеников Его, Андрей, брат Симона Петра, говорит Ему:
JOHN|6|9|здесь есть у одного мальчика пять хлебов ячменных и две рыбки; но что это для такого множества?
JOHN|6|10|Иисус сказал: велите им возлечь. Было же на том месте много травы. Итак возлегло людей числом около пяти тысяч.
JOHN|6|11|Иисус, взяв хлебы и воздав благодарение, роздал ученикам, а ученики возлежавшим, также и рыбы, сколько кто хотел.
JOHN|6|12|И когда насытились, то сказал ученикам Своим: соберите оставшиеся куски, чтобы ничего не пропало.
JOHN|6|13|И собрали, и наполнили двенадцать коробов кусками от пяти ячменных хлебов, оставшимися у тех, которые ели.
JOHN|6|14|Тогда люди, видевшие чудо, сотворенное Иисусом, сказали: это истинно Тот Пророк, Которому должно придти в мир.
JOHN|6|15|Иисус же, узнав, что хотят придти, нечаянно взять его и сделать царем, опять удалился на гору один.
JOHN|6|16|Когда же настал вечер, то ученики Его сошли к морю
JOHN|6|17|и, войдя в лодку, отправились на ту сторону моря, в Капернаум. Становилось темно, а Иисус не приходил к ним.
JOHN|6|18|Дул сильный ветер, и море волновалось.
JOHN|6|19|Проплыв около двадцати пяти или тридцати стадий, они увидели Иисуса, идущего по морю и приближающегося к лодке, и испугались.
JOHN|6|20|Но Он сказал им: это Я; не бойтесь.
JOHN|6|21|Они хотели принять Его в лодку; и тотчас лодка пристала к берегу, куда плыли.
JOHN|6|22|На другой день народ, стоявший по ту сторону моря, видел, что там, кроме одной лодки, в которую вошли ученики Его, иной не было, и что Иисус не входил в лодку с учениками Своими, а отплыли одни ученики Его.
JOHN|6|23|Между тем пришли из Тивериады другие лодки близко к тому месту, где ели хлеб по благословении Господнем.
JOHN|6|24|Итак, когда народ увидел, что тут нет Иисуса, ни учеников Его, то вошли в лодки и приплыли в Капернаум, ища Иисуса.
JOHN|6|25|И, найдя Его на той стороне моря, сказали Ему: Равви! когда Ты сюда пришел?
JOHN|6|26|Иисус сказал им в ответ: истинно, истинно говорю вам: вы ищете Меня не потому, что видели чудеса, но потому, что ели хлеб и насытились.
JOHN|6|27|Старайтесь не о пище тленной, но о пище, пребывающей в жизнь вечную, которую даст вам Сын Человеческий, ибо на Нем положил печать [Свою] Отец, Бог.
JOHN|6|28|Итак сказали Ему: что нам делать, чтобы творить дела Божии?
JOHN|6|29|Иисус сказал им в ответ: вот дело Божие, чтобы вы веровали в Того, Кого Он послал.
JOHN|6|30|На это сказали Ему: какое же Ты дашь знамение, чтобы мы увидели и поверили Тебе? что Ты делаешь?
JOHN|6|31|Отцы наши ели манну в пустыне, как написано: хлеб с неба дал им есть.
JOHN|6|32|Иисус же сказал им: истинно, истинно говорю вам: не Моисей дал вам хлеб с неба, а Отец Мой дает вам истинный хлеб с небес.
JOHN|6|33|Ибо хлеб Божий есть тот, который сходит с небес и дает жизнь миру.
JOHN|6|34|На это сказали Ему: Господи! подавай нам всегда такой хлеб.
JOHN|6|35|Иисус же сказал им: Я есмь хлеб жизни; приходящий ко Мне не будет алкать, и верующий в Меня не будет жаждать никогда.
JOHN|6|36|Но Я сказал вам, что вы и видели Меня, и не веруете.
JOHN|6|37|Все, что дает Мне Отец, ко Мне придет; и приходящего ко Мне не изгоню вон,
JOHN|6|38|ибо Я сошел с небес не для того, чтобы творить волю Мою, но волю пославшего Меня Отца.
JOHN|6|39|Воля же пославшего Меня Отца есть та, чтобы из того, что Он Мне дал, ничего не погубить, но все то воскресить в последний день.
JOHN|6|40|Воля Пославшего Меня есть та, чтобы всякий, видящий Сына и верующий в Него, имел жизнь вечную; и Я воскрешу его в последний день.
JOHN|6|41|Возроптали на Него Иудеи за то, что Он сказал: Я есмь хлеб, сшедший с небес.
JOHN|6|42|И говорили: не Иисус ли это, сын Иосифов, Которого отца и Мать мы знаем? Как же говорит Он: я сшел с небес?
JOHN|6|43|Иисус сказал им в ответ: не ропщите между собою.
JOHN|6|44|Никто не может придти ко Мне, если не привлечет его Отец, пославший Меня; и Я воскрешу его в последний день.
JOHN|6|45|У пророков написано: и будут все научены Богом. Всякий, слышавший от Отца и научившийся, приходит ко Мне.
JOHN|6|46|Это не то, чтобы кто видел Отца, кроме Того, Кто есть от Бога; Он видел Отца.
JOHN|6|47|Истинно, истинно говорю вам: верующий в Меня имеет жизнь вечную.
JOHN|6|48|Я есмь хлеб жизни.
JOHN|6|49|Отцы ваши ели манну в пустыне и умерли;
JOHN|6|50|хлеб же, сходящий с небес, таков, что ядущий его не умрет.
JOHN|6|51|Я хлеб живый, сшедший с небес; ядущий хлеб сей будет жить вовек; хлеб же, который Я дам, есть Плоть Моя, которую Я отдам за жизнь мира.
JOHN|6|52|Тогда Иудеи стали спорить между собою, говоря: как Он может дать нам есть Плоть Свою?
JOHN|6|53|Иисус же сказал им: истинно, истинно говорю вам: если не будете есть Плоти Сына Человеческого и пить Крови Его, то не будете иметь в себе жизни.
JOHN|6|54|Ядущий Мою Плоть и пиющий Мою Кровь имеет жизнь вечную, и Я воскрешу его в последний день.
JOHN|6|55|Ибо Плоть Моя истинно есть пища, и Кровь Моя истинно есть питие.
JOHN|6|56|Ядущий Мою Плоть и пиющий Мою Кровь пребывает во Мне, и Я в нем.
JOHN|6|57|Как послал Меня живый Отец, и Я живу Отцем, [так] и ядущий Меня жить будет Мною.
JOHN|6|58|Сей–то есть хлеб, сшедший с небес. Не так, как отцы ваши ели манну и умерли: ядущий хлеб сей жить будет вовек.
JOHN|6|59|Сие говорил Он в синагоге, уча в Капернауме.
JOHN|6|60|Многие из учеников Его, слыша то, говорили: какие странные слова! кто может это слушать?
JOHN|6|61|Но Иисус, зная Сам в Себе, что ученики Его ропщут на то, сказал им: это ли соблазняет вас?
JOHN|6|62|Что ж, если увидите Сына Человеческого восходящего [туда], где был прежде?
JOHN|6|63|Дух животворит; плоть не пользует нимало. Слова, которые говорю Я вам, суть дух и жизнь.
JOHN|6|64|Но есть из вас некоторые неверующие. Ибо Иисус от начала знал, кто суть неверующие и кто предаст Его.
JOHN|6|65|И сказал: для того–то и говорил Я вам, что никто не может придти ко Мне, если то не дано будет ему от Отца Моего.
JOHN|6|66|С этого времени многие из учеников Его отошли от Него и уже не ходили с Ним.
JOHN|6|67|Тогда Иисус сказал двенадцати: не хотите ли и вы отойти?
JOHN|6|68|Симон Петр отвечал Ему: Господи! к кому нам идти? Ты имеешь глаголы вечной жизни:
JOHN|6|69|и мы уверовали и познали, что Ты Христос, Сын Бога живаго.
JOHN|6|70|Иисус отвечал им: не двенадцать ли вас избрал Я? но один из вас диавол.
JOHN|6|71|Это говорил Он об Иуде Симонове Искариоте, ибо сей хотел предать Его, будучи один из двенадцати.
JOHN|7|1|После сего Иисус ходил по Галилее, ибо по Иудее не хотел ходить, потому что Иудеи искали убить Его.
JOHN|7|2|Приближался праздник Иудейский – поставление кущей.
JOHN|7|3|Тогда братья Его сказали Ему: выйди отсюда и пойди в Иудею, чтобы и ученики Твои видели дела, которые Ты делаешь.
JOHN|7|4|Ибо никто не делает чего–либо втайне, и ищет сам быть известным. Если Ты творишь такие дела, то яви Себя миру.
JOHN|7|5|Ибо и братья Его не веровали в Него.
JOHN|7|6|На это Иисус сказал им: Мое время еще не настало, а для вас всегда время.
JOHN|7|7|Вас мир не может ненавидеть, а Меня ненавидит, потому что Я свидетельствую о нем, что дела его злы.
JOHN|7|8|Вы пойдите на праздник сей; а Я еще не пойду на сей праздник, потому что Мое время еще не исполнилось.
JOHN|7|9|Сие сказав им, остался в Галилее.
JOHN|7|10|Но когда пришли братья Его, тогда и Он пришел на праздник не явно, а как бы тайно.
JOHN|7|11|Иудеи же искали Его на празднике и говорили: где Он?
JOHN|7|12|И много толков было о Нем в народе: одни говорили, что Он добр; а другие говорили: нет, но обольщает народ.
JOHN|7|13|Впрочем никто не говорил о Нем явно, боясь Иудеев.
JOHN|7|14|Но в половине уже праздника вошел Иисус в храм и учил.
JOHN|7|15|И дивились Иудеи, говоря: как Он знает Писания, не учившись?
JOHN|7|16|Иисус, отвечая им, сказал: Мое учение – не Мое, но Пославшего Меня;
JOHN|7|17|кто хочет творить волю Его, тот узнает о сем учении, от Бога ли оно, или Я Сам от Себя говорю.
JOHN|7|18|Говорящий сам от себя ищет славы себе; а Кто ищет славы Пославшему Его, Тот истинен, и нет неправды в Нем.
JOHN|7|19|Не дал ли вам Моисей закона? и никто из вас не поступает по закону. За что ищете убить Меня?
JOHN|7|20|Народ сказал в ответ: не бес ли в Тебе? кто ищет убить Тебя?
JOHN|7|21|Иисус, продолжая речь, сказал им: одно дело сделал Я, и все вы дивитесь.
JOHN|7|22|Моисей дал вам обрезание – хотя оно не от Моисея, но от отцов, – и в субботу вы обрезываете человека.
JOHN|7|23|Если в субботу принимает человек обрезание, чтобы не был нарушен закон Моисеев, – на Меня ли негодуете за то, что Я всего человека исцелил в субботу?
JOHN|7|24|Не судите по наружности, но судите судом праведным.
JOHN|7|25|Тут некоторые из Иерусалимлян говорили: не Тот ли это, Которого ищут убить?
JOHN|7|26|Вот, Он говорит явно, и ничего не говорят Ему: не удостоверились ли начальники, что Он подлинно Христос?
JOHN|7|27|Но мы знаем Его, откуда Он; Христос же когда придет, никто не будет знать, откуда Он.
JOHN|7|28|Тогда Иисус возгласил в храме, уча и говоря: и знаете Меня, и знаете, откуда Я; и Я пришел не Сам от Себя, но истинен Пославший Меня, Которого вы не знаете.
JOHN|7|29|Я знаю Его, потому что Я от Него, и Он послал Меня.
JOHN|7|30|И искали схватить Его, но никто не наложил на Него руки, потому что еще не пришел час Его.
JOHN|7|31|Многие же из народа уверовали в Него и говорили: когда придет Христос, неужели сотворит больше знамений, нежели сколько Сей сотворил?
JOHN|7|32|Услышали фарисеи такие толки о Нем в народе, и послали фарисеи и первосвященники служителей – схватить Его.
JOHN|7|33|Иисус же сказал им: еще недолго быть Мне с вами, и пойду к Пославшему Меня;
JOHN|7|34|будете искать Меня, и не найдете; и где буду Я, [туда] вы не можете придти.
JOHN|7|35|При сем Иудеи говорили между собою: куда Он хочет идти, так что мы не найдем Его? Не хочет ли Он идти в Еллинское рассеяние и учить Еллинов?
JOHN|7|36|Что значат сии слова, которые Он сказал: будете искать Меня, и не найдете; и где буду Я, [туда] вы не можете придти?
JOHN|7|37|В последний же великий день праздника стоял Иисус и возгласил, говоря: кто жаждет, иди ко Мне и пей.
JOHN|7|38|Кто верует в Меня, у того, как сказано в Писании, из чрева потекут реки воды живой.
JOHN|7|39|Сие сказал Он о Духе, Которого имели принять верующие в Него: ибо еще не было на них Духа Святаго, потому что Иисус еще не был прославлен.
JOHN|7|40|Многие из народа, услышав сии слова, говорили: Он точно пророк.
JOHN|7|41|Другие говорили: это Христос. А иные говорили: разве из Галилеи Христос придет?
JOHN|7|42|Не сказано ли в Писании, что Христос придет от семени Давидова и из Вифлеема, из того места, откуда был Давид?
JOHN|7|43|Итак произошла о Нем распря в народе.
JOHN|7|44|Некоторые из них хотели схватить Его; но никто не наложил на Него рук.
JOHN|7|45|Итак служители возвратились к первосвященникам и фарисеям, и сии сказали им: для чего вы не привели Его?
JOHN|7|46|Служители отвечали: никогда человек не говорил так, как Этот Человек.
JOHN|7|47|Фарисеи сказали им: неужели и вы прельстились?
JOHN|7|48|Уверовал ли в Него кто из начальников, или из фарисеев?
JOHN|7|49|Но этот народ невежда в законе, проклят он.
JOHN|7|50|Никодим, приходивший к Нему ночью, будучи один из них, говорит им:
JOHN|7|51|судит ли закон наш человека, если прежде не выслушают его и не узнают, что он делает?
JOHN|7|52|На это сказали ему: и ты не из Галилеи ли? рассмотри и увидишь, что из Галилеи не приходит пророк.
JOHN|7|53|И разошлись все по домам.
JOHN|8|1|Иисус же пошел на гору Елеонскую.
JOHN|8|2|А утром опять пришел в храм, и весь народ шел к Нему. Он сел и учил их.
JOHN|8|3|Тут книжники и фарисеи привели к Нему женщину, взятую в прелюбодеянии, и, поставив ее посреди,
JOHN|8|4|сказали Ему: Учитель! эта женщина взята в прелюбодеянии;
JOHN|8|5|а Моисей в законе заповедал нам побивать таких камнями: Ты что скажешь?
JOHN|8|6|Говорили же это, искушая Его, чтобы найти что–нибудь к обвинению Его. Но Иисус, наклонившись низко, писал перстом на земле, не обращая на них внимания.
JOHN|8|7|Когда же продолжали спрашивать Его, Он, восклонившись, сказал им: кто из вас без греха, первый брось на нее камень.
JOHN|8|8|И опять, наклонившись низко, писал на земле.
JOHN|8|9|Они же, услышав [то] и будучи обличаемы совестью, стали уходить один за другим, начиная от старших до последних; и остался один Иисус и женщина, стоящая посреди.
JOHN|8|10|Иисус, восклонившись и не видя никого, кроме женщины, сказал ей: женщина! где твои обвинители? никто не осудил тебя?
JOHN|8|11|Она отвечала: никто, Господи. Иисус сказал ей: и Я не осуждаю тебя; иди и впредь не греши.
JOHN|8|12|Опять говорил Иисус [к народу] и сказал им: Я свет миру; кто последует за Мною, тот не будет ходить во тьме, но будет иметь свет жизни.
JOHN|8|13|Тогда фарисеи сказали Ему: Ты Сам о Себе свидетельствуешь, свидетельство Твое не истинно.
JOHN|8|14|Иисус сказал им в ответ: если Я и Сам о Себе свидетельствую, свидетельство Мое истинно; потому что Я знаю, откуда пришел и куда иду; а вы не знаете, откуда Я и куда иду.
JOHN|8|15|Вы судите по плоти; Я не сужу никого.
JOHN|8|16|А если и сужу Я, то суд Мой истинен, потому что Я не один, но Я и Отец, пославший Меня.
JOHN|8|17|А и в законе вашем написано, что двух человек свидетельство истинно.
JOHN|8|18|Я Сам свидетельствую о Себе, и свидетельствует о Мне Отец, пославший Меня.
JOHN|8|19|Тогда сказали Ему: где Твой Отец? Иисус отвечал: вы не знаете ни Меня, ни Отца Моего; если бы вы знали Меня, то знали бы и Отца Моего.
JOHN|8|20|Сии слова говорил Иисус у сокровищницы, когда учил в храме; и никто не взял Его, потому что еще не пришел час Его.
JOHN|8|21|Опять сказал им Иисус: Я отхожу, и будете искать Меня, и умрете во грехе вашем. Куда Я иду, [туда] вы не можете придти.
JOHN|8|22|Тут Иудеи говорили: неужели Он убьет Сам Себя, что говорит: "куда Я иду, вы не можете придти"?
JOHN|8|23|Он сказал им: вы от нижних, Я от вышних; вы от мира сего, Я не от сего мира.
JOHN|8|24|Потому Я и сказал вам, что вы умрете во грехах ваших; ибо если не уверуете, что это Я, то умрете во грехах ваших.
JOHN|8|25|Тогда сказали Ему: кто же Ты? Иисус сказал им: от начала Сущий, как и говорю вам.
JOHN|8|26|Много имею говорить и судить о вас; но Пославший Меня есть истинен, и что Я слышал от Него, то и говорю миру.
JOHN|8|27|Не поняли, что Он говорил им об Отце.
JOHN|8|28|Итак Иисус сказал им: когда вознесете Сына Человеческого, тогда узнаете, что это Я и что ничего не делаю от Себя, но как научил Меня Отец Мой, так и говорю.
JOHN|8|29|Пославший Меня есть со Мною; Отец не оставил Меня одного, ибо Я всегда делаю то, что Ему угодно.
JOHN|8|30|Когда Он говорил это, многие уверовали в Него.
JOHN|8|31|Тогда сказал Иисус к уверовавшим в Него Иудеям: если пребудете в слове Моем, то вы истинно Мои ученики,
JOHN|8|32|и познаете истину, и истина сделает вас свободными.
JOHN|8|33|Ему отвечали: мы семя Авраамово и не были рабами никому никогда; как же Ты говоришь: сделаетесь свободными?
JOHN|8|34|Иисус отвечал им: истинно, истинно говорю вам: всякий, делающий грех, есть раб греха.
JOHN|8|35|Но раб не пребывает в доме вечно; сын пребывает вечно.
JOHN|8|36|Итак, если Сын освободит вас, то истинно свободны будете.
JOHN|8|37|Знаю, что вы семя Авраамово; однако ищете убить Меня, потому что слово Мое не вмещается в вас.
JOHN|8|38|Я говорю то, что видел у Отца Моего; а вы делаете то, что видели у отца вашего.
JOHN|8|39|Сказали Ему в ответ: отец наш есть Авраам. Иисус сказал им: если бы вы были дети Авраама, то дела Авраамовы делали бы.
JOHN|8|40|А теперь ищете убить Меня, Человека, сказавшего вам истину, которую слышал от Бога: Авраам этого не делал.
JOHN|8|41|Вы делаете дела отца вашего. На это сказали Ему: мы не от любодеяния рождены; одного Отца имеем, Бога.
JOHN|8|42|Иисус сказал им: если бы Бог был Отец ваш, то вы любили бы Меня, потому что Я от Бога исшел и пришел; ибо Я не Сам от Себя пришел, но Он послал Меня.
JOHN|8|43|Почему вы не понимаете речи Моей? Потому что не можете слышать слова Моего.
JOHN|8|44|Ваш отец диавол; и вы хотите исполнять похоти отца вашего. Он был человекоубийца от начала и не устоял в истине, ибо нет в нем истины. Когда говорит он ложь, говорит свое, ибо он лжец и отец лжи.
JOHN|8|45|А как Я истину говорю, то не верите Мне.
JOHN|8|46|Кто из вас обличит Меня в неправде? Если же Я говорю истину, почему вы не верите Мне?
JOHN|8|47|Кто от Бога, тот слушает слова Божии. Вы потому не слушаете, что вы не от Бога.
JOHN|8|48|На это Иудеи отвечали и сказали Ему: не правду ли мы говорим, что Ты Самарянин и что бес в Тебе?
JOHN|8|49|Иисус отвечал: во Мне беса нет; но Я чту Отца Моего, а вы бесчестите Меня.
JOHN|8|50|Впрочем Я не ищу Моей славы: есть Ищущий и Судящий.
JOHN|8|51|Истинно, истинно говорю вам: кто соблюдет слово Мое, тот не увидит смерти вовек.
JOHN|8|52|Иудеи сказали Ему: теперь узнали мы, что бес в Тебе. Авраам умер и пророки, а Ты говоришь: кто соблюдет слово Мое, тот не вкусит смерти вовек.
JOHN|8|53|Неужели Ты больше отца нашего Авраама, который умер? и пророки умерли: чем Ты Себя делаешь?
JOHN|8|54|Иисус отвечал: если Я Сам Себя славлю, то слава Моя ничто. Меня прославляет Отец Мой, о Котором вы говорите, что Он Бог ваш.
JOHN|8|55|И вы не познали Его, а Я знаю Его; и если скажу, что не знаю Его, то буду подобный вам лжец. Но Я знаю Его и соблюдаю слово Его.
JOHN|8|56|Авраам, отец ваш, рад был увидеть день Мой; и увидел и возрадовался.
JOHN|8|57|На это сказали Ему Иудеи: Тебе нет еще пятидесяти лет, – и Ты видел Авраама?
JOHN|8|58|Иисус сказал им: истинно, истинно говорю вам: прежде нежели был Авраам, Я есмь.
JOHN|8|59|Тогда взяли каменья, чтобы бросить на Него; но Иисус скрылся и вышел из храма, пройдя посреди них, и пошел далее.
JOHN|9|1|И, проходя, увидел человека, слепого от рождения.
JOHN|9|2|Ученики Его спросили у Него: Равви! кто согрешил, он или родители его, что родился слепым?
JOHN|9|3|Иисус отвечал: не согрешил ни он, ни родители его, но [это для] [того], чтобы на нем явились дела Божии.
JOHN|9|4|Мне должно делать дела Пославшего Меня, доколе есть день; приходит ночь, когда никто не может делать.
JOHN|9|5|Доколе Я в мире, Я свет миру.
JOHN|9|6|Сказав это, Он плюнул на землю, сделал брение из плюновения и помазал брением глаза слепому,
JOHN|9|7|и сказал ему: пойди, умойся в купальне Силоам, что значит: посланный. Он пошел и умылся, и пришел зрячим.
JOHN|9|8|Тут соседи и видевшие прежде, что он был слеп, говорили: не тот ли это, который сидел и просил милостыни?
JOHN|9|9|Иные говорили: это он, а иные: похож на него. Он же говорил: это я.
JOHN|9|10|Тогда спрашивали у него: как открылись у тебя глаза?
JOHN|9|11|Он сказал в ответ: Человек, называемый Иисус, сделал брение, помазал глаза мои и сказал мне: пойди на купальню Силоам и умойся. Я пошел, умылся и прозрел.
JOHN|9|12|Тогда сказали ему: где Он? Он отвечал: не знаю.
JOHN|9|13|Повели сего бывшего слепца к фарисеям.
JOHN|9|14|А была суббота, когда Иисус сделал брение и отверз ему очи.
JOHN|9|15|Спросили его также и фарисеи, как он прозрел. Он сказал им: брение положил Он на мои глаза, и я умылся, и вижу.
JOHN|9|16|Тогда некоторые из фарисеев говорили: не от Бога Этот Человек, потому что не хранит субботы. Другие говорили: как может человек грешный творить такие чудеса? И была между ними распря.
JOHN|9|17|Опять говорят слепому: ты что скажешь о Нем, потому что Он отверз тебе очи? Он сказал: это пророк.
JOHN|9|18|Тогда Иудеи не поверили, что он был слеп и прозрел, доколе не призвали родителей сего прозревшего
JOHN|9|19|и спросили их: это ли сын ваш, о котором вы говорите, что родился слепым? как же он теперь видит?
JOHN|9|20|Родители его сказали им в ответ: мы знаем, что это сын наш и что он родился слепым,
JOHN|9|21|а как теперь видит, не знаем, или кто отверз ему очи, мы не знаем. Сам в совершенных летах; самого спросите; пусть сам о себе скажет.
JOHN|9|22|Так отвечали родители его, потому что боялись Иудеев; ибо Иудеи сговорились уже, чтобы, кто признает Его за Христа, того отлучать от синагоги.
JOHN|9|23|Посему–то родители его и сказали: он в совершенных летах; самого спросите.
JOHN|9|24|Итак, вторично призвали человека, который был слеп, и сказали ему: воздай славу Богу; мы знаем, что Человек Тот грешник.
JOHN|9|25|Он сказал им в ответ: грешник ли Он, не знаю; одно знаю, что я был слеп, а теперь вижу.
JOHN|9|26|Снова спросили его: что сделал Он с тобою? как отверз твои очи?
JOHN|9|27|Отвечал им: я уже сказал вам, и вы не слушали; что еще хотите слышать? или и вы хотите сделаться Его учениками?
JOHN|9|28|Они же укорили его и сказали: ты ученик Его, а мы Моисеевы ученики.
JOHN|9|29|Мы знаем, что с Моисеем говорил Бог; Сего же не знаем, откуда Он.
JOHN|9|30|Человек [прозревший] сказал им в ответ: это и удивительно, что вы не знаете, откуда Он, а Он отверз мне очи.
JOHN|9|31|Но мы знаем, что грешников Бог не слушает; но кто чтит Бога и творит волю Его, того слушает.
JOHN|9|32|От века не слыхано, чтобы кто отверз очи слепорожденному.
JOHN|9|33|Если бы Он не был от Бога, не мог бы творить ничего.
JOHN|9|34|Сказали ему в ответ: во грехах ты весь родился, и ты ли нас учишь? И выгнали его вон.
JOHN|9|35|Иисус, услышав, что выгнали его вон, и найдя его, сказал ему: ты веруешь ли в Сына Божия?
JOHN|9|36|Он отвечал и сказал: а кто Он, Господи, чтобы мне веровать в Него?
JOHN|9|37|Иисус сказал ему: и видел ты Его, и Он говорит с тобою.
JOHN|9|38|Он же сказал: верую, Господи! И поклонился Ему.
JOHN|9|39|И сказал Иисус: на суд пришел Я в мир сей, чтобы невидящие видели, а видящие стали слепы.
JOHN|9|40|Услышав это, некоторые из фарисеев, бывших с Ним, сказали Ему: неужели и мы слепы?
JOHN|9|41|Иисус сказал им: если бы вы были слепы, то не имели бы [на] [себе] греха; но как вы говорите, что видите, то грех остается на вас.
JOHN|10|1|Истинно, истинно говорю вам: кто не дверью входит во двор овчий, но перелазит инде, тот вор и разбойник;
JOHN|10|2|а входящий дверью есть пастырь овцам.
JOHN|10|3|Ему придверник отворяет, и овцы слушаются голоса его, и он зовет своих овец по имени и выводит их.
JOHN|10|4|И когда выведет своих овец, идет перед ними; а овцы за ним идут, потому что знают голос его.
JOHN|10|5|За чужим же не идут, но бегут от него, потому что не знают чужого голоса.
JOHN|10|6|Сию притчу сказал им Иисус; но они не поняли, что такое Он говорил им.
JOHN|10|7|Итак, опять Иисус сказал им: истинно, истинно говорю вам, что Я дверь овцам.
JOHN|10|8|Все, сколько их ни приходило предо Мною, суть воры и разбойники; но овцы не послушали их.
JOHN|10|9|Я есмь дверь: кто войдет Мною, тот спасется, и войдет, и выйдет, и пажить найдет.
JOHN|10|10|Вор приходит только для того, чтобы украсть, убить и погубить. Я пришел для того, чтобы имели жизнь и имели с избытком.
JOHN|10|11|Я есмь пастырь добрый: пастырь добрый полагает жизнь свою за овец.
JOHN|10|12|А наемник, не пастырь, которому овцы не свои, видит приходящего волка, и оставляет овец, и бежит; и волк расхищает овец, и разгоняет их.
JOHN|10|13|А наемник бежит, потому что наемник, и нерадит об овцах.
JOHN|10|14|Я есмь пастырь добрый; и знаю Моих, и Мои знают Меня.
JOHN|10|15|Как Отец знает Меня, [так] и Я знаю Отца; и жизнь Мою полагаю за овец.
JOHN|10|16|Есть у Меня и другие овцы, которые не сего двора, и тех надлежит Мне привести: и они услышат голос Мой, и будет одно стадо и один Пастырь.
JOHN|10|17|Потому любит Меня Отец, что Я отдаю жизнь Мою, чтобы опять принять ее.
JOHN|10|18|Никто не отнимает ее у Меня, но Я Сам отдаю ее. Имею власть отдать ее и власть имею опять принять ее. Сию заповедь получил Я от Отца Моего.
JOHN|10|19|От этих слов опять произошла между Иудеями распря.
JOHN|10|20|Многие из них говорили: Он одержим бесом и безумствует; что слушаете Его?
JOHN|10|21|Другие говорили: это слова не бесноватого; может ли бес отверзать очи слепым?
JOHN|10|22|Настал же тогда в Иерусалиме [праздник] обновления, и была зима.
JOHN|10|23|И ходил Иисус в храме, в притворе Соломоновом.
JOHN|10|24|Тут Иудеи обступили Его и говорили Ему: долго ли Тебе держать нас в недоумении? если Ты Христос, скажи нам прямо.
JOHN|10|25|Иисус отвечал им: Я сказал вам, и не верите; дела, которые творю Я во имя Отца Моего, они свидетельствуют о Мне.
JOHN|10|26|Но вы не верите, ибо вы не из овец Моих, как Я сказал вам.
JOHN|10|27|Овцы Мои слушаются голоса Моего, и Я знаю их; и они идут за Мною.
JOHN|10|28|И Я даю им жизнь вечную, и не погибнут вовек; и никто не похитит их из руки Моей.
JOHN|10|29|Отец Мой, Который дал Мне их, больше всех; и никто не может похитить их из руки Отца Моего.
JOHN|10|30|Я и Отец – одно.
JOHN|10|31|Тут опять Иудеи схватили каменья, чтобы побить Его.
JOHN|10|32|Иисус отвечал им: много добрых дел показал Я вам от Отца Моего; за которое из них хотите побить Меня камнями?
JOHN|10|33|Иудеи сказали Ему в ответ: не за доброе дело хотим побить Тебя камнями, но за богохульство и за то, что Ты, будучи человек, делаешь Себя Богом.
JOHN|10|34|Иисус отвечал им: не написано ли в законе вашем: Я сказал: вы боги?
JOHN|10|35|Если Он назвал богами тех, к которым было слово Божие, и не может нарушиться Писание, –
JOHN|10|36|Тому ли, Которого Отец освятил и послал в мир, вы говорите: богохульствуешь, потому что Я сказал: Я Сын Божий?
JOHN|10|37|Если Я не творю дел Отца Моего, не верьте Мне;
JOHN|10|38|а если творю, то, когда не верите Мне, верьте делам Моим, чтобы узнать и поверить, что Отец во Мне и Я в Нем.
JOHN|10|39|Тогда опять искали схватить Его; но Он уклонился от рук их,
JOHN|10|40|и пошел опять за Иордан, на то место, где прежде крестил Иоанн, и остался там.
JOHN|10|41|Многие пришли к Нему и говорили, что Иоанн не сотворил никакого чуда, но все, что сказал Иоанн о Нем, было истинно.
JOHN|10|42|И многие там уверовали в Него.
JOHN|11|1|Был болен некто Лазарь из Вифании, из селения, [где жили] Мария и Марфа, сестра ее.
JOHN|11|2|Мария же, которой брат Лазарь был болен, была [та], которая помазала Господа миром и отерла ноги Его волосами своими.
JOHN|11|3|Сестры послали сказать Ему: Господи! вот, кого Ты любишь, болен.
JOHN|11|4|Иисус, услышав [то], сказал: эта болезнь не к смерти, но к славе Божией, да прославится через нее Сын Божий.
JOHN|11|5|Иисус же любил Марфу и сестру ее и Лазаря.
JOHN|11|6|Когда же услышал, что он болен, то пробыл два дня на том месте, где находился.
JOHN|11|7|После этого сказал ученикам: пойдем опять в Иудею.
JOHN|11|8|Ученики сказали Ему: Равви! давно ли Иудеи искали побить Тебя камнями, и Ты опять идешь туда?
JOHN|11|9|Иисус отвечал: не двенадцать ли часов во дне? кто ходит днем, тот не спотыкается, потому что видит свет мира сего;
JOHN|11|10|а кто ходит ночью, спотыкается, потому что нет света с ним.
JOHN|11|11|Сказав это, говорит им потом: Лазарь, друг наш, уснул; но Я иду разбудить его.
JOHN|11|12|Ученики Его сказали: Господи! если уснул, то выздоровеет.
JOHN|11|13|Иисус говорил о смерти его, а они думали, что Он говорит о сне обыкновенном.
JOHN|11|14|Тогда Иисус сказал им прямо: Лазарь умер;
JOHN|11|15|и радуюсь за вас, что Меня не было там, дабы вы уверовали; но пойдем к нему.
JOHN|11|16|Тогда Фома, иначе называемый Близнец, сказал ученикам: пойдем и мы умрем с ним.
JOHN|11|17|Иисус, придя, нашел, что он уже четыре дня в гробе.
JOHN|11|18|Вифания же была близ Иерусалима, стадиях в пятнадцати;
JOHN|11|19|и многие из Иудеев пришли к Марфе и Марии утешать их [в] [печали] о брате их.
JOHN|11|20|Марфа, услышав, что идет Иисус, пошла навстречу Ему; Мария же сидела дома.
JOHN|11|21|Тогда Марфа сказала Иисусу: Господи! если бы Ты был здесь, не умер бы брат мой.
JOHN|11|22|Но и теперь знаю, что чего Ты попросишь у Бога, даст Тебе Бог.
JOHN|11|23|Иисус говорит ей: воскреснет брат твой.
JOHN|11|24|Марфа сказала Ему: знаю, что воскреснет в воскресение, в последний день.
JOHN|11|25|Иисус сказал ей: Я есмь воскресение и жизнь; верующий в Меня, если и умрет, оживет.
JOHN|11|26|И всякий, живущий и верующий в Меня, не умрет вовек. Веришь ли сему?
JOHN|11|27|Она говорит Ему: так, Господи! я верую, что Ты Христос, Сын Божий, грядущий в мир.
JOHN|11|28|Сказав это, пошла и позвала тайно Марию, сестру свою, говоря: Учитель здесь и зовет тебя.
JOHN|11|29|Она, как скоро услышала, поспешно встала и пошла к Нему.
JOHN|11|30|Иисус еще не входил в селение, но был на том месте, где встретила Его Марфа.
JOHN|11|31|Иудеи, которые были с нею в доме и утешали ее, видя, что Мария поспешно встала и вышла, пошли за нею, полагая, что она пошла на гроб – плакать там.
JOHN|11|32|Мария же, придя туда, где был Иисус, и увидев Его, пала к ногам Его и сказала Ему: Господи! если бы Ты был здесь, не умер бы брат мой.
JOHN|11|33|Иисус, когда увидел ее плачущую и пришедших с нею Иудеев плачущих, Сам восскорбел духом и возмутился
JOHN|11|34|и сказал: где вы положили его? Говорят Ему: Господи! пойди и посмотри.
JOHN|11|35|Иисус прослезился.
JOHN|11|36|Тогда Иудеи говорили: смотри, как Он любил его.
JOHN|11|37|А некоторые из них сказали: не мог ли Сей, отверзший очи слепому, сделать, чтобы и этот не умер?
JOHN|11|38|Иисус же, опять скорбя внутренно, приходит ко гробу. То была пещера, и камень лежал на ней.
JOHN|11|39|Иисус говорит: отнимите камень. Сестра умершего, Марфа, говорит Ему: Господи! уже смердит; ибо четыре дня, как он во гробе.
JOHN|11|40|Иисус говорит ей: не сказал ли Я тебе, что, если будешь веровать, увидишь славу Божию?
JOHN|11|41|Итак отняли камень [от пещеры], где лежал умерший. Иисус же возвел очи к небу и сказал: Отче! благодарю Тебя, что Ты услышал Меня.
JOHN|11|42|Я и знал, что Ты всегда услышишь Меня; но сказал [сие] для народа, здесь стоящего, чтобы поверили, что Ты послал Меня.
JOHN|11|43|Сказав это, Он воззвал громким голосом: Лазарь! иди вон.
JOHN|11|44|И вышел умерший, обвитый по рукам и ногам погребальными пеленами, и лице его обвязано было платком. Иисус говорит им: развяжите его, пусть идет.
JOHN|11|45|Тогда многие из Иудеев, пришедших к Марии и видевших, что сотворил Иисус, уверовали в Него.
JOHN|11|46|А некоторые из них пошли к фарисеям и сказали им, что сделал Иисус.
JOHN|11|47|Тогда первосвященники и фарисеи собрали совет и говорили: что нам делать? Этот Человек много чудес творит.
JOHN|11|48|Если оставим Его так, то все уверуют в Него, и придут Римляне и овладеют и местом нашим и народом.
JOHN|11|49|Один же из них, некто Каиафа, будучи на тот год первосвященником, сказал им: вы ничего не знаете,
JOHN|11|50|и не подумаете, что лучше нам, чтобы один человек умер за людей, нежели чтобы весь народ погиб.
JOHN|11|51|Сие же он сказал не от себя, но, будучи на тот год первосвященником, предсказал, что Иисус умрет за народ,
JOHN|11|52|и не только за народ, но чтобы и рассеянных чад Божиих собрать воедино.
JOHN|11|53|С этого дня положили убить Его.
JOHN|11|54|Посему Иисус уже не ходил явно между Иудеями, а пошел оттуда в страну близ пустыни, в город, называемый Ефраим, и там оставался с учениками Своими.
JOHN|11|55|Приближалась Пасха Иудейская, и многие из всей страны пришли в Иерусалим перед Пасхою, чтобы очиститься.
JOHN|11|56|Тогда искали Иисуса и, стоя в храме, говорили друг другу: как вы думаете? не придет ли Он на праздник?
JOHN|11|57|Первосвященники же и фарисеи дали приказание, что если кто узнает, где Он будет, то объявил бы, дабы взять Его.
JOHN|12|1|За шесть дней до Пасхи пришел Иисус в Вифанию, где был Лазарь умерший, которого Он воскресил из мертвых.
JOHN|12|2|Там приготовили Ему вечерю, и Марфа служила, и Лазарь был одним из возлежавших с Ним.
JOHN|12|3|Мария же, взяв фунт нардового чистого драгоценного мира, помазала ноги Иисуса и отерла волосами своими ноги Его; и дом наполнился благоуханием от мира.
JOHN|12|4|Тогда один из учеников Его, Иуда Симонов Искариот, который хотел предать Его, сказал:
JOHN|12|5|Для чего бы не продать это миро за триста динариев и не раздать нищим?
JOHN|12|6|Сказал же он это не потому, чтобы заботился о нищих, но потому что был вор. Он имел [при себе денежный] ящик и носил, что туда опускали.
JOHN|12|7|Иисус же сказал: оставьте ее; она сберегла это на день погребения Моего.
JOHN|12|8|Ибо нищих всегда имеете с собою, а Меня не всегда.
JOHN|12|9|Многие из Иудеев узнали, что Он там, и пришли не только для Иисуса, но чтобы видеть и Лазаря, которого Он воскресил из мертвых.
JOHN|12|10|Первосвященники же положили убить и Лазаря,
JOHN|12|11|потому что ради него многие из Иудеев приходили и веровали в Иисуса.
JOHN|12|12|На другой день множество народа, пришедшего на праздник, услышав, что Иисус идет в Иерусалим,
JOHN|12|13|взяли пальмовые ветви, вышли навстречу Ему и восклицали: осанна! благословен грядущий во имя Господне, Царь Израилев!
JOHN|12|14|Иисус же, найдя молодого осла, сел на него, как написано:
JOHN|12|15|Не бойся, дщерь Сионова! се, Царь твой грядет, сидя на молодом осле.
JOHN|12|16|Ученики Его сперва не поняли этого; но когда прославился Иисус, тогда вспомнили, что так было о Нем написано, и это сделали Ему.
JOHN|12|17|Народ, бывший с Ним прежде, свидетельствовал, что Он вызвал из гроба Лазаря и воскресил его из мертвых.
JOHN|12|18|Потому и встретил Его народ, ибо слышал, что Он сотворил это чудо.
JOHN|12|19|Фарисеи же говорили между собою: видите ли, что не успеваете ничего? весь мир идет за Ним.
JOHN|12|20|Из пришедших на поклонение в праздник были некоторые Еллины.
JOHN|12|21|Они подошли к Филиппу, который был из Вифсаиды Галилейской, и просили его, говоря: господин! нам хочется видеть Иисуса.
JOHN|12|22|Филипп идет и говорит о том Андрею; и потом Андрей и Филипп сказывают о том Иисусу.
JOHN|12|23|Иисус же сказал им в ответ: пришел час прославиться Сыну Человеческому.
JOHN|12|24|Истинно, истинно говорю вам: если пшеничное зерно, пав в землю, не умрет, то останется одно; а если умрет, то принесет много плода.
JOHN|12|25|Любящий душу свою погубит ее; а ненавидящий душу свою в мире сем сохранит ее в жизнь вечную.
JOHN|12|26|Кто Мне служит, Мне да последует; и где Я, там и слуга Мой будет. И кто Мне служит, того почтит Отец Мой.
JOHN|12|27|Душа Моя теперь возмутилась; и что Мне сказать? Отче! избавь Меня от часа сего! Но на сей час Я и пришел.
JOHN|12|28|Отче! прославь имя Твое. Тогда пришел с неба глас: и прославил и еще прославлю.
JOHN|12|29|Народ, стоявший и слышавший [то], говорил: это гром; а другие говорили: Ангел говорил Ему.
JOHN|12|30|Иисус на это сказал: не для Меня был глас сей, но для народа.
JOHN|12|31|Ныне суд миру сему; ныне князь мира сего изгнан будет вон.
JOHN|12|32|И когда Я вознесен буду от земли, всех привлеку к Себе.
JOHN|12|33|Сие говорил Он, давая разуметь, какою смертью Он умрет.
JOHN|12|34|Народ отвечал Ему: мы слышали из закона, что Христос пребывает вовек; как же Ты говоришь, что должно вознесену быть Сыну Человеческому? кто Этот Сын Человеческий?
JOHN|12|35|Тогда Иисус сказал им: еще на малое время свет есть с вами; ходите, пока есть свет, чтобы не объяла вас тьма: а ходящий во тьме не знает, куда идет.
JOHN|12|36|Доколе свет с вами, веруйте в свет, да будете сынами света. Сказав это, Иисус отошел и скрылся от них.
JOHN|12|37|Столько чудес сотворил Он пред ними, и они не веровали в Него,
JOHN|12|38|да сбудется слово Исаии пророка: Господи! кто поверил слышанному от нас? и кому открылась мышца Господня?
JOHN|12|39|Потому не могли они веровать, что, как еще сказал Исаия,
JOHN|12|40|народ сей ослепил глаза свои и окаменил сердце свое, да не видят глазами, и не уразумеют сердцем, и не обратятся, чтобы Я исцелил их.
JOHN|12|41|Сие сказал Исаия, когда видел славу Его и говорил о Нем.
JOHN|12|42|Впрочем и из начальников многие уверовали в Него; но ради фарисеев не исповедывали, чтобы не быть отлученными от синагоги,
JOHN|12|43|ибо возлюбили больше славу человеческую, нежели славу Божию.
JOHN|12|44|Иисус же возгласил и сказал: верующий в Меня не в Меня верует, но в Пославшего Меня.
JOHN|12|45|И видящий Меня видит Пославшего Меня.
JOHN|12|46|Я свет пришел в мир, чтобы всякий верующий в Меня не оставался во тьме.
JOHN|12|47|И если кто услышит Мои слова и не поверит, Я не сужу его, ибо Я пришел не судить мир, но спасти мир.
JOHN|12|48|Отвергающий Меня и не принимающий слов Моих имеет судью себе: слово, которое Я говорил, оно будет судить его в последний день.
JOHN|12|49|Ибо Я говорил не от Себя; но пославший Меня Отец, Он дал Мне заповедь, что сказать и что говорить.
JOHN|12|50|И Я знаю, что заповедь Его есть жизнь вечная. Итак, что Я говорю, говорю, как сказал Мне Отец.
JOHN|13|1|Перед праздником Пасхи Иисус, зная, что пришел час Его перейти от мира сего к Отцу, [явил делом, что], возлюбив Своих сущих в мире, до конца возлюбил их.
JOHN|13|2|И во время вечери, когда диавол уже вложил в сердце Иуде Симонову Искариоту предать Его,
JOHN|13|3|Иисус, зная, что Отец все отдал в руки Его, и что Он от Бога исшел и к Богу отходит,
JOHN|13|4|встал с вечери, снял [с Себя верхнюю] одежду и, взяв полотенце, препоясался.
JOHN|13|5|Потом влил воды в умывальницу и начал умывать ноги ученикам и отирать полотенцем, которым был препоясан.
JOHN|13|6|Подходит к Симону Петру, и тот говорит Ему: Господи! Тебе ли умывать мои ноги?
JOHN|13|7|Иисус сказал ему в ответ: что Я делаю, теперь ты не знаешь, а уразумеешь после.
JOHN|13|8|Петр говорит Ему: не умоешь ног моих вовек. Иисус отвечал ему: если не умою тебя, не имеешь части со Мною.
JOHN|13|9|Симон Петр говорит Ему: Господи! не только ноги мои, но и руки и голову.
JOHN|13|10|Иисус говорит ему: омытому нужно только ноги умыть, потому что чист весь; и вы чисты, но не все.
JOHN|13|11|Ибо знал Он предателя Своего, потому [и] сказал: не все вы чисты.
JOHN|13|12|Когда же умыл им ноги и надел одежду Свою, то, возлегши опять, сказал им: знаете ли, что Я сделал вам?
JOHN|13|13|Вы называете Меня Учителем и Господом, и правильно говорите, ибо Я точно то.
JOHN|13|14|Итак, если Я, Господь и Учитель, умыл ноги вам, то и вы должны умывать ноги друг другу.
JOHN|13|15|Ибо Я дал вам пример, чтобы и вы делали то же, что Я сделал вам.
JOHN|13|16|Истинно, истинно говорю вам: раб не больше господина своего, и посланник не больше пославшего его.
JOHN|13|17|Если это знаете, блаженны вы, когда исполняете.
JOHN|13|18|Не о всех вас говорю; Я знаю, которых избрал. Но да сбудется Писание: ядущий со Мною хлеб поднял на Меня пяту свою.
JOHN|13|19|Теперь сказываю вам, прежде нежели [то] сбылось, дабы, когда сбудется, вы поверили, что это Я.
JOHN|13|20|Истинно, истинно говорю вам: принимающий того, кого Я пошлю, Меня принимает; а принимающий Меня принимает Пославшего Меня.
JOHN|13|21|Сказав это, Иисус возмутился духом, и засвидетельствовал, и сказал: истинно, истинно говорю вам, что один из вас предаст Меня.
JOHN|13|22|Тогда ученики озирались друг на друга, недоумевая, о ком Он говорит.
JOHN|13|23|Один же из учеников Его, которого любил Иисус, возлежал у груди Иисуса.
JOHN|13|24|Ему Симон Петр сделал знак, чтобы спросил, кто это, о котором говорит.
JOHN|13|25|Он, припав к груди Иисуса, сказал Ему: Господи! кто это?
JOHN|13|26|Иисус отвечал: тот, кому Я, обмакнув кусок хлеба, подам. И, обмакнув кусок, подал Иуде Симонову Искариоту.
JOHN|13|27|И после сего куска вошел в него сатана. Тогда Иисус сказал ему: что делаешь, делай скорее.
JOHN|13|28|Но никто из возлежавших не понял, к чему Он это сказал ему.
JOHN|13|29|А как у Иуды был ящик, то некоторые думали, что Иисус говорит ему: купи, что нам нужно к празднику, или чтобы дал что–нибудь нищим.
JOHN|13|30|Он, приняв кусок, тотчас вышел; а была ночь.
JOHN|13|31|Когда он вышел, Иисус сказал: ныне прославился Сын Человеческий, и Бог прославился в Нем.
JOHN|13|32|Если Бог прославился в Нем, то и Бог прославит Его в Себе, и вскоре прославит Его.
JOHN|13|33|Дети! недолго уже быть Мне с вами. Будете искать Меня, и, как сказал Я Иудеям, что, куда Я иду, вы не можете придти, [так] и вам говорю теперь.
JOHN|13|34|Заповедь новую даю вам, да любите друг друга; как Я возлюбил вас, [так] и вы да любите друг друга.
JOHN|13|35|По тому узнают все, что вы Мои ученики, если будете иметь любовь между собою.
JOHN|13|36|Симон Петр сказал Ему: Господи! куда Ты идешь? Иисус отвечал ему: куда Я иду, ты не можешь теперь за Мною идти, а после пойдешь за Мною.
JOHN|13|37|Петр сказал Ему: Господи! почему я не могу идти за Тобою теперь? я душу мою положу за Тебя.
JOHN|13|38|Иисус отвечал ему: душу твою за Меня положишь? истинно, истинно говорю тебе: не пропоет петух, как отречешься от Меня трижды.
JOHN|14|1|Да не смущается сердце ваше; веруйте в Бога, и в Меня веруйте.
JOHN|14|2|В доме Отца Моего обителей много. А если бы не так, Я сказал бы вам: Я иду приготовить место вам.
JOHN|14|3|И когда пойду и приготовлю вам место, приду опять и возьму вас к Себе, чтобы и вы были, где Я.
JOHN|14|4|А куда Я иду, вы знаете, и путь знаете.
JOHN|14|5|Фома сказал Ему: Господи! не знаем, куда идешь; и как можем знать путь?
JOHN|14|6|Иисус сказал ему: Я есмь путь и истина и жизнь; никто не приходит к Отцу, как только через Меня.
JOHN|14|7|Если бы вы знали Меня, то знали бы и Отца Моего. И отныне знаете Его и видели Его.
JOHN|14|8|Филипп сказал Ему: Господи! покажи нам Отца, и довольно для нас.
JOHN|14|9|Иисус сказал ему: столько времени Я с вами, и ты не знаешь Меня, Филипп? Видевший Меня видел Отца; как же ты говоришь, покажи нам Отца?
JOHN|14|10|Разве ты не веришь, что Я в Отце и Отец во Мне? Слова, которые говорю Я вам, говорю не от Себя; Отец, пребывающий во Мне, Он творит дела.
JOHN|14|11|Верьте Мне, что Я в Отце и Отец во Мне; а если не так, то верьте Мне по самым делам.
JOHN|14|12|Истинно, истинно говорю вам: верующий в Меня, дела, которые творю Я, и он сотворит, и больше сих сотворит, потому что Я к Отцу Моему иду.
JOHN|14|13|И если чего попросите у Отца во имя Мое, то сделаю, да прославится Отец в Сыне.
JOHN|14|14|Если чего попросите во имя Мое, Я то сделаю.
JOHN|14|15|Если любите Меня, соблюдите Мои заповеди.
JOHN|14|16|И Я умолю Отца, и даст вам другого Утешителя, да пребудет с вами вовек,
JOHN|14|17|Духа истины, Которого мир не может принять, потому что не видит Его и не знает Его; а вы знаете Его, ибо Он с вами пребывает и в вас будет.
JOHN|14|18|Не оставлю вас сиротами; приду к вам.
JOHN|14|19|Еще немного, и мир уже не увидит Меня; а вы увидите Меня, ибо Я живу, и вы будете жить.
JOHN|14|20|В тот день узнаете вы, что Я в Отце Моем, и вы во Мне, и Я в вас.
JOHN|14|21|Кто имеет заповеди Мои и соблюдает их, тот любит Меня; а кто любит Меня, тот возлюблен будет Отцем Моим; и Я возлюблю его и явлюсь ему Сам.
JOHN|14|22|Иуда – не Искариот – говорит Ему: Господи! что это, что Ты хочешь явить Себя нам, а не миру?
JOHN|14|23|Иисус сказал ему в ответ: кто любит Меня, тот соблюдет слово Мое; и Отец Мой возлюбит его, и Мы придем к нему и обитель у него сотворим.
JOHN|14|24|Нелюбящий Меня не соблюдает слов Моих; слово же, которое вы слышите, не есть Мое, но пославшего Меня Отца.
JOHN|14|25|Сие сказал Я вам, находясь с вами.
JOHN|14|26|Утешитель же, Дух Святый, Которого пошлет Отец во имя Мое, научит вас всему и напомнит вам все, что Я говорил вам.
JOHN|14|27|Мир оставляю вам, мир Мой даю вам; не так, как мир дает, Я даю вам. Да не смущается сердце ваше и да не устрашается.
JOHN|14|28|Вы слышали, что Я сказал вам: иду от вас и приду к вам. Если бы вы любили Меня, то возрадовались бы, что Я сказал: иду к Отцу; ибо Отец Мой более Меня.
JOHN|14|29|И вот, Я сказал вам [о том], прежде нежели сбылось, дабы вы поверили, когда сбудется.
JOHN|14|30|Уже немного Мне говорить с вами; ибо идет князь мира сего, и во Мне не имеет ничего.
JOHN|14|31|Но чтобы мир знал, что Я люблю Отца и, как заповедал Мне Отец, так и творю: встаньте, пойдем отсюда.
JOHN|15|1|Я есмь истинная виноградная лоза, а Отец Мой – виноградарь.
JOHN|15|2|Всякую у Меня ветвь, не приносящую плода, Он отсекает; и всякую, приносящую плод, очищает, чтобы более принесла плода.
JOHN|15|3|Вы уже очищены через слово, которое Я проповедал вам.
JOHN|15|4|Пребудьте во Мне, и Я в вас. Как ветвь не может приносить плода сама собою, если не будет на лозе: так и вы, если не будете во Мне.
JOHN|15|5|Я есмь лоза, а вы ветви; кто пребывает во Мне, и Я в нем, тот приносит много плода; ибо без Меня не можете делать ничего.
JOHN|15|6|Кто не пребудет во Мне, извергнется вон, как ветвь, и засохнет; а такие [ветви] собирают и бросают в огонь, и они сгорают.
JOHN|15|7|Если пребудете во Мне и слова Мои в вас пребудут, то, чего ни пожелаете, просите, и будет вам.
JOHN|15|8|Тем прославится Отец Мой, если вы принесете много плода и будете Моими учениками.
JOHN|15|9|Как возлюбил Меня Отец, и Я возлюбил вас; пребудьте в любви Моей.
JOHN|15|10|Если заповеди Мои соблюдете, пребудете в любви Моей, как и Я соблюл заповеди Отца Моего и пребываю в Его любви.
JOHN|15|11|Сие сказал Я вам, да радость Моя в вас пребудет и радость ваша будет совершенна.
JOHN|15|12|Сия есть заповедь Моя, да любите друг друга, как Я возлюбил вас.
JOHN|15|13|Нет больше той любви, как если кто положит душу свою за друзей своих.
JOHN|15|14|Вы друзья Мои, если исполняете то, что Я заповедую вам.
JOHN|15|15|Я уже не называю вас рабами, ибо раб не знает, что делает господин его; но Я назвал вас друзьями, потому что сказал вам все, что слышал от Отца Моего.
JOHN|15|16|Не вы Меня избрали, а Я вас избрал и поставил вас, чтобы вы шли и приносили плод, и чтобы плод ваш пребывал, дабы, чего ни попросите от Отца во имя Мое, Он дал вам.
JOHN|15|17|Сие заповедаю вам, да любите друг друга.
JOHN|15|18|Если мир вас ненавидит, знайте, что Меня прежде вас возненавидел.
JOHN|15|19|Если бы вы были от мира, то мир любил бы свое; а как вы не от мира, но Я избрал вас от мира, потому ненавидит вас мир.
JOHN|15|20|Помните слово, которое Я сказал вам: раб не больше господина своего. Если Меня гнали, будут гнать и вас; если Мое слово соблюдали, будут соблюдать и ваше.
JOHN|15|21|Но все то сделают вам за имя Мое, потому что не знают Пославшего Меня.
JOHN|15|22|Если бы Я не пришел и не говорил им, то не имели бы греха; а теперь не имеют извинения во грехе своем.
JOHN|15|23|Ненавидящий Меня ненавидит и Отца моего.
JOHN|15|24|Если бы Я не сотворил между ними дел, каких никто другой не делал, то не имели бы греха; а теперь и видели, и возненавидели и Меня и Отца Моего.
JOHN|15|25|Но да сбудется слово, написанное в законе их: возненавидели Меня напрасно.
JOHN|15|26|Когда же приидет Утешитель, Которого Я пошлю вам от Отца, Дух истины, Который от Отца исходит, Он будет свидетельствовать о Мне;
JOHN|15|27|а также и вы будете свидетельствовать, потому что вы сначала со Мною.
JOHN|16|1|Сие сказал Я вам, чтобы вы не соблазнились.
JOHN|16|2|Изгонят вас из синагог; даже наступает время, когда всякий, убивающий вас, будет думать, что он тем служит Богу.
JOHN|16|3|Так будут поступать, потому что не познали ни Отца, ни Меня.
JOHN|16|4|Но Я сказал вам сие для того, чтобы вы, когда придет то время вспомнили, что Я сказывал вам о том; не говорил же сего вам сначала, потому что был с вами.
JOHN|16|5|А теперь иду к Пославшему Меня, и никто из вас не спрашивает Меня: куда идешь?
JOHN|16|6|Но от того, что Я сказал вам это, печалью исполнилось сердце ваше.
JOHN|16|7|Но Я истину говорю вам: лучше для вас, чтобы Я пошел; ибо, если Я не пойду, Утешитель не приидет к вам; а если пойду, то пошлю Его к вам,
JOHN|16|8|и Он, придя, обличит мир о грехе и о правде и о суде:
JOHN|16|9|о грехе, что не веруют в Меня;
JOHN|16|10|о правде, что Я иду к Отцу Моему, и уже не увидите Меня;
JOHN|16|11|о суде же, что князь мира сего осужден.
JOHN|16|12|Еще многое имею сказать вам; но вы теперь не можете вместить.
JOHN|16|13|Когда же приидет Он, Дух истины, то наставит вас на всякую истину: ибо не от Себя говорить будет, но будет говорить, что услышит, и будущее возвестит вам.
JOHN|16|14|Он прославит Меня, потому что от Моего возьмет и возвестит вам.
JOHN|16|15|Все, что имеет Отец, есть Мое; потому Я сказал, что от Моего возьмет и возвестит вам.
JOHN|16|16|Вскоре вы не увидите Меня, и опять вскоре увидите Меня, ибо Я иду к Отцу.
JOHN|16|17|Тут [некоторые] из учеников Его сказали один другому: что это Он говорит нам: вскоре не увидите Меня, и опять вскоре увидите Меня, и: Я иду к Отцу?
JOHN|16|18|Итак они говорили: что это говорит Он: "вскоре"? Не знаем, что говорит.
JOHN|16|19|Иисус, уразумев, что хотят спросить Его, сказал им: о том ли спрашиваете вы один другого, что Я сказал: вскоре не увидите Меня, и опять вскоре увидите Меня?
JOHN|16|20|Истинно, истинно говорю вам: вы восплачете и возрыдаете, а мир возрадуется; вы печальны будете, но печаль ваша в радость будет.
JOHN|16|21|Женщина, когда рождает, терпит скорбь, потому что пришел час ее; но когда родит младенца, уже не помнит скорби от радости, потому что родился человек в мир.
JOHN|16|22|Так и вы теперь имеете печаль; но Я увижу вас опять, и возрадуется сердце ваше, и радости вашей никто не отнимет у вас;
JOHN|16|23|и в тот день вы не спросите Меня ни о чем. Истинно, истинно говорю вам: о чем ни попросите Отца во имя Мое, даст вам.
JOHN|16|24|Доныне вы ничего не просили во имя Мое; просите, и получите, чтобы радость ваша была совершенна.
JOHN|16|25|Доселе Я говорил вам притчами; но наступает время, когда уже не буду говорить вам притчами, но прямо возвещу вам об Отце.
JOHN|16|26|В тот день будете просить во имя Мое, и не говорю вам, что Я буду просить Отца о вас:
JOHN|16|27|ибо Сам Отец любит вас, потому что вы возлюбили Меня и уверовали, что Я исшел от Бога.
JOHN|16|28|Я исшел от Отца и пришел в мир; и опять оставляю мир и иду к Отцу.
JOHN|16|29|Ученики Его сказали Ему: вот, теперь Ты прямо говоришь, и притчи не говоришь никакой.
JOHN|16|30|Теперь видим, что Ты знаешь все и не имеешь нужды, чтобы кто спрашивал Тебя. Посему веруем, что Ты от Бога исшел.
JOHN|16|31|Иисус отвечал им: теперь веруете?
JOHN|16|32|Вот, наступает час, и настал уже, что вы рассеетесь каждый в свою [сторону] и Меня оставите одного; но Я не один, потому что Отец со Мною.
JOHN|16|33|Сие сказал Я вам, чтобы вы имели во Мне мир. В мире будете иметь скорбь; но мужайтесь: Я победил мир.
JOHN|17|1|После сих слов Иисус возвел очи Свои на небо и сказал: Отче! пришел час, прославь Сына Твоего, да и Сын Твой прославит Тебя,
JOHN|17|2|так как Ты дал Ему власть над всякою плотью, да всему, что Ты дал Ему, даст Он жизнь вечную.
JOHN|17|3|Сия же есть жизнь вечная, да знают Тебя, единого истинного Бога, и посланного Тобою Иисуса Христа.
JOHN|17|4|Я прославил Тебя на земле, совершил дело, которое Ты поручил Мне исполнить.
JOHN|17|5|И ныне прославь Меня Ты, Отче, у Тебя Самого славою, которую Я имел у Тебя прежде бытия мира.
JOHN|17|6|Я открыл имя Твое человекам, которых Ты дал Мне от мира; они были Твои, и Ты дал их Мне, и они сохранили слово Твое.
JOHN|17|7|Ныне уразумели они, что все, что Ты дал Мне, от Тебя есть,
JOHN|17|8|ибо слова, которые Ты дал Мне, Я передал им, и они приняли, и уразумели истинно, что Я исшел от Тебя, и уверовали, что Ты послал Меня.
JOHN|17|9|Я о них молю: не о всем мире молю, но о тех, которых Ты дал Мне, потому что они Твои.
JOHN|17|10|И все Мое Твое, и Твое Мое; и Я прославился в них.
JOHN|17|11|Я уже не в мире, но они в мире, а Я к Тебе иду. Отче Святый! соблюди их во имя Твое, [тех], которых Ты Мне дал, чтобы они были едино, как и Мы.
JOHN|17|12|Когда Я был с ними в мире, Я соблюдал их во имя Твое; тех, которых Ты дал Мне, Я сохранил, и никто из них не погиб, кроме сына погибели, да сбудется Писание.
JOHN|17|13|Ныне же к Тебе иду, и сие говорю в мире, чтобы они имели в себе радость Мою совершенную.
JOHN|17|14|Я передал им слово Твое; и мир возненавидел их, потому что они не от мира, как и Я не от мира.
JOHN|17|15|Не молю, чтобы Ты взял их из мира, но чтобы сохранил их от зла.
JOHN|17|16|Они не от мира, как и Я не от мира.
JOHN|17|17|Освяти их истиною Твоею; слово Твое есть истина.
JOHN|17|18|Как Ты послал Меня в мир, [так] и Я послал их в мир.
JOHN|17|19|И за них Я посвящаю Себя, чтобы и они были освящены истиною.
JOHN|17|20|Не о них же только молю, но и о верующих в Меня по слову их,
JOHN|17|21|да будут все едино, как Ты, Отче, во Мне, и Я в Тебе, [так] и они да будут в Нас едино, – да уверует мир, что Ты послал Меня.
JOHN|17|22|И славу, которую Ты дал Мне, Я дал им: да будут едино, как Мы едино.
JOHN|17|23|Я в них, и Ты во Мне; да будут совершены воедино, и да познает мир, что Ты послал Меня и возлюбил их, как возлюбил Меня.
JOHN|17|24|Отче! которых Ты дал Мне, хочу, чтобы там, где Я, и они были со Мною, да видят славу Мою, которую Ты дал Мне, потому что возлюбил Меня прежде основания мира.
JOHN|17|25|Отче праведный! и мир Тебя не познал; а Я познал Тебя, и сии познали, что Ты послал Меня.
JOHN|17|26|И Я открыл им имя Твое и открою, да любовь, которою Ты возлюбил Меня, в них будет, и Я в них.
JOHN|18|1|Сказав сие, Иисус вышел с учениками Своими за поток Кедрон, где был сад, в который вошел Сам и ученики Его.
JOHN|18|2|Знал же это место и Иуда, предатель Его, потому что Иисус часто собирался там с учениками Своими.
JOHN|18|3|Итак Иуда, взяв отряд [воинов] и служителей от первосвященников и фарисеев, приходит туда с фонарями и светильниками и оружием.
JOHN|18|4|Иисус же, зная все, что с Ним будет, вышел и сказал им: кого ищете?
JOHN|18|5|Ему отвечали: Иисуса Назорея. Иисус говорит им: это Я. Стоял же с ними и Иуда, предатель Его.
JOHN|18|6|И когда сказал им: это Я, они отступили назад и пали на землю.
JOHN|18|7|Опять спросил их: кого ищете? Они сказали: Иисуса Назорея.
JOHN|18|8|Иисус отвечал: Я сказал вам, что это Я; итак, если Меня ищете, оставьте их, пусть идут,
JOHN|18|9|да сбудется слово, реченное Им: из тех, которых Ты Мне дал, Я не погубил никого.
JOHN|18|10|Симон же Петр, имея меч, извлек его, и ударил первосвященнического раба, и отсек ему правое ухо. Имя рабу было Малх.
JOHN|18|11|Но Иисус сказал Петру: вложи меч в ножны; неужели Мне не пить чаши, которую дал Мне Отец?
JOHN|18|12|Тогда воины и тысяченачальник и служители Иудейские взяли Иисуса и связали Его,
JOHN|18|13|и отвели Его сперва к Анне, ибо он был тесть Каиафе, который был на тот год первосвященником.
JOHN|18|14|Это был Каиафа, который подал совет Иудеям, что лучше одному человеку умереть за народ.
JOHN|18|15|За Иисусом следовали Симон Петр и другой ученик; ученик же сей был знаком первосвященнику и вошел с Иисусом во двор первосвященнический.
JOHN|18|16|А Петр стоял вне за дверями. Потом другой ученик, который был знаком первосвященнику, вышел, и сказал придвернице, и ввел Петра.
JOHN|18|17|Тут раба придверница говорит Петру: и ты не из учеников ли Этого Человека? Он сказал: нет.
JOHN|18|18|Между тем рабы и служители, разведя огонь, потому что было холодно, стояли и грелись. Петр также стоял с ними и грелся.
JOHN|18|19|Первосвященник же спросил Иисуса об учениках Его и об учении Его.
JOHN|18|20|Иисус отвечал ему: Я говорил явно миру; Я всегда учил в синагоге и в храме, где всегда Иудеи сходятся, и тайно не говорил ничего.
JOHN|18|21|Что спрашиваешь Меня? спроси слышавших, что Я говорил им; вот, они знают, что Я говорил.
JOHN|18|22|Когда Он сказал это, один из служителей, стоявший близко, ударил Иисуса по щеке, сказав: так отвечаешь Ты первосвященнику?
JOHN|18|23|Иисус отвечал ему: если Я сказал худо, покажи, что худо; а если хорошо, что ты бьешь Меня?
JOHN|18|24|Анна послал Его связанного к первосвященнику Каиафе.
JOHN|18|25|Симон же Петр стоял и грелся. Тут сказали ему: не из учеников ли Его и ты? Он отрекся и сказал: нет.
JOHN|18|26|Один из рабов первосвященнических, родственник тому, которому Петр отсек ухо, говорит: не я ли видел тебя с Ним в саду?
JOHN|18|27|Петр опять отрекся; и тотчас запел петух.
JOHN|18|28|От Каиафы повели Иисуса в преторию. Было утро; и они не вошли в преторию, чтобы не оскверниться, но чтобы [можно было] есть пасху.
JOHN|18|29|Пилат вышел к ним и сказал: в чем вы обвиняете Человека Сего?
JOHN|18|30|Они сказали ему в ответ: если бы Он не был злодей, мы не предали бы Его тебе.
JOHN|18|31|Пилат сказал им: возьмите Его вы, и по закону вашему судите Его. Иудеи сказали ему: нам не позволено предавать смерти никого, –
JOHN|18|32|да сбудется слово Иисусово, которое сказал Он, давая разуметь, какою смертью Он умрет.
JOHN|18|33|Тогда Пилат опять вошел в преторию, и призвал Иисуса, и сказал Ему: Ты Царь Иудейский?
JOHN|18|34|Иисус отвечал ему: от себя ли ты говоришь это, или другие сказали тебе о Мне?
JOHN|18|35|Пилат отвечал: разве я Иудей? Твой народ и первосвященники предали Тебя мне; что Ты сделал?
JOHN|18|36|Иисус отвечал: Царство Мое не от мира сего; если бы от мира сего было Царство Мое, то служители Мои подвизались бы за Меня, чтобы Я не был предан Иудеям; но ныне Царство Мое не отсюда.
JOHN|18|37|Пилат сказал Ему: итак Ты Царь? Иисус отвечал: ты говоришь, что Я Царь. Я на то родился и на то пришел в мир, чтобы свидетельствовать о истине; всякий, кто от истины, слушает гласа Моего.
JOHN|18|38|Пилат сказал Ему: что есть истина? И, сказав это, опять вышел к Иудеям и сказал им: я никакой вины не нахожу в Нем.
JOHN|18|39|Есть же у вас обычай, чтобы я одного отпускал вам на Пасху; хотите ли, отпущу вам Царя Иудейского?
JOHN|18|40|Тогда опять закричали все, говоря: не Его, но Варавву. Варавва же был разбойник.
JOHN|19|1|Тогда Пилат взял Иисуса и [велел] бить Его.
JOHN|19|2|И воины, сплетши венец из терна, возложили Ему на голову, и одели Его в багряницу,
JOHN|19|3|и говорили: радуйся, Царь Иудейский! и били Его по ланитам.
JOHN|19|4|Пилат опять вышел и сказал им: вот, я вывожу Его к вам, чтобы вы знали, что я не нахожу в Нем никакой вины.
JOHN|19|5|Тогда вышел Иисус в терновом венце и в багрянице. И сказал им [Пилат]: се, Человек!
JOHN|19|6|Когда же увидели Его первосвященники и служители, то закричали: распни, распни Его! Пилат говорит им: возьмите Его вы, и распните; ибо я не нахожу в Нем вины.
JOHN|19|7|Иудеи отвечали ему: мы имеем закон, и по закону нашему Он должен умереть, потому что сделал Себя Сыном Божиим.
JOHN|19|8|Пилат, услышав это слово, больше убоялся.
JOHN|19|9|И опять вошел в преторию и сказал Иисусу: откуда Ты? Но Иисус не дал ему ответа.
JOHN|19|10|Пилат говорит Ему: мне ли не отвечаешь? не знаешь ли, что я имею власть распять Тебя и власть имею отпустить Тебя?
JOHN|19|11|Иисус отвечал: ты не имел бы надо Мною никакой власти, если бы не было дано тебе свыше; посему более греха на том, кто предал Меня тебе.
JOHN|19|12|С этого [времени] Пилат искал отпустить Его. Иудеи же кричали: если отпустишь Его, ты не друг кесарю; всякий, делающий себя царем, противник кесарю.
JOHN|19|13|Пилат, услышав это слово, вывел вон Иисуса и сел на судилище, на месте, называемом Лифостротон, а по–еврейски Гаввафа.
JOHN|19|14|Тогда была пятница перед Пасхою, и час шестый. И сказал [Пилат] Иудеям: се, Царь ваш!
JOHN|19|15|Но они закричали: возьми, возьми, распни Его! Пилат говорит им: Царя ли вашего распну? Первосвященники отвечали: нет у нас царя, кроме кесаря.
JOHN|19|16|Тогда наконец он предал Его им на распятие. И взяли Иисуса и повели.
JOHN|19|17|И, неся крест Свой, Он вышел на место, называемое Лобное, по–еврейски Голгофа;
JOHN|19|18|там распяли Его и с Ним двух других, по ту и по другую сторону, а посреди Иисуса.
JOHN|19|19|Пилат же написал и надпись, и поставил на кресте. Написано было: Иисус Назорей, Царь Иудейский.
JOHN|19|20|Эту надпись читали многие из Иудеев, потому что место, где был распят Иисус, было недалеко от города, и написано было по–еврейски, по–гречески, по–римски.
JOHN|19|21|Первосвященники же Иудейские сказали Пилату: не пиши: Царь Иудейский, но что Он говорил: Я Царь Иудейский.
JOHN|19|22|Пилат отвечал: что я написал, то написал.
JOHN|19|23|Воины же, когда распяли Иисуса, взяли одежды Его и разделили на четыре части, каждому воину по части, и хитон; хитон же был не сшитый, а весь тканый сверху.
JOHN|19|24|Итак сказали друг другу: не станем раздирать его, а бросим о нем жребий, чей будет, – да сбудется реченное в Писании: разделили ризы Мои между собою и об одежде Моей бросали жребий. Так поступили воины.
JOHN|19|25|При кресте Иисуса стояли Матерь Его и сестра Матери Его, Мария Клеопова, и Мария Магдалина.
JOHN|19|26|Иисус, увидев Матерь и ученика тут стоящего, которого любил, говорит Матери Своей: Жено! се, сын Твой.
JOHN|19|27|Потом говорит ученику: се, Матерь твоя! И с этого времени ученик сей взял Ее к себе.
JOHN|19|28|После того Иисус, зная, что уже все совершилось, да сбудется Писание, говорит: жажду.
JOHN|19|29|Тут стоял сосуд, полный уксуса. [Воины], напоив уксусом губку и наложив на иссоп, поднесли к устам Его.
JOHN|19|30|Когда же Иисус вкусил уксуса, сказал: совершилось! И, преклонив главу, предал дух.
JOHN|19|31|Но так как [тогда] была пятница, то Иудеи, дабы не оставить тел на кресте в субботу, – ибо та суббота была день великий, – просили Пилата, чтобы перебить у них голени и снять их.
JOHN|19|32|Итак пришли воины, и у первого перебили голени, и у другого, распятого с Ним.
JOHN|19|33|Но, придя к Иисусу, как увидели Его уже умершим, не перебили у Него голеней,
JOHN|19|34|но один из воинов копьем пронзил Ему ребра, и тотчас истекла кровь и вода.
JOHN|19|35|И видевший засвидетельствовал, и истинно свидетельство его; он знает, что говорит истину, дабы вы поверили.
JOHN|19|36|Ибо сие произошло, да сбудется Писание: кость Его да не сокрушится.
JOHN|19|37|Также и в другом [месте] Писание говорит: воззрят на Того, Которого пронзили.
JOHN|19|38|После сего Иосиф из Аримафеи – ученик Иисуса, но тайный из страха от Иудеев, – просил Пилата, чтобы снять тело Иисуса; и Пилат позволил. Он пошел и снял тело Иисуса.
JOHN|19|39|Пришел также и Никодим, – приходивший прежде к Иисусу ночью, – и принес состав из смирны и алоя, литр около ста.
JOHN|19|40|Итак они взяли тело Иисуса и обвили его пеленами с благовониями, как обыкновенно погребают Иудеи.
JOHN|19|41|На том месте, где Он распят, был сад, и в саду гроб новый, в котором еще никто не был положен.
JOHN|19|42|Там положили Иисуса ради пятницы Иудейской, потому что гроб был близко.
JOHN|20|1|В первый же [день] недели Мария Магдалина приходит ко гробу рано, когда было еще темно, и видит, что камень отвален от гроба.
JOHN|20|2|Итак, бежит и приходит к Симону Петру и к другому ученику, которого любил Иисус, и говорит им: унесли Господа из гроба, и не знаем, где положили Его.
JOHN|20|3|Тотчас вышел Петр и другой ученик, и пошли ко гробу.
JOHN|20|4|Они побежали оба вместе; но другой ученик бежал скорее Петра, и пришел ко гробу первый.
JOHN|20|5|И, наклонившись, увидел лежащие пелены; но не вошел [во гроб].
JOHN|20|6|Вслед за ним приходит Симон Петр, и входит во гроб, и видит одни пелены лежащие,
JOHN|20|7|и плат, который был на главе Его, не с пеленами лежащий, но особо свитый на другом месте.
JOHN|20|8|Тогда вошел и другой ученик, прежде пришедший ко гробу, и увидел, и уверовал.
JOHN|20|9|Ибо они еще не знали из Писания, что Ему надлежало воскреснуть из мертвых.
JOHN|20|10|Итак ученики опять возвратились к себе.
JOHN|20|11|А Мария стояла у гроба и плакала. И, когда плакала, наклонилась во гроб,
JOHN|20|12|и видит двух Ангелов, в белом одеянии сидящих, одного у главы и другого у ног, где лежало тело Иисуса.
JOHN|20|13|И они говорят ей: жена! что ты плачешь? Говорит им: унесли Господа моего, и не знаю, где положили Его.
JOHN|20|14|Сказав сие, обратилась назад и увидела Иисуса стоящего; но не узнала, что это Иисус.
JOHN|20|15|Иисус говорит ей: жена! что ты плачешь? кого ищешь? Она, думая, что это садовник, говорит Ему: господин! если ты вынес Его, скажи мне, где ты положил Его, и я возьму Его.
JOHN|20|16|Иисус говорит ей: Мария! Она, обратившись, говорит Ему: Раввуни! – что значит: Учитель!
JOHN|20|17|Иисус говорит ей: не прикасайся ко Мне, ибо Я еще не восшел к Отцу Моему; а иди к братьям Моим и скажи им: восхожу к Отцу Моему и Отцу вашему, и к Богу Моему и Богу вашему.
JOHN|20|18|Мария Магдалина идет и возвещает ученикам, [что] видела Господа и [что] Он это сказал ей.
JOHN|20|19|В тот же первый день недели вечером, когда двери [дома], где собирались ученики Его, были заперты из опасения от Иудеев, пришел Иисус, и стал посреди, и говорит им: мир вам!
JOHN|20|20|Сказав это, Он показал им руки и ноги и ребра Свои. Ученики обрадовались, увидев Господа.
JOHN|20|21|Иисус же сказал им вторично: мир вам! как послал Меня Отец, [так] и Я посылаю вас.
JOHN|20|22|Сказав это, дунул, и говорит им: примите Духа Святаго.
JOHN|20|23|Кому простите грехи, тому простятся; на ком оставите, на том останутся.
JOHN|20|24|Фома же, один из двенадцати, называемый Близнец, не был тут с ними, когда приходил Иисус.
JOHN|20|25|Другие ученики сказали ему: мы видели Господа. Но он сказал им: если не увижу на руках Его ран от гвоздей, и не вложу перста моего в раны от гвоздей, и не вложу руки моей в ребра Его, не поверю.
JOHN|20|26|После восьми дней опять были в доме ученики Его, и Фома с ними. Пришел Иисус, когда двери были заперты, стал посреди них и сказал: мир вам!
JOHN|20|27|Потом говорит Фоме: подай перст твой сюда и посмотри руки Мои; подай руку твою и вложи в ребра Мои; и не будь неверующим, но верующим.
JOHN|20|28|Фома сказал Ему в ответ: Господь мой и Бог мой!
JOHN|20|29|Иисус говорит ему: ты поверил, потому что увидел Меня; блаженны невидевшие и уверовавшие.
JOHN|20|30|Много сотворил Иисус пред учениками Своими и других чудес, о которых не писано в книге сей.
JOHN|20|31|Сие же написано, дабы вы уверовали, что Иисус есть Христос, Сын Божий, и, веруя, имели жизнь во имя Его.
JOHN|21|1|После того опять явился Иисус ученикам Своим при море Тивериадском. Явился же так:
JOHN|21|2|были вместе Симон Петр, и Фома, называемый Близнец, и Нафанаил из Каны Галилейской, и сыновья Зеведеевы, и двое других из учеников Его.
JOHN|21|3|Симон Петр говорит им: иду ловить рыбу. Говорят ему: идем и мы с тобою. Пошли и тотчас вошли в лодку, и не поймали в ту ночь ничего.
JOHN|21|4|А когда уже настало утро, Иисус стоял на берегу; но ученики не узнали, что это Иисус.
JOHN|21|5|Иисус говорит им: дети! есть ли у вас какая пища? Они отвечали Ему: нет.
JOHN|21|6|Он же сказал им: закиньте сеть по правую сторону лодки, и поймаете. Они закинули, и уже не могли вытащить [сети] от множества рыбы.
JOHN|21|7|Тогда ученик, которого любил Иисус, говорит Петру: это Господь. Симон же Петр, услышав, что это Господь, опоясался одеждою, – ибо он был наг, – и бросился в море.
JOHN|21|8|А другие ученики приплыли в лодке, – ибо недалеко были от земли, локтей около двухсот, – таща сеть с рыбою.
JOHN|21|9|Когда же вышли на землю, видят разложенный огонь и на нем лежащую рыбу и хлеб.
JOHN|21|10|Иисус говорит им: принесите рыбы, которую вы теперь поймали.
JOHN|21|11|Симон Петр пошел и вытащил на землю сеть, наполненную большими рыбами, [которых было] сто пятьдесят три; и при таком множестве не прорвалась сеть.
JOHN|21|12|Иисус говорит им: придите, обедайте. Из учеников же никто не смел спросить Его: кто Ты?, зная, что это Господь.
JOHN|21|13|Иисус приходит, берет хлеб и дает им, также и рыбу.
JOHN|21|14|Это уже в третий раз явился Иисус ученикам Своим по воскресении Своем из мертвых.
JOHN|21|15|Когда же они обедали, Иисус говорит Симону Петру: Симон Ионин! любишь ли ты Меня больше, нежели они? [Петр] говорит Ему: так, Господи! Ты знаешь, что я люблю Тебя. [Иисус] говорит ему: паси агнцев Моих.
JOHN|21|16|Еще говорит ему в другой раз: Симон Ионин! любишь ли ты Меня? [Петр] говорит Ему: так, Господи! Ты знаешь, что я люблю Тебя. [Иисус] говорит ему: паси овец Моих.
JOHN|21|17|Говорит ему в третий раз: Симон Ионин! любишь ли ты Меня? Петр опечалился, что в третий раз спросил его: любишь ли Меня? и сказал Ему: Господи! Ты все знаешь; Ты знаешь, что я люблю Тебя. Иисус говорит ему: паси овец Моих.
JOHN|21|18|Истинно, истинно говорю тебе: когда ты был молод, то препоясывался сам и ходил, куда хотел; а когда состаришься, то прострешь руки твои, и другой препояшет тебя, и поведет, куда не хочешь.
JOHN|21|19|Сказал же это, давая разуметь, какою смертью [Петр] прославит Бога. И, сказав сие, говорит ему: иди за Мною.
JOHN|21|20|Петр же, обратившись, видит идущего за ним ученика, которого любил Иисус и который на вечери, приклонившись к груди Его, сказал: Господи! кто предаст Тебя?
JOHN|21|21|Его увидев, Петр говорит Иисусу: Господи! а он что?
JOHN|21|22|Иисус говорит ему: если Я хочу, чтобы он пребыл, пока приду, что тебе [до того]? ты иди за Мною.
JOHN|21|23|И пронеслось это слово между братиями, что ученик тот не умрет. Но Иисус не сказал ему, что не умрет, но: если Я хочу, чтобы он пребыл, пока приду, что тебе [до того]?
JOHN|21|24|Сей ученик и свидетельствует о сем, и написал сие; и знаем, что истинно свидетельство его.
JOHN|21|25|Многое и другое сотворил Иисус; но, если бы писать о том подробно, то, думаю, и самому миру не вместить бы написанных книг. Аминь.
