2CHR|1|1|大卫 的儿子 所罗门 巩固他的国度；耶和华－他的上帝与他同在，使他极其尊大。
2CHR|1|2|所罗门 吩咐全 以色列 ，就是千夫长、百夫长、审判官、全 以色列 的众领袖和族长前来。
2CHR|1|3|所罗门 率领全会众往 基遍 的丘坛去，因那里有上帝的会幕，就是耶和华的仆人 摩西 在旷野所造的。
2CHR|1|4|只是上帝的约柜， 大卫 已经从 基列．耶琳 接到他所预备的地方，因他曾在 耶路撒冷 为约柜支搭了帐幕，
2CHR|1|5|把 户珥 的孙子， 乌利 的儿子 比撒列 所造的铜坛摆在 基遍 耶和华的会幕前。 所罗门 和会众求告耶和华。
2CHR|1|6|所罗门 上到耶和华面前会幕的铜坛那里，在坛上献一千祭牲为燔祭。
2CHR|1|7|当夜，上帝向 所罗门 显现，对他说：“你愿我赐你什么，你可以求。”
2CHR|1|8|所罗门 对上帝说：“你曾向我父亲 大卫 大施慈爱，使我接续他作王。
2CHR|1|9|耶和华上帝啊，现在求你实现向我父亲 大卫 所应许的话；因你立我作这百姓的王，他们如同地上的尘沙那样多。
2CHR|1|10|现在，求你赐我智慧聪明，好在这百姓面前出入；不然，谁能判断你这么多的百姓呢？”
2CHR|1|11|上帝对 所罗门 说：“你有这心意，不求资财、丰富、尊荣，也不求灭绝恨你之人的性命，又不求长寿；我既立你作我百姓的王，你只求智慧聪明，好审判我的百姓，
2CHR|1|12|我必赐你智慧聪明，也必赐你资财、丰富、尊荣，在你以前的列王未曾有过，在你以后也不会再有。”
2CHR|1|13|于是， 所罗门 从 基遍 丘坛会幕前回到 耶路撒冷 ，治理 以色列 。
2CHR|1|14|所罗门 聚集战车骑兵；他有一千四百辆战车，一万二千名骑兵，安置在屯车城，在 耶路撒冷 的王那里。
2CHR|1|15|王在 耶路撒冷 使金银多如石头，香柏木多如 谢非拉 的桑树。
2CHR|1|16|所罗门 的马是从 埃及 和 科威 运来的，是王的商人按着定价从 科威 买来的。
2CHR|1|17|他们从 埃及 进口战车，每辆六百舍客勒银子，马每匹一百五十舍客勒； 赫 人众王和 亚兰 诸王的战车和马，也是经由他们的手出口的。
2CHR|2|1|所罗门 吩咐要为耶和华的名建造殿宇，又为自己的王国建造宫殿。
2CHR|2|2|所罗门 征召七万名扛抬的，八万个在山上凿石头的人，三千六百个监工。
2CHR|2|3|所罗门 派人去见 推罗 王 希兰 ，说：“你曾运香柏木给我父亲 大卫 建造宫殿居住，请你也这样待我。
2CHR|2|4|看哪，我要为耶和华－我上帝的名建造殿宇，分别为圣献给他，在他面前烧芬芳的香，经常献供饼，每早晚、安息日、初一，以及耶和华－我们上帝所定的节期献燔祭。这是 以色列 人永远的定例。
2CHR|2|5|我所要建造的殿宇宏大，因为我们的上帝至大，超乎众神。
2CHR|2|6|天和天上的天，尚且不足他居住，谁能为他建造殿宇呢？我是谁，能为他建造殿宇吗？不过在他面前烧香而已！
2CHR|2|7|现在请你派一个巧匠来，就是善用金、银、铜、铁，和紫色、朱红色、蓝色线做工，并精于雕刻之工的巧匠，与跟我一起在 犹大 和 耶路撒冷 、我父亲 大卫 所预备的巧匠一同做工；
2CHR|2|8|又请你从 黎巴嫩 运香柏木、松木、檀香木到我这里来，因我知道你的仆人擅长砍伐 黎巴嫩 的树木。看哪，我的仆人必帮助你的仆人，
2CHR|2|9|好为我预备许多的木料，因我要建造的殿宇高大出奇。
2CHR|2|10|看哪，我必给你仆人，就是砍伐树木的伐木工，二万歌珥压碎的小麦 ，二万歌珥大麦，二万罢特酒，二万罢特油。”
2CHR|2|11|推罗 王 希兰 写信回答 所罗门 说：“耶和华因为爱他的百姓，所以立你作他们的王。”
2CHR|2|12|又说：“创造天和地的耶和华－ 以色列 的上帝是应当称颂的！他赐给 大卫 王一个有智慧的儿子，使他有见识，有聪明，可以为耶和华建造殿宇，又为自己的王国建造宫殿。
2CHR|2|13|“现在我派一个精巧聪明的人去，他是我的师父 户兰 ，
2CHR|2|14|是 但 支派一个妇人的儿子，父亲是 推罗 人。他善用金、银、铜、铁、石、木，和紫色、蓝色、细麻和朱红色线制造各物，并精于雕刻，又能设计各样交给他做的图案。我派这人与你的巧匠和你父亲－我主 大卫 的巧匠一同做工。
2CHR|2|15|我主所说的小麦、大麦、酒、油，请运来给众仆人。
2CHR|2|16|我们必照你所需用的，从 黎巴嫩 砍伐树木，扎成筏子，浮海运到 约帕 ；你可以从那里运到 耶路撒冷 。”
2CHR|2|17|所罗门 仿照他父亲 大卫 数点所有在 以色列 地寄居的外邦人，共有十五万三千六百名。
2CHR|2|18|他叫其中的七万人作扛抬，八万人在山上凿石头，三千六百人监督百姓工作。
2CHR|3|1|所罗门 在 耶路撒冷 开工建造耶和华的殿，就在耶和华向他父亲 大卫 显现的 摩利亚山 上， 耶布斯 人 阿珥楠 的禾场， 大卫 指定的地方。
2CHR|3|2|所罗门 作王第四年二月初二 开工建造。
2CHR|3|3|所罗门 所建筑的上帝殿的根基是这样：长六十肘，宽二十肘，都按着古时的尺寸。
2CHR|3|4|前面的 走廊长二十肘，与殿的宽度一样，高一百二十肘；里面贴上纯金。
2CHR|3|5|大殿的墙都用松木板遮蔽，又贴上纯金，上面刻着棕树和链子。
2CHR|3|6|他用宝石装饰这殿，使殿华美；金子都是 巴瓦音 的金子。
2CHR|3|7|他用金子贴殿和殿的栋梁、门槛、墙壁、门扇；墙上刻着基路伯。
2CHR|3|8|他建造至圣所，长二十肘，与殿的宽度一样，宽二十肘，都贴上纯金，共用了六百他连得金子。
2CHR|3|9|金的钉子重五十舍客勒。楼房都贴上金子。
2CHR|3|10|他又在至圣所用雕刻的手艺造两个基路伯，包上金子。
2CHR|3|11|两个基路伯的翅膀共长二十肘。这基路伯的一个翅膀长五肘，挨着殿这边的墙；另一个翅膀也长五肘，与那基路伯翅膀相接。
2CHR|3|12|那基路伯的一个翅膀长五肘，挨着殿那边的墙；另一个翅膀也长五肘，与这基路伯的翅膀相接。
2CHR|3|13|这两个基路伯张开翅膀，共长二十肘，用脚站立，脸面向殿。
2CHR|3|14|他又用蓝色、紫色、朱红色线和细麻织幔子，在其上绣基路伯。
2CHR|3|15|他在殿前造了两根柱子，高三十五肘；柱子上面的柱顶高五肘。
2CHR|3|16|他造链子在内殿里，安在柱顶上，又做一百个石榴，安在链子上。
2CHR|3|17|他把两根柱子立在殿前，一根在右边，一根在左边；右边的起名叫 雅斤 ，左边的起名叫 波阿斯 。
2CHR|4|1|他造一座铜坛，长二十肘，宽二十肘，高十肘。
2CHR|4|2|他又铸一个铜海，周围是圆的，直径十肘，高五肘，用绳子量周围是三十肘。
2CHR|4|3|铜海下面的周围有牛的样式，有十肘，绕着铜海；牛有两行，是造铜海的时候铸上去的。
2CHR|4|4|铜海安在十二头铜牛上：三头向北，三头向西，三头向南，三头向东。铜海安在牛上，牛尾都向内。
2CHR|4|5|铜海厚一掌，边如杯边，像百合花，容量是三千罢特。
2CHR|4|6|他又造十个盆：五个放在右边，五个放在左边，作洗涤之用。献燔祭所用之物都洗在盆内；但铜海是为祭司洗涤用的。
2CHR|4|7|他照所定的样式造十个金灯台，放在殿里：五个在右边，五个在左边。
2CHR|4|8|他造十张桌子，放在殿里：五张在右边，五张在左边。他又造一百个金碗。
2CHR|4|9|他建造祭司院和大院，以及院门，门扇包上铜。
2CHR|4|10|他把铜海安在殿的右边，就是东南边。
2CHR|4|11|户兰 又造了盆、铲子和盘子。这样， 户兰 为 所罗门 王做完了上帝殿的工：
2CHR|4|12|两根柱子和柱子顶上两个如碗的柱顶，以及盖着如碗柱顶的两个网子；
2CHR|4|13|四百个石榴，安在两个网子上，每网两行石榴，盖着柱子上面两个如碗的柱顶。
2CHR|4|14|他造盆座，又造其上的盆；
2CHR|4|15|铜海和其下的十二头牛；
2CHR|4|16|盆、铲子、肉叉。巧匠 户兰 给 所罗门 王为耶和华殿造的这一切器皿都是用磨亮的铜，
2CHR|4|17|是王在 约旦 平原、 疏割 和 撒利但 中间的泥巴地铸成的。
2CHR|4|18|所罗门 造这一切器皿，数量很多，铜的重量无法计算。
2CHR|4|19|所罗门 又为上帝的殿造了各样的器皿：金坛和献供饼的供桌；
2CHR|4|20|纯金的灯台和灯盏，可以照定例点在内殿前；
2CHR|4|21|灯台上的花和灯盏，以及灯剪，都是金的，而且是纯金的；
2CHR|4|22|纯金的钳子、盘子、勺子、火盆。至于殿门和至圣所的门扇，以及殿的门扇，都是金的。
2CHR|5|1|所罗门 王做完了耶和华殿一切的工，就把他父亲 大卫 分别为圣的金银和一切器皿都带来，放在上帝殿的库房里。
2CHR|5|2|于是， 所罗门 召集 以色列 的长老、各支派的领袖和 以色列 人的族长到 耶路撒冷 ，要把耶和华的约柜从 大卫城 ，就是 锡安 ，接上来。
2CHR|5|3|在七月节期的时候，所有的 以色列 人都聚集到王那里。
2CHR|5|4|以色列 众长老一来到， 利未 人就抬起约柜。
2CHR|5|5|祭司和 利未 人将约柜请上来，又把会幕和会幕一切的圣器皿都带上来。
2CHR|5|6|所罗门 王和聚集到他那里的 以色列 全会众都在约柜前献牛羊为祭，多得不可胜数，无法计算。
2CHR|5|7|祭司将耶和华的约柜请进内殿，就是至圣所，安置在两个基路伯的翅膀底下约柜自己的地方。
2CHR|5|8|基路伯张开翅膀在约柜上面的地方，从上面遮住约柜和抬柜的杠。
2CHR|5|9|这杠很长，从内殿前的约柜可以看见杠头，从外面却看不见。这杠直到今日还在那里。
2CHR|5|10|约柜里没有别的，只有两块石版，就是 以色列 人出 埃及 ，耶和华与他们立约的时候， 摩西 在 何烈山 所放的。
2CHR|5|11|当时，所有在那里的祭司，不论哪个班次供职的，都使自己分别为圣。祭司从圣所出来的时候，
2CHR|5|12|所有歌唱的 利未 人， 亚萨 、 希幔 、 耶杜顿 ，和他们的众儿子、众弟兄都穿细麻布衣服，站在祭坛的东边敲钹，鼓瑟，弹琴，和他们一起的还有一百二十个吹号的祭司。
2CHR|5|13|吹号的、歌唱的都合一齐声，赞美称谢耶和华。他们配合号筒、铙钹和其他乐器，扬声赞美耶和华： “耶和华本为善， 他的慈爱永远长存！” 那时，耶和华的殿充满了云彩。
2CHR|5|14|祭司因云彩的缘故不能站立供职，因为耶和华的荣光充满了上帝的殿。
2CHR|6|1|那时， 所罗门 说： “耶和华曾说要住在幽暗之处。
2CHR|6|2|我为你建了一座雄伟的殿宇， 作为你永远居住的地方。”
2CHR|6|3|王转过脸来为 以色列 全会众祝福， 以色列 全会众都站立。
2CHR|6|4|所罗门 说：“耶和华－ 以色列 的上帝是应当称颂的！因他亲口向我父 大卫 应许的，也亲手成就了；他曾说：
2CHR|6|5|‘自从那日我领我百姓出 埃及 地以来，我未曾在 以色列 各支派中选择一城，在那里为我的名建造殿宇，也未曾拣选一人作我百姓 以色列 的君王。
2CHR|6|6|但我选择 耶路撒冷 ，使我的名留在那里，又拣选 大卫 治理我的百姓 以色列 。’
2CHR|6|7|我父 大卫 的心意是要为耶和华－ 以色列 上帝的名建殿。
2CHR|6|8|耶和华却对我父 大卫 说：‘你有心为我的名建殿，这心意是好的；
2CHR|6|9|但你不可建殿，惟有你亲生的儿子才可为我的名建殿。’
2CHR|6|10|现在耶和华实现了他所应许的话，使我接续我父 大卫 坐 以色列 的王位，正如耶和华所说的，我也为耶和华－ 以色列 上帝的名建造了这殿。
2CHR|6|11|我将约柜安置在那里，柜内有耶和华的约，就是他与 以色列 人所立的约。”
2CHR|6|12|所罗门 当着 以色列 全会众，站在耶和华的坛前，举起手来。
2CHR|6|13|所罗门 曾造一个铜台，长五肘，宽五肘，高三肘，放在院中。他站在台上，当着 以色列 全会众双膝跪下，向天举手，
2CHR|6|14|说：“耶和华－ 以色列 的上帝啊，天上地下没有神明可与你相比！你向那些尽心行在你面前的仆人守约施慈爱，
2CHR|6|15|这约是你向你仆人 大卫 守的，是你应许他的。你亲口应许，亲手成就，正如今日一样。
2CHR|6|16|耶和华－ 以色列 的上帝啊，你向你仆人我父 大卫 应许说：‘你的子孙若谨慎自己的行为，遵行我的律法，像你在我面前所行的，就不断有人在我面前坐 以色列 的王位。’现在求你信守这话。
2CHR|6|17|耶和华－ 以色列 的上帝啊，现在求你成就向你仆人 大卫 所应许的话。
2CHR|6|18|“上帝果真与世人同住在地上吗？看哪，天和天上的天尚且不足容纳你，何况我所建的这殿呢？
2CHR|6|19|惟求耶和华－我的上帝垂顾仆人的祷告祈求，俯听仆人在你面前的祈祷呼求。
2CHR|6|20|愿你的眼目昼夜看顾这殿，就是你应许立为你名的居所；求你垂听祷告，你仆人向此处的祷告。
2CHR|6|21|你仆人和你百姓 以色列 向此处祈祷的时候，求你从天上你的居所垂听，垂听而赦免。
2CHR|6|22|“人若得罪邻舍，有人强迫他，要他起誓，他来到这殿，在你的坛前起誓，
2CHR|6|23|求你从天上垂听、处理，向你的仆人施行审判，定恶人有罪，照他所行的报应在他头上；定义人为义，照他的义赏赐他。
2CHR|6|24|“你的百姓 以色列 若得罪你，败在仇敌面前，却又归向你，宣认你的名，在这殿里向你祈求祷告，
2CHR|6|25|求你从天上垂听，赦免你百姓 以色列 的罪，使他们归回你赐给他们和他们列祖之地。
2CHR|6|26|“你的百姓若得罪了你，你使天闭塞不下雨；他们若向此处祷告，宣认你的名，因你的惩罚而离开他们的罪，
2CHR|6|27|求你在天上垂听，赦免你仆人你百姓 以色列 的罪，将当行的善道教导他们，并降雨在你的地，就是你赐给你百姓为业之地。
2CHR|6|28|“这地若有饥荒、瘟疫、焚风 、霉烂、蝗虫、蚂蚱，或有仇敌围困这地的城门，无论遭遇什么灾祸疾病，
2CHR|6|29|你的百姓 以色列 ，或众人或一人，自觉灾祸困苦，向这殿举手，无论祈求什么，祷告什么，
2CHR|6|30|求你从天上你的居所垂听赦免。因为你知道人心，惟有你知道世人的心，求你照各人所行的一切待他们，
2CHR|6|31|使他们在你赐给我们列祖的土地上一生一世敬畏你，遵行你的道。
2CHR|6|32|“论到不属你百姓 以色列 的外邦人，若为你的大名和大能的手，以及伸出来的膀臂，从远方而来，来向这殿祷告，
2CHR|6|33|求你从天上你的居所垂听，照着外邦人向你所求的一切而行，使地上万民都认识你的名，敬畏你，像你的百姓 以色列 一样，又使他们知道我所建造的是称为你名下的殿。
2CHR|6|34|“你的百姓若奉你的派遣出去，无论往何处与仇敌争战，他们若向你所选择的这城和我为你名所建造的殿祷告，
2CHR|6|35|求你从天上垂听他们的祷告祈求，为他们伸张正义。
2CHR|6|36|“你的百姓若得罪你，因为没有人不犯罪，你向他们发怒，把他们交在仇敌面前，掳他们的人把他们带到或远或近之地；
2CHR|6|37|他们若在被掳之地那里回心转意，在被掳之地悔改，向你恳求说：‘我们有罪了，我们悖逆了，我们作恶了’；
2CHR|6|38|他们若在被掳之地尽心尽性归向你，又向自己的地，就是你赐给他们列祖的地和你所选择的城，以及我为你名所建造的这殿祷告，
2CHR|6|39|求你从天上你的居所垂听他们的祷告祈求，为他们伸张正义，赦免你的百姓向你犯的罪。
2CHR|6|40|我的上帝啊，现在求你睁眼看，侧耳听在此处所献的祷告。
2CHR|6|41|“耶和华上帝啊，现在求你兴起， 与你有能力的约柜同入安歇之所。 耶和华上帝啊，愿你的祭司披上救恩， 愿你的圣民蒙福欢乐。
2CHR|6|42|耶和华上帝啊，求你不要厌弃你的受膏者， 要记得向你仆人 大卫 所施的慈爱。”
2CHR|7|1|所罗门 祈祷完毕，就有火从天降下来，烧尽燔祭和祭物。耶和华的荣光充满了殿；
2CHR|7|2|因耶和华的荣光充满了耶和华的殿，所以祭司不能进耶和华的殿。
2CHR|7|3|那火降下、耶和华的荣光在殿上的时候， 以色列 众人看见，就在石板地俯伏敬拜，称谢耶和华： “耶和华本为善， 他的慈爱永远长存！”
2CHR|7|4|王和众百姓在耶和华面前献祭。
2CHR|7|5|所罗门 王献二万二千头牛，十二万只羊为祭。这样，王和众百姓为上帝的殿行了奉献之礼。
2CHR|7|6|祭司各供其职侍立， 利未 人拿着耶和华的乐器，就是 大卫 王所造、为要颂赞耶和华的乐器，因他的慈爱永远长存；他们为 大卫 的赞美诗奏乐；祭司在众人面前吹号， 以色列 众人都站立。
2CHR|7|7|所罗门 因他所造的铜坛容不下燔祭、素祭和脂肪，就将耶和华殿前院子的中间分别为圣，在那里献燔祭和平安祭牲的脂肪。
2CHR|7|8|那时 所罗门 守节七日，从 哈马口 直到 埃及 溪谷的 以色列 众人都与他同在一起，成了一个极其盛大的会。
2CHR|7|9|第八日他们举行严肃会，行奉献坛的礼七日，守节七日。
2CHR|7|10|七月二十三日，王差遣百姓回自己的帐棚去；他们为耶和华向 大卫 和 所罗门 ，以及他百姓 以色列 所施的恩惠，心里都欢喜快乐。
2CHR|7|11|所罗门 建完了耶和华的殿和王宫；在耶和华的殿和王宫的工程上，凡他心中所要做的，都顺利做成了。
2CHR|7|12|夜间耶和华向 所罗门 显现，对他说：“我已听了你的祷告，也选择这地方归我作献祭的殿宇。
2CHR|7|13|我若使天闭塞不下雨，或使蝗虫吃这地的出产，或降瘟疫在我子民中，
2CHR|7|14|这称为我名下的子民，若是谦卑自己，祷告，寻求我的面，转离他们的恶行，我必从天上垂听，赦免他们的罪，医治他们的地。
2CHR|7|15|我必睁眼看，侧耳听在此处所献的祷告。
2CHR|7|16|现在我已选择这殿，分别为圣，使我的名永在其中；我的眼、我的心也必时常在那里。
2CHR|7|17|你若行在我面前，效法你父 大卫 所行的，遵行我一切所吩咐你的，谨守我的律例典章，
2CHR|7|18|我就必坚固你国度的王位，正如我与你父 大卫 所立的约，说：‘你的子孙必不断有人治理 以色列 。’
2CHR|7|19|“倘若你们转去，离弃我摆在你们面前的律例诫命，去事奉别神，敬拜它们，
2CHR|7|20|我就必把 以色列 人从我赐给他们的地上连根拔起，也必从我面前舍弃那为我名所分别为圣的殿，使它在万民中成为笑柄，被人讥诮。
2CHR|7|21|这殿虽然崇高，将来凡经过的人必惊讶说：‘耶和华为何向这地和这殿如此行呢？’
2CHR|7|22|人必说：‘因为此地的人离弃领他们祖先出 埃及 地的耶和华－他们的上帝，去亲近别神，敬拜事奉它们，所以耶和华使这一切灾祸临到他们。’”
2CHR|8|1|所罗门 建造耶和华的殿和王宫，用了二十年才完成。
2CHR|8|2|所罗门 修筑 希兰 送给他的城镇，使 以色列 人住在那里。
2CHR|8|3|所罗门 往 哈马．琐巴 去，攻取了那地方。
2CHR|8|4|所罗门 建造旷野的 达莫 ，建造 哈马 一切的储货城，
2CHR|8|5|又建造 上伯．和仑 、 下伯．和仑 ，成为有墙、门、闩的堡垒城。
2CHR|8|6|所罗门 建造 巴拉 和一切的储货城、战车城、战马城，以及他所想要建造的，在 耶路撒冷 、 黎巴嫩 ，和自己所治理全国中的一切建设。
2CHR|8|7|至于所有剩下的百姓，不属 以色列 的 赫 人、 亚摩利 人、 比利洗 人、 希未 人、 耶布斯 人，
2CHR|8|8|那些 以色列 人在当地不能灭尽的人， 所罗门 征召他们剩下的后代服劳役，直到今日。
2CHR|8|9|惟有 以色列 人， 所罗门 不使他们当奴仆做工，而是作他的战士、军官、战车长、骑兵长。
2CHR|8|10|这些是 所罗门 王的监工，共有二百五十名百姓的监工。
2CHR|8|11|所罗门 把法老的女儿迁出 大卫城 ，上到他为她建造的宫里，因 所罗门 说：“耶和华约柜所到之处都是圣地，所以我的妻子不可住在 以色列 王 大卫 的宫里。”
2CHR|8|12|那时， 所罗门 在走廊前他所筑的耶和华的坛上，向耶和华献燔祭，
2CHR|8|13|又遵照 摩西 的吩咐，在安息日、初一，以及每年在除酵节、七七节、住棚节三个节期，献每日所当献上的祭。
2CHR|8|14|所罗门 照着他父亲 大卫 所定的条例，分派祭司的班次，担任他们的职务，又分派 利未 人的任务，负责颂赞，并在祭司面前做每日当做的事，又派门口的守卫按着班次看守各门，因为神人 大卫 是这样吩咐的。
2CHR|8|15|王对众祭司和 利未 人的吩咐，无论是管理库房或任何事务，他们都不违背。
2CHR|8|16|所罗门 所有的工作都准备就绪，从立耶和华殿的根基直到完工的日子。耶和华的殿就完成了。
2CHR|8|17|那时， 所罗门 往 以东 地海岸的 以旬．迦别 和 以禄 去。
2CHR|8|18|希兰 派他的臣仆，把船只和熟悉航海的仆人送到 所罗门 那里。他们同 所罗门 的仆人到了 俄斐 ，从那里得了四百五十他连得金子，运到 所罗门 王那里。
2CHR|9|1|示巴 女王听见 所罗门 的名声，就来到 耶路撒冷 ，要用难题考问 所罗门 。她带着很多的随从，有骆驼驮着香料、许多金子和宝石。她来到 所罗门 那里，向他提出心中所有的问题。
2CHR|9|2|所罗门 回答了她所有的问题，没有一个问题太难，是 所罗门 不能向她解答的。
2CHR|9|3|示巴 女王看见 所罗门 的智慧和他所建造的宫殿，
2CHR|9|4|席上的食物，坐着的群臣，侍立的仆人和他们的服装，司酒长和他们的服装，以及他上耶和华殿的台阶 ，就诧异得神不守舍。
2CHR|9|5|她对王说：“我在本国所听到的话，论到你的事和你的智慧是真的！
2CHR|9|6|我本来不信那些话，及至我来亲眼看见了，看哪，人所告诉我的，还不及你丰富智慧的一半，超过我所听见的传闻。
2CHR|9|7|你的人是有福的！你这些常侍立在你面前、听你智慧话的仆人是有福的！
2CHR|9|8|耶和华－你的上帝是应当称颂的！他喜爱你，使你坐他的王位，为耶和华－你的上帝作王；因为你的上帝爱 以色列 ，要永远坚立它，所以立你作他们的王，使你秉公行义。”
2CHR|9|9|于是 示巴 女王把一百二十他连得金子、极多的香料和宝石送给 所罗门 王；从来没有像 示巴 女王送给 所罗门 王那么多的香料。
2CHR|9|10|希兰 的仆人和 所罗门 的仆人也从 俄斐 运了金子来，又运了檀香木和宝石来。
2CHR|9|11|王用檀香木为耶和华的殿和王宫做阶梯，又为歌唱的人做琴瑟； 犹大 地从来没有见过这样的。
2CHR|9|12|所罗门 王除了回赠 示巴 女王所带来的，凡她所提出的一切要求， 所罗门 王都送给她。于是女王和她臣仆转回，到本国去了。
2CHR|9|13|所罗门 每年所得的金子，重六百六十六他连得，
2CHR|9|14|另外还有从商人和贸易所收到的，以及 阿拉伯 诸王和各地的省长进贡给 所罗门 的金银。
2CHR|9|15|所罗门 王用锤出来的金子打成二百面盾牌，每面盾牌用六百舍客勒锤出来的金子；
2CHR|9|16|又用锤出来的金子打成三百面小盾牌，每面小盾牌用三百舍客勒金子。王把它们放在 黎巴嫩林宫 里。
2CHR|9|17|王又制造一个大的象牙宝座，包上纯金。
2CHR|9|18|宝座有六层台阶，又有金脚凳，与宝座相连。座位之处两旁有扶手，靠近扶手有两只狮子站立。
2CHR|9|19|六层台阶上有十二只狮子站立，分站左边和右边；任何国度都没有这样做的。
2CHR|9|20|所罗门 王一切的饮器都是金的， 黎巴嫩林宫 里所有的器皿都是纯金的。在 所罗门 的日子，银子算不了什么。
2CHR|9|21|因王的船只与 希兰 的仆人一同往 他施 去， 他施 船只每三年一次把金、银、象牙、猿猴、孔雀 运回来。
2CHR|9|22|所罗门 王的财宝与智慧胜过地上的众王。
2CHR|9|23|地上的众王都求见 所罗门 的面，要听上帝放在他心里的智慧。
2CHR|9|24|他们各带贡物，就是银器、金器、衣服、兵器、香料、马、骡子，每年都有一定的数量。
2CHR|9|25|所罗门 拥有给战车和马用的四千个棚子，还有一万二千名骑兵，安置在屯车城，在 耶路撒冷 的王那里。
2CHR|9|26|所罗门 统管诸王，从 大河 到 非利士 人的地，直到 埃及 的边界。
2CHR|9|27|王在 耶路撒冷 使银子多如石头，香柏木多如 谢非拉 的桑树。
2CHR|9|28|有人从 埃及 和各国为 所罗门 把马匹运来。
2CHR|9|29|所罗门 其余的事，自始至终，不都写在 拿单 先知的书上和 示罗 人 亚希雅 的《预言书》上，以及 易多 先见论 尼八 儿子 耶罗波安 的《默示书》上吗？
2CHR|9|30|所罗门 在 耶路撒冷 作全 以色列 的王四十年。
2CHR|9|31|所罗门 与他祖先同睡，葬在他父亲 大卫 的城里，他儿子 罗波安 接续他作王。
2CHR|10|1|罗波安 往 示剑 去，因 以色列 众人都到了 示剑 ，要立他作王。
2CHR|10|2|尼八 的儿子 耶罗波安 先前躲避 所罗门 王，逃往 埃及 ，住在那里；他听见这事，就从 埃及 回来。
2CHR|10|3|以色列 人派人去请他来。 耶罗波安 就和 以色列 众人来，与 罗波安 谈话，说：
2CHR|10|4|“你父亲使我们负重轭，现在求你减轻你父亲所加给我们的苦工和重轭，我们就服事你。”
2CHR|10|5|罗波安 对他们说：“过三天再来见我吧！”百姓就走了。
2CHR|10|6|罗波安 的父亲 所罗门 在世的时候，有侍立在他面前的长者， 罗波安 王和他们商议，说：“你们出个主意，好把话带回给这百姓。”
2CHR|10|7|他们对他说：“王若恩待这百姓，使他们喜悦，跟他们说好话，他们就永远作王的仆人了。”
2CHR|10|8|王不采纳长者给他出的主意，却和那些与他一同长大、在他面前侍立的年轻人商议。
2CHR|10|9|他对他们说：“这百姓对我说：‘你父亲使我们负重轭，求你减轻一些。’你们出个什么主意，我们好把话带回给他们。”
2CHR|10|10|那些与他一同长大的年轻人对他说：“这些百姓对王说：‘你父亲使我们负重轭，求你给我们减轻一些。’王要对他们如此说：‘我的小指头比我父亲的腰还粗呢！
2CHR|10|11|我父亲使你们负重轭，现在我必使你们负更重的轭！我父亲用鞭子惩罚你们，我却要用蝎子！’”
2CHR|10|12|耶罗波安 和众百姓遵照王所说“你们第三天再来见我”的话，第三天来到 罗波安 那里。
2CHR|10|13|王严厉地回答他们。 罗波安 王不采纳长者所出的主意，
2CHR|10|14|却照着年轻人所出的主意对他们说：“我 使你们负重轭，我必使你们负更重的轭！我父亲用鞭子惩罚你们，我却要用蝎子！”
2CHR|10|15|王不依从百姓，因这事件是出于上帝，为要应验耶和华藉 示罗 人 亚希雅 对 尼八 的儿子 耶罗波安 所说的话。
2CHR|10|16|以色列 众人见王不依从他们，百姓就回覆王说： “我们在 大卫 中有什么分呢？ 我们在 耶西 的儿子中没有产业！ 以色列 啊，各回自己的帐棚去吧！ 大卫 啊，现在你顾自己的家吧！” 于是， 以色列 众人都回自己的帐棚去了；
2CHR|10|17|至于住 犹大 城镇的 以色列 人， 罗波安 仍作他们的王。
2CHR|10|18|罗波安 王派监管劳役的 哈多兰 去， 以色列 人用石头打他，他就死了。 罗波安 王急忙上车，逃回 耶路撒冷 去了。
2CHR|10|19|这样， 以色列 背叛 大卫 家，直到今日。
2CHR|11|1|罗波安 来到 耶路撒冷 ，召集 犹大 家和 便雅悯 家，共十八万人，都是精选的战士，要与 以色列 争战，好将国夺回再归自己。
2CHR|11|2|但耶和华的话临到神人 示玛雅 ，说：
2CHR|11|3|“你去告诉 所罗门 的儿子 犹大 王 罗波安 和住 犹大 、 便雅悯 的 以色列 众人，说：
2CHR|11|4|‘耶和华如此说：你们不可上去与你们的弟兄争战。各自回家去吧！因为这事是出于我。’”众人就听从耶和华的话回去，不去与 耶罗波安 争战。
2CHR|11|5|罗波安 住在 耶路撒冷 ，在 犹大 为防御修筑城镇，
2CHR|11|6|他修筑 伯利恒 、 以坦 、 提哥亚 、
2CHR|11|7|伯．夙 、 梭哥 、 亚杜兰 、
2CHR|11|8|迦特 、 玛利沙 、 西弗 、
2CHR|11|9|亚多莱音 、 拉吉 、 亚西加 、
2CHR|11|10|琐拉 、 亚雅仑 、 希伯仑 。这都是 犹大 和 便雅悯 的坚固城。
2CHR|11|11|罗波安 又巩固这些堡垒，在其中安置军官，储备粮食、油和酒。
2CHR|11|12|他在各城里预备盾牌和枪，使城极其坚固。 犹大 和 便雅悯 都归了他。
2CHR|11|13|全 以色列 的祭司和 利未 人都从四方来归 罗波安 。
2CHR|11|14|利未 人放弃他们的郊野和产业，来到 犹大 与 耶路撒冷 ，因为 耶罗波安 和他的儿子拒绝他们，不许他们担任祭司事奉耶和华。
2CHR|11|15|耶罗波安 为丘坛，为山羊鬼魔，为自己所造的牛犊设立祭司。
2CHR|11|16|以色列 各支派中，凡立定心意寻求耶和华－ 以色列 上帝的，都随从 利未 人来到 耶路撒冷 献祭给耶和华－他们列祖的上帝。
2CHR|11|17|这就巩固了 犹大 王国，使 所罗门 的儿子 罗波安 强盛三年，因为这三年他们遵行 大卫 和 所罗门 的道。
2CHR|11|18|罗波安 娶 大卫 儿子 耶利末 的女儿 玛哈拉 为妻，又娶 耶西 儿子 以利押 的女儿 亚比孩 为妻，
2CHR|11|19|从她生了几个儿子，就是 耶乌施 、 示玛利雅 和 撒罕 。
2CHR|11|20|后来他又娶 押沙龙 的女儿 玛迦 ，从她生了 亚比雅 、 亚太 、 细撒 和 示罗密 。
2CHR|11|21|罗波安 有十八个妻和六十个妾，生了二十八个儿子，六十个女儿；他却爱 押沙龙 的女儿 玛迦 ，过于爱其他的妻妾。
2CHR|11|22|罗波安 立 玛迦 的儿子 亚比雅 作太子，在他兄弟中为首，因为要立他作王。
2CHR|11|23|罗波安 办事精明，把他众儿子分散在 犹大 和 便雅悯 全地各坚固城里，赐他们大量的粮食，又给他们娶许多妻子。
2CHR|12|1|罗波安 的王国稳固，他强盛的时候就离弃耶和华的律法，全 以色列 都跟从他。
2CHR|12|2|罗波安 王第五年， 埃及 王 示撒 上来攻打 耶路撒冷 ，因为他们背叛了耶和华。
2CHR|12|3|示撒 带着一千二百辆战车，六万名骑兵，以及跟随他从 埃及 出来的 路比 人、 苏基 人和 古实 人的军队，多得不可胜数。
2CHR|12|4|他攻取了 犹大 的坚固城，来到 耶路撒冷 。
2CHR|12|5|那时， 犹大 的领袖因为 示撒 的缘故聚集在 耶路撒冷 ，有先知 示玛雅 去见 罗波安 和众领袖，对他们说：“耶和华如此说：‘你们离弃了我，所以我也离弃你们，把你们交在 示撒 手里。’”
2CHR|12|6|于是 以色列 的领袖和王都谦卑说：“耶和华是公义的。”
2CHR|12|7|耶和华见他们谦卑，耶和华的话就临到 示玛雅 ，说：“他们既谦卑，我必不灭绝他们；我要使他们暂时得拯救，不藉着 示撒 的手将我的怒气倒在 耶路撒冷 。
2CHR|12|8|然而他们必作 示撒 的仆人，好叫他们知道，服事我与服事地上邦国有何分别。”
2CHR|12|9|于是， 埃及 王 示撒 上来攻取 耶路撒冷 ，夺了耶和华殿和王宫里的宝物，尽都带走，又夺走 所罗门 制造的金盾牌。
2CHR|12|10|罗波安 王制造铜盾牌代替那些金盾牌，交给看守王宫宫门的护卫长看管。
2CHR|12|11|每逢王进耶和华的殿，护卫兵就来，举起这些盾牌；随后仍将盾牌送回护卫室。
2CHR|12|12|王谦卑的时候，耶和华的怒气就转消了，不全然灭尽，并且在 犹大 中，情况也有好转。
2CHR|12|13|罗波安 王自强，在 耶路撒冷 作王。他登基的时候年四十一岁，在 耶路撒冷 ，就是耶和华从 以色列 众支派中所选择立他名的城，作王十七年。 罗波安 的母亲名叫 拿玛 ，是 亚扪 人。
2CHR|12|14|罗波安 行恶，因他没有立定心意寻求耶和华。
2CHR|12|15|罗波安 的事迹，自始至终不都写在 示玛雅 先知和 易多 先见的《史记》上吗？ 罗波安 与 耶罗波安 时常交战。
2CHR|12|16|罗波安 与他祖先同睡，葬在 大卫城 ，他的儿子 亚比雅 接续他作王。
2CHR|13|1|耶罗波安 王十八年， 亚比雅 登基作 犹大 王，
2CHR|13|2|在 耶路撒冷 作王三年。他母亲名叫 米该亚 ，是 基比亚 人 乌列 的女儿 。 亚比雅 常与 耶罗波安 交战。
2CHR|13|3|有一次 亚比雅 率领四十万精选的士兵出战，他们都是勇敢的战士； 耶罗波安 也率领八十万精选的大能勇士，迎着 亚比雅 摆阵。
2CHR|13|4|亚比雅 站在 以法莲 山区中的 洗玛脸山 上，说：“ 耶罗波安 和 以色列 众人哪，要听我说！
2CHR|13|5|耶和华－ 以色列 的上帝曾立盐约，将 以色列 国永远赐给 大卫 和他的子孙，你们不知道吗？
2CHR|13|6|但 大卫 儿子 所罗门 的臣仆、 尼八 的儿子 耶罗波安 起来背叛他的主人。
2CHR|13|7|有些无赖的歹徒聚集跟从他，逞强攻击 所罗门 的儿子 罗波安 ；那时 罗波安 还年轻，心志软弱，不能抵挡他们。
2CHR|13|8|“现在你们说要抗拒 大卫 子孙手下所治理的耶和华的国，你们的人数众多，你们那里又有 耶罗波安 为你们所造当作神明的金牛犊。
2CHR|13|9|你们不是驱逐耶和华的祭司 亚伦 的后裔和 利未 人吗？不是照着外邦人的恶俗为自己立祭司吗？无论何人牵一头公牛犊、七只公绵羊将自己分别出来，就可作虚无神明的祭司。
2CHR|13|10|至于我们，耶和华是我们的上帝，我们并没有离弃他。我们有事奉耶和华的祭司，都是 亚伦 的后裔，并有 利未 人各尽其职。
2CHR|13|11|他们每日早晚向耶和华献燔祭，烧芬芳的香，又在纯金的 供桌上摆供饼，每晚点燃金灯台上的灯盏，因为我们遵守耶和华－我们上帝的命令，但你们却离弃了他。
2CHR|13|12|看哪，率领我们的是上帝，又有他的祭司拿号向你们吹出响声。 以色列 人哪，不要与耶和华－你们列祖的上帝争战，因你们必不能得胜。”
2CHR|13|13|耶罗波安 却在 犹大 人的后头设伏兵。这样， 以色列 人在 犹大 人的前头，伏兵在 犹大 人的后头。
2CHR|13|14|犹大 人转过来，看哪，前后都有战事，就呼求耶和华，祭司也吹号。
2CHR|13|15|于是 犹大 人呐喊。 犹大 人呐喊的时候，上帝就击打 耶罗波安 和 以色列 众人，使他们败在 亚比雅 与 犹大 人面前。
2CHR|13|16|以色列 人在 犹大 人面前逃跑，上帝将他们交在 犹大 人手里。
2CHR|13|17|亚比雅 和他的军兵大大击杀 以色列 人， 以色列 人被杀仆倒的精兵有五十万。
2CHR|13|18|那时， 以色列 人被制伏了。 犹大 人得胜，因为他们倚靠耶和华－他们列祖的上帝。
2CHR|13|19|亚比雅 追赶 耶罗波安 ，攻取了他的几座城，就是 伯特利 和所属的乡镇 ， 耶沙拿 和所属的乡镇， 以法拉音 和所属的乡镇。
2CHR|13|20|亚比雅 在世的时候， 耶罗波安 不再强盛；耶和华击打他，他就死了。
2CHR|13|21|亚比雅 却渐渐强盛。他娶了十四个妻妾，生了二十二个儿子，十六个女儿。
2CHR|13|22|亚比雅 其余的事和他的言行都写在 易多 先知的评传上。
2CHR|14|1|亚比雅 与他祖先同睡，葬在 大卫城 ，他的儿子 亚撒 接续他作王。 亚撒 在位期间，国中太平十年。
2CHR|14|2|亚撒 行耶和华－他上帝眼中看为善为正的事，
2CHR|14|3|除掉外邦的祭坛和丘坛，打碎柱像，砍下 亚舍拉 ，
2CHR|14|4|吩咐 犹大 人寻求耶和华－他们列祖的上帝，遵行他的律法和诫命，
2CHR|14|5|又在 犹大 各城镇除掉丘坛和香坛。在他治理下，国中太平。
2CHR|14|6|他在 犹大 建造了几座坚固城。那些年间，国中太平，没有战争，因为耶和华赐他平安。
2CHR|14|7|他对 犹大 人说：“我们要建造这些城镇，四围筑墙，盖城楼，安门，做闩；地仍属于我们，因为我们寻求耶和华－我们的上帝；我们寻求他，他就赐我们四境平安。”于是他们建造城镇，诸事亨通。
2CHR|14|8|亚撒 的军兵，出自 犹大 拿盾牌拿枪的三十万人，出自 便雅悯 拿小盾牌拉弓的二十八万人；这些全都是大能的勇士。
2CHR|14|9|古实 人 谢拉 率领一百万军兵，三百辆战车，出来攻击 犹大 人，到了 玛利沙 。
2CHR|14|10|亚撒 出去迎战，在 玛利沙 的 洗法谷 彼此摆阵。
2CHR|14|11|亚撒 呼求耶和华－他的上帝说：“耶和华啊，在强弱之间，惟有你能帮助。耶和华－我们的上帝啊，求你帮助我们，因为我们仰赖你，奉你的名来抵挡这大军。耶和华啊，你是我们的上帝，不要让人胜过你。”
2CHR|14|12|于是耶和华击打 古实 人，使他们败在 亚撒 和 犹大 人面前， 古实 人就逃跑了。
2CHR|14|13|亚撒 和跟随他的军兵追赶他们，直到 基拉耳 。 古实 人被杀的很多，无法复原，因为他们在耶和华与他军兵面前被击溃。 犹大 人夺了许多财物，
2CHR|14|14|又攻打 基拉耳 四围一切的城镇；城中的人都惧怕耶和华。 犹大 人掳掠了一切的城镇，因其中的财物很多，
2CHR|14|15|又毁坏了群畜的圈，夺取许多的羊和骆驼，就回 耶路撒冷 去了。
2CHR|15|1|上帝的灵临到 俄德 的儿子 亚撒利雅 。
2CHR|15|2|他出来迎接 亚撒 ，对他说：“ 亚撒 ， 犹大 和 便雅悯 众人哪，要听我说：你们若顺从耶和华，耶和华必与你们同在；你们若寻求他，就必寻见；你们若离弃他，他必离弃你们。
2CHR|15|3|以色列 人不信真神，没有训诲的祭司，也没有律法，已经许多日子了。
2CHR|15|4|但他们在急难的时候归向耶和华－ 以色列 的上帝，寻求他，他就被他们寻见。
2CHR|15|5|那时，出入的人不得平安，各地的居民都遭大乱；
2CHR|15|6|他们被破坏殆尽，这国攻击那国，这城攻击那城，因为上帝用各样灾难扰乱他们。
2CHR|15|7|现在你们要刚强，不要手软，因你们所行的必得赏赐。”
2CHR|15|8|亚撒 听见这些话和 俄德 先知的预言，就壮起胆来，在 犹大 和 便雅悯 全地，以及 以法莲 山区所夺的各城，把其中的可憎之物尽都除掉，又在耶和华殿的走廊前重新修筑耶和华的坛。
2CHR|15|9|他又召集 犹大 和 便雅悯 众人，以及他们中间寄居的 以法莲 人、 玛拿西 人、 西缅 人。有许多 以色列 人归顺 亚撒 ，因为他们看见耶和华－他的上帝与他同在。
2CHR|15|10|亚撒 作王第十五年三月，他们都聚集在 耶路撒冷 。
2CHR|15|11|那日他们从所取的掳物中，将七百头牛和七千只羊献给耶和华。
2CHR|15|12|他们立约，要尽心尽性寻求耶和华－他们列祖的上帝。
2CHR|15|13|凡不寻求耶和华－ 以色列 上帝的，无论大小、男女，必被处死。
2CHR|15|14|他们就大声欢呼，吹号吹角，向耶和华起誓。
2CHR|15|15|犹大 众人为所起的誓欢喜，因他们尽心起誓，尽意寻求耶和华，耶和华就被他们寻见，且赐他们四境平安。
2CHR|15|16|亚撒 王甚至废了他祖母 玛迦 太后的位，因 玛迦 造了可憎的 亚舍拉 。 亚撒 砍下她的偶像，捣得粉碎，在 汲沦溪 边烧了，
2CHR|15|17|只是丘坛还没有从 以色列 中废去，然而 亚撒 一生有纯正的心。
2CHR|15|18|亚撒 将他父亲所分别为圣与自己所分别为圣的金银和器皿都奉到上帝的殿里。
2CHR|15|19|亚撒 作王直到第三十五年，都没有战事。
2CHR|16|1|亚撒 作王第三十六年， 以色列 王 巴沙 上来攻击 犹大 ，修筑 拉玛 ，不许人从 犹大 王 亚撒 那里出入。
2CHR|16|2|于是 亚撒 从耶和华殿和王宫的府库里拿出金银来，送给住在 大马士革 的 亚兰 王 便．哈达 ，说：
2CHR|16|3|“你父曾与我父立约，我与你也要这样立约。看哪，我把金银送给你，请你废掉你与 以色列 王 巴沙 所立的约，使他从我这里撤退。”
2CHR|16|4|便．哈达 听从了 亚撒 王，就派遣他的军官去攻打 以色列 的城镇。他们攻下了 以云 、 但 、 亚伯．玛音 和 拿弗他利 一切的储货城。
2CHR|16|5|巴沙 听见了，就停工不修筑 拉玛 ，任由他的工程停止。
2CHR|16|6|于是 亚撒 王率领 犹大 众人，运走 巴沙 修筑 拉玛 所用的石头和木料，用以修筑 迦巴 和 米斯巴 。
2CHR|16|7|那时， 哈拿尼 先见来见 犹大 王 亚撒 ，对他说：“因你仰赖 亚兰 王，没有仰赖耶和华－你的上帝，所以 亚兰 王的军兵逃脱了你的手。
2CHR|16|8|古实 人和 路比 人的军队不是非常强大吗？他们的战车骑兵不是极多吗？只因你仰赖耶和华，他就将他们交在你手里。
2CHR|16|9|因为耶和华的眼目遍察全地，要坚固向他存纯正之心的人。你在这事上行得愚昧；因此，以后你必有战争。”
2CHR|16|10|亚撒 恼恨先见，为了这事向他发怒，将他囚在监里。那时 亚撒 也虐待一些百姓。
2CHR|16|11|亚撒 自始至终的事迹，看哪，都写在《犹大和以色列诸王记》上。
2CHR|16|12|亚撒 作王三十九年的时候患了脚疾，非常严重。他生病的时候没有求耶和华，只求医生。
2CHR|16|13|他作王四十一年死了，与他祖先同睡，
2CHR|16|14|葬在 大卫城 自己所凿的坟墓里。人把他放在床上，床上堆满各样馨香的香料，就是按做香的作法调和的香料，又为他生一堆大火志哀。
2CHR|17|1|亚撒 的儿子 约沙法 接续他作王，奋勇自强，防备 以色列 。
2CHR|17|2|他安置军兵在 犹大 一切坚固城里，又安置驻军在 犹大 地和他父亲 亚撒 所得 以法莲 的城镇中。
2CHR|17|3|耶和华与 约沙法 同在，因为他行他祖先 大卫 从前所行的道，不去寻求诸 巴力 ，
2CHR|17|4|只寻求他父亲的上帝，遵行他的诫命，不效法 以色列 人的行为。
2CHR|17|5|所以耶和华坚定 约沙法 手中的国， 犹大 众人给他进贡； 约沙法 大有财富和尊荣。
2CHR|17|6|他乐意遵行耶和华的道，并且从 犹大 再次除掉一切丘坛和 亚舍拉 。
2CHR|17|7|他作王第三年，差遣官员 便．亥伊勒 、 俄巴底 、 撒迦利雅 、 拿坦业 、 米该亚 往 犹大 各城去教导百姓。
2CHR|17|8|跟他们一同去的有 利未 人 示玛雅 、 尼探雅 、 西巴第雅 、 亚撒黑 、 示米拉末 、 约拿单 、 亚多尼雅 、 多比雅 、 驼．巴多尼雅 ；跟他们一同的又有 以利沙玛 和 约兰 二位祭司。
2CHR|17|9|他们在 犹大 教导，带着耶和华的律法书，走遍 犹大 各城教导百姓。
2CHR|17|10|犹大 四围地上的邦国都惧怕耶和华，不敢与 约沙法 争战。
2CHR|17|11|有些 非利士 人送礼物，进贡银子给 约沙法 。 阿拉伯 人也送他七千七百只公绵羊，七千七百只公山羊。
2CHR|17|12|约沙法 日渐强大，他在 犹大 建造堡垒和储货城。
2CHR|17|13|他在 犹大 城镇中有许多工程，在 耶路撒冷 又有战士，就是大能的勇士。
2CHR|17|14|他们按着父家的数目如下： 犹大 族的千夫长以 押拿 为首，率领三十万大能的勇士；
2CHR|17|15|其次是 约哈难 千夫长，率领二十八万；
2CHR|17|16|其次是 细基利 的儿子 亚玛斯雅 ，他是一个自愿奉献给耶和华的人，率领二十万大能的勇士。
2CHR|17|17|便雅悯 族有大能的勇士 以利雅大 ，率领二十万拿弓箭和盾牌的人；
2CHR|17|18|其次是 约萨拔 ，率领十八万预备打仗的人。
2CHR|17|19|这些都是伺候王的，还有王在全 犹大 的坚固城所安置的不在其内。
2CHR|18|1|约沙法 大有财富和尊荣，他与 亚哈 结亲。
2CHR|18|2|过了几年，他下到 撒玛利亚 去见 亚哈 ； 亚哈 为他和跟从他的人宰了许多牛羊，劝他一同上去攻打 基列 的 拉末 。
2CHR|18|3|以色列 王 亚哈 问 犹大 王 约沙法 说：“你肯同我去攻打 基列 的 拉末 吗？”他回答说：“你我不分彼此，我的军队就是你的军队，我们必与你一同去争战。”
2CHR|18|4|约沙法 对 以色列 王说：“请你先求问耶和华的话。”
2CHR|18|5|于是 以色列 王召集先知四百人，问他们说：“我可以上去攻打 基列 的 拉末 吗？还是不要上去呢？”他们说：“可以上去，因为上帝必将那城交在王的手里。”
2CHR|18|6|约沙法 说：“这里还有没有耶和华的先知，我们好求问他呢？”
2CHR|18|7|以色列 王对 约沙法 说：“还有一个人，是 音拉 的儿子 米该雅 ，我们可以托他求问耶和华。只是我真的很恨他，因为他对我说预言，从不说吉言，总是说凶信。” 约沙法 说：“请王不要这么说。”
2CHR|18|8|以色列 王就召了一个官员来，说：“你快去，把 音拉 的儿子 米该雅 召来。”
2CHR|18|9|以色列 王和 犹大 王 约沙法 在 撒玛利亚 城门前的禾场，各穿朝服，坐在宝座上，所有的先知都在他们面前说预言。
2CHR|18|10|基拿拿 的儿子 西底家 为自己造了铁角，说：“耶和华如此说：‘你要用这些角抵触 亚兰 人，直到将他们灭尽。’”
2CHR|18|11|所有的先知也都这样预言说：“可以上 基列 的 拉末 去，必然得胜，因为耶和华必将那城交在王的手中。”
2CHR|18|12|那去召 米该雅 的使者对他说：“看哪，众先知都异口同声向王说吉言，你也跟他们说一样的话，说吉言吧！”
2CHR|18|13|米该雅 说：“我指着永生的耶和华起誓，我的上帝说什么，我就说什么。”
2CHR|18|14|米该雅 来到王那里，王问他：“ 米该雅 啊，我们可以上去攻打 基列 的 拉末 吗？还是不要上去呢？”他说：“可以上去，必然得胜，敌人必交在你们手里。”
2CHR|18|15|王对他说：“我要你发誓多少次，你才会奉耶和华的名向我说实话呢？”
2CHR|18|16|米该雅 说：“我看见 以色列 众人散布在山上，如同没有牧人的羊群一般。耶和华说：‘这些人没有主人，他们可以平安地各自回家去。’”
2CHR|18|17|以色列 王对 约沙法 说：“我岂没有告诉你，这人对我说预言，从不说吉言，只说凶信吗？”
2CHR|18|18|米该雅 说：“因此你们要听耶和华的话！我看见耶和华坐在宝座上，天上的万军侍立在他左右。
2CHR|18|19|耶和华 说：‘谁去引诱 以色列 王 亚哈 上 基列 的 拉末 去阵亡呢？’这个这样说，那个那样说。
2CHR|18|20|随后有一个灵出来，站在耶和华面前，说：‘我去引诱他。’耶和华问他：‘用什么方法呢？’
2CHR|18|21|他说：‘我要出去，在他众先知的口中成为谎言的灵。’耶和华说：‘这样，你去引诱他，必能成功。你出去，照样做吧！’
2CHR|18|22|现在，看哪，耶和华使谎言的灵入了你的这些先知的口，并且耶和华已经宣告要降祸于你。”
2CHR|18|23|基拿拿 的儿子 西底家 前来打 米该雅 一巴掌，说：“耶和华的灵从哪里离开我向你说话呢？”
2CHR|18|24|米该雅 说：“看哪，你进入严密的内室躲藏的那日，就必看见。”
2CHR|18|25|以色列 王说：“把 米该雅 带走，交回给 亚们 市长和 约阿施 王子。
2CHR|18|26|你们要说：‘王如此说：把这个人关在监狱里，使他受苦，吃不饱喝不足，直等到我平安回来。’”
2CHR|18|27|米该雅 说：“你若真的能平安回来，那就是耶和华没有藉我说话了。”他又说：“众百姓啊，你们都要听！”
2CHR|18|28|以色列 王和 犹大 王 约沙法 上 基列 的 拉末 去。
2CHR|18|29|以色列 王对 约沙法 说：“我要改装上阵，你可以仍穿王服。”于是 以色列 王改装，他们上阵去了。
2CHR|18|30|亚兰 王吩咐他的战车长说：“你们不要与他们的大将或小兵交战，只要单单攻击 以色列 王。”
2CHR|18|31|那些战车长看见 约沙法 就说：“这一定是 以色列 王！”他们转过去与他交战。 约沙法 一呼喊，耶和华就帮助他，上帝使他们转离他。
2CHR|18|32|战车长见他不是 以色列 王，就转身不追他了。
2CHR|18|33|有一人开弓，并不知情，箭恰巧射入 以色列 王铠甲的缝里。王对驾车的说：“我受重伤了，你掉过车来，载我离开战场！”
2CHR|18|34|那日，战况越来越猛， 以色列 王勉强站在战车上，面对 亚兰 人，直到傍晚。日落的时候，王就死了。
2CHR|19|1|犹大 王 约沙法 平安回 耶路撒冷 ，到自己的宫里。
2CHR|19|2|哈拿尼 的儿子 耶户 先见出来迎接 约沙法 王，对他说：“你怎么可以帮助恶人，爱那恨耶和华的人呢？因此耶和华的愤怒临到你了。
2CHR|19|3|然而你还有善行，因你从国中除掉 亚舍拉 ，立定心意寻求上帝。”
2CHR|19|4|约沙法 住在 耶路撒冷 ，以后又出巡民间，从 别是巴 直到 以法莲 山区，引导百姓归向耶和华－他们列祖的上帝。
2CHR|19|5|他在国中，在 犹大 一切坚固城设立审判官，各城都是如此。
2CHR|19|6|他对审判官说：“你们应当谨慎所做的事，因为你们审判不是为人，而是为耶和华。在审判的事上，他必与你们同在。
2CHR|19|7|现在，你们应当敬畏耶和华，谨慎办事，因为耶和华－我们的上帝没有不义，不看人的情面，也不受贿赂。”
2CHR|19|8|约沙法 从 利未 人和祭司，以及 以色列 族长中，也委派人在 耶路撒冷 为耶和华施行审判，为 耶路撒冷 的居民听讼断案 。
2CHR|19|9|约沙法 吩咐他们说：“你们当这样，以敬畏耶和华、诚实和纯正的心办事。
2CHR|19|10|你们住在各城的弟兄，若有争讼的案件呈到你们这里，或为流血，或犯律法、诫命、律例、典章，你们要警戒他们，免得他们得罪耶和华，以致愤怒临到你们和你们的弟兄；你们当这样行，就没有罪了。
2CHR|19|11|看哪，凡属耶和华的事，有 亚玛利雅 祭司长管理你们；凡属王的事，有 犹大 家的领袖 以实玛利 的儿子 西巴第雅 管理你们；在你们面前有 利未 人作官长。你们应当壮胆办事，愿耶和华与善人同在。”
2CHR|20|1|此后， 摩押 人和 亚扪 人，连同一些 米乌尼 人 来攻击 约沙法 。
2CHR|20|2|有人来报告 约沙法 说：“从海的那边， 以东 有大军来攻击你，看哪，他们在 哈洗逊．他玛 ，就是 隐．基底 。”
2CHR|20|3|约沙法 惧怕，就定意寻求耶和华，在全 犹大 宣告禁食。
2CHR|20|4|于是 犹大 人聚集，求耶和华帮助，甚至他们从 犹大 各城前来寻求耶和华。
2CHR|20|5|约沙法 站在 犹大 和 耶路撒冷 的会众中，在耶和华殿新的院子前，
2CHR|20|6|说：“耶和华－我们列祖的上帝啊，你不是天上的上帝吗？你不是万邦万国的主宰吗？在你手中有大能大力，无人能抵挡你。
2CHR|20|7|我们的上帝啊，你不是曾在你百姓 以色列 面前驱逐这地的居民，将这地赐给你朋友 亚伯拉罕 的后裔永远为业吗？
2CHR|20|8|他们住在这地，又为你的名建造圣所，说：
2CHR|20|9|‘若有祸患临到我们，或刀兵的惩罚，或瘟疫饥荒，我们在急难的时候，站在这殿前向你呼求，你必垂听并且拯救，因为你的名在这殿里。’
2CHR|20|10|现在，看哪， 以色列 人出 埃及 地的时候，你不容许 以色列 人侵犯 亚扪 人、 摩押 人和 西珥山 人， 以色列 人就离开他们，不灭绝他们。
2CHR|20|11|看哪，他们这样回报我们，要来驱逐我们离开你赐给我们为业之地。
2CHR|20|12|我们的上帝啊，你不惩罚他们吗？因为我们无力抵挡这来攻击我们的大军。我们不知道该怎么做，我们的眼目单仰望你。”
2CHR|20|13|犹大 众人和他们的孩童、妻子、儿女都站在耶和华面前。
2CHR|20|14|那时，耶和华的灵在会众中临到 利未 人 亚萨 的后裔 雅哈悉 ，他是 玛探雅 的玄孙， 耶利 的曾孙， 比拿雅 的孙子， 撒迦利雅 的儿子。
2CHR|20|15|他说：“ 犹大 众人、 耶路撒冷 的居民和 约沙法 王啊，你们要留心听，耶和华对你们如此说：‘不要因这大军恐惧惊惶，因为胜败不在乎你们，而是在乎上帝。
2CHR|20|16|明日你们要下去迎敌；看哪，他们从 洗斯坡 上来，你们必在 耶鲁伊勒 旷野前的谷口遇见他们。
2CHR|20|17|犹大 和 耶路撒冷 人哪，这次你们不要争战，要摆阵站着，看耶和华为你们施行拯救。不要恐惧，也不要惊惶。明日当出去迎敌，因为耶和华与你们同在。’”
2CHR|20|18|约沙法 屈身，脸伏于地， 犹大 众人和 耶路撒冷 的居民也俯伏在耶和华面前，敬拜耶和华。
2CHR|20|19|哥辖 子孙和 可拉 子孙的 利未 人都起来，用极大的声音赞美耶和华－ 以色列 的上帝。
2CHR|20|20|清晨，众人早起往 提哥亚 的旷野去。出去的时候， 约沙法 站着说：“ 犹大 人和 耶路撒冷 的居民哪，要听我说：信靠耶和华－你们的上帝就必站立得稳；信赖他的先知就必亨通。”
2CHR|20|21|约沙法 与百姓商议，就设立歌唱的人，颂赞耶和华，使他们穿上圣洁的礼服，走在军队前赞美耶和华： “当称谢耶和华， 因他的慈爱永远长存！”
2CHR|20|22|他们开始唱歌赞美的时候，耶和华派伏兵击杀那来攻击 犹大 的 亚扪 人、 摩押 人和 西珥山 人，他们就被打败了。
2CHR|20|23|亚扪 人和 摩押 人起来，击杀住 西珥山 的人，把他们灭尽；灭尽住 西珥山 的人之后，他们又彼此自相击杀。
2CHR|20|24|犹大 人来到旷野的了望楼，向那大军观看，看哪，遍地都是尸体，没有一个逃脱的。
2CHR|20|25|约沙法 和他的百姓就来收取掠物，找到许多牲畜 、财物、衣服 和珍宝。他们取掠物归为己有，直到无法携带；因为掠物太多，他们足足收取了三日。
2CHR|20|26|第四日，众人聚集在 比拉迦谷 ，在那里称颂耶和华；因此那地方名叫 比拉迦谷 ，直到今日。
2CHR|20|27|在 约沙法 率领下， 犹大 人和 耶路撒冷 人都欢欢喜喜地回 耶路撒冷 ，耶和华使他们因战胜仇敌而喜乐。
2CHR|20|28|他们弹琴、鼓瑟、吹号来到 耶路撒冷 ，进了耶和华的殿。
2CHR|20|29|地上所有的邦国听见耶和华打败 以色列 的仇敌，就都惧怕上帝。
2CHR|20|30|这样， 约沙法 的国得享太平，因为上帝赐他四境平安。
2CHR|20|31|约沙法 作 犹大 王，登基的时候年三十五岁，在 耶路撒冷 作王二十五年。他母亲名叫 阿苏巴 ，是 示利希 的女儿。
2CHR|20|32|约沙法 效法他父亲 亚撒 所行的道，不偏离左右，行耶和华眼中看为正的事。
2CHR|20|33|只是丘坛还没有废去，百姓也没有立定心意归向他们列祖的上帝。
2CHR|20|34|约沙法 其余的事，看哪，自始至终都写在 哈拿尼 的儿子 耶户 的书上，这些事也记载在《以色列诸王记》上。
2CHR|20|35|此后， 犹大 王 约沙法 与 以色列 王 亚哈谢 结盟； 亚哈谢 多行恶事。
2CHR|20|36|他们合伙造船要往 他施 去，就在 以旬．迦别 造船。
2CHR|20|37|玛利沙 人 多大瓦 的儿子 以利以谢 向 约沙法 预言说：“因你与 亚哈谢 结盟，耶和华必破坏你所造的。”后来那些船果然毁坏，不能往 他施 去了。
2CHR|21|1|约沙法 与他祖先同睡，与他祖先同葬在 大卫城 ，他的儿子 约兰 接续他作王。
2CHR|21|2|约兰 有几个兄弟，就是 约沙法 的儿子 亚撒利雅 、 耶歇 、 撒迦利雅 、 亚撒列夫 、 米迦勒 、 示法提雅 ；这些都是 以色列 王 约沙法 的儿子。
2CHR|21|3|他们的父亲把许多礼物，金银财宝和 犹大 的坚固城赐给他们，却把国赐给 约兰 ，因为他是长子。
2CHR|21|4|约兰 起来治理他父亲的国，奋勇自强，用刀杀了他所有的兄弟和 以色列 的几个领袖。
2CHR|21|5|约兰 登基的时候年三十二岁，在 耶路撒冷 作王八年。
2CHR|21|6|他行 以色列 诸王的道，正如 亚哈 家所行的，因他娶了 亚哈 的女儿为妻，行耶和华眼中看为恶的事。
2CHR|21|7|耶和华却因自己与 大卫 所立的约，不肯灭绝 大卫 的家，要照他所应许的，永远赐灯光给 大卫 和他的子孙。
2CHR|21|8|约兰 在位期间， 以东 背叛，自己立王治理他们，脱离 犹大 的权势。
2CHR|21|9|约兰 就率领他的军官和所有的战车过去。他夜间起来，攻打围困他的 以东 人和战车长。
2CHR|21|10|这样， 以东 背叛，脱离 犹大 的权势，直到今日。那时， 立拿 也背叛了，脱离它的权势，因为 约兰 离弃耶和华－他列祖的上帝。
2CHR|21|11|他又在 犹大 山岭 建造丘坛，使 耶路撒冷 的居民行淫，诱惑 犹大 。
2CHR|21|12|以利亚 先知写信给 约兰 说：“耶和华－你祖先 大卫 的上帝如此说：‘因为你不行你父 约沙法 和 犹大 王 亚撒 的道，
2CHR|21|13|反而行 以色列 诸王的道，使 犹大 和 耶路撒冷 居民行淫，像 亚哈 家行淫一样，又杀了你父家比你好的那些兄弟。
2CHR|21|14|看哪，耶和华必降大灾于你的百姓和你的妻妾、儿女，以及你一切所有的。
2CHR|21|15|至于你，你必患许多的病 ，你的肠子也必生许多的病，日渐沉重，直到肠子坠落下来。’”
2CHR|21|16|耶和华激发 非利士 人和靠近 古实 人的 阿拉伯 人的心来攻击 约兰 。
2CHR|21|17|他们上来攻击 犹大 ，侵入境内，掳掠了王宫里所有的财物和他的妻妾、儿女，除了他的小儿子 约哈斯 之外，没有留下一个儿子。
2CHR|21|18|这一切事以后，耶和华击打 约兰 ，使他的肠子患不能医治的病。
2CHR|21|19|这病缠绵日久，过了二年，肠子坠落下来，他就病重而死。他的百姓没有为他生火志哀，像从前为他祖先生火一样。
2CHR|21|20|约兰 登基的时候年三十二岁，在 耶路撒冷 作王八年。他逝世无人思慕，众人把他葬在 大卫城 ，只是不在列王的坟墓里。
2CHR|22|1|耶路撒冷 的居民立 约兰 的小儿子 亚哈谢 接续他作王，因为跟随 阿拉伯 人来攻营的军兵把 亚哈谢 所有的兄长都杀了； 犹大 王 约兰 的儿子 亚哈谢 就作了王。
2CHR|22|2|亚哈谢 登基的时候年四十二岁 ，在 耶路撒冷 作王一年。他母亲名叫 亚她利雅 ，是 暗利 的孙女。
2CHR|22|3|亚哈谢 也行 亚哈 家的道，因为他母亲给他主谋，使他行恶。
2CHR|22|4|他行耶和华眼中看为恶的事，像 亚哈 家一样；因他父亲死后，他们给他主谋，使他败坏。
2CHR|22|5|他也听从他们的计谋，与 以色列 王 亚哈 的儿子 约兰 同往 基列 的 拉末 去，与 亚兰 王 哈薛 交战。 亚兰 人打伤了 约兰 ，
2CHR|22|6|他回到 耶斯列 ，医治在 拉末 与 亚兰 王 哈薛 打仗时被击打所受的伤。 约兰 的儿子 犹大 王 亚哈谢 因为 亚哈 的儿子 约兰 病了，就下到 耶斯列 看望他。
2CHR|22|7|亚哈谢 去见 约兰 而遇害，这是出乎上帝；因为他一到就同 约兰 出去攻击 宁示 的孙子 耶户 ；这 耶户 是耶和华所膏，使他剪除 亚哈 家的。
2CHR|22|8|耶户 向 亚哈 家施行惩罚的时候，遇见 犹大 的众领袖和 亚哈谢 的侄子们正服事 亚哈谢 ，就把他们都杀了。
2CHR|22|9|亚哈谢 躲在 撒玛利亚 ， 耶户 寻找他，众人把他拿住，送到 耶户 那里，就杀了他。他们把他埋葬，因他们说，他是那尽心寻求耶和华之 约沙法 的儿子。这样， 亚哈谢 的家无力保住国权。
2CHR|22|10|亚哈谢 的母亲 亚她利雅 见她儿子死了，就起来剿灭 犹大 王室所有的后裔。
2CHR|22|11|但王的女儿 约示巴 将 亚哈谢 的儿子 约阿施 从那被杀的王子中偷出来，把他和他的奶妈藏在卧房里。 约示巴 是 约兰 王的女儿， 亚哈谢 的妹妹，祭司 耶何耶大 的妻子。她藏了 约阿施 ，躲避 亚她利雅 ，免受杀害。
2CHR|22|12|亚她利雅 治理这地的时候， 约阿施 和他们一同在上帝殿里藏了六年。
2CHR|23|1|第七年， 耶何耶大 奋勇自强，叫了 耶罗罕 的儿子 亚撒利雅 、 约哈难 的儿子 以实玛利 、 俄备得 的儿子 亚撒利雅 、 亚大雅 的儿子 玛西雅 ，和 细基利 的儿子 以利沙法 等众百夫长，与他们立约。
2CHR|23|2|他们走遍 犹大 ，从 犹大 各城召集 利未 人和 以色列 的众族长到 耶路撒冷 来。
2CHR|23|3|全会众在上帝殿里与王立约。 耶何耶大 对他们说：“看哪，王的儿子必作王，正如耶和华指着 大卫 子孙所应许的。
2CHR|23|4|你们要这样做：在安息日值班的祭司和 利未 人，三分之一要把守各门，
2CHR|23|5|三分之一要在王宫，三分之一要在 根基门 ；众百姓都要在耶和华殿的院内。
2CHR|23|6|除了祭司和供职的 利未 人之外，不准别人进耶和华的殿；只有他们可以进去，因为他们是神圣的。众百姓都要遵守耶和华所吩咐的。
2CHR|23|7|利未 人要手中各拿兵器，四围保护王；凡擅自进殿的，要被处死。王出入的时候，你们当跟随他。”
2CHR|23|8|利未 人和 犹大 众人都照着 耶何耶大 祭司一切所吩咐的去做，各带自己的人，无论安息日值班或不值班的都来，因为 耶何耶大 祭司不许他们下班。
2CHR|23|9|耶何耶大 祭司就把上帝殿里所藏 大卫 王的枪和大小盾牌交给百夫长，
2CHR|23|10|又分派众百姓手中各拿兵器，在祭坛和殿那里，从殿南到殿北，站在王的四围；
2CHR|23|11|他们领 约阿施 出来，给他戴上冠冕，把律法书交给他，立他作王。 耶何耶大 和他的儿子们膏他，他们说：“愿王万岁！”
2CHR|23|12|亚她利雅 听见百姓奔走赞美王的声音，就进耶和华的殿，到百姓那里。
2CHR|23|13|她观看，看哪，王站在殿门的柱旁，百夫长和号手在王旁边，国中的众百姓都欢乐吹号，又有歌唱的人用乐器领人歌唱赞美。 亚她利雅 就撕裂衣服，喊着说：“反了！反了！”
2CHR|23|14|耶何耶大 祭司带领管军兵的百夫长出来，对他们说：“把她从行列之间赶出去，凡跟随她的必用刀杀死！”因为祭司说：“不可在耶和华殿里杀她。”
2CHR|23|15|他们就下手拿住她；她进入通往王宫的 马门 ，他们就在那里把她杀了。
2CHR|23|16|耶何耶大 与众百姓，又与王立约，要作耶和华的子民。
2CHR|23|17|于是众百姓到 巴力 庙去，拆毁了庙，打碎祭坛和偶像，又在坛前把 巴力 的祭司 玛坦 杀了。
2CHR|23|18|耶何耶大 派官员在 利未 家的祭司手下看守耶和华的殿，他们是 大卫 所分派的，在耶和华殿中照 摩西 律法上所写，献燔祭给耶和华，又按 大卫 所定的，欢乐歌唱。
2CHR|23|19|耶何耶大 又设立守卫把守耶和华殿的各门，无论因何事而不洁净的人，都不准进去。
2CHR|23|20|他又率领百夫长和贵族，与民间的官长，以及国中的众百姓，请王从耶和华的殿下来，由 上门 正中进入王宫，使王坐在国度的王位上。
2CHR|23|21|国中的众百姓都欢乐，合城也都平静。他们已将 亚她利雅 用刀杀了。
2CHR|24|1|约阿施 登基的时候年方七岁，在 耶路撒冷 作王四十年。他母亲名叫 西比亚 ，是 别是巴 人。
2CHR|24|2|耶何耶大 祭司在世的日子， 约阿施 行耶和华眼中看为正的事。
2CHR|24|3|耶何耶大 为他娶了两个妻子，他生儿育女。
2CHR|24|4|此后， 约阿施 有心重修耶和华的殿，
2CHR|24|5|就召集祭司和 利未 人，吩咐他们说：“你们要往 犹大 各城去，向 以色列 众人征收银子，按每年的需要整修你们上帝的殿；你们要急速办理这事。”但 利未 人没有急速办理。
2CHR|24|6|王召了 耶何耶大 祭司长来，对他说：“从前耶和华的仆人 摩西 ，为法柜的帐幕与 以色列 会众所定的捐献，你为何不叫 利未 人照这例向 犹大 和 耶路撒冷 征收呢？”
2CHR|24|7|因为那恶妇 亚她利雅 的儿子们曾拆毁上帝的殿，又用耶和华殿中分别为圣的物供奉诸 巴力 。
2CHR|24|8|于是王下令造一个柜子，放在耶和华殿的门外，
2CHR|24|9|又通告 犹大 和 耶路撒冷 ，要将上帝仆人 摩西 在旷野所吩咐 以色列 的捐献送来给耶和华。
2CHR|24|10|众领袖和百姓都欢欢喜喜带捐献来，投入柜中，直到投满。
2CHR|24|11|利未 人见银子多了，把柜子抬到王所派的官长面前；这时王的书记和祭司长的助手就会来把柜子倒空，然后放回原处。日日都是这样做，积蓄的银子很多。
2CHR|24|12|王与 耶何耶大 把银子交给耶和华殿里办事的人，他们就雇了石匠、木匠重修耶和华的殿，又雇了铁匠、铜匠整修耶和华的殿。
2CHR|24|13|工人做工，修理工程在他们手中渐渐完成，他们将上帝的殿修理得如同从前一样，非常坚固。
2CHR|24|14|他们做完了，就把多余的银子拿到王与 耶何耶大 面前，用以制造耶和华殿供奉所用的器皿和调羹，以及金银的器皿。 耶何耶大 在世的日子，众人经常在耶和华殿里献燔祭。
2CHR|24|15|耶何耶大 年纪老迈，日子满足而死，死的时候年一百三十岁。
2CHR|24|16|众人把他与列王同葬在 大卫城 ，因为他在 以色列 中为上帝和他的殿做了美善的事。
2CHR|24|17|耶何耶大 死后， 犹大 的众领袖来叩拜王，那时王就听了他们。
2CHR|24|18|他们离弃耶和华－他们列祖上帝的殿，去事奉 亚舍拉 和偶像；因他们这罪，就有愤怒临到 犹大 和 耶路撒冷 。
2CHR|24|19|但上帝仍差遣先知到他们那里，引导他们归向耶和华。先知警戒他们，他们却不肯听。
2CHR|24|20|那时，上帝的灵感动 耶何耶大 的儿子 撒迦利亚 祭司，他就站在上面，对百姓说：“上帝如此说：‘你们为何干犯耶和华的诫命，以致不得亨通呢？因为你们离弃耶和华，所以他也离弃你们。’”
2CHR|24|21|众人谋害 撒迦利亚 ，照着王的吩咐，在耶和华殿的院内用石头打死他。
2CHR|24|22|这样， 约阿施 王不记念 撒迦利亚 的父亲 耶何耶大 向自己所施的恩，杀了他的儿子。 撒迦利亚 临死的时候说：“愿耶和华鉴察伸冤！”
2CHR|24|23|年底的时候， 亚兰 的军兵上来攻击 约阿施 ，来到 犹大 和 耶路撒冷 ，杀了百姓中的众领袖，把所掠取的财物全送到 大马士革 王那里。
2CHR|24|24|亚兰 的军兵虽只来了一小队人，耶和华却将极大的军队交在他们手里；因为 犹大 人离弃耶和华－他们列祖的上帝，所以 亚兰 人惩罚 约阿施 。
2CHR|24|25|亚兰 人离开 约阿施 的时候，他患重病 ；他的臣仆背叛他，要报 耶何耶大 祭司儿子 的流血之仇，在床上杀了他。他就死了，葬在 大卫城 ，只是不葬在列王的坟墓里。
2CHR|24|26|背叛他的是 亚扪 妇人 示米押 的儿子 撒拔 和 摩押 妇人 示米利 的儿子 约萨拔 。
2CHR|24|27|至于他的儿子们和他所受的众多警戒，以及他重修上帝殿的事，看哪，都写在《列王评传》上。他的儿子 亚玛谢 接续他作王。
2CHR|25|1|亚玛谢 登基的时候年二十五岁，在 耶路撒冷 作王二十九年。他母亲名叫 约耶但 ，是 耶路撒冷 人。
2CHR|25|2|亚玛谢 行耶和华眼中看为正的事，只是没有纯正的心。
2CHR|25|3|他的王国一巩固，就把杀他父王的臣仆杀了，
2CHR|25|4|却没有处死他们的儿子，这是照 摩西 律法书上耶和华所吩咐的说：“不可因子杀父，也不可因父杀子，各人要为自己的罪而死。”
2CHR|25|5|亚玛谢 召集 犹大 人，按着父家为全 犹大 和 便雅悯 设立千夫长、百夫长，又数点人数，从二十岁以上，能拿枪拿盾牌出去打仗的精兵共有三十万；
2CHR|25|6|又用一百他连得银子，从 以色列 招募了十万大能的勇士。
2CHR|25|7|有一个神人来见 亚玛谢 ，对他说：“王啊，不要带领 以色列 的军兵与你同去，因为耶和华不和 以色列 ，和任何 以法莲 的子孙同在。
2CHR|25|8|你若一定要去，就奋勇作战吧！但上帝必使你败在敌人面前，因为上帝能助人得胜，也能使人落败。”
2CHR|25|9|亚玛谢 问神人：“我给了 以色列 军队的那一百他连得银子怎么样呢？”神人回答：“耶和华会把比这些更多的赐给你。”
2CHR|25|10|于是 亚玛谢 把那从 以法莲 来的军兵分别出来，叫他们到自己的地方去。他们非常恼怒 犹大 ，气愤地回自己的地方去了。
2CHR|25|11|亚玛谢 壮起胆来，率领他的军队到 盐谷 ，杀了一万 西珥 人。
2CHR|25|12|犹大 人又生擒了一万人，把他们带到 西拉 山顶上，从 西拉 山顶扔下去，把他们全都摔碎了。
2CHR|25|13|但 亚玛谢 所打发回去、不许一同出征的那些军兵劫掠 犹大 各城，从 撒玛利亚 直到 伯．和仑 ，杀了三千人，抢了许多财物。
2CHR|25|14|亚玛谢 击杀 以东 人回来以后，他把 西珥 人的神像带回，立为自己的神明，在它们面前叩拜烧香。
2CHR|25|15|耶和华的怒气向 亚玛谢 发作，差派一个先知去见他，对他说：“这些神明不能救自己的百姓脱离你的手，你为何寻求它们呢？”
2CHR|25|16|先知与王说话的时候，王对他说：“难道我们立你作王的谋士吗？你住口吧！为何要挨打呢？”先知就止住了，却说：“我知道上帝已定意要消灭你，因为你行这事，不听从我的劝戒。”
2CHR|25|17|犹大 王 亚玛谢 经商议后，就派人去见 耶户 的孙子， 约哈斯 的儿子 以色列 王 约阿施 ，说：“来，让我们面对面较量吧！”
2CHR|25|18|以色列 王 约阿施 派人去见 犹大 王 亚玛谢 ，说：“ 黎巴嫩 的蒺藜派人去见 黎巴嫩 的香柏树，说：‘将你的女儿嫁给我的儿子。’但有一只野兽经过 黎巴嫩 ，把蒺藜践踏了。
2CHR|25|19|你说，看哪，你打败了 以东 ，就心高气傲，以此为荣。现在，你待在家里算了吧，为何要惹祸使自己和 犹大 一同败亡呢？”
2CHR|25|20|亚玛谢 却不肯听从。这是出乎上帝，好将他们交在敌人手里，因为他们寻求 以东 的神明。
2CHR|25|21|于是 以色列 王 约阿施 上来，在 犹大 的 伯．示麦 与 犹大 王 亚玛谢 面对面较量。
2CHR|25|22|犹大 败在 以色列 面前，他们逃跑，各人逃回自己的帐棚去了。
2CHR|25|23|以色列 王 约阿施 在 伯．示麦 擒住 约哈斯 的孙子， 约阿施 的儿子 犹大 王 亚玛谢 ，把他带到 耶路撒冷 ，又拆毁 耶路撒冷 的城墙，从 以法莲门 直到 角门 共四百肘。
2CHR|25|24|他带着 俄别．以东 所看守上帝殿里的一切金银和器皿，与王宫里的财宝，又带着人质，回 撒玛利亚 去了。
2CHR|25|25|约哈斯 的儿子 以色列 王 约阿施 死后， 犹大 王 约阿施 的儿子 亚玛谢 又活了十五年。
2CHR|25|26|亚玛谢 其余的事，自始至终，看哪，不都写在《犹大和以色列诸王记》上吗？
2CHR|25|27|自从 亚玛谢 离弃耶和华之后，在 耶路撒冷 有人背叛他，他就逃往 拉吉 ；他们却派人追到 拉吉 ，在那里杀了他。
2CHR|25|28|有人用马将他驮回，把他与祖先一同葬在 犹大 的城 。
2CHR|26|1|犹大 众百姓立 乌西雅 接续他父亲 亚玛谢 作王，那时他年十六岁。
2CHR|26|2|亚玛谢 王与他祖先同睡之后， 乌西雅 收复 以禄 回归 犹大 ，又重新修建。
2CHR|26|3|乌西雅 登基的时候年十六岁，在 耶路撒冷 作王五十二年。他母亲名叫 耶可利雅 ，是 耶路撒冷 人。
2CHR|26|4|乌西雅 行耶和华眼中看为正的事，效法他父亲 亚玛谢 一切所行的。
2CHR|26|5|撒迦利亚 是一个通晓上帝默示的人 ，他在世的日子， 乌西雅 定意寻求上帝； 乌西雅 寻求耶和华的日子，上帝使他亨通。
2CHR|26|6|他出去攻击 非利士 人，拆毁了 迦特 、 雅比尼 和 亚实突 的城墙，又在 非利士 人中，在 亚实突 境内建筑城镇。
2CHR|26|7|上帝帮助他攻击 非利士 人和住在 姑珥．巴力 的 阿拉伯 人，以及 米乌尼 人。
2CHR|26|8|米乌尼 人 向 乌西雅 进贡。他的名声传到 埃及 ，因他非常强盛。
2CHR|26|9|乌西雅 在 耶路撒冷 的 角门 和 谷门 ，以及城墙转角之处建筑城楼，非常坚固。
2CHR|26|10|他在旷野建筑了望楼，又挖了许多井，因为他在 谢非拉 和平原有很多牲畜。他在山区和肥沃的土地雇用耕种田地和修整葡萄园的人，因为他喜爱土地。
2CHR|26|11|乌西雅 又有军兵，照书记 耶利 和官长 玛西雅 所数点的，在王的一个将军 哈拿尼雅 手下，分队出战。
2CHR|26|12|族长和大能勇士的总数共二千六百人，
2CHR|26|13|他们手下的军兵共三十万七千五百人，都大有能力，善于作战，帮助王攻击仇敌。
2CHR|26|14|乌西雅 为全军预备盾牌、头盔、铠甲、枪、弓和甩石的机弦，
2CHR|26|15|又在 耶路撒冷 叫巧匠设计机器，安在城楼和角楼上，用以射箭，投掷大石。 乌西雅 的名声传到远方，因为他得了非凡的帮助，极其强盛。
2CHR|26|16|乌西雅 既强盛，就心高气傲，以致败坏。他干犯耶和华－他的上帝，进耶和华的殿，要在香坛上烧香。
2CHR|26|17|亚撒利雅 祭司率领八十名勇敢的耶和华的祭司，跟随他进去。
2CHR|26|18|他们阻止 乌西雅 王，对他说：“ 乌西雅 啊，给耶和华烧香不是你的事，而是 亚伦 子孙的事，他们是分别为圣来烧香的祭司。你出圣殿吧！因为你犯了罪，耶和华上帝必不使你得尊荣。”
2CHR|26|19|乌西雅 发怒，手拿香炉要烧香。他在耶和华殿中香坛旁向众祭司发怒的时候，他的额头在众祭司面前忽然长出痲疯 。
2CHR|26|20|亚撒利雅 祭司长和众祭司转向他，看哪，他的额头长出痲疯，就催他离开那里；他自己也急速出去，因为耶和华降灾于他。
2CHR|26|21|乌西雅 王患痲疯直到死的那日；他因为染上痲疯，就住在隔离的行宫里，与耶和华的殿隔绝。他儿子 约坦 管理王的家，治理这地的百姓。
2CHR|26|22|乌西雅 其余的事，自始至终， 亚摩斯 的儿子 以赛亚 先知都记录下来。
2CHR|26|23|乌西雅 与他祖先同睡，与他祖先同葬在田间的王陵；因为人说，他是长痲疯的。他的儿子 约坦 接续他作王。
2CHR|27|1|约坦 登基的时候年二十五岁，在 耶路撒冷 作王十六年。他母亲名叫 耶路沙 ，是 撒督 的女儿。
2CHR|27|2|约坦 行耶和华眼中看为正的事，效法他父亲 乌西雅 一切所行的，只是他不入耶和华的殿。百姓仍旧行败坏的事。
2CHR|27|3|约坦 建造耶和华殿的 上门 ，在 俄斐勒 城墙上有很多建设，
2CHR|27|4|又在 犹大 山区建造城镇，在树林中建筑营寨和了望楼。
2CHR|27|5|约坦 与 亚扪 人的王打仗，胜了他们。那年 亚扪 人向他进贡一百他连得银子，一万歌珥小麦，一万歌珥大麦；第二年、第三年 亚扪 人也这样做。
2CHR|27|6|约坦 日渐强盛，因为他在耶和华－他上帝面前行正道。
2CHR|27|7|约坦 其余的事和一切战役，以及他的行为，看哪，都写在《以色列和犹大列王记》上。
2CHR|27|8|他登基的时候年二十五岁，在 耶路撒冷 作王十六年。
2CHR|27|9|约坦 与他祖先同睡，葬在 大卫城 ，他儿子 亚哈斯 接续他作王。
2CHR|28|1|亚哈斯 登基的时候年二十岁，在 耶路撒冷 作王十六年。他不像他祖先 大卫 行耶和华眼中看为正的事，
2CHR|28|2|却行 以色列 诸王的道，又铸造诸 巴力 的像，
2CHR|28|3|照着耶和华从 以色列 人面前赶出的外邦人所行可憎的事，在 欣嫩子谷 烧香，用火焚烧他的儿女，
2CHR|28|4|又在丘坛上、山冈上、各青翠树下献祭烧香。
2CHR|28|5|耶和华－他的上帝将他交在 亚兰 王手里。 亚兰 王打败他，从他掳走了许多人，带到 大马士革 去。上帝又将他交在 以色列 王手里， 以色列 王向他大行杀戮。
2CHR|28|6|利玛利 的儿子 比加 一日之内在 犹大 杀了十二万人，都是勇士，因为他们离弃了耶和华－他们列祖的上帝。
2CHR|28|7|有一个叫 细基利 的 以法莲 勇士，杀了 玛西雅 王子、 押斯利甘 宫廷总管和 以利加拿 宰相。
2CHR|28|8|以色列 人掳了他们的弟兄，连妇人带儿女共二十万，又掠取了许多财物，把这些掠物带到 撒玛利亚 去。
2CHR|28|9|但那里有耶和华的一个先知，名叫 俄德 ，出来迎接往 撒玛利亚 去的军兵，对他们说：“看哪，耶和华－你们列祖的上帝恼怒 犹大 人，将他们交在你们手里，你们竟怒气冲天，向他们大行杀戮。
2CHR|28|10|如今你们又有意强逼 犹大 人和 耶路撒冷 人作你们的奴婢，你们岂不是也得罪了耶和华－你们的上帝吗？
2CHR|28|11|现在你们当听我说，要将从你们弟兄中掳来的释放回去，因耶和华的烈怒已临到你们了。”
2CHR|28|12|于是， 以法莲 人的几个领袖，就是 约哈难 的儿子 亚撒利雅 、 米实利末 的儿子 比利家 、 沙龙 的儿子 耶希西家 、 哈得莱 的儿子 亚玛撒 ，起来拦阻从战场上回来的人，
2CHR|28|13|对他们说：“你们不可把这些被掳的人带到这里，因我们已经得罪耶和华了。你们还想加增我们的罪恶过犯吗？因为我们的罪过深重，已经有烈怒临到 以色列 了。”
2CHR|28|14|于是带兵器的人将掳来的人口和掠取的财物都留在众领袖和全会众面前。
2CHR|28|15|以上提名的那些人就起来，照顾被掳的人；其中凡赤身的，就从所掠取的财物中拿出衣服和鞋来，给他们穿，又给他们吃喝，用膏抹他们；其中凡软弱的，就使他们骑驴，送到棕树城 耶利哥 他们弟兄那里。然后，他们就回 撒玛利亚 去了。
2CHR|28|16|那时， 亚哈斯 王派人去求 亚述 诸王 来帮助他，
2CHR|28|17|因为 以东 人又来攻击 犹大 ，掳掠俘虏。
2CHR|28|18|非利士 人也来侵占 谢非拉 和 犹大 的 尼革夫 的城镇，攻取了 伯．示麦 、 亚雅仑 、 基低罗 、 梭哥 和所属的乡镇、 亭拿 和所属的乡镇、 瑾锁 和所属的乡镇，就住在那里。
2CHR|28|19|因为 以色列 王 亚哈斯 在 犹大 放肆，大大干犯耶和华，所以耶和华使 犹大 卑微。
2CHR|28|20|亚述 王 提革拉．毗列色 来攻击他，不帮助他，反倒欺负他。
2CHR|28|21|亚哈斯 从耶和华殿里和王宫中，以及众领袖家中取财宝送给 亚述 王，也无济于事。
2CHR|28|22|这 亚哈斯 王在急难的时候，越发得罪耶和华。
2CHR|28|23|他向那攻击他的 大马士革 的神明献祭，说：“因为 亚兰 王的神明帮助他们，我也要向这些神明献祭，好让它们帮助我。”但那些神明却使他和全 以色列 败亡。
2CHR|28|24|亚哈斯 聚集上帝殿里的器皿，把上帝殿里的器皿都打碎了，并且封锁耶和华殿的门，又在 耶路撒冷 各处的转角为自己建筑祭坛。
2CHR|28|25|他在 犹大 各城建立丘坛，向别神烧香，惹耶和华－他列祖的上帝发怒。
2CHR|28|26|亚哈斯 其余的事和他一切的行为，自始至终，看哪，都写在《犹大和以色列诸王记》上。
2CHR|28|27|亚哈斯 与他祖先同睡，葬在 耶路撒冷 城里，却没有送入 以色列 诸王的坟墓。他的儿子 希西家 接续他作王。
2CHR|29|1|希西家 登基的时候年二十五岁，在 耶路撒冷 作王二十九年。他母亲名叫 亚比雅 ，是 撒迦利雅 的女儿。
2CHR|29|2|希西家 行耶和华眼中看为正的事，效法他祖先 大卫 一切所行的。
2CHR|29|3|元年正月，他开了耶和华殿的门，重新整修。
2CHR|29|4|他召祭司和 利未 人来，聚集在东边的广场，
2CHR|29|5|对他们说：“ 利未 人哪，当听我说：现在你们要将自己分别为圣，又将耶和华－你们列祖上帝的殿分别为圣，从圣所中除去污秽之物。
2CHR|29|6|因我们的祖先犯了罪，行耶和华－我们上帝眼中看为恶的事，离弃他，转脸背向耶和华的居所。
2CHR|29|7|他们又封锁走廊的门，吹灭灯火，不在圣所中向 以色列 的上帝烧香，或献燔祭。
2CHR|29|8|耶和华的愤怒临到 犹大 和 耶路撒冷 ，使他们恐惧，令人惊骇，使人嗤笑，正如你们亲眼所见的。
2CHR|29|9|看哪，我们的祖宗倒在刀下，我们的妻子儿女也为此被掳掠。
2CHR|29|10|现在我心中有意与耶和华－ 以色列 的上帝立约，好使他的烈怒转离我们。
2CHR|29|11|我的众子啊，现在不要懈怠；因为耶和华拣选你们站在他面前事奉他，作他的仆人，向他烧香。”
2CHR|29|12|于是， 利未 人起来，当中有 哥辖 的子孙， 亚玛赛 的儿子 玛哈 、 亚撒利雅 的儿子 约珥 ； 米拉利 的子孙， 亚伯底 的儿子 基士 、 耶哈利勒 的儿子 亚撒利雅 ； 革顺 人， 薪玛 的儿子 约亚 、 约亚 的儿子 伊甸 ；
2CHR|29|13|以利撒反 的子孙 申利 和 耶利 ； 亚萨 的子孙， 撒迦利雅 和 玛探雅 ；
2CHR|29|14|希幔 的子孙 耶歇 和 示每 ； 耶杜顿 的子孙 示玛雅 和 乌薛 。
2CHR|29|15|他们聚集他们的弟兄，将自己分别为圣，照着耶和华的话和王的吩咐，进去洁净耶和华的殿。
2CHR|29|16|祭司进入耶和华的内殿要洁净殿，把耶和华殿中所发现一切污秽之物都搬出去，搬到耶和华殿的院子，由 利未 人接走，搬出去到外头的 汲沦溪 。
2CHR|29|17|从正月初一开始分别为圣，初八就来到耶和华殿的走廊。他们又用了八日使耶和华的殿分别为圣，到正月十六日才完成。
2CHR|29|18|于是，他们到里面去见 希西家 王，说：“我们已将耶和华的全殿和燔祭坛，以及坛的一切器皿、供饼的供桌，与供桌的一切器皿都洁净了；
2CHR|29|19|并且连 亚哈斯 王在位犯罪的时候所废弃的器皿，我们也都预备齐全，分别为圣，看哪，它们都在耶和华的祭坛前。”
2CHR|29|20|希西家 王清早起来，召集城里的领袖都上耶和华的殿。
2CHR|29|21|他们牵了七头公牛，七只公羊，七只羔羊，七只公山羊，要为国、为殿、为 犹大 作赎罪祭。王吩咐 亚伦 的子孙众祭司在耶和华的坛上献祭。
2CHR|29|22|他们宰了公牛，祭司将血接来，洒在坛上；他们宰了公羊，把血洒在坛上，又宰了羔羊，也把血洒在坛上。
2CHR|29|23|他们把那些作赎罪祭的公山羊牵到王和会众面前，按手在公山羊上。
2CHR|29|24|祭司宰了羊，将血献在坛上作赎罪祭，为全 以色列 赎罪，因为王吩咐要为全 以色列 献上燔祭和赎罪祭。
2CHR|29|25|王又派 利未 人在耶和华殿中敲钹，鼓瑟，弹琴，正如 大卫 和王的先见 迦得 ，以及 拿单 先知所吩咐的，就是耶和华藉先知所吩咐的。
2CHR|29|26|利未 人拿 大卫 的乐器，祭司拿号，一同站立。
2CHR|29|27|希西家 吩咐在坛上献燔祭，开始献燔祭的时候，他们就唱赞美耶和华的歌，吹号，并用 以色列 王 大卫 的乐器伴奏。
2CHR|29|28|全会众都敬拜，歌唱的歌唱，吹号的吹号，如此直到燔祭献完了。
2CHR|29|29|献完了祭，王和所有在场跟随他的人都俯伏敬拜。
2CHR|29|30|希西家 王与众领袖吩咐 利未 人用 大卫 和 亚萨 先见的诗词颂赞耶和华，他们欢欢喜喜地颂赞，低头敬拜。
2CHR|29|31|希西家 回应说：“如今你们既承接圣职归耶和华，就要前来把祭物和感谢祭奉到耶和华的殿里。”会众就奉上祭物和感谢祭，凡甘心乐意的也奉上燔祭。
2CHR|29|32|会众所奉的燔祭数目如下：七十头公牛，一百只公羊，二百只羔羊，这些全都是要作燔祭献给耶和华的；
2CHR|29|33|又有分别为圣之物，就是六百头公牛，三千只绵羊。
2CHR|29|34|但祭司太少，不能剥尽所有燔祭牲的皮，所以他们的弟兄 利未 人帮助他们，直等献祭的事完毕，直到其他的祭司也分别为圣了；因 利未 人以正直的心分别为圣，胜过祭司。
2CHR|29|35|燔祭和平安祭牲的脂肪，以及与燔祭同献的浇酒祭很多。这样，耶和华殿中的事务俱都齐备了。
2CHR|29|36|希西家 和众百姓都因上帝为百姓所预备的而喜乐，因为这事办得很迅速。
2CHR|30|1|希西家 派人去见 以色列 和 犹大 众人，又写信给 以法莲 和 玛拿西 人，要他们到 耶路撒冷 耶和华的殿，向耶和华－ 以色列 的上帝守逾越节，
2CHR|30|2|因为王和众领袖，以及 耶路撒冷 全会众已经商议，要在二月份守逾越节。
2CHR|30|3|那时他们不能守，因为分别为圣的祭司不够，百姓也还没有聚集在 耶路撒冷 。
2CHR|30|4|这事在王与全会众眼中都看为合宜。
2CHR|30|5|于是他们下令，通告全 以色列 ，从 别是巴 直到 但 ，吩咐百姓都来，在 耶路撒冷 向耶和华－ 以色列 的上帝守逾越节，因为他们已经许久没有照所写的守这节了 。
2CHR|30|6|信差遵着王命，拿着王和众领袖所发的信，送达全 以色列 和 犹大 ，说：“ 以色列 人哪，当转向耶和华－ 亚伯拉罕 、 以撒 、 以色列 的上帝，好叫他转向你们这些脱离 亚述 诸王之手的余民。
2CHR|30|7|不要效法你们的祖先和你们的弟兄；他们干犯耶和华－他们列祖的上帝，以致耶和华使他们令人惊骇，正如你们所见的。
2CHR|30|8|现在，不要像你们祖先硬着颈项，只要归顺耶和华，进入他的圣所，就是永远成圣的居所，又要事奉耶和华－你们的上帝，好使他的烈怒转离你们。
2CHR|30|9|你们若转向耶和华，你们的弟兄和儿女必在掳掠他们的人面前蒙怜悯，得以归回这地，因为耶和华－你们的上帝有恩惠，有怜悯。你们若转向他，他必不会转脸不顾你们。”
2CHR|30|10|信差从这城跑到那城，传遍了 以法莲 和 玛拿西 之地，直到 西布伦 ；那里的人却戏笑他们，讥诮他们。
2CHR|30|11|然而 亚设 、 玛拿西 、 西布伦 中也有人谦卑自己，来到 耶路撒冷 。
2CHR|30|12|上帝也按手在 犹大 人身上，使他们一心遵行王与众领袖照着耶和华的话所发的命令。
2CHR|30|13|二月时，许多百姓聚集在 耶路撒冷 ，成为一个盛大的会，要守除酵节。
2CHR|30|14|他们起来，把 耶路撒冷 的祭坛和烧香的坛尽都除去，扔在 汲沦溪 中。
2CHR|30|15|二月十四日，他们宰了逾越节的羔羊。祭司与 利未 人觉得惭愧，就使自己分别为圣，把燔祭奉到耶和华的殿中。
2CHR|30|16|他们遵照神人 摩西 的律法，按定例站在自己的地方；祭司从 利未 人手里接过血来，洒出去。
2CHR|30|17|会众中有许多人尚未分别为圣，所以 利未 人为所有不洁的人宰逾越节的羔羊，使他们归耶和华为圣。
2CHR|30|18|从 以法莲 、 玛拿西 、 以萨迦 、 西布伦 来的许多百姓尚未自洁，他们却吃逾越节的羔羊，不合所写的条例。 希西家 为他们祷告说：“求至善的耶和华饶恕
2CHR|30|19|那凡专心寻求上帝耶和华－他列祖的上帝，却未照圣所洁净礼自洁的人。”
2CHR|30|20|耶和华应允 希西家 ，医治了百姓。
2CHR|30|21|在 耶路撒冷 的 以色列 人守除酵节七日，大大喜乐。 利未 人和祭司为耶和华演奏响亮的乐器，天天颂赞耶和华。
2CHR|30|22|希西家 慰劳所有精通礼仪，事奉耶和华的 利未 人。于是众人吃节期的筵席七日，又献平安祭，并且称谢耶和华－他们列祖的上帝。
2CHR|30|23|全会众商议，要再守节七日；于是他们欢欢喜喜地又守节七日。
2CHR|30|24|犹大 王 希西家 赐给会众一千头公牛，七千只羊；众领袖也赐给会众一千头公牛，一万只羊，并有许多祭司将自己分别为圣。
2CHR|30|25|犹大 全会众、祭司、 利未 人和从 以色列 来的全会众，以及那些从 以色列 地来的和住在 犹大 的寄居的人，尽都喜乐。
2CHR|30|26|这样，在 耶路撒冷 大有喜乐，因自从 以色列 王 大卫 的儿子 所罗门 以来，在 耶路撒冷 从未有过这样的喜乐。
2CHR|30|27|那时，祭司和 利未 人起来，为百姓祝福。他们的声音蒙上帝垂听，他们的祷告达到他天上的圣所。
2CHR|31|1|这一切事都完毕以后，在那里的 以色列 众人就到 犹大 的城镇，打碎柱像，砍断 亚舍拉 ，又在 犹大 、 便雅悯 、 以法莲 、 玛拿西 遍地把丘坛和祭坛完全拆毁。于是 以色列 众人各回各城，各归自己产业的地去了。
2CHR|31|2|希西家 分派祭司和 利未 人的班次，使祭司和 利未 人照各自的班次，按各自的职分献燔祭和平安祭，又在耶和华殿 的门内事奉，称谢颂赞耶和华。
2CHR|31|3|王又从自己的产业中分出一份来作燔祭，就是早晚的燔祭，和安息日、初一，以及节期的燔祭，都是按耶和华律法上所记载的。
2CHR|31|4|他又吩咐住 耶路撒冷 的百姓将祭司和 利未 人所应得的份给他们，使他们坚守耶和华的律法。
2CHR|31|5|命令一出， 以色列 人就把初熟的五谷、新酒、新油、蜜和田地的出产多多送来；他们把各样出产的十分之一大量送来。
2CHR|31|6|住 犹大 各城的 以色列 人和 犹大 人也将牛羊的十分之一，以及分别为圣归耶和华－他们上帝之物，就是十分取一之物，尽都送来，积成一堆一堆；
2CHR|31|7|他们从三月开始堆积，到七月才完成。
2CHR|31|8|希西家 和众领袖来，看见这些堆积物，就称颂耶和华，又为耶和华的百姓 以色列 祝福。
2CHR|31|9|希西家 向祭司和 利未 人查问这些堆积物。
2CHR|31|10|撒督 家的 亚撒利雅 祭司长告诉他说：“自从礼物开始送到耶和华的殿以来，我们不但吃饱，而且剩下的很多；因为耶和华赐福给他的百姓，所剩下的才这样丰盛。”
2CHR|31|11|希西家 吩咐要在耶和华殿里预备仓房，他们就预备了。
2CHR|31|12|他们诚心将礼物，十分取一之物，就是分别为圣之物，都搬入仓内。 利未 人 歌楠雅 主管这事，他的兄弟 示每 是副主管。
2CHR|31|13|耶歇 、 亚撒细雅 、 拿哈 、 亚撒黑 、 耶利摩 、 约撒拔 、 以列 、 伊斯玛基雅 、 玛哈 、 比拿雅 都是督办，在 歌楠雅 和他兄弟 示每 的手下，是 希西家 王和管理上帝殿的 亚撒利雅 所委派的。
2CHR|31|14|守东门的 利未 人 音拿 的儿子 可利 ，掌管献给上帝的甘心祭，发放献给耶和华的礼物和至圣的物。
2CHR|31|15|在祭司的各城里，在他手下忠心协助他的有 伊甸 、 (王民)雅(王民) 、 耶书亚 、 示玛雅 、 亚玛利雅 、 示迦尼雅 ，都按着班次分给他们的弟兄，无论大小，
2CHR|31|16|不论是否登录在家谱，凡三岁以上的男丁，每日进耶和华殿、按班次供职事奉的，都分给他，
2CHR|31|17|也发放给按父家登录在家谱的祭司；又按班次职任分给二十岁以上的 利未 人，
2CHR|31|18|又按家谱的登记，分给他们的小孩、妻子、儿女，给全体会众；因为他们忠诚，将自己分别为圣。
2CHR|31|19|住在各城郊野 亚伦 的子孙、按名受委任的人，要把应得的份给祭司中所有的男丁和载入家谱的 利未 人。
2CHR|31|20|希西家 在全 犹大 都这样办理，在耶和华－他上帝面前行良善、正直、忠诚的事。
2CHR|31|21|凡他所行的，无论是开始办上帝殿的事，是遵律法守诫命，是寻求他的上帝，他都尽心去做，无不亨通。
2CHR|32|1|在这些虔诚的事以后， 亚述 王 西拿基立 来侵犯 犹大 ，围困坚固城，想要攻破它们。
2CHR|32|2|希西家 见 西拿基立 来，定意要攻打 耶路撒冷 ，
2CHR|32|3|就与领袖和勇士商议，塞住城外的泉源；他们都帮助他。
2CHR|32|4|于是许多百姓聚集，塞住一切泉源，以及国中流通的小河，说：“ 亚述 诸王来，为何让他们得着许多水呢？”
2CHR|32|5|希西家 奋勇自强，修筑所有毁坏的城墙，升高城楼，又在城外筑另一片城墙，坚固 大卫城 的 米罗 ，制造许多兵器和盾牌。
2CHR|32|6|他设立军事将领管理百姓，召集他们在城门的广场，勉励他们，说：
2CHR|32|7|“你们当刚强壮胆，不要因 亚述 王和跟随他的大军恐惧惊慌，因为与我们同在的，比与他们同在的更大。
2CHR|32|8|与他们同在的是血肉之臂，但与我们同在的是耶和华－我们的上帝，他必帮助我们，为我们争战。”百姓因 犹大 王 希西家 的话就得到鼓励。
2CHR|32|9|此后， 亚述 王 西拿基立 和跟随他的全军攻打 拉吉 ，派臣仆到 耶路撒冷 见 犹大 王 希西家 和所有在 耶路撒冷 的 犹大 人，说：
2CHR|32|10|“ 亚述 王 西拿基立 如此说：‘你们倚靠什么，还留在 耶路撒冷 受困吗？
2CHR|32|11|希西家 说：耶和华－我们的上帝必救我们脱离 亚述 王的手，这不是诱惑你们，使你们受饥渴而死吗？
2CHR|32|12|希西家 岂不是将耶和华的丘坛和祭坛废去，并且吩咐 犹大 与 耶路撒冷 的人说：你们当在一个坛前敬拜，在其上烧香吗？
2CHR|32|13|我与我祖先向列邦民族所行的，你们岂不知道吗？列邦的神明何尝能救自己的国脱离我的手呢？
2CHR|32|14|我祖先所灭的那些国的神明，有谁能救自己的百姓脱离我的手呢？难道你们的上帝能救你们脱离我的手吗？
2CHR|32|15|现在，不要让 希西家 这样欺骗你们，诱惑你们，也不要相信他，因为没有一国一邦的神明能救自己的百姓脱离我的手和我祖先的手，你们的上帝也绝不能救你们脱离我的手。’”
2CHR|32|16|西拿基立 的臣仆还说了一些话来毁谤耶和华上帝和他的仆人 希西家 。
2CHR|32|17|西拿基立 也写信毁谤耶和华－ 以色列 的上帝，说：“列邦的神明既不能救自己的百姓脱离我的手， 希西家 的上帝也不能救他的百姓脱离我的手。”
2CHR|32|18|亚述 王的臣仆用 犹大 话向 耶路撒冷 城墙上的百姓大声呼喊，要恐吓他们，扰乱他们，以便取城。
2CHR|32|19|他们谈论 耶路撒冷 的上帝，如同谈论世上人手所造的神明一样。
2CHR|32|20|希西家 王和 亚摩斯 的儿子 以赛亚 先知为此祷告，向天呼求。
2CHR|32|21|耶和华就差遣一个使者进入 亚述 王的营中，把所有大能的勇士、官长和将领尽都灭了。 亚述 王满面羞愧地回到本国，进了他神明的庙中，他几个亲生的儿子在那里用刀杀了他。
2CHR|32|22|这样，耶和华救 希西家 和 耶路撒冷 的居民脱离 亚述 王 西拿基立 的手，也脱离一切仇敌的手，又赐他们四境平安 。
2CHR|32|23|有许多人到 耶路撒冷 将供物献与耶和华，又将宝物送给 犹大 王 希西家 。自此之后， 希西家 在列国人的眼中受人尊崇。
2CHR|32|24|那些日子， 希西家 病得要死，就向耶和华祷告，耶和华应允他，赐他一个预兆。
2CHR|32|25|希西家 却没有照他所蒙的恩回报，因他心里骄傲，所以愤怒要临到他，临到 犹大 和 耶路撒冷 。
2CHR|32|26|但 希西家 和 耶路撒冷 的居民为了心里骄傲，就一同谦卑，以致耶和华的愤怒在 希西家 的日子没有临到他们。
2CHR|32|27|希西家 大有财富和尊荣，他为自己建造府库，收藏金银、宝石、香料、盾牌和各样的宝器，
2CHR|32|28|又建造仓房，收藏五谷、新酒和新的油，又为各类牲畜盖棚立圈，
2CHR|32|29|并且为自己建立城镇，也拥有许多的羊群牛群，因为上帝赐他极多的财产。
2CHR|32|30|这 希西家 也塞住 基训 的上源，引水直下，流在 大卫城 的西边。 希西家 所行的事尽都亨通。
2CHR|32|31|但当 巴比伦 诸侯差遣使者来见 希西家 ，询问国中所发生的奇事时，上帝离开他，要考验他，好知道他心里的一切。
2CHR|32|32|希西家 其余的事和他的善行，看哪，都写在 亚摩斯 的儿子 以赛亚 先知的《默示书》上和《犹大和以色列诸王记》上。
2CHR|32|33|希西家 与他祖先同睡，葬在 大卫 子孙陵墓的斜坡上。他死的时候， 犹大 众人和 耶路撒冷 的居民都向他致敬。他的儿子 玛拿西 接续他作王。
2CHR|33|1|玛拿西 登基的时候年十二岁，在 耶路撒冷 作王五十五年。
2CHR|33|2|他行耶和华眼中看为恶的事，效法耶和华在 以色列 人面前赶出的列国那些可憎的事。
2CHR|33|3|他重新建筑他父亲 希西家 所拆毁的丘坛，为诸 巴力 筑坛，造 亚舍拉 ，又敬拜天上的万象，事奉它们。
2CHR|33|4|他在耶和华殿中筑坛，耶和华曾指着这殿说：“我的名必永远在 耶路撒冷 。”
2CHR|33|5|他在耶和华殿的两个院子为天上的万象筑坛，
2CHR|33|6|并在 欣嫩子谷 使他的儿子经火，又观星象，行法术，行邪术，求问招魂的和行巫术的，多行耶和华眼中看为恶的事，惹他发怒。
2CHR|33|7|他在上帝殿内立雕刻的偶像；上帝曾对 大卫 和他儿子 所罗门 说：“我在 以色列 众支派中所选择的 耶路撒冷 和这殿，必立我的名，直到永远。
2CHR|33|8|只要 以色列 人谨守遵行我藉 摩西 吩咐他们的一切律法、律例、典章，我就不再使他们的脚挪移，离开我所赐给他们列祖之土地。”
2CHR|33|9|玛拿西 引诱 犹大 和 耶路撒冷 的居民行恶，比耶和华在 以色列 人面前所灭的列国更严重。
2CHR|33|10|耶和华警戒 玛拿西 和他的百姓，他们却不听。
2CHR|33|11|所以耶和华使 亚述 王的将领来攻击他们，用手铐铐住 玛拿西 ，用铜链锁住他，把他带到 巴比伦 去。
2CHR|33|12|他在急难的时候恳求耶和华－他的上帝，并在他列祖的上帝面前极其谦卑。
2CHR|33|13|他祈祷耶和华，耶和华就应允他，垂听他的祷告，使他归回 耶路撒冷 ，仍坐王位。 玛拿西 这才知道惟独耶和华是上帝。
2CHR|33|14|此后， 玛拿西 在 大卫城 外，从谷内 基训 西边直到 鱼门 口，建筑城墙，环绕 俄斐勒 ；这墙建得很高。他又在 犹大 各坚固城内设立将领。
2CHR|33|15|他除掉外邦人的神像与耶和华殿中的偶像，又将他在耶和华殿的山上和 耶路撒冷 所筑的各坛都拆毁，抛在城外。
2CHR|33|16|他重修耶和华的祭坛，在坛上献平安祭和感谢祭，并吩咐 犹大 人事奉耶和华－ 以色列 的上帝。
2CHR|33|17|百姓却仍在丘坛上献祭，不过，他们只献给耶和华－他们的上帝。
2CHR|33|18|玛拿西 其余的事和他向上帝的祷告，以及先见奉耶和华－ 以色列 上帝的名警戒他的话，看哪，都在《以色列诸王记》上。
2CHR|33|19|他的祷告，上帝怎样应允他，他未谦卑以前的一切罪愆过犯，以及在何处建筑丘坛，设立 亚舍拉 和雕刻的偶像，看哪，都写在 何赛 的书上。
2CHR|33|20|玛拿西 与他祖先同睡，葬在自己的宫中，他儿子 亚们 接续他作王。
2CHR|33|21|亚们 登基的时候年二十二岁，在 耶路撒冷 作王二年。
2CHR|33|22|他行耶和华眼中看为恶的事，效法他父亲 玛拿西 所行的，祭祀他父亲 玛拿西 所雕刻的一切偶像，事奉它们，
2CHR|33|23|但他不像他父亲 玛拿西 在耶和华面前那样谦卑下来。这 亚们 的罪越犯越大。
2CHR|33|24|他的臣仆背叛他，在宫里杀了他。
2CHR|33|25|但这地的百姓杀了所有背叛 亚们 王的人；这地的百姓立他儿子 约西亚 接续他作王。
2CHR|34|1|约西亚 登基的时候年八岁，在 耶路撒冷 作王三十一年。
2CHR|34|2|他行耶和华眼中看为正的事，行他祖先 大卫 所行的道，不偏左右。
2CHR|34|3|他作王第八年，尚且年轻，就寻求他祖先 大卫 的上帝。到了十二年，他开始洁净 犹大 和 耶路撒冷 ，除掉丘坛、 亚舍拉 、雕刻的像和铸造的像。
2CHR|34|4|众人在他面前拆毁诸 巴力 的坛，砍断坛上高高的香坛，又把 亚舍拉 和雕刻的像，以及铸造的像打碎成灰，撒在向偶像献祭之人的坟上，
2CHR|34|5|把祭司的骸骨烧在他们的坛上，洁净了 犹大 和 耶路撒冷 。
2CHR|34|6|他又在 玛拿西 、 以法莲 、 西缅 、 拿弗他利 各城和四围的废墟 ，
2CHR|34|7|拆毁祭坛，把 亚舍拉 和雕刻的像打碎成灰，砍断 以色列 全地所有的香坛。于是他回 耶路撒冷 去了。
2CHR|34|8|约西亚 王十八年，这地和殿洁净了之后，他派 亚萨利雅 的儿子 沙番 、 玛西雅 市长、 约哈斯 的儿子 约亚 史官去整修耶和华－他上帝的殿。
2CHR|34|9|他们去见 希勒家 大祭司，把奉到上帝殿的银子交给他；这银子是看守殿门的 利未 人从 玛拿西 、 以法莲 ，和 以色列 所有幸存的人，以及 犹大 、 便雅悯 众人和 耶路撒冷 的居民收来的。
2CHR|34|10|他们把这银子交给耶和华殿里督工的，由他们转交整修耶和华殿的工匠，
2CHR|34|11|就是交给木匠和石匠，好为 犹大 王所毁坏的殿，买凿成的石头和作钩子与栋梁的木料。
2CHR|34|12|这些人办事诚实，管理他们的是 利未 人 米拉利 的子孙 雅哈 和 俄巴底 ，又有 哥辖 人 撒迦利亚 和 米书兰 ；还有所有善于奏乐的 利未 人。
2CHR|34|13|他们监督扛抬的人，督导一切做各样工的人。 利未 人中也有作书记、官员、守卫的。
2CHR|34|14|他们把奉到耶和华殿的银子运出来的时候， 希勒家 祭司发现了耶和华藉 摩西 所传的律法书。
2CHR|34|15|希勒家 对 沙番 书记说：“我在耶和华殿里发现了律法书。” 希勒家 把书递给 沙番 。
2CHR|34|16|沙番 把书拿到王那里，又把这事回覆王说：“凡交给仆人的手所办的事，他们都办好了。
2CHR|34|17|耶和华殿里所发现的银子已经倒出来，交在督工和工匠的手里了。”
2CHR|34|18|沙番 书记又向王报告说：“ 希勒家 祭司递给我一卷书。” 沙番 就在王面前朗读那书。
2CHR|34|19|王听见律法的话，就撕裂衣服。
2CHR|34|20|王吩咐 希勒家 与 沙番 的儿子 亚希甘 、 米迦 的儿子 亚比顿 、 沙番 书记和王的臣仆 亚撒雅 ，说：
2CHR|34|21|“你们去，以所发现这书上的话，为我、为 以色列 和 犹大 幸存的人求问耶和华；因为我们的祖先没有遵守耶和华的话，没有照这书上所记的一切去做，耶和华的烈怒就倒在我们身上。”
2CHR|34|22|于是， 希勒家 和王的人 都去见 户勒大 女先知，她是掌管礼服的 沙龙 的妻子， 沙龙 是 哈斯拉 的孙子， 特瓦 的儿子。 户勒大 住在 耶路撒冷 第二区。他们向她说明来意。
2CHR|34|23|她对他们说：“耶和华－ 以色列 的上帝如此说：‘你们可以回覆那派你们来见我的人说，
2CHR|34|24|耶和华如此说：看哪，我必照着在 犹大 王面前所读那书上记载的一切诅咒，降祸于这地方和其上的居民。
2CHR|34|25|因为他们离弃我，向别神烧香，用他们手所做的一切惹我发怒，所以我的愤怒必倒在这地方，总不止息。’
2CHR|34|26|然而，派你们来求问耶和华的 犹大 王，你们要这样回覆他：‘耶和华－ 以色列 的上帝如此说：至于你所听见的话，
2CHR|34|27|就是听见我指着这地方和其上居民所说的话，你的心就软化，在我面前谦卑下来，撕裂衣服，向我哭泣，因此我应允你。这是耶和华说的。
2CHR|34|28|看哪，我必使你归到你祖先那里，平安地进入坟墓，我要降于这地方和其上居民的一切灾祸，你不会亲眼看见。’”他们就去把这话回覆王。
2CHR|34|29|王派人召集 犹大 和 耶路撒冷 的众长老来。
2CHR|34|30|王和 犹大 众人、 耶路撒冷 的居民、祭司、 利未 人，以及所有的百姓，无论大小，都一同上到耶和华的殿去；王把殿里所发现的约书上面一切的话读给他们听。
2CHR|34|31|王站在自己的位上，在耶和华面前立约，要尽心尽性跟从耶和华，遵守他的诫命、法度、律例，实行这书上所记这约的话；
2CHR|34|32|又使所有住 耶路撒冷 和 便雅悯 的人都服从这约。于是 耶路撒冷 的居民都遵行上帝，就是他们列祖之上帝的约。
2CHR|34|33|约西亚 从 以色列 各处把一切可憎之物尽都除掉，使 以色列 境内的人都事奉耶和华－他们的上帝。 约西亚 在世的日子，众人都跟从耶和华－他们列祖的上帝，总不离开。
2CHR|35|1|约西亚 在 耶路撒冷 向耶和华守逾越节。正月十四日，他们宰了逾越节的羔羊。
2CHR|35|2|王分派祭司各尽其职，又勉励他们办耶和华殿中的事。
2CHR|35|3|他对那归耶和华为圣、教导 以色列 众人的 利未 人说：“你们将圣约柜安放在 以色列 王 大卫 儿子 所罗门 建造的殿里，不必再用肩扛抬。现在你们要服事耶和华－你们的上帝和他的百姓 以色列 。
2CHR|35|4|你们应当按着父家，照着班次，遵照 以色列 王 大卫 和他儿子 所罗门 所写的，预备自己。
2CHR|35|5|要按着你们百姓的弟兄、父家的班次，侍立在圣所；每父家的班次中要有几个 利未 人。
2CHR|35|6|要宰逾越节的羔羊，将自己分别为圣，为你们的弟兄预备，好遵守耶和华藉 摩西 所吩咐的话。”
2CHR|35|7|约西亚 从群畜中赐给所有在场的百姓，三万只小绵羊和小山羊，三千头牛，作逾越节的祭物；这些都是出自王的产业。
2CHR|35|8|约西亚 的众领袖也乐意把祭牲给百姓、祭司和 利未 人；管理上帝殿的 希勒家 、 撒迦利亚 、 耶歇 ，把二千六百只羔羊和三百头牛给祭司作逾越节的祭物。
2CHR|35|9|利未 人的族长 歌楠雅 和他两个兄弟 示玛雅 、 拿坦业 ，与 哈沙比雅 、 耶利 、 约撒拔 ，把五千只羔羊和五百头牛给 利未 人作逾越节的祭物。
2CHR|35|10|这样，事奉的工作都安排好了，照王所吩咐的，祭司站在自己的位上， 利未 人按着班次侍立。
2CHR|35|11|他们宰了逾越节的羔羊，祭司从他们手里接过血来 洒出去； 利未 人剥皮，
2CHR|35|12|把燔祭拿走，再按着父家的班次分给众百姓，照 摩西 书上所写的献给耶和华；献牛也是这样。
2CHR|35|13|他们按着常例，用火烤逾越节的羔羊。至于其他的圣物，他们用盆，用锅，用釜煮了，速速地送给众百姓。
2CHR|35|14|然后他们为自己和祭司预备祭物，因为作祭司的 亚伦 子孙献燔祭和脂肪，直到晚上。所以 利未 人为自己和作祭司的 亚伦 子孙预备。
2CHR|35|15|歌唱的 亚萨 子孙，照着 大卫 、 亚萨 、 希幔 和王的先见 耶杜顿 所吩咐的，站在自己的位上。守门的看守各门，不用离开他们的职守，因为他们的弟兄 利未 人给他们预备。
2CHR|35|16|当日，一切供奉耶和华、守逾越节，以及在耶和华坛上献燔祭的事，都照 约西亚 王的吩咐预备好了。
2CHR|35|17|那时，在场的 以色列 人都守逾越节，又守除酵节七日。
2CHR|35|18|自从 撒母耳 先知的日子以来，在 以色列 中没有守过这样的逾越节， 以色列 诸王也没有守过像 约西亚 、祭司、 利未 人、所有住 犹大 和 以色列 的人，以及 耶路撒冷 居民所守的逾越节。
2CHR|35|19|这逾越节是 约西亚 作王十八年时守的。
2CHR|35|20|约西亚 为殿做完这一切事以后， 埃及 王 尼哥 上来，要攻打靠近 幼发拉底河 的 迦基米施 ； 约西亚 出去迎击他。
2CHR|35|21|他派使者来见 约西亚 ，说：“ 犹大 王啊，我跟你有什么相干呢？我今日来不是要攻打你，而是要攻打与我争战之家，并且上帝吩咐我从速行事。你不要干预与我同在的上帝，免得他毁灭你。”
2CHR|35|22|约西亚 却不转脸离开他，反而改装要与他打仗。他不听从上帝藉 尼哥 的口所说的话，就来到 米吉多 平原争战。
2CHR|35|23|弓箭手射中 约西亚 王。王对他的臣仆说：“我受了重伤，你们载我离开战场吧！”
2CHR|35|24|他的臣仆扶他下了战车，上了他的副座车，送他到 耶路撒冷 。他就死了，葬在他祖先的坟墓里。全 犹大 和 耶路撒冷 都哀悼 约西亚 。
2CHR|35|25|耶利米 为 约西亚 作哀歌，所有歌唱的男女也唱哀歌，追悼 约西亚 ，直到今日。他们在 以色列 中以此为定例；看哪，这些哀歌写在《哀歌书》上。
2CHR|35|26|约西亚 其余的事和他遵照耶和华律法上所记而行的善事，
2CHR|35|27|以及他自始至终所行的，看哪，都写在《以色列和犹大列王记》上。
2CHR|36|1|这地的百姓立 约西亚 的儿子 约哈斯 在 耶路撒冷 接续他父亲作王。
2CHR|36|2|约哈斯 登基的时候年二十三岁，在 耶路撒冷 作王三个月。
2CHR|36|3|埃及 王在 耶路撒冷 废了他，又罚这地一百他连得银子，一他连得金子。
2CHR|36|4|埃及 王 尼哥 立 约哈斯 的哥哥 以利雅敬 作 犹大 和 耶路撒冷 的王，给他改名叫 约雅敬 。 尼哥 却将他的弟弟 约哈斯 带到 埃及 去。
2CHR|36|5|约雅敬 登基的时候年二十五岁，在 耶路撒冷 作王十一年。他行耶和华－他上帝眼中看为恶的事。
2CHR|36|6|巴比伦 王 尼布甲尼撒 上来攻击他，用铜链锁着他，要把他带到 巴比伦 去。
2CHR|36|7|尼布甲尼撒 又将耶和华殿里的一些器皿带到 巴比伦 ，放在 巴比伦 自己的宫里 。
2CHR|36|8|约雅敬 其余的事和他所行可憎的事，以及发生在他身上的事，看哪，都写在《以色列和犹大列王记》上，他儿子 约雅斤 接续他作王。
2CHR|36|9|约雅斤 登基的时候年八岁 ，在 耶路撒冷 作王三个月十天，他行耶和华眼中看为恶的事。
2CHR|36|10|过了一年， 尼布甲尼撒 王差遣人将 约雅斤 和耶和华殿里宝贵的器皿带到 巴比伦 ，然后立 约雅斤 的叔父 西底家 作 犹大 和 耶路撒冷 的王。
2CHR|36|11|西底家 登基的时候年二十一岁，在 耶路撒冷 作王十一年。
2CHR|36|12|他行耶和华－他上帝眼中看为恶的事，没有谦卑听从 耶利米 先知所传达耶和华的话。
2CHR|36|13|尼布甲尼撒 王曾叫他指着上帝起誓，他却背叛，硬着颈项，内心顽固，不归向耶和华－ 以色列 的上帝。
2CHR|36|14|众祭司长和百姓也多多犯罪，效法列国一切可憎的事，玷污耶和华在 耶路撒冷 分别为圣的殿。
2CHR|36|15|耶和华－他们列祖的上帝因为爱惜自己的百姓和居所，一再差遣使者去警戒他们。
2CHR|36|16|他们却嘲笑上帝的使者，藐视他的话，讥诮他的先知，以致耶和华向他的百姓大发烈怒，甚至无法可救。
2CHR|36|17|所以，耶和华使 迦勒底 人的王来攻击他们，在他们圣殿里用刀杀了他们的壮丁，不怜悯他们的少男少女、老人长者。耶和华把所有的人都交在他手里。
2CHR|36|18|他把上帝殿里一切的大小器皿与耶和华殿里的财宝，以及王和众领袖的财宝，全都带到 巴比伦 去。
2CHR|36|19|迦勒底 人焚烧了上帝的殿，拆毁 耶路撒冷 的城墙，用火烧了城里所有的宫殿，毁坏了城里一切宝贵的器皿。
2CHR|36|20|凡脱离刀剑的幸存者， 迦勒底 王都掳到 巴比伦 去，作他和他子孙的仆婢，直到 波斯 国兴起。
2CHR|36|21|这就应验耶和华藉 耶利米 的口所说的话：地得享安息；在荒凉的日子，地就守安息，直到满了七十年。
2CHR|36|22|波斯 王 居鲁士 元年，耶和华为要应验藉 耶利米 的口所说的话，就激发 波斯 王 居鲁士 的心，使他下诏书通告全国，说：
2CHR|36|23|“ 波斯 王 居鲁士 如此说：耶和华－天上的上帝已将地上万国赐给我，又委派我在 犹大 的 耶路撒冷 为他建造殿宇。你们中间凡作他子民的可以上去，愿耶和华－他的上帝与他同在。”
