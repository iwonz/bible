JUDE|1|1|Iudas Iesu Christi servus frater autem Iacobi his qui in Deo Patre dilectis et Iesu Christo conservatis vocatis
JUDE|1|2|misericordia vobis et pax et caritas adimpleatur
JUDE|1|3|carissimi omnem sollicitudinem faciens scribendi vobis de communi vestra salute necesse habui scribere vobis deprecans supercertari semel traditae sanctis fidei
JUDE|1|4|subintroierunt enim quidam homines qui olim praescripti sunt in hoc iudicium impii Dei nostri gratiam transferentes in luxuriam et solum Dominatorem et Dominum nostrum Iesum Christum negantes
JUDE|1|5|commonere autem vos volo scientes semel omnia quoniam Iesus populum de terra Aegypti salvans secundo eos qui non crediderunt perdidit
JUDE|1|6|angelos vero qui non servaverunt suum principatum sed dereliquerunt suum domicilium in iudicium magni diei vinculis aeternis sub caligine reservavit
JUDE|1|7|sicut Sodoma et Gomorra et finitimae civitates simili modo exfornicatae et abeuntes post carnem alteram factae sunt exemplum ignis aeterni poenam sustinentes
JUDE|1|8|similiter et hii carnem quidem maculant dominationem autem spernunt maiestates autem blasphemant
JUDE|1|9|cum Michahel archangelus cum diabolo disputans altercaretur de Mosi corpore non est ausus iudicium inferre blasphemiae sed dixit imperet tibi Dominus
JUDE|1|10|hii autem quaecumque quidem ignorant blasphemant quaecumque autem naturaliter tamquam muta animalia norunt in his corrumpuntur
JUDE|1|11|vae illis quia via Cain abierunt et errore Balaam mercede effusi sunt et contradictione Core perierunt
JUDE|1|12|hii sunt in epulis suis maculae convivantes sine timore semet ipsos pascentes nubes sine aqua quae a ventis circumferuntur arbores autumnales infructuosae bis mortuae eradicatae
JUDE|1|13|fluctus feri maris despumantes suas confusiones sidera errantia quibus procella tenebrarum in aeternum servata est
JUDE|1|14|prophetavit autem et his septimus ab Adam Enoc dicens ecce venit Dominus in sanctis milibus suis
JUDE|1|15|facere iudicium contra omnes et arguere omnes impios de omnibus operibus impietatis eorum quibus impie egerunt et de omnibus duris quae locuti sunt contra eum peccatores impii
JUDE|1|16|hii sunt murmuratores querellosi secundum desideria sua ambulantes et os illorum loquitur superba mirantes personas quaestus causa
JUDE|1|17|vos autem carissimi memores estote verborum quae praedicta sunt ab apostolis Domini nostri Iesu Christi
JUDE|1|18|quia dicebant vobis quoniam in novissimo tempore venient inlusores secundum sua desideria ambulantes impietatum
JUDE|1|19|hii sunt qui segregant animales Spiritum non habentes
JUDE|1|20|vos autem carissimi superaedificantes vosmet ipsos sanctissimae vestrae fidei in Spiritu Sancto orantes
JUDE|1|21|ipsos vos in dilectione Dei servate
JUDE|1|22|et hos quidem arguite iudicatos
JUDE|1|23|illos vero salvate de igne rapientes aliis autem miseremini in timore odientes et eam quae carnalis est maculatam tunicam
JUDE|1|24|ei autem qui potest vos conservare sine peccato et constituere ante conspectum gloriae suae inmaculatos in exultatione
JUDE|1|25|soli Deo salvatori nostro per Iesum Christum Dominum nostrum gloria magnificentia imperium et potestas ante omne saeculum et nunc et in omnia saecula amen
