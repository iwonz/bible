3JOHN|1|1|我作长老的写信给亲爱的 该犹 ，就是我真心所爱的。
3JOHN|1|2|亲爱的，我愿你事事安宁，身体健康，正如你的心神安宁一样。
3JOHN|1|3|我非常欢喜，有弟兄到这里来，证实你对真理的忠诚，就是你按着真理而行。
3JOHN|1|4|我听见我的儿女按真理而行，我的欢喜没有比这个更大的。
3JOHN|1|5|亲爱的，你对弟兄，特别是对作客旅的弟兄所做的都是忠诚的。
3JOHN|1|6|他们在教会面前证实了你的爱；你若以对得起上帝的方式，为他们送行就好了；
3JOHN|1|7|因为他们是为基督的名 出外，并没有从未信的人接受什么。
3JOHN|1|8|所以，我们应当接待这样的人，好让我们与他们在真理上成为同工。
3JOHN|1|9|我曾写过一些东西给教会，但他们中间那好作领袖的 丢特腓 不接纳我们。
3JOHN|1|10|为此，我若去，要提起他所做的事，就是他用恶言攻击我们，还不满足，他自己不接纳弟兄，有人愿意接纳，他还阻止，并且把接纳弟兄的人赶出教会。
3JOHN|1|11|亲爱的，不要效法恶，只要效法善。行善的人属乎上帝；行恶的人未曾见过上帝。
3JOHN|1|12|低米丢 行善，有众人给他作见证，又有真理给他作见证，就是我们也给他作见证，你知道我们的见证是真的。
3JOHN|1|13|我还有许多事要写给你，却不愿意用笔墨来写给你，
3JOHN|1|14|但盼望很快见到你，我们好面对面谈论。
3JOHN|1|15|愿你平安！朋友们都向你问安。请你替我按著名字一一向朋友们问安。
