JOEL|1|1|耶和华的话临到 毗土珥 的儿子 约珥 。
JOEL|1|2|老年人哪，当听这话； 这地所有的居民哪，要侧耳而听。 在你们的日子， 或你们祖先的日子， 曾发生过这样的事吗？
JOEL|1|3|你们要将这事传与子， 子传与孙， 孙传与后代。
JOEL|1|4|剪虫吃剩的，蝗虫来吃； 蝗虫吃剩的，蝻子来吃； 蝻子吃剩的，蚂蚱 来吃。
JOEL|1|5|醉酒的人哪，要清醒，要哭泣； 好酒的人哪，都要为甜酒哀号， 因为酒从你们的口中断绝了。
JOEL|1|6|有一队蝗虫 ，强盛且不可数， 上来侵犯我的地； 它的牙齿如狮子的牙齿， 如母狮的大牙。
JOEL|1|7|它毁坏我的葡萄树， 撕裂我的无花果树， 剥光又丢弃，使枝条露白。
JOEL|1|8|你要像童女腰束麻布， 为她年少时的丈夫哀号。
JOEL|1|9|耶和华的殿中断绝素祭和浇酒祭， 事奉耶和华的祭司都悲哀。
JOEL|1|10|田荒凉，地悲哀； 因为五谷毁坏， 新酒枯竭， 新的油也缺乏。
JOEL|1|11|农夫啊，要惭愧； 修整葡萄园的啊，你们要哀号； 因为大麦、小麦与田间的庄稼全都毁了。
JOEL|1|12|葡萄树枯干， 无花果树衰残， 石榴树、棕树、苹果树， 田野一切的树木都枯干； 众人的喜乐尽都消逝。
JOEL|1|13|祭司啊，当束上麻布痛哭； 事奉祭坛的啊，要哀号； 事奉我上帝的啊，你们要来，披上麻布过夜， 因为在你们上帝的殿中不再有素祭和浇酒祭了。
JOEL|1|14|你们要使禁食的日子分别为圣， 宣告严肃会， 召集长老和这地所有的居民 来到耶和华－你们上帝的殿， 向耶和华哀求。
JOEL|1|15|哀哉，这日子！ 因为耶和华的日子临近， 好像毁灭从全能者来到。
JOEL|1|16|粮食不是在我们眼前断绝了吗？ 欢喜快乐不是从我们上帝的殿中止息了吗？
JOEL|1|17|种子在土块下朽烂， 仓荒凉，廪破坏， 因为五谷枯干了。
JOEL|1|18|牲畜哀鸣， 牛群混乱，因无草场， 羊群也受苦。
JOEL|1|19|耶和华啊，我向你求告， 因为有火吞噬野地的草场， 火焰烧尽田野的树木。
JOEL|1|20|田野的走兽切慕你， 因为溪水干涸， 火吞噬了野地的草场。
JOEL|2|1|你们要在 锡安 吹角， 在我的圣山发出警报。 这地所有的居民要发颤， 因为耶和华的日子快到， 已经临近了。
JOEL|2|2|那是黑暗、阴森的日子， 是密云、乌黑的日子， 如同黎明笼罩山岭。 有一队蝗虫，又大又强， 自古以来没有像这样的， 以后直到万代也必没有。
JOEL|2|3|它们前面有火吞噬， 后面有火焰烧尽。 它们未到以前，地如 伊甸园 ， 过去以后，却成了荒凉的旷野， 没有一样能躲避它们。
JOEL|2|4|它们形状如马， 奔跑如战马。
JOEL|2|5|响声如战车在山顶上跳动， 如火焰吞噬碎秸， 好像强大的军队摆阵备战。
JOEL|2|6|在它们面前，万民伤恸， 脸都变色。
JOEL|2|7|它们如勇士奔跑， 如战士攀登城墙， 各行于自己的道路， 不乱队伍；
JOEL|2|8|它们并不彼此推挤， 各行于自己的大道， 冲过防御 ， 并不停止。
JOEL|2|9|它们蹦上城， 跳上墙， 爬上房屋， 从窗户进来，如同盗贼。
JOEL|2|10|在它们面前， 地动天摇， 日月昏暗， 星宿无光。
JOEL|2|11|耶和华在他的军旅前出声， 他的队伍庞大， 遵行他命令的强盛。 耶和华的日子大而可畏， 谁能当得起呢？
JOEL|2|12|然而你们现在要禁食，哭泣，哀号， 一心归向我。 这是耶和华说的。
JOEL|2|13|你们要撕裂心肠， 不要撕裂衣服。 归向耶和华－你们的上帝， 因为他有恩惠，有怜悯， 不轻易发怒， 有丰盛的慈爱， 并且会改变心意， 不降那灾难。
JOEL|2|14|谁知道他也许会回心转意，留下余福， 就是献给耶和华－你们上帝的素祭和浇酒祭。
JOEL|2|15|你们要在 锡安 吹角， 使禁食的日子分别为圣， 宣告严肃会。
JOEL|2|16|聚集百姓，使会众自洁； 召集老年人， 聚集孩童和在母怀吃奶的； 使新郎出内室， 新娘离开洞房。
JOEL|2|17|事奉耶和华的祭司 要在走廊和祭坛间哭泣，说： “耶和华啊，求你顾惜你的百姓， 不要使你的产业受羞辱， 在列国中成为笑柄。 为何让人在万民中说 ‘他们的上帝在哪里’呢？”
JOEL|2|18|耶和华为自己的地发热心， 怜悯他的百姓。
JOEL|2|19|耶和华应允他的百姓说： “看哪，我要赏赐你们五谷、新酒和新的油， 使你们饱足， 我必不再使你们受列国的羞辱。
JOEL|2|20|我要使北方来的队伍远离你们， 将他们赶到干旱荒芜之地： 前队赶入东海， 后队赶入西海； 臭气上升，恶臭腾空。 耶和华果然行了大事！
JOEL|2|21|“土地啊，不要惧怕， 要欢喜快乐， 因为耶和华行了大事。
JOEL|2|22|田野的走兽啊，不要惧怕， 因为旷野的草已生长， 树木结果， 无花果树、葡萄树也都效力 。
JOEL|2|23|“ 锡安 的民哪，你们要欢喜， 要因耶和华－你们的上帝快乐； 因他赏赐你们合宜的秋雨 ， 为你们降下甘霖， 秋雨和春雨，和先前一样。
JOEL|2|24|“禾场充满五谷， 池中漫溢新酒和新的油。
JOEL|2|25|我差遣到你们中间的大军队， 就是蝗虫、蝻子、蚂蚱、剪虫， 那些年间所吃的，我要补还给你们。
JOEL|2|26|“你们必吃得饱足， 赞美耶和华－你们上帝的名， 他为你们行了奇妙的事。 我的百姓不致羞愧，直到永远。
JOEL|2|27|你们必知道我是在 以色列 中， 又知道我是耶和华－你们的上帝，没有别的。 我的百姓不致羞愧，直到永远。”
JOEL|2|28|“以后，我要将我的灵浇灌凡有血肉之躯的。 你们的儿女要说预言， 你们的老人要做异梦， 你们的少年要见异象。
JOEL|2|29|在那些日子， 我要将我的灵浇灌我的仆人和婢女。
JOEL|2|30|“我要在天上地下显出奇事，有血，有火，有烟柱。
JOEL|2|31|太阳要变为黑暗，月亮要变为血，这都在耶和华大而可畏的日子未到以前。
JOEL|2|32|那时，凡求告耶和华名的就必得救；因为照耶和华所说的，在 锡安山 ，在 耶路撒冷 将有逃脱的人。凡耶和华所召的 ，都在余民之列。”
JOEL|3|1|“看哪，在那些日子，到那个时候，我使 犹大 和 耶路撒冷 被掳之人归回的时候，
JOEL|3|2|我要聚集万民，带他们下到 约沙法谷 去，在那里我要为我百姓，我产业 以色列 的缘故，向万民施行审判；因为他们把我的百姓分散到列国，瓜分了我的土地，
JOEL|3|3|为我的百姓抽签，以男孩换取妓女，为喝酒卖掉女孩。
JOEL|3|4|“ 推罗 、 西顿 和 非利士 四境的人哪，你们与我何干？你们要报复我吗？若要报复我，我必使报应速速归到你们头上。
JOEL|3|5|你们夺取我的金银，把我珍贵的宝物带入你们的庙宇 ，
JOEL|3|6|并将 犹大 人和 耶路撒冷 人卖给 希腊 人 ，使他们远离自己的疆土。
JOEL|3|7|看哪，我必激发他们离开你们把他们卖去的地方，又必使报应归到你们头上。
JOEL|3|8|我要将你们的儿女卖到 犹大 人手中，他们必转卖给远方的国家 示巴 人。这是耶和华说的。”
JOEL|3|9|当在列国中宣告： 预备打仗， 激发勇士， 使所有战士上前来。
JOEL|3|10|要将犁头打成刀剑， 镰刀打成戈矛； 弱者要说：“我是勇士。”
JOEL|3|11|四围的列国啊， 要速速前来， 一同聚集。 耶和华啊， 求你使你的勇士降临。
JOEL|3|12|列国都当兴起， 上到 约沙法谷 ； 因为我必坐在那里， 审判四围的列国。
JOEL|3|13|挥镰刀吧！因为庄稼熟了； 来踩踏吧！因为醡酒池满了。 酒池已经满溢， 因为他们的罪恶甚大。
JOEL|3|14|在 断定谷 有许多许多的人， 因为耶和华的日子临近 断定谷 了。
JOEL|3|15|日月昏暗， 星宿无光。
JOEL|3|16|耶和华必从 锡安 吼叫， 从 耶路撒冷 出声， 天地就震动。 耶和华却要作他百姓的避难所， 作 以色列 人的保障。
JOEL|3|17|你们就知道我是耶和华－你们的上帝， 我住在 锡安 －我的圣山。 耶路撒冷 必成为圣； 陌生人不再从其中经过。
JOEL|3|18|在那日，大山要滴甜酒， 小山要流奶， 犹大 的溪河都有水流出； 必有泉源从耶和华的殿中流出， 滋润 什亭谷 。
JOEL|3|19|埃及 必定荒凉， 以东 成为荒凉的旷野， 因为他们向 犹大 人行残暴， 又因他们在本地流无辜人的血。
JOEL|3|20|但 犹大 必存到永远， 耶路撒冷 必存到万代。
JOEL|3|21|我要免除 流人血的罪， 是先前未曾免除的， 耶和华居住在 锡安 。
