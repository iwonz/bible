1KGS|1|1|大卫 王年纪老迈，虽然盖着外袍，仍不够暖和。
1KGS|1|2|臣仆对他说：“不如为我主我王找一个年轻的少女，侍立在王面前，照顾王，睡在王的怀中，好使我主我王得暖。”
1KGS|1|3|于是他们在 以色列 全境寻找美貌的少女，找到了一个 书念 女子 亚比煞 ，带到王那里。
1KGS|1|4|这少女极其美貌，她照顾王，伺候王，王却没有与她亲近。
1KGS|1|5|那时， 哈及 的儿子 亚多尼雅 妄自尊大，说：“我要作王”，就为自己预备座车、骑兵，又派五十人在他前头奔跑。
1KGS|1|6|他父亲从来没有责怪他，说：“你为何这么做？”他非常俊美，生在 押沙龙 之后。
1KGS|1|7|亚多尼雅 与 洗鲁雅 的儿子 约押 和 亚比亚他 祭司商议；他们就顺从 亚多尼雅 ，帮助他。
1KGS|1|8|但 撒督 祭司、 耶何耶大 的儿子 比拿雅 、 拿单 先知、 示每 、 利以 ，以及 大卫 自己的勇士 都不顺从 亚多尼雅 。
1KGS|1|9|亚多尼雅 在 隐．罗结 旁 琐希列 磐石那里献牛羊、肥犊为祭，请了他的众兄弟，就是王的众儿子，以及所有作王臣仆的 犹大 人。
1KGS|1|10|但他没有邀请 拿单 先知、 比拿雅 和勇士们，以及他的弟弟 所罗门 。
1KGS|1|11|拿单 对 所罗门 的母亲 拔示巴 说：“ 哈及 的儿子 亚多尼雅 作王了，你没有听见吗？我们的主 大卫 却不知道。
1KGS|1|12|现在，来，我给你出个主意，好保全你和你儿子 所罗门 的性命。
1KGS|1|13|你去，进到 大卫 王那里，对他说：‘我主我王啊，你不是曾向使女起誓说：你儿子 所罗门 必接续我作王，他必坐在我的王位上吗？ 亚多尼雅 怎么作了王呢？’
1KGS|1|14|看哪，你还在那里与王说话的时候，我会随后进去，证实你的话。”
1KGS|1|15|拔示巴 进入内室，到王那里。那时，王很老了， 书念 女子 亚比煞 正伺候着王。
1KGS|1|16|拔示巴 向王屈身下拜，王说：“你要什么？”
1KGS|1|17|她对王说：“我主啊，你曾向使女指着耶和华－你的上帝起誓：‘你儿子 所罗门 必接续我作王，他必坐在我的王位上。’
1KGS|1|18|现在，看哪， 亚多尼雅 作王了，你 ，我主我王却不知道。
1KGS|1|19|他献许多牛羊、肥犊为祭，请了王的众儿子和 亚比亚他 祭司，以及 约押 元帅，他却没有请王的仆人 所罗门 。
1KGS|1|20|但你 ，我主我王啊， 以色列 众人的眼目都仰望你，等你告诉他们，在我主我王之后谁坐你的王位。
1KGS|1|21|若不然，我主我王与祖先同睡的时候，我和我儿子 所罗门 必列为罪犯了。”
1KGS|1|22|看哪， 拔示巴 还与王说话的时候， 拿单 先知也进来了。
1KGS|1|23|有人奏告王说：“看哪， 拿单 先知来了。” 拿单 进到王面前，脸伏于地，向王叩拜。
1KGS|1|24|拿单 说：“我主我王，你果真说过‘ 亚多尼雅 必接续我作王，他要坐在我的王位上’吗？
1KGS|1|25|他今日下去，献了许多牛羊、肥犊为祭，请了王的众儿子和军官们，以及 亚比亚他 祭司；看哪，他们正在 亚多尼雅 面前吃喝，说：‘ 亚多尼雅 王万岁！’
1KGS|1|26|至于我，就是你的仆人，和 撒督 祭司、 耶何耶大 的儿子 比拿雅 、王的仆人 所罗门 ，他都没有请。
1KGS|1|27|这事果真出于我主我王吗？王却没有告诉仆人们，在我主我王之后谁坐你的王位。”
1KGS|1|28|大卫 王回答说：“召 拔示巴 到我这里来。” 拔示巴 就来，站在王面前。
1KGS|1|29|王起誓说：“我指着救我性命脱离一切苦难的永生的耶和华起誓。
1KGS|1|30|我既然指着耶和华－ 以色列 的上帝向你起誓说：你儿子 所罗门 必接续我作王，他必继承我坐在我的王位上，我今日必这样做。”
1KGS|1|31|于是， 拔示巴 屈身，脸伏于地，向王叩拜，说：“我主 大卫 王万岁！”
1KGS|1|32|大卫 王又说：“召 撒督 祭司、 拿单 先知、 耶何耶大 的儿子 比拿雅 到我这里来！”他们就都来到王面前。
1KGS|1|33|王对他们说：“要带领你们主的仆人，让我儿子 所罗门 骑我自己的骡子，送他下到 基训 。
1KGS|1|34|在那里， 撒督 祭司和 拿单 先知要膏他作 以色列 的王；你们也要吹角，说：‘ 所罗门 王万岁！’
1KGS|1|35|你们要跟随他上来，使他坐在我的王位上，他要接续我作王。我已立他作 以色列 和 犹大 的君王。”
1KGS|1|36|耶何耶大 的儿子 比拿雅 回应王说：“阿们！愿耶和华－我主我王的上帝这样说。
1KGS|1|37|耶和华怎样与我主我王同在，愿他照样与 所罗门 同在，使他的王位比我主 大卫 王的王位更大。”
1KGS|1|38|于是， 撒督 祭司、 拿单 先知、 耶何耶大 的儿子 比拿雅 ，以及 基利提 人和 比利提 人都下去，让 所罗门 骑上 大卫 王的骡子，送他到 基训 。
1KGS|1|39|撒督 祭司从帐幕中取了盛膏油的角来，膏 所罗门 。他们就吹角，众百姓都说：“ 所罗门 王万岁！”
1KGS|1|40|众百姓跟随他上来，吹着笛，大大欢呼，地被他们的声音震裂。
1KGS|1|41|亚多尼雅 和所有的宾客刚吃完，听见这声音； 约押 听见角声就说：“城中为何有这响声呢？”
1KGS|1|42|他正说话的时候，看哪， 亚比亚他 祭司的儿子 约拿单 来了。 亚多尼雅 说：“进来吧！你是个贤明的人，必是来报好消息的。”
1KGS|1|43|约拿单 回答 亚多尼雅 说：“我们的主 大卫 王已经立 所罗门 为王了！
1KGS|1|44|王派 撒督 祭司、 拿单 先知、 耶何耶大 的儿子 比拿雅 ，以及 基利提 人和 比利提 人和 所罗门 一起去，叫他骑上王的骡子。
1KGS|1|45|撒督 祭司和 拿单 先知已经在 基训 膏他作王了。他们从那里欢呼着上来，城都震动，这就是你们所听见的声音。
1KGS|1|46|所罗门 也已经登上国度的王位了。
1KGS|1|47|王的臣仆也来为我们的主 大卫 王祝福，说：‘愿上帝使 所罗门 的名比你的名更尊荣，使他的王位比你的王位更大。’王在床上屈身敬拜，
1KGS|1|48|王也这样说：‘耶和华－ 以色列 的上帝是应当称颂的，因他今日赏赐一个人坐在我的王位上，我也亲眼看见了。’”
1KGS|1|49|亚多尼雅 所有的宾客都战兢，起来，各走各路去了。
1KGS|1|50|亚多尼雅 惧怕 所罗门 ，就起来，去抓住祭坛的翘角。
1KGS|1|51|有人告诉 所罗门 说：“看哪， 亚多尼雅 惧怕 所罗门 王。看哪，他抓住祭坛的翘角，说：‘愿 所罗门 王先向我起誓，必不用刀杀死仆人。’”
1KGS|1|52|所罗门 说：“他若作贤明的人，连一根头发也不致落在地上；他若作恶，必要死亡。”
1KGS|1|53|于是 所罗门 王派人叫 亚多尼雅 从坛上下来，他就来向 所罗门 王下拜。 所罗门 对他说：“你回家去吧！”
1KGS|2|1|大卫 的死期临近了，就吩咐他儿子 所罗门 说：
1KGS|2|2|“我要走世人必走的路了。你当刚强，作大丈夫，
1KGS|2|3|遵守耶和华－你上帝所吩咐的，照着 摩西 律法上所写的行耶和华的道，谨守他的律例、诫命、典章、法度，好让你无论做什么，不拘往何处去，尽都亨通。
1KGS|2|4|耶和华必成就他所说关于我的话，说：‘你的子孙若谨慎自己的行为，尽心尽意凭信实行在我面前，就不断有人坐 以色列 的王位。’
1KGS|2|5|你也知道 洗鲁雅 的儿子 约押 向我所做的事，他对付 以色列 的两个元帅， 尼珥 的儿子 押尼珥 和 益帖 的儿子 亚玛撒 ，杀了他们。他在太平之时，如同战争一般，流这二人的血，把这战争的血染了他腰间束的带和脚上穿的鞋。
1KGS|2|6|所以你要照你的智慧去做，不让他白发安然下阴间。
1KGS|2|7|你当恩待 基列 人 巴西莱 的众儿子，请他们常与你同席吃饭，因为我躲避你哥哥 押沙龙 的时候，他们亲近我。
1KGS|2|8|看哪，在你这里有来自 巴户琳 的 便雅悯 人， 基拉 的儿子 示每 。我到 玛哈念 去的那日，他用狠毒的言语咒骂我。后来他却下 约旦河 迎接我，我就指着耶和华向他起誓说：‘我必不用刀杀死你。’
1KGS|2|9|但现在你不要以他为无罪。你是有智慧的人，必知道怎样待他，使他白发流血下阴间。”
1KGS|2|10|大卫 与他祖先同睡，葬在 大卫城 。
1KGS|2|11|大卫 作 以色列 王四十年：在 希伯仑 作王七年，在 耶路撒冷 作王三十三年。
1KGS|2|12|所罗门 坐他父亲 大卫 的王位，他的国度非常稳固。
1KGS|2|13|哈及 的儿子 亚多尼雅 到 所罗门 的母亲 拔示巴 那里， 拔示巴 问他说：“你是为平安来的吗？”他说：“为平安来的。”
1KGS|2|14|他又说：“我有话对你说。” 拔示巴 说：“你说吧。”
1KGS|2|15|亚多尼雅 说：“你知道这国原是归我的，全 以色列 也都期望我作王。然而，这国反归了我兄弟，因这国归了他是出乎耶和华。
1KGS|2|16|现在我有一件事求你，请你不要推辞。” 拔示巴 对他说：“你说吧。”
1KGS|2|17|他说：“求你请 所罗门 王把 书念 女子 亚比煞 赐我为妻，因他必不拒绝你。”
1KGS|2|18|拔示巴 说：“好，我必为你对王提说。”
1KGS|2|19|于是， 拔示巴 来到 所罗门 王那里，要为 亚多尼雅 说话。王起来迎接，向她下拜，然后坐在自己的位上，又为王的母亲设一座位，她就坐在王的右边。
1KGS|2|20|拔示巴 说：“我要向你提出一个小小的请求，请你不要回绝我。”王对她说：“母亲，请提出来，我必不回绝你。”
1KGS|2|21|拔示巴 说：“请你把 书念 女子 亚比煞 赐给你哥哥 亚多尼雅 为妻。”
1KGS|2|22|所罗门 王回答母亲说：“为何替 亚多尼雅 求 书念 女子 亚比煞 呢？可以为他求王国吧！他是我的兄长，不但为他，也为 亚比亚他 祭司和 洗鲁雅 的儿子 约押 求吧！ ”
1KGS|2|23|所罗门 王指着耶和华起誓说：“ 亚多尼雅 讲这话是自己送命，不然，愿上帝重重惩罚我。
1KGS|2|24|耶和华坚立我，使我坐在父亲 大卫 的王位上，照着他所应许的为我建立家室；现在我指着永生的耶和华起誓， 亚多尼雅 今日必被处死。”
1KGS|2|25|于是 所罗门 王派 耶何耶大 的儿子 比拿雅 去击杀 亚多尼雅 ，他就死了。
1KGS|2|26|王对 亚比亚他 祭司说：“你回 亚拿突 归自己的田地去吧！你本是该死的，但因你在我父亲 大卫 面前抬过主耶和华的约柜，又与我父亲同受一切苦难，所以我今日不杀死你。”
1KGS|2|27|所罗门 就革除 亚比亚他 ，不让他作耶和华的祭司。这就应验了耶和华在 示罗 论 以利 家所说的话。
1KGS|2|28|虽然 约押 没有拥护 押沙龙 ，却拥护了 亚多尼雅 ；这消息传到 约押 那里，他就逃到耶和华的帐幕，抓住祭坛的翘角。
1KGS|2|29|有人告诉 所罗门 王：“ 约押 逃到耶和华的帐幕，看哪，他在祭坛的旁边。” 所罗门 就派 耶何耶大 的儿子 比拿雅 ，说：“去，杀了他。”
1KGS|2|30|比拿雅 来到耶和华的帐幕，对 约押 说：“王这样吩咐：‘你出来吧！’”他说：“不，我要死在这里。” 比拿雅 就去回覆王，说：“ 约押 这样说，他这样回答我。”
1KGS|2|31|王对他说：“你可以照着他的话去做，杀了他，把他葬了，好叫 约押 流无辜人血的罪不归在我和我的父家。
1KGS|2|32|耶和华必使 约押 的血归到他自己头上，因为他击杀两个比他又公义又良善的人，就是 尼珥 的儿子 以色列 的元帅 押尼珥 和 益帖 的儿子 犹大 的元帅 亚玛撒 ，用刀杀了他们，我父亲 大卫 却不知道。
1KGS|2|33|这二人的血必归到 约押 和他后裔头上，直到永远；惟有 大卫 和他的后裔，以及他的家与王位，必从耶和华那里得平安，直到永远。”
1KGS|2|34|于是 耶何耶大 的儿子 比拿雅 上去，击杀 约押 ，杀死他，把他葬在旷野 约押 自己的家里。
1KGS|2|35|王就立 耶何耶大 的儿子 比拿雅 作元帅，代替 约押 ，又使 撒督 祭司代替 亚比亚他 。
1KGS|2|36|王派人召 示每 来，对他说：“你要在 耶路撒冷 为自己建造房屋，住在那里，不可从那里出来到任何地方去。
1KGS|2|37|你当确实知道，你何日出来过 汲沦溪 ，就必定死！你的血必归到自己头上。”
1KGS|2|38|示每 对王说：“这话很好！我主我王怎样说，仆人必照样做。”于是 示每 住在 耶路撒冷 许多日子。
1KGS|2|39|过了三年， 示每 的两个奴仆逃到 玛迦 的儿子 迦特 王 亚吉 那里去。有人告诉 示每 说：“看哪，你的奴仆在 迦特 。”
1KGS|2|40|示每 起来，备上驴，往 迦特 到 亚吉 那里去找他的奴仆，从 迦特 带他的奴仆回来。
1KGS|2|41|有人告诉 所罗门 ：“ 示每 出 耶路撒冷 到 迦特 去，又回来了。”
1KGS|2|42|王就派人召 示每 来，对他说：“我岂不是叫你指着耶和华起誓，并且警告你说‘你当确实知道，你何日出来到任何地方去，就必定死’吗？你也对我说：‘这话很好，我必听从。’
1KGS|2|43|你为何不遵守你对耶和华的誓言和我吩咐你的命令呢？”
1KGS|2|44|王又对 示每 说：“你向我父亲 大卫 所做的一切恶事，你自己心里都知道，耶和华必使你的罪恶归到你自己的头上。
1KGS|2|45|但 所罗门 王必蒙福， 大卫 的王位必在耶和华面前坚立，直到永远。”
1KGS|2|46|于是王吩咐 耶何耶大 的儿子 比拿雅 ，他就出去，击杀 示每 ， 示每 就死了。这样，国度在 所罗门 的手中巩固了。
1KGS|3|1|所罗门 与 埃及 王法老结亲，娶了法老的女儿，接她进入 大卫城 ，直等到建完了自己的宫和耶和华的殿，以及 耶路撒冷 周围的城墙。
1KGS|3|2|当那些日子，百姓仍在丘坛献祭，因为还没有为耶和华的名建殿。
1KGS|3|3|所罗门 爱耶和华，遵行他父亲 大卫 的律例，只是还在丘坛献祭烧香。
1KGS|3|4|所罗门 王到 基遍 ，在那里献祭，因为 基遍 有极大的丘坛。 所罗门 在那坛上献了一千祭牲为燔祭。
1KGS|3|5|在 基遍 ，耶和华夜间在梦中向 所罗门 显现；上帝说：“你愿我赐你什么，你可以求。”
1KGS|3|6|所罗门 说：“你曾向你仆人我父亲 大卫 大施慈爱，因为他用忠信、公义、正直的心行在你面前。你又为他存留大慈爱，赐他一个儿子坐在他的王位上，正如今日一样。
1KGS|3|7|现在，耶和华－我的上帝啊，你使仆人接续我父亲 大卫 作王；但我是幼小的孩子，不知道应当怎样出入。
1KGS|3|8|仆人住在你拣选的百姓中，这百姓之多，多得不可点，不可算。
1KGS|3|9|所以求你赐仆人善于了解的心，可以判断你的百姓，辨别是非。不然，谁能判断你这么多的百姓呢？”
1KGS|3|10|所罗门 因为求这事，就蒙主喜悦。
1KGS|3|11|上帝对他说：“你既然求这事，不为自己求寿、求富，也不求灭绝你仇敌的性命，只求能明辨，可以听讼，
1KGS|3|12|看哪，我会照你的话去做，看哪，我会赐你智慧和明辨的心，在你以前没有像你的，在你以后也没有兴起像你的。
1KGS|3|13|你没有求的，我也赐给你，就是富足、尊荣，使你在世一切的日子，列王中没有一个能比你的。
1KGS|3|14|你若遵行我的道，谨守我的律例、诫命，正如你父亲 大卫 所行的，我必使你长寿。”
1KGS|3|15|所罗门 醒了，看哪，是个梦。他就来到 耶路撒冷 ，站在耶和华的约柜前，献燔祭和平安祭，又为众臣仆摆设宴席。
1KGS|3|16|那时，有两个妓女来，站在王面前。
1KGS|3|17|一个妇人说：“我主啊，我和这妇人同住一屋。她在屋子里的时候，我生了一个孩子。
1KGS|3|18|我生了以后第三天，这妇人也生了。我们是一起的，屋子里除了我们二人之外，再没有别人在屋子里。
1KGS|3|19|夜间，这妇人的儿子死了，因为她压在她的儿子身上。
1KGS|3|20|她半夜起来，趁你使女睡着的时候，从我旁边把我儿子抱走，放在她怀里，又把她死的儿子放在我怀里。
1KGS|3|21|清早，我起来要给我的儿子吃奶，看哪，他死了；早晨我仔细察看他，看哪，他不是我所生的儿子。”
1KGS|3|22|另一个妇人说：“不！我的儿子是活的，你的儿子是死的。”但这一个说：“不！你的儿子是死的，我的儿子是活的。”她们就在王面前争吵。
1KGS|3|23|王说：“这妇人说：‘这是我的儿子，他是活的，你的儿子是死的。’那妇人说：‘不！你的儿子是死的，我的儿子是活的。’”
1KGS|3|24|王就说：“给我拿刀来！”人就把刀拿到王面前来。
1KGS|3|25|王说：“把活孩子劈成两半，一半给这妇人，一半给那妇人。”
1KGS|3|26|活孩子的母亲为自己的儿子心急如焚，对王说：“求我主把活孩子给那妇人吧，万不可杀死他！”那妇人说：“这孩子也不归我，也不归你，你们就劈了吧！”
1KGS|3|27|王回应说：“把活孩子给这妇人，万不可杀死他，因为这妇人是他的母亲。”
1KGS|3|28|全 以色列 听见王这样判断，就都敬畏王，因为他们看见他心中有上帝的智慧，能够断案。
1KGS|4|1|所罗门 作全 以色列 的王。
1KGS|4|2|这些是他的官员： 撒督 的儿子 亚撒利雅 作祭司，
1KGS|4|3|示沙 的两个儿子 以利何烈 、 亚希亚 作书记， 亚希律 的儿子 约沙法 作史官，
1KGS|4|4|耶何耶大 的儿子 比拿雅 作元帅， 撒督 和 亚比亚他 作祭司，
1KGS|4|5|拿单 的儿子 亚撒利雅 作宰相， 拿单 的儿子 撒布得 作祭司和王的顾问，
1KGS|4|6|亚希煞 作管家， 亚比大 的儿子 亚多尼兰 掌管服劳役的工人。
1KGS|4|7|所罗门 在全 以色列 有十二个官员，供给王和王室的食物，每年各人供给一个月。
1KGS|4|8|这些是他们的名字：在 以法莲 山区有 便．户珥 ；
1KGS|4|9|在 玛迦斯 、 沙宾 、 伯．示麦 、 以伦．伯．哈南 有 便．底甲 ；
1KGS|4|10|在 亚鲁泊 有 便．希悉 ，他管理 梭哥 和 希弗 全地；
1KGS|4|11|在 多珥 山冈 有 便．亚比拿达 ，他娶了 所罗门 的女儿 她法 为妻；
1KGS|4|12|在 他纳 和 米吉多 ，以及靠近 撒拉他拿 、 耶斯列 下边的 伯．善 全地，从 伯．善 到 亚伯．米何拉 直到 约缅 的另一边有 亚希律 的儿子 巴拿 ；
1KGS|4|13|在 基列 的 拉末 有 便．基别 ，他管理在 基列 的 玛拿西 子孙 睚珥 的城镇， 巴珊 的 亚珥歌伯 地的六十座大城，各有城墙和铜闩；
1KGS|4|14|在 玛哈念 有 易多 的儿子 亚希拿达 ；
1KGS|4|15|在 拿弗他利 有 亚希玛斯 ，他也娶了 所罗门 的一个女儿 巴实抹 为妻；
1KGS|4|16|在 亚设 和 亚禄 有 户筛 的儿子 巴拿 ；
1KGS|4|17|在 以萨迦 有 帕路亚 的儿子 约沙法 ；
1KGS|4|18|在 便雅悯 有 以拉 的儿子 示每 ；
1KGS|4|19|在 基列 地，就是 亚摩利 王 西宏 和 巴珊 王 噩 之地，有 乌利 的儿子 基别 ，他一个官员管理这地 。
1KGS|4|20|犹大 人和 以色列 人如同海边的沙那样多，都吃喝快乐。
1KGS|4|21|所罗门 统治诸国，从 大河 到 非利士 地，直到 埃及 的边界。 所罗门 在世的日子，这些国都向他进贡，服事他。
1KGS|4|22|所罗门 每日所用的食物：三十歌珥细面，六十歌珥粗面，
1KGS|4|23|十头肥牛，二十头草场的牛，一百只羊，还有鹿、羚羊、麃子，以及肥禽。
1KGS|4|24|所罗门 管理整个 大河 西边，从 提弗萨 直到 迦萨 ，以及 大河 西边的诸王，属他的四境尽都平安。
1KGS|4|25|所罗门 在世的日子，从 但 到 别是巴 ， 犹大 和 以色列 各人都在自己的葡萄树下和无花果树下安然居住。
1KGS|4|26|所罗门 拥有给战车用的四万个 马棚，还有一万二千名骑兵。
1KGS|4|27|这些官员各按自己的月份供给 所罗门 王，以及一切与他同席之人的食物，一无所缺。
1KGS|4|28|他们各按其分，把给马与快马吃的大麦和干草送到指定的地方去。
1KGS|4|29|上帝赐给 所罗门 极大的智慧和聪明，以及宽阔的心，如同海边的沙。
1KGS|4|30|所罗门 的智慧超过所有东方人的智慧，和 埃及 人一切的智慧。
1KGS|4|31|他的智慧胜过万人，胜过 以斯拉 人 以探 ，以及 玛曷 的儿子 希幔 、 甲各 、 达大 。他的名声传遍四围的列国。
1KGS|4|32|他作箴言三千句，诗歌一千零五首。
1KGS|4|33|他讲论草木，从 黎巴嫩 的香柏树直到墙上长的牛膝草，又讲论飞禽、走兽、爬行动物和鱼类。
1KGS|4|34|地上凡曾听过他智慧的君王，都派人来；万民都有人来听 所罗门 的智慧。
1KGS|5|1|推罗 王 希兰 是 大卫 平生的好友。 希兰 听见 以色列 人膏 所罗门 接续他父亲作王，就派臣仆到他那里。
1KGS|5|2|所罗门 也派人到 希兰 那里，说：
1KGS|5|3|“你知道我父亲 大卫 因四围的战争，不能为耶和华－他上帝的名建殿，直等到耶和华使仇敌都服在他脚下。
1KGS|5|4|现在耶和华－我的上帝使我四围太平，没有仇敌，没有灾祸。
1KGS|5|5|看哪，我吩咐要为耶和华－我上帝的名建殿，是照耶和华向我父亲 大卫 说的：‘我必使你儿子接续你，坐你的王位，他必为我的名建殿。’
1KGS|5|6|现在，请吩咐人在 黎巴嫩 为我砍伐香柏木，我的仆人必帮助你的仆人。至于你仆人的工钱，我必照你所定的给你。你知道，在我们中间没有人像 西顿 人那样擅长砍伐树木。”
1KGS|5|7|希兰 听见 所罗门 的话，就很高兴，说：“今日耶和华是应当称颂的，因为他赐给 大卫 一个有智慧的儿子，治理这众多的百姓。”
1KGS|5|8|希兰 送信给 所罗门 ，说：“你派人向我所提的那事，我已听见了；论到香柏木和松木，我必照你一切的心愿去做。
1KGS|5|9|我的仆人必把这木料从 黎巴嫩 运到海里，我会把它们扎成筏子浮在海上，运到你告诉我的地方，在那里拆开，你就可以收取；你也要照我的心愿做，把食物给我的家。”
1KGS|5|10|于是 希兰 照 所罗门 的心愿，给他香柏木和松木；
1KGS|5|11|所罗门 给 希兰 二万歌珥麦子，二十歌珥 捣成的油，作他家的食物。 所罗门 每年都是这样给 希兰 。
1KGS|5|12|耶和华照着所应许的赐智慧给 所罗门 。 希兰 与 所罗门 和平相处，二人彼此立约。
1KGS|5|13|所罗门 王从全 以色列 挑取服劳役的人，征来的人有三万，
1KGS|5|14|派他们轮流每月一万人上 黎巴嫩 去；一个月在 黎巴嫩 ，两个月在家里。 亚多尼兰 管理他们。
1KGS|5|15|所罗门 有七万扛抬的，八万在山上凿石头的。
1KGS|5|16|此外， 所罗门 有三千三百个监督工作的官长，监管百姓做工。
1KGS|5|17|王下令，他们就凿出又大又贵重的石头来，用以立殿的根基。
1KGS|5|18|所罗门 的工匠和 希兰 的工匠，以及 迦巴勒 人，把石头凿好，预备了木料和石头来建殿。
1KGS|6|1|以色列 人出 埃及 地后四百八十年， 所罗门 作 以色列 王第四年西弗月，就是二月，他开工建造耶和华的殿。
1KGS|6|2|所罗门 王为耶和华所建的殿，长六十肘，宽二十肘，高三十肘。
1KGS|6|3|殿的正堂前走廊长二十肘，与殿的宽度一样，殿前宽十肘；
1KGS|6|4|他为殿做了有框嵌壁式的窗户。
1KGS|6|5|靠着殿墙，围着外殿和内殿的墙，周围建造了厢房；
1KGS|6|6|下层宽五肘，中层宽六肘，第三层宽七肘。他在殿墙的周围造坎，免得梁木插入殿墙里。
1KGS|6|7|殿是用山中凿成的石头建的，所以建殿的时候，锤子、斧子和别样铁器的响声都没有听见。
1KGS|6|8|在殿右边当中的厢房有门，可以从螺旋梯上到中层，再从中层上到第三层。
1KGS|6|9|所罗门 完成殿的建造。他用香柏木作梁木和横板，遮盖殿顶。
1KGS|6|10|靠着整个殿所造的厢房，每层高五肘，香柏木的梁板搁在殿的墙坎上。
1KGS|6|11|耶和华的话临到 所罗门 ，说：
1KGS|6|12|“论到你所建的这殿，你若遵行我的律例，谨守我的典章，遵从我的一切诫命，行在其中，我必向你应验我所应许你父亲 大卫 的话。
1KGS|6|13|我必住在 以色列 人中间，并不丢弃我的百姓 以色列 。”
1KGS|6|14|所罗门 完成殿的建造。
1KGS|6|15|他用香柏木板建造殿的内墙，从殿的地到墙顶 都贴上木板，又用松木板铺地。
1KGS|6|16|他在殿的后部建了一间内殿，长二十肘，从地到墙 用香柏木板，作为至圣所。
1KGS|6|17|殿，就在内殿的前面 ，长四十肘。
1KGS|6|18|殿里一点石头都不显露，一概用香柏木遮蔽；香柏木上刻着野瓜和绽开的花。
1KGS|6|19|他在殿的中间预备内殿，在那里安放耶和华的约柜。
1KGS|6|20|内殿 长二十肘，宽二十肘，高二十肘，都贴上纯金。他又用香柏木做坛。
1KGS|6|21|所罗门 用纯金贴殿内，又用金链子挂在内殿前，内殿也贴上金子。
1KGS|6|22|整个殿都贴上金子，直到贴满；内殿前的整个坛，也都包上金子。
1KGS|6|23|他在内殿里用橄榄木做两个基路伯，各高十肘。
1KGS|6|24|这基路伯的一个翅膀长五肘，另一个翅膀长五肘，从一个翅膀尖到另一个翅膀尖共有十肘；
1KGS|6|25|第二个基路伯也是十肘；两个基路伯的尺寸、形状都一样。
1KGS|6|26|这一个基路伯高十肘，第二个基路伯也是如此。
1KGS|6|27|他把两个基路伯安在内殿中间。基路伯的翅膀是张开的，这基路伯的一个翅膀挨着这边的墙，第二个基路伯的一个翅膀挨着那边的墙，向内的两个翅膀在殿中间彼此相接。
1KGS|6|28|二基路伯都包上金子。
1KGS|6|29|殿周围的墙上全都刻着基路伯、棕树和绽开的花，内外都是如此。
1KGS|6|30|殿的地板都贴上金子，内外都是如此。
1KGS|6|31|他用橄榄木制造内殿的入口、门楣和五边形的门柱。
1KGS|6|32|在橄榄木做的两门扇上刻着基路伯、棕树和绽开的花，都贴上金子。基路伯和棕树上也洒上金子。
1KGS|6|33|他又为外殿的入口，用橄榄木制造门柱，是四边形的。
1KGS|6|34|他用松木做两扇门。这一扇有两叶摺叠，第二扇也有两叶 摺叠。
1KGS|6|35|上面刻着基路伯、棕树和绽开的花，雕刻物都均匀地贴上金子。
1KGS|6|36|他又用三层凿成的石头、香柏木一层建造内院。
1KGS|6|37|所罗门 在位第四年西弗月，立了耶和华殿的根基。
1KGS|6|38|到十一年布勒月，就是八月，殿和一切属殿的都按着样式造成。他建殿共用了七年。
1KGS|7|1|所罗门 为自己建造宫殿，十三年方才建成整座宫殿。
1KGS|7|2|他建造 黎巴嫩林宫 ，长一百肘，宽五十肘，高三十肘，有四行香柏木柱，柱上有香柏木横梁；
1KGS|7|3|厢房以上覆盖着香柏木，在四十五根柱子之上，每行十五根。
1KGS|7|4|窗户有三排，三排的窗与窗相对。
1KGS|7|5|所有的门和门柱都有四方形的框，共有三行，彼此相对。
1KGS|7|6|他建造有柱子的厅，长五十肘，宽三十肘。在这前面有走廊，前面有柱子和顶盖 。
1KGS|7|7|他又建造一个有座位的厅，就是审判厅，他在那里审判；这厅的地板从这边到那边都铺上香柏木。
1KGS|7|8|厅后面的院内有 所罗门 自己住的宫殿，都用同样的建造方式。 所罗门 又为所娶法老的女儿建造一座宫，建造方式与这厅一样。
1KGS|7|9|建造这一切所用的石头都是贵重的，按着尺寸凿成，用锯子里外锯齐；从根基直到房檐，从外头直到大院，都是如此。
1KGS|7|10|根基是贵重的大石头，有长十肘的，有长八肘的；
1KGS|7|11|上面有香柏木和按着尺寸凿成的贵重石头。
1KGS|7|12|大院周围有凿成的石头三层、香柏木板一层，都照耶和华殿的内院和殿的走廊的样式。
1KGS|7|13|所罗门 王派人从 推罗 把 户兰 接来。
1KGS|7|14|他是 拿弗他利 支派中一个寡妇的儿子，父亲是 推罗 人，是作铜匠的。 户兰 满有智慧、聪明、技能，善作各样的铜器。他来到 所罗门 王那里，为王做一切的工。
1KGS|7|15|户兰 制造两根铜柱，一根高十八肘，第二根柱子用绳子量，周围是十二肘 ；
1KGS|7|16|他做了两个柱顶安在柱上，是用铜铸造的，一个柱顶高五肘，第二个柱顶也高五肘。
1KGS|7|17|柱子顶上有装饰的网子和编成的链子，一个柱顶有七个，第二个柱顶也有七个。
1KGS|7|18|他做了柱子 ，第一根柱子的柱顶上，周围有两行网子在柱子 上面遮盖柱顶，第二根柱顶也是这样做。
1KGS|7|19|走廊柱子顶上的柱顶高四肘，刻着百合花。
1KGS|7|20|两根柱子上面有柱顶，柱顶靠近网子的圆凸面上，有石榴的行列环绕着，共二百个，第二个柱顶也是如此。
1KGS|7|21|他把两根柱子立在殿的走廊前：右边立一根，起名叫 雅斤 ；左边立一根，起名叫 波阿斯 。
1KGS|7|22|柱顶上刻着百合花。这样，柱子的工程就完毕了。
1KGS|7|23|他又铸一个铜海，周围是圆的，直径十肘，高五肘，用绳子量周围是三十肘。
1KGS|7|24|铜海边缘下面的周围有野瓜的形状，每肘十个，共两行，绕着铜海，是造铜海的时候铸上去的。
1KGS|7|25|铜海安在十二头铜牛上：三头向北，三头向西，三头向南，三头向东。铜海安在牛上，牛尾都向内。
1KGS|7|26|铜海厚一掌，边如杯边，像百合花，容量是二千罢特。
1KGS|7|27|他用铜制造十个盆座，每座长四肘，宽四肘，高三肘。
1KGS|7|28|铜座的造法是这样：周围各有嵌边，嵌边装在框架中。
1KGS|7|29|装在框架中的嵌边上有狮子和牛，以及基路伯。框架上有小座，狮子和牛的上面和下面有锤成的花纹浮雕。
1KGS|7|30|每座有四个铜轮和铜轴，它有四个支架在盆以下，这些支架是铸成的，各边都有花纹。
1KGS|7|31|它的口在柱顶里，向上高一肘，口是圆的，做法如座一样，直径是一肘半，口上也有雕工。嵌边是方形的，不是圆的。
1KGS|7|32|四个轮子在嵌边以下，轮轴与座相连，每轮高一肘半。
1KGS|7|33|轮的样式如同车的轮子；轴、辋、辐、毂都是铸成的。
1KGS|7|34|每个座四边有四个盆形的支架，这些支架是与座从一整块铸成的。
1KGS|7|35|座顶有圆架，高半肘；座顶有支柱和嵌边，是与座从一整块铸成的。
1KGS|7|36|他在支柱和嵌边上，每个空处刻上基路伯、狮子和棕树，周围有花纹。
1KGS|7|37|他按照这样的做法造了十个盆座，它们的铸法、尺寸、样式全都相同。
1KGS|7|38|他又造十个铜盆，每盆的容量四十罢特，直径四肘。在十个座上，每座安设一盆。
1KGS|7|39|他把五个安置在殿的右边，五个安置在殿的左边，又把铜海安置在殿的右旁，在东南边。
1KGS|7|40|户兰 又造了盆、铲子和盘子。这样， 户兰 为 所罗门 王做完了耶和华殿一切的工：
1KGS|7|41|两根柱子和柱子顶上两个如碗的柱顶，以及盖着如碗柱顶的两个网子；
1KGS|7|42|四百个石榴，安在两个网子上，每网两行石榴，盖着柱子上面两个如碗的柱顶；
1KGS|7|43|十个盆座和其上的十个盆；
1KGS|7|44|铜海和其下的十二头牛；
1KGS|7|45|盆、铲子、盘子。 户兰 给 所罗门 王为耶和华殿造的这一切器皿都是用光亮的铜，
1KGS|7|46|是王在 约旦 平原、 疏割 和 撒拉但 中间的泥巴地铸成的。
1KGS|7|47|所罗门 允许这一切器皿不过秤，因为所用的铜太多，重量无法计算。
1KGS|7|48|所罗门 又为耶和华的殿造了各样的器皿：金坛和献供饼的金供桌；
1KGS|7|49|内殿前的纯金灯台，右边五个，左边五个，以及其上的花、灯盏、灯剪，都是金的；
1KGS|7|50|纯金的杯、钳子、盘子、勺子 、火盆，以及圣殿的最里面，就是至圣所的门枢和外殿的门枢，都是金的。
1KGS|7|51|所罗门 王做完了耶和华殿一切的工，就把他父亲 大卫 分别为圣的金银和器皿都带来，放在耶和华殿的库房里。
1KGS|8|1|那时， 所罗门 召集 以色列 的长老、各支派的领袖和 以色列 人的族长到 耶路撒冷 ， 所罗门 王那里，要把耶和华的约柜从 大卫城 ，就是 锡安 ，接上来。
1KGS|8|2|以他念月，就是七月，在节期时，所有的 以色列 人都聚集到 所罗门 王那里。
1KGS|8|3|以色列 众长老一来到，祭司就抬起约柜。
1KGS|8|4|祭司和 利未 人将耶和华的约柜请上来，又把会幕和会幕一切的圣器皿都带上来。
1KGS|8|5|所罗门 王和聚集到他那里的 以色列 全会众一同在约柜前献牛羊为祭，多得不可胜数，无法计算。
1KGS|8|6|祭司将耶和华的约柜请进内殿，就是至圣所，安置在两个基路伯的翅膀底下约柜的地方。
1KGS|8|7|基路伯张开翅膀在约柜上面的地方，从上面遮住约柜和抬柜的杠。
1KGS|8|8|这杠很长，从内殿前的圣所可以看见杠头，从外面却看不见。这杠直到今日还在那里。
1KGS|8|9|约柜里没有别的，只有两块石版，就是 以色列 人出 埃及 地，耶和华与他们立约的时候， 摩西 在 何烈山 放在那里的。
1KGS|8|10|祭司从圣所出来的时候，有云充满耶和华的殿，
1KGS|8|11|祭司因云彩的缘故不能站立供职，因为耶和华的荣光充满了耶和华的殿。
1KGS|8|12|那时， 所罗门 说： “耶和华曾说要住在幽暗之处 。
1KGS|8|13|我的确为你建了一座雄伟的殿宇， 作为你永远居住的地方。”
1KGS|8|14|王转过脸来为 以色列 全会众祝福， 以色列 全会众都站立。
1KGS|8|15|所罗门 说：“耶和华－ 以色列 的上帝是应当称颂的！因他亲口向我父 大卫 应许的，也亲手成就了；他曾说：
1KGS|8|16|‘自从那日我领我百姓 以色列 出 埃及 以来，我未曾在 以色列 各支派中选择一城，在那里为我的名建造殿宇，但我拣选 大卫 治理我的百姓 以色列 。’
1KGS|8|17|我父 大卫 的心意是要为耶和华－ 以色列 上帝的名建殿。
1KGS|8|18|耶和华却对我父 大卫 说：‘你有心为我的名建殿，这心意是好的；
1KGS|8|19|但你不可建殿，惟有你亲生的儿子才可为我的名建殿。’
1KGS|8|20|现在耶和华实现了他所应许的话，使我接续我父 大卫 坐 以色列 的王位，正如耶和华所说的，我也为耶和华－ 以色列 上帝的名建造了这殿。
1KGS|8|21|我也在那里为约柜预备一处。约柜那里有耶和华的约，就是他领我们列祖出 埃及 地的时候，与他们所立的约。”
1KGS|8|22|所罗门 当着 以色列 全会众，站在耶和华的坛前，向天举手，
1KGS|8|23|说：“耶和华－ 以色列 的上帝啊，天上地下没有神明可与你相比！你向那些尽心行在你面前的仆人守约施慈爱，
1KGS|8|24|这约是你向你仆人 大卫 守的，是你应许他的。你亲口应许，亲手成就，正如今日一样。
1KGS|8|25|耶和华－ 以色列 的上帝啊，你向你仆人我父 大卫 应许说：‘你的子孙若谨慎自己的行为，在我面前行事像你所行的一样，就不断有人在我面前坐 以色列 的王位。’现在求你信守这话。
1KGS|8|26|以色列 的上帝啊，现在求你成就向你仆人我父 大卫 所应许的话。
1KGS|8|27|“上帝果真住在地上吗？看哪，天和天上的天尚且不足容纳你，何况我所建的这殿呢？
1KGS|8|28|惟求耶和华－我的上帝垂顾仆人的祷告祈求，俯听仆人今日在你面前的祈祷呼求。
1KGS|8|29|愿你的眼目昼夜看顾这殿，就是你说要作为你名的居所；求你垂听祷告，你仆人向此处的祷告。
1KGS|8|30|你仆人和你百姓 以色列 向此处祈祷的时候，求你在你天上的居所垂听，垂听而赦免。
1KGS|8|31|“人若得罪邻舍，有人强迫他，要他起誓，他来到这殿，在你的坛前起誓，
1KGS|8|32|求你在天上垂听、处理，向你的仆人施行审判，定恶人有罪，照他所行的报应在他头上；定义人为义，照他的义赏赐他。
1KGS|8|33|“你的百姓 以色列 若得罪你，败在仇敌面前，却又归向你，宣认你的名，在这殿里向你祈求祷告，
1KGS|8|34|求你在天上垂听，赦免你百姓 以色列 的罪，使他们归回你赐给他们列祖的地。
1KGS|8|35|“你的百姓若得罪了你，你使天闭塞不下雨；他们若向此处祷告，宣认你的名，因你的惩罚而离开他们的罪，
1KGS|8|36|求你在天上垂听，赦免你仆人你百姓 以色列 的罪，将当行的善道教导他们，并降雨在你的地，就是你赐给你百姓为业之地。
1KGS|8|37|“这地若有饥荒、瘟疫、焚风 、霉烂、蝗虫、蚂蚱，或有仇敌围困这地的 城门，无论遭遇什么灾祸疾病，
1KGS|8|38|你的百姓 以色列 ，或众人或一人，内心知道有祸，向这殿举手，无论祈求什么，祷告什么，
1KGS|8|39|求你在天上你的居所垂听、赦免、处理。因为你知道人心，惟有你知道世人的心，求你照各人所行的一切待他们，
1KGS|8|40|使他们在你赐给我们列祖的土地上一生一世敬畏你。
1KGS|8|41|“论到不属你百姓 以色列 的外邦人，若为你的名从远方而来，
1KGS|8|42|他们因听见你的大名和大能的手，以及伸出来的膀臂，来向这殿祷告，
1KGS|8|43|求你在天上你的居所垂听，照着外邦人向你所求的一切而行，使地上万民都认识你的名，敬畏你，像你的百姓 以色列 一样，又使他们知道我所建造的是称为你名下的殿。
1KGS|8|44|“你的百姓若奉你的派遣出去，无论往何处与仇敌争战，他们若向耶和华所选择的城，以及我为你名所建造的这殿祷告，
1KGS|8|45|求你在天上垂听他们的祷告祈求，为他们伸张正义。
1KGS|8|46|“你的百姓若得罪你，因为没有人不犯罪，你向他们发怒，把他们交在仇敌面前，掳他们的人把他们带到仇敌之地，或远或近，
1KGS|8|47|他们若在被掳之地那里回心转意，在掳掠者之地悔改，向你恳求说：‘我们有罪了，我们悖逆了，我们作恶了’；
1KGS|8|48|他们若在掳他们的仇敌之地尽心尽性归向你，又向自己的地，就是你赐给他们列祖的地和你所选择的城，以及我为你名所建造的这殿祷告，
1KGS|8|49|求你在天上你的居所垂听他们的祷告祈求，为他们伸张正义，
1KGS|8|50|饶恕得罪你的子民，赦免他们向你所犯一切的过犯，使他们在掳他们的人面前蒙怜悯。
1KGS|8|51|因为他们是你的子民，你的产业，是你从 埃及 ，从铁炉中领出来的。
1KGS|8|52|愿你的眼目看顾仆人和你百姓 以色列 的祈求；他们无论何时向你呼求，愿你垂听。
1KGS|8|53|主耶和华啊，你将他们从地上万民中分别出来作你的产业，是照着你领我们列祖出 埃及 的时候，藉你仆人 摩西 所应许的。”
1KGS|8|54|所罗门 在耶和华的坛前屈膝跪着，向天举手；他在耶和华面前祷告祈求完毕的时候，就起来，
1KGS|8|55|站着，大声为 以色列 全会众祝福，说：
1KGS|8|56|“耶和华是应当称颂的！因为他照着一切所应许的赐平安给他的百姓 以色列 ，凡藉他仆人 摩西 应许赐福的话，一句都没有落空。
1KGS|8|57|愿耶和华－我们的上帝与我们同在，像与我们列祖同在一样，不撇下我们，不丢弃我们，
1KGS|8|58|使我们的心归向他，遵行他一切的道，谨守他吩咐我们列祖的诫命、律例、典章。
1KGS|8|59|愿我在耶和华面前祈求的这些话，昼夜靠近耶和华－我们的上帝，好让他每日为他仆人和他百姓 以色列 伸张正义，
1KGS|8|60|使地上的万民都知道惟独耶和华是上帝，没有别的了。
1KGS|8|61|所以你们当向耶和华－我们的上帝存纯正的心，遵行他的律例，谨守他的诫命，如同今日一样。”
1KGS|8|62|王和全 以色列 一同在耶和华面前献祭。
1KGS|8|63|所罗门 向耶和华献平安祭，二万二千头牛，十二万只羊。这样，王和全 以色列 为耶和华的殿行了奉献之礼。
1KGS|8|64|当日，王因耶和华殿前的铜坛太小，容不下燔祭、素祭和平安祭牲的脂肪，就将耶和华殿前院子的中间分别为圣，在那里献燔祭、素祭和平安祭牲的脂肪。
1KGS|8|65|那时 所罗门 守节，从 哈马口 直到 埃及 溪谷的 以色列 众人都与他同在一起，成了一个盛大的会，在耶和华－我们的上帝面前七日又七日，共十四日。
1KGS|8|66|第八日，王遣散百姓；他们都为王祝福。他们为耶和华向他仆人 大卫 和他百姓 以色列 所施的一切恩惠都心中喜乐，愉快地各回自己的帐棚去了。
1KGS|9|1|所罗门 建造耶和华的殿和王宫，以及一切所想要建造的都完毕了，
1KGS|9|2|耶和华第二次向 所罗门 显现，如先前在 基遍 向他显现一样。
1KGS|9|3|耶和华对他说：“我已听了你在我面前的祷告和祈求，将你所建的这殿分别为圣，使我的名永远立在那里；我的眼、我的心也必时常在那里。
1KGS|9|4|你若以纯正的心和正直行在我面前，效法你父 大卫 所行的，遵行我一切所吩咐你的，谨守我的律例典章，
1KGS|9|5|我就必坚固你在 以色列 国度的王位，直到永远，正如我应许你父 大卫 说：‘你的子孙必不断有人坐 以色列 的王位。’
1KGS|9|6|倘若你们和你们的子孙转去不跟从我，不守我摆在你们面前的诫命律例，去事奉别神，敬拜它们，
1KGS|9|7|我就必把 以色列 从我赐给他们的地上剪除，也必从我面前舍弃那为我名所分别为圣的殿，使 以色列 在万民中成为笑柄，被人讥诮。
1KGS|9|8|这殿虽然崇高 ，将来凡经过的人必惊讶，嗤笑，说：‘耶和华为何向这地和这殿如此行呢？’
1KGS|9|9|人必说：‘因为此地的人离弃领他们祖先出 埃及 地的耶和华－他们的上帝，去亲近别神，敬拜事奉它们，所以耶和华使这一切灾祸临到他们。’”
1KGS|9|10|所罗门 建造耶和华殿和王宫这两座殿宇，用了二十年才完成。
1KGS|9|11|推罗 王 希兰 曾照 所罗门 所要的资助他香柏木、松木和金子， 所罗门 王就把 加利利 地的二十座城给了 希兰 。
1KGS|9|12|希兰 从 推罗 出来，察看 所罗门 给他的城镇，看不顺眼，
1KGS|9|13|就说：“我兄啊，你给我的是什么城镇呢？”他就给这些城镇起名叫 迦步勒 地，直到今日。
1KGS|9|14|希兰 曾给 所罗门 一百二十他连得金子。
1KGS|9|15|所罗门 王挑取服劳役的工人，为要建造耶和华的殿、自己的宫、 米罗 、 耶路撒冷 的城墙、 夏琐 、 米吉多 和 基色 。
1KGS|9|16|先前 埃及 王法老上来攻取 基色 ，用火焚烧，杀了城内居住的 迦南 人，把城赐给他的女儿，就是 所罗门 的妻子，作为嫁妆。
1KGS|9|17|所罗门 建造 基色 、 下伯．和仑 、
1KGS|9|18|巴拉 ，和位于境内旷野的 达莫 。
1KGS|9|19|所罗门 建造一切的储货城、战车城、战马城，以及他所想要建造的，在 耶路撒冷 、 黎巴嫩 和自己治理全国中的一切建设。
1KGS|9|20|至于所有剩下的百姓，不属 以色列 人的 亚摩利 人、 赫 人、 比利洗 人、 希未 人、 耶布斯 人，
1KGS|9|21|那些 以色列 人在当地不能灭尽的人， 所罗门 征召他们剩下的后代作服劳役的奴仆，直到今日。
1KGS|9|22|惟有 以色列 人， 所罗门 不使他们作奴仆，而是作他的战士、臣仆、官长、军官、战车长、骑兵长。
1KGS|9|23|这些是 所罗门 工程的五百五十个监工，他们在百姓中监管作工的人。
1KGS|9|24|法老的女儿从 大卫城 上到 所罗门 为她建造的宫里。那时， 所罗门 才建造 米罗 。
1KGS|9|25|所罗门 每年三次在他为耶和华所筑的坛上献燔祭和平安祭，又在耶和华面前的坛上烧香。这样，他完成了建殿。
1KGS|9|26|所罗门 王在 以东 地 红海 边，靠近 以禄 的 以旬．迦别 制造船只。
1KGS|9|27|希兰 派他的仆人，就是熟悉航海的船员，与 所罗门 的仆人一同坐船航海。
1KGS|9|28|他们到了 俄斐 ，从那里得了四百二十他连得金子，运到 所罗门 王那里。
1KGS|10|1|示巴 女王听见 所罗门 因耶和华的名所得的名声，就来要用难题考问 所罗门 。
1KGS|10|2|她带着很多的随从来到 耶路撒冷 ，有骆驼驮着香料、极多金子和宝石。她来到 所罗门 那里，向他提出心中所有的问题。
1KGS|10|3|所罗门 回答了她所有的问题，没有一个问题太难，王不能向她解答的。
1KGS|10|4|示巴 女王看见 所罗门 一切的智慧，和他所建造的宫殿，
1KGS|10|5|席上的食物，坐着的群臣，侍立的仆人，他们的服装，和他的司酒长，以及他在耶和华殿里所献的燔祭 ，就诧异得神不守舍。
1KGS|10|6|她对王说：“我在本国所听到的话，论到你的事和你的智慧是真的！
1KGS|10|7|我本来不信那些话，及至我来亲眼看见了，看哪，人所告诉我的还不到一半，你的智慧和你的福分超过我所听见的传闻。
1KGS|10|8|你的人 是有福的！你这些仆人常侍立在你面前、听你智慧的话是有福的！
1KGS|10|9|耶和华－你的上帝是应当称颂的！他喜爱你，使你坐 以色列 的王位，因为他永远爱 以色列 ，所以立你作王，使你秉公行义。”
1KGS|10|10|于是， 示巴 女王把一百二十他连得金子、极多的香料和宝石送给 所罗门 王；送来的香料，从来没有像 示巴 女王送给他的那么多。
1KGS|10|11|希兰 的船只也从 俄斐 运了金子来，又从 俄斐 运了许多檀香木和宝石来。
1KGS|10|12|王用檀香木为耶和华的殿和王宫做栏杆，又为歌唱的人做琴瑟。以后再没有这样的檀香木运进来，也再没有人见过，直到如今。
1KGS|10|13|所罗门 王除了照自己的厚意馈赠 示巴 女王之外，凡她所提出的一切要求， 所罗门 王都送给她。于是女王和她臣仆转回，到本国去了。
1KGS|10|14|所罗门 每年所得的金子，重六百六十六他连得；
1KGS|10|15|另外还有来自商人 和做生意的商品，以及 阿拉伯 诸王和各地省长的。
1KGS|10|16|所罗门 王用锤出来的金子打成二百面盾牌，每面盾牌用六百舍客勒金子；
1KGS|10|17|又用锤出来的金子打成三百面小盾牌，每面小盾牌用三弥那金子。王把它们放在 黎巴嫩林宫 里。
1KGS|10|18|王又制造一个大的象牙宝座，包上纯金。
1KGS|10|19|宝座有六层台阶，座的后背是圆的，座位之处两旁有扶手，靠近扶手有两只狮子站立。
1KGS|10|20|六层台阶上有十二只狮子站立，分站左边和右边；任何国度都没有这样做的。
1KGS|10|21|所罗门 王一切的饮器都是金的， 黎巴嫩林宫 里所有的器皿都是纯金的。在 所罗门 的日子，银子算不了什么。
1KGS|10|22|王有 他施 船只与 希兰 的船只一同航海， 他施 船只每三年一次把金、银、象牙、猿猴、孔雀 运回来。
1KGS|10|23|所罗门 王的财宝与智慧胜过地上的众王。
1KGS|10|24|全地都求见 所罗门 的面，要听上帝放在他心里的智慧。
1KGS|10|25|他们各带贡物，就是银器、金器、衣服、兵器、香料、马、骡子，每年都有一定的数量。
1KGS|10|26|所罗门 聚集战车骑兵；他有一千四百辆战车，一万二千名骑兵，安置在屯车城，在 耶路撒冷 的王那里。
1KGS|10|27|王在 耶路撒冷 使银子多如石头，香柏木多如 谢非拉 的桑树。
1KGS|10|28|所罗门 的马是从 埃及 和 科威 运来的，是王的商人按着定价从 科威 买来的。
1KGS|10|29|从 埃及 进口的战车，每辆六百舍客勒银子，马每匹一百五十舍客勒； 赫 人众王和 亚兰 诸王的战车和马，也是经由他们的手出口的。
1KGS|11|1|所罗门 王在法老的女儿之外，又宠爱许多外邦女子，就是 摩押 女子、 亚扪 女子、 以东 女子、 西顿 女子、 赫 人女子。
1KGS|11|2|论到这些国的人，耶和华曾吩咐 以色列 人说：“你们不可跟他们通婚，他们也不可跟你们在一起，因为他们一定会诱惑你们的心去随从他们的神明。” 所罗门 却为了爱，紧紧跟从他们。
1KGS|11|3|所罗门 娶七百个公主，三百个妃嫔。这些妻妾诱惑他的心。
1KGS|11|4|所罗门 年老的时候，他的妻妾诱惑他的心去随从别神，不像他父亲 大卫 以纯正的心顺服耶和华－他的上帝。
1KGS|11|5|所罗门 随从 西顿 人的女神 亚斯她录 和 亚扪 人可憎的 米勒公 。
1KGS|11|6|所罗门 行耶和华眼中看为恶的事，不像他父亲 大卫 专心顺从耶和华。
1KGS|11|7|那时， 所罗门 为 摩押 可憎的 基抹 和 亚扪 人可憎的 摩洛 ，在 耶路撒冷 对面的山上建造丘坛。
1KGS|11|8|他为所有的妻妾，就是那些向自己神明烧香献祭的外邦女子，也是这样做。
1KGS|11|9|耶和华向 所罗门 发怒，因为他的心偏离了向他显现两次的耶和华－ 以色列 的上帝。
1KGS|11|10|耶和华曾吩咐他这件事，不可随从别神，他却没有遵守耶和华所吩咐的。
1KGS|11|11|所以耶和华对他说：“你既然是这样，不遵守我所吩咐你守的约和律例，我必定把国度撕裂离开你，将它赐给你的大臣。
1KGS|11|12|然而，因你父亲 大卫 的缘故，我不在你的日子行这事，而要从你儿子的手中撕裂这国。
1KGS|11|13|只是我不撕裂全国，却要因我仆人 大卫 和我所选择的 耶路撒冷 ，保留一个支派给你的儿子。”
1KGS|11|14|耶和华使 以东 人 哈达 兴起，作 所罗门 的敌人；他是 以东 王的后裔。
1KGS|11|15|大卫 在 以东 的时候， 约押 元帅上去埋葬阵亡的人，杀了 以东 所有的男丁。
1KGS|11|16|约押 和 以色列 众人在 以东 住了六个月，直到把 以东 的男丁尽都剪除。
1KGS|11|17|那时 哈达 还是幼童；他和他父亲的臣仆，以及几个 以东 人逃往 埃及 。
1KGS|11|18|他们从 米甸 起行，到了 巴兰 ，再从 巴兰 带着几个人来到 埃及 ，到 埃及 王法老那里。法老给他房屋，吩咐给他粮食，又把地赐给他。
1KGS|11|19|哈达 在法老眼前大蒙恩宠，法老就把王后 答比匿 的妹妹嫁给他。
1KGS|11|20|答比匿 的妹妹给 哈达 生了一个儿子，叫 基努拔 。 答比匿 使 基努拔 在法老的宫里断奶， 基努拔 就与法老的众子一同住在法老的宫里。
1KGS|11|21|哈达 在 埃及 听见 大卫 与他祖先同睡， 约押 元帅也死了，就对法老说：“请你让我走，我要回本国去。”
1KGS|11|22|法老对他说：“你在我这里有什么缺乏？看哪，你竟想要回你本国去！”他说：“我没有缺乏什么，只是恳求王准我回去。”
1KGS|11|23|上帝又使 以利亚大 的儿子 利逊 兴起，作 所罗门 的敌人。他曾逃避主人 琐巴 王 哈大底谢 。
1KGS|11|24|大卫 击杀 琐巴 人的时候， 利逊 召集了一群人，自己作他们的领袖。他们往 大马士革 ，住在那里，在 大马士革 建立王国。
1KGS|11|25|所罗门 活着的时候，除了 哈达 为患之外， 利逊 也作 以色列 的敌人。他憎恨 以色列 ，作了 亚兰 人的王。
1KGS|11|26|尼八 的儿子 耶罗波安 也举起手来攻击王。他是 所罗门 的臣仆， 以法莲 支派的 洗利达 人；他母亲是个寡妇，名叫 洗鲁阿 。
1KGS|11|27|他举手攻击王是因先前 所罗门 建造 米罗 ，修补他父亲 大卫城 缺口的这件事。
1KGS|11|28|耶罗波安 是个大有才能的人。 所罗门 见这青年殷勤，就派他监管 约瑟 家所有服劳役的工人。
1KGS|11|29|那时， 耶罗波安 出了 耶路撒冷 ， 示罗 人 亚希雅 先知在路上遇见他； 亚希雅 身上穿着一件新衣。田野中只有他们二人，没有其他的人。
1KGS|11|30|亚希雅 拿起穿在自己身上的新衣，把它撕成十二片，
1KGS|11|31|对 耶罗波安 说：“你可以拿十片。耶和华－ 以色列 的上帝如此说：‘看哪，我必从 所罗门 手里撕裂这国，把十个支派赐给你。
1KGS|11|32|我因我仆人 大卫 和我在 以色列 众支派中所选择的 耶路撒冷城 的缘故，仍为 所罗门 留一个支派。
1KGS|11|33|因为他们 离弃我，敬拜 西顿 人的女神 亚斯她录 、 摩押 的神明 基抹 和 亚扪 人的神明 米勒公 ，没有像他父亲 大卫 一样遵从我的道，行我眼中看为正的事，守我的律例典章。
1KGS|11|34|但我不从他手里夺走整个国家，却使他在活着的日子作君王，是因我所拣选的仆人 大卫 遵守我的诫命律例。
1KGS|11|35|我必从他儿子手里将王国夺走，赐给你十个支派，
1KGS|11|36|只留一个支派给他的儿子，使我仆人 大卫 在我所选择立我名的 耶路撒冷城 那里，在我面前常有灯光。
1KGS|11|37|我选你，使你照你心里一切所愿的作王，成为 以色列 的王。
1KGS|11|38|你若听从我一切所吩咐你的，遵行我的道，行我眼中看为正的事，谨守我的律例诫命，像我仆人 大卫 所行的，我就与你同在，为你立坚固的家，像我为 大卫 所立的一样，将 以色列 赐给你。
1KGS|11|39|我必因这事使 大卫 的后裔遭受患难，但不是永远的。’”
1KGS|11|40|所罗门 想要杀 耶罗波安 ， 耶罗波安 起身逃往 埃及 。他到了 埃及 王 示撒 那里，就住在 埃及 ，直到 所罗门 死了。
1KGS|11|41|所罗门 其余的事，凡他所做的和他的智慧，不都写在《所罗门记》上吗？
1KGS|11|42|所罗门 在 耶路撒冷 作全 以色列 的王四十年。
1KGS|11|43|所罗门 与他祖先同睡，葬在他父亲 大卫 的城里，他儿子 罗波安 接续他作王。
1KGS|12|1|罗波安 往 示剑 去，因 以色列 众人都到了 示剑 ，要立他作王。
1KGS|12|2|尼八 的儿子 耶罗波安 先前躲避 所罗门 王，逃往 埃及 ，住在那里。他还在 埃及 ，听见了这事 ，
1KGS|12|3|以色列 人派人去请他来。 耶罗波安 就和 以色列 全会众来，与 罗波安 谈话，说：
1KGS|12|4|“你父亲使我们负重轭，现在求你减轻你父亲所加给我们的苦工和重轭，我们就服事你。”
1KGS|12|5|罗波安 对他们说：“你们走吧，过三天再来见我。”百姓就走了。
1KGS|12|6|罗波安 的父亲 所罗门 在世的日子，有侍立在他面前的长者， 罗波安 王和他们商议，说：“你们出个主意，好把话带回给这百姓。”
1KGS|12|7|他们对他说：“现在王若像仆人一样服事这百姓，用好话回覆他们，他们就永远作王的仆人了。”
1KGS|12|8|王不采纳长者给他出的主意，却和那些与他一同长大、在他面前侍立的年轻人商议。
1KGS|12|9|他对他们说：“这百姓对我说：‘你父亲使我们负重轭，求你减轻一些。’你们出个什么主意，我们好把话带回给他们。”
1KGS|12|10|那些与他一同长大的年轻人对他说：“这百姓对王说：‘你父亲使我们负重轭，求你给我们减轻一些。’王要对他们如此说：‘我的小指头比我父亲的腰还粗呢！
1KGS|12|11|我父亲使你们负重轭，现在我必使你们负更重的轭！我父亲用鞭子惩罚你们，我要用蝎子惩罚你们！’”
1KGS|12|12|耶罗波安 和众百姓遵照王所说“你们第三天再来见我”的话，第三天来到 罗波安 那里。
1KGS|12|13|王严厉地回答百姓，不采纳长者给他出的主意。
1KGS|12|14|他照着年轻人所出的主意对他们说：“我父亲使你们负重轭，我必使你们负更重的轭！我父亲用鞭子惩罚你们，我却要用蝎子惩罚你们！”
1KGS|12|15|王不依从百姓，因这事件是出于耶和华，为要应验耶和华藉 示罗 人 亚希雅 对 尼八 的儿子 耶罗波安 所说的话。
1KGS|12|16|以色列 众人见王不依从他们，百姓就回话给王，说： “我们在 大卫 中有什么份呢？ 我们在 耶西 的儿子中没有产业！ 以色列 啊，回你的帐棚去吧！ 大卫 啊，现在你顾自己的家吧！” 于是， 以色列 人都回自己的帐棚去了；
1KGS|12|17|至于住 犹大 城镇的 以色列 人， 罗波安 仍作他们的王。
1KGS|12|18|罗波安 王派监管劳役的 亚多兰 去， 以色列 众人用石头打他，他就死了。 罗波安 王急忙上车，逃回 耶路撒冷 去了。
1KGS|12|19|这样， 以色列 背叛 大卫 家，直到今日。
1KGS|12|20|以色列 众人听见 耶罗波安 回来了，就派人去请他到会众那里，立他作全 以色列 的王。除了 犹大 支派，没有跟从 大卫 家的。
1KGS|12|21|罗波安 来到 耶路撒冷 ，召集了 犹大 全家和 便雅悯 支派的人共十八万，都是精选的战士，要与 以色列 家打仗，好将王国夺回，归 所罗门 的儿子 罗波安 。
1KGS|12|22|但上帝的话临到神人 示玛雅 ，说：
1KGS|12|23|“你去告诉 所罗门 的儿子 犹大 王 罗波安 ， 犹大 和 便雅悯 全家，以及其余的百姓，说：
1KGS|12|24|‘耶和华如此说：你们不可上去与你们的弟兄 以色列 人打仗。你们各自回家去吧！因为这事是出于我。’”众人就听从耶和华的话，遵照耶和华的话回去了。
1KGS|12|25|耶罗波安 在 以法莲 山区建了 示剑 ，住在其中，又从 示剑 出去，建了 毗努伊勒 。
1KGS|12|26|耶罗波安 心里说：“现在，这国恐怕仍会归 大卫 家；
1KGS|12|27|这百姓若上 耶路撒冷 去，在耶和华的殿里献祭，他们的心必归向他们的主 犹大 王 罗波安 。他们会杀了我，仍归 犹大 王 罗波安 。”
1KGS|12|28|耶罗波安 王就筹划，铸造了两个金牛犊，对众百姓说：“你们上 耶路撒冷 去实在够久了。 以色列 啊，看哪，这是领你出 埃及 地的神明。”
1KGS|12|29|他把一个安置在 伯特利 ，另一个安置在 但 。
1KGS|12|30|这事使百姓陷入罪里，因为他们甚至到 但 去拜那牛犊。
1KGS|12|31|耶罗波安 在一些丘坛建神殿，立不属 利未 人的平民百姓为祭司。
1KGS|12|32|耶罗波安 定八月十五日为节期，像在 犹大 的节期一样，自己上坛献祭。他在 伯特利 这样做，向他所铸的牛犊献祭，又把他所立丘坛的祭司安置在 伯特利 。
1KGS|12|33|他在八月十五日，就是他自己心中所定的月份，在 伯特利 上到自己所造的祭坛；他为 以色列 人定了一个节期，亲自上坛烧香。
1KGS|13|1|看哪，有一个神人遵照耶和华的话从 犹大 来到 伯特利 。 耶罗波安 正站在坛旁烧香；
1KGS|13|2|神人遵照耶和华的话向坛呼叫，说：“坛哪，坛哪！耶和华如此说：‘看哪， 大卫 家必生一个儿子，名叫 约西亚 ，他必将在你上面烧香的丘坛祭司，宰杀在你上面，人的骨头也必烧在你上面。’”
1KGS|13|3|当日，神人设个预兆，说：“这是耶和华说的预兆：‘看哪，这坛必破裂，坛上的灰必倾倒出来。’”
1KGS|13|4|耶罗波安 王听见神人向 伯特利 的坛呼叫的话，就从坛上伸手，说：“拿住他！”王向神人所伸的手却萎缩了，不能弯回。
1KGS|13|5|坛也破裂了，坛上的灰倾倒出来，正如神人遵照耶和华的话所设的预兆。
1KGS|13|6|王对神人说：“请你为我祷告，向耶和华－你的上帝恳求恩惠，使我的手复原。”于是神人向耶和华恳求，王的手就复原了，如平常一样。
1KGS|13|7|王对神人说：“请你跟我回宫，让你恢复心力，我必给你赏赐。”
1KGS|13|8|神人对王说：“你就是把你一半的王宫给我，我也不跟你进去，也不在这地方吃饭喝水，
1KGS|13|9|因为耶和华的话这样吩咐我说：‘不可吃饭喝水，也不可从你去的原路回来。’”
1KGS|13|10|于是神人从别的路回去，不从他到 伯特利 来的原路回去。
1KGS|13|11|有一个老先知住在 伯特利 ，他的儿子来，把神人当日在 伯特利 所做的一切事和他向王所说的话，都告诉了父亲。
1KGS|13|12|父亲对他们说：“神人从哪条路去了呢？”他的儿子都看到 从 犹大 来的神人所去的路。
1KGS|13|13|老先知吩咐儿子说：“你们为我备驴。”他们备好了驴，他就骑上，
1KGS|13|14|去追神人，遇见神人坐在橡树底下，就对他说：“你是不是从 犹大 来的神人？”他说：“是我。”
1KGS|13|15|老先知对他说：“请你跟我一起回家吃饭。”
1KGS|13|16|神人说：“我不能跟你回去，与你同行，也不能在这地方跟你一起吃饭喝水，
1KGS|13|17|因为有耶和华的话吩咐我说：‘你在那里不可吃饭喝水，也不可从你去的原路回来。’”
1KGS|13|18|老先知对他说：“我也是先知，和你一样。有天使遵照耶和华的话对我说：‘你去带他一同回你的家，给他吃饭喝水。’”老先知在欺骗他。
1KGS|13|19|于是神人跟老先知回去，在他家里吃饭喝水。
1KGS|13|20|他们坐席的时候，耶和华的话临到那带神人回来的先知，
1KGS|13|21|他就对从 犹大 来的神人宣告说：“耶和华如此说：‘你既违背耶和华的指示，不遵守耶和华－你上帝的命令，
1KGS|13|22|反倒回来，在耶和华禁止你吃饭喝水的地方吃了饭喝了水，因此你的尸体必不得葬在你祖先的坟墓里。’”
1KGS|13|23|神人吃喝完了，老先知为他带回来的先知备驴。
1KGS|13|24|神人就去了，在路上有只狮子遇见他，把他咬死。他的尸体倒在路上，驴站在尸体旁边，狮子也站在尸体旁边。
1KGS|13|25|看哪，有人经过，看见尸体倒在路上，狮子站在尸体旁边，就来到老先知所住的城里述说这事。
1KGS|13|26|那带神人回来的先知听见了，就说：“这是那违背了耶和华指示的神人，所以耶和华把他交给狮子；狮子撕裂他，咬死他，正如耶和华对他说的话。”
1KGS|13|27|老先知吩咐他儿子说：“你们为我备驴。”他们就备了驴。
1KGS|13|28|他去了，发现神人的尸体倒在路上，驴和狮子站在尸体旁边，狮子却没有吃尸体，也没有撕裂驴。
1KGS|13|29|老先知把神人的尸体抬起，驮在驴上，带回自己的城里，要为他哀哭，为他安葬。
1KGS|13|30|老先知把尸体葬在自己的坟里，为他哀哭，说：“哀哉！我的弟兄啊！”
1KGS|13|31|安葬之后，老先知对他儿子说：“我死了，你们要把我葬在神人所葬的坟里，使我的尸骨在他的尸骨旁边，
1KGS|13|32|因为他遵照耶和华的话，指着 伯特利 的坛和 撒玛利亚 各城丘坛神殿所宣告的话必定应验。”
1KGS|13|33|这事以后， 耶罗波安 仍不离开他的恶道，立平民百姓为丘坛的祭司；凡愿意的，他都分别为圣，立为丘坛的祭司。
1KGS|13|34|这事使 耶罗波安 的家陷入罪里，甚至他的家被剪除，从地面上消灭了。
1KGS|14|1|那时， 耶罗波安 的儿子 亚比雅 病了。
1KGS|14|2|耶罗波安 对他的妻子说：“你起来改装，使人认不出你是 耶罗波安 的妻子。你往 示罗 去，看哪，那里有先知 亚希雅 ，他曾告诉我说，你必作这百姓的王。
1KGS|14|3|现在你手里要带十个饼、几个薄饼和一瓶蜜到他那里去，他必告诉你，孩子会怎样。”
1KGS|14|4|耶罗波安 的妻子就照样做，起身往 示罗 去，到了 亚希雅 的家。 亚希雅 因年纪老迈，两眼发直，不能看见。
1KGS|14|5|耶和华对 亚希雅 说：“看哪， 耶罗波安 的妻子来问你她儿子的事，因她儿子病了，你当如此如此告诉她。她进来的时候会扮成别的妇人。”
1KGS|14|6|她刚进门， 亚希雅 听见她的脚步声，就说：“ 耶罗波安 的妻子，进来吧！你为何扮成别的妇人呢？我奉差遣将凶信告诉你。
1KGS|14|7|你回去告诉 耶罗波安 说：‘耶和华－ 以色列 的上帝如此说：我从百姓中提拔了你，立你作我百姓 以色列 的君王，
1KGS|14|8|将 大卫 家的国撕裂，赐给你，你却不效法我仆人 大卫 ，遵守我的诫命，全心顺从我，行我眼中看为正的事。
1KGS|14|9|你反倒行恶，比在你之前所有的人更严重；你离开了我，为自己立了别神，铸了偶像，惹我发怒，将我丢在背后。
1KGS|14|10|因此，看哪，我必使灾祸临到 耶罗波安 的家，把属 耶罗波安 的男丁，无论是奴役的、自由的，都从 以色列 中剪除。我必除灭 耶罗波安 的家，如同人扫除粪土，直到消灭。
1KGS|14|11|凡属 耶罗波安 的人，死在城中的必被狗吃，死在田野的必被空中的鸟吃。这是耶和华说的。’
1KGS|14|12|你起身回家去吧！你的脚一进城，孩子就死了。
1KGS|14|13|以色列 众人必为他哀哭，为他安葬。凡属 耶罗波安 的人，只有他可以葬入坟墓，因为在 耶罗波安 的家中，只有他向耶和华－ 以色列 的上帝表现出好的行为。
1KGS|14|14|耶和华必另立一王治理 以色列 ，这一天，他必剪除 耶罗波安 的家；什么时候呢？现在就是了。
1KGS|14|15|耶和华必击打 以色列 ，使他们摇动，像水中的芦苇一样，又将他们从耶和华赐给他们列祖的美地上拔出来，分散在 大河 那边，因为他们造了 亚舍拉 ，惹耶和华发怒。
1KGS|14|16|因 耶罗波安 所犯的罪，又因他使 以色列 陷入罪里，耶和华必将 以色列 交出来。”
1KGS|14|17|耶罗波安 的妻子起身回去，到了 得撒 ，刚到门槛，孩子就死了。
1KGS|14|18|以色列 众人为他安葬，为他哀哭，正如耶和华藉他仆人 亚希雅 先知所说的话。
1KGS|14|19|耶罗波安 其余的事，他怎样打仗，怎样作王，看哪，都写在《以色列诸王记》上。
1KGS|14|20|耶罗波安 作王二十二年，就与他祖先同睡，他儿子 拿答 接续他作王。
1KGS|14|21|所罗门 的儿子 罗波安 作 犹大 王。他登基的时候年四十一岁，在 耶路撒冷 ，就是耶和华从 以色列 众支派中所选择立他名的城，作王十七年。 罗波安 的母亲名叫 拿玛 ，是 亚扪 人。
1KGS|14|22|犹大 人行耶和华眼中看为恶的事，以所犯的罪惹动他的妒忌，比他们的祖先所犯的一切更严重。
1KGS|14|23|因为他们在各高冈上，各青翠树下筑丘坛，立柱像和 亚舍拉 。
1KGS|14|24|国中也有男的庙妓。他们效法耶和华在 以色列 人面前所赶出的外邦人，行一切可憎恶的事。
1KGS|14|25|罗波安 王第五年， 埃及 王 示撒 上来攻打 耶路撒冷 ，
1KGS|14|26|夺了耶和华殿和王宫里的宝物，尽都带走，又夺走 所罗门 制造的一切金盾牌。
1KGS|14|27|罗波安 王制造铜盾牌代替那些金盾牌，交给看守王宫宫门的护卫长看管。
1KGS|14|28|每逢王进耶和华的殿，护卫兵就举起这些盾牌；随后仍将盾牌送回护卫室。
1KGS|14|29|罗波安 其余的事，凡他所做的，不都写在《犹大列王记》上吗？
1KGS|14|30|罗波安 与 耶罗波安 时常交战。
1KGS|14|31|罗波安 与他祖先同睡，与他祖先同葬在 大卫城 。他母亲名叫 拿玛 ，是 亚扪 人，他儿子 亚比央 接续他作王。
1KGS|15|1|尼八 的儿子 耶罗波安 王十八年， 亚比央 登基作 犹大 王，
1KGS|15|2|在 耶路撒冷 作王三年。他母亲名叫 玛迦 ，是 押沙龙 的女儿。
1KGS|15|3|亚比央 行他父亲从前所犯一切的罪，他的心不像他曾祖父 大卫 以纯正的心顺服耶和华－他的上帝。
1KGS|15|4|然而耶和华－他的上帝因 大卫 的缘故，仍使大卫在 耶路撒冷 有灯光，立他儿子接续他作王，又坚立 耶路撒冷 。
1KGS|15|5|因为 大卫 除了 赫 人 乌利亚 那件事，都行耶和华眼中看为正的事，一生没有违背耶和华一切所吩咐的。
1KGS|15|6|罗波安 在世的日子常与 耶罗波安 交战。
1KGS|15|7|亚比央 其余的事，凡他所做的，不都写在《犹大列王记》上吗？ 亚比央 常与 耶罗波安 交战。
1KGS|15|8|亚比央 与他祖先同睡，葬在 大卫城 ，他儿子 亚撒 接续他作王。
1KGS|15|9|以色列 王 耶罗波安 第二十年， 亚撒 登基作 犹大 王，
1KGS|15|10|在 耶路撒冷 作王四十一年。他祖母名叫 玛迦 ，是 押沙龙 的女儿。
1KGS|15|11|亚撒 效法他的高祖父 大卫 行耶和华眼中看为正的事，
1KGS|15|12|从国中除去男的庙妓，又除掉他祖先所造的一切偶像。
1KGS|15|13|他甚至废了他祖母 玛迦 太后的位，因 玛迦 造了可憎的 亚舍拉 。 亚撒 砍下她的偶像，在 汲沦溪 边烧了，
1KGS|15|14|只是丘坛还没有废去。 亚撒 一生向耶和华存纯正的心。
1KGS|15|15|亚撒 将他父亲所分别为圣与自己所分别为圣的金银和器皿都奉到耶和华的殿里。
1KGS|15|16|亚撒 和 以色列 王 巴沙 在世的日子常常交战。
1KGS|15|17|以色列 王 巴沙 上来攻击 犹大 ，修筑 拉玛 ，不许人从 犹大 王 亚撒 那里出入。
1KGS|15|18|于是 亚撒 把耶和华殿和王宫府库里所剩下的金银都交在他臣仆手中，派他们到住在 大马士革 的 亚兰 王，就是 希旬 的孙子， 他伯利门 的儿子 便．哈达 那里去，说：
1KGS|15|19|“你父曾与我父立约，我与你也要这样立约。看哪，我把金银送给你作礼物，请你废掉你与 以色列 王 巴沙 所立的约，使他从我这里撤退。”
1KGS|15|20|便．哈达 听从了 亚撒 王，就派遣他的军官去攻打 以色列 的城镇，攻下了 以云 、 但 、 亚伯．伯．玛迦 、全 基尼烈 、 拿弗他利 全地。
1KGS|15|21|巴沙 听见了，就停工不修筑 拉玛 ，仍住在 得撒 。
1KGS|15|22|于是 亚撒 王向 犹大 众人宣布，不准任何人推辞，吩咐他们运走 巴沙 修筑 拉玛 所用的石头和木料。 亚撒 王用它们来修筑 便雅悯 的 迦巴 和 米斯巴 。
1KGS|15|23|亚撒 其余的事，他英勇的事迹，凡他所做的，以及他所建筑的城镇，不都写在《犹大列王记》上吗？只是 亚撒 年老的时候患有脚疾。
1KGS|15|24|亚撒 与他祖先同睡，与他祖先同葬在 大卫城 ，他儿子 约沙法 接续他作王。
1KGS|15|25|犹大 王 亚撒 第二年， 耶罗波安 的儿子 拿答 登基作 以色列 王二年，
1KGS|15|26|拿答 行耶和华眼中看为恶的事，行他父亲所行的道，犯他父亲使 以色列 陷入罪里的那罪。
1KGS|15|27|以萨迦 人 亚希雅 的儿子 巴沙 背叛 拿答 ，在 非利士 人的 基比顿 杀了他，那时 拿答 和 以色列 众人正围困 基比顿 。
1KGS|15|28|犹大 王 亚撒 第三年， 巴沙 杀了 拿答 ，篡了他的位。
1KGS|15|29|巴沙 一作王就杀了 耶罗波安 全家， 耶罗波安 家凡有气息的，一个也没有留下，都杀灭了，正如耶和华藉他仆人 示罗 人 亚希雅 所说的话。
1KGS|15|30|这是因为 耶罗波安 所犯的罪，他使 以色列 陷入罪里，激怒了耶和华－ 以色列 的上帝。
1KGS|15|31|拿答 其余的事，凡他所做的，不都写在《以色列诸王记》上吗？
1KGS|15|32|亚撒 和 以色列 王 巴沙 在世的日子常常交战。
1KGS|15|33|犹大 王 亚撒 第三年， 亚希雅 的儿子 巴沙 在 得撒 登基，作全 以色列 的王二十四年。
1KGS|15|34|他行耶和华眼中看为恶的事，行 耶罗波安 所行的道，犯他使 以色列 陷入罪里的那罪。
1KGS|16|1|耶和华的话临到 哈拿尼 的儿子 耶户 ，责备 巴沙 说：
1KGS|16|2|“我既从尘埃中提拔你，立你作我百姓 以色列 的君王，你竟行 耶罗波安 所行的道，使我的百姓 以色列 陷入罪里，以他们的罪惹我发怒，
1KGS|16|3|看哪，我必除尽 巴沙 和他的家，使你的家像 尼八 的儿子 耶罗波安 的家一样。
1KGS|16|4|凡属 巴沙 的人，死在城中的必被狗吃，死在田野的必被空中的鸟吃。”
1KGS|16|5|巴沙 其余的事，凡他所做的和他英勇的事迹，不都写在《以色列诸王记》上吗？
1KGS|16|6|巴沙 与他祖先同睡，葬在 得撒 ，他儿子 以拉 接续他作王。
1KGS|16|7|耶和华的话临到 哈拿尼 的儿子 耶户 先知，责备 巴沙 和他的家，因他行耶和华眼中看为恶的一切事，以他手所做的惹耶和华发怒，像 耶罗波安 的家一样，又因他杀了 耶罗波安 全家。
1KGS|16|8|犹大 王 亚撒 第二十六年， 巴沙 的儿子 以拉 在 得撒 登基，作 以色列 王二年。
1KGS|16|9|他的大臣 心利 ，就是管理他一半战车的军官背叛他。当他在 得撒 ，在王宫的管家 亚杂 家里喝醉的时候，
1KGS|16|10|心利 进去击杀他，把他杀死，篡了他的位。这是 犹大 王 亚撒 第二十七年的事。
1KGS|16|11|心利 一坐上王位就杀了 巴沙 全家，连他的亲属和朋友，一个男丁也没有留下。
1KGS|16|12|心利 灭绝 巴沙 全家，正如耶和华藉 耶户 先知责备 巴沙 的话。
1KGS|16|13|这是因为 巴沙 和他儿子 以拉 的一切罪，就是他们使 以色列 陷入罪里的那罪，以虚无的神明 惹耶和华－ 以色列 的上帝发怒。
1KGS|16|14|以拉 其余的事，凡他所做的，不都写在《以色列诸王记》上吗？
1KGS|16|15|犹大 王 亚撒 第二十七年， 心利 在 得撒 作王七日。那时军兵正安营围攻 非利士 人的 基比顿 。
1KGS|16|16|军兵在营中听说 心利 已经背叛，杀了王， 以色列 众人当日就在营中立 暗利 元帅作 以色列 王。
1KGS|16|17|暗利 率领 以色列 众人，从 基比顿 上去，围困 得撒 。
1KGS|16|18|心利 见城被攻陷，就进了王宫的堡垒，放火焚烧宫殿，自焚而死。
1KGS|16|19|这是因为他犯罪，行耶和华眼中看为恶的事，行 耶罗波安 所行的道，犯他使 以色列 陷入罪里的那罪。
1KGS|16|20|心利 其余的事和他背叛的事，不都写在《以色列诸王记》上吗？
1KGS|16|21|那时， 以色列 百姓分为两半：一半随从 基纳 的儿子 提比尼 ，要拥立他作王；另一半随从 暗利 。
1KGS|16|22|但随从 暗利 的百姓胜过随从 基纳 儿子 提比尼 的百姓。 提比尼 死了， 暗利 就作了王。
1KGS|16|23|犹大 王 亚撒 第三十一年， 暗利 登基作 以色列 王十二年；他在 得撒 作王六年。
1KGS|16|24|暗利 用二他连得银子向 撒玛 买了 撒玛利亚山 ，在山上建城，按着山的原主 撒玛 的名，给所建的城起名叫 撒玛利亚 。
1KGS|16|25|暗利 行耶和华眼中看为恶的事，比他以前所有的王作恶更严重。
1KGS|16|26|因为他行了 尼八 的儿子 耶罗波安 所行的道，犯他使 以色列 陷入罪里的那罪，以虚无的神明惹耶和华－ 以色列 的上帝发怒。
1KGS|16|27|暗利 其余的事，他所做的和所显出的英勇事迹，不都写在《以色列诸王记》上吗？
1KGS|16|28|暗利 与他祖先同睡，葬在 撒玛利亚 ，他儿子 亚哈 接续他作王。
1KGS|16|29|犹大 王 亚撒 第三十八年， 暗利 的儿子 亚哈 登基作 以色列 王。 暗利 的儿子 亚哈 在 撒玛利亚 作 以色列 王二十二年。
1KGS|16|30|暗利 的儿子 亚哈 行耶和华眼中看为恶的事，比他以前所有的王更严重。
1KGS|16|31|他犯了 尼八 的儿子 耶罗波安 所犯的罪，还当作是小事，又娶了 西顿 王 谒巴力 的女儿 耶洗别 为妻，去事奉 巴力 ，敬拜它，
1KGS|16|32|又在 撒玛利亚 建 巴力庙 ，在庙里为 巴力 筑坛。
1KGS|16|33|亚哈 又造 亚舍拉 ，他所做的惹耶和华－ 以色列 的上帝发怒，比他以前所有的 以色列 王更严重。
1KGS|16|34|亚哈 的日子， 伯特利 人 希伊勒 重修 耶利哥 。立根基的时候，他丧了长子 亚比兰 ；安门的时候，他丧了幼子 西割 ，正如耶和华藉 嫩 的儿子 约书亚 所说的话。
1KGS|17|1|住在 基列 的 提斯比 人 以利亚 对 亚哈 说：“我指着所事奉永生的耶和华－ 以色列 的上帝起誓，这几年我若不祷告，必不降露水，也不下雨。”
1KGS|17|2|耶和华的话临到 以利亚 ，说：
1KGS|17|3|“你离开这里往东去，躲在 约旦河 东边的 基立溪 旁。
1KGS|17|4|你要喝那溪里的水，我已吩咐乌鸦在那里供养你。”
1KGS|17|5|于是 以利亚 去了，他遵照耶和华的话做，去住在 约旦河 东的 基立溪 旁。
1KGS|17|6|乌鸦早上给他叼饼和肉来，晚上也有饼和肉，他又喝溪里的水。
1KGS|17|7|过了些日子溪水干了，因为雨没有下在地上。
1KGS|17|8|耶和华的话临到他，说：
1KGS|17|9|“你起身到 西顿 的 撒勒法 去，住在那里，看哪，我已吩咐那里的一个寡妇供养你。”
1KGS|17|10|以利亚 就起身往 撒勒法 去。他到了城门，看哪，有一个寡妇在那里捡柴。 以利亚 呼唤她说：“请你用器皿取点水来给我喝。”
1KGS|17|11|她去取水的时候， 以利亚 又呼唤她说：“请你手里也拿点饼来给我。”
1KGS|17|12|她说：“我指着永生的耶和华－你的上帝起誓，我没有饼，坛内只有一把面，瓶里只有一点油。看哪，我去找两根柴，带回家为我和我儿子做饼。我们吃了，就等死吧！”
1KGS|17|13|以利亚 对她说：“不要怕！你去照你所说的做吧！只要先为我做一个小饼，拿来给我，然后为你和你的儿子做饼；
1KGS|17|14|因为耶和华－ 以色列 的上帝如此说：‘坛内的面必不用尽，瓶里的油必不短缺，直到耶和华使雨降在地上的日子。’”
1KGS|17|15|妇人就照 以利亚 的话去做。她和 以利亚 ，以及她家中的人，吃了许多日子。
1KGS|17|16|坛内的面果然没有用尽，瓶里的油也不短缺，正如耶和华藉 以利亚 所说的话。
1KGS|17|17|这事以后，那妇人，就是那家的女主人，她的儿子病了，病得很重，甚至没有气息。
1KGS|17|18|妇人对 以利亚 说：“神人哪，我跟你有什么关系，你竟到我这里来，使上帝记起我的罪，以致我的儿子死了呢？”
1KGS|17|19|以利亚 对她说：“把你儿子交给我。” 以利亚 就从妇人怀中接过孩子来，抱到他所住的顶楼，放在自己的床上。
1KGS|17|20|他求告耶和华说：“耶和华－我的上帝啊，我寄居在这寡妇的家里，你却降祸于她，使她的儿子死了吗？”
1KGS|17|21|以利亚 三次伏在孩子的身上，求告耶和华说：“耶和华－我的上帝啊，求你使这孩子的生命归回给他吧！”
1KGS|17|22|耶和华听了 以利亚 的呼求，孩子的生命归回给他，他就活了。
1KGS|17|23|以利亚 把孩子从楼上抱下来，进了房间交给他母亲，说：“看，你的儿子活了！”
1KGS|17|24|妇人对 以利亚 说：“现在我知道你是神人，耶和华藉你口所说的话是真的。”
1KGS|18|1|过了许多日子，到了第三年，耶和华的话临到 以利亚 ，说：“你去，让 亚哈 看见你，我要降雨在地面上。”
1KGS|18|2|以利亚 就去，要让 亚哈 见到他。那时， 撒玛利亚 的饥荒非常严重。
1KGS|18|3|亚哈 召来他的管家 俄巴底 。 俄巴底 非常敬畏耶和华。
1KGS|18|4|耶洗别 杀耶和华先知的时候， 俄巴底 把一百个先知藏了，每五十人藏在一个洞里，拿饼和水供养他们。
1KGS|18|5|亚哈 对 俄巴底 说：“我们要走遍这地，到一切水泉旁和一切溪边，或者能找到青草，可以救活马和骡子，免得丧失一些牲畜。”
1KGS|18|6|于是二人分地巡查， 亚哈 独自走一路， 俄巴底 独自走另一路。
1KGS|18|7|俄巴底 在路上时，看哪， 以利亚 遇见他。 俄巴底 认出他来，就脸伏于地，说：“你是我主 以利亚 吗？”
1KGS|18|8|以利亚 对他说：“我是。你去，告诉你主人说：‘看哪， 以利亚 在这里。’”
1KGS|18|9|俄巴底 说：“仆人犯了什么罪，你竟要把我交在 亚哈 手里，使他杀我呢？
1KGS|18|10|我指着永生的耶和华－你的上帝起誓，无论哪一邦哪一国，我主都派人去找你。若他们说：‘不在这里’，他就叫那邦那国的人起誓说，他们实在找不到你。
1KGS|18|11|现在你说：‘你去告诉你主人说，看哪， 以利亚 在这里’；
1KGS|18|12|恐怕我一离开你，耶和华的灵就把你提到我所不知道的地方去。这样，我去告诉 亚哈 ，他若找不到你，就必杀我。仆人是自幼敬畏耶和华的。
1KGS|18|13|耶洗别 杀耶和华先知的时候，我把耶和华的一百个先知藏了，每五十人藏在一个洞里，拿饼和水供养他们，难道没有人把我做的这事告诉我主吗？
1KGS|18|14|现在你说：‘你去告诉你主人说，看哪， 以利亚 在这里’，他一定会杀我。”
1KGS|18|15|以利亚 说：“我指着所事奉永生的万军之耶和华起誓，我今日要让 亚哈 见到我。”
1KGS|18|16|于是 俄巴底 去迎见 亚哈 ，告诉他这事。 亚哈 就去见 以利亚 。
1KGS|18|17|亚哈 见了 以利亚 ，就说：“真的是你吗？你这使 以色列 遭殃的人！”
1KGS|18|18|以利亚 说：“使 以色列 遭殃的不是我，而是你和你的父家，因为你们离弃耶和华的诫命 ，去随从 巴力 。
1KGS|18|19|现在你要派人去召集 以色列 众人，以及 耶洗别 所供养的四百五十个 巴力 的先知和四百个 亚舍拉 的先知，叫他们都上 迦密山 到我这里来。”
1KGS|18|20|亚哈 就派人到 以色列 众人那里，召集先知上 迦密山 。
1KGS|18|21|以利亚 近前来对众百姓说：“你们心持二意要到几时呢？如果耶和华是上帝，就当顺从耶和华；如果是 巴力 ，就当顺从 巴力 。”百姓一言不答。
1KGS|18|22|以利亚 对百姓说：“作耶和华先知的只剩下我一个； 巴力 的先知却有四百五十人。
1KGS|18|23|请给我们两头牛犊， 巴力 的先知可以为自己挑选一头牛犊，切成小块，放在柴上，不要点火；我也预备一头牛犊放在柴上，也不点火。
1KGS|18|24|你们求告你们神明的名，我也求告耶和华的名。那应允祷告降火的就是上帝。”众百姓回答说：“好主意。”
1KGS|18|25|以利亚 对 巴力 的先知说：“因为你们人多，先挑选一头牛犊，预备好了，求告你们神明的名，却不要点火。”
1KGS|18|26|他们把所给他们的牛犊预备好了，从早晨到中午，求告 巴力 的名说：“ 巴力 啊，求你应允我们！”却没有声音，也没有回应。他们就在所筑的坛四围蹦跳。
1KGS|18|27|到了正午， 以利亚 嘲笑他们，说：“大声求告吧！因为它是神明，它或许在默想，或许正忙着 ，或许在路上，或许在睡觉，它该醒过来了。”
1KGS|18|28|他们大声求告，按着他们的仪式，用刀枪刺割自己，直到浑身流血。
1KGS|18|29|中午过去了，他们狂呼乱叫，直到献晚祭的时候，却没有声音，没有回应的，也没有理睬的。
1KGS|18|30|以利亚 对众百姓说：“你们到我这里来。”众百姓就到他那里，他把那已经毁坏了的耶和华的坛修好。
1KGS|18|31|以利亚 按照 雅各 子孙支派的数目，取了十二块石头；耶和华的话曾临到 雅各 ，说：“你的名要叫 以色列 。”
1KGS|18|32|以利亚 用这些石头为耶和华的名筑一座坛，在坛的四围挖沟，可容纳二细亚谷种。
1KGS|18|33|他又在坛上摆好了柴，把牛犊切成小块放在柴上，说：“你们用四个桶盛满水，倒在燔祭和柴上。”
1KGS|18|34|他又说：“倒第二次。”他们就倒第二次。他又说：“倒第三次。”他们就倒第三次。
1KGS|18|35|水流到坛的四围，沟里也满了水。
1KGS|18|36|到了献晚祭的时候，先知 以利亚 近前来，说：“耶和华－ 亚伯拉罕 、 以撒 、 以色列 的上帝啊，求你今日使人知道你是 以色列 的上帝，我是你的仆人，我遵照你的话做这一切事。
1KGS|18|37|求你应允我，耶和华啊，应允我，使这百姓知道你－耶和华是上帝，是你叫他们回心转意的。”
1KGS|18|38|于是，耶和华降下火来，烧尽燔祭、木柴、石头、尘土，又烧干了沟里的水。
1KGS|18|39|众百姓看见了，就脸伏于地，说：“耶和华是上帝！耶和华是上帝！”
1KGS|18|40|以利亚 对他们说：“拿住 巴力 的先知，不让任何人逃走！”众人就拿住他们。 以利亚 带他们到 基顺河 边，在那里杀了他们。
1KGS|18|41|以利亚 对 亚哈 说：“你现在可以上去吃喝，因为有暴雨的响声了。”
1KGS|18|42|亚哈 就上去吃喝。 以利亚 上了 迦密山 顶，屈身在地，把脸伏在两膝之中。
1KGS|18|43|他对仆人说：“你上去，向海观看。”仆人就上去观看，说：“没有什么。” 以利亚 说：“你再去。”如此七次。
1KGS|18|44|第七次，仆人说：“看哪，有一小片云从海里上来，好像人的手掌那么大。” 以利亚 说：“你上去告诉 亚哈 ，当套车下去，免得被雨阻挡。”
1KGS|18|45|霎时间，天因风云黑暗，降下大雨。 亚哈 就坐上车，往 耶斯列 去了。
1KGS|18|46|耶和华的手按在 以利亚 身上，他就束上腰，奔在 亚哈 前头，一路到 耶斯列 。
1KGS|19|1|亚哈 把 以利亚 一切所做的和他用刀杀众先知的事都告诉 耶洗别 。
1KGS|19|2|耶洗别 就派使者到 以利亚 那里，说：“明日约这时候，我若不使你的性命像那些人的性命一样，愿神明重重惩罚我。”
1KGS|19|3|以利亚 害怕 ，就起来逃命，到了 犹大 的 别是巴 ，把仆人留在那里。
1KGS|19|4|他自己在旷野走了一日的路程，来到一棵罗腾 树下，就坐在那里求死，说：“耶和华啊，现在够了！求你取我的性命吧，因为我不比我的祖先好。”
1KGS|19|5|他躺在罗腾树下睡着了。看哪，有一个天使拍他，对他说：“起来吃吧！”
1KGS|19|6|他观看，看哪，头旁有烧热的石头烤的饼和一壶水，他就吃了喝了，又再躺下。
1KGS|19|7|耶和华的使者回来，第二次拍他，说：“起来吃吧！因为你要走的路很远。”
1KGS|19|8|他就起来吃了喝了，仗着这饮食的力走了四十昼夜，到了上帝的山，就是 何烈山 。
1KGS|19|9|他在那里进了一个洞，在洞中过夜。看哪，耶和华的话临到他，说：“ 以利亚 ，你在这里做什么？”
1KGS|19|10|他说：“我为耶和华－万军之上帝大发热心，因为 以色列 人背弃了你的约，毁坏了你的坛，用刀杀了你的先知，只剩下我一人，他们还要追杀我。”
1KGS|19|11|耶和华说：“你出来站在山上，在耶和华面前。”看哪，耶和华从那里经过。在耶和华面前有烈风大作，山崩石裂，耶和华却不在风中；风后有地震，耶和华也不在其中；
1KGS|19|12|地震后有火，耶和华也不在火中；火以后，有轻微细小的声音。
1KGS|19|13|以利亚 听见，就用外衣蒙脸，出来站在洞口。听啊，有声音向他说：“ 以利亚 ，你在这里做什么？”
1KGS|19|14|他说：“我为耶和华－万军之上帝大发热心，因为 以色列 人背弃了你的约，毁坏了你的坛，用刀杀了你的先知，只剩下我一人，他们还要追杀我。”
1KGS|19|15|耶和华对他说：“去吧，从原路回去，往 大马士革 的旷野去。到了那里，你要膏 哈薛 作 亚兰 王，
1KGS|19|16|又膏 宁示 的孙子 耶户 作 以色列 王，并膏 亚伯．米何拉 人 沙法 的儿子 以利沙 作先知接续你。
1KGS|19|17|将来逃过 哈薛 之刀的，必被 耶户 所杀；逃过 耶户 之刀的，必被 以利沙 所杀。
1KGS|19|18|但我在 以色列 中留下七千人，是未曾向 巴力 屈膝，未曾亲吻 巴力 的。”
1KGS|19|19|于是， 以利亚 离开那里走了，遇见 沙法 的儿子 以利沙 ；他正在耕田，在他前头有十二对牛，自己赶着第十二对。 以利亚 经过他，把自己的外衣搭在他身上。
1KGS|19|20|以利沙 就离开牛，跑到 以利亚 那里，说：“请你让我先与父母吻别，然后我就跟随你。” 以利亚 对他说：“因我对你所做的事，你去吧，然后回来。 ”
1KGS|19|21|以利沙 离开他回去，宰了一对牛，用套牛的器具煮肉给百姓吃，随后就起身跟随 以利亚 ，服事他。
1KGS|20|1|亚兰 王 便．哈达 召集他的全军，率领三十二个王，带着马和战车，上来围困 撒玛利亚 ，要攻打它。
1KGS|20|2|他派使者进城到 以色列 王 亚哈 那里，对他说：“ 便．哈达 如此说：
1KGS|20|3|‘你的金银都要归我，你妻妾儿女中最美的也要归我。’”
1KGS|20|4|以色列 王回答说：“我主我王啊，就照着你的话，我和我所有的都归你。”
1KGS|20|5|使者又来说：“ 便．哈达 如此说：‘我已派人到你那里，要你把你的金银、妻妾、儿女都归我。’
1KGS|20|6|但明日约在这时候，我还要派臣仆到你那里，搜查你的家和你仆人的家，你眼中一切所喜爱的都由他们的手拿走。”
1KGS|20|7|以色列 王召了国内所有的长老来，说：“你们要知道，看哪，这人是来找麻烦的！他派人到我这里来，要我的妻妾、儿女和金银，我并没有拒绝他。”
1KGS|20|8|所有的长老和众百姓对王说：“不要听从他，也不要答应他。”
1KGS|20|9|以色列 王对 便．哈达 的使者说：“你们告诉我主我王说：‘王头一次派人向仆人所要的一切，仆人都依从，但这事我不能依从。’”使者就去回覆 便．哈达 。
1KGS|20|10|便．哈达 又派人到 亚哈 那里，说：“ 撒玛利亚 的尘土若足够跟从我的军兵每人手拿一把，愿神明重重惩罚我！”
1KGS|20|11|以色列 王回答说：“你们告诉他说，‘刚束上腰带的，不要像已卸下的那样夸口。’”
1KGS|20|12|便．哈达 和诸王正在帐幕里喝酒，听见这话，就对他臣仆说：“摆阵吧！”他们就摆阵攻城。
1KGS|20|13|看哪，一个先知靠近 以色列 王 亚哈 ，说：“耶和华如此说：‘这一大群人你看见了吗？看哪，今日我必把他们交在你手里，你就知道我是耶和华。’”
1KGS|20|14|亚哈 说：“藉着谁呢？”他说：“耶和华如此说：‘藉着跟从省长的年轻人。’” 亚哈 说：“谁要开战呢？”他说：“你！”
1KGS|20|15|于是 亚哈 数点跟从省长的年轻人，共二百三十二名，然后又数点 以色列 的众军兵，共七千名。
1KGS|20|16|中午，他们出了城； 便．哈达 和帮助他的三十二个王正在帐幕里畅饮。
1KGS|20|17|跟从省长的年轻人先出城。 便．哈达 派人去，他们回报说：“有人从 撒玛利亚 出来了。”
1KGS|20|18|他说：“他们若为求和出来，要活捉他们，若为打仗出来，也要活捉他们。”
1KGS|20|19|跟从省长的年轻人，和跟随他们的军兵，都出了城，
1KGS|20|20|各人遇见敌人就击杀。 亚兰 人逃跑， 以色列 人追赶他们； 亚兰 王 便．哈达 骑着马和骑兵一同逃跑。
1KGS|20|21|以色列 王出城攻击 马和战车，大大击杀 亚兰 人。
1KGS|20|22|那先知靠近 以色列 王，对他说：“去吧，你当自强，看清楚，也要知道你所要做的事，因为再过一年， 亚兰 王会上来攻击你。”
1KGS|20|23|亚兰 王的臣仆对他说：“他们的神是山神，所以他们胜过我们。但在平原与他们打仗，我们一定胜过他们。
1KGS|20|24|王当做这样的事，把诸王革去，派军官代替他们，
1KGS|20|25|又照着王丧失军兵的数目，再招募一支军队，马补马，车补车。然后在平原与他们打仗，我们一定胜过他们。”王就听臣仆的话，照样去做。
1KGS|20|26|过了一年， 便．哈达 果然召集 亚兰 人上 亚弗 去，要与 以色列 人打仗。
1KGS|20|27|以色列 人也召集军兵，预备食物，去迎战 亚兰 人。 以色列 人对着他们安营，好像两小群的山羊； 亚兰 人却布满了地面。
1KGS|20|28|有神人靠近，对 以色列 王说：“耶和华如此说：‘ 亚兰 人既说我－耶和华是山神，不是平原之神，我必将这一大群人全都交在你手中，你们就知道我是耶和华。’”
1KGS|20|29|以色列 人与 亚兰 人相对安营七日，到第七日两军开战。那一日 以色列 人杀了 亚兰 的十万步兵，
1KGS|20|30|其余的都逃向 亚弗 ，到了城里，城墙倒塌，压死了剩下的二万七千人。 便．哈达 也逃入城内，藏在严密的内室里。
1KGS|20|31|他的臣仆对他说：“看哪，我们听说 以色列 家的王都是仁慈的王；让我们腰束麻布，头套绳索，出去到 以色列 王那里，也许他会存留王的性命。”
1KGS|20|32|于是他们腰束麻布，头套绳索，来到 以色列 王那里，说：“王的仆人 便．哈达 说：‘求王饶我一命。’” 亚哈 说：“他还活着吗？他是我的兄弟。”
1KGS|20|33|这些人正在探测吉凶，就立即抓住他的话说：“ 便．哈达 是王的兄弟！”王说：“你们去请他来。” 便．哈达 出来到王那里，王就请他上车。
1KGS|20|34|便．哈达 对王说：“我父从你父那里所夺的城镇，我必归还给你。你可以在 大马士革 为你自己设立街市，像我父在 撒玛利亚 所设立的一样。” 亚哈 说：“我照此立约，放你回去。”王就与他立约，放了他。
1KGS|20|35|有一个人是先知的门徒，遵照耶和华的话对他同伴说：“你打我吧！”那人不肯打他。
1KGS|20|36|他就对那人说：“你既不听从耶和华的话，看哪，你一离开我，必有狮子咬死你。”那人一离开他，果然遇见狮子，把他咬死了。
1KGS|20|37|先知的门徒又遇见一个人，对他说：“你打我吧！”那人就打他，把他打伤。
1KGS|20|38|那先知就去了，用头巾蒙眼，改了装，在路旁等候王。
1KGS|20|39|王从那里经过，他向王呼叫说：“仆人出战的时候，看哪，有人转过来，带了一个人到我这里来，说：‘你要看守这人，若他真的失踪了，你的性命必代替他的性命，否则，你就要交出一他连得银子来。’
1KGS|20|40|仆人正在到处忙碌的时候，那人就不见了。” 以色列 王对他说：“你自己决定了，就必照样判你。”
1KGS|20|41|他急忙除掉蒙眼的头巾， 以色列 王就认出他是一个先知。
1KGS|20|42|他对王说：“耶和华如此说：‘因你把我决定要消灭的人从你手中放走，所以你的命必代替他的命，你的百姓必代替他的百姓。’”
1KGS|20|43|于是 以色列 王生气，忧闷地回 撒玛利亚 ，到自己的宫去了。
1KGS|21|1|这些事以后，又有一事。 耶斯列 人 拿伯 在 耶斯列 有一个葡萄园，靠近 撒玛利亚 ， 亚哈 王的宫。
1KGS|21|2|亚哈 对 拿伯 说：“把你的葡萄园给我作菜园，因为它靠近我的宫，我就把更好的葡萄园换给你。你若要银子，我就按着价钱给你。”
1KGS|21|3|拿伯 对 亚哈 说：“耶和华不准我把我祖先留下的产业给你。”
1KGS|21|4|亚哈 因 耶斯列 人 拿伯 说“我不把我祖先留下的产业给你”，就生气，忧闷地回宫，躺在床上，脸转向内，也不吃饭。
1KGS|21|5|耶洗别 王后来对他说：“你为什么心里这样生气，不吃饭呢？”
1KGS|21|6|他对王后说：“我向 耶斯列 人 拿伯 说：‘把你的葡萄园按价钱卖给我，或是你愿意，我可以把别的葡萄园换给你。’他却说：‘我不把我的葡萄园给你。’”
1KGS|21|7|耶洗别 王后对王说：“你现在是不是治理 以色列 国呢？只管起来，心里畅畅快快地吃饭，我会把 耶斯列 人 拿伯 的葡萄园给你。”
1KGS|21|8|于是王后以 亚哈 的名义写信，盖上王的印，把信送给那些与 拿伯 同城居住的长老和贵族。
1KGS|21|9|她在信上写着说：“你们当宣告禁食，叫 拿伯 坐在百姓的高位上，
1KGS|21|10|又叫两个无赖坐在 拿伯 对面，作证告他说：‘你诅咒了上帝和王。’然后把他拉出去用石头打死。”
1KGS|21|11|那些与 拿伯 同城居住的长老和贵族，照 耶洗别 送给他们的信去做。正如她送的信上所写，
1KGS|21|12|他们宣告禁食，叫 拿伯 坐在百姓的高位上。
1KGS|21|13|有两个无赖来，坐在 拿伯 对面。无赖当着百姓作证告他说：“ 拿伯 诅咒上帝和王了！”众人就把他拉到城外，用石头打他，他就死了。
1KGS|21|14|于是他们派人到 耶洗别 那里，说：“ 拿伯 被石头打死了。”
1KGS|21|15|耶洗别 听见 拿伯 被石头打死，就对 亚哈 说：“你起来，去取得 耶斯列 人 拿伯 不肯出价卖给你的葡萄园吧！因为 拿伯 不在了，他已经死了。”
1KGS|21|16|亚哈 听见 拿伯 死了，就起来，下去要取得 耶斯列 人 拿伯 的葡萄园。
1KGS|21|17|耶和华的话临到 提斯比 人 以利亚 ，说：
1KGS|21|18|“你起来，去见在 撒玛利亚 的 以色列 王 亚哈 。看哪，他下去要取得 拿伯 的葡萄园，他正在那园里。
1KGS|21|19|你要对他说：‘耶和华如此说：你杀了人，还要取得他的产业吗？’又要对他说：‘耶和华如此说：狗在何处舔 拿伯 的血，狗也必在何处舔你的血。’”
1KGS|21|20|亚哈 对 以利亚 说：“我的仇敌啊，你找到我了吗？”他说：“我找到你了。因为你出卖自己，行了耶和华眼中看为恶的事。
1KGS|21|21|耶和华说：‘看哪，我必使灾祸临到你，把你除灭。 以色列 中凡属 亚哈 的男丁，无论是奴役的、自由的，我都要剪除。
1KGS|21|22|我必使你的家像 尼八 的儿子 耶罗波安 的家，又像 亚希雅 的儿子 巴沙 的家，因为你惹我发怒，又使 以色列 陷入罪里。’
1KGS|21|23|论到 耶洗别 ，耶和华说：‘狗必在 耶斯列 的城郭 吃 耶洗别 。
1KGS|21|24|凡属 亚哈 的人，死在城中的必被狗吃，死在田野的必被空中的鸟吃。’”
1KGS|21|25|（只是从来没有像 亚哈 的，因他受 耶洗别 王后的唆使，出卖自己，行了耶和华眼中看为恶的事。
1KGS|21|26|他行了最可憎的事，随从偶像，正如耶和华在 以色列 人面前赶出的 亚摩利 人所行的一切。）
1KGS|21|27|亚哈 听见这些话，就撕裂衣服，禁食，贴身穿着麻布，也睡在麻布上，沮丧地走来走去。
1KGS|21|28|耶和华的话临到 提斯比 人 以利亚 ，说：
1KGS|21|29|“ 亚哈 在我面前这样谦卑，你看见了吗？因为他在我面前谦卑，所以在他的日子，我不降这祸；到他儿子的时候，我必降这祸于他的家。”
1KGS|22|1|亚兰 和 以色列 之间连续三年没有战争。
1KGS|22|2|到了第三年， 犹大 王 约沙法 下去见 以色列 王。
1KGS|22|3|以色列 王对臣仆说：“你们不知道 基列 的 拉末 是属我们的吗？我们岂可不采取行动，把它从 亚兰 王手里夺回来呢？”
1KGS|22|4|亚哈 问 约沙法 说：“你肯同我去攻打 基列 的 拉末 吗？” 约沙法 对 以色列 王说：“你我不分彼此，我的军队就是你的军队，我的马就是你的马。”
1KGS|22|5|约沙法 对 以色列 王说：“请你先求问耶和华的话。”
1KGS|22|6|于是 以色列 王召集先知，约有四百人，问他们说：“我可以上去攻打 基列 的 拉末 吗？还是不要上去呢？”他们说：“可以上去，因为主必将那城交在王的手里。”
1KGS|22|7|约沙法 说：“这里还有没有耶和华的先知，我们好求问他呢？”
1KGS|22|8|以色列 王对 约沙法 说：“还有一个人，是 音拉 的儿子 米该雅 ，我们可以托他求问耶和华。只是我真的很恨他，因为他对我说预言，从不说吉言，总是说凶信。” 约沙法 说：“请王不要这么说。”
1KGS|22|9|以色列 王召了一个官员来，说：“你快去，把 音拉 的儿子 米该雅 召来。”
1KGS|22|10|以色列 王和 犹大 王 约沙法 在 撒玛利亚 城门前的禾场，各穿朝服，坐在宝座上，所有的先知都在他们面前说预言。
1KGS|22|11|基拿拿 的儿子 西底家 造了铁角，说：“耶和华如此说：‘你要用这些角抵触 亚兰 人，直到将他们灭尽。’”
1KGS|22|12|所有的先知也都这样预言说：“可以上 基列 的 拉末 去，必然得胜，因为耶和华必将那城交在王的手中。”
1KGS|22|13|那去召 米该雅 的使者对他说：“看哪，众先知都异口同声向王说吉言，你也跟他们说一样的话，说吉言吧！”
1KGS|22|14|米该雅 说：“我指着永生的耶和华起誓，耶和华向我说什么，我就说什么。”
1KGS|22|15|米该雅 来到王那里，王问他：“ 米该雅 ，我们可以上去攻打 基列 的 拉末 吗？还是不要上去呢？”他对王说：“你可以上去，必然得胜，耶和华必将那城交在王的手中。”
1KGS|22|16|王对他说：“我要你发誓多少次，你才会奉耶和华的名向我说实话呢？”
1KGS|22|17|米该雅 说：“我看见 以色列 众人散布在山上，如同没有牧人的羊群一般。耶和华说：‘这些人没有主人，他们可以平安地各自回家去。’”
1KGS|22|18|以色列 王对 约沙法 说：“我岂没有告诉你，这人对我说预言，从不说吉言，只说凶信吗？”
1KGS|22|19|米该雅 说：“因此你要听耶和华的话！我看见耶和华坐在宝座上，天上的万军侍立在他左右。
1KGS|22|20|耶和华说：‘谁去引诱 亚哈 上 基列 的 拉末 去阵亡呢？’这个这样说，那个那样说。
1KGS|22|21|随后有一个灵出来，站在耶和华面前，说：‘我去引诱他。’
1KGS|22|22|耶和华问他：‘用什么方法呢？’他说：‘我要出去，在他众先知的口中成为谎言的灵。’耶和华说：‘这样，你去引诱他，必能成功。你出去，照样做吧！’
1KGS|22|23|现在，看哪，耶和华使谎言的灵入了你所有的这些先知的口，并且耶和华已经宣告要降祸于你。”
1KGS|22|24|基拿拿 的儿子 西底家 前来，打 米该雅 一巴掌，说：“耶和华的灵从哪里离开我向你说话呢？”
1KGS|22|25|米该雅 说：“看哪，你进入严密的内室躲藏的那日，就必看见。”
1KGS|22|26|以色列 王说：“把 米该雅 带走，交回给 亚们 市长和 约阿施 王子。
1KGS|22|27|你们要说：‘王如此说，把这个人关在监狱里，使他受苦，吃不饱喝不足，直等到我平安回来。’”
1KGS|22|28|米该雅 说：“你若真的能平安回来，那就是耶和华没有藉我说这话了。”他又说：“众百姓啊，你们都要听！”
1KGS|22|29|以色列 王和 犹大 王 约沙法 上 基列 的 拉末 去。
1KGS|22|30|以色列 王对 约沙法 说：“我要改装上阵，你可以仍穿王袍。” 以色列 王就改装上阵去了。
1KGS|22|31|亚兰 王吩咐他的三十二个战车长说：“你们不要与他们的大将或小兵交战，只要单单攻击 以色列 王。”
1KGS|22|32|那些战车长看见 约沙法 就说：“这一定是 以色列 王！”他们转过去与他交战， 约沙法 就呼喊起来。
1KGS|22|33|战车长见他不是 以色列 王，就转身不追他了。
1KGS|22|34|有一人开弓，并不知情，箭恰巧射入 以色列 王铠甲的缝里。王对驾车的说：“我受重伤了，你掉过车来，载我离开战场！”
1KGS|22|35|那日，战况越来越猛，有人扶着王站在战车上，面对 亚兰 人。到了傍晚，王就死了，血从伤处流入车底。
1KGS|22|36|约在日落的时候，有喊声传遍军中，说：“大家各归本城，各归本地吧！”
1KGS|22|37|王死了，人把他送到 撒玛利亚 ，葬在 撒玛利亚 。
1KGS|22|38|他们在 撒玛利亚 的水池旁洗他的车，有狗来舔他的血，有妓女在那里洗澡，正如耶和华所说的话。
1KGS|22|39|亚哈 其余的事，凡他所做的、他所修造的象牙宫和所建筑的一切城镇，不都写在《以色列诸王记》上吗？
1KGS|22|40|亚哈 与他祖先同睡，他儿子 亚哈谢 接续他作王。
1KGS|22|41|以色列 王 亚哈 第四年， 亚撒 的儿子 约沙法 登基作 犹大 王。
1KGS|22|42|约沙法 登基的时候年三十五岁，在 耶路撒冷 作王二十五年。他母亲名叫 阿苏巴 ，是 示利希 的女儿。
1KGS|22|43|约沙法 效法他父亲 亚撒 所行的道，不偏离左右，行耶和华眼中看为正的事。只是丘坛还没有废去，百姓仍在那里献祭烧香。
1KGS|22|44|约沙法 与 以色列 王和平相处。
1KGS|22|45|约沙法 其余的事和他所行的英勇事迹，以及他的战役，不都写在《犹大列王记》上吗？
1KGS|22|46|约沙法 把他父亲 亚撒 的日子所剩下男的庙妓都从国中除去了。
1KGS|22|47|那时 以东 没有立王，由总督治理。
1KGS|22|48|约沙法 造了 他施 船只，要往 俄斐 去，把金子运来，却没有启航，因为船在 以旬．迦别 毁坏了。
1KGS|22|49|亚哈 的儿子 亚哈谢 对 约沙法 说：“让我的仆人和你的仆人坐船同去吧！” 约沙法 却不肯。
1KGS|22|50|约沙法 与他祖先同睡，与他祖先同葬在 大卫城 ，他儿子 约兰 接续他作王。
1KGS|22|51|犹大 王 约沙法 第十七年， 亚哈 的儿子 亚哈谢 在 撒玛利亚 登基作 以色列 王；他作 以色列 王二年。
1KGS|22|52|他行耶和华眼中看为恶的事，行他父母的道，又行 尼八 的儿子 耶罗波安 的道，使 以色列 陷入罪里。
1KGS|22|53|他事奉 巴力 ，敬拜它，惹耶和华－ 以色列 的上帝发怒，正如他父亲一切所行的。
