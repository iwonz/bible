EZRA|1|1|in anno primo Cyri regis Persarum ut conpleretur verbum Domini ex ore Hieremiae suscitavit Dominus spiritum Cyri regis Persarum et transduxit vocem in universo regno suo etiam per scripturam dicens
EZRA|1|2|haec dicit Cyrus rex Persarum omnia regna terrae dedit mihi Dominus Deus caeli et ipse praecepit mihi ut aedificarem ei domum in Hierusalem quae est in Iudaea
EZRA|1|3|quis est in vobis de universo populo eius sit Deus illius cum ipso ascendat Hierusalem quae est in Iudaea et aedificet domum Domini Dei Israhel ipse est Deus qui est in Hierusalem
EZRA|1|4|et omnes reliqui in cunctis locis ubicumque habitant adiuvent eum viri de loco suo argento et auro et substantia et pecoribus excepto quod voluntarie offerunt templo Dei quod est in Hierusalem
EZRA|1|5|et surrexerunt principes patrum de Iuda et Beniamin et sacerdotes et Levitae omnis cuius suscitavit Deus spiritum ut ascenderent ad aedificandum templum Domini quod erat in Hierusalem
EZRA|1|6|universique qui erant in circuitu adiuverunt manus eorum in vasis argenteis et aureis in substantia in iumentis in supellectili exceptis his quae sponte obtulerunt
EZRA|1|7|rex quoque Cyrus protulit vasa templi Domini quae tulerat Nabuchodonosor de Hierusalem et posuerat ea in templo dei sui
EZRA|1|8|protulit autem ea Cyrus rex Persarum per manum Mitridatis filii Gazabar et adnumeravit ea Sasabassar principi Iudae
EZRA|1|9|et hic est numerus eorum fialae aureae triginta fialae argenteae mille cultri viginti novem scyphi aurei triginta
EZRA|1|10|scyphi argentei secundi quadringenti decem vasa alia mille
EZRA|1|11|omnia vasa aurea et argentea quinque milia quadringenta universa tulit Sasabassar cum his qui ascendebant de transmigratione Babylonis in Hierusalem
EZRA|2|1|hii sunt autem filii provinciae qui ascenderunt de captivitate quam transtulerat Nabuchodonosor rex Babylonis in Babylonem et reversi sunt in Hierusalem et Iudam unusquisque in civitatem suam
EZRA|2|2|qui venerunt cum Zorobabel Hiesua Neemia Saraia Rahelaia Mardochai Belsan Mesphar Beguai Reum Baana numerus virorum populi Israhel
EZRA|2|3|filii Pharos duo milia centum septuaginta duo
EZRA|2|4|filii Sephetia trecenti septuaginta duo
EZRA|2|5|filii Area septingenti septuaginta quinque
EZRA|2|6|filii Phaethmoab filiorum Iosue Ioab duo milia octingenti duodecim
EZRA|2|7|filii Helam mille ducenti quinquaginta quattuor
EZRA|2|8|filii Zeththua nongenti quadraginta quinque
EZRA|2|9|filii Zacchai septingenti sexaginta
EZRA|2|10|filii Bani sescenti quadraginta duo
EZRA|2|11|filii Bebai sescenti viginti tres
EZRA|2|12|filii Azgad mille ducenti viginti duo
EZRA|2|13|filii Adonicam sescenti sexaginta sex
EZRA|2|14|filii Beguai duo milia quinquaginta sex
EZRA|2|15|filii Adin quadringenti quinquaginta quattuor
EZRA|2|16|filii Ater qui erant ex Hiezechia nonaginta octo
EZRA|2|17|filii Besai trecenti viginti tres
EZRA|2|18|filii Iora centum duodecim
EZRA|2|19|filii Asom ducenti viginti tres
EZRA|2|20|filii Gebbar nonaginta quinque
EZRA|2|21|filii Bethleem centum viginti tres
EZRA|2|22|viri Netupha quinquaginta sex
EZRA|2|23|viri Anathoth centum viginti octo
EZRA|2|24|filii Azmaveth quadraginta duo
EZRA|2|25|filii Cariathiarim Caephira et Beroth septingenti quadraginta tres
EZRA|2|26|filii Arama et Gaba sescenti viginti unus
EZRA|2|27|viri Machmas centum viginti duo
EZRA|2|28|viri Bethel et Gai ducenti viginti tres
EZRA|2|29|filii Nebo quinquaginta duo
EZRA|2|30|filii Megbis centum quinquaginta sex
EZRA|2|31|filii Helam alterius mille ducenti quinquaginta quattuor
EZRA|2|32|filii Arim trecenti viginti
EZRA|2|33|filii Lod Adid et Ono septingenti viginti quinque
EZRA|2|34|filii Hiericho trecenti quadraginta quinque
EZRA|2|35|filii Sennaa tria milia sescenti triginta
EZRA|2|36|sacerdotes filii Idaia in domo Hiesue nongenti septuaginta tres
EZRA|2|37|filii Emmer mille quinquaginta duo
EZRA|2|38|filii Phessur mille ducenti quadraginta septem
EZRA|2|39|filii Arim mille decem et septem
EZRA|2|40|Levitae filii Hiesue et Cedmihel filiorum Odevia septuaginta quattuor
EZRA|2|41|cantores filii Asaph centum viginti octo
EZRA|2|42|filii ianitorum filii Sellum filii Ater filii Telmon filii Accub filii Atita filii Sobai universi centum triginta novem
EZRA|2|43|Nathinnei filii Sia filii Asupha filii Tebbaoth
EZRA|2|44|filii Ceros filii Siaa filii Phadon
EZRA|2|45|filii Levana filii Agaba filii Accub
EZRA|2|46|filii Agab filii Selmai filii Anan
EZRA|2|47|filii Gaddel filii Gaer filii Rahaia
EZRA|2|48|filii Rasin filii Nechoda filii Gazem
EZRA|2|49|filii Aza filii Phasea filii Besee
EZRA|2|50|filii Asenaa filii Munim filii Nephusim
EZRA|2|51|filii Becbuc filii Acupha filii Arur
EZRA|2|52|filii Besluth filii Maida filii Arsa
EZRA|2|53|filii Bercos filii Sisara filii Thema
EZRA|2|54|filii Nasia filii Atupha
EZRA|2|55|filii servorum Salomonis filii Sotei filii Suphereth filii Pharuda
EZRA|2|56|filii Iala filii Dercon filii Gedel
EZRA|2|57|filii Saphatia filii Athil filii Phocereth qui erant de Asebaim filii Ammi
EZRA|2|58|omnes Nathinnei et filii servorum Salomonis trecenti nonaginta duo
EZRA|2|59|et hii qui ascenderunt de Thelmela Thelarsa Cherub et Don et Mer et non potuerunt indicare domum patrum suorum et semen suum utrum ex Israhel essent
EZRA|2|60|filii Delaia filii Tobia filii Necoda sescenti quinquaginta duo
EZRA|2|61|et de filiis sacerdotum filii Obia filii Accos filii Berzellai qui accepit de filiabus Berzellai Galaditis uxorem et vocatus est nomine eorum
EZRA|2|62|hii quaesierunt scripturam genealogiae suae et non invenerunt et eiecti sunt de sacerdotio
EZRA|2|63|et dixit Athersatha eis ut non comederent de sancto sanctorum donec surgeret sacerdos doctus atque perfectus
EZRA|2|64|omnis multitudo quasi unus quadraginta duo milia trecenti sexaginta
EZRA|2|65|exceptis servis eorum et ancillis qui erant septem milia trecenti triginta septem et in ipsis cantores atque cantrices ducentae
EZRA|2|66|equi eorum septingenti triginta sex muli eorum ducenti quadraginta quinque
EZRA|2|67|cameli eorum quadringenti triginta quinque asini eorum sex milia septingenti viginti
EZRA|2|68|et de principibus patrum cum ingrederentur templum Domini quod est in Hierusalem sponte obtulerunt in domum Dei ad extruendam eam in loco suo
EZRA|2|69|secundum vires suas dederunt in inpensas operis auri solidos sexaginta milia et mille argenti minas quinque milia et vestes sacerdotales centum
EZRA|2|70|habitaverunt ergo sacerdotes et Levitae et de populo et cantores et ianitores et Nathinnei in urbibus suis universusque Israhel in civitatibus suis
EZRA|3|1|iamque venerat mensis septimus et erant filii Israhel in civitatibus suis congregatus est ergo populus quasi vir unus in Hierusalem
EZRA|3|2|et surrexit Iosue filius Iosedech et fratres eius sacerdotes et Zorobabel filius Salathihel et fratres eius et aedificaverunt altare Dei Israhel ut offerrent in eo holocaustomata sicut scriptum est in lege Mosi viri Dei
EZRA|3|3|conlocaverunt autem altare super bases suas deterrentibus eos per circuitum populis terrarum et obtulerunt super illud holocaustum Domino mane et vespere
EZRA|3|4|feceruntque sollemnitatem tabernaculorum sicut scriptum est et holocaustum diebus singulis per ordinem secundum praeceptum opus diei in die suo
EZRA|3|5|et post haec holocaustum iuge tam in kalendis quam in universis sollemnitatibus Domini quae erant consecratae et in omnibus in quibus ultro offerebatur munus Deo
EZRA|3|6|a primo die mensis septimi coeperunt offerre holocaustum Domino porro templum Dei fundatum necdum erat
EZRA|3|7|dederunt autem pecunias latomis et cementariis cibum quoque et potum et oleum Sidoniis Tyriisque ut deferrent ligna cedrina de Libano ad mare Ioppes iuxta quod praeceperat Cyrus rex Persarum eis
EZRA|3|8|anno autem secundo adventus eorum ad templum Dei in Hierusalem mense secundo coeperunt Zorobabel filius Salathihel et Iosue filius Iosedech et reliqui de fratribus eorum sacerdotes et Levitae et omnes qui venerant de captivitate in Hierusalem et constituerunt Levitas a viginti annis et supra ut urguerent opus Domini
EZRA|3|9|stetitque Iosue filii eius et fratres eius Cedmihel et filii eius et filii Iuda quasi unus ut instarent super eos qui faciebant opus in templo Dei filii Enadad filii eorum et fratres eorum Levitae
EZRA|3|10|fundato igitur a cementariis templo Domini steterunt sacerdotes in ornatu suo cum tubis et Levitae filii Asaph in cymbalis ut laudarent Deum per manus David regis Israhel
EZRA|3|11|et concinebant in hymnis et confessione Domino quoniam bonus quoniam in aeternum misericordia eius super Israhel omnis quoque populus vociferabatur clamore magno in laudando Dominum eo quod fundatum esset templum Domini
EZRA|3|12|plurimi etiam de sacerdotibus et Levitis et principes patrum seniores qui viderant templum prius cum fundatum esset et hoc templum in oculis eorum flebant voce magna et multi vociferantes in laetitia elevabant vocem
EZRA|3|13|nec poterat quisquam agnoscere vocem clamoris laetantium et vocem fletus populi commixtim enim populus vociferabatur clamore magno et vox audiebatur procul
EZRA|4|1|audierunt autem hostes Iudae et Beniamin quia filii captivitatis aedificarent templum Domino Deo Israhel
EZRA|4|2|et accedentes ad Zorobabel et ad principes patrum dixerunt eis aedificemus vobiscum quia ita ut vos quaerimus Deum vestrum ecce nos immolamus victimas ex diebus Asoraddan regis Assur qui adduxit nos huc
EZRA|4|3|et dixit eis Zorobabel et Iosue et reliqui principes patrum Israhel non est vobis et nobis ut aedificemus domum Deo nostro sed nos ipsi soli aedificabimus Domino Deo nostro sicut praecepit nobis rex Cyrus rex Persarum
EZRA|4|4|factum est igitur ut populus terrae inpediret manus populi Iudae et turbaret eos in aedificando
EZRA|4|5|conduxerunt quoque adversum eos consiliatores ut destruerent consilium eorum omnibus diebus Cyri regis Persarum et usque ad regnum Darii regis Persarum
EZRA|4|6|in regno autem Asueri principio regni eius scripserunt accusationem adversum habitatores Iudae et Hierusalem
EZRA|4|7|et in diebus Artarxersis scripsit Beselam Mitridatis et Tabel et reliqui qui erant in consilio eorum ad Artarxersen regem Persarum epistula autem accusationis scripta erat syriace et legebatur sermone syro
EZRA|4|8|Reum Beelteem et Samsai scriba scripserunt epistulam unam de Hierusalem Artarxersi regi huiuscemodi
EZRA|4|9|Reum Beelteem et Samsai scriba et reliqui consiliatores eorum Dinei et Apharsathei Terphalei Apharsei Erchuei Babylonii Susannechei Deaei Aelamitae
EZRA|4|10|et ceteri de gentibus quas transtulit Asennaphar magnus et gloriosus et habitare eas fecit in civitatibus Samariae et in reliquis regionibus trans Flumen in pace
EZRA|4|11|hoc est exemplar epistulae quam miserunt ad eum Artarxersi regi servi tui viri qui sunt trans Fluvium salutem dicunt
EZRA|4|12|notum sit regi quia Iudaei qui ascenderunt a te ad nos venerunt in Hierusalem civitatem rebellem et pessimam quam aedificant extruentes muros eius et parietes conponentes
EZRA|4|13|nunc igitur notum sit regi quia si civitas illa aedificata fuerit et muri eius instaurati tributum et vectigal et annuos reditus non dabunt et usque ad reges haec noxa perveniet
EZRA|4|14|nos ergo memores salis quod in palatio comedimus et quia laesiones regis videre nefas ducimus idcirco misimus et nuntiavimus regi
EZRA|4|15|ut recenseas in libris historiarum patrum tuorum et invenies scriptum in commentariis et scies quoniam urbs illa urbs rebellis est et nocens regibus et provinciis et bella concitant in ea ex diebus antiquis quam ob rem et civitas ipsa destructa est
EZRA|4|16|nuntiamus nos regi quoniam si civitas illa aedificata fuerit et muri ipsius instaurati possessionem trans Fluvium non habebis
EZRA|4|17|verbum misit rex ad Reum Beelteem et Samsai scribam et ad reliquos qui erant in consilio eorum habitatores Samariae et ceteris trans Fluvium salutem dicens et pacem
EZRA|4|18|accusationem quam misistis ad nos manifeste lecta est coram me
EZRA|4|19|et a me praeceptum est et recensuerunt inveneruntque quoniam civitas illa a diebus antiquis adversum reges rebellat et seditiones et proelia concitantur in ea
EZRA|4|20|nam et reges fortissimi fuerunt in Hierusalem qui et dominati sunt omni regioni quae trans Fluvium est tributum quoque et vectigal et reditus accipiebant
EZRA|4|21|nunc ergo audite sententiam ut prohibeatis viros illos et urbs illa non aedificetur donec si forte a me iussum fuerit
EZRA|4|22|videte ne neglegenter hoc impleatis et paulatim crescat malum contra reges
EZRA|4|23|itaque exemplum edicti Artarxersis regis lectum est coram Reum et Samsai scriba et consiliariis eorum et abierunt festini in Hierusalem ad Iudaeos et prohibuerunt eos in brachio et robore
EZRA|4|24|tunc intermissum est opus domus Dei in Hierusalem et non fiebat usque ad annum secundum regni Darii regis Persarum
EZRA|5|1|prophetaverunt autem Aggeus propheta et Zaccharias filius Addo prophetantes ad Iudaeos qui erant in Iudaea et Hierusalem in nomine Dei Israhel
EZRA|5|2|tunc surrexerunt Zorobabel filius Salathihel et Iosue filius Iosedech et coeperunt aedificare templum Dei in Hierusalem et cum eis prophetae Dei adiuvantes eos
EZRA|5|3|in ipso tempore venit ad eos Tatannai qui erat dux trans Flumen et Starbuzannai et consiliarii eorum sicque dixerunt eis quis dedit vobis consilium ut domum hanc aedificaretis et muros hos instauraretis
EZRA|5|4|ad quod respondimus eis quae essent nomina hominum auctorum illius aedificationis
EZRA|5|5|oculus autem Dei eorum factus est super senes Iudaeorum et non potuerunt inhibere eos placuitque ut res ad Darium referretur et tunc satisfacerent adversus accusationem illam
EZRA|5|6|exemplar epistulae quam misit Tatannai dux regionis trans Flumen et Starbuzannai et consiliatores eius Apharsacei qui erant trans Flumen ad Darium regem
EZRA|5|7|sermo quem miserant ei sic scriptus erat Dario regi pax omnis
EZRA|5|8|notum sit regi isse nos ad Iudaeam provinciam ad domum Dei magni quae aedificatur lapide inpolito et ligna ponuntur in parietibus opusque illud diligenter extruitur et crescit in manibus eorum
EZRA|5|9|interrogavimus ergo senes illos et ita diximus eis quis dedit vobis potestatem ut domum hanc aedificaretis et muros instauraretis
EZRA|5|10|sed et nomina eorum quaesivimus ab eis ut nuntiaremus tibi quae scripsimus nomina virorum qui sunt principes in eis
EZRA|5|11|huiuscemodi autem sermonem responderunt nobis dicentes nos sumus servi Dei caeli et terrae et aedificamus templum quod erat extructum ante hos annos multos quodque rex Israhel magnus aedificaverat et extruxerat
EZRA|5|12|postquam autem ad iracundiam provocaverunt patres nostri Deum caeli et tradidit eos in manu Nabuchodonosor regis Babylonis Chaldei domum quoque hanc destruxit et populum eius transtulit in Babylonem
EZRA|5|13|anno autem primo Cyri regis Babylonis Cyrus rex proposuit edictum ut domus Dei aedificaretur
EZRA|5|14|nam et vasa templi Dei aurea et argentea quae Nabuchodonosor tulerat de templo quod erat in Hierusalem et asportaverat ea in templum Babylonis protulit Cyrus rex de templo Babylonis et data sunt Sasabassar vocabulo quem et principem constituit
EZRA|5|15|dixitque ei haec vasa tolle et vade et pone ea in templo quod est in Hierusalem et domus Dei aedificetur in loco suo
EZRA|5|16|tunc itaque Sasabassar ille venit et posuit fundamenta templi Dei in Hierusalem et ex eo tempore usque nunc aedificatur et necdum conpletum est
EZRA|5|17|nunc ergo si videtur regi bonum recenseat in bibliotheca regis quae est in Babylone utrumnam a Cyro rege iussum sit ut aedificaretur domus Dei in Hierusalem et voluntatem regis super hac re mittat ad nos
EZRA|6|1|tunc Darius rex praecepit et recensuerunt in bibliotheca librorum qui erant repositi in Babylone
EZRA|6|2|et inventum est in Ecbathanis quod est castrum in Madena provincia volumen unum talisque scriptus erat in eo commentarius
EZRA|6|3|anno primo Cyri regis Cyrus rex decrevit ut domus Dei quae est in Hierusalem aedificaretur in loco ubi immolent hostias et ut ponant fundamenta subportantia altitudinem cubitorum sexaginta et latitudinem cubitorum sexaginta
EZRA|6|4|ordines de lapidibus inpolitis tres et sic ordines de lignis novis sumptus autem de domo regis dabuntur
EZRA|6|5|sed et vasa templi Dei aurea et argentea quae Nabuchodonosor tulerat de templo Hierusalem et adtulerat ea in Babylonem reddantur et referantur in templo Hierusalem in locum suum quae et posita sunt in templo Dei
EZRA|6|6|nunc ergo Tatannai dux regionis quae est trans Flumen Starbuzannai et consiliarii vestri Apharsacei qui estis trans Flumen procul recedite ab illis
EZRA|6|7|et dimittite fieri templum Dei illud a duce Iudaeorum et a senioribus eorum domum Dei illam aedificent in loco suo
EZRA|6|8|sed et a me praeceptum est quid oporteat fieri a presbyteris Iudaeorum illis ut aedificetur domus Dei scilicet ut de arca regis id est de tributis quae dantur de regione trans Flumen studiose sumptus dentur viris illis ne inpediatur opus
EZRA|6|9|quod si necesse fuerit et vitulos et agnos et hedos in holocaustum Deo caeli frumentum sal vinum et oleum secundum ritum sacerdotum qui sunt in Hierusalem detur eis per dies singulos ne sit in aliquo querimonia
EZRA|6|10|et offerant oblationes Deo caeli orentque pro vita regis et filiorum eius
EZRA|6|11|a me ergo positum est decretum ut omnis homo qui hanc mutaverit iussionem tollatur lignum de domo ipsius et erigatur et configatur in eo domus autem eius publicetur
EZRA|6|12|Deus autem qui habitare fecit nomen suum ibi dissipet omnia regna et populum qui extenderit manum suam ut repugnet et dissipet domum Dei illam quae est in Hierusalem ego Darius statui decretum quod studiose impleri volo
EZRA|6|13|igitur Tatannai dux regionis trans Flumen et Starbuzannai et consiliarii eius secundum quod praeceperat Darius rex sic diligenter exsecuti sunt
EZRA|6|14|seniores autem Iudaeorum aedificabant et prosperabantur iuxta prophetiam Aggei prophetae et Zacchariae filii Addo et aedificaverunt et construxerunt iubente Deo Israhel et iubente Cyro et Dario et Artarxerse regibus Persarum
EZRA|6|15|et conpleverunt domum Dei istam usque ad diem tertium mensis adar qui est annus sextus regni Darii regis
EZRA|6|16|fecerunt autem filii Israhel sacerdotes et Levitae et reliqui filiorum transmigrationis dedicationem domus Dei in gaudio
EZRA|6|17|et obtulerunt in dedicationem domus Dei vitulos centum arietes ducentos agnos quadringentos hircos caprarum pro peccato totius Israhel duodecim iuxta numerum tribuum Israhel
EZRA|6|18|et statuerunt sacerdotes in ordinibus suis et Levitas in vicibus suis super opera Dei in Hierusalem sicut scriptum est in libro Mosi
EZRA|6|19|fecerunt autem filii transmigrationis pascha quartadecima die mensis primi
EZRA|6|20|purificati enim fuerant sacerdotes et Levitae quasi unus omnes mundi ad immolandum pascha universis filiis transmigrationis et fratribus suis sacerdotibus et sibi
EZRA|6|21|et comederunt filii Israhel qui reversi fuerant de transmigratione et omnis qui se separaverat a coinquinatione gentium terrae ad eos ut quaererent Dominum Deum Israhel
EZRA|6|22|et fecerunt sollemnitatem azymorum septem diebus in laetitia quoniam laetificaverat eos Dominus et converterat cor regis Assur ad eos ut adiuvaret manus eorum in opere domus Domini Dei Israhel
EZRA|7|1|post haec autem verba in regno Artarxersis regis Persarum Ezras filius Saraiae filii Azariae filii Helciae
EZRA|7|2|filii Sellum filii Sadoc filii Achitob
EZRA|7|3|filii Amariae filii Azariae filii Maraioth
EZRA|7|4|filii Zaraiae filii Ozi filii Bocci
EZRA|7|5|filii Abisue filii Finees filii Eleazar filii Aaron sacerdotis ab initio
EZRA|7|6|ipse Ezras ascendit de Babylone et ipse scriba velox in lege Mosi quam dedit Dominus Deus Israhel et dedit ei rex secundum manum Domini Dei eius super eum omnem petitionem eius
EZRA|7|7|et ascenderunt de filiis Israhel et de filiis sacerdotum et de filiis Levitarum et de cantoribus et de ianitoribus et de Nathinneis in Hierusalem anno septimo Artarxersis regis
EZRA|7|8|et venerunt in Hierusalem mense quinto ipse est annus septimus regis
EZRA|7|9|quia in primo die mensis primi coepit ascendere de Babylone et in primo mensis quinti venit in Hierusalem iuxta manum Dei sui bonam super se
EZRA|7|10|Ezras enim paravit cor suum ut investigaret legem Domini et faceret et doceret in Israhel praeceptum et iudicium
EZRA|7|11|hoc est autem exemplar epistulae edicti quod dedit rex Artarxersis Ezrae sacerdoti scribae erudito in sermonibus et praeceptis Domini et caerimoniis eius in Israhel
EZRA|7|12|Artarxersis rex regum Ezrae sacerdoti scribae legis Dei caeli doctissimo salutem
EZRA|7|13|a me decretum est ut cuicumque placuerit in regno meo de populo Israhel et de sacerdotibus eius et de Levitis ire in Hierusalem tecum vadat
EZRA|7|14|a facie enim regis et septem consiliatorum eius missus es ut visites Iudaeam et Hierusalem in lege Dei tui quae est in manu tua
EZRA|7|15|et ut feras argentum et aurum quod rex et consiliatores eius sponte obtulerunt Deo Israhel cuius in Hierusalem tabernaculum est
EZRA|7|16|et omne argentum et aurum quodcumque inveneris in universa provincia Babylonis et populus offerre voluerit et de sacerdotibus qui sponte obtulerint domui Dei sui quae est in Hierusalem
EZRA|7|17|libere accipe et studiose eme de hac pecunia vitulos arietes agnos et sacrificia et libamina eorum et offer ea super altare templi Dei vestri quod est in Hierusalem
EZRA|7|18|sed et si quid tibi et fratribus tuis placuerit de reliquo argento et auro ut faciatis iuxta voluntatem Dei vestri facite
EZRA|7|19|vasa quoque quae dantur tibi in ministerium domus Dei tui trade in conspectu Dei Hierusalem
EZRA|7|20|sed et cetera quibus opus fuerit in domo Dei tui quantumcumque necesse est ut expendas dabis de thesauro et de fisco regis
EZRA|7|21|et a me ego Artarxersis rex statui atque decrevi omnibus custodibus arcae publicae qui sunt trans Flumen ut quodcumque petierit a vobis Ezras sacerdos scriba legis Dei caeli absque mora detis
EZRA|7|22|usque ad argenti talenta centum et usque ad frumenti choros centum et usque ad vini batos centum et usque ad batos olei centum sal vero absque mensura
EZRA|7|23|omne quod ad ritum Dei caeli pertinet tribuatur diligenter in domo Dei caeli ne forte irascatur contra regnum regis et filiorum eius
EZRA|7|24|vobisque notum facimus de universis sacerdotibus et Levitis cantoribus ianitoribus Nathinneis et ministris domus Dei huius ut vectigal et tributum et annonas non habeatis potestatem inponendi super eos
EZRA|7|25|tu autem Ezras secundum sapientiam Dei tui quae est in manu tua constitue iudices et praesides ut iudicent omni populo qui est trans Flumen his videlicet qui noverunt legem Dei tui sed et inperitos docete libere
EZRA|7|26|et omnis qui non fecerit legem Dei tui et legem regis diligenter iudicium erit de eo sive in mortem sive in exilium sive in condemnationem substantiae eius vel certe in carcerem
EZRA|7|27|benedictus Dominus Deus patrum nostrorum qui dedit hoc in corde regis ut glorificaret domum Domini quae est in Hierusalem
EZRA|7|28|et in me inclinavit misericordiam coram rege et consiliatoribus eius et universis principibus regis potentibus et ego confortatus manu Domini Dei mei quae erat in me congregavi de Israhel principes qui ascenderent mecum
EZRA|8|1|hii sunt ergo principes familiarum et genealogia eorum qui ascenderunt mecum in regno Artarxersis regis de Babylone
EZRA|8|2|de filiis Finees Gersom de filiis Ithamar Danihel de filiis David Attus
EZRA|8|3|de filiis Secheniae et de filiis Pharos Zaccharias et cum eo numerati sunt viri centum quinquaginta
EZRA|8|4|de filiis Phaethmoab Helioenai filius Zareae et cum eo ducenti viri
EZRA|8|5|de filiis Secheniae filius Hiezihel et cum eo trecenti viri
EZRA|8|6|de filiis Adden Abeth filius Ionathan et cum eo quinquaginta viri
EZRA|8|7|de filiis Helam Isaias filius Athaliae et cum eo septuaginta viri
EZRA|8|8|de filiis Saphatiae Zebedia filius Michahel et cum eo octoginta viri
EZRA|8|9|de filiis Ioab Obedia filius Iehihel et cum eo ducenti decem et octo viri
EZRA|8|10|de filiis Selomith filius Iosphiae et cum eo centum sexaginta viri
EZRA|8|11|de filiis Bebai Zaccharias filius Bebai et cum eo viginti octo viri
EZRA|8|12|de filiis Ezgad Iohanan filius Eccetan et cum eo centum decem viri
EZRA|8|13|de filiis Adonicam qui erant novissimi et haec nomina eorum Helifeleth et Heihel et Samaias et cum eis sexaginta viri
EZRA|8|14|de filiis Beggui Uthai et Zacchur et cum eo septuaginta viri
EZRA|8|15|congregavi autem eos ad fluvium qui decurrit ad Ahavva et mansimus ibi diebus tribus quaesivique in populo et in sacerdotibus de filiis Levi et non inveni ibi
EZRA|8|16|itaque misi Heliezer et Arihel et Semeam et Helnathan et Iarib et alterum Helnathan et Nathan et Zacchariam et Mesolam principes et Ioarib et Helnathan sapientes
EZRA|8|17|et misi eos ad Heddo qui est primus in Casphiae loco et posui in ore eorum verba quae loquerentur ad Addom et ad fratres eius Nathinneos in loco Casphiae ut adducerent nobis ministros domus Dei nostri
EZRA|8|18|et adduxerunt nobis per manum Dei nostri bonam super nos virum doctissimum de filiis Moolli filii Levi filii Israhel et Sarabiam et filios eius et fratres eius decem et octo
EZRA|8|19|et Asabiam et cum eo Isaiam de filiis Merari fratres eius et filios eius viginti
EZRA|8|20|et de Nathinneis quos dederat David et principes ad ministeria Levitarum Nathinneos ducentos viginti omnes hii suis nominibus vocabantur
EZRA|8|21|et praedicavi ibi ieiunium iuxta fluvium Ahavva ut adfligeremur coram Domino Deo nostro et peteremus ab eo viam rectam nobis et filiis nostris universaeque substantiae nostrae
EZRA|8|22|erubui enim petere regem auxilium et equites qui defenderent nos ab inimico in via quia dixeramus regi manus Dei nostri est super omnes qui quaerunt eum in bonitate et imperium eius et fortitudo eius et furor super omnes qui derelinquunt eum
EZRA|8|23|ieiunavimus autem et rogavimus Deum nostrum pro hoc et evenit nobis prospere
EZRA|8|24|et separavi de principibus sacerdotum duodecim Sarabian Asabian et cum eis de fratribus eorum decem
EZRA|8|25|adpendique eis argentum et aurum et vasa consecrata domus Dei nostri quae obtulerat rex et consiliatores eius et principes eius universusque Israhel eorum qui inventi fuerant
EZRA|8|26|et adpendi in manibus eorum argenti talenta sescenta quinquaginta et vasa argentea centum auri centum talenta
EZRA|8|27|et crateras aureos viginti qui habebant solidos millenos et vasa aeris fulgentis optimi duo pulchra ut aurum
EZRA|8|28|et dixi eis vos sancti Domini et vasa sancta et argentum et aurum quod sponte oblatum est Domino Deo patrum vestrorum
EZRA|8|29|vigilate et custodite donec adpendatis coram principibus sacerdotum et Levitarum et ducibus familiarum Israhel in Hierusalem et thesaurum domus Domini
EZRA|8|30|susceperunt autem sacerdotes et Levitae pondus argenti et auri et vasorum ut deferrent in Hierusalem in domum Dei nostri
EZRA|8|31|promovimus ergo a flumine Ahavva duodecimo die mensis primi ut pergeremus Hierusalem et manus Dei nostri fuit super nos et liberavit nos de manu inimici et insidiatoris in via
EZRA|8|32|et venimus Hierusalem et mansimus ibi diebus tribus
EZRA|8|33|die autem quarta adpensum est argentum et aurum et vasa in domo Dei nostri per manum Meremoth filii Uriae sacerdotis et cum eo Eleazar filius Finees cumque eis Iozaded filius Iosue et Noadaia filius Bennoi Levitae
EZRA|8|34|iuxta numerum et pondus omnium descriptumque est omne pondus in tempore illo
EZRA|8|35|sed et qui venerant de captivitate filii transmigrationis obtulerunt holocaustomata Deo Israhel vitulos duodecim pro omni Israhel arietes nonaginta sex agnos septuaginta septem hircos pro peccato duodecim omnia in holocaustum Domino
EZRA|8|36|dederunt autem edicta regis satrapis qui erant de conspectu regis et ducibus trans Flumen et elevaverunt populum et domum Dei
EZRA|9|1|postquam autem haec conpleta sunt accesserunt ad me principes dicentes non est separatus populus Israhel et sacerdotes et Levitae a populis terrarum et de abominationibus eorum Chananei videlicet et Hetthei et Ferezei et Iebusei et Ammanitarum et Moabitarum et Aegyptiorum et Amorreorum
EZRA|9|2|tulerunt enim de filiabus eorum sibi et filiis suis et commiscuerunt semen sanctum cum populis terrarum manus etiam principum et magistratuum fuit in transgressione hac prima
EZRA|9|3|cumque audissem sermonem istum scidi pallium meum et tunicam et evelli capillos capitis mei et barbae et sedi maerens
EZRA|9|4|convenerunt autem ad me omnes qui timebant verbum Dei Israhel pro transgressione eorum qui de captivitate venerant et ego sedebam tristis usque ad sacrificium vespertinum
EZRA|9|5|et in sacrificio vespertino surrexi de adflictione mea et scisso pallio et tunica curvavi genua mea et expandi manus meas ad Dominum Deum meum
EZRA|9|6|et dixi Deus meus confundor et erubesco levare Deus meus faciem meam ad te quoniam iniquitates nostrae multiplicatae sunt super caput et delicta nostra creverunt usque in caelum
EZRA|9|7|a diebus patrum nostrorum sed et nos ipsi peccavimus granditer usque ad diem hanc et in iniquitatibus nostris traditi sumus ipsi et reges nostri et sacerdotes nostri in manum regum terrarum in gladium in captivitatem in rapinam et in confusionem vultus sicut et die hac
EZRA|9|8|et nunc quasi parum et ad momentum facta est deprecatio nostra apud Dominum Deum nostrum ut dimitterentur nobis reliquiae et daretur paxillus in loco sancto eius et inluminaret oculos nostros Deus noster et daret nobis vitam modicam in servitute nostra
EZRA|9|9|quia servi sumus et in servitute nostra non dereliquit nos Deus noster et inclinavit super nos misericordiam coram rege Persarum ut daret nobis vitam et sublimaret domum Dei nostri et extrueret solitudines eius et daret nobis sepem in Iuda et in Hierusalem
EZRA|9|10|et nunc quid dicemus Deus noster post haec quia dereliquimus mandata tua
EZRA|9|11|quae praecepisti in manu servorum tuorum prophetarum dicens terram ad quam vos ingredimini ut possideatis eam terra inmunda est iuxta inmunditiam populorum ceterarumque terrarum abominationibus eorum qui repleverunt eam ab ore usque ad os in coinquinatione sua
EZRA|9|12|nunc ergo filias vestras ne detis filiis eorum et filias eorum non accipiatis filiis vestris et non quaeratis pacem eorum et prosperitatem eorum usque in aeternum ut confortemini et comedatis quae bona sunt terrae et heredes habeatis filios vestros usque in saeculum
EZRA|9|13|et post omnia quae venerunt super nos in operibus nostris pessimis et in delicto nostro magno quia tu Deus noster liberasti nos de iniquitate nostra et dedisti nobis salutem sicut est hodie
EZRA|9|14|ut non converteremur et irrita faceremus mandata tua neque matrimonia iungeremus cum populis abominationum istarum numquid iratus es nobis usque ad consummationem ne dimitteres nobis reliquias et salutem
EZRA|9|15|Domine Deus Israhel iustus tu quoniam derelicti sumus qui salvaremur sicut die hac ecce coram te sumus in delicto nostro non enim stari potest coram te super hoc
EZRA|10|1|sic ergo orante Ezra et inplorante eo et flente et iacente ante templum Dei collectus est ad eum de Israhel coetus grandis nimis virorum et mulierum puerorumque et flevit populus multo fletu
EZRA|10|2|et respondit Sechenia filius Iehihel de filiis Helam et dixit Ezrae nos praevaricati sumus in Deum nostrum et duximus uxores alienigenas de populis terrae et nunc si est paenitentia Israhel super hoc
EZRA|10|3|percutiamus foedus cum Deo nostro ut proiciamus universas uxores et eos qui de his nati sunt iuxta voluntatem Domini et eorum qui timent praeceptum Dei nostri secundum legem fiat
EZRA|10|4|surge tuum est decernere nosque erimus tecum confortare et fac
EZRA|10|5|surrexit ergo Ezras et adiuravit principes sacerdotum Levitarum et omnem Israhel ut facerent secundum verbum hoc et iuraverunt
EZRA|10|6|et surrexit Ezras ante domum Dei et abiit ad cubiculum Iohanan filii Eliasib et ingressus est illuc panem non comedit et aquam non bibit lugebat enim in transgressione eorum qui de captivitate venerant
EZRA|10|7|et missa est vox in Iuda et in Hierusalem omnibus filiis transmigrationis ut congregarentur in Hierusalem
EZRA|10|8|et omnis qui non venerit in tribus diebus iuxta consilium principum et seniorum auferetur universa substantia eius et ipse abicietur de coetu transmigrationis
EZRA|10|9|convenerunt igitur omnes viri Iuda et Beniamin in Hierusalem tribus diebus ipse est mensis nonus vicesimo die mensis et sedit omnis populus in platea domus Dei trementes pro peccato et pluviis
EZRA|10|10|et surrexit Ezras sacerdos et dixit ad eos vos transgressi estis et duxistis uxores alienigenas ut adderetis super delictum Israhel
EZRA|10|11|et nunc date confessionem Domino Deo patrum vestrorum et facite placitum eius et separamini a populis terrae et ab uxoribus alienigenis
EZRA|10|12|et respondit universa multitudo dixitque voce magna iuxta verbum tuum ad nos sic fiat
EZRA|10|13|verumtamen quia populus multus est et tempus pluviae et non sustinemus stare foris et opus non est diei unius vel duorum vehementer quippe peccavimus in sermone isto
EZRA|10|14|constituantur principes in universa multitudine et omnes in civitatibus nostris qui duxerunt uxores alienigenas veniant in temporibus statutis et cum his seniores per civitatem et civitatem et iudices eius donec avertatur ira Dei nostri a nobis super peccato hoc
EZRA|10|15|igitur Ionathan filius Asahel et Iaazia filius Thecuae steterunt super hoc et Mesollam et Sebethai Levites adiuverunt eos
EZRA|10|16|feceruntque sic filii transmigrationis et abierunt Ezras sacerdos et viri principes familiarum in domum patrum suorum et omnes per nomina sua et sederunt in die primo mensis decimi ut quaererent rem
EZRA|10|17|et consummati sunt omnes viri qui duxerant uxores alienigenas usque ad diem primam mensis primi
EZRA|10|18|et inventi sunt de filiis sacerdotum qui duxerant uxores alienigenas de filiis Iosue filii Iosedech et fratres eius Maasia et Eliezer et Iarib et Godolia
EZRA|10|19|et dederunt manus suas ut eicerent uxores suas et pro delicto suo arietem de ovibus offerrent
EZRA|10|20|et de filiis Emmer Anani et Zebedia
EZRA|10|21|et de filiis Erim Masia et Helia et Semeia et Hiehihel et Ozias
EZRA|10|22|et de filiis Phessur Helioenai Maasia Ismahel Nathanahel Iozabeth et Elasa
EZRA|10|23|et de filiis Levitarum Iozabeth et Semei et Celaia ipse est Calita Phataia Iuda et Eliezer
EZRA|10|24|et de cantoribus Eliasub et de ianitoribus Sellum et Telem et Uri
EZRA|10|25|et ex Israhel de filiis Pharos Remia et Ezia et Melchia et Miamin et Eliezer et Melchia et Banea
EZRA|10|26|et de filiis Helam Mathania Zaccharias et Hiehil et Abdi et Irimoth et Helia
EZRA|10|27|et de filiis Zethua Helioenai Eliasib Mathania et Ierimuth et Zabeth et Aziza
EZRA|10|28|et de filiis Bebai Iohanan Anania Zabbai Athalai
EZRA|10|29|et de filiis Bani Mosollam et Melluch et Adaia Iasub et Saal et Ramoth
EZRA|10|30|et de filiis Phaethmoab Edna et Chalal Banaias Maasias Mathanias Beselehel et Bennui et Manasse
EZRA|10|31|et de filiis Erem Eliezer Iesue Melchias Semeias Symeon
EZRA|10|32|Beniamin Maloch Samarias
EZRA|10|33|de filiis Asom Matthanai Matthetha Zabed Elipheleth Iermai Manasse Semei
EZRA|10|34|de filiis Bani Maaddi Amram et Huhel
EZRA|10|35|Baneas et Badaias Cheiliau
EZRA|10|36|Vannia Marimuth et Eliasib
EZRA|10|37|Matthanias Mathanai et Iasi
EZRA|10|38|et Bani et Bennui Semei
EZRA|10|39|et Salmias et Nathan et Adaias
EZRA|10|40|Mechnedabai Sisai Sarai
EZRA|10|41|Ezrel et Selemau Semeria
EZRA|10|42|Sellum Amaria Ioseph
EZRA|10|43|de filiis Nebu Iaihel Matthathias Zabed Zabina Ieddu et Iohel Banaia
EZRA|10|44|omnes hii acceperunt uxores alienigenas et fuerunt ex eis mulieres quae pepererant filios
