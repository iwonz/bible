ESTH|1|1|這事發生在 亞哈隨魯 的時代， 亞哈隨魯 從 印度 直到 古實 統治一百二十七個省，
ESTH|1|2|就是 亞哈隨魯 王在 書珊 城堡中坐國度王位的那些日子。
ESTH|1|3|他在位第三年，為所有官員和臣僕擺設宴席，有 波斯 和 瑪代 的權貴，各省的貴族與領袖在他面前。
ESTH|1|4|他把他榮耀國度的豐富和他偉大威嚴的尊貴給他們看了許多日子，共一百八十天。
ESTH|1|5|這些日子滿了，王又為所有住 書珊 城堡的百姓，無論大小，在御花園的院子裏擺設宴席七日。
ESTH|1|6|院子裏有白色棉和藍色線，用細麻繩、紫色繩繫在白玉石柱的銀環上，又有金銀的床榻擺在紅、白、黃、黑大理石鑲嵌的地上。
ESTH|1|7|用金器皿盛酒，有很多不同的器皿，照王的厚意提供豐富的御酒。
ESTH|1|8|飲酒有規定，不准勉強人 ，因為王吩咐宮裏所有的臣宰，讓人各隨己意。
ESTH|1|9|瓦實提 王后在 亞哈隨魯 王的宮內也為婦女擺設宴席。
ESTH|1|10|第七日， 亞哈隨魯 王飲酒，心中快樂，就吩咐在他面前侍立的七個太監 米戶幔 、 比斯他 、 哈波拿 、 比革他 、 亞拔他 、 西達 、 甲迦 ，
ESTH|1|11|請 瓦實提 王后頭戴王后的冠冕到王面前，讓各民族和官員觀看她的美貌，因為她容貌美麗。
ESTH|1|12|瓦實提 王后卻不肯遵照太監所傳的王命前來，所以王非常憤怒，怒火中燒。
ESTH|1|13|按王的常規，辦事必先詢問知例明法的人。那時，王詢問通達時務的智慧人，
ESTH|1|14|就是在王左右常見王面、在國中坐高位的 波斯 和 瑪代 的七個大臣， 甲示拿 、 示達 、 押瑪他 、 他施斯 、 米力 、 瑪西拿 、 米慕干 ：
ESTH|1|15|「 瓦實提 王后不遵照太監所傳的王命，照例應當怎樣辦理呢？」
ESTH|1|16|米慕干 在王和眾官長面前回答說：「 瓦實提 王后這事，不但得罪王，並且有害於 亞哈隨魯 王各省的臣民。
ESTH|1|17|因為王后這事必傳到眾婦人那裏，她們就會藐視自己的丈夫，說：『 亞哈隨魯 王吩咐 瓦實提 王后到王面前，她卻不來。』
ESTH|1|18|今日 波斯 和 瑪代 的眾夫人聽見王后這事，必向王所有的官長照樣說，如此必造成無數的藐視和憤怒。
ESTH|1|19|王若以為好，請降諭旨，寫在 波斯 和 瑪代 人的條例中，永不更改，不准 瓦實提 再到 亞哈隨魯 王面前，把她王后的位分賜給比她更好的妃子。
ESTH|1|20|王的諭旨一傳遍全國，國土縱然遼闊，凡作妻子的，無論丈夫是尊貴或卑賤，都必尊敬他。」
ESTH|1|21|王和眾官長都以這話為美，王就照 米慕干 的建議去做。
ESTH|1|22|王下詔書，用各省的文字、各族的語言通知各省，使凡作丈夫的在家中作主，各說本地的語言 。
ESTH|2|1|這些事以後， 亞哈隨魯 王的憤怒平息，就想起 瓦實提 和她所做的，以及自己怎樣降旨辦她。
ESTH|2|2|於是王的侍臣對王說：「請派人為王尋找美貌的少女；
ESTH|2|3|請王派官員在國中各省招聚所有美貌的少女到 書珊 城堡的女院，交給王所派掌管女子的太監 希該 ，給她們香膏塗抹。
ESTH|2|4|王眼中看為好的女子可以立為王后，代替 瓦實提 。」王以這話為美，就照樣做。
ESTH|2|5|書珊 城堡中有一個 猶太 人名叫 末底改 ，是 便雅憫 人 基士 的曾孫， 示每 的孫子， 睚珥 的兒子。
ESTH|2|6|從前 巴比倫 王 尼布甲尼撒 把 猶大 王 耶哥尼雅 和百姓從 耶路撒冷 擄來， 末底改 也在被擄的人當中。
ESTH|2|7|末底改 撫養他叔叔的女兒 哈大沙 ，就是 以斯帖 ，因為她沒有父母。這女子容貌美麗；她父母死了， 末底改 收她為自己的女兒。
ESTH|2|8|王的諭旨和敕令傳出之後，許多女子被招聚到 書珊 城堡，交給掌管女子的 希該 ； 以斯帖 也被送入王宮，交給 希該 。
ESTH|2|9|希該 眼中寵愛 以斯帖 ，就恩待她，急忙給她塗抹的香膏和當得的份，又從王宮裏挑選七個宮女來服事她，使她和她的宮女搬入女院上好的房屋。
ESTH|2|10|以斯帖 未曾將自己的籍貫宗族告訴人，因為 末底改 囑咐她不可叫人知道。
ESTH|2|11|末底改 天天在女院前徘徊，要知道 以斯帖 是否平安，過得如何。
ESTH|2|12|眾女子照例先塗抹身體十二個月：六個月用沒藥油，六個月用香料和塗抹的香膏。滿了日期，每個女子挨次進去朝見 亞哈隨魯 王。
ESTH|2|13|女子進去朝見王是這樣：從女院到王宮的時候，凡她所要的都必給她帶進去。
ESTH|2|14|晚上她進去，次日回到另一個女院，交給掌管妃嬪的太監 沙甲 。除非王喜愛她，再提名召她，她就不再進去見王。
ESTH|2|15|末底改 的叔叔 亞比孩 的女兒，就是 末底改 收為自己女兒的 以斯帖 ，按次序要進去朝見王的時候，除了掌管女子的太監 希該 所分派給她的，她別無所求。凡看見 以斯帖 的都喜歡她。
ESTH|2|16|亞哈隨魯 王第七年十月，就是提別月， 以斯帖 被引入宮中朝見王。
ESTH|2|17|王愛 以斯帖 過於眾女子，她在王面前蒙寵愛勝過眾少女。王把王后的冠冕戴在她頭上，立她為王后，代替 瓦實提 。
ESTH|2|18|王為所有的官長和臣僕擺設大宴席，稱為 以斯帖 的宴席，又豁免各省的租稅，並照王的厚意大頒賞賜。
ESTH|2|19|第二次招聚少女的時候， 末底改 坐在朝門。
ESTH|2|20|以斯帖 遵照 末底改 所囑咐的，沒有將籍貫宗族告訴人； 以斯帖 照 末底改 的吩咐去做，正如受他撫養的時候一樣。
ESTH|2|21|那時候， 末底改 坐在朝門，王有兩個守門的太監， 辟探 和 提列 ，惱恨 亞哈隨魯 王，想要下手害他。
ESTH|2|22|末底改 知道了這件事，就告訴 以斯帖 王后。 以斯帖 以 末底改 的名向王報告。
ESTH|2|23|這事經過查究後發現是真的，二人就被掛在木頭上。這事在王面前記錄在史籍上。
ESTH|3|1|這些事以後， 亞哈隨魯 王使 亞甲 人 哈米大他 的兒子 哈曼 尊大，提升了他，叫他的爵位超過所有與他同朝的官長。
ESTH|3|2|在朝門，王所有的臣僕都跪拜 哈曼 ，因為王如此吩咐，但 末底改 不跪不拜。
ESTH|3|3|在朝門，王的臣僕對 末底改 說：「你為何違背王的命令呢？」
ESTH|3|4|他們天天勸他，他還是不聽，他們就告訴 哈曼 ，要看 末底改 的事是否站得住，因他已經告訴他們自己是 猶太 人。
ESTH|3|5|哈曼 見 末底改 不跪不拜，就非常憤怒。
ESTH|3|6|有人把 末底改 的宗族告訴 哈曼 。 哈曼 看下手只害 末底改 一人是小事，還圖謀要滅絕 亞哈隨魯 王全國所有的 猶太 人，就是 末底改 的宗族。
ESTH|3|7|亞哈隨魯 王十二年正月，就是尼散月，人在 哈曼 面前抽普珥，普珥即籤，要定何月何日；抽到了十二月，就是亞達月。
ESTH|3|8|哈曼 對 亞哈隨魯 王說：「有一民族散居在王國各省的民族中，與眾不同；他們的律例與萬民的律例不同，也不守王的律例，所以容留他們對王無益。
ESTH|3|9|王若以為好，請下諭旨滅絕他們，我就捐一萬他連得銀子交給管財政的人，納入王的府庫。」
ESTH|3|10|於是王從自己手上摘下戒指給 猶太 人的仇敵， 亞甲 人 哈米大他 的兒子 哈曼 。
ESTH|3|11|王對 哈曼 說：「這銀子賜給你，這民族也交給你，可以照你眼中看為好的待他們。」
ESTH|3|12|正月十三日，王的一些書記受召而來，照著 哈曼 一切所吩咐的，用各省的文字、各族的語言，奉 亞哈隨魯 王的名寫諭旨，又用王的戒指蓋印，傳給王的總督、各省的省長，以及各族的領袖。
ESTH|3|13|詔書由信差傳到王的各省，限令一日之內，就是在十二月，亞達月十三日，把所有的 猶太 人，無論老少婦女孩子，全然剪除，殺戮滅絕，並搶奪他們的財產。
ESTH|3|14|這諭旨的抄本以敕令的方式在各省頒佈，通知各族，預備等候那日。
ESTH|3|15|信差奉王的命令急忙起行，敕令傳遍了 書珊 城堡。王同 哈曼 坐下飲酒， 書珊 城堡卻陷入慌亂中。
ESTH|4|1|末底改 知道所發生的這一切事，就撕裂衣服，披麻蒙灰，在城中行走，痛哭哀號。
ESTH|4|2|他到了朝門前就停住腳步，因為穿麻衣的不可進朝門。
ESTH|4|3|王的諭旨和敕令所到的各省各處， 猶太 人都極其悲哀，禁食哭泣哀號，許多人躺在麻布和爐灰中。
ESTH|4|4|以斯帖 王后的宮女和太監來把這事告訴 以斯帖 ，她非常憂愁，就送衣服給 末底改 穿，要他脫下身上的麻衣，他卻不肯接受。
ESTH|4|5|以斯帖 把王所派伺候她的一個太監 哈他革 召來，吩咐他去見 末底改 ，要知道到底發生了甚麼事，為何如此。
ESTH|4|6|於是 哈他革 出來，到朝門前的廣場見 末底改 。
ESTH|4|7|末底改 把自己遭遇的一切，以及 哈曼 為滅絕 猶太 人答應捐入王庫的銀數都告訴了他；
ESTH|4|8|又把那傳遍 書珊 、要滅絕 猶太 人的諭旨抄本交給 哈他革 ，要他給 以斯帖 看，並向她說明，囑咐她去晉見王，向王懇求，為本族的人在王面前請命。
ESTH|4|9|哈他革 回來，把 末底改 的話告訴 以斯帖 。
ESTH|4|10|以斯帖 吩咐 哈他革 去見 末底改 ，說：
ESTH|4|11|「王所有的臣僕和各省的百姓都知道有一個定例，若未奉召見，擅入內院見王的，無論男女必被處死；除非王向他伸出金杖，不得存活。但我沒有被召進去見王已經有三十天了。」
ESTH|4|12|他們把 以斯帖 的話告訴 末底改 。
ESTH|4|13|末底改 託人回覆 以斯帖 說：「你不要自己以為在王宮裏強過任何 猶太 人，得以倖免。
ESTH|4|14|此時你若閉口不言， 猶太 人必從別處得解脫，蒙拯救；你和你父家必致滅亡。焉知你得了王后的位分不是為現今的機會嗎？」
ESTH|4|15|以斯帖 吩咐人回覆 末底改 說：
ESTH|4|16|「你當去召集 書珊 所有的 猶太 人，為我禁食三晝三夜，不吃不喝；我和我的宮女也要這樣禁食。然後我違例去晉見王，我若死就死吧！」
ESTH|4|17|於是 末底改 照 以斯帖 一切所吩咐的去做。
ESTH|5|1|第三日， 以斯帖 穿上朝服，站立在王宮的內院，對著王宮。王在殿裏坐在寶座上，對著殿的門。
ESTH|5|2|王見 以斯帖 王后站在院內，她在王的眼中得恩寵，王向她伸出手中的金杖。 以斯帖 往前去摸杖頭。
ESTH|5|3|王對她說：「 以斯帖 王后啊，你要甚麼？無論你求甚麼，就是國的一半也必賜給你。」
ESTH|5|4|以斯帖 說：「王若以為好，請王帶著 哈曼 今日赴我為王預備的宴席。」
ESTH|5|5|王說：「叫 哈曼 速速照 以斯帖 的話去做。」於是王帶著 哈曼 赴 以斯帖 所預備的宴席。
ESTH|5|6|在宴席喝酒的時候，王又對 以斯帖 說：「你要甚麼，必賜給你；無論你求甚麼，就是國的一半也必給你。」
ESTH|5|7|以斯帖 回答說：「我所要的、我所求的，嗯......。
ESTH|5|8|我若在王眼前蒙恩，王若願意賜我所要的，准我所求的，就請王和 哈曼 再赴我為你們預備的宴席。明日我必照王的話去做。」
ESTH|5|9|那日 哈曼 心中快樂，歡歡喜喜地出來。但是當他看見 末底改 在朝門不站起來，也不因他動一下，就滿心惱怒 末底改 。
ESTH|5|10|哈曼 忍著氣回家，叫人請他的一些朋友和他妻子 細利斯 來。
ESTH|5|11|哈曼 將他的榮華富貴、眾多的兒女，和王使他尊大、提升他高過官長和臣僕的事，都述說給他們聽。
ESTH|5|12|哈曼 又說：「 以斯帖 王后預備宴席，除了我之外不許別人隨王赴席。明日王后又請我隨王赴席。
ESTH|5|13|只是每當我看見 猶太 人 末底改 坐在朝門，這一切對我就都毫無意義了。」
ESTH|5|14|他的妻子 細利斯 和他所有的朋友對他說：「叫人做一個五十肘高的木架，早晨求王把 末底改 掛在其上，然後你可以歡歡喜喜隨王赴席。」 哈曼 認為這話很好，就叫人做了木架。
ESTH|6|1|那夜王睡不著覺，吩咐人取歷史書，就是史籍，念給他聽，
ESTH|6|2|發現書上寫著：王有兩個守門的太監 辟探 和 提列 ，想要下手害 亞哈隨魯 王， 末底改 告發了這件事。
ESTH|6|3|王說：「 末底改 做了這事，有沒有賜給他甚麼尊榮或高位呢？」伺候王的臣僕說：「沒有賜給他甚麼。」
ESTH|6|4|王說：「誰在院子裏？」那時 哈曼 正進入王宮的外院，要請王把 末底改 掛在他所預備的木架上。
ESTH|6|5|王的臣僕對他說：「看哪， 哈曼 站在院子裏。」王說：「叫他進來。」
ESTH|6|6|哈曼 就進去。王對他說：「王所喜愛要賜尊榮的人，當如何待他呢？」 哈曼 心裏說：「王所喜愛要賜尊榮的人，除了我，還有誰呢？」
ESTH|6|7|哈曼 就對王說：「王所喜愛要賜尊榮的人，
ESTH|6|8|當把王所穿的王袍拿來，牽了戴冠的御馬，
ESTH|6|9|把王袍和御馬都交給王一個極尊貴的大臣，吩咐人把王袍給王所喜愛要賜尊榮的人穿上，領他騎著御馬走遍城裏的廣場，在他面前宣告：『王所喜愛要賜尊榮的人，就是這樣待他。』」
ESTH|6|10|王對 哈曼 說：「你速速把這王袍和御馬，照你所說的，向坐在朝門的 猶太 人 末底改 去做。凡你所說的，一樣都不可缺。」
ESTH|6|11|於是 哈曼 把王袍給 末底改 穿上，領他騎著御馬走遍城裏的廣場，在他面前宣告：「王所喜愛要賜尊榮的人，就是這樣待他。」
ESTH|6|12|末底改 仍回到朝門， 哈曼 卻憂憂悶悶地蒙著頭，急忙回家去了。
ESTH|6|13|哈曼 把所遭遇的一切都說給他妻子 細利斯 和他所有的朋友聽。他的智囊團和他的妻子 細利斯 對他說：「你在 末底改 面前開始敗落；他既是 猶太 人，你必不能勝過他，終必在他面前敗落。」
ESTH|6|14|他們正跟 哈曼 說話的時候，王的幾位太監來了，催 哈曼 快去赴 以斯帖 所預備的宴席。
ESTH|7|1|王帶著 哈曼 來赴 以斯帖 王后的宴席。
ESTH|7|2|第二天在宴席喝酒的時候，王又對 以斯帖 說：「 以斯帖 王后啊，你要甚麼，必賜給你；無論你求甚麼，就是國的一半也必給你。」
ESTH|7|3|以斯帖 王后回答說：「王啊，我若在你眼前蒙恩，王若以為好，我所要的，是王把我的性命賜給我；我所求的，是求我的本族。
ESTH|7|4|因為我和我的本族被出賣了，要被剪除，殺戮，滅絕。我們若被賣為奴為婢，我就閉口不言；但我們的痛苦比起王的損失，算不得甚麼 。」
ESTH|7|5|亞哈隨魯 王問 以斯帖 王后說：「擅敢起意如此行的是誰？這人在哪裏呢？」
ESTH|7|6|以斯帖 說：「仇人敵人就是這惡人 哈曼 ！」 哈曼 在王和王后面前非常驚惶。
ESTH|7|7|王大怒，起來離開酒席往御花園去了。 哈曼 見王定意要加罪於他，就留下來求 以斯帖 王后救他的命。
ESTH|7|8|王從御花園回到酒席廳，見 哈曼 伏在 以斯帖 所靠的榻上；王說：「他竟敢在宮內、在我面前凌辱王后嗎？」這話一出王口， 哈曼 的臉就被蒙住了。
ESTH|7|9|有一個伺候王名叫 哈波拿 的太監說：「看哪， 哈曼 還為那報告給王、救王有功的 末底改 做了一個五十肘高的木架，現今立在 哈曼 的家裏。」王說：「把 哈曼 掛在木架上。」
ESTH|7|10|於是 哈曼 被掛在他為 末底改 所預備的木架上；王的憤怒才平息了。
ESTH|8|1|那日， 亞哈隨魯 王把 猶太 人的仇敵 哈曼 的家產賜給 以斯帖 王后。 末底改 也來到王面前，因為 以斯帖 已經告訴王， 末底改 跟她是甚麼關係。
ESTH|8|2|王摘下自己的戒指，就是從 哈曼 取回的，給了 末底改 。 以斯帖 派 末底改 管理 哈曼 的家產。
ESTH|8|3|以斯帖 又在王面前求情，俯伏在他腳前，流淚哀求他阻止 亞甲 人 哈曼 害 猶太 人的惡謀。
ESTH|8|4|王向 以斯帖 伸出金杖， 以斯帖 就起來，站在王面前，
ESTH|8|5|說：「王若以為好，我若在王面前蒙恩，王若認為合宜，我若在王眼前得喜悅，請王下諭旨，廢除 亞甲 人 哈米大他 的兒子 哈曼 設謀，要殺滅王各省的 猶太 人所頒的詔書。
ESTH|8|6|我何忍見我本族的人受害？何忍見我同宗的人被滅呢？」
ESTH|8|7|亞哈隨魯 王對 以斯帖 王后和 猶太 人 末底改 說：「因為 哈曼 要下手害 猶太 人，看哪，我已把他的家產賜給 以斯帖 ，也把 哈曼 掛在木架上了。
ESTH|8|8|你們可以照你們看為好的，奉王的名寫諭旨給 猶太 人，用王的戒指蓋印；因為奉王的名所寫、用王的戒指蓋印的諭旨是不能廢除的。」
ESTH|8|9|三月，就是西彎月二十三日，當時王的一些書記受召而來，按著 末底改 所吩咐的，用各省的文字、各族的語言，以及 猶太 人的文字語言寫諭旨，傳給那從 印度 直到 古實 一百二十七省的 猶太 人，以及總督、省長和領袖。
ESTH|8|10|末底改 奉 亞哈隨魯 王的名寫諭旨，用王的戒指蓋印，交給信差們騎上御用的王室快馬去頒佈。
ESTH|8|11|王准各城各鎮的 猶太 人在一日之內，在十二月，就是亞達月的十三日聚集，在 亞哈隨魯 王的各省保護自己的性命，剪除，殺戮，滅絕那要攻擊 猶太 人的各省各族所有的軍隊，以及他們的妻子兒女，奪取他們的財產為掠物。
ESTH|8|12|
ESTH|8|13|這諭旨的抄本以敕令的方式在各省頒佈，通知各族，使 猶太 人預備等候那日，好在仇敵身上報仇。
ESTH|8|14|於是騎御用快馬的信差奉王命催促，急忙起行；敕令傳遍了 書珊 城堡。
ESTH|8|15|末底改 穿著藍色白色的朝服，頭戴大金冠冕，又穿紫色細麻布的外袍，從王面前出來； 書珊城 充滿了歡樂的呼聲。
ESTH|8|16|猶太 人有光榮，歡喜快樂，得享尊貴。
ESTH|8|17|王的諭旨和敕令所到的各省各城， 猶太 人都歡喜快樂，擺設宴席，以那日為吉日。國中許多民族的人因懼怕 猶太 人，就自稱為 猶太 人。
ESTH|9|1|十二月，就是亞達月十三日，王的諭旨和敕令要執行的那一日， 猶太 人的仇敵盼望制伏他們，但 猶太 人反倒制伏了恨他們的人。
ESTH|9|2|猶太 人在 亞哈隨魯 王各省的城裏聚集，下手擊殺那些要害他們的人。沒有人能在他們面前站立得住，因為各民族都懼怕他們。
ESTH|9|3|各省的領袖、總督、省長，和辦理王事務的人，因懼怕 末底改 ，就都幫助 猶太 人。
ESTH|9|4|末底改 在朝中為大，名聲傳遍各省； 末底改 這人的權勢日漸擴大。
ESTH|9|5|猶太 人用刀擊殺所有的仇敵，殺滅他們，隨意待那些恨他們的人。
ESTH|9|6|在 書珊 城堡中， 猶太 人殺滅了五百人。
ESTH|9|7|他們殺了 巴珊大他 、 達分 、 亞斯帕他 、
ESTH|9|8|破拉他 、 亞大利雅 、 亞利大他 、
ESTH|9|9|帕瑪斯他 、 亞利賽 、 亞利代 、 瓦耶撒他 ；
ESTH|9|10|這十人都是 哈米大他 的孫子， 猶太 人的仇敵 哈曼 的兒子。 猶太 人卻沒有下手奪取財物。
ESTH|9|11|那日， 書珊 城堡中被殺的人數呈報到王面前。
ESTH|9|12|王對 以斯帖 王后說：「 猶太 人在 書珊 城堡中殺滅了五百人，又殺了 哈曼 的十個兒子，在王其餘的各省不知如何。你要甚麼，必賜給你；你還求甚麼，也必為你成就。」
ESTH|9|13|以斯帖 說：「王若以為好，求你允准 書珊 的 猶太 人，明日也照今日的諭旨去做，並把 哈曼 十個兒子的屍體掛在木架上。」
ESTH|9|14|王允准這麼做。敕令傳遍 書珊 ， 哈曼 十個兒子的屍體被掛了起來。
ESTH|9|15|亞達月十四日，在 書珊 的 猶太 人又聚集，在 書珊 殺了三百人，卻沒有下手奪取財物。
ESTH|9|16|亞達月十三日，在王各省其餘的 猶太 人也都聚集，保護自己的性命，擺脫仇敵得享平安。他們殺了七萬五千個恨他們的人，卻沒有下手奪取財物；十四日他們休息，以這日為設宴歡樂的日子。
ESTH|9|17|
ESTH|9|18|但 書珊 的 猶太 人卻在十三日、十四日聚集；十五日休息，以這日為設宴歡樂的日子。
ESTH|9|19|所以住在無城牆的鄉村的 猶太 人，都以亞達月十四日為設宴歡樂的吉日，彼此餽送禮物。
ESTH|9|20|末底改 記錄這些事，寫信給 亞哈隨魯 王各省遠近所有的 猶太 人，
ESTH|9|21|吩咐他們每年守亞達月十四、十五兩日，
ESTH|9|22|以這兩日為 猶太 人擺脫仇敵得享平安、轉憂為喜、轉悲為樂的吉日，並在這兩日設宴歡樂，彼此餽送禮物，賙濟窮人。
ESTH|9|23|於是， 猶太 人照 末底改 所寫給他們的，把開始所做的作為遵守的定例。
ESTH|9|24|因為 猶太 人的仇敵 亞甲 人 哈米大他 的兒子 哈曼 設謀要殺害 猶太 人，抽普珥，普珥即籤，為要殺盡滅絕他們；
ESTH|9|25|但這陰謀 到了王面前，王卻降旨使 哈曼 謀害 猶太 人的惡事歸到他自己的頭上，他和他的眾子都被掛在木架上。
ESTH|9|26|所以 猶太 人照著普珥這名字稱這兩日為普珥日。他們因這信上一切的話，又因所看見所遇見的事，
ESTH|9|27|就規定自己與後裔，以及歸化他們的人，每年按所寫的、按時守這兩日，永久不廢。
ESTH|9|28|各省各城、世世代代、家家戶戶都記念並守這兩日，使這普珥日在 猶太 人中不可廢掉，在他們後裔中也永不遺忘。
ESTH|9|29|亞比孩 的女兒 以斯帖 王后和 猶太 人 末底改 以全權寫第二封信，堅立這普珥日，
ESTH|9|30|送信給 亞哈隨魯 王國中一百二十七省所有的 猶太 人，祝他們平安和安穩，
ESTH|9|31|勸他們遵照 猶太 人 末底改 和 以斯帖 王后所規定的，按時守這普珥日，並照著 猶太 人為自己與後裔所規定的，禁食與哀求。
ESTH|9|32|以斯帖 規定了守普珥日的條例，這事也記錄在書上。
ESTH|10|1|亞哈隨魯 王向國中和海島的人徵稅。
ESTH|10|2|他以權柄能力所做的一切，以及他使 末底改 尊大、提升他的事，豈不都寫在 瑪代 和 波斯 王的史籍上嗎？
ESTH|10|3|猶太 人 末底改 作 亞哈隨魯 王的宰相，在 猶太 人中為大，得許多弟兄的喜悅，為本族的人爭取福利，為他所有的後代謀求幸福。
