1THESS|1|1|Paul, Silas and Timothy, To the church of the Thessalonians in God the Father and the Lord Jesus Christ: Grace and peace to you.
1THESS|1|2|We always thank God for all of you, mentioning you in our prayers.
1THESS|1|3|We continually remember before our God and Father your work produced by faith, your labor prompted by love, and your endurance inspired by hope in our Lord Jesus Christ.
1THESS|1|4|For we know, brothers loved by God, that he has chosen you,
1THESS|1|5|because our gospel came to you not simply with words, but also with power, with the Holy Spirit and with deep conviction. You know how we lived among you for your sake.
1THESS|1|6|You became imitators of us and of the Lord; in spite of severe suffering, you welcomed the message with the joy given by the Holy Spirit.
1THESS|1|7|And so you became a model to all the believers in Macedonia and Achaia.
1THESS|1|8|The Lord's message rang out from you not only in Macedonia and Achaia--your faith in God has become known everywhere. Therefore we do not need to say anything about it,
1THESS|1|9|for they themselves report what kind of reception you gave us. They tell how you turned to God from idols to serve the living and true God,
1THESS|1|10|and to wait for his Son from heaven, whom he raised from the dead--Jesus, who rescues us from the coming wrath.
1THESS|2|1|You know, brothers, that our visit to you was not a failure.
1THESS|2|2|We had previously suffered and been insulted in Philippi, as you know, but with the help of our God we dared to tell you his gospel in spite of strong opposition.
1THESS|2|3|For the appeal we make does not spring from error or impure motives, nor are we trying to trick you.
1THESS|2|4|On the contrary, we speak as men approved by God to be entrusted with the gospel. We are not trying to please men but God, who tests our hearts.
1THESS|2|5|You know we never used flattery, nor did we put on a mask to cover up greed--God is our witness.
1THESS|2|6|We were not looking for praise from men, not from you or anyone else.
1THESS|2|7|As apostles of Christ we could have been a burden to you, but we were gentle among you, like a mother caring for her little children.
1THESS|2|8|We loved you so much that we were delighted to share with you not only the gospel of God but our lives as well, because you had become so dear to us.
1THESS|2|9|Surely you remember, brothers, our toil and hardship; we worked night and day in order not to be a burden to anyone while we preached the gospel of God to you.
1THESS|2|10|You are witnesses, and so is God, of how holy, righteous and blameless we were among you who believed.
1THESS|2|11|For you know that we dealt with each of you as a father deals with his own children,
1THESS|2|12|encouraging, comforting and urging you to live lives worthy of God, who calls you into his kingdom and glory.
1THESS|2|13|And we also thank God continually because, when you received the word of God, which you heard from us, you accepted it not as the word of men, but as it actually is, the word of God, which is at work in you who believe.
1THESS|2|14|For you, brothers, became imitators of God's churches in Judea, which are in Christ Jesus: You suffered from your own countrymen the same things those churches suffered from the Jews,
1THESS|2|15|who killed the Lord Jesus and the prophets and also drove us out. They displease God and are hostile to all men
1THESS|2|16|in their effort to keep us from speaking to the Gentiles so that they may be saved. In this way they always heap up their sins to the limit. The wrath of God has come upon them at last.
1THESS|2|17|But, brothers, when we were torn away from you for a short time (in person, not in thought), out of our intense longing we made every effort to see you.
1THESS|2|18|For we wanted to come to you--certainly I, Paul, did, again and again--but Satan stopped us.
1THESS|2|19|For what is our hope, our joy, or the crown in which we will glory in the presence of our Lord Jesus when he comes? Is it not you?
1THESS|2|20|Indeed, you are our glory and joy.
1THESS|3|1|So when we could stand it no longer, we thought it best to be left by ourselves in Athens.
1THESS|3|2|We sent Timothy, who is our brother and God's fellow worker in spreading the gospel of Christ, to strengthen and encourage you in your faith,
1THESS|3|3|so that no one would be unsettled by these trials. You know quite well that we were destined for them.
1THESS|3|4|In fact, when we were with you, we kept telling you that we would be persecuted. And it turned out that way, as you well know.
1THESS|3|5|For this reason, when I could stand it no longer, I sent Timothy to find out about your faith. I was afraid that in some way the tempter might have tempted you and our efforts might have been useless.
1THESS|3|6|But Timothy has just now come to us from you and has brought good news about your faith and love. He has told us that you always have pleasant memories of us and that you long to see us, just as we also long to see you.
1THESS|3|7|Therefore, brothers, in all our distress and persecution we were encouraged about you because of your faith.
1THESS|3|8|For now we really live, since you are standing firm in the Lord.
1THESS|3|9|How can we thank God enough for you in return for all the joy we have in the presence of our God because of you?
1THESS|3|10|Night and day we pray most earnestly that we may see you again and supply what is lacking in your faith.
1THESS|3|11|Now may our God and Father himself and our Lord Jesus clear the way for us to come to you.
1THESS|3|12|May the Lord make your love increase and overflow for each other and for everyone else, just as ours does for you.
1THESS|3|13|May he strengthen your hearts so that you will be blameless and holy in the presence of our God and Father when our Lord Jesus comes with all his holy ones.
1THESS|4|1|Finally, brothers, we instructed you how to live in order to please God, as in fact you are living. Now we ask you and urge you in the Lord Jesus to do this more and more.
1THESS|4|2|For you know what instructions we gave you by the authority of the Lord Jesus.
1THESS|4|3|It is God's will that you should be sanctified: that you should avoid sexual immorality;
1THESS|4|4|that each of you should learn to control his own body in a way that is holy and honorable,
1THESS|4|5|not in passionate lust like the heathen, who do not know God;
1THESS|4|6|and that in this matter no one should wrong his brother or take advantage of him. The Lord will punish men for all such sins, as we have already told you and warned you.
1THESS|4|7|For God did not call us to be impure, but to live a holy life.
1THESS|4|8|Therefore, he who rejects this instruction does not reject man but God, who gives you his Holy Spirit.
1THESS|4|9|Now about brotherly love we do not need to write to you, for you yourselves have been taught by God to love each other.
1THESS|4|10|And in fact, you do love all the brothers throughout Macedonia. Yet we urge you, brothers, to do so more and more.
1THESS|4|11|Make it your ambition to lead a quiet life, to mind your own business and to work with your hands, just as we told you,
1THESS|4|12|so that your daily life may win the respect of outsiders and so that you will not be dependent on anybody.
1THESS|4|13|Brothers, we do not want you to be ignorant about those who fall asleep, or to grieve like the rest of men, who have no hope.
1THESS|4|14|We believe that Jesus died and rose again and so we believe that God will bring with Jesus those who have fallen asleep in him.
1THESS|4|15|According to the Lord's own word, we tell you that we who are still alive, who are left till the coming of the Lord, will certainly not precede those who have fallen asleep.
1THESS|4|16|For the Lord himself will come down from heaven, with a loud command, with the voice of the archangel and with the trumpet call of God, and the dead in Christ will rise first.
1THESS|4|17|After that, we who are still alive and are left will be caught up together with them in the clouds to meet the Lord in the air. And so we will be with the Lord forever.
1THESS|4|18|Therefore encourage each other with these words.
1THESS|5|1|Now, brothers, about times and dates we do not need to write to you,
1THESS|5|2|for you know very well that the day of the Lord will come like a thief in the night.
1THESS|5|3|While people are saying, "Peace and safety," destruction will come on them suddenly, as labor pains on a pregnant woman, and they will not escape.
1THESS|5|4|But you, brothers, are not in darkness so that this day should surprise you like a thief.
1THESS|5|5|You are all sons of the light and sons of the day. We do not belong to the night or to the darkness.
1THESS|5|6|So then, let us not be like others, who are asleep, but let us be alert and self-controlled.
1THESS|5|7|For those who sleep, sleep at night, and those who get drunk, get drunk at night.
1THESS|5|8|But since we belong to the day, let us be self-controlled, putting on faith and love as a breastplate, and the hope of salvation as a helmet.
1THESS|5|9|For God did not appoint us to suffer wrath but to receive salvation through our Lord Jesus Christ.
1THESS|5|10|He died for us so that, whether we are awake or asleep, we may live together with him.
1THESS|5|11|Therefore encourage one another and build each other up, just as in fact you are doing.
1THESS|5|12|Now we ask you, brothers, to respect those who work hard among you, who are over you in the Lord and who admonish you.
1THESS|5|13|Hold them in the highest regard in love because of their work. Live in peace with each other.
1THESS|5|14|And we urge you, brothers, warn those who are idle, encourage the timid, help the weak, be patient with everyone.
1THESS|5|15|Make sure that nobody pays back wrong for wrong, but always try to be kind to each other and to everyone else.
1THESS|5|16|Be joyful always;
1THESS|5|17|pray continually;
1THESS|5|18|give thanks in all circumstances, for this is God's will for you in Christ Jesus.
1THESS|5|19|Do not put out the Spirit's fire;
1THESS|5|20|do not treat prophecies with contempt.
1THESS|5|21|Test everything. Hold on to the good.
1THESS|5|22|Avoid every kind of evil.
1THESS|5|23|May God himself, the God of peace, sanctify you through and through. May your whole spirit, soul and body be kept blameless at the coming of our Lord Jesus Christ.
1THESS|5|24|The one who calls you is faithful and he will do it.
1THESS|5|25|Brothers, pray for us.
1THESS|5|26|Greet all the brothers with a holy kiss.
1THESS|5|27|I charge you before the Lord to have this letter read to all the brothers.
1THESS|5|28|The grace of our Lord Jesus Christ be with you.
