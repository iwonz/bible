JOEL|1|1|The word of the LORD that came to Joel son of Pethuel.
JOEL|1|2|Hear this, you elders; listen, all who live in the land. Has anything like this ever happened in your days or in the days of your forefathers?
JOEL|1|3|Tell it to your children, and let your children tell it to their children, and their children to the next generation.
JOEL|1|4|What the locust swarm has left the great locusts have eaten; what the great locusts have left the young locusts have eaten; what the young locusts have left other locusts have eaten.
JOEL|1|5|Wake up, you drunkards, and weep! Wail, all you drinkers of wine; wail because of the new wine, for it has been snatched from your lips.
JOEL|1|6|A nation has invaded my land, powerful and without number; it has the teeth of a lion, the fangs of a lioness.
JOEL|1|7|It has laid waste my vines and ruined my fig trees. It has stripped off their bark and thrown it away, leaving their branches white.
JOEL|1|8|Mourn like a virgin in sackcloth grieving for the husband of her youth.
JOEL|1|9|Grain offerings and drink offerings are cut off from the house of the LORD. The priests are in mourning, those who minister before the LORD.
JOEL|1|10|The fields are ruined, the ground is dried up; the grain is destroyed, the new wine is dried up, the oil fails.
JOEL|1|11|Despair, you farmers, wail, you vine growers; grieve for the wheat and the barley, because the harvest of the field is destroyed.
JOEL|1|12|The vine is dried up and the fig tree is withered; the pomegranate, the palm and the apple tree- all the trees of the field-are dried up. Surely the joy of mankind is withered away.
JOEL|1|13|Put on sackcloth, O priests, and mourn; wail, you who minister before the altar. Come, spend the night in sackcloth, you who minister before my God; for the grain offerings and drink offerings are withheld from the house of your God.
JOEL|1|14|Declare a holy fast; call a sacred assembly. Summon the elders and all who live in the land to the house of the LORD your God, and cry out to the LORD.
JOEL|1|15|Alas for that day! For the day of the LORD is near; it will come like destruction from the Almighty.
JOEL|1|16|Has not the food been cut off before our very eyes- joy and gladness from the house of our God?
JOEL|1|17|The seeds are shriveled beneath the clods. The storehouses are in ruins, the granaries have been broken down, for the grain has dried up.
JOEL|1|18|How the cattle moan! The herds mill about because they have no pasture; even the flocks of sheep are suffering.
JOEL|1|19|To you, O LORD, I call, for fire has devoured the open pastures and flames have burned up all the trees of the field.
JOEL|1|20|Even the wild animals pant for you; the streams of water have dried up and fire has devoured the open pastures.
JOEL|2|1|Blow the trumpet in Zion; sound the alarm on my holy hill. Let all who live in the land tremble, for the day of the LORD is coming. It is close at hand-
JOEL|2|2|a day of darkness and gloom, a day of clouds and blackness. Like dawn spreading across the mountains a large and mighty army comes, such as never was of old nor ever will be in ages to come.
JOEL|2|3|Before them fire devours, behind them a flame blazes. Before them the land is like the garden of Eden, behind them, a desert waste- nothing escapes them.
JOEL|2|4|They have the appearance of horses; they gallop along like cavalry.
JOEL|2|5|With a noise like that of chariots they leap over the mountaintops, like a crackling fire consuming stubble, like a mighty army drawn up for battle.
JOEL|2|6|At the sight of them, nations are in anguish; every face turns pale.
JOEL|2|7|They charge like warriors; they scale walls like soldiers. They all march in line, not swerving from their course.
JOEL|2|8|They do not jostle each other; each marches straight ahead. They plunge through defenses without breaking ranks.
JOEL|2|9|They rush upon the city; they run along the wall. They climb into the houses; like thieves they enter through the windows.
JOEL|2|10|Before them the earth shakes, the sky trembles, the sun and moon are darkened, and the stars no longer shine.
JOEL|2|11|The LORD thunders at the head of his army; his forces are beyond number, and mighty are those who obey his command. The day of the LORD is great; it is dreadful. Who can endure it?
JOEL|2|12|"Even now," declares the LORD, "return to me with all your heart, with fasting and weeping and mourning."
JOEL|2|13|Rend your heart and not your garments. Return to the LORD your God, for he is gracious and compassionate, slow to anger and abounding in love, and he relents from sending calamity.
JOEL|2|14|Who knows? He may turn and have pity and leave behind a blessing- grain offerings and drink offerings for the LORD your God.
JOEL|2|15|Blow the trumpet in Zion, declare a holy fast, call a sacred assembly.
JOEL|2|16|Gather the people, consecrate the assembly; bring together the elders, gather the children, those nursing at the breast. Let the bridegroom leave his room and the bride her chamber.
JOEL|2|17|Let the priests, who minister before the LORD, weep between the temple porch and the altar. Let them say, "Spare your people, O LORD. Do not make your inheritance an object of scorn, a byword among the nations. Why should they say among the peoples, 'Where is their God?'"
JOEL|2|18|Then the LORD will be jealous for his land and take pity on his people.
JOEL|2|19|The LORD will reply to them: "I am sending you grain, new wine and oil, enough to satisfy you fully; never again will I make you an object of scorn to the nations.
JOEL|2|20|"I will drive the northern army far from you, pushing it into a parched and barren land, with its front columns going into the eastern sea and those in the rear into the western sea. And its stench will go up; its smell will rise." Surely he has done great things.
JOEL|2|21|Be not afraid, O land; be glad and rejoice. Surely the LORD has done great things.
JOEL|2|22|Be not afraid, O wild animals, for the open pastures are becoming green. The trees are bearing their fruit; the fig tree and the vine yield their riches.
JOEL|2|23|Be glad, O people of Zion, rejoice in the LORD your God, for he has given you the autumn rains in righteousness. He sends you abundant showers, both autumn and spring rains, as before.
JOEL|2|24|The threshing floors will be filled with grain; the vats will overflow with new wine and oil.
JOEL|2|25|"I will repay you for the years the locusts have eaten- the great locust and the young locust, the other locusts and the locust swarm - my great army that I sent among you.
JOEL|2|26|You will have plenty to eat, until you are full, and you will praise the name of the LORD your God, who has worked wonders for you; never again will my people be shamed.
JOEL|2|27|Then you will know that I am in Israel, that I am the LORD your God, and that there is no other; never again will my people be shamed.
JOEL|2|28|"And afterward, I will pour out my Spirit on all people. Your sons and daughters will prophesy, your old men will dream dreams, your young men will see visions.
JOEL|2|29|Even on my servants, both men and women, I will pour out my Spirit in those days.
JOEL|2|30|I will show wonders in the heavens and on the earth, blood and fire and billows of smoke.
JOEL|2|31|The sun will be turned to darkness and the moon to blood before the coming of the great and dreadful day of the LORD.
JOEL|2|32|And everyone who calls on the name of the LORD will be saved; for on Mount Zion and in Jerusalem there will be deliverance, as the LORD has said, among the survivors whom the LORD calls.
JOEL|3|1|"In those days and at that time, when I restore the fortunes of Judah and Jerusalem,
JOEL|3|2|I will gather all nations and bring them down to the Valley of Jehoshaphat. There I will enter into judgment against them concerning my inheritance, my people Israel, for they scattered my people among the nations and divided up my land.
JOEL|3|3|They cast lots for my people and traded boys for prostitutes; they sold girls for wine that they might drink.
JOEL|3|4|"Now what have you against me, O Tyre and Sidon and all you regions of Philistia? Are you repaying me for something I have done? If you are paying me back, I will swiftly and speedily return on your own heads what you have done.
JOEL|3|5|For you took my silver and my gold and carried off my finest treasures to your temples.
JOEL|3|6|You sold the people of Judah and Jerusalem to the Greeks, that you might send them far from their homeland.
JOEL|3|7|"See, I am going to rouse them out of the places to which you sold them, and I will return on your own heads what you have done.
JOEL|3|8|I will sell your sons and daughters to the people of Judah, and they will sell them to the Sabeans, a nation far away." The LORD has spoken.
JOEL|3|9|Proclaim this among the nations: Prepare for war! Rouse the warriors! Let all the fighting men draw near and attack.
JOEL|3|10|Beat your plowshares into swords and your pruning hooks into spears. Let the weakling say, "I am strong!"
JOEL|3|11|Come quickly, all you nations from every side, and assemble there. Bring down your warriors, O LORD!
JOEL|3|12|"Let the nations be roused; let them advance into the Valley of Jehoshaphat, for there I will sit to judge all the nations on every side.
JOEL|3|13|Swing the sickle, for the harvest is ripe. Come, trample the grapes, for the winepress is full and the vats overflow- so great is their wickedness!"
JOEL|3|14|Multitudes, multitudes in the valley of decision! For the day of the LORD is near in the valley of decision.
JOEL|3|15|The sun and moon will be darkened, and the stars no longer shine.
JOEL|3|16|The LORD will roar from Zion and thunder from Jerusalem; the earth and the sky will tremble. But the LORD will be a refuge for his people, a stronghold for the people of Israel.
JOEL|3|17|"Then you will know that I, the LORD your God, dwell in Zion, my holy hill. Jerusalem will be holy; never again will foreigners invade her.
JOEL|3|18|"In that day the mountains will drip new wine, and the hills will flow with milk; all the ravines of Judah will run with water. A fountain will flow out of the LORD's house and will water the valley of acacias.
JOEL|3|19|But Egypt will be desolate, Edom a desert waste, because of violence done to the people of Judah, in whose land they shed innocent blood.
JOEL|3|20|Judah will be inhabited forever and Jerusalem through all generations.
JOEL|3|21|Their bloodguilt, which I have not pardoned, I will pardon." The LORD dwells in Zion!
