JONAH|1|1|І було слово Господнє до Йони, Аміттаєвого сина, таке:
JONAH|1|2|Устань, іди до Ніневії, великого міста, і проповідуй проти нього, бо їхнє зло прийшло перед лице Моє.
JONAH|1|3|І встав Йона, щоб утекти до Таршішу з-перед Господнього лиця. І зійшов він до Яфи, і знайшов корабля, що йшов до Таршішу, і дав заплату його, і ввійшов у нього, щоб відплисти з ними до Таршішу з-перед Господнього лиця.
JONAH|1|4|А Господь кинув сильного вітра на море, і знялася на морі велика буря, і вже думали, що корабель буде розбитий.
JONAH|1|5|І налякалися моряки, і кликали кожен до своїх богів, і викидали ті речі, що були на кораблі, до моря, щоб полегшити себе. А Йона зійшов до споду корабля, і ліг, і заснув.
JONAH|1|6|І приступив до нього керівник корабля, та й сказав йому: Чого ти спиш? Уставай, заклич до свого Бога, може згадає цей Бог про нас, і ми не згинемо.
JONAH|1|7|І сказали вони один до одного: Ідіть, і киньмо жеребки, та й пізнаємо, через кого нам оце лихо. І кинули вони жеребки, і впав жеребок на Йону.
JONAH|1|8|І сказали до нього: Об'яви ж нам, через що нам це лихо? Яке твоє зайняття, і звідки ти йдеш? Який твій край, і з якого ти народу?
JONAH|1|9|І сказав він до них: Я єврей, і боюся я Господа, Небесного Бога, що вчинив море та суходіл.
JONAH|1|10|І налякалися ті люди великим страхом, і сказали до нього: Що це ти наробив? Бо ці люди довідалися, що він утікає з-перед Господнього лиця, бо він це їм об'явив.
JONAH|1|11|І вони сказали до нього: Що ми зробимо тобі, щоб утихомирилось море, щоб не заливало нас? Бо море бушувало все більше.
JONAH|1|12|І сказав він до них: Візьміть мене, і киньте мене до моря, і втихомириться море перед вами; бо я знаю, що через мене оця велика буря на вас.
JONAH|1|13|І міцно гребли ці люди, щоб дістатися до суходолу, та не могли, бо море бушувало все більш проти них.
JONAH|1|14|І вони кликнули до Господа та й сказали: О Господи, нехай же не згинемо ми за душу цього чоловіка, і не давай на нас неповинної крови, бо Ти, Господи, чиниш, як бажаєш!
JONAH|1|15|І підняли вони Йону, і кинули його до моря, і спинилося море від своєї лютости.
JONAH|1|16|І налякалися ці люди Господа великим страхом, і приносили Господеві жертви, і складали обітниці.
JONAH|1|17|(2-1) І призначив Господь велику рибу, щоб вона проковтнула Йону. І був Йона в середині цієї риби три дні та три ночі.
JONAH|2|1|(2-2) І молився Йона до Господа, Бога свого, з утроби тієї риби,
JONAH|2|2|(2-3) та й казав: Я кликав з нещастя свого до Господа, і відповідь дав Він мені, із нутра шеолу кричав я, і почув Ти мій голос!
JONAH|2|3|(2-4) І Ти кинув мене в глибочінь, у серце моря, і потік оточив був мене. Усі хвилі Твої та буруни Твої надо мною пройшли.
JONAH|2|4|(2-5) І сказав я: Я вигнаний з-перед очей Твоїх, проте ще побачу я храм Твій святий.
JONAH|2|5|(2-6) Вода аж по душу мене обгорнула, безодня мене оточила, очерет обвиває кругом мою голову!
JONAH|2|6|(2-7) Я зійшов аж до споду гори, а земля її засуви стали за мною навіки! Та підіймеш із ями життя моє, Господи, Боже Ти мій!
JONAH|2|7|(2-8) Як у мені омлівала душа моя, Господа я спогадав, і молитва моя ця до Тебе долинула, до храму святого Твого!
JONAH|2|8|(2-9) Ті, що тримаються марних божків, свого Милосердного кидають.
JONAH|2|9|(2-10) А я голосною подякою принесу Тобі жертву, про що присягав я, те виконаю. Спасіння у Господа!
JONAH|2|10|(2-11) І Господь звелів рибі, і вона викинула Йону на суходіл.
JONAH|3|1|І було Господнє слово до Йони вдруге таке:
JONAH|3|2|Устань, іди до Ніневії, великого міста, і проповідуй на нього те слово, що Я говорив був тобі!
JONAH|3|3|І Йона встав, і пішов до Ніневії за Господнім словом. А Ніневія була місто велике-превелике, на три дні ходи.
JONAH|3|4|І зачав Йона ходити по місті, на один день ходи, і проповідував і казав: Ще сорок день, і Ніневія буде зруйнована!
JONAH|3|5|І ніневітяни ввірували в Бога, і оголосили піст, і позодягали верети, від найбільшого з них аж до найменшого.
JONAH|3|6|І дійшло це слово до царя Ніневії, і він устав зо свого трону, і скинув плаща свого з себе, і покрився веретою, та й сів на попелі.
JONAH|3|7|І він звелів кликнути й сказати в Ніневії з наказу царя та його вельмож, говорячи: Нехай не покуштують нічого ані людина, ані худоба, худоба велика чи худоба дрібна, нехай вони не пасуться, і нехай не п'ють води!
JONAH|3|8|І нехай покриваються веретами та людина й та худоба, і нехай сильно кличуть до Бога, і нехай кожен зверне з своєї дороги та від насильства, що в їхніх руках.
JONAH|3|9|Хто знає, може Бог обернеться й пожалує, і відвернеться з жару гніву Свого, і ми не погинемо!
JONAH|3|10|І побачив Бог їхні вчинки, що звернули зо своєї злої дороги, і пожалував Бог щодо того лиха, про яке говорив, що їм учинить, і не вчинив.
JONAH|4|1|І було це для Йони на досаду, досаду велику, і він запалився.
JONAH|4|2|І молився він до Господа та й казав: О Господи, чи ж не це моє слово, поки я ще був на своїй землі? Тому я перед тим утік до Таршішу, бо я знав, що Ти Бог милостивий та милосердий, довготерпеливий та многомилостивий, і Ти жалкуєш за зло.
JONAH|4|3|А тепер, Господи, візьми мою душу від мене, бо краще мені смерть від мого життя!
JONAH|4|4|А Господь відказав: Чи слушно ти запалився?
JONAH|4|5|І вийшов Йона з міста, і сів від сходу міста, і поставив собі там куреня, і сів під ним у тіні, аж поки побачить, що буде в місті.
JONAH|4|6|І виростив Бог рицинового куща, і він вигнався понад Йону, щоб бути тінню над його головою, щоб урятувати його від його досади. І втішився Йона від цього рицинового куща великою радістю.
JONAH|4|7|А при сході зірниці другого дня призначив Бог червяка, і він підточив рицинового куща, і той усох.
JONAH|4|8|І сталося, як сонце зійшло, то призначив Бог східнього гарячого вітра, і вдарило сонце на Йонину голову, і він зомлів. І він жадав, щоб йому померти, і казав: Краще мені смерть від мого життя!
JONAH|4|9|І промовив Бог до Йони: Чи слушно запалився ти за рициновий кущ? А той відказав: Дуже розлютився я, аж на смерть!
JONAH|4|10|І сказав Господь: Ти змилувався над рициновим кущем, над яким не трудився, і не плекав його, який виріс за одну ніч, і за одну ніч згинув.
JONAH|4|11|А Я не змилувався б над Ніневією, цим великим містом, що в ньому більше дванадцяти десятисячок люда, які не вміють розрізняти правиці своєї від своєї лівиці, та численна худоба?
