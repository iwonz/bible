EZRA|1|1|波斯 王 居鲁士 元年，耶和华为要应验藉 耶利米 的口所说的话，就激发 波斯 王 居鲁士 的心，使他下诏书通告全国，说：
EZRA|1|2|“ 波斯 王 居鲁士 如此说：耶和华天上的上帝已将地上万国赐给我，又委派我在 犹大 的 耶路撒冷 为他建造殿宇。
EZRA|1|3|你们中间凡作他子民的，可以上 犹大 的 耶路撒冷 去，重建耶和华－ 以色列 上帝的殿，他是在 耶路撒冷 的上帝；愿上帝与这人同在。
EZRA|1|4|凡存留的人，无论寄居何处，那地的人要用金银、财物、牲畜帮助他，还要为 耶路撒冷 上帝的殿甘心献上礼物。”
EZRA|1|5|于是， 犹大 和 便雅悯 的族长、祭司、 利未 人，凡是心被上帝感动的人都起来，要上 耶路撒冷 去建造耶和华的殿。
EZRA|1|6|四围所有的人都拿银器 、金子、财物、牲畜、珍宝支持他们 ，此外还有甘心献的一切礼物 。
EZRA|1|7|居鲁士 王也把耶和华殿的器皿拿出来，这些器皿是 尼布甲尼撒 从 耶路撒冷 掠取，放在自己神明庙中的。
EZRA|1|8|波斯 王 居鲁士 派 米提利达 司库把这些器皿拿出来，点交给 犹大 的领袖 设巴萨 。
EZRA|1|9|它们的数目如下：金盘三十个，银盘一千个，刀二十九把，
EZRA|1|10|金碗三十个，备用银碗四百一十个，其他器皿一千件。
EZRA|1|11|金银器皿共有五千四百件。被掳的人从 巴比伦 上 耶路撒冷 的时候， 设巴萨 把这一切都带了上来。
EZRA|2|1|这些是从被掳之地上来的省民， 巴比伦 王 尼布甲尼撒 把他们掳到 巴比伦 ，他们重返 耶路撒冷 和 犹大 ，各归本城。
EZRA|2|2|他们是同 所罗巴伯 、 耶书亚 、 尼希米 、 西莱雅 、 利来雅 、 末底改 、 必珊 、 米斯拔 、 比革瓦伊 、 利宏 、 巴拿 一起回来的。 以色列 百姓的人数如下：
EZRA|2|3|巴录 的子孙二千一百七十二名；
EZRA|2|4|示法提雅 的子孙三百七十二名；
EZRA|2|5|亚拉 的子孙七百七十五名；
EZRA|2|6|巴哈．摩押 的后裔，就是 耶书亚 和 约押 的子孙二千八百一十二名；
EZRA|2|7|以拦 的子孙一千二百五十四名；
EZRA|2|8|萨土 的子孙九百四十五名；
EZRA|2|9|萨改 的子孙七百六十名；
EZRA|2|10|巴尼 的子孙六百四十二名；
EZRA|2|11|比拜 的子孙六百二十三名；
EZRA|2|12|押甲 的子孙一千二百二十二名；
EZRA|2|13|亚多尼干 的子孙六百六十六名；
EZRA|2|14|比革瓦伊 的子孙二千零五十六名；
EZRA|2|15|亚丁 的子孙四百五十四名；
EZRA|2|16|亚特 的后裔，就是 希西家 的子孙九十八名；
EZRA|2|17|比赛 的子孙三百二十三名；
EZRA|2|18|约拉 的子孙一百一十二名；
EZRA|2|19|哈顺 的子孙二百二十三名；
EZRA|2|20|吉罢珥 人九十五名；
EZRA|2|21|伯利恒 人一百二十三名；
EZRA|2|22|尼陀法 人五十六名；
EZRA|2|23|亚拿突 人一百二十八名；
EZRA|2|24|亚斯玛弗 人四十二名；
EZRA|2|25|基列．耶琳 人、 基非拉 人、 比录 人共七百四十三名；
EZRA|2|26|拉玛 人和 迦巴 人共六百二十一名；
EZRA|2|27|默玛 人一百二十二名；
EZRA|2|28|伯特利 人和 艾 人共二百二十三名；
EZRA|2|29|尼波 人五十二名；
EZRA|2|30|末必 人一百五十六名；
EZRA|2|31|另一个 以拦 的子孙一千二百五十四名；
EZRA|2|32|哈琳 的子孙三百二十名；
EZRA|2|33|罗德 人、 哈第 人、 阿挪 人共七百二十五名；
EZRA|2|34|耶利哥 人三百四十五名；
EZRA|2|35|西拿 人三千六百三十名。
EZRA|2|36|祭司： 耶书亚 家 耶大雅 的子孙九百七十三名；
EZRA|2|37|音麦 的子孙一千零五十二名；
EZRA|2|38|巴施户珥 的子孙一千二百四十七名；
EZRA|2|39|哈琳 的子孙一千零一十七名。
EZRA|2|40|利未 人： 何达威雅 的后裔，就是 耶书亚 和 甲篾 的子孙七十四名。
EZRA|2|41|歌唱的： 亚萨 的子孙一百二十八名。
EZRA|2|42|门口的守卫： 沙龙 的子孙、 亚特 的子孙、 达们 的子孙、 亚谷 的子孙、 哈底大 的子孙、 朔拜 的子孙，共一百三十九名。
EZRA|2|43|殿役： 西哈 的子孙、 哈苏巴 的子孙、 答巴俄 的子孙、
EZRA|2|44|基绿 的子孙、 西亚 的子孙、 巴顿 的子孙、
EZRA|2|45|利巴拿 的子孙、 哈迦巴 的子孙、 亚谷 的子孙、
EZRA|2|46|哈甲 的子孙、 萨买 的子孙、 哈难 的子孙、
EZRA|2|47|吉德 的子孙、 迦哈 的子孙、 利亚雅 的子孙、
EZRA|2|48|利汛 的子孙、 尼哥大 的子孙、 迦散 的子孙、
EZRA|2|49|乌撒 的子孙、 巴西亚 的子孙、 比赛 的子孙、
EZRA|2|50|押拿 的子孙、 米乌宁 的子孙、 尼普心 的子孙、
EZRA|2|51|巴卜 的子孙、 哈古巴 的子孙、 哈忽 的子孙、
EZRA|2|52|巴洗律 的子孙、 米希大 的子孙、 哈沙 的子孙、
EZRA|2|53|巴柯 的子孙、 西西拉 的子孙、 答玛 的子孙、
EZRA|2|54|尼细亚 的子孙、 哈提法 的子孙。
EZRA|2|55|所罗门 仆人的后裔： 琐太 的子孙、 琐斐列 的子孙、 比路大 的子孙、
EZRA|2|56|雅拉 的子孙、 达昆 的子孙、 吉德 的子孙、
EZRA|2|57|示法提雅 的子孙、 哈替 的子孙、 玻黑列．哈斯巴音 的子孙、 亚米 的子孙。
EZRA|2|58|殿役和 所罗门 仆人的后裔共三百九十二名。
EZRA|2|59|从 特．米拉 、 特．哈萨 、 基绿 、 亚顿 、 音麦 上来，不能证明他们的父系家族和后裔是否属 以色列 的如下：
EZRA|2|60|第莱雅 的子孙、 多比雅 的子孙、 尼哥大 的子孙，共六百五十二名。
EZRA|2|61|祭司中， 哈巴雅 的子孙、 哈哥斯 的子孙、 巴西莱 的子孙， 巴西莱 因为娶了 基列 人 巴西莱 的女儿为妻，所以就以此为名。
EZRA|2|62|这些人在族谱之中寻查自己的谱系，却寻不着，因此算为不洁，不得作祭司。
EZRA|2|63|省长对他们说，不可吃至圣的物，直到有会用乌陵和土明的祭司兴起来。
EZRA|2|64|全会众共有四万二千三百六十名。
EZRA|2|65|此外，还有他们的仆婢七千三百三十七名，又有歌唱的男女二百名。
EZRA|2|66|他们有七百三十六匹马，二百四十五匹骡子，
EZRA|2|67|四百三十五匹骆驼，六千七百二十匹驴。
EZRA|2|68|有些族长到了 耶路撒冷 耶和华的殿，为上帝的殿甘心献上礼物，要在原有的根基上重新建造。
EZRA|2|69|他们量力捐入工程的库房，有六万一千达利克 金子，五千弥那银子，以及一百件祭司的礼服。
EZRA|2|70|于是祭司、 利未 人、百姓中的一些人、歌唱的、门口的守卫、殿役，各住在自己的城里； 以色列 众人都住在自己的城里。
EZRA|3|1|到了七月， 以色列 人住在自己的城里；那时他们如同一人，聚集在 耶路撒冷 。
EZRA|3|2|约萨达 的儿子 耶书亚 和他的弟兄众祭司，以及 撒拉铁 的儿子 所罗巴伯 和他的弟兄，都起来建筑 以色列 上帝的坛，要照神人 摩西 律法书上所写的，在坛上献燔祭。
EZRA|3|3|他们在原有的根基上筑坛，因为他们惧怕邻邦民族，又在其上向耶和华早晚献燔祭，
EZRA|3|4|并照律法书上所写的守住棚节，按数照例每日献所当献的燔祭。
EZRA|3|5|此后，他们献常献的燔祭，并在初一和耶和华一切分别为圣的节期献祭，又向耶和华献各人的甘心祭。
EZRA|3|6|从七月初一起，虽然耶和华殿的根基尚未立定，他们开始向耶和华献燔祭。
EZRA|3|7|他们把银子给石匠、木匠，把粮食、酒、油给 西顿 人、 推罗 人，好将香柏树从 黎巴嫩 浮海运到 约帕 ，是照 波斯 王 居鲁士 所允准他们的。
EZRA|3|8|他们到了 耶路撒冷 上帝殿的第二年，二月的时候， 撒拉铁 的儿子 所罗巴伯 ， 约萨达 的儿子 耶书亚 和其余的弟兄，就是祭司和 利未 人，以及所有被掳归回 耶路撒冷 的人，就开工建造；他们派二十岁以上的 利未 人，监督建造耶和华殿的工作。
EZRA|3|9|于是 何达威雅 的后裔，就是 耶书亚 和他的子孙与弟兄、 甲篾 和他的子孙，他们和 利未 人 希拿达 的子孙与弟兄，都起来如同一人，监督那些在上帝殿里做工的人。
EZRA|3|10|工匠立耶和华殿根基的时候，祭司穿礼服吹号， 利未 人 亚萨 的子孙敲钹，都照 以色列 王 大卫 亲手所定的，站着赞美耶和华。
EZRA|3|11|他们彼此唱和，赞美称谢耶和华： “他本为善， 他向 以色列 永施慈爱。” 他们赞美耶和华的时候，众百姓大声呼喊，因为耶和华殿的根基已经立定。
EZRA|3|12|然而有许多祭司、 利未 人和族长，就是见过先前那殿的老年人，现在亲眼看见这殿立了根基，就大声哭号，也有许多人大声欢呼，
EZRA|3|13|百姓不能分辨欢呼的声音或哭号的声音，因为百姓大声呼喊，声音连远处都可听到。
EZRA|4|1|犹大 和 便雅悯 的敌人听说被掳归回的人为耶和华－ 以色列 的上帝建造殿宇，
EZRA|4|2|就去见 所罗巴伯 和族长，对他们说：“请让我们与你们一同建造，因为我们也与你们一样寻求你们的上帝。自从 亚述 王 以撒．哈顿 带我们上这地的日子以来，我们常向上帝献祭。”
EZRA|4|3|但 所罗巴伯 、 耶书亚 和其余 以色列 的族长对他们说：“我们建造上帝的殿与你们无关，因为我们要照 波斯 王 居鲁士 所吩咐的，自己为耶和华－ 以色列 的上帝协力建造。”
EZRA|4|4|那地的人就在 犹大 百姓建造的时候，使他们的手发软，扰乱他们。
EZRA|4|5|从 波斯 王 居鲁士 年间，直到 波斯 王 大流士 在位的时候，那些人贿赂谋士，要破坏他们的计划。
EZRA|4|6|亚哈随鲁 在位，他的国度刚开始的时候，他们上书控告 犹大 和 耶路撒冷 的居民。
EZRA|4|7|亚达薛西 年间， 比施兰 、 米特利达 、 他别 和他们 的同僚上书奏告 波斯 王 亚达薛西 。奏文是用 亚兰 文写的，以 亚兰 文呈上。
EZRA|4|8|利宏 省长、 伸帅 书记也上奏 亚达薛西 王，控告 耶路撒冷 如下
EZRA|4|9|（那时， 利宏 省长、 伸帅 书记和他们其余的同僚，法官、官员、军官、 波斯 官员 、 亚基卫 人、 巴比伦 人，和 书珊迦 人，就是 以拦 人 ，
EZRA|4|10|以及被 亚斯那巴 大人迁移、安置在 撒玛利亚城 和 大河 西边一带地方其余的人。现在 ，
EZRA|4|11|这是他们上奏 亚达薛西 王奏文的抄本）：“ 河西 的臣仆上奏 亚达薛西 王，现在
EZRA|4|12|请王知道，从王那里上到我们这里的 犹太 人，已经抵达 耶路撒冷 。他们正在重建这反叛恶劣的城，已经完成了城墙，正要修复根基。
EZRA|4|13|如今请王知道，这城若再建造，城墙完工，他们就不再进贡、纳粮、缴税，王的国库必受亏损。
EZRA|4|14|如今，我们吃的盐既然全是宫廷的盐，就不忍见王吃亏，因此奏告于王，
EZRA|4|15|请王考察先王史籍，必会在史籍上查知这城是反叛的城，对列王和各省有害；自古以来，城中常有悖逆的事，因此这城曾被拆毁。
EZRA|4|16|我们谨奏王知，这城若再建造，城墙完工， 河西 之地王就无份了。”
EZRA|4|17|那时王谕覆 利宏 省长、 伸帅 书记和他们其余的同僚，就是住 撒玛利亚 和 河西 一带地方的人，说：“愿你们平安。现在
EZRA|4|18|你们所呈给我们的奏本，已经清楚地在我面前读了。
EZRA|4|19|我已下令考查，得知这城自古以来果然背叛列王，其中常有反叛悖逆的事。
EZRA|4|20|也曾有强大的君王治理 耶路撒冷 ，统管 河西 全地，人就给他们进贡、纳粮、缴税。
EZRA|4|21|现在你们要下令叫这些人停工，使这城不得建造，等到我再降旨。
EZRA|4|22|你们当谨慎办这事，不可迟延，何必让损害加重，使王受亏损呢？”
EZRA|4|23|亚达薛西 王上谕的抄本在 利宏 和 伸帅 书记，以及他们的同僚面前宣读，他们就急忙往 耶路撒冷 去见 犹太 人，用势力和强权叫他们停工。
EZRA|4|24|于是，在 耶路撒冷 上帝殿的工程就停止了，直停到 波斯 王 大流士 第二年。
EZRA|5|1|那时， 哈该 先知和 易多 的孙子 撒迦利亚 ，两个先知奉 以色列 上帝的名向 犹大 和 耶路撒冷 的 犹太 人说预言。
EZRA|5|2|于是 撒拉铁 的儿子 所罗巴伯 和 约萨达 的儿子 耶书亚 起来，开始建造 耶路撒冷 上帝的殿，有上帝的先知在那里帮助他们。
EZRA|5|3|当时 河西 的 达乃 总督和 示他．波斯乃 ，以及他们的同僚来对 犹太 人这样说：“谁降旨让你们建造这殿，完成这建筑呢？”
EZRA|5|4|于是我们告诉他们建造这建筑物的人叫什么名字。
EZRA|5|5|但上帝的眼目看顾 犹太 人的长老，以致没有人叫他们停工，直到奏文上告 大流士 ，得着他对这事的回谕。
EZRA|5|6|这是 河西 的 达乃 总督和 示他．波斯乃 ，以及他们的同僚，就是住 河西 的官员 ，上书奏告 大流士 王的抄本，
EZRA|5|7|他们上书给王的奏文，其中写着：“愿 大流士 王诸事平安。
EZRA|5|8|请王知道，我们往 犹大 省去，到了至大上帝的殿。这殿是用凿成的石头建造的，梁木插入墙内。这项工程进行迅速，在他们手中顺利。
EZRA|5|9|于是我们问那些长老，对他们这样说：‘谁降旨让你们建造这殿，完成这建筑呢？’
EZRA|5|10|我们又问他们的名字，要记下他们领袖的名字，奏告于王。
EZRA|5|11|他们这样回答我们说：‘我们是天和地之上帝的仆人，重建多年前所建造的殿，就是 以色列 一位伟大的君王建造完成的。
EZRA|5|12|但因我们祖先惹天上的上帝发怒，上帝把他们交在 迦勒底 人 巴比伦 王 尼布甲尼撒 的手中，他就拆毁这殿，又把百姓掳到 巴比伦 。
EZRA|5|13|然而 巴比伦 王 居鲁士 元年，他降旨允准建造上帝的这殿。
EZRA|5|14|上帝殿中的金银器皿，就是 尼布甲尼撒 从 耶路撒冷 殿中掠取带到 巴比伦 庙里的， 居鲁士 王从 巴比伦 庙里取出来，交给派为省长，名叫 设巴萨 的，
EZRA|5|15|对他说：可以将这些器皿带去，放在 耶路撒冷 的殿中，在原处建造上帝的殿。
EZRA|5|16|于是那位 设巴萨 来建立 耶路撒冷 上帝殿的根基。但从那时直到如今，这殿尚未修建完毕。’
EZRA|5|17|现在，王若以为好，请查阅 巴比伦 王的档案库，看 居鲁士 王有没有降旨允准在 耶路撒冷 建造上帝的殿。请降旨指示我们王对这件事的心意。”
EZRA|6|1|于是 大流士 王降旨，要寻察典籍库，就是在 巴比伦 藏档案之处；
EZRA|6|2|在 玛代 省 亚马他城 的宫内寻得一卷，其中这样写着，“纪录如下：
EZRA|6|3|居鲁士 王元年，王降旨论到在 耶路撒冷 上帝的殿，要建造这殿作为献祭之处，坚固它的根基。殿高六十肘，宽六十肘，
EZRA|6|4|要用三层凿成的石头，一层木头 ，经费可出于王的库房。
EZRA|6|5|至于上帝殿的金银器皿，就是 尼布甲尼撒 从 耶路撒冷 的殿中掠取带到 巴比伦 的，必须归还，带回 耶路撒冷 的殿中，各按原处放在上帝的殿里。”
EZRA|6|6|“现在， 河西 的 达乃 总督和 示他．波斯乃 ，以及他们的同僚，就是住 河西 的官员，你们当远离那里。
EZRA|6|7|不要拦阻这上帝殿的工作，任由 犹太 人的省长和长老在原处建造上帝的这殿。
EZRA|6|8|我又降旨，吩咐你们为建造上帝的殿当向 犹太 人的长老这样行：从王的财产中，由 河西 所缴纳的贡银，迅速支付这些人，免得工程停顿。
EZRA|6|9|他们向天上的上帝献燔祭所需用的公牛犊、公绵羊、小绵羊，以及麦子、盐、酒、油，都要照 耶路撒冷 祭司的话，每日供给他们，不得有误；
EZRA|6|10|好叫他们献馨香的祭给天上的上帝，又为王和王众子的寿命祈祷。
EZRA|6|11|我再降旨，无论谁更改这命令，必从他房屋中拆出一根梁木，把他举起，悬在其上，又使他的房屋为此成为粪堆。
EZRA|6|12|任何王或百姓若伸手更改这命令，拆毁在 耶路撒冷 上帝的这殿，愿那立他名在那里的上帝将他们灭绝。我 大流士 降这谕旨，你们要速速遵行。”
EZRA|6|13|于是， 河西 的 达乃 总督和 示他．波斯乃 ，以及他们的同僚，急速遵行 大流士 王所颁的命令。
EZRA|6|14|犹太 人的长老因 哈该 先知和 易多 的孙子 撒迦利亚 的预言，就建造这殿，凡事顺利。他们遵照 以色列 上帝的命令和 波斯 王 居鲁士 、 大流士 、 亚达薛西 的谕旨，建造完毕。
EZRA|6|15|大流士 王第六年，亚达月初三，这殿完工了。
EZRA|6|16|以色列 人、祭司和 利未 人，以及其余被掳归回的人都欢欢喜喜地为上帝的这殿行奉献礼。
EZRA|6|17|他们为这上帝殿的奉献礼献了一百头公牛，二百只公绵羊，四百只小绵羊，又照 以色列 支派的数目献十二只公山羊，作 以色列 众人的赎罪祭。
EZRA|6|18|他们派祭司按着班次， 利未 人也按着班次在 耶路撒冷 事奉上帝，正如 摩西 律法书上所写的。
EZRA|6|19|正月十四日，被掳归回的人守逾越节。
EZRA|6|20|祭司和 利未 人一同自洁，他们全都洁净了。 利未 人为被掳归回的众人和他们的弟兄众祭司，并为自己宰逾越节的羔羊。
EZRA|6|21|从被掳之地归回的 以色列 人，并所有归附他们、除掉这地外邦人的污秽、寻求耶和华－ 以色列 上帝的人，都吃这羔羊。
EZRA|6|22|他们欢欢喜喜地守除酵节七日，因为耶和华使他们欢喜。耶和华又使 亚述 王的心转向他们，坚固他们的手，去做上帝－ 以色列 上帝殿的工。
EZRA|7|1|这些事以后， 波斯 王 亚达薛西 在位的时候，有个人叫 以斯拉 ，他是 西莱雅 的儿子， 西莱雅 是 亚撒利雅 的儿子， 亚撒利雅 是 希勒家 的儿子，
EZRA|7|2|希勒家 是 沙龙 的儿子， 沙龙 是 撒督 的儿子， 撒督 是 亚希突 的儿子，
EZRA|7|3|亚希突 是 亚玛利雅 的儿子， 亚玛利雅 是 亚撒利雅 的儿子， 亚撒利雅 是 米拉约 的儿子，
EZRA|7|4|米拉约 是 西拉希雅 的儿子， 西拉希雅 是 乌西 的儿子， 乌西 是 布基 的儿子，
EZRA|7|5|布基 是 亚比书 的儿子， 亚比书 是 非尼哈 的儿子， 非尼哈 是 以利亚撒 的儿子， 以利亚撒 是 亚伦 大祭司的儿子。
EZRA|7|6|这 以斯拉 从 巴比伦 上来，他是一个文士，精通耶和华－ 以色列 上帝所赐 摩西 的律法。王允准他一切所求的，因为耶和华－他上帝的手帮助他。
EZRA|7|7|亚达薛西 王第七年，有些 以色列 人、一些祭司、 利未 人、歌唱的、门口的守卫、殿役，上 耶路撒冷 去。
EZRA|7|8|王第七年五月， 以斯拉 到了 耶路撒冷 。
EZRA|7|9|正月初一，他从 巴比伦 起程，五月初一就到了 耶路撒冷 ，因为他上帝施恩的手帮助他。
EZRA|7|10|以斯拉 立志考究遵行耶和华的律法，又将律例典章教导 以色列 人。
EZRA|7|11|亚达薛西 王赐给精通耶和华诫命和 以色列 律例的文士 以斯拉 祭司的谕旨，抄本如下：
EZRA|7|12|“诸王之王 亚达薛西 ，达于精通天上之上帝律法的 以斯拉 祭司文士等等：现在
EZRA|7|13|住在我国中的 以色列 百姓、祭司、 利未 人，凡愿意上 耶路撒冷 去的，我降旨准他们与你同去。
EZRA|7|14|既然王与七个谋士派你去，照你手中上帝的律法视察 犹大 和 耶路撒冷 的景况；
EZRA|7|15|你又带着王和谋士乐意献给住 耶路撒冷 、 以色列 上帝的金银，
EZRA|7|16|和你在 巴比伦 全省所得的一切金银，以及百姓、祭司甘心献给 耶路撒冷 他们上帝殿的礼物，
EZRA|7|17|那么，你就当用这银子急速买公牛、公绵羊、小绵羊，和同献的素祭、浇酒祭，献在 耶路撒冷 你们上帝殿的坛上。
EZRA|7|18|剩下的金银，你和你的弟兄看怎样好，就怎样用，但总要遵照你们上帝的旨意。
EZRA|7|19|你要带着交托给你、在上帝殿中事奉用的器皿，到 耶路撒冷 上帝面前。
EZRA|7|20|你上帝殿里若再有需用的经费，是你负责供应的，可以从王的宝库里支取。
EZRA|7|21|“我 亚达薛西 王又降旨达于 河西 所有的司库：‘精通天上之上帝律法的 以斯拉 祭司文士无论向你们要什么，你们要速速办理，
EZRA|7|22|直至一百他连得银子，一百柯珥 麦子，一百罢特酒，一百罢特油，盐不限其数。
EZRA|7|23|凡天上之上帝所吩咐的，当为天上之上帝的殿切实办理。何必使愤怒临到王和王众子的国呢？
EZRA|7|24|我再吩咐你们：至于任何祭司、 利未 人、歌唱的、门口的守卫和殿役，以及在上帝的这殿事奉的人，不可要求他们进贡，纳粮，缴税。’
EZRA|7|25|“你， 以斯拉 啊，要照着你上帝赐你的智慧，指派所有明白你上帝律法的人作官长、审判官，治理 河西 所有的百姓，教导不明白上帝律法的人。
EZRA|7|26|凡不遵行你上帝律法和王命令的人，当速速定他的罪，或处死，或充军，或抄家，或囚禁。”
EZRA|7|27|以斯拉 说：“耶和华－我们列祖的上帝是应当称颂的！因他使王起这心愿，使 耶路撒冷 耶和华的殿得荣耀，
EZRA|7|28|他又在王和谋士，以及王所有大能的军官面前施恩于我。我因耶和华－我上帝的手的帮助，得以坚强，从 以色列 中召集领袖，与我一同上来。”
EZRA|8|1|这些是 亚达薛西 王在位的时候，同我从 巴比伦 上来的族长和他们的家谱：
EZRA|8|2|属 非尼哈 的子孙有 革顺 ；属 以他玛 的子孙有 但以理 ；属 大卫 的子孙有 哈突 ；
EZRA|8|3|属 示迦尼 的子孙；属 巴录 的子孙有 撒迦利亚 ，同着他按家谱计算，男丁一百五十人；
EZRA|8|4|属 巴哈．摩押 的子孙有 西拉希雅 的儿子 以利约乃 ，同着他有男丁二百人；
EZRA|8|5|属 萨土 的子孙有 雅哈悉 的儿子 示迦尼 ，同着他有男丁三百人；
EZRA|8|6|属 亚丁 的子孙有 约拿单 的儿子 以别 ，同着他有男丁五十人；
EZRA|8|7|属 以拦 的子孙有 亚他利雅 的儿子 耶筛亚 ，同着他有男丁七十人；
EZRA|8|8|属 示法提雅 的子孙有 米迦勒 的儿子 西巴第雅 ，同着他有男丁八十人；
EZRA|8|9|属 约押 的子孙有 耶歇 的儿子 俄巴底亚 ，同着他有男丁二百一十八人；
EZRA|8|10|属 巴尼 的子孙有 约细斐 的儿子 示罗密 ，同着他有男丁一百六十人；
EZRA|8|11|属 比拜 的子孙有 比拜 的儿子 撒迦利亚 ，同着他有男丁二十八人；
EZRA|8|12|属 押甲 的子孙有 哈加坦 的儿子 约哈难 ，同着他有男丁一百一十人；
EZRA|8|13|属 亚多尼干 的子孙，就是晚到的，他们的名字是 以利法列 、 耶利 、 示玛雅 ，同着他们有男丁六十人；
EZRA|8|14|属 比革瓦伊 的子孙有 乌太 和 撒刻 ，同着他们有男丁七十人。
EZRA|8|15|我召集这些人在流入 亚哈瓦 的河旁边，我们在那里扎营三日。我查看百姓和祭司，发现并没有 利未 人在那里，
EZRA|8|16|就派人到 以利以谢 、 亚列 、 示玛雅 、 以利拿单 、 雅立 、 以利拿单 、 拿单 、 撒迦利亚 、 米书兰 等领袖，以及 约雅立 和 以利拿单 教师那里。
EZRA|8|17|我吩咐他们往 迦西斐雅 地方去见那里的领袖 易多 ，又告诉他们当向 易多 和他的弟兄，就是 迦西斐雅 那地方的殿役说什么话，好为我们上帝的殿带事奉的人来。
EZRA|8|18|蒙我们上帝施恩的手帮助我们，他们在 以色列 的曾孙， 利未 的孙子， 抹利 的后裔中带了一个精明的人来，就是 示利比 ，还有他的众子与兄弟共十八人。
EZRA|8|19|另外，还有 哈沙比雅 ，同着他有 米拉利 的子孙 耶筛亚 ，以及他的众子和兄弟共二十人。
EZRA|8|20|从前 大卫 和众领袖派殿役服事 利未 人，现在从这殿役中也带了二百二十人来，全都是按名指定的。
EZRA|8|21|那时，我在 亚哈瓦河 边宣告禁食，为要在我们上帝面前刻苦己心，求他使我们和我们的孩子，以及一切所有的，都得平坦的道路。
EZRA|8|22|我以求王拨步兵骑兵帮助我们抵挡路上的仇敌为羞愧，因我们曾对王说：“我们上帝施恩的手必帮助凡寻求他的，但他的能力和愤怒必攻击凡离弃他的。”
EZRA|8|23|我们为此禁食祈求我们的上帝，他就应允我们。
EZRA|8|24|我分派十二位祭司长，就是 示利比 、 哈沙比雅 和与他们一起的兄弟十人，
EZRA|8|25|把王和谋士、军官，并在那里的 以色列 众人为我们上帝殿所献的金银和器皿，都秤了交给他们。
EZRA|8|26|我秤了交在他们手中的有六百五十他连得银子，一百他连得银器，一百他连得金子，
EZRA|8|27|二十个金碗，值一千达利克，上等光亮的铜器皿两个，珍贵如金。
EZRA|8|28|我对他们说：“你们归耶和华为圣，器皿也归为圣；金银是甘心献给耶和华－你们列祖之上帝的。
EZRA|8|29|你们要警醒看守，直到你们在祭司长和 利未 族长，以及 以色列 的各族长面前，在 耶路撒冷 耶和华殿的库房内，把这些过了秤。”
EZRA|8|30|于是，祭司和 利未 人把秤过的金银和器皿接过来，要带到 耶路撒冷 我们上帝的殿里。
EZRA|8|31|正月十二日，我们从 亚哈瓦河 边起行，要往 耶路撒冷 去。我们上帝的手保佑我们，救我们脱离仇敌和路上埋伏之人的手。
EZRA|8|32|我们到了 耶路撒冷 ，在那里住了三日。
EZRA|8|33|第四日，金银和器皿都在我们上帝的殿里过了秤，交在 乌利亚 的儿子 米利末 祭司的手中。同着他的有 非尼哈 的儿子 以利亚撒 ，还有 利未 人 耶书亚 的儿子 约撒拔 和 宾内 的儿子 挪亚底 。
EZRA|8|34|那时，这一切都点过秤过了，重量全写在册上。
EZRA|8|35|从被掳之地归回的人向 以色列 的上帝献燔祭，为 以色列 众人献十二头公牛，九十六只公绵羊，七十七只小绵羊，又献十二只公山羊作赎罪祭，这些全都是献给耶和华的燔祭。
EZRA|8|36|被掳归回的人把王的谕旨交给王的总督与 河西 的省长，他们就支助百姓和上帝的殿。
EZRA|9|1|这些事完成以后，众领袖来接近我，说：“ 以色列 百姓、祭司和 利未 人没有弃绝 迦南 人、 赫 人、 比利洗 人、 耶布斯 人、 亚扪 人、 摩押 人、 埃及 人和 亚摩利 人等列邦民族所行可憎的事。
EZRA|9|2|因他们为自己和儿子娶了这些外邦女子，以致圣洁的种籽和列邦民族混杂，而且领袖和官长在这事上是罪魁。”
EZRA|9|3|我一听见这事，就撕裂衣服和外袍，拔了头发和胡须，惊惶地坐着。
EZRA|9|4|凡为 以色列 上帝言语战兢的人，都因被掳归回之人所犯的罪，聚集到我这里来。我惊惶地坐着，直到献晚祭的时候。
EZRA|9|5|献晚祭的时候我从愁烦中起来，穿着撕裂的衣服和外袍，双膝跪下，向耶和华－我的上帝举手，
EZRA|9|6|说： “我的上帝啊，我抱愧蒙羞，不敢向你－我的上帝仰面，因为我们的罪孽多到灭顶，我们的罪恶滔天。
EZRA|9|7|从我们祖先的日子直到今日，我们的罪恶深重；因我们的罪孽，我们和君王、祭司都交在邻国诸王的手中，被杀害，掳掠，抢夺，脸上蒙羞，正如今日的景况。
EZRA|9|8|现在耶和华－我们的上帝暂且向我们施恩，为我们留下一些残存之民，使我们如钉子钉在他的圣所，好让我们的上帝光照我们的眼目，使我们在受辖制之中稍微复兴。
EZRA|9|9|我们是奴仆，然而在受辖制之中，我们的上帝没有丢弃我们，在 波斯 诸王面前向我们施恩，叫我们复兴，能重建我们上帝的殿，修补毁坏之处，使我们在 犹大 和 耶路撒冷 有城墙。
EZRA|9|10|“我们的上帝啊，既然如此，现在我们还有什么话可说呢？因为我们离弃了你的诫命，
EZRA|9|11|就是你藉你仆人众先知所吩咐的，说：‘你们要去得为业之地是污秽之地，因列邦民族的污秽和可憎的事，叫这地从这边到那边都充满了污秽。
EZRA|9|12|现在，不可把你们的女儿嫁给他们的儿子，也不可为你们的儿子娶他们的女儿，永不可求他们的平安和他们的利益，这样你们就可以强盛，吃这地的美物，并把这地留给你们的子孙永远为业。’
EZRA|9|13|我们因自己的恶行和大罪，遭遇这一切的事，但你－我们的上帝惩罚我们轻于我们罪所当得的，又为我们留下这些残存之民。
EZRA|9|14|我们岂可再违背你的诫命，与行这些可憎之事的民族结亲呢？若我们这样行，你岂不向我们发怒，将我们灭绝，以致没有一个余民或残存之民吗？
EZRA|9|15|耶和华－ 以色列 的上帝啊，你是公义的，我们才能剩下这些残存之民，正如今日的景况。看哪，我们在你面前有罪恶，因此无人能在你面前站立得住。”
EZRA|10|1|以斯拉 祷告，认罪，哭泣，俯伏在上帝殿前的时候，有 以色列 中的男女和孩童聚集到 以斯拉 那里，成了一个盛大的会，百姓无不痛哭。
EZRA|10|2|以拦 的子孙， 耶歇 的儿子 示迦尼 对 以斯拉 说：“我们娶了这地的外邦女子，干犯了我们的上帝，然而现在 以色列 人在这事上还有指望。
EZRA|10|3|现在，我们要与我们的上帝立约，送走所有的妻子和她们所生的，照着主和那些因我们上帝诫命战兢之人所议定的，按律法去行。
EZRA|10|4|起来，这是你当办的事，我们必支持你，你当奋勇而行。”
EZRA|10|5|以斯拉 就起来，叫祭司长和 利未 人，以及 以色列 众人起誓，要照这话去做；他们就起了誓。
EZRA|10|6|以斯拉 从上帝殿前起来，进入 以利亚实 的儿子 约哈难 的屋里，到了那里不吃饭，也不喝水，为被掳归回之人所犯的罪悲伤。
EZRA|10|7|他们通告 犹大 和 耶路撒冷 ，叫所有被掳归回的人聚集在 耶路撒冷 。
EZRA|10|8|凡不遵照领袖和长老所议定，三日之内不来的，就必毁坏他所有的财产，把他从被掳归回之人的会中开除。
EZRA|10|9|于是， 犹大 和 便雅悯 众人三日之内都聚集在 耶路撒冷 。那时是九月，那月的二十日，众百姓坐在上帝殿前的广场，因这事，又因下大雨，就都战抖。
EZRA|10|10|以斯拉 祭司站起来，对他们说：“你们有罪了，因为你们娶了外邦女子，增添 以色列 的罪恶。
EZRA|10|11|现在当向耶和华－你们列祖的上帝认罪，遵行他的旨意，离开这地的百姓和外邦女子。”
EZRA|10|12|全会众大声回答说：“好！我们必照着你的话去做。
EZRA|10|13|只是百姓众多，又逢大雨的季节，我们没有气力站在外面；这也不是一两天可以办完的事，因我们在这事上犯了大罪。
EZRA|10|14|让我们的领袖代表全会众留在那里。我们城镇中凡娶外邦女子的，当按所定的日期，会同本城的长老和审判官前来，直到办完这事，上帝的烈怒转离我们 。”
EZRA|10|15|惟有 亚撒黑 的儿子 约拿单 ， 特瓦 的儿子 雅哈谢 反对这事，并有 米书兰 和 利未 人 沙比太 支持他们。
EZRA|10|16|被掳归回的人就如此做了。 以斯拉 祭司按着父家指名选派一些族长 。十月初一，他们一同坐下来查办这事，
EZRA|10|17|到正月初一，才查清所有娶外邦女子的人数。
EZRA|10|18|在祭司中查出娶外邦女子的： 耶书亚 的子孙中，有 约萨达 的儿子，和他兄弟 玛西雅 、 以利以谢 、 雅立 、 基大利 ，
EZRA|10|19|他们承诺要送走他们的妻子。他们因有罪，就献羊群中的一只公绵羊赎罪；
EZRA|10|20|音麦 的子孙中，有 哈拿尼 、 西巴第雅 ；
EZRA|10|21|哈琳 的子孙中，有 玛西雅 、 以利雅 、 示玛雅 、 耶歇 、 乌西雅 ；
EZRA|10|22|巴施户珥 的子孙中，有 以利约乃 、 玛西雅 、 以实玛利 、 拿坦业 、 约撒拔 、 以利亚萨 。
EZRA|10|23|利未 人中，有 约撒拔 、 示每 、 基拉雅 ， 基拉雅 就是 基利他 ，还有 毗他希雅 、 犹大 、 以利以谢 。
EZRA|10|24|歌唱的人中有 以利亚实 。门口的守卫中，有 沙龙 、 提联 、 乌利 。
EZRA|10|25|以色列 人 巴录 的子孙中，有 拉米 、 耶西雅 、 玛基雅 、 米雅民 、 以利亚撒 、 玛基雅 、 比拿雅 。
EZRA|10|26|以拦 的子孙中，有 玛他尼 、 撒迦利亚 、 耶歇 、 押底 、 耶列末 、 以利雅 。
EZRA|10|27|萨土 的子孙中，有 以利约乃 、 以利亚实 、 玛他尼 、 耶列末 、 撒拔 、 亚西撒 。
EZRA|10|28|比拜 的子孙中，有 约哈难 、 哈拿尼雅 、 萨拜 、 亚勒 。
EZRA|10|29|巴尼 的子孙中，有 米书兰 、 玛鹿 、 亚大雅 、 雅述 、 示押 、 拉末 。
EZRA|10|30|巴哈．摩押 的子孙中，有 阿底拿 、 基拉 、 比拿雅 、 玛西雅 、 玛他尼 、 比撒列 、 宾内 、 玛拿西 。
EZRA|10|31|哈琳 的子孙中，有 以利以谢 、 伊示雅 、 玛基雅 、 示玛雅 、 西缅 、
EZRA|10|32|便雅悯 、 玛鹿 、 示玛利雅 。
EZRA|10|33|哈顺 的子孙中，有 玛特乃 、 玛达他 、 撒拔 、 以利法列 、 耶利买 、 玛拿西 、 示每 。
EZRA|10|34|巴尼 的子孙中，有 玛玳 、 暗兰 、 乌益 、
EZRA|10|35|比拿雅 、 比底雅 、 基禄 、
EZRA|10|36|瓦尼雅 、 米利末 、 以利亚实 、
EZRA|10|37|玛他尼 、 玛特乃 、 雅扫 、
EZRA|10|38|巴尼 、 宾内 、 示每 、
EZRA|10|39|示利米雅 、 拿单 、 亚大雅 、
EZRA|10|40|玛拿底拜 、 沙赛 、 沙赖 、
EZRA|10|41|亚萨利 、 示利米雅 、 示玛利雅 、
EZRA|10|42|沙龙 、 亚玛利雅 、 约瑟 。
EZRA|10|43|尼波 的子孙中，有 耶利 、 玛他提雅 、 撒拔 、 西比拿 、 雅玳 、 约珥 、 比拿雅 。
EZRA|10|44|这些人全都娶了外邦女子，其中也有生了儿女的 。
