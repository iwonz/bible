NEH|1|1|The words of Nehemiah the son of Hachaliah. And it came to pass in the month Chisleu, in the twentieth year, as I was in Shushan the palace,
NEH|1|2|That Hanani, one of my brethren, came, he and certain men of Judah; and I asked them concerning the Jews that had escaped, which were left of the captivity, and concerning Jerusalem.
NEH|1|3|And they said unto me, The remnant that are left of the captivity there in the province are in great affliction and reproach: the wall of Jerusalem also is broken down, and the gates thereof are burned with fire.
NEH|1|4|And it came to pass, when I heard these words, that I sat down and wept, and mourned certain days, and fasted, and prayed before the God of heaven,
NEH|1|5|And said, I beseech thee, O LORD God of heaven, the great and terrible God, that keepeth covenant and mercy for them that love him and observe his commandments:
NEH|1|6|Let thine ear now be attentive, and thine eyes open, that thou mayest hear the prayer of thy servant, which I pray before thee now, day and night, for the children of Israel thy servants, and confess the sins of the children of Israel, which we have sinned against thee: both I and my father's house have sinned.
NEH|1|7|We have dealt very corruptly against thee, and have not kept the commandments, nor the statutes, nor the judgments, which thou commandedst thy servant Moses.
NEH|1|8|Remember, I beseech thee, the word that thou commandedst thy servant Moses, saying, If ye transgress, I will scatter you abroad among the nations:
NEH|1|9|But if ye turn unto me, and keep my commandments, and do them; though there were of you cast out unto the uttermost part of the heaven, yet will I gather them from thence, and will bring them unto the place that I have chosen to set my name there.
NEH|1|10|Now these are thy servants and thy people, whom thou hast redeemed by thy great power, and by thy strong hand.
NEH|1|11|O LORD, I beseech thee, let now thine ear be attentive to the prayer of thy servant, and to the prayer of thy servants, who desire to fear thy name: and prosper, I pray thee, thy servant this day, and grant him mercy in the sight of this man. For I was the king's cupbearer.
NEH|2|1|And it came to pass in the month Nisan, in the twentieth year of Artaxerxes the king, that wine was before him: and I took up the wine, and gave it unto the king. Now I had not been beforetime sad in his presence.
NEH|2|2|Wherefore the king said unto me, Why is thy countenance sad, seeing thou art not sick? this is nothing else but sorrow of heart. Then I was very sore afraid,
NEH|2|3|And said unto the king, Let the king live for ever: why should not my countenance be sad, when the city, the place of my fathers' sepulchres, lieth waste, and the gates thereof are consumed with fire?
NEH|2|4|Then the king said unto me, For what dost thou make request? So I prayed to the God of heaven.
NEH|2|5|And I said unto the king, If it please the king, and if thy servant have found favour in thy sight, that thou wouldest send me unto Judah, unto the city of my fathers' sepulchres, that I may build it.
NEH|2|6|And the king said unto me, (the queen also sitting by him,) For how long shall thy journey be? and when wilt thou return? So it pleased the king to send me; and I set him a time.
NEH|2|7|Moreover I said unto the king, If it please the king, let letters be given me to the governors beyond the river, that they may convey me over till I come into Judah;
NEH|2|8|And a letter unto Asaph the keeper of the king's forest, that he may give me timber to make beams for the gates of the palace which appertained to the house, and for the wall of the city, and for the house that I shall enter into. And the king granted me, according to the good hand of my God upon me.
NEH|2|9|Then I came to the governors beyond the river, and gave them the king's letters. Now the king had sent captains of the army and horsemen with me.
NEH|2|10|When Sanballat the Horonite, and Tobiah the servant, the Ammonite, heard of it, it grieved them exceedingly that there was come a man to seek the welfare of the children of Israel.
NEH|2|11|So I came to Jerusalem, and was there three days.
NEH|2|12|And I arose in the night, I and some few men with me; neither told I any man what my God had put in my heart to do at Jerusalem: neither was there any beast with me, save the beast that I rode upon.
NEH|2|13|And I went out by night by the gate of the valley, even before the dragon well, and to the dung port, and viewed the walls of Jerusalem, which were broken down, and the gates thereof were consumed with fire.
NEH|2|14|Then I went on to the gate of the fountain, and to the king's pool: but there was no place for the beast that was under me to pass.
NEH|2|15|Then went I up in the night by the brook, and viewed the wall, and turned back, and entered by the gate of the valley, and so returned.
NEH|2|16|And the rulers knew not whither I went, or what I did; neither had I as yet told it to the Jews, nor to the priests, nor to the nobles, nor to the rulers, nor to the rest that did the work.
NEH|2|17|Then said I unto them, Ye see the distress that we are in, how Jerusalem lieth waste, and the gates thereof are burned with fire: come, and let us build up the wall of Jerusalem, that we be no more a reproach.
NEH|2|18|Then I told them of the hand of my God which was good upon me; as also the king's words that he had spoken unto me. And they said, Let us rise up and build. So they strengthened their hands for this good work.
NEH|2|19|But when Sanballat the Horonite, and Tobiah the servant, the Ammonite, and Geshem the Arabian, heard it, they laughed us to scorn, and despised us, and said, What is this thing that ye do? will ye rebel against the king?
NEH|2|20|Then answered I them, and said unto them, The God of heaven, he will prosper us; therefore we his servants will arise and build: but ye have no portion, nor right, nor memorial, in Jerusalem.
NEH|3|1|Then Eliashib the high priest rose up with his brethren the priests, and they builded the sheep gate; they sanctified it, and set up the doors of it; even unto the tower of Meah they sanctified it, unto the tower of Hananeel.
NEH|3|2|And next unto him builded the men of Jericho. And next to them builded Zaccur the son of Imri.
NEH|3|3|But the fish gate did the sons of Hassenaah build, who also laid the beams thereof, and set up the doors thereof, the locks thereof, and the bars thereof.
NEH|3|4|And next unto them repaired Meremoth the son of Urijah, the son of Koz. And next unto them repaired Meshullam the son of Berechiah, the son of Meshezabeel. And next unto them repaired Zadok the son of Baana.
NEH|3|5|And next unto them the Tekoites repaired; but their nobles put not their necks to the work of their LORD.
NEH|3|6|Moreover the old gate repaired Jehoiada the son of Paseah, and Meshullam the son of Besodeiah; they laid the beams thereof, and set up the doors thereof, and the locks thereof, and the bars thereof.
NEH|3|7|And next unto them repaired Melatiah the Gibeonite, and Jadon the Meronothite, the men of Gibeon, and of Mizpah, unto the throne of the governor on this side the river.
NEH|3|8|Next unto him repaired Uzziel the son of Harhaiah, of the goldsmiths. Next unto him also repaired Hananiah the son of one of the apothecaries, and they fortified Jerusalem unto the broad wall.
NEH|3|9|And next unto them repaired Rephaiah the son of Hur, the ruler of the half part of Jerusalem.
NEH|3|10|And next unto them repaired Jedaiah the son of Harumaph, even over against his house. And next unto him repaired Hattush the son of Hashabniah.
NEH|3|11|Malchijah the son of Harim, and Hashub the son of Pahathmoab, repaired the other piece, and the tower of the furnaces.
NEH|3|12|And next unto him repaired Shallum the son of Halohesh, the ruler of the half part of Jerusalem, he and his daughters.
NEH|3|13|The valley gate repaired Hanun, and the inhabitants of Zanoah; they built it, and set up the doors thereof, the locks thereof, and the bars thereof, and a thousand cubits on the wall unto the dung gate.
NEH|3|14|But the dung gate repaired Malchiah the son of Rechab, the ruler of part of Bethhaccerem; he built it, and set up the doors thereof, the locks thereof, and the bars thereof.
NEH|3|15|But the gate of the fountain repaired Shallun the son of Colhozeh, the ruler of part of Mizpah; he built it, and covered it, and set up the doors thereof, the locks thereof, and the bars thereof, and the wall of the pool of Siloah by the king's garden, and unto the stairs that go down from the city of David.
NEH|3|16|After him repaired Nehemiah the son of Azbuk, the ruler of the half part of Bethzur, unto the place over against the sepulchres of David, and to the pool that was made, and unto the house of the mighty.
NEH|3|17|After him repaired the Levites, Rehum the son of Bani. Next unto him repaired Hashabiah, the ruler of the half part of Keilah, in his part.
NEH|3|18|After him repaired their brethren, Bavai the son of Henadad, the ruler of the half part of Keilah.
NEH|3|19|And next to him repaired Ezer the son of Jeshua, the ruler of Mizpah, another piece over against the going up to the armoury at the turning of the wall.
NEH|3|20|After him Baruch the son of Zabbai earnestly repaired the other piece, from the turning of the wall unto the door of the house of Eliashib the high priest.
NEH|3|21|After him repaired Meremoth the son of Urijah the son of Koz another piece, from the door of the house of Eliashib even to the end of the house of Eliashib.
NEH|3|22|And after him repaired the priests, the men of the plain.
NEH|3|23|After him repaired Benjamin and Hashub over against their house. After him repaired Azariah the son of Maaseiah the son of Ananiah by his house.
NEH|3|24|After him repaired Binnui the son of Henadad another piece, from the house of Azariah unto the turning of the wall, even unto the corner.
NEH|3|25|Palal the son of Uzai, over against the turning of the wall, and the tower which lieth out from the king's high house, that was by the court of the prison. After him Pedaiah the son of Parosh.
NEH|3|26|Moreover the Nethinims dwelt in Ophel, unto the place over against the water gate toward the east, and the tower that lieth out.
NEH|3|27|After them the Tekoites repaired another piece, over against the great tower that lieth out, even unto the wall of Ophel.
NEH|3|28|From above the horse gate repaired the priests, every one over against his house.
NEH|3|29|After them repaired Zadok the son of Immer over against his house. After him repaired also Shemaiah the son of Shechaniah, the keeper of the east gate.
NEH|3|30|After him repaired Hananiah the son of Shelemiah, and Hanun the sixth son of Zalaph, another piece. After him repaired Meshullam the son of Berechiah over against his chamber.
NEH|3|31|After him repaired Malchiah the goldsmith's son unto the place of the Nethinims, and of the merchants, over against the gate Miphkad, and to the going up of the corner.
NEH|3|32|And between the going up of the corner unto the sheep gate repaired the goldsmiths and the merchants.
NEH|4|1|But it came to pass, that when Sanballat heard that we builded the wall, he was wroth, and took great indignation, and mocked the Jews.
NEH|4|2|And he spake before his brethren and the army of Samaria, and said, What do these feeble Jews? will they fortify themselves? will they sacrifice? will they make an end in a day? will they revive the stones out of the heaps of the rubbish which are burned?
NEH|4|3|Now Tobiah the Ammonite was by him, and he said, Even that which they build, if a fox go up, he shall even break down their stone wall.
NEH|4|4|Hear, O our God; for we are despised: and turn their reproach upon their own head, and give them for a prey in the land of captivity:
NEH|4|5|And cover not their iniquity, and let not their sin be blotted out from before thee: for they have provoked thee to anger before the builders.
NEH|4|6|So built we the wall; and all the wall was joined together unto the half thereof: for the people had a mind to work.
NEH|4|7|But it came to pass, that when Sanballat, and Tobiah, and the Arabians, and the Ammonites, and the Ashdodites, heard that the walls of Jerusalem were made up, and that the breaches began to be stopped, then they were very wroth,
NEH|4|8|And conspired all of them together to come and to fight against Jerusalem, and to hinder it.
NEH|4|9|Nevertheless we made our prayer unto our God, and set a watch against them day and night, because of them.
NEH|4|10|And Judah said, The strength of the bearers of burdens is decayed, and there is much rubbish; so that we are not able to build the wall.
NEH|4|11|And our adversaries said, They shall not know, neither see, till we come in the midst among them, and slay them, and cause the work to cease.
NEH|4|12|And it came to pass, that when the Jews which dwelt by them came, they said unto us ten times, From all places whence ye shall return unto us they will be upon you.
NEH|4|13|Therefore set I in the lower places behind the wall, and on the higher places, I even set the people after their families with their swords, their spears, and their bows.
NEH|4|14|And I looked, and rose up, and said unto the nobles, and to the rulers, and to the rest of the people, Be not ye afraid of them: remember the LORD, which is great and terrible, and fight for your brethren, your sons, and your daughters, your wives, and your houses.
NEH|4|15|And it came to pass, when our enemies heard that it was known unto us, and God had brought their counsel to nought, that we returned all of us to the wall, every one unto his work.
NEH|4|16|And it came to pass from that time forth, that the half of my servants wrought in the work, and the other half of them held both the spears, the shields, and the bows, and the habergeons; and the rulers were behind all the house of Judah.
NEH|4|17|They which builded on the wall, and they that bare burdens, with those that laded, every one with one of his hands wrought in the work, and with the other hand held a weapon.
NEH|4|18|For the builders, every one had his sword girded by his side, and so builded. And he that sounded the trumpet was by me.
NEH|4|19|And I said unto the nobles, and to the rulers, and to the rest of the people, The work is great and large, and we are separated upon the wall, one far from another.
NEH|4|20|In what place therefore ye hear the sound of the trumpet, resort ye thither unto us: our God shall fight for us.
NEH|4|21|So we laboured in the work: and half of them held the spears from the rising of the morning till the stars appeared.
NEH|4|22|Likewise at the same time said I unto the people, Let every one with his servant lodge within Jerusalem, that in the night they may be a guard to us, and labour on the day.
NEH|4|23|So neither I, nor my brethren, nor my servants, nor the men of the guard which followed me, none of us put off our clothes, saving that every one put them off for washing.
NEH|5|1|And there was a great cry of the people and of their wives against their brethren the Jews.
NEH|5|2|For there were that said, We, our sons, and our daughters, are many: therefore we take up corn for them, that we may eat, and live.
NEH|5|3|Some also there were that said, We have mortgaged our lands, vineyards, and houses, that we might buy corn, because of the dearth.
NEH|5|4|There were also that said, We have borrowed money for the king's tribute, and that upon our lands and vineyards.
NEH|5|5|Yet now our flesh is as the flesh of our brethren, our children as their children: and, lo, we bring into bondage our sons and our daughters to be servants, and some of our daughters are brought unto bondage already: neither is it in our power to redeem them; for other men have our lands and vineyards.
NEH|5|6|And I was very angry when I heard their cry and these words.
NEH|5|7|Then I consulted with myself, and I rebuked the nobles, and the rulers, and said unto them, Ye exact usury, every one of his brother. And I set a great assembly against them.
NEH|5|8|And I said unto them, We after our ability have redeemed our brethren the Jews, which were sold unto the heathen; and will ye even sell your brethren? or shall they be sold unto us? Then held they their peace, and found nothing to answer.
NEH|5|9|Also I said, It is not good that ye do: ought ye not to walk in the fear of our God because of the reproach of the heathen our enemies?
NEH|5|10|I likewise, and my brethren, and my servants, might exact of them money and corn: I pray you, let us leave off this usury.
NEH|5|11|Restore, I pray you, to them, even this day, their lands, their vineyards, their oliveyards, and their houses, also the hundredth part of the money, and of the corn, the wine, and the oil, that ye exact of them.
NEH|5|12|Then said they, We will restore them, and will require nothing of them; so will we do as thou sayest. Then I called the priests, and took an oath of them, that they should do according to this promise.
NEH|5|13|Also I shook my lap, and said, So God shake out every man from his house, and from his labour, that performeth not this promise, even thus be he shaken out, and emptied. And all the congregation said, Amen, and praised the LORD. And the people did according to this promise.
NEH|5|14|Moreover from the time that I was appointed to be their governor in the land of Judah, from the twentieth year even unto the two and thirtieth year of Artaxerxes the king, that is, twelve years, I and my brethren have not eaten the bread of the governor.
NEH|5|15|But the former governors that had been before me were chargeable unto the people, and had taken of them bread and wine, beside forty shekels of silver; yea, even their servants bare rule over the people: but so did not I, because of the fear of God.
NEH|5|16|Yea, also I continued in the work of this wall, neither bought we any land: and all my servants were gathered thither unto the work.
NEH|5|17|Moreover there were at my table an hundred and fifty of the Jews and rulers, beside those that came unto us from among the heathen that are about us.
NEH|5|18|Now that which was prepared for me daily was one ox and six choice sheep; also fowls were prepared for me, and once in ten days store of all sorts of wine: yet for all this required not I the bread of the governor, because the bondage was heavy upon this people.
NEH|5|19|Think upon me, my God, for good, according to all that I have done for this people.
NEH|6|1|Now it came to pass when Sanballat, and Tobiah, and Geshem the Arabian, and the rest of our enemies, heard that I had builded the wall, and that there was no breach left therein; (though at that time I had not set up the doors upon the gates;)
NEH|6|2|That Sanballat and Geshem sent unto me, saying, Come, let us meet together in some one of the villages in the plain of Ono. But they thought to do me mischief.
NEH|6|3|And I sent messengers unto them, saying, I am doing a great work, so that I cannot come down: why should the work cease, whilst I leave it, and come down to you?
NEH|6|4|Yet they sent unto me four times after this sort; and I answered them after the same manner.
NEH|6|5|Then sent Sanballat his servant unto me in like manner the fifth time with an open letter in his hand;
NEH|6|6|Wherein was written, It is reported among the heathen, and Gashmu saith it, that thou and the Jews think to rebel: for which cause thou buildest the wall, that thou mayest be their king, according to these words.
NEH|6|7|And thou hast also appointed prophets to preach of thee at Jerusalem, saying, There is a king in Judah: and now shall it be reported to the king according to these words. Come now therefore, and let us take counsel together.
NEH|6|8|Then I sent unto him, saying, There are no such things done as thou sayest, but thou feignest them out of thine own heart.
NEH|6|9|For they all made us afraid, saying, Their hands shall be weakened from the work, that it be not done. Now therefore, O God, strengthen my hands.
NEH|6|10|Afterward I came unto the house of Shemaiah the son of Delaiah the son of Mehetabeel, who was shut up; and he said, Let us meet together in the house of God, within the temple, and let us shut the doors of the temple: for they will come to slay thee; yea, in the night will they come to slay thee.
NEH|6|11|And I said, Should such a man as I flee? and who is there, that, being as I am, would go into the temple to save his life? I will not go in.
NEH|6|12|And, lo, I perceived that God had not sent him; but that he pronounced this prophecy against me: for Tobiah and Sanballat had hired him.
NEH|6|13|Therefore was he hired, that I should be afraid, and do so, and sin, and that they might have matter for an evil report, that they might reproach me.
NEH|6|14|My God, think thou upon Tobiah and Sanballat according to these their works, and on the prophetess Noadiah, and the rest of the prophets, that would have put me in fear.
NEH|6|15|So the wall was finished in the twenty and fifth day of the month Elul, in fifty and two days.
NEH|6|16|And it came to pass, that when all our enemies heard thereof, and all the heathen that were about us saw these things, they were much cast down in their own eyes: for they perceived that this work was wrought of our God.
NEH|6|17|Moreover in those days the nobles of Judah sent many letters unto Tobiah, and the letters of Tobiah came unto them.
NEH|6|18|For there were many in Judah sworn unto him, because he was the son in law of Shechaniah the son of Arah; and his son Johanan had taken the daughter of Meshullam the son of Berechiah.
NEH|6|19|Also they reported his good deeds before me, and uttered my words to him. And Tobiah sent letters to put me in fear.
NEH|7|1|Now it came to pass, when the wall was built, and I had set up the doors, and the porters and the singers and the Levites were appointed,
NEH|7|2|That I gave my brother Hanani, and Hananiah the ruler of the palace, charge over Jerusalem: for he was a faithful man, and feared God above many.
NEH|7|3|And I said unto them, Let not the gates of Jerusalem be opened until the sun be hot; and while they stand by, let them shut the doors, and bar them: and appoint watches of the inhabitants of Jerusalem, every one in his watch, and every one to be over against his house.
NEH|7|4|Now the city was large and great: but the people were few therein, and the houses were not builded.
NEH|7|5|And my God put into mine heart to gather together the nobles, and the rulers, and the people, that they might be reckoned by genealogy. And I found a register of the genealogy of them which came up at the first, and found written therein,
NEH|7|6|These are the children of the province, that went up out of the captivity, of those that had been carried away, whom Nebuchadnezzar the king of Babylon had carried away, and came again to Jerusalem and to Judah, every one unto his city;
NEH|7|7|Who came with Zerubbabel, Jeshua, Nehemiah, Azariah, Raamiah, Nahamani, Mordecai, Bilshan, Mispereth, Bigvai, Nehum, Baanah. The number, I say, of the men of the people of Israel was this;
NEH|7|8|The children of Parosh, two thousand an hundred seventy and two.
NEH|7|9|The children of Shephatiah, three hundred seventy and two.
NEH|7|10|The children of Arah, six hundred fifty and two.
NEH|7|11|The children of Pahathmoab, of the children of Jeshua and Joab, two thousand and eight hundred and eighteen.
NEH|7|12|The children of Elam, a thousand two hundred fifty and four.
NEH|7|13|The children of Zattu, eight hundred forty and five.
NEH|7|14|The children of Zaccai, seven hundred and threescore.
NEH|7|15|The children of Binnui, six hundred forty and eight.
NEH|7|16|The children of Bebai, six hundred twenty and eight.
NEH|7|17|The children of Azgad, two thousand three hundred twenty and two.
NEH|7|18|The children of Adonikam, six hundred threescore and seven.
NEH|7|19|The children of Bigvai, two thousand threescore and seven.
NEH|7|20|The children of Adin, six hundred fifty and five.
NEH|7|21|The children of Ater of Hezekiah, ninety and eight.
NEH|7|22|The children of Hashum, three hundred twenty and eight.
NEH|7|23|The children of Bezai, three hundred twenty and four.
NEH|7|24|The children of Hariph, an hundred and twelve.
NEH|7|25|The children of Gibeon, ninety and five.
NEH|7|26|The men of Bethlehem and Netophah, an hundred fourscore and eight.
NEH|7|27|The men of Anathoth, an hundred twenty and eight.
NEH|7|28|The men of Bethazmaveth, forty and two.
NEH|7|29|The men of Kirjathjearim, Chephirah, and Beeroth, seven hundred forty and three.
NEH|7|30|The men of Ramah and Gaba, six hundred twenty and one.
NEH|7|31|The men of Michmas, an hundred and twenty and two.
NEH|7|32|The men of Bethel and Ai, an hundred twenty and three.
NEH|7|33|The men of the other Nebo, fifty and two.
NEH|7|34|The children of the other Elam, a thousand two hundred fifty and four.
NEH|7|35|The children of Harim, three hundred and twenty.
NEH|7|36|The children of Jericho, three hundred forty and five.
NEH|7|37|The children of Lod, Hadid, and Ono, seven hundred twenty and one.
NEH|7|38|The children of Senaah, three thousand nine hundred and thirty.
NEH|7|39|The priests: the children of Jedaiah, of the house of Jeshua, nine hundred seventy and three.
NEH|7|40|The children of Immer, a thousand fifty and two.
NEH|7|41|The children of Pashur, a thousand two hundred forty and seven.
NEH|7|42|The children of Harim, a thousand and seventeen.
NEH|7|43|The Levites: the children of Jeshua, of Kadmiel, and of the children of Hodevah, seventy and four.
NEH|7|44|The singers: the children of Asaph, an hundred forty and eight.
NEH|7|45|The porters: the children of Shallum, the children of Ater, the children of Talmon, the children of Akkub, the children of Hatita, the children of Shobai, an hundred thirty and eight.
NEH|7|46|The Nethinims: the children of Ziha, the children of Hashupha, the children of Tabbaoth,
NEH|7|47|The children of Keros, the children of Sia, the children of Padon,
NEH|7|48|The children of Lebana, the children of Hagaba, the children of Shalmai,
NEH|7|49|The children of Hanan, the children of Giddel, the children of Gahar,
NEH|7|50|The children of Reaiah, the children of Rezin, the children of Nekoda,
NEH|7|51|The children of Gazzam, the children of Uzza, the children of Phaseah,
NEH|7|52|The children of Besai, the children of Meunim, the children of Nephishesim,
NEH|7|53|The children of Bakbuk, the children of Hakupha, the children of Harhur,
NEH|7|54|The children of Bazlith, the children of Mehida, the children of Harsha,
NEH|7|55|The children of Barkos, the children of Sisera, the children of Tamah,
NEH|7|56|The children of Neziah, the children of Hatipha.
NEH|7|57|The children of Solomon's servants: the children of Sotai, the children of Sophereth, the children of Perida,
NEH|7|58|The children of Jaala, the children of Darkon, the children of Giddel,
NEH|7|59|The children of Shephatiah, the children of Hattil, the children of Pochereth of Zebaim, the children of Amon.
NEH|7|60|All the Nethinims, and the children of Solomon's servants, were three hundred ninety and two.
NEH|7|61|And these were they which went up also from Telmelah, Telharesha, Cherub, Addon, and Immer: but they could not shew their father's house, nor their seed, whether they were of Israel.
NEH|7|62|The children of Delaiah, the children of Tobiah, the children of Nekoda, six hundred forty and two.
NEH|7|63|And of the priests: the children of Habaiah, the children of Koz, the children of Barzillai, which took one of the daughters of Barzillai the Gileadite to wife, and was called after their name.
NEH|7|64|These sought their register among those that were reckoned by genealogy, but it was not found: therefore were they, as polluted, put from the priesthood.
NEH|7|65|And the Tirshatha said unto them, that they should not eat of the most holy things, till there stood up a priest with Urim and Thummim.
NEH|7|66|The whole congregation together was forty and two thousand three hundred and threescore,
NEH|7|67|Beside their manservants and their maidservants, of whom there were seven thousand three hundred thirty and seven: and they had two hundred forty and five singing men and singing women.
NEH|7|68|Their horses, seven hundred thirty and six: their mules, two hundred forty and five:
NEH|7|69|Their camels, four hundred thirty and five: six thousand seven hundred and twenty asses.
NEH|7|70|And some of the chief of the fathers gave unto the work. The Tirshatha gave to the treasure a thousand drams of gold, fifty basons, five hundred and thirty priests' garments.
NEH|7|71|And some of the chief of the fathers gave to the treasure of the work twenty thousand drams of gold, and two thousand and two hundred pound of silver.
NEH|7|72|And that which the rest of the people gave was twenty thousand drams of gold, and two thousand pound of silver, and threescore and seven priests' garments.
NEH|7|73|So the priests, and the Levites, and the porters, and the singers, and some of the people, and the Nethinims, and all Israel, dwelt in their cities; and when the seventh month came, the children of Israel were in their cities.
NEH|8|1|And all the people gathered themselves together as one man into the street that was before the water gate; and they spake unto Ezra the scribe to bring the book of the law of Moses, which the LORD had commanded to Israel.
NEH|8|2|And Ezra the priest brought the law before the congregation both of men and women, and all that could hear with understanding, upon the first day of the seventh month.
NEH|8|3|And he read therein before the street that was before the water gate from the morning until midday, before the men and the women, and those that could understand; and the ears of all the people were attentive unto the book of the law.
NEH|8|4|And Ezra the scribe stood upon a pulpit of wood, which they had made for the purpose; and beside him stood Mattithiah, and Shema, and Anaiah, and Urijah, and Hilkiah, and Maaseiah, on his right hand; and on his left hand, Pedaiah, and Mishael, and Malchiah, and Hashum, and Hashbadana, Zechariah, and Meshullam.
NEH|8|5|And Ezra opened the book in the sight of all the people; (for he was above all the people;) and when he opened it, all the people stood up:
NEH|8|6|And Ezra blessed the LORD, the great God. And all the people answered, Amen, Amen, with lifting up their hands: and they bowed their heads, and worshipped the LORD with their faces to the ground.
NEH|8|7|Also Jeshua, and Bani, and Sherebiah, Jamin, Akkub, Shabbethai, Hodijah, Maaseiah, Kelita, Azariah, Jozabad, Hanan, Pelaiah, and the Levites, caused the people to understand the law: and the people stood in their place.
NEH|8|8|So they read in the book in the law of God distinctly, and gave the sense, and caused them to understand the reading.
NEH|8|9|And Nehemiah, which is the Tirshatha, and Ezra the priest the scribe, and the Levites that taught the people, said unto all the people, This day is holy unto the LORD your God; mourn not, nor weep. For all the people wept, when they heard the words of the law.
NEH|8|10|Then he said unto them, Go your way, eat the fat, and drink the sweet, and send portions unto them for whom nothing is prepared: for this day is holy unto our LORD: neither be ye sorry; for the joy of the LORD is your strength.
NEH|8|11|So the Levites stilled all the people, saying, Hold your peace, for the day is holy; neither be ye grieved.
NEH|8|12|And all the people went their way to eat, and to drink, and to send portions, and to make great mirth, because they had understood the words that were declared unto them.
NEH|8|13|And on the second day were gathered together the chief of the fathers of all the people, the priests, and the Levites, unto Ezra the scribe, even to understand the words of the law.
NEH|8|14|And they found written in the law which the LORD had commanded by Moses, that the children of Israel should dwell in booths in the feast of the seventh month:
NEH|8|15|And that they should publish and proclaim in all their cities, and in Jerusalem, saying, Go forth unto the mount, and fetch olive branches, and pine branches, and myrtle branches, and palm branches, and branches of thick trees, to make booths, as it is written.
NEH|8|16|So the people went forth, and brought them, and made themselves booths, every one upon the roof of his house, and in their courts, and in the courts of the house of God, and in the street of the water gate, and in the street of the gate of Ephraim.
NEH|8|17|And all the congregation of them that were come again out of the captivity made booths, and sat under the booths: for since the days of Jeshua the son of Nun unto that day had not the children of Israel done so. And there was very great gladness.
NEH|8|18|Also day by day, from the first day unto the last day, he read in the book of the law of God. And they kept the feast seven days; and on the eighth day was a solemn assembly, according unto the manner.
NEH|9|1|Now in the twenty and fourth day of this month the children of Israel were assembled with fasting, and with sackclothes, and earth upon them.
NEH|9|2|And the seed of Israel separated themselves from all strangers, and stood and confessed their sins, and the iniquities of their fathers.
NEH|9|3|And they stood up in their place, and read in the book of the law of the LORD their God one fourth part of the day; and another fourth part they confessed, and worshipped the LORD their God.
NEH|9|4|Then stood up upon the stairs, of the Levites, Jeshua, and Bani, Kadmiel, Shebaniah, Bunni, Sherebiah, Bani, and Chenani, and cried with a loud voice unto the LORD their God.
NEH|9|5|Then the Levites, Jeshua, and Kadmiel, Bani, Hashabniah, Sherebiah, Hodijah, Shebaniah, and Pethahiah, said, Stand up and bless the LORD your God for ever and ever: and blessed be thy glorious name, which is exalted above all blessing and praise.
NEH|9|6|Thou, even thou, art LORD alone; thou hast made heaven, the heaven of heavens, with all their host, the earth, and all things that are therein, the seas, and all that is therein, and thou preservest them all; and the host of heaven worshippeth thee.
NEH|9|7|Thou art the LORD the God, who didst choose Abram, and broughtest him forth out of Ur of the Chaldees, and gavest him the name of Abraham;
NEH|9|8|And foundest his heart faithful before thee, and madest a covenant with him to give the land of the Canaanites, the Hittites, the Amorites, and the Perizzites, and the Jebusites, and the Girgashites, to give it, I say, to his seed, and hast performed thy words; for thou art righteous:
NEH|9|9|And didst see the affliction of our fathers in Egypt, and heardest their cry by the Red sea;
NEH|9|10|And shewedst signs and wonders upon Pharaoh, and on all his servants, and on all the people of his land: for thou knewest that they dealt proudly against them. So didst thou get thee a name, as it is this day.
NEH|9|11|And thou didst divide the sea before them, so that they went through the midst of the sea on the dry land; and their persecutors thou threwest into the deeps, as a stone into the mighty waters.
NEH|9|12|Moreover thou leddest them in the day by a cloudy pillar; and in the night by a pillar of fire, to give them light in the way wherein they should go.
NEH|9|13|Thou camest down also upon mount Sinai, and spakest with them from heaven, and gavest them right judgments, and true laws, good statutes and commandments:
NEH|9|14|And madest known unto them thy holy sabbath, and commandedst them precepts, statutes, and laws, by the hand of Moses thy servant:
NEH|9|15|And gavest them bread from heaven for their hunger, and broughtest forth water for them out of the rock for their thirst, and promisedst them that they should go in to possess the land which thou hadst sworn to give them.
NEH|9|16|But they and our fathers dealt proudly, and hardened their necks, and hearkened not to thy commandments,
NEH|9|17|And refused to obey, neither were mindful of thy wonders that thou didst among them; but hardened their necks, and in their rebellion appointed a captain to return to their bondage: but thou art a God ready to pardon, gracious and merciful, slow to anger, and of great kindness, and forsookest them not.
NEH|9|18|Yea, when they had made them a molten calf, and said, This is thy God that brought thee up out of Egypt, and had wrought great provocations;
NEH|9|19|Yet thou in thy manifold mercies forsookest them not in the wilderness: the pillar of the cloud departed not from them by day, to lead them in the way; neither the pillar of fire by night, to shew them light, and the way wherein they should go.
NEH|9|20|Thou gavest also thy good spirit to instruct them, and withheldest not thy manna from their mouth, and gavest them water for their thirst.
NEH|9|21|Yea, forty years didst thou sustain them in the wilderness, so that they lacked nothing; their clothes waxed not old, and their feet swelled not.
NEH|9|22|Moreover thou gavest them kingdoms and nations, and didst divide them into corners: so they possessed the land of Sihon, and the land of the king of Heshbon, and the land of Og king of Bashan.
NEH|9|23|Their children also multipliedst thou as the stars of heaven, and broughtest them into the land, concerning which thou hadst promised to their fathers, that they should go in to possess it.
NEH|9|24|So the children went in and possessed the land, and thou subduedst before them the inhabitants of the land, the Canaanites, and gavest them into their hands, with their kings, and the people of the land, that they might do with them as they would.
NEH|9|25|And they took strong cities, and a fat land, and possessed houses full of all goods, wells digged, vineyards, and oliveyards, and fruit trees in abundance: so they did eat, and were filled, and became fat, and delighted themselves in thy great goodness.
NEH|9|26|Nevertheless they were disobedient, and rebelled against thee, and cast thy law behind their backs, and slew thy prophets which testified against them to turn them to thee, and they wrought great provocations.
NEH|9|27|Therefore thou deliveredst them into the hand of their enemies, who vexed them: and in the time of their trouble, when they cried unto thee, thou heardest them from heaven; and according to thy manifold mercies thou gavest them saviours, who saved them out of the hand of their enemies.
NEH|9|28|But after they had rest, they did evil again before thee: therefore leftest thou them in the land of their enemies, so that they had the dominion over them: yet when they returned, and cried unto thee, thou heardest them from heaven; and many times didst thou deliver them according to thy mercies;
NEH|9|29|And testifiedst against them, that thou mightest bring them again unto thy law: yet they dealt proudly, and hearkened not unto thy commandments, but sinned against thy judgments, (which if a man do, he shall live in them;) and withdrew the shoulder, and hardened their neck, and would not hear.
NEH|9|30|Yet many years didst thou forbear them, and testifiedst against them by thy spirit in thy prophets: yet would they not give ear: therefore gavest thou them into the hand of the people of the lands.
NEH|9|31|Nevertheless for thy great mercies' sake thou didst not utterly consume them, nor forsake them; for thou art a gracious and merciful God.
NEH|9|32|Now therefore, our God, the great, the mighty, and the terrible God, who keepest covenant and mercy, let not all the trouble seem little before thee, that hath come upon us, on our kings, on our princes, and on our priests, and on our prophets, and on our fathers, and on all thy people, since the time of the kings of Assyria unto this day.
NEH|9|33|Howbeit thou art just in all that is brought upon us; for thou hast done right, but we have done wickedly:
NEH|9|34|Neither have our kings, our princes, our priests, nor our fathers, kept thy law, nor hearkened unto thy commandments and thy testimonies, wherewith thou didst testify against them.
NEH|9|35|For they have not served thee in their kingdom, and in thy great goodness that thou gavest them, and in the large and fat land which thou gavest before them, neither turned they from their wicked works.
NEH|9|36|Behold, we are servants this day, and for the land that thou gavest unto our fathers to eat the fruit thereof and the good thereof, behold, we are servants in it:
NEH|9|37|And it yieldeth much increase unto the kings whom thou hast set over us because of our sins: also they have dominion over our bodies, and over our cattle, at their pleasure, and we are in great distress.
NEH|9|38|And because of all this we make a sure covenant, and write it; and our princes, Levites, and priests, seal unto it.
NEH|10|1|Now those that sealed were, Nehemiah, the Tirshatha, the son of Hachaliah, and Zidkijah,
NEH|10|2|Seraiah, Azariah, Jeremiah,
NEH|10|3|Pashur, Amariah, Malchijah,
NEH|10|4|Hattush, Shebaniah, Malluch,
NEH|10|5|Harim, Meremoth, Obadiah,
NEH|10|6|Daniel, Ginnethon, Baruch,
NEH|10|7|Meshullam, Abijah, Mijamin,
NEH|10|8|Maaziah, Bilgai, Shemaiah: these were the priests.
NEH|10|9|And the Levites: both Jeshua the son of Azaniah, Binnui of the sons of Henadad, Kadmiel;
NEH|10|10|And their brethren, Shebaniah, Hodijah, Kelita, Pelaiah, Hanan,
NEH|10|11|Micha, Rehob, Hashabiah,
NEH|10|12|Zaccur, Sherebiah, Shebaniah,
NEH|10|13|Hodijah, Bani, Beninu.
NEH|10|14|The chief of the people; Parosh, Pahathmoab, Elam, Zatthu, Bani,
NEH|10|15|Bunni, Azgad, Bebai,
NEH|10|16|Adonijah, Bigvai, Adin,
NEH|10|17|Ater, Hizkijah, Azzur,
NEH|10|18|Hodijah, Hashum, Bezai,
NEH|10|19|Hariph, Anathoth, Nebai,
NEH|10|20|Magpiash, Meshullam, Hezir,
NEH|10|21|Meshezabeel, Zadok, Jaddua,
NEH|10|22|Pelatiah, Hanan, Anaiah,
NEH|10|23|Hoshea, Hananiah, Hashub,
NEH|10|24|Hallohesh, Pileha, Shobek,
NEH|10|25|Rehum, Hashabnah, Maaseiah,
NEH|10|26|And Ahijah, Hanan, Anan,
NEH|10|27|Malluch, Harim, Baanah.
NEH|10|28|And the rest of the people, the priests, the Levites, the porters, the singers, the Nethinims, and all they that had separated themselves from the people of the lands unto the law of God, their wives, their sons, and their daughters, every one having knowledge, and having understanding;
NEH|10|29|They clave to their brethren, their nobles, and entered into a curse, and into an oath, to walk in God's law, which was given by Moses the servant of God, and to observe and do all the commandments of the LORD our Lord, and his judgments and his statutes;
NEH|10|30|And that we would not give our daughters unto the people of the land, not take their daughters for our sons:
NEH|10|31|And if the people of the land bring ware or any victuals on the sabbath day to sell, that we would not buy it of them on the sabbath, or on the holy day: and that we would leave the seventh year, and the exaction of every debt.
NEH|10|32|Also we made ordinances for us, to charge ourselves yearly with the third part of a shekel for the service of the house of our God;
NEH|10|33|For the shewbread, and for the continual meat offering, and for the continual burnt offering, of the sabbaths, of the new moons, for the set feasts, and for the holy things, and for the sin offerings to make an atonement for Israel, and for all the work of the house of our God.
NEH|10|34|And we cast the lots among the priests, the Levites, and the people, for the wood offering, to bring it into the house of our God, after the houses of our fathers, at times appointed year by year, to burn upon the altar of the LORD our God, as it is written in the law:
NEH|10|35|And to bring the firstfruits of our ground, and the firstfruits of all fruit of all trees, year by year, unto the house of the LORD:
NEH|10|36|Also the firstborn of our sons, and of our cattle, as it is written in the law, and the firstlings of our herds and of our flocks, to bring to the house of our God, unto the priests that minister in the house of our God:
NEH|10|37|And that we should bring the firstfruits of our dough, and our offerings, and the fruit of all manner of trees, of wine and of oil, unto the priests, to the chambers of the house of our God; and the tithes of our ground unto the Levites, that the same Levites might have the tithes in all the cities of our tillage.
NEH|10|38|And the priest the son of Aaron shall be with the Levites, when the Levites take tithes: and the Levites shall bring up the tithe of the tithes unto the house of our God, to the chambers, into the treasure house.
NEH|10|39|For the children of Israel and the children of Levi shall bring the offering of the corn, of the new wine, and the oil, unto the chambers, where are the vessels of the sanctuary, and the priests that minister, and the porters, and the singers: and we will not forsake the house of our God.
NEH|11|1|And the rulers of the people dwelt at Jerusalem: the rest of the people also cast lots, to bring one of ten to dwell in Jerusalem the holy city, and nine parts to dwell in other cities.
NEH|11|2|And the people blessed all the men, that willingly offered themselves to dwell at Jerusalem.
NEH|11|3|Now these are the chief of the province that dwelt in Jerusalem: but in the cities of Judah dwelt every one in his possession in their cities, to wit, Israel, the priests, and the Levites, and the Nethinims, and the children of Solomon's servants.
NEH|11|4|And at Jerusalem dwelt certain of the children of Judah, and of the children of Benjamin. Of the children of Judah; Athaiah the son of Uzziah, the son of Zechariah, the son of Amariah, the son of Shephatiah, the son of Mahalaleel, of the children of Perez;
NEH|11|5|And Maaseiah the son of Baruch, the son of Colhozeh, the son of Hazaiah, the son of Adaiah, the son of Joiarib, the son of Zechariah, the son of Shiloni.
NEH|11|6|All the sons of Perez that dwelt at Jerusalem were four hundred threescore and eight valiant men.
NEH|11|7|And these are the sons of Benjamin; Sallu the son of Meshullam, the son of Joed, the son of Pedaiah, the son of Kolaiah, the son of Maaseiah, the son of Ithiel, the son of Jesaiah.
NEH|11|8|And after him Gabbai, Sallai, nine hundred twenty and eight.
NEH|11|9|And Joel the son of Zichri was their overseer: and Judah the son of Senuah was second over the city.
NEH|11|10|Of the priests: Jedaiah the son of Joiarib, Jachin.
NEH|11|11|Seraiah the son of Hilkiah, the son of Meshullam, the son of Zadok, the son of Meraioth, the son of Ahitub, was the ruler of the house of God.
NEH|11|12|And their brethren that did the work of the house were eight hundred twenty and two: and Adaiah the son of Jeroham, the son of Pelaliah, the son of Amzi, the son of Zechariah, the son of Pashur, the son of Malchiah.
NEH|11|13|And his brethren, chief of the fathers, two hundred forty and two: and Amashai the son of Azareel, the son of Ahasai, the son of Meshillemoth, the son of Immer,
NEH|11|14|And their brethren, mighty men of valour, an hundred twenty and eight: and their overseer was Zabdiel, the son of one of the great men.
NEH|11|15|Also of the Levites: Shemaiah the son of Hashub, the son of Azrikam, the son of Hashabiah, the son of Bunni;
NEH|11|16|And Shabbethai and Jozabad, of the chief of the Levites, had the oversight of the outward business of the house of God.
NEH|11|17|And Mattaniah the son of Micha, the son of Zabdi, the son of Asaph, was the principal to begin the thanksgiving in prayer: and Bakbukiah the second among his brethren, and Abda the son of Shammua, the son of Galal, the son of Jeduthun.
NEH|11|18|All the Levites in the holy city were two hundred fourscore and four.
NEH|11|19|Moreover the porters, Akkub, Talmon, and their brethren that kept the gates, were an hundred seventy and two.
NEH|11|20|And the residue of Israel, of the priests, and the Levites, were in all the cities of Judah, every one in his inheritance.
NEH|11|21|But the Nethinims dwelt in Ophel: and Ziha and Gispa were over the Nethinims.
NEH|11|22|The overseer also of the Levites at Jerusalem was Uzzi the son of Bani, the son of Hashabiah, the son of Mattaniah, the son of Micha. Of the sons of Asaph, the singers were over the business of the house of God.
NEH|11|23|For it was the king's commandment concerning them, that a certain portion should be for the singers, due for every day.
NEH|11|24|And Pethahiah the son of Meshezabeel, of the children of Zerah the son of Judah, was at the king's hand in all matters concerning the people.
NEH|11|25|And for the villages, with their fields, some of the children of Judah dwelt at Kirjatharba, and in the villages thereof, and at Dibon, and in the villages thereof, and at Jekabzeel, and in the villages thereof,
NEH|11|26|And at Jeshua, and at Moladah, and at Bethphelet,
NEH|11|27|And at Hazarshual, and at Beersheba, and in the villages thereof,
NEH|11|28|And at Ziklag, and at Mekonah, and in the villages thereof,
NEH|11|29|And at Enrimmon, and at Zareah, and at Jarmuth,
NEH|11|30|Zanoah, Adullam, and in their villages, at Lachish, and the fields thereof, at Azekah, and in the villages thereof. And they dwelt from Beersheba unto the valley of Hinnom.
NEH|11|31|The children also of Benjamin from Geba dwelt at Michmash, and Aija, and Bethel, and in their villages.
NEH|11|32|And at Anathoth, Nob, Ananiah,
NEH|11|33|Hazor, Ramah, Gittaim,
NEH|11|34|Hadid, Zeboim, Neballat,
NEH|11|35|Lod, and Ono, the valley of craftsmen.
NEH|11|36|And of the Levites were divisions in Judah, and in Benjamin.
NEH|12|1|Now these are the priests and the Levites that went up with Zerubbabel the son of Shealtiel, and Jeshua: Seraiah, Jeremiah, Ezra,
NEH|12|2|Amariah, Malluch, Hattush,
NEH|12|3|Shechaniah, Rehum, Meremoth,
NEH|12|4|Iddo, Ginnetho, Abijah,
NEH|12|5|Miamin, Maadiah, Bilgah,
NEH|12|6|Shemaiah, and Joiarib, Jedaiah,
NEH|12|7|Sallu, Amok, Hilkiah, Jedaiah. These were the chief of the priests and of their brethren in the days of Jeshua.
NEH|12|8|Moreover the Levites: Jeshua, Binnui, Kadmiel, Sherebiah, Judah, and Mattaniah, which was over the thanksgiving, he and his brethren.
NEH|12|9|Also Bakbukiah and Unni, their brethren, were over against them in the watches.
NEH|12|10|And Jeshua begat Joiakim, Joiakim also begat Eliashib, and Eliashib begat Joiada,
NEH|12|11|And Joiada begat Jonathan, and Jonathan begat Jaddua.
NEH|12|12|And in the days of Joiakim were priests, the chief of the fathers: of Seraiah, Meraiah; of Jeremiah, Hananiah;
NEH|12|13|Of Ezra, Meshullam; of Amariah, Jehohanan;
NEH|12|14|Of Melicu, Jonathan; of Shebaniah, Joseph;
NEH|12|15|Of Harim, Adna; of Meraioth, Helkai;
NEH|12|16|Of Iddo, Zechariah; of Ginnethon, Meshullam;
NEH|12|17|Of Abijah, Zichri; of Miniamin, of Moadiah, Piltai:
NEH|12|18|Of Bilgah, Shammua; of Shemaiah, Jehonathan;
NEH|12|19|And of Joiarib, Mattenai; of Jedaiah, Uzzi;
NEH|12|20|Of Sallai, Kallai; of Amok, Eber;
NEH|12|21|Of Hilkiah, Hashabiah; of Jedaiah, Nethaneel.
NEH|12|22|The Levites in the days of Eliashib, Joiada, and Johanan, and Jaddua, were recorded chief of the fathers: also the priests, to the reign of Darius the Persian.
NEH|12|23|The sons of Levi, the chief of the fathers, were written in the book of the chronicles, even until the days of Johanan the son of Eliashib.
NEH|12|24|And the chief of the Levites: Hashabiah, Sherebiah, and Jeshua the son of Kadmiel, with their brethren over against them, to praise and to give thanks, according to the commandment of David the man of God, ward over against ward.
NEH|12|25|Mattaniah, and Bakbukiah, Obadiah, Meshullam, Talmon, Akkub, were porters keeping the ward at the thresholds of the gates.
NEH|12|26|These were in the days of Joiakim the son of Jeshua, the son of Jozadak, and in the days of Nehemiah the governor, and of Ezra the priest, the scribe.
NEH|12|27|And at the dedication of the wall of Jerusalem they sought the Levites out of all their places, to bring them to Jerusalem, to keep the dedication with gladness, both with thanksgivings, and with singing, with cymbals, psalteries, and with harps.
NEH|12|28|And the sons of the singers gathered themselves together, both out of the plain country round about Jerusalem, and from the villages of Netophathi;
NEH|12|29|Also from the house of Gilgal, and out of the fields of Geba and Azmaveth: for the singers had builded them villages round about Jerusalem.
NEH|12|30|And the priests and the Levites purified themselves, and purified the people, and the gates, and the wall.
NEH|12|31|Then I brought up the princes of Judah upon the wall, and appointed two great companies of them that gave thanks, whereof one went on the right hand upon the wall toward the dung gate:
NEH|12|32|And after them went Hoshaiah, and half of the princes of Judah,
NEH|12|33|And Azariah, Ezra, and Meshullam,
NEH|12|34|Judah, and Benjamin, and Shemaiah, and Jeremiah,
NEH|12|35|And certain of the priests' sons with trumpets; namely, Zechariah the son of Jonathan, the son of Shemaiah, the son of Mattaniah, the son of Michaiah, the son of Zaccur, the son of Asaph:
NEH|12|36|And his brethren, Shemaiah, and Azarael, Milalai, Gilalai, Maai, Nethaneel, and Judah, Hanani, with the musical instruments of David the man of God, and Ezra the scribe before them.
NEH|12|37|And at the fountain gate, which was over against them, they went up by the stairs of the city of David, at the going up of the wall, above the house of David, even unto the water gate eastward.
NEH|12|38|And the other company of them that gave thanks went over against them, and I after them, and the half of the people upon the wall, from beyond the tower of the furnaces even unto the broad wall;
NEH|12|39|And from above the gate of Ephraim, and above the old gate, and above the fish gate, and the tower of Hananeel, and the tower of Meah, even unto the sheep gate: and they stood still in the prison gate.
NEH|12|40|So stood the two companies of them that gave thanks in the house of God, and I, and the half of the rulers with me:
NEH|12|41|And the priests; Eliakim, Maaseiah, Miniamin, Michaiah, Elioenai, Zechariah, and Hananiah, with trumpets;
NEH|12|42|And Maaseiah, and Shemaiah, and Eleazar, and Uzzi, and Jehohanan, and Malchijah, and Elam, and Ezer. And the singers sang loud, with Jezrahiah their overseer.
NEH|12|43|Also that day they offered great sacrifices, and rejoiced: for God had made them rejoice with great joy: the wives also and the children rejoiced: so that the joy of Jerusalem was heard even afar off.
NEH|12|44|And at that time were some appointed over the chambers for the treasures, for the offerings, for the firstfruits, and for the tithes, to gather into them out of the fields of the cities the portions of the law for the priests and Levites: for Judah rejoiced for the priests and for the Levites that waited.
NEH|12|45|And both the singers and the porters kept the ward of their God, and the ward of the purification, according to the commandment of David, and of Solomon his son.
NEH|12|46|For in the days of David and Asaph of old there were chief of the singers, and songs of praise and thanksgiving unto God.
NEH|12|47|And all Israel in the days of Zerubbabel, and in the days of Nehemiah, gave the portions of the singers and the porters, every day his portion: and they sanctified holy things unto the Levites; and the Levites sanctified them unto the children of Aaron.
NEH|13|1|On that day they read in the book of Moses in the audience of the people; and therein was found written, that the Ammonite and the Moabite should not come into the congregation of God for ever;
NEH|13|2|Because they met not the children of Israel with bread and with water, but hired Balaam against them, that he should curse them: howbeit our God turned the curse into a blessing.
NEH|13|3|Now it came to pass, when they had heard the law, that they separated from Israel all the mixed multitude.
NEH|13|4|And before this, Eliashib the priest, having the oversight of the chamber of the house of our God, was allied unto Tobiah:
NEH|13|5|And he had prepared for him a great chamber, where aforetime they laid the meat offerings, the frankincense, and the vessels, and the tithes of the corn, the new wine, and the oil, which was commanded to be given to the Levites, and the singers, and the porters; and the offerings of the priests.
NEH|13|6|But in all this time was not I at Jerusalem: for in the two and thirtieth year of Artaxerxes king of Babylon came I unto the king, and after certain days obtained I leave of the king:
NEH|13|7|And I came to Jerusalem, and understood of the evil that Eliashib did for Tobiah, in preparing him a chamber in the courts of the house of God.
NEH|13|8|And it grieved me sore: therefore I cast forth all the household stuff to Tobiah out of the chamber.
NEH|13|9|Then I commanded, and they cleansed the chambers: and thither brought I again the vessels of the house of God, with the meat offering and the frankincense.
NEH|13|10|And I perceived that the portions of the Levites had not been given them: for the Levites and the singers, that did the work, were fled every one to his field.
NEH|13|11|Then contended I with the rulers, and said, Why is the house of God forsaken? And I gathered them together, and set them in their place.
NEH|13|12|Then brought all Judah the tithe of the corn and the new wine and the oil unto the treasuries.
NEH|13|13|And I made treasurers over the treasuries, Shelemiah the priest, and Zadok the scribe, and of the Levites, Pedaiah: and next to them was Hanan the son of Zaccur, the son of Mattaniah: for they were counted faithful, and their office was to distribute unto their brethren.
NEH|13|14|Remember me, O my God, concerning this, and wipe not out my good deeds that I have done for the house of my God, and for the offices thereof.
NEH|13|15|In those days saw I in Judah some treading wine presses on the sabbath, and bringing in sheaves, and lading asses; as also wine, grapes, and figs, and all manner of burdens, which they brought into Jerusalem on the sabbath day: and I testified against them in the day wherein they sold victuals.
NEH|13|16|There dwelt men of Tyre also therein, which brought fish, and all manner of ware, and sold on the sabbath unto the children of Judah, and in Jerusalem.
NEH|13|17|Then I contended with the nobles of Judah, and said unto them, What evil thing is this that ye do, and profane the sabbath day?
NEH|13|18|Did not your fathers thus, and did not our God bring all this evil upon us, and upon this city? yet ye bring more wrath upon Israel by profaning the sabbath.
NEH|13|19|And it came to pass, that when the gates of Jerusalem began to be dark before the sabbath, I commanded that the gates should be shut, and charged that they should not be opened till after the sabbath: and some of my servants set I at the gates, that there should no burden be brought in on the sabbath day.
NEH|13|20|So the merchants and sellers of all kind of ware lodged without Jerusalem once or twice.
NEH|13|21|Then I testified against them, and said unto them, Why lodge ye about the wall? if ye do so again, I will lay hands on you. From that time forth came they no more on the sabbath.
NEH|13|22|And I commanded the Levites that they should cleanse themselves, and that they should come and keep the gates, to sanctify the sabbath day. Remember me, O my God, concerning this also, and spare me according to the greatness of thy mercy.
NEH|13|23|In those days also saw I Jews that had married wives of Ashdod, of Ammon, and of Moab:
NEH|13|24|And their children spake half in the speech of Ashdod, and could not speak in the Jews' language, but according to the language of each people.
NEH|13|25|And I contended with them, and cursed them, and smote certain of them, and plucked off their hair, and made them swear by God, saying, Ye shall not give your daughters unto their sons, nor take their daughters unto your sons, or for yourselves.
NEH|13|26|Did not Solomon king of Israel sin by these things? yet among many nations was there no king like him, who was beloved of his God, and God made him king over all Israel: nevertheless even him did outlandish women cause to sin.
NEH|13|27|Shall we then hearken unto you to do all this great evil, to transgress against our God in marrying strange wives?
NEH|13|28|And one of the sons of Joiada, the son of Eliashib the high priest, was son in law to Sanballat the Horonite: therefore I chased him from me.
NEH|13|29|Remember them, O my God, because they have defiled the priesthood, and the covenant of the priesthood, and of the Levites.
NEH|13|30|Thus cleansed I them from all strangers, and appointed the wards of the priests and the Levites, every one in his business;
NEH|13|31|And for the wood offering, at times appointed, and for the firstfruits. Remember me, O my God, for good.
