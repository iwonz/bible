JOSH|1|1|Et factum est, ut post mortem Moysi servi Domini loqueretur Dominus ad Iosue filium Nun ministrum Moysi et diceret ei:
JOSH|1|2|" Moyses servus meus mortuus est; nunc igitur surge et transi Iordanem istum, tu et omnis populus iste, in terram, quam ego dabo filiis Israel.
JOSH|1|3|Omnem locum, quem calcaverit vestigium pedis vestri, vobis tradidi, sicut locutus sum Moysi.
JOSH|1|4|A deserto et Libano isto usque ad fluvium magnum Euphraten, omnis terra Hetthaeorum usque ad mare Magnum contra solis occasum erit terminus vester.
JOSH|1|5|Nullus tibi poterit resistere cunctis diebus vitae tuae: sicut fui cum Moyse, ero et tecum; non dimittam nec derelinquam te.
JOSH|1|6|Confortare et esto robustus; tu enim sorte divides populo huic terram, pro qua iuravi patribus suis, ut traderem eam illis.
JOSH|1|7|Confortare tantum et esto robustus valde, ut custodias et facias iuxta omnem legem, quam praecepit tibi Moyses servus meus. Ne declines ab ea ad dexteram vel ad sinistram, ut prospereris in omnibus, ad quaecumque perrexeris.
JOSH|1|8|Non recedat hoc volumen legis de ore tuo, sed meditaberis in eo diebus ac noctibus, ut custodias et facias iuxta omnia, quae scripta sunt in eo: tunc optime diriges viam tuam et tunc prosperaberis.
JOSH|1|9|Nonne praecepi tibi: Confortare et esto robustus, noli metuere et noli timere, quoniam tecum est Dominus Deus tuus in omnibus, ad quaecumque perrexeris?".
JOSH|1|10|Praecepitque Iosue praefectis populi dicens: " Transite per medium castrorum et imperate populo ac dicite:
JOSH|1|11|Praeparate vobis cibaria, quoniam post diem tertium transibitis Iordanem hunc et intrabitis ad possidendam terram, quam Dominus Deus vester daturus est vobis ".
JOSH|1|12|Rubenitis quoque et Gaditis et dimidiae tribui Manasse ait:
JOSH|1|13|" Mementote sermonis, quem praecepit vobis Moyses famulus Domini dicens: "Dominus Deus vester dedit vobis requiem et terram hanc".
JOSH|1|14|Uxores vestrae et filii ac iumenta manebunt in terra, quam tradidit vobis Moyses trans Iordanem; vos autem transibitis armati ante fratres vestros, omnes viri fortes, et adiuvabitis eos,
JOSH|1|15|donec det requiem Dominus fratribus vestris, sicut et vobis dedit, et possideant ipsi quoque terram, quam Dominus Deus vester daturus est eis. Et sic revertemini in terram possessionis vestrae et habitabitis in ea, quam vobis dedit Moyses famulus Domini trans Iordanem contra solis ortum.
JOSH|1|16|Responderuntque ad Iosue atque dixerunt: " Omnia, quae praecepisti nobis, faciemus et, quocumque miseris, ibimus.
JOSH|1|17|Sicut oboedivimus in cunctis Moysi, ita oboediemus et tibi; tantum sit Dominus Deus tuus tecum, sicut fuit cum Moyse.
JOSH|1|18|Quicumque contradixerit ori tuo et non oboedierit cunctis sermonibus, quos praeceperis ei, moriatur; tu tantum confortare et viriliter age ".
JOSH|2|1|Misit ergo Iosue filius Nun de Settim duos viros exploratores in abscondito et dixit eis; "Ite et considerate terram urbemque Iericho ". Qui pergentes ingressi sunt domum mulieris meretricis nomine Rahab et quieverunt ibi.
JOSH|2|2|Nuntiatumque est regi Iericho et dictum: " Ecce viri ingressi sunt huc per noctem de filiis Israel, ut explorarent terram ".
JOSH|2|3|Misitque rex Iericho ad Rahab dicens: " Educ viros, qui venerunt ad te et ingressi sunt domum tuam; exploratores quippe sunt et omnem terram considerare venerunt ".
JOSH|2|4|Tollensque mulier viros abscondit et ait: " Fateor, venerunt ad me, sed nesciebam unde essent;
JOSH|2|5|cumque porta clauderetur in tenebris, et illi pariter exierunt, nescio quo abierunt. Persequimini cito et comprehendetis eos ".
JOSH|2|6|Ipsa autem fecit ascendere viros in solarium domus suae operuitque eos lini stipula, quae ibi erat.
JOSH|2|7|Hi autem, qui missi fuerant, secuti sunt eos per viam, quae ducit ad vadum Iordanis; illisque egressis, statim porta clausa est.
JOSH|2|8|Necdum obdormierant qui latebant, et ecce mulier ascendit ad eos et ait:
JOSH|2|9|" Novi quod tradiderit Dominus vobis terram, et irruit in nos terror vester, et elanguerunt omnes habitatores terrae coram vobis.
JOSH|2|10|Audivimus enim quod siccaverit Dominus aquas maris Rubri ad vestrum introitum, quando egressi estis ex Aegypto, et quae feceritis duobus Amorraeorum regibus, qui erant trans Iordanem, Sehon et Og, quos interfecistis.
JOSH|2|11|Et haec audientes pertimuimus, et elanguit cor nostrum, nec remansit in nobis spiritus ad introitum vestrum; Dominus enim Deus vester ipse est Deus in caelo sursum et in terra deorsum.
JOSH|2|12|Nunc ergo iurate mihi per Dominum, ut, quomodo ego feci vobiscum misericordiam, ita et vos faciatis cum domo patris mei detisque mihi signum verum,
JOSH|2|13|ut salvetis patrem meum et matrem, fratres ac sorores meas et omnia, quae eorum sunt, et eruatis animas nostras de morte ".
JOSH|2|14|Qui responderunt ei: " Anima nostra sit pro vobis in mortem, si tamen non prodideris; cumque tradiderit nobis Dominus terram, faciemus in te misericordiam et veritatem ".
JOSH|2|15|Demisit ergo eos per funem de fenestra; domus enim eius haerebat muro, et in muro habitabat.
JOSH|2|16|Dixitque ad eos: " Ad montana pergite, ne forte occurrant vobis persecutores, ibique latete diebus tribus, donec redeant; et postea ibitis per viam vestram.
JOSH|2|17|Qui dixerunt ad eam: " Innoxii erimus a iuramento hoc, quo adiurasti nos,
JOSH|2|18|si, ingredientibus nobis terram, signum fuerit funiculus iste coccineus, et ligaveris eum in fenestra, per quam nos demisisti, et patrem tuum ac matrem fratresque et omnem cognationem tuam congregaveris in domum tuam.
JOSH|2|19|Qui ostium domus tuae egressus fuerit, sanguis ipsius erit in caput eius, et nos erimus innoxii; cunctorum autem sanguis, qui tecum fuerint in domo, redundabit in caput nostrum, si eos aliquis tetigerit.
JOSH|2|20|Quod si prodideris hoc verbum, erimus mundi ab hoc iuramento, quo adiurasti nos ".
JOSH|2|21|Et illa respondit: " Sicut locuti estis, ita fiat ". Dimittensque eos, ut pergerent, appendit funiculum coccineum in fenestra.
JOSH|2|22|Illi vero ambulantes pervenerunt ad montana et manserunt ibi tres dies, donec reverterentur, qui fuerant persecuti; quaerentes enim per omnem viam non reppererunt eos.
JOSH|2|23|Duo viri reversi sunt et descenderunt de monte et, transmisso Iordane, venerunt ad Iosue filium Nun narraveruntque ei omnia, quae acciderant sibi,
JOSH|2|24|atque dixerunt: " Tradidit Dominus in manus nostras omnem terram, et timore prostrati sunt cuncti habitatores eius in conspectu nostro ".
JOSH|3|1|Igitur Iosue de nocte consur gens movit castra. Egredientes que de Settim venerunt ad Iordanem, ipse et omnes filii Israel; et morati sunt ibi, antequam transirent.
JOSH|3|2|Tribus diebus evolutis, transierunt praefecti per castrorum medium
JOSH|3|3|et praeceperunt populo: " Quando videritis arcam foederis Domini Dei vestri et sacerdotes stirpis leviticae portantes eam, vos quoque consurgite et sequimini eam
JOSH|3|4|- sitque inter vos et arcam spatium cubitorum duum fere milium, et cavete, ne appropinquetis ad eam - ut sciatis per quam viam ingrediamini, quia prius non ambulastis per eam ".
JOSH|3|5|Dixitque Iosue ad populum: " Sanctificamini; cras enim faciet Dominus inter vos mirabilia ".
JOSH|3|6|Et ait ad sacerdotes: " Tollite arcam foederis et praecedite populum ". Qui tulerunt et ambulaverunt ante eos.
JOSH|3|7|Dixitque Dominus ad Iosue: " Hodie incipiam exaltare te coram omni Israel, ut sciant quod, sicut cum Moyse fui, ita et tecum sim.
JOSH|3|8|Tu autem praecipe sacerdotibus, qui portant arcam foederis, et dic eis: Cum veneritis ad oram aquae Iordanis, state in Iordane".
JOSH|3|9|Dixitque Iosue ad filios Israel: " Accedite huc et audite verba Domini Dei vestri ".
JOSH|3|10|Et rursum: " In hoc, inquit, scietis quod Deus vivens in medio vestri est et disperdet in conspectu vestro Chananaeum et Hetthaeum, Hevaeum et Pherezaeum, Gergesaeum quoque et Amorraeum et Iebusaeum.
JOSH|3|11|Ecce arca foederis Domini omnis terrae antecedet vos per Iordanem.
JOSH|3|12|Parate duodecim viros de tribubus Israel, singulos per singulas tribus;
JOSH|3|13|et cum posuerint vestigia pedum suorum sacerdotes, qui portant arcam Domini Dei universae terrae, in aquis Iordanis, aquae, quae inferiores sunt, decurrent, quae autem desuper veniunt, in una mole consistent ".
JOSH|3|14|Igitur egressus est populus de tabernaculis suis, ut transiret Iordanem; et sacerdotes, qui portabant arcam foederis, pergebant ante eum.
JOSH|3|15|Veneruntque usque ad Iordanem et, pedibus eorum in ora aquae tinctis - Iordanis autem omnes ripas alvei sui toto tempore messis impleverat -
JOSH|3|16|steterunt aquae desuper descendentes in loco uno instar molis procul valde apud urbem, quae vocatur Adam, ex latere Sarthan; quae autem inferiores erant, in mare Arabae, quod est mare Salsissimum, descenderunt, usquequo omnino deficerent.
JOSH|3|17|Populus autem incedebat contra Iericho, et sacerdotes, qui portabant arcam foederis Domini, stabant super siccam humum in medio Iordanis firmiter, donec omnis Israel compleret per arentem alveum transitum Iordanis.
JOSH|4|1|Quibus transgressis, dixit Dominus ad Iosue:
JOSH|4|2|" Sumite vobis de populo duodecim viros singulos per singulas tribus
JOSH|4|3|et praecipite eis, ut tollant de medio Iordanis alveo, ubi firmiter steterunt sacerdotum pedes, duodecim lapides; quos portabitis vobiscum et ponetis in loco castrorum, ubi fixeritis hac nocte tentoria ".
JOSH|4|4|Vocavitque Iosue duodecim viros, quos elegerat de filiis Israel, singulos de tribubus singulis,
JOSH|4|5|et ait ad eos: " Ite ante arcam Domini Dei vestri ad Iordanis medium et portate singuli singulos lapides in umeris vestris, iuxta numerum tribuum filiorum Israel,
JOSH|4|6|ut sit hoc signum inter vos. Quando interrogaverint vos filii vestri cras dicentes: "Quid sibi volunt isti lapides?",
JOSH|4|7|respondebitis eis: Defecerunt aquae Iordanis ante arcam foederis Domini, cum transiret eum; idcirco positi sunt lapides isti in monumentum filiis Israel usque in aeternum ".
JOSH|4|8|Fecerunt ergo filii Israel, sicut eis praecepit Iosue, portantes de medio Iordanis alveo duodecim lapides, ut ei Dominus imperarat, iuxta numerum tribuum filiorum Israel, usque ad locum, in quo castrametati sunt; ibique posuerunt eos.
JOSH|4|9|Alios quoque duodecim lapides posuit Iosue in medio Iordanis alveo, ubi steterunt sacerdotes, qui portabant arcam foederis; et sunt ibi usque in praesentem diem.
JOSH|4|10|Sacerdotes autem, qui portabant arcam, stabant in Iordanis medio, donec omnia complerentur, quae Iosue ut loqueretur ad populum praeceperat Dominus secundum omnia, quae dixerat ei Moyses. Festinavitque populus et transiit.
JOSH|4|11|Cumque transissent omnes, transivit et arca Domini; sacerdotesque pergebant ante populum.
JOSH|4|12|Filii quoque Ruben et Gad et dimidia tribus Manasse armati praecedebant filios Israel, sicut eis praeceperat Moyses;
JOSH|4|13|quadraginta fere milia expeditorum ad pugnam incedebant coram Domino in campestria Iericho.
JOSH|4|14|In illo die magnificavit Dominus Iosue coram omni Israel, ut timerent eum, sicut timuerant Moysen, omnibus diebus vitae suae.
JOSH|4|15|Dixitque ad eum:
JOSH|4|16|" Praecipe sacerdotibus, qui portant arcam testimonii, ut ascendant de Iordane ".
JOSH|4|17|Qui praecepit eis dicens: " Ascendite de Iordane ".
JOSH|4|18|Cumque ascendissent portantes arcam foederis Domini et siccam humum calcare coepissent, reversae sunt aquae in alveum suum et fluebant sicut ante super omnes ripas suas.
JOSH|4|19|Populus autem ascendit de Iordane decimo die mensis primi, et castrametati sunt in Galgalis, in termino orientali Iericho.
JOSH|4|20|Duodecim quoque lapides, quos de Iordanis alveo sumpserant, posuit Iosue in Galgalis.
JOSH|4|21|Et dixit ad filios Israel: " Quando interrogaverint filii vestri cras patres suos et dixerint eis: "Quid sibi volunt isti lapides?",
JOSH|4|22|docebitis eos atque dicetis: Per arentem alveum transivit Israel Iordanem istum,
JOSH|4|23|siccante Domino Deo vestro aquas eius in conspectu vestro, donec transiretis,
JOSH|4|24|sicut fecerat prius in mari Rubro, quod siccavit coram nobis, donec transiremus,
JOSH|4|25|ut cognoscant omnes terrarum populi fortissimam Domini manum, et ut vos timeatis Dominum Deum vestrum omni tempore ".
JOSH|5|1|Postquam ergo audierunt om nes reges Amorraeorum, qui ha bitabant trans Iordanem ad occidentalem plagam, et cuncti reges Chanaan, qui propinqua possidebant Magno mari loca, quod siccasset Dominus fluenta Iordanis coram filiis Israel, donec transirent, dissolutum est cor eorum, et non remansit in eis spiritus coram filiis Israel.
JOSH|5|2|Eo tempore ait Dominus ad Iosue: " Fac tibi cultros lapideos et circumcide iterum secundo filios Israel ".
JOSH|5|3|Fecit, quod iusserat Dominus, et circumcidit filios Israel in colle Praeputiorum.
JOSH|5|4|Haec autem causa est secundae circumcisionis: omnis populus, qui egressus est ex Aegypto, generis masculini, universi bellatores viri mortui sunt in deserto in via;
JOSH|5|5|qui omnes circumcisi erant. Populus autem, qui natus est in deserto, incircumcisus fuit.
JOSH|5|6|Per quadraginta enim annos ambulabant filii Israel, donec consumerentur omnes homines bellatores, qui non audierant vocem Domini, et quibus iuraverat, ut non ostenderet eis terram, super qua iuraverat patribus eorum, ut daret illis terram lacte et melle manantem.
JOSH|5|7|Horum filii in locum successerunt patrum et circumcisi sunt a Iosue, quia, sicut nati fuerant, in praeputio erant, nec eos in via aliquis circumciderat.
JOSH|5|8|Postquam autem omnes circumcisi sunt, manserunt in eodem castrorum loco, donec sanarentur.
JOSH|5|9|Dixitque Dominus ad Iosue: " Hodie abstuli opprobrium Aegypti a vobis ". Vocatumque est nomen loci illius Galgala usque in praesentem diem.
JOSH|5|10|Manseruntque filii Israel in Galgalis et fecerunt Pascha quarta decima die mensis ad vesperum in campestribus Iericho;
JOSH|5|11|et comederunt de frugibus terrae a die altero, azymos panes et polentam hoc ipso die.
JOSH|5|12|Defecitque manna a die sequenti, postquam comederunt de frugibus terrae, nec usi sunt ultra cibo illo filii Israel, sed comederunt de frugibus terrae Chanaan in anno illo.
JOSH|5|13|Cum autem esset Iosue in agro urbis Iericho, levavit oculos et vidit virum stantem contra se et evaginatum tenentem gladium; perrexitque ad eum et ait: " Noster es an adversariorum? ".
JOSH|5|14|Qui respondit: " Nequaquam, sed sum princeps exercitus Domini et nunc veni ".
JOSH|5|15|Cecidit Iosue pronus in terram et adorans ait: " Quid Dominus meus loquitur ad servum suum? ".
JOSH|5|16|Et dixit princeps exercitus Domini ad Iosue: " Solve calceamentum de pedibus tuis; locus enim, in quo stas, sanctus est ". Fecitque Iosue, ut sibi fuerat imperatum.
JOSH|6|1|Iericho autem erat munita et clausa coram filiis Israel, et nul lus egredi audebat aut ingredi.
JOSH|6|2|Dixitque Dominus ad Iosue: " Ecce dedi in manu tua Iericho et regem eius omnesque fortes viros.
JOSH|6|3|Circuite urbem cuncti bellatores semel per diem: sic facietis sex diebus.
JOSH|6|4|Septem sacerdotes portabunt septem bucinas, cornua arietum, ante arcam foederis. Die autem septimo septies circuibitis civitatem, et sacerdotes clangent bucinis.
JOSH|6|5|Cumque insonuerit vox tubae longior et in auribus vestris increpuerit, conclamabit omnis populus vociferatione maxima, et muri funditus corruent civitatis; ingredienturque singuli per locum, contra quem steterint ".
JOSH|6|6|Vocavit ergo Iosue filius Nun sacerdotes et dixit ad eos: " Tollite arcam foederis, et septem alii sacerdotes tollant septem bucinas et incedant ante arcam Domini ".
JOSH|6|7|Ad populum quoque ait: " Vadite et circuite civitatem, et viri armati praecedant arcam Domini ".
JOSH|6|8|Cumque Iosue verba finisset, septem sacerdotes septem bucinis clangebant ante arcam foederis Domini,
JOSH|6|9|omnisque armatus exercitus praecedebat sacerdotes clangentes, reliquum vulgus arcam sequebatur, ac bucinis omnia concrepabant.
JOSH|6|10|Praeceperat autem Iosue populo dicens: " Non clamabitis, nec audietur vox vestra, neque ullus sermo ex ore vestro egredietur, donec veniat dies, in quo dicam vobis: Clamate et vociferamini ".
JOSH|6|11|Circuivit ergo arca Domini civitatem per diem, et reversi in castra pernoctaverunt ibi.
JOSH|6|12|Igitur, Iosue de nocte consurgente, tulerunt sacerdotes arcam Domini,
JOSH|6|13|et septem ex eis septem bucinas, cornua arietum, praecedebantque arcam Domini ambulantes atque clangentes, et armatus populus ibat ante eos; vulgus autem reliquum sequebatur arcam, bucinis personantibus.
JOSH|6|14|Circuieruntque civitatem secundo die semel et reversi sunt in castra; sic fecerunt sex diebus.
JOSH|6|15|Die autem septimo, diluculo consurgentes circuierunt urbem eodem modo septies; in illo die tantum circuierunt urbem septies.
JOSH|6|16|Cumque septimo circuitu clangerent bucinis sacerdotes, dixit Iosue ad populum: " Vociferamini! Tradidit enim vobis Dominus civitatem.
JOSH|6|17|Sitque civitas anathema, ipsa et omnia, quae in ea sunt, Domino; sola Rahab meretrix vivat cum universis, qui cum ea in domo sunt: abscondit enim nuntios, quos direximus.
JOSH|6|18|Vos autem cavete, ne de anathemate quippiam auferatis et sitis praevaricationis rei, et omnia castra Israel anathema sint atque turbentur.
JOSH|6|19|Quidquid auri et argenti fuerit et vasorum aeneorum ac ferri, Domino consecretur repositum in thesauris eius ".
JOSH|6|20|Igitur, omni vociferante populo et clangentibus tubis, postquam in aures multitudinis vox sonitusque increpuit, muri ilico corruerunt; et ascendit unusquisque per locum, qui contra se erat, ceperuntque civitatem.
JOSH|6|21|Et interfecerunt omnia, quae erant in ea, a viro usque ad mulierem, ab infante usque ad senem; boves quoque et oves et asinos in ore gladii percusserunt.
JOSH|6|22|Duobus autem viris, qui exploratores missi fuerant, dixit Iosue: " Ingredimini domum mulieris meretricis et producite eam et omnia, quae illius sunt, sicut illi iuramento firmastis ".
JOSH|6|23|Ingressique iuvenes eduxerunt Rahab et parentes eius, fratres quoque et cunctam supellectilem ac cognationem illius et extra castra Israel manere fecerunt.
JOSH|6|24|Urbem autem et omnia, quae erant in ea, succenderunt, absque argento et auro et vasis aeneis ac ferro, quae in aerarium domus Domini consecrarunt.
JOSH|6|25|Rahab vero meretricem et domum patris eius et omnia, quae habebat, fecit Iosue vivere; et habitavit in medio Israel usque in praesentem diem, eo quod absconderit nuntios, quos miserat Iosue, ut explorarent Iericho.In tempore illo imprecatus est Iosue dicens:
JOSH|6|26|"Maledictus vir coram Domino, qui suscitaverit et aedificaverit civitatem Iericho; in primogenito suo fundamenta illius faciet et in novissimo liberorum ponet portas eius ".
JOSH|6|27|Fuit ergo Dominus cum Iosue, et nomen eius in omni terra vulgatum est.
JOSH|7|1|Filii autem Israel praevaricati sunt mandatum et usurpaverunt de anathemate: nam Achan filius Charmi filii Zabdi filii Zarae de tribu Iudae tulit aliquid de anathemate. Iratusque est Dominus contra filios Israel.
JOSH|7|2|Cumque mitteret Iosue de Iericho viros contra Hai, quae est iuxta Bethaven ad orientalem plagam oppidi Bethel, dixit eis: " Ascendite et explorate terram ". Qui praecepta complentes exploraverunt Hai
JOSH|7|3|et reversi dixerunt ei: " Non ascendat omnis populus, sed duo vel tria milia virorum pergant et deleant civitatem. Noli vexare omnem populum contra hostes paucissimos ".
JOSH|7|4|Ascenderunt ergo tria fere milia pugnatorum, qui statim terga verterunt coram viris urbis Hai,
JOSH|7|5|qui percusserunt ex eis circiter triginta et sex homines persecutique sunt eos de porta usque ad Sabarim et percusserunt eos in descensu; pertimuitque cor populi et instar aquae liquefactum est.
JOSH|7|6|Iosue vero scidit vestimenta sua et cecidit pronus in terram coram arca Domini usque ad vesperum, tam ipse quam omnes senes Israel; miseruntque pulverem super capita sua.
JOSH|7|7|Et dixit Iosue: " Heu, Domine Deus, quid voluisti traducere populum istum Iordanem fluvium, ut traderes nos in manus Amorraei et perderes? Utinam mansissemus trans Iordanem!
JOSH|7|8|Quaeso, Domine, quid dicam videns Israelem hostibus suis terga vertentem?
JOSH|7|9|Audient Chananaei et omnes habitatores terrae ac pariter conglobati circumdabunt nos atque delebunt nomen nostrum de terra. Et quid facies magno nomini tuo? ".
JOSH|7|10|Dixitque Dominus ad Iosue: " Surge! Cur iaces pronus in terra?
JOSH|7|11|Peccavit Israel et praevaricatus est pactum meum, quod mandaveram eis; tuleruntque de anathemate et furati sunt atque mentiti et absconderunt inter vasa sua.
JOSH|7|12|Nec poterunt filii Israel stare ante hostes suos eosque fugient, quia facti sunt anathema; non ero ultra vobiscum, donec conteratis anathema de medio vestri.
JOSH|7|13|Surge! Sanctifica populum et dic eis: Sanctificamini in crastinum. Haec enim dicit Dominus, Deus Israel: Anathema in medio tui est, Israel! Non poteris stare coram hostibus tuis, donec auferatis anathema de medio vestri.
JOSH|7|14|Accedetisque mane singuli per tribus vestras; et quamcumque tribum Dominus designaverit, accedet per cognationes suas et cognatio per domos domusque per viros:
JOSH|7|15|et quicumque ille in hoc facinore fuerit deprehensus, comburetur igni cum omnibus, quae ipsius sunt, quoniam praevaricatus est pactum Domini et fecit nefas in Israel ".
JOSH|7|16|Surgens itaque Iosue mane applicuit Israel per tribus suas, et inventa est tribus Iudae.
JOSH|7|17|Quae cum iuxta familias suas esset oblata, inventa est familia Zarae; illam quoque per domos offerens repperit Zabdi.
JOSH|7|18|Cuius domum in singulos dividens viros invenit Achan filium Charmi filii Zabdi filii Zarae de tribu Iudae.
JOSH|7|19|Et ait Iosue ad Achan: " Fili mi, da gloriam Domino, Deo Israel, et confitere atque indica mihi quid feceris; ne abscondas ".
JOSH|7|20|Responditque Achan Iosue et dixit ei: " Vere ego peccavi Domino, Deo Israel, et sic et sic feci:
JOSH|7|21|Vidi enim inter spolia pallium de Sennaar valde bonum et ducentos siclos argenti regulamque auream quinquaginta siclorum; et concupiscens abstuli et abscondi in terra contra medium tabernaculi mei argentumque subter ".
JOSH|7|22|Misit ergo Iosue ministros, qui currentes ad tabernaculum illius reppererunt cuncta abscondita in eodem loco et argentum simul;
JOSH|7|23|auferentesque de tentorio tulerunt ea ad Iosue et ad omnes filios Israel proieceruntque ante Dominum.
JOSH|7|24|Tollens itaque Iosue Achan filium Zarae argentumque et pallium et auream regulam filiosque eius et filias, boves et asinos et oves ipsumque tabernaculum et cunctam supellectilem - et omnis Israel cum eo - duxerunt eos ad vallem Achor,
JOSH|7|25|ubi dixit Iosue: " Quia turbasti nos, exturbet te Dominus in die hac ". Lapidavitque eum omnis Israel; et cuncta, quae illius erant, igne consumpta sunt.
JOSH|7|26|Congregaverunt quoque super eum acervum magnum lapidum, qui permanet usque in praesentem diem. Et aversus est furor Domini ab eis; vocatumque est nomen loci illius vallis Achor usque hodie.
JOSH|8|1|Dixit autem Dominus ad Iosue: " Ne timeas neque formides; tol le tecum omnem multitudinem pugnatorum et consurgens ascende in oppidum Hai: ecce tradidi in manu tua regem eius et populum urbemque et terram eius.
JOSH|8|2|Faciesque urbi Hai et regi eius, sicut fecisti Iericho et regi illius; praedam vero et omnia animantia diripietis vobis. Pone insidias urbi post eam ".
JOSH|8|3|Surrexitque Iosue et omnis exercitus bellatorum cum eo, ut ascenderent in Hai; et electa triginta milia virorum fortium misit nocte
JOSH|8|4|praecepitque eis dicens: "Collocamini in insidiis post civitatem nec longius recedatis ab illa; et eritis omnes parati.
JOSH|8|5|Ego autem et reliqua multitudo, quae mecum est, accedemus ex adverso contra urbem; cumque exierint contra nos sicut ante, fugiemus et terga vertemus,
JOSH|8|6|donec persequentes ab urbe longius protrahantur: putabunt enim nos fugere sicut prius.
JOSH|8|7|Nobis ergo fugientibus et illis sequentibus, consurgetis de insidiis et capietis civitatem; tradetque eam Dominus Deus vester in manus vestras.
JOSH|8|8|Cumque ceperitis, succendite eam; secundum verbum Domini facietis. Ecce mandavi vobis".
JOSH|8|9|Dimisitque eos, et perrexerunt ad insidiarum locum sederuntque inter Bethel et Hai ad occidentalem plagam urbis Hai. Iosue autem nocte illa in medio mansit populi.
JOSH|8|10|Surgensque diluculo recensuit populum et ascendit cum senioribus in fronte exercitus.
JOSH|8|11|Cumque omnes pugnatores cum eo ascendissent et appropinquassent civitati, steterunt ad septentrionalem urbis plagam, inter quam et eos vallis media erat.
JOSH|8|12|Et elegit fere quinque milia viros et posuit in insidiis inter Bethel et Hai ex occidentali parte eiusdem civitatis.
JOSH|8|13|Et posuit populus tota castra, quae erant in aquilone urbis, et agmen extremum ad occidentalem plagam urbis. Abiit ergo Iosue nocte illa et stetit in vallis medio.
JOSH|8|14|Quod cum vidisset rex Hai, festinavit mane et egressus est cum omni exercitu civitatis direxitque aciem contra Arabam ignorans quod post tergum laterent insidiae.
JOSH|8|15|Iosue vero et omnis Israel cesserunt loco simulantes metum et fugientes per solitudinis viam.
JOSH|8|16|Et convocatus est totus populus, qui erat in civitate, ad persequendum eos, et persecuti sunt eos. Cumque recessissent a civitate,
JOSH|8|17|et ne unus quidem in urbe Hai remansisset, qui non persequeretur Israel, et apertam urbem reliquissent,
JOSH|8|18|dixit Dominus ad Iosue: "Leva acinacem, quod in manu tua est, contra urbem Hai, quoniam tibi tradam eam ".
JOSH|8|19|Cumque elevasset acinacem ex adverso civitatis, insidiae, quae latebant, surrexerunt confestim et currentes ad civitatem ceperunt et cito succenderunt eam.
JOSH|8|20|Viri autem civitatis, qui persequebantur Iosue, respicientes et videntes fumum urbis ad caelum usque conscendere, non potuerunt ultra huc illucque diffugere, praesertim cum hi, qui simulaverant fugam et tendebant ad solitudinem, contra persequentes conversi essent.
JOSH|8|21|Vidensque Iosue et omnis Israel quod capta esset civitas, et fumus urbis ascenderet, reversi percusserunt viros Hai.
JOSH|8|22|Siquidem et illi, qui ceperant et succenderant civitatem, egressi sunt ex urbe in occursum eorum et hostes medios habuerunt. Cum ergo ex utraque parte adversarii caederentur, ita ut nullus de tanta multitudine salvaretur,
JOSH|8|23|regem quoque urbis Hai apprehenderunt viventem et obtulerunt Iosue.
JOSH|8|24|Igitur, omnibus habitatoribus Hai interfectis, qui Israelem ad deserta tendentem fuerant persecuti, et in eodem loco gladio corruentibus, reversi filii Israel percusserunt civitatem ore gladii.
JOSH|8|25|Erant autem, qui in eo die conciderant, a viro usque ad mulierem duodecim milia hominum omnes urbis Hai.
JOSH|8|26|Iosue vero non contraxit manum, quam in sublime porrexerat tenens acinacem, donec interficerentur omnes habitatores Hai.
JOSH|8|27|Iumenta tantum et praedam civitatis diviserunt sibi filii Israel, sicut praeceperat Dominus Iosue.
JOSH|8|28|Qui succendit urbem et fecit eam tumulum sempiternum, desolationem usque in praesentem diem.
JOSH|8|29|Regem quoque eius suspendit in ligno usque ad vesperum; et ad solis occasum praecepit Iosue, et deposuerunt cadaver eius de ligno proieceruntque in ipso introitu portae civitatis, congesto super eum magno acervo lapidum, qui permanet usque in praesentem diem.
JOSH|8|30|Tunc aedificavit Iosue altare Domino, Deo Israel, in monte Hebal,
JOSH|8|31|sicut praeceperat Moyses famulus Domini filiis Israel, et scriptum est in volumine legis Moysi, altare de lapidibus impolitis, quos ferrum non tetigit. Et obtulerunt super eo holocausta Domino immolaveruntque pacificas victimas.
JOSH|8|32|Et scripsit ibi super lapides exemplar legis Moysi, quod ille scripserat coram filiis Israel.
JOSH|8|33|Omnis autem populus et maiores natu praefectique ac iudices stabant ex utraque parte arcae in conspectu sacerdotum levitici generis, qui portabant arcam foederis Domini, ut advena ita et indigena. Media eorum pars iuxta montem Garizim et media iuxta montem Hebal, sicut praeceperat Moyses famulus Domini ad benedicendum populo Israel primum;
JOSH|8|34|post haec legit omnia verba legis, benedictionem et maledictionem, secundum cuncta, quae scripta erant in legis volumine.
JOSH|8|35|Nihil ex his, quae Moyses iusserat, omisit legere, sed universa replicavit coram omni congregatione Israel, mulieribus ac parvulis et advenis, qui inter eos morabantur.
JOSH|9|1|Quibus auditis, cuncti reges, qui trans Iordanem versabantur in montanis et in Sephela, in omni litore maris Magni, hi quoque, qui habitabant usque ad Libanum, Hetthaeus et Amorraeus, Chananaeus, Pherezaeus et Hevaeus et Iebusaeus
JOSH|9|2|congregati sunt pariter, ut pugnarent contra Iosue et Israel uno animo eademque sententia.
JOSH|9|3|At hi, qui habitabant in Gabaon, audientes cuncta, quae fecerat Iosue Iericho et Hai,
JOSH|9|4|et callide cogitantes tulerunt sibi cibaria, saccos veteres asinis imponentes et utres vinarios vetustos, scissos atque consutos,
JOSH|9|5|calceamentaque perantiqua, quae ad indicium vetustatis pittaciis consuta erant, induti veteribus vestimentis; panes quoque, quos portabant ob viaticum, duri erant et in frusta comminuti.
JOSH|9|6|Perrexeruntque ad Iosue, qui tunc morabatur in castris Galgalae, et dixerunt ei atque omni simul Israeli: " De terra longinqua venimus pactum vobiscum facere cupientes ". Responderuntque viri Israel ad Hevaeos atque dixerunt:
JOSH|9|7|" Ne forte in medio nostri habitetis, et non possimus foedus inire vobiscum ".
JOSH|9|8|At illi ad Iosue: " Servi, inquiunt, tui sumus ". Quibus Iosue ait: " Quinam estis et unde venistis? ".
JOSH|9|9|Responderunt: " De terra longinqua valde venerunt servi tui in nomine Domini Dei tui; audivimus enim famam potentiae eius, cuncta, quae fecit in Aegypto
JOSH|9|10|et duobus Amorraeorum regibus trans Iordanem, Sehon regi Hesebon et Og regi Basan, qui erat in Astharoth.
JOSH|9|11|Dixeruntque nobis seniores et omnes habitatores terrae nostrae: Tollite in manibus cibaria in viam et occurrite eis ac dicite: Servi vestri sumus; foedus inite nobiscum".
JOSH|9|12|En panes: quando egressi sumus de domibus nostris, ut veniremus ad vos, calidos sumpsimus; nunc sicci facti sunt et vetustate nimia comminuti.
JOSH|9|13|Utres vini novos implevimus, nunc rupti sunt et soluti; vestes et calceamenta, quibus induimur et quae habemus in pedibus, ob longitudinem largioris viae trita sunt et paene consumpta ".
JOSH|9|14|Susceperunt igitur viri de cibariis eorum et os Domini non interrogaverunt.
JOSH|9|15|Fecitque Iosue cum eis pacem et, inito foedere, pollicitus est quod viverent; principes quoque coetus iuraverunt eis.
JOSH|9|16|Post dies autem tres initi foederis, audierunt quod in vicino et inter eos habitarent.
JOSH|9|17|Moveruntque castra filii Israel et venerunt ad civitates eorum die tertio, quarum haec vocabula sunt: Gabaon et Cephira et Beroth et Cariathiarim;
JOSH|9|18|et non percusserunt eos filii Israel, eo quod iurassent eis principes coetus in nomine Domini, Dei Israel. Murmuravit itaque omnis coetus contra principes,
JOSH|9|19|qui responderunt eis: "Iuravimus illis in nomine Domini, Dei Israel, et idcirco non possumus eos contingere.
JOSH|9|20|Sed hoc faciemus eis: reserventur quidem, ut vivant, ne contra nos ira Domini concitetur, si peieraverimus;
JOSH|9|21|sed sic vivant, ut in usus universae multitudinis ligna caedant aquasque comportent ".Quibus haec loquentibus,
JOSH|9|22|vocavit Gabaonitas Iosue et dixit eis: " Cur nos decipere fraude voluistis, ut diceretis: "Procul valde habitamus a vobis", cum in medio nostri sitis?
JOSH|9|23|Itaque sub maledictione eritis, et non deficiet de stirpe vestra servus ligna caedens aquasque comportans in domum Dei mei".
JOSH|9|24|Qui responderunt: " Nuntiatum est nobis servis tuis, quod mandasset Dominus Deus tuus Moysi servo suo, ut traderet vobis omnem terram et disperderet cunctos habitatores eius; timuimus igitur valde pro animabus nostris, vestro terrore compulsi, et hoc consilium inivimus.
JOSH|9|25|Nunc autem in manu tua sumus: quod tibi bonum et rectum videtur, fac nobis ".
JOSH|9|26|Fecit ergo Iosue, ut dixerat, et liberavit eos de manu filiorum Israel, ut non occiderentur.
JOSH|9|27|Decrevitque in illo die esse eos in ministerium cuncti populi et altaris Domini caedentes ligna et aquas comportantes usque in praesens tempus pro loco, quem Dominus elegisset.
JOSH|10|1|Quae cum audisset Adonise dec rex Ierusalem, quod scili cet cepisset Iosue Hai et subvertisset eam - sicut enim fecerat Iericho et regi eius, sic fecit Hai et regi illius - et quod pacem fecissent Gabaonitae cum Israel et essent in medio eorum,
JOSH|10|2|timuerunt valde. Urbs enim magna erat Gabaon, sicut una regalium civitatum, et maior oppido Hai, omnesque viri eius bellatores fortissimi.
JOSH|10|3|Misit ergo Adonisedec rex Ierusalem ad Oham regem Hebron et ad Pharam regem Ierimoth, ad Iaphia quoque regem Lachis et ad Dabir regem Eglon dicens:
JOSH|10|4|" Ascendite ad me et ferte praesidium, ut expugnemus Gabaon, quia fecit pacem cum Iosue et filiis Israel ".
JOSH|10|5|Congregati igitur ascenderunt quinque reges Amorraeorum: rex Ierusalem, rex Hebron, rex Ierimoth, rex Lachis, rex Eglon simul cum exercitibus suis; et castrametati sunt circa Gabaon oppugnantes eam.
JOSH|10|6|Habitatores autem Gabaon miserunt ad Iosue, qui tunc morabatur in castris apud Galgalam, et dixerunt ei: " Ne retrahas manus tuas ab auxilio servorum tuorum! Ascende cito et libera nos ferque praesidium: convenerunt enim adversum nos omnes reges Amorraeorum, qui habitant in montanis ".
JOSH|10|7|Ascenditque Iosue de Galgalis, et omnis exercitus bellatorum cum eo, viri fortissimi.
JOSH|10|8|Dixitque Dominus ad Iosue: "Ne timeas eos! In manus enim tuas tradidi illos; nullus tibi ex eis resistere poterit ".
JOSH|10|9|Irruit itaque Iosue super eos repente tota ascendens nocte de Galgalis,
JOSH|10|10|et conturbavit eos Dominus a facie Israel; contrivitque plaga magna in Gabaon ac persecutus est per viam ascensus Bethoron et percussit usque Azeca et Maceda.
JOSH|10|11|Cumque fugerent filios Israel et essent in descensu Bethoron, Dominus misit super eos lapides magnos de caelo usque Azeca, et mortui sunt multo plures lapidibus grandinis, quam quos gladio percusserant filii Israel.
JOSH|10|12|Tunc locutus est Iosue Domino in die, qua tradidit Amorraeum in conspectu filiorum Israel, dixitque coram Israel: Sol, in Gabaon ne movearis,et luna, in valle Aialon ".
JOSH|10|13|Steteruntque sol et luna,donec ulcisceretur se gens de inimicis suis.Nonne scriptum est hoc in libro Iusti? Stetit itaque sol in medio caeli et non festinavit occumbere spatio unius fere diei.
JOSH|10|14|Non fuit antea et postea sicut dies illa, oboediente Domino voci hominis, quia Dominus pugnavit pro Israel.
JOSH|10|15|Reversusque est Iosue cum omni Israel in castra Galgalae.
JOSH|10|16|Fugerant autem quinque reges et se absconderant in spelunca urbis Maceda.
JOSH|10|17|Nuntiatumque est Iosue quod inventi essent quinque reges latentes in spelunca urbis Maceda.
JOSH|10|18|Qui praecepit: " Volvite saxa ingentia ad os speluncae et ponite viros, qui clausos custodiant.
JOSH|10|19|Vos autem nolite stare, sed persequimini hostes et extremos quoque fugientium caedite; ne dimittatis eos urbium suarum intrare praesidia, quia tradidit eos Dominus Deus vester in manus vestras ".
JOSH|10|20|Caesis igitur adversariis plaga maxima usque ad internecionem, ut reliquiae tantum ex eis effugere possent in civitates munitas,
JOSH|10|21|reversus est omnis exercitus ad Iosue in Maceda ad castra, sani et integri; nullusque contra filios Israel mutire ausus est.
JOSH|10|22|Praecepitque Iosue dicens: " Aperite os speluncae et producite ad me quinque reges, qui in ea latitant ".
JOSH|10|23|Feceruntque sic et eduxerunt ad eum quinque reges de spelunca: regem Ierusalem, regem Hebron, regem Ierimoth, regem Lachis, regem Eglon.
JOSH|10|24|Cumque educti essent ad eum, vocavit omnes viros Israel et ait ad principes exercitus, qui secum erant: "Accedite et ponite pedes super colla regum istorum". Qui cum accessissent et subiectorum colla pedibus calcarent,
JOSH|10|25|rursum ait ad eos: " Nolite timere nec paveatis; confortamini et estote robusti! Sic enim faciet Dominus cunctis hostibus vestris, adversum quos dimicatis ".
JOSH|10|26|Percussitque Iosue et interfecit eos atque suspendit super quinque ligna; fueruntque suspensi usque ad vesperum.
JOSH|10|27|Cumque occumberet sol, praecepit Iosue, ut deponerent eos de lignis; et depositos proiecerunt in speluncam, in qua latuerant, et posuerunt super os eius saxa ingentia, quae permanent usque in praesens.
JOSH|10|28|Eodem quoque die Macedam cepit Iosue et percussit eam in ore gladii regemque illius interfecit et omnes habitatores eius; non dimisit in ea ullas reliquias fecitque regi Maceda, sicut fecerat regi Iericho.
JOSH|10|29|Transivit cum omni Israel de Maceda in Lobna et pugnabat contra eam.
JOSH|10|30|Quam tradidit Dominus cum rege suo in manu Israel, percusseruntque urbem in ore gladii et omnes habitatores eius; non dimiserunt in ea ullas reliquias feceruntque regi Lobna, sicut fecerant regi Iericho.
JOSH|10|31|De Lobna transivit Iosue in Lachis cum omni Israel et, exercitu per gyrum disposito, oppugnabat eam.
JOSH|10|32|Tradiditque Dominus Lachis in manu Israel, qui cepit eam die altero; atque percussit in ore gladii omnemque animam, quae fuerat in ea, sicut fecerat Lobna.
JOSH|10|33|Eo tempore ascendit Horam rex Gazer, ut auxiliaretur Lachis; quem percussit Iosue cum omni populo eius usque ad internecionem.
JOSH|10|34|Transivitque de Lachis in Eglon cum omni Israel et circumdedit
JOSH|10|35|atque expugnavit eam eadem die percussitque in ore gladii omnes animas, quae erant in ea, iuxta omnia, quae fecerat Lachis.
JOSH|10|36|Ascendit quoque cum omni Israel de Eglon in Hebron et pugnavit contra eam.
JOSH|10|37|Cepitque eam et percussit in ore gladii, regem quoque eius et omnia oppida eius universasque animas, quae ibi fuerant commoratae; non reliquit ullas reliquias: sicut fecerat Eglon, sic fecit et Hebron, cuncta, quae in ea repperit, consumens gladio.
JOSH|10|38|Inde reversus cum omni Israel in Dabir oppugnavit
JOSH|10|39|et cepit eam; regem quoque eius et omnia oppida eius percussit in ore gladii; non dimisit in ea ullas reliquias: sicut fecerat Hebron et Lobna et regibus earum, sic fecit Dabir et regi illius.
JOSH|10|40|Percussit itaque Iosue omnem terram: montanam et Nageb atque Sephelam et declivia cum regibus suis; non dimisit in ea ullas reliquias, sed omne, quod spirare poterat, interfecit, sicut praeceperat Dominus, Deus Israel.
JOSH|10|41|Et percussit eos a Cadesbarne usque Gazam, omnem terram Gosen usque Gabaon,
JOSH|10|42|universosque reges et regiones eorum uno cepit impetu; Dominus enim, Deus Israel, pugnabat pro Israel.
JOSH|10|43|Reversusque est Iosue cum omni Israel ad locum castrorum in Galgala.
JOSH|11|1|Quae cum audisset Iabin rex Asor, misit ad Iobab regem Madon et ad regern Semeron atque ad regem Achsaph,
JOSH|11|2|ad reges quoque aquilonis, qui habitabant in montanis et in Araba contra meridiem Chenereth, in Sephela quoque et in regionibus Dor iuxta mare,
JOSH|11|3|Chananaeum in oriente et occidente, et Amorraeum atque Hetthaeum ac Pherezaeum et Iebusaeum in montanis, Hevaeum quoque, qui habitabat ad radices Hermon in terra Maspha.
JOSH|11|4|Egressique sunt omnes cum turmis suis, populus multus nimis sicut arena, quae est in litore maris, equi quoque et currus immensae multitudinis;
JOSH|11|5|conveneruntque omnes reges isti et castrametati sunt in unum ad aquas Merom, ut pugnarent contra Israel.
JOSH|11|6|Dixitque Dominus ad Iosue: "Ne timeas eos! Cras enim hac eadem hora ego tradam omnes istos occisos in conspectu Israel: equos eorum subnervabis et currus igne combures ".
JOSH|11|7|Venitque Iosue et omnis exercitus cum eo adversus illos ad aquas Merom subito, et irruerunt super eos.
JOSH|11|8|Tradiditque illos Dominus in manu Israel; qui percusserunt eos et persecuti sunt usque ad Sidonem magnam et Maserephoth in occidente campumque Maspha in oriente. Ita percussit omnes, ut nullas dimitteret ex eis reliquias;
JOSH|11|9|fecit sicut praeceperat ei Dominus: equos eorum subnervavit currusque combussit.
JOSH|11|10|Reversusque tempore illo cepit Asor et regem eius percussit gladio. Asor enim antiquitus inter omnia regna haec principatum tenebat.
JOSH|11|11|Percussitque omnes animas, quae ibidem morabantur; non dimisit in ea ullas reliquias, sed usque ad internecionem universa vastavit ipsamque urbem peremit incendio.
JOSH|11|12|Et omnes per circuitum civitates regesque earum cepit, percussit atque delevit, sicut praeceperat Moyses famulus Domini.
JOSH|11|13|Urbes tantum, quae erant in tumulis earum sitae, non succendit Israel; unam Asor solam Iosue flamma consumpsit.
JOSH|11|14|Omnemque praedam istarum urbium ac iumenta diviserunt sibi filii Israel, cunctis hominibus interfectis; nullum vivum reliquerunt.
JOSH|11|15|Sicut praeceperat Dominus Moysi servo suo, ita praecepit Moyses Iosue, et ille universa complevit; non praeteriit de universis mandatis ne unum quidem verbum, quod iusserat Dominus Moysi.
JOSH|11|16|Cepit itaque Iosue omnem terram hanc, montanam et Nageb terramque Gosen et Sephelam et Arabam montemque Israel et campestria eius,
JOSH|11|17|a monte Calvo, qui ascendit Seir, usque Baalgad in planitie Libani subter montem Hermon; omnes reges eorum cepit, percussit et occidit.
JOSH|11|18|Multo tempore pugnavit Iosue contra reges istos.
JOSH|11|19|Non fuit civitas, quae foedus iniret cum filiis Israel, praeter Hevaeum, qui habitabat in Gabaon: omnes bellando cepit.
JOSH|11|20|Domini enim sententia fuerat, ut indurarentur corda eorum, et pugnarent contra Israel et caderent et non mererentur ullam clementiam ac perirent, sicut praeceperat Dominus Moysi.
JOSH|11|21|In tempore illo venit Iosue et interfecit Enacim de montanis Hebron et Dabir et Anab et de omni monte Iudae et Israel urbesque eorum delevit.
JOSH|11|22|Non reliquit ullum de stirpe Enacim in terra filiorum Israel, absque civitatibus Gaza et Geth et Azoto, in quibus solis relicti sunt.
JOSH|11|23|Cepit ergo Iosue omnem terram, sicut locutus est Dominus ad Moysen, et tradidit eam in possessionem filiis Israel secundum partes et tribus suas; quievitque terra a proeliis.
JOSH|12|1|Hi sunt reges, quos percusserunt filii Israel et possederunt terram eorum trans Iordanem ad solis ortum, a torrente Arnon usque ad montem Hermon et omnem orientalem plagam Arabae.
JOSH|12|2|Sehon rex Amorraeorum, qui habitavit in Hesebon, dominatus est ab Aroer, quae sita est super ripam torrentis Arnon, et a media parte vallis et in dimidia parte Galaad usque ad torrentem Iaboc, qui est terminus filiorum Ammon;
JOSH|12|3|et in Araba usque ad mare Chenereth in oriente et usque ad mare Arabae, quod est mare Salsissimum, ad orientalem plagam in via, quae ducit Bethiesimoth, et in australi parte, quae iacet ad radices Phasga.
JOSH|12|4|Terminus Og regis Basan de reliquiis Raphaim, qui habitavit in Astharoth et in Edrai,
JOSH|12|5|et dominatus est in monte Hermon et in Salcha atque in universa Basan usque ad terminos Gesuri et Maachathi et in dimidia parte Galaad usque ad terminos Sehon regis Hesebon.
JOSH|12|6|Moyses famulus Domini et filii Israel percusserunt eos; tradiditque terram eorum Moyses in possessionem Rubenitis et Gaditis et dimidiae tribui Manasse.
JOSH|12|7|Hi sunt reges terrae, quos percussit Iosue et filii Israel trans Iordanem ad occidentalem plagam, a Baalgad in campo Libani usque ad montem Calvum, qui ascendit in Seir; tradiditque eam Iosue in possessionem tribubus Israel, singulis partes suas,
JOSH|12|8|tam in montanis quam in Sephela, in Araba et in declivibus et in solitudine ac in Nageb; Hetthaeus fuit et Amorraeus, Chananaeus et Pherezaeus, Hevaeus et Iebusaeus:
JOSH|12|9|rex Iericho unus, rex Hai, quae est ex latere Bethel, unus,
JOSH|12|10|rex Ierusalem unus, rex Hebron unus,
JOSH|12|11|rex Ierimoth unus, rex Lachis unus,
JOSH|12|12|rex Eglon unus, rex Gazer unus,
JOSH|12|13|rex Dabir unus, rex Gader unus,
JOSH|12|14|rex Horma unus, rex Arad unus,
JOSH|12|15|rex Lobna unus, rex Odollam unus,
JOSH|12|16|rex Maceda unus, rex Bethel unus,
JOSH|12|17|rex Thapphua unus, rex Opher unus,
JOSH|12|18|rex Aphec unus, rex Saron unus,
JOSH|12|19|rex Madon unus, rex Asor unus,
JOSH|12|20|rex Semeron unus, rex Achsaph unus,
JOSH|12|21|rex Thanach unus, rex Mageddo unus,
JOSH|12|22|rex Cedes unus, rex Iecnaam Carmeli unus,
JOSH|12|23|rex Dor et provinciae Dor unus, rex gentium Galgal unus,
JOSH|12|24|rex Thersa unus: omnes reges triginta unus.
JOSH|13|1|Iosue senex provectaeque aetatis erat, et dixit Dominus ad eum: " Senuisti et longaevus es; terraque latissima adhuc superest, quae necdum occupata est.
JOSH|13|2|Omnis videlicet Galilaea, regio Philisthim et universa Gesuri,
JOSH|13|3|a fluvio Sihor, qui est ad orientem Aegypti, usque ad terminos Accaron contra aquilonem, terra Chananaea, quae in quinque principes Philisthim dividitur, Gazaeos et Azotios, Ascalonitas, Getthaeos et Accaronitas ac Hevaei
JOSH|13|4|meridie; et omnis terra Chanaan de Ara Sidoniorum usque Apheca et terminos Amorraei;
JOSH|13|5|et terra Gibliorum et omnis Libanus in oriente a Baalgad sub monte Hermon usque ad introitum Emath,
JOSH|13|6|omnes, qui habitant in monte a Libano usque ad Maserephoth in occidente, universi Sidonii. Ego sum qui delebo eos a facie filiorum Israel. Sorte tantum distribue terram Israel in hereditatem, sicut praecepi tibi.
JOSH|13|7|Et nunc divide terram hanc in possessionem novem tribubus et dimidiae tribui Manasse ".
JOSH|13|8|Cum qua Ruben et Gad possederunt terram, quam tradidit eis Moyses famulus Domini trans fluenta Iordanis ad orientalem plagam:
JOSH|13|9|ab Aroer, quae sita est in ripa torrentis Arnon, et civitate in vallis medio, universaque campestria Medaba usque Dibon;
JOSH|13|10|et cunctas civitates Sehon regis Amorraei, qui regnavit in Hesebon, usque ad terminos filiorum Ammon;
JOSH|13|11|et Galaad ac terminos Gesuri et Maachathi omnemque montem Hermon et universam Basan usque Salcha,
JOSH|13|12|omne regnum Og in Basan, qui regnavit in Astharoth et Edrai - ipse fuit de reliquiis Raphaim C; percussitque eos Moyses atque delevit.
JOSH|13|13|Non autem disperdiderunt filii Israel Gesuri et Maachathi, et habitaverunt in medio Israel usque in praesentem diem.
JOSH|13|14|Tribui tantum Levi non dedit possessionem, sed sacrificia Domini, Dei Israel: ipsa est eius hereditas, sicut locutus est illi.
JOSH|13|15|Dedit ergo Moyses possessionem tribui filiorum Ruben iuxta cognationes suas.
JOSH|13|16|Fuitque terminus eorum ab Aroer, quae sita est in ripa torrentis Arnon, et a civitate in valle eiusdem torrentis media, et universa planities usque Medaba,
JOSH|13|17|Hesebon cunctaque oppida eius, quae sunt in campestribus: Dibon et Bamothbaal et Bethbaalmeon
JOSH|13|18|et Iasa et Cademoth et Mephaath,
JOSH|13|19|Cariathaim et Sabama et Serethsahar in monte convallis,
JOSH|13|20|Bethphegor et declivia Phasga et Bethiesimoth
JOSH|13|21|et omnes urbes campestres universumque regnum Sehon regis Amorraei, qui regnavit in Hesebon, quem percussit Moyses, ipsum et principes Madian, Evi et Recem et Sur et Hur et Rebe, duces Sehon habitatores terrae.
JOSH|13|22|Et Balaam filium Beor hariolum occiderunt filii Israel gladio cum ceteris interfectis.
JOSH|13|23|Factusque est terminus filiorum Ruben Iordanis fluvius. Haec est possessio Rubenitarum per cognationes suas, urbes et viculi earum.
JOSH|13|24|Deditque Moyses tribui Gad, filiis Gad, per cognationes suas possessionem, cuius hic est
JOSH|13|25|terminus: Iazer et omnes civitates Galaad dimidiaque pars terrae filiorum Ammon usque ad Aroer, quae est contra Rabba;
JOSH|13|26|et ab Hesebon usque Ramothmaspha et Betonim et a Mahanaim usque ad terminos Lodabar,
JOSH|13|27|in valle quoque Betharan et Bethnemra et Succoth et Saphon, reliqua pars regni Sehon regis Hesebon; Iordanis et terminus usque ad extremam partem maris Chenereth trans Iordanem ad orientalem plagam.
JOSH|13|28|Haec est possessio filiorum Gad per familias suas, civitates et villae earum.
JOSH|13|29|Dedit Moyses et dimidiae tribui filiorum Manasse, iuxta cognationes suas possessionem:
JOSH|13|30|Manasse, a Mahanaim universam Basan, cunctum regnum Og regis Basan omnesque vicos Iair, qui sunt in Basan, sexaginta oppida;
JOSH|13|31|et dimidiam partem Galaad et Astharoth et Edrai, urbes regni Og in Basan, filiis Machir filii Manasse, dimidiae parti filiorum Machir, iuxta cognationes suas.
JOSH|13|32|Hanc possessionem divisit Moyses in campestribus Moab trans Iordanem contra Iericho ad orientalem plagam.
JOSH|13|33|Tribui autem Levi non dedit possessionem, quoniam Dominus, Deus Israel, ipse est possessio eius, ut locutus est illi.
JOSH|14|1|Hoc est, quod hereditave runt filii Israel in terra Cha naan, quod dederunt eis Eleazar sacerdos et Iosue filius Nun et principes familiarum tribuum Israel,
JOSH|14|2|sorte omnia dividentes, sicut praeceperat Dominus in manu Moysi, novem tribubus et dimidiae tribui.
JOSH|14|3|Duabus enim tribubus et dimidiae dederat Moyses trans Iordanem possessionem, absque Levitis, quibus nihil dedit inter fratres suos;
JOSH|14|4|sed sunt filii Ioseph in duas divisi tribus, Manasse et Ephraim, nec acceperunt Levitae aliam in terra partem, nisi urbes ad habitandum et suburbana earum ad alenda iumenta et pecora sua.
JOSH|14|5|Sicut praeceperat Dominus Moysi, ita fecerunt filii Israel et diviserunt terram.
JOSH|14|6|Accesserunt itaque filii Iudae ad Iosue in Galgala, locutusque est ad eum Chaleb filius Iephonne Cenezaeus: " Nosti quid locutus sit Dominus ad Moysen hominem Dei de me et te in Cadesbarne.
JOSH|14|7|Quadraginta annorum eram, quando me misit Moyses famulus Domini de Cadesbarne, ut considerarem terram; nuntiavique ei quod mihi verum videbatur.
JOSH|14|8|Fratres autem mei, qui ascenderant mecum, dissolverunt cor populi, et nihilominus ego adimplevi, ut sequerer Dominum Deum meum.
JOSH|14|9|Iuravitque Moyses in die illo dicens: "Terra, quam calcavit pes tuus, erit possessio tua et filiorum tuorum in aeternum, quia adimplevisti, ut sequereris Dominum Deum meum".
JOSH|14|10|Concessit ergo Dominus vitam mihi, sicut pollicitus est, usque in praesentem diem. Quadraginta et quinque anni sunt ex quo locutus est Dominus verbum istud ad Moysen, quando ambulabat Israel per solitudinem; hodie octoginta quinque annorum sum,
JOSH|14|11|sic valens ut eo valebam tempore, quando ad explorandum missus sum; illius in me temporis fortitudo usque hodie perseverat tam ad bellandum quam ad gradiendum.
JOSH|14|12|Da ergo mihi montem istum, quem pollicitus est Dominus die illo, te quoque audiente quod Enacim ibi sunt et urbes magnae atque munitae; si forte sit Dominus mecum, et potuero delere eos, sicut promisit mihi ".
JOSH|14|13|Benedixitque ei Iosue et tradidit Hebron in possessionem;
JOSH|14|14|atque ex eo fuit Hebron Chaleb filio Iephonne Cenezaeo usque in praesentem diem, quia adimplevit, ut sequeretur Dominum, Deum Israel.
JOSH|14|15|Nomen Hebron antea vocabatur Cariatharbe (id est civitas Arbe), hominis maximi inter Enacim. Et terra cessavit a proeliis.
JOSH|15|1|Sors tribus filiorum Iudae per cognationes suas ista fuit: usque ad terminum Edom, ad desertum Sin contra Nageb, usque ad extremam partem australis plagae.
JOSH|15|2|Terminus eius meridionalis a summitate maris Salsissimi et a lingua eius, quae respicit meridiem.
JOSH|15|3|Egrediturque contra ascensum Acrabbim et pertransit in Sin ascenditque in meridie Cadesbarne et pervenit in Esron ascendens ad Addar et vertitur in Carca;
JOSH|15|4|atque inde pertransiens in Asemona pervenit ad torrentem Aegypti; eruntque exitus eius ad mare Magnum: hic erit vobis finis meridianae plagae.
JOSH|15|5|Ab oriente vero terminus erit mare Salsissimum usque ad extrema Iordanis. Terminus aquilonis a lingua maris et ab extremis Iordanis
JOSH|15|6|ascendit in Bethagla et transit ab aquilone Betharaba ascendens ad lapidem Boen filii Ruben
JOSH|15|7|et ascendens ad Dabir de valle Achor et contra aquilonem vergens ad Galiloth (hi sunt circuli), qui sunt ex adverso ascensionis Adommim, quae est ab australi parte torrentis, transit ad aquas, quae vocantur fons Solis, et erunt exitus eius ad fontem Rogel.
JOSH|15|8|Ascenditque per convallem Benennom ex latere Iebusaei ad meridiem - haec est Ierusalem - et inde se erigens ad verticem montis, qui est contra vallem Ennom ad occidentem in extrema parte vallis Raphaim contra aquilonem;
JOSH|15|9|pertransitque a vertice montis usque ad fontem aquae Nephtoa et pervenit usque ad vicos montis Ephron inclinaturque in Baala, quae est Cariathiarim.
JOSH|15|10|Et vergit de Baala contra occidentem usque ad montem Seir transitque iuxta latus montis Iarim ad aquilonem - id est Cheslon - et descendit in Bethsames transitque in Thamna
JOSH|15|11|et pervenit ad latus septentrionale Accaron inclinaturque in Sechron et transit montem Baala pervenitque in Iebneel et finitur mari. Terminus occidentalis est mare Magnum.
JOSH|15|12|Hi sunt termini filiorum Iudae per circuitum in cognationibus suis.
JOSH|15|13|Chaleb vero filio Iephonne dedit partem in medio filiorum Iudae, sicut praeceperat Dominus Iosue: Cariatharbe (id est civitas Arbe), patris Enac, ipsa est Hebron.
JOSH|15|14|Delevitque ex ea Chaleb tres filios Enac: Sesai et Ahiman et Tholmai de stirpe Enac.
JOSH|15|15|Atque inde conscendens venit ad habitatores Dabir, quae prius vocabatur Cariathsepher (id est civitas Litterarum).
JOSH|15|16|Dixitque Chaleb: " Qui percusserit Cariathsepher et ceperit eam, dabo illi Axam filiam meam uxorem ".
JOSH|15|17|Cepitque eam Othoniel filius Cenez frater Chaleb, deditque ei Axam filiam suam uxorem.
JOSH|15|18|Quae cum veniret, suasit viro suo, ut peteret a patre suo agrum; descenditque de asino. Cui Chaleb: " Quid habes? ", inquit.
JOSH|15|19|At illa respondit: " Da mihi benedictionem. Terram Nageb arentem dedisti mihi; iunge et irriguam ". Dedit itaque ei Chaleb irriguum superius et inferius.
JOSH|15|20|Haec est possessio tribus filiorum Iudae per cognationes suas.
JOSH|15|21|Erantque civitates ab extremis partibus filiorum Iudae iuxta terminos Edom in Nageb: Cabseel et Eder et Iagur
JOSH|15|22|et Cina et Dimona et Adada
JOSH|15|23|et Cades et Asor et Iethnan,
JOSH|15|24|Ziph et Telem et Baloth
JOSH|15|25|et Asorhadatta et Carioth, Esron - haec est Asor -
JOSH|15|26|Amam et Sama et Molada
JOSH|15|27|et Asargadda et Hasemon et Bethphelet
JOSH|15|28|et Asarsual et Bersabee et Baziothia,
JOSH|15|29|Baala et Iim et Esem
JOSH|15|30|et Eltholad et Cesil et Horma
JOSH|15|31|et Siceleg et Madmena et Sensenna
JOSH|15|32|et Lebaoth et Selim et Enremmon: omnes civitates viginti novem et villae earum.
JOSH|15|33|In campestribus vero: Esthaol et Saraa et Asena
JOSH|15|34|et Zanoa et Engannim, Thapphua et Enaim,
JOSH|15|35|Ierimoth et Odollam, Socho et Azeca
JOSH|15|36|et Saarim et Adithaim et Gedera et Gederothaim: urbes quattuordecim et villae earum.
JOSH|15|37|Sanan et Hadasa et Magdalgad
JOSH|15|38|et Delean et Maspha et Iecethel,
JOSH|15|39|Lachis et Bascath et Eglon
JOSH|15|40|et Chebbon et Lehemas et Cethlis
JOSH|15|41|et Gederoth, Bethdagon et Naama et Maceda: civitates sedecim et villae earum.
JOSH|15|42|Lobna et Ether et Asan
JOSH|15|43|et Iephtha et Esna et Nesib
JOSH|15|44|et Ceila et Achzib et Maresa: civitates novem et villae earum.
JOSH|15|45|Accaron cum filiabus et villulis suis;
JOSH|15|46|ab Accaron usque ad mare: omnia, quae sunt ad latus Azoti, et viculos eorum,
JOSH|15|47|Azotus cum filiabus et villulis suis, Gaza cum filiabus et villulis suis usque ad torrentem Aegypti, et mare Magnum terminus.
JOSH|15|48|Et in monte: Samir et Iether et Socho
JOSH|15|49|et Danna et Cariathsenna - haec est Dabir -
JOSH|15|50|et Anab et Esthemo et Anim
JOSH|15|51|et Gosen et Helon et Gilo: civitates undecim et villae earum.
JOSH|15|52|Arab et Duma et Esaan
JOSH|15|53|et Ianum et Beththapphua et Apheca
JOSH|15|54|et Ammatha et Cariatharbe - haec est Hebron - et Sior: civitates novem et villae earum.
JOSH|15|55|Maon et Carmel et Ziph et Iutta
JOSH|15|56|et Iezrahel et Iucadam et Zanoa,
JOSH|15|57|Accain, Gabaa et Thamna: civitates decem et villae earum.
JOSH|15|58|Halhul, Bethsur et Gedor
JOSH|15|59|et Mareth et Bethanoth et Eltecon: civitates sex et villae earum. Thecue et Ephratha - haec est Bethlehem - et Phegor et Etam et Culon et Tatam et Sores et Carem et Gallim et Bether et Manahath: civitates undecim et villae earum.
JOSH|15|60|Cariathbaal - haec est Cariathiarim (urbs Silvarum) - et Arebba: civitates duae et villae earum.
JOSH|15|61|In deserto: Betharaba, Meddin et Sachacha
JOSH|15|62|et Nebsan et civitas Salis et Engaddi: civitates sex et villae earum.
JOSH|15|63|Iebusaeum autem habitatorem Ierusalem non potuerunt filii Iudae delere; habitavitque Iebusaeus cum filiis Iudae in Ierusalem usque in praesentem diem.
JOSH|16|1|Cecidit quoque sors filiorum Ioseph ab Iordane contra Ie richo et aquas eius ab oriente, solitudo, quae ascendit de Iericho ad montem Bethel
JOSH|16|2|et egreditur de Bethel Luz transitque per terminum Arachitarum in Ataroth
JOSH|16|3|et descendit ad occidentem ad terminum Iephlethi usque ad terminos Bethoron inferioris et Gazer; finiunturque regiones eius mari Magno.
JOSH|16|4|Hereditaverunt illas filii Ioseph Manasses et Ephraim.
JOSH|16|5|Et factus est terminus filiorum Ephraim per cognationes suas et possessio eorum contra orientem Atarothaddar usque Bethoron superiorem;
JOSH|16|6|egrediunturque confinia in mare, Machmethath vero aquilonem respicit et vertitur terminus contra orientem in Thanathselo et pertransit ab oriente Ianoe.
JOSH|16|7|Descenditque de Ianoe in Ataroth et Naaratha et pervenit in Iericho et egreditur ad Iordanem.
JOSH|16|8|De Thapphua pertransit terminus ad occidentem ad torrentem Cana, suntque egressus eius in mare: haec est possessio tribus filiorum Ephraim per familias suas,
JOSH|16|9|urbesque separatae filiis Ephraim in medio possessionis filiorum Manasse, omnes urbes et villae earum.
JOSH|16|10|Et non interfecerunt filii Ephraim Chananaeum, qui habitabat in Gazer; habitavitque Chananaeus in medio Ephraim usque in diem hanc et factus est tributarius.
JOSH|17|1|Cecidit autem sors tribui Manasse - ipse est enim pri mogenitus Ioseph C; Machir primogenito Manasse patri Galaad, quia fuit vir pugnator, accepit in possessionem Galaad et Basan.
JOSH|17|2|Et reliqui filiorum Manasse acceperunt iuxta familias suas: filii Abiezer et filii Helec et filii Asriel et filii Sechem et filii Hepher et filii Semida: isti sunt filii Manasse filii Ioseph, mares per cognationes suas.
JOSH|17|3|Salphaad vero filio Hepher filii Galaad filii Machir filii Manasse non erant filii, sed solae filiae, quarum ista sunt nomina: Maala et Noa, Hegla et Melcha et Thersa.
JOSH|17|4|Veneruntque in conspectu Eleazari sacerdotis et Iosue filii Nun et principum dicentes: " Dominus praecepit per manum Moysi, ut daretur nobis possessio in medio fratrum nostrorum ". Deditque eis iuxta imperium Domini possessionem in medio fratrum patris earum.
JOSH|17|5|Et ceciderunt funiculi Manasse decem, absque terra Galaad et Basan trans Iordanem.
JOSH|17|6|Filiae enim Manasse acceperunt hereditatem in medio filiorum eius. Terra autem Galaad cecidit in sortem filiorum Manasse, qui reliqui erant.
JOSH|17|7|Fuitque terminus Manasse ab Aser: Machmethath, quae respicit Sichem et egreditur ad dextram in Iasib apud fontem Thapphuae.
JOSH|17|8|Etenim in sorte Manasse ceciderat terra Thapphuae; Thapphua autem ipsa, quae est iuxta terminos Manasse, fuit filiis Ephraim.
JOSH|17|9|Descenditque terminus ad torrentem Cana. In meridie torrentis civitates sunt Ephraim in medio urbium Manasse. Terminus Manasse est ab aquilone torrentis, et exitus eius pergit ad mare,
JOSH|17|10|ita ut ab austro sit possessio Ephraim et ab aquilone Manasse, et utramque claudat mare, et attingunt tribum Aser ab aquilone et tribum Issachar ab oriente.
JOSH|17|11|Fuitque hereditas Manasse in Issachar et in Aser: Bethsan et filiae eius et Ieblaam cum filiabus suis et habitatores Dor cum filiabus suis, habitatores quoque Endor cum filiabus suis; similiterque habitatores Thanach cum filiabus suis et habitatores Mageddo cum filiabus suis et tertia pars regionis Nopheth.
JOSH|17|12|Nec potuerunt filii Manasse has occupare civitates, sed Chananaeus permansit in terra ista.
JOSH|17|13|Postquam autem convaluerunt filii Israel, subiecerunt Chananaeos et fecerunt sibi tributarios nec expulerunt eos.
JOSH|17|14|Locutique sunt filii Ioseph ad Iosue atque dixerunt: " Quare dedisti mihi possessionem sortis et funiculi unius, cum sim tantae multitudinis et benedixerit mihi Dominus? ".
JOSH|17|15|Ad quos Iosue ait: " Si populus multus es, ascende in silvam et succide tibi spatia in terra Pherezaei et Raphaim, quia angusta est tibi possessio montis Ephraim ".
JOSH|17|16|Cui responderunt filii Ioseph: " Montana non sufficiunt nobis, et ferreis curribus utuntur omnes Chananaei, qui habitant in terra campestri, Bethsan cum filiabus suis et illi, qui sunt in planitie Iezrahel ".
JOSH|17|17|Dixitque Iosue ad domum Ioseph, Ephraim et Manasse: "Populus multus es et magnae fortitudinis; non habebis sortem unam,
JOSH|17|18|sed transibis ad montem et succides tibi atque purgabis ad habitandum spatia; et poteris ultra procedere cum subverteris Chananaeum, qui ferreos habet currus et est fortis ".
JOSH|18|1|Congregatique sunt omnes filii Israel in Silo ibique fixe runt tabernaculum conventus, et fuit eis terra subiecta.
JOSH|18|2|Remanserant autem filiorum Israel septem tribus, quae necdum acceperant possessiones suas.
JOSH|18|3|Ad quos Iosue ait: " Usquequo marcetis ignavia et non intratis ad possidendam terram, quam Dominus, Deus patrum vestrorum,dedit vobis?
JOSH|18|4|Eligite de singulis tribubus ternos viros, ut mittam eos, et surgant atque circumeant terram et describant eam iuxta numerum uniuscuiusque multitudinis referantque ad me, quod descripserint.
JOSH|18|5|Dividite vobis terram in septem partes: Iudas sit in terminis suis in australi plaga, et domus Ioseph in aquilone.
JOSH|18|6|Reliquam terram in septem partes describite; et huc afferetis ad me, ut coram Domino Deo nostro mittam vobis hic sortem,
JOSH|18|7|quia non est inter vos pars Levitarum, sed sacerdotium Domini est eorum hereditas. Gad autem et Ruben et dimidia tribus Manasse iam acceperant possessiones suas trans Iordanem ad orientalem plagam, quas dedit eis Moyses famulus Domini ".
JOSH|18|8|Cumque surrexissent viri, ut pergerent ad describendam terram, praecepit eis Iosue dicens: "Circuite terram et describite eam ac revertimini ad me, ut hic coram Domino in Silo mittam vobis sortem ".
JOSH|18|9|Itaque perrexerunt et lustrantes terram secundum urbes in septem partes diviserunt scribentes in volumine; reversique sunt ad Iosue in castra Silo.
JOSH|18|10|Qui misit eis sortes coram Domino in Silo divisitque ibi terram filiis Israel secundum partes eorum.
JOSH|18|11|Et ascendit sors prima filiorum Beniamin per familias suas, ut possiderent terram inter filios Iudae et filios Ioseph.
JOSH|18|12|Fuitque terminus eorum contra aquilonem a Iordane pergens iuxta latus Iericho septentrionalis plagae et inde contra occidentem ad montana conscendens et perveniens in solitudinem Bethaven;
JOSH|18|13|atque pertransiens iuxta Luzam ad meridiem - ipsa est Bethel - descendit in Atarothaddar in montem, qui est ad meridiem Bethoron inferioris,
JOSH|18|14|et inclinatur vergens contra mare ad meridiem a monte, qui respicit Bethoron contra meridiem; suntque exitus eius in Cariathbaal, quae vocatur et Cariathiarim, urbem filiorum Iudae. Haec est plaga ad occidentem.
JOSH|18|15|In plaga autem ad meridiem, ex parte Cariathiarim egreditur terminus in Gasim et pervenit usque ad fontem aquarum Nephtoa
JOSH|18|16|descenditque in extremam partem montis, qui respicit vallem Benennom et est contra septentrionalem plagam in extrema parte vallis Raphaim; descenditque in vallem Ennom, iuxta latus Iebusaei ad austrum, et pervenit ad fontem Rogel
JOSH|18|17|transiens ad aquilonem et egrediens ad Ensemes (id est fontem Solis). Et pertransit usque ad Galiloth (hi sunt circuli), qui sunt e regione ascensus Adommim, descenditque ad Abenboen (id est lapidem Boen) filii Ruben
JOSH|18|18|et pertransit ex latere aquilonis Betharaba descenditque in Arabam.
JOSH|18|19|Et praetergreditur contra aquilonem Bethagla; suntque exitus eius contra linguam maris Salsissimi ab aquilone in fine Iordanis. Haec est australis plaga.
JOSH|18|20|Iordanis autem est terminus ab oriente. Haec est possessio filiorum Beniamin per terminos suos in circuitu secundum familias suas.
JOSH|18|21|Fueruntque civitates eius: Iericho et Bethagla et Ameccasis
JOSH|18|22|et Betharaba et Semaraim et Bethel
JOSH|18|23|et Avim et Phara et Ophra,
JOSH|18|24|Capharemona et Ophni et Gabaa: civitates duodecim et villae earum.
JOSH|18|25|Gabaon et Rama et Beroth
JOSH|18|26|et Maspha et Cephira et Mosa
JOSH|18|27|et Recem, Iaraphel et Tharala
JOSH|18|28|et Sela, Eleph et Iebus, quae est Ierusalem, Gabaath et Cariath: civitates quattuordecim et villae earum. Haec est possessio filiorum Beniamin iuxta familias suas.
JOSH|19|1|Et egressa est sors secunda fi liorum Simeon per cognatio nes suas; fuitque hereditas
JOSH|19|2|eorum in medio possessionis filiorum Iudae. Bersabee et Sama et Molada
JOSH|19|3|et Asarsual et Bala et Esem
JOSH|19|4|et Eltholad et Bethul et Horma
JOSH|19|5|et Siceleg et Bethmarchaboth et Asarsusa
JOSH|19|6|et Bethlebaoth et Sarohen: civitates tredecim et villae earum.
JOSH|19|7|Ain et Remmon et Ethar et Asan: civitates quattuor et villae earum.
JOSH|19|8|Omnes viculi per circuitum urbium istarum usque ad Baalathbeer, Ramathnageb: haec est hereditas filiorum Simeon iuxta cognationes suas.
JOSH|19|9|Sumpta est de funiculo filiorum Iudae, quia maior erat; et idcirco possederunt filii Simeon in medio hereditatis eorum.
JOSH|19|10|Ceciditque sors tertia filiorum Zabulon per cognationes suas. Et factus est terminus possessionis eorum usque Sarid
JOSH|19|11|ascenditque contra occidentem et Merala et pervenit in Debbaseth usque ad torrentem, qui est contra Iecnaam,
JOSH|19|12|et revertitur de Sarid contra orientem in fines Ceseleththabor et egreditur ad Dabereth ascenditque contra Iaphia.
JOSH|19|13|Et inde pertransit usque ad orientalem plagam Gethhepher, Etthacasin et egreditur in Remmon et inclinatur in Noa;
JOSH|19|14|et vergit ad aquilonem ad Hanathon. Suntque egressus eius vallis Iephthael;
JOSH|19|15|et Cateth et Naalol et Semeron et Iedala et Bethlehem: civitates duodecim et villae earum.
JOSH|19|16|Haec est hereditas tribus filiorum Zabulon per cognationes suas, urbes et viculi earum.
JOSH|19|17|Issachar egressa est sors quarta per cognationes suas.
JOSH|19|18|Fuitque eius hereditas Iezrahel et Chasaloth et Sunam
JOSH|19|19|et Hapharaim et Seon et Anaharath
JOSH|19|20|et Rabbith et Cesion et Abes
JOSH|19|21|et Rameth et Engannim et Enhadda et Bethpheses.
JOSH|19|22|Et pervenit terminus eius usque Thabor et Sehesima et Bethsames; suntque exitus eius ad Iordanem; civitates sedecim et villae earum.
JOSH|19|23|Haec est possessio filiorum Issachar per cognationes suas, urbes et viculi earum.
JOSH|19|24|Ceciditque sors quinta tribui filiorum Aser per cognationes suas.
JOSH|19|25|Fuitque terminus eorum Helcath et Chali et Beten et Achsaph
JOSH|19|26|et Elmelech et Amaad et Masal et pervenit usque ad Carmelum in occidente et ad Sihorlabanath;
JOSH|19|27|ac revertitur contra orientem in Bethdagon et pertransit usque Zabulon et vallem Iephthael contra aquilonem in Bethemec et Neiel. Egrediturque ad laevam Chabul
JOSH|19|28|et Abran et Rohob et Hamon et Cana usque ad Sidonem magnam
JOSH|19|29|revertiturque in Rama usque ad civitatem munitissimam Tyrum et revertitur in Hosa; suntque exitus eius in mare; Mahaleb, Achazib
JOSH|19|30|et Amma et Aphec et Rohob: civitates viginti duae et villae earum.
JOSH|19|31|Haec est possessio filiorum Aser per cognationes suas, urbes et viculi earum.
JOSH|19|32|Filiorum Nephthali sexta sors cecidit per familias suas.
JOSH|19|33|Et coepit terminus de Heleph et de quercu in Saananim et Adamineceb et Iebnael usque Lecum et egressus eius usque ad Iordanem;
JOSH|19|34|revertiturque terminus contra occidentem in Aznotthabor atque inde egreditur in Hucoc et attingit Zabulon contra meridiem et Aser contra occidentem et Iordanem contra ortum solis;
JOSH|19|35|civitates munitissimae Assedim, Ser et Ammath, Reccath et Chenereth
JOSH|19|36|et Edema et Rama, Asor
JOSH|19|37|et Cedes et Edrai et Enasor,
JOSH|19|38|Ieron et Magdalel, Horem et Bethanath et Bethsames: civitates decem et novem et villae earum.
JOSH|19|39|Haec est possessio tribus filiorum Nephthali per cognationes suas, urbes et viculi earum.
JOSH|19|40|Tribui filiorum Dan per familias suas egressa est sors septima.
JOSH|19|41|Et fuit terminus possessionis eius Saraa et Esthaol et Hirsemes (id est civitas Solis)
JOSH|19|42|et Selebin et Aialon et Iethela
JOSH|19|43|et Elon et Thamna et Accaron
JOSH|19|44|et Elthece et Gebbethon et Baalath
JOSH|19|45|et Iud et Benebarach et Gethremmon
JOSH|19|46|et Meiarcon et Areccon cum termino, qui respicit Ioppen.
JOSH|19|47|Et terminus filiorum Dan effugit ab eis. Ascenderuntque filii Dan et pugnaverunt contra Lesem ceperuntque eam; et percusserunt in ore gladii ac possederunt et habitaverunt in ea, vocantes Lesemdan ex nomine Dan patris sui.
JOSH|19|48|Haec est possessio tribus filiorum Dan per cognationes suas, urbes et viculi earum.
JOSH|19|49|Cumque complessent terram sorte dividere singulis per tribus suas, dederunt filii Israel possessionem Iosue filio Nun in medio sui,
JOSH|19|50|iuxta praeceptum Domini, urbem quam postulavit: Thamnathsare in monte Ephraim. Et aedificavit civitatem habitavitque in ea.
JOSH|19|51|Hae sunt possessiones, quas sorte diviserunt Eleazar sacerdos et Iosue filius Nun et principes familiarum tribuum filiorum Israel in Silo coram Domino ad ostium tabernaculi conventus; compleveruntque partiri terram.
JOSH|20|1|Et locutus est Dominus ad Iosue dicens: " Loquere filiis Israel et dic eis:
JOSH|20|2|Separate vobis urbes fugitivorum, de quibus locutus sum ad vos per manum Moysi,
JOSH|20|3|ut confugiat ad eas, quicumque animam percusserit per errorem nescius, et possit evadere iram proximi, qui ultor est sanguinis.
JOSH|20|4|Cum ad unam harum confugerit civitatum, stabit ante portam civitatis et loquetur senioribus urbis illius ea, quae se comprobent innocentem; sicque suscipient eum et dabunt ei locum ad habitandum.
JOSH|20|5|Cumque ultor sanguinis eum fuerit persecutus, non tradent in manus eius, quia ignorans percussit proximum suum nec ante biduum triduumve eius probatur inimicus.
JOSH|20|6|Et habitabit in civitate illa, donec stet ante coetum ad iudicium, causam reddens facti sui, donec moriatur sacerdos magnus, qui fuerit in illo tempore. Tunc revertetur homicida et ingredietur civitatem suam et domum suam, de qua fugerat ".
JOSH|20|7|Decreveruntque Cedes in Galilaea montis Nephthali et Sichem in monte Ephraim et Cariatharbe - ipsa est Hebron - in monte Iudae;
JOSH|20|8|et trans Iordanem contra orientalem plagam Iericho statuerunt Bosor, quae sita est in campestri solitudine de tribu Ruben, et Ramoth in Galaad de tribu Gad et Golan in Basan de tribu Manasse.
JOSH|20|9|Hae civitates constitutae sunt cunctis filiis Israel et advenis, qui habitant inter eos, ut fugeret ad eas, qui animam nescius percussisset et non moreretur in manu proximi effusum sanguinem vindicare cupientis, donec staret ante populum expositurus causam suam.
JOSH|21|1|Accesseruntque principes familiarum Levi ad Eleazarum sacerdotem et Iosue filium Nun et ad duces cognationum per singulas tribus filiorum Israel
JOSH|21|2|locutique sunt ad eos in Silo terrae Chanaan atque dixerunt: " Dominus praecepit per manum Moysi, ut darentur nobis urbes ad habitandum et suburbana earum ad alenda iumenta ".
JOSH|21|3|Dederuntque filii Israel Levitis de possessionibus suis, iuxta imperium Domini, civitates illas et suburbana earum.
JOSH|21|4|Egressaque est sors in familias Caath: et acceperunt filii Aaron sacerdotis de tribubus Iudae et Simeon et Beniamin civitates tredecim.
JOSH|21|5|Et reliqui filiorum Caath, id est Levitae, acceperunt de tribubus Ephraim et Dan et dimidia tribu Manasse civitates decem.
JOSH|21|6|Porro filiis Gerson egressa est sors, ut acciperent de tribubus Issachar et Aser et Nephthali dimidiaque tribu Manasse in Basan civitates numero tredecim.
JOSH|21|7|Et filiis Merari per cognationes suas de tribubus Ruben et Gad et Zabulon urbes duodecim.
JOSH|21|8|Dederuntque filii Israel Levitis civitates illas et suburbana earum, sicut praecepit Dominus per manum Moysi, singulis sorte tribuentes.
JOSH|21|9|De tribubus filiorum Iudae et Simeon dederunt civitates, quarum ista sunt nomina,
JOSH|21|10|filiis Aaron ex familiis Caath levitici generis - prima enim sors illis egressa est C:
JOSH|21|11|Cariatharbe (id est civitas Arbe), patris Enac, quae vocatur Hebron, in monte Iudae et suburbana eius per circuitum.
JOSH|21|12|Agros vero et villas eius dederant Chaleb filio Iephonne ad possidendum.
JOSH|21|13|Dederunt ergo filiis Aaron sacerdotis Hebron confugii civitatem ac suburbana eius et Lobnam cum suburbanis suis
JOSH|21|14|et Iether et Esthemo
JOSH|21|15|et Helon et Dabir
JOSH|21|16|et Ain et Iutta et Bethsames cum suburbanis suis: civitates novem de tribubus illis duabus.
JOSH|21|17|De tribu autem Beniamin Gabaon et Gabaa
JOSH|21|18|et Anathoth et Almath cum suburbanis suis: civitates quattuor.
JOSH|21|19|Omnes simul civitates filiorum Aaron sacerdotis tredecim cum suburbanis suis.
JOSH|21|20|Reliquis vero ex familiis filiorum Caath Levitis haec est data possessio:
JOSH|21|21|de tribu Ephraim urbs confugii Sichem cum suburbanis suis in monte Ephraim et Gazer
JOSH|21|22|et Cibsaim et Bethoron cum suburbanis suis: civitates quattuor.
JOSH|21|23|De tribu quoque Dan Elthece et Gebbethon
JOSH|21|24|et Aialon et Gethremmon cum suburbanis suis: civitates quattuor.
JOSH|21|25|Porro de dimidia tribu Manasse Thanach et Gethremmon cum suburbanis suis: civitates duae.
JOSH|21|26|Omnes civitates decem et suburbana earum datae sunt filiis Caath inferioris gradus.
JOSH|21|27|Filiis quoque Gerson levitici generis dederunt de dimidia tribu Manasse confugii civitatem Golan in Basan et Astharoth cum suburbanis suis: civitates duas.
JOSH|21|28|Porro de tribu Issachar Cesion et Dabereth
JOSH|21|29|et Iaramoth et Engannim cum suburbanis suis: civitates quattuor.
JOSH|21|30|De tribu autem Aser Masal et Abdon
JOSH|21|31|et Helcath et Rohob cum suburbanis suis: civitates quattuor.
JOSH|21|32|De tribu quoque Nephthali civitas confugii Cedes in Galilaea et Ammothdor et Carthan cum suburbanis suis: civitates tres.
JOSH|21|33|Omnes urbes familiarum Gerson tredecim cum suburbanis suis.
JOSH|21|34|Filiis autem Merari Levitis inferioris gradus per familias suas data est de tribu Zabulon Iecnaam et Cartha
JOSH|21|35|et Remmon et Naalol: civitates quattuor cum suburbanis suis.
JOSH|21|36|De tribu Ruben ultra Iordanem contra Iericho civitas refugii Bosor in solitudine planitiei et Iasa
JOSH|21|37|et Cademoth et Mephaath: civitates quattuor cum suburbanis suis.
JOSH|21|38|Et de tribu Gad civitas confugii Ramoth in Galaad et Mahanaim
JOSH|21|39|et Hesebon et Iazer: civitates quattuor cum suburbanis suis.
JOSH|21|40|Omnes urbes filiorum Merari per familias reliquas de cognationibus Levitarum duodecim.
JOSH|21|41|Itaque universae civitates Levitarum in medio possessionis filiorum Israel fuerunt quadraginta octo
JOSH|21|42|cum suburbanis suis, singulae cum suburbanis suis in circuitu.
JOSH|21|43|Deditque Dominus Israeli omnem terram, quam traditurum se patribus eorum iuraverat, et possederunt illam atque habitaverunt in ea.
JOSH|21|44|Deditque Dominus eis requiem secundum omnia, quae iuraverat patribus eorum, nullusque eis hostium resistere ausus est, sed cunctos in eorum dicionem redegit.
JOSH|21|45|Ne unum quidem verbum bonum, quod locutus est ad domum Israel, irritum fuit, sed rebus expleta sunt omnia.
JOSH|22|1|Tunc vocavit Iosue Rubenitas et Gaditas et dimidiam tribum Manasse
JOSH|22|2|dixitque ad eos: "Fecistis omnia, quae vobis praecepit Moyses famulus Domini; mihi quoque in omnibus, quae praecepi vobis, oboedistis
JOSH|22|3|nec reliquistis fratres vestros hoc longo tempore usque in praesentem diem custodientes imperium Domini Dei vestri.
JOSH|22|4|Quia igitur dedit Dominus Deus vester fratribus vestris quietem ac pacem, sicut eis pollicitus est, revertimini nunc et ite in tabernacula vestra et in terram possessionis, quam tradidit vobis Moyses famulus Domini trans Iordanem;
JOSH|22|5|ita dumtaxat ut custodiatis attente et opere compleatis mandatum et legem, quam praecepit vobis Moyses servus Domini, ut diligatis Dominum Deum vestrum et ambuletis in omnibus viis eius et observetis mandata illius adhaereatisque ei ac serviatis in omni corde et in omni anima vestra ".
JOSH|22|6|Benedixitque eis Iosue et dimisit eos, qui reversi sunt in tabernacula sua.
JOSH|22|7|Dimidiae autem tribui Manasse possessionem Moyses dederat in Basan; et idcirco mediae, quae superfuit, dedit Iosue sortem inter ceteros fratres suos trans Iordanem ad occidentalem eius plagam. Cumque dimitteret eos in tabernacula sua et benedixisset illis,
JOSH|22|8|dixit ad eos: "Cum multis divitiis revertimini ad sedes vestras, cum argento et auro, aere ac ferro et veste multiplici; dividite praedam hostium cum fratribus vestris ".
JOSH|22|9|Reversique sunt et abierunt filii Ruben et filii Gad et dimidia tribus Manasse a filiis Israel de Silo, quae sita est in Chanaan, ut intrarent Galaad terram possessionis suae, quam obtinuerant iuxta imperium Domini in manu Moysi.
JOSH|22|10|Cumque venissent ad circulos Iordanis in terra Chanaan, aedificaverunt iuxta Iordanem altare ingens aspectu.
JOSH|22|11|Cum audissent filii Israel aedificasse filios Ruben et Gad et dimidiam tribum Manasse altare e regione terrae Chanaan ad Iordanis circulos ex adverso filiorum Israel,
JOSH|22|12|convenerunt omnes in Silo, ut ascenderent et dimicarent contra eos.
JOSH|22|13|Et interim miserunt ad illos in terram Galaad Phinees filium Eleazari sacerdotem
JOSH|22|14|et decem principes cum eo, singulos de tribubus, unusquisque erat caput familiae in cognationibus Israel.
JOSH|22|15|Qui venerunt ad filios Ruben et Gad et dimidiam tribum Manasse in terram Galaad dixeruntque ad eos:
JOSH|22|16|" Haec mandat omnis coetus Domini: Quae est ista transgressio? Cur reliquistis Dominum, Deum Israel, aedificantes vobis altare sacrilegum et a cultu illius recedentes?
JOSH|22|17|An parum vobis est peccatum Phegor, et usque in praesentem diem macula huius sceleris in nobis permanet, et facta est plaga in coetu Domini?
JOSH|22|18|Et vos hodie reliquistis Dominum, et factum est ut rebellaretis contra Dominum; et cras in universum coetum Israel eius ira desaeviet.
JOSH|22|19|Quod si putatis immundam esse terram possessionis vestrae, transite ad terram possessionis Domini, in qua habitaculum Domini est, et habitate inter nos; tantum ut contra Dominum non rebelletis nec nos rebellare faciatis aedificantes altare praeter altare Domini Dei nostri.
JOSH|22|20|Nonne Achan filius Zarae praeteriit mandatum Domini de anathemate, et super omnem coetum Israel ira Domini incubuit? Et ille erat unus homo; atque utinam solus perisset in scelere suo! ".
JOSH|22|21|Responderuntque filii Ruben et Gad et dimidia tribus Manasse principibus legationis Israel:
JOSH|22|22|" Fortissimus Deus Dominus, fortissimus Deus Dominus ipse novit, et Israel simul intelleget: si rebellionis, si praevaricationis animo contra Dominum hoc altare construximus, non salvet nos, sed puniat in praesenti;
JOSH|22|23|et si ea mente fecimus, ut recedamus a Domino et holocausta et oblationes et pacificas victimas super eo imponeremus, Dominus ipse quaerat et iudicet;
JOSH|22|24|et si non ea magis sollicitudine et cogitatione fecimus hoc dicentes: Cras dicent filii vestri filiis nostris: "Quid vobis et Domino, Deo Israel?
JOSH|22|25|Terminum posuit Dominus inter nos et vos, o filii Ruben et filii Gad, Iordanem fluvium, et idcirco partem non habetis in Domino"; et per hanc occasionem avertent filii vestri filios nostros a timore Domini. Putavimus itaque melius
JOSH|22|26|et diximus: Exstruamus nobis altare non in holocausta neque ad victimas offerendas,
JOSH|22|27|sed in testimonium inter nos et vos et sobolem nostram vestramque progeniem, ut serviamus Domino, et iuris nostri sit offerre holocausta et victimas et pacificas hostias, et nequaquam dicant cras filii vestri filiis nostris: "Non est vobis pars in Domino".
JOSH|22|28|Quod si voluerint dicere, respondebunt eis: "Ecce similitudo altaris Domini, quam fecerunt patres nostri non in holocausta neque in sacrificia, sed in testimonium inter nos et vos".
JOSH|22|29|Absit a nobis hoc scelus, ut recedamus a Domino et eius vestigia relinquamus, exstructo altari ad holocausta et oblationes et victimas offerendas, praeter altare Domini Dei nostri, quod est ante habitaculum eius ".
JOSH|22|30|Quibus auditis, Phinees sacerdos et principes legationis Israel, qui erant cum eo, placati sunt et verba filiorum Ruben et Gad et dimidiae tribus Manasse libentissime susceperunt;
JOSH|22|31|dixitque Phinees filius Eleazar sacerdos ad eos: " Nunc scimus quod nobiscum sit Dominus, quoniam alieni estis a praevaricatione hac et liberastis filios Israel de manu Domini ".
JOSH|22|32|Reversusque est cum principibus a filiis Ruben et Gad de terra Galaad in terram Chanaan ad filios Israel et rettulit eis.
JOSH|22|33|Placuitque sermo cunctis audientibus, et laudaverunt Deum filii Israel; et nequaquam ultra dixerunt, ut ascenderent contra eos in bellum et delerent terram, in qua habitabant filii Ruben et Gad.
JOSH|22|34|Vocaveruntque filii Ruben et filii Gad altare, quod exstruxerant, Testem; dixerunt enim: " Testis est inter nos quod Dominus ipse sit Deus.
JOSH|23|1|Evoluto autem multo tem pore, postquam pacem Do minus dederat Israeli ab omnibus in gyro nationibus et Iosue iam longaevo et persenilis aetatis,
JOSH|23|2|vocavit Iosue omnem Israelem maioresque natu et principes ac iudices et praefectos dixitque ad eos: " Ego senui et progressioris aetatis sum,
JOSH|23|3|vosque vidistis omnia, quae fecerit Dominus Deus vester cunctis nationibus istis, quomodo pro vobis ipse pugnaverit.
JOSH|23|4|Videte, sorte divisi vobis gentes, quae supersunt, in possessionem tribuum vestrarum, sicut omnes, quas delevi, a Iordane usque ad mare Magnum in occidente.
JOSH|23|5|Dominus Deus vester disperdet eas et auferet a facie vestra, et possidebitis terram eorum, sicut vobis pollicitus est.
JOSH|23|6|Tantum confortamini, ut custodiatis cuncta, quae scripta sunt in volumine legis Moysi, et non declinetis ab eis nec ad dexteram nec ad sinistram;
JOSH|23|7|ne conveniatis cum gentibus, quae inter vos residuae sunt, et iuretis in nomine deorum earum et serviatis eis et adoretis illos;
JOSH|23|8|sed adhaereatis Domino Deo vestro, quod fecistis usque in diem hanc.
JOSH|23|9|Et expulit Dominus in conspectu vestro gentes magnas et robustissimas, et nullus vobis resistere potuit:
JOSH|23|10|unus e vobis persequitur hostium mille viros, quia Dominus Deus vester pro vobis ipse pugnat, sicut pollicitus est;
JOSH|23|11|hoc tantum diligentissime praecavete, ut diligatis Dominum Deum vestrum.
JOSH|23|12|Quod si volueritis gentium harum, quae inter vos residuae sunt, erroribus adhaerere et cum eis miscere conubia atque amicitias copulare,
JOSH|23|13|iam nunc scitote quod Dominus Deus vester non eas deleat ante faciem vestram; sed sint vobis in rete, foveam ac laqueum et flagellum ex latere vestro, et spinae in oculis vestris, donec vos disperdat de terra hac optima, quam tradidit vobis.
JOSH|23|14|En ego hodie ingredior viam universae terrae; et toto animo cognoscetis quod de omnibus verbis bonis, quae Dominus Deus vester locutus est vobis, non praeterierit ne unum quidem incassum.
JOSH|23|15|Sicut ergo implevit opere, quod promisit, et prospera cuncta venerunt, sic adducet super vos quidquid malorum comminatus est, donec vos disperdat de terra hac optima, quam tradidit vobis.
JOSH|23|16|Si praeterieritis pactum Domini Dei vestri, quod mandavit vobis, et servieritis diis alienis et adoraveritis eos, consurget in vos furor Domini, et cito peribitis ab hac terra optima, quam tradidit vobis ".
JOSH|24|1|Congregavitque Iosue omnes tribus Israel in Sichem et vocavit maiores natu ac principes et iudices et praefectos, steteruntque in conspectu Dei;
JOSH|24|2|et ad totum populum sic locutus est: " Haec dicit Dominus, Deus Israel: Trans fluvium habitaverunt patres vestri ab initio, Thare pater Abraham et Nachor, servieruntque diis alienis.
JOSH|24|3|Tuli ergo patrem vestrum Abraham de Mesopotamiae finibus et adduxi eum per totam terram Chanaan multiplicavique semen eius.
JOSH|24|4|Et dedi ei Isaac illique rursum dedi Iacob et Esau; e quibus Esau dedi montem Seir ad possidendum, Iacob vero et filii eius descenderunt in Aegyptum.
JOSH|24|5|Misique Moysen et Aaron et percussi Aegyptum signis, quae feci in medio eius, et postea eduxi vos.
JOSH|24|6|Eduxique patres vestros de Aegypto, et venistis ad mare. Persecutique sunt Aegyptii patres vestros cum curribus et equitatu usque ad mare Rubrum.
JOSH|24|7|Clamaverunt autem ad Dominum, qui posuit tenebras inter vos et Aegyptios et adduxit super eos mare et operuit illos. Viderunt oculi vestri, quae in Aegypto fecerim; et habitastis in solitudine multo tempore.
JOSH|24|8|Et introduxi vos ad terram Amorraei, qui habitabat trans Iordanem; cumque pugnarent contra vos, tradidi eos in manus vestras, et occupastis terram eorum atque interfecistis illos.
JOSH|24|9|Surrexit autem Balac filius Sephor rex Moab et pugnavit contra Israelem; misitque et vocavit Balaam filium Beor, ut malediceret vobis.
JOSH|24|10|Et ego nolui audire eum, sed e contrario benedixit vobis, et liberavi vos de manu eius.
JOSH|24|11|Transistisque Iordanem et venistis ad Iericho; pugnaveruntque contra vos viri civitatis illius, Amorraeus et Pherezaeus et Chananaeus et Hetthaeus et Gergesaeus et Hevaeus et Iebusaeus; et tradidi illos in manus vestras.
JOSH|24|12|Misique ante vos crabrones, et eiecerunt eos coram vobis - duos reges Amorraeorum - non in gladio nec in arcu tuo.
JOSH|24|13|Dedique vobis terram, de qua non laborastis, et urbes, quas non aedificastis, et habitatis in eis, vineas et oliveta, quae non plantastis, et manducatis ex eis.
JOSH|24|14|Nunc ergo timete Dominum et servite ei perfecto corde atque verissimo; et auferte deos, quibus servierunt patres vestri in Mesopotamia et in Aegypto, ac servite Domino.
JOSH|24|15|Sin autem malum vobis videtur, ut Domino serviatis, eligite vobis hodie, cui servire vultis, utrum diis, quibus servierunt patres vestri in Mesopotamia, an diis Amorraeorum, in quorum terra habitatis. Ego autem et domus mea serviemus Domino ".
JOSH|24|16|Responditque populus et ait: " Absit a nobis, ut relinquamus Dominum et serviamus diis alienis.
JOSH|24|17|Dominus Deus noster ipse eduxit nos et patres nostros de terra Aegypti, de domo servitutis; fecitque videntibus nobis signa ingentia et custodivit nos in omni via, per quam ambulavimus, et in cunctis populis, per quos transivimus;
JOSH|24|18|et eiecit universas gentes, Amorraeum habitatorem terrae, quam nos intravimus. Serviemus igitur etiam nos Domino, quia ipse est Deus noster.
JOSH|24|19|Dixitque Iosue ad populum: " Non poteritis servire Domino. Deus enim sanctus et Deus aemulator est nec ignoscet sceleribus vestris atque peccatis.
JOSH|24|20|Si dimiseritis Dominum et servieritis diis alienis, convertet se et affliget vos atque subvertet, postquam vobis praestiterit bona ".
JOSH|24|21|Dixitque populus ad Iosue: " Nequaquam, sed Domino serviemus ".
JOSH|24|22|Et Iosue ad populum: " Testes, inquit, vos estis contra vos quia ipsi elegeritis vobis Dominum, ut serviatis ei ". Responderuntque: " Testes ".
JOSH|24|23|" Nunc ergo, ait, auferte deos alienos de medio vestri et inclinate corda vestra ad Dominum, Deum Israel".
JOSH|24|24|Dixitque populus ad Iosue: "Domino Deo nostro serviemus; oboedientes erimus praeceptis eius ".
JOSH|24|25|Percussit igitur Iosue in die illo foedus populo et proposuit ei praecepta atque iudicia in Sichem.
JOSH|24|26|Scripsitque verba haec in volumine legis Dei; et tulit lapidem pergrandem posuitque eum ibi subter quercum, quae erat in sanctuario Domini,
JOSH|24|27|et dixit ad omnem populum: " En lapis iste erit adversus vos in testimonium quia audivit omnia verba Domini, quae locutus est inter nos, ne forte postea negare velitis et mentiri Domino Deo vestro ".
JOSH|24|28|Dimisitque populum, singulos in possessionem suam.
JOSH|24|29|Et post haec mortuus est Iosue filius Nun, servus Domini, centum decem annorum.
JOSH|24|30|Sepelieruntque eum in finibus possessionis suae in Thamnathsare, quae sita est in monte Ephraim a septentrionali parte montis Gaas.
JOSH|24|31|Servivitque Israel Domino cunctis diebus Iosue et seniorum, qui longo vixerunt tempore post Iosue et qui noverunt omnia opera Domini, quae fecerat Israel.
JOSH|24|32|Ossa quoque Ioseph, quae tulerant filii Israel de Aegypto, sepelierunt in Sichem, in parte agri, quem emerat Iacob a filiis Hemmor patris Sichem centum argenteis, et fuit in possessionem filiorum Ioseph.
JOSH|24|33|Eleazar quoque filius Aaron mortuus est; et sepelierunt eum in Gabaa Phinees filii eius, quae data est ei in monte Ephraim.
