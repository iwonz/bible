NAH|1|1|The burden of Nineveh. The book of the vision of Nahum the Elkoshite.
NAH|1|2|God is jealous, and the LORD revengeth; the LORD revengeth, and is furious; the LORD will take vengeance on his adversaries, and he reserveth wrath for his enemies.
NAH|1|3|The LORD is slow to anger, and great in power, and will not at all acquit the wicked: the LORD hath his way in the whirlwind and in the storm, and the clouds are the dust of his feet.
NAH|1|4|He rebuketh the sea, and maketh it dry, and drieth up all the rivers: Bashan languisheth, and Carmel, and the flower of Lebanon languisheth.
NAH|1|5|The mountains quake at him, and the hills melt, and the earth is burned at his presence, yea, the world, and all that dwell therein.
NAH|1|6|Who can stand before his indignation? and who can abide in the fierceness of his anger? his fury is poured out like fire, and the rocks are thrown down by him.
NAH|1|7|The LORD is good, a strong hold in the day of trouble; and he knoweth them that trust in him.
NAH|1|8|But with an overrunning flood he will make an utter end of the place thereof, and darkness shall pursue his enemies.
NAH|1|9|What do ye imagine against the LORD? he will make an utter end: affliction shall not rise up the second time.
NAH|1|10|For while they be folden together as thorns, and while they are drunken as drunkards, they shall be devoured as stubble fully dry.
NAH|1|11|There is one come out of thee, that imagineth evil against the LORD, a wicked counsellor.
NAH|1|12|Thus saith the LORD; Though they be quiet, and likewise many, yet thus shall they be cut down, when he shall pass through. Though I have afflicted thee, I will afflict thee no more.
NAH|1|13|For now will I break his yoke from off thee, and will burst thy bonds in sunder.
NAH|1|14|And the LORD hath given a commandment concerning thee, that no more of thy name be sown: out of the house of thy gods will I cut off the graven image and the molten image: I will make thy grave; for thou art vile.
NAH|1|15|Behold upon the mountains the feet of him that bringeth good tidings, that publisheth peace! O Judah, keep thy solemn feasts, perform thy vows: for the wicked shall no more pass through thee; he is utterly cut off.
NAH|2|1|He that dasheth in pieces is come up before thy face: keep the munition, watch the way, make thy loins strong, fortify thy power mightily.
NAH|2|2|For the LORD hath turned away the excellency of Jacob, as the excellency of Israel: for the emptiers have emptied them out, and marred their vine branches.
NAH|2|3|The shield of his mighty men is made red, the valiant men are in scarlet: the chariots shall be with flaming torches in the day of his preparation, and the fir trees shall be terribly shaken.
NAH|2|4|The chariots shall rage in the streets, they shall justle one against another in the broad ways: they shall seem like torches, they shall run like the lightnings.
NAH|2|5|He shall recount his worthies: they shall stumble in their walk; they shall make haste to the wall thereof, and the defence shall be prepared.
NAH|2|6|The gates of the rivers shall be opened, and the palace shall be dissolved.
NAH|2|7|And Huzzab shall be led away captive, she shall be brought up, and her maids shall lead her as with the voice of doves, tabering upon their breasts.
NAH|2|8|But Nineveh is of old like a pool of water: yet they shall flee away. Stand, stand, shall they cry; but none shall look back.
NAH|2|9|Take ye the spoil of silver, take the spoil of gold: for there is none end of the store and glory out of all the pleasant furniture.
NAH|2|10|She is empty, and void, and waste: and the heart melteth, and the knees smite together, and much pain is in all loins, and the faces of them all gather blackness.
NAH|2|11|Where is the dwelling of the lions, and the feedingplace of the young lions, where the lion, even the old lion, walked, and the lion's whelp, and none made them afraid?
NAH|2|12|The lion did tear in pieces enough for his whelps, and strangled for his lionesses, and filled his holes with prey, and his dens with ravin.
NAH|2|13|Behold, I am against thee, saith the LORD of hosts, and I will burn her chariots in the smoke, and the sword shall devour thy young lions: and I will cut off thy prey from the earth, and the voice of thy messengers shall no more be heard.
NAH|3|1|Woe to the bloody city! it is all full of lies and robbery; the prey departeth not;
NAH|3|2|The noise of a whip, and the noise of the rattling of the wheels, and of the pransing horses, and of the jumping chariots.
NAH|3|3|The horseman lifteth up both the bright sword and the glittering spear: and there is a multitude of slain, and a great number of carcases; and there is none end of their corpses; they stumble upon their corpses:
NAH|3|4|Because of the multitude of the whoredoms of the wellfavoured harlot, the mistress of witchcrafts, that selleth nations through her whoredoms, and families through her witchcrafts.
NAH|3|5|Behold, I am against thee, saith the LORD of hosts; and I will discover thy skirts upon thy face, and I will shew the nations thy nakedness, and the kingdoms thy shame.
NAH|3|6|And I will cast abominable filth upon thee, and make thee vile, and will set thee as a gazingstock.
NAH|3|7|And it shall come to pass, that all they that look upon thee shall flee from thee, and say, Nineveh is laid waste: who will bemoan her? whence shall I seek comforters for thee?
NAH|3|8|Art thou better than populous No, that was situate among the rivers, that had the waters round about it, whose rampart was the sea, and her wall was from the sea?
NAH|3|9|Ethiopia and Egypt were her strength, and it was infinite; Put and Lubim were thy helpers.
NAH|3|10|Yet was she carried away, she went into captivity: her young children also were dashed in pieces at the top of all the streets: and they cast lots for her honourable men, and all her great men were bound in chains.
NAH|3|11|Thou also shalt be drunken: thou shalt be hid, thou also shalt seek strength because of the enemy.
NAH|3|12|All thy strong holds shall be like fig trees with the firstripe figs: if they be shaken, they shall even fall into the mouth of the eater.
NAH|3|13|Behold, thy people in the midst of thee are women: the gates of thy land shall be set wide open unto thine enemies: the fire shall devour thy bars.
NAH|3|14|Draw thee waters for the siege, fortify thy strong holds: go into clay, and tread the morter, make strong the brickkiln.
NAH|3|15|There shall the fire devour thee; the sword shall cut thee off, it shall eat thee up like the cankerworm: make thyself many as the cankerworm, make thyself many as the locusts.
NAH|3|16|Thou hast multiplied thy merchants above the stars of heaven: the cankerworm spoileth, and fleeth away.
NAH|3|17|Thy crowned are as the locusts, and thy captains as the great grasshoppers, which camp in the hedges in the cold day, but when the sun ariseth they flee away, and their place is not known where they are.
NAH|3|18|Thy shepherds slumber, O king of Assyria: thy nobles shall dwell in the dust: thy people is scattered upon the mountains, and no man gathereth them.
NAH|3|19|There is no healing of thy bruise; thy wound is grievous: all that hear the bruit of thee shall clap the hands over thee: for upon whom hath not thy wickedness passed continually?
