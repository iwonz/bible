EPH|1|1|奉上帝旨意作基督耶穌使徒的 保羅 ，寫信給在 以弗所 的 眾聖徒，就是在基督耶穌裏忠心的人。
EPH|1|2|願恩惠、平安 從我們的父上帝和主耶穌基督歸給你們！
EPH|1|3|願頌讚歸給我們主耶穌基督的父上帝。他在基督裏曾把天上各樣屬靈的福氣賜給我們。
EPH|1|4|因為他從創世以前，在基督裏揀選了我們，使我們在他面前成為聖潔，沒有瑕疵，滿有愛心。
EPH|1|5|他按著自己旨意所喜悅的 ，預定我們藉著耶穌基督得兒子的名分，
EPH|1|6|使他榮耀的恩典得到稱讚；這恩典是他在愛子裏白白賜給我們的。
EPH|1|7|我們藉著這愛子的血得蒙救贖，過犯得以赦免，這是照他豐富的恩典，
EPH|1|8|充充足足地賞給我們的。他以諸般的智慧聰明，
EPH|1|9|照自己在基督裏所立定的美意，使我們知道他旨意的奧祕，
EPH|1|10|要照著所安排的，在時機成熟的時候，使天上、地上、一切所有的，都在基督裏面同歸於一。
EPH|1|11|我們也在他裏面得了基業；這原是那位隨己意行萬事的上帝照著自己的旨意所預定的，
EPH|1|12|為要使我們，這些首先把希望寄託在基督裏的人，頌讚他的榮耀。
EPH|1|13|在基督裏你們聽見真理的道，就是那使你們得救的福音，你們也信了他，就受了所應許的聖靈為印記。
EPH|1|14|這聖靈是我們得基業的憑據，直等到上帝的子民得救贖，使他的榮耀得到稱讚。
EPH|1|15|因此，我既然聽見你們對主耶穌有信心，對眾聖徒有愛心，
EPH|1|16|就不住地為你們感謝上帝，禱告的時候常常提到你們，
EPH|1|17|求我們主耶穌基督的上帝，榮耀的父，把那賜人智慧和啟示的靈賜給你們，使你們真正認識他，
EPH|1|18|照亮你們心中的眼睛，使你們知道他呼召你們來得的指望是甚麼，他在聖徒中所得榮耀的基業是何等豐盛，
EPH|1|19|並知道他向我們這些信的人所顯的能力是何等浩大，這是照他的大能大力運行的。
EPH|1|20|這大能曾運行在基督身上，使他從死人中復活，又使他在天上坐在自己的右邊，
EPH|1|21|遠超越一切執政的、掌權的、有權能的、統治的和一切有名號的；不但是今世的，連來世的也都超越了。
EPH|1|22|上帝使萬有服在他的腳下，又使他為了教會作萬有之首；
EPH|1|23|教會是他的身體，是那充滿萬有者所充滿的。
EPH|2|1|從前，你們因著自己的過犯罪惡而死了。
EPH|2|2|那時，你們在過犯罪惡中生活，隨從今世的風俗，順服空中掌權者的領袖，就是現今在悖逆的人心中運行的邪靈。
EPH|2|3|我們從前也都生活在他們當中，放縱肉體的私慾，隨著肉體和心中的意念去做，和別人一樣，生來就是該受懲罰的人。
EPH|2|4|然而，上帝有豐富的憐憫，因著他愛我們的大愛，
EPH|2|5|竟在我們因過犯而死了的時候，使我們與基督一同活過來—可見你們得救是本乎恩—
EPH|2|6|他又使我們在基督耶穌裏與他一同復活，一同坐在天上，
EPH|2|7|為要把他極豐富的恩典，就是他在基督耶穌裏向我們所施的恩慈，顯明給後來的世代。
EPH|2|8|你們得救是本乎恩，也因著信；這並不是出於自己，而是上帝所賜的；
EPH|2|9|也不是出於行為，免得有人自誇。
EPH|2|10|我們是他所造之物，在基督耶穌裏創造的，為要使我們行善，就是上帝早已預備好要我們做的。
EPH|2|11|所以，你們要記得：從前你們按肉體是外邦人，是「沒受割禮的」；這名字是那些憑人手在肉身上「受割禮的人」所取的。
EPH|2|12|要記得那時候，你們與基督無關，與 以色列 選民團體隔絕，在所應許的約上是局外人，而且在世上沒有指望，沒有上帝。
EPH|2|13|從前你們是遠離上帝的人，如今卻在基督耶穌裏，靠著他的血，已經得以親近了。
EPH|2|14|因為他自己是我們的和平 ，使雙方合而為一，拆毀了中間隔絕的牆，而且以自己的身體終止了冤仇，
EPH|2|15|廢掉那記在律法上的規條，為要使兩方藉著自己造成一個新人，促成了和平；
EPH|2|16|既在十字架上消滅了冤仇，就藉這十字架使雙方歸為一體，與上帝和好，
EPH|2|17|並且來傳和平的福音給你們遠處的人，也傳和平給那些近處的人，
EPH|2|18|因為我們雙方藉著他，在同一位聖靈裏得以進到父面前。
EPH|2|19|這樣，你們不再是外人或客旅，是與聖徒同國，是上帝家裏的人了，
EPH|2|20|被建造在使徒和先知的根基上，而基督耶穌自己為房角石，
EPH|2|21|靠著他整座房子連接得緊湊，漸漸成為在主裏的聖殿。
EPH|2|22|你們也靠他同被建造，成為上帝藉著聖靈居住的所在。
EPH|3|1|因此，我— 保羅 為你們外邦人作了基督耶穌 囚徒的，替你們祈禱 。
EPH|3|2|想你們必曾聽見上帝賜恩給我，把關切你們的職分託付我，
EPH|3|3|用啟示讓我知道福音的奧祕，正如我以前略略寫過的。
EPH|3|4|你們讀了，就會知道我深深了解基督的奧祕；
EPH|3|5|這奧祕在以前的世代沒有讓人知道，像如今藉著聖靈向他的聖使徒和先知啟示一樣，
EPH|3|6|就是外邦人在基督耶穌裏，藉著福音，得以同為後嗣，同為一體，同為蒙應許的人。
EPH|3|7|我作了這福音的僕役，是照著上帝的恩賜，是照他運行的大能賜給我的。
EPH|3|8|雖然我比眾聖徒中最小的還小，他還賜我這恩典，讓我把基督那測不透的豐富傳給外邦人，
EPH|3|9|又使眾人都明白 甚麼是歷代以來隱藏在創造萬物之上帝裏的奧祕，
EPH|3|10|為要在現今藉著教會使天上執政的、掌權的知道上帝百般的智慧。
EPH|3|11|這是照著上帝在我們主基督耶穌裏所完成的永恆的計劃。
EPH|3|12|我們因信耶穌 ，就在他裏面放膽無懼，滿有自信地進到上帝面前。
EPH|3|13|所以我求你們，不要因我為你們所受的患難喪膽；這原是你們的光榮。
EPH|3|14|因此，我在父面前屈膝—
EPH|3|15|天上地上的各家都是從他得名的－
EPH|3|16|為要他按著他豐盛的榮耀，藉著他的靈，使你們內心的力量剛強起來；
EPH|3|17|又要他使基督因著你們的信住在你們心裏，使你們既在愛中生根立基，
EPH|3|18|能夠和眾聖徒一同明白基督的愛是何等的長、闊、高、深，並知道這愛是超過人的知識所能測度的，為要使你們充滿上帝一切的豐盛。
EPH|3|19|
EPH|3|20|上帝能照著運行在我們心裏的大能充充足足地成就一切，超過我們所求所想的。
EPH|3|21|願他在教會中，並在基督耶穌裏，得著榮耀，直到世世代代，永永遠遠。阿們！
EPH|4|1|我為主作囚徒的勸你們，既然蒙召，行事為人就要與你們所蒙的呼召相稱。
EPH|4|2|凡事要謙虛、溫柔、忍耐，用愛心互相寬容，
EPH|4|3|以和平彼此聯繫，竭力保持聖靈所賜的合一。
EPH|4|4|身體只有一個，聖靈只有一位，正如你們蒙召，是為同有一個指望而蒙召，
EPH|4|5|一主，一信，一洗，
EPH|4|6|一上帝－就是萬人之父，超越萬有之上，貫通萬有，在萬有之中。
EPH|4|7|我們每個人蒙恩都是照基督所量給每個人的恩賜。
EPH|4|8|所以有話說： 「他升上高天的時候，擄掠了俘虜， 將各樣的恩賜賞給人。」
EPH|4|9|既說「他升上」，豈不是指他曾降到地底下嗎？
EPH|4|10|那降下的，就是高升遠超越諸天之上的，為要充滿萬有。
EPH|4|11|他所賜的有使徒，有先知，有傳福音的，有牧者和教師，
EPH|4|12|為要裝備聖徒，做事奉的工作，建立基督的身體，
EPH|4|13|直等到我們眾人在信仰上同歸於一，認識上帝的兒子，得以長大成人，達到基督完全長成的身量。
EPH|4|14|這樣，我們不再作小孩子，中了人的詭計和欺騙的法術，被一切邪說之風搖動，飄來飄去。
EPH|4|15|我們反而要用愛心說誠實話，各方面向著基督長進，連於元首基督，
EPH|4|16|靠著他全身都連接得緊湊，百節各按各職，照著各體的功用彼此相助，使身體漸漸增長，在愛中建立自己。
EPH|4|17|所以我這樣說，且在主裏鄭重地說，你們行事為人，不要再像外邦人存虛妄的心而活。
EPH|4|18|他們心地昏昧，因自己無知，心裏剛硬而與上帝所賜的生命隔絕了。
EPH|4|19|既然他們已經麻木，就放縱情慾，貪婪地行種種污穢的事。
EPH|4|20|但你們從基督學的不是這樣。
EPH|4|21|如果你們聽過他的道，領了他的教，因為真理就在耶穌裏，
EPH|4|22|你們要脫去從前的行為，脫去舊我；這舊我是因私慾的迷惑而漸漸敗壞的。
EPH|4|23|你們要把自己的心志更新，
EPH|4|24|並且穿上新我；這新我是照著上帝的形像造的，有從真理來的公義和聖潔。
EPH|4|25|所以，你們要棄絕謊言，每個人要與鄰舍說誠實話，因為我們是互為肢體。
EPH|4|26|即使生氣也不要犯罪；不可含怒到日落，
EPH|4|27|不可給魔鬼留地步。
EPH|4|28|偷竊的，不要再偷；總要勤勞，親手 做正當的事，這樣才可以把自己有的，分給有缺乏的人。
EPH|4|29|一句壞話也不可出口，只要隨著需要說造就人的好話，讓聽見的人得益處。
EPH|4|30|不要使上帝的聖靈擔憂，你們原是受了他的印記，等候得救贖的日子來到。
EPH|4|31|一切苦毒、憤怒、惱恨、嚷鬧、毀謗，和一切的惡毒都要從你們中間除掉。
EPH|4|32|要仁慈相待，存憐憫的心，彼此饒恕，正如上帝在基督裏饒恕了你們一樣。
EPH|5|1|所以，作為蒙慈愛的兒女，你們該效法上帝。
EPH|5|2|要憑愛心行事，正如基督愛我們，為我們捨了自己，當作馨香的供物和祭物獻給上帝。
EPH|5|3|至於淫亂和一切污穢，或是貪婪，在你們中間連提都不可，這才合乎聖徒的體統。
EPH|5|4|淫詞、妄語和粗俗的俏皮話都不合宜；總要說感謝的話。
EPH|5|5|要確實知道，無論是淫亂的，是污穢的，是貪心的（貪心的就是拜偶像的），在基督和上帝的國裏都得不到基業。
EPH|5|6|不要被人虛浮的話欺騙了，因這些事，上帝的憤怒必臨到那些悖逆的人。
EPH|5|7|所以，不要與他們同夥。
EPH|5|8|從前你們是暗昧的，但如今在主裏面是光明的，行事為人要像光明的子女—
EPH|5|9|光明所結的果子就是一切的良善、公義、誠實。
EPH|5|10|總要察驗甚麼是主所喜悅的事。
EPH|5|11|那暗昧無益的事，不可參與，倒要把這種事揭發出來。
EPH|5|12|因為，他們暗中所做的，就是連提起來都是可恥的。
EPH|5|13|凡被光所照明的都顯露出來，
EPH|5|14|因為使一切顯露出來的就是光。所以有話說： 「你這睡著的人醒過來吧！ 要從死人中復活， 基督要光照你了。」
EPH|5|15|你們要謹慎行事，不要像無知的人，要像智慧的人。
EPH|5|16|要把握時機 ，因為現今的世代邪惡。
EPH|5|17|不要作糊塗人，要明白主的旨意如何。
EPH|5|18|不要醉酒，酒能使人放蕩；要被聖靈充滿。
EPH|5|19|要用詩篇、讚美詩、靈歌彼此對說，口唱心和地讚美主。
EPH|5|20|凡事要奉我們主耶穌基督的名常常感謝父上帝。
EPH|5|21|要存敬畏基督的心彼此順服。
EPH|5|22|作妻子的，你們要順服自己的丈夫，如同順服主。
EPH|5|23|因為丈夫是妻子的頭，如同基督是教會的頭；他又是這身體的救主。
EPH|5|24|教會怎樣順服基督，妻子也要怎樣凡事順服丈夫。
EPH|5|25|作丈夫的，你們要愛自己的妻子，正如基督愛教會，為教會捨己，
EPH|5|26|以水藉著道把教會洗淨，使她成為聖潔，
EPH|5|27|好獻給自己，作榮耀的教會，毫無玷污、皺紋等類的缺陷，而是聖潔沒有瑕疵的。
EPH|5|28|丈夫也應當照樣愛妻子，如同愛自己的身體；愛妻子就是愛自己了。
EPH|5|29|從來沒有人恨惡自己的身體，總是保養愛惜，正像基督待教會一樣，
EPH|5|30|因我們是他身體的肢體。
EPH|5|31|「為這個緣故，人要離開父母，與妻子結合，二人成為一體。」
EPH|5|32|這是極大的奧祕，而我是指基督和教會說的。
EPH|5|33|然而，你們每個人都要愛妻子，如同愛自己一樣；妻子也要敬重她的丈夫。
EPH|6|1|作兒女的，你們要在主裏 聽從父母，這是理所當然的。
EPH|6|2|當孝敬父母，使你得福，在世長壽。這是第一條帶應許的誡命。
EPH|6|3|
EPH|6|4|作父親的，你們不要激怒兒女，但要照著主的教導和勸戒養育他們。
EPH|6|5|作僕人的，你們要懼怕戰兢，用誠實的心聽從你們肉身的主人，好像聽從基督一般；
EPH|6|6|不要只在人的眼前這樣做，像僅是討人的喜歡，而是作基督的僕人，從心裏遵行上帝的旨意，
EPH|6|7|甘心服侍，好像服侍主，不像服侍人，
EPH|6|8|因為知道每個人所做的善事，不論是為奴的或是自主的，都必按所做的從主得到賞賜。
EPH|6|9|作主人的，你們待僕人也是一樣，不要威嚇他們，因為知道他們和你們在天上同有一位主，他並不偏待人。
EPH|6|10|最後，你們要靠著主，依賴他的大能大力作剛強的人。
EPH|6|11|要穿戴上帝所賜的全副軍裝，好抵擋魔鬼的詭計。
EPH|6|12|因為我們的爭戰並不是對抗有血有肉的人，而是對抗那些執政的、掌權的、管轄這幽暗世界的，以及天空靈界的惡魔。
EPH|6|13|所以，要拿起上帝所賜的全副軍裝，好在邪惡的日子能抵擋仇敵，並且完成了一切後還能站立得住。
EPH|6|14|所以，要站穩了，用真理當作帶子束腰，用公義當作護心鏡遮胸，
EPH|6|15|又用和平的福音當作預備走路的鞋穿在腳上。
EPH|6|16|此外，要拿信德當作盾牌，用來撲滅那惡者一切燒著的箭。
EPH|6|17|要戴上救恩的頭盔，拿著聖靈的寶劍—就是上帝的道。
EPH|6|18|要靠著聖靈，隨時多方禱告祈求，並要為此警醒不倦，為眾聖徒祈求。
EPH|6|19|也要為我祈求，讓我有口才，能放膽開口講明福音的奧祕，
EPH|6|20|我為這福音的奧祕作了帶鐵鏈的使者，讓我能照著當盡的本分放膽宣講。
EPH|6|21|今有親愛、忠心服事主的弟兄 推基古 ，為了你們也明白我的事情和我的景況，他會讓你們知道一切的事。
EPH|6|22|我特意打發他到你們那裏去，好讓你們知道我們的情況，又讓他安慰你們的心。
EPH|6|23|願平安 、慈愛、信心從父上帝和主耶穌基督歸給弟兄們。
EPH|6|24|願所有恆心愛我們主耶穌基督的人都蒙恩惠。
