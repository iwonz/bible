1JOHN|1|1|Quod fuit ab initio, quod audi vimus, quod vidimus oculis no stris, quod perspeximus, et manus nostrae contrectaverunt de verbo vitae
1JOHN|1|2|- et vita apparuit, et vidimus et testamur et annuntiamus vobis vitam aeternam, quae erat coram Patre et apparuit nobis -
1JOHN|1|3|quod vidimus et audivimus, annuntiamus et vobis, ut et vos communionem habeatis nobiscum. Communio autem nostra est cum Patre et cum Filio eius Iesu Christo.
1JOHN|1|4|Et haec scribimus nos, ut gaudium nostrum sit plenum.
1JOHN|1|5|Et haec est annuntiatio, quam audivimus ab eo et annuntiamus vobis, quoniam Deus lux est, et tenebrae in eo non sunt ullae.
1JOHN|1|6|Si dixerimus quoniam communionem habemus cum eo, et in tenebris ambulamus, mentimur et non facimus veritatem;
1JOHN|1|7|si autem in luce ambulemus, sicut ipse est in luce, communionem habemus ad invicem, et sanguis Iesu Filii eius mundat nos ab omni peccato.
1JOHN|1|8|Si dixerimus quoniam peccatum non habemus, nosmetipsos seducimus, et veritas in nobis non est.
1JOHN|1|9|Si confiteamur peccata nostra, fidelis est et iustus, ut remittat nobis peccata et emundet nos ab omni iniustitia.
1JOHN|1|10|Si dixerimus quoniam non peccavimus, mendacem facimus eum, et verbum eius non est in nobis.
1JOHN|2|1|Filioli mei, haec scribo vobis, ut non peccetis. Sed si quis pecca verit, advocatum habemus ad Patrem, Iesum Christum iustum;
1JOHN|2|2|et ipse est propitiatio pro peccatis nostris, non pro nostris autem tantum sed etiam pro totius mundi.
1JOHN|2|3|Et in hoc cognoscimus quoniam novimus eum: si mandata eius servemus.
1JOHN|2|4|Qui dicit: " Novi eum ", et mandata eius non servat, mendax est, et in isto veritas non est;
1JOHN|2|5|qui autem servat verbum eius, vere in hoc caritas Dei consummata est. In hoc cognoscimus quoniam in ipso sumus.
1JOHN|2|6|Qui dicit se in ipso manere, debet, sicut ille ambulavit, et ipse ambulare.
1JOHN|2|7|Carissimi, non mandatum novum scribo vobis sed mandatum vetus, quod habuistis ab initio: mandatum vetus est verbum, quod audistis.
1JOHN|2|8|Verumtamen mandatum novum scribo vobis, quod est verum in ipso et in vobis, quoniam tenebrae transeunt, et lumen verum iam lucet.
1JOHN|2|9|Qui dicit se in luce esse, et fratrem suum odit, in tenebris est usque adhuc.
1JOHN|2|10|Qui diligit fratrem suum, in lumine manet, et scandalum ei non est;
1JOHN|2|11|qui autem odit fratrem suum, in tenebris est et in tenebris ambulat et nescit quo vadat, quoniam tenebrae obcaecaverunt oculos eius.
1JOHN|2|12|Scribo vobis, filioli: Remissa sunt vobis peccata propter nomen eius.
1JOHN|2|13|Scribo vobis, patres: Nostis eum, qui ab initio est. Scribo vobis, adulescentes: Vicistis Malignum.
1JOHN|2|14|Scripsi vobis, parvuli: Nostis Patrem. Scripsi vobis, patres: Nostis eum, qui ab initio est. Scripsi vobis, adulescentes: Fortes estis, et verbum Dei in vobis manet, et vicistis Malignum.
1JOHN|2|15|Nolite diligere mundum neque ea, quae in mundo sunt. Si quis diligit mundum, non est caritas Patris in eo;
1JOHN|2|16|quoniam omne, quod est in mundo, concupiscentia carnis et concupiscentia oculorum et iactantia divitiarum, non est ex Patre, sed ex mundo est.
1JOHN|2|17|Et mundus transit, et concupiscentia eius; qui autem facit voluntatem Dei, manet in aeternum.
1JOHN|2|18|Filioli, novissima hora est; et sicut audistis quia antichristus venit, ita nunc antichristi multi adsunt, unde cognoscimus quoniam novissima hora est.
1JOHN|2|19|Ex nobis prodierunt, sed non erant ex nobis, nam si fuissent ex nobis, permansissent nobiscum; sed ut manifestaretur quoniam illi omnes non sunt ex nobis.
1JOHN|2|20|Sed vos unctionem habetis a Sancto et scitis omnes.
1JOHN|2|21|Non scripsi vobis quasi nescientibus veritatem sed quasi scientibus eam, et quoniam omne mendacium ex veritate non est.
1JOHN|2|22|Quis est mendax, nisi is qui negat quoniam Iesus est Christus? Hic est antichristus, qui negat Patrem et Filium.
1JOHN|2|23|Omnis, qui negat Filium, nec Patrem habet; qui confitetur Filium, et Patrem habet.
1JOHN|2|24|Vos, quod audistis ab initio, in vobis permaneat; si in vobis permanserit, quod ab initio audistis, et vos in Filio et in Patre manebitis.
1JOHN|2|25|Et haec est repromissio, quam ipse pollicitus est nobis: vitam aeternam.
1JOHN|2|26|Haec scripsi vobis de eis, qui seducunt vos.
1JOHN|2|27|Et vos, unctionem, quam accepistis ab eo, manet in vobis, et non necesse habetis, ut aliquis doceat vos; sed sicut unctio ipsius docet vos de omnibus, et verum est, et non est mendacium, et, sicut docuit vos, manetis in eo.
1JOHN|2|28|Et nunc, filioli, manete in eo, ut, cum apparuerit, habeamus fiduciam et non confundamur ab eo in adventu eius.
1JOHN|2|29|Si scitis quoniam iustus est, scitote quoniam et omnis, qui facit iustitiam, ex ipso natus est.
1JOHN|3|1|Videte qualem caritatem dedit nobis Pater, ut filii Dei nomine mur, et sumus! Propter hoc mundus non cognoscit nos, quia non cognovit eum.
1JOHN|3|2|Carissimi, nunc filii Dei sumus, et nondum manifestatum est quid erimus; scimus quoniam, cum ipse apparuerit, similes ei erimus, quoniam videbimus eum, sicuti est.
1JOHN|3|3|Et omnis, qui habet spem hanc in eo, purificat se, sicut ille purus est.
1JOHN|3|4|Omnis, qui facit peccatum, et iniquitatem facit, quia peccatum est iniquitas.
1JOHN|3|5|Et scitis quoniam ille apparuit, ut peccata tolleret, et peccatum in eo non est.
1JOHN|3|6|Omnis, qui in eo manet, non peccat; omnis, qui peccat, non vidit eum nec novit eum.
1JOHN|3|7|Filioli, nemo vos seducat. Qui facit iustitiam, iustus est, sicut ille iustus est;
1JOHN|3|8|qui facit peccatum, ex Diabolo est, quoniam a principio Diabolus peccat. Propter hoc apparuit Filius Dei, ut dissolvat opera Diaboli.
1JOHN|3|9|Omnis, qui natus est ex Deo, peccatum non facit, quoniam semen ipsius in eo manet; et non potest peccare, quoniam ex Deo natus est.
1JOHN|3|10|In hoc manifesti sunt filii Dei et filii Diaboli: omnis, qui non facit iustitiam, non est ex Deo, et qui non diligit fratrem suum.
1JOHN|3|11|Quoniam haec est annuntiatio, quam audistis ab initio, ut diligamus alterutrum.
1JOHN|3|12|Non sicut Cain: ex Maligno erat et occidit fratrem suum. Et propter quid occidit eum? Quoniam opera eius maligna erant, fratris autem eius iusta.
1JOHN|3|13|Nolite mirari, fratres, si odit vos mundus.
1JOHN|3|14|Nos scimus quoniam transivimus de morte in vitam, quoniam diligimus fratres; qui non diligit, manet in morte.
1JOHN|3|15|Omnis, qui odit fratrem suum, homicida est, et scitis quoniam omnis homicida non habet vitam aeternam in semetipso manentem.
1JOHN|3|16|In hoc novimus caritatem, quoniam ille pro nobis animam suam posuit; et nos debemus pro fratribus animas ponere.
1JOHN|3|17|Qui habuerit substantiam mundi et viderit fratrem suum necesse habere et clauserit viscera sua ab eo, quomodo caritas Dei manet in eo?
1JOHN|3|18|Filioli, non diligamus verbo nec lingua sed in opere et veritate.
1JOHN|3|19|In hoc cognoscemus quoniam ex veritate sumus, et in conspectu eius placabimus corda nostra,
1JOHN|3|20|quoniam si reprehenderit nos cor, maior est Deus corde nostro et cognoscit omnia.
1JOHN|3|21|Carissimi, si cor nostrum non reprehenderit nos, fiduciam habemus ad Deum
1JOHN|3|22|et, quodcumque petierimus, accipimus ab eo, quoniam mandata eius custodimus et ea, quae sunt placita coram eo, facimus.
1JOHN|3|23|Et hoc est mandatum eius, ut credamus nomini Filii eius Iesu Christi et diligamus alterutrum, sicut dedit mandatum nobis.
1JOHN|3|24|Et, qui servat mandata eius, in ipso manet, et ipse in eo; et in hoc cognoscimus quoniam manet in nobis, ex Spiritu, quem nobis dedit.
1JOHN|4|1|Carissimi, nolite omni spiritui credere, sed probate spiritus si ex Deo sint, quoniam multi pseudoprophetae prodierunt in mundum.
1JOHN|4|2|In hoc cognoscitis Spiritum Dei: omnis spiritus, qui confitetur Iesum Christum in carne venisse, ex Deo est.
1JOHN|4|3|Et omnis spiritus, qui non confitetur Iesum, ex Deo non est; et hoc est antichristi, quod audistis quoniam venit, et nunc iam in mundo est.
1JOHN|4|4|Vos ex Deo estis, filioli, et vicistis eos, quoniam maior est, qui in vobis est, quam qui in mundo.
1JOHN|4|5|Ipsi ex mundo sunt; ideo ex mundo loquuntur, et mundus eos audit.
1JOHN|4|6|Nos ex Deo sumus. Qui cognoscit Deum, audit nos; qui non est ex Deo, non audit nos. Ex hoc cognoscimus Spiritum veritatis et spiritum erroris.
1JOHN|4|7|Carissimi, diligamus invicem, quoniam caritas ex Deo est; et omnis, qui diligit, ex Deo natus est et cognoscit Deum.
1JOHN|4|8|Qui non diligit, non cognovit Deum, quoniam Deus caritas est.
1JOHN|4|9|In hoc apparuit caritas Dei in nobis, quoniam Filium suum unigenitum misit Deus in mundum, ut vivamus per eum.
1JOHN|4|10|In hoc est caritas, non quasi nos dilexerimus Deum, sed quoniam ipse dilexit nos et misit Filium suum propitiationem pro peccatis nostris.
1JOHN|4|11|Carissimi, si sic Deus dilexit nos, et nos debemus alterutrum diligere.
1JOHN|4|12|Deum nemo vidit umquam; si diligamus invicem, Deus in nobis manet, et caritas eius in nobis consummata est.
1JOHN|4|13|In hoc cognoscimus quoniam in ipso manemus, et ipse in nobis, quoniam de Spiritu suo dedit nobis.
1JOHN|4|14|Et nos vidimus et testificamur quoniam Pater misit Filium salvatorem mundi.
1JOHN|4|15|Quisque confessus fuerit: " Iesus est Filius Dei ", Deus in ipso manet, et ipse in Deo.
1JOHN|4|16|Et nos, qui credidimus, novimus caritatem, quam habet Deus in nobis. Deus caritas est; et, qui manet in caritate, in Deo manet, et Deus in eo manet.
1JOHN|4|17|In hoc consummata est caritas nobiscum, ut fiduciam habeamus in die iudicii; quia sicut ille est, et nos sumus in hoc mundo.
1JOHN|4|18|Timor non est in caritate, sed perfecta caritas foras mittit timorem, quoniam timor poenam habet; qui autem timet, non est consummatus in caritate.
1JOHN|4|19|Nos diligimus, quoniam ipse prior dilexit nos.
1JOHN|4|20|Si quis dixerit: " Diligo Deum ", et fratrem suum oderit, mendax est; qui enim non diligit fratrem suum, quem videt, Deum, quem non videt, non potest diligere.
1JOHN|4|21|Et hoc mandatum habemus ab eo, ut, qui diligit Deum, diligat et fratrem suum.
1JOHN|5|1|Omnis, qui credit quoniam Iesus est Christus, ex Deo natus est; et omnis, qui diligit Deum, qui genuit, diligit et eum, qui natus est ex eo.
1JOHN|5|2|In hoc cognoscimus quoniam diligimus natos Dei, cum Deum diligamus et mandata eius faciamus.
1JOHN|5|3|Haec est enim caritas Dei, ut mandata eius servemus; et mandata eius gravia non sunt,
1JOHN|5|4|quoniam omne, quod natum est ex Deo, vincit mundum; et haec est victoria, quae vicit mundum: fides nostra.
1JOHN|5|5|Quis est qui vincit mundum, nisi qui credit quoniam Iesus est Filius Dei?
1JOHN|5|6|Hic est, qui venit per aquam et sanguinem, Iesus Christus; non in aqua solum sed in aqua et in sanguine. Et Spiritus est, qui testificatur, quoniam Spiritus est veritas.
1JOHN|5|7|Quia tres sunt, qui testificantur:
1JOHN|5|8|Spiritus et aqua et sanguis; et hi tres in unum sunt.
1JOHN|5|9|Si testimonium hominum accipimus, testimonium Dei maius est, quoniam hoc est testimonium Dei, quia testificatus est de Filio suo.
1JOHN|5|10|Qui credit in Filium Dei, habet testimonium in se. Qui non credit Deo, mendacem facit eum, quoniam non credidit in testimonium, quod testificatus est Deus de Filio suo.
1JOHN|5|11|Et hoc est testimonium, quoniam vitam aeternam dedit nobis Deus, et haec vita in Filio eius est.
1JOHN|5|12|Qui habet Filium, habet vitam; qui non habet Filium Dei, vitam non habet.
1JOHN|5|13|Haec scripsi vobis, ut sciatis quoniam vitam habetis aeternam, qui creditis in nomen Filii Dei.
1JOHN|5|14|Et haec est fiducia, quam habemus ad eum, quia si quid petierimus secundum voluntatem eius, audit nos.
1JOHN|5|15|Et si scimus quoniam audit nos, quidquid petierimus, scimus quoniam habemus petitiones, quas postulavimus ab eo.
1JOHN|5|16|Si quis videt fratrem suum peccare peccatum non ad mortem, petet, et dabit ei Deus vitam, peccantibus non ad mortem. Est peccatum ad mortem; non pro illo dico, ut roget.
1JOHN|5|17|Omnis iniustitia peccatum est, et est peccatum non ad mortem.
1JOHN|5|18|Scimus quoniam omnis, qui natus est ex Deo, non peccat, sed ille, qui genitus est ex Deo, conservat eum, et Malignus non tangit eum.
1JOHN|5|19|Scimus quoniam ex Deo sumus, et mundus totus in Maligno positus est.
1JOHN|5|20|Et scimus quoniam Filius Dei venit et dedit nobis sensum, ut cognoscamus eum, qui verus est; et sumus in eo, qui verus est, in Filio eius Iesu Christo. Hic est qui verus est, Deus et vita aeterna.
1JOHN|5|21|Filioli, custodite vos a simulacris!
