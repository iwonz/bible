ZEPH|1|1|Слово Господне, которое было к Софонии, сыну Хусия, сыну Годолии, сыну Амории, сыну Езекии, во дни Иосии, сына Амонова, царя Иудейского.
ZEPH|1|2|Все истреблю с лица земли, говорит Господь:
ZEPH|1|3|истреблю людей и скот, истреблю птиц небесных и рыб морских, и соблазны вместе с нечестивыми; истреблю людей с лица земли, говорит Господь.
ZEPH|1|4|И простру руку Мою на Иудею и на всех жителей Иерусалима: истреблю с места сего остатки Ваала, имя жрецов со священниками,
ZEPH|1|5|и тех, которые на кровлях поклоняются воинству небесному, и тех поклоняющихся, которые клянутся Господом и клянутся царем своим,
ZEPH|1|6|и тех, которые отступили от Господа, не искали Господа и не вопрошали о Нем.
ZEPH|1|7|Умолкни пред лицем Господа Бога! ибо близок день Господень: уже приготовил Господь жертвенное заклание, назначил, кого позвать.
ZEPH|1|8|И будет в день жертвы Господней: Я посещу князей и сыновей царя и всех, одевающихся в одежду иноплеменников;
ZEPH|1|9|посещу в тот день всех, которые перепрыгивают через порог, которые дом Господа своего наполняют насилием и обманом.
ZEPH|1|10|И будет в тот день, говорит Господь, вопль у ворот рыбных и рыдание у других ворот и великое разрушение на холмах.
ZEPH|1|11|Рыдайте, жители нижней части города, ибо исчезнет весь торговый народ и истреблены будут обремененные серебром.
ZEPH|1|12|И будет в то время: Я со светильником осмотрю Иерусалим и накажу тех, которые сидят на дрожжах своих и говорят в сердце своем: "не делает Господь ни добра, ни зла".
ZEPH|1|13|И обратятся богатства их в добычу и домы их – в запустение; они построят домы, а жить в них не будут, насадят виноградники, а вина из них не будут пить.
ZEPH|1|14|Близок великий день Господа, близок, и очень поспешает: уже слышен голос дня Господня; горько возопиет тогда и самый храбрый!
ZEPH|1|15|День гнева – день сей, день скорби и тесноты, день опустошения и разорения, день тьмы и мрака, день облака и мглы,
ZEPH|1|16|день трубы и бранного крика против укрепленных городов и высоких башен.
ZEPH|1|17|И Я стесню людей, и они будут ходить, как слепые, потому что они согрешили против Господа, и разметана будет кровь их, как прах, и плоть их – как помет.
ZEPH|1|18|Ни серебро их, ни золото их не может спасти их в день гнева Господа, и огнем ревности Его пожрана будет вся эта земля, ибо истребление, и притом внезапное, совершит Он над всеми жителями земли.
ZEPH|2|1|Исследуйте себя внимательно, исследуйте, народ необузданный,
ZEPH|2|2|доколе не пришло определение – день пролетит как мякина – доколе не пришел на вас пламенный гнев Господень, доколе не наступил для вас день ярости Господней.
ZEPH|2|3|Взыщите Господа, все смиренные земли, исполняющие законы Его; взыщите правду, взыщите смиренномудрие; может быть, вы укроетесь в день гнева Господня.
ZEPH|2|4|Ибо Газа будет покинута и Аскалон опустеет, Азот будет выгнан среди дня и Екрон искоренится.
ZEPH|2|5|Горе жителям приморской страны, народу Критскому! Слово Господне на вас, Хананеи, земля Филистимская! Я истреблю тебя, и не будет у тебя жителей, –
ZEPH|2|6|и будет приморская страна пастушьим овчарником и загоном для скота.
ZEPH|2|7|И достанется этот край остаткам дома Иудина, и будут пасти там, и в домах Аскалона будут вечером отдыхать, ибо Господь Бог их посетит их и возвратит плен их.
ZEPH|2|8|Слышал Я поношение Моава и ругательства сынов Аммоновых, как они издевались над Моим народом и величались на пределах его.
ZEPH|2|9|Посему, живу Я! говорит Господь Саваоф, Бог Израилев: Моав будет, как Содом, и сыны Аммона будут, как Гоморра, достоянием крапивы, соляною рытвиною, пустынею навеки; остаток народа Моего возьмет их в добычу, и уцелевшие из людей Моих получат их в наследие.
ZEPH|2|10|Это им за высокомерие их, за то, что они издевались и величались над народом Господа Саваофа.
ZEPH|2|11|Страшен будет для них Господь, ибо истребит всех богов земли, и Ему будут поклоняться, каждый со своего места, все острова народов.
ZEPH|2|12|И вы, Ефиопляне, избиты будете мечом Моим.
ZEPH|2|13|И прострет Он руку Свою на север, и уничтожит Ассура, и обратит Ниневию в развалины, в место сухое, как пустыня,
ZEPH|2|14|и покоиться будут среди нее стада и всякого рода животные; пеликан и еж будут ночевать в резных украшениях ее; голос их будет раздаваться в окнах, разрушение обнаружится на дверных столбах, ибо не станет на них кедровой обшивки.
ZEPH|2|15|Вот чем будет город торжествующий, живущий беспечно, говорящий в сердце своем: "я, и нет иного кроме меня". Как он стал развалиною, логовищем для зверей! Всякий, проходя мимо него, посвищет и махнет рукою.
ZEPH|3|1|Горе городу нечистому и оскверненному, притеснителю!
ZEPH|3|2|Не слушает голоса, не принимает наставления, на Господа не уповает, к Богу своему не приближается.
ZEPH|3|3|Князья его посреди него – рыкающие львы, судьи его – вечерние волки, не оставляющие до утра ни одной кости.
ZEPH|3|4|Пророки его – люди легкомысленные, вероломные; священники его оскверняют святыню, попирают закон.
ZEPH|3|5|Господь праведен посреди него, не делает неправды, каждое утро являет суд Свой неизменно; но беззаконник не знает стыда.
ZEPH|3|6|Я истребил народы, разрушены твердыни их; пустыми сделал улицы их, так что никто уже не ходит по ним; разорены города их: нет ни одного человека, нет жителей.
ZEPH|3|7|Я говорил: "бойся только Меня, принимай наставление!" и не будет истреблено жилище его, и не постигнет его зло, какое Я постановил о нем; а они прилежно старались портить все свои действия.
ZEPH|3|8|Итак ждите Меня, говорит Господь, до того дня, когда Я восстану для опустошения, ибо Мною определено собрать народы, созвать царства, чтобы излить на них негодование Мое, всю ярость гнева Моего; ибо огнем ревности Моей пожрана будет вся земля.
ZEPH|3|9|Тогда опять Я дам народам уста чистые, чтобы все призывали имя Господа и служили Ему единодушно.
ZEPH|3|10|Из заречных стран Ефиопии поклонники Мои, дети рассеянных Моих, принесут Мне дары.
ZEPH|3|11|В тот день ты не будешь срамить себя всякими поступками твоими, какими ты грешил против Меня, ибо тогда Я удалю из среды твоей тщеславящихся твоею знатностью, и не будешь более превозноситься на святой горе Моей.
ZEPH|3|12|Но оставлю среди тебя народ смиренный и простой, и они будут уповать на имя Господне.
ZEPH|3|13|Остатки Израиля не будут делать неправды, не станут говорить лжи, и не найдется в устах их языка коварного, ибо сами будут пастись и покоиться, и никто не потревожит их.
ZEPH|3|14|Ликуй, дщерь Сиона! торжествуй, Израиль! веселись и радуйся от всего сердца, дщерь Иерусалима!
ZEPH|3|15|Отменил Господь приговор над тобою, прогнал врага твоего! Господь, царь Израилев, посреди тебя: уже более не увидишь зла.
ZEPH|3|16|В тот день скажут Иерусалиму: "не бойся", и Сиону: "да не ослабевают руки твои!"
ZEPH|3|17|Господь Бог твой среди тебя, Он силен спасти тебя; возвеселится о тебе радостью, будет милостив по любви Своей, будет торжествовать о тебе с ликованием.
ZEPH|3|18|Сетующих о торжественных празднествах Я соберу: твои они, на них тяготеет поношение.
ZEPH|3|19|Вот, Я стесню всех притеснителей твоих в то время и спасу хромлющее, и соберу рассеянное, и приведу их в почет и именитость на всей этой земле поношения их.
ZEPH|3|20|В то время приведу вас и тогда же соберу вас, ибо сделаю вас именитыми и почетными между всеми народами земли, когда возвращу плен ваш перед глазами вашими, говорит Господь.
