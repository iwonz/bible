NAH|1|1|An oracle concerning Nineveh. The book of the vision of Nahum of Elkosh.
NAH|1|2|The LORD is a jealous and avenging God; the LORD is avenging and wrathful; the LORD takes vengeance on his adversaries and keeps wrath for his enemies.
NAH|1|3|The LORD is slow to anger and great in power, and the LORD will by no means clear the guilty. His way is in whirlwind and storm, and the clouds are the dust of his feet.
NAH|1|4|He rebukes the sea and makes it dry; he dries up all the rivers; Bashan and Carmel wither; the bloom of Lebanon withers.
NAH|1|5|The mountains quake before him; the hills melt; the earth heaves before him, the world and all who dwell in it.
NAH|1|6|Who can stand before his indignation? Who can endure the heat of his anger? His wrath is poured out like fire, and the rocks are broken into pieces by him.
NAH|1|7|The LORD is good, a stronghold in the day of trouble; he knows those who take refuge in him.
NAH|1|8|But with an overflowing flood he will make a complete end of the adversaries, and will pursue his enemies into darkness.
NAH|1|9|What do you plot against the LORD? He will make a complete end; trouble will not rise up a second time.
NAH|1|10|For they are like entangled thorns, like drunkards as they drink; they are consumed like stubble fully dried.
NAH|1|11|From you came one who plotted evil against the LORD, a worthless counselor.
NAH|1|12|Thus says the LORD, "Though they are at full strength and many, they will be cut down and pass away. Though I have afflicted you, I will afflict you no more.
NAH|1|13|And now I will break his yoke from off you and will burst your bonds apart."
NAH|1|14|The LORD has given commandment about you: "No more shall your name be perpetuated; from the house of your gods I will cut off the carved image and the metal image. I will make your grave, for you are vile."
NAH|1|15|Behold, upon the mountains, the feet of him who brings good news, who publishes peace! Keep your feasts, O Judah; fulfill your vows, for never again shall the worthless pass through you; he is utterly cut off.
NAH|2|1|The scatterer has come up against you. Man the ramparts; watch the road; dress for battle; collect all your strength.
NAH|2|2|For the LORD is restoring the majesty of Jacob as the majesty of Israel, for plunderers have plundered them and ruined their branches.
NAH|2|3|The shield of his mighty men is red; his soldiers are clothed in scarlet. The chariots come with flashing metal on the day he musters them; the cypress spears are brandished.
NAH|2|4|The chariots race madly through the streets; they rush to and fro through the squares; they gleam like torches; they dart like lightning.
NAH|2|5|He remembers his officers; they stumble as they go, they hasten to the wall; the siege tower is set up.
NAH|2|6|The river gates are opened; the palace melts away;
NAH|2|7|its mistress is stripped; she is carried off, her slave girls lamenting, moaning like doves and beating their breasts.
NAH|2|8|Nineveh is like a pool whose waters run away. "Halt! Halt!" they cry, but none turns back.
NAH|2|9|Plunder the silver, plunder the gold! There is no end of the treasure or of the wealth of all precious things.
NAH|2|10|Desolate! Desolation and ruin! Hearts melt and knees tremble; anguish is in all loins; all faces grow pale!
NAH|2|11|Where is the lions' den, the feeding place of the young lions, where the lion and lioness went, where his cubs were, with none to disturb?
NAH|2|12|The lion tore enough for his cubs and strangled prey for his lionesses; he filled his caves with prey and his dens with torn flesh.
NAH|2|13|Behold, I am against you, declares the LORD of hosts, and I will burn your chariots in smoke, and the sword shall devour your young lions. I will cut off your prey from the earth, and the voice of your messengers shall no longer be heard.
NAH|3|1|Woe to the bloody city, all full of lies and plunder- no end to the prey!
NAH|3|2|The crack of the whip, and rumble of the wheel, galloping horse and bounding chariot!
NAH|3|3|Horsemen charging, flashing sword and glittering spear, hosts of slain, heaps of corpses, dead bodies without end- they stumble over the bodies!
NAH|3|4|And all for the countless whorings of the prostitute, graceful and of deadly charms, who betrays nations with her whorings, and peoples with her charms.
NAH|3|5|Behold, I am against you, declares the LORD of hosts, and will lift up your skirts over your face; and I will make nations look at your nakedness and kingdoms at your shame.
NAH|3|6|I will throw filth at you and treat you with contempt and make you a spectacle.
NAH|3|7|And all who look at you will shrink from you and say, Wasted is Nineveh; who will grieve for her? Where shall I seek comforters for you?
NAH|3|8|Are you better than Thebes that sat by the Nile, with water around her, her rampart a sea, and water her wall?
NAH|3|9|Cush was her strength; Egypt too, and that without limit; Put and the Libyans were her helpers.
NAH|3|10|Yet she became an exile; she went into captivity; her infants were dashed in pieces at the head of every street; for her honored men lots were cast, and all her great men were bound in chains.
NAH|3|11|You also will be drunken; you will go into hiding; you will seek a refuge from the enemy.
NAH|3|12|All your fortresses are like fig trees with first-ripe figs- if shaken they fall into the mouth of the eater.
NAH|3|13|Behold, your troops are women in your midst. The gates of your land are wide open to your enemies; fire has devoured your bars.
NAH|3|14|Draw water for the siege; strengthen your forts; go into the clay; tread the mortar; take hold of the brick mold!
NAH|3|15|There will the fire devour you; the sword will cut you off. It will devour you like the locust. Multiply yourselves like the locust; multiply like the grasshopper!
NAH|3|16|You increased your merchants more than the stars of the heavens. The locust spreads its wings and flies away.
NAH|3|17|Your princes are like grasshoppers, your scribes like clouds of locusts settling on the fences in a day of cold- when the sun rises, they fly away; no one knows where they are.
NAH|3|18|Your shepherds are asleep, O king of Assyria; your nobles slumber. Your people are scattered on the mountains with none to gather them.
NAH|3|19|There is no easing your hurt; your wound is grievous. All who hear the news about you clap their hands over you. For upon whom has not come your unceasing evil?
