AMOS|1|1|Слова Амоса, що був між вівчарями з Текої, які він бачив на Ізраїля за днів Уззійї, Юдиного царя, та за днів Єровоама, Йоашового сина, Ізраїлевого царя, за два роки перед землетрусом.
AMOS|1|2|І він проказав: Загримить із Сіону Господь, і з Єрусалиму Свій голос подасть, і впадуть пасовища пастуші в жалобу та всохне вершина Кармелу!
AMOS|1|3|Так говорить Господь: За три переступи Дамаску й за чотири цього не прощу: за те, що вони молотили Ґілеада ціпами залізними.
AMOS|1|4|І пошлю Я огонь на дім Хазаїла, і пожере він палати Бен-Гадада.
AMOS|1|5|І зламаю засува Дамаску, і мешканця витну з долини Авен, і того, хто держатиме берло з Бет-Едене, і арамський народ піде в Кір на вигнання, говорить Господь.
AMOS|1|6|Так говорить Господь: За три переступи Аззи й за чотири цього не прощу: що всіх гнали в полон, щоб віддати Едомові.
AMOS|1|7|І пошлю Я огонь на мур Ґази, і поїсть він палати її.
AMOS|1|8|І мешканця витну з Ашдоду, і берлодержця з Ашкелону, і зверну Свою руку на Екрон, і вигинуть рештки филистимлян, говорить Господь.
AMOS|1|9|Так говорить Господь: За три переступи Тиру й за чотири цього не прощу: за те, що він видав усіх на вигнання в Едом, і не пам'ятав заповіту братів.
AMOS|1|10|І пошлю Я огонь на мур Тиру, і пожере він палати його!
AMOS|1|11|Так говорить Господь: За три переступи Едому й за чотири цього не прощу: за те, що мечем він гнав брата свого, і знищив своє милосердя, свій гнів завжди стеріг, а лютість свою пильнував повсякчасно.
AMOS|1|12|І пошлю Я огонь до Теману і пожере він палати Боцри!
AMOS|1|13|Так говорить Господь: За три переступи Аммонових синів й за чотири цього не прощу: за те, що пороли ґілеадських вагітних, щоб поширити границі свої!
AMOS|1|14|І огонь запалю Я на мурі Рабби, і пожере він палати її, із криком в день бою, із вихром в день бурі.
AMOS|1|15|І піде їхній цар на вигнання, він і князі його разом, говорить Господь.
AMOS|2|1|Так говорить Господь: За три переступи Моава й за чотири цього не прощу: за те, що спалив на вапно кості едомського царя!
AMOS|2|2|І пошлю Я огонь на Моава, і пожере він палати Керіййоту, і загине Моав серед галасу, серед крику, при голосі рога.
AMOS|2|3|І витну суддю з-серед нього, а з ним позабиваю князів його всіх, говорить Господь.
AMOS|2|4|Так говорить Господь: За три прогріхи Юди й за чотири цього не прощу: за те, що повідкидали Господній Закон, і постанов Його не стерегли, і що на манівці їх звели їхні лжебоги, за якими пішли їхні батьки.
AMOS|2|5|І пошлю Я на Юду огонь, і пожере він палати Єрусалиму!
AMOS|2|6|Так говорить Господь: За три переступи Ізраїлеві й за чотири цього не прощу: за те, що за срібло вони продають справедливого, а за чоботи вбогого!
AMOS|2|7|Вони топчуть у земному поросі голову бідних, а дорогу сумирних викривлюють. А син й його батько вчащають до однієї блудниці, щоб святе Моє Ймення зневажити.
AMOS|2|8|І вони стелять одіж заставлену, щоб півлежати при кожному жертівнику, і п'ють в домі Бога свого вино від покараних.
AMOS|2|9|І Я вигубив був з-перед них Аморея, що його височінь, як високий той кедр, і він міцний, як дуб. Та Я плід його знищив згори, а здолу коріння його.
AMOS|2|10|А вас Я був вивів із краю єгипетського, і сорок років провадив пустинею вас, щоб ви Край аморейський успадкували.
AMOS|2|11|І пророків Я збуджував з ваших синів, а з ваших юнців назореїв. Хіба ж то не так, синове Ізраїлеві? говорить Господь.
AMOS|2|12|А ви назореїв поїли вином, а пророкам наказували й говорили: Не пророкуйте!
AMOS|2|13|Отож Я потисну на вас, як тисне снопами наповнений віз,
AMOS|2|14|і згине й в моторного втеча, і потужний не втримає сили своєї, а лицар свого життя не врятує.
AMOS|2|15|І не встоїть із лука стрілець, і своїми ногами прудкий не втече, і верхівець не врятує свого життя.
AMOS|2|16|І наймужніший з лицарства нагим утече того дня, говорить Господь.
AMOS|3|1|Послухайте слова того, що Господь говорив проти вас, синове Ізраїлеві, на ввесь оцей рід, що його Я підніс був із краю єгипетського, промовляючи:
AMOS|3|2|Тільки вас Я пізнав зо всіх родів землі, тому вас навіщу за всі ваші провини!
AMOS|3|3|Чи йдуть двоє разом, якщо не умовились?
AMOS|3|4|Чи реве в лісі лев, як нема йому здобичі? Чи левчук видає голос свій із своєї нори, якщо він не зловив?
AMOS|3|5|Чи впаде на землі пташка в сітку, як немає сільця? Чи підійметься сітка з землі, як нічого не зловить?
AMOS|3|6|Чи в місті засурмлять у сурму, а народ не тремтітиме? Чи станеться в місті нещастя, що його не Господь допустив?
AMOS|3|7|Бо не чинить нічого Господь Бог, не виявивши таємниці Своєї Своїм рабам пророкам.
AMOS|3|8|Лев зареве, хто того не злякається? Господь Бог заговорить, хто пророкувати не буде?
AMOS|3|9|Розголосіть над палацами в Ашдоді, і над палатами в краї єгипетському, та й скажіть: Позбирайтеся на горах Самарії, і побачте велике збентеження в ній, та утиск у ній!
AMOS|3|10|І правдиво не вміють робити вони, говорить Господь, насильство громадять та грабунок в палатах своїх.
AMOS|3|11|Тому так Господь Бог промовляє: Ворог обляже навколо цієї землі, і скине із тебе він силу твою, і пограбовані будуть палати твої.
AMOS|3|12|Так говорить Господь: Як часом рятує пастух з пащі лев'ячої дві коліні, або пипку вуха, так будуть врятовані діти Ізраїлеві, що сидять в Самарії в закуточку ліжка, та на адамашку постелі.
AMOS|3|13|Послухайте ви та й засвідчіть ув Якововім домі, говорить Господь Бог, Бог Саваот.
AMOS|3|14|Бо в той день, коли Я покараю Ізраїля за провини його, то Я покараю за жертівники Бет-Елу, і будуть відрубані роги жертівника, і на землю попадають.
AMOS|3|15|І Я розіб'ю дім зимовий разом з домом літнім, і загинуть доми із слонової кости, і не стане багато домів, говорить Господь.
AMOS|4|1|Послухайте слова оцього, корови башанські, які на горі самарійській, що тиснете бідних, торощите вбогих, що своїм хазяям ви говорите: Принеси, і ми будемо пити!
AMOS|4|2|Присягав Господь Бог Своєю святістю, що ось дні настають на вас, і будуть тягти вас гаками, а ваших нащадків гачками для ловлення риби!
AMOS|4|3|І ви повиходите виломами, кожна окремо собі, і кинетеся до Хермону, говорить Господь.
AMOS|4|4|Прийдіть до Бет-Елу й грішіть, до Ґілґалу примножте грішити. І свої жертви приносьте щоранку, на три дні ваші десятини.
AMOS|4|5|І з димом пустіть жертву вдячну квасну, і сповістіть добровільні дарунки, розголосіть, бо ви любите так, синове Ізраїлеві, говорить Господь Бог.
AMOS|4|6|І тому Я вам дав чистоту зубів по всіх ваших містах, і брак хліба по всіх ваших місцях, та ви не вернулись до Мене, говорить Господь...
AMOS|4|7|І Я стримав вам дощ за три місяці перед жнивами, і дощ посилав на одне місто, а на друге місто не посилав; одна ділянка була побита дощем, а ділянка, на яку не пустив Я дощу, висихала.
AMOS|4|8|І два-три міста рушали до міста одного напитись води, але не насичувались, та ви не вернулись до Мене, говорить Господь...
AMOS|4|9|Я бив вас посухою та зеленячкою, сарана жерла безліч ваших садків й виноградників ваших, і ваших фіґовниць та ваших олив, та ви не вернулись до Мене, говорить Господь...
AMOS|4|10|Я на вас посилав моровицю, немов на Єгипет, мечем побивав ваших хлопців, полонячи разом і коней у вас, підіймав до ніздер сморід ваших таборів, та ви не вернулись до Мене, говорить Господь...
AMOS|4|11|Я винищив вас, як Содом та Гоморру Бог винищив, і ви стали, немов головешка, з пожару врятована, та ви не вернулись до Мене, говорить Господь...
AMOS|4|12|Тому то зроблю тобі так, о Ізраїлю, а що Я зроблю тобі це, приготуйся, Ізраїлю, до зустрічі Бога свого!
AMOS|4|13|Бо це Той, що вформовує гори, і що створює вітра, що людині показує задум її, що робить зірницю темнотою, і ступає по згір'ях землі, Господь Бог Саваот Йому Ймення!
AMOS|5|1|Послухайте слова цього, що я ним голосіння підношу за вас, о доме Ізраїлів!
AMOS|5|2|Упала, і більше не встане та діва Ізраїлева! Вона кинена на свою землю, немає, хто звів би її!
AMOS|5|3|Бо так Господь Бог промовляє: Місто, що виходило тисячею, позоставить лиш сотню, а те, що виходило сотнею, позоставить десятку для дому Ізраїля.
AMOS|5|4|Бо так промовляє Господь до дому Ізраїлевого: Наверніться до Мене й живіть!
AMOS|5|5|І не звертайтеся до Бет-Елу, і до Ґілґалу не приходьте, а через Беер-Шеву не переходьте, бо на вигнання Ґілґал конче піде, і марнотою стане Бет-Ел.
AMOS|5|6|Наверніться до Господа, і будете жити, щоб Він не ввійшов, як огонь до Йосипового дому, і буде він жерти, та не буде кому погасити в Бет-Елі,
AMOS|5|7|вони змінюють суд на полин, і кидають правду на землю.
AMOS|5|8|Той, хто Волосожара й Оріона створив, Хто смертну темноту зміняє на ранок, а день затемняє на ніч, хто прикликує воду морську й виливає її на поверхню землі, Господь Ймення Йому!
AMOS|5|9|Він наводить погибіль на сильного, і прийде погибіль твердині!
AMOS|5|10|Вони ненавидять того, хто у брамі картає, і обриджують тим, хто говорить правдиве.
AMOS|5|11|Тому, що нужденного топчете ви, і дарунки збіжеві берете від нього, що ви набудували будинків із каменя тесаного, то сидіти не будете в них; понасаджували винограду улюбленого, та не будете пити із нього вина!
AMOS|5|12|Бо Я знаю про ваші численні провини і про ваші великі гріхи: тиснете ви справедливого, берете ви підкупа та викривляєте право убогих у брамі.
AMOS|5|13|Тому то розумний мовчить цього часу, бо це час лихий.
AMOS|5|14|Шукайте добра, а не зла, щоб вам жити, і буде із вами Господь, Бог Саваот, так, як кажете ви.
AMOS|5|15|Ненавидьте зло й покохайте добро, і правосуддя поставте у брамі, може змилується Господь, Бог Саваот над решткою Йосипа.
AMOS|5|16|Тому так промовляє Господь, Бог Саваот, Вседержитель: На майданах усіх голосіння, на всіх вулицях крики: ой, ой! І покличуть хліборобів на жалобу, і голосільниць, що вміють плачливі пісні,
AMOS|5|17|і стане ридання по всіх виноградниках, бо Я перейду серед тебе, говорить Господь!
AMOS|5|18|Горе тим, що жадають Господнього дня, нащо це вам день Господній? Він не світло, а темрява!
AMOS|5|19|Це так, коли хто утікає від лева, і ведмідь спотикає його! І він убігає до дому, і оперся своєю рукою об стіну, аж гадюка кусає його...
AMOS|5|20|Чи ж не є день Господній темнота, а не світло, і хіба він не темний, і сяйва немає у ньому?
AMOS|5|21|Зненавидів Я, обридив Собі ваші свята, і не нюхаю жертов ваших зборів...
AMOS|5|22|І коли принесете Мені цілопалення та хлібні жертви свої, Я Собі не вподобаю їх, а на мирні жертви ваші із ситих баранів не погляну...
AMOS|5|23|Усунь же від Мене пісень своїх гук, і не почую Я рокоту гусел твоїх,
AMOS|5|24|і хай тече правосуддя, немов та вода, а справедливість як сильний потік!
AMOS|5|25|Чи ж жертви та хлібні приноси за тих сорок літ на пустині Мені ви приносили, доме Ізраїлів?
AMOS|5|26|Ви ж носили Саккута, свойого царя, та Кевана, свої виображення, зорю ваших богів, що собі поробили.
AMOS|5|27|Тому Я вас вижену геть за Дамаск, говорить Господь, що Бог Саваот Йому Ймення!
AMOS|6|1|Горе безпечним на Сіоні, тим, хто надіється на самарійськую гору, тим шляхетним першого з народів, до яких прибуває Ізраїлів дім!
AMOS|6|2|Перейдіть до Калне та й побачте, і звідти підіть до Гамату великого, і зійдіть до Ґату филистимлян! Чи ліпші вони від цих царств? Чи їхня границя більша за вашу границю?
AMOS|6|3|День нещастя вважаєте ви за далекий, а час насильства зближаєте!
AMOS|6|4|Ви вилежуєтеся на ложах з слонової кости і вивалюєтесь на постелях своїх, і їсте баранів із отари та ситих телят із обори.
AMOS|6|5|Під гусла співаєте ви, мов Давид, ви музичні знаряддя собі видумляєте.
AMOS|6|6|Ви вино попиваєте чашами, і намащуєтесь добірною оливою, і над спустошенням Йосипа не вболіваєте.
AMOS|6|7|Тому вони підуть тепер на вигнання на чолі полонених, і перестане крик випещених.
AMOS|6|8|Господь присягнув був Своєю душею, говорить Господь, Бог Саваот: Пишнотою Якова бриджу, і палати його Я ненавиджу, і видам те місто та все, що є в ньому.
AMOS|6|9|І буде, якщо десять люда зостануться в домі одному, то й вони повмирають.
AMOS|6|10|І його візьме родич та й спалить його, щоб винести кості із дому, і скаже до того, хто буде в середині дому: Чи ще є хто з тобою? А той відповість: Вже немає нікого! і скаже той: Тихше, бо не згадується Ймення Господа!
AMOS|6|11|Бо Господь ось накаже, і ворог розіб'є великий той дім на відламки, а дім малий на тріски.
AMOS|6|12|Чи бігають коні по скелі? Чи хто виоре море худобою? Таж ви суд обернули на гіркість, а плід справедливости на полин!
AMOS|6|13|Ви марнотою тішитеся та говорите: Хіба ж ми не власною силою набули собі роги?
AMOS|6|14|Бо ось Я поставлю народ проти вас, доме Ізраїлів, каже Господь, Бог Саваот, і вони вас потиснуть ізвідти, де йдуть до Гамату, аж до степового потоку!
AMOS|7|1|Господь Бог учинив, що я бачив таке: Ось Він утворив сарану, коли почала виростати отава, і ось отава як по сінокосі царському!
AMOS|7|2|І сталось, як вона вже пожерла траву на землі, я сказав: Господи, Боже, прости! Як же Яків устояти може, бо такий він малий?
AMOS|7|3|І Господь пожалів був про те. Не станеться це, промовив Господь.
AMOS|7|4|Господь Бог учинив, що я бачив таке: Ось Господь Бог покликав судитись огнем, і пожер той велику безодню, і частку пожер.
AMOS|7|5|І сказав я: О, Господи, Боже, спини! Як же Яків устояти може, бо такий він малий?
AMOS|7|6|І Господь пожалів був про те. Не станеться й це! сказав Господь Бог!
AMOS|7|7|І Він знов учинив, що я бачив таке: Ось на мурі стрімкому стоїть Господь Бог, а в руці Його висок.
AMOS|7|8|І промовив до мене Господь: Що ти бачиш, Амосе? А я відказав: Виска. І промовив Господь: Ось Я цього виска покладу посеред народу Мого, Ізраїля, уже більше йому не прощу!
AMOS|7|9|І спустошіють жертовні підгірки Ісакові, і поруйновані будуть святині Ізраїлеві, і Я стану з мечем на дім Єровоамів.
AMOS|7|10|І послав Амація, священик Бет-Елу, до Єровоама, царя Ізраїлевого, кажучи: Амос змовлюється на тебе серед Ізраїлевого дому, не може земля змістити всіх його слів!
AMOS|7|11|Бо так говорить Амос: Єровоам помре від меча, а Ізраїль конче піде на вигнання з своєї землі!
AMOS|7|12|І сказав Амація до Амоса: Ясновидче, іди, утікай собі до Юдиного краю, і їж там хліб, і там пророкуй.
AMOS|7|13|А в Бет-Елі вже більше не будеш пророкувати, бо він святиня царя та дім царства.
AMOS|7|14|І відповів Амос і сказав до Амації: Я не пророк, і не син я пророків, я пастух та оброблювач диких фіґовниць.
AMOS|7|15|І взяв мене Господь від отари, і промовив до мене Господь: Іди, пророкуй Моєму народові Ізраїлеві!
AMOS|7|16|А тепер послухай Господнього слова: Ти кажеш: Не будеш пророкувати на Ізраїля, і не будеш проповідувати на Ісаків дім.
AMOS|7|17|Тому так промовляє Господь: Твоя жінка в місті буде блудлива, і сини твої та дочки твої попадають від меча, а земля твоя буде поділена шнуром, і ти помреш на нечистій землі, а Ізраїль конче піде на вигнання з своєї землі!
AMOS|8|1|Господь Бог учинив, що я бачив таке: Ось кіш доспілих плодів.
AMOS|8|2|І сказав Він: Що бачиш, Амосе? А я відказав: Кіш доспілих плодів. І промовив до мене Господь: Доспів кінець Моєму народові Ізраїлеві, уже більше йому не прощу!
AMOS|8|3|І обернуться пісні в палатах на зойк того дня, говорить Господь Бог: буде трупів багато, бо ворог на кожному місці накидає їх!
AMOS|8|4|Послухайте це, ви, що топчете бідного, і що прагнете винищити всіх убогих з землі,
AMOS|8|5|кажучи: Коли то мине новомісяччя, щоб нам збіжжя продати? і субота, щоб нам відчинити збіжеві комори? Щоб зменшити ефу, і щоб шекля побільшити, і щоб викривляти обманну вагу,
AMOS|8|6|щоб купувати за срібло нужденних, а вбогого за взуття, і попродати послід збіжевий?
AMOS|8|7|Господь присягнув славою Якова: Не забуду ніколи усіх їхніх вчинків!
AMOS|8|8|Чи не затрясеться від цього земля, і всі мешканці її не впадуть у жалобу? Вся вона захвилюється, мов та Ріка, і бурхливо поплине й обнизиться знов, немов річка Єгипту.
AMOS|8|9|І станеться в день той, говорить Господь Бог, і вчиню захід сонця опівдні, і для землі серед світлого дня воно стемніє.
AMOS|8|10|І оберну ваші свята в жалобу, а всі ваші пісні в голосіння, і на всі стегна спроваджу верету, а на всякую голову лисину, і вчиню це, немов та жалоба по одинакові, кінець же отого, немов гіркий день!
AMOS|8|11|Ось дні настають, говорить Господь Бог, і голод пошлю Я на землю, не голод на хліб, і не спрагу на воду, але спрагу почути Господні слова!
AMOS|8|12|І будуть ходити від моря до моря, і з півночі до сходу блукатимуть, щоб знайти слово Господа, та не знайдуть його!
AMOS|8|13|Того дня будуть мліти від спраги вродливі дівчата та хлопці,
AMOS|8|14|що клянуться гріхом самарійським та кажуть: Як живий твій Бог, Дане, і як жива дорога до Беер-Шеви! Та вони всі попадають, і більше не встануть...
AMOS|9|1|Я бачив Господа, що стояв над жертівником, і Він сказав: Удар но по маковиці цих воріт, щоб затряслися пороги, і порозбивай їх на всіх їхніх головах, а їхній останок заб'ю Я мечем. Не втече їм втікач, і гонець не врятується в них!
AMOS|9|2|Якщо б закопались вони до шеолу, то й звідти рука Моя їх забере, і якщо б піднялися на небо, то й звідти їх скину!
AMOS|9|3|А якщо б поховались вони на верховині Кармелу, звідти вишукаю й заберу їх, а якщо на дні моря вони поховаються з-перед очей Моїх, то й там Я гадюці звелю, і вона їх покусає!
AMOS|9|4|А якщо вони підуть в полон перед своїми ворогами, то й там накажу Я мечеві і він їх повбиває, і на них Я зверну Своє око на зле, а не на добре.
AMOS|9|5|Бо коли Господь Бог Саваот доторкнеться землі, то розтане вона, і в жалобу впадуть всі мешканці її. І вся вона вийде, немов та Ріка, і мов річка Єгипту обнизиться.
AMOS|9|6|Він будує на небі чертоги Свої, а Свій небозвід заклав над землею, воду морську Він кличе, і виливає її на поверхню землі, Господь Йому Ймення!
AMOS|9|7|Хіба ж ви, Ізраїлеві сини, Мені не такі, як сини етіоплян? говорить Господь. Хіба ж не Ізраїля вивів Я з краю єгипетського, а филистимлян з Кафтору, а Арама із Кіру?
AMOS|9|8|Ось очі Господа Бога на грішне це царство, і з поверхні землі його вигублю, та вигублюючи, не погублю дому Якового, говорить Господь.
AMOS|9|9|Бо ось Я звелів, і серед народів усіх пересію Ізраїлів дім, як пересівається решетом, і жодне зеренце на землю не випаде!
AMOS|9|10|Упадуть усі грішні народу Мого від меча, що говорять: Не досягне до нас і не стріне оце нас нещастя!
AMOS|9|11|Того дня Я поставлю упалу Давидову скинію і проломи в ній загороджу, і поставлю руїни його, і відбудую його, як за днів стародавніх,
AMOS|9|12|щоб решту Едому посіли вони, і всі ті народи, що в них кликалося Моє Ймення, говорить Господь, Який чинить оце.
AMOS|9|13|Ось дні настають, говорить Господь, і орач із женцем зустрінеться, а топтач винограду із сіячем, і гори закрапають виноградовим соком, а всі взгір'я добром потечуть.
AMOS|9|14|І долю народу Свого, Ізраїля, Я поверну, і побудую міста попустошені, і осядуть вони, і засадять вони виноградники, й питимуть їхнє вино, і порозводять садки, і будуть їсти їхній овоч.
AMOS|9|15|І Я посаджу їх на їхній землі, і не будуть їх більш виривати з своєї землі, яку Я їм дав, говорить Господь, Бог твій!
