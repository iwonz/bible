ACTS|1|1|In my former book, Theophilus, I wrote about all that Jesus began to do and to teach
ACTS|1|2|until the day he was taken up to heaven, after giving instructions through the Holy Spirit to the apostles he had chosen.
ACTS|1|3|After his suffering, he showed himself to these men and gave many convincing proofs that he was alive. He appeared to them over a period of forty days and spoke about the kingdom of God.
ACTS|1|4|On one occasion, while he was eating with them, he gave them this command: "Do not leave Jerusalem, but wait for the gift my Father promised, which you have heard me speak about.
ACTS|1|5|For John baptized with water, but in a few days you will be baptized with the Holy Spirit."
ACTS|1|6|So when they met together, they asked him, "Lord, are you at this time going to restore the kingdom to Israel?"
ACTS|1|7|He said to them: "It is not for you to know the times or dates the Father has set by his own authority.
ACTS|1|8|But you will receive power when the Holy Spirit comes on you; and you will be my witnesses in Jerusalem, and in all Judea and Samaria, and to the ends of the earth."
ACTS|1|9|After he said this, he was taken up before their very eyes, and a cloud hid him from their sight.
ACTS|1|10|They were looking intently up into the sky as he was going, when suddenly two men dressed in white stood beside them.
ACTS|1|11|"Men of Galilee," they said, "why do you stand here looking into the sky? This same Jesus, who has been taken from you into heaven, will come back in the same way you have seen him go into heaven."
ACTS|1|12|Then they returned to Jerusalem from the hill called the Mount of Olives, a Sabbath day's walk from the city.
ACTS|1|13|When they arrived, they went upstairs to the room where they were staying. Those present were Peter, John, James and Andrew; Philip and Thomas, Bartholomew and Matthew; James son of Alphaeus and Simon the Zealot, and Judas son of James.
ACTS|1|14|They all joined together constantly in prayer, along with the women and Mary the mother of Jesus, and with his brothers.
ACTS|1|15|In those days Peter stood up among the believers (a group numbering about a hundred and twenty)
ACTS|1|16|and said, "Brothers, the Scripture had to be fulfilled which the Holy Spirit spoke long ago through the mouth of David concerning Judas, who served as guide for those who arrested Jesus--
ACTS|1|17|he was one of our number and shared in this ministry."
ACTS|1|18|(With the reward he got for his wickedness, Judas bought a field; there he fell headlong, his body burst open and all his intestines spilled out.
ACTS|1|19|Everyone in Jerusalem heard about this, so they called that field in their language Akeldama, that is, Field of Blood.)
ACTS|1|20|"For," said Peter, "it is written in the book of Psalms, "'May his place be deserted; let there be no one to dwell in it,' and, "'May another take his place of leadership.'
ACTS|1|21|Therefore it is necessary to choose one of the men who have been with us the whole time the Lord Jesus went in and out among us,
ACTS|1|22|beginning from John's baptism to the time when Jesus was taken up from us. For one of these must become a witness with us of his resurrection."
ACTS|1|23|So they proposed two men: Joseph called Barsabbas (also known as Justus) and Matthias.
ACTS|1|24|Then they prayed, "Lord, you know everyone's heart. Show us which of these two you have chosen
ACTS|1|25|to take over this apostolic ministry, which Judas left to go where he belongs."
ACTS|1|26|Then they cast lots, and the lot fell to Matthias; so he was added to the eleven apostles.
ACTS|2|1|When the day of Pentecost came, they were all together in one place.
ACTS|2|2|Suddenly a sound like the blowing of a violent wind came from heaven and filled the whole house where they were sitting.
ACTS|2|3|They saw what seemed to be tongues of fire that separated and came to rest on each of them.
ACTS|2|4|All of them were filled with the Holy Spirit and began to speak in other tongues as the Spirit enabled them.
ACTS|2|5|Now there were staying in Jerusalem God-fearing Jews from every nation under heaven.
ACTS|2|6|When they heard this sound, a crowd came together in bewilderment, because each one heard them speaking in his own language.
ACTS|2|7|Utterly amazed, they asked: "Are not all these men who are speaking Galileans?
ACTS|2|8|Then how is it that each of us hears them in his own native language?
ACTS|2|9|Parthians, Medes and Elamites; residents of Mesopotamia, Judea and Cappadocia, Pontus and Asia,
ACTS|2|10|Phrygia and Pamphylia, Egypt and the parts of Libya near Cyrene; visitors from Rome
ACTS|2|11|(both Jews and converts to Judaism); Cretans and Arabs--we hear them declaring the wonders of God in our own tongues!"
ACTS|2|12|Amazed and perplexed, they asked one another, "What does this mean?"
ACTS|2|13|Some, however, made fun of them and said, "They have had too much wine. "
ACTS|2|14|Then Peter stood up with the Eleven, raised his voice and addressed the crowd: "Fellow Jews and all of you who live in Jerusalem, let me explain this to you; listen carefully to what I say.
ACTS|2|15|These men are not drunk, as you suppose. It's only nine in the morning!
ACTS|2|16|No, this is what was spoken by the prophet Joel:
ACTS|2|17|"'In the last days, God says, I will pour out my Spirit on all people. Your sons and daughters will prophesy, your young men will see visions, your old men will dream dreams.
ACTS|2|18|Even on my servants, both men and women, I will pour out my Spirit in those days, and they will prophesy.
ACTS|2|19|I will show wonders in the heaven above and signs on the earth below, blood and fire and billows of smoke.
ACTS|2|20|The sun will be turned to darkness and the moon to blood before the coming of the great and glorious day of the Lord.
ACTS|2|21|And everyone who calls on the name of the Lord will be saved.'
ACTS|2|22|"Men of Israel, listen to this: Jesus of Nazareth was a man accredited by God to you by miracles, wonders and signs, which God did among you through him, as you yourselves know.
ACTS|2|23|This man was handed over to you by God's set purpose and foreknowledge; and you, with the help of wicked men, put him to death by nailing him to the cross.
ACTS|2|24|But God raised him from the dead, freeing him from the agony of death, because it was impossible for death to keep its hold on him.
ACTS|2|25|David said about him: "'I saw the Lord always before me. Because he is at my right hand, I will not be shaken.
ACTS|2|26|Therefore my heart is glad and my tongue rejoices; my body also will live in hope,
ACTS|2|27|because you will not abandon me to the grave, nor will you let your Holy One see decay.
ACTS|2|28|You have made known to me the paths of life; you will fill me with joy in your presence.'
ACTS|2|29|"Brothers, I can tell you confidently that the patriarch David died and was buried, and his tomb is here to this day.
ACTS|2|30|But he was a prophet and knew that God had promised him on oath that he would place one of his descendants on his throne.
ACTS|2|31|Seeing what was ahead, he spoke of the resurrection of the Christ, that he was not abandoned to the grave, nor did his body see decay.
ACTS|2|32|God has raised this Jesus to life, and we are all witnesses of the fact.
ACTS|2|33|Exalted to the right hand of God, he has received from the Father the promised Holy Spirit and has poured out what you now see and hear.
ACTS|2|34|For David did not ascend to heaven, and yet he said, "'The Lord said to my Lord: "Sit at my right hand
ACTS|2|35|until I make your enemies a footstool for your feet."'
ACTS|2|36|"Therefore let all Israel be assured of this: God has made this Jesus, whom you crucified, both Lord and Christ."
ACTS|2|37|When the people heard this, they were cut to the heart and said to Peter and the other apostles, "Brothers, what shall we do?"
ACTS|2|38|Peter replied, "Repent and be baptized, every one of you, in the name of Jesus Christ for the forgiveness of your sins. And you will receive the gift of the Holy Spirit.
ACTS|2|39|The promise is for you and your children and for all who are far off--for all whom the Lord our God will call."
ACTS|2|40|With many other words he warned them; and he pleaded with them, "Save yourselves from this corrupt generation."
ACTS|2|41|Those who accepted his message were baptized, and about three thousand were added to their number that day.
ACTS|2|42|They devoted themselves to the apostles' teaching and to the fellowship, to the breaking of bread and to prayer.
ACTS|2|43|Everyone was filled with awe, and many wonders and miraculous signs were done by the apostles.
ACTS|2|44|All the believers were together and had everything in common.
ACTS|2|45|Selling their possessions and goods, they gave to anyone as he had need.
ACTS|2|46|Every day they continued to meet together in the temple courts. They broke bread in their homes and ate together with glad and sincere hearts,
ACTS|2|47|praising God and enjoying the favor of all the people. And the Lord added to their number daily those who were being saved.
ACTS|3|1|One day Peter and John were going up to the temple at the time of prayer--at three in the afternoon.
ACTS|3|2|Now a man crippled from birth was being carried to the temple gate called Beautiful, where he was put every day to beg from those going into the temple courts.
ACTS|3|3|When he saw Peter and John about to enter, he asked them for money.
ACTS|3|4|Peter looked straight at him, as did John. Then Peter said, "Look at us!"
ACTS|3|5|So the man gave them his attention, expecting to get something from them.
ACTS|3|6|Then Peter said, "Silver or gold I do not have, but what I have I give you. In the name of Jesus Christ of Nazareth, walk."
ACTS|3|7|Taking him by the right hand, he helped him up, and instantly the man's feet and ankles became strong.
ACTS|3|8|He jumped to his feet and began to walk. Then he went with them into the temple courts, walking and jumping, and praising God.
ACTS|3|9|When all the people saw him walking and praising God,
ACTS|3|10|they recognized him as the same man who used to sit begging at the temple gate called Beautiful, and they were filled with wonder and amazement at what had happened to him.
ACTS|3|11|While the beggar held on to Peter and John, all the people were astonished and came running to them in the place called Solomon's Colonnade.
ACTS|3|12|When Peter saw this, he said to them: "Men of Israel, why does this surprise you? Why do you stare at us as if by our own power or godliness we had made this man walk?
ACTS|3|13|The God of Abraham, Isaac and Jacob, the God of our fathers, has glorified his servant Jesus. You handed him over to be killed, and you disowned him before Pilate, though he had decided to let him go.
ACTS|3|14|You disowned the Holy and Righteous One and asked that a murderer be released to you.
ACTS|3|15|You killed the author of life, but God raised him from the dead. We are witnesses of this.
ACTS|3|16|By faith in the name of Jesus, this man whom you see and know was made strong. It is Jesus' name and the faith that comes through him that has given this complete healing to him, as you can all see.
ACTS|3|17|"Now, brothers, I know that you acted in ignorance, as did your leaders.
ACTS|3|18|But this is how God fulfilled what he had foretold through all the prophets, saying that his Christ would suffer.
ACTS|3|19|Repent, then, and turn to God, so that your sins may be wiped out, that times of refreshing may come from the Lord,
ACTS|3|20|and that he may send the Christ, who has been appointed for you--even Jesus.
ACTS|3|21|He must remain in heaven until the time comes for God to restore everything, as he promised long ago through his holy prophets.
ACTS|3|22|For Moses said, 'The Lord your God will raise up for you a prophet like me from among your own people; you must listen to everything he tells you.
ACTS|3|23|Anyone who does not listen to him will be completely cut off from among his people.'
ACTS|3|24|"Indeed, all the prophets from Samuel on, as many as have spoken, have foretold these days.
ACTS|3|25|And you are heirs of the prophets and of the covenant God made with your fathers. He said to Abraham, 'Through your offspring all peoples on earth will be blessed.'
ACTS|3|26|When God raised up his servant, he sent him first to you to bless you by turning each of you from your wicked ways."
ACTS|4|1|The priests and the captain of the temple guard and the Sadducees came up to Peter and John while they were speaking to the people.
ACTS|4|2|They were greatly disturbed because the apostles were teaching the people and proclaiming in Jesus the resurrection of the dead.
ACTS|4|3|They seized Peter and John, and because it was evening, they put them in jail until the next day.
ACTS|4|4|But many who heard the message believed, and the number of men grew to about five thousand.
ACTS|4|5|The next day the rulers, elders and teachers of the law met in Jerusalem.
ACTS|4|6|Annas the high priest was there, and so were Caiaphas, John, Alexander and the other men of the high priest's family.
ACTS|4|7|They had Peter and John brought before them and began to question them: "By what power or what name did you do this?"
ACTS|4|8|Then Peter, filled with the Holy Spirit, said to them: "Rulers and elders of the people!
ACTS|4|9|If we are being called to account today for an act of kindness shown to a cripple and are asked how he was healed,
ACTS|4|10|then know this, you and all the people of Israel: It is by the name of Jesus Christ of Nazareth, whom you crucified but whom God raised from the dead, that this man stands before you healed.
ACTS|4|11|He is "'the stone you builders rejected, which has become the capstone. '
ACTS|4|12|Salvation is found in no one else, for there is no other name under heaven given to men by which we must be saved."
ACTS|4|13|When they saw the courage of Peter and John and realized that they were unschooled, ordinary men, they were astonished and they took note that these men had been with Jesus.
ACTS|4|14|But since they could see the man who had been healed standing there with them, there was nothing they could say.
ACTS|4|15|So they ordered them to withdraw from the Sanhedrin and then conferred together.
ACTS|4|16|"What are we going to do with these men?" they asked. "Everybody living in Jerusalem knows they have done an outstanding miracle, and we cannot deny it.
ACTS|4|17|But to stop this thing from spreading any further among the people, we must warn these men to speak no longer to anyone in this name."
ACTS|4|18|Then they called them in again and commanded them not to speak or teach at all in the name of Jesus.
ACTS|4|19|But Peter and John replied, "Judge for yourselves whether it is right in God's sight to obey you rather than God.
ACTS|4|20|For we cannot help speaking about what we have seen and heard."
ACTS|4|21|After further threats they let them go. They could not decide how to punish them, because all the people were praising God for what had happened.
ACTS|4|22|For the man who was miraculously healed was over forty years old.
ACTS|4|23|On their release, Peter and John went back to their own people and reported all that the chief priests and elders had said to them.
ACTS|4|24|When they heard this, they raised their voices together in prayer to God. "Sovereign Lord," they said, "you made the heaven and the earth and the sea, and everything in them.
ACTS|4|25|You spoke by the Holy Spirit through the mouth of your servant, our father David: "'Why do the nations rage and the peoples plot in vain?
ACTS|4|26|The kings of the earth take their stand and the rulers gather together against the Lord and against his Anointed One. '
ACTS|4|27|Indeed Herod and Pontius Pilate met together with the Gentiles and the people of Israel in this city to conspire against your holy servant Jesus, whom you anointed.
ACTS|4|28|They did what your power and will had decided beforehand should happen.
ACTS|4|29|Now, Lord, consider their threats and enable your servants to speak your word with great boldness.
ACTS|4|30|Stretch out your hand to heal and perform miraculous signs and wonders through the name of your holy servant Jesus."
ACTS|4|31|After they prayed, the place where they were meeting was shaken. And they were all filled with the Holy Spirit and spoke the word of God boldly.
ACTS|4|32|All the believers were one in heart and mind. No one claimed that any of his possessions was his own, but they shared everything they had.
ACTS|4|33|With great power the apostles continued to testify to the resurrection of the Lord Jesus, and much grace was upon them all.
ACTS|4|34|There were no needy persons among them. For from time to time those who owned lands or houses sold them, brought the money from the sales
ACTS|4|35|and put it at the apostles' feet, and it was distributed to anyone as he had need.
ACTS|4|36|Joseph, a Levite from Cyprus, whom the apostles called Barnabas (which means Son of Encouragement),
ACTS|4|37|sold a field he owned and brought the money and put it at the apostles' feet.
ACTS|5|1|Now a man named Ananias, together with his wife Sapphira, also sold a piece of property.
ACTS|5|2|With his wife's full knowledge he kept back part of the money for himself, but brought the rest and put it at the apostles' feet.
ACTS|5|3|Then Peter said, "Ananias, how is it that Satan has so filled your heart that you have lied to the Holy Spirit and have kept for yourself some of the money you received for the land?
ACTS|5|4|Didn't it belong to you before it was sold? And after it was sold, wasn't the money at your disposal? What made you think of doing such a thing? You have not lied to men but to God."
ACTS|5|5|When Ananias heard this, he fell down and died. And great fear seized all who heard what had happened.
ACTS|5|6|Then the young men came forward, wrapped up his body, and carried him out and buried him.
ACTS|5|7|About three hours later his wife came in, not knowing what had happened.
ACTS|5|8|Peter asked her, "Tell me, is this the price you and Ananias got for the land?Yes," she said, "that is the price."
ACTS|5|9|Peter said to her, "How could you agree to test the Spirit of the Lord? Look! The feet of the men who buried your husband are at the door, and they will carry you out also."
ACTS|5|10|At that moment she fell down at his feet and died. Then the young men came in and, finding her dead, carried her out and buried her beside her husband.
ACTS|5|11|Great fear seized the whole church and all who heard about these events.
ACTS|5|12|The apostles performed many miraculous signs and wonders among the people. And all the believers used to meet together in Solomon's Colonnade.
ACTS|5|13|No one else dared join them, even though they were highly regarded by the people.
ACTS|5|14|Nevertheless, more and more men and women believed in the Lord and were added to their number.
ACTS|5|15|As a result, people brought the sick into the streets and laid them on beds and mats so that at least Peter's shadow might fall on some of them as he passed by.
ACTS|5|16|Crowds gathered also from the towns around Jerusalem, bringing their sick and those tormented by evil spirits, and all of them were healed.
ACTS|5|17|Then the high priest and all his associates, who were members of the party of the Sadducees, were filled with jealousy.
ACTS|5|18|They arrested the apostles and put them in the public jail.
ACTS|5|19|But during the night an angel of the Lord opened the doors of the jail and brought them out.
ACTS|5|20|"Go, stand in the temple courts," he said, "and tell the people the full message of this new life."
ACTS|5|21|At daybreak they entered the temple courts, as they had been told, and began to teach the people.
ACTS|5|22|When the high priest and his associates arrived, they called together the Sanhedrin--the full assembly of the elders of Israel--and sent to the jail for the apostles. But on arriving at the jail, the officers did not find them there. So they went back and reported,
ACTS|5|23|"We found the jail securely locked, with the guards standing at the doors; but when we opened them, we found no one inside."
ACTS|5|24|On hearing this report, the captain of the temple guard and the chief priests were puzzled, wondering what would come of this.
ACTS|5|25|Then someone came and said, "Look! The men you put in jail are standing in the temple courts teaching the people."
ACTS|5|26|At that, the captain went with his officers and brought the apostles. They did not use force, because they feared that the people would stone them.
ACTS|5|27|Having brought the apostles, they made them appear before the Sanhedrin to be questioned by the high priest.
ACTS|5|28|"We gave you strict orders not to teach in this name," he said. "Yet you have filled Jerusalem with your teaching and are determined to make us guilty of this man's blood."
ACTS|5|29|Peter and the other apostles replied: "We must obey God rather than men!
ACTS|5|30|The God of our fathers raised Jesus from the dead--whom you had killed by hanging him on a tree.
ACTS|5|31|God exalted him to his own right hand as Prince and Savior that he might give repentance and forgiveness of sins to Israel.
ACTS|5|32|We are witnesses of these things, and so is the Holy Spirit, whom God has given to those who obey him."
ACTS|5|33|When they heard this, they were furious and wanted to put them to death.
ACTS|5|34|But a Pharisee named Gamaliel, a teacher of the law, who was honored by all the people, stood up in the Sanhedrin and ordered that the men be put outside for a little while.
ACTS|5|35|Then he addressed them: "Men of Israel, consider carefully what you intend to do to these men.
ACTS|5|36|Some time ago Theudas appeared, claiming to be somebody, and about four hundred men rallied to him. He was killed, all his followers were dispersed, and it all came to nothing.
ACTS|5|37|After him, Judas the Galilean appeared in the days of the census and led a band of people in revolt. He too was killed, and all his followers were scattered.
ACTS|5|38|Therefore, in the present case I advise you: Leave these men alone! Let them go! For if their purpose or activity is of human origin, it will fail.
ACTS|5|39|But if it is from God, you will not be able to stop these men; you will only find yourselves fighting against God."
ACTS|5|40|His speech persuaded them. They called the apostles in and had them flogged. Then they ordered them not to speak in the name of Jesus, and let them go.
ACTS|5|41|The apostles left the Sanhedrin, rejoicing because they had been counted worthy of suffering disgrace for the Name.
ACTS|5|42|Day after day, in the temple courts and from house to house, they never stopped teaching and proclaiming the good news that Jesus is the Christ.
ACTS|6|1|In those days when the number of disciples was increasing, the Grecian Jews among them complained against the Hebraic Jews because their widows were being overlooked in the daily distribution of food.
ACTS|6|2|So the Twelve gathered all the disciples together and said, "It would not be right for us to neglect the ministry of the word of God in order to wait on tables.
ACTS|6|3|Brothers, choose seven men from among you who are known to be full of the Spirit and wisdom. We will turn this responsibility over to them
ACTS|6|4|and will give our attention to prayer and the ministry of the word."
ACTS|6|5|This proposal pleased the whole group. They chose Stephen, a man full of faith and of the Holy Spirit; also Philip, Procorus, Nicanor, Timon, Parmenas, and Nicolas from Antioch, a convert to Judaism.
ACTS|6|6|They presented these men to the apostles, who prayed and laid their hands on them.
ACTS|6|7|So the word of God spread. The number of disciples in Jerusalem increased rapidly, and a large number of priests became obedient to the faith.
ACTS|6|8|Now Stephen, a man full of God's grace and power, did great wonders and miraculous signs among the people.
ACTS|6|9|Opposition arose, however, from members of the Synagogue of the Freedmen (as it was called)--Jews of Cyrene and Alexandria as well as the provinces of Cilicia and Asia. These men began to argue with Stephen,
ACTS|6|10|but they could not stand up against his wisdom or the Spirit by whom he spoke.
ACTS|6|11|Then they secretly persuaded some men to say, "We have heard Stephen speak words of blasphemy against Moses and against God."
ACTS|6|12|So they stirred up the people and the elders and the teachers of the law. They seized Stephen and brought him before the Sanhedrin.
ACTS|6|13|They produced false witnesses, who testified, "This fellow never stops speaking against this holy place and against the law.
ACTS|6|14|For we have heard him say that this Jesus of Nazareth will destroy this place and change the customs Moses handed down to us."
ACTS|6|15|All who were sitting in the Sanhedrin looked intently at Stephen, and they saw that his face was like the face of an angel.
ACTS|7|1|Then the high priest asked him, "Are these charges true?"
ACTS|7|2|To this he replied: "Brothers and fathers, listen to me! The God of glory appeared to our father Abraham while he was still in Mesopotamia, before he lived in Haran.
ACTS|7|3|'Leave your country and your people,' God said, 'and go to the land I will show you.'
ACTS|7|4|"So he left the land of the Chaldeans and settled in Haran. After the death of his father, God sent him to this land where you are now living.
ACTS|7|5|He gave him no inheritance here, not even a foot of ground. But God promised him that he and his descendants after him would possess the land, even though at that time Abraham had no child.
ACTS|7|6|God spoke to him in this way: 'Your descendants will be strangers in a country not their own, and they will be enslaved and mistreated four hundred years.
ACTS|7|7|But I will punish the nation they serve as slaves,' God said, 'and afterward they will come out of that country and worship me in this place.'
ACTS|7|8|Then he gave Abraham the covenant of circumcision. And Abraham became the father of Isaac and circumcised him eight days after his birth. Later Isaac became the father of Jacob, and Jacob became the father of the twelve patriarchs.
ACTS|7|9|"Because the patriarchs were jealous of Joseph, they sold him as a slave into Egypt. But God was with him
ACTS|7|10|and rescued him from all his troubles. He gave Joseph wisdom and enabled him to gain the goodwill of Pharaoh king of Egypt; so he made him ruler over Egypt and all his palace.
ACTS|7|11|"Then a famine struck all Egypt and Canaan, bringing great suffering, and our fathers could not find food.
ACTS|7|12|When Jacob heard that there was grain in Egypt, he sent our fathers on their first visit.
ACTS|7|13|On their second visit, Joseph told his brothers who he was, and Pharaoh learned about Joseph's family.
ACTS|7|14|After this, Joseph sent for his father Jacob and his whole family, seventy-five in all.
ACTS|7|15|Then Jacob went down to Egypt, where he and our fathers died.
ACTS|7|16|Their bodies were brought back to Shechem and placed in the tomb that Abraham had bought from the sons of Hamor at Shechem for a certain sum of money.
ACTS|7|17|"As the time drew near for God to fulfill his promise to Abraham, the number of our people in Egypt greatly increased.
ACTS|7|18|Then another king, who knew nothing about Joseph, became ruler of Egypt.
ACTS|7|19|He dealt treacherously with our people and oppressed our forefathers by forcing them to throw out their newborn babies so that they would die.
ACTS|7|20|"At that time Moses was born, and he was no ordinary child. For three months he was cared for in his father's house.
ACTS|7|21|When he was placed outside, Pharaoh's daughter took him and brought him up as her own son.
ACTS|7|22|Moses was educated in all the wisdom of the Egyptians and was powerful in speech and action.
ACTS|7|23|"When Moses was forty years old, he decided to visit his fellow Israelites.
ACTS|7|24|He saw one of them being mistreated by an Egyptian, so he went to his defense and avenged him by killing the Egyptian.
ACTS|7|25|Moses thought that his own people would realize that God was using him to rescue them, but they did not.
ACTS|7|26|The next day Moses came upon two Israelites who were fighting. He tried to reconcile them by saying, 'Men, you are brothers; why do you want to hurt each other?'
ACTS|7|27|"But the man who was mistreating the other pushed Moses aside and said, 'Who made you ruler and judge over us?
ACTS|7|28|Do you want to kill me as you killed the Egyptian yesterday?'
ACTS|7|29|When Moses heard this, he fled to Midian, where he settled as a foreigner and had two sons.
ACTS|7|30|"After forty years had passed, an angel appeared to Moses in the flames of a burning bush in the desert near Mount Sinai.
ACTS|7|31|When he saw this, he was amazed at the sight. As he went over to look more closely, he heard the Lord's voice:
ACTS|7|32|'I am the God of your fathers, the God of Abraham, Isaac and Jacob.' Moses trembled with fear and did not dare to look.
ACTS|7|33|"Then the Lord said to him, 'Take off your sandals; the place where you are standing is holy ground.
ACTS|7|34|I have indeed seen the oppression of my people in Egypt. I have heard their groaning and have come down to set them free. Now come, I will send you back to Egypt.'
ACTS|7|35|"This is the same Moses whom they had rejected with the words, 'Who made you ruler and judge?' He was sent to be their ruler and deliverer by God himself, through the angel who appeared to him in the bush.
ACTS|7|36|He led them out of Egypt and did wonders and miraculous signs in Egypt, at the Red Sea and for forty years in the desert.
ACTS|7|37|"This is that Moses who told the Israelites, 'God will send you a prophet like me from your own people.'
ACTS|7|38|He was in the assembly in the desert, with the angel who spoke to him on Mount Sinai, and with our fathers; and he received living words to pass on to us.
ACTS|7|39|"But our fathers refused to obey him. Instead, they rejected him and in their hearts turned back to Egypt.
ACTS|7|40|They told Aaron, 'Make us gods who will go before us. As for this fellow Moses who led us out of Egypt--we don't know what has happened to him!'
ACTS|7|41|That was the time they made an idol in the form of a calf. They brought sacrifices to it and held a celebration in honor of what their hands had made.
ACTS|7|42|But God turned away and gave them over to the worship of the heavenly bodies. This agrees with what is written in the book of the prophets: "'Did you bring me sacrifices and offerings forty years in the desert, O house of Israel?
ACTS|7|43|You have lifted up the shrine of Molech and the star of your god Rephan, the idols you made to worship. Therefore I will send you into exile' beyond Babylon.
ACTS|7|44|"Our forefathers had the tabernacle of the Testimony with them in the desert. It had been made as God directed Moses, according to the pattern he had seen.
ACTS|7|45|Having received the tabernacle, our fathers under Joshua brought it with them when they took the land from the nations God drove out before them. It remained in the land until the time of David,
ACTS|7|46|who enjoyed God's favor and asked that he might provide a dwelling place for the God of Jacob.
ACTS|7|47|But it was Solomon who built the house for him.
ACTS|7|48|"However, the Most High does not live in houses made by men. As the prophet says:
ACTS|7|49|"'Heaven is my throne, and the earth is my footstool. What kind of house will you build for me? says the Lord. Or where will my resting place be?
ACTS|7|50|Has not my hand made all these things?'
ACTS|7|51|"You stiff-necked people, with uncircumcised hearts and ears! You are just like your fathers: You always resist the Holy Spirit!
ACTS|7|52|Was there ever a prophet your fathers did not persecute? They even killed those who predicted the coming of the Righteous One. And now you have betrayed and murdered him--
ACTS|7|53|you who have received the law that was put into effect through angels but have not obeyed it."
ACTS|7|54|When they heard this, they were furious and gnashed their teeth at him.
ACTS|7|55|But Stephen, full of the Holy Spirit, looked up to heaven and saw the glory of God, and Jesus standing at the right hand of God.
ACTS|7|56|"Look," he said, "I see heaven open and the Son of Man standing at the right hand of God."
ACTS|7|57|At this they covered their ears and, yelling at the top of their voices, they all rushed at him,
ACTS|7|58|dragged him out of the city and began to stone him. Meanwhile, the witnesses laid their clothes at the feet of a young man named Saul.
ACTS|7|59|While they were stoning him, Stephen prayed, "Lord Jesus, receive my spirit."
ACTS|7|60|Then he fell on his knees and cried out, "Lord, do not hold this sin against them." When he had said this, he fell asleep.
ACTS|8|1|And Saul was there, giving approval to his death.
ACTS|8|2|On that day a great persecution broke out against the church at Jerusalem, and all except the apostles were scattered throughout Judea and Samaria. Godly men buried Stephen and mourned deeply for him.
ACTS|8|3|But Saul began to destroy the church. Going from house to house, he dragged off men and women and put them in prison.
ACTS|8|4|Those who had been scattered preached the word wherever they went.
ACTS|8|5|Philip went down to a city in Samaria and proclaimed the Christ there.
ACTS|8|6|When the crowds heard Philip and saw the miraculous signs he did, they all paid close attention to what he said.
ACTS|8|7|With shrieks, evil spirits came out of many, and many paralytics and cripples were healed.
ACTS|8|8|So there was great joy in that city.
ACTS|8|9|Now for some time a man named Simon had practiced sorcery in the city and amazed all the people of Samaria. He boasted that he was someone great,
ACTS|8|10|and all the people, both high and low, gave him their attention and exclaimed, "This man is the divine power known as the Great Power."
ACTS|8|11|They followed him because he had amazed them for a long time with his magic.
ACTS|8|12|But when they believed Philip as he preached the good news of the kingdom of God and the name of Jesus Christ, they were baptized, both men and women.
ACTS|8|13|Simon himself believed and was baptized. And he followed Philip everywhere, astonished by the great signs and miracles he saw.
ACTS|8|14|When the apostles in Jerusalem heard that Samaria had accepted the word of God, they sent Peter and John to them.
ACTS|8|15|When they arrived, they prayed for them that they might receive the Holy Spirit,
ACTS|8|16|because the Holy Spirit had not yet come upon any of them; they had simply been baptized into the name of the Lord Jesus.
ACTS|8|17|Then Peter and John placed their hands on them, and they received the Holy Spirit.
ACTS|8|18|When Simon saw that the Spirit was given at the laying on of the apostles' hands, he offered them money
ACTS|8|19|and said, "Give me also this ability so that everyone on whom I lay my hands may receive the Holy Spirit."
ACTS|8|20|Peter answered: "May your money perish with you, because you thought you could buy the gift of God with money!
ACTS|8|21|You have no part or share in this ministry, because your heart is not right before God.
ACTS|8|22|Repent of this wickedness and pray to the Lord. Perhaps he will forgive you for having such a thought in your heart.
ACTS|8|23|For I see that you are full of bitterness and captive to sin."
ACTS|8|24|Then Simon answered, "Pray to the Lord for me so that nothing you have said may happen to me."
ACTS|8|25|When they had testified and proclaimed the word of the Lord, Peter and John returned to Jerusalem, preaching the gospel in many Samaritan villages.
ACTS|8|26|Now an angel of the Lord said to Philip, "Go south to the road--the desert road--that goes down from Jerusalem to Gaza."
ACTS|8|27|So he started out, and on his way he met an Ethiopian eunuch, an important official in charge of all the treasury of Candace, queen of the Ethiopians. This man had gone to Jerusalem to worship,
ACTS|8|28|and on his way home was sitting in his chariot reading the book of Isaiah the prophet.
ACTS|8|29|The Spirit told Philip, "Go to that chariot and stay near it."
ACTS|8|30|Then Philip ran up to the chariot and heard the man reading Isaiah the prophet. "Do you understand what you are reading?" Philip asked.
ACTS|8|31|"How can I," he said, "unless someone explains it to me?" So he invited Philip to come up and sit with him.
ACTS|8|32|The eunuch was reading this passage of Scripture: "He was led like a sheep to the slaughter, and as a lamb before the shearer is silent, so he did not open his mouth.
ACTS|8|33|In his humiliation he was deprived of justice. Who can speak of his descendants? For his life was taken from the earth."
ACTS|8|34|The eunuch asked Philip, "Tell me, please, who is the prophet talking about, himself or someone else?"
ACTS|8|35|Then Philip began with that very passage of Scripture and told him the good news about Jesus.
ACTS|8|36|As they traveled along the road, they came to some water and the eunuch said, "Look, here is water. Why shouldn't I be baptized?"
ACTS|8|37|See Footnote
ACTS|8|38|And he gave orders to stop the chariot. Then both Philip and the eunuch went down into the water and Philip baptized him.
ACTS|8|39|When they came up out of the water, the Spirit of the Lord suddenly took Philip away, and the eunuch did not see him again, but went on his way rejoicing.
ACTS|8|40|Philip, however, appeared at Azotus and traveled about, preaching the gospel in all the towns until he reached Caesarea.
ACTS|9|1|Meanwhile, Saul was still breathing out murderous threats against the Lord's disciples. He went to the high priest
ACTS|9|2|and asked him for letters to the synagogues in Damascus, so that if he found any there who belonged to the Way, whether men or women, he might take them as prisoners to Jerusalem.
ACTS|9|3|As he neared Damascus on his journey, suddenly a light from heaven flashed around him.
ACTS|9|4|He fell to the ground and heard a voice say to him, "Saul, Saul, why do you persecute me?"
ACTS|9|5|"Who are you, Lord?" Saul asked.
ACTS|9|6|"I am Jesus, whom you are persecuting," he replied. "Now get up and go into the city, and you will be told what you must do."
ACTS|9|7|The men traveling with Saul stood there speechless; they heard the sound but did not see anyone.
ACTS|9|8|Saul got up from the ground, but when he opened his eyes he could see nothing. So they led him by the hand into Damascus.
ACTS|9|9|For three days he was blind, and did not eat or drink anything.
ACTS|9|10|In Damascus there was a disciple named Ananias. The Lord called to him in a vision, "Ananias!Yes, Lord," he answered.
ACTS|9|11|The Lord told him, "Go to the house of Judas on Straight Street and ask for a man from Tarsus named Saul, for he is praying.
ACTS|9|12|In a vision he has seen a man named Ananias come and place his hands on him to restore his sight."
ACTS|9|13|"Lord," Ananias answered, "I have heard many reports about this man and all the harm he has done to your saints in Jerusalem.
ACTS|9|14|And he has come here with authority from the chief priests to arrest all who call on your name."
ACTS|9|15|But the Lord said to Ananias, "Go! This man is my chosen instrument to carry my name before the Gentiles and their kings and before the people of Israel.
ACTS|9|16|I will show him how much he must suffer for my name."
ACTS|9|17|Then Ananias went to the house and entered it. Placing his hands on Saul, he said, "Brother Saul, the Lord--Jesus, who appeared to you on the road as you were coming here--has sent me so that you may see again and be filled with the Holy Spirit."
ACTS|9|18|Immediately, something like scales fell from Saul's eyes, and he could see again. He got up and was baptized,
ACTS|9|19|and after taking some food, he regained his strength.
ACTS|9|20|Saul spent several days with the disciples in Damascus. At once he began to preach in the synagogues that Jesus is the Son of God.
ACTS|9|21|All those who heard him were astonished and asked, "Isn't he the man who raised havoc in Jerusalem among those who call on this name? And hasn't he come here to take them as prisoners to the chief priests?"
ACTS|9|22|Yet Saul grew more and more powerful and baffled the Jews living in Damascus by proving that Jesus is the Christ.
ACTS|9|23|After many days had gone by, the Jews conspired to kill him,
ACTS|9|24|but Saul learned of their plan. Day and night they kept close watch on the city gates in order to kill him.
ACTS|9|25|But his followers took him by night and lowered him in a basket through an opening in the wall.
ACTS|9|26|When he came to Jerusalem, he tried to join the disciples, but they were all afraid of him, not believing that he really was a disciple.
ACTS|9|27|But Barnabas took him and brought him to the apostles. He told them how Saul on his journey had seen the Lord and that the Lord had spoken to him, and how in Damascus he had preached fearlessly in the name of Jesus.
ACTS|9|28|So Saul stayed with them and moved about freely in Jerusalem, speaking boldly in the name of the Lord.
ACTS|9|29|He talked and debated with the Grecian Jews, but they tried to kill him.
ACTS|9|30|When the brothers learned of this, they took him down to Caesarea and sent him off to Tarsus.
ACTS|9|31|Then the church throughout Judea, Galilee and Samaria enjoyed a time of peace. It was strengthened; and encouraged by the Holy Spirit, it grew in numbers, living in the fear of the Lord.
ACTS|9|32|As Peter traveled about the country, he went to visit the saints in Lydda.
ACTS|9|33|There he found a man named Aeneas, a paralytic who had been bedridden for eight years.
ACTS|9|34|"Aeneas," Peter said to him, "Jesus Christ heals you. Get up and take care of your mat." Immediately Aeneas got up.
ACTS|9|35|All those who lived in Lydda and Sharon saw him and turned to the Lord.
ACTS|9|36|In Joppa there was a disciple named Tabitha (which, when translated, is Dorcas ), who was always doing good and helping the poor.
ACTS|9|37|About that time she became sick and died, and her body was washed and placed in an upstairs room.
ACTS|9|38|Lydda was near Joppa; so when the disciples heard that Peter was in Lydda, they sent two men to him and urged him, "Please come at once!"
ACTS|9|39|Peter went with them, and when he arrived he was taken upstairs to the room. All the widows stood around him, crying and showing him the robes and other clothing that Dorcas had made while she was still with them.
ACTS|9|40|Peter sent them all out of the room; then he got down on his knees and prayed. Turning toward the dead woman, he said, "Tabitha, get up." She opened her eyes, and seeing Peter she sat up.
ACTS|9|41|He took her by the hand and helped her to her feet. Then he called the believers and the widows and presented her to them alive.
ACTS|9|42|This became known all over Joppa, and many people believed in the Lord.
ACTS|9|43|Peter stayed in Joppa for some time with a tanner named Simon.
ACTS|10|1|At Caesarea there was a man named Cornelius, a centurion in what was known as the Italian Regiment.
ACTS|10|2|He and all his family were devout and God-fearing; he gave generously to those in need and prayed to God regularly.
ACTS|10|3|One day at about three in the afternoon he had a vision. He distinctly saw an angel of God, who came to him and said, "Cornelius!"
ACTS|10|4|Cornelius stared at him in fear. "What is it, Lord?" he asked.
ACTS|10|5|The angel answered, "Your prayers and gifts to the poor have come up as a memorial offering before God. Now send men to Joppa to bring back a man named Simon who is called Peter.
ACTS|10|6|He is staying with Simon the tanner, whose house is by the sea."
ACTS|10|7|When the angel who spoke to him had gone, Cornelius called two of his servants and a devout soldier who was one of his attendants.
ACTS|10|8|He told them everything that had happened and sent them to Joppa.
ACTS|10|9|About noon the following day as they were on their journey and approaching the city, Peter went up on the roof to pray.
ACTS|10|10|He became hungry and wanted something to eat, and while the meal was being prepared, he fell into a trance.
ACTS|10|11|He saw heaven opened and something like a large sheet being let down to earth by its four corners.
ACTS|10|12|It contained all kinds of four-footed animals, as well as reptiles of the earth and birds of the air.
ACTS|10|13|Then a voice told him, "Get up, Peter. Kill and eat."
ACTS|10|14|"Surely not, Lord!" Peter replied. "I have never eaten anything impure or unclean."
ACTS|10|15|The voice spoke to him a second time, "Do not call anything impure that God has made clean."
ACTS|10|16|This happened three times, and immediately the sheet was taken back to heaven.
ACTS|10|17|While Peter was wondering about the meaning of the vision, the men sent by Cornelius found out where Simon's house was and stopped at the gate.
ACTS|10|18|They called out, asking if Simon who was known as Peter was staying there.
ACTS|10|19|While Peter was still thinking about the vision, the Spirit said to him, "Simon, three men are looking for you.
ACTS|10|20|So get up and go downstairs. Do not hesitate to go with them, for I have sent them."
ACTS|10|21|Peter went down and said to the men, "I'm the one you're looking for. Why have you come?"
ACTS|10|22|The men replied, "We have come from Cornelius the centurion. He is a righteous and God-fearing man, who is respected by all the Jewish people. A holy angel told him to have you come to his house so that he could hear what you have to say."
ACTS|10|23|Then Peter invited the men into the house to be his guests.
ACTS|10|24|The next day Peter started out with them, and some of the brothers from Joppa went along. The following day he arrived in Caesarea. Cornelius was expecting them and had called together his relatives and close friends.
ACTS|10|25|As Peter entered the house, Cornelius met him and fell at his feet in reverence.
ACTS|10|26|But Peter made him get up. "Stand up," he said, "I am only a man myself."
ACTS|10|27|Talking with him, Peter went inside and found a large gathering of people.
ACTS|10|28|He said to them: "You are well aware that it is against our law for a Jew to associate with a Gentile or visit him. But God has shown me that I should not call any man impure or unclean.
ACTS|10|29|So when I was sent for, I came without raising any objection. May I ask why you sent for me?"
ACTS|10|30|Cornelius answered: "Four days ago I was in my house praying at this hour, at three in the afternoon. Suddenly a man in shining clothes stood before me
ACTS|10|31|and said, 'Cornelius, God has heard your prayer and remembered your gifts to the poor.
ACTS|10|32|Send to Joppa for Simon who is called Peter. He is a guest in the home of Simon the tanner, who lives by the sea.'
ACTS|10|33|So I sent for you immediately, and it was good of you to come. Now we are all here in the presence of God to listen to everything the Lord has commanded you to tell us."
ACTS|10|34|Then Peter began to speak: "I now realize how true it is that God does not show favoritism
ACTS|10|35|but accepts men from every nation who fear him and do what is right.
ACTS|10|36|You know the message God sent to the people of Israel, telling the good news of peace through Jesus Christ, who is Lord of all.
ACTS|10|37|You know what has happened throughout Judea, beginning in Galilee after the baptism that John preached--
ACTS|10|38|how God anointed Jesus of Nazareth with the Holy Spirit and power, and how he went around doing good and healing all who were under the power of the devil, because God was with him.
ACTS|10|39|"We are witnesses of everything he did in the country of the Jews and in Jerusalem. They killed him by hanging him on a tree,
ACTS|10|40|but God raised him from the dead on the third day and caused him to be seen.
ACTS|10|41|He was not seen by all the people, but by witnesses whom God had already chosen--by us who ate and drank with him after he rose from the dead.
ACTS|10|42|He commanded us to preach to the people and to testify that he is the one whom God appointed as judge of the living and the dead.
ACTS|10|43|All the prophets testify about him that everyone who believes in him receives forgiveness of sins through his name."
ACTS|10|44|While Peter was still speaking these words, the Holy Spirit came on all who heard the message.
ACTS|10|45|The circumcised believers who had come with Peter were astonished that the gift of the Holy Spirit had been poured out even on the Gentiles.
ACTS|10|46|For they heard them speaking in tongues and praising God.
ACTS|10|47|Then Peter said, "Can anyone keep these people from being baptized with water? They have received the Holy Spirit just as we have."
ACTS|10|48|So he ordered that they be baptized in the name of Jesus Christ. Then they asked Peter to stay with them for a few days.
ACTS|11|1|The apostles and the brothers throughout Judea heard that the Gentiles also had received the word of God.
ACTS|11|2|So when Peter went up to Jerusalem, the circumcised believers criticized him
ACTS|11|3|and said, "You went into the house of uncircumcised men and ate with them."
ACTS|11|4|Peter began and explained everything to them precisely as it had happened:
ACTS|11|5|"I was in the city of Joppa praying, and in a trance I saw a vision. I saw something like a large sheet being let down from heaven by its four corners, and it came down to where I was.
ACTS|11|6|I looked into it and saw four-footed animals of the earth, wild beasts, reptiles, and birds of the air.
ACTS|11|7|Then I heard a voice telling me, 'Get up, Peter. Kill and eat.'
ACTS|11|8|"I replied, 'Surely not, Lord! Nothing impure or unclean has ever entered my mouth.'
ACTS|11|9|"The voice spoke from heaven a second time, 'Do not call anything impure that God has made clean.'
ACTS|11|10|This happened three times, and then it was all pulled up to heaven again.
ACTS|11|11|"Right then three men who had been sent to me from Caesarea stopped at the house where I was staying.
ACTS|11|12|The Spirit told me to have no hesitation about going with them. These six brothers also went with me, and we entered the man's house.
ACTS|11|13|He told us how he had seen an angel appear in his house and say, 'Send to Joppa for Simon who is called Peter.
ACTS|11|14|He will bring you a message through which you and all your household will be saved.'
ACTS|11|15|"As I began to speak, the Holy Spirit came on them as he had come on us at the beginning.
ACTS|11|16|Then I remembered what the Lord had said: 'John baptized with water, but you will be baptized with the Holy Spirit.'
ACTS|11|17|So if God gave them the same gift as he gave us, who believed in the Lord Jesus Christ, who was I to think that I could oppose God?"
ACTS|11|18|When they heard this, they had no further objections and praised God, saying, "So then, God has granted even the Gentiles repentance unto life."
ACTS|11|19|Now those who had been scattered by the persecution in connection with Stephen traveled as far as Phoenicia, Cyprus and Antioch, telling the message only to Jews.
ACTS|11|20|Some of them, however, men from Cyprus and Cyrene, went to Antioch and began to speak to Greeks also, telling them the good news about the Lord Jesus.
ACTS|11|21|The Lord's hand was with them, and a great number of people believed and turned to the Lord.
ACTS|11|22|News of this reached the ears of the church at Jerusalem, and they sent Barnabas to Antioch.
ACTS|11|23|When he arrived and saw the evidence of the grace of God, he was glad and encouraged them all to remain true to the Lord with all their hearts.
ACTS|11|24|He was a good man, full of the Holy Spirit and faith, and a great number of people were brought to the Lord.
ACTS|11|25|Then Barnabas went to Tarsus to look for Saul,
ACTS|11|26|and when he found him, he brought him to Antioch. So for a whole year Barnabas and Saul met with the church and taught great numbers of people. The disciples were called Christians first at Antioch.
ACTS|11|27|During this time some prophets came down from Jerusalem to Antioch.
ACTS|11|28|One of them, named Agabus, stood up and through the Spirit predicted that a severe famine would spread over the entire Roman world. (This happened during the reign of Claudius.)
ACTS|11|29|The disciples, each according to his ability, decided to provide help for the brothers living in Judea.
ACTS|11|30|This they did, sending their gift to the elders by Barnabas and Saul.
ACTS|12|1|It was about this time that King Herod arrested some who belonged to the church, intending to persecute them.
ACTS|12|2|He had James, the brother of John, put to death with the sword.
ACTS|12|3|When he saw that this pleased the Jews, he proceeded to seize Peter also. This happened during the Feast of Unleavened Bread.
ACTS|12|4|After arresting him, he put him in prison, handing him over to be guarded by four squads of four soldiers each. Herod intended to bring him out for public trial after the Passover.
ACTS|12|5|So Peter was kept in prison, but the church was earnestly praying to God for him.
ACTS|12|6|The night before Herod was to bring him to trial, Peter was sleeping between two soldiers, bound with two chains, and sentries stood guard at the entrance.
ACTS|12|7|Suddenly an angel of the Lord appeared and a light shone in the cell. He struck Peter on the side and woke him up. "Quick, get up!" he said, and the chains fell off Peter's wrists.
ACTS|12|8|Then the angel said to him, "Put on your clothes and sandals." And Peter did so. "Wrap your cloak around you and follow me," the angel told him.
ACTS|12|9|Peter followed him out of the prison, but he had no idea that what the angel was doing was really happening; he thought he was seeing a vision.
ACTS|12|10|They passed the first and second guards and came to the iron gate leading to the city. It opened for them by itself, and they went through it. When they had walked the length of one street, suddenly the angel left him.
ACTS|12|11|Then Peter came to himself and said, "Now I know without a doubt that the Lord sent his angel and rescued me from Herod's clutches and from everything the Jewish people were anticipating."
ACTS|12|12|When this had dawned on him, he went to the house of Mary the mother of John, also called Mark, where many people had gathered and were praying.
ACTS|12|13|Peter knocked at the outer entrance, and a servant girl named Rhoda came to answer the door.
ACTS|12|14|When she recognized Peter's voice, she was so overjoyed she ran back without opening it and exclaimed, "Peter is at the door!"
ACTS|12|15|"You're out of your mind," they told her. When she kept insisting that it was so, they said, "It must be his angel."
ACTS|12|16|But Peter kept on knocking, and when they opened the door and saw him, they were astonished.
ACTS|12|17|Peter motioned with his hand for them to be quiet and described how the Lord had brought him out of prison. "Tell James and the brothers about this," he said, and then he left for another place.
ACTS|12|18|In the morning, there was no small commotion among the soldiers as to what had become of Peter.
ACTS|12|19|After Herod had a thorough search made for him and did not find him, he cross-examined the guards and ordered that they be executed.
ACTS|12|20|Then Herod went from Judea to Caesarea and stayed there a while. He had been quarreling with the people of Tyre and Sidon; they now joined together and sought an audience with him. Having secured the support of Blastus, a trusted personal servant of the king, they asked for peace, because they depended on the king's country for their food supply.
ACTS|12|21|On the appointed day Herod, wearing his royal robes, sat on his throne and delivered a public address to the people.
ACTS|12|22|They shouted, "This is the voice of a god, not of a man."
ACTS|12|23|Immediately, because Herod did not give praise to God, an angel of the Lord struck him down, and he was eaten by worms and died.
ACTS|12|24|But the word of God continued to increase and spread.
ACTS|12|25|When Barnabas and Saul had finished their mission, they returned from Jerusalem, taking with them John, also called Mark.
ACTS|13|1|In the church at Antioch there were prophets and teachers: Barnabas, Simeon called Niger, Lucius of Cyrene, Manaen (who had been brought up with Herod the tetrarch) and Saul.
ACTS|13|2|While they were worshiping the Lord and fasting, the Holy Spirit said, "Set apart for me Barnabas and Saul for the work to which I have called them."
ACTS|13|3|So after they had fasted and prayed, they placed their hands on them and sent them off.
ACTS|13|4|The two of them, sent on their way by the Holy Spirit, went down to Seleucia and sailed from there to Cyprus.
ACTS|13|5|When they arrived at Salamis, they proclaimed the word of God in the Jewish synagogues. John was with them as their helper.
ACTS|13|6|They traveled through the whole island until they came to Paphos. There they met a Jewish sorcerer and false prophet named Bar-Jesus,
ACTS|13|7|who was an attendant of the proconsul, Sergius Paulus. The proconsul, an intelligent man, sent for Barnabas and Saul because he wanted to hear the word of God.
ACTS|13|8|But Elymas the sorcerer (for that is what his name means) opposed them and tried to turn the proconsul from the faith.
ACTS|13|9|Then Saul, who was also called Paul, filled with the Holy Spirit, looked straight at Elymas and said,
ACTS|13|10|"You are a child of the devil and an enemy of everything that is right! You are full of all kinds of deceit and trickery. Will you never stop perverting the right ways of the Lord?
ACTS|13|11|Now the hand of the Lord is against you. You are going to be blind, and for a time you will be unable to see the light of the sun."
ACTS|13|12|Immediately mist and darkness came over him, and he groped about, seeking someone to lead him by the hand. When the proconsul saw what had happened, he believed, for he was amazed at the teaching about the Lord.
ACTS|13|13|From Paphos, Paul and his companions sailed to Perga in Pamphylia, where John left them to return to Jerusalem.
ACTS|13|14|From Perga they went on to Pisidian Antioch. On the Sabbath they entered the synagogue and sat down.
ACTS|13|15|After the reading from the Law and the Prophets, the synagogue rulers sent word to them, saying, "Brothers, if you have a message of encouragement for the people, please speak."
ACTS|13|16|Standing up, Paul motioned with his hand and said: "Men of Israel and you Gentiles who worship God, listen to me!
ACTS|13|17|The God of the people of Israel chose our fathers; he made the people prosper during their stay in Egypt, with mighty power he led them out of that country,
ACTS|13|18|he endured their conduct for about forty years in the desert,
ACTS|13|19|he overthrew seven nations in Canaan and gave their land to his people as their inheritance.
ACTS|13|20|All this took about 450 years.
ACTS|13|21|"After this, God gave them judges until the time of Samuel the prophet. Then the people asked for a king, and he gave them Saul son of Kish, of the tribe of Benjamin, who ruled forty years.
ACTS|13|22|After removing Saul, he made David their king. He testified concerning him: 'I have found David son of Jesse a man after my own heart; he will do everything I want him to do.'
ACTS|13|23|"From this man's descendants God has brought to Israel the Savior Jesus, as he promised.
ACTS|13|24|Before the coming of Jesus, John preached repentance and baptism to all the people of Israel.
ACTS|13|25|As John was completing his work, he said: 'Who do you think I am? I am not that one. No, but he is coming after me, whose sandals I am not worthy to untie.'
ACTS|13|26|"Brothers, children of Abraham, and you God-fearing Gentiles, it is to us that this message of salvation has been sent.
ACTS|13|27|The people of Jerusalem and their rulers did not recognize Jesus, yet in condemning him they fulfilled the words of the prophets that are read every Sabbath.
ACTS|13|28|Though they found no proper ground for a death sentence, they asked Pilate to have him executed.
ACTS|13|29|When they had carried out all that was written about him, they took him down from the tree and laid him in a tomb.
ACTS|13|30|But God raised him from the dead,
ACTS|13|31|and for many days he was seen by those who had traveled with him from Galilee to Jerusalem. They are now his witnesses to our people.
ACTS|13|32|"We tell you the good news: What God promised our fathers
ACTS|13|33|he has fulfilled for us, their children, by raising up Jesus. As it is written in the second Psalm: "'You are my Son; today I have become your Father. '
ACTS|13|34|The fact that God raised him from the dead, never to decay, is stated in these words: "'I will give you the holy and sure blessings promised to David.'
ACTS|13|35|So it is stated elsewhere: "'You will not let your Holy One see decay.'
ACTS|13|36|"For when David had served God's purpose in his own generation, he fell asleep; he was buried with his fathers and his body decayed.
ACTS|13|37|But the one whom God raised from the dead did not see decay.
ACTS|13|38|"Therefore, my brothers, I want you to know that through Jesus the forgiveness of sins is proclaimed to you.
ACTS|13|39|Through him everyone who believes is justified from everything you could not be justified from by the law of Moses.
ACTS|13|40|Take care that what the prophets have said does not happen to you:
ACTS|13|41|"'Look, you scoffers, wonder and perish, for I am going to do something in your days that you would never believe, even if someone told you.'"
ACTS|13|42|As Paul and Barnabas were leaving the synagogue, the people invited them to speak further about these things on the next Sabbath.
ACTS|13|43|When the congregation was dismissed, many of the Jews and devout converts to Judaism followed Paul and Barnabas, who talked with them and urged them to continue in the grace of God.
ACTS|13|44|On the next Sabbath almost the whole city gathered to hear the word of the Lord.
ACTS|13|45|When the Jews saw the crowds, they were filled with jealousy and talked abusively against what Paul was saying.
ACTS|13|46|Then Paul and Barnabas answered them boldly: "We had to speak the word of God to you first. Since you reject it and do not consider yourselves worthy of eternal life, we now turn to the Gentiles.
ACTS|13|47|For this is what the Lord has commanded us: "'I have made you a light for the Gentiles, that you may bring salvation to the ends of the earth.'"
ACTS|13|48|When the Gentiles heard this, they were glad and honored the word of the Lord; and all who were appointed for eternal life believed.
ACTS|13|49|The word of the Lord spread through the whole region.
ACTS|13|50|But the Jews incited the God-fearing women of high standing and the leading men of the city. They stirred up persecution against Paul and Barnabas, and expelled them from their region.
ACTS|13|51|So they shook the dust from their feet in protest against them and went to Iconium.
ACTS|13|52|And the disciples were filled with joy and with the Holy Spirit.
ACTS|14|1|At Iconium Paul and Barnabas went as usual into the Jewish synagogue. There they spoke so effectively that a great number of Jews and Gentiles believed.
ACTS|14|2|But the Jews who refused to believe stirred up the Gentiles and poisoned their minds against the brothers.
ACTS|14|3|So Paul and Barnabas spent considerable time there, speaking boldly for the Lord, who confirmed the message of his grace by enabling them to do miraculous signs and wonders.
ACTS|14|4|The people of the city were divided; some sided with the Jews, others with the apostles.
ACTS|14|5|There was a plot afoot among the Gentiles and Jews, together with their leaders, to mistreat them and stone them.
ACTS|14|6|But they found out about it and fled to the Lycaonian cities of Lystra and Derbe and to the surrounding country,
ACTS|14|7|where they continued to preach the good news.
ACTS|14|8|In Lystra there sat a man crippled in his feet, who was lame from birth and had never walked.
ACTS|14|9|He listened to Paul as he was speaking. Paul looked directly at him, saw that he had faith to be healed
ACTS|14|10|and called out, "Stand up on your feet!" At that, the man jumped up and began to walk.
ACTS|14|11|When the crowd saw what Paul had done, they shouted in the Lycaonian language, "The gods have come down to us in human form!"
ACTS|14|12|Barnabas they called Zeus, and Paul they called Hermes because he was the chief speaker.
ACTS|14|13|The priest of Zeus, whose temple was just outside the city, brought bulls and wreaths to the city gates because he and the crowd wanted to offer sacrifices to them.
ACTS|14|14|But when the apostles Barnabas and Paul heard of this, they tore their clothes and rushed out into the crowd, shouting:
ACTS|14|15|"Men, why are you doing this? We too are only men, human like you. We are bringing you good news, telling you to turn from these worthless things to the living God, who made heaven and earth and sea and everything in them.
ACTS|14|16|In the past, he let all nations go their own way.
ACTS|14|17|Yet he has not left himself without testimony: He has shown kindness by giving you rain from heaven and crops in their seasons; he provides you with plenty of food and fills your hearts with joy."
ACTS|14|18|Even with these words, they had difficulty keeping the crowd from sacrificing to them.
ACTS|14|19|Then some Jews came from Antioch and Iconium and won the crowd over. They stoned Paul and dragged him outside the city, thinking he was dead.
ACTS|14|20|But after the disciples had gathered around him, he got up and went back into the city. The next day he and Barnabas left for Derbe.
ACTS|14|21|They preached the good news in that city and won a large number of disciples. Then they returned to Lystra, Iconium and Antioch,
ACTS|14|22|strengthening the disciples and encouraging them to remain true to the faith. "We must go through many hardships to enter the kingdom of God," they said.
ACTS|14|23|Paul and Barnabas appointed elders for them in each church and, with prayer and fasting, committed them to the Lord, in whom they had put their trust.
ACTS|14|24|After going through Pisidia, they came into Pamphylia,
ACTS|14|25|and when they had preached the word in Perga, they went down to Attalia.
ACTS|14|26|From Attalia they sailed back to Antioch, where they had been committed to the grace of God for the work they had now completed.
ACTS|14|27|On arriving there, they gathered the church together and reported all that God had done through them and how he had opened the door of faith to the Gentiles.
ACTS|14|28|And they stayed there a long time with the disciples.
ACTS|15|1|Some men came down from Judea to Antioch and were teaching the brothers: "Unless you are circumcised, according to the custom taught by Moses, you cannot be saved."
ACTS|15|2|This brought Paul and Barnabas into sharp dispute and debate with them. So Paul and Barnabas were appointed, along with some other believers, to go up to Jerusalem to see the apostles and elders about this question.
ACTS|15|3|The church sent them on their way, and as they traveled through Phoenicia and Samaria, they told how the Gentiles had been converted. This news made all the brothers very glad.
ACTS|15|4|When they came to Jerusalem, they were welcomed by the church and the apostles and elders, to whom they reported everything God had done through them.
ACTS|15|5|Then some of the believers who belonged to the party of the Pharisees stood up and said, "The Gentiles must be circumcised and required to obey the law of Moses."
ACTS|15|6|The apostles and elders met to consider this question.
ACTS|15|7|After much discussion, Peter got up and addressed them: "Brothers, you know that some time ago God made a choice among you that the Gentiles might hear from my lips the message of the gospel and believe.
ACTS|15|8|God, who knows the heart, showed that he accepted them by giving the Holy Spirit to them, just as he did to us.
ACTS|15|9|He made no distinction between us and them, for he purified their hearts by faith.
ACTS|15|10|Now then, why do you try to test God by putting on the necks of the disciples a yoke that neither we nor our fathers have been able to bear?
ACTS|15|11|No! We believe it is through the grace of our Lord Jesus that we are saved, just as they are."
ACTS|15|12|The whole assembly became silent as they listened to Barnabas and Paul telling about the miraculous signs and wonders God had done among the Gentiles through them.
ACTS|15|13|When they finished, James spoke up: "Brothers, listen to me.
ACTS|15|14|Simon has described to us how God at first showed his concern by taking from the Gentiles a people for himself.
ACTS|15|15|The words of the prophets are in agreement with this, as it is written:
ACTS|15|16|"'After this I will return and rebuild David's fallen tent. Its ruins I will rebuild, and I will restore it,
ACTS|15|17|that the remnant of men may seek the Lord, and all the Gentiles who bear my name, says the Lord, who does these things'
ACTS|15|18|that have been known for ages.
ACTS|15|19|"It is my judgment, therefore, that we should not make it difficult for the Gentiles who are turning to God.
ACTS|15|20|Instead we should write to them, telling them to abstain from food polluted by idols, from sexual immorality, from the meat of strangled animals and from blood.
ACTS|15|21|For Moses has been preached in every city from the earliest times and is read in the synagogues on every Sabbath."
ACTS|15|22|Then the apostles and elders, with the whole church, decided to choose some of their own men and send them to Antioch with Paul and Barnabas. They chose Judas (called Barsabbas) and Silas, two men who were leaders among the brothers.
ACTS|15|23|With them they sent the following letter: The apostles and elders, your brothers, To the Gentile believers in Antioch, Syria and Cilicia: Greetings.
ACTS|15|24|We have heard that some went out from us without our authorization and disturbed you, troubling your minds by what they said.
ACTS|15|25|So we all agreed to choose some men and send them to you with our dear friends Barnabas and Paul--
ACTS|15|26|men who have risked their lives for the name of our Lord Jesus Christ.
ACTS|15|27|Therefore we are sending Judas and Silas to confirm by word of mouth what we are writing.
ACTS|15|28|It seemed good to the Holy Spirit and to us not to burden you with anything beyond the following requirements:
ACTS|15|29|You are to abstain from food sacrificed to idols, from blood, from the meat of strangled animals and from sexual immorality. You will do well to avoid these things. Farewell.
ACTS|15|30|The men were sent off and went down to Antioch, where they gathered the church together and delivered the letter.
ACTS|15|31|The people read it and were glad for its encouraging message.
ACTS|15|32|Judas and Silas, who themselves were prophets, said much to encourage and strengthen the brothers.
ACTS|15|33|After spending some time there, they were sent off by the brothers with the blessing of peace to return to those who had sent them.
ACTS|15|34|See Footnote
ACTS|15|35|But Paul and Barnabas remained in Antioch, where they and many others taught and preached the word of the Lord.
ACTS|15|36|Some time later Paul said to Barnabas, "Let us go back and visit the brothers in all the towns where we preached the word of the Lord and see how they are doing."
ACTS|15|37|Barnabas wanted to take John, also called Mark, with them,
ACTS|15|38|but Paul did not think it wise to take him, because he had deserted them in Pamphylia and had not continued with them in the work.
ACTS|15|39|They had such a sharp disagreement that they parted company. Barnabas took Mark and sailed for Cyprus,
ACTS|15|40|but Paul chose Silas and left, commended by the brothers to the grace of the Lord.
ACTS|15|41|He went through Syria and Cilicia, strengthening the churches.
ACTS|16|1|He came to Derbe and then to Lystra, where a disciple named Timothy lived, whose mother was a Jewess and a believer, but whose father was a Greek.
ACTS|16|2|The brothers at Lystra and Iconium spoke well of him.
ACTS|16|3|Paul wanted to take him along on the journey, so he circumcised him because of the Jews who lived in that area, for they all knew that his father was a Greek.
ACTS|16|4|As they traveled from town to town, they delivered the decisions reached by the apostles and elders in Jerusalem for the people to obey.
ACTS|16|5|So the churches were strengthened in the faith and grew daily in numbers.
ACTS|16|6|Paul and his companions traveled throughout the region of Phrygia and Galatia, having been kept by the Holy Spirit from preaching the word in the province of Asia.
ACTS|16|7|When they came to the border of Mysia, they tried to enter Bithynia, but the Spirit of Jesus would not allow them to.
ACTS|16|8|So they passed by Mysia and went down to Troas.
ACTS|16|9|During the night Paul had a vision of a man of Macedonia standing and begging him, "Come over to Macedonia and help us."
ACTS|16|10|After Paul had seen the vision, we got ready at once to leave for Macedonia, concluding that God had called us to preach the gospel to them.
ACTS|16|11|From Troas we put out to sea and sailed straight for Samothrace, and the next day on to Neapolis.
ACTS|16|12|From there we traveled to Philippi, a Roman colony and the leading city of that district of Macedonia. And we stayed there several days.
ACTS|16|13|On the Sabbath we went outside the city gate to the river, where we expected to find a place of prayer. We sat down and began to speak to the women who had gathered there.
ACTS|16|14|One of those listening was a woman named Lydia, a dealer in purple cloth from the city of Thyatira, who was a worshiper of God. The Lord opened her heart to respond to Paul's message.
ACTS|16|15|When she and the members of her household were baptized, she invited us to her home. "If you consider me a believer in the Lord," she said, "come and stay at my house." And she persuaded us.
ACTS|16|16|Once when we were going to the place of prayer, we were met by a slave girl who had a spirit by which she predicted the future. She earned a great deal of money for her owners by fortune-telling.
ACTS|16|17|This girl followed Paul and the rest of us, shouting, "These men are servants of the Most High God, who are telling you the way to be saved."
ACTS|16|18|She kept this up for many days. Finally Paul became so troubled that he turned around and said to the spirit, "In the name of Jesus Christ I command you to come out of her!" At that moment the spirit left her.
ACTS|16|19|When the owners of the slave girl realized that their hope of making money was gone, they seized Paul and Silas and dragged them into the marketplace to face the authorities.
ACTS|16|20|They brought them before the magistrates and said, "These men are Jews, and are throwing our city into an uproar
ACTS|16|21|by advocating customs unlawful for us Romans to accept or practice."
ACTS|16|22|The crowd joined in the attack against Paul and Silas, and the magistrates ordered them to be stripped and beaten.
ACTS|16|23|After they had been severely flogged, they were thrown into prison, and the jailer was commanded to guard them carefully.
ACTS|16|24|Upon receiving such orders, he put them in the inner cell and fastened their feet in the stocks.
ACTS|16|25|About midnight Paul and Silas were praying and singing hymns to God, and the other prisoners were listening to them.
ACTS|16|26|Suddenly there was such a violent earthquake that the foundations of the prison were shaken. At once all the prison doors flew open, and everybody's chains came loose.
ACTS|16|27|The jailer woke up, and when he saw the prison doors open, he drew his sword and was about to kill himself because he thought the prisoners had escaped.
ACTS|16|28|But Paul shouted, "Don't harm yourself! We are all here!"
ACTS|16|29|The jailer called for lights, rushed in and fell trembling before Paul and Silas.
ACTS|16|30|He then brought them out and asked, "Sirs, what must I do to be saved?"
ACTS|16|31|They replied, "Believe in the Lord Jesus, and you will be saved--you and your household."
ACTS|16|32|Then they spoke the word of the Lord to him and to all the others in his house.
ACTS|16|33|At that hour of the night the jailer took them and washed their wounds; then immediately he and all his family were baptized.
ACTS|16|34|The jailer brought them into his house and set a meal before them; he was filled with joy because he had come to believe in God--he and his whole family.
ACTS|16|35|When it was daylight, the magistrates sent their officers to the jailer with the order: "Release those men."
ACTS|16|36|The jailer told Paul, "The magistrates have ordered that you and Silas be released. Now you can leave. Go in peace."
ACTS|16|37|But Paul said to the officers: "They beat us publicly without a trial, even though we are Roman citizens, and threw us into prison. And now do they want to get rid of us quietly? No! Let them come themselves and escort us out."
ACTS|16|38|The officers reported this to the magistrates, and when they heard that Paul and Silas were Roman citizens, they were alarmed.
ACTS|16|39|They came to appease them and escorted them from the prison, requesting them to leave the city.
ACTS|16|40|After Paul and Silas came out of the prison, they went to Lydia's house, where they met with the brothers and encouraged them. Then they left.
ACTS|17|1|When they had passed through Amphipolis and Apollonia, they came to Thessalonica, where there was a Jewish synagogue.
ACTS|17|2|As his custom was, Paul went into the synagogue, and on three Sabbath days he reasoned with them from the Scriptures,
ACTS|17|3|explaining and proving that the Christ had to suffer and rise from the dead. "This Jesus I am proclaiming to you is the Christ, "he said.
ACTS|17|4|Some of the Jews were persuaded and joined Paul and Silas, as did a large number of God-fearing Greeks and not a few prominent women.
ACTS|17|5|But the Jews were jealous; so they rounded up some bad characters from the marketplace, formed a mob and started a riot in the city. They rushed to Jason's house in search of Paul and Silas in order to bring them out to the crowd.
ACTS|17|6|But when they did not find them, they dragged Jason and some other brothers before the city officials, shouting: "These men who have caused trouble all over the world have now come here,
ACTS|17|7|and Jason has welcomed them into his house. They are all defying Caesar's decrees, saying that there is another king, one called Jesus."
ACTS|17|8|When they heard this, the crowd and the city officials were thrown into turmoil.
ACTS|17|9|Then they made Jason and the others post bond and let them go.
ACTS|17|10|As soon as it was night, the brothers sent Paul and Silas away to Berea. On arriving there, they went to the Jewish synagogue.
ACTS|17|11|Now the Bereans were of more noble character than the Thessalonians, for they received the message with great eagerness and examined the Scriptures every day to see if what Paul said was true.
ACTS|17|12|Many of the Jews believed, as did also a number of prominent Greek women and many Greek men.
ACTS|17|13|When the Jews in Thessalonica learned that Paul was preaching the word of God at Berea, they went there too, agitating the crowds and stirring them up.
ACTS|17|14|The brothers immediately sent Paul to the coast, but Silas and Timothy stayed at Berea.
ACTS|17|15|The men who escorted Paul brought him to Athens and then left with instructions for Silas and Timothy to join him as soon as possible.
ACTS|17|16|While Paul was waiting for them in Athens, he was greatly distressed to see that the city was full of idols.
ACTS|17|17|So he reasoned in the synagogue with the Jews and the God-fearing Greeks, as well as in the marketplace day by day with those who happened to be there.
ACTS|17|18|A group of Epicurean and Stoic philosophers began to dispute with him. Some of them asked, "What is this babbler trying to say?" Others remarked, "He seems to be advocating foreign gods." They said this because Paul was preaching the good news about Jesus and the resurrection.
ACTS|17|19|Then they took him and brought him to a meeting of the Areopagus, where they said to him, "May we know what this new teaching is that you are presenting?
ACTS|17|20|You are bringing some strange ideas to our ears, and we want to know what they mean."
ACTS|17|21|(All the Athenians and the foreigners who lived there spent their time doing nothing but talking about and listening to the latest ideas.)
ACTS|17|22|Paul then stood up in the meeting of the Areopagus and said: "Men of Athens! I see that in every way you are very religious.
ACTS|17|23|For as I walked around and looked carefully at your objects of worship, I even found an altar with this inscription:|sc TO AN UNKNOWN GOD. Now what you worship as something unknown I am going to proclaim to you.
ACTS|17|24|"The God who made the world and everything in it is the Lord of heaven and earth and does not live in temples built by hands.
ACTS|17|25|And he is not served by human hands, as if he needed anything, because he himself gives all men life and breath and everything else.
ACTS|17|26|From one man he made every nation of men, that they should inhabit the whole earth; and he determined the times set for them and the exact places where they should live.
ACTS|17|27|God did this so that men would seek him and perhaps reach out for him and find him, though he is not far from each one of us.
ACTS|17|28|'For in him we live and move and have our being.' As some of your own poets have said, 'We are his offspring.'
ACTS|17|29|"Therefore since we are God's offspring, we should not think that the divine being is like gold or silver or stone--an image made by man's design and skill.
ACTS|17|30|In the past God overlooked such ignorance, but now he commands all people everywhere to repent.
ACTS|17|31|For he has set a day when he will judge the world with justice by the man he has appointed. He has given proof of this to all men by raising him from the dead."
ACTS|17|32|When they heard about the resurrection of the dead, some of them sneered, but others said, "We want to hear you again on this subject."
ACTS|17|33|At that, Paul left the Council.
ACTS|17|34|A few men became followers of Paul and believed. Among them was Dionysius, a member of the Areopagus, also a woman named Damaris, and a number of others.
ACTS|18|1|After this, Paul left Athens and went to Corinth.
ACTS|18|2|There he met a Jew named Aquila, a native of Pontus, who had recently come from Italy with his wife Priscilla, because Claudius had ordered all the Jews to leave Rome. Paul went to see them,
ACTS|18|3|and because he was a tentmaker as they were, he stayed and worked with them.
ACTS|18|4|Every Sabbath he reasoned in the synagogue, trying to persuade Jews and Greeks.
ACTS|18|5|When Silas and Timothy came from Macedonia, Paul devoted himself exclusively to preaching, testifying to the Jews that Jesus was the Christ.
ACTS|18|6|But when the Jews opposed Paul and became abusive, he shook out his clothes in protest and said to them, "Your blood be on your own heads! I am clear of my responsibility. From now on I will go to the Gentiles."
ACTS|18|7|Then Paul left the synagogue and went next door to the house of Titius Justus, a worshiper of God.
ACTS|18|8|Crispus, the synagogue ruler, and his entire household believed in the Lord; and many of the Corinthians who heard him believed and were baptized.
ACTS|18|9|One night the Lord spoke to Paul in a vision: "Do not be afraid; keep on speaking, do not be silent.
ACTS|18|10|For I am with you, and no one is going to attack and harm you, because I have many people in this city."
ACTS|18|11|So Paul stayed for a year and a half, teaching them the word of God.
ACTS|18|12|While Gallio was proconsul of Achaia, the Jews made a united attack on Paul and brought him into court.
ACTS|18|13|"This man," they charged, "is persuading the people to worship God in ways contrary to the law."
ACTS|18|14|Just as Paul was about to speak, Gallio said to the Jews, "If you Jews were making a complaint about some misdemeanor or serious crime, it would be reasonable for me to listen to you.
ACTS|18|15|But since it involves questions about words and names and your own law--settle the matter yourselves. I will not be a judge of such things."
ACTS|18|16|So he had them ejected from the court.
ACTS|18|17|Then they all turned on Sosthenes the synagogue ruler and beat him in front of the court. But Gallio showed no concern whatever.
ACTS|18|18|Paul stayed on in Corinth for some time. Then he left the brothers and sailed for Syria, accompanied by Priscilla and Aquila. Before he sailed, he had his hair cut off at Cenchrea because of a vow he had taken.
ACTS|18|19|They arrived at Ephesus, where Paul left Priscilla and Aquila. He himself went into the synagogue and reasoned with the Jews.
ACTS|18|20|When they asked him to spend more time with them, he declined.
ACTS|18|21|But as he left, he promised, "I will come back if it is God's will." Then he set sail from Ephesus.
ACTS|18|22|When he landed at Caesarea, he went up and greeted the church and then went down to Antioch.
ACTS|18|23|After spending some time in Antioch, Paul set out from there and traveled from place to place throughout the region of Galatia and Phrygia, strengthening all the disciples.
ACTS|18|24|Meanwhile a Jew named Apollos, a native of Alexandria, came to Ephesus. He was a learned man, with a thorough knowledge of the Scriptures.
ACTS|18|25|He had been instructed in the way of the Lord, and he spoke with great fervor and taught about Jesus accurately, though he knew only the baptism of John.
ACTS|18|26|He began to speak boldly in the synagogue. When Priscilla and Aquila heard him, they invited him to their home and explained to him the way of God more adequately.
ACTS|18|27|When Apollos wanted to go to Achaia, the brothers encouraged him and wrote to the disciples there to welcome him. On arriving, he was a great help to those who by grace had believed.
ACTS|18|28|For he vigorously refuted the Jews in public debate, proving from the Scriptures that Jesus was the Christ.
ACTS|19|1|While Apollos was at Corinth, Paul took the road through the interior and arrived at Ephesus. There he found some disciples
ACTS|19|2|and asked them, "Did you receive the Holy Spirit when you believed?" They answered, "No, we have not even heard that there is a Holy Spirit."
ACTS|19|3|So Paul asked, "Then what baptism did you receive?John's baptism," they replied.
ACTS|19|4|Paul said, "John's baptism was a baptism of repentance. He told the people to believe in the one coming after him, that is, in Jesus."
ACTS|19|5|On hearing this, they were baptized into the name of the Lord Jesus.
ACTS|19|6|When Paul placed his hands on them, the Holy Spirit came on them, and they spoke in tongues and prophesied.
ACTS|19|7|There were about twelve men in all.
ACTS|19|8|Paul entered the synagogue and spoke boldly there for three months, arguing persuasively about the kingdom of God.
ACTS|19|9|But some of them became obstinate; they refused to believe and publicly maligned the Way. So Paul left them. He took the disciples with him and had discussions daily in the lecture hall of Tyrannus.
ACTS|19|10|This went on for two years, so that all the Jews and Greeks who lived in the province of Asia heard the word of the Lord.
ACTS|19|11|God did extraordinary miracles through Paul,
ACTS|19|12|so that even handkerchiefs and aprons that had touched him were taken to the sick, and their illnesses were cured and the evil spirits left them.
ACTS|19|13|Some Jews who went around driving out evil spirits tried to invoke the name of the Lord Jesus over those who were demon-possessed. They would say, "In the name of Jesus, whom Paul preaches, I command you to come out."
ACTS|19|14|Seven sons of Sceva, a Jewish chief priest, were doing this.
ACTS|19|15|One day the evil spirit answered them, "Jesus I know, and I know about Paul, but who are you?"
ACTS|19|16|Then the man who had the evil spirit jumped on them and overpowered them all. He gave them such a beating that they ran out of the house naked and bleeding.
ACTS|19|17|When this became known to the Jews and Greeks living in Ephesus, they were all seized with fear, and the name of the Lord Jesus was held in high honor.
ACTS|19|18|Many of those who believed now came and openly confessed their evil deeds.
ACTS|19|19|A number who had practiced sorcery brought their scrolls together and burned them publicly. When they calculated the value of the scrolls, the total came to fifty thousand drachmas.
ACTS|19|20|In this way the word of the Lord spread widely and grew in power.
ACTS|19|21|After all this had happened, Paul decided to go to Jerusalem, passing through Macedonia and Achaia. "After I have been there," he said, "I must visit Rome also."
ACTS|19|22|He sent two of his helpers, Timothy and Erastus, to Macedonia, while he stayed in the province of Asia a little longer.
ACTS|19|23|About that time there arose a great disturbance about the Way.
ACTS|19|24|A silversmith named Demetrius, who made silver shrines of Artemis, brought in no little business for the craftsmen.
ACTS|19|25|He called them together, along with the workmen in related trades, and said: "Men, you know we receive a good income from this business.
ACTS|19|26|And you see and hear how this fellow Paul has convinced and led astray large numbers of people here in Ephesus and in practically the whole province of Asia. He says that man-made gods are no gods at all.
ACTS|19|27|There is danger not only that our trade will lose its good name, but also that the temple of the great goddess Artemis will be discredited, and the goddess herself, who is worshiped throughout the province of Asia and the world, will be robbed of her divine majesty."
ACTS|19|28|When they heard this, they were furious and began shouting: "Great is Artemis of the Ephesians!"
ACTS|19|29|Soon the whole city was in an uproar. The people seized Gaius and Aristarchus, Paul's traveling companions from Macedonia, and rushed as one man into the theater.
ACTS|19|30|Paul wanted to appear before the crowd, but the disciples would not let him.
ACTS|19|31|Even some of the officials of the province, friends of Paul, sent him a message begging him not to venture into the theater.
ACTS|19|32|The assembly was in confusion: Some were shouting one thing, some another. Most of the people did not even know why they were there.
ACTS|19|33|The Jews pushed Alexander to the front, and some of the crowd shouted instructions to him. He motioned for silence in order to make a defense before the people.
ACTS|19|34|But when they realized he was a Jew, they all shouted in unison for about two hours: "Great is Artemis of the Ephesians!"
ACTS|19|35|The city clerk quieted the crowd and said: "Men of Ephesus, doesn't all the world know that the city of Ephesus is the guardian of the temple of the great Artemis and of her image, which fell from heaven?
ACTS|19|36|Therefore, since these facts are undeniable, you ought to be quiet and not do anything rash.
ACTS|19|37|You have brought these men here, though they have neither robbed temples nor blasphemed our goddess.
ACTS|19|38|If, then, Demetrius and his fellow craftsmen have a grievance against anybody, the courts are open and there are proconsuls. They can press charges.
ACTS|19|39|If there is anything further you want to bring up, it must be settled in a legal assembly.
ACTS|19|40|As it is, we are in danger of being charged with rioting because of today's events. In that case we would not be able to account for this commotion, since there is no reason for it."
ACTS|19|41|After he had said this, he dismissed the assembly.
ACTS|20|1|When the uproar had ended, Paul sent for the disciples and, after encouraging them, said good-by and set out for Macedonia.
ACTS|20|2|He traveled through that area, speaking many words of encouragement to the people, and finally arrived in Greece,
ACTS|20|3|where he stayed three months. Because the Jews made a plot against him just as he was about to sail for Syria, he decided to go back through Macedonia.
ACTS|20|4|He was accompanied by Sopater son of Pyrrhus from Berea, Aristarchus and Secundus from Thessalonica, Gaius from Derbe, Timothy also, and Tychicus and Trophimus from the province of Asia.
ACTS|20|5|These men went on ahead and waited for us at Troas.
ACTS|20|6|But we sailed from Philippi after the Feast of Unleavened Bread, and five days later joined the others at Troas, where we stayed seven days.
ACTS|20|7|On the first day of the week we came together to break bread. Paul spoke to the people and, because he intended to leave the next day, kept on talking until midnight.
ACTS|20|8|There were many lamps in the upstairs room where we were meeting.
ACTS|20|9|Seated in a window was a young man named Eutychus, who was sinking into a deep sleep as Paul talked on and on. When he was sound asleep, he fell to the ground from the third story and was picked up dead.
ACTS|20|10|Paul went down, threw himself on the young man and put his arms around him. "Don't be alarmed," he said. "He's alive!"
ACTS|20|11|Then he went upstairs again and broke bread and ate. After talking until daylight, he left.
ACTS|20|12|The people took the young man home alive and were greatly comforted.
ACTS|20|13|We went on ahead to the ship and sailed for Assos, where we were going to take Paul aboard. He had made this arrangement because he was going there on foot.
ACTS|20|14|When he met us at Assos, we took him aboard and went on to Mitylene.
ACTS|20|15|The next day we set sail from there and arrived off Kios. The day after that we crossed over to Samos, and on the following day arrived at Miletus.
ACTS|20|16|Paul had decided to sail past Ephesus to avoid spending time in the province of Asia, for he was in a hurry to reach Jerusalem, if possible, by the day of Pentecost.
ACTS|20|17|From Miletus, Paul sent to Ephesus for the elders of the church.
ACTS|20|18|When they arrived, he said to them: "You know how I lived the whole time I was with you, from the first day I came into the province of Asia.
ACTS|20|19|I served the Lord with great humility and with tears, although I was severely tested by the plots of the Jews.
ACTS|20|20|You know that I have not hesitated to preach anything that would be helpful to you but have taught you publicly and from house to house.
ACTS|20|21|I have declared to both Jews and Greeks that they must turn to God in repentance and have faith in our Lord Jesus.
ACTS|20|22|"And now, compelled by the Spirit, I am going to Jerusalem, not knowing what will happen to me there.
ACTS|20|23|I only know that in every city the Holy Spirit warns me that prison and hardships are facing me.
ACTS|20|24|However, I consider my life worth nothing to me, if only I may finish the race and complete the task the Lord Jesus has given me--the task of testifying to the gospel of God's grace.
ACTS|20|25|"Now I know that none of you among whom I have gone about preaching the kingdom will ever see me again.
ACTS|20|26|Therefore, I declare to you today that I am innocent of the blood of all men.
ACTS|20|27|For I have not hesitated to proclaim to you the whole will of God.
ACTS|20|28|Keep watch over yourselves and all the flock of which the Holy Spirit has made you overseers. Be shepherds of the church of God, which he bought with his own blood.
ACTS|20|29|I know that after I leave, savage wolves will come in among you and will not spare the flock.
ACTS|20|30|Even from your own number men will arise and distort the truth in order to draw away disciples after them.
ACTS|20|31|So be on your guard! Remember that for three years I never stopped warning each of you night and day with tears.
ACTS|20|32|"Now I commit you to God and to the word of his grace, which can build you up and give you an inheritance among all those who are sanctified.
ACTS|20|33|I have not coveted anyone's silver or gold or clothing.
ACTS|20|34|You yourselves know that these hands of mine have supplied my own needs and the needs of my companions.
ACTS|20|35|In everything I did, I showed you that by this kind of hard work we must help the weak, remembering the words the Lord Jesus himself said: 'It is more blessed to give than to receive.'"
ACTS|20|36|When he had said this, he knelt down with all of them and prayed.
ACTS|20|37|They all wept as they embraced him and kissed him.
ACTS|20|38|What grieved them most was his statement that they would never see his face again. Then they accompanied him to the ship.
ACTS|21|1|After we had torn ourselves away from them, we put out to sea and sailed straight to Cos. The next day we went to Rhodes and from there to Patara.
ACTS|21|2|We found a ship crossing over to Phoenicia, went on board and set sail.
ACTS|21|3|After sighting Cyprus and passing to the south of it, we sailed on to Syria. We landed at Tyre, where our ship was to unload its cargo.
ACTS|21|4|Finding the disciples there, we stayed with them seven days. Through the Spirit they urged Paul not to go on to Jerusalem.
ACTS|21|5|But when our time was up, we left and continued on our way. All the disciples and their wives and children accompanied us out of the city, and there on the beach we knelt to pray.
ACTS|21|6|After saying good-by to each other, we went aboard the ship, and they returned home.
ACTS|21|7|We continued our voyage from Tyre and landed at Ptolemais, where we greeted the brothers and stayed with them for a day.
ACTS|21|8|Leaving the next day, we reached Caesarea and stayed at the house of Philip the evangelist, one of the Seven.
ACTS|21|9|He had four unmarried daughters who prophesied.
ACTS|21|10|After we had been there a number of days, a prophet named Agabus came down from Judea.
ACTS|21|11|Coming over to us, he took Paul's belt, tied his own hands and feet with it and said, "The Holy Spirit says, 'In this way the Jews of Jerusalem will bind the owner of this belt and will hand him over to the Gentiles.'"
ACTS|21|12|When we heard this, we and the people there pleaded with Paul not to go up to Jerusalem.
ACTS|21|13|Then Paul answered, "Why are you weeping and breaking my heart? I am ready not only to be bound, but also to die in Jerusalem for the name of the Lord Jesus."
ACTS|21|14|When he would not be dissuaded, we gave up and said, "The Lord's will be done."
ACTS|21|15|After this, we got ready and went up to Jerusalem.
ACTS|21|16|Some of the disciples from Caesarea accompanied us and brought us to the home of Mnason, where we were to stay. He was a man from Cyprus and one of the early disciples.
ACTS|21|17|When we arrived at Jerusalem, the brothers received us warmly.
ACTS|21|18|The next day Paul and the rest of us went to see James, and all the elders were present.
ACTS|21|19|Paul greeted them and reported in detail what God had done among the Gentiles through his ministry.
ACTS|21|20|When they heard this, they praised God. Then they said to Paul: "You see, brother, how many thousands of Jews have believed, and all of them are zealous for the law.
ACTS|21|21|They have been informed that you teach all the Jews who live among the Gentiles to turn away from Moses, telling them not to circumcise their children or live according to our customs.
ACTS|21|22|What shall we do? They will certainly hear that you have come,
ACTS|21|23|so do what we tell you. There are four men with us who have made a vow.
ACTS|21|24|Take these men, join in their purification rites and pay their expenses, so that they can have their heads shaved. Then everybody will know there is no truth in these reports about you, but that you yourself are living in obedience to the law.
ACTS|21|25|As for the Gentile believers, we have written to them our decision that they should abstain from food sacrificed to idols, from blood, from the meat of strangled animals and from sexual immorality."
ACTS|21|26|The next day Paul took the men and purified himself along with them. Then he went to the temple to give notice of the date when the days of purification would end and the offering would be made for each of them.
ACTS|21|27|When the seven days were nearly over, some Jews from the province of Asia saw Paul at the temple. They stirred up the whole crowd and seized him,
ACTS|21|28|shouting, "Men of Israel, help us! This is the man who teaches all men everywhere against our people and our law and this place. And besides, he has brought Greeks into the temple area and defiled this holy place."
ACTS|21|29|(They had previously seen Trophimus the Ephesian in the city with Paul and assumed that Paul had brought him into the temple area.)
ACTS|21|30|The whole city was aroused, and the people came running from all directions. Seizing Paul, they dragged him from the temple, and immediately the gates were shut.
ACTS|21|31|While they were trying to kill him, news reached the commander of the Roman troops that the whole city of Jerusalem was in an uproar.
ACTS|21|32|He at once took some officers and soldiers and ran down to the crowd. When the rioters saw the commander and his soldiers, they stopped beating Paul.
ACTS|21|33|The commander came up and arrested him and ordered him to be bound with two chains. Then he asked who he was and what he had done.
ACTS|21|34|Some in the crowd shouted one thing and some another, and since the commander could not get at the truth because of the uproar, he ordered that Paul be taken into the barracks.
ACTS|21|35|When Paul reached the steps, the violence of the mob was so great he had to be carried by the soldiers.
ACTS|21|36|The crowd that followed kept shouting, "Away with him!"
ACTS|21|37|As the soldiers were about to take Paul into the barracks, he asked the commander, "May I say something to you?"
ACTS|21|38|"Do you speak Greek?" he replied. "Aren't you the Egyptian who started a revolt and led four thousand terrorists out into the desert some time ago?"
ACTS|21|39|Paul answered, "I am a Jew, from Tarsus in Cilicia, a citizen of no ordinary city. Please let me speak to the people."
ACTS|21|40|Having received the commander's permission, Paul stood on the steps and motioned to the crowd. When they were all silent, he said to them in Aramaic:
ACTS|22|1|"Brothers and fathers, listen now to my defense."
ACTS|22|2|When they heard him speak to them in Aramaic, they became very quiet.
ACTS|22|3|Then Paul said: "I am a Jew, born in Tarsus of Cilicia, but brought up in this city. Under Gamaliel I was thoroughly trained in the law of our fathers and was just as zealous for God as any of you are today.
ACTS|22|4|I persecuted the followers of this Way to their death, arresting both men and women and throwing them into prison,
ACTS|22|5|as also the high priest and all the Council can testify. I even obtained letters from them to their brothers in Damascus, and went there to bring these people as prisoners to Jerusalem to be punished.
ACTS|22|6|"About noon as I came near Damascus, suddenly a bright light from heaven flashed around me.
ACTS|22|7|I fell to the ground and heard a voice say to me, 'Saul! Saul! Why do you persecute me?'
ACTS|22|8|"'Who are you, Lord?' I asked.
ACTS|22|9|"'I am Jesus of Nazareth, whom you are persecuting,' he replied. My companions saw the light, but they did not understand the voice of him who was speaking to me.
ACTS|22|10|"'What shall I do, Lord?' I asked.
ACTS|22|11|"'Get up,' the Lord said, 'and go into Damascus. There you will be told all that you have been assigned to do.' My companions led me by the hand into Damascus, because the brilliance of the light had blinded me.
ACTS|22|12|"A man named Ananias came to see me. He was a devout observer of the law and highly respected by all the Jews living there.
ACTS|22|13|He stood beside me and said, 'Brother Saul, receive your sight!' And at that very moment I was able to see him.
ACTS|22|14|"Then he said: 'The God of our fathers has chosen you to know his will and to see the Righteous One and to hear words from his mouth.
ACTS|22|15|You will be his witness to all men of what you have seen and heard.
ACTS|22|16|And now what are you waiting for? Get up, be baptized and wash your sins away, calling on his name.'
ACTS|22|17|"When I returned to Jerusalem and was praying at the temple, I fell into a trance
ACTS|22|18|and saw the Lord speaking. 'Quick!' he said to me. 'Leave Jerusalem immediately, because they will not accept your testimony about me.'
ACTS|22|19|"'Lord,' I replied, 'these men know that I went from one synagogue to another to imprison and beat those who believe in you.
ACTS|22|20|And when the blood of your martyr Stephen was shed, I stood there giving my approval and guarding the clothes of those who were killing him.'
ACTS|22|21|"Then the Lord said to me, 'Go; I will send you far away to the Gentiles.'"
ACTS|22|22|The crowd listened to Paul until he said this. Then they raised their voices and shouted, "Rid the earth of him! He's not fit to live!"
ACTS|22|23|As they were shouting and throwing off their cloaks and flinging dust into the air,
ACTS|22|24|the commander ordered Paul to be taken into the barracks. He directed that he be flogged and questioned in order to find out why the people were shouting at him like this.
ACTS|22|25|As they stretched him out to flog him, Paul said to the centurion standing there, "Is it legal for you to flog a Roman citizen who hasn't even been found guilty?"
ACTS|22|26|When the centurion heard this, he went to the commander and reported it. "What are you going to do?" he asked. "This man is a Roman citizen."
ACTS|22|27|The commander went to Paul and asked, "Tell me, are you a Roman citizen?Yes, I am," he answered.
ACTS|22|28|Then the commander said, "I had to pay a big price for my citizenship.But I was born a citizen," Paul replied.
ACTS|22|29|Those who were about to question him withdrew immediately. The commander himself was alarmed when he realized that he had put Paul, a Roman citizen, in chains.
ACTS|22|30|The next day, since the commander wanted to find out exactly why Paul was being accused by the Jews, he released him and ordered the chief priests and all the Sanhedrin to assemble. Then he brought Paul and had him stand before them.
ACTS|23|1|Paul looked straight at the Sanhedrin and said, "My brothers, I have fulfilled my duty to God in all good conscience to this day."
ACTS|23|2|At this the high priest Ananias ordered those standing near Paul to strike him on the mouth.
ACTS|23|3|Then Paul said to him, "God will strike you, you whitewashed wall! You sit there to judge me according to the law, yet you yourself violate the law by commanding that I be struck!"
ACTS|23|4|Those who were standing near Paul said, "You dare to insult God's high priest?"
ACTS|23|5|Paul replied, "Brothers, I did not realize that he was the high priest; for it is written: 'Do not speak evil about the ruler of your people.'"
ACTS|23|6|Then Paul, knowing that some of them were Sadducees and the others Pharisees, called out in the Sanhedrin, "My brothers, I am a Pharisee, the son of a Pharisee. I stand on trial because of my hope in the resurrection of the dead."
ACTS|23|7|When he said this, a dispute broke out between the Pharisees and the Sadducees, and the assembly was divided.
ACTS|23|8|(The Sadducees say that there is no resurrection, and that there are neither angels nor spirits, but the Pharisees acknowledge them all.)
ACTS|23|9|There was a great uproar, and some of the teachers of the law who were Pharisees stood up and argued vigorously. "We find nothing wrong with this man," they said. "What if a spirit or an angel has spoken to him?"
ACTS|23|10|The dispute became so violent that the commander was afraid Paul would be torn to pieces by them. He ordered the troops to go down and take him away from them by force and bring him into the barracks.
ACTS|23|11|The following night the Lord stood near Paul and said, "Take courage! As you have testified about me in Jerusalem, so you must also testify in Rome."
ACTS|23|12|The next morning the Jews formed a conspiracy and bound themselves with an oath not to eat or drink until they had killed Paul.
ACTS|23|13|More than forty men were involved in this plot.
ACTS|23|14|They went to the chief priests and elders and said, "We have taken a solemn oath not to eat anything until we have killed Paul.
ACTS|23|15|Now then, you and the Sanhedrin petition the commander to bring him before you on the pretext of wanting more accurate information about his case. We are ready to kill him before he gets here."
ACTS|23|16|But when the son of Paul's sister heard of this plot, he went into the barracks and told Paul.
ACTS|23|17|Then Paul called one of the centurions and said, "Take this young man to the commander; he has something to tell him."
ACTS|23|18|So he took him to the commander. The centurion said, "Paul, the prisoner, sent for me and asked me to bring this young man to you because he has something to tell you."
ACTS|23|19|The commander took the young man by the hand, drew him aside and asked, "What is it you want to tell me?"
ACTS|23|20|He said: "The Jews have agreed to ask you to bring Paul before the Sanhedrin tomorrow on the pretext of wanting more accurate information about him.
ACTS|23|21|Don't give in to them, because more than forty of them are waiting in ambush for him. They have taken an oath not to eat or drink until they have killed him. They are ready now, waiting for your consent to their request."
ACTS|23|22|The commander dismissed the young man and cautioned him, "Don't tell anyone that you have reported this to me."
ACTS|23|23|Then he called two of his centurions and ordered them, "Get ready a detachment of two hundred soldiers, seventy horsemen and two hundred spearmen to go to Caesarea at nine tonight.
ACTS|23|24|Provide mounts for Paul so that he may be taken safely to Governor Felix."
ACTS|23|25|He wrote a letter as follows:
ACTS|23|26|Claudius Lysias, To His Excellency, Governor Felix: Greetings.
ACTS|23|27|This man was seized by the Jews and they were about to kill him, but I came with my troops and rescued him, for I had learned that he is a Roman citizen.
ACTS|23|28|I wanted to know why they were accusing him, so I brought him to their Sanhedrin.
ACTS|23|29|I found that the accusation had to do with questions about their law, but there was no charge against him that deserved death or imprisonment.
ACTS|23|30|When I was informed of a plot to be carried out against the man, I sent him to you at once. I also ordered his accusers to present to you their case against him.
ACTS|23|31|So the soldiers, carrying out their orders, took Paul with them during the night and brought him as far as Antipatris.
ACTS|23|32|The next day they let the cavalry go on with him, while they returned to the barracks.
ACTS|23|33|When the cavalry arrived in Caesarea, they delivered the letter to the governor and handed Paul over to him.
ACTS|23|34|The governor read the letter and asked what province he was from. Learning that he was from Cilicia,
ACTS|23|35|he said, "I will hear your case when your accusers get here." Then he ordered that Paul be kept under guard in Herod's palace.
ACTS|24|1|Five days later the high priest Ananias went down to Caesarea with some of the elders and a lawyer named Tertullus, and they brought their charges against Paul before the governor.
ACTS|24|2|When Paul was called in, Tertullus presented his case before Felix: "We have enjoyed a long period of peace under you, and your foresight has brought about reforms in this nation.
ACTS|24|3|Everywhere and in every way, most excellent Felix, we acknowledge this with profound gratitude.
ACTS|24|4|But in order not to weary you further, I would request that you be kind enough to hear us briefly.
ACTS|24|5|"We have found this man to be a troublemaker, stirring up riots among the Jews all over the world. He is a ringleader of the Nazarene sect
ACTS|24|6|and even tried to desecrate the temple; so we seized him.
ACTS|24|7|See Footnote
ACTS|24|8|By examining him yourself you will be able to learn the truth about all these charges we are bringing against him."
ACTS|24|9|The Jews joined in the accusation, asserting that these things were true.
ACTS|24|10|When the governor motioned for him to speak, Paul replied: "I know that for a number of years you have been a judge over this nation; so I gladly make my defense.
ACTS|24|11|You can easily verify that no more than twelve days ago I went up to Jerusalem to worship.
ACTS|24|12|My accusers did not find me arguing with anyone at the temple, or stirring up a crowd in the synagogues or anywhere else in the city.
ACTS|24|13|And they cannot prove to you the charges they are now making against me.
ACTS|24|14|However, I admit that I worship the God of our fathers as a follower of the Way, which they call a sect. I believe everything that agrees with the Law and that is written in the Prophets,
ACTS|24|15|and I have the same hope in God as these men, that there will be a resurrection of both the righteous and the wicked.
ACTS|24|16|So I strive always to keep my conscience clear before God and man.
ACTS|24|17|"After an absence of several years, I came to Jerusalem to bring my people gifts for the poor and to present offerings.
ACTS|24|18|I was ceremonially clean when they found me in the temple courts doing this. There was no crowd with me, nor was I involved in any disturbance.
ACTS|24|19|But there are some Jews from the province of Asia, who ought to be here before you and bring charges if they have anything against me.
ACTS|24|20|Or these who are here should state what crime they found in me when I stood before the Sanhedrin--
ACTS|24|21|unless it was this one thing I shouted as I stood in their presence: 'It is concerning the resurrection of the dead that I am on trial before you today.'"
ACTS|24|22|Then Felix, who was well acquainted with the Way, adjourned the proceedings. "When Lysias the commander comes," he said, "I will decide your case."
ACTS|24|23|He ordered the centurion to keep Paul under guard but to give him some freedom and permit his friends to take care of his needs.
ACTS|24|24|Several days later Felix came with his wife Drusilla, who was a Jewess. He sent for Paul and listened to him as he spoke about faith in Christ Jesus.
ACTS|24|25|As Paul discoursed on righteousness, self-control and the judgment to come, Felix was afraid and said, "That's enough for now! You may leave. When I find it convenient, I will send for you."
ACTS|24|26|At the same time he was hoping that Paul would offer him a bribe, so he sent for him frequently and talked with him.
ACTS|24|27|When two years had passed, Felix was succeeded by Porcius Festus, but because Felix wanted to grant a favor to the Jews, he left Paul in prison.
ACTS|25|1|Three days after arriving in the province, Festus went up from Caesarea to Jerusalem,
ACTS|25|2|where the chief priests and Jewish leaders appeared before him and presented the charges against Paul.
ACTS|25|3|They urgently requested Festus, as a favor to them, to have Paul transferred to Jerusalem, for they were preparing an ambush to kill him along the way.
ACTS|25|4|Festus answered, "Paul is being held at Caesarea, and I myself am going there soon.
ACTS|25|5|Let some of your leaders come with me and press charges against the man there, if he has done anything wrong."
ACTS|25|6|After spending eight or ten days with them, he went down to Caesarea, and the next day he convened the court and ordered that Paul be brought before him.
ACTS|25|7|When Paul appeared, the Jews who had come down from Jerusalem stood around him, bringing many serious charges against him, which they could not prove.
ACTS|25|8|Then Paul made his defense: "I have done nothing wrong against the law of the Jews or against the temple or against Caesar."
ACTS|25|9|Festus, wishing to do the Jews a favor, said to Paul, "Are you willing to go up to Jerusalem and stand trial before me there on these charges?"
ACTS|25|10|Paul answered: "I am now standing before Caesar's court, where I ought to be tried. I have not done any wrong to the Jews, as you yourself know very well.
ACTS|25|11|If, however, I am guilty of doing anything deserving death, I do not refuse to die. But if the charges brought against me by these Jews are not true, no one has the right to hand me over to them. I appeal to Caesar!"
ACTS|25|12|After Festus had conferred with his council, he declared: "You have appealed to Caesar. To Caesar you will go!"
ACTS|25|13|A few days later King Agrippa and Bernice arrived at Caesarea to pay their respects to Festus.
ACTS|25|14|Since they were spending many days there, Festus discussed Paul's case with the king. He said: "There is a man here whom Felix left as a prisoner.
ACTS|25|15|When I went to Jerusalem, the chief priests and elders of the Jews brought charges against him and asked that he be condemned.
ACTS|25|16|"I told them that it is not the Roman custom to hand over any man before he has faced his accusers and has had an opportunity to defend himself against their charges.
ACTS|25|17|When they came here with me, I did not delay the case, but convened the court the next day and ordered the man to be brought in.
ACTS|25|18|When his accusers got up to speak, they did not charge him with any of the crimes I had expected.
ACTS|25|19|Instead, they had some points of dispute with him about their own religion and about a dead man named Jesus who Paul claimed was alive.
ACTS|25|20|I was at a loss how to investigate such matters; so I asked if he would be willing to go to Jerusalem and stand trial there on these charges.
ACTS|25|21|When Paul made his appeal to be held over for the Emperor's decision, I ordered him held until I could send him to Caesar."
ACTS|25|22|Then Agrippa said to Festus, "I would like to hear this man myself." He replied, "Tomorrow you will hear him."
ACTS|25|23|The next day Agrippa and Bernice came with great pomp and entered the audience room with the high ranking officers and the leading men of the city. At the command of Festus, Paul was brought in.
ACTS|25|24|Festus said: "King Agrippa, and all who are present with us, you see this man! The whole Jewish community has petitioned me about him in Jerusalem and here in Caesarea, shouting that he ought not to live any longer.
ACTS|25|25|I found he had done nothing deserving of death, but because he made his appeal to the Emperor I decided to send him to Rome.
ACTS|25|26|But I have nothing definite to write to His Majesty about him. Therefore I have brought him before all of you, and especially before you, King Agrippa, so that as a result of this investigation I may have something to write.
ACTS|25|27|For I think it is unreasonable to send on a prisoner without specifying the charges against him."
ACTS|26|1|Then Agrippa said to Paul, "You have permission to speak for yourself." So Paul motioned with his hand and began his defense:
ACTS|26|2|"King Agrippa, I consider myself fortunate to stand before you today as I make my defense against all the accusations of the Jews,
ACTS|26|3|and especially so because you are well acquainted with all the Jewish customs and controversies. Therefore, I beg you to listen to me patiently.
ACTS|26|4|"The Jews all know the way I have lived ever since I was a child, from the beginning of my life in my own country, and also in Jerusalem.
ACTS|26|5|They have known me for a long time and can testify, if they are willing, that according to the strictest sect of our religion, I lived as a Pharisee.
ACTS|26|6|And now it is because of my hope in what God has promised our fathers that I am on trial today.
ACTS|26|7|This is the promise our twelve tribes are hoping to see fulfilled as they earnestly serve God day and night. O king, it is because of this hope that the Jews are accusing me.
ACTS|26|8|Why should any of you consider it incredible that God raises the dead?
ACTS|26|9|"I too was convinced that I ought to do all that was possible to oppose the name of Jesus of Nazareth.
ACTS|26|10|And that is just what I did in Jerusalem. On the authority of the chief priests I put many of the saints in prison, and when they were put to death, I cast my vote against them.
ACTS|26|11|Many a time I went from one synagogue to another to have them punished, and I tried to force them to blaspheme. In my obsession against them, I even went to foreign cities to persecute them.
ACTS|26|12|"On one of these journeys I was going to Damascus with the authority and commission of the chief priests.
ACTS|26|13|About noon, O king, as I was on the road, I saw a light from heaven, brighter than the sun, blazing around me and my companions.
ACTS|26|14|We all fell to the ground, and I heard a voice saying to me in Aramaic, 'Saul, Saul, why do you persecute me? It is hard for you to kick against the goads.'
ACTS|26|15|"Then I asked, 'Who are you, Lord?'
ACTS|26|16|"'I am Jesus, whom you are persecuting,' the Lord replied. 'Now get up and stand on your feet. I have appeared to you to appoint you as a servant and as a witness of what you have seen of me and what I will show you.
ACTS|26|17|I will rescue you from your own people and from the Gentiles. I am sending you to them
ACTS|26|18|to open their eyes and turn them from darkness to light, and from the power of Satan to God, so that they may receive forgiveness of sins and a place among those who are sanctified by faith in me.'
ACTS|26|19|"So then, King Agrippa, I was not disobedient to the vision from heaven.
ACTS|26|20|First to those in Damascus, then to those in Jerusalem and in all Judea, and to the Gentiles also, I preached that they should repent and turn to God and prove their repentance by their deeds.
ACTS|26|21|That is why the Jews seized me in the temple courts and tried to kill me.
ACTS|26|22|But I have had God's help to this very day, and so I stand here and testify to small and great alike. I am saying nothing beyond what the prophets and Moses said would happen--
ACTS|26|23|that the Christ would suffer and, as the first to rise from the dead, would proclaim light to his own people and to the Gentiles."
ACTS|26|24|At this point Festus interrupted Paul's defense. "You are out of your mind, Paul!" he shouted. "Your great learning is driving you insane."
ACTS|26|25|"I am not insane, most excellent Festus," Paul replied. "What I am saying is true and reasonable.
ACTS|26|26|The king is familiar with these things, and I can speak freely to him. I am convinced that none of this has escaped his notice, because it was not done in a corner.
ACTS|26|27|King Agrippa, do you believe the prophets? I know you do."
ACTS|26|28|Then Agrippa said to Paul, "Do you think that in such a short time you can persuade me to be a Christian?"
ACTS|26|29|Paul replied, "Short time or long--I pray God that not only you but all who are listening to me today may become what I am, except for these chains."
ACTS|26|30|The king rose, and with him the governor and Bernice and those sitting with them.
ACTS|26|31|They left the room, and while talking with one another, they said, "This man is not doing anything that deserves death or imprisonment."
ACTS|26|32|Agrippa said to Festus, "This man could have been set free if he had not appealed to Caesar."
ACTS|27|1|When it was decided that we would sail for Italy, Paul and some other prisoners were handed over to a centurion named Julius, who belonged to the Imperial Regiment.
ACTS|27|2|We boarded a ship from Adramyttium about to sail for ports along the coast of the province of Asia, and we put out to sea. Aristarchus, a Macedonian from Thessalonica, was with us.
ACTS|27|3|The next day we landed at Sidon; and Julius, in kindness to Paul, allowed him to go to his friends so they might provide for his needs.
ACTS|27|4|From there we put out to sea again and passed to the lee of Cyprus because the winds were against us.
ACTS|27|5|When we had sailed across the open sea off the coast of Cilicia and Pamphylia, we landed at Myra in Lycia.
ACTS|27|6|There the centurion found an Alexandrian ship sailing for Italy and put us on board.
ACTS|27|7|We made slow headway for many days and had difficulty arriving off Cnidus. When the wind did not allow us to hold our course, we sailed to the lee of Crete, opposite Salmone.
ACTS|27|8|We moved along the coast with difficulty and came to a place called Fair Havens, near the town of Lasea.
ACTS|27|9|Much time had been lost, and sailing had already become dangerous because by now it was after the Fast. So Paul warned them,
ACTS|27|10|"Men, I can see that our voyage is going to be disastrous and bring great loss to ship and cargo, and to our own lives also."
ACTS|27|11|But the centurion, instead of listening to what Paul said, followed the advice of the pilot and of the owner of the ship.
ACTS|27|12|Since the harbor was unsuitable to winter in, the majority decided that we should sail on, hoping to reach Phoenix and winter there. This was a harbor in Crete, facing both southwest and northwest.
ACTS|27|13|When a gentle south wind began to blow, they thought they had obtained what they wanted; so they weighed anchor and sailed along the shore of Crete.
ACTS|27|14|Before very long, a wind of hurricane force, called the "northeaster," swept down from the island.
ACTS|27|15|The ship was caught by the storm and could not head into the wind; so we gave way to it and were driven along.
ACTS|27|16|As we passed to the lee of a small island called Cauda, we were hardly able to make the lifeboat secure.
ACTS|27|17|When the men had hoisted it aboard, they passed ropes under the ship itself to hold it together. Fearing that they would run aground on the sandbars of Syrtis, they lowered the sea anchor and let the ship be driven along.
ACTS|27|18|We took such a violent battering from the storm that the next day they began to throw the cargo overboard.
ACTS|27|19|On the third day, they threw the ship's tackle overboard with their own hands.
ACTS|27|20|When neither sun nor stars appeared for many days and the storm continued raging, we finally gave up all hope of being saved.
ACTS|27|21|After the men had gone a long time without food, Paul stood up before them and said: "Men, you should have taken my advice not to sail from Crete; then you would have spared yourselves this damage and loss.
ACTS|27|22|But now I urge you to keep up your courage, because not one of you will be lost; only the ship will be destroyed.
ACTS|27|23|Last night an angel of the God whose I am and whom I serve stood beside me
ACTS|27|24|and said, 'Do not be afraid, Paul. You must stand trial before Caesar; and God has graciously given you the lives of all who sail with you.'
ACTS|27|25|So keep up your courage, men, for I have faith in God that it will happen just as he told me.
ACTS|27|26|Nevertheless, we must run aground on some island."
ACTS|27|27|On the fourteenth night we were still being driven across the Adriatic Sea, when about midnight the sailors sensed they were approaching land.
ACTS|27|28|They took soundings and found that the water was a hundred and twenty feet deep. A short time later they took soundings again and found it was ninety feet deep.
ACTS|27|29|Fearing that we would be dashed against the rocks, they dropped four anchors from the stern and prayed for daylight.
ACTS|27|30|In an attempt to escape from the ship, the sailors let the lifeboat down into the sea, pretending they were going to lower some anchors from the bow.
ACTS|27|31|Then Paul said to the centurion and the soldiers, "Unless these men stay with the ship, you cannot be saved."
ACTS|27|32|So the soldiers cut the ropes that held the lifeboat and let it fall away.
ACTS|27|33|Just before dawn Paul urged them all to eat. "For the last fourteen days," he said, "you have been in constant suspense and have gone without food--you haven't eaten anything.
ACTS|27|34|Now I urge you to take some food. You need it to survive. Not one of you will lose a single hair from his head."
ACTS|27|35|After he said this, he took some bread and gave thanks to God in front of them all. Then he broke it and began to eat.
ACTS|27|36|They were all encouraged and ate some food themselves.
ACTS|27|37|Altogether there were 276 of us on board.
ACTS|27|38|When they had eaten as much as they wanted, they lightened the ship by throwing the grain into the sea.
ACTS|27|39|When daylight came, they did not recognize the land, but they saw a bay with a sandy beach, where they decided to run the ship aground if they could.
ACTS|27|40|Cutting loose the anchors, they left them in the sea and at the same time untied the ropes that held the rudders. Then they hoisted the foresail to the wind and made for the beach.
ACTS|27|41|But the ship struck a sandbar and ran aground. The bow stuck fast and would not move, and the stern was broken to pieces by the pounding of the surf.
ACTS|27|42|The soldiers planned to kill the prisoners to prevent any of them from swimming away and escaping.
ACTS|27|43|But the centurion wanted to spare Paul's life and kept them from carrying out their plan. He ordered those who could swim to jump overboard first and get to land.
ACTS|27|44|The rest were to get there on planks or on pieces of the ship. In this way everyone reached land in safety.
ACTS|28|1|Once safely on shore, we found out that the island was called Malta.
ACTS|28|2|The islanders showed us unusual kindness. They built a fire and welcomed us all because it was raining and cold.
ACTS|28|3|Paul gathered a pile of brushwood and, as he put it on the fire, a viper, driven out by the heat, fastened itself on his hand.
ACTS|28|4|When the islanders saw the snake hanging from his hand, they said to each other, "This man must be a murderer; for though he escaped from the sea, Justice has not allowed him to live."
ACTS|28|5|But Paul shook the snake off into the fire and suffered no ill effects.
ACTS|28|6|The people expected him to swell up or suddenly fall dead, but after waiting a long time and seeing nothing unusual happen to him, they changed their minds and said he was a god.
ACTS|28|7|There was an estate nearby that belonged to Publius, the chief official of the island. He welcomed us to his home and for three days entertained us hospitably.
ACTS|28|8|His father was sick in bed, suffering from fever and dysentery. Paul went in to see him and, after prayer, placed his hands on him and healed him.
ACTS|28|9|When this had happened, the rest of the sick on the island came and were cured.
ACTS|28|10|They honored us in many ways and when we were ready to sail, they furnished us with the supplies we needed.
ACTS|28|11|After three months we put out to sea in a ship that had wintered in the island. It was an Alexandrian ship with the figurehead of the twin gods Castor and Pollux.
ACTS|28|12|We put in at Syracuse and stayed there three days.
ACTS|28|13|From there we set sail and arrived at Rhegium. The next day the south wind came up, and on the following day we reached Puteoli.
ACTS|28|14|There we found some brothers who invited us to spend a week with them. And so we came to Rome.
ACTS|28|15|The brothers there had heard that we were coming, and they traveled as far as the Forum of Appius and the Three Taverns to meet us. At the sight of these men Paul thanked God and was encouraged.
ACTS|28|16|When we got to Rome, Paul was allowed to live by himself, with a soldier to guard him.
ACTS|28|17|Three days later he called together the leaders of the Jews. When they had assembled, Paul said to them: "My brothers, although I have done nothing against our people or against the customs of our ancestors, I was arrested in Jerusalem and handed over to the Romans.
ACTS|28|18|They examined me and wanted to release me, because I was not guilty of any crime deserving death.
ACTS|28|19|But when the Jews objected, I was compelled to appeal to Caesar--not that I had any charge to bring against my own people.
ACTS|28|20|For this reason I have asked to see you and talk with you. It is because of the hope of Israel that I am bound with this chain."
ACTS|28|21|They replied, "We have not received any letters from Judea concerning you, and none of the brothers who have come from there has reported or said anything bad about you.
ACTS|28|22|But we want to hear what your views are, for we know that people everywhere are talking against this sect."
ACTS|28|23|They arranged to meet Paul on a certain day, and came in even larger numbers to the place where he was staying. From morning till evening he explained and declared to them the kingdom of God and tried to convince them about Jesus from the Law of Moses and from the Prophets.
ACTS|28|24|Some were convinced by what he said, but others would not believe.
ACTS|28|25|They disagreed among themselves and began to leave after Paul had made this final statement: "The Holy Spirit spoke the truth to your forefathers when he said through Isaiah the prophet:
ACTS|28|26|"'Go to this people and say, "You will be ever hearing but never understanding; you will be ever seeing but never perceiving."
ACTS|28|27|For this people's heart has become calloused; they hardly hear with their ears, and they have closed their eyes. Otherwise they might see with their eyes, hear with their ears, understand with their hearts and turn, and I would heal them.'
ACTS|28|28|"Therefore I want you to know that God's salvation has been sent to the Gentiles, and they will listen!"
ACTS|28|29|See Footnote
ACTS|28|30|For two whole years Paul stayed there in his own rented house and welcomed all who came to see him.
ACTS|28|31|Boldly and without hindrance he preached the kingdom of God and taught about the Lord Jesus Christ.
