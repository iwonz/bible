GEN|1|1|In the beginning God created the heavens and the earth.
GEN|1|2|Now the earth was formless and empty, darkness was over the surface of the deep, and the Spirit of God was hovering over the waters.
GEN|1|3|And God said, "Let there be light," and there was light.
GEN|1|4|God saw that the light was good, and he separated the light from the darkness.
GEN|1|5|God called the light "day," and the darkness he called "night." And there was evening, and there was morning-the first day.
GEN|1|6|And God said, "Let there be an expanse between the waters to separate water from water."
GEN|1|7|So God made the expanse and separated the water under the expanse from the water above it. And it was so.
GEN|1|8|God called the expanse "sky." And there was evening, and there was morning-the second day.
GEN|1|9|And God said, "Let the water under the sky be gathered to one place, and let dry ground appear." And it was so.
GEN|1|10|God called the dry ground "land," and the gathered waters he called "seas." And God saw that it was good.
GEN|1|11|Then God said, "Let the land produce vegetation: seed-bearing plants and trees on the land that bear fruit with seed in it, according to their various kinds." And it was so.
GEN|1|12|The land produced vegetation: plants bearing seed according to their kinds and trees bearing fruit with seed in it according to their kinds. And God saw that it was good.
GEN|1|13|And there was evening, and there was morning-the third day.
GEN|1|14|And God said, "Let there be lights in the expanse of the sky to separate the day from the night, and let them serve as signs to mark seasons and days and years,
GEN|1|15|and let them be lights in the expanse of the sky to give light on the earth." And it was so.
GEN|1|16|God made two great lights-the greater light to govern the day and the lesser light to govern the night. He also made the stars.
GEN|1|17|God set them in the expanse of the sky to give light on the earth,
GEN|1|18|to govern the day and the night, and to separate light from darkness. And God saw that it was good.
GEN|1|19|And there was evening, and there was morning-the fourth day.
GEN|1|20|And God said, "Let the water teem with living creatures, and let birds fly above the earth across the expanse of the sky."
GEN|1|21|So God created the great creatures of the sea and every living and moving thing with which the water teems, according to their kinds, and every winged bird according to its kind. And God saw that it was good.
GEN|1|22|God blessed them and said, "Be fruitful and increase in number and fill the water in the seas, and let the birds increase on the earth."
GEN|1|23|And there was evening, and there was morning-the fifth day.
GEN|1|24|And God said, "Let the land produce living creatures according to their kinds: livestock, creatures that move along the ground, and wild animals, each according to its kind." And it was so.
GEN|1|25|God made the wild animals according to their kinds, the livestock according to their kinds, and all the creatures that move along the ground according to their kinds. And God saw that it was good.
GEN|1|26|Then God said, "Let us make man in our image, in our likeness, and let them rule over the fish of the sea and the birds of the air, over the livestock, over all the earth, and over all the creatures that move along the ground."
GEN|1|27|So God created man in his own image, in the image of God he created him; male and female he created them.
GEN|1|28|God blessed them and said to them, "Be fruitful and increase in number; fill the earth and subdue it. Rule over the fish of the sea and the birds of the air and over every living creature that moves on the ground."
GEN|1|29|Then God said, "I give you every seed-bearing plant on the face of the whole earth and every tree that has fruit with seed in it. They will be yours for food.
GEN|1|30|And to all the beasts of the earth and all the birds of the air and all the creatures that move on the ground-everything that has the breath of life in it-I give every green plant for food." And it was so.
GEN|1|31|God saw all that he had made, and it was very good. And there was evening, and there was morning-the sixth day.
GEN|2|1|Thus the heavens and the earth were completed in all their vast array.
GEN|2|2|By the seventh day God had finished the work he had been doing; so on the seventh day he rested from all his work.
GEN|2|3|And God blessed the seventh day and made it holy, because on it he rested from all the work of creating that he had done.
GEN|2|4|This is the account of the heavens and the earth when they were created. When the LORD God made the earth and the heavens-
GEN|2|5|and no shrub of the field had yet appeared on the earth and no plant of the field had yet sprung up, for the LORD God had not sent rain on the earth and there was no man to work the ground,
GEN|2|6|but streams came up from the earth and watered the whole surface of the ground-
GEN|2|7|the LORD God formed the man from the dust of the ground and breathed into his nostrils the breath of life, and the man became a living being.
GEN|2|8|Now the LORD God had planted a garden in the east, in Eden; and there he put the man he had formed.
GEN|2|9|And the LORD God made all kinds of trees grow out of the ground-trees that were pleasing to the eye and good for food. In the middle of the garden were the tree of life and the tree of the knowledge of good and evil.
GEN|2|10|A river watering the garden flowed from Eden; from there it was separated into four headwaters.
GEN|2|11|The name of the first is the Pishon; it winds through the entire land of Havilah, where there is gold.
GEN|2|12|(The gold of that land is good; aromatic resin and onyx are also there.)
GEN|2|13|The name of the second river is the Gihon; it winds through the entire land of Cush.
GEN|2|14|The name of the third river is the Tigris; it runs along the east side of Asshur. And the fourth river is the Euphrates.
GEN|2|15|The LORD God took the man and put him in the Garden of Eden to work it and take care of it.
GEN|2|16|And the LORD God commanded the man, "You are free to eat from any tree in the garden;
GEN|2|17|but you must not eat from the tree of the knowledge of good and evil, for when you eat of it you will surely die."
GEN|2|18|The LORD God said, "It is not good for the man to be alone. I will make a helper suitable for him."
GEN|2|19|Now the LORD God had formed out of the ground all the beasts of the field and all the birds of the air. He brought them to the man to see what he would name them; and whatever the man called each living creature, that was its name.
GEN|2|20|So the man gave names to all the livestock, the birds of the air and all the beasts of the field. But for Adam no suitable helper was found.
GEN|2|21|So the LORD God caused the man to fall into a deep sleep; and while he was sleeping, he took one of the man's ribs and closed up the place with flesh.
GEN|2|22|Then the LORD God made a woman from the rib he had taken out of the man, and he brought her to the man.
GEN|2|23|The man said, "This is now bone of my bones and flesh of my flesh; she shall be called 'woman, 'for she was taken out of man."
GEN|2|24|For this reason a man will leave his father and mother and be united to his wife, and they will become one flesh.
GEN|2|25|The man and his wife were both naked, and they felt no shame.
GEN|3|1|Now the serpent was more crafty than any of the wild animals the LORD God had made. He said to the woman, "Did God really say, 'You must not eat from any tree in the garden'?"
GEN|3|2|The woman said to the serpent, "We may eat fruit from the trees in the garden,
GEN|3|3|but God did say, 'You must not eat fruit from the tree that is in the middle of the garden, and you must not touch it, or you will die.'"
GEN|3|4|"You will not surely die," the serpent said to the woman.
GEN|3|5|"For God knows that when you eat of it your eyes will be opened, and you will be like God, knowing good and evil."
GEN|3|6|When the woman saw that the fruit of the tree was good for food and pleasing to the eye, and also desirable for gaining wisdom, she took some and ate it. She also gave some to her husband, who was with her, and he ate it.
GEN|3|7|Then the eyes of both of them were opened, and they realized they were naked; so they sewed fig leaves together and made coverings for themselves.
GEN|3|8|Then the man and his wife heard the sound of the LORD God as he was walking in the garden in the cool of the day, and they hid from the LORD God among the trees of the garden.
GEN|3|9|But the LORD God called to the man, "Where are you?"
GEN|3|10|He answered, "I heard you in the garden, and I was afraid because I was naked; so I hid."
GEN|3|11|And he said, "Who told you that you were naked? Have you eaten from the tree that I commanded you not to eat from?"
GEN|3|12|The man said, "The woman you put here with me-she gave me some fruit from the tree, and I ate it."
GEN|3|13|Then the LORD God said to the woman, "What is this you have done?" The woman said, "The serpent deceived me, and I ate."
GEN|3|14|So the LORD God said to the serpent, "Because you have done this, "Cursed are you above all the livestock and all the wild animals! You will crawl on your belly and you will eat dust all the days of your life.
GEN|3|15|And I will put enmity between you and the woman, and between your offspring and hers; he will crush your head, and you will strike his heel."
GEN|3|16|To the woman he said, "I will greatly increase your pains in childbearing; with pain you will give birth to children. Your desire will be for your husband, and he will rule over you."
GEN|3|17|To Adam he said, "Because you listened to your wife and ate from the tree about which I commanded you, 'You must not eat of it,'"Cursed is the ground because of you; through painful toil you will eat of it all the days of your life.
GEN|3|18|It will produce thorns and thistles for you, and you will eat the plants of the field.
GEN|3|19|By the sweat of your brow you will eat your food until you return to the ground, since from it you were taken; for dust you are and to dust you will return."
GEN|3|20|Adam named his wife Eve, because she would become the mother of all the living.
GEN|3|21|The LORD God made garments of skin for Adam and his wife and clothed them.
GEN|3|22|And the LORD God said, "The man has now become like one of us, knowing good and evil. He must not be allowed to reach out his hand and take also from the tree of life and eat, and live forever."
GEN|3|23|So the LORD God banished him from the Garden of Eden to work the ground from which he had been taken.
GEN|3|24|After he drove the man out, he placed on the east side of the Garden of Eden cherubim and a flaming sword flashing back and forth to guard the way to the tree of life.
GEN|4|1|Adam lay with his wife Eve, and she became pregnant and gave birth to Cain. She said, "With the help of the LORD I have brought forth a man."
GEN|4|2|Later she gave birth to his brother Abel. Now Abel kept flocks, and Cain worked the soil.
GEN|4|3|In the course of time Cain brought some of the fruits of the soil as an offering to the LORD.
GEN|4|4|But Abel brought fat portions from some of the firstborn of his flock. The LORD looked with favor on Abel and his offering,
GEN|4|5|but on Cain and his offering he did not look with favor. So Cain was very angry, and his face was downcast.
GEN|4|6|Then the LORD said to Cain, "Why are you angry? Why is your face downcast?
GEN|4|7|If you do what is right, will you not be accepted? But if you do not do what is right, sin is crouching at your door; it desires to have you, but you must master it."
GEN|4|8|Now Cain said to his brother Abel, "Let's go out to the field." And while they were in the field, Cain attacked his brother Abel and killed him.
GEN|4|9|Then the LORD said to Cain, "Where is your brother Abel?I don't know," he replied. "Am I my brother's keeper?"
GEN|4|10|The LORD said, "What have you done? Listen! Your brother's blood cries out to me from the ground.
GEN|4|11|Now you are under a curse and driven from the ground, which opened its mouth to receive your brother's blood from your hand.
GEN|4|12|When you work the ground, it will no longer yield its crops for you. You will be a restless wanderer on the earth."
GEN|4|13|Cain said to the LORD, "My punishment is more than I can bear.
GEN|4|14|Today you are driving me from the land, and I will be hidden from your presence; I will be a restless wanderer on the earth, and whoever finds me will kill me."
GEN|4|15|But the LORD said to him, "Not so; if anyone kills Cain, he will suffer vengeance seven times over." Then the LORD put a mark on Cain so that no one who found him would kill him.
GEN|4|16|So Cain went out from the LORD's presence and lived in the land of Nod, east of Eden.
GEN|4|17|Cain lay with his wife, and she became pregnant and gave birth to Enoch. Cain was then building a city, and he named it after his son Enoch.
GEN|4|18|To Enoch was born Irad, and Irad was the father of Mehujael, and Mehujael was the father of Methushael, and Methushael was the father of Lamech.
GEN|4|19|Lamech married two women, one named Adah and the other Zillah.
GEN|4|20|Adah gave birth to Jabal; he was the father of those who live in tents and raise livestock.
GEN|4|21|His brother's name was Jubal; he was the father of all who play the harp and flute.
GEN|4|22|Zillah also had a son, Tubal-Cain, who forged all kinds of tools out of bronze and iron. Tubal-Cain's sister was Naamah.
GEN|4|23|Lamech said to his wives, "Adah and Zillah, listen to me; wives of Lamech, hear my words. I have killed a man for wounding me, a young man for injuring me.
GEN|4|24|If Cain is avenged seven times, then Lamech seventy-seven times."
GEN|4|25|Adam lay with his wife again, and she gave birth to a son and named him Seth, saying, "God has granted me another child in place of Abel, since Cain killed him."
GEN|4|26|Seth also had a son, and he named him Enosh. At that time men began to call on the name of the LORD.
GEN|5|1|This is the written account of Adam's line. When God created man, he made him in the likeness of God.
GEN|5|2|He created them male and female and blessed them. And when they were created, he called them "man. "
GEN|5|3|When Adam had lived 130 years, he had a son in his own likeness, in his own image; and he named him Seth.
GEN|5|4|After Seth was born, Adam lived 800 years and had other sons and daughters.
GEN|5|5|Altogether, Adam lived 930 years, and then he died.
GEN|5|6|When Seth had lived 105 years, he became the father of Enosh.
GEN|5|7|And after he became the father of Enosh, Seth lived 807 years and had other sons and daughters.
GEN|5|8|Altogether, Seth lived 912 years, and then he died.
GEN|5|9|When Enosh had lived 90 years, he became the father of Kenan.
GEN|5|10|And after he became the father of Kenan, Enosh lived 815 years and had other sons and daughters.
GEN|5|11|Altogether, Enosh lived 905 years, and then he died.
GEN|5|12|When Kenan had lived 70 years, he became the father of Mahalalel.
GEN|5|13|And after he became the father of Mahalalel, Kenan lived 840 years and had other sons and daughters.
GEN|5|14|Altogether, Kenan lived 910 years, and then he died.
GEN|5|15|When Mahalalel had lived 65 years, he became the father of Jared.
GEN|5|16|And after he became the father of Jared, Mahalalel lived 830 years and had other sons and daughters.
GEN|5|17|Altogether, Mahalalel lived 895 years, and then he died.
GEN|5|18|When Jared had lived 162 years, he became the father of Enoch.
GEN|5|19|And after he became the father of Enoch, Jared lived 800 years and had other sons and daughters.
GEN|5|20|Altogether, Jared lived 962 years, and then he died.
GEN|5|21|When Enoch had lived 65 years, he became the father of Methuselah.
GEN|5|22|And after he became the father of Methuselah, Enoch walked with God 300 years and had other sons and daughters.
GEN|5|23|Altogether, Enoch lived 365 years.
GEN|5|24|Enoch walked with God; then he was no more, because God took him away.
GEN|5|25|When Methuselah had lived 187 years, he became the father of Lamech.
GEN|5|26|And after he became the father of Lamech, Methuselah lived 782 years and had other sons and daughters.
GEN|5|27|Altogether, Methuselah lived 969 years, and then he died.
GEN|5|28|When Lamech had lived 182 years, he had a son.
GEN|5|29|He named him Noah and said, "He will comfort us in the labor and painful toil of our hands caused by the ground the LORD has cursed."
GEN|5|30|After Noah was born, Lamech lived 595 years and had other sons and daughters.
GEN|5|31|Altogether, Lamech lived 777 years, and then he died.
GEN|5|32|After Noah was 500 years old, he became the father of Shem, Ham and Japheth.
GEN|6|1|When men began to increase in number on the earth and daughters were born to them,
GEN|6|2|the sons of God saw that the daughters of men were beautiful, and they married any of them they chose.
GEN|6|3|Then the LORD said, "My Spirit will not contend with man forever, for he is mortal; his days will be a hundred and twenty years."
GEN|6|4|The Nephilim were on the earth in those days-and also afterward-when the sons of God went to the daughters of men and had children by them. They were the heroes of old, men of renown.
GEN|6|5|The LORD saw how great man's wickedness on the earth had become, and that every inclination of the thoughts of his heart was only evil all the time.
GEN|6|6|The LORD was grieved that he had made man on the earth, and his heart was filled with pain.
GEN|6|7|So the LORD said, "I will wipe mankind, whom I have created, from the face of the earth-men and animals, and creatures that move along the ground, and birds of the air-for I am grieved that I have made them."
GEN|6|8|But Noah found favor in the eyes of the LORD.
GEN|6|9|This is the account of Noah. Noah was a righteous man, blameless among the people of his time, and he walked with God.
GEN|6|10|Noah had three sons: Shem, Ham and Japheth.
GEN|6|11|Now the earth was corrupt in God's sight and was full of violence.
GEN|6|12|God saw how corrupt the earth had become, for all the people on earth had corrupted their ways.
GEN|6|13|So God said to Noah, "I am going to put an end to all people, for the earth is filled with violence because of them. I am surely going to destroy both them and the earth.
GEN|6|14|So make yourself an ark of cypress wood; make rooms in it and coat it with pitch inside and out.
GEN|6|15|This is how you are to build it: The ark is to be 450 feet long, 75 feet wide and 45 feet high.
GEN|6|16|Make a roof for it and finish the ark to within 18 inches of the top. Put a door in the side of the ark and make lower, middle and upper decks.
GEN|6|17|I am going to bring floodwaters on the earth to destroy all life under the heavens, every creature that has the breath of life in it. Everything on earth will perish.
GEN|6|18|But I will establish my covenant with you, and you will enter the ark-you and your sons and your wife and your sons' wives with you.
GEN|6|19|You are to bring into the ark two of all living creatures, male and female, to keep them alive with you.
GEN|6|20|Two of every kind of bird, of every kind of animal and of every kind of creature that moves along the ground will come to you to be kept alive.
GEN|6|21|You are to take every kind of food that is to be eaten and store it away as food for you and for them."
GEN|6|22|Noah did everything just as God commanded him.
GEN|7|1|The LORD then said to Noah, "Go into the ark, you and your whole family, because I have found you righteous in this generation.
GEN|7|2|Take with you seven of every kind of clean animal, a male and its mate, and two of every kind of unclean animal, a male and its mate,
GEN|7|3|and also seven of every kind of bird, male and female, to keep their various kinds alive throughout the earth.
GEN|7|4|Seven days from now I will send rain on the earth for forty days and forty nights, and I will wipe from the face of the earth every living creature I have made."
GEN|7|5|And Noah did all that the LORD commanded him.
GEN|7|6|Noah was six hundred years old when the floodwaters came on the earth.
GEN|7|7|And Noah and his sons and his wife and his sons' wives entered the ark to escape the waters of the flood.
GEN|7|8|Pairs of clean and unclean animals, of birds and of all creatures that move along the ground,
GEN|7|9|male and female, came to Noah and entered the ark, as God had commanded Noah.
GEN|7|10|And after the seven days the floodwaters came on the earth.
GEN|7|11|In the six hundredth year of Noah's life, on the seventeenth day of the second month-on that day all the springs of the great deep burst forth, and the floodgates of the heavens were opened.
GEN|7|12|And rain fell on the earth forty days and forty nights.
GEN|7|13|On that very day Noah and his sons, Shem, Ham and Japheth, together with his wife and the wives of his three sons, entered the ark.
GEN|7|14|They had with them every wild animal according to its kind, all livestock according to their kinds, every creature that moves along the ground according to its kind and every bird according to its kind, everything with wings.
GEN|7|15|Pairs of all creatures that have the breath of life in them came to Noah and entered the ark.
GEN|7|16|The animals going in were male and female of every living thing, as God had commanded Noah. Then the LORD shut him in.
GEN|7|17|For forty days the flood kept coming on the earth, and as the waters increased they lifted the ark high above the earth.
GEN|7|18|The waters rose and increased greatly on the earth, and the ark floated on the surface of the water.
GEN|7|19|They rose greatly on the earth, and all the high mountains under the entire heavens were covered.
GEN|7|20|The waters rose and covered the mountains to a depth of more than twenty feet.,
GEN|7|21|Every living thing that moved on the earth perished-birds, livestock, wild animals, all the creatures that swarm over the earth, and all mankind.
GEN|7|22|Everything on dry land that had the breath of life in its nostrils died.
GEN|7|23|Every living thing on the face of the earth was wiped out; men and animals and the creatures that move along the ground and the birds of the air were wiped from the earth. Only Noah was left, and those with him in the ark.
GEN|7|24|The waters flooded the earth for a hundred and fifty days.
GEN|8|1|But God remembered Noah and all the wild animals and the livestock that were with him in the ark, and he sent a wind over the earth, and the waters receded.
GEN|8|2|Now the springs of the deep and the floodgates of the heavens had been closed, and the rain had stopped falling from the sky.
GEN|8|3|The water receded steadily from the earth. At the end of the hundred and fifty days the water had gone down,
GEN|8|4|and on the seventeenth day of the seventh month the ark came to rest on the mountains of Ararat.
GEN|8|5|The waters continued to recede until the tenth month, and on the first day of the tenth month the tops of the mountains became visible.
GEN|8|6|After forty days Noah opened the window he had made in the ark
GEN|8|7|and sent out a raven, and it kept flying back and forth until the water had dried up from the earth.
GEN|8|8|Then he sent out a dove to see if the water had receded from the surface of the ground.
GEN|8|9|But the dove could find no place to set its feet because there was water over all the surface of the earth; so it returned to Noah in the ark. He reached out his hand and took the dove and brought it back to himself in the ark.
GEN|8|10|He waited seven more days and again sent out the dove from the ark.
GEN|8|11|When the dove returned to him in the evening, there in its beak was a freshly plucked olive leaf! Then Noah knew that the water had receded from the earth.
GEN|8|12|He waited seven more days and sent the dove out again, but this time it did not return to him.
GEN|8|13|By the first day of the first month of Noah's six hundred and first year, the water had dried up from the earth. Noah then removed the covering from the ark and saw that the surface of the ground was dry.
GEN|8|14|By the twenty-seventh day of the second month the earth was completely dry.
GEN|8|15|Then God said to Noah,
GEN|8|16|"Come out of the ark, you and your wife and your sons and their wives.
GEN|8|17|Bring out every kind of living creature that is with you-the birds, the animals, and all the creatures that move along the ground-so they can multiply on the earth and be fruitful and increase in number upon it."
GEN|8|18|So Noah came out, together with his sons and his wife and his sons' wives.
GEN|8|19|All the animals and all the creatures that move along the ground and all the birds-everything that moves on the earth-came out of the ark, one kind after another.
GEN|8|20|Then Noah built an altar to the LORD and, taking some of all the clean animals and clean birds, he sacrificed burnt offerings on it.
GEN|8|21|The LORD smelled the pleasing aroma and said in his heart: "Never again will I curse the ground because of man, even though every inclination of his heart is evil from childhood. And never again will I destroy all living creatures, as I have done.
GEN|8|22|"As long as the earth endures, seedtime and harvest, cold and heat, summer and winter, day and night will never cease."
GEN|9|1|Then God blessed Noah and his sons, saying to them, "Be fruitful and increase in number and fill the earth.
GEN|9|2|The fear and dread of you will fall upon all the beasts of the earth and all the birds of the air, upon every creature that moves along the ground, and upon all the fish of the sea; they are given into your hands.
GEN|9|3|Everything that lives and moves will be food for you. Just as I gave you the green plants, I now give you everything.
GEN|9|4|"But you must not eat meat that has its lifeblood still in it.
GEN|9|5|And for your lifeblood I will surely demand an accounting. I will demand an accounting from every animal. And from each man, too, I will demand an accounting for the life of his fellow man.
GEN|9|6|"Whoever sheds the blood of man, by man shall his blood be shed; for in the image of God has God made man.
GEN|9|7|As for you, be fruitful and increase in number; multiply on the earth and increase upon it."
GEN|9|8|Then God said to Noah and to his sons with him:
GEN|9|9|"I now establish my covenant with you and with your descendants after you
GEN|9|10|and with every living creature that was with you-the birds, the livestock and all the wild animals, all those that came out of the ark with you-every living creature on earth.
GEN|9|11|I establish my covenant with you: Never again will all life be cut off by the waters of a flood; never again will there be a flood to destroy the earth."
GEN|9|12|And God said, "This is the sign of the covenant I am making between me and you and every living creature with you, a covenant for all generations to come:
GEN|9|13|I have set my rainbow in the clouds, and it will be the sign of the covenant between me and the earth.
GEN|9|14|Whenever I bring clouds over the earth and the rainbow appears in the clouds,
GEN|9|15|I will remember my covenant between me and you and all living creatures of every kind. Never again will the waters become a flood to destroy all life.
GEN|9|16|Whenever the rainbow appears in the clouds, I will see it and remember the everlasting covenant between God and all living creatures of every kind on the earth."
GEN|9|17|So God said to Noah, "This is the sign of the covenant I have established between me and all life on the earth."
GEN|9|18|The sons of Noah who came out of the ark were Shem, Ham and Japheth. (Ham was the father of Canaan.)
GEN|9|19|These were the three sons of Noah, and from them came the people who were scattered over the earth.
GEN|9|20|Noah, a man of the soil, proceeded to plant a vineyard.
GEN|9|21|When he drank some of its wine, he became drunk and lay uncovered inside his tent.
GEN|9|22|Ham, the father of Canaan, saw his father's nakedness and told his two brothers outside.
GEN|9|23|But Shem and Japheth took a garment and laid it across their shoulders; then they walked in backward and covered their father's nakedness. Their faces were turned the other way so that they would not see their father's nakedness.
GEN|9|24|When Noah awoke from his wine and found out what his youngest son had done to him,
GEN|9|25|he said, "Cursed be Canaan! The lowest of slaves will he be to his brothers."
GEN|9|26|He also said, "Blessed be the LORD, the God of Shem! May Canaan be the slave of Shem.
GEN|9|27|May God extend the territory of Japheth; may Japheth live in the tents of Shem, and may Canaan be his slave."
GEN|9|28|After the flood Noah lived 350 years.
GEN|9|29|Altogether, Noah lived 950 years, and then he died.
GEN|10|1|This is the account of Shem, Ham and Japheth, Noah's sons, who themselves had sons after the flood. The Japhethites
GEN|10|2|The sons of Japheth: Gomer, Magog, Madai, Javan, Tubal, Meshech and Tiras.
GEN|10|3|The sons of Gomer: Ashkenaz, Riphath and Togarmah.
GEN|10|4|The sons of Javan: Elishah, Tarshish, the Kittim and the Rodanim.
GEN|10|5|(From these the maritime peoples spread out into their territories by their clans within their nations, each with its own language.) The Hamites
GEN|10|6|The sons of Ham: Cush, Mizraim, Put and Canaan.
GEN|10|7|The sons of Cush: Seba, Havilah, Sabtah, Raamah and Sabteca. The sons of Raamah: Sheba and Dedan.
GEN|10|8|Cush was the father of Nimrod, who grew to be a mighty warrior on the earth.
GEN|10|9|He was a mighty hunter before the LORD; that is why it is said, "Like Nimrod, a mighty hunter before the LORD."
GEN|10|10|The first centers of his kingdom were Babylon, Erech, Akkad and Calneh, in Shinar.
GEN|10|11|From that land he went to Assyria, where he built Nineveh, Rehoboth Ir, Calah
GEN|10|12|and Resen, which is between Nineveh and Calah; that is the great city.
GEN|10|13|Mizraim was the father of the Ludites, Anamites, Lehabites, Naphtuhites,
GEN|10|14|Pathrusites, Casluhites (from whom the Philistines came) and Caphtorites.
GEN|10|15|Canaan was the father of Sidon his firstborn, and of the Hittites,
GEN|10|16|Jebusites, Amorites, Girgashites,
GEN|10|17|Hivites, Arkites, Sinites,
GEN|10|18|Arvadites, Zemarites and Hamathites. Later the Canaanite clans scattered
GEN|10|19|and the borders of Canaan reached from Sidon toward Gerar as far as Gaza, and then toward Sodom, Gomorrah, Admah and Zeboiim, as far as Lasha.
GEN|10|20|These are the sons of Ham by their clans and languages, in their territories and nations. The Semites
GEN|10|21|Sons were also born to Shem, whose older brother was Japheth; Shem was the ancestor of all the sons of Eber.
GEN|10|22|The sons of Shem: Elam, Asshur, Arphaxad, Lud and Aram.
GEN|10|23|The sons of Aram: Uz, Hul, Gether and Meshech.
GEN|10|24|Arphaxad was the father of Shelah, and Shelah the father of Eber.
GEN|10|25|Two sons were born to Eber: One was named Peleg, because in his time the earth was divided; his brother was named Joktan.
GEN|10|26|Joktan was the father of Almodad, Sheleph, Hazarmaveth, Jerah,
GEN|10|27|Hadoram, Uzal, Diklah,
GEN|10|28|Obal, Abimael, Sheba,
GEN|10|29|Ophir, Havilah and Jobab. All these were sons of Joktan.
GEN|10|30|The region where they lived stretched from Mesha toward Sephar, in the eastern hill country.
GEN|10|31|These are the sons of Shem by their clans and languages, in their territories and nations.
GEN|10|32|These are the clans of Noah's sons, according to their lines of descent, within their nations. From these the nations spread out over the earth after the flood.
GEN|11|1|Now the whole world had one language and a common speech.
GEN|11|2|As men moved eastward, they found a plain in Shinar and settled there.
GEN|11|3|They said to each other, "Come, let's make bricks and bake them thoroughly." They used brick instead of stone, and tar for mortar.
GEN|11|4|Then they said, "Come, let us build ourselves a city, with a tower that reaches to the heavens, so that we may make a name for ourselves and not be scattered over the face of the whole earth."
GEN|11|5|But the LORD came down to see the city and the tower that the men were building.
GEN|11|6|The LORD said, "If as one people speaking the same language they have begun to do this, then nothing they plan to do will be impossible for them.
GEN|11|7|Come, let us go down and confuse their language so they will not understand each other."
GEN|11|8|So the LORD scattered them from there over all the earth, and they stopped building the city.
GEN|11|9|That is why it was called Babel -because there the LORD confused the language of the whole world. From there the LORD scattered them over the face of the whole earth.
GEN|11|10|This is the account of Shem. Two years after the flood, when Shem was 100 years old, he became the father of Arphaxad.
GEN|11|11|And after he became the father of Arphaxad, Shem lived 500 years and had other sons and daughters.
GEN|11|12|When Arphaxad had lived 35 years, he became the father of Shelah.
GEN|11|13|And after he became the father of Shelah, Arphaxad lived 403 years and had other sons and daughters.
GEN|11|14|When Shelah had lived 30 years, he became the father of Eber.
GEN|11|15|And after he became the father of Eber, Shelah lived 403 years and had other sons and daughters.
GEN|11|16|When Eber had lived 34 years, he became the father of Peleg.
GEN|11|17|And after he became the father of Peleg, Eber lived 430 years and had other sons and daughters.
GEN|11|18|When Peleg had lived 30 years, he became the father of Reu.
GEN|11|19|And after he became the father of Reu, Peleg lived 209 years and had other sons and daughters.
GEN|11|20|When Reu had lived 32 years, he became the father of Serug.
GEN|11|21|And after he became the father of Serug, Reu lived 207 years and had other sons and daughters.
GEN|11|22|When Serug had lived 30 years, he became the father of Nahor.
GEN|11|23|And after he became the father of Nahor, Serug lived 200 years and had other sons and daughters.
GEN|11|24|When Nahor had lived 29 years, he became the father of Terah.
GEN|11|25|And after he became the father of Terah, Nahor lived 119 years and had other sons and daughters.
GEN|11|26|After Terah had lived 70 years, he became the father of Abram, Nahor and Haran.
GEN|11|27|This is the account of Terah. Terah became the father of Abram, Nahor and Haran. And Haran became the father of Lot.
GEN|11|28|While his father Terah was still alive, Haran died in Ur of the Chaldeans, in the land of his birth.
GEN|11|29|Abram and Nahor both married. The name of Abram's wife was Sarai, and the name of Nahor's wife was Milcah; she was the daughter of Haran, the father of both Milcah and Iscah.
GEN|11|30|Now Sarai was barren; she had no children.
GEN|11|31|Terah took his son Abram, his grandson Lot son of Haran, and his daughter-in-law Sarai, the wife of his son Abram, and together they set out from Ur of the Chaldeans to go to Canaan. But when they came to Haran, they settled there.
GEN|11|32|Terah lived 205 years, and he died in Haran.
GEN|12|1|The LORD had said to Abram, "Leave your country, your people and your father's household and go to the land I will show you.
GEN|12|2|"I will make you into a great nation and I will bless you; I will make your name great, and you will be a blessing.
GEN|12|3|I will bless those who bless you, and whoever curses you I will curse; and all peoples on earth will be blessed through you."
GEN|12|4|So Abram left, as the LORD had told him; and Lot went with him. Abram was seventy-five years old when he set out from Haran.
GEN|12|5|He took his wife Sarai, his nephew Lot, all the possessions they had accumulated and the people they had acquired in Haran, and they set out for the land of Canaan, and they arrived there.
GEN|12|6|Abram traveled through the land as far as the site of the great tree of Moreh at Shechem. At that time the Canaanites were in the land.
GEN|12|7|The LORD appeared to Abram and said, "To your offspring I will give this land." So he built an altar there to the LORD, who had appeared to him.
GEN|12|8|From there he went on toward the hills east of Bethel and pitched his tent, with Bethel on the west and Ai on the east. There he built an altar to the LORD and called on the name of the LORD.
GEN|12|9|Then Abram set out and continued toward the Negev.
GEN|12|10|Now there was a famine in the land, and Abram went down to Egypt to live there for a while because the famine was severe.
GEN|12|11|As he was about to enter Egypt, he said to his wife Sarai, "I know what a beautiful woman you are.
GEN|12|12|When the Egyptians see you, they will say, 'This is his wife.' Then they will kill me but will let you live.
GEN|12|13|Say you are my sister, so that I will be treated well for your sake and my life will be spared because of you."
GEN|12|14|When Abram came to Egypt, the Egyptians saw that she was a very beautiful woman.
GEN|12|15|And when Pharaoh's officials saw her, they praised her to Pharaoh, and she was taken into his palace.
GEN|12|16|He treated Abram well for her sake, and Abram acquired sheep and cattle, male and female donkeys, menservants and maidservants, and camels.
GEN|12|17|But the LORD inflicted serious diseases on Pharaoh and his household because of Abram's wife Sarai.
GEN|12|18|So Pharaoh summoned Abram. "What have you done to me?" he said. "Why didn't you tell me she was your wife?
GEN|12|19|Why did you say, 'She is my sister,' so that I took her to be my wife? Now then, here is your wife. Take her and go!"
GEN|12|20|Then Pharaoh gave orders about Abram to his men, and they sent him on his way, with his wife and everything he had.
GEN|13|1|So Abram went up from Egypt to the Negev, with his wife and everything he had, and Lot went with him.
GEN|13|2|Abram had become very wealthy in livestock and in silver and gold.
GEN|13|3|From the Negev he went from place to place until he came to Bethel, to the place between Bethel and Ai where his tent had been earlier
GEN|13|4|and where he had first built an altar. There Abram called on the name of the LORD.
GEN|13|5|Now Lot, who was moving about with Abram, also had flocks and herds and tents.
GEN|13|6|But the land could not support them while they stayed together, for their possessions were so great that they were not able to stay together.
GEN|13|7|And quarreling arose between Abram's herdsmen and the herdsmen of Lot. The Canaanites and Perizzites were also living in the land at that time.
GEN|13|8|So Abram said to Lot, "Let's not have any quarreling between you and me, or between your herdsmen and mine, for we are brothers.
GEN|13|9|Is not the whole land before you? Let's part company. If you go to the left, I'll go to the right; if you go to the right, I'll go to the left."
GEN|13|10|Lot looked up and saw that the whole plain of the Jordan was well watered, like the garden of the LORD, like the land of Egypt, toward Zoar. (This was before the LORD destroyed Sodom and Gomorrah.)
GEN|13|11|So Lot chose for himself the whole plain of the Jordan and set out toward the east. The two men parted company:
GEN|13|12|Abram lived in the land of Canaan, while Lot lived among the cities of the plain and pitched his tents near Sodom.
GEN|13|13|Now the men of Sodom were wicked and were sinning greatly against the LORD.
GEN|13|14|The LORD said to Abram after Lot had parted from him, "Lift up your eyes from where you are and look north and south, east and west.
GEN|13|15|All the land that you see I will give to you and your offspring forever.
GEN|13|16|I will make your offspring like the dust of the earth, so that if anyone could count the dust, then your offspring could be counted.
GEN|13|17|Go, walk through the length and breadth of the land, for I am giving it to you."
GEN|13|18|So Abram moved his tents and went to live near the great trees of Mamre at Hebron, where he built an altar to the LORD.
GEN|14|1|At this time Amraphel king of Shinar, Arioch king of Ellasar, Kedorlaomer king of Elam and Tidal king of Goiim
GEN|14|2|went to war against Bera king of Sodom, Birsha king of Gomorrah, Shinab king of Admah, Shemeber king of Zeboiim, and the king of Bela (that is, Zoar).
GEN|14|3|All these latter kings joined forces in the Valley of Siddim (the Salt Sea ).
GEN|14|4|For twelve years they had been subject to Kedorlaomer, but in the thirteenth year they rebelled.
GEN|14|5|In the fourteenth year, Kedorlaomer and the kings allied with him went out and defeated the Rephaites in Ashteroth Karnaim, the Zuzites in Ham, the Emites in Shaveh Kiriathaim
GEN|14|6|and the Horites in the hill country of Seir, as far as El Paran near the desert.
GEN|14|7|Then they turned back and went to En Mishpat (that is, Kadesh), and they conquered the whole territory of the Amalekites, as well as the Amorites who were living in Hazazon Tamar.
GEN|14|8|Then the king of Sodom, the king of Gomorrah, the king of Admah, the king of Zeboiim and the king of Bela (that is, Zoar) marched out and drew up their battle lines in the Valley of Siddim
GEN|14|9|against Kedorlaomer king of Elam, Tidal king of Goiim, Amraphel king of Shinar and Arioch king of Ellasar-four kings against five.
GEN|14|10|Now the Valley of Siddim was full of tar pits, and when the kings of Sodom and Gomorrah fled, some of the men fell into them and the rest fled to the hills.
GEN|14|11|The four kings seized all the goods of Sodom and Gomorrah and all their food; then they went away.
GEN|14|12|They also carried off Abram's nephew Lot and his possessions, since he was living in Sodom.
GEN|14|13|One who had escaped came and reported this to Abram the Hebrew. Now Abram was living near the great trees of Mamre the Amorite, a brother of Eshcol and Aner, all of whom were allied with Abram.
GEN|14|14|When Abram heard that his relative had been taken captive, he called out the 318 trained men born in his household and went in pursuit as far as Dan.
GEN|14|15|During the night Abram divided his men to attack them and he routed them, pursuing them as far as Hobah, north of Damascus.
GEN|14|16|He recovered all the goods and brought back his relative Lot and his possessions, together with the women and the other people.
GEN|14|17|After Abram returned from defeating Kedorlaomer and the kings allied with him, the king of Sodom came out to meet him in the Valley of Shaveh (that is, the King's Valley).
GEN|14|18|Then Melchizedek king of Salem brought out bread and wine. He was priest of God Most High,
GEN|14|19|and he blessed Abram, saying, "Blessed be Abram by God Most High, Creator of heaven and earth.
GEN|14|20|And blessed be God Most High, who delivered your enemies into your hand." Then Abram gave him a tenth of everything.
GEN|14|21|The king of Sodom said to Abram, "Give me the people and keep the goods for yourself."
GEN|14|22|But Abram said to the king of Sodom, "I have raised my hand to the LORD, God Most High, Creator of heaven and earth, and have taken an oath
GEN|14|23|that I will accept nothing belonging to you, not even a thread or the thong of a sandal, so that you will never be able to say, 'I made Abram rich.'
GEN|14|24|I will accept nothing but what my men have eaten and the share that belongs to the men who went with me-to Aner, Eshcol and Mamre. Let them have their share."
GEN|15|1|After this, the word of the LORD came to Abram in a vision: "Do not be afraid, Abram. I am your shield, your very great reward. "
GEN|15|2|But Abram said, "O Sovereign LORD, what can you give me since I remain childless and the one who will inherit my estate is Eliezer of Damascus?"
GEN|15|3|And Abram said, "You have given me no children; so a servant in my household will be my heir."
GEN|15|4|Then the word of the LORD came to him: "This man will not be your heir, but a son coming from your own body will be your heir."
GEN|15|5|He took him outside and said, "Look up at the heavens and count the stars-if indeed you can count them." Then he said to him, "So shall your offspring be."
GEN|15|6|Abram believed the LORD, and he credited it to him as righteousness.
GEN|15|7|He also said to him, "I am the LORD, who brought you out of Ur of the Chaldeans to give you this land to take possession of it."
GEN|15|8|But Abram said, "O Sovereign LORD, how can I know that I will gain possession of it?"
GEN|15|9|So the LORD said to him, "Bring me a heifer, a goat and a ram, each three years old, along with a dove and a young pigeon."
GEN|15|10|Abram brought all these to him, cut them in two and arranged the halves opposite each other; the birds, however, he did not cut in half.
GEN|15|11|Then birds of prey came down on the carcasses, but Abram drove them away.
GEN|15|12|As the sun was setting, Abram fell into a deep sleep, and a thick and dreadful darkness came over him.
GEN|15|13|Then the LORD said to him, "Know for certain that your descendants will be strangers in a country not their own, and they will be enslaved and mistreated four hundred years.
GEN|15|14|But I will punish the nation they serve as slaves, and afterward they will come out with great possessions.
GEN|15|15|You, however, will go to your fathers in peace and be buried at a good old age.
GEN|15|16|In the fourth generation your descendants will come back here, for the sin of the Amorites has not yet reached its full measure."
GEN|15|17|When the sun had set and darkness had fallen, a smoking firepot with a blazing torch appeared and passed between the pieces.
GEN|15|18|On that day the LORD made a covenant with Abram and said, "To your descendants I give this land, from the river of Egypt to the great river, the Euphrates-
GEN|15|19|the land of the Kenites, Kenizzites, Kadmonites,
GEN|15|20|Hittites, Perizzites, Rephaites,
GEN|15|21|Amorites, Canaanites, Girgashites and Jebusites."
GEN|16|1|Now Sarai, Abram's wife, had borne him no children. But she had an Egyptian maidservant named Hagar;
GEN|16|2|so she said to Abram, "The LORD has kept me from having children. Go, sleep with my maidservant; perhaps I can build a family through her." Abram agreed to what Sarai said.
GEN|16|3|So after Abram had been living in Canaan ten years, Sarai his wife took her Egyptian maidservant Hagar and gave her to her husband to be his wife.
GEN|16|4|He slept with Hagar, and she conceived. When she knew she was pregnant, she began to despise her mistress.
GEN|16|5|Then Sarai said to Abram, "You are responsible for the wrong I am suffering. I put my servant in your arms, and now that she knows she is pregnant, she despises me. May the LORD judge between you and me."
GEN|16|6|"Your servant is in your hands," Abram said. "Do with her whatever you think best." Then Sarai mistreated Hagar; so she fled from her.
GEN|16|7|The angel of the LORD found Hagar near a spring in the desert; it was the spring that is beside the road to Shur.
GEN|16|8|And he said, "Hagar, servant of Sarai, where have you come from, and where are you going?I'm running away from my mistress Sarai," she answered.
GEN|16|9|Then the angel of the LORD told her, "Go back to your mistress and submit to her."
GEN|16|10|The angel added, "I will so increase your descendants that they will be too numerous to count."
GEN|16|11|The angel of the LORD also said to her: "You are now with child and you will have a son. You shall name him Ishmael, for the LORD has heard of your misery.
GEN|16|12|He will be a wild donkey of a man; his hand will be against everyone and everyone's hand against him, and he will live in hostility toward all his brothers."
GEN|16|13|She gave this name to the LORD who spoke to her: "You are the God who sees me," for she said, "I have now seen the One who sees me."
GEN|16|14|That is why the well was called Beer Lahai Roi; it is still there, between Kadesh and Bered.
GEN|16|15|So Hagar bore Abram a son, and Abram gave the name Ishmael to the son she had borne.
GEN|16|16|Abram was eighty-six years old when Hagar bore him Ishmael.
GEN|17|1|When Abram was ninety-nine years old, the LORD appeared to him and said, "I am God Almighty; walk before me and be blameless.
GEN|17|2|I will confirm my covenant between me and you and will greatly increase your numbers."
GEN|17|3|Abram fell facedown, and God said to him,
GEN|17|4|"As for me, this is my covenant with you: You will be the father of many nations.
GEN|17|5|No longer will you be called Abram; your name will be Abraham, for I have made you a father of many nations.
GEN|17|6|I will make you very fruitful; I will make nations of you, and kings will come from you.
GEN|17|7|I will establish my covenant as an everlasting covenant between me and you and your descendants after you for the generations to come, to be your God and the God of your descendants after you.
GEN|17|8|The whole land of Canaan, where you are now an alien, I will give as an everlasting possession to you and your descendants after you; and I will be their God."
GEN|17|9|Then God said to Abraham, "As for you, you must keep my covenant, you and your descendants after you for the generations to come.
GEN|17|10|This is my covenant with you and your descendants after you, the covenant you are to keep: Every male among you shall be circumcised.
GEN|17|11|You are to undergo circumcision, and it will be the sign of the covenant between me and you.
GEN|17|12|For the generations to come every male among you who is eight days old must be circumcised, including those born in your household or bought with money from a foreigner-those who are not your offspring.
GEN|17|13|Whether born in your household or bought with your money, they must be circumcised. My covenant in your flesh is to be an everlasting covenant.
GEN|17|14|Any uncircumcised male, who has not been circumcised in the flesh, will be cut off from his people; he has broken my covenant."
GEN|17|15|God also said to Abraham, "As for Sarai your wife, you are no longer to call her Sarai; her name will be Sarah.
GEN|17|16|I will bless her and will surely give you a son by her. I will bless her so that she will be the mother of nations; kings of peoples will come from her."
GEN|17|17|Abraham fell facedown; he laughed and said to himself, "Will a son be born to a man a hundred years old? Will Sarah bear a child at the age of ninety?"
GEN|17|18|And Abraham said to God, "If only Ishmael might live under your blessing!"
GEN|17|19|Then God said, "Yes, but your wife Sarah will bear you a son, and you will call him Isaac. I will establish my covenant with him as an everlasting covenant for his descendants after him.
GEN|17|20|And as for Ishmael, I have heard you: I will surely bless him; I will make him fruitful and will greatly increase his numbers. He will be the father of twelve rulers, and I will make him into a great nation.
GEN|17|21|But my covenant I will establish with Isaac, whom Sarah will bear to you by this time next year."
GEN|17|22|When he had finished speaking with Abraham, God went up from him.
GEN|17|23|On that very day Abraham took his son Ishmael and all those born in his household or bought with his money, every male in his household, and circumcised them, as God told him.
GEN|17|24|Abraham was ninety-nine years old when he was circumcised,
GEN|17|25|and his son Ishmael was thirteen;
GEN|17|26|Abraham and his son Ishmael were both circumcised on that same day.
GEN|17|27|And every male in Abraham's household, including those born in his household or bought from a foreigner, was circumcised with him.
GEN|18|1|The LORD appeared to Abraham near the great trees of Mamre while he was sitting at the entrance to his tent in the heat of the day.
GEN|18|2|Abraham looked up and saw three men standing nearby. When he saw them, he hurried from the entrance of his tent to meet them and bowed low to the ground.
GEN|18|3|He said, "If I have found favor in your eyes, my lord, do not pass your servant by.
GEN|18|4|Let a little water be brought, and then you may all wash your feet and rest under this tree.
GEN|18|5|Let me get you something to eat, so you can be refreshed and then go on your way-now that you have come to your servant.Very well," they answered, "do as you say."
GEN|18|6|So Abraham hurried into the tent to Sarah. "Quick," he said, "get three seahs of fine flour and knead it and bake some bread."
GEN|18|7|Then he ran to the herd and selected a choice, tender calf and gave it to a servant, who hurried to prepare it.
GEN|18|8|He then brought some curds and milk and the calf that had been prepared, and set these before them. While they ate, he stood near them under a tree.
GEN|18|9|"Where is your wife Sarah?" they asked him. "There, in the tent," he said.
GEN|18|10|Then the LORD said, "I will surely return to you about this time next year, and Sarah your wife will have a son." Now Sarah was listening at the entrance to the tent, which was behind him.
GEN|18|11|Abraham and Sarah were already old and well advanced in years, and Sarah was past the age of childbearing.
GEN|18|12|So Sarah laughed to herself as she thought, "After I am worn out and my master is old, will I now have this pleasure?"
GEN|18|13|Then the LORD said to Abraham, "Why did Sarah laugh and say, 'Will I really have a child, now that I am old?'
GEN|18|14|Is anything too hard for the LORD? I will return to you at the appointed time next year and Sarah will have a son."
GEN|18|15|Sarah was afraid, so she lied and said, "I did not laugh." But he said, "Yes, you did laugh."
GEN|18|16|When the men got up to leave, they looked down toward Sodom, and Abraham walked along with them to see them on their way.
GEN|18|17|Then the LORD said, "Shall I hide from Abraham what I am about to do?
GEN|18|18|Abraham will surely become a great and powerful nation, and all nations on earth will be blessed through him.
GEN|18|19|For I have chosen him, so that he will direct his children and his household after him to keep the way of the LORD by doing what is right and just, so that the LORD will bring about for Abraham what he has promised him."
GEN|18|20|Then the LORD said, "The outcry against Sodom and Gomorrah is so great and their sin so grievous
GEN|18|21|that I will go down and see if what they have done is as bad as the outcry that has reached me. If not, I will know."
GEN|18|22|The men turned away and went toward Sodom, but Abraham remained standing before the LORD.
GEN|18|23|Then Abraham approached him and said: "Will you sweep away the righteous with the wicked?
GEN|18|24|What if there are fifty righteous people in the city? Will you really sweep it away and not spare the place for the sake of the fifty righteous people in it?
GEN|18|25|Far be it from you to do such a thing-to kill the righteous with the wicked, treating the righteous and the wicked alike. Far be it from you! Will not the Judge of all the earth do right?"
GEN|18|26|The LORD said, "If I find fifty righteous people in the city of Sodom, I will spare the whole place for their sake."
GEN|18|27|Then Abraham spoke up again: "Now that I have been so bold as to speak to the Lord, though I am nothing but dust and ashes,
GEN|18|28|what if the number of the righteous is five less than fifty? Will you destroy the whole city because of five people?If I find forty-five there," he said, "I will not destroy it."
GEN|18|29|Once again he spoke to him, "What if only forty are found there?" He said, "For the sake of forty, I will not do it."
GEN|18|30|Then he said, "May the Lord not be angry, but let me speak. What if only thirty can be found there?" He answered, "I will not do it if I find thirty there."
GEN|18|31|Abraham said, "Now that I have been so bold as to speak to the Lord, what if only twenty can be found there?" He said, "For the sake of twenty, I will not destroy it."
GEN|18|32|Then he said, "May the Lord not be angry, but let me speak just once more. What if only ten can be found there?" He answered, "For the sake of ten, I will not destroy it."
GEN|18|33|When the LORD had finished speaking with Abraham, he left, and Abraham returned home.
GEN|19|1|The two angels arrived at Sodom in the evening, and Lot was sitting in the gateway of the city. When he saw them, he got up to meet them and bowed down with his face to the ground.
GEN|19|2|"My lords," he said, "please turn aside to your servant's house. You can wash your feet and spend the night and then go on your way early in the morning.No," they answered, "we will spend the night in the square."
GEN|19|3|But he insisted so strongly that they did go with him and entered his house. He prepared a meal for them, baking bread without yeast, and they ate.
GEN|19|4|Before they had gone to bed, all the men from every part of the city of Sodom-both young and old-surrounded the house.
GEN|19|5|They called to Lot, "Where are the men who came to you tonight? Bring them out to us so that we can have sex with them."
GEN|19|6|Lot went outside to meet them and shut the door behind him
GEN|19|7|and said, "No, my friends. Don't do this wicked thing.
GEN|19|8|Look, I have two daughters who have never slept with a man. Let me bring them out to you, and you can do what you like with them. But don't do anything to these men, for they have come under the protection of my roof."
GEN|19|9|"Get out of our way," they replied. And they said, "This fellow came here as an alien, and now he wants to play the judge! We'll treat you worse than them." They kept bringing pressure on Lot and moved forward to break down the door.
GEN|19|10|But the men inside reached out and pulled Lot back into the house and shut the door.
GEN|19|11|Then they struck the men who were at the door of the house, young and old, with blindness so that they could not find the door.
GEN|19|12|The two men said to Lot, "Do you have anyone else here-sons-in-law, sons or daughters, or anyone else in the city who belongs to you? Get them out of here,
GEN|19|13|because we are going to destroy this place. The outcry to the LORD against its people is so great that he has sent us to destroy it."
GEN|19|14|So Lot went out and spoke to his sons-in-law, who were pledged to marry his daughters. He said, "Hurry and get out of this place, because the LORD is about to destroy the city!" But his sons-in-law thought he was joking.
GEN|19|15|With the coming of dawn, the angels urged Lot, saying, "Hurry! Take your wife and your two daughters who are here, or you will be swept away when the city is punished."
GEN|19|16|When he hesitated, the men grasped his hand and the hands of his wife and of his two daughters and led them safely out of the city, for the LORD was merciful to them.
GEN|19|17|As soon as they had brought them out, one of them said, "Flee for your lives! Don't look back, and don't stop anywhere in the plain! Flee to the mountains or you will be swept away!"
GEN|19|18|But Lot said to them, "No, my lords, please!
GEN|19|19|Your servant has found favor in your eyes, and you have shown great kindness to me in sparing my life. But I can't flee to the mountains; this disaster will overtake me, and I'll die.
GEN|19|20|Look, here is a town near enough to run to, and it is small. Let me flee to it-it is very small, isn't it? Then my life will be spared."
GEN|19|21|He said to him, "Very well, I will grant this request too; I will not overthrow the town you speak of.
GEN|19|22|But flee there quickly, because I cannot do anything until you reach it." (That is why the town was called Zoar. )
GEN|19|23|By the time Lot reached Zoar, the sun had risen over the land.
GEN|19|24|Then the LORD rained down burning sulfur on Sodom and Gomorrah-from the LORD out of the heavens.
GEN|19|25|Thus he overthrew those cities and the entire plain, including all those living in the cities-and also the vegetation in the land.
GEN|19|26|But Lot's wife looked back, and she became a pillar of salt.
GEN|19|27|Early the next morning Abraham got up and returned to the place where he had stood before the LORD.
GEN|19|28|He looked down toward Sodom and Gomorrah, toward all the land of the plain, and he saw dense smoke rising from the land, like smoke from a furnace.
GEN|19|29|So when God destroyed the cities of the plain, he remembered Abraham, and he brought Lot out of the catastrophe that overthrew the cities where Lot had lived.
GEN|19|30|Lot and his two daughters left Zoar and settled in the mountains, for he was afraid to stay in Zoar. He and his two daughters lived in a cave.
GEN|19|31|One day the older daughter said to the younger, "Our father is old, and there is no man around here to lie with us, as is the custom all over the earth.
GEN|19|32|Let's get our father to drink wine and then lie with him and preserve our family line through our father."
GEN|19|33|That night they got their father to drink wine, and the older daughter went in and lay with him. He was not aware of it when she lay down or when she got up.
GEN|19|34|The next day the older daughter said to the younger, "Last night I lay with my father. Let's get him to drink wine again tonight, and you go in and lie with him so we can preserve our family line through our father."
GEN|19|35|So they got their father to drink wine that night also, and the younger daughter went and lay with him. Again he was not aware of it when she lay down or when she got up.
GEN|19|36|So both of Lot's daughters became pregnant by their father.
GEN|19|37|The older daughter had a son, and she named him Moab; he is the father of the Moabites of today.
GEN|19|38|The younger daughter also had a son, and she named him Ben-Ammi; he is the father of the Ammonites of today.
GEN|20|1|Now Abraham moved on from there into the region of the Negev and lived between Kadesh and Shur. For a while he stayed in Gerar,
GEN|20|2|and there Abraham said of his wife Sarah, "She is my sister." Then Abimelech king of Gerar sent for Sarah and took her.
GEN|20|3|But God came to Abimelech in a dream one night and said to him, "You are as good as dead because of the woman you have taken; she is a married woman."
GEN|20|4|Now Abimelech had not gone near her, so he said, "Lord, will you destroy an innocent nation?
GEN|20|5|Did he not say to me, 'She is my sister,' and didn't she also say, 'He is my brother'? I have done this with a clear conscience and clean hands."
GEN|20|6|Then God said to him in the dream, "Yes, I know you did this with a clear conscience, and so I have kept you from sinning against me. That is why I did not let you touch her.
GEN|20|7|Now return the man's wife, for he is a prophet, and he will pray for you and you will live. But if you do not return her, you may be sure that you and all yours will die."
GEN|20|8|Early the next morning Abimelech summoned all his officials, and when he told them all that had happened, they were very much afraid.
GEN|20|9|Then Abimelech called Abraham in and said, "What have you done to us? How have I wronged you that you have brought such great guilt upon me and my kingdom? You have done things to me that should not be done."
GEN|20|10|And Abimelech asked Abraham, "What was your reason for doing this?"
GEN|20|11|Abraham replied, "I said to myself, 'There is surely no fear of God in this place, and they will kill me because of my wife.'
GEN|20|12|Besides, she really is my sister, the daughter of my father though not of my mother; and she became my wife.
GEN|20|13|And when God had me wander from my father's household, I said to her, 'This is how you can show your love to me: Everywhere we go, say of me, "He is my brother."'"
GEN|20|14|Then Abimelech brought sheep and cattle and male and female slaves and gave them to Abraham, and he returned Sarah his wife to him.
GEN|20|15|And Abimelech said, "My land is before you; live wherever you like."
GEN|20|16|To Sarah he said, "I am giving your brother a thousand shekels of silver. This is to cover the offense against you before all who are with you; you are completely vindicated."
GEN|20|17|Then Abraham prayed to God, and God healed Abimelech, his wife and his slave girls so they could have children again,
GEN|20|18|for the LORD had closed up every womb in Abimelech's household because of Abraham's wife Sarah.
GEN|21|1|Now the LORD was gracious to Sarah as he had said, and the LORD did for Sarah what he had promised.
GEN|21|2|Sarah became pregnant and bore a son to Abraham in his old age, at the very time God had promised him.
GEN|21|3|Abraham gave the name Isaac to the son Sarah bore him.
GEN|21|4|When his son Isaac was eight days old, Abraham circumcised him, as God commanded him.
GEN|21|5|Abraham was a hundred years old when his son Isaac was born to him.
GEN|21|6|Sarah said, "God has brought me laughter, and everyone who hears about this will laugh with me."
GEN|21|7|And she added, "Who would have said to Abraham that Sarah would nurse children? Yet I have borne him a son in his old age."
GEN|21|8|The child grew and was weaned, and on the day Isaac was weaned Abraham held a great feast.
GEN|21|9|But Sarah saw that the son whom Hagar the Egyptian had borne to Abraham was mocking,
GEN|21|10|and she said to Abraham, "Get rid of that slave woman and her son, for that slave woman's son will never share in the inheritance with my son Isaac."
GEN|21|11|The matter distressed Abraham greatly because it concerned his son.
GEN|21|12|But God said to him, "Do not be so distressed about the boy and your maidservant. Listen to whatever Sarah tells you, because it is through Isaac that your offspring will be reckoned.
GEN|21|13|I will make the son of the maidservant into a nation also, because he is your offspring."
GEN|21|14|Early the next morning Abraham took some food and a skin of water and gave them to Hagar. He set them on her shoulders and then sent her off with the boy. She went on her way and wandered in the desert of Beersheba.
GEN|21|15|When the water in the skin was gone, she put the boy under one of the bushes.
GEN|21|16|Then she went off and sat down nearby, about a bowshot away, for she thought, "I cannot watch the boy die." And as she sat there nearby, she began to sob.
GEN|21|17|God heard the boy crying, and the angel of God called to Hagar from heaven and said to her, "What is the matter, Hagar? Do not be afraid; God has heard the boy crying as he lies there.
GEN|21|18|Lift the boy up and take him by the hand, for I will make him into a great nation."
GEN|21|19|Then God opened her eyes and she saw a well of water. So she went and filled the skin with water and gave the boy a drink.
GEN|21|20|God was with the boy as he grew up. He lived in the desert and became an archer.
GEN|21|21|While he was living in the Desert of Paran, his mother got a wife for him from Egypt.
GEN|21|22|At that time Abimelech and Phicol the commander of his forces said to Abraham, "God is with you in everything you do.
GEN|21|23|Now swear to me here before God that you will not deal falsely with me or my children or my descendants. Show to me and the country where you are living as an alien the same kindness I have shown to you."
GEN|21|24|Abraham said, "I swear it."
GEN|21|25|Then Abraham complained to Abimelech about a well of water that Abimelech's servants had seized.
GEN|21|26|But Abimelech said, "I don't know who has done this. You did not tell me, and I heard about it only today."
GEN|21|27|So Abraham brought sheep and cattle and gave them to Abimelech, and the two men made a treaty.
GEN|21|28|Abraham set apart seven ewe lambs from the flock,
GEN|21|29|and Abimelech asked Abraham, "What is the meaning of these seven ewe lambs you have set apart by themselves?"
GEN|21|30|He replied, "Accept these seven lambs from my hand as a witness that I dug this well."
GEN|21|31|So that place was called Beersheba, because the two men swore an oath there.
GEN|21|32|After the treaty had been made at Beersheba, Abimelech and Phicol the commander of his forces returned to the land of the Philistines.
GEN|21|33|Abraham planted a tamarisk tree in Beersheba, and there he called upon the name of the LORD, the Eternal God.
GEN|21|34|And Abraham stayed in the land of the Philistines for a long time.
GEN|22|1|Some time later God tested Abraham. He said to him, "Abraham!Here I am," he replied.
GEN|22|2|Then God said, "Take your son, your only son, Isaac, whom you love, and go to the region of Moriah. Sacrifice him there as a burnt offering on one of the mountains I will tell you about."
GEN|22|3|Early the next morning Abraham got up and saddled his donkey. He took with him two of his servants and his son Isaac. When he had cut enough wood for the burnt offering, he set out for the place God had told him about.
GEN|22|4|On the third day Abraham looked up and saw the place in the distance.
GEN|22|5|He said to his servants, "Stay here with the donkey while I and the boy go over there. We will worship and then we will come back to you."
GEN|22|6|Abraham took the wood for the burnt offering and placed it on his son Isaac, and he himself carried the fire and the knife. As the two of them went on together,
GEN|22|7|Isaac spoke up and said to his father Abraham, "Father?Yes, my son?" Abraham replied. "The fire and wood are here," Isaac said, "but where is the lamb for the burnt offering?"
GEN|22|8|Abraham answered, "God himself will provide the lamb for the burnt offering, my son." And the two of them went on together.
GEN|22|9|When they reached the place God had told him about, Abraham built an altar there and arranged the wood on it. He bound his son Isaac and laid him on the altar, on top of the wood.
GEN|22|10|Then he reached out his hand and took the knife to slay his son.
GEN|22|11|But the angel of the LORD called out to him from heaven, "Abraham! Abraham!Here I am," he replied.
GEN|22|12|"Do not lay a hand on the boy," he said. "Do not do anything to him. Now I know that you fear God, because you have not withheld from me your son, your only son."
GEN|22|13|Abraham looked up and there in a thicket he saw a ram caught by its horns. He went over and took the ram and sacrificed it as a burnt offering instead of his son.
GEN|22|14|So Abraham called that place The LORD Will Provide. And to this day it is said, "On the mountain of the LORD it will be provided."
GEN|22|15|The angel of the LORD called to Abraham from heaven a second time
GEN|22|16|and said, "I swear by myself, declares the LORD, that because you have done this and have not withheld your son, your only son,
GEN|22|17|I will surely bless you and make your descendants as numerous as the stars in the sky and as the sand on the seashore. Your descendants will take possession of the cities of their enemies,
GEN|22|18|and through your offspring all nations on earth will be blessed, because you have obeyed me."
GEN|22|19|Then Abraham returned to his servants, and they set off together for Beersheba. And Abraham stayed in Beersheba.
GEN|22|20|Some time later Abraham was told, "Milcah is also a mother; she has borne sons to your brother Nahor:
GEN|22|21|Uz the firstborn, Buz his brother, Kemuel (the father of Aram),
GEN|22|22|Kesed, Hazo, Pildash, Jidlaph and Bethuel."
GEN|22|23|Bethuel became the father of Rebekah. Milcah bore these eight sons to Abraham's brother Nahor.
GEN|22|24|His concubine, whose name was Reumah, also had sons: Tebah, Gaham, Tahash and Maacah.
GEN|23|1|Sarah lived to be a hundred and twenty-seven years old.
GEN|23|2|She died at Kiriath Arba (that is, Hebron) in the land of Canaan, and Abraham went to mourn for Sarah and to weep over her.
GEN|23|3|Then Abraham rose from beside his dead wife and spoke to the Hittites. He said,
GEN|23|4|"I am an alien and a stranger among you. Sell me some property for a burial site here so I can bury my dead."
GEN|23|5|The Hittites replied to Abraham,
GEN|23|6|"Sir, listen to us. You are a mighty prince among us. Bury your dead in the choicest of our tombs. None of us will refuse you his tomb for burying your dead."
GEN|23|7|Then Abraham rose and bowed down before the people of the land, the Hittites.
GEN|23|8|He said to them, "If you are willing to let me bury my dead, then listen to me and intercede with Ephron son of Zohar on my behalf
GEN|23|9|so he will sell me the cave of Machpelah, which belongs to him and is at the end of his field. Ask him to sell it to me for the full price as a burial site among you."
GEN|23|10|Ephron the Hittite was sitting among his people and he replied to Abraham in the hearing of all the Hittites who had come to the gate of his city.
GEN|23|11|"No, my lord," he said. "Listen to me; I give you the field, and I give you the cave that is in it. I give it to you in the presence of my people. Bury your dead."
GEN|23|12|Again Abraham bowed down before the people of the land
GEN|23|13|and he said to Ephron in their hearing, "Listen to me, if you will. I will pay the price of the field. Accept it from me so I can bury my dead there."
GEN|23|14|Ephron answered Abraham,
GEN|23|15|"Listen to me, my lord; the land is worth four hundred shekels of silver, but what is that between me and you? Bury your dead."
GEN|23|16|Abraham agreed to Ephron's terms and weighed out for him the price he had named in the hearing of the Hittites: four hundred shekels of silver, according to the weight current among the merchants.
GEN|23|17|So Ephron's field in Machpelah near Mamre-both the field and the cave in it, and all the trees within the borders of the field-was deeded
GEN|23|18|to Abraham as his property in the presence of all the Hittites who had come to the gate of the city.
GEN|23|19|Afterward Abraham buried his wife Sarah in the cave in the field of Machpelah near Mamre (which is at Hebron) in the land of Canaan.
GEN|23|20|So the field and the cave in it were deeded to Abraham by the Hittites as a burial site.
GEN|24|1|Abraham was now old and well advanced in years, and the LORD had blessed him in every way.
GEN|24|2|He said to the chief servant in his household, the one in charge of all that he had, "Put your hand under my thigh.
GEN|24|3|I want you to swear by the LORD, the God of heaven and the God of earth, that you will not get a wife for my son from the daughters of the Canaanites, among whom I am living,
GEN|24|4|but will go to my country and my own relatives and get a wife for my son Isaac."
GEN|24|5|The servant asked him, "What if the woman is unwilling to come back with me to this land? Shall I then take your son back to the country you came from?"
GEN|24|6|"Make sure that you do not take my son back there," Abraham said.
GEN|24|7|"The LORD, the God of heaven, who brought me out of my father's household and my native land and who spoke to me and promised me on oath, saying, 'To your offspring I will give this land'-he will send his angel before you so that you can get a wife for my son from there.
GEN|24|8|If the woman is unwilling to come back with you, then you will be released from this oath of mine. Only do not take my son back there."
GEN|24|9|So the servant put his hand under the thigh of his master Abraham and swore an oath to him concerning this matter.
GEN|24|10|Then the servant took ten of his master's camels and left, taking with him all kinds of good things from his master. He set out for Aram Naharaim and made his way to the town of Nahor.
GEN|24|11|He had the camels kneel down near the well outside the town; it was toward evening, the time the women go out to draw water.
GEN|24|12|Then he prayed, "O LORD, God of my master Abraham, give me success today, and show kindness to my master Abraham.
GEN|24|13|See, I am standing beside this spring, and the daughters of the townspeople are coming out to draw water.
GEN|24|14|May it be that when I say to a girl, 'Please let down your jar that I may have a drink,' and she says, 'Drink, and I'll water your camels too'-let her be the one you have chosen for your servant Isaac. By this I will know that you have shown kindness to my master."
GEN|24|15|Before he had finished praying, Rebekah came out with her jar on her shoulder. She was the daughter of Bethuel son of Milcah, who was the wife of Abraham's brother Nahor.
GEN|24|16|The girl was very beautiful, a virgin; no man had ever lain with her. She went down to the spring, filled her jar and came up again.
GEN|24|17|The servant hurried to meet her and said, "Please give me a little water from your jar."
GEN|24|18|"Drink, my lord," she said, and quickly lowered the jar to her hands and gave him a drink.
GEN|24|19|After she had given him a drink, she said, "I'll draw water for your camels too, until they have finished drinking."
GEN|24|20|So she quickly emptied her jar into the trough, ran back to the well to draw more water, and drew enough for all his camels.
GEN|24|21|Without saying a word, the man watched her closely to learn whether or not the LORD had made his journey successful.
GEN|24|22|When the camels had finished drinking, the man took out a gold nose ring weighing a beka and two gold bracelets weighing ten shekels.
GEN|24|23|Then he asked, "Whose daughter are you? Please tell me, is there room in your father's house for us to spend the night?"
GEN|24|24|She answered him, "I am the daughter of Bethuel, the son that Milcah bore to Nahor."
GEN|24|25|And she added, "We have plenty of straw and fodder, as well as room for you to spend the night."
GEN|24|26|Then the man bowed down and worshiped the LORD,
GEN|24|27|saying, "Praise be to the LORD, the God of my master Abraham, who has not abandoned his kindness and faithfulness to my master. As for me, the LORD has led me on the journey to the house of my master's relatives."
GEN|24|28|The girl ran and told her mother's household about these things.
GEN|24|29|Now Rebekah had a brother named Laban, and he hurried out to the man at the spring.
GEN|24|30|As soon as he had seen the nose ring, and the bracelets on his sister's arms, and had heard Rebekah tell what the man said to her, he went out to the man and found him standing by the camels near the spring.
GEN|24|31|"Come, you who are blessed by the LORD," he said. "Why are you standing out here? I have prepared the house and a place for the camels."
GEN|24|32|So the man went to the house, and the camels were unloaded. Straw and fodder were brought for the camels, and water for him and his men to wash their feet.
GEN|24|33|Then food was set before him, but he said, "I will not eat until I have told you what I have to say.Then tell us," Laban said.
GEN|24|34|So he said, "I am Abraham's servant.
GEN|24|35|The LORD has blessed my master abundantly, and he has become wealthy. He has given him sheep and cattle, silver and gold, menservants and maidservants, and camels and donkeys.
GEN|24|36|My master's wife Sarah has borne him a son in her old age, and he has given him everything he owns.
GEN|24|37|And my master made me swear an oath, and said, 'You must not get a wife for my son from the daughters of the Canaanites, in whose land I live,
GEN|24|38|but go to my father's family and to my own clan, and get a wife for my son.'
GEN|24|39|"Then I asked my master, 'What if the woman will not come back with me?'
GEN|24|40|"He replied, 'The LORD, before whom I have walked, will send his angel with you and make your journey a success, so that you can get a wife for my son from my own clan and from my father's family.
GEN|24|41|Then, when you go to my clan, you will be released from my oath even if they refuse to give her to you-you will be released from my oath.'
GEN|24|42|"When I came to the spring today, I said, 'O LORD, God of my master Abraham, if you will, please grant success to the journey on which I have come.
GEN|24|43|See, I am standing beside this spring; if a maiden comes out to draw water and I say to her, "Please let me drink a little water from your jar,"
GEN|24|44|and if she says to me, "Drink, and I'll draw water for your camels too," let her be the one the LORD has chosen for my master's son.'
GEN|24|45|"Before I finished praying in my heart, Rebekah came out, with her jar on her shoulder. She went down to the spring and drew water, and I said to her, 'Please give me a drink.'
GEN|24|46|"She quickly lowered her jar from her shoulder and said, 'Drink, and I'll water your camels too.' So I drank, and she watered the camels also.
GEN|24|47|"I asked her, 'Whose daughter are you?'"She said, 'The daughter of Bethuel son of Nahor, whom Milcah bore to him.'"Then I put the ring in her nose and the bracelets on her arms,
GEN|24|48|and I bowed down and worshiped the LORD. I praised the LORD, the God of my master Abraham, who had led me on the right road to get the granddaughter of my master's brother for his son.
GEN|24|49|Now if you will show kindness and faithfulness to my master, tell me; and if not, tell me, so I may know which way to turn."
GEN|24|50|Laban and Bethuel answered, "This is from the LORD; we can say nothing to you one way or the other.
GEN|24|51|Here is Rebekah; take her and go, and let her become the wife of your master's son, as the LORD has directed."
GEN|24|52|When Abraham's servant heard what they said, he bowed down to the ground before the LORD.
GEN|24|53|Then the servant brought out gold and silver jewelry and articles of clothing and gave them to Rebekah; he also gave costly gifts to her brother and to her mother.
GEN|24|54|Then he and the men who were with him ate and drank and spent the night there. When they got up the next morning, he said, "Send me on my way to my master."
GEN|24|55|But her brother and her mother replied, "Let the girl remain with us ten days or so; then you may go."
GEN|24|56|But he said to them, "Do not detain me, now that the LORD has granted success to my journey. Send me on my way so I may go to my master."
GEN|24|57|Then they said, "Let's call the girl and ask her about it."
GEN|24|58|So they called Rebekah and asked her, "Will you go with this man?I will go," she said.
GEN|24|59|So they sent their sister Rebekah on her way, along with her nurse and Abraham's servant and his men.
GEN|24|60|And they blessed Rebekah and said to her, "Our sister, may you increase to thousands upon thousands; may your offspring possess the gates of their enemies."
GEN|24|61|Then Rebekah and her maids got ready and mounted their camels and went back with the man. So the servant took Rebekah and left.
GEN|24|62|Now Isaac had come from Beer Lahai Roi, for he was living in the Negev.
GEN|24|63|He went out to the field one evening to meditate, and as he looked up, he saw camels approaching.
GEN|24|64|Rebekah also looked up and saw Isaac. She got down from her camel
GEN|24|65|and asked the servant, "Who is that man in the field coming to meet us?He is my master," the servant answered. So she took her veil and covered herself.
GEN|24|66|Then the servant told Isaac all he had done.
GEN|24|67|Isaac brought her into the tent of his mother Sarah, and he married Rebekah. So she became his wife, and he loved her; and Isaac was comforted after his mother's death.
GEN|25|1|Abraham took another wife, whose name was Keturah.
GEN|25|2|She bore him Zimran, Jokshan, Medan, Midian, Ishbak and Shuah.
GEN|25|3|Jokshan was the father of Sheba and Dedan; the descendants of Dedan were the Asshurites, the Letushites and the Leummites.
GEN|25|4|The sons of Midian were Ephah, Epher, Hanoch, Abida and Eldaah. All these were descendants of Keturah.
GEN|25|5|Abraham left everything he owned to Isaac.
GEN|25|6|But while he was still living, he gave gifts to the sons of his concubines and sent them away from his son Isaac to the land of the east.
GEN|25|7|Altogether, Abraham lived a hundred and seventy-five years.
GEN|25|8|Then Abraham breathed his last and died at a good old age, an old man and full of years; and he was gathered to his people.
GEN|25|9|His sons Isaac and Ishmael buried him in the cave of Machpelah near Mamre, in the field of Ephron son of Zohar the Hittite,
GEN|25|10|the field Abraham had bought from the Hittites. There Abraham was buried with his wife Sarah.
GEN|25|11|After Abraham's death, God blessed his son Isaac, who then lived near Beer Lahai Roi.
GEN|25|12|This is the account of Abraham's son Ishmael, whom Sarah's maidservant, Hagar the Egyptian, bore to Abraham.
GEN|25|13|These are the names of the sons of Ishmael, listed in the order of their birth: Nebaioth the firstborn of Ishmael, Kedar, Adbeel, Mibsam,
GEN|25|14|Mishma, Dumah, Massa,
GEN|25|15|Hadad, Tema, Jetur, Naphish and Kedemah.
GEN|25|16|These were the sons of Ishmael, and these are the names of the twelve tribal rulers according to their settlements and camps.
GEN|25|17|Altogether, Ishmael lived a hundred and thirty-seven years. He breathed his last and died, and he was gathered to his people.
GEN|25|18|His descendants settled in the area from Havilah to Shur, near the border of Egypt, as you go toward Asshur. And they lived in hostility toward all their brothers.
GEN|25|19|This is the account of Abraham's son Isaac. Abraham became the father of Isaac,
GEN|25|20|and Isaac was forty years old when he married Rebekah daughter of Bethuel the Aramean from Paddan Aram and sister of Laban the Aramean.
GEN|25|21|Isaac prayed to the LORD on behalf of his wife, because she was barren. The LORD answered his prayer, and his wife Rebekah became pregnant.
GEN|25|22|The babies jostled each other within her, and she said, "Why is this happening to me?" So she went to inquire of the LORD.
GEN|25|23|The LORD said to her, "Two nations are in your womb, and two peoples from within you will be separated; one people will be stronger than the other, and the older will serve the younger."
GEN|25|24|When the time came for her to give birth, there were twin boys in her womb.
GEN|25|25|The first to come out was red, and his whole body was like a hairy garment; so they named him Esau.
GEN|25|26|After this, his brother came out, with his hand grasping Esau's heel; so he was named Jacob. Isaac was sixty years old when Rebekah gave birth to them.
GEN|25|27|The boys grew up, and Esau became a skillful hunter, a man of the open country, while Jacob was a quiet man, staying among the tents.
GEN|25|28|Isaac, who had a taste for wild game, loved Esau, but Rebekah loved Jacob.
GEN|25|29|Once when Jacob was cooking some stew, Esau came in from the open country, famished.
GEN|25|30|He said to Jacob, "Quick, let me have some of that red stew! I'm famished!" (That is why he was also called Edom. )
GEN|25|31|Jacob replied, "First sell me your birthright."
GEN|25|32|"Look, I am about to die," Esau said. "What good is the birthright to me?"
GEN|25|33|But Jacob said, "Swear to me first." So he swore an oath to him, selling his birthright to Jacob.
GEN|25|34|Then Jacob gave Esau some bread and some lentil stew. He ate and drank, and then got up and left. So Esau despised his birthright.
GEN|26|1|Now there was a famine in the land-besides the earlier famine of Abraham's time-and Isaac went to Abimelech king of the Philistines in Gerar.
GEN|26|2|The LORD appeared to Isaac and said, "Do not go down to Egypt; live in the land where I tell you to live.
GEN|26|3|Stay in this land for a while, and I will be with you and will bless you. For to you and your descendants I will give all these lands and will confirm the oath I swore to your father Abraham.
GEN|26|4|I will make your descendants as numerous as the stars in the sky and will give them all these lands, and through your offspring all nations on earth will be blessed,
GEN|26|5|because Abraham obeyed me and kept my requirements, my commands, my decrees and my laws."
GEN|26|6|So Isaac stayed in Gerar.
GEN|26|7|When the men of that place asked him about his wife, he said, "She is my sister," because he was afraid to say, "She is my wife." He thought, "The men of this place might kill me on account of Rebekah, because she is beautiful."
GEN|26|8|When Isaac had been there a long time, Abimelech king of the Philistines looked down from a window and saw Isaac caressing his wife Rebekah.
GEN|26|9|So Abimelech summoned Isaac and said, "She is really your wife! Why did you say, 'She is my sister'?" Isaac answered him, "Because I thought I might lose my life on account of her."
GEN|26|10|Then Abimelech said, "What is this you have done to us? One of the men might well have slept with your wife, and you would have brought guilt upon us."
GEN|26|11|So Abimelech gave orders to all the people: "Anyone who molests this man or his wife shall surely be put to death."
GEN|26|12|Isaac planted crops in that land and the same year reaped a hundredfold, because the LORD blessed him.
GEN|26|13|The man became rich, and his wealth continued to grow until he became very wealthy.
GEN|26|14|He had so many flocks and herds and servants that the Philistines envied him.
GEN|26|15|So all the wells that his father's servants had dug in the time of his father Abraham, the Philistines stopped up, filling them with earth.
GEN|26|16|Then Abimelech said to Isaac, "Move away from us; you have become too powerful for us."
GEN|26|17|So Isaac moved away from there and encamped in the Valley of Gerar and settled there.
GEN|26|18|Isaac reopened the wells that had been dug in the time of his father Abraham, which the Philistines had stopped up after Abraham died, and he gave them the same names his father had given them.
GEN|26|19|Isaac's servants dug in the valley and discovered a well of fresh water there.
GEN|26|20|But the herdsmen of Gerar quarreled with Isaac's herdsmen and said, "The water is ours!" So he named the well Esek, because they disputed with him.
GEN|26|21|Then they dug another well, but they quarreled over that one also; so he named it Sitnah.
GEN|26|22|He moved on from there and dug another well, and no one quarreled over it. He named it Rehoboth, saying, "Now the LORD has given us room and we will flourish in the land."
GEN|26|23|From there he went up to Beersheba.
GEN|26|24|That night the LORD appeared to him and said, "I am the God of your father Abraham. Do not be afraid, for I am with you; I will bless you and will increase the number of your descendants for the sake of my servant Abraham."
GEN|26|25|Isaac built an altar there and called on the name of the LORD. There he pitched his tent, and there his servants dug a well.
GEN|26|26|Meanwhile, Abimelech had come to him from Gerar, with Ahuzzath his personal adviser and Phicol the commander of his forces.
GEN|26|27|Isaac asked them, "Why have you come to me, since you were hostile to me and sent me away?"
GEN|26|28|They answered, "We saw clearly that the LORD was with you; so we said, 'There ought to be a sworn agreement between us'-between us and you. Let us make a treaty with you
GEN|26|29|that you will do us no harm, just as we did not molest you but always treated you well and sent you away in peace. And now you are blessed by the LORD."
GEN|26|30|Isaac then made a feast for them, and they ate and drank.
GEN|26|31|Early the next morning the men swore an oath to each other. Then Isaac sent them on their way, and they left him in peace.
GEN|26|32|That day Isaac's servants came and told him about the well they had dug. They said, "We've found water!"
GEN|26|33|He called it Shibah, and to this day the name of the town has been Beersheba.
GEN|26|34|When Esau was forty years old, he married Judith daughter of Beeri the Hittite, and also Basemath daughter of Elon the Hittite.
GEN|26|35|They were a source of grief to Isaac and Rebekah.
GEN|27|1|When Isaac was old and his eyes were so weak that he could no longer see, he called for Esau his older son and said to him, "My son.Here I am," he answered.
GEN|27|2|Isaac said, "I am now an old man and don't know the day of my death.
GEN|27|3|Now then, get your weapons-your quiver and bow-and go out to the open country to hunt some wild game for me.
GEN|27|4|Prepare me the kind of tasty food I like and bring it to me to eat, so that I may give you my blessing before I die."
GEN|27|5|Now Rebekah was listening as Isaac spoke to his son Esau. When Esau left for the open country to hunt game and bring it back,
GEN|27|6|Rebekah said to her son Jacob, "Look, I overheard your father say to your brother Esau,
GEN|27|7|'Bring me some game and prepare me some tasty food to eat, so that I may give you my blessing in the presence of the LORD before I die.'
GEN|27|8|Now, my son, listen carefully and do what I tell you:
GEN|27|9|Go out to the flock and bring me two choice young goats, so I can prepare some tasty food for your father, just the way he likes it.
GEN|27|10|Then take it to your father to eat, so that he may give you his blessing before he dies."
GEN|27|11|Jacob said to Rebekah his mother, "But my brother Esau is a hairy man, and I'm a man with smooth skin.
GEN|27|12|What if my father touches me? I would appear to be tricking him and would bring down a curse on myself rather than a blessing."
GEN|27|13|His mother said to him, "My son, let the curse fall on me. Just do what I say; go and get them for me."
GEN|27|14|So he went and got them and brought them to his mother, and she prepared some tasty food, just the way his father liked it.
GEN|27|15|Then Rebekah took the best clothes of Esau her older son, which she had in the house, and put them on her younger son Jacob.
GEN|27|16|She also covered his hands and the smooth part of his neck with the goatskins.
GEN|27|17|Then she handed to her son Jacob the tasty food and the bread she had made.
GEN|27|18|He went to his father and said, "My father.Yes, my son," he answered. "Who is it?"
GEN|27|19|Jacob said to his father, "I am Esau your firstborn. I have done as you told me. Please sit up and eat some of my game so that you may give me your blessing."
GEN|27|20|Isaac asked his son, "How did you find it so quickly, my son?The LORD your God gave me success," he replied.
GEN|27|21|Then Isaac said to Jacob, "Come near so I can touch you, my son, to know whether you really are my son Esau or not."
GEN|27|22|Jacob went close to his father Isaac, who touched him and said, "The voice is the voice of Jacob, but the hands are the hands of Esau."
GEN|27|23|He did not recognize him, for his hands were hairy like those of his brother Esau; so he blessed him.
GEN|27|24|"Are you really my son Esau?" he asked. "I am," he replied.
GEN|27|25|Then he said, "My son, bring me some of your game to eat, so that I may give you my blessing." Jacob brought it to him and he ate; and he brought some wine and he drank.
GEN|27|26|Then his father Isaac said to him, "Come here, my son, and kiss me."
GEN|27|27|So he went to him and kissed him. When Isaac caught the smell of his clothes, he blessed him and said, "Ah, the smell of my son is like the smell of a field that the LORD has blessed.
GEN|27|28|May God give you of heaven's dew and of earth's richness- an abundance of grain and new wine.
GEN|27|29|May nations serve you and peoples bow down to you. Be lord over your brothers, and may the sons of your mother bow down to you. May those who curse you be cursed and those who bless you be blessed."
GEN|27|30|After Isaac finished blessing him and Jacob had scarcely left his father's presence, his brother Esau came in from hunting.
GEN|27|31|He too prepared some tasty food and brought it to his father. Then he said to him, "My father, sit up and eat some of my game, so that you may give me your blessing."
GEN|27|32|His father Isaac asked him, "Who are you?I am your son," he answered, "your firstborn, Esau."
GEN|27|33|Isaac trembled violently and said, "Who was it, then, that hunted game and brought it to me? I ate it just before you came and I blessed him-and indeed he will be blessed!"
GEN|27|34|When Esau heard his father's words, he burst out with a loud and bitter cry and said to his father, "Bless me-me too, my father!"
GEN|27|35|But he said, "Your brother came deceitfully and took your blessing."
GEN|27|36|Esau said, "Isn't he rightly named Jacob? He has deceived me these two times: He took my birthright, and now he's taken my blessing!" Then he asked, "Haven't you reserved any blessing for me?"
GEN|27|37|Isaac answered Esau, "I have made him lord over you and have made all his relatives his servants, and I have sustained him with grain and new wine. So what can I possibly do for you, my son?"
GEN|27|38|Esau said to his father, "Do you have only one blessing, my father? Bless me too, my father!" Then Esau wept aloud.
GEN|27|39|His father Isaac answered him, "Your dwelling will be away from the earth's richness, away from the dew of heaven above.
GEN|27|40|You will live by the sword and you will serve your brother. But when you grow restless, you will throw his yoke from off your neck."
GEN|27|41|Esau held a grudge against Jacob because of the blessing his father had given him. He said to himself, "The days of mourning for my father are near; then I will kill my brother Jacob."
GEN|27|42|When Rebekah was told what her older son Esau had said, she sent for her younger son Jacob and said to him, "Your brother Esau is consoling himself with the thought of killing you.
GEN|27|43|Now then, my son, do what I say: Flee at once to my brother Laban in Haran.
GEN|27|44|Stay with him for a while until your brother's fury subsides.
GEN|27|45|When your brother is no longer angry with you and forgets what you did to him, I'll send word for you to come back from there. Why should I lose both of you in one day?"
GEN|27|46|Then Rebekah said to Isaac, "I'm disgusted with living because of these Hittite women. If Jacob takes a wife from among the women of this land, from Hittite women like these, my life will not be worth living."
GEN|28|1|So Isaac called for Jacob and blessed him and commanded him: "Do not marry a Canaanite woman.
GEN|28|2|Go at once to Paddan Aram, to the house of your mother's father Bethuel. Take a wife for yourself there, from among the daughters of Laban, your mother's brother.
GEN|28|3|May God Almighty bless you and make you fruitful and increase your numbers until you become a community of peoples.
GEN|28|4|May he give you and your descendants the blessing given to Abraham, so that you may take possession of the land where you now live as an alien, the land God gave to Abraham."
GEN|28|5|Then Isaac sent Jacob on his way, and he went to Paddan Aram, to Laban son of Bethuel the Aramean, the brother of Rebekah, who was the mother of Jacob and Esau.
GEN|28|6|Now Esau learned that Isaac had blessed Jacob and had sent him to Paddan Aram to take a wife from there, and that when he blessed him he commanded him, "Do not marry a Canaanite woman,"
GEN|28|7|and that Jacob had obeyed his father and mother and had gone to Paddan Aram.
GEN|28|8|Esau then realized how displeasing the Canaanite women were to his father Isaac;
GEN|28|9|so he went to Ishmael and married Mahalath, the sister of Nebaioth and daughter of Ishmael son of Abraham, in addition to the wives he already had.
GEN|28|10|Jacob left Beersheba and set out for Haran.
GEN|28|11|When he reached a certain place, he stopped for the night because the sun had set. Taking one of the stones there, he put it under his head and lay down to sleep.
GEN|28|12|He had a dream in which he saw a stairway resting on the earth, with its top reaching to heaven, and the angels of God were ascending and descending on it.
GEN|28|13|There above it stood the LORD, and he said: "I am the LORD, the God of your father Abraham and the God of Isaac. I will give you and your descendants the land on which you are lying.
GEN|28|14|Your descendants will be like the dust of the earth, and you will spread out to the west and to the east, to the north and to the south. All peoples on earth will be blessed through you and your offspring.
GEN|28|15|I am with you and will watch over you wherever you go, and I will bring you back to this land. I will not leave you until I have done what I have promised you."
GEN|28|16|When Jacob awoke from his sleep, he thought, "Surely the LORD is in this place, and I was not aware of it."
GEN|28|17|He was afraid and said, "How awesome is this place! This is none other than the house of God; this is the gate of heaven."
GEN|28|18|Early the next morning Jacob took the stone he had placed under his head and set it up as a pillar and poured oil on top of it.
GEN|28|19|He called that place Bethel, though the city used to be called Luz.
GEN|28|20|Then Jacob made a vow, saying, "If God will be with me and will watch over me on this journey I am taking and will give me food to eat and clothes to wear
GEN|28|21|so that I return safely to my father's house, then the LORD will be my God
GEN|28|22|and this stone that I have set up as a pillar will be God's house, and of all that you give me I will give you a tenth."
GEN|29|1|Then Jacob continued on his journey and came to the land of the eastern peoples.
GEN|29|2|There he saw a well in the field, with three flocks of sheep lying near it because the flocks were watered from that well. The stone over the mouth of the well was large.
GEN|29|3|When all the flocks were gathered there, the shepherds would roll the stone away from the well's mouth and water the sheep. Then they would return the stone to its place over the mouth of the well.
GEN|29|4|Jacob asked the shepherds, "My brothers, where are you from?We're from Haran," they replied.
GEN|29|5|He said to them, "Do you know Laban, Nahor's grandson?Yes, we know him," they answered.
GEN|29|6|Then Jacob asked them, "Is he well?Yes, he is," they said, "and here comes his daughter Rachel with the sheep."
GEN|29|7|"Look," he said, "the sun is still high; it is not time for the flocks to be gathered. Water the sheep and take them back to pasture."
GEN|29|8|"We can't," they replied, "until all the flocks are gathered and the stone has been rolled away from the mouth of the well. Then we will water the sheep."
GEN|29|9|While he was still talking with them, Rachel came with her father's sheep, for she was a shepherdess.
GEN|29|10|When Jacob saw Rachel daughter of Laban, his mother's brother, and Laban's sheep, he went over and rolled the stone away from the mouth of the well and watered his uncle's sheep.
GEN|29|11|Then Jacob kissed Rachel and began to weep aloud.
GEN|29|12|He had told Rachel that he was a relative of her father and a son of Rebekah. So she ran and told her father.
GEN|29|13|As soon as Laban heard the news about Jacob, his sister's son, he hurried to meet him. He embraced him and kissed him and brought him to his home, and there Jacob told him all these things.
GEN|29|14|Then Laban said to him, "You are my own flesh and blood." After Jacob had stayed with him for a whole month,
GEN|29|15|Laban said to him, "Just because you are a relative of mine, should you work for me for nothing? Tell me what your wages should be."
GEN|29|16|Now Laban had two daughters; the name of the older was Leah, and the name of the younger was Rachel.
GEN|29|17|Leah had weak eyes, but Rachel was lovely in form, and beautiful.
GEN|29|18|Jacob was in love with Rachel and said, "I'll work for you seven years in return for your younger daughter Rachel."
GEN|29|19|Laban said, "It's better that I give her to you than to some other man. Stay here with me."
GEN|29|20|So Jacob served seven years to get Rachel, but they seemed like only a few days to him because of his love for her.
GEN|29|21|Then Jacob said to Laban, "Give me my wife. My time is completed, and I want to lie with her."
GEN|29|22|So Laban brought together all the people of the place and gave a feast.
GEN|29|23|But when evening came, he took his daughter Leah and gave her to Jacob, and Jacob lay with her.
GEN|29|24|And Laban gave his servant girl Zilpah to his daughter as her maidservant.
GEN|29|25|When morning came, there was Leah! So Jacob said to Laban, "What is this you have done to me? I served you for Rachel, didn't I? Why have you deceived me?"
GEN|29|26|Laban replied, "It is not our custom here to give the younger daughter in marriage before the older one.
GEN|29|27|Finish this daughter's bridal week; then we will give you the younger one also, in return for another seven years of work."
GEN|29|28|And Jacob did so. He finished the week with Leah, and then Laban gave him his daughter Rachel to be his wife.
GEN|29|29|Laban gave his servant girl Bilhah to his daughter Rachel as her maidservant.
GEN|29|30|Jacob lay with Rachel also, and he loved Rachel more than Leah. And he worked for Laban another seven years.
GEN|29|31|When the LORD saw that Leah was not loved, he opened her womb, but Rachel was barren.
GEN|29|32|Leah became pregnant and gave birth to a son. She named him Reuben, for she said, "It is because the LORD has seen my misery. Surely my husband will love me now."
GEN|29|33|She conceived again, and when she gave birth to a son she said, "Because the LORD heard that I am not loved, he gave me this one too." So she named him Simeon.
GEN|29|34|Again she conceived, and when she gave birth to a son she said, "Now at last my husband will become attached to me, because I have borne him three sons." So he was named Levi.
GEN|29|35|She conceived again, and when she gave birth to a son she said, "This time I will praise the LORD." So she named him Judah. Then she stopped having children.
GEN|30|1|When Rachel saw that she was not bearing Jacob any children, she became jealous of her sister. So she said to Jacob, "Give me children, or I'll die!"
GEN|30|2|Jacob became angry with her and said, "Am I in the place of God, who has kept you from having children?"
GEN|30|3|Then she said, "Here is Bilhah, my maidservant. Sleep with her so that she can bear children for me and that through her I too can build a family."
GEN|30|4|So she gave him her servant Bilhah as a wife. Jacob slept with her,
GEN|30|5|and she became pregnant and bore him a son.
GEN|30|6|Then Rachel said, "God has vindicated me; he has listened to my plea and given me a son." Because of this she named him Dan.
GEN|30|7|Rachel's servant Bilhah conceived again and bore Jacob a second son.
GEN|30|8|Then Rachel said, "I have had a great struggle with my sister, and I have won." So she named him Naphtali.
GEN|30|9|When Leah saw that she had stopped having children, she took her maidservant Zilpah and gave her to Jacob as a wife.
GEN|30|10|Leah's servant Zilpah bore Jacob a son.
GEN|30|11|Then Leah said, "What good fortune!" So she named him Gad.
GEN|30|12|Leah's servant Zilpah bore Jacob a second son.
GEN|30|13|Then Leah said, "How happy I am! The women will call me happy." So she named him Asher.
GEN|30|14|During wheat harvest, Reuben went out into the fields and found some mandrake plants, which he brought to his mother Leah. Rachel said to Leah, "Please give me some of your son's mandrakes."
GEN|30|15|But she said to her, "Wasn't it enough that you took away my husband? Will you take my son's mandrakes too?Very well," Rachel said, "he can sleep with you tonight in return for your son's mandrakes."
GEN|30|16|So when Jacob came in from the fields that evening, Leah went out to meet him. "You must sleep with me," she said. "I have hired you with my son's mandrakes." So he slept with her that night.
GEN|30|17|God listened to Leah, and she became pregnant and bore Jacob a fifth son.
GEN|30|18|Then Leah said, "God has rewarded me for giving my maidservant to my husband." So she named him Issachar.
GEN|30|19|Leah conceived again and bore Jacob a sixth son.
GEN|30|20|Then Leah said, "God has presented me with a precious gift. This time my husband will treat me with honor, because I have borne him six sons." So she named him Zebulun.
GEN|30|21|Some time later she gave birth to a daughter and named her Dinah.
GEN|30|22|Then God remembered Rachel; he listened to her and opened her womb.
GEN|30|23|She became pregnant and gave birth to a son and said, "God has taken away my disgrace."
GEN|30|24|She named him Joseph, and said, "May the LORD add to me another son."
GEN|30|25|After Rachel gave birth to Joseph, Jacob said to Laban, "Send me on my way so I can go back to my own homeland.
GEN|30|26|Give me my wives and children, for whom I have served you, and I will be on my way. You know how much work I've done for you."
GEN|30|27|But Laban said to him, "If I have found favor in your eyes, please stay. I have learned by divination that the LORD has blessed me because of you."
GEN|30|28|He added, "Name your wages, and I will pay them."
GEN|30|29|Jacob said to him, "You know how I have worked for you and how your livestock has fared under my care.
GEN|30|30|The little you had before I came has increased greatly, and the LORD has blessed you wherever I have been. But now, when may I do something for my own household?"
GEN|30|31|"What shall I give you?" he asked. "Don't give me anything," Jacob replied. "But if you will do this one thing for me, I will go on tending your flocks and watching over them:
GEN|30|32|Let me go through all your flocks today and remove from them every speckled or spotted sheep, every dark-colored lamb and every spotted or speckled goat. They will be my wages.
GEN|30|33|And my honesty will testify for me in the future, whenever you check on the wages you have paid me. Any goat in my possession that is not speckled or spotted, or any lamb that is not dark-colored, will be considered stolen."
GEN|30|34|"Agreed," said Laban. "Let it be as you have said."
GEN|30|35|That same day he removed all the male goats that were streaked or spotted, and all the speckled or spotted female goats (all that had white on them) and all the dark-colored lambs, and he placed them in the care of his sons.
GEN|30|36|Then he put a three-day journey between himself and Jacob, while Jacob continued to tend the rest of Laban's flocks.
GEN|30|37|Jacob, however, took fresh-cut branches from poplar, almond and plane trees and made white stripes on them by peeling the bark and exposing the white inner wood of the branches.
GEN|30|38|Then he placed the peeled branches in all the watering troughs, so that they would be directly in front of the flocks when they came to drink. When the flocks were in heat and came to drink,
GEN|30|39|they mated in front of the branches. And they bore young that were streaked or speckled or spotted.
GEN|30|40|Jacob set apart the young of the flock by themselves, but made the rest face the streaked and dark-colored animals that belonged to Laban. Thus he made separate flocks for himself and did not put them with Laban's animals.
GEN|30|41|Whenever the stronger females were in heat, Jacob would place the branches in the troughs in front of the animals so they would mate near the branches,
GEN|30|42|but if the animals were weak, he would not place them there. So the weak animals went to Laban and the strong ones to Jacob.
GEN|30|43|In this way the man grew exceedingly prosperous and came to own large flocks, and maidservants and menservants, and camels and donkeys.
GEN|31|1|Jacob heard that Laban's sons were saying, "Jacob has taken everything our father owned and has gained all this wealth from what belonged to our father."
GEN|31|2|And Jacob noticed that Laban's attitude toward him was not what it had been.
GEN|31|3|Then the LORD said to Jacob, "Go back to the land of your fathers and to your relatives, and I will be with you."
GEN|31|4|So Jacob sent word to Rachel and Leah to come out to the fields where his flocks were.
GEN|31|5|He said to them, "I see that your father's attitude toward me is not what it was before, but the God of my father has been with me.
GEN|31|6|You know that I've worked for your father with all my strength,
GEN|31|7|yet your father has cheated me by changing my wages ten times. However, God has not allowed him to harm me.
GEN|31|8|If he said, 'The speckled ones will be your wages,' then all the flocks gave birth to speckled young; and if he said, 'The streaked ones will be your wages,' then all the flocks bore streaked young.
GEN|31|9|So God has taken away your father's livestock and has given them to me.
GEN|31|10|"In breeding season I once had a dream in which I looked up and saw that the male goats mating with the flock were streaked, speckled or spotted.
GEN|31|11|The angel of God said to me in the dream, 'Jacob.' I answered, 'Here I am.'
GEN|31|12|And he said, 'Look up and see that all the male goats mating with the flock are streaked, speckled or spotted, for I have seen all that Laban has been doing to you.
GEN|31|13|I am the God of Bethel, where you anointed a pillar and where you made a vow to me. Now leave this land at once and go back to your native land.'"
GEN|31|14|Then Rachel and Leah replied, "Do we still have any share in the inheritance of our father's estate?
GEN|31|15|Does he not regard us as foreigners? Not only has he sold us, but he has used up what was paid for us.
GEN|31|16|Surely all the wealth that God took away from our father belongs to us and our children. So do whatever God has told you."
GEN|31|17|Then Jacob put his children and his wives on camels,
GEN|31|18|and he drove all his livestock ahead of him, along with all the goods he had accumulated in Paddan Aram, to go to his father Isaac in the land of Canaan.
GEN|31|19|When Laban had gone to shear his sheep, Rachel stole her father's household gods.
GEN|31|20|Moreover, Jacob deceived Laban the Aramean by not telling him he was running away.
GEN|31|21|So he fled with all he had, and crossing the River, he headed for the hill country of Gilead.
GEN|31|22|On the third day Laban was told that Jacob had fled.
GEN|31|23|Taking his relatives with him, he pursued Jacob for seven days and caught up with him in the hill country of Gilead.
GEN|31|24|Then God came to Laban the Aramean in a dream at night and said to him, "Be careful not to say anything to Jacob, either good or bad."
GEN|31|25|Jacob had pitched his tent in the hill country of Gilead when Laban overtook him, and Laban and his relatives camped there too.
GEN|31|26|Then Laban said to Jacob, "What have you done? You've deceived me, and you've carried off my daughters like captives in war.
GEN|31|27|Why did you run off secretly and deceive me? Why didn't you tell me, so I could send you away with joy and singing to the music of tambourines and harps?
GEN|31|28|You didn't even let me kiss my grandchildren and my daughters good-by. You have done a foolish thing.
GEN|31|29|I have the power to harm you; but last night the God of your father said to me, 'Be careful not to say anything to Jacob, either good or bad.'
GEN|31|30|Now you have gone off because you longed to return to your father's house. But why did you steal my gods?"
GEN|31|31|Jacob answered Laban, "I was afraid, because I thought you would take your daughters away from me by force.
GEN|31|32|But if you find anyone who has your gods, he shall not live. In the presence of our relatives, see for yourself whether there is anything of yours here with me; and if so, take it." Now Jacob did not know that Rachel had stolen the gods.
GEN|31|33|So Laban went into Jacob's tent and into Leah's tent and into the tent of the two maidservants, but he found nothing. After he came out of Leah's tent, he entered Rachel's tent.
GEN|31|34|Now Rachel had taken the household gods and put them inside her camel's saddle and was sitting on them. Laban searched through everything in the tent but found nothing.
GEN|31|35|Rachel said to her father, "Don't be angry, my lord, that I cannot stand up in your presence; I'm having my period." So he searched but could not find the household gods.
GEN|31|36|Jacob was angry and took Laban to task. "What is my crime?" he asked Laban. "What sin have I committed that you hunt me down?
GEN|31|37|Now that you have searched through all my goods, what have you found that belongs to your household? Put it here in front of your relatives and mine, and let them judge between the two of us.
GEN|31|38|"I have been with you for twenty years now. Your sheep and goats have not miscarried, nor have I eaten rams from your flocks.
GEN|31|39|I did not bring you animals torn by wild beasts; I bore the loss myself. And you demanded payment from me for whatever was stolen by day or night.
GEN|31|40|This was my situation: The heat consumed me in the daytime and the cold at night, and sleep fled from my eyes.
GEN|31|41|It was like this for the twenty years I was in your household. I worked for you fourteen years for your two daughters and six years for your flocks, and you changed my wages ten times.
GEN|31|42|If the God of my father, the God of Abraham and the Fear of Isaac, had not been with me, you would surely have sent me away empty-handed. But God has seen my hardship and the toil of my hands, and last night he rebuked you."
GEN|31|43|Laban answered Jacob, "The women are my daughters, the children are my children, and the flocks are my flocks. All you see is mine. Yet what can I do today about these daughters of mine, or about the children they have borne?
GEN|31|44|Come now, let's make a covenant, you and I, and let it serve as a witness between us."
GEN|31|45|So Jacob took a stone and set it up as a pillar.
GEN|31|46|He said to his relatives, "Gather some stones." So they took stones and piled them in a heap, and they ate there by the heap.
GEN|31|47|Laban called it Jegar Sahadutha, and Jacob called it Galeed.
GEN|31|48|Laban said, "This heap is a witness between you and me today." That is why it was called Galeed.
GEN|31|49|It was also called Mizpah, because he said, "May the LORD keep watch between you and me when we are away from each other.
GEN|31|50|If you mistreat my daughters or if you take any wives besides my daughters, even though no one is with us, remember that God is a witness between you and me."
GEN|31|51|Laban also said to Jacob, "Here is this heap, and here is this pillar I have set up between you and me.
GEN|31|52|This heap is a witness, and this pillar is a witness, that I will not go past this heap to your side to harm you and that you will not go past this heap and pillar to my side to harm me.
GEN|31|53|May the God of Abraham and the God of Nahor, the God of their father, judge between us." So Jacob took an oath in the name of the Fear of his father Isaac.
GEN|31|54|He offered a sacrifice there in the hill country and invited his relatives to a meal. After they had eaten, they spent the night there.
GEN|31|55|Early the next morning Laban kissed his grandchildren and his daughters and blessed them. Then he left and returned home.
GEN|32|1|Jacob also went on his way, and the angels of God met him.
GEN|32|2|When Jacob saw them, he said, "This is the camp of God!" So he named that place Mahanaim.
GEN|32|3|Jacob sent messengers ahead of him to his brother Esau in the land of Seir, the country of Edom.
GEN|32|4|He instructed them: "This is what you are to say to my master Esau: 'Your servant Jacob says, I have been staying with Laban and have remained there till now.
GEN|32|5|I have cattle and donkeys, sheep and goats, menservants and maidservants. Now I am sending this message to my lord, that I may find favor in your eyes.'"
GEN|32|6|When the messengers returned to Jacob, they said, "We went to your brother Esau, and now he is coming to meet you, and four hundred men are with him."
GEN|32|7|In great fear and distress Jacob divided the people who were with him into two groups, and the flocks and herds and camels as well.
GEN|32|8|He thought, "If Esau comes and attacks one group, the group that is left may escape."
GEN|32|9|Then Jacob prayed, "O God of my father Abraham, God of my father Isaac, O LORD, who said to me, 'Go back to your country and your relatives, and I will make you prosper,'
GEN|32|10|I am unworthy of all the kindness and faithfulness you have shown your servant. I had only my staff when I crossed this Jordan, but now I have become two groups.
GEN|32|11|Save me, I pray, from the hand of my brother Esau, for I am afraid he will come and attack me, and also the mothers with their children.
GEN|32|12|But you have said, 'I will surely make you prosper and will make your descendants like the sand of the sea, which cannot be counted.'"
GEN|32|13|He spent the night there, and from what he had with him he selected a gift for his brother Esau:
GEN|32|14|two hundred female goats and twenty male goats, two hundred ewes and twenty rams,
GEN|32|15|thirty female camels with their young, forty cows and ten bulls, and twenty female donkeys and ten male donkeys.
GEN|32|16|He put them in the care of his servants, each herd by itself, and said to his servants, "Go ahead of me, and keep some space between the herds."
GEN|32|17|He instructed the one in the lead: "When my brother Esau meets you and asks, 'To whom do you belong, and where are you going, and who owns all these animals in front of you?'
GEN|32|18|then you are to say, 'They belong to your servant Jacob. They are a gift sent to my lord Esau, and he is coming behind us.'"
GEN|32|19|He also instructed the second, the third and all the others who followed the herds: "You are to say the same thing to Esau when you meet him.
GEN|32|20|And be sure to say, 'Your servant Jacob is coming behind us.'" For he thought, "I will pacify him with these gifts I am sending on ahead; later, when I see him, perhaps he will receive me."
GEN|32|21|So Jacob's gifts went on ahead of him, but he himself spent the night in the camp.
GEN|32|22|That night Jacob got up and took his two wives, his two maidservants and his eleven sons and crossed the ford of the Jabbok.
GEN|32|23|After he had sent them across the stream, he sent over all his possessions.
GEN|32|24|So Jacob was left alone, and a man wrestled with him till daybreak.
GEN|32|25|When the man saw that he could not overpower him, he touched the socket of Jacob's hip so that his hip was wrenched as he wrestled with the man.
GEN|32|26|Then the man said, "Let me go, for it is daybreak." But Jacob replied, "I will not let you go unless you bless me."
GEN|32|27|The man asked him, "What is your name?Jacob," he answered.
GEN|32|28|Then the man said, "Your name will no longer be Jacob, but Israel, because you have struggled with God and with men and have overcome."
GEN|32|29|Jacob said, "Please tell me your name." But he replied, "Why do you ask my name?" Then he blessed him there.
GEN|32|30|So Jacob called the place Peniel, saying, "It is because I saw God face to face, and yet my life was spared."
GEN|32|31|The sun rose above him as he passed Peniel, and he was limping because of his hip.
GEN|32|32|Therefore to this day the Israelites do not eat the tendon attached to the socket of the hip, because the socket of Jacob's hip was touched near the tendon.
GEN|33|1|Jacob looked up and there was Esau, coming with his four hundred men; so he divided the children among Leah, Rachel and the two maidservants.
GEN|33|2|He put the maidservants and their children in front, Leah and her children next, and Rachel and Joseph in the rear.
GEN|33|3|He himself went on ahead and bowed down to the ground seven times as he approached his brother.
GEN|33|4|But Esau ran to meet Jacob and embraced him; he threw his arms around his neck and kissed him. And they wept.
GEN|33|5|Then Esau looked up and saw the women and children. "Who are these with you?" he asked. Jacob answered, "They are the children God has graciously given your servant."
GEN|33|6|Then the maidservants and their children approached and bowed down.
GEN|33|7|Next, Leah and her children came and bowed down. Last of all came Joseph and Rachel, and they too bowed down.
GEN|33|8|Esau asked, "What do you mean by all these droves I met?To find favor in your eyes, my lord," he said.
GEN|33|9|But Esau said, "I already have plenty, my brother. Keep what you have for yourself."
GEN|33|10|"No, please!" said Jacob. "If I have found favor in your eyes, accept this gift from me. For to see your face is like seeing the face of God, now that you have received me favorably.
GEN|33|11|Please accept the present that was brought to you, for God has been gracious to me and I have all I need." And because Jacob insisted, Esau accepted it.
GEN|33|12|Then Esau said, "Let us be on our way; I'll accompany you."
GEN|33|13|But Jacob said to him, "My lord knows that the children are tender and that I must care for the ewes and cows that are nursing their young. If they are driven hard just one day, all the animals will die.
GEN|33|14|So let my lord go on ahead of his servant, while I move along slowly at the pace of the droves before me and that of the children, until I come to my lord in Seir."
GEN|33|15|Esau said, "Then let me leave some of my men with you.But why do that?" Jacob asked. "Just let me find favor in the eyes of my lord."
GEN|33|16|So that day Esau started on his way back to Seir.
GEN|33|17|Jacob, however, went to Succoth, where he built a place for himself and made shelters for his livestock. That is why the place is called Succoth.
GEN|33|18|After Jacob came from Paddan Aram, he arrived safely at the city of Shechem in Canaan and camped within sight of the city.
GEN|33|19|For a hundred pieces of silver, he bought from the sons of Hamor, the father of Shechem, the plot of ground where he pitched his tent.
GEN|33|20|There he set up an altar and called it El Elohe Israel.
GEN|34|1|Now Dinah, the daughter Leah had borne to Jacob, went out to visit the women of the land.
GEN|34|2|When Shechem son of Hamor the Hivite, the ruler of that area, saw her, he took her and violated her.
GEN|34|3|His heart was drawn to Dinah daughter of Jacob, and he loved the girl and spoke tenderly to her.
GEN|34|4|And Shechem said to his father Hamor, "Get me this girl as my wife."
GEN|34|5|When Jacob heard that his daughter Dinah had been defiled, his sons were in the fields with his livestock; so he kept quiet about it until they came home.
GEN|34|6|Then Shechem's father Hamor went out to talk with Jacob.
GEN|34|7|Now Jacob's sons had come in from the fields as soon as they heard what had happened. They were filled with grief and fury, because Shechem had done a disgraceful thing in Israel by lying with Jacob's daughter-a thing that should not be done.
GEN|34|8|But Hamor said to them, "My son Shechem has his heart set on your daughter. Please give her to him as his wife.
GEN|34|9|Intermarry with us; give us your daughters and take our daughters for yourselves.
GEN|34|10|You can settle among us; the land is open to you. Live in it, trade in it, and acquire property in it."
GEN|34|11|Then Shechem said to Dinah's father and brothers, "Let me find favor in your eyes, and I will give you whatever you ask.
GEN|34|12|Make the price for the bride and the gift I am to bring as great as you like, and I'll pay whatever you ask me. Only give me the girl as my wife."
GEN|34|13|Because their sister Dinah had been defiled, Jacob's sons replied deceitfully as they spoke to Shechem and his father Hamor.
GEN|34|14|They said to them, "We can't do such a thing; we can't give our sister to a man who is not circumcised. That would be a disgrace to us.
GEN|34|15|We will give our consent to you on one condition only: that you become like us by circumcising all your males.
GEN|34|16|Then we will give you our daughters and take your daughters for ourselves. We'll settle among you and become one people with you.
GEN|34|17|But if you will not agree to be circumcised, we'll take our sister and go."
GEN|34|18|Their proposal seemed good to Hamor and his son Shechem.
GEN|34|19|The young man, who was the most honored of all his father's household, lost no time in doing what they said, because he was delighted with Jacob's daughter.
GEN|34|20|So Hamor and his son Shechem went to the gate of their city to speak to their fellow townsmen.
GEN|34|21|"These men are friendly toward us," they said. "Let them live in our land and trade in it; the land has plenty of room for them. We can marry their daughters and they can marry ours.
GEN|34|22|But the men will consent to live with us as one people only on the condition that our males be circumcised, as they themselves are.
GEN|34|23|Won't their livestock, their property and all their other animals become ours? So let us give our consent to them, and they will settle among us."
GEN|34|24|All the men who went out of the city gate agreed with Hamor and his son Shechem, and every male in the city was circumcised.
GEN|34|25|Three days later, while all of them were still in pain, two of Jacob's sons, Simeon and Levi, Dinah's brothers, took their swords and attacked the unsuspecting city, killing every male.
GEN|34|26|They put Hamor and his son Shechem to the sword and took Dinah from Shechem's house and left.
GEN|34|27|The sons of Jacob came upon the dead bodies and looted the city where their sister had been defiled.
GEN|34|28|They seized their flocks and herds and donkeys and everything else of theirs in the city and out in the fields.
GEN|34|29|They carried off all their wealth and all their women and children, taking as plunder everything in the houses.
GEN|34|30|Then Jacob said to Simeon and Levi, "You have brought trouble on me by making me a stench to the Canaanites and Perizzites, the people living in this land. We are few in number, and if they join forces against me and attack me, I and my household will be destroyed."
GEN|34|31|But they replied, "Should he have treated our sister like a prostitute?"
GEN|35|1|Then God said to Jacob, "Go up to Bethel and settle there, and build an altar there to God, who appeared to you when you were fleeing from your brother Esau."
GEN|35|2|So Jacob said to his household and to all who were with him, "Get rid of the foreign gods you have with you, and purify yourselves and change your clothes.
GEN|35|3|Then come, let us go up to Bethel, where I will build an altar to God, who answered me in the day of my distress and who has been with me wherever I have gone."
GEN|35|4|So they gave Jacob all the foreign gods they had and the rings in their ears, and Jacob buried them under the oak at Shechem.
GEN|35|5|Then they set out, and the terror of God fell upon the towns all around them so that no one pursued them.
GEN|35|6|Jacob and all the people with him came to Luz (that is, Bethel) in the land of Canaan.
GEN|35|7|There he built an altar, and he called the place El Bethel, because it was there that God revealed himself to him when he was fleeing from his brother.
GEN|35|8|Now Deborah, Rebekah's nurse, died and was buried under the oak below Bethel. So it was named Allon Bacuth.
GEN|35|9|After Jacob returned from Paddan Aram, God appeared to him again and blessed him.
GEN|35|10|God said to him, "Your name is Jacob, but you will no longer be called Jacob; your name will be Israel. "So he named him Israel.
GEN|35|11|And God said to him, "I am God Almighty; be fruitful and increase in number. A nation and a community of nations will come from you, and kings will come from your body.
GEN|35|12|The land I gave to Abraham and Isaac I also give to you, and I will give this land to your descendants after you."
GEN|35|13|Then God went up from him at the place where he had talked with him.
GEN|35|14|Jacob set up a stone pillar at the place where God had talked with him, and he poured out a drink offering on it; he also poured oil on it.
GEN|35|15|Jacob called the place where God had talked with him Bethel.
GEN|35|16|Then they moved on from Bethel. While they were still some distance from Ephrath, Rachel began to give birth and had great difficulty.
GEN|35|17|And as she was having great difficulty in childbirth, the midwife said to her, "Don't be afraid, for you have another son."
GEN|35|18|As she breathed her last-for she was dying-she named her son Ben-Oni. But his father named him Benjamin.
GEN|35|19|So Rachel died and was buried on the way to Ephrath (that is, Bethlehem).
GEN|35|20|Over her tomb Jacob set up a pillar, and to this day that pillar marks Rachel's tomb.
GEN|35|21|Israel moved on again and pitched his tent beyond Migdal Eder.
GEN|35|22|While Israel was living in that region, Reuben went in and slept with his father's concubine Bilhah, and Israel heard of it. Jacob had twelve sons:
GEN|35|23|The sons of Leah: Reuben the firstborn of Jacob, Simeon, Levi, Judah, Issachar and Zebulun.
GEN|35|24|The sons of Rachel: Joseph and Benjamin.
GEN|35|25|The sons of Rachel's maidservant Bilhah: Dan and Naphtali.
GEN|35|26|The sons of Leah's maidservant Zilpah: Gad and Asher. These were the sons of Jacob, who were born to him in Paddan Aram.
GEN|35|27|Jacob came home to his father Isaac in Mamre, near Kiriath Arba (that is, Hebron), where Abraham and Isaac had stayed.
GEN|35|28|Isaac lived a hundred and eighty years.
GEN|35|29|Then he breathed his last and died and was gathered to his people, old and full of years. And his sons Esau and Jacob buried him.
GEN|36|1|This is the account of Esau (that is, Edom).
GEN|36|2|Esau took his wives from the women of Canaan: Adah daughter of Elon the Hittite, and Oholibamah daughter of Anah and granddaughter of Zibeon the Hivite-
GEN|36|3|also Basemath daughter of Ishmael and sister of Nebaioth.
GEN|36|4|Adah bore Eliphaz to Esau, Basemath bore Reuel,
GEN|36|5|and Oholibamah bore Jeush, Jalam and Korah. These were the sons of Esau, who were born to him in Canaan.
GEN|36|6|Esau took his wives and sons and daughters and all the members of his household, as well as his livestock and all his other animals and all the goods he had acquired in Canaan, and moved to a land some distance from his brother Jacob.
GEN|36|7|Their possessions were too great for them to remain together; the land where they were staying could not support them both because of their livestock.
GEN|36|8|So Esau (that is, Edom) settled in the hill country of Seir.
GEN|36|9|This is the account of Esau the father of the Edomites in the hill country of Seir.
GEN|36|10|These are the names of Esau's sons: Eliphaz, the son of Esau's wife Adah, and Reuel, the son of Esau's wife Basemath.
GEN|36|11|The sons of Eliphaz: Teman, Omar, Zepho, Gatam and Kenaz.
GEN|36|12|Esau's son Eliphaz also had a concubine named Timna, who bore him Amalek. These were grandsons of Esau's wife Adah.
GEN|36|13|The sons of Reuel: Nahath, Zerah, Shammah and Mizzah. These were grandsons of Esau's wife Basemath.
GEN|36|14|The sons of Esau's wife Oholibamah daughter of Anah and granddaughter of Zibeon, whom she bore to Esau: Jeush, Jalam and Korah.
GEN|36|15|These were the chiefs among Esau's descendants: The sons of Eliphaz the firstborn of Esau: Chiefs Teman, Omar, Zepho, Kenaz,
GEN|36|16|Korah, Gatam and Amalek. These were the chiefs descended from Eliphaz in Edom; they were grandsons of Adah.
GEN|36|17|The sons of Esau's son Reuel: Chiefs Nahath, Zerah, Shammah and Mizzah. These were the chiefs descended from Reuel in Edom; they were grandsons of Esau's wife Basemath.
GEN|36|18|The sons of Esau's wife Oholibamah: Chiefs Jeush, Jalam and Korah. These were the chiefs descended from Esau's wife Oholibamah daughter of Anah.
GEN|36|19|These were the sons of Esau (that is, Edom), and these were their chiefs.
GEN|36|20|These were the sons of Seir the Horite, who were living in the region: Lotan, Shobal, Zibeon, Anah,
GEN|36|21|Dishon, Ezer and Dishan. These sons of Seir in Edom were Horite chiefs.
GEN|36|22|The sons of Lotan: Hori and Homam. Timna was Lotan's sister.
GEN|36|23|The sons of Shobal: Alvan, Manahath, Ebal, Shepho and Onam.
GEN|36|24|The sons of Zibeon: Aiah and Anah. This is the Anah who discovered the hot springs in the desert while he was grazing the donkeys of his father Zibeon.
GEN|36|25|The children of Anah: Dishon and Oholibamah daughter of Anah.
GEN|36|26|The sons of Dishon: Hemdan, Eshban, Ithran and Keran.
GEN|36|27|The sons of Ezer: Bilhan, Zaavan and Akan.
GEN|36|28|The sons of Dishan: Uz and Aran.
GEN|36|29|These were the Horite chiefs: Lotan, Shobal, Zibeon, Anah,
GEN|36|30|Dishon, Ezer and Dishan. These were the Horite chiefs, according to their divisions, in the land of Seir.
GEN|36|31|These were the kings who reigned in Edom before any Israelite king reigned:
GEN|36|32|Bela son of Beor became king of Edom. His city was named Dinhabah.
GEN|36|33|When Bela died, Jobab son of Zerah from Bozrah succeeded him as king.
GEN|36|34|When Jobab died, Husham from the land of the Temanites succeeded him as king.
GEN|36|35|When Husham died, Hadad son of Bedad, who defeated Midian in the country of Moab, succeeded him as king. His city was named Avith.
GEN|36|36|When Hadad died, Samlah from Masrekah succeeded him as king.
GEN|36|37|When Samlah died, Shaul from Rehoboth on the river succeeded him as king.
GEN|36|38|When Shaul died, Baal-Hanan son of Acbor succeeded him as king.
GEN|36|39|When Baal-Hanan son of Acbor died, Hadad succeeded him as king. His city was named Pau, and his wife's name was Mehetabel daughter of Matred, the daughter of Me-Zahab.
GEN|36|40|These were the chiefs descended from Esau, by name, according to their clans and regions: Timna, Alvah, Jetheth,
GEN|36|41|Oholibamah, Elah, Pinon,
GEN|36|42|Kenaz, Teman, Mibzar,
GEN|36|43|Magdiel and Iram. These were the chiefs of Edom, according to their settlements in the land they occupied. This was Esau the father of the Edomites.
GEN|37|1|Jacob lived in the land where his father had stayed, the land of Canaan.
GEN|37|2|This is the account of Jacob. Joseph, a young man of seventeen, was tending the flocks with his brothers, the sons of Bilhah and the sons of Zilpah, his father's wives, and he brought their father a bad report about them.
GEN|37|3|Now Israel loved Joseph more than any of his other sons, because he had been born to him in his old age; and he made a richly ornamented robe for him.
GEN|37|4|When his brothers saw that their father loved him more than any of them, they hated him and could not speak a kind word to him.
GEN|37|5|Joseph had a dream, and when he told it to his brothers, they hated him all the more.
GEN|37|6|He said to them, "Listen to this dream I had:
GEN|37|7|We were binding sheaves of grain out in the field when suddenly my sheaf rose and stood upright, while your sheaves gathered around mine and bowed down to it."
GEN|37|8|His brothers said to him, "Do you intend to reign over us? Will you actually rule us?" And they hated him all the more because of his dream and what he had said.
GEN|37|9|Then he had another dream, and he told it to his brothers. "Listen," he said, "I had another dream, and this time the sun and moon and eleven stars were bowing down to me."
GEN|37|10|When he told his father as well as his brothers, his father rebuked him and said, "What is this dream you had? Will your mother and I and your brothers actually come and bow down to the ground before you?"
GEN|37|11|His brothers were jealous of him, but his father kept the matter in mind.
GEN|37|12|Now his brothers had gone to graze their father's flocks near Shechem,
GEN|37|13|and Israel said to Joseph, "As you know, your brothers are grazing the flocks near Shechem. Come, I am going to send you to them.Very well," he replied.
GEN|37|14|So he said to him, "Go and see if all is well with your brothers and with the flocks, and bring word back to me." Then he sent him off from the Valley of Hebron. When Joseph arrived at Shechem,
GEN|37|15|a man found him wandering around in the fields and asked him, "What are you looking for?"
GEN|37|16|He replied, "I'm looking for my brothers. Can you tell me where they are grazing their flocks?"
GEN|37|17|"They have moved on from here," the man answered. "I heard them say, 'Let's go to Dothan.'" So Joseph went after his brothers and found them near Dothan.
GEN|37|18|But they saw him in the distance, and before he reached them, they plotted to kill him.
GEN|37|19|"Here comes that dreamer!" they said to each other.
GEN|37|20|"Come now, let's kill him and throw him into one of these cisterns and say that a ferocious animal devoured him. Then we'll see what comes of his dreams."
GEN|37|21|When Reuben heard this, he tried to rescue him from their hands. "Let's not take his life," he said.
GEN|37|22|"Don't shed any blood. Throw him into this cistern here in the desert, but don't lay a hand on him." Reuben said this to rescue him from them and take him back to his father.
GEN|37|23|So when Joseph came to his brothers, they stripped him of his robe-the richly ornamented robe he was wearing-
GEN|37|24|and they took him and threw him into the cistern. Now the cistern was empty; there was no water in it.
GEN|37|25|As they sat down to eat their meal, they looked up and saw a caravan of Ishmaelites coming from Gilead. Their camels were loaded with spices, balm and myrrh, and they were on their way to take them down to Egypt.
GEN|37|26|Judah said to his brothers, "What will we gain if we kill our brother and cover up his blood?
GEN|37|27|Come, let's sell him to the Ishmaelites and not lay our hands on him; after all, he is our brother, our own flesh and blood." His brothers agreed.
GEN|37|28|So when the Midianite merchants came by, his brothers pulled Joseph up out of the cistern and sold him for twenty shekels of silver to the Ishmaelites, who took him to Egypt.
GEN|37|29|When Reuben returned to the cistern and saw that Joseph was not there, he tore his clothes.
GEN|37|30|He went back to his brothers and said, "The boy isn't there! Where can I turn now?"
GEN|37|31|Then they got Joseph's robe, slaughtered a goat and dipped the robe in the blood.
GEN|37|32|They took the ornamented robe back to their father and said, "We found this. Examine it to see whether it is your son's robe."
GEN|37|33|He recognized it and said, "It is my son's robe! Some ferocious animal has devoured him. Joseph has surely been torn to pieces."
GEN|37|34|Then Jacob tore his clothes, put on sackcloth and mourned for his son many days.
GEN|37|35|All his sons and daughters came to comfort him, but he refused to be comforted. "No," he said, "in mourning will I go down to the grave to my son." So his father wept for him.
GEN|37|36|Meanwhile, the Midianites sold Joseph in Egypt to Potiphar, one of Pharaoh's officials, the captain of the guard.
GEN|38|1|At that time, Judah left his brothers and went down to stay with a man of Adullam named Hirah.
GEN|38|2|There Judah met the daughter of a Canaanite man named Shua. He married her and lay with her;
GEN|38|3|she became pregnant and gave birth to a son, who was named Er.
GEN|38|4|She conceived again and gave birth to a son and named him Onan.
GEN|38|5|She gave birth to still another son and named him Shelah. It was at Kezib that she gave birth to him.
GEN|38|6|Judah got a wife for Er, his firstborn, and her name was Tamar.
GEN|38|7|But Er, Judah's firstborn, was wicked in the LORD's sight; so the LORD put him to death.
GEN|38|8|Then Judah said to Onan, "Lie with your brother's wife and fulfill your duty to her as a brother-in-law to produce offspring for your brother."
GEN|38|9|But Onan knew that the offspring would not be his; so whenever he lay with his brother's wife, he spilled his semen on the ground to keep from producing offspring for his brother.
GEN|38|10|What he did was wicked in the LORD's sight; so he put him to death also.
GEN|38|11|Judah then said to his daughter-in-law Tamar, "Live as a widow in your father's house until my son Shelah grows up." For he thought, "He may die too, just like his brothers." So Tamar went to live in her father's house.
GEN|38|12|After a long time Judah's wife, the daughter of Shua, died. When Judah had recovered from his grief, he went up to Timnah, to the men who were shearing his sheep, and his friend Hirah the Adullamite went with him.
GEN|38|13|When Tamar was told, "Your father-in-law is on his way to Timnah to shear his sheep,"
GEN|38|14|she took off her widow's clothes, covered herself with a veil to disguise herself, and then sat down at the entrance to Enaim, which is on the road to Timnah. For she saw that, though Shelah had now grown up, she had not been given to him as his wife.
GEN|38|15|When Judah saw her, he thought she was a prostitute, for she had covered her face.
GEN|38|16|Not realizing that she was his daughter-in-law, he went over to her by the roadside and said, "Come now, let me sleep with you.And what will you give me to sleep with you?" she asked.
GEN|38|17|"I'll send you a young goat from my flock," he said. "Will you give me something as a pledge until you send it?" she asked.
GEN|38|18|He said, "What pledge should I give you?Your seal and its cord, and the staff in your hand," she answered. So he gave them to her and slept with her, and she became pregnant by him.
GEN|38|19|After she left, she took off her veil and put on her widow's clothes again.
GEN|38|20|Meanwhile Judah sent the young goat by his friend the Adullamite in order to get his pledge back from the woman, but he did not find her.
GEN|38|21|He asked the men who lived there, "Where is the shrine prostitute who was beside the road at Enaim?There hasn't been any shrine prostitute here," they said.
GEN|38|22|So he went back to Judah and said, "I didn't find her. Besides, the men who lived there said, 'There hasn't been any shrine prostitute here.'"
GEN|38|23|Then Judah said, "Let her keep what she has, or we will become a laughingstock. After all, I did send her this young goat, but you didn't find her."
GEN|38|24|About three months later Judah was told, "Your daughter-in-law Tamar is guilty of prostitution, and as a result she is now pregnant." Judah said, "Bring her out and have her burned to death!"
GEN|38|25|As she was being brought out, she sent a message to her father-in-law. "I am pregnant by the man who owns these," she said. And she added, "See if you recognize whose seal and cord and staff these are."
GEN|38|26|Judah recognized them and said, "She is more righteous than I, since I wouldn't give her to my son Shelah." And he did not sleep with her again.
GEN|38|27|When the time came for her to give birth, there were twin boys in her womb.
GEN|38|28|As she was giving birth, one of them put out his hand; so the midwife took a scarlet thread and tied it on his wrist and said, "This one came out first."
GEN|38|29|But when he drew back his hand, his brother came out, and she said, "So this is how you have broken out!" And he was named Perez.
GEN|38|30|Then his brother, who had the scarlet thread on his wrist, came out and he was given the name Zerah.
GEN|39|1|Now Joseph had been taken down to Egypt. Potiphar, an Egyptian who was one of Pharaoh's officials, the captain of the guard, bought him from the Ishmaelites who had taken him there.
GEN|39|2|The LORD was with Joseph and he prospered, and he lived in the house of his Egyptian master.
GEN|39|3|When his master saw that the LORD was with him and that the LORD gave him success in everything he did,
GEN|39|4|Joseph found favor in his eyes and became his attendant. Potiphar put him in charge of his household, and he entrusted to his care everything he owned.
GEN|39|5|From the time he put him in charge of his household and of all that he owned, the LORD blessed the household of the Egyptian because of Joseph. The blessing of the LORD was on everything Potiphar had, both in the house and in the field.
GEN|39|6|So he left in Joseph's care everything he had; with Joseph in charge, he did not concern himself with anything except the food he ate. Now Joseph was well-built and handsome,
GEN|39|7|and after a while his master's wife took notice of Joseph and said, "Come to bed with me!"
GEN|39|8|But he refused. "With me in charge," he told her, "my master does not concern himself with anything in the house; everything he owns he has entrusted to my care.
GEN|39|9|No one is greater in this house than I am. My master has withheld nothing from me except you, because you are his wife. How then could I do such a wicked thing and sin against God?"
GEN|39|10|And though she spoke to Joseph day after day, he refused to go to bed with her or even be with her.
GEN|39|11|One day he went into the house to attend to his duties, and none of the household servants was inside.
GEN|39|12|She caught him by his cloak and said, "Come to bed with me!" But he left his cloak in her hand and ran out of the house.
GEN|39|13|When she saw that he had left his cloak in her hand and had run out of the house,
GEN|39|14|she called her household servants. "Look," she said to them, "this Hebrew has been brought to us to make sport of us! He came in here to sleep with me, but I screamed.
GEN|39|15|When he heard me scream for help, he left his cloak beside me and ran out of the house."
GEN|39|16|She kept his cloak beside her until his master came home.
GEN|39|17|Then she told him this story: "That Hebrew slave you brought us came to me to make sport of me.
GEN|39|18|But as soon as I screamed for help, he left his cloak beside me and ran out of the house."
GEN|39|19|When his master heard the story his wife told him, saying, "This is how your slave treated me," he burned with anger.
GEN|39|20|Joseph's master took him and put him in prison, the place where the king's prisoners were confined. But while Joseph was there in the prison,
GEN|39|21|the LORD was with him; he showed him kindness and granted him favor in the eyes of the prison warden.
GEN|39|22|So the warden put Joseph in charge of all those held in the prison, and he was made responsible for all that was done there.
GEN|39|23|The warden paid no attention to anything under Joseph's care, because the LORD was with Joseph and gave him success in whatever he did.
GEN|40|1|Some time later, the cupbearer and the baker of the king of Egypt offended their master, the king of Egypt.
GEN|40|2|Pharaoh was angry with his two officials, the chief cupbearer and the chief baker,
GEN|40|3|and put them in custody in the house of the captain of the guard, in the same prison where Joseph was confined.
GEN|40|4|The captain of the guard assigned them to Joseph, and he attended them. After they had been in custody for some time,
GEN|40|5|each of the two men-the cupbearer and the baker of the king of Egypt, who were being held in prison-had a dream the same night, and each dream had a meaning of its own.
GEN|40|6|When Joseph came to them the next morning, he saw that they were dejected.
GEN|40|7|So he asked Pharaoh's officials who were in custody with him in his master's house, "Why are your faces so sad today?"
GEN|40|8|"We both had dreams," they answered, "but there is no one to interpret them." Then Joseph said to them, "Do not interpretations belong to God? Tell me your dreams."
GEN|40|9|So the chief cupbearer told Joseph his dream. He said to him, "In my dream I saw a vine in front of me,
GEN|40|10|and on the vine were three branches. As soon as it budded, it blossomed, and its clusters ripened into grapes.
GEN|40|11|Pharaoh's cup was in my hand, and I took the grapes, squeezed them into Pharaoh's cup and put the cup in his hand."
GEN|40|12|"This is what it means," Joseph said to him. "The three branches are three days.
GEN|40|13|Within three days Pharaoh will lift up your head and restore you to your position, and you will put Pharaoh's cup in his hand, just as you used to do when you were his cupbearer.
GEN|40|14|But when all goes well with you, remember me and show me kindness; mention me to Pharaoh and get me out of this prison.
GEN|40|15|For I was forcibly carried off from the land of the Hebrews, and even here I have done nothing to deserve being put in a dungeon."
GEN|40|16|When the chief baker saw that Joseph had given a favorable interpretation, he said to Joseph, "I too had a dream: On my head were three baskets of bread.
GEN|40|17|In the top basket were all kinds of baked goods for Pharaoh, but the birds were eating them out of the basket on my head."
GEN|40|18|"This is what it means," Joseph said. "The three baskets are three days.
GEN|40|19|Within three days Pharaoh will lift off your head and hang you on a tree. And the birds will eat away your flesh."
GEN|40|20|Now the third day was Pharaoh's birthday, and he gave a feast for all his officials. He lifted up the heads of the chief cupbearer and the chief baker in the presence of his officials:
GEN|40|21|He restored the chief cupbearer to his position, so that he once again put the cup into Pharaoh's hand,
GEN|40|22|but he hanged the chief baker, just as Joseph had said to them in his interpretation.
GEN|40|23|The chief cupbearer, however, did not remember Joseph; he forgot him.
GEN|41|1|When two full years had passed, Pharaoh had a dream: He was standing by the Nile,
GEN|41|2|when out of the river there came up seven cows, sleek and fat, and they grazed among the reeds.
GEN|41|3|After them, seven other cows, ugly and gaunt, came up out of the Nile and stood beside those on the riverbank.
GEN|41|4|And the cows that were ugly and gaunt ate up the seven sleek, fat cows. Then Pharaoh woke up.
GEN|41|5|He fell asleep again and had a second dream: Seven heads of grain, healthy and good, were growing on a single stalk.
GEN|41|6|After them, seven other heads of grain sprouted-thin and scorched by the east wind.
GEN|41|7|The thin heads of grain swallowed up the seven healthy, full heads. Then Pharaoh woke up; it had been a dream.
GEN|41|8|In the morning his mind was troubled, so he sent for all the magicians and wise men of Egypt. Pharaoh told them his dreams, but no one could interpret them for him.
GEN|41|9|Then the chief cupbearer said to Pharaoh, "Today I am reminded of my shortcomings.
GEN|41|10|Pharaoh was once angry with his servants, and he imprisoned me and the chief baker in the house of the captain of the guard.
GEN|41|11|Each of us had a dream the same night, and each dream had a meaning of its own.
GEN|41|12|Now a young Hebrew was there with us, a servant of the captain of the guard. We told him our dreams, and he interpreted them for us, giving each man the interpretation of his dream.
GEN|41|13|And things turned out exactly as he interpreted them to us: I was restored to my position, and the other man was hanged. "
GEN|41|14|So Pharaoh sent for Joseph, and he was quickly brought from the dungeon. When he had shaved and changed his clothes, he came before Pharaoh.
GEN|41|15|Pharaoh said to Joseph, "I had a dream, and no one can interpret it. But I have heard it said of you that when you hear a dream you can interpret it."
GEN|41|16|"I cannot do it," Joseph replied to Pharaoh, "but God will give Pharaoh the answer he desires."
GEN|41|17|Then Pharaoh said to Joseph, "In my dream I was standing on the bank of the Nile,
GEN|41|18|when out of the river there came up seven cows, fat and sleek, and they grazed among the reeds.
GEN|41|19|After them, seven other cows came up-scrawny and very ugly and lean. I had never seen such ugly cows in all the land of Egypt.
GEN|41|20|The lean, ugly cows ate up the seven fat cows that came up first.
GEN|41|21|But even after they ate them, no one could tell that they had done so; they looked just as ugly as before. Then I woke up.
GEN|41|22|"In my dreams I also saw seven heads of grain, full and good, growing on a single stalk.
GEN|41|23|After them, seven other heads sprouted-withered and thin and scorched by the east wind.
GEN|41|24|The thin heads of grain swallowed up the seven good heads. I told this to the magicians, but none could explain it to me."
GEN|41|25|Then Joseph said to Pharaoh, "The dreams of Pharaoh are one and the same. God has revealed to Pharaoh what he is about to do.
GEN|41|26|The seven good cows are seven years, and the seven good heads of grain are seven years; it is one and the same dream.
GEN|41|27|The seven lean, ugly cows that came up afterward are seven years, and so are the seven worthless heads of grain scorched by the east wind: They are seven years of famine.
GEN|41|28|"It is just as I said to Pharaoh: God has shown Pharaoh what he is about to do.
GEN|41|29|Seven years of great abundance are coming throughout the land of Egypt,
GEN|41|30|but seven years of famine will follow them. Then all the abundance in Egypt will be forgotten, and the famine will ravage the land.
GEN|41|31|The abundance in the land will not be remembered, because the famine that follows it will be so severe.
GEN|41|32|The reason the dream was given to Pharaoh in two forms is that the matter has been firmly decided by God, and God will do it soon.
GEN|41|33|"And now let Pharaoh look for a discerning and wise man and put him in charge of the land of Egypt.
GEN|41|34|Let Pharaoh appoint commissioners over the land to take a fifth of the harvest of Egypt during the seven years of abundance.
GEN|41|35|They should collect all the food of these good years that are coming and store up the grain under the authority of Pharaoh, to be kept in the cities for food.
GEN|41|36|This food should be held in reserve for the country, to be used during the seven years of famine that will come upon Egypt, so that the country may not be ruined by the famine."
GEN|41|37|The plan seemed good to Pharaoh and to all his officials.
GEN|41|38|So Pharaoh asked them, "Can we find anyone like this man, one in whom is the spirit of God?"
GEN|41|39|Then Pharaoh said to Joseph, "Since God has made all this known to you, there is no one so discerning and wise as you.
GEN|41|40|You shall be in charge of my palace, and all my people are to submit to your orders. Only with respect to the throne will I be greater than you."
GEN|41|41|So Pharaoh said to Joseph, "I hereby put you in charge of the whole land of Egypt."
GEN|41|42|Then Pharaoh took his signet ring from his finger and put it on Joseph's finger. He dressed him in robes of fine linen and put a gold chain around his neck.
GEN|41|43|He had him ride in a chariot as his second-in-command, and men shouted before him, "Make way!" Thus he put him in charge of the whole land of Egypt.
GEN|41|44|Then Pharaoh said to Joseph, "I am Pharaoh, but without your word no one will lift hand or foot in all Egypt."
GEN|41|45|Pharaoh gave Joseph the name Zaphenath-Paneah and gave him Asenath daughter of Potiphera, priest of On, to be his wife. And Joseph went throughout the land of Egypt.
GEN|41|46|Joseph was thirty years old when he entered the service of Pharaoh king of Egypt. And Joseph went out from Pharaoh's presence and traveled throughout Egypt.
GEN|41|47|During the seven years of abundance the land produced plentifully.
GEN|41|48|Joseph collected all the food produced in those seven years of abundance in Egypt and stored it in the cities. In each city he put the food grown in the fields surrounding it.
GEN|41|49|Joseph stored up huge quantities of grain, like the sand of the sea; it was so much that he stopped keeping records because it was beyond measure.
GEN|41|50|Before the years of famine came, two sons were born to Joseph by Asenath daughter of Potiphera, priest of On.
GEN|41|51|Joseph named his firstborn Manasseh and said, "It is because God has made me forget all my trouble and all my father's household."
GEN|41|52|The second son he named Ephraim and said, "It is because God has made me fruitful in the land of my suffering."
GEN|41|53|The seven years of abundance in Egypt came to an end,
GEN|41|54|and the seven years of famine began, just as Joseph had said. There was famine in all the other lands, but in the whole land of Egypt there was food.
GEN|41|55|When all Egypt began to feel the famine, the people cried to Pharaoh for food. Then Pharaoh told all the Egyptians, "Go to Joseph and do what he tells you."
GEN|41|56|When the famine had spread over the whole country, Joseph opened the storehouses and sold grain to the Egyptians, for the famine was severe throughout Egypt.
GEN|41|57|And all the countries came to Egypt to buy grain from Joseph, because the famine was severe in all the world.
GEN|42|1|When Jacob learned that there was grain in Egypt, he said to his sons, "Why do you just keep looking at each other?"
GEN|42|2|He continued, "I have heard that there is grain in Egypt. Go down there and buy some for us, so that we may live and not die."
GEN|42|3|Then ten of Joseph's brothers went down to buy grain from Egypt.
GEN|42|4|But Jacob did not send Benjamin, Joseph's brother, with the others, because he was afraid that harm might come to him.
GEN|42|5|So Israel's sons were among those who went to buy grain, for the famine was in the land of Canaan also.
GEN|42|6|Now Joseph was the governor of the land, the one who sold grain to all its people. So when Joseph's brothers arrived, they bowed down to him with their faces to the ground.
GEN|42|7|As soon as Joseph saw his brothers, he recognized them, but he pretended to be a stranger and spoke harshly to them. "Where do you come from?" he asked. "From the land of Canaan," they replied, "to buy food."
GEN|42|8|Although Joseph recognized his brothers, they did not recognize him.
GEN|42|9|Then he remembered his dreams about them and said to them, "You are spies! You have come to see where our land is unprotected."
GEN|42|10|"No, my lord," they answered. "Your servants have come to buy food.
GEN|42|11|We are all the sons of one man. Your servants are honest men, not spies."
GEN|42|12|"No!" he said to them. "You have come to see where our land is unprotected."
GEN|42|13|But they replied, "Your servants were twelve brothers, the sons of one man, who lives in the land of Canaan. The youngest is now with our father, and one is no more."
GEN|42|14|Joseph said to them, "It is just as I told you: You are spies!
GEN|42|15|And this is how you will be tested: As surely as Pharaoh lives, you will not leave this place unless your youngest brother comes here.
GEN|42|16|Send one of your number to get your brother; the rest of you will be kept in prison, so that your words may be tested to see if you are telling the truth. If you are not, then as surely as Pharaoh lives, you are spies!"
GEN|42|17|And he put them all in custody for three days.
GEN|42|18|On the third day, Joseph said to them, "Do this and you will live, for I fear God:
GEN|42|19|If you are honest men, let one of your brothers stay here in prison, while the rest of you go and take grain back for your starving households.
GEN|42|20|But you must bring your youngest brother to me, so that your words may be verified and that you may not die." This they proceeded to do.
GEN|42|21|They said to one another, "Surely we are being punished because of our brother. We saw how distressed he was when he pleaded with us for his life, but we would not listen; that's why this distress has come upon us."
GEN|42|22|Reuben replied, "Didn't I tell you not to sin against the boy? But you wouldn't listen! Now we must give an accounting for his blood."
GEN|42|23|They did not realize that Joseph could understand them, since he was using an interpreter.
GEN|42|24|He turned away from them and began to weep, but then turned back and spoke to them again. He had Simeon taken from them and bound before their eyes.
GEN|42|25|Joseph gave orders to fill their bags with grain, to put each man's silver back in his sack, and to give them provisions for their journey. After this was done for them,
GEN|42|26|they loaded their grain on their donkeys and left.
GEN|42|27|At the place where they stopped for the night one of them opened his sack to get feed for his donkey, and he saw his silver in the mouth of his sack.
GEN|42|28|"My silver has been returned," he said to his brothers. "Here it is in my sack." Their hearts sank and they turned to each other trembling and said, "What is this that God has done to us?"
GEN|42|29|When they came to their father Jacob in the land of Canaan, they told him all that had happened to them. They said,
GEN|42|30|"The man who is lord over the land spoke harshly to us and treated us as though we were spying on the land.
GEN|42|31|But we said to him, 'We are honest men; we are not spies.
GEN|42|32|We were twelve brothers, sons of one father. One is no more, and the youngest is now with our father in Canaan.'
GEN|42|33|"Then the man who is lord over the land said to us, 'This is how I will know whether you are honest men: Leave one of your brothers here with me, and take food for your starving households and go.
GEN|42|34|But bring your youngest brother to me so I will know that you are not spies but honest men. Then I will give your brother back to you, and you can trade in the land.'"
GEN|42|35|As they were emptying their sacks, there in each man's sack was his pouch of silver! When they and their father saw the money pouches, they were frightened.
GEN|42|36|Their father Jacob said to them, "You have deprived me of my children. Joseph is no more and Simeon is no more, and now you want to take Benjamin. Everything is against me!"
GEN|42|37|Then Reuben said to his father, "You may put both of my sons to death if I do not bring him back to you. Entrust him to my care, and I will bring him back."
GEN|42|38|But Jacob said, "My son will not go down there with you; his brother is dead and he is the only one left. If harm comes to him on the journey you are taking, you will bring my gray head down to the grave in sorrow."
GEN|43|1|Now the famine was still severe in the land.
GEN|43|2|So when they had eaten all the grain they had brought from Egypt, their father said to them, "Go back and buy us a little more food."
GEN|43|3|But Judah said to him, "The man warned us solemnly, 'You will not see my face again unless your brother is with you.'
GEN|43|4|If you will send our brother along with us, we will go down and buy food for you.
GEN|43|5|But if you will not send him, we will not go down, because the man said to us, 'You will not see my face again unless your brother is with you.'"
GEN|43|6|Israel asked, "Why did you bring this trouble on me by telling the man you had another brother?"
GEN|43|7|They replied, "The man questioned us closely about ourselves and our family. 'Is your father still living?' he asked us. 'Do you have another brother?' We simply answered his questions. How were we to know he would say, 'Bring your brother down here'?"
GEN|43|8|Then Judah said to Israel his father, "Send the boy along with me and we will go at once, so that we and you and our children may live and not die.
GEN|43|9|I myself will guarantee his safety; you can hold me personally responsible for him. If I do not bring him back to you and set him here before you, I will bear the blame before you all my life.
GEN|43|10|As it is, if we had not delayed, we could have gone and returned twice."
GEN|43|11|Then their father Israel said to them, "If it must be, then do this: Put some of the best products of the land in your bags and take them down to the man as a gift-a little balm and a little honey, some spices and myrrh, some pistachio nuts and almonds.
GEN|43|12|Take double the amount of silver with you, for you must return the silver that was put back into the mouths of your sacks. Perhaps it was a mistake.
GEN|43|13|Take your brother also and go back to the man at once.
GEN|43|14|And may God Almighty grant you mercy before the man so that he will let your other brother and Benjamin come back with you. As for me, if I am bereaved, I am bereaved."
GEN|43|15|So the men took the gifts and double the amount of silver, and Benjamin also. They hurried down to Egypt and presented themselves to Joseph.
GEN|43|16|When Joseph saw Benjamin with them, he said to the steward of his house, "Take these men to my house, slaughter an animal and prepare dinner; they are to eat with me at noon."
GEN|43|17|The man did as Joseph told him and took the men to Joseph's house.
GEN|43|18|Now the men were frightened when they were taken to his house. They thought, "We were brought here because of the silver that was put back into our sacks the first time. He wants to attack us and overpower us and seize us as slaves and take our donkeys."
GEN|43|19|So they went up to Joseph's steward and spoke to him at the entrance to the house.
GEN|43|20|"Please, sir," they said, "we came down here the first time to buy food.
GEN|43|21|But at the place where we stopped for the night we opened our sacks and each of us found his silver-the exact weight-in the mouth of his sack. So we have brought it back with us.
GEN|43|22|We have also brought additional silver with us to buy food. We don't know who put our silver in our sacks."
GEN|43|23|"It's all right," he said. "Don't be afraid. Your God, the God of your father, has given you treasure in your sacks; I received your silver." Then he brought Simeon out to them.
GEN|43|24|The steward took the men into Joseph's house, gave them water to wash their feet and provided fodder for their donkeys.
GEN|43|25|They prepared their gifts for Joseph's arrival at noon, because they had heard that they were to eat there.
GEN|43|26|When Joseph came home, they presented to him the gifts they had brought into the house, and they bowed down before him to the ground.
GEN|43|27|He asked them how they were, and then he said, "How is your aged father you told me about? Is he still living?"
GEN|43|28|They replied, "Your servant our father is still alive and well." And they bowed low to pay him honor.
GEN|43|29|As he looked about and saw his brother Benjamin, his own mother's son, he asked, "Is this your youngest brother, the one you told me about?" And he said, "God be gracious to you, my son."
GEN|43|30|Deeply moved at the sight of his brother, Joseph hurried out and looked for a place to weep. He went into his private room and wept there.
GEN|43|31|After he had washed his face, he came out and, controlling himself, said, "Serve the food."
GEN|43|32|They served him by himself, the brothers by themselves, and the Egyptians who ate with him by themselves, because Egyptians could not eat with Hebrews, for that is detestable to Egyptians.
GEN|43|33|The men had been seated before him in the order of their ages, from the firstborn to the youngest; and they looked at each other in astonishment.
GEN|43|34|When portions were served to them from Joseph's table, Benjamin's portion was five times as much as anyone else's. So they feasted and drank freely with him.
GEN|44|1|Now Joseph gave these instructions to the steward of his house: "Fill the men's sacks with as much food as they can carry, and put each man's silver in the mouth of his sack.
GEN|44|2|Then put my cup, the silver one, in the mouth of the youngest one's sack, along with the silver for his grain." And he did as Joseph said.
GEN|44|3|As morning dawned, the men were sent on their way with their donkeys.
GEN|44|4|They had not gone far from the city when Joseph said to his steward, "Go after those men at once, and when you catch up with them, say to them, 'Why have you repaid good with evil?
GEN|44|5|Isn't this the cup my master drinks from and also uses for divination? This is a wicked thing you have done.'"
GEN|44|6|When he caught up with them, he repeated these words to them.
GEN|44|7|But they said to him, "Why does my lord say such things? Far be it from your servants to do anything like that!
GEN|44|8|We even brought back to you from the land of Canaan the silver we found inside the mouths of our sacks. So why would we steal silver or gold from your master's house?
GEN|44|9|If any of your servants is found to have it, he will die; and the rest of us will become my lord's slaves."
GEN|44|10|"Very well, then," he said, "let it be as you say. Whoever is found to have it will become my slave; the rest of you will be free from blame."
GEN|44|11|Each of them quickly lowered his sack to the ground and opened it.
GEN|44|12|Then the steward proceeded to search, beginning with the oldest and ending with the youngest. And the cup was found in Benjamin's sack.
GEN|44|13|At this, they tore their clothes. Then they all loaded their donkeys and returned to the city.
GEN|44|14|Joseph was still in the house when Judah and his brothers came in, and they threw themselves to the ground before him.
GEN|44|15|Joseph said to them, "What is this you have done? Don't you know that a man like me can find things out by divination?"
GEN|44|16|"What can we say to my lord?" Judah replied. "What can we say? How can we prove our innocence? God has uncovered your servants' guilt. We are now my lord's slaves-we ourselves and the one who was found to have the cup."
GEN|44|17|But Joseph said, "Far be it from me to do such a thing! Only the man who was found to have the cup will become my slave. The rest of you, go back to your father in peace."
GEN|44|18|Then Judah went up to him and said: "Please, my lord, let your servant speak a word to my lord. Do not be angry with your servant, though you are equal to Pharaoh himself.
GEN|44|19|My lord asked his servants, 'Do you have a father or a brother?'
GEN|44|20|And we answered, 'We have an aged father, and there is a young son born to him in his old age. His brother is dead, and he is the only one of his mother's sons left, and his father loves him.'
GEN|44|21|"Then you said to your servants, 'Bring him down to me so I can see him for myself.'
GEN|44|22|And we said to my lord, 'The boy cannot leave his father; if he leaves him, his father will die.'
GEN|44|23|But you told your servants, 'Unless your youngest brother comes down with you, you will not see my face again.'
GEN|44|24|When we went back to your servant my father, we told him what my lord had said.
GEN|44|25|"Then our father said, 'Go back and buy a little more food.'
GEN|44|26|But we said, 'We cannot go down. Only if our youngest brother is with us will we go. We cannot see the man's face unless our youngest brother is with us.'
GEN|44|27|"Your servant my father said to us, 'You know that my wife bore me two sons.
GEN|44|28|One of them went away from me, and I said, "He has surely been torn to pieces." And I have not seen him since.
GEN|44|29|If you take this one from me too and harm comes to him, you will bring my gray head down to the grave in misery.'
GEN|44|30|"So now, if the boy is not with us when I go back to your servant my father and if my father, whose life is closely bound up with the boy's life,
GEN|44|31|sees that the boy isn't there, he will die. Your servants will bring the gray head of our father down to the grave in sorrow.
GEN|44|32|Your servant guaranteed the boy's safety to my father. I said, 'If I do not bring him back to you, I will bear the blame before you, my father, all my life!'
GEN|44|33|"Now then, please let your servant remain here as my lord's slave in place of the boy, and let the boy return with his brothers.
GEN|44|34|How can I go back to my father if the boy is not with me? No! Do not let me see the misery that would come upon my father."
GEN|45|1|Then Joseph could no longer control himself before all his attendants, and he cried out, "Have everyone leave my presence!" So there was no one with Joseph when he made himself known to his brothers.
GEN|45|2|And he wept so loudly that the Egyptians heard him, and Pharaoh's household heard about it.
GEN|45|3|Joseph said to his brothers, "I am Joseph! Is my father still living?" But his brothers were not able to answer him, because they were terrified at his presence.
GEN|45|4|Then Joseph said to his brothers, "Come close to me." When they had done so, he said, "I am your brother Joseph, the one you sold into Egypt!
GEN|45|5|And now, do not be distressed and do not be angry with yourselves for selling me here, because it was to save lives that God sent me ahead of you.
GEN|45|6|For two years now there has been famine in the land, and for the next five years there will not be plowing and reaping.
GEN|45|7|But God sent me ahead of you to preserve for you a remnant on earth and to save your lives by a great deliverance.
GEN|45|8|"So then, it was not you who sent me here, but God. He made me father to Pharaoh, lord of his entire household and ruler of all Egypt.
GEN|45|9|Now hurry back to my father and say to him, 'This is what your son Joseph says: God has made me lord of all Egypt. Come down to me; don't delay.
GEN|45|10|You shall live in the region of Goshen and be near me-you, your children and grandchildren, your flocks and herds, and all you have.
GEN|45|11|I will provide for you there, because five years of famine are still to come. Otherwise you and your household and all who belong to you will become destitute.'
GEN|45|12|"You can see for yourselves, and so can my brother Benjamin, that it is really I who am speaking to you.
GEN|45|13|Tell my father about all the honor accorded me in Egypt and about everything you have seen. And bring my father down here quickly."
GEN|45|14|Then he threw his arms around his brother Benjamin and wept, and Benjamin embraced him, weeping.
GEN|45|15|And he kissed all his brothers and wept over them. Afterward his brothers talked with him.
GEN|45|16|When the news reached Pharaoh's palace that Joseph's brothers had come, Pharaoh and all his officials were pleased.
GEN|45|17|Pharaoh said to Joseph, "Tell your brothers, 'Do this: Load your animals and return to the land of Canaan,
GEN|45|18|and bring your father and your families back to me. I will give you the best of the land of Egypt and you can enjoy the fat of the land.'
GEN|45|19|"You are also directed to tell them, 'Do this: Take some carts from Egypt for your children and your wives, and get your father and come.
GEN|45|20|Never mind about your belongings, because the best of all Egypt will be yours.'"
GEN|45|21|So the sons of Israel did this. Joseph gave them carts, as Pharaoh had commanded, and he also gave them provisions for their journey.
GEN|45|22|To each of them he gave new clothing, but to Benjamin he gave three hundred shekels of silver and five sets of clothes.
GEN|45|23|And this is what he sent to his father: ten donkeys loaded with the best things of Egypt, and ten female donkeys loaded with grain and bread and other provisions for his journey.
GEN|45|24|Then he sent his brothers away, and as they were leaving he said to them, "Don't quarrel on the way!"
GEN|45|25|So they went up out of Egypt and came to their father Jacob in the land of Canaan.
GEN|45|26|They told him, "Joseph is still alive! In fact, he is ruler of all Egypt." Jacob was stunned; he did not believe them.
GEN|45|27|But when they told him everything Joseph had said to them, and when he saw the carts Joseph had sent to carry him back, the spirit of their father Jacob revived.
GEN|45|28|And Israel said, "I'm convinced! My son Joseph is still alive. I will go and see him before I die."
GEN|46|1|So Israel set out with all that was his, and when he reached Beersheba, he offered sacrifices to the God of his father Isaac.
GEN|46|2|And God spoke to Israel in a vision at night and said, "Jacob! Jacob!Here I am," he replied.
GEN|46|3|"I am God, the God of your father," he said. "Do not be afraid to go down to Egypt, for I will make you into a great nation there.
GEN|46|4|I will go down to Egypt with you, and I will surely bring you back again. And Joseph's own hand will close your eyes."
GEN|46|5|Then Jacob left Beersheba, and Israel's sons took their father Jacob and their children and their wives in the carts that Pharaoh had sent to transport him.
GEN|46|6|They also took with them their livestock and the possessions they had acquired in Canaan, and Jacob and all his offspring went to Egypt.
GEN|46|7|He took with him to Egypt his sons and grandsons and his daughters and granddaughters-all his offspring.
GEN|46|8|These are the names of the sons of Israel (Jacob and his descendants) who went to Egypt: Reuben the firstborn of Jacob.
GEN|46|9|The sons of Reuben: Hanoch, Pallu, Hezron and Carmi.
GEN|46|10|The sons of Simeon: Jemuel, Jamin, Ohad, Jakin, Zohar and Shaul the son of a Canaanite woman.
GEN|46|11|The sons of Levi: Gershon, Kohath and Merari.
GEN|46|12|The sons of Judah: Er, Onan, Shelah, Perez and Zerah (but Er and Onan had died in the land of Canaan). The sons of Perez: Hezron and Hamul.
GEN|46|13|The sons of Issachar: Tola, Puah, Jashub and Shimron.
GEN|46|14|The sons of Zebulun: Sered, Elon and Jahleel.
GEN|46|15|These were the sons Leah bore to Jacob in Paddan Aram, besides his daughter Dinah. These sons and daughters of his were thirty-three in all.
GEN|46|16|The sons of Gad: Zephon, Haggi, Shuni, Ezbon, Eri, Arodi and Areli.
GEN|46|17|The sons of Asher: Imnah, Ishvah, Ishvi and Beriah. Their sister was Serah. The sons of Beriah: Heber and Malkiel.
GEN|46|18|These were the children born to Jacob by Zilpah, whom Laban had given to his daughter Leah-sixteen in all.
GEN|46|19|The sons of Jacob's wife Rachel: Joseph and Benjamin.
GEN|46|20|In Egypt, Manasseh and Ephraim were born to Joseph by Asenath daughter of Potiphera, priest of On.
GEN|46|21|The sons of Benjamin: Bela, Beker, Ashbel, Gera, Naaman, Ehi, Rosh, Muppim, Huppim and Ard.
GEN|46|22|These were the sons of Rachel who were born to Jacob-fourteen in all.
GEN|46|23|The son of Dan: Hushim.
GEN|46|24|The sons of Naphtali: Jahziel, Guni, Jezer and Shillem.
GEN|46|25|These were the sons born to Jacob by Bilhah, whom Laban had given to his daughter Rachel-seven in all.
GEN|46|26|All those who went to Egypt with Jacob-those who were his direct descendants, not counting his sons' wives-numbered sixty-six persons.
GEN|46|27|With the two sons who had been born to Joseph in Egypt, the members of Jacob's family, which went to Egypt, were seventy in all.
GEN|46|28|Now Jacob sent Judah ahead of him to Joseph to get directions to Goshen. When they arrived in the region of Goshen,
GEN|46|29|Joseph had his chariot made ready and went to Goshen to meet his father Israel. As soon as Joseph appeared before him, he threw his arms around his father and wept for a long time.
GEN|46|30|Israel said to Joseph, "Now I am ready to die, since I have seen for myself that you are still alive."
GEN|46|31|Then Joseph said to his brothers and to his father's household, "I will go up and speak to Pharaoh and will say to him, 'My brothers and my father's household, who were living in the land of Canaan, have come to me.
GEN|46|32|The men are shepherds; they tend livestock, and they have brought along their flocks and herds and everything they own.'
GEN|46|33|When Pharaoh calls you in and asks, 'What is your occupation?'
GEN|46|34|you should answer, 'Your servants have tended livestock from our boyhood on, just as our fathers did.' Then you will be allowed to settle in the region of Goshen, for all shepherds are detestable to the Egyptians."
GEN|47|1|Joseph went and told Pharaoh, "My father and brothers, with their flocks and herds and everything they own, have come from the land of Canaan and are now in Goshen."
GEN|47|2|He chose five of his brothers and presented them before Pharaoh.
GEN|47|3|Pharaoh asked the brothers, "What is your occupation?Your servants are shepherds," they replied to Pharaoh, "just as our fathers were."
GEN|47|4|They also said to him, "We have come to live here awhile, because the famine is severe in Canaan and your servants' flocks have no pasture. So now, please let your servants settle in Goshen."
GEN|47|5|Pharaoh said to Joseph, "Your father and your brothers have come to you,
GEN|47|6|and the land of Egypt is before you; settle your father and your brothers in the best part of the land. Let them live in Goshen. And if you know of any among them with special ability, put them in charge of my own livestock."
GEN|47|7|Then Joseph brought his father Jacob in and presented him before Pharaoh. After Jacob blessed Pharaoh,
GEN|47|8|Pharaoh asked him, "How old are you?"
GEN|47|9|And Jacob said to Pharaoh, "The years of my pilgrimage are a hundred and thirty. My years have been few and difficult, and they do not equal the years of the pilgrimage of my fathers."
GEN|47|10|Then Jacob blessed Pharaoh and went out from his presence.
GEN|47|11|So Joseph settled his father and his brothers in Egypt and gave them property in the best part of the land, the district of Rameses, as Pharaoh directed.
GEN|47|12|Joseph also provided his father and his brothers and all his father's household with food, according to the number of their children.
GEN|47|13|There was no food, however, in the whole region because the famine was severe; both Egypt and Canaan wasted away because of the famine.
GEN|47|14|Joseph collected all the money that was to be found in Egypt and Canaan in payment for the grain they were buying, and he brought it to Pharaoh's palace.
GEN|47|15|When the money of the people of Egypt and Canaan was gone, all Egypt came to Joseph and said, "Give us food. Why should we die before your eyes? Our money is used up."
GEN|47|16|"Then bring your livestock," said Joseph. "I will sell you food in exchange for your livestock, since your money is gone."
GEN|47|17|So they brought their livestock to Joseph, and he gave them food in exchange for their horses, their sheep and goats, their cattle and donkeys. And he brought them through that year with food in exchange for all their livestock.
GEN|47|18|When that year was over, they came to him the following year and said, "We cannot hide from our lord the fact that since our money is gone and our livestock belongs to you, there is nothing left for our lord except our bodies and our land.
GEN|47|19|Why should we perish before your eyes-we and our land as well? Buy us and our land in exchange for food, and we with our land will be in bondage to Pharaoh. Give us seed so that we may live and not die, and that the land may not become desolate."
GEN|47|20|So Joseph bought all the land in Egypt for Pharaoh. The Egyptians, one and all, sold their fields, because the famine was too severe for them. The land became Pharaoh's,
GEN|47|21|and Joseph reduced the people to servitude, from one end of Egypt to the other.
GEN|47|22|However, he did not buy the land of the priests, because they received a regular allotment from Pharaoh and had food enough from the allotment Pharaoh gave them. That is why they did not sell their land.
GEN|47|23|Joseph said to the people, "Now that I have bought you and your land today for Pharaoh, here is seed for you so you can plant the ground.
GEN|47|24|But when the crop comes in, give a fifth of it to Pharaoh. The other four-fifths you may keep as seed for the fields and as food for yourselves and your households and your children."
GEN|47|25|"You have saved our lives," they said. "May we find favor in the eyes of our lord; we will be in bondage to Pharaoh."
GEN|47|26|So Joseph established it as a law concerning land in Egypt-still in force today-that a fifth of the produce belongs to Pharaoh. It was only the land of the priests that did not become Pharaoh's.
GEN|47|27|Now the Israelites settled in Egypt in the region of Goshen. They acquired property there and were fruitful and increased greatly in number.
GEN|47|28|Jacob lived in Egypt seventeen years, and the years of his life were a hundred and forty-seven.
GEN|47|29|When the time drew near for Israel to die, he called for his son Joseph and said to him, "If I have found favor in your eyes, put your hand under my thigh and promise that you will show me kindness and faithfulness. Do not bury me in Egypt,
GEN|47|30|but when I rest with my fathers, carry me out of Egypt and bury me where they are buried.I will do as you say," he said.
GEN|47|31|"Swear to me," he said. Then Joseph swore to him, and Israel worshiped as he leaned on the top of his staff.
GEN|48|1|Some time later Joseph was told, "Your father is ill." So he took his two sons Manasseh and Ephraim along with him.
GEN|48|2|When Jacob was told, "Your son Joseph has come to you," Israel rallied his strength and sat up on the bed.
GEN|48|3|Jacob said to Joseph, "God Almighty appeared to me at Luz in the land of Canaan, and there he blessed me
GEN|48|4|and said to me, 'I am going to make you fruitful and will increase your numbers. I will make you a community of peoples, and I will give this land as an everlasting possession to your descendants after you.'
GEN|48|5|"Now then, your two sons born to you in Egypt before I came to you here will be reckoned as mine; Ephraim and Manasseh will be mine, just as Reuben and Simeon are mine.
GEN|48|6|Any children born to you after them will be yours; in the territory they inherit they will be reckoned under the names of their brothers.
GEN|48|7|As I was returning from Paddan, to my sorrow Rachel died in the land of Canaan while we were still on the way, a little distance from Ephrath. So I buried her there beside the road to Ephrath" (that is, Bethlehem).
GEN|48|8|When Israel saw the sons of Joseph, he asked, "Who are these?"
GEN|48|9|"They are the sons God has given me here," Joseph said to his father. Then Israel said, "Bring them to me so I may bless them."
GEN|48|10|Now Israel's eyes were failing because of old age, and he could hardly see. So Joseph brought his sons close to him, and his father kissed them and embraced them.
GEN|48|11|Israel said to Joseph, "I never expected to see your face again, and now God has allowed me to see your children too."
GEN|48|12|Then Joseph removed them from Israel's knees and bowed down with his face to the ground.
GEN|48|13|And Joseph took both of them, Ephraim on his right toward Israel's left hand and Manasseh on his left toward Israel's right hand, and brought them close to him.
GEN|48|14|But Israel reached out his right hand and put it on Ephraim's head, though he was the younger, and crossing his arms, he put his left hand on Manasseh's head, even though Manasseh was the firstborn.
GEN|48|15|Then he blessed Joseph and said, "May the God before whom my fathers Abraham and Isaac walked, the God who has been my shepherd all my life to this day,
GEN|48|16|the Angel who has delivered me from all harm -may he bless these boys. May they be called by my name and the names of my fathers Abraham and Isaac, and may they increase greatly upon the earth."
GEN|48|17|When Joseph saw his father placing his right hand on Ephraim's head he was displeased; so he took hold of his father's hand to move it from Ephraim's head to Manasseh's head.
GEN|48|18|Joseph said to him, "No, my father, this one is the firstborn; put your right hand on his head."
GEN|48|19|But his father refused and said, "I know, my son, I know. He too will become a people, and he too will become great. Nevertheless, his younger brother will be greater than he, and his descendants will become a group of nations."
GEN|48|20|He blessed them that day and said, "In your name will Israel pronounce this blessing: 'May God make you like Ephraim and Manasseh.'" So he put Ephraim ahead of Manasseh.
GEN|48|21|Then Israel said to Joseph, "I am about to die, but God will be with you and take you back to the land of your fathers.
GEN|48|22|And to you, as one who is over your brothers, I give the ridge of land I took from the Amorites with my sword and my bow."
GEN|49|1|Then Jacob called for his sons and said: "Gather around so I can tell you what will happen to you in days to come.
GEN|49|2|"Assemble and listen, sons of Jacob; listen to your father Israel.
GEN|49|3|"Reuben, you are my firstborn, my might, the first sign of my strength, excelling in honor, excelling in power.
GEN|49|4|Turbulent as the waters, you will no longer excel, for you went up onto your father's bed, onto my couch and defiled it.
GEN|49|5|"Simeon and Levi are brothers- their swords are weapons of violence.
GEN|49|6|Let me not enter their council, let me not join their assembly, for they have killed men in their anger and hamstrung oxen as they pleased.
GEN|49|7|Cursed be their anger, so fierce, and their fury, so cruel! I will scatter them in Jacob and disperse them in Israel.
GEN|49|8|"Judah, your brothers will praise you; your hand will be on the neck of your enemies; your father's sons will bow down to you.
GEN|49|9|You are a lion's cub, O Judah; you return from the prey, my son. Like a lion he crouches and lies down, like a lioness-who dares to rouse him?
GEN|49|10|The scepter will not depart from Judah, nor the ruler's staff from between his feet, until he comes to whom it belongs and the obedience of the nations is his.
GEN|49|11|He will tether his donkey to a vine, his colt to the choicest branch; he will wash his garments in wine, his robes in the blood of grapes.
GEN|49|12|His eyes will be darker than wine, his teeth whiter than milk.
GEN|49|13|"Zebulun will live by the seashore and become a haven for ships; his border will extend toward Sidon.
GEN|49|14|"Issachar is a rawboned donkey lying down between two saddlebags.
GEN|49|15|When he sees how good is his resting place and how pleasant is his land, he will bend his shoulder to the burden and submit to forced labor.
GEN|49|16|"Dan will provide justice for his people as one of the tribes of Israel.
GEN|49|17|Dan will be a serpent by the roadside, a viper along the path, that bites the horse's heels so that its rider tumbles backward.
GEN|49|18|"I look for your deliverance, O LORD.
GEN|49|19|"Gad will be attacked by a band of raiders, but he will attack them at their heels.
GEN|49|20|"Asher's food will be rich; he will provide delicacies fit for a king.
GEN|49|21|"Naphtali is a doe set free that bears beautiful fawns.
GEN|49|22|"Joseph is a fruitful vine, a fruitful vine near a spring, whose branches climb over a wall.
GEN|49|23|With bitterness archers attacked him; they shot at him with hostility.
GEN|49|24|But his bow remained steady, his strong arms stayed limber, because of the hand of the Mighty One of Jacob, because of the Shepherd, the Rock of Israel,
GEN|49|25|because of your father's God, who helps you, because of the Almighty, who blesses you with blessings of the heavens above, blessings of the deep that lies below, blessings of the breast and womb.
GEN|49|26|Your father's blessings are greater than the blessings of the ancient mountains, than the bounty of the age-old hills. Let all these rest on the head of Joseph, on the brow of the prince among his brothers.
GEN|49|27|"Benjamin is a ravenous wolf; in the morning he devours the prey, in the evening he divides the plunder."
GEN|49|28|All these are the twelve tribes of Israel, and this is what their father said to them when he blessed them, giving each the blessing appropriate to him.
GEN|49|29|Then he gave them these instructions: "I am about to be gathered to my people. Bury me with my fathers in the cave in the field of Ephron the Hittite,
GEN|49|30|the cave in the field of Machpelah, near Mamre in Canaan, which Abraham bought as a burial place from Ephron the Hittite, along with the field.
GEN|49|31|There Abraham and his wife Sarah were buried, there Isaac and his wife Rebekah were buried, and there I buried Leah.
GEN|49|32|The field and the cave in it were bought from the Hittites. "
GEN|49|33|When Jacob had finished giving instructions to his sons, he drew his feet up into the bed, breathed his last and was gathered to his people.
GEN|50|1|Joseph threw himself upon his father and wept over him and kissed him.
GEN|50|2|Then Joseph directed the physicians in his service to embalm his father Israel. So the physicians embalmed him,
GEN|50|3|taking a full forty days, for that was the time required for embalming. And the Egyptians mourned for him seventy days.
GEN|50|4|When the days of mourning had passed, Joseph said to Pharaoh's court, "If I have found favor in your eyes, speak to Pharaoh for me. Tell him,
GEN|50|5|'My father made me swear an oath and said, "I am about to die; bury me in the tomb I dug for myself in the land of Canaan." Now let me go up and bury my father; then I will return.'"
GEN|50|6|Pharaoh said, "Go up and bury your father, as he made you swear to do."
GEN|50|7|So Joseph went up to bury his father. All Pharaoh's officials accompanied him-the dignitaries of his court and all the dignitaries of Egypt-
GEN|50|8|besides all the members of Joseph's household and his brothers and those belonging to his father's household. Only their children and their flocks and herds were left in Goshen.
GEN|50|9|Chariots and horsemen also went up with him. It was a very large company.
GEN|50|10|When they reached the threshing floor of Atad, near the Jordan, they lamented loudly and bitterly; and there Joseph observed a seven-day period of mourning for his father.
GEN|50|11|When the Canaanites who lived there saw the mourning at the threshing floor of Atad, they said, "The Egyptians are holding a solemn ceremony of mourning." That is why that place near the Jordan is called Abel Mizraim.
GEN|50|12|So Jacob's sons did as he had commanded them:
GEN|50|13|They carried him to the land of Canaan and buried him in the cave in the field of Machpelah, near Mamre, which Abraham had bought as a burial place from Ephron the Hittite, along with the field.
GEN|50|14|After burying his father, Joseph returned to Egypt, together with his brothers and all the others who had gone with him to bury his father.
GEN|50|15|When Joseph's brothers saw that their father was dead, they said, "What if Joseph holds a grudge against us and pays us back for all the wrongs we did to him?"
GEN|50|16|So they sent word to Joseph, saying, "Your father left these instructions before he died:
GEN|50|17|'This is what you are to say to Joseph: I ask you to forgive your brothers the sins and the wrongs they committed in treating you so badly.' Now please forgive the sins of the servants of the God of your father." When their message came to him, Joseph wept.
GEN|50|18|His brothers then came and threw themselves down before him. "We are your slaves," they said.
GEN|50|19|But Joseph said to them, "Don't be afraid. Am I in the place of God?
GEN|50|20|You intended to harm me, but God intended it for good to accomplish what is now being done, the saving of many lives.
GEN|50|21|So then, don't be afraid. I will provide for you and your children." And he reassured them and spoke kindly to them.
GEN|50|22|Joseph stayed in Egypt, along with all his father's family. He lived a hundred and ten years
GEN|50|23|and saw the third generation of Ephraim's children. Also the children of Makir son of Manasseh were placed at birth on Joseph's knees.
GEN|50|24|Then Joseph said to his brothers, "I am about to die. But God will surely come to your aid and take you up out of this land to the land he promised on oath to Abraham, Isaac and Jacob."
GEN|50|25|And Joseph made the sons of Israel swear an oath and said, "God will surely come to your aid, and then you must carry my bones up from this place."
GEN|50|26|So Joseph died at the age of a hundred and ten. And after they embalmed him, he was placed in a coffin in Egypt.
