ZECH|1|1|in mense octavo in anno secundo Darii factum est verbum Domini ad Zacchariam filium Barachiae filium Addo prophetam dicens
ZECH|1|2|iratus est Dominus super patres vestros iracundia
ZECH|1|3|et dices ad eos haec dicit Dominus exercituum convertimini ad me ait Dominus exercituum et convertar ad vos dicit Dominus exercituum
ZECH|1|4|ne sitis sicut patres vestri ad quos clamabant prophetae priores dicentes haec dicit Dominus exercituum convertimini de viis vestris malis et cogitationibus vestris pessimis et non audierunt neque adtenderunt ad me dicit Dominus
ZECH|1|5|patres vestri ubi sunt et prophetae numquid in sempiternum vivent
ZECH|1|6|verumtamen verba mea et legitima mea quae mandavi servis meis prophetis numquid non conprehenderunt patres vestros et conversi sunt et dixerunt sicut cogitavit Dominus exercituum facere nobis secundum vias nostras et secundum adinventiones nostras fecit nobis
ZECH|1|7|in die vicesima et quarta undecimo mense sabath in anno secundo Darii factum est verbum Domini ad Zacchariam filium Barachiae filium Addo prophetam dicens
ZECH|1|8|vidi per noctem et ecce vir ascendens super equum rufum et ipse stabat inter myrteta quae erant in profundo et post eum equi rufi varii et albi
ZECH|1|9|et dixi quid sunt isti domine mi et dixit ad me angelus qui loquebatur in me ego ostendam tibi quid sint haec
ZECH|1|10|et respondit vir qui stabat inter myrteta et dixit isti sunt quos misit Dominus ut perambularent terram
ZECH|1|11|et responderunt angelo Domini qui stabat inter myrteta et dixerunt perambulavimus terram et ecce omnis terra habitatur et quiescit
ZECH|1|12|et respondit angelus Domini et dixit Domine exercituum usquequo tu non misereberis Hierusalem et urbium Iuda quibus iratus es iste septuagesimus annus est
ZECH|1|13|et respondit Dominus angelo qui loquebatur in me verba bona verba consolatoria
ZECH|1|14|et dixit ad me angelus qui loquebatur in me clama dicens haec dicit Dominus exercituum zelatus sum Hierusalem et Sion zelo magno
ZECH|1|15|et ira magna ego irascor super gentes opulentas quia ego iratus sum parum ipsi vero adiuverunt in malum
ZECH|1|16|propterea haec dicit Dominus revertar ad Hierusalem in misericordiis domus mea aedificabitur in ea ait Dominus exercituum et perpendiculum extendetur super Hierusalem
ZECH|1|17|adhuc clama dicens haec dicit Dominus exercituum adhuc affluent civitates meae bonis et consolabitur Dominus adhuc Sion et eliget adhuc Hierusalem
ZECH|1|18|et levavi oculos meos et vidi et ecce quattuor cornua
ZECH|1|19|et dixi ad angelum qui loquebatur in me quid sunt haec et dixit ad me haec sunt cornua quae ventilaverunt Iudam et Israhel et Hierusalem
ZECH|1|20|et ostendit mihi Dominus quattuor fabros
ZECH|1|21|et dixi quid isti veniunt facere qui ait dicens haec sunt cornua quae ventilaverunt Iudam per singulos viros et nemo eorum levavit caput suum et venerunt isti deterrere ea ut deiciant cornua gentium quae levaverunt cornu super terram Iuda ut dispergerent eam
ZECH|2|1|et levavi oculos meos et vidi et ecce vir et in manu eius funiculus mensorum
ZECH|2|2|et dixi quo tu vadis et dixit ad me ut metiar Hierusalem et videam quanta sit latitudo eius et quanta longitudo eius
ZECH|2|3|et ecce angelus qui loquebatur in me egrediebatur et angelus alius egrediebatur in occursum eius
ZECH|2|4|et dixit ad eum curre loquere ad puerum istum dicens absque muro habitabitur Hierusalem prae multitudine hominum et iumentorum in medio eius
ZECH|2|5|et ego ero ei ait Dominus murus ignis in circuitu et in gloria ero in medio eius
ZECH|2|6|o o fugite de terra aquilonis dicit Dominus quoniam in quattuor ventos caeli dispersi vos dicit Dominus
ZECH|2|7|o Sion fuge quae habitas apud filiam Babylonis
ZECH|2|8|quia haec dicit Dominus exercituum post gloriam misit me ad gentes quae spoliaverunt vos qui enim tetigerit vos tangit pupillam oculi eius
ZECH|2|9|quia ecce ego levo manum meam super eos et erunt praedae his qui serviebant sibi et cognoscetis quia Dominus exercituum misit me
ZECH|2|10|lauda et laetare filia Sion quia ecce ego venio et habitabo in medio tui ait Dominus
ZECH|2|11|et adplicabuntur gentes multae ad Dominum in die illa et erunt mihi in populum et habitabo in medio tui et scies quia Dominus exercituum misit me ad te
ZECH|2|12|et possidebit Dominus Iudam partem suam in terra sanctificata et eliget adhuc Hierusalem
ZECH|2|13|sileat omnis caro a facie Domini quia consurrexit de habitaculo sancto suo
ZECH|3|1|et ostendit mihi Iesum sacerdotem magnum stantem coram angelo Domini et Satan stabat a dextris eius ut adversaretur ei
ZECH|3|2|et dixit Dominus ad Satan increpet Dominus in te Satan et increpet Dominus in te qui elegit Hierusalem numquid non iste torris est erutus de igne
ZECH|3|3|et Iesus erat indutus vestibus sordidis et stabat ante faciem angeli
ZECH|3|4|qui respondit et ait ad eos qui stabant coram se dicens auferte vestimenta sordida ab eo et dixit ad eum ecce abstuli a te iniquitatem tuam et indui te mutatoriis
ZECH|3|5|et dixit ponite cidarim mundam super caput eius et posuerunt cidarim mundam super caput eius et induerunt eum vestibus et angelus Domini stabat
ZECH|3|6|et contestabatur angelus Domini Iesum dicens
ZECH|3|7|haec dicit Dominus exercituum si in viis meis ambulaveris et custodiam meam custodieris tu quoque iudicabis domum meam et custodies atria mea et dabo tibi ambulantes de his qui nunc hic adsistunt
ZECH|3|8|audi Iesu sacerdos magne tu et amici tui qui habitant coram te quia viri portendentes sunt ecce enim ego adducam servum meum orientem
ZECH|3|9|quia ecce lapis quem dedi coram Iesu super lapidem unum septem oculi sunt ecce ego celabo sculpturam eius ait Dominus exercituum et auferam iniquitatem terrae illius in die una
ZECH|3|10|in die illa dicit Dominus exercituum vocabit vir amicum suum subter vineam et subter ficum
ZECH|4|1|et reversus est angelus qui loquebatur in me et suscitavit me quasi virum qui suscitatur de somno suo
ZECH|4|2|et dixit ad me quid tu vides et dixi vidi et ecce candelabrum aureum totum et lampas eius super caput ipsius et septem lucernae eius super illud septem et septem infusoria lucernis quae erant super caput illius
ZECH|4|3|et duae olivae super illud una a dextris lampadis et una a sinistris eius
ZECH|4|4|et respondi et aio ad angelum qui loquebatur in me dicens quid sunt haec domine mi
ZECH|4|5|et respondit angelus qui loquebatur in me et dixit ad me numquid nescis quid sunt haec et dixi non domine mi
ZECH|4|6|et respondit et ait ad me dicens hoc est verbum Domini ad Zorobabel dicens non in exercitu nec in robore sed in spiritu meo dicit Dominus exercituum
ZECH|4|7|quis tu mons magne coram Zorobabel in planum et educet lapidem primarium et exaequabit gratiam gratiae eius
ZECH|4|8|et factum est verbum Domini ad me dicens
ZECH|4|9|manus Zorobabel fundaverunt domum istam et manus eius perficient eam et scietis quia Dominus exercituum misit me ad vos
ZECH|4|10|quis enim despexit dies parvos et laetabuntur et videbunt lapidem stagneum in manu Zorobabel septem isti oculi Domini qui discurrunt in universa terra
ZECH|4|11|et respondi et dixi ad eum quid sunt duae olivae istae ad dextram candelabri et ad sinistram eius
ZECH|4|12|et respondi secundo et dixi ad eum quid sunt duae spicae olivarum quae sunt iuxta duo rostra aurea in quibus sunt suffusoria ex auro
ZECH|4|13|et ait ad me dicens numquid nescis quid sunt haec et dixi non domine
ZECH|4|14|et dixit isti duo filii olei qui adsistunt Dominatori universae terrae
ZECH|5|1|et conversus sum et levavi oculos meos et vidi et ecce volumen volans
ZECH|5|2|et dixit ad me quid tu vides et dixi ego video volumen volans longitudo eius viginti cubitorum et latitudo eius decem cubitorum
ZECH|5|3|et dixit ad me haec est maledictio quae egreditur super faciem omnis terrae quia omnis fur sicut ibi scriptum est iudicabitur et omnis iurans ex hoc similiter iudicabitur
ZECH|5|4|educam illud dicit Dominus exercituum et veniet ad domum furis et ad domum iurantis in nomine meo mendaciter et commorabitur in medio domus eius et consumet eam et ligna eius et lapides eius
ZECH|5|5|et egressus est angelus qui loquebatur in me et dixit ad me leva oculos tuos et vide quid est hoc quod egreditur
ZECH|5|6|et dixi quidnam est et ait haec est amphora egrediens et dixit haec est oculus eorum in universa terra
ZECH|5|7|et ecce talentum plumbi portabatur et ecce mulier una sedens in medio amphorae
ZECH|5|8|et dixit haec est impietas et proiecit eam in medio amphorae et misit massam plumbeam in os eius
ZECH|5|9|et levavi oculos meos et vidi et ecce duae mulieres egredientes et spiritus in alis earum et habebant alas quasi alas milvi et levaverunt amphoram inter terram et caelum
ZECH|5|10|et dixi ad angelum qui loquebatur in me quo istae deferunt amphoram
ZECH|5|11|et dixit ad me ut aedificetur ei domus in terra Sennaar et stabiliatur et ponatur ibi super basem suam
ZECH|6|1|et conversus sum et levavi oculos meos et vidi et ecce quattuor quadrigae egredientes de medio duorum montium et montes montes aerei
ZECH|6|2|in quadriga prima equi rufi et in quadriga secunda equi nigri
ZECH|6|3|et in quadriga tertia equi albi et in quadriga quarta equi varii fortes
ZECH|6|4|et respondi et dixi ad angelum qui loquebatur in me quid sunt haec domine mi
ZECH|6|5|et respondit angelus et ait ad me isti sunt quattuor venti caeli qui egrediuntur ut stent coram Dominatore omnis terrae
ZECH|6|6|in quo erant equi nigri egrediebantur in terra aquilonis et albi egressi sunt post eos et varii egressi sunt ad terram austri
ZECH|6|7|qui autem erant robustissimi exierunt et quaerebant ire et discurrere per omnem terram et dixit ite perambulate terram et perambulaverunt terram
ZECH|6|8|et vocavit me et locutus est ad me dicens ecce qui egrediuntur in terram aquilonis requiescere fecerunt spiritum meum in terra aquilonis
ZECH|6|9|et factum est verbum Domini ad me dicens
ZECH|6|10|sume a transmigratione ab Oldai et a Tobia et ab Idaia et venies tu in die illa et intrabis domum Iosiae filii Sofoniae qui venerunt de Babylone
ZECH|6|11|et sumes argentum et aurum et facies coronas et pones in capite Iesu filii Iosedech sacerdotis magni
ZECH|6|12|et loqueris ad eum dicens haec ait Dominus exercituum dicens ecce vir Oriens nomen eius et subter eum orietur et aedificabit templum Domino
ZECH|6|13|et ipse extruet templum Domino et ipse portabit gloriam et sedebit et dominabitur super solio suo et erit sacerdos super solio suo et consilium pacis erit inter duos illos
ZECH|6|14|et coronae erunt Helem et Tobiae et Idaiae et Hen filio Sofoniae memoriale in templo Domini
ZECH|6|15|et qui procul sunt venient et aedificabunt in templo Domini et scietis quia Dominus exercituum misit me ad vos erit autem hoc si auditu audieritis vocem Domini Dei vestri
ZECH|7|1|et factum est in anno quarto Darii regis factum est verbum Domini ad Zacchariam in quarta mensis noni qui est casleu
ZECH|7|2|et miserunt ad domum Dei Sarasar et Rogomelech et viri qui erant cum eo ad deprecandam faciem Domini
ZECH|7|3|ut dicerent sacerdotibus domus Domini exercituum et prophetis loquentes numquid flendum mihi est in mense quinto vel sanctificare me debeo sicuti feci iam multis annis
ZECH|7|4|et factum est verbum Domini exercituum ad me dicens
ZECH|7|5|loquere ad omnem populum terrae et ad sacerdotes dicens cum ieiunaretis et plangeretis in quinto et septimo per hos septuaginta annos numquid ieiunium ieiunastis mihi
ZECH|7|6|et cum comedistis et cum bibistis numquid non vobis comedistis et vobismet ipsis bibistis
ZECH|7|7|numquid non sunt verba quae locutus est Dominus in manu prophetarum priorum cum adhuc Hierusalem habitaretur et esset opulenta ipsa et urbes in circuitu eius et ad austrum et in campestribus habitaretur
ZECH|7|8|et factum est verbum Domini ad Zacchariam dicens
ZECH|7|9|haec ait Dominus exercituum dicens iudicium verum iudicate et misericordiam et miserationes facite unusquisque cum fratre suo
ZECH|7|10|et viduam et pupillum et advenam et pauperem nolite calumniari et malum vir fratri suo non cogitet in corde suo
ZECH|7|11|et noluerunt adtendere et verterunt scapulam recedentem et aures suas adgravaverunt ne audirent
ZECH|7|12|et cor suum posuerunt adamantem ne audirent legem et verba quae misit Dominus exercituum in spiritu suo per manum prophetarum priorum et facta est indignatio magna a Domino exercituum
ZECH|7|13|et factum est sicut locutus est et non audierunt sic clamabunt et non exaudiam dicit Dominus exercituum
ZECH|7|14|et dispersi eos per omnia regna quae nesciunt et terra desolata est ab eis eo quod non esset transiens et revertens et posuerunt terram desiderabilem in desertum
ZECH|8|1|et factum est verbum Domini exercituum dicens
ZECH|8|2|haec dicit Dominus exercituum zelatus sum Sion zelo magno et indignatione magna zelatus sum eam
ZECH|8|3|haec dicit Dominus exercituum reversus sum ad Sion et habitabo in medio Hierusalem et vocabitur Hierusalem civitas veritatis et mons Domini exercituum mons sanctificatus
ZECH|8|4|haec dicit Dominus exercituum adhuc habitabunt senes et anus in plateis Hierusalem et viri baculus in manu eius prae multitudine dierum
ZECH|8|5|et plateae civitatis conplebuntur infantibus et puellis ludentibus in plateis eius
ZECH|8|6|haec dicit Dominus exercituum si difficile videbitur in oculis reliquiarum populi huius in diebus illis numquid in oculis meis difficile erit dicit Dominus exercituum
ZECH|8|7|haec dicit Dominus exercituum ecce ego salvabo populum meum de terra orientis et de terra occasus solis
ZECH|8|8|et adducam eos et habitabunt in medio Hierusalem et erunt mihi in populum et ego ero eis in Deum in veritate et iustitia
ZECH|8|9|haec dicit Dominus exercituum confortentur manus vestrae qui auditis in diebus his sermones istos per os prophetarum in die qua fundata est domus Domini exercituum ut templum aedificaretur
ZECH|8|10|siquidem ante dies illos merces hominum non erat nec merces iumentorum erat neque introeunti et exeunti erat pax prae tribulatione et dimisi omnes homines unumquemque contra proximum suum
ZECH|8|11|nunc autem non iuxta dies priores ego faciam reliquiis populi huius dicit Dominus exercituum
ZECH|8|12|sed semen pacis erit vinea dabit fructum suum et terra dabit germen suum et caeli dabunt rorem suum et possidere faciam reliquias populi huius universa haec
ZECH|8|13|et erit sicut eratis maledictio in gentibus domus Iuda et domus Israhel sic salvabo vos et eritis benedictio nolite timere confortentur manus vestrae
ZECH|8|14|quia haec dicit Dominus exercituum sicut cogitavi ut adfligerem vos cum ad iracundiam provocassent patres vestri me dicit Dominus
ZECH|8|15|et non sum misertus sic conversus cogitavi in diebus istis ut benefaciam Hierusalem et domui Iuda nolite timere
ZECH|8|16|haec sunt ergo verba quae facietis loquimini veritatem unusquisque cum proximo suo veritatem et iudicium pacis iudicate in portis vestris
ZECH|8|17|et unusquisque malum contra amicum suum ne cogitetis in cordibus vestris et iuramentum mendax ne diligatis omnia enim haec sunt quae odi dicit Dominus
ZECH|8|18|et factum est verbum Domini exercituum ad me dicens
ZECH|8|19|haec dicit Dominus exercituum ieiunium quarti et ieiunium quinti et ieiunium septimi et ieiunium decimi erit domui Iuda in gaudium et in laetitiam et in sollemnitates praeclaras veritatem tantum et pacem diligite
ZECH|8|20|haec dicit Dominus exercituum usquequo veniant populi et habitent in civitatibus multis
ZECH|8|21|et vadant habitatores unus ad alterum dicentes eamus et deprecemur faciem Domini et quaeramus Dominum exercituum vadam etiam ego
ZECH|8|22|et venient populi multi et gentes robustae ad quaerendum Dominum exercituum in Hierusalem et deprecandam faciem Domini
ZECH|8|23|haec dicit Dominus exercituum in diebus illis in quibus adprehendent decem homines ex omnibus linguis gentium et adprehendent fimbriam viri iudaei dicentes ibimus vobiscum audivimus enim quoniam Deus vobiscum est
ZECH|9|1|onus verbi Domini in terra Adrach et Damasci requiei eius quia Domini est oculus hominis et omnium tribuum Israhel
ZECH|9|2|Emath quoque in terminis eius et Tyrus et Sidon adsumpserunt quippe sibi sapientiam valde
ZECH|9|3|et aedificavit Tyrus munitionem suam et coacervavit argentum quasi humum et aurum ut lutum platearum
ZECH|9|4|ecce Dominus possidebit eam et percutiet in mari fortitudinem eius et haec igni devorabitur
ZECH|9|5|videbit Ascalon et timebit et Gaza et dolebit nimis et Accaron quoniam confusa est spes eius et peribit rex de Gaza et Ascalon non habitabitur
ZECH|9|6|et sedebit separator in Azoto et disperdam superbiam Philisthinorum
ZECH|9|7|et auferam sanguinem eius de ore eius et abominationes eius de medio dentium eius et relinquetur etiam ipse Deo nostro et erit quasi dux in Iuda et Accaron quasi Iebuseus
ZECH|9|8|et circumdabo domum meam ex his qui militant mihi euntes et revertentes et non transibit super eos ultra exactor quia nunc vidi in oculis meis
ZECH|9|9|exulta satis filia Sion iubila filia Hierusalem ecce rex tuus veniet tibi iustus et salvator ipse pauper et ascendens super asinum et super pullum filium asinae
ZECH|9|10|et disperdam quadrigam ex Ephraim et equum de Hierusalem et dissipabitur arcus belli et loquetur pacem gentibus et potestas eius a mari usque ad mare et a fluminibus usque ad fines terrae
ZECH|9|11|tu quoque in sanguine testamenti tui emisisti vinctos tuos de lacu in quo non est aqua
ZECH|9|12|convertimini ad munitionem vincti spei hodie quoque adnuntians duplicia reddam tibi
ZECH|9|13|quoniam extendi mihi Iudam quasi arcum implevi Ephraim et suscitabo filios tuos Sion super filios tuos Graecia et ponam te quasi gladium fortium
ZECH|9|14|et Dominus Deus super eos videbitur et exibit ut fulgur iaculum eius et Dominus Deus in tuba canet et vadet in turbine austri
ZECH|9|15|Dominus exercituum proteget eos et devorabunt et subicient lapidibus fundae et bibentes inebriabuntur quasi vino et replebuntur ut fialae et quasi cornua altaris
ZECH|9|16|et salvabit eos Dominus Deus eorum in die illa ut gregem populi sui quia lapides sancti elevantur super terram eius
ZECH|9|17|quid enim bonum eius est et quid pulchrum eius nisi frumentum electorum et vinum germinans virgines
ZECH|10|1|petite a Domino pluviam in tempore serotino et Dominus faciet nives et pluviam imbris dabit eis singulis herbam in agro
ZECH|10|2|quia simulacra locuta sunt inutile et divini viderunt mendacium et somniatores frustra locuti sunt vane consolabantur idcirco abducti sunt quasi grex adfligentur quia non est eis pastor
ZECH|10|3|super pastores iratus est furor meus et super hircos visitabo quia visitavit Dominus exercituum gregem suum domum Iuda et posuit eos quasi equum gloriae suae in bello
ZECH|10|4|ex ipso angulus ex ipso paxillus ex ipso arcus proelii ex ipso egredietur omnis exactor simul
ZECH|10|5|et erunt quasi fortes conculcantes lutum viarum in proelio et bellabunt quia Dominus cum eis et confundentur ascensores equorum
ZECH|10|6|et confortabo domum Iuda et domum Ioseph salvabo et convertam eos quia miserebor eorum et erunt sicut fuerunt quando non proieceram eos ego enim Dominus Deus eorum et exaudiam eos
ZECH|10|7|et erunt quasi fortes Ephraim et laetabitur cor eorum quasi a vino et filii eorum videbunt et laetabuntur et exultabit cor eorum in Domino
ZECH|10|8|sibilabo eis et congregabo illos quia redemi eos et multiplicabo eos sicut ante fuerant multiplicati
ZECH|10|9|et seminabo eos in populis et de longe recordabuntur mei et vivent cum filiis suis et revertentur
ZECH|10|10|et reducam eos de terra Aegypti et de Assyriis congregabo eos et ad terram Galaad et Libani adducam eos et non invenietur eis locus
ZECH|10|11|et transibit in maris freto et percutiet in mari fluctus et confundentur omnia profunda Fluminis et humiliabitur superbia Assur et sceptrum Aegypti recedet
ZECH|10|12|confortabo eos in Domino et in nomine eius ambulabunt dicit Dominus
ZECH|11|1|aperi Libane portas tuas et comedat ignis cedros tuas
ZECH|11|2|ulula abies quia cecidit cedrus quoniam magnifici vastati sunt ululate quercus Basan quoniam succisus est saltus munitus
ZECH|11|3|vox ululatus pastorum quia vastata est magnificentia eorum vox rugitus leonum quoniam vastata est superbia Iordanis
ZECH|11|4|haec dicit Dominus Deus meus pasce pecora occisionis
ZECH|11|5|quae qui possederant occidebant et non dolebant et vendebant ea dicentes benedictus Dominus divites facti sumus et pastores eorum non parcebant eis
ZECH|11|6|et ego non parcam ultra super habitantes terram dicit Dominus ecce ego tradam homines unumquemque in manu proximi sui et in manu regis sui et concident terram et non eruam de manu eorum
ZECH|11|7|et pascam pecus occisionis propter hoc o pauperes gregis et adsumpsi mihi duas virgas unam vocavi Decorem et alteram vocavi Funiculos et pavi gregem
ZECH|11|8|et succidi tres pastores in mense uno et contracta est anima mea in eis siquidem anima eorum variavit in me
ZECH|11|9|et dixi non pascam vos quod moritur moriatur et quod succiditur succidatur et reliqui vorent unusquisque carnem proximi sui
ZECH|11|10|et tuli virgam meam quae vocabatur Decus et abscidi eam ut irritum facerem foedus meum quod percussi cum omnibus populis
ZECH|11|11|et in irritum deductum est in die illa et cognoverunt sic pauperes gregis qui custodiunt mihi quia verbum Domini est
ZECH|11|12|et dixi ad eos si bonum est in oculis vestris adferte mercedem meam et si non quiescite et adpenderunt mercedem meam triginta argenteos
ZECH|11|13|et dixit Dominus ad me proice illud ad statuarium decorum pretium quod adpretiatus sum ab eis et tuli triginta argenteos et proieci illos in domo Domini ad statuarium
ZECH|11|14|et praecidi virgam meam secundam quae appellabatur Funiculus ut dissolverem germanitatem inter Iudam et inter Israhel
ZECH|11|15|et dixit Dominus ad me adhuc sume tibi vasa pastoris stulti
ZECH|11|16|quia ecce ego suscitabo pastorem in terra qui derelicta non visitabit dispersum non quaeret et contritum non sanabit et id quod stat non enutriet et carnes pinguium comedet et ungulas eorum dissolvet
ZECH|11|17|o pastor et idolum derelinquens gregem gladius super brachium eius et super oculum dextrum eius brachium eius ariditate siccabitur et oculus dexter eius tenebrescens obscurabitur
ZECH|12|1|onus verbi Domini super Israhel dixit Dominus extendens caelum et fundans terram et fingens spiritum hominis in eo
ZECH|12|2|ecce ego ponam Hierusalem superliminare crapulae omnibus populis in circuitu sed et Iuda erit in obsidione contra Hierusalem
ZECH|12|3|et erit in die illa ponam Hierusalem lapidem oneris cunctis populis omnes qui levabunt eam concisione lacerabuntur et colligentur adversum eam omnia regna terrae
ZECH|12|4|in die illa dicit Dominus percutiam omnem equum in stuporem et ascensorem eius in amentiam et super domum Iuda aperiam oculos meos et omnem equum populorum percutiam in caecitate
ZECH|12|5|et dicent duces Iuda in corde suo confortentur mihi habitatores Hierusalem in Domino exercituum Deo eorum
ZECH|12|6|in die illo ponam duces Iuda sicut caminum ignis in lignis et sicut facem ignis in faeno et devorabunt ad dextram et ad sinistram omnes populos in circuitu et habitabitur Hierusalem rursum in loco suo in Hierusalem
ZECH|12|7|et salvabit Dominus tabernacula Iuda sicut in principio ut non magnifice glorietur domus David et gloria habitantium Hierusalem contra Iudam
ZECH|12|8|in die illo proteget Dominus habitatores Hierusalem et erit qui offenderit ex eis in die illa quasi David et domus David quasi Dei sicut angelus Domini in conspectu eius
ZECH|12|9|et erit in die illa quaeram conterere omnes gentes quae veniunt contra Hierusalem
ZECH|12|10|et effundam super domum David et super habitatores Hierusalem spiritum gratiae et precum et aspicient ad me quem confixerunt et plangent eum planctu quasi super unigenitum et dolebunt super eum ut doleri solet in morte primogeniti
ZECH|12|11|in die illa magnus erit planctus in Hierusalem sicut planctus Adadremmon in campo Mageddon
ZECH|12|12|et planget terra familiae et familiae seorsum familiae domus David seorsum et mulieres eorum seorsum
ZECH|12|13|familiae domus Nathan seorsum et mulieres eorum seorsum familiae domus Levi seorsum et mulieres eorum seorsum familiae Semei seorsum et mulieres eorum seorsum
ZECH|12|14|omnes familiae reliquae familiae et familiae seorsum et mulieres eorum seorsum
ZECH|13|1|in die illa erit fons patens domus David et habitantibus Hierusalem in ablutionem peccatoris et menstruatae
ZECH|13|2|et erit in die illa dicit Dominus exercituum disperdam nomina idolorum de terra et non memorabuntur ultra et prophetas et spiritum inmundum auferam de terra
ZECH|13|3|et erit cum prophetaverit quispiam ultra dicent ei pater eius et mater eius qui genuerunt eum non vives quia mendacium locutus es in nomine Domini et configent eum pater eius et mater eius genitores eius cum prophetaverit
ZECH|13|4|et erit in die illa confundentur prophetae unusquisque ex visione sua cum prophetaverit nec operientur pallio saccino ut mentiantur
ZECH|13|5|sed dicet non sum propheta homo agricola ego sum quoniam Adam exemplum meum ab adulescentia mea
ZECH|13|6|et dicetur ei quid sunt plagae istae in medio manuum tuarum et dicet his plagatus sum in domo eorum qui diligebant me
ZECH|13|7|framea suscitare super pastorem meum et super virum coherentem mihi dicit Dominus exercituum percute pastorem et dispergantur oves et convertam manum meam ad parvulos
ZECH|13|8|et erunt in omni terra dicit Dominus partes duae in ea disperdentur et deficient et tertia pars relinquetur in ea
ZECH|13|9|et ducam tertiam partem per ignem et uram eas sicut uritur argentum et probabo eos sicut probatur aurum ipse vocabit nomen meum et ego exaudiam eum dicam populus meus es et ipse dicet Dominus Deus meus
ZECH|14|1|ecce dies veniunt Domini et dividentur spolia tua in medio tui
ZECH|14|2|et congregabo omnes gentes ad Hierusalem in proelium et capietur civitas et vastabuntur domus et mulieres violabuntur et egredietur media pars civitatis in captivitatem et reliquum populi non auferetur ex urbe
ZECH|14|3|et egredietur Dominus et proeliabitur contra gentes illas sicut proeliatus est in die certaminis
ZECH|14|4|et stabunt pedes eius in die illa super montem Olivarum qui est contra Hierusalem ad orientem et scindetur mons Olivarum ex media parte sui ad orientem et occidentem praerupto grandi valde et separabitur medium montis ad aquilonem et medium eius ad meridiem
ZECH|14|5|et fugietis ad vallem montium meorum quoniam coniungetur vallis montium usque ad proximum et fugietis sicut fugistis a facie terraemotus in diebus Oziae regis Iuda et veniet Dominus Deus meus omnesque sancti cum eo
ZECH|14|6|et erit in die illa non erit lux sed frigus et gelu
ZECH|14|7|et erit dies una quae nota est Domino non dies neque nox et in tempore vesperae erit lux
ZECH|14|8|et erit in die illa exibunt aquae vivae de Hierusalem medium earum ad mare orientale et medium earum ad mare novissimum in aestate et in hieme erunt
ZECH|14|9|et erit Dominus rex super omnem terram in die illa erit Dominus unus et erit nomen eius unum
ZECH|14|10|et revertetur omnis terra usque ad desertum de colle Remmon ad austrum Hierusalem et exaltabitur et habitabit in loco suo a porta Beniamin usque ad locum portae Prioris usque ad portam Angulorum et a turre Ananehel usque ad torcularia regis
ZECH|14|11|et habitabunt in ea et anathema non erit amplius sed sedebit Hierusalem secura
ZECH|14|12|et haec erit plaga qua percutiet Dominus omnes gentes quae pugnaverunt adversus Hierusalem tabescet caro uniuscuiusque stantis super pedes suos et oculi eius contabescent in foraminibus suis et lingua eorum contabescet in ore suo
ZECH|14|13|in die illo erit tumultus Domini magnus in eis et adprehendet vir manum proximi sui et conseretur manus eius super manum proximi sui
ZECH|14|14|sed et Iudas pugnabit adversus Hierusalem et congregabuntur divitiae omnium gentium in circuitu aurum et argentum et vestes multae satis
ZECH|14|15|et sic erit ruina equi et muli cameli et asini et omnium iumentorum quae fuerint in castris illis sicut ruina haec
ZECH|14|16|et omnes qui reliqui fuerint de universis gentibus quae venerint contra Hierusalem ascendent ab anno in annum ut adorent regem Dominum exercituum et celebrent festivitatem tabernaculorum
ZECH|14|17|et erit qui non ascenderit de familiis terrae ad Hierusalem ut adoret regem Dominum exercituum non erit super eos imber
ZECH|14|18|quod si et familia Aegypti non ascenderit et non venerit nec super eos erit sed erit ruina qua percutiet Dominus omnes gentes quae non ascenderint ad celebrandam festivitatem tabernaculorum
ZECH|14|19|hoc erit peccatum Aegypti et hoc peccatum omnium gentium quae non ascenderint ad celebrandam festivitatem tabernaculorum
ZECH|14|20|in die illo erit quod super frenum equi est sanctum Domino et erunt lebetes in domo Domini quasi fialae coram altari
ZECH|14|21|et erit omnis lebes in Hierusalem et in Iuda sanctificatus Domino exercituum et venient omnes immolantes et sument ex eis et coquent in eis et non erit mercator ultra in domo Domini exercituum in die illo
