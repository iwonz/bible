RUTH|1|1|І сталось за часу, коли судді судили, то був голод у Краю. І пішов був чоловік з Юдиного Віфлеєму мешкати в моавських полях, він і жінка та двоє синів його.
RUTH|1|2|А ім'я тому чоловікові Елімелех, а ім'я жінці його Ноомі; і ім'я двох синів його Махлон і Кілйон, ефратяни з Віфлеєму Юдиного. І прийшли вони на моавські поля, та й залишилися.
RUTH|1|3|І помер Елімелех, муж Ноомі, і зосталася вона та два їхні сини.
RUTH|1|4|І взяли вони собі за жінок моавітянок, ім'я одній Орпа, а ім'я другій Рут. І сиділи вони там близько десяти літ.
RUTH|1|5|І повмирали й вони обоє, Махлон та Кілйон. І позосталася та жінка по двох дітях своїх та по чоловікові своєму.
RUTH|1|6|І встала вона та невістки її, і вернулися з моавських піль, бо почула на моавському полі, що Господь згадав про народ Свій, даючи їм хліба.
RUTH|1|7|І вийшла вона з того місця, де була там, та обидві невістки з нею, та й пішли дорогою, щоб вернутися до Юдиного краю.
RUTH|1|8|І сказала Ноомі до двох своїх невісток: Ідіть, верніться кожна до дому своєї матері. І нехай Господь зробить із вами милість, як ви зробили з померлими та зо мною.
RUTH|1|9|Нехай Господь дасть вам, і ви знайдете відпочинок кожна в домі свого мужа! І вона поцілувала їх, а вони підняли свій голос та плакали.
RUTH|1|10|І вони сказали до неї: Ні, з тобою ми вернемось до народу твого!
RUTH|1|11|А Ноомі сказала: Вертайтеся, дочки мої, чого ви підете зо мною? Чи я маю ще в утробі своїй синів, а вони стануть вам за чоловіків?
RUTH|1|12|Верніться, дочки мої, ідіть, бо я занадто стара, щоб бути для мужа. А коли б я й сказала: Маю надію, і коли б цієї ночі була з мужем, і також породила синів,
RUTH|1|13|чи ж ви чекали б їх, аж поки повиростають? Чи ж ви зв'язалися б з ними, щоб не бути замужем? Ні, дочки мої, бо мені значно гірше, як вам, бо Господня рука знайшла мене.
RUTH|1|14|І підняли вони голос свій, і заплакали ще. І поцілувала Орпа свою свекруху, а Рут пригорнулася до неї.
RUTH|1|15|І сказала Ноомі: Ось зовиця твоя вернулася до народу свого та до богів своїх, вернися й ти за зовицею своєю!
RUTH|1|16|А Рут відказала: Не силуй мене, щоб я покинула тебе, щоб я вернулася від тебе, бо куди підеш ти, туди піду й я, а де житимеш ти, там житиму й я. Народ твій буде мій народ, а Бог твій мій Бог.
RUTH|1|17|Де помреш ти, там помру й я, і там буду похована. Нехай Господь зробить мені так, і так нехай додасть, і тільки смерть розлучить мене з тобою.
RUTH|1|18|І побачила Ноомі, що вона настоює йти за нею, і перестала вговорювати її.
RUTH|1|19|І пішли вони вдвох, аж прийшли до Віфлеєму. І сталося, коли вони входили до Віфлеєму, то зашуміло все місто про них, і говорили: Чи це Ноомі?
RUTH|1|20|А вона сказала їм: Не кличте мене: Ноомі, кличте мене: Мара, бо велику гіркоту зробив мені Всемогутній.
RUTH|1|21|Я заможною пішла була, та порожньою вернув мене Господь. Чого кличете мене: Ноомі, коли Господь свідчив проти мене, а Всемогутній послав мені горе?
RUTH|1|22|І вернулася Ноомі та з нею моавітянка Рут, невістка її, що верталася з моавських піль. І прийшли вони до Віфлеєму на початку жнив ячменю.
RUTH|2|1|А Ноомі мала родича свого чоловіка, мужа багатого, з Елімелехового роду, а ім'я йому Боаз.
RUTH|2|2|І сказала моавітянка Рут до Ноомі: Піду но я на поле, і назбираю колосся за тим, у кого в очах знайду милість. А та їй сказала: Іди, моя дочко!
RUTH|2|3|І пішла вона, і прийшла та й збирала за женцями. А припадок навів її на ділянку поля Боаза, що з Елімелехового роду.
RUTH|2|4|Аж ось прийшов із Віфлеєму Боаз, та й сказав до женців: Господь з вами! А вони відказали йому: Нехай поблагословить тебе Господь!
RUTH|2|5|І сказав Боаз до слуги свого, поставленого над женцями: Чия це дівчина?
RUTH|2|6|І відповів той слуга, поставлений над женцями, і сказав: Дівчина моавітянка вона, що вернулася з Ноомі з моавських піль.
RUTH|2|7|А вона сказала: Нехай я збиратиму, та назбираю між снопами за женцями! І прийшла вона, і стала від самого ранку й аж дотепер; а вдома вона була мало.
RUTH|2|8|І сказав Боаз до Рут: Ото чуєш, дочко моя, не ходи збирати на іншому полі, і не йди звідси, і так пристань до моїх дівчат.
RUTH|2|9|Доглядай цього поля, де будуть жати, і ти підеш за ними. Ось я наказав слугам не займати тебе. А як спрагнеш, то підеш до начинь, та й нап'єшся з того, що поначерпують слуги!
RUTH|2|10|І впала вона на обличчя своє, та й вклонилася до землі, і сказала йому: Чому знайшла я милість в очах твоїх, що ти прихилився до мене, хоч я чужа?
RUTH|2|11|І відповів Боаз і сказав їй: Докладно розповіджено мені все, що зробила ти з своєю свекрухою по смерті твого чоловіка, і ти кинула батька свого й матір свою та край свого народження, і пішла до народу, якого не знала вчора-позавчора.
RUTH|2|12|Нехай Господь заплатить за чин твій, і нехай буде нагорода твоя повна від Господа, Бога Ізраїлевого, що ти прийшла сховатися під крильми Його!
RUTH|2|13|А вона сказала: Нехай я знайду милість в очах твоїх, пане мій, бо ти потішив мене, і говорив до серця своєї невільниці. А я не є навіть як одна з твоїх невільниць!
RUTH|2|14|І сказав їй Боаз у час їди: Підійди сюди, та з'їж хліба й замочи у квасі шматок свій. І сіла вона збоку женців, а він подав їй праженого зерна. І їла вона й наситилася, і ще й позоставила.
RUTH|2|15|І встала вона збирати. А Боаз наказав слугам своїм, говорячи: І між снопами нехай збирає, і не кривдьте її.
RUTH|2|16|І також конче киньте їй зо снопів, і позоставте, і буде вона збирати, а ви не лайте її.
RUTH|2|17|І збирала вона на полі аж до вечора, і вимолотила те, що назбирала, і було близько ефи ячменю.
RUTH|2|18|І понесла вона, і ввійшла до міста, і її свекруха побачила, що вона назбирала. А вона вийняла, і дала їй, що позоставила по своїй їжі.
RUTH|2|19|І сказала їй свекруха її: Де ти збирала сьогодні, і де ти робила? Нехай буде благословенний, хто прийняв тебе! І вона розповіла своїй свекрусі, у кого працювала, та й сказала: Ім'я того чоловіка, що я сьогодні робила в нього, Боаз.
RUTH|2|20|І сказала Ноомі до невістки своєї: Благословенний він у Господа, що не позбавив милости своєї ані живих, ані померлих. І сказала їй Ноомі: Близький нам той чоловік, він із наших родичів.
RUTH|2|21|І сказала моавітянка Рут: Він також сказав мені: Пристань до моїх слуг, аж поки не скінчать моїх жнив.
RUTH|2|22|І сказала Ноомі до своєї невістки Рут: Добре, дочко моя, що ти вийдеш з його служницями, щоб не чіпали тебе на іншому полі.
RUTH|2|23|І вона пристала до Боазових служниць, щоб збирати аж до закінчення жнив ячменю та жнив пшениці. І вона жила з своєю свекрухою.
RUTH|3|1|І сказала їй свекруха її Ноомі: Дочко моя, ось я пошукаю для тебе місця спочинку, що буде добре тобі.
RUTH|3|2|А тепер ось Боаз, наш родич, що була ти з його служницями, ось він цієї ночі буде віяти ячмінь на току.
RUTH|3|3|А ти вмийся, і намастися, і надягни на себе кращу одежу свою, та й зійди на тік. Але не показуйся на очі тому чоловікові, аж поки він не скінчить їсти та пити.
RUTH|3|4|І станеться, коли він ляже, то ти зауваж те місце, де він лежить. І ти прийдеш, і відкриєш приніжжя його та й ляжеш, а він скаже тобі, що маєш робити.
RUTH|3|5|А та відказала до неї: Усе, що ти кажеш мені, я зроблю.
RUTH|3|6|І зійшла вона на тік, і зробила все, як наказала їй свекруха її.
RUTH|3|7|А Боаз з'їв та випив, та й стало весело йому на серці, і прийшов він покластися біля копиці. А вона тихо прийшла, і відкрила його приніжжя та й лягла.
RUTH|3|8|І сталося опівночі, і затремтів той чоловік, та й звівся, аж ось жінка лежить у приніжжі його!
RUTH|3|9|І він сказав: Хто ти? А вона відказала: Я невільниця твоя Рут. Простягни ж крило над своєю невільницею, бо ти мій родич.
RUTH|3|10|А він сказав: Благословенна ти в Господа, дочко моя! Твоя остання ласка до мене ліпша від першої, що не пішла ти за юнаками, чи вони бідні, чи вони багаті.
RUTH|3|11|А тепер, дочко моя, не бійся! Усе, що скажеш, я зроблю тобі, бо все місто народу мого знає, що ти жінка чеснотна!
RUTH|3|12|А тепер справді, що я родич, та є родич ще, ближчий від мене.
RUTH|3|13|Ночуй цю ніч, а ранком, якщо він викупить тебе добре, нехай викупить. А якщо він не схоче викупити тебе, то викуплю тебе я, як живий Господь! Лежи тут аж до ранку.
RUTH|3|14|І лежала вона у приніжжі його аж до ранку, і встала, перше ніж можна розпізнати один одного. А він сказав: Нехай не пізнають, що жінка приходила на тік.
RUTH|3|15|І він сказав: Дай хустку, що на тобі, і подерж її. І держала вона її, а він відміряв шість мір ячменю, і поклав на неї, та й пішов до міста.
RUTH|3|16|А вона прийшла до своєї свекрухи. А та сказала: Як справа, дочко моя? А вона розповіла їй усе, що зробив їй той чоловік.
RUTH|3|17|І сказала: Ці шість мір ячменю він дав мені, бо сказав: Не приходь порожньо до своєї свекрухи.
RUTH|3|18|А та сказала: Почекай, моя дочко, аж поки довідаєшся, як випаде справа, бо той чоловік не заспокоїться, доки не викінчить цієї справи сьогодні.
RUTH|4|1|А Боаз прийшов до брами, та й сів там. Аж ось проходить родич, про якого говорив був Боаз. І він сказав йому: Зайди сюди, послухай, і сядь отут! І той зайшов і сів.
RUTH|4|2|А Боаз узяв десять мужа зо старших того міста та й сказав: Сідайте тут! І вони посідали.
RUTH|4|3|І сказав він до родича: Ділянку поля, що нашого брата Елімелеха, продала Ноомі, яка вернулася з моавського поля.
RUTH|4|4|А я постановив: Подам тобі до ушей твоїх, говорячи: Купи при тих, що сидять тут, та при старших мого народу. Якщо викупиш викупи, а якщо не викупиш скажи мені, і нехай я знаю, бо окрім тебе нема кому викупити, а я за тобою. А той сказав: Я викуплю.
RUTH|4|5|І сказав Боаз: Того дня, коли набудеш поле з руки Ноомі, то набудеш також моавитянку Рут, жінку померлого, щоб поставити ім'я померлому на наділі його.
RUTH|4|6|А родич сказав: Не можу я викупити собі, щоб не понищити свого наділу. Викупи собі мого викупа, бо я не можу викупити.
RUTH|4|7|А оце було колись серед Ізраїля на викуп, і на заміну, і на ствердження кожної справи: чоловік здіймав сандалю свою, і давав своєму ближньому, і це було свідоцтвом серед Ізраїля.
RUTH|4|8|І сказав родич до Боаза: Купи собі! І зняв свою сандалю.
RUTH|4|9|І сказав Боаз до старших та до всього народу: Ви свідки сьогодні, що я набув усе, що Елімелехове, і все, що Кілйонове та Махлонове з руки Ноомі.
RUTH|4|10|А також моавітянку Рут, Махлонову жінку, набув я собі за жінку, щоб поставити ім'я померлому на спадкові його, і не буде знищене ім'я померлого між братами його та з брами його місця. Ви сьогодні свідки на це!
RUTH|4|11|І сказав увесь народ, що були в брамі, та старші, свідки: Нехай дасть Господь цю жінку, що входить до дому твого, як Рахиль та як Лію, що вони обидві збудували Ізраїлів дім. І розбагатій в Ефраті, і здобуть собі славне ім'я в Віфлеємі.
RUTH|4|12|А з насіння, що Господь дасть тобі від цієї молодої жінки, нехай стане дім твій, як дім Переца, що Тамар породила була Юді.
RUTH|4|13|І взяв Боаз Рут, і вона стала йому за жінку. І він увійшов до неї, а Господь дав їй вагітність, і вона породила сина.
RUTH|4|14|І сказали жінки до Ноомі: Благословенний Господь, що не позбавив тебе сьогодні родича! І буде славним ім'я його серед Ізраїля.
RUTH|4|15|І він буде тобі потішителем душі та на виживлення твоєї сивини, бо породила його твоя невістка, що любить тебе, що ліпша тобі за сімох синів.
RUTH|4|16|І взяла Ноомі ту дитину, і поклала її на коліна свої, і була їй за няньку.
RUTH|4|17|А сусідки назвали ім'я йому, говорячи: Народився син для Ноомі! І назвали ім'я йому: Овед. А він батько Єссея, Давидового батька.
RUTH|4|18|А оце Перецові нащадки: Перец породив Гецрона,
RUTH|4|19|а Гецрон породив Рама, а Рам породив Аммінадава,
RUTH|4|20|а Аммінадав породив Нахшона, а Нахшон породив Салмона;
RUTH|4|21|а Салмон породив Боаза, а Боаз породив Оведа;
RUTH|4|22|а Овед породив Єссея, а Єссей породив Давида.
