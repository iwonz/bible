HOS|1|1|Слово Господне, которое было к Осии, сыну Беериину, во дни Озии, Иоафама, Ахаза, Езекии, царей Иудейских, и во дни Иеровоама, сына Иоасова, царя Израильского.
HOS|1|2|Начало слова Господня к Осии. И сказал Господь Осии: иди, возьми себе жену блудницу и детей блуда; ибо сильно блудодействует земля сия, отступив от Господа.
HOS|1|3|И пошел он и взял Гомерь, дочь Дивлаима; и она зачала и родила ему сына.
HOS|1|4|И Господь сказал ему: нареки ему имя Изреель, потому что еще немного пройдет, и Я взыщу кровь Изрееля с дома Ииуева, и положу конец царству дома Израилева,
HOS|1|5|и будет в тот день, Я сокрушу лук Израилев в долине Изреель.
HOS|1|6|И зачала еще, и родила дочь, и Он сказал ему: нареки ей имя Лорухама; ибо Я уже не буду более миловать дома Израилева, чтобы прощать им.
HOS|1|7|А дом Иудин помилую и спасу их в Господе Боге их, спасу их ни луком, ни мечом, ни войною, ни конями и всадниками.
HOS|1|8|И, откормив грудью Непомилованную, она зачала, и родила сына.
HOS|1|9|И сказал Он: нареки ему имя Лоамми, потому что вы не Мой народ, и Я не буду вашим [Богом].
HOS|1|10|Но будет число сынов Израилевых как песок морской, которого нельзя ни измерить, ни исчислить; и там, где говорили им: "вы не Мой народ", будут говорить им: "вы сыны Бога живаго".
HOS|1|11|И соберутся сыны Иудины и сыны Израилевы вместе, и поставят себе одну главу, и выйдут из земли [переселения]; ибо велик день Изрееля!
HOS|2|1|Говорите братьям вашим: "Мой народ", и сестрам вашим: "Помилованная".
HOS|2|2|Судитесь с вашею матерью, судитесь; ибо она не жена Моя, и Я не муж ее; пусть она удалит блуд от лица своего и прелюбодеяние от грудей своих,
HOS|2|3|дабы Я не разоблачил ее донага и не выставил ее, как в день рождения ее, не сделал ее пустынею, не обратил ее в землю сухую и не уморил ее жаждою.
HOS|2|4|И детей ее не помилую, потому что они дети блуда.
HOS|2|5|Ибо блудодействовала мать их и осрамила себя зачавшая их; ибо говорила: "пойду за любовниками моими, которые дают мне хлеб и воду, шерсть и лен, елей и напитки".
HOS|2|6|За то вот, Я загорожу путь ее тернами и обнесу ее оградою, и она не найдет стезей своих,
HOS|2|7|и погонится за любовниками своими, но не догонит их, и будет искать их, но не найдет, и скажет: "пойду я, и возвращусь к первому мужу моему; ибо тогда лучше было мне, нежели теперь".
HOS|2|8|А не знала она, что Я, Я давал ей хлеб и вино и елей и умножил у нее серебро и золото, из которого сделали [истукана] Ваала.
HOS|2|9|За то Я возьму назад хлеб Мой в его время и вино Мое в его пору и отниму шерсть и лен Мой, чем покрывается нагота ее.
HOS|2|10|И ныне открою срамоту ее пред глазами любовников ее, и никто не исторгнет ее из руки Моей.
HOS|2|11|И прекращу у нее всякое веселье, праздники ее и новомесячия ее, и субботы ее, и все торжества ее.
HOS|2|12|И опустошу виноградные лозы ее и смоковницы ее, о которых она говорит: "это у меня подарки, которые надарили мне любовники мои"; и Я превращу их в лес, и полевые звери поедят их.
HOS|2|13|И накажу ее за дни служения Ваалам, когда она кадила им и, украсив себя серьгами и ожерельями, ходила за любовниками своими, а Меня забывала, говорит Господь.
HOS|2|14|Посему вот, и Я увлеку ее, приведу ее в пустыню, и буду говорить к сердцу ее.
HOS|2|15|И дам ей оттуда виноградники ее и долину Ахор, в преддверие надежды; и она будет петь там, как во дни юности своей и как в день выхода своего из земли Египетской.
HOS|2|16|И будет в тот день, говорит Господь, ты будешь звать Меня: "муж мой", и не будешь более звать Меня: "Ваали".
HOS|2|17|И удалю имена Ваалов от уст ее, и не будут более вспоминаемы имена их.
HOS|2|18|И заключу в то время для них союз с полевыми зверями и с птицами небесными, и с пресмыкающимися по земле; и лук, и меч, и войну истреблю от земли той, и дам им жить в безопасности.
HOS|2|19|И обручу тебя Мне навек, и обручу тебя Мне в правде и суде, в благости и милосердии.
HOS|2|20|И обручу тебя Мне в верности, и ты познаешь Господа.
HOS|2|21|И будет в тот день, Я услышу, говорит Господь, услышу небо, и оно услышит землю,
HOS|2|22|и земля услышит хлеб и вино и елей; а сии услышат Изреель.
HOS|2|23|И посею ее для Себя на земле, и помилую Непомилованную, и скажу не Моему народу: "ты Мой народ", а он скажет: "Ты мой Бог!"
HOS|3|1|И сказал мне Господь: иди еще и полюби женщину, любимую мужем, но прелюбодействующую, подобно тому, как любит Господь сынов Израилевых, а они обращаются к другим богам и любят виноградные лепешки их.
HOS|3|2|И приобрел я ее себе за пятнадцать сребренников и за хомер ячменя и полхомера ячменя
HOS|3|3|и сказал ей: много дней оставайся у меня; не блуди, и не будь с другим; так же и я буду для тебя.
HOS|3|4|Ибо долгое время сыны Израилевы будут оставаться без царя и без князя и без жертвы, без жертвенника, без ефода и терафима.
HOS|3|5|После того обратятся сыны Израилевы и взыщут Господа Бога своего и Давида, царя своего, и будут благоговеть пред Господом и благостью Его в последние дни.
HOS|4|1|Слушайте слово Господне, сыны Израилевы; ибо суд у Господа с жителями сей земли, потому что нет ни истины, ни милосердия, ни Богопознания на земле.
HOS|4|2|Клятва и обман, убийство и воровство и прелюбодейство крайне распространились, и кровопролитие следует за кровопролитием.
HOS|4|3|За то восплачет земля сия, и изнемогут все, живущие на ней, со зверями полевыми и птицами небесными, даже и рыбы морские погибнут.
HOS|4|4|Но никто не спорь, никто не обличай другого; и твой народ – как спорящие со священником.
HOS|4|5|И ты падешь днем, и пророк падет с тобою ночью, и истреблю матерь твою.
HOS|4|6|Истреблен будет народ Мой за недостаток ведения: так как ты отверг ведение, то и Я отвергну тебя от священнодействия предо Мною; и как ты забыл закон Бога твоего то и Я забуду детей твоих.
HOS|4|7|Чем больше они умножаются, тем больше грешат против Меня; славу их обращу в бесславие.
HOS|4|8|Грехами народа Моего кормятся они, и к беззаконию его стремится душа их.
HOS|4|9|И что будет с народом, то и со священником; и накажу его по путям его, и воздам ему по делам его.
HOS|4|10|Будут есть, и не насытятся; будут блудить, и не размножатся; ибо оставили служение Господу.
HOS|4|11|Блуд, вино и напитки завладели сердцем их.
HOS|4|12|Народ Мой вопрошает свое дерево и жезл его дает ему ответ; ибо дух блуда ввел их в заблуждение, и, блудодействуя, они отступили от Бога своего.
HOS|4|13|На вершинах гор они приносят жертвы и на холмах совершают каждение под дубом и тополем и теревинфом, потому что хороша от них тень; поэтому любодействуют дочери ваши и прелюбодействуют невестки ваши.
HOS|4|14|Я оставлю наказывать дочерей ваших, когда они блудодействуют, и невесток ваших, когда они прелюбодействуют, потому что вы сами на стороне блудниц и с любодейцами приносите жертвы, а невежественный народ гибнет.
HOS|4|15|Если ты, Израиль, блудодействуешь, то пусть не грешил бы Иуда; и не ходите в Галгал, и не восходите в Беф–Авен, и не клянитесь: "жив Господь!"
HOS|4|16|Ибо как упрямая телица, упорен стал Израиль; посему будет ли теперь Господь пасти их, как агнцев на пространном пастбище?
HOS|4|17|Привязался к идолам Ефрем; оставь его!
HOS|4|18|Отвратительно пьянство их, совершенно предались блудодеянию; князья их любят постыдное.
HOS|4|19|Охватит их ветер своими крыльями, и устыдятся они жертв своих.
HOS|5|1|Слушайте это, священники, и внимайте, дом Израилев, и приклоните ухо, дом царя; ибо вам будет суд, потому что вы были западнею в Массифе и сетью, раскинутою на Фаворе.
HOS|5|2|Глубоко погрязли они в распутстве; но Я накажу всех их.
HOS|5|3|Ефрема Я знаю, и Израиль не сокрыт от Меня; ибо ты блудодействуешь, Ефрем, и Израиль осквернился.
HOS|5|4|Дела их не допускают их обратиться к Богу своему, ибо дух блуда внутри них, и Господа они не познали.
HOS|5|5|И гордость Израиля унижена в глазах их; и Израиль и Ефрем падут от нечестия своего; падет и Иуда с ними.
HOS|5|6|С овцами своими и волами своими пойдут искать Господа и не найдут Его: Он удалился от них.
HOS|5|7|Господу они изменили, потому что родили чужих детей; ныне новый месяц поест их с их имуществом.
HOS|5|8|Вострубите рогом в Гиве, трубою в Раме; возглашайте в Беф–Авене: "за тобою, Вениамин!"
HOS|5|9|Ефрем сделается пустынею в день наказания; между коленами Израилевыми Я возвестил это.
HOS|5|10|Вожди Иудины стали подобны передвигающим межи: изолью на них гнев Мой, как воду.
HOS|5|11|Угнетен Ефрем, поражен судом; ибо захотел ходить вслед суетных.
HOS|5|12|И буду как моль для Ефрема и как червь для дома Иудина.
HOS|5|13|И увидел Ефрем болезнь свою, и Иуда – свою рану, и пошел Ефрем к Ассуру, и послал к царю Иареву; но он не может исцелить вас, и не излечит вас от раны.
HOS|5|14|Ибо Я как лев для Ефрема и как скимен для дома Иудина; Я, Я растерзаю, и уйду; унесу, и никто не спасет.
HOS|5|15|Пойду, возвращусь в Мое место, доколе они не признают себя виновными и не взыщут лица Моего.
HOS|6|1|В скорби своей они с раннего утра будут искать Меня и говорить: "пойдем и возвратимся к Господу! ибо Он уязвил – и Он исцелит нас, поразил – и перевяжет наши раны;
HOS|6|2|оживит нас через два дня, в третий день восставит нас, и мы будем жить пред лицем Его.
HOS|6|3|Итак познаем, будем стремиться познать Господа; как утренняя заря – явление Его, и Он придет к нам, как дождь, как поздний дождь оросит землю".
HOS|6|4|Что сделаю тебе, Ефрем? что сделаю тебе, Иуда? благочестие ваше, как утренний туман и как роса, скоро исчезающая.
HOS|6|5|Посему Я поражал через пророков и бил их словами уст Моих, и суд Мой, как восходящий свет.
HOS|6|6|Ибо Я милости хочу, а не жертвы, и Боговедения более, нежели всесожжений.
HOS|6|7|Они же, подобно Адаму, нарушили завет и там изменили Мне.
HOS|6|8|Галаад – город нечестивцев, запятнанный кровью.
HOS|6|9|Как разбойники подстерегают человека, так сборище священников убивают на пути в Сихем и совершают мерзости.
HOS|6|10|В доме Израиля Я вижу ужасное; там блудодеяние у Ефрема, осквернился Израиль.
HOS|6|11|И тебе, Иуда, назначена жатва, когда Я возвращу плен народа Моего.
HOS|7|1|Когда Я врачевал Израиля, открылась неправда Ефрема и злодейство Самарии: ибо они поступают лживо; и входит вор, и разбойник грабит по улицам.
HOS|7|2|Не помышляют они в сердце своем, что Я помню все злодеяния их; теперь окружают их дела их; они пред лицем Моим.
HOS|7|3|Злодейством своим они увеселяют царя и обманами своими – князей.
HOS|7|4|Все они пылают прелюбодейством, как печь, растопленная пекарем, который перестает поджигать ее, когда замесит тесто и оно вскиснет.
HOS|7|5|"День нашего царя!" [говорят] князья, разгоряченные до болезни вином, а он протягивает руку свою к кощунам.
HOS|7|6|Ибо они коварством своим делают сердце свое подобным печи: пекарь их спит всю ночь, а утром она горит, как пылающий огонь.
HOS|7|7|Все они распалены, как печь, и пожирают судей своих; все цари их падают, и никто из них не взывает ко Мне.
HOS|7|8|Ефрем смешался с народами, Ефрем стал, как неповороченный хлеб.
HOS|7|9|Чужие пожирали силу его и он не замечал; седина покрыла его, а он не знает.
HOS|7|10|И гордость Израиля унижена в глазах их и при всем том они не обратились к Господу Богу своему и не взыскали Его.
HOS|7|11|И стал Ефрем, как глупый голубь, без сердца: зовут Египтян, идут в Ассирию.
HOS|7|12|Когда они пойдут, Я закину на них сеть Мою; как птиц небесных низвергну их; накажу их, как слышало собрание их.
HOS|7|13|Горе им, что они удалились от Меня; гибель им, что они отпали от Меня! Я спасал их, а они ложь говорили на Меня.
HOS|7|14|И не взывали ко Мне сердцем своим, когда вопили на ложах своих; собираются из–за хлеба и вина, а от Меня удаляются.
HOS|7|15|Я вразумлял [их] и укреплял мышцы их, а они умышляли злое против Меня.
HOS|7|16|Они обращались, но не к Всевышнему, стали – как неверный лук; падут от меча князья их за дерзость языка своего; это будет посмеянием над ними в земле Египетской.
HOS|8|1|Трубу к устам твоим! Как орел [налетит] на дом Господень за то, что они нарушили завет Мой и преступили закон Мой!
HOS|8|2|Ко Мне будут взывать: "Боже мой! мы познали Тебя, мы – Израиль".
HOS|8|3|Отверг Израиль доброе; враг будет преследовать его.
HOS|8|4|Поставляли царей сами, без Меня; ставили князей, но без Моего ведома; из серебра своего и золота своего сделали для себя идолов: оттуда гибель.
HOS|8|5|Оставил тебя телец твой, Самария! воспылал гнев Мой на них; доколе не могут они очиститься?
HOS|8|6|Ибо и он – дело Израиля: художник сделал его, и потому он не бог; в куски обратится телец Самарийский!
HOS|8|7|Так как они сеяли ветер, то и пожнут бурю: хлеба на корню не будет у него; зерно не даст муки; а если и даст, то чужие проглотят ее.
HOS|8|8|Поглощен Израиль; теперь они будут среди народов как негодный сосуд.
HOS|8|9|Они пошли к Ассуру, как дикий осел, одиноко бродящий; Ефрем приобретал подарками расположение к себе.
HOS|8|10|Хотя они и посылали дары к народам, но скоро Я соберу их, и они начнут страдать от бремени царя князей;
HOS|8|11|ибо много жертвенников настроил Ефрем для греха, – ко греху послужили ему эти жертвенники.
HOS|8|12|Написал Я ему важные законы Мои, но они сочтены им как бы чужие.
HOS|8|13|В жертвоприношениях Мне они приносят мясо и едят его; Господу неугодны они; ныне Он вспомнит нечестие их и накажет их за грехи их: они возвратятся в Египет.
HOS|8|14|Забыл Израиль Создателя своего и устроил капища, и Иуда настроил много укрепленных городов; но Я пошлю огонь на города его, и пожрет чертоги его.
HOS|9|1|Не радуйся, Израиль, до восторга, как [другие] народы, ибо ты блудодействуешь, удалившись от Бога твоего: любишь блудодейные дары на всех гумнах.
HOS|9|2|Гумно и точило не будут питать их, и [надежда] на виноградный сок обманет их.
HOS|9|3|Не будут они жить на земле Господней: Ефрем возвратится в Египет, и в Ассирии будут есть нечистое.
HOS|9|4|Не будут возливать Господу вина, и неугодны Ему будут жертвы их; они будут для них, как хлеб похоронный: все, которые будут есть его, осквернятся, ибо хлеб их – для души их, а в дом Господень он не войдет.
HOS|9|5|Что будете делать в день торжества и в день праздника Господня?
HOS|9|6|Ибо вот, они уйдут по причине опустошения; Египет соберет их, Мемфис похоронит их; драгоценностями их из серебра завладеет крапива, колючий терн будет в шатрах их.
HOS|9|7|Пришли дни посещения, пришли дни воздаяния; да узнает Израиль, что глуп прорицатель, безумен выдающий себя за вдохновенного, по причине множества беззаконий твоих и великой враждебности.
HOS|9|8|Ефрем – страж подле Бога моего; пророк – сеть птицелова на всех путях его; соблазн в доме Бога его.
HOS|9|9|Глубоко упали они, развратились, как во дни Гивы; Он вспомнит нечестие их, накажет их за грехи их.
HOS|9|10|Как виноград в пустыне, Я нашел Израиля; как первую ягоду на смоковнице, в первое время ее, увидел Я отцов ваших, – но они пошли к Ваал–Фегору и предались постыдному, и сами стали мерзкими, как те, которых возлюбили.
HOS|9|11|У Ефремлян, как птица улетит слава: ни рождения, ни беременности, ни зачатия [не будет].
HOS|9|12|А хотя бы они и воспитали детей своих, отниму их; ибо горе им, когда удалюсь от них!
HOS|9|13|Ефрем, как Я видел его до Тира, насажден на прекрасной местности; однако Ефрем выведет детей своих к убийце.
HOS|9|14|Дай им, Господи: что Ты дашь им? дай им утробу нерождающую и сухие сосцы.
HOS|9|15|Все зло их в Галгале: там Я возненавидел их за злые дела их; изгоню их из дома Моего, не буду больше любить их; все князья их – отступники.
HOS|9|16|Поражен Ефрем; иссох корень их, – не будут приносить они плода, а если и будут рождать, Я умерщвлю вожделенный плод утробы их.
HOS|9|17|Отвергнет их Бог мой, потому что они не послушались Его, и будут скитальцами между народами.
HOS|10|1|Израиль – ветвистый виноград, умножает для себя плод: чем более у него плодов, тем более умножает жертвенники; чем лучше земля у него, тем более украшают они кумиры.
HOS|10|2|Разделилось сердце их, за то они и будут наказаны: Он разрушит жертвенники их, сокрушит кумиры их.
HOS|10|3|Теперь они говорят: "нет у нас царя, ибо мы не убоялись Господа; а царь, – что он нам сделает?"
HOS|10|4|Говорят слова [пустые], клянутся ложно, заключают союзы; за то явится суд над ними, как ядовитая трава на бороздах поля.
HOS|10|5|За тельца Беф–Авена вострепещут жители Самарии; восплачет о нем народ его, и жрецы его, радовавшиеся о нем, будут плакать о славе его, потому что она отойдет от него.
HOS|10|6|И сам он отнесен будет в Ассирию, в дар царю Иареву; постыжен будет Ефрем, и посрамится Израиль от замысла своего.
HOS|10|7|Исчезнет в Самарии царь ее, как пена на поверхности воды.
HOS|10|8|И истреблены будут высоты Авена, грех Израиля; терние и волчцы вырастут на жертвенниках их, и скажут они горам: "покройте нас", и холмам: "падите на нас".
HOS|10|9|Больше, нежели во дни Гивы, грешил ты, Израиль; там они устояли; война в Гаваоне против сынов нечестия не постигла их.
HOS|10|10|По желанию Моему накажу их, и соберутся против них народы, и они будут связаны за двойное преступление их.
HOS|10|11|Ефрем – обученная телица, привычная к молотьбе, и Я Сам возложу ярмо на тучную шею его; на Ефреме будут верхом ездить, Иуда будет пахать, Иаков будет боронить.
HOS|10|12|Сейте себе в правду, и пожнете милость; распахивайте у себя новину, ибо время взыскать Господа, чтобы Он, когда придет, дождем пролил на вас правду.
HOS|10|13|Вы возделывали нечестие, пожинаете беззаконие, едите плод лжи, потому что ты надеялся на путь твой, на множество ратников твоих.
HOS|10|14|И произойдет смятение в народе твоем, и все твердыни твои будут разрушены, как Салман разрушил Бет–Арбел в день брани: мать была убита с детьми.
HOS|10|15|Вот что причинит вам Вефиль за крайнее нечестие ваше.
HOS|11|1|На заре погибнет царь Израилев! Когда Израиль был юн, Я любил его и из Египта вызвал сына Моего.
HOS|11|2|Звали их, а они уходили прочь от лица их: приносили жертву Ваалам и кадили истуканам.
HOS|11|3|Я Сам приучал Ефрема ходить, носил его на руках Своих, а они не сознавали, что Я врачевал их.
HOS|11|4|Узами человеческими влек Я их, узами любви, и был для них как бы поднимающий ярмо с челюстей их, и ласково подкладывал пищу им.
HOS|11|5|Не возвратится он в Египет, но Ассур – он будет царем его, потому что они не захотели обратиться [ко Мне].
HOS|11|6|И падет меч на города его, и истребит затворы его, и пожрет их за умыслы их.
HOS|11|7|Народ Мой закоснел в отпадении от Меня, и хотя призывают его к горнему, он не возвышается единодушно.
HOS|11|8|Как поступлю с тобою, Ефрем? как предам тебя, Израиль? Поступлю ли с тобою, как с Адамою, сделаю ли тебе, что Севоиму? Повернулось во Мне сердце Мое, возгорелась вся жалость Моя!
HOS|11|9|Не сделаю по ярости гнева Моего, не истреблю Ефрема, ибо Я Бог, а не человек; среди тебя Святый; Я не войду в город.
HOS|11|10|Вслед Господа пойдут они; как лев, Он даст глас Свой, даст глас Свой, и встрепенутся к Нему сыны с запада,
HOS|11|11|встрепенутся из Египта, как птицы, и из земли Ассирийской, как голуби, и вселю их в домы их, говорит Господь.
HOS|11|12|Окружил Меня Ефрем ложью и дом Израилев лукавством; Иуда держался еще Бога и верен был со святыми.
HOS|12|1|Ефрем пасет ветер и гоняется за восточным ветром, каждый день умножает ложь и разорение; заключают они союз с Ассуром, и в Египет отвозится елей.
HOS|12|2|Но и с Иудою у Господа суд и Он посетит Иакова по путям его, воздаст ему по делам его.
HOS|12|3|Еще во чреве матери запинал он брата своего, а возмужав боролся с Богом.
HOS|12|4|Он боролся с Ангелом – и превозмог; плакал и умолял Его; в Вефиле Он нашел нас и там говорил с нами.
HOS|12|5|А Господь есть Бог Саваоф; Сущий (Иегова) – имя Его.
HOS|12|6|Обратись и ты к Богу твоему; наблюдай милость и суд и уповай на Бога твоего всегда.
HOS|12|7|Хананеянин с неверными весами в руке любит обижать;
HOS|12|8|и Ефрем говорит: "однако я разбогател; накопил себе имущества, хотя во всех моих трудах не найдут ничего незаконного, что было бы грехом".
HOS|12|9|А Я, Господь Бог твой от самой земли Египетской, опять поселю тебя в кущах, как во дни праздника.
HOS|12|10|Я говорил к пророкам, и умножал видения, и чрез пророков употреблял притчи.
HOS|12|11|Если Галаад сделался Авеном, то они стали суетны, в Галгалах заколали в жертву тельцов, и жертвенники их стояли как груды камней на межах поля.
HOS|12|12|Убежал Иаков на поля Сирийские, и служил Израиль за жену, и за жену стерег [овец].
HOS|12|13|Чрез пророка вывел Господь Израиля из Египта, и чрез пророка Он охранял его.
HOS|12|14|Сильно раздражил Ефрем [Господа] и за то кровь его оставит на нем, и поношение его обратит Господь на него.
HOS|13|1|Когда Ефрем говорил, все трепетали. Он был высок в Израиле; но сделался виновным через Ваала, и погиб.
HOS|13|2|И ныне прибавили они ко греху: сделали для себя литых истуканов из серебра своего, по понятию своему, – полная работа художников, – и говорят они приносящим жертву людям: "целуйте тельцов!"
HOS|13|3|За то они будут как утренний туман, как роса, скоро исчезающая, как мякина, свеваемая с гумна, и как дым из трубы.
HOS|13|4|Но Я – Господь Бог твой от земли Египетской, – и ты не должен знать другого бога, кроме Меня, и нет спасителя, кроме Меня.
HOS|13|5|Я признал тебя в пустыне, в земле жаждущей.
HOS|13|6|Имея пажити, они были сыты; а когда насыщались, то превозносилось сердце их, и потому они забывали Меня.
HOS|13|7|И Я буду для них как лев, как скимен буду подстерегать при дороге.
HOS|13|8|Буду нападать на них, как лишенная детей медведица, и раздирать вместилище сердца их, и поедать их там, как львица; полевые звери будут терзать их.
HOS|13|9|Погубил ты себя, Израиль, ибо только во Мне опора твоя.
HOS|13|10|Где царь твой теперь? Пусть он спасет тебя во всех городах твоих! Где судьи твои, о которых говорил ты: "дай нам царя и начальников"?
HOS|13|11|И Я дал тебе царя во гневе Моем, и отнял в негодовании Моем.
HOS|13|12|Связано в узел беззаконие Ефрема, сбережен его грех.
HOS|13|13|Муки родильницы постигнут его; он – сын неразумный, иначе не стоял бы долго в положении рождающихся детей.
HOS|13|14|От власти ада Я искуплю их, от смерти избавлю их. Смерть! где твое жало? ад! где твоя победа? Раскаяния в том не будет у Меня.
HOS|13|15|Хотя [Ефрем] плодовит между братьями, но придет восточный ветер, поднимется ветер Господень из пустыни, и иссохнет родник его, и иссякнет источник его; он опустошит сокровищницу всех драгоценных сосудов.
HOS|14|1|Опустошена будет Самария, потому что восстала против Бога своего; от меча падут они; младенцы их будут разбиты, и беременные их будут рассечены.
HOS|14|2|Обратись, Израиль, к Господу Богу твоему; ибо ты упал от нечестия твоего.
HOS|14|3|Возьмите с собою [молитвенные] слова и обратитесь к Господу; говорите Ему: "отними всякое беззаконие и прими во благо, и мы принесем жертву уст наших.
HOS|14|4|Ассур не будет уже спасать нас; не станем садиться на коня и не будем более говорить изделию рук наших: боги наши; потому что у Тебя милосердие для сирот".
HOS|14|5|Уврачую отпадение их, возлюблю их по благоволению; ибо гнев Мой отвратился от них.
HOS|14|6|Я буду росою для Израиля; он расцветет, как лилия, и пустит корни свои, как Ливан.
HOS|14|7|Расширятся ветви его, и будет красота его, как маслины, и благоухание от него, как от Ливана.
HOS|14|8|Возвратятся сидевшие под тенью его, будут изобиловать хлебом, и расцветут, как виноградная лоза, славны будут, как вино Ливанское.
HOS|14|9|"Что мне еще за дело до идолов?" – скажет Ефрем. – Я услышу его и призрю на него; Я буду как зеленеющий кипарис; от Меня будут тебе плоды.
HOS|14|10|Кто мудр, чтобы разуметь это? кто разумен, чтобы познать это? Ибо правы пути Господни, и праведники ходят по ним, а беззаконные падут на них.
