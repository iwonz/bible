NEH|1|1|哈迦利亚 的儿子 尼希米 的言语如下： 亚达薛西 王二十年基斯流月，我在 书珊 城堡中。
NEH|1|2|那时，我有一个兄弟 哈拿尼 ，同几个人从 犹大 来。我问他们那些被掳归回、剩下残存的 犹太 人和 耶路撒冷 的情况。
NEH|1|3|他们对我说：“那些被掳归回剩下的余民在 犹大 省那里遭大难，受凌辱； 耶路撒冷 的城墙被拆毁，城门被火焚烧。”
NEH|1|4|我听见这话，就坐下哭泣，悲哀几日，在天上的上帝面前禁食祈祷，
NEH|1|5|说：“唉，耶和华－天上大而可畏的上帝，向爱你、守你诫命的人守约施慈爱的上帝啊，
NEH|1|6|愿你睁眼看，侧耳听你仆人今日昼夜在你面前，为你众仆人 以色列 人的祈祷，承认我们 以色列 人向你所犯的罪；我与我父家都犯了罪。
NEH|1|7|我们向你所行的非常败坏，没有遵守你吩咐你仆人 摩西 的诫命、律例、典章。
NEH|1|8|求你记念所吩咐你仆人 摩西 的话，说：‘你们若犯罪，我就把你们分散在万民中；
NEH|1|9|但你们若归向我，谨守遵行我的诫命，你们被赶散的人虽在天涯，我也必从那里将他们召集回来，带到我所选择立为我名居所的地方。’
NEH|1|10|他们是你的仆人和你的百姓，是你用大力和大能的手所救赎的。
NEH|1|11|唉，主啊，求你侧耳听你仆人的祈祷，听喜爱敬畏你名众仆人的祈祷，使你仆人今日亨通，在这人面前蒙恩。” 我是王的酒政。
NEH|2|1|亚达薛西 王二十年尼散月，酒摆在王面前 ，我拿起酒来奉给王。我在王面前从来没有愁容。
NEH|2|2|王对我说：“你既没有病，为什么面带愁容呢？这不是别的，必是你心中愁烦。”于是我非常惧怕。
NEH|2|3|我对王说：“愿王万岁！我祖先坟墓所在的那城荒凉，城门被火焚烧，我岂能面无愁容呢？”
NEH|2|4|王对我说：“你想求什么？”于是我向天上的上帝祈祷。
NEH|2|5|我对王说：“王若以为好，仆人若在王面前蒙宠爱，求王差遣我往 犹大 ，到我祖先坟墓所在的那城去，我好重新建造。”
NEH|2|6|那时王后坐在王的旁边，王对我说：“你要去多久？几时回来？”王看这事为好，就派我去。我给王定了日期。
NEH|2|7|我又对王说：“王若以为好，求王赐我诏书，通知 河西 的省长准我经过，直到 犹大 ；
NEH|2|8|又赐诏书，通知管理王园林的 亚萨 ，叫他给我木材，作为殿的营楼之门、城墙，和我自己要住的房屋的横梁。”王就允准我，因为我上帝施恩的手帮助我。
NEH|2|9|王派了军官和骑兵护送我。我到了 河西 的省长那里，将王的诏书交给他们。
NEH|2|10|和伦 人 参巴拉 和作臣仆的 亚扪 人 多比雅 ，听见有人来为 以色列 人争取利益，就很恼怒。
NEH|2|11|我到了 耶路撒冷 ，在那里停留了三天。
NEH|2|12|夜间我和跟随我的几个人起来；但上帝感动我心要为 耶路撒冷 做的事，我并没有告诉人。只有我自己骑的牲口，没有别的牲口在我那里。
NEH|2|13|当夜，我出了 谷门 ，往 野狗泉 去，到了 粪厂门 ，察看 耶路撒冷 的城墙，城墙被拆毁，城门被火焚烧。
NEH|2|14|我又往前，到了 泉门 ，又到 王池 ，但所骑的牲口没有地方可以过去。
NEH|2|15|于是我夜间沿溪而上，察看城墙，又转身进入 谷门 ，就回来了。
NEH|2|16|我往哪里去，我做什么事，官长都不知道。我也没有告诉 犹大 人、祭司、贵族、官长和其余做工的人。
NEH|2|17|以后，我对他们说：“我们所遭的难， 耶路撒冷 怎样荒凉，城门被火焚烧，你们都看见了。来吧，让我们重建 耶路撒冷 的城墙，免得再受凌辱！”
NEH|2|18|我告诉他们我上帝施恩的手怎样帮助我，以及王向我所说的话。他们就说：“我们起来建造吧！”于是他们使自己的手坚强，做这美好的工作。
NEH|2|19|但 和伦 人 参巴拉 、作臣仆的 亚扪 人 多比雅 和 阿拉伯 人 基善 听见就嗤笑我们，藐视我们，说：“你们所做的这事是什么呢？要背叛王吗？”
NEH|2|20|我回答他们的话，对他们说：“天上的上帝必使我们亨通。我们作他仆人的，要起来建造；你们却在 耶路撒冷 无份、无权、无名号 。”
NEH|3|1|那时， 以利亚实 大祭司和他的弟兄众祭司起来建立 羊门 ，将门分别为圣，安立门扇，直到 哈米亚楼 。他们又将它分别为圣，直到 哈楠业楼 。
NEH|3|2|在他旁边建造的是 耶利哥 人。在他旁边建造的是 音利 的儿子 撒刻 。
NEH|3|3|哈西拿 的子孙建立 鱼门 ，架横梁、安门扇，装闩和锁。
NEH|3|4|在他们旁边修造的是 哈哥斯 的孙子， 乌利亚 的儿子 米利末 。在他们旁边修造的是 米示萨别 的孙子， 比利迦 的儿子 米书兰 。在他们旁边修造的是 巴拿 的儿子 撒督 。
NEH|3|5|在他们旁边修造的是 提哥亚 人；但是他们的贵族不用肩 扛他们主人的工作。
NEH|3|6|巴西亚 的儿子 耶何耶大 与 比所玳 的儿子 米书兰 修造 古门 ，架横梁，安门扇，装闩和锁。
NEH|3|7|在他们旁边修造的是 基遍 人 米拉提 、 米伦 人 雅顿 、 基遍 人，和 河西 总督所管的 米斯巴 人。
NEH|3|8|在他旁边修造的是 哈海雅 的儿子 乌薛 银匠。在他旁边修造的是做香料的 哈拿尼雅 。他们修复 耶路撒冷 ，直到 宽墙 。
NEH|3|9|在他们旁边修造的是管理 耶路撒冷 城区的一半、 户珥 的儿子 利法雅 。
NEH|3|10|在他们旁边的是 哈路抹 的儿子 耶大雅 在自己房屋的对面修造。在他旁边修造的是 哈沙尼 的儿子 哈突 。
NEH|3|11|哈琳 的儿子 玛基雅 和 巴哈．摩押 的儿子 哈述 修造下一段和 炉楼 。
NEH|3|12|在他旁边修造的是管理 耶路撒冷 城区的另一半、 哈罗黑 的儿子 沙龙 和他的女儿们。
NEH|3|13|哈嫩 和 撒挪亚 的居民修造 谷门 ；他们立门，安门扇，装闩和锁，又修造城墙一千肘，直到 粪厂门 。
NEH|3|14|管理 伯．哈基琳 区、 利甲 的儿子 玛基雅 修造 粪厂门 ；他立门，安门扇，装闩和锁。
NEH|3|15|管理 米斯巴 区、 各．荷西 的儿子 沙仑 修造 泉门 ；他立门，盖门顶，安门扇，装闩和锁，又修造靠近王的花园 西罗亚池 的城墙，直到那从 大卫城 下来的台阶。
NEH|3|16|接续他修造的是管理 伯．夙 区的一半、 押卜 的儿子 尼希米 ，直到 大卫 坟地的对面，又到人造池，到达勇士的房屋。
NEH|3|17|接续他修造的是 利未 人 巴尼 的儿子 利宏 。在他旁边的是管理 基伊拉 区一半的 哈沙比雅 为本区修造。
NEH|3|18|接续他修造的是他们弟兄中管理 基伊拉 区的另一半、 希拿达 的儿子 宾内 。
NEH|3|19|在他旁边的是管理 米斯巴 、 耶书亚 的儿子 以谢珥 修造武库的上坡对面、城墙转弯处的那一段。
NEH|3|20|接续他的是 萨拜 的儿子 巴录 竭力修造下一段，从转弯处，直到 以利亚实 大祭司的府门。
NEH|3|21|接续他的是 哈哥斯 的孙子， 乌利亚 的儿子 米利末 修造下一段，从 以利亚实 的府门，直到 以利亚实 府的尽头。
NEH|3|22|接续他修造的是住平原的祭司。
NEH|3|23|接续他的是 便雅悯 与 哈述 在自己房屋的对面修造。接续他的是 亚难尼 的孙子， 玛西雅 的儿子 亚撒利雅 在自己房屋的旁边修造。
NEH|3|24|接续他的是 希拿达 的儿子 宾内 修造下一段，从 亚撒利雅 的房屋直到转弯处，又到城角。
NEH|3|25|乌赛 的儿子 巴拉 修造转弯处的对面和靠近护卫院、王宫上层凸出来的城楼。接续他的是 巴录 的儿子 毗大雅 ，
NEH|3|26|（殿役住在 俄斐勒 ，直到朝东 水门 的对面和凸出来的城楼。）
NEH|3|27|接续他的是 提哥亚 人又修造一段，对着那凸出来的大城楼，直到 俄斐勒 的城墙。
NEH|3|28|从 马门 往上，祭司各在自己房屋的对面修造。
NEH|3|29|接续他的是 音麦 的儿子 撒督 在自己房屋的对面修造。接续他修造的是 东门 的守卫、 示迦尼 的儿子 示玛雅 。
NEH|3|30|接续他的是 示利米雅 的儿子 哈拿尼雅 和 萨拉 的第六个儿子 哈嫩 修造下一段。接续他的是 比利迦 的儿子 米书兰 在自己房屋的对面修造。
NEH|3|31|接续他的是 玛基雅 银匠修造，直到殿役和商人的房屋，对着 集合门 ，直到角楼。
NEH|3|32|银匠与商人在角楼和 羊门 之间修造。
NEH|4|1|参巴拉 听见我们建造城墙就发怒，非常恼恨，并嗤笑 犹太 人。
NEH|4|2|他对他的弟兄和 撒玛利亚 的军兵说：“这些软弱的 犹太 人做什么呢？要为自己重建吗 ？要献祭吗？要一日完工吗？要使土堆里火烧过的石头再有用吗？”
NEH|4|3|亚扪 人 多比雅 在一旁说：“他们所修造的石墙，就是狐狸上去也必崩裂。”
NEH|4|4|我们的上帝啊，求你垂听，因为我们被藐视。求你使他们的毁谤归于他们自己头上，使他们在被掳之地成为掠物。
NEH|4|5|不要遮掩他们的罪孽，不要使他们的罪恶从你面前涂去，因为他们在修造的人前面惹你发怒。
NEH|4|6|这样，我们修造城墙，整个城墙就连接起来，到一半高，因为百姓一心做工。
NEH|4|7|参巴拉 、 多比雅 、 阿拉伯 人、 亚扪 人和 亚实突 人听见 耶路撒冷 城墙正在修造，破裂的地方开始进行修补，就非常愤怒。
NEH|4|8|大家同谋要来攻打 耶路撒冷 ，使城混乱。
NEH|4|9|然而，我们向我们的上帝祷告，又因他们的缘故，就派人站岗，昼夜防备他们。
NEH|4|10|但 犹大 有话说： “扛抬的人力气衰弱， 瓦砾太多， 我们自己不可能 建造城墙。”
NEH|4|11|我们的敌人说：“趁他们不知道，看不见的时候，我们进入他们中间，杀了他们，使工作停止。”
NEH|4|12|那靠近敌人居住的 犹太 人十次从各处来见我们，说：“你们必须回到我们那里。”
NEH|4|13|我叫百姓站在城墙后边低洼的空处，使百姓各按宗族站着，拿刀、拿枪、拿弓。
NEH|4|14|我察看了，就起来对贵族、官长和其余的百姓说：“不要怕他们！当记得主是大而可畏的。你们要为你们的弟兄、儿女、妻子、家园争战。”
NEH|4|15|仇敌听见我们知道了他们的计谋，上帝也破坏他们的计谋，我们就都回到城墙那里，各做各的工。
NEH|4|16|从那日起，我的仆人一半做工，一半拿枪、拿盾牌、拿弓、穿铠甲，官长都站在 犹大 全家的后边。
NEH|4|17|他们建造城墙；扛抬材料的人扛抬的时候，一手做工，一手拿兵器。
NEH|4|18|建造的人都腰间佩刀建造，吹角的人在我旁边。
NEH|4|19|我对贵族、官长和其余的百姓说：“这工程浩大，范围辽阔，我们在城墙上彼此相离很远。
NEH|4|20|你们一听见角声在哪里，就聚集到我们那里去。我们的上帝必为我们争战。”
NEH|4|21|于是，我们做这工程，一半的人拿枪，从天亮直到星宿出现的时候。
NEH|4|22|那时，我又对百姓说：“各人和他的仆人当在 耶路撒冷 过夜，好为我们夜间守卫，白昼做工。”
NEH|4|23|这样，我和弟兄仆人，以及跟从我的卫兵都不脱衣服，各人打水时 也拿着自己的兵器。
NEH|5|1|百姓和他们的妻子大大呼号，埋怨他们的弟兄 犹太 人。
NEH|5|2|有的说：“我们和儿女人口众多，必须得粮食吃，才能活下去。”
NEH|5|3|有的说：“我们典押了田地、葡萄园、房屋，才得粮食充饥。”
NEH|5|4|有的说：“我们借了钱付田地和葡萄园的税给王。
NEH|5|5|现在，我们的身体与我们弟兄的身体是一样的，我们的儿女与他们的儿女没有差别。看哪，我们却要迫使儿女作人的奴婢。我们有些女儿已被抢走了，我们却无能为力，因为我们的田地和葡萄园已经归了别人。”
NEH|5|6|我听见他们的呼号和这些话，就非常愤怒。
NEH|5|7|我心里作了决定，就斥责贵族和官长，对他们说：“你们各人借钱给弟兄，竟然索取利息！”于是我召开大会攻击他们。
NEH|5|8|我对他们说：“我们已尽力赎回我们的弟兄，就是卖到列国的 犹太 人；你们还要卖弟兄，让我们去买回来吗？”他们就静默不语，无话可答。
NEH|5|9|我又说：“你们做的这事不对！你们行事不是应该敬畏我们的上帝，免得列国我们的仇敌毁谤我们吗？
NEH|5|10|我和我的弟兄仆人也要把银钱粮食借给百姓，大家都当免除利息。
NEH|5|11|就在今日，你们要把他们的田地、葡萄园、橄榄园、房屋，以及向他们所取银钱的利息 、粮食、新酒和新油都归还他们。”
NEH|5|12|贵族和官长说：“我们必归还，不再向他们索取，必照你所说的去做。”我就召了祭司来，叫贵族和官长起誓，必照这话去做。
NEH|5|13|我也抖着胸前的衣袋，说：“凡不实行这话的，愿上帝照样抖他离开他的家和他劳碌得来的，直到抖空了。”全会众都说：“阿们！”又赞美耶和华。百姓就照着这话去做。
NEH|5|14|自从我奉派作 犹大 地省长的那日，就是从 亚达薛西 王二十年直到三十二年，共十二年之久，我与我弟兄都没有吃省长的俸禄。
NEH|5|15|在我以前的省长加重百姓的负担，向百姓索取粮食和酒，以及四十舍客勒银子 ，甚至他们的仆人也辖制百姓，但我因敬畏上帝不这样做。
NEH|5|16|我也努力修造城墙。我们并没有购置田地，我所有的仆人也都聚集在那里做工。
NEH|5|17|除了从四围列国来的人以外，有 犹太 人和官长一百五十人与我同席。
NEH|5|18|每日预备一头公牛，六只肥羊，又为我预备飞禽；每十日一次多多预备各样的酒。虽然如此，我并不索取省长的俸禄，因为这百姓负的劳役很重。
NEH|5|19|我的上帝啊，求你记念我为这百姓所做的一切，施恩于我。
NEH|6|1|参巴拉 、 多比雅 、 阿拉伯 人 基善 和我们其余的仇敌听见我已经建造了城墙，没有破裂之处在其中，那时我还没有在城门安门扇；
NEH|6|2|参巴拉 和 基善 就派人来见我，说：“请你来，我们在 阿挪 平原的村庄见面。”其实，他们想要害我。
NEH|6|3|于是我派使者到他们那里，说：“我正在进行大的工程，不能下去。我怎么能离开，下去见你们，而让工程停顿呢？”
NEH|6|4|他们这样派人来见我四次，我都用这话回答他们。
NEH|6|5|参巴拉 第五次同样派仆人来见我，手里拿着未封的信，
NEH|6|6|信上写着：“列国中有风声， 基善 也说，你和 犹太 人谋反，所以你建造城墙。据说，你要作他们的王，
NEH|6|7|并且你派先知在 耶路撒冷 指着你宣讲说，‘在 犹大 有王。’如今这些话必传给王知，现在请你来，我们一起商议。”
NEH|6|8|我就派人到他那里，说：“你所说的这些事，一概没有，是你心里捏造的。”
NEH|6|9|他们全都要使我们惧怕，说：“他们的手必软弱，不能工作，以致不能完工。”现在，求你坚固我的手。
NEH|6|10|我到了 米希大别 的孙子， 第来雅 的儿子 示玛雅 家里；那时，他闭门不出。他说：“我们可以在上帝的殿里，就在殿的中间会面，锁住殿门，因为他们要来杀你，要在夜里来杀你。”
NEH|6|11|我说：“像我这样的人岂会逃跑呢？像我这样的人岂能进入殿里保全生命呢？我不进去！”
NEH|6|12|我看清楚了，看哪，上帝并没有派他，是他自己说预言攻击我，是 多比雅 和 参巴拉 收买了他；
NEH|6|13|收买他的目的是要叫我惧怕，依从他犯罪，留下一个坏名声，好让他们毁谤我。
NEH|6|14|我的上帝啊，求你记得 多比雅 、 参巴拉 、 挪亚底 女先知和其余的先知，因他们行这些事，要叫我惧怕。
NEH|6|15|以禄月二十五日，城墙修完了，共修了五十二天。
NEH|6|16|我们所有的仇敌听见了，四围的列国就惧怕，愁眉不展，因为他们知道这工作得以完成，是出于我们的上帝。
NEH|6|17|而且，在那些日子， 犹大 的贵族屡次寄信给 多比雅 ， 多比雅 也回信给他们。
NEH|6|18|在 犹大 有许多人与 多比雅 结盟，因为他是 亚拉 的儿子 示迦尼 的女婿，并且他的儿子 约哈难 娶了 比利迦 的儿子 米书兰 的女儿。
NEH|6|19|他们也在我面前说 多比雅 的好话，又把我的话传给他。 多比雅 常寄信来，要叫我惧怕。
NEH|7|1|城墙修完，我安了门扇，门口的守卫、歌唱的和 利未 人都已派定。
NEH|7|2|我吩咐我的兄弟 哈拿尼 和城堡的官长 哈拿尼雅 管理 耶路撒冷 ，因为 哈拿尼雅 是一个忠信的人，敬畏上帝过于众人。
NEH|7|3|我对他们说：“等到太阳热的时候才可开 耶路撒冷 的城门；要派 耶路撒冷 的居民，各按班次在自己房屋的前面站岗。他们还在站岗的时候，就要关门上闩。”
NEH|7|4|城又宽又大，城中的百姓却稀少，房屋也还没有建造。
NEH|7|5|我的上帝感动我的心，我就召集贵族、官长和百姓，要登记家谱。我找到第一次上来之人的家谱，发现上面写着：
NEH|7|6|这些是从被掳之地上来的省民， 巴比伦 王 尼布甲尼撒 把他们掳去，他们重返 耶路撒冷 和 犹大 ，各归本城。
NEH|7|7|他们是同 所罗巴伯 、 耶书亚 、 尼希米 、 亚撒利雅 、 拉米 、 拿哈玛尼 、 末底改 、 必珊 、 米斯毗列 、 比革瓦伊 、 尼宏 、 巴拿 一起回来的。 以色列 百姓的人数如下：
NEH|7|8|巴录 的子孙二千一百七十二名；
NEH|7|9|示法提雅 的子孙三百七十二名；
NEH|7|10|亚拉 的子孙六百五十二名；
NEH|7|11|巴哈．摩押 的后裔，就是 耶书亚 和 约押 的子孙二千八百一十八名；
NEH|7|12|以拦 的子孙一千二百五十四名；
NEH|7|13|萨土 的子孙八百四十五名；
NEH|7|14|萨改 的子孙七百六十名；
NEH|7|15|宾内 的子孙六百四十八名；
NEH|7|16|比拜 的子孙六百二十八名；
NEH|7|17|押甲 的子孙二千三百二十二名；
NEH|7|18|亚多尼干 的子孙六百六十七名；
NEH|7|19|比革瓦伊 的子孙二千零六十七名；
NEH|7|20|亚丁 的子孙六百五十五名；
NEH|7|21|亚特 的后裔，就是 希西家 的子孙九十八名；
NEH|7|22|哈顺 的子孙三百二十八名；
NEH|7|23|比赛 的子孙三百二十四名；
NEH|7|24|哈拉 的子孙一百一十二名；
NEH|7|25|基遍 人九十五名；
NEH|7|26|伯利恒 人和 尼陀法 人共一百八十八名；
NEH|7|27|亚拿突 人一百二十八名；
NEH|7|28|伯．亚斯玛弗 人四十二名；
NEH|7|29|基列．耶琳 人、 基非拉 人、 比录 人共七百四十三名；
NEH|7|30|拉玛 人和 迦巴 人共六百二十一名；
NEH|7|31|默玛 人一百二十二名；
NEH|7|32|伯特利 人和 艾 人共一百二十三名；
NEH|7|33|别的 尼波 人五十二名；
NEH|7|34|另一个 以拦 子孙一千二百五十四名；
NEH|7|35|哈琳 的子孙三百二十名；
NEH|7|36|耶利哥 人三百四十五名；
NEH|7|37|罗德 人、 哈第 人、 阿挪 人共七百二十一名；
NEH|7|38|西拿 人三千九百三十名。
NEH|7|39|祭司： 耶书亚 家， 耶大雅 的子孙九百七十三名；
NEH|7|40|音麦 的子孙一千零五十二名；
NEH|7|41|巴施户珥 的子孙一千二百四十七名；
NEH|7|42|哈琳 的子孙一千零一十七名。
NEH|7|43|利未 人： 何达威 的后裔，就是 耶书亚 和 甲篾 的子孙七十四名。
NEH|7|44|歌唱的： 亚萨 的子孙一百四十八名。
NEH|7|45|门口的守卫： 沙龙 的子孙、 亚特 的子孙、 达们 的子孙、 亚谷 的子孙、 哈底大 的子孙、 朔拜 的子孙，共一百三十八名。
NEH|7|46|殿役： 西哈 的子孙、 哈苏巴 的子孙、 答巴俄 的子孙、
NEH|7|47|基绿 的子孙、 西亚 的子孙、 巴顿 的子孙、
NEH|7|48|利巴拿 的子孙、 哈迦巴 的子孙、 萨买 的子孙、
NEH|7|49|哈难 的子孙、 吉德 的子孙、 迦哈 的子孙、
NEH|7|50|利亚雅 的子孙、 利汛 的子孙、 尼哥大 的子孙、
NEH|7|51|迦散 的子孙、 乌撒 的子孙、 巴西亚 的子孙、
NEH|7|52|比赛 的子孙、 米乌宁 的子孙、 尼普心 的子孙、
NEH|7|53|巴卜 的子孙、 哈古巴 的子孙、 哈忽 的子孙、
NEH|7|54|巴洗律 的子孙、 米希大 的子孙、 哈沙 的子孙、
NEH|7|55|巴柯 的子孙、 西西拉 的子孙、 答玛 的子孙、
NEH|7|56|尼细亚 的子孙、 哈提法 的子孙。
NEH|7|57|所罗门 仆人的后裔： 琐太 的子孙、 琐斐列 的子孙、 比路大 的子孙、
NEH|7|58|雅拉 的子孙、 达昆 的子孙、 吉德 的子孙、
NEH|7|59|示法提雅 的子孙、 哈替 的子孙、 玻黑列．哈斯巴音 的子孙、 亚们 的子孙。
NEH|7|60|殿役和 所罗门 仆人的后裔共三百九十二名。
NEH|7|61|从 特．米拉 、 特．哈萨 、 基绿 、 亚顿 、 音麦 上来，不能证明他们的父系家族和后裔是否属 以色列 的如下：
NEH|7|62|第莱雅 的子孙、 多比雅 的子孙、 尼哥大 的子孙，共六百四十二名。
NEH|7|63|祭司中， 哈巴雅 的子孙、 哈哥斯 的子孙、 巴西莱 的子孙， 巴西莱 因为娶了 基列 人 巴西莱 的女儿为妻，所以就以此为名。
NEH|7|64|这些人在族谱之中寻查自己的谱系，却寻不着，因此算为不洁，不得作祭司。
NEH|7|65|省长对他们说，不可吃至圣的物，直到有会用乌陵和土明的祭司兴起来。
NEH|7|66|全会众共有四万二千三百六十名。
NEH|7|67|此外，还有他们的仆婢七千三百三十七名，又有歌唱的男女二百四十五名。
NEH|7|68|他们有七百三十六匹马，二百四十五匹骡子，
NEH|7|69|四百三十五匹骆驼，六千七百二十匹驴。
NEH|7|70|有些族长为工程捐助。省长捐入库房中的有一千达利克 金子，五十个碗，五百三十件祭司的礼服。
NEH|7|71|有些族长捐入工程的库房，有二万达利克金子，二千二百弥那银子。
NEH|7|72|其余百姓所捐的有二万达利克金子，二千弥那银子，六十七件祭司的礼服。
NEH|7|73|于是祭司、 利未 人、门口的守卫、歌唱的、百姓中的一些人、殿役，并 以色列 众人，都住在自己的城里。 到了七月， 以色列 人住在自己的城里。
NEH|8|1|那时，众百姓如同一人聚集在 水门 前的广场，请 以斯拉 文士将耶和华吩咐 以色列 的 摩西 的律法书带来。
NEH|8|2|七月初一， 以斯拉 祭司将律法书带到听了能明白的男女会众面前。
NEH|8|3|他在 水门 前的广场，从清早到中午，在男女和能明白的人面前读这律法书，众百姓都侧耳而听。
NEH|8|4|以斯拉 文士站在为这事特制的木台上。站在他旁边的有 玛他提雅 、 示玛 、 亚奈雅 、 乌利亚 和 希勒家 ；站在他右边的有 玛西雅 ；站在他左边的有 毗大雅 、 米沙利 、 玛基雅 、 哈顺 、 哈拔大拿 、 撒迦利亚 和 米书兰 。
NEH|8|5|以斯拉 站在上面，在众百姓眼前展开这书。他一展开，众百姓都站起来。
NEH|8|6|以斯拉 称颂耶和华至大的上帝，众百姓都举手应声说：“阿们！阿们！”他们低头，俯伏在地，敬拜耶和华。
NEH|8|7|耶书亚 、 巴尼 、 示利比 、 雅悯 、 亚谷 、 沙比太 、 荷第雅 、 玛西雅 、 基利他 、 亚撒利雅 、 约撒拔 、 哈难 、 毗莱雅 和 利未 人使百姓明白律法；百姓都站在自己的地方。
NEH|8|8|他们清清楚楚地念上帝的律法书，讲明意思，使百姓明白所念的。
NEH|8|9|尼希米 省长、 以斯拉 祭司文士，和教导百姓的 利未 人对众百姓说：“今日是耶和华－你们上帝的圣日，不要悲哀，也不要哭泣。”这是因为众百姓听见律法书上的话都哭了。
NEH|8|10|尼希米 对他们说：“你们去吃肥美的，喝甘甜的，有不能预备的就分给他，因为今日是我们主的圣日。你们不要忧愁，因靠耶和华而得的喜乐是你们的力量。”
NEH|8|11|于是 利未 人叫众百姓安静，说：“安静，因今日是圣日，不要忧愁。”
NEH|8|12|众百姓去吃喝，也分给别人，都大大喜乐，因为他们明白所教导他们的话。
NEH|8|13|次日，众百姓的族长、祭司和 利未 人都聚集到 以斯拉 文士那里，要明白律法书上的话。
NEH|8|14|他们发现律法书上写着，耶和华藉 摩西 吩咐 以色列 人要在七月的节期中住在棚里，
NEH|8|15|并要在各城和 耶路撒冷 传扬宣告说：“你们当出去，上山，把橄榄树、野橄榄树、番石榴树、棕树和各样茂密树的枝子取来，照着所写的搭棚。”
NEH|8|16|于是百姓出去，取了树枝来，各人在自己的房顶上，院子里，上帝殿的院内， 水门 的广场，和 以法莲门 的广场搭棚。
NEH|8|17|从被掳之地归回的全会众就搭棚，住在棚里。从 嫩 的儿子 约书亚 的时候直到这日， 以色列 人没有这样行。他们都大大喜乐。
NEH|8|18|从第一天直到末一天， 以斯拉 天天朗读上帝的律法书。他们守节七日，第八日照例有严肃会。
NEH|9|1|这月二十四日， 以色列 人聚集禁食，他们披麻蒙灰。
NEH|9|2|以色列 的后裔与所有的外邦人分别出来，站着承认自己的罪和祖先的罪孽。
NEH|9|3|那日的四分之一，他们站在自己的地方念耶和华－他们上帝的律法书，又在那日的四分之一认罪，敬拜耶和华－他们的上帝。
NEH|9|4|耶书亚 、 巴尼 、 甲篾 、 示巴尼 、 布尼 、 示利比 、 巴尼 、 基拿尼 站在 利未 人的台阶上，大声哀求耶和华－他们的上帝。
NEH|9|5|利未 人 耶书亚 、 甲篾 、 巴尼 、 哈沙尼 、 示利比 、 荷第雅 、 示巴尼 、 毗他希雅 说：“起来，称颂耶和华－你们的上帝，永世无尽：‘你荣耀之名是应当称颂的，超乎一切称颂和赞美。
NEH|9|6|“‘你，惟独你是耶和华！你造了天和天上的天，以及天上的万象，地和地上的万物，海和海中所有的；一切的生命全都是你赏赐的。天军都敬拜你。
NEH|9|7|你是耶和华上帝，曾拣选 亚伯兰 ，领他出 迦勒底 的 吾珥 ，给他改名叫 亚伯拉罕 。
NEH|9|8|你发现他在你面前心里忠诚，就与他立约，要把 迦南 人、 赫 人、 亚摩利 人、 比利洗 人、 耶布斯 人、 革迦撒 人之地赐给他的后裔，并且你也实现了你的话，因为你是公义的。
NEH|9|9|“‘你曾看见我们祖先在 埃及 所受的困苦，垂听他们在 红海 边的哀求，
NEH|9|10|施行神迹奇事在法老和他所有臣仆，以及他国中众百姓身上，因为你知道他们向我们祖先行事狂傲。你也得了名声，正如今日一样。
NEH|9|11|你在我们祖先面前把海分开，使他们走过海中干地，将追赶他们的人抛在深海，如石头抛在大水中。
NEH|9|12|白昼你用云柱引导他们，黑夜你用火柱照亮他们当行的路。
NEH|9|13|你降临在 西奈山 ，从天上与他们说话，赐给他们正直的典章、真实的律法、美好的律例与诫命，
NEH|9|14|又使他们知道你的圣安息日，并藉你仆人 摩西 传给他们诫命、律例、律法。
NEH|9|15|你从天上赐下粮食给他们充饥，使水从磐石流出给他们解渴。你吩咐他们进去，得你起誓应许要赐给他们的地。
NEH|9|16|“‘但我们的祖先行事狂傲，硬着颈项不听从你的诫命。
NEH|9|17|他们不肯顺从，也不记念你在他们中间所行的奇事，竟硬着颈项，居心悖逆，自立领袖，要回 埃及 他们为奴之地 。但你是乐意饶恕人，有恩惠，有怜悯，不轻易发怒，有丰盛慈爱的上帝，并没有丢弃他们。
NEH|9|18|他们虽然为自己铸了一头牛犊，说，这就是领你出 埃及 的神明，因而犯了亵渎的大罪，
NEH|9|19|你还是有丰富的怜悯，不把他们丢弃在旷野。白昼，云柱不离开他们，仍引导他们行路；黑夜，火柱仍照亮他们当行的路。
NEH|9|20|你赐下你良善的灵教导他们，没有收回吗哪不给他们吃，仍赐水给他们解渴。
NEH|9|21|在旷野四十年，你养育他们，他们一无所缺，衣服没有穿破，脚也没有肿。
NEH|9|22|你将列国和诸民族交给他们，把那些角落分给他们，他们就得了 西宏 之地，就是 希实本 王之地，和 巴珊 王 噩 之地。
NEH|9|23|你使他们的子孙多如天上的星，带他们到你对他们祖先说要进去得为业之地。
NEH|9|24|这样，这些子孙进去得了那地。你在他们面前制伏那地的居民 迦南 人，把 迦南 人和他们的君王，以及那地的民族，都交在他们手里，让他们任意处置。
NEH|9|25|他们得了坚固的城镇、肥沃的土地，取了装满各样美物的房屋、挖成的水井、葡萄园、橄榄园，以及许多果树。他们就吃了，而且饱足，身体肥胖，因你的大恩活得快乐。
NEH|9|26|“‘然而，他们不顺从，竟背叛你，将你的律法丢在背后，又杀害那些劝他们回转归向你的众先知，犯了亵渎的大罪。
NEH|9|27|所以你将他们交在敌人的手中，敌人就折磨他们。他们遭难的时候哀求你，你就从天上垂听，照你丰富的怜悯赐给他们拯救者，救他们脱离敌人的手。
NEH|9|28|但他们得享太平之后，又在你面前行恶，所以你丢弃他们，交在仇敌的手中，仇敌就辖制他们；然而他们转回哀求你，你就从天上垂听，屡次照你的怜悯拯救他们，
NEH|9|29|你警戒他们，要使他们归顺你的律法。他们却行事狂傲，不听从你的诫命，干犯你的典章，人若遵行就必因此存活。他们顽梗地扭转肩头，硬着颈项，不肯听从。
NEH|9|30|但你多年宽容他们，又以你的灵藉众先知劝戒他们，他们仍不侧耳而听，所以你将他们交在列邦民族的手中。
NEH|9|31|然而因你丰富的怜悯，你不全然灭绝他们，也不丢弃他们，因为你是有恩惠、有怜悯的上帝。
NEH|9|32|“‘现在，我们的上帝啊，你是至大、至能、至可畏、守约施慈爱的上帝；我们的君王、官长、祭司、先知、祖先和你的众百姓，从 亚述 诸王的时候直到今日所遭遇的一切苦难，求你不要看为小事。
NEH|9|33|在一切临到我们的事上，你是公义的，因为你所行的是信实，我们所做的是邪恶。
NEH|9|34|我们的君王、官长、祭司、祖先都不遵守你的律法，不听从你的诫命和你警戒他们的话。
NEH|9|35|他们在本国领受你大恩的时候，在你所赐给他们这广大肥沃之地不事奉你，也不转离他们的恶行。
NEH|9|36|看哪，我们今日成了奴仆！你赐给我们祖先享受土产和美物的地，看哪，我们在这地上竟作了奴仆！
NEH|9|37|这地许多的出产都归了诸王，就是你因我们的罪派来辖制我们的。他们任意辖制我们的身体和牲畜，我们遭了大难。’”
NEH|9|38|因这一切，我们立确实的约，写在册上。我们的领袖、 利未 人和祭司都用了印。
NEH|10|1|用印的是 哈迦利亚 的儿子 尼希米 省长、 西底家 ；
NEH|10|2|还有 西莱雅 、 亚撒利雅 、 耶利米 、
NEH|10|3|巴施户珥 、 亚玛利雅 、 玛基雅 、
NEH|10|4|哈突 、 示巴尼 、 玛鹿 、
NEH|10|5|哈琳 、 米利末 、 俄巴底亚 、
NEH|10|6|但以理 、 近顿 、 巴录 、
NEH|10|7|米书兰 、 亚比雅 、 米雅民 、
NEH|10|8|玛西亚 、 璧该 、 示玛雅 等祭司；
NEH|10|9|又有 利未 人 亚散尼 的儿子 耶书亚 、 希拿达 的子孙 宾内 、 甲篾 ，
NEH|10|10|他们的弟兄 示巴尼 、 荷第雅 、 基利他 、 毗莱雅 、 哈难 、
NEH|10|11|米迦 、 利合 、 哈沙比雅 、
NEH|10|12|撒刻 、 示利比 、 示巴尼 、
NEH|10|13|荷第雅 、 巴尼 、 比尼努 ；
NEH|10|14|还有百姓中的领袖 巴录 、 巴哈．摩押 、 以拦 、 萨土 、 巴尼 、
NEH|10|15|布尼 、 押甲 、 比拜 、
NEH|10|16|亚多尼雅 、 比革瓦伊 、 亚丁 、
NEH|10|17|亚特 、 希西家 、 押朔 、
NEH|10|18|荷第雅 、 哈顺 、 比赛 、
NEH|10|19|哈拉 、 亚拿突 、 尼拜 、
NEH|10|20|抹比押 、 米书兰 、 希悉 、
NEH|10|21|米示萨别 、 撒督 、 押杜亚 、
NEH|10|22|毗拉提 、 哈难 、 亚奈雅 、
NEH|10|23|何细亚 、 哈拿尼雅 、 哈述 、
NEH|10|24|哈罗黑 、 毗利哈 、 朔百 、
NEH|10|25|利宏 、 哈沙拿 、 玛西雅 、
NEH|10|26|亚希雅 、 哈难 、 亚难 、
NEH|10|27|玛鹿 、 哈琳 、 巴拿 。
NEH|10|28|其余的百姓、祭司、 利未 人、门口的守卫、歌唱的、殿役，所有与邻邦民族分别出来、归服上帝律法的，以及他们的妻子、儿女，凡有知识、能明白的，
NEH|10|29|都随从他们贵族的弟兄发咒起誓，要遵行上帝藉他仆人 摩西 所赐的律法，谨守遵行耶和华－我们主的一切诫命、典章、律例。
NEH|10|30|我们不把我们的女儿嫁给这地的居民，也不为我们的儿子娶他们的女儿。
NEH|10|31|这地的民族若在安息日，或什么圣日，带了货物或粮食来卖，我们必不买。每逢第七年必不耕种，凡欠我们债的必不追讨。
NEH|10|32|我们又为自己定例，每年各人捐献三分之一舍客勒，作为我们上帝殿之用：
NEH|10|33|为供饼、常献的素祭和燔祭，安息日、初一、节期所献的祭和圣物， 以色列 的赎罪祭，以及我们上帝殿里一切工作之用。
NEH|10|34|我们的祭司、 利未 人和百姓都抽签，每年按父家定期将奉献的木柴带到我们上帝的殿里，照着律法上所写的，烧在耶和华－我们上帝的坛上。
NEH|10|35|每年我们又将地上初熟的土产和各样树上初熟的果子，都奉到耶和华的殿里。
NEH|10|36|我们又照律法上所写的，将我们头胎的儿子和首生的牛羊都奉到我们上帝的殿，交给在上帝殿里供职的祭司；
NEH|10|37|并将初熟麦子所磨的面和举祭、各样树上的果子、新酒与新油奉给祭司，收在我们上帝殿的库房里，又把我们土地所产的十分之一奉给 利未 人，因 利未 人在我们一切城镇的土产中当取十分之一。
NEH|10|38|利未 人取十分之一的时候， 亚伦 的子孙中当有一个祭司与 利未 人同在。 利未 人也当从十分之一中取十分之一，奉到我们上帝的殿，收在库房的仓里。
NEH|10|39|因 以色列 人和 利未 人要把礼物，就是五谷、新酒和新油，带到收存圣所器皿的仓里，供职的祭司、门口的守卫、歌唱的都在那里。我们绝不会不顾我们上帝的殿。
NEH|11|1|百姓的领袖住在 耶路撒冷 。其余的百姓抽签，每十人中选一人来住在圣城 耶路撒冷 ，另外九人住在别的城镇。
NEH|11|2|凡甘心乐意住在 耶路撒冷 的，百姓都为他们祝福。
NEH|11|3|以色列 人、祭司、 利未 人、殿役和 所罗门 仆人的后裔都住在 犹大 的城镇，各在自己城内的地业中。本省的领袖住在 耶路撒冷 的如下：
NEH|11|4|住在 耶路撒冷 的有一些 犹大 人和 便雅悯 人。 犹大 人中有 法勒斯 的子孙 亚他雅 ； 亚他雅 是 乌西雅 的儿子， 乌西雅 是 撒迦利雅 的儿子， 撒迦利雅 是 亚玛利雅 的儿子， 亚玛利雅 是 示法提雅 的儿子， 示法提雅 是 玛勒列 的儿子；
NEH|11|5|又有 玛西雅 ； 玛西雅 是 巴录 的儿子， 巴录 是 谷．何西 的儿子， 谷．何西 是 哈赛雅 的儿子， 哈赛雅 是 亚大雅 的儿子， 亚大雅 是 约雅立 的儿子， 约雅立 是 撒迦利雅 的儿子， 撒迦利雅 是 示罗尼 的儿子；
NEH|11|6|住在 耶路撒冷 所有 法勒斯 的子孙共四百六十八名，都是勇士。
NEH|11|7|便雅悯 人中有 撒路 ； 撒路 是 米书兰 的儿子， 米书兰 是 约叶 的儿子， 约叶 是 毗大雅 的儿子， 毗大雅 是 哥赖雅 的儿子， 哥赖雅 是 玛西雅 的儿子， 玛西雅 是 以铁 的儿子， 以铁 是 耶筛亚 的儿子；
NEH|11|8|其次有 迦拜 、 撒来 ，共九百二十八名。
NEH|11|9|细基利 的儿子 约珥 是他们的长官； 哈西努亚 的儿子 犹大 是 耶路撒冷 的副长官。
NEH|11|10|祭司中有 约雅立 的儿子 耶大雅 ，又有 雅斤 ，
NEH|11|11|还有管理上帝殿的 西莱雅 ； 西莱雅 是 希勒家 的儿子， 希勒家 是 米书兰 的儿子， 米书兰 是 撒督 的儿子， 撒督 是 米拉约 的儿子， 米拉约 是 亚希突 的儿子；
NEH|11|12|还有他们的弟兄在殿里供职的，共八百二十二名；又有 亚大雅 ； 亚大雅 是 耶罗罕 的儿子， 耶罗罕 是 毗拉利 的儿子， 毗拉利 是 暗洗 的儿子， 暗洗 是 撒迦利亚 的儿子， 撒迦利亚 是 巴施户珥 的儿子， 巴施户珥 是 玛基雅 的儿子；
NEH|11|13|还有他的弟兄作族长的，共二百四十二名；又有 亚玛帅 ； 亚玛帅 是 亚萨列 的儿子， 亚萨列 是 亚哈赛 的儿子， 亚哈赛 是 米实利末 的儿子， 米实利末 是 音麦 的儿子；
NEH|11|14|还有他们的弟兄，大能的勇士共一百二十八名； 哈基多琳 的儿子 撒巴第业 是他们的长官。
NEH|11|15|利未 人中有 示玛雅 ； 示玛雅 是 哈述 的儿子， 哈述 是 押利甘 的儿子， 押利甘 是 哈沙比雅 的儿子， 哈沙比雅 是 布尼 的儿子；
NEH|11|16|又有 利未 人的族长 沙比太 和 约撒拔 管理上帝殿外面的事务；
NEH|11|17|祈祷的时候， 玛他尼 是主礼，开始称谢； 玛他尼 是 米迦 的儿子， 米迦 是 撒底 的儿子， 撒底 是 亚萨 的儿子；又有 玛他尼 弟兄中的 八布迦 为副；还有 押大 ； 押大 是 沙母亚 的儿子， 沙母亚 是 加拉 的儿子， 加拉 是 耶杜顿 的儿子；
NEH|11|18|在圣城所有的 利未 人共二百八十四名。
NEH|11|19|门口的守卫是 亚谷 和 达们 ，以及他们的弟兄，看守各门，共一百七十二名。
NEH|11|20|其余的 以色列 人、祭司、 利未 人都住在 犹大 一切的城镇，各在自己的地业中。
NEH|11|21|殿役却住在 俄斐勒 ； 西哈 和 基斯帕 管理他们。
NEH|11|22|在 耶路撒冷 ， 利未 人的长官，管理上帝殿事务的是歌唱者 亚萨 的子孙 乌西 ； 乌西 是 巴尼 的儿子， 巴尼 是 哈沙比雅 的儿子， 哈沙比雅 是 玛他尼 的儿子， 玛他尼 是 米迦 的儿子。
NEH|11|23|王为歌唱者下命令，确定他们每日当办的事 。
NEH|11|24|犹大 的儿子 谢拉 的子孙， 米示萨别 的儿子 毗他希雅 辅助王办理百姓一切的事。
NEH|11|25|至于村庄和所属的田地，有 犹大 人住在 基列．亚巴 和所属的乡镇 、 底本 和所属的乡镇、 叶甲薛 和所属的村庄、
NEH|11|26|耶书亚 、 摩拉大 、 伯．帕列 、
NEH|11|27|哈萨．书亚 、 别是巴 和所属的乡镇、
NEH|11|28|洗革拉 、 米哥拿 和所属的乡镇、
NEH|11|29|隐．临门 、 琐拉 、 耶末 、
NEH|11|30|撒挪亚 、 亚杜兰 和属它们的村庄、 拉吉 和所属的田地、 亚西加 和所属的乡镇；他们所住的地方是从 别是巴 直到 欣嫩谷 。
NEH|11|31|便雅悯 人从 迦巴 起，住在 密抹 、 亚雅 、 伯特利 和所属的乡镇、
NEH|11|32|亚拿突 、 挪伯 、 亚难雅 、
NEH|11|33|夏琐 、 拉玛 、 基他音 、
NEH|11|34|哈第 、 洗编 、 尼八拉 、
NEH|11|35|罗德 、 阿挪 、 革．夏纳欣 。
NEH|11|36|在 犹大 地区的 利未 人中，有些已归属 便雅悯 。
NEH|12|1|这些是同 撒拉铁 的儿子 所罗巴伯 以及 耶书亚 一起上来的祭司和 利未 人： 西莱雅 、 耶利米 、 以斯拉 、
NEH|12|2|亚玛利雅 、 玛鹿 、 哈突 、
NEH|12|3|示迦尼 、 利宏 、 米利末 、
NEH|12|4|易多 、 近顿 、 亚比雅 、
NEH|12|5|米雅民 、 玛底雅 、 璧迦 、
NEH|12|6|示玛雅 、 约雅立 、 耶大雅 、
NEH|12|7|撒路 、 亚木 、 希勒家 、 耶大雅 ；这些人在 耶书亚 的时代作祭司和他们弟兄的领袖。
NEH|12|8|利未 人有 耶书亚 、 宾内 、 甲篾 、 示利比 、 犹大 、 玛他尼 ； 玛他尼 和他的弟兄负责赞美诗歌。
NEH|12|9|他们的弟兄 八布迦 和 乌尼 按照班次站在他们的对面。
NEH|12|10|耶书亚 生 约雅金 ， 约雅金 生 以利亚实 ， 以利亚实 生 耶何耶大 ，
NEH|12|11|耶何耶大 生 约拿单 ， 约拿单 生 押杜亚 。
NEH|12|12|在 约雅金 的时代，祭司作族长的， 西莱雅 族有 米拉雅 ， 耶利米 族有 哈拿尼雅 ，
NEH|12|13|以斯拉 族有 米书兰 ， 亚玛利雅 族有 约哈难 ，
NEH|12|14|米利古 族有 约拿单 ， 示巴尼 族有 约瑟 ，
NEH|12|15|哈琳 族有 押拿 ， 米拉约 族有 希勒恺 ，
NEH|12|16|易多 族有 撒迦利亚 ， 近顿 族有 米书兰 ，
NEH|12|17|亚比雅 族有 细基利 ， 米拿民 族， 摩亚底 族有 毗勒太 ，
NEH|12|18|璧迦 族有 沙母亚 ， 示玛雅 族有 约拿单 ，
NEH|12|19|约雅立 族有 玛特乃 ， 耶大雅 族有 乌西 ，
NEH|12|20|撒来 族有 加莱 ， 亚木 族有 希伯 ，
NEH|12|21|希勒家 族有 哈沙比雅 ， 耶大雅 族有 拿坦业 。
NEH|12|22|在 以利亚实 、 耶何耶大 、 约哈难 、 押杜亚 的时代， 利未 人的族长都记在册上，祭司也一样，直到 波斯 王 大流士 在位的时候。
NEH|12|23|利未 人作族长的记在史籍上，一直记到 以利亚实 的儿子 约哈难 的时代。
NEH|12|24|利未 人的族长是 哈沙比雅 、 示利比 、 甲篾 的儿子 耶书亚 ，他们的弟兄站在他们的对面，照神人 大卫 的命令按着班次赞美称谢。
NEH|12|25|玛他尼 、 八布迦 、 俄巴底亚 、 米书兰 、 达们 、 亚谷 是门口的守卫，在库房的门口站岗。
NEH|12|26|这些人都在 约撒达 的孙子， 耶书亚 的儿子 约雅金 和 尼希米 省长，以及 以斯拉 祭司文士的时代供职。
NEH|12|27|为 耶路撒冷 城墙行奉献礼的时候，众人把各处的 利未 人召到 耶路撒冷 ，要以称谢、歌唱、敲钹、鼓瑟、弹琴，喜乐地行奉献礼。
NEH|12|28|歌唱的人从 耶路撒冷 的周围聚集，从 尼陀法 人的村庄、
NEH|12|29|伯．吉甲 ，以及 迦巴 和 亚斯玛弗 的田地而来；因为歌唱的人在 耶路撒冷 四围为自己建立了村庄。
NEH|12|30|祭司和 利未 人就洁净自己，也洁净百姓，以及城门和城墙。
NEH|12|31|我带 犹大 的领袖上城墙，把称谢的人分为两大队，在城墙上往右边的 粪厂门 行进，
NEH|12|32|在他们后面行进的有 何沙雅 与 犹大 一半的领袖，
NEH|12|33|又有 亚撒利雅 、 以斯拉 、 米书兰 、
NEH|12|34|犹大 、 便雅悯 、 示玛雅 、 耶利米 。
NEH|12|35|还有祭司的子孙，吹号的有 撒迦利亚 ； 撒迦利亚 是 约拿单 的儿子， 约拿单 是 示玛雅 的儿子， 示玛雅 是 玛他尼 的儿子， 玛他尼 是 米该亚 的儿子， 米该亚 是 撒刻 的儿子， 撒刻 是 亚萨 的儿子；
NEH|12|36|又有 撒迦利亚 的弟兄 示玛雅 、 亚撒利 、 米拉莱 、 基拉莱 、 玛艾 、 拿坦业 、 犹大 、 哈拿尼 ，各拿着神人 大卫 的乐器，由 以斯拉 文士在前面引领。
NEH|12|37|他们经过 泉门 往前，登 大卫城 的台阶，上城墙的斜坡，从 大卫 宫殿之上，直到朝东的 水门 。
NEH|12|38|第二队称谢的人要往反方向而行。我和一半的百姓在城墙上跟随他们，从 炉楼 之上，直到 宽墙 ；
NEH|12|39|又过了 以法莲门 、 古门 、 鱼门 、 哈楠业楼 、 哈米亚楼 ，直到 羊门 ，就在 护卫门 站住。
NEH|12|40|于是，这两队称谢的人连同我和一半跟随我的官长，站在上帝的殿里。
NEH|12|41|还有 以利亚金 、 玛西雅 、 米拿民 、 米该亚 、 以利约乃 、 撒迦利亚 、 哈楠尼亚 等吹号的祭司；
NEH|12|42|又有 玛西雅 、 示玛雅 、 以利亚撒 、 乌西 、 约哈难 、 玛基雅 、 以拦 和 以谢 。歌唱的大声唱歌，有 伊斯拉希雅 作指挥。
NEH|12|43|那日，众人献上丰盛的祭物，并且欢乐，因为上帝使他们大大欢乐，连妇女带孩童也都欢乐，甚至从远处都可听到 耶路撒冷 的欢声。
NEH|12|44|当日，有些人受派管理库房，把举祭、初熟之物，和所取的十一奉献，按各城的田地，照律法所定，归给祭司和 利未 人的份，都收在库房里。 犹大 人因祭司和 利未 人供职就欢乐。
NEH|12|45|祭司和 利未 人遵守上帝所吩咐的，守洁净礼。歌唱的和门口的守卫照着 大卫 和他儿子 所罗门 的命令也如此行。
NEH|12|46|古时，在 大卫 和 亚萨 的日子，有歌唱者的指挥，也有赞美称谢上帝的诗歌。
NEH|12|47|在 所罗巴伯 和 尼希米 的时代， 以色列 众人把歌唱者和门口的守卫每日当得的份供给他们，又把给 利未 人的分别出来； 利未 人又把给 亚伦 子孙的分别出来。
NEH|13|1|在那日，百姓听到人朗读 摩西 的律法书，发现书上写着， 亚扪 人和 摩押 人永不可入上帝的会；
NEH|13|2|因为他们没有拿食物和水来迎接 以色列 人，却雇了 巴兰 诅咒他们，但我们的上帝使那诅咒变为祝福。
NEH|13|3|以色列 人听见这律法，就与所有不同族群的人分别出来。
NEH|13|4|在这之前，与 多比雅 结亲的 以利亚实 祭司，受派管理我们上帝殿中的库房，
NEH|13|5|为 多比雅 预备了一间大屋子，就是从前收存素祭、乳香、器皿，和照例供给 利未 人、歌唱者、门口守卫的五谷、新酒和新油的十分之一，以及归祭司之举祭的屋子。
NEH|13|6|当这一切事发生的时候，我不在 耶路撒冷 ，因为 巴比伦 王 亚达薛西 三十二年，我回到王那里。过了多日，我又向王告假。
NEH|13|7|我来到 耶路撒冷 ，才知道 以利亚实 为 多比雅 所做、在上帝殿的院内为他预备屋子的那件恶事。
NEH|13|8|我非常愤怒，就把 多比雅 的一切家具都从屋子里抛出去。
NEH|13|9|我又吩咐人洁净这屋子，然后将上帝殿的器皿、素祭和乳香搬回那里。
NEH|13|10|我发现 利未 人当得的份无人供给他们，甚至供职的 利未 人与歌唱的都各奔回自己的田地去了。
NEH|13|11|我就斥责官长说：“你们为何不顾上帝的殿呢？”于是我召集 利未 人，使他们在自己的岗位上供职。
NEH|13|12|犹大 众人就把五谷、新酒和新油的十分之一送入库房。
NEH|13|13|我派 示利米雅 祭司、 撒督 文士和 利未 人 毗大雅 作司库管理库房，副手是 哈难 ； 哈难 是 撒刻 的儿子， 撒刻 是 玛他尼 的儿子；这些人都是忠实的，他们的职务是分派他们弟兄所当得的份。
NEH|13|14|我的上帝啊，求你因这事记念我，不要涂去我为上帝的殿与其中的礼仪所献的忠心。
NEH|13|15|那些日子，我在 犹大 见有人在安息日踹醡酒池，搬运禾捆驮在驴上，又把酒、葡萄、无花果和各样的担子在安息日扛入 耶路撒冷 ，我就在他们卖食物的那日警戒他们。
NEH|13|16|有一些住在城里的 推罗 人也把鱼和各样货物运进来，甚至在 耶路撒冷 ，在安息日卖给 犹大 人。
NEH|13|17|我就斥责 犹大 的贵族，对他们说：“你们怎么会做这恶事干犯安息日呢！
NEH|13|18|你们祖先岂不是这样做，以致我们的上帝使一切灾祸临到我们和这城吗？你们竟干犯安息日，使愤怒越发临到 以色列 ！”
NEH|13|19|安息日前一日黄昏的时候，我吩咐人把 耶路撒冷 城门锁上；我又吩咐，不过安息日不准开门。我也派几个仆人在城门口站岗，免得有人在安息日挑担子进城。
NEH|13|20|于是商人和贩卖各样货物的人，有一两次在 耶路撒冷 城外过夜。
NEH|13|21|我警告他们说：“你们为何在城墙前过夜呢？若再这样，我必下手办你们。”从此以后，他们在安息日就不再来了。
NEH|13|22|我吩咐 利未 人洁净自己来守城门，使安息日分别为圣。我的上帝啊，求你因这事记念我，照你丰盛的慈爱怜悯我。
NEH|13|23|那些日子，我又看见 犹太 人娶了 亚实突 、 亚扪 和 摩押 的女子为妻。
NEH|13|24|他们的儿女，一半说 亚实突 话，或其他种族的方言，不会说 犹大 话。
NEH|13|25|我就斥责他们，诅咒他们，打了他们几个人，拔下他们的胡须，叫他们指着上帝起誓：“你们不可把自己的女儿嫁给外邦人的儿子，也不可为自己和儿子娶他们的女儿。
NEH|13|26|以色列 王 所罗门 不也在这样的事上犯罪吗？在许多国家中并没有一位王像他，蒙他上帝喜爱，上帝立他作王治理全 以色列 。然而，连他也被外邦女子引诱犯罪。
NEH|13|27|我们岂能听凭你们行这一切大恶，娶外邦女子干犯我们的上帝呢？”
NEH|13|28|以利亚实 大祭司的孙子， 耶何耶大 的一个儿子是 和伦 人 参巴拉 的女婿，我就把他从我这里赶出去。
NEH|13|29|我的上帝啊，求你记得他们的罪，因为他们玷污了祭司的职分，违背祭司和 利未 人的约。
NEH|13|30|这样，我洁净他们，使他们脱离属外邦人的一切；我又分派祭司和 利未 人的班次，使他们各尽其职，
NEH|13|31|按定期奉献木柴和初熟的土产。我的上帝啊，求你记念我，施恩于我。
