HEB|1|1|Багато разів і багатьма способами в давнину промовляв був Бог до отців через пророків,
HEB|1|2|а в останні ці дні промовляв Він до нас через Сина, що Його настановив за Наслідника всього, що Ним і віки Він створив.
HEB|1|3|Він був сяєвом слави та образом істоти Його, тримав усе словом сили Своєї, учинив Собою очищення наших гріхів, і засів на правиці величности на висоті.
HEB|1|4|Він остільки був ліпший понад Анголів, оскільки славніше за них успадкував Ім'я.
HEB|1|5|Кому бо коли з Анголів Він промовив: Ти Мій Син, Я сьогодні Тебе породив! І знову: Я буду Йому за Отця, а Він Мені буде за Сина!
HEB|1|6|І коли знов Він уводить на світ Перворідного, то говорить: І нехай Йому вклоняться всі Анголи Божі.
HEB|1|7|А про Анголів Він говорить: Ти чиниш духів Анголами Своїми, а палючий огонь Своїми слугами.
HEB|1|8|А про Сина: Престол Твій, о Боже, навік віку; берло Твого царювання берло праведности.
HEB|1|9|Ти полюбив праведність, а беззаконня зненавидів; через це намастив Тебе, Боже, Твій Бог оливою радости більше, ніж друзів Твоїх.
HEB|1|10|І: Ти, Господи, землю колись заклав, а небо то чин Твоїх рук.
HEB|1|11|Загинуть вони, а Ти будеш стояти, всі вони, як той одяг, постаріють.
HEB|1|12|Як одежу, їх зміниш, і минуться вони, а Ти завжди Той Самий, і роки Твої не закінчаться!
HEB|1|13|Кому з Анголів Він промовив коли: Сядь праворуч Мене, доки не покладу Я Твоїх ворогів підніжком ногам Твоїм!
HEB|1|14|Чи не всі вони духи служебні, що їх посилають на службу для тих, хто має спасіння вспадкувати?
HEB|2|1|Через це подобає нам більше вважати на почуте, щоб ми не відпали коли.
HEB|2|2|Коли бо те слово, що сказали його Анголи, було певне, а всякий переступ та непослух прийняли справедливу заплату,
HEB|2|3|то як ми втечемо, коли ми не дбали про таке велике спасіння? Воно проповідувалося спочатку від Господа, ствердилося нам через тих, хто почув,
HEB|2|4|коли Бог був засвідчив ознаками й чудами, і різними силами та обдаруванням Духом Святим із волі Своєї.
HEB|2|5|Бо Він не піддав Анголам світ майбутній, що про нього говоримо.
HEB|2|6|Але хтось десь засвідчив був, кажучи: Що є чоловік, що Ти пам'ятаєш про нього, і син людський, якого відвідуєш?
HEB|2|7|Ти його вчинив мало меншим від Анголів, і честю й величністю Ти вінчаєш його, і поставив його над ділами рук Своїх,
HEB|2|8|усе піддав Ти під ноги йому! А коли Він піддав йому все, то не залишив нічого йому непідданого. А тепер ще не бачимо, щоб піддане було йому все.
HEB|2|9|Але бачимо Ісуса, мало чим уменшеним від Анголів, що за перетерплення смерти Він увінчаний честю й величністю, щоб за благодаттю Божою смерть скуштувати за всіх.
HEB|2|10|Бо належало, щоб Той, що все ради Нього й усе від Нього, Хто до слави привів багато синів, Провідника їхнього спасіння вчинив досконалим через страждання.
HEB|2|11|Бо Хто освячує, і ті, хто освячується усі від Одного. З цієї причини не соромиться Він звати братами їх, кажучи:
HEB|2|12|Сповіщу про Ім'я Твоє браттям Своїм, буду хвалити Тебе серед Церкви!
HEB|2|13|І ще: На Нього я буду надіятися! І ще: Ото Я та діти, яких Бог Мені дав.
HEB|2|14|А що діти стали спільниками тіла та крови, то й Він став учасником їхнім, щоб смертю знищити того, хто має владу смерти, цебто диявола,
HEB|2|15|та визволити тих усіх, хто все життя страхом смерти тримався в неволі.
HEB|2|16|Бо приймає Він не Анголів, але Авраамове насіння.
HEB|2|17|Тому мусів бути Він у всьому подібний братам, щоб стати милостивим та вірним Первосвящеником у Божих справах, для вблагання за гріхи людей.
HEB|2|18|Бо в чому був Сам постраждав, випробовуваний, у тому Він може й випробовуваним помогти.
HEB|3|1|Отож, святі брати, учасники небесного покликання, уважайте на Апостола й Первосвященика нашого ісповідання, Ісуса,
HEB|3|2|що вірний Тому, Хто настановив Його, як був і Мойсей у всім домі Його,
HEB|3|3|бо гідний Він вищої слави понад Мойсея, поскільки будівничий має більшу честь, аніж дім.
HEB|3|4|Усякий бо дім хтось будує, а Той, хто все збудував, то Бог.
HEB|3|5|І Мойсей вірний був у всім домі Його, як слуга, на свідоцтво того, що сказати повинно було.
HEB|3|6|Христос же, як Син, у Його домі. А дім Його ми, коли тільки відвагу й похвалу надії додержимо певними аж до кінця.
HEB|3|7|Тому то, як каже Дух Святий: Сьогодні, як голос Його ви почуєте,
HEB|3|8|не робіть затверділими ваших сердець, як під час нарікань, за дня випробовування на пустині,
HEB|3|9|де Мене випробовували отці ваші, Мене випробовували, і бачили працю Мою сорок років.
HEB|3|10|Через це Я розгнівався був на той рід і сказав: Постійно вони блудять серцем, вони не пізнали доріг Моїх,
HEB|3|11|тому Я присягнув був у гніві Своїм, що вони до Мого відпочинку не ввійдуть!
HEB|3|12|Стережіться, брати, щоб у комусь із вас не було злого серця невірства, що воно відступало б від Бога Живого!
HEB|3|13|Але кожного дня заохочуйте один одного, доки зветься Сьогодні, щоб запеклим не став котрий з вас через підступ гріха.
HEB|3|14|Бо ми стали учасниками Христа, коли тільки почате життя ми затримаємо певним аж до кінця,
HEB|3|15|аж поки говориться: Сьогодні, як голос Його ви почуєте, не робіть затверділими ваших сердець, як під час нарікань!
HEB|3|16|Котрі бо, почувши, розгнівали Бога? Чи не всі, хто з Єгипту вийшов з Мойсеєм?
HEB|3|17|На кого ж Він гнівався був сорок років? Хіба не на тих, хто згрішив, що їхні кості в пустині полягли?
HEB|3|18|Проти кого Він був присягався, що не ввійдуть вони до Його відпочинку, як не проти неслухняних?
HEB|3|19|І ми бачимо, що вони не змогли ввійти за невірство.
HEB|4|1|Отже, біймося, коли зостається обітниця входу до Його відпочинку, щоб не виявилось, що хтось із вас опізнився.
HEB|4|2|Бо Євангелія була звіщена нам, як і тим. Але не принесло пожитку їм слово почуте, бо воно не злучилося з вірою слухачів.
HEB|4|3|Бо до Його відпочинку входимо ми, що ввірували, як Він провістив: Я присяг був у гніві Своїм, що до місця Мого відпочинку не ввійдуть вони, хоч діла Його були вчинені від закладин світу.
HEB|4|4|Бо колись про день сьомий сказав Він отак: І Бог відпочив сьомого дня від усієї праці Своєї.
HEB|4|5|А ще тут: До Мого відпочинку не ввійдуть вони!
HEB|4|6|Коли ж залишається ото, що деякі ввійдуть до нього, а ті, кому Євангелія була перше звіщена, не ввійшли за непослух,
HEB|4|7|то ще призначає Він деякий день, сьогодні, бо через Давида говорить по такім довгім часі, як вище вже сказано: Сьогодні, як голос Його ви почуєте, не робіть затверділими ваших сердець!
HEB|4|8|Бо коли б Ісус Навин дав їм відпочинок, то про інший день не казав би по цьому.
HEB|4|9|Отож, людові Божому залишається суботство, спочинок.
HEB|4|10|Хто бо ввійшов був у Його відпочинок, то й той відпочив від учинків своїх, як і Бог від Своїх.
HEB|4|11|Отож, попильнуймо ввійти до того відпочинку, щоб ніхто не потрапив у непослух за прикладом тим.
HEB|4|12|Бо Боже Слово живе та діяльне, гостріше від усякого меча обосічного, проходить воно аж до поділу душі й духа, суглобів та мозків, і спосібне судити думки та наміри серця.
HEB|4|13|І немає створіння, щоб сховалось перед Ним, але все наге та відкрите перед очима Його, Йому дамо звіт!
HEB|4|14|Отож, мавши великого Первосвященика, що небо перейшов, Ісуса, Сина Божого, тримаймося ісповідання нашого!
HEB|4|15|Бо ми маємо не такого Первосвященика, що не міг би співчувати слабостям нашим, але випробуваного в усьому, подібно до нас, окрім гріха.
HEB|4|16|Отож, приступаймо з відвагою до престолу благодаті, щоб прийняти милість та для своєчасної допомоги знайти благодать.
HEB|5|1|Кожен бо первосвященик, що з-між людей вибирається, настановляється для людей на служіння Богові, щоб приносити дари та жертви за гріхи,
HEB|5|2|і щоб міг співчувати недосвідченим та заблудженим, бо й сам він перейнятий слабістю.
HEB|5|3|І тому він повинен як за людей, так само й за себе самого приносити жертви за гріхи.
HEB|5|4|А чести цієї ніхто не бере сам собою, а покликаний Богом, як і Аарон.
HEB|5|5|Так і Христос, не Сам Він прославив Себе, щоб Первосвящеником стати, а Той, що до Нього сказав: Ти Мій Син, Я сьогодні Тебе породив.
HEB|5|6|Як і на іншому місці говорить: Ти Священик навіки за чином Мелхиседековим.
HEB|5|7|Він за днів тіла Свого з голосінням великим та слізьми приніс був благання й молитви до Того, хто від смерти Його міг спасти, і був вислуханий за побожність Свою.
HEB|5|8|І хоч Сином Він був, проте навчився послуху з того, що вистраждав був.
HEB|5|9|А вдосконалившися, Він для всіх, хто слухняний Йому, спричинився для вічного спасіння,
HEB|5|10|і від Бога був названий Первосвящеником за чином Мелхиседековим.
HEB|5|11|Про це нам би треба багато казати, та висловити важко його, бо нездібні ви стали, щоб слухати.
HEB|5|12|Ви бо за віком повинні б бути вчителями, але ви потребуєте ще, щоб хтось вас навчав перших початків Божого Слова. І ви стали такими, яким потрібне молоко, а не страва тверда.
HEB|5|13|Бо хто молока вживає, той недосвідчений у слові правди, бо він немовля.
HEB|5|14|А страва тверда для дорослих, що мають чуття, привчені звичкою розрізняти добро й зло.
HEB|6|1|Тому полишімо початки науки Христа, та й звернімося до досконалости, і не кладімо знову засади покаяння від мертвих учинків та про віру в Бога,
HEB|6|2|науки про хрищення, про покладання рук, про воскресіння мертвих та вічний суд.
HEB|6|3|Зробимо й це, коли Бог дозволить.
HEB|6|4|Не можна бо тих, що раз просвітились були, і скуштували небесного дару, і стали причасниками Духа Святого,
HEB|6|5|і скуштували доброго Божого Слова та сили майбутнього віку,
HEB|6|6|та й відпали, знов відновляти покаянням, коли вдруге вони розпинають у собі Сина Божого та зневажають.
HEB|6|7|Бо земля, що п'є дощ, який падає часто на неї, і родить рослини, добрі для тих, хто їх і вирощує, вона благословення від Бога приймає.
HEB|6|8|Але та, що приносить терня й будяччя, непотрібна вона та близька до прокляття, а кінець її спалення.
HEB|6|9|Та ми сподіваємось, любі, кращого про вас, що спасіння тримаєтеся, хоч говоримо й так.
HEB|6|10|Та не є Бог несправедливий, щоб забути діло ваше та працю любови, яку показали в Ім'я Його ви, що святим послужили та служите.
HEB|6|11|Ми ж бажаємо, щоб кожен із вас виявляв таку саму завзятість на певність надії аж до кінця,
HEB|6|12|щоб ви не розлінились, але переймали від тих, хто обітниці вспадковує вірою та терпеливістю.
HEB|6|13|Бо Бог, обітницю давши Авраамові, як не міг ніким вищим поклястися, поклявся Сам Собою,
HEB|6|14|говорячи: Поблагословити Я конче тебе поблагословлю, та розмножити розмножу тебе!
HEB|6|15|І, терплячи довго отак, Авраам одержав обітницю.
HEB|6|16|Бо люди клянуться вищим, і клятва на ствердження кінчає всяку їхню суперечку.
HEB|6|17|Тому й Бог, хотівши переважно показати спадкоємцям обітниці незмінність волі Своєї, учинив те при помочі клятви,
HEB|6|18|щоб у двох тих незмінних речах, що в них не можна сказати неправди Богові, мали потіху міцну ми, хто прибіг прийняти надію, що лежить перед нами,
HEB|6|19|що вони для душі як котвиця, міцна та безпечна, що аж до середини входить за заслону,
HEB|6|20|куди, як предтеча, за нас увійшов був Ісус, ставши навіки Первосвящеником за чином Мелхиседековим.
HEB|7|1|Бо цей Мелхиседек, цар Салиму, священик Бога Всевишнього, що був стрів Авраама, як той вертався по поразці царів, і його поблагословив.
HEB|7|2|Авраам відділив йому й десятину від усього, найперше бо він визначає цар правди, а потім цар Салиму, цебто цар миру.
HEB|7|3|Він без батька, без матері, без родоводу, не мав ані початку днів, ані кінця життя, уподобився Божому Сину, пробуває священиком завжди.
HEB|7|4|Побачте ж, який він великий, що йому й десятину з добичі найліпшої дав патріярх Авраам!
HEB|7|5|Ті з синів Левієвих, що священство приймають, мають заповідь брати за Законом десятину з народу, цебто з братів своїх, хоч і вийшли вони з Авраамових стегон.
HEB|7|6|Але цей, що не походить з їхнього роду, десятину одержав від Авраама, і поблагословив того, хто обітницю мав.
HEB|7|7|І без усякої суперечки більший меншого благословляє.
HEB|7|8|І тут люди смертельні беруть десятину, а там той, про якого засвідчується, що живе.
HEB|7|9|І, щоб сказати отак, через Авраама і Левій, що бере десятини, дав сам десятини.
HEB|7|10|Бо ще в батькових стегнах він був, коли стрів його Мелхиседек.
HEB|7|11|Отож, коли б досконалість була через священство левитське, бо люди Закона одержали з ним, то яка ще потреба була, щоб Інший Священик повстав за чином Мелхиседековим, а не зватися за чином Аароновим?
HEB|7|12|Коли бо священство зміняється, то з потреби буває переміна й Закону.
HEB|7|13|Бо Той, що про Нього говориться це, належав до іншого племени, з якого ніхто не ставав був до жертівника.
HEB|7|14|Бож відомо, що Господь наш походить від Юди, а про це плем'я, про священство його, нічого Мойсей не сказав.
HEB|7|15|І ще більше відомо, коли повстає на подобу Мелхиседека Інший Священик,
HEB|7|16|що був не за законом тілесної заповіді, але з сили незнищального життя.
HEB|7|17|Бо свідчить: Ти Священик навіки за чином Мелхиседековим.
HEB|7|18|Попередня бо заповідь відкладається через неміч її та некорисність.
HEB|7|19|Бо не вдосконалив нічого Закон. Запроваджена ж краща надія, що нею ми наближуємось до Бога.
HEB|7|20|І поскільки воно не без клятви,
HEB|7|21|вони бо без клятви були священиками, Цей же з клятвою через Того, Хто говорить до Нього: Клявся Господь і не буде Він каятися: Ти Священик навіки за чином Мелхиседековим,
HEB|7|22|то постільки Ісус став запорукою кращого Заповіту!
HEB|7|23|І багато було їх священиків, бо смерть боронила лишатися їм,
HEB|7|24|але Цей, що навіки лишається, безперестанне Священство Він має.
HEB|7|25|Тому може Він завжди й спасати тих, хто через Нього до Бога приходить, бо Він завжди живий, щоб за них заступитись.
HEB|7|26|Отакий бо потрібний нам Первосвященик: святий, незлобивий, невинний, відлучений від грішників, що вищий над небеса,
HEB|7|27|що потреби не має щодня, як ті первосвященики, перше приносити жертви за власні гріхи, а потому за людські гріхи, бо Він це раз назавжди вчинив, принісши Самого Себе.
HEB|7|28|Закон бо людей ставить первосвящениками, що немочі мають, але слово клятви, що воно за Законом, ставить Сина, Який досконалий навіки!
HEB|8|1|Головна ж річ у тому, про що я говорю: маємо Первосвященика, що засів на небесах, по правиці престолу величности,
HEB|8|2|що Він Священнослужитель святині й правдивої скинії, що її збудував був Господь, а не людина.
HEB|8|3|Усякий бо первосвященик настановляється, щоб приносити дари та жертви, а тому було треба, щоб і Цей щось мав, що принести.
HEB|8|4|Бо коли б на землі перебував, то не був би Він священиком, бо тут пробувають священики, що дари приносять за Законом.
HEB|8|5|Вони служать образові й тіні небесного, як Мойсеєві сказано, коли мав докінчити скинію: Дивись бо, сказав, зроби все за зразком, що тобі на горі був показаний!
HEB|8|6|А тепер одержав Він краще служіння, поскільки Він посередник і кращого заповіту, який на кращих обітницях був узаконений.
HEB|8|7|Бо коли б отой перший був бездоганний, не шукалося б місця для другого.
HEB|8|8|Бо їм докоряючи, каже: Ото дні надходять, говорить Господь, коли з домом Ізраїля й з Юдиним домом Я складу Заповіта Нового,
HEB|8|9|не за заповітом, що його Я склав був з отцями їхніми дня, коли взяв їх за руку, щоб вивести їх із землі єгипетської. А що вони не залишилися в Моїм заповіті, то й Я їх покинув, говорить Господь!
HEB|8|10|Оце Заповіт, що його Я складу по тих днях із домом Ізраїлевим, говорить Господь: Покладу Я Закони Свої в їхні думки, і на їхніх серцях напишу їх, і буду їм Богом, вони ж будуть народом Моїм!
HEB|8|11|І кожен не буде навчати свого ближнього, і кожен брата свого, промовляючи: Пізнай Господа! Усі бо вони будуть знати Мене від малого та аж до великого з них!
HEB|8|12|Буду бо Я милостивий до їхніх неправд, і їхніх гріхів не згадаю Я більш!
HEB|8|13|Коли ж каже Новий Заповіт, то тим назвав перший старим. А що порохнявіє й старіє, те близьке до зотління.
HEB|9|1|Мав же і перший заповіт постанови богослужби та світську святиню.
HEB|9|2|Була бо уряджена перша скинія, яка зветься святиня, а в ній був свічник, і стіл, і жертвенні хліби.
HEB|9|3|А за другою заслоною скинія, що зветься Святеє Святих.
HEB|9|4|Мала вона золоту кадильницю й ковчега заповіту, усюди обкутого золотом, а в нім золота посудина з манною, і розцвіле жезло Ааронове та таблиці заповіту.
HEB|9|5|А над ним херувими слави, що затінювали престола благодаті, про що говорити докладно тепер не потрібно.
HEB|9|6|При такому ж урядженні до першої скинії входили завжди священики, правлячи служби Богові,
HEB|9|7|а до другої раз на рік сам первосвященик, не без крови, яку він приносить за себе й за людські провини.
HEB|9|8|Святий Дух виявляє оцим, що ще не відкрита дорога в святиню, коли ще стоїть перша скинія.
HEB|9|9|Вона образ для часу теперішнього, за якого приносяться дари та жертви, що того не можуть вдосконалити, щодо сумління того, хто служить,
HEB|9|10|що тільки в потравах та в напоях, та в різних обмиваннях, в уставах тілесних, установлено їх аж до часу направи.
HEB|9|11|Але Христос, Первосвященик майбутнього доброго, прийшов із більшою й досконалішою скинією, нерукотворною, цебто не цього втворення,
HEB|9|12|і не з кров'ю козлів та телят, але з власною кров'ю увійшов до святині один раз, та й набув вічне відкуплення.
HEB|9|13|Бо коли кров козлів та телят та попіл із ялівок, як покропить нечистих, освячує їх на очищення тіла,
HEB|9|14|скільки ж більш кров Христа, що Себе непорочного Богу приніс Святим Духом, очистить наше сумління від мертвих учинків, щоб служити нам Богові Живому!
HEB|9|15|Тому Він Посередник Нового Заповіту, щоб через смерть, що була для відкуплення від переступів, учинених за першого заповіту, покликані прийняли обітницю вічного спадку.
HEB|9|16|Бо де заповіт, там має відбутися смерть заповітника,
HEB|9|17|заповіт бо важливий по мертвих, бо нічого не варт він, як живе заповітник.
HEB|9|18|Тому й перший заповіт освячений був не без крови:
HEB|9|19|Коли бо Мойсей сповістив був усі заповіді за Законом усьому народові, він узяв кров козлів та телят із водою й червоною вовною та з ісопом, та й покропив і саму оту книгу, і людей,
HEB|9|20|проказуючи: Це кров заповіту, що його наказав для вас Бог!
HEB|9|21|Так само і скинію, і ввесь посуд служебний покропив він кров'ю.
HEB|9|22|І майже все за Законом кров'ю очищується, а без пролиття крови не має відпущення.
HEB|9|23|Отож, треба було, щоб образи небесного очищалися цими, а небесне саме кращими від оцих жертвами.
HEB|9|24|Бо Христос увійшов не в рукотворну святиню, що була на взір правдивої, але в саме небо, щоб з'явитись тепер перед Божим лицем за нас,
HEB|9|25|і не тому, щоб часто приносити в жертву Себе, як первосвященик увіходить у святиню кожнорічно із кров'ю чужою,
HEB|9|26|бо інакше Він мусів би часто страждати ще від закладин світу, а тепер Він з'явився один раз на схилку віків, щоб власною жертвою знищити гріх.
HEB|9|27|І як людям призначено вмерти один раз, потім же суд,
HEB|9|28|так і Христос один раз був у жертву принесений, щоб понести гріхи багатьох, і не в справі гріха другий раз з'явитися тим, хто чекає Його на спасіння.
HEB|10|1|Бо Закон, мавши тільки тінь майбутнього добра, а не самий образ речей, тими самими жертвами, що завжди щороку приносяться, не може ніколи вдосконалити тих, хто приступає.
HEB|10|2|Інакше вони перестали б приноситись, бо ті, хто служить, очищені раз, уже б не мали жадної свідомости гріхів.
HEB|10|3|Але в них спомин про гріхи буває щороку,
HEB|10|4|бо тож неможливе, щоб кров биків та козлів здіймала гріхи!
HEB|10|5|Тому то, входячи в світ, Він говорить: Жертви й приношення Ти не схотів, але тіло Мені приготував.
HEB|10|6|Цілопалення й жертви покутної Ти не жадав.
HEB|10|7|Тоді Я сказав: Ось іду, в звої книжки про Мене написано, щоб волю чинити Твою, Боже!
HEB|10|8|Він вище сказав, що жертви й приносу, та цілопалення й жертви покутної, які за Законом приносяться, Ти не жадав і Собі не вподобав.
HEB|10|9|Потому сказав: Ось іду, щоб волю Твою чинити, Боже. Відміняє Він перше, щоб друге поставити.
HEB|10|10|У цій волі ми освячені жертвоприношенням тіла Ісуса Христа один раз.
HEB|10|11|І кожен священик щоденно стоїть, служачи, і часто приносить жертви ті самі, що ніколи не можуть зняти гріхів.
HEB|10|12|А Він за гріхи світу приніс жертву один раз, і назавжди по Божій правиці засів,
HEB|10|13|далі чекаючи, аж вороги Його будуть покладені за підніжка Його ніг.
HEB|10|14|Бо жертвоприношенням одним вдосконалив Він тих, хто освячується.
HEB|10|15|Свідкує ж і Дух Святий нам, як говорить:
HEB|10|16|Оце заповіт, що його по цих днях встановляю Я з ними, говорить Господь, Закони вої Я дам в їхні серця, і в їхніх думках напишу їх.
HEB|10|17|А їхніх гріхів та несправедливостей їхніх Я більш не згадаю!
HEB|10|18|А де їхнє відпущення, там нема вже жертвоприношення за гріхи.
HEB|10|19|Отож, браття, ми маємо відвагу входити до святині кров'ю Ісусовою,
HEB|10|20|новою й живою дорогою, яку нам обновив Він через завісу, цебто через тіло Своє,
HEB|10|21|маємо й Великого Священика над домом Божим,
HEB|10|22|то приступімо з щирим серцем, у повноті віри, окропивши серця від сумління лукавого та обмивши тіла чистою водою!
HEB|10|23|Тримаймо непохитне визнання надії, вірний бо Той, Хто обіцяв.
HEB|10|24|І уважаймо один за одним для заохоти до любови й до добрих учинків.
HEB|10|25|Не кидаймо збору свого, як то звичай у деяких, але заохочуймося, і тим більше, скільки більше ви бачите, що зближається день той.
HEB|10|26|Бо як ми грішимо самовільно, одержавши пізнання правди, то вже за гріхи не знаходиться жертви,
HEB|10|27|а страшливе якесь сподівання суду та гнів палючий, що має пожерти противників.
HEB|10|28|Хто відкидає Закона Мойсея, такий немилосердно вмирає при двох чи трьох свідках,
HEB|10|29|скільки ж більшої муки, додумуєтеся? заслуговує той, хто потоптав Сина Божого, і хто кров заповіту, що нею освячений, за звичайну вважав, і хто Духа благодаті зневажив!
HEB|10|30|Бо знаємо Того, Хто сказав: Мені помста належить, Я відплачу, говорить Господь. І ще: Господь буде судити народа Свого!
HEB|10|31|Страшна річ упасти в руки Бога Живого!
HEB|10|32|Згадайте ж про перші дні ваші, як ви просвітилися й витерпіли запеклу боротьбу страждань.
HEB|10|33|Ви були то видовищем зневаги й знущання, то були учасниками тих, що жили так.
HEB|10|34|Ви бо страждали й з ув'язненими, і грабунок свого майна прийняли з потіхою, відаючи, що маєте в небі для себе майно неминуще та краще.
HEB|10|35|Тож не відкидайте відваги своєї, бо має велику нагороду вона.
HEB|10|36|Бо вам терпеливість потрібна, щоб Божу волю вчинити й прийняти обітницю.
HEB|10|37|Бо ще мало, дуже мало, і Той, хто має прийти, прийде й баритись не буде!
HEB|10|38|А праведний житиме вірою. І: Коли захитається він, то душа Моя його не вподобає.
HEB|10|39|Ми ж не з тих, хто хитається на загибіль, але віруємо на спасіння душі.
HEB|11|1|А віра то підстава сподіваного, доказ небаченого.
HEB|11|2|Бо нею засвідчені старші були.
HEB|11|3|Вірою ми розуміємо, що віки Словом Божим збудовані, так що з невидимого сталось видиме.
HEB|11|4|Вірою Авель приніс Богові жертву кращу, як Каїн; нею засвідчений був, що він праведний, як Бог свідчив про дари його; нею, і вмерши, він ще промовляє.
HEB|11|5|Вірою Енох був перенесений на небо, щоб не бачити смерти; і його не знайшли, бо Бог переніс його. Бо раніш, як його перенесено, він був засвідчений, що Богові він догодив.
HEB|11|6|Догодити ж без віри не можна. І той, хто до Бога приходить, мусить вірувати, що Він є, а тим, хто шукає Його, Він дає нагороду.
HEB|11|7|Вірою Ной, як дістав був об'явлення про те, чого ще не бачив, побоявшись, зробив ковчега, щоб дім свій спасти; нею світ засудив він, і став спадкоємцем праведности, що з віри вона.
HEB|11|8|Вірою Авраам, покликаний на місце, яке мав прийняти в спадщину, послухався та й пішов, не відаючи, куди йде.
HEB|11|9|Вірою він перебував на Землі Обіцяній, як на чужій, і проживав у наметах з Ісаком та Яковом, співспадкоємцями тієї ж обітниці,
HEB|11|10|бо чекав він міста, що має підвалини, що Бог його будівничий та творець.
HEB|11|11|Вірою й Сара сама дістала силу прийняти насіння, і породила понад час свого віку, бо вірним вважала Того, Хто обітницю дав.
HEB|11|12|Тому й від одного, та ще змертвілого, народилось так багато, як зорі небесні й пісок незчисленний край моря.
HEB|11|13|Усі вони повмирали за вірою, не одержавши обітниць, але здалека бачили їх, і повітали, і вірували в них, та визнавали, що вони на землі чужаниці й приходьки.
HEB|11|14|Бо ті, що говорять таке, виявляють, що шукають батьківщини.
HEB|11|15|І коли б вони пам'ятали ту, що вийшли з неї, то мали б були час повернутись.
HEB|11|16|Та бажають вони тепер кращої, цебто небесної, тому й Бог не соромиться їх, щоб звати Себе їхнім Богом, бо Він приготував їм місто.
HEB|11|17|Вірою Авраам, випробовуваний, привів був на жертву Ісака, і, мавши обітницю, приніс однородженого,
HEB|11|18|що йому було сказано: В Ісакові буде насіння тобі.
HEB|11|19|Бо він розумів, що Бог має силу й воскресити з мертвих, тому й одержав його на прообраз.
HEB|11|20|Вірою в майбутнє поблагословив Ісак Якова та Ісава.
HEB|11|21|Вірою Яків, умираючи, поблагословив кожного сина Йосипового, і схилився на верх свого жезла.
HEB|11|22|Вірою Йосип, умираючи, згадав про вихід синів Ізраїлевих та про кості свої заповів.
HEB|11|23|Вірою Мойсей, як родився, переховувався батьками своїми три місяці, бо вони бачили, що гарне дитя, і не злякались наказу царевого.
HEB|11|24|Вірою Мойсей, коли виріс, відрікся зватися сином дочки фараонової.
HEB|11|25|Він хотів краще страждати з народом Божим, аніж мати дочасну гріховну потіху.
HEB|11|26|Він наругу Христову вважав за більше багатство, ніж скарби єгипетські, бо він озирався на Божу нагороду.
HEB|11|27|Вірою він покинув Єгипет, не злякавшися гніву царевого, бо він був непохитний, як той, хто Невидимого бачить.
HEB|11|28|Вірою справив він Пасху й покроплення крови, щоб їх не торкнувся той, хто погубив первороджених.
HEB|11|29|Вірою вони перейшли Червоне море, немов суходолом, на що спокусившись єгиптяни, потопились.
HEB|11|30|Вірою впали єрихонські мури по семиденнім обходженні їх.
HEB|11|31|Вірою блудниця Рахав не згинула з невірними, коли з миром прийняла вивідувачів.
HEB|11|32|І що ще скажу? Бо не стане часу мені, щоб оповідати про Гедеона, Варака, Самсона, Ефтая, Давида й Самуїла та про пророків,
HEB|11|33|що вірою царства побивали, правду чинили, одержували обітниці, пащі левам загороджували,
HEB|11|34|силу огненну гасили, утікали від вістря меча, зміцнялись від слабости, хоробрі були на війні, обертали в розтіч полки чужоземців;
HEB|11|35|жінки діставали померлих своїх із воскресіння; а інші бували скатовані, не прийнявши визволення, щоб отримати краще воскресіння;
HEB|11|36|а інші дізнали наруги та рани, а також кайдани й в'язниці.
HEB|11|37|Камінням побиті бували, допитувані, перепилювані, умирали, зарубані мечем, тинялися в овечих та козячих шкурах, збідовані, засумовані, витерпілі.
HEB|11|38|Ті, що світ не вартий був їх, тинялися по пустинях та горах, і по печерах та проваллях земних.
HEB|11|39|І всі вони, одержавши засвідчення вірою, обітниці не прийняли,
HEB|11|40|бо Бог передбачив щось краще про нас, щоб вони не без нас досконалість одержали.
HEB|12|1|Тож і ми, мавши навколо себе велику таку хмару свідків, скиньмо всякий тягар та гріх, що обплутує нас, та й біжім з терпеливістю до боротьби, яка перед нами,
HEB|12|2|дивлячись на Ісуса, на Начальника й Виконавця віри, що замість радости, яка була перед Ним, перетерпів хреста, не звертавши уваги на сором, і сів по правиці престолу Божого.
HEB|12|3|Тож подумайте про Того, хто перетерпів такий перекір проти Себе від грішних, щоб ви не знемоглись, і не впали на душах своїх.
HEB|12|4|Ви ще не змагались до крови, борючись проти гріха,
HEB|12|5|і забули нагад, що говорить до вас, як синів: Мій сину, не нехтуй Господньої кари, і не знемагай, коли Він докоряє тобі.
HEB|12|6|Бо Господь, кого любить, того Він карає, і б'є кожного сина, якого приймає!
HEB|12|7|Коли терпите кару, то робить Бог вам, як синам. Хіба є такий син, що батько його не карає?
HEB|12|8|А коли ви без кари, що спільна для всіх, то ви діти з перелюбу, а не сини.
HEB|12|9|А до того, ми мали батьків, що карали наше тіло, і боялися їх, то чи ж не далеко більше повинні коритися ми Отцеві духів, щоб жити?
HEB|12|10|Ті нас за короткого часу карали, як їм до вподоби було, Цей же на користь, щоб ми стали учасниками Його святости.
HEB|12|11|Усяка кара в теперішній час не здається потіхою, але смутком, та згодом для навчених нею приносить мирний плід праведности!
HEB|12|12|Тому то опущені руки й коліна знеможені випростуйте,
HEB|12|13|і чиніть прості стежки ногам вашим, щоб кульгаве не збочило, але краще виправилось.
HEB|12|14|Пильнуйте про мир зо всіма, і про святість, без якої ніхто не побачить Господа.
HEB|12|15|Дивіться, щоб хто не зостався без Божої благодаті, щоб не виріс який гіркий корінь і не наробив непокою, і щоб багато-хто не опоганились тим.
HEB|12|16|Щоб не був хто блудник чи безбожник, немов той Ісав, що своє перворідство віддав за поживу саму.
HEB|12|17|Бо знаєте ви, що й після, як схотів він успадкувати благословення, відкинутий був, не знайшов бо був можливости до покаяння, хоч його із слізьми шукав.
HEB|12|18|Бо ви не приступили до гори дотикальної та до палючого огню, і до хмари, і до темряви, та до бурі,
HEB|12|19|і до сурмового звуку, і до голосу слів, що його ті, хто чув, просили, щоб більше не мовилось слово до них.
HEB|12|20|Не могли бо вони того витримати, що наказано: Коли й звірина до гори доторкнеться, то буде камінням побита.
HEB|12|21|І таке страшне те видіння було, що Мойсей проказав: Я боюся й тремчу!...
HEB|12|22|Але ви приступили до гори Сіонської, і до міста Бога Живого, до Єрусалиму небесного, і до десятків тисяч Анголів,
HEB|12|23|і до Церкви первороджених, на небі написаних, і до Судді всіх до Бога, і до духів удосконалених праведників,
HEB|12|24|і до Посередника Нового Заповіту до Ісуса, і до покроплення крови, що краще промовляє, як Авелева.
HEB|12|25|Глядіть, не відвертайтеся від того, хто промовляє. Бо як не повтікали вони, що зреклися того, хто звіщав на землі, то тим більше ми, якщо зрікаємся Того, Хто з неба звіщає,
HEB|12|26|що голос Його захитав тоді землю, а тепер обіцяв та каже: Ще раз захитаю не тільки землею, але й небом.
HEB|12|27|А ще раз визначає заміну захитаного, як створеного, щоб зосталися ті, хто непохитний.
HEB|12|28|Отож ми, що приймаємо царство непохитне, нехай маємо благодать, що нею приємно служитимемо Богові з побожністю й зо страхом.
HEB|12|29|Бо наш Бог то палючий огонь!
HEB|13|1|Братолюбство нехай пробуває між вами!
HEB|13|2|Не забувайте любови до приходнів, бо деякі нею, навіть не відаючи, гостинно були прийняли Анголів.
HEB|13|3|Пам'ятайте про в'язнів, немов із ними були б ви пов'язані, про тих, хто страждає, як такі, що й самі ви знаходитесь в тілі.
HEB|13|4|Нехай буде в усіх чесний шлюб та ложе непорочне, а блудників та перелюбів судитиме Бог.
HEB|13|5|Будьте життям не грошолюбні, задовольняйтеся тим, що маєте. Сам бо сказав: Я тебе не покину, ані не відступлюся від тебе!
HEB|13|6|Тому то ми сміливо говоримо: Господь мені помічник, і я не злякаюсь нікого: що зробить людина мені?
HEB|13|7|Спогадуйте наставників ваших, що вам говорили Слово Боже; і, дивлячися на кінець їхнього життя, переймайте їхню віру.
HEB|13|8|Ісус Христос учора, і сьогодні, і навіки Той Самий!
HEB|13|9|Не захоплюйтеся всілякими та чужими науками. Бо річ добра зміцняти серця благодаттю, а не стравами, що користи від них не одержали ті, хто за ними ходив.
HEB|13|10|Маємо жертівника, що від нього годуватися права не мають ті, хто скинії служить,
HEB|13|11|бо котрих звірят кров первосвященик уносить до святині за гріхи, тих м'ясо палиться поза табором,
HEB|13|12|тому то Ісус, щоб кров'ю Своєю людей освятити, постраждав поза брамою.
HEB|13|13|Тож виходьмо до Нього поза табір, і наругу Його понесімо,
HEB|13|14|бо постійного міста не маємо тут, а шукаємо майбутнього!
HEB|13|15|Отож, завжди приносьмо Богові жертву хвали, цебто плід уст, що Ім'я Його славлять.
HEB|13|16|Не забувайте ж і про доброчинність та спільність, бо жертви такі вгодні Богові.
HEB|13|17|Слухайтесь ваших наставників та коріться їм, вони бо пильнують душ ваших, як ті, хто має здати справу. Нехай вони роблять це з радістю, а не зідхаючи, бо це для вас не корисне.
HEB|13|18|Моліться за нас, бо надіємося, що ми маємо добре сумління, бо хочемо добре в усьому поводитись.
HEB|13|19|А надто прошу це робити, щоб швидше до вас мене вернено.
HEB|13|20|Бог же миру, що з мертвих підняв великого Пастиря вівцям кров'ю вічного заповіту, Господа нашого Ісуса,
HEB|13|21|нехай вас удосконалить у кожному доброму ділі, щоб волю чинити Його, чинячи в вас любе перед лицем Його через Ісуса Христа, Якому слава на віки вічні. Амінь.
HEB|13|22|Благаю ж вас, браття, прийміть слово потіхи, бо коротко я написав вам.
HEB|13|23|Знайте, що наш брат Тимофій вже випущений, і я з ним; коли незабаром він прийде, я вас побачу.
HEB|13|24|Вітайте всіх ваших наставників та всіх святих. Вітають вас ті, хто в Італії.
HEB|13|25|Благодать зо всіма вами! Амінь.
