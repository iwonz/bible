MAL|1|1|耶和华的话，藉 玛拉基 传给 以色列 的默示。
MAL|1|2|耶和华说：“我曾爱你们。”你们却说：“你在何事上爱我们呢？”耶和华说：“ 以扫 不是 雅各 的哥哥吗？我却爱 雅各 ，
MAL|1|3|恶 以扫 ，使他的山岭荒凉，把他的地业交给旷野的野狗。”
MAL|1|4|以东 若说：“我们虽被毁坏，却要重建荒废之处。”万军之耶和华如此说：“任他们建造，我必拆毁；人必称他们为‘邪恶之境’，为‘耶和华永远恼怒之民’。”
MAL|1|5|你们必亲眼看见，你们要说：“耶和华在 以色列 疆界之外必尊为大！”
MAL|1|6|万军之耶和华对你们说：“儿子孝敬父亲，仆人敬畏主人；我既为父亲，孝敬我的在哪里呢？我既为主人，敬畏我的在哪里呢？你们这些藐视我名的祭司啊！”你们却说：“我们在何事上藐视你的名呢？”
MAL|1|7|“你们将不洁净的食物献在我的祭坛上，却说：‘我们在何事上使你不洁净呢？’你们说，耶和华的供桌是可藐视的。
MAL|1|8|你们将瞎眼的献为祭物，这不算为恶吗？将瘸腿的、有病的献上，这不算为恶吗？那么，请把这些献给你的省长，他岂会悦纳你 ，岂会抬举你呢？这是万军之耶和华说的。”
MAL|1|9|现在我劝你们要恳求上帝，好让他施恩给我们。这事既出于你们的手，他岂会抬举你们任何人呢？这是万军之耶和华说的。
MAL|1|10|万军之耶和华说：“甚愿你们中间有人把殿的门 关上，免得你们徒然在我坛上烧火。我不喜欢你们，也不从你们手中悦纳供物。”
MAL|1|11|万军之耶和华说：“从日出之地到日落之处，我的名在列国中必尊为大。在各处，人必奉我的名烧香，献洁净的供物，因为我的名在列国中必尊为大。
MAL|1|12|你们却亵渎我的名，说：‘主的供桌是不洁净的，供桌上的果子和食物是可藐视的。’
MAL|1|13|你们又说：‘看哪，这些事何等烦琐！’并嗤之以鼻 。这是万军之耶和华说的。你们把抢来的、瘸腿的、有病的拿来献上为祭，我岂能从你们手中悦纳它呢？这是耶和华说的。
MAL|1|14|行诡诈的人是可诅咒的！他的群畜中虽有公羊，他许了愿，却将有残疾的献给主。因我是大君王，我的名在列国中是可畏的。这是万军之耶和华说的。”
MAL|2|1|现在，众祭司啊，这诫命是给你们的。
MAL|2|2|万军之耶和华说：“你们若不听，不放在心上，不将荣耀归给我的名，我就使诅咒临到你们，使你们的福分变为诅咒；其实我已经诅咒了你们的福分，因你们不把诫命放在心上。
MAL|2|3|看哪，我要斥责你们的后裔，把粪抹在你们脸上，就是你们祭牲 的粪。人要把你们和粪一起抬出去，
MAL|2|4|你们就知道我颁这诫命给你们，使我与 利未 所立的约可以常存。这是万军之耶和华说的。
MAL|2|5|我曾与他立生命和平安的约。我将这两样赐给他，使他存敬畏的心；他就敬畏我，惧怕我的名。
MAL|2|6|真实的训诲在他口中，他的嘴唇中没有不义。他以平安和正直与我同行，使许多人回转离开罪孽。
MAL|2|7|祭司的嘴唇当守护知识，人也当从他口中寻求训诲，因为他是万军之耶和华的使者。
MAL|2|8|你们却偏离正道，使许多人在这训诲上绊跌。你们破坏了我与 利未 人所立的约。这是万军之耶和华说的。
MAL|2|9|所以我使你们被众百姓藐视，看为卑贱；因你们不遵守我的道，在律法上看人的情面 。”
MAL|2|10|我们岂不都有一位父吗？岂不是一位上帝创造了我们吗？为何互相行诡诈，亵渎了上帝与我们列祖所立的约呢？
MAL|2|11|犹大 行事诡诈，在 以色列 和 耶路撒冷 中行了可憎的事；因为 犹大 人亵渎耶和华所喜爱的圣殿，娶外邦神明的女子为妻。
MAL|2|12|凡做这事的，无论是清醒的 或回应的，即使献供物给万军之耶和华，耶和华也要将他从 雅各 的帐棚中剪除。
MAL|2|13|你们又再做这样的事，使哭泣和叹息的眼泪遮盖耶和华的祭坛，以致耶和华不再理会那供物，也不喜欢从你们的手中收纳。
MAL|2|14|你们还说：“这是为什么呢？”因为耶和华在你和你年轻时所娶的妻之间作证。她虽是你的配偶，你誓约 的妻，你却背弃她。
MAL|2|15|一个人如果还剩下一点灵性，他不会这么做。这人在寻找什么呢？上帝的后裔！ 当谨守你们的灵性，谁也不可背弃年轻时所娶的妻。
MAL|2|16|耶和华－ 以色列 的上帝说：“我恨恶休妻的事和衣服外面披上暴力的人。所以当谨守你们的心，不可行诡诈。这是万军之耶和华说的。”
MAL|2|17|你们用言语使耶和华厌烦，却说：“我们在何事上使他厌烦呢？”因为你们说：“凡行恶的，耶和华看为善，并且喜爱他们；”又说：“公平的上帝在哪里呢？”
MAL|3|1|万军之耶和华说：“看哪，我要差遣我的使者在我前面预备道路。你们所寻求的主必忽然来到他的殿；立约的使者，就是你们所仰慕的，看哪，快要来到。”
MAL|3|2|他来的日子，谁能当得起呢？他显现的时候，谁能立得住呢？因为他如炼金匠的火，如漂洗者的碱。
MAL|3|3|他必坐下如炼净银子的人，必洁净 利未 人，熬炼他们像金银一样；他们就凭公义献供物给耶和华。
MAL|3|4|那时， 犹大 和 耶路撒冷 所献的供物必蒙耶和华悦纳，仿佛古时之日、上古之年。
MAL|3|5|万军之耶和华说：“我必临近你们，施行审判。我必速速作见证，警戒那些行邪术的、犯奸淫的、起假誓的、剥削雇工工钱的、欺压孤儿寡妇的、屈枉寄居者的和不敬畏我的人。”
MAL|3|6|“我－耶和华是不改变的；所以， 雅各 的子孙啊，你们不致灭亡。
MAL|3|7|从你们祖先的日子以来，你们就偏离我的律例而不遵守。现在你们要转向我，我就转向你们。这是万军之耶和华说的。你们却说：‘我们如何转向呢？’
MAL|3|8|人岂可抢夺上帝呢？你们竟抢夺我！你们却说：‘我们在何事上抢夺你呢？’其实就是在你们当纳的十分之一奉献和当献的供物上。
MAL|3|9|因你们全国上下都抢夺我的供物，诅咒就临到你们身上。
MAL|3|10|你们要将当纳的十分之一全然送入仓库，使我家有粮，以此试试我，是否为你们敞开天上的窗户，倾福与你们，甚至无处可容。这是万军之耶和华说的。
MAL|3|11|我必为你们斥责蝗虫 ，不容它毁坏你们的土产。你们田间的葡萄树，果实未熟以先也不会掉落。这是万军之耶和华说的。
MAL|3|12|万国必称你们为有福的，因你们必成为喜乐之地。这是万军之耶和华说的。”
MAL|3|13|耶和华说：“你们用话顶撞我。”你们却说：“我们说了什么话顶撞你呢？”
MAL|3|14|你们说：“事奉上帝是枉然，我们遵守上帝所吩咐的，在万军之耶和华面前哀痛而行，有什么益处呢？
MAL|3|15|现在，我们称狂傲的人为有福，并且行恶的人得以建立；他们虽然试探上帝，却得以逃脱。”
MAL|3|16|那时，敬畏耶和华的人彼此谈论，耶和华侧耳而听，且有纪念册在他面前，记录那敬畏耶和华、思念他名的人。
MAL|3|17|万军之耶和华说：“在我所定的日子，他们必属我，是我宝贵的产业。我必怜悯他们，如同人怜悯那服侍他的儿子。
MAL|3|18|那时你们必再一次 看出义人和恶人，事奉上帝和不事奉上帝的人有何差别。”
MAL|4|1|万军之耶和华说：“看哪，那日临近，势如烧着的火炉，凡狂傲的和行恶的都如碎秸，在那日被烧尽，根与枝条无一存留。
MAL|4|2|但是，对你们敬畏我名的人，必有公义的太阳出现，其光线 有医治的能力。你们必出来跳跃如圈里的牛犊。
MAL|4|3|你们必践踏恶人；在我所定的日子，他们必成为你们脚掌下的灰尘。这是万军之耶和华说的。
MAL|4|4|“你们当记念我仆人 摩西 的律法，就是我在 何烈山 为 以色列 众人所吩咐他的律例典章。
MAL|4|5|“看哪，耶和华大而可畏之日未到以前，我要差遣 以利亚 先知到你们那里去。
MAL|4|6|他必使父亲的心转向儿女，儿女的心转向父亲，免得我来诅咒这地。”
