2COR|1|1|Павло, з волі Божої апостол Христа Ісуса, та брат Тимофій, до Божої Церкви в Коринті, з усіма святими в цілій Ахаї,
2COR|1|2|благодать вам і мир від Бога Отця нашого й Господа Ісуса Христа!
2COR|1|3|Благословенний Бог і Отець Господа нашого Ісуса Христа, Отець милосердя й Бог потіхи всілякої,
2COR|1|4|що в усякій скорботі Він нас потішає, щоб змогли потішати й ми тих, що в усякій скорботі знаходяться, тією потіхою, якою потішує Бог нас самих.
2COR|1|5|Бо поскільки намножуються в нас терпіння Христові, так через Христа й потішення наше намножується.
2COR|1|6|Бо як терпимо скорботи, то на вашу потіху й спасіння; коли потішаємось, то на вашу потіху в терпінні тих самих страждань, які терпимо й ми.
2COR|1|7|А наша надія певна про вас, бо ми знаємо, що ви спільники як у терпіннях, так само і в потісі.
2COR|1|8|Бо не хочемо, браття, щоб не відали ви про нашу скорботу, що в Азії трапилась нам, бо над міру й над силу були ми обтяжені, так що ми не надіялися навіть жити.
2COR|1|9|Та самі ми в собі мали присуд на смерть, щоб нам не покладати надії на себе, а на Бога, що воскрешує мертвих,
2COR|1|10|що від смерти такої нас визволив і визволяє, і на Нього й покладаємося, що й ще визволить Він,
2COR|1|11|як поможете разом і ви молитвою за нас, щоб за дар ласки, що нам виявлений багатьма, багато-хто дяку складали за нас.
2COR|1|12|Бо це нам хвала, свідчення нашого сумління, що в святості й чистості Божій, не в тілесній мудрості, але в Божій благодаті жили ми на світі, особливо ж у вас.
2COR|1|13|Бо іншого вам ми не пишемо, тільки те, що читаєте та розумієте, а сподіваюсь, що ви й до кінця зрозумієте,
2COR|1|14|як частинно нас ви й зрозуміли, що ми вам похвала, як і ви нам, у день Господа нашого Ісуса.
2COR|1|15|І з певністю цією хотів я давніше прибути до вас, щоб мали ви благодать удруге,
2COR|1|16|і через вас перейти в Македонію, а з Македонії знову прибути до вас, а ви щоб в Юдею мене відпровадили.
2COR|1|17|Маючи задум такий, чи я чинив легковажно? Чи те, що задумую, за тілом задумую, щоб було в мене і Так, так, і Ні, ні?
2COR|1|18|Але вірний Бог, що наше слово до вас не було Так і Ні.
2COR|1|19|Бо Син Божий Ісус Христос, що ми Його вам проповідували, я й Силуан, і Тимофій, не був Так і Ні, але в Нім було Так.
2COR|1|20|Скільки бо Божих обітниць, то в Ньому Так, і в Ньому Амінь, Богові на славу через нас.
2COR|1|21|А Той, Хто нас із вами в Христа утверджує, і Хто нас намастив, то Бог,
2COR|1|22|Який і назнаменував нас, і в наші серця дав завдаток Духа.
2COR|1|23|А я кличу Бога на свідка на душу мою, що я, щадячи вас, не прийшов у Коринт дотепер,
2COR|1|24|не тому, ніби ми беремо владу над вашою вірою, але вашої радости помічники ми, бо ви встояли вірою!
2COR|2|1|А я постановив у собі те, щоб до вас не прийти знов у смутку.
2COR|2|2|Бо коли я засмучую вас, то хто той, хто потішить мене, як не той, кого я засмутив?
2COR|2|3|І це саме писав я до вас, щоб, прийшовши, я смутку не мав би від тих, що від них мені тішитися належало, про всіх вас бувши певний, що радість моя то радість усіх вас!
2COR|2|4|Бо з великого горя та з туги сердечної я написав вам з рясними слізьми не на те, щоб були ви засмучені, але щоб пізнали любов, що в мене її пребагато до вас!
2COR|2|5|А як хто засмутив, не мене засмутив, а почасти щоб не пригнітити і всіх вас.
2COR|2|6|Досить такому карання того, що від багатьох,
2COR|2|7|через те навпаки, краще простити й потішити, щоб смуток великий його не пожер.
2COR|2|8|Через те вас благаю: зміцніть до нього любов!
2COR|2|9|Бо на це я й писав, щоб пізнати ваш досвід, чи в усім ви слухняні.
2COR|2|10|А кому ви прощаєте що, тому й я; бо й я, як простив що кому, то кому я простив, зробив те через вас від Особи Христа,
2COR|2|11|щоб нас сатана не перехитрував, відомі бо нам його задуми!
2COR|2|12|А коли я прийшов до Троади звіщати Христову Євангелію, і були двері для мене відчинені в Господі,
2COR|2|13|не мав я спокою для духа свого, бо я не знайшов був свого брата Тита; але, попрощавшися з ними, я пішов в Македонію.
2COR|2|14|А Богові подяка, що Він постійно чинить нас переможцями в Христі, і запашність знання про Себе через нас виявляє на всякому місці!
2COR|2|15|Ми бо для Бога Христова запашність серед тих, хто спасається, і тих, які гинуть,
2COR|2|16|для одних бо смертельна запашність на смерть, а для других запашність життєва в життя. І хто здатен на це?
2COR|2|17|Бо ми не такі, як багато-хто, що Боже Слово фальшують, але ми провіщаємо, як із щирости, як від Бога, перед Богом, у Христі!
2COR|3|1|Чи нам знов зачинати доручувати самих себе? Чи ми потребуємо, як дехто, листів доручальних до вас чи від вас?
2COR|3|2|Ви наш лист, написаний у наших серцях, якого всі люди знають і читають!
2COR|3|3|Виявляєте ви, що ви лист Христів, нами вислужений, що написаний не чорнилом, але Духом Бога Живого, не на таблицях камінних, але на тілесних таблицях серця.
2COR|3|4|Таку ж певність до Бога ми маємо через Христа,
2COR|3|5|не тому, що ми здібні помислити щось із себе, як від себе, але наша здібність від Бога.
2COR|3|6|І Він нас зробив бути здатними служителями Нового Заповіту, не букви, а духа, бо буква вбиває, а дух оживляє.
2COR|3|7|Коли ж служіння смерті, вирізане на каменях буквами, було таке славне, що Ізраїлеві сини не могли дивитись на обличчя Мойсея, через славу минущу обличчя його,
2COR|3|8|скільки ж більш буде в славі те служіння духа!
2COR|3|9|Бо як служіння осуду слава, то служіння праведности тим більше багате на славу!
2COR|3|10|Не прославилося бо прославлене, у цій частині, ради слави, що вона переважує,
2COR|3|11|бо коли славне те, що минає, то багато більш у славі те, що триває!
2COR|3|12|Тож, мавши надію таку, ми вживаємо великої сміливости,
2COR|3|13|а не як Мойсей, що покривало клав на обличчя своє, щоб Ізраїлеві сини не дивилися на кінець того, що минає.
2COR|3|14|Але засліпилися їхні думки, бо те саме покривало аж до сьогодні лишилось незняте в читанні Старого Заповіту, бо зникає воно Христом.
2COR|3|15|Але аж до сьогодні, як читають Мойсея, на їхньому серці лежить покривало,
2COR|3|16|коли ж вони навернуться до Господа, тоді покривало здіймається.
2COR|3|17|Господь же то Дух, а де Дух Господній, там воля.
2COR|3|18|Ми ж відкритим обличчям, як у дзеркало, дивимося всі на славу Господню, і зміняємося в той же образ від слави на славу, як від Духа Господнього.
2COR|4|1|Ось тому, мавши за милосердям Божим таке служіння, ми не тратимо відваги,
2COR|4|2|але ми відреклися тайного сорому, не ходячи в хитрості та не перекручуючи Божого Слова, але з'явленням правди доручуємо себе кожному сумлінню людському перед Богом.
2COR|4|3|Коли ж наша Євангелія й закрита, то закрита для тих, хто гине,
2COR|4|4|для невіруючих, яким бог цього віку засліпив розум, щоб для них не засяяло світло Євангелії слави Христа, а Він образ Божий.
2COR|4|5|Бо ми не себе самих проповідуємо, але Христа Ісуса, Господа, ми ж самі раби ваші ради Ісуса.
2COR|4|6|Бо Бог, що звелів був світлу засяяти з темряви, у серцях наших засяяв, щоб просвітити нам знання слави Божої в Особі Христовій.
2COR|4|7|А ми маємо скарб цей у посудинах глиняних, щоб велич сили була Божа, а не від нас.
2COR|4|8|У всьому нас тиснуть, та не потиснені ми; ми в важких обставинах, але не впадаємо в розпач.
2COR|4|9|Переслідують нас, але ми не полишені; ми повалені, та не погублені.
2COR|4|10|Ми завсіди носимо в тілі мертвість Ісусову, щоб з'явилося в нашому тілі й життя Ісусове.
2COR|4|11|Бо завсіди нас, що живемо, віддають на смерть за Ісуса, щоб з'явилось Ісусове в нашому смертельному тілі.
2COR|4|12|Тому то смерть діє в нас, а життя у вас.
2COR|4|13|Та мавши того ж духа віри, за написаним: Вірував я, через те говорив, і ми віруємо, тому то й говоримо,
2COR|4|14|знавши, що Той, Хто воскресив Господа Ісуса, воскресить з Ісусом і нас, і поставить із вами.
2COR|4|15|Усе бо для вас, щоб благодать, розмножена через багатьох, збагатила подяку на Божу славу.
2COR|4|16|Через те ми відваги не тратимо, бо хоч нищиться зовнішній наш чоловік, зате день-у-день відновляється внутрішній.
2COR|4|17|Бо теперішнє легке наше горе достачає для нас у безмірнім багатстві славу вічної ваги,
2COR|4|18|коли ми не дивимося на видиме, а на невидиме. Бо видиме дочасне, невидиме ж вічне!
2COR|5|1|Знаємо бо, коли земний мешкальний намет наш зруйнується, то маємо будівлю від Бога на небі, дім нерукотворний та вічний.
2COR|5|2|Тому то й зідхаємо, бажаючи приодягтися будівлею нашею, що з неба,
2COR|5|3|коли б тільки й одягнені ми не знайшлися нагі!
2COR|5|4|Бо ми, знаходячися в цьому наметі, зідхаємо під тягарем, бо не хочемо роздягтися, але одягтися, щоб смертне пожерлось життям.
2COR|5|5|А Той, Хто на це саме й створив нас, то Бог, що й дав нам завдаток Духа.
2COR|5|6|Отож, бувши відважні постійно, та знаючи, що, мавши дім у тілі, ми не перебуваємо в домі Господньому,
2COR|5|7|бо ходимо вірою, а не видінням,
2COR|5|8|ми ж відважні, і бажаємо краще покинути дім тіла й мати дім у Господа.
2COR|5|9|Тому ми й пильнуємо, чи зостаємося в домі тіла, чи виходимо з дому, бути Йому любими.
2COR|5|10|Бо мусимо всі ми з'явитися перед судовим престолом Христовим, щоб кожен прийняв згідно з тим, що в тілі робив він, чи добре, чи лихе.
2COR|5|11|Отже, відаючи страх Господній, ми людей переконуємо, а Богові явні; але маю надію, що й у ваших сумліннях ми явні.
2COR|5|12|Бо не знову себе ми доручуємо вам, але даємо вам привід хвалитися нами, щоб мали ви що проти тих, що хваляться обличчям, а не серцем.
2COR|5|13|Коли бо ми з розуму сходимо, то Богові, коли ж при здоровому розумі, то для вас.
2COR|5|14|Бо Христова любов спонукує нас, що думають так, що коли вмер Один за всіх, то всі померли.
2COR|5|15|А вмер Він за всіх, щоб ті, хто живе, не жили вже для себе самих, а для Того, Хто за них був умер і воскрес.
2COR|5|16|Через те відтепер ми нікого не знаємо за тілом; коли ж і знали за тілом Христа, то тепер ми не знаємо вже!
2COR|5|17|Тому то, коли хто в Христі, той створіння нове, стародавнє минуло, ото сталось нове!
2COR|5|18|Усе ж від Бога, що нас примирив із Собою Ісусом Христом і дав нам служіння примирення,
2COR|5|19|бо Бог у Христі примирив світ із Собою Самим, не зважавши на їхні провини, і поклав у нас слово примирення.
2COR|5|20|Оце ми як посли замість Христа, ніби Бог благає через нас, благаємо замість Христа: примиріться з Богом!
2COR|5|21|Бо Того, Хто не відав гріха, Він учинив за нас гріхом, щоб стали ми Божою правдою в Нім!
2COR|6|1|А ми, як співробітники, благаємо, щоб ви Божої благодаті не брали надармо.
2COR|6|2|Бо каже: Приємного часу почув Я тебе, і поміг Я тобі в день спасіння! Ось тепер час приємний, ось тепер день спасіння!
2COR|6|3|Ні в чому ніякого спотикання не робимо, щоб служіння було бездоганне,
2COR|6|4|а в усьому себе виявляємо, як служителів Божих, у великім терпінні, у скорботах, у бідах, у тіснотах,
2COR|6|5|у вдарах, у в'язницях, у розрухах, у працях, у недосипаннях, у постах,
2COR|6|6|у чистості, у розумі, у лагідності, у добрості, у Дусі Святім, у нелицемірній любові,
2COR|6|7|у слові істини, у силі Божій, зо зброєю правди в правиці й лівиці,
2COR|6|8|через славу й безчестя, через ганьбу й хвалу, як обманці, але ми правдиві;
2COR|6|9|як незнані, та познані, як умираючі, та ось ми живі; як карані, та не забиті;
2COR|6|10|як сумні, але завжди веселі; як убогі, але багатьох ми збагачуємо; як ті, що нічого не мають, але всім володіємо.
2COR|6|11|Уста наші відкрились до вас, коринтяни, серце наше розширене!
2COR|6|12|У нас вам не тісно, але тісно вам у ваших серцях!
2COR|6|13|Такою ж відплатою говорю, немов дітям розширені будьте й ви!
2COR|6|14|До чужого ярма не впрягайтесь з невірними; бо що спільного між праведністю та беззаконням, або яка спільність у світла з темрявою?
2COR|6|15|Яка згода в Христа з белійяаром? Або яка частка вірного з невірним?
2COR|6|16|Або яка згода поміж Божим храмом та ідолами? Бо ви храм Бога Живого, як Бог прорік: Поселюсь серед них і ходитиму, і буду їм Богом, а вони будуть народом Моїм!
2COR|6|17|Вийдіть тому з-поміж них та й відлучіться, каже Господь, і не торкайтесь нечистого, і Я вас прийму,
2COR|6|18|і буду Я вам за Отця, а ви за синів і дочок Мені будете, говорить Господь Вседержитель!
2COR|7|1|Отож, мої любі, мавши ці обітниці, очистьмо себе від усякої нечисти тіла та духа, і творімо святиню у Божім страху!
2COR|7|2|Дайте місце для нас! Ми нікого не скривдили, нікого не зіпсували, нікого не ошукали!
2COR|7|3|Говорю не на осуд, бо я перед тим був сказав, що ви в серцях наших, щоб нам із вами чи померти чи жити.
2COR|7|4|У мене велика сміливість до вас, велика мені похвала з вас, я повний потіхи, збагачаюся радістю при всякому нашому горі.
2COR|7|5|Бо коли ми прийшли в Македонію, тіло наше не мало спочинку ніякого, у всьому бідуючи: назовні бої, страхіття всередині.
2COR|7|6|Але Бог, що тішить принижених, потішив нас приходом Тита,
2COR|7|7|і не тільки його прибуттям, а й потішенням, що ним він потішився з вас, коли розповідав нам про вашу журбу, про ваш смуток, про вашу горливість до мене, так що я більше тішився.
2COR|7|8|Коли я й засмутив вас листом, то не каюся, хоч і каявся був, бо бачу, що той лист засмутив вас, хоч і часово.
2COR|7|9|Я радію тепер не тому, що ви засмутились, а що ви засмутилися на покаяння, бо ви засмутились для Бога, щоб ні в чому не мати втрати від нас.
2COR|7|10|Бо смуток для Бога чинить каяття на спасіння, а про нього не жалуємо, а смуток світський чинить смерть.
2COR|7|11|Бо ось саме це, що ви засмутились для Бога, яку пильність велику воно вам зробило, яку оборону, яке обурення, який страх, яке бажання, яку горливість, яку помсту! Ви в усім показали, що чисті ви в справі.
2COR|7|12|А коли я й писав вам, то не через того, хто кривдить, і не через покривдженого, а щоб виявилася для вас наша пильність про вас перед Богом.
2COR|7|13|Тому то потіхою вашою втішились ми, а ще більше зраділи ми радістю Тита, що ви всі заспокоїли духа його.
2COR|7|14|Бо коли я про вас йому чим похвалився, то не осоромився; але як ми вам говорили все правду, так і наша хвала перед Титом правдива була!
2COR|7|15|І серце його прихильніше до вас, коли згадує він про покору всіх вас, як його прийняли ви були зо страхом і тремтінням.
2COR|7|16|Отож, тішуся я, що можу покластись у всьому на вас!
2COR|8|1|Повідомляємо ж вас, браття, про Божу благодать, що дана Церквам македонським,
2COR|8|2|що серед великого досвіду горя вони мають радість рясну, і глибоке їхнє убозтво збагатилось багатством їхньої щирости;
2COR|8|3|бо вони добровільні в міру сил своїх, і над силу, засвідчую,
2COR|8|4|із ревним благанням вони нас просили, щоб ми прийняли дар та спільність служіння святим.
2COR|8|5|І не так, як надіялись ми, але віддали себе перш Господеві та нам із волі Божої,
2COR|8|6|щоб ми благали Тита, щоб він, як був перше зачав, так і скінчив би в вас оце добре діло.
2COR|8|7|А ви, як у всім, збагачуєтесь: вірою, і словом, і розумом, і всякою пильністю, і вашою любов'ю до нас, щоб збагачувались ви і в благодаті оцій.
2COR|8|8|Не кажу це, як наказа, але пильністю інших досвідчую щирість любови й вашої.
2COR|8|9|Бо ви знаєте благодать Господа нашого Ісуса Христа, Який, бувши багатий, збіднів ради вас, щоб ви збагатились Його убозтвом.
2COR|8|10|І раду даю вам про це, бо це вам на пожиток, що не тільки чинили, але перші ви стали й бажати з минулого року.
2COR|8|11|А тепер закінчіть роботу, щоб ви, як горливо бажали, так і виконали б у міру можности.
2COR|8|12|Бо коли є охота, то приємна вона згідно з тим, що хто має, а не з тим, чого хто не має.
2COR|8|13|Хай не буде для інших полегша, а тягар для вас, але рівність для всіх.
2COR|8|14|Часу теперішнього ваш достаток нехай нестаткові їхньому допоможе, щоб і їхній достаток був на ваш нестаток, щоб рівність була,
2COR|8|15|як написано: Хто мав багато, той не мав зайвини, а хто мало, не мав недостачі.
2COR|8|16|Та Богові дяка, що Він таку пильність про вас дав у Титове серце,
2COR|8|17|бо благання прийняв він, але, бувши горливий, удався до вас добровільно.
2COR|8|18|А з ним разом послали ми брата, якого по всіх Церквах хвалять за Євангелію,
2COR|8|19|і не тільки оце, але вибраний був від Церков бути товаришем нашим у дорозі для благодаті тієї, якій служимо ми на хвалу Самого Господа,
2COR|8|20|остерігаючись того, щоб хто не дорікав нам цим достатком, що ним служимо ми,
2COR|8|21|дбаючи про добро не тільки перед Богом, але й перед людьми.
2COR|8|22|А ми з ними послали були брата нашого, про пильність якого ми часто досвідчувались у речах багатьох, який ще пильніший тепер через велике довір'я до вас.
2COR|8|23|Щодо Тита, то він мій товариш, а ваш співробітник; щождо наших братів вони посланці від Церков, вони слава Христова!
2COR|8|24|Отож, дайте їм доказа своєї любови й нашого хваління вас перед Церквами!
2COR|9|1|А про службу святим мені зайво писати до вас,
2COR|9|2|бо відаю вашу охоту, і нею хвалюся за вас македонянам, що Ахая готова з минулого року, а ваша ревність заохотила багатьох.
2COR|9|3|А я послав братів, щоб моя похвала, щодо вас, не даремна була в цім випадкові, але, як казав, щоб були ви приготовані,
2COR|9|4|щоб, коли македоняни прийдуть зо мною та знайдуть, що ви неготові, щоб не осоромитись нам не кажемо вам у цій речі.
2COR|9|5|Отож, я надумався, що треба вблагати братів, щоб пішли перше до вас та приготували заздалегідь оголошений ваш щедрий дар, щоб був він приготований, як щедрий дар, а не річ примусова.
2COR|9|6|А до цього кажу: Хто скупо сіє, той скупо й жатиме, а хто сіє щедро, той щедро й жатиме!
2COR|9|7|Нехай кожен дає, як серце йому призволяє, не в смутку й не з примусу, бо Бог любить того, хто з радістю дає!
2COR|9|8|А Бог має силу всякою благодаттю вас збагатити, щоб ви, мавши завжди в усьому всілякий достаток, збагачувалися всяким добрим учинком,
2COR|9|9|як написано: Розсипав та вбогим роздав, Його справедливість триває навіки!
2COR|9|10|А Той, Хто насіння дає сіячеві та хліб на поживу, нехай дасть і примножить ваше насіння, і нехай Він зростить плоди праведности вашої,
2COR|9|11|щоб усім ви збагачувались на всіляку щирість, яка через нас чинить Богові дяку.
2COR|9|12|Бо діло служіння цього не тільки виповнює недостачі святих, але й багатіє багатьма подяками Богові.
2COR|9|13|Досвідченням цього служіння вони хвалять Бога за послух Христовій Євангелії, що ви визнаєте її, та за щирість учасництва з ними й усіма,
2COR|9|14|вони за вас моляться й тужать по вас із-за дуже великої Божої благодаті на вас.
2COR|9|15|Дяка Богові за невимовний дар Його!
2COR|10|1|А я сам, Павло, благаю вас лагідністю й ласкавістю Христовою; я, коли присутній слухняний між вами, а не бувши між вами сміливий я супроти вас.
2COR|10|2|І благаю, щоб я, прибувши, не осмілився надією, що нею я думаю сміливим бути проти деяких, що про нас вони гадають, ніби ми поступаєм за тілом.
2COR|10|3|Бо ходячи в тілі, не за тілом воюємо ми,
2COR|10|4|зброя бо нашого воювання не тілесна, але міцна Богом на зруйнування твердинь, ми руйнуємо задуми,
2COR|10|5|і всяке винесення, що підіймається проти пізнання Бога, і полонимо всяке знання на послух Христові,
2COR|10|6|і покарати ми готові всякий непослух, коли здійсниться послух ваш.
2COR|10|7|Чи на обличчя ви дивитеся? Як хто певний про себе, що Христовий він, нехай думає знов по собі, що як сам він Христовий, так само Христові й ми.
2COR|10|8|Бо коли б я ще більш став хвалитися нашою владою, яку дав нам Господь на збудування, а не на зруйнування ваше, то не осоромлюсь.
2COR|10|9|Та щоб не здавалось, ніби хочу лякати вас листами.
2COR|10|10|Бо листи його кажуть важкі та міцні, але особисто присутній слабий, а мова його незначна,
2COR|10|11|такий нехай знає оце, що які ми на слові в листах, неприсутніми бувши, такі ми й на ділі, присутніми бувши.
2COR|10|12|Бо не сміємо вважати себе чи рівняти до інших, що самі себе хвалять, вони нерозумно самі себе міряють собою, і рівняють з собою себе.
2COR|10|13|Ми ж не будем хвалитись над міру, а в міру мірила, що його Бог призначив на міру для нас, щоб і до нас досягти.
2COR|10|14|Бо ми не розтягуємося над міру, ніби не досягли ми до вас, бо ми досягли аж до вас із Євангелією Христовою.
2COR|10|15|Ми не хвалимось над міру у чужих працях, але маємо надію, що як буде рости ваша віра, то за нашим мірилом сильно звеличимося ми між вами,
2COR|10|16|щоб і в дальших за вами країнах звіщати Євангелію, а не хвалитись готовим, як це чужі твердять.
2COR|10|17|А хто хвалиться, нехай хвалиться в Господі!
2COR|10|18|Бо достойний не той, хто сам себе хвалить, але кого хвалить Господь!
2COR|11|1|О, коли б потерпіли ви трохи безумство моє! Але й терпите ви мене.
2COR|11|2|Бо пильную про вас пильністю Божою, заручив бо я вас одному чоловікові, щоб Христові привести вас чистою дівою.
2COR|11|3|Та боюсь я, як змій звів був Єву лукавством своїм, щоб так не попсувалися ваші думки, і ви не вхилилися від простоти й чистости, що в Христі.
2COR|11|4|Коли бо хто прийде й зачне проповідувати про Ісуса іншого, про якого ми не проповідували, або приймете іншого Духа, якого ви не прийняли, або іншу Євангелію, якої ви не прийняли, то радо терпіли б ви те!
2COR|11|5|Та думаю я, що нічим не лишаюсь позад передніших апостолів.
2COR|11|6|Хоч і неук я словом, але не знанням, та всюди в усьому ми виявлені поміж вами.
2COR|11|7|Чи я гріх учинив, себе впокоряючи, щоб підвищити вас, бо я Божу Євангелію благовістив для вас дармо?
2COR|11|8|Оббирав я інші Церкви, приймаючи плату для служіння вам. А коли я прийшов до вас і терпів недостачу, то нікого я не обтяжив.
2COR|11|9|Бо мій нестаток поповнили брати, що прийшли з Македонії; і в усьому беріг я себе, щоб не бути для вас тягарем, і збережу.
2COR|11|10|Як правда Христова в мені, так оця похвала не замовчана буде про мене в країнах Ахаї.
2COR|11|11|Для чого? Тому, що я вас не люблю? Відомо те Богові!
2COR|11|12|А що я роблю, те й робитиму, щоб відтяти причину для тих, хто шукає причини, щоб у тому, чим хваляться, показались такі, як і ми.
2COR|11|13|Такі бо фальшиві апостоли, лукаві робітники, що підроблюються на Христових апостолів.
2COR|11|14|І не дивно, бо сам сатана прикидається анголом світла!
2COR|11|15|Отож, не велика це річ, якщо й слуги його прикидаються слугами правди. Буде їхній кінець згідно з учинками їхніми!
2COR|11|16|Знову кажу: хай ніхто не вважає мене за безумного! А як ні, то прийміть мене бодай як безумного, щоб хоч трохи й я похвалився!
2COR|11|17|А що я кажу, не кажу того в Господі, але ніби в безумстві у цій частині хвали.
2COR|11|18|Через те ж, що тілом багато-хто хваляться, то й я похвалюся.
2COR|11|19|Бо ви терпите радо безумних, самі мудрими бувши.
2COR|11|20|Бо ви терпите, коли вас хто неволить, коли хто об'їдає, коли хто обдирає, коли хто підвищується, коли хто по щоках вас б'є.
2COR|11|21|На безчестя кажу, що ми ніби стратили сили. Коли хто відважиться чим, то скажу нерозумно відважуюся й я.
2COR|11|22|Євреї вони? То й я. Ізраїльтяни вони? То й я. Насіння вони Авраамове? То й я!
2COR|11|23|Слуги Христові вони? Говорю нерозумне: більш я! Я був більш у працях, у ранах над міру, частіш у в'язницях, часто при смерті.
2COR|11|24|Від євреїв п'ять раз я прийняв був по сорок ударів без одного,
2COR|11|25|тричі киями бито мене, один раз мене каменували, тричі розбивсь корабель, ніч і день я пробув у глибочині морській;
2COR|11|26|у мандрівках я часто бував, бував у небезпеках на річках, у небезпеках розбійничих, у небезпеках свого народу, у небезпеках поган, у небезпеках по містах, у небезпеках на пустині, у небезпеках на морі, у небезпеках між братами фальшивими,
2COR|11|27|у виснажуванні та в праці, часто в недосипанні, у голоді й спразі, часто в пості, у холоді та в наготі.
2COR|11|28|Окрім зовнішнього, налягають на мене денні повинності й журба про всі Церкви.
2COR|11|29|Хто слабує, а я не слабую? Хто спокушується, а я не палюся?
2COR|11|30|Коли треба хвалитись, то неміччю я похвалюся.
2COR|11|31|Знає Бог і Отець Господа нашого Ісуса Христа, а Він благословенний навіки, що я не говорю неправди.
2COR|11|32|У Дамаску намісник царя Арети стеріг місто Дамаск, щоб схопити мене,
2COR|11|33|але по мурі мене спущено в коші віконцем, і я з рук його втік!
2COR|12|1|Не корисно хвалитись мені, бо я прийду до видінь і об'явлень Господніх.
2COR|12|2|Я знаю чоловіка в Христі, що він чотирнадцять років тому чи в тілі, не знаю, чи без тіла, не знаю, знає Бог був узятий до третього неба.
2COR|12|3|І чоловіка я знаю такого, чи в тілі, чи без тіла, не знаю, знає Бог,
2COR|12|4|що до раю був узятий, і чув він слова невимовні, що не можна людині їх висловити.
2COR|12|5|Отаким похвалюся, а собою хвалитись не буду, хіба тільки своїми немочами.
2COR|12|6|Бо коли я захочу хвалитись, то безумний не буду, бо правду казатиму; але стримуюсь я, щоб про мене хто більш не подумав, ніж бачить у мені або чує від мене.
2COR|12|7|А щоб я через пребагато об'явлень не величався, то дано мені в тіло колючку, посланця сатани, щоб бив в обличчя мене, щоб я не величався.
2COR|12|8|Про нього три рази благав я Господа, щоб він відступився від мене.
2COR|12|9|І сказав Він мені: Досить тобі Моєї благодаті, бо сила Моя здійснюється в немочі. Отож, краще я буду хвалитись своїми немочами, щоб сила Христова вселилася в мене.
2COR|12|10|Тому любо мені перебувати в недугах, у прикростях, у бідах, у переслідуваннях, в утисках через Христа. Коли бо я слабий, тоді я сильний.
2COR|12|11|Хвалячися, я став нерозумний, до того мене ви примусили. Бо хвалити мене мали б ви, бо ні в чому я не залишився позад від найперших апостолів, хоч я й ніщо.
2COR|12|12|А ознаки апостола виявилися між вами в усякім терпінні, у знаменах і чудах та в силах.
2COR|12|13|Що бо є, що ним ви понизилися більше від інших Церков? Хіба те, що я сам тягарем вам не був? Даруйте мені цю провину!
2COR|12|14|Ось утретє готовий прийти я до вас, і не буду для вас тягарем, не шукаю бо вашого я, тільки вас. Не діти повинні збирати маєток батькам, але дітям батьки.
2COR|12|15|Я ж з охотою витрачуся й себе витрачу за душі ваші, хоч що більше люблю вас, то менше я люблений.
2COR|12|16|Та нехай буде так, тягара я на вас не поклав, але, бувши хитрий, я лукавством від вас брав.
2COR|12|17|Чи я використовував вас через когось із тих, кого до вас посилав?
2COR|12|18|Ублагав я був Тита, і з ним послав брата. Чи Тит використав вас чим? Хіба ми ходили не в одному дусі? Хіба не одними стопами?
2COR|12|19|Чи ви знову не думаєте, що виправдуємось перед вами? Перед Богом, у Христі ми говоримо, а все, любі, на вашу будову!
2COR|12|20|Я ж боюся, щоб, прийшовши, не знайшов вас такими, якими не хочу, і щоб мене не знайшли ви таким, якого не хочете, хай не будуть між вами суперечка, заздрість, гніви, обмани, свари, нашепти, пихи, безладдя,
2COR|12|21|щоб знову, коли я прийду, не принизив мене поміж вами мій Бог, і щоб мені не оплакувати багатьох, що перше згрішили були, і не покаялися в нечистості, і в перелюбі, і в розпусті, що коїли їх.
2COR|13|1|Оце втретє до вас я йду. Кожна справа хай станеться вироком двох чи трьох свідків.
2COR|13|2|Попереджував я й попередую, як у вас був удруге, так тепер неприсутній, отих, що згрішили перед тим, і всіх інших, що коли прийду знову, то я не помилую,
2COR|13|3|через те, що шукаєте доказу, що в мені промовляє Христос, Який не безсилий до вас, але сильний у вас.
2COR|13|4|Бо хоч Він був і розп'ятий в немочі, та живий із сили Божої. Так і ми, хоча немічні в Нім, та з Ним будемо жити з Божої сили у вас.
2COR|13|5|Випробовуйте самих себе, чи ви в вірі, пізнавайте самих себе. Хіба ви не знаєте самих себе, що Ісус Христос у вас? Хіба тільки, що ви не такі, якими мали б бути.
2COR|13|6|Але маю надію, що пізнаєте ви, що ми такі, якими мали б бути.
2COR|13|7|І ми молимо Бога, щоб ви не чинили ніякого лиха, не для того, щоб виявились ми досвідчені, а щоб учинили ви добре, а ми будем немов негідні.
2COR|13|8|Бо нічого не можемо ми проти правди, а за правду.
2COR|13|9|Ми тішимося, коли ми слабі, а ви сильні. Про це й молимось щоб були досконалими ви!
2COR|13|10|Ось тому то, відсутній, пишу це, щоб прийшовши, не мав я вчинити суворо за владою, якої Господь мені дав на будування, а не на руйнування.
2COR|13|11|А накінець, браття, радійте, удосконалюйтесь, тіштеся, будьте однодумні, майте мир, і Бог любови та миру буде з вами!
2COR|13|12|Вітайте один одного святим поцілунком!
2COR|13|13|(13-12) Усі святі вас вітають!
2COR|13|14|(13-13) Благодать Господа нашого Ісуса Христа, і любов Бога й Отця, і причастя Святого Духа нехай буде зо всіма вами! Амінь.
