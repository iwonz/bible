NAH|1|1|Пророцтво на Ніневію. Книга видіння елкошейця Наума.
NAH|1|2|Палкий Бог, і мстивий Господь, Господь мстивий та лютий, Господь мстивий до тих, хто Його ненавидить, і пам'ятає про кривду Своїх ворогів.
NAH|1|3|Господь довготерпеливий і великої потуги, та очистити винного Він не очистить. Господь у бурі та в вихрі дорога Його, а хмара від стіп Його курява.
NAH|1|4|Як загнівається Він на море, то сушить його, і всі ріки висушує, в'яне Башан та Кармел, і в'яне та квітка Лівану.
NAH|1|5|Гори тремтять перед Ним, а підгірки топніють, перед обличчям Його трясеться земля та вселенна, та всі її мешканці.
NAH|1|6|Хто встоїть перед гнівом Його, і хто стане у полум'ї люті Його? Його шал виливається, мов той огонь, і розпадаються скелі від Нього!
NAH|1|7|Добрий Господь, пристановище Він у день утиску, і знає Він тих, хто на Нього надіється!
NAH|1|8|Але в зливі навальній Він зробить кінця між Його заколотниками, і ворогів зажене у темноту.
NAH|1|9|Що ви думаєте проти Господа? Бо Він зробить кінця, не постане два рази насильство.
NAH|1|10|Бо вони переплутані, наче той терен, і повпивались, немов би вином, вони будуть пожерті зовсім, мов солома суха!
NAH|1|11|З тебе вийшов задумуючий проти Господа лихо, радник нікчемний.
NAH|1|12|Так говорить Господь: Хоч були б найсильніші і дуже численні, та постинані будуть вони, та й минуться! І хоч Я тебе мучив, та мучити більше тебе вже не буду!
NAH|1|13|А тепер Я зламаю ярмо його, яке на тобі, і пута твої позриваю.
NAH|1|14|І накаже на тебе, Ашшуре, Господь: Більш не буде вже сіятися з твого ймення! З дому бога твого Я боввана та ідола витну, зроблю тобі гроба із них, бо ти став легковажений.
NAH|1|15|(2-1) Ось на горах ноги благовісника, що звіщає про мир: Святкуй, Юдо, свята свої, виконуй присяги свої, бо більше не буде нікчемний ходити по тобі, він витятий ввесь!
NAH|2|1|(2-2) На тебе йде розпорошувач, твердині свої стережи, виглядай на дорогу, зміцняй свої стегна, міцно скріпи свою потугу,
NAH|2|2|(2-3) бо верне Господь велич Якова, як велич Ізраїля, що їхні спустошителі поруйнували, і понищили їхні виноградні галузки.
NAH|2|3|(2-4) Щит хоробрих його зачервонений, вояки в кармазині; блищить сталь у день зброєння їхнього на колесницях, хвилюються ратища.
NAH|2|4|(2-5) Колесниці шалено по вулицях мчать, по майданах гуркочуть, їхній вид немов полум'я те смолоскипів, літають вони, як ті блискавки.
NAH|2|5|(2-6) Він згадає шляхетних своїх, та спіткнуться вони у ході своїй; вони поспішають на мури її, і поставлена міцно будівля облоги.
NAH|2|6|(2-7) Брами річок відчиняються, а палата руйнується.
NAH|2|7|(2-8) І постановлено: буде оголена, відведеться в полон, а рабині її голоситимуть, мов ті голубки, що воркують на персах своїх.
NAH|2|8|(2-9) І Ніневія як саджавка водна, що води її відпливають. Стійте, стійте! Та немає нікого, хто б їх завернув!
NAH|2|9|(2-10) Розграбовуйте срібло, розграбовуйте золото, немає кінця наготовленому, багатству коштовних речей.
NAH|2|10|(2-11) Знищення та зруйнування й спустошення буде... І серце розтопиться, і ноги дрижатимуть, і корчі по крижах усіх, а обличчя їх всіх на червоно розпаляться.
NAH|2|11|(2-12) Де леговище левів, і для левчуків пасовище, що там ходив лев та левиця, та левеня, і ніхто не лякав?
NAH|2|12|(2-13) Лев грабував для своїх молодят і душив для левиць своїх він, і печери свої переповнював здобиччю, а лігва свої награбованим.
NAH|2|13|(2-14) Ось Я проти тебе, говорить Господь Саваот, і попалю серед диму твої колесниці, а твоїх левчуків поїсть меч, і повитинаю з землі грабування твої, і вже не почується голос твого посла.
NAH|3|1|Горе місту цьому кровожерному, воно все неправда, воно повне насилля, грабіж не виходить із нього!
NAH|3|2|Чути свист батога, гуркіт колеса, і чвал коней, і колеснична гуркотнява,
NAH|3|3|і гін верхівця, і полум'я меча, і блиск ратища, і багато побитих, і мертвих велике число, і трупу немає кінця, і спотикатимуться об їхній труп,
NAH|3|4|це за многоту блудодійства розпусниці, привабно ласкавої, вправної в чарах, що народи за блуд свій вона продавала, а роди за чари свої.
NAH|3|5|Ось Я проти тебе, говорить Господь Саваот, і подолка твого підійму на обличчя твоє, і покажу Я твій сором народам, а царствам твій стид!
NAH|3|6|І кину на тебе огиди, і погордженою вчиню Я тебе, і зроблю Я тебе, мов позорище!
NAH|3|7|І станеться, кожен, хто вгледить тебе, від тебе втече та й прокаже: Пограбована Ніневія! Хто висловить їй співчуття? Звідки буду шукати тобі потішителів?
NAH|3|8|Чи краща ти від Но-Амона, що сидить серед рік, вода коло нього, що вал його море, від моря його мур?
NAH|3|9|Етіопія сила його, і Єгипет, і не має кінця. Пут та лівійці були тобі в поміч,
NAH|3|10|та й він на вигнання пішов, у полон... А діти його порозбивані на роздоріжжі всіх вулиць, і кидали жереб про славних його, й всі вельможі його у кайдани закуті.
NAH|3|11|Уп'єшся і ти, будеш схована, твердині від ворога будеш шукати і ти!
NAH|3|12|Всі фортеці твої, мов ті фіґи з доспілими овочами: коли затрясуться, то падають в уста того, хто їх їсть.
NAH|3|13|Ось народ твій немов ті жінки серед тебе: вони повідчиняють твоїм ворогам брами краю твого, огонь пожере твої засуви.
NAH|3|14|Води на облогу собі набери, твердині свої позміцняй, увійди до болота та в глині топчись, форму на цеглу візьми міцно в руку.
NAH|3|15|Там огонь тебе з'їсть, посіче тебе меч, пожеруть тебе, наче та гусінь. Стань численна, як гусінь, стань численна, немов сарана,
NAH|3|16|понамножуй купців своїх більше від зірок небесних, але гусінь та знищить тебе й полетить!
NAH|3|17|Вельможні твої немов та сарана, гетьмани твої мов мошва, що гніздиться по стінах в день холоду, але сонце засвітить і вони помандрують, і не пізнане буде те місце, де вони пробували.
NAH|3|18|Твої пастирі, царю асирійський, поснули, лежать вельможі твої, твій народ розпорошивсь по горах, і немає кому позбирати його.
NAH|3|19|Нема ліку для лиха твого, рана твоя невигойна! Всі, що звістку про тебе почують, заплещуть у долоні на тебе, бо над ким твоє зло не ходило постійно?
