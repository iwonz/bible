1CHR|1|1|Адам 121, Сиф 8352, Енош 583,
1CHR|1|2|Кенан 7018, Магалел'їл 4111, Яред 3382,
1CHR|1|3|Енох 2585, Метушелах 4968, Ламех 3929,
1CHR|1|4|Ной 5146, Сим 8035, Хам 2526 та Яфет 3315.
1CHR|1|5|Сини 1121 Яфетові 3315: Ґомер 1586, і Маґоґ 4031, і Мадай 4074, і Яван 3120, і Тувал 8422, і Мешех 4902, і Тірас 8494.
1CHR|1|6|А сини 1121 Ґомерові 1586: Ашкеназ 813 і Діфат 7384, і Тоґарма 8425.
1CHR|1|7|А сини 1121 Яванові 3120: Еліша 473 й Таршіша 8659, кіттяни 3794 й роданяни 1721.
1CHR|1|8|Сини 1121 Хамові 2526: Куш 3568 і Міцраїм 4714, Пут 6316 і Ханаан 3667.
1CHR|1|9|А сини 1121 Кушеві 3568: Шева 5434, і Хавіла 2341, і Савта 5454, і Раама 7484, і Савтеха 5455. А сини 1121 Рамині 7484: Шева 7614 й Дедан 1719.
1CHR|1|10|А Куш 3568 породив 3205 8804 Німрода 5248, він зачав 2490 8689 бути велетом 1368 на землі 776.
1CHR|1|11|А Міцраїм 4714 породив 3205 8804 лудян 3866, і анам'ян 6047, і легав'ян 3853, і нафтух'ян 5320,
1CHR|1|12|і патрусян 6625, і каслух'ян 3695, що вийшли 3318 8804 звідти филистимляни 6430, і кафторян 3732.
1CHR|1|13|А Ханаан породив Сидона, свого первородженого, і Хета,
1CHR|1|14|і євусеянина, і амореянина, і ґірґашеянина,
1CHR|1|15|і хіввеянина, і аркеянина, і сінеянина,
1CHR|1|16|і арвадянина, і цемарянина, і хаматянина.
1CHR|1|17|Сини Симові: Елам, і Ашшур, і Арпахшад, і Луд, і Арам. Сини Арамові: і Уц, і Хул, і Ґетер, і Мешех.
1CHR|1|18|А Арпахшад породив Шалаха, а Шалах породив Евера.
1CHR|1|19|А Еверові народилося двоє синів, ім'я одному Пелеґ, бо за його днів була поділена земля, а ім'я брата його Йоктан.
1CHR|1|20|А Йоктан породив Алмодада, і Шелефа, і Хацармавета, і Єраха,
1CHR|1|21|і Гадорама, і Узала, і Діклу,
1CHR|1|22|і Евала, і Авімаїла, і Шеву,
1CHR|1|23|і Офіра, і Хавілу, і Йовава, усі вони сини Йоктанові.
1CHR|1|24|Сим, Арпахшад, Шелах,
1CHR|1|25|Пелеґ, Реу,
1CHR|1|26|Серуґ, Нахор, Терах,
1CHR|1|27|Аврам, він же Авраам.
1CHR|1|28|Сини Авраамові: Ісак та Ізмаїл.
1CHR|1|29|Оце їхні нащадки: первороджений Ізмаїлів Невайот, і Кедар, і Адбеїл, і Мівсам,
1CHR|1|30|Мішма, і Дума, Масса, Хадад, і Тема,
1CHR|1|31|Єтур, Нафіш, і Кедема, оце вони сини Ізмаїлові.
1CHR|1|32|А сини Кетури, Авраамової наложниці: вона породила Зімрана, і Йокшана, і Медана, і Мідіяна, і Їшбака, і Шуаха. А Йокшанові сини: Шева й Дедан.
1CHR|1|33|А Мідіянові сини: Ефа, і Ефер, і Ханох, і Авіда, і Елдаа, ці всі сини Кетури.
1CHR|1|34|А Авраам породив Ісака. Ісакові сини: Ісав і Ізраїль.
1CHR|1|35|Ісавові сини: Еліфаз, Реуїл, і Єуш, і Йалам, і Кора.
1CHR|1|36|Сини Еліфазові: Теман і Омар, Цефі й Ґатам, Кеназ і Тімна, і Амалик.
1CHR|1|37|Сини Реуїлові: Нахат, Зерах, Шамма й Мізза.
1CHR|1|38|А сини Сеїрові: Лотан, і Шовал, і Ців'он, і Ана, і Дішон, і Ецер, і Дішан.
1CHR|1|39|А сини Лотанові: Хорі, і Гомам, і Ахот, Лотан, Тімна.
1CHR|1|40|Сини Шовалові: Ал'ян, і Манахат, і Евал, Шефі, і Онам. А сини Ців'онові: Айя й Ана.
1CHR|1|41|А сини Анині: Дішон. А сини Дішонові: Хамран, і Ешбан, і Їтран, і Керан.
1CHR|1|42|Сини Ецерові: Білган, і Зааван, Яакан. Сини Дішонові: Уц та Аран.
1CHR|1|43|А оце царі, що царювали в Едомовому краї перед зацарюванням царя в Ізраїлевих синів: Бела, Беорів син, а ім'я його міста Дінгава.
1CHR|1|44|І помер Бела, а замість нього зацарював Йовав, Зерахів син з Боцри.
1CHR|1|45|І помер Йовав, а замість нього зацарював Хушам із краю теманянина.
1CHR|1|46|І помер Хушам, а замість нього зацарював Гадад, Бедадів син, що побив був Мідіяна на Моавському полі, а ім'я місту його Авіт.
1CHR|1|47|І помер Гадад, а замість нього зацарював Самла з Масреки.
1CHR|1|48|І помер Самла, а замість нього зацарював Саул з Рехевот-Ганнагару.
1CHR|1|49|І помер Саул, а замість нього зацарював Баал-Ханан, син Ахборів.
1CHR|1|50|І помер Баал-Ханан, а замість нього зацарював Гадад, а ім'я його міста Раї, а ім'я жінки його Мегетав'їл, дочка Матреда, дочки Ме-Загавової.
1CHR|1|51|І помер Гадад. І були потому провідники Едому: провідник Тімна, провідник Ал'я, провідник Єтет,
1CHR|1|52|провідник Оголівама, провідник Ела, провідник Пінон,
1CHR|1|53|провідник Кеназ, провідник Теман, провідник Мівцар,
1CHR|1|54|провідник Маґдіїл, провідник Ірам, оце провідники Едому.
1CHR|2|1|Оце Ізраїлеві сини: Рувим, Симеон, Левій, і Юда, Іссахар, і Завулон,
1CHR|2|2|Дан, Йосип, Веніямин, Нефталим, Ґад і Асир.
1CHR|2|3|Юдині сини: Ер, і Онан, і Шела, троє народилися йому від ханаанеянки Бат-Шуї. І був Ер, Юдин первороджений, нечестивий в очах Господа, і Він забив його.
1CHR|2|4|А Тамар, невістка його, породила йому Переца та Зеваха, усіх Юдиних синів п'ятеро.
1CHR|2|5|Сини Перецові: Хецрон та Хамул.
1CHR|2|6|А сини Зерахові: Зімрі, і Етан, і Геман, і Калкол, і Дера, усіх їх п'ятеро.
1CHR|2|7|А Кармієві сини: Ахар, що напровадив біду на Ізраїля, що спроневірився в заклятті.
1CHR|2|8|А сини Етанові: Азарія.
1CHR|2|9|А сини Хецронові, що народилися йому: Єрахмеїл, і Рам, і Келувай.
1CHR|2|10|А Рам породив Аммінадава, а Аммінадав породив Нахшона, начальника синів Юдиних.
1CHR|2|11|А Нахшон породив Салму, а Салма породив Боаза,
1CHR|2|12|а Боаз породив Оведа, а Овед породив Єссея.
1CHR|2|13|А Єссей породив свого первородженого Еліава, і Авінадава другого, і Шім'у третього,
1CHR|2|14|Натаніїла четвертого, Раддая п'ятого,
1CHR|2|15|Оцема шостого, Давида сьомого.
1CHR|2|16|А їхні сестри: Церуя й Авідаїл. А Церуїні сини: Авшай, і Йоав, і Аса-Ел, усіх троє.
1CHR|2|17|А Авіґаїл породила Амасу, а батько Амасин їшмеелянин Єтер.
1CHR|2|18|А Калев, Хецронів син, породив зо своєю жінкою Азувою та з Еріот дітей. А оце сини її: Єшер, і Шовав, і Ардон.
1CHR|2|19|І померла Азува, а Калев узяв собі Ефрату, і вона породила йому Хура.
1CHR|2|20|А Хур породив Урі, а Урі породив Бецаліїла.
1CHR|2|21|А потому прийшов Хецрон до дочки Махіра, Ґілеадового батька, і він узяв її, а він був віку шостидесяти років, і вона породила йому Сеґува.
1CHR|2|22|А Сеґув породив Яіра, і він мав двадцять і три місті в ґілеадському краї.
1CHR|2|23|Але Ґешур та Арам забрали від них Яірові оселі, Кенат та залежні від нього міста, шістдесят міст. Усе це сини Махіра, Ґілеадового батька.
1CHR|2|24|А по Хецроновій смерті прийшов Калев до Єфрати, і Хецронова жінка Авійя породила йому Ашхура, батька Текої.
1CHR|2|25|А сини Єрахмеїла, Хецронового первородженого, були: первороджений Рам, і Буна, і Орен, і Оцем, Ахійя.
1CHR|2|26|І була в Єрахмеїла інша жінка, а ім'я їй Атара, вона мати Онама.
1CHR|2|27|А сини Рама, Єрахмеїлового первородженого, були: Маац, і Ямін, і Екер.
1CHR|2|28|А сини Онамові були: Шаммай, і Яда. А сини Шаммая: Надав та Авішур.
1CHR|2|29|А ім'я Авішуровій жінці Авіхаїл, і вона породила йому Ахбана та Моліда.
1CHR|2|30|А сини Надавові: Селед та Аппаїм, а Селед помер без дітей.
1CHR|2|31|А сини Аппаїмові: Їш'ї. А сини Їш'ї: Шешан. А сини Шешанові: Ахлай.
1CHR|2|32|А сини Яди, Шаммаєвого брата: Єтер і Йонатан. І помер Єтер без дітей.
1CHR|2|33|А Йонатанові сини: Пелет, і Заза, оце були сини Єрахмеїлові.
1CHR|2|34|А в Шешана не було синів, а тільки дочки. Був у Шешана раб єгиптянин, а ім'я йому Ярха.
1CHR|2|35|І дав Шешан рабові своєму Ярсі свою дочку за жінку, і вона породила йому Аттая.
1CHR|2|36|А Аттай породив Натана, а Натан породив Завада,
1CHR|2|37|А Завад породив Ефлала, а Ефлал породив Оведа.
1CHR|2|38|А Овед породив Єгу, а Єгу породив Азарію,
1CHR|2|39|а Азарія породив Хелеца, а Хелец породив Ел'асу.
1CHR|2|40|А Ел'аса породив Сісмая, а Сісмай породив Шаллума.
1CHR|2|41|А Шаллум породив Єкамію, а Єкамія породив Елішаму.
1CHR|2|42|А сини Калева, Єрахмеїлового брата: Меша, його первороджений, він батько Зіфа. І сини Мареші, Хевронового батька.
1CHR|2|43|А Хевронові сини: Корах, і Таппуах, і Рекем, і Шама.
1CHR|2|44|А Шама породив Рахама, Єракеамового батька, а Рекем породив Шаммая.
1CHR|2|45|А сини Шаммаєві: Маон, а Маон був основник Бет-Цуру.
1CHR|2|46|А Ефа, наложниця Калева, породила Харана, і Моцу, і Ґазеза. А Харан породив Ґазеза.
1CHR|2|47|А сини Єгдаєві: Реґем, і Йотам, і Ґешан, і Фелет, і Ефа, і Шааф.
1CHR|2|48|Калевова наложниця Мааха породила Шевера та Тірхату.
1CHR|2|49|І породила вона Шаафа, батька Мадманни, Шеву, батька Махбени, та батька Ґів'и. А дочка Калевова Ахса.
1CHR|2|50|Оце були сини Калева, сина Гура, первородженого Ефрати: Шовал, батько Кір'ят-Єаріму,
1CHR|2|51|Салма, батько Віфлеєма, Гареф, батько Бе-Ґадеру.
1CHR|2|52|У Шовала, батька Кір'ят-Єаріму, були сини: Гарое, Хаці-Гамменухот.
1CHR|2|53|А роди Кір'ят-Єаріма: їтряни, путяни, шуматяни, мішраяни, від них пішли цор'атяни та єштауляни.
1CHR|2|54|Сини Салмині: Бет-Лехем, і нетофаляни, Атрот, Бет-Йоав, і хаці-гаммонахтяни, цоряни.
1CHR|2|55|А роди писарів, мешканців Ябецу, тір'атяни, шім'атяни, сухатяни, вони кіняни, що походять від Хамата, батька Бет-Рехавового.
1CHR|3|1|А оце були Давидові сини, що народилися йому в Хевроні: первороджений Амнон, від їзреелітянки Ахіноам; другий Даниїл, від кармелітянки Авіґаїл;
1CHR|3|2|третій Авесалом, син Маахи, дочки Талмая, царя ґешурського; четвертий Адонійя, син Хаґґіт;
1CHR|3|3|п'ятий Шефатія, від Авітал; шостий Їтреам, від жінки його Еґли;
1CHR|3|4|шестеро народжено йому в Хевроні. І царював він там сім років і шість місяців, а тридцять і три роки царював в Єрусалимі.
1CHR|3|5|А оці народилися йому в Єрусалимі: Шім'а, і Шовав, і Натан, і Соломон, четверо від Вірсавії, Амміїлової дочки,
1CHR|3|6|і Ївхар, і Елішама, і Еліфалет,
1CHR|3|7|і Ноґаг, і Нефеґ, і Яфія,
1CHR|3|8|і Елішама, і Еліяда, і Еліфелет, дев'ятеро.
1CHR|3|9|Усе це Давидові сини, окрім синів наложниць та сестри їх Тамари.
1CHR|3|10|А син Соломонів Рехав'ам, його син Авійя, його син Аса, його син Йосафат,
1CHR|3|11|його син Йорам, його син Ахазія, його син Йоаш,
1CHR|3|12|його син Амація, його син Азарія, його син Йотам,
1CHR|3|13|його син Ахаз, його син Хізкійя, його син Манасія,
1CHR|3|14|його син Амон, його син Йосія.
1CHR|3|15|А сини Йосії: первороджений Йоханан, другий Єгояким, третій Седекія, четвертий Шаллум.
1CHR|3|16|А сини Єгоякимові: Єхонія син його, та син його Седекія.
1CHR|3|17|А сини Єхонії: Ассір, Шеал'тіїл, син його,
1CHR|3|18|і Малкірам, і Педая, і Шен'аццар, Єкам'я, Гошама, і Недав'я.
1CHR|3|19|А сини Педаї: Зоровавель і Шім'ї. А сини Зоровавеля: Мешуллам, і Хананія, і сестра їхня Шеломіт,
1CHR|3|20|і Хашува, і Огел, і Верех'я, і Хасад'я, Юшав-Хесед, п'ятеро.
1CHR|3|21|А сини Хананії: Пелатія та Єшая, сини Рефаї, сини Арнонові, сини Овадії, сини Шеханії.
1CHR|3|22|А сини Шеханії: Шемая. А сини Шемаї: Хаттиш, і Їґ'ал, і Баріах, і Неарія, і Шафат, шестеро.
1CHR|3|23|А сини Неарії: Ел'йоенай, і Хізкійя, і Азрікам, троє.
1CHR|3|24|А сини Ел'йоенаєві: Годав'я, і Ел'яшів, і Пелая, і Аккув, і Йоханан, і Делая, і Анані, семеро.
1CHR|4|1|Сини Юдині: Перец, Хецрон, і Кармі, і Хур, і Шовал.
1CHR|4|2|А Реая, син Шовалів, породив Яхата, а Яхат породив Ахумая та Лахада, оце роди цор'атян.
1CHR|4|3|А оці Аві-Етамові: Їзреел, і Їшма, і Їдбаш, а ім'я їхній сестрі Гаццелелпоні.
1CHR|4|4|А Пенуїл батько Ґедора, а Езер батько Хуші. Оце сини Хура, Єфремового первородженого, батька Віфлеєму.
1CHR|4|5|А в Ашхура, батька Текої, були дві жінки: Хел'а та Наара.
1CHR|4|6|І породила йому Наара Ахуззама, і Хефера, і Темені, і Ахаштарі, оце сини Наарині.
1CHR|4|7|А сини Хел'ині: Церет, і Цохар, і Етнан.
1CHR|4|8|А Коц породив Анува, і Гаццовеву, і роди Ахархела, сина Гарумового.
1CHR|4|9|А Ябец був поважаний більше від своїх братів, і мати його назвала йому ім'я Ябец, говорячи: Я породила його в болісті.
1CHR|4|10|кликнув Ябец до Бога Ізраїлевого, говорячи: Коли б Ти, благословляючи, поблагословив мене, і побільшив границю мою, і рука Твоя була зо мною, і зробив охорону від лиха, щоб не засмучувати мене! І Бог послав, чого він просив.
1CHR|4|11|А Келув, брат Шухи, породив Мехіра, він батько Ештона.
1CHR|4|12|А Ештон породив Бет-Рафу, і Пасеаха, і Техінну, батька міста Нахаша. Це люди Рехи.
1CHR|4|13|А сини Кеназа: Отніїл та Серая. А сини Отніїлові: Хатат.
1CHR|4|14|А Меонотай породив Офру, а Серая породив Яава, батька Ремісничої Долини, бо вони були ремісники.
1CHR|4|15|А сини Калева, Єфуннеєвого сина: Іру, Ела та Наам. А Елин син Кеназ.
1CHR|4|16|А сини Єгаллел'їлові: Зіф і Зіфа, Тір'я й Асар'їл.
1CHR|4|17|А сини Езри: Єтер, і Меред, і Ефер, і Ялон. А оце сини Біт'ї, фараонової дочки, що взяв Меред; і вона зачала й породила Мір'яма, і Шаммая, і Їшбаха, батька Ештемої.
1CHR|4|18|А жінка його юдеянка породила Єреда, батька Ґедору, і Хевера, батька Сохо, і Єкутіїла, батька Заноаха.
1CHR|4|19|А сини жінки Годійї, сестри Нахама, батька ґарм'янина Кеїли та маахатянина Ештемоа,
1CHR|4|20|а сини Симеонові: Амнон, і Рінна, Бен-Ханан, і Тілон. А сини Їш'ї: Зохет та Бен-Зохет.
1CHR|4|21|Сини Шели, Юдиного сина: Ер, батько Лехи, і Лада, батько Мареші, і роди дому робітників віссону, з дому Ашбеа.
1CHR|4|22|І Йокін, і люди Козеви, і Йоаш, і Сараф, що володіли Моавом, і Яшуві-Лехем. Та це справи стародавні.
1CHR|4|23|Вони були ганчарі, і замешкували садки та городи; вони жили там у царя для його роботи.
1CHR|4|24|Сини Симеонові: Немуїл, і Ямім, Ярів, Зерах, Саул,
1CHR|4|25|його син Шаллум, його син Мівсам, його син Мішма.
1CHR|4|26|А сини Мішми: Хаммуїл син його, його син Заккур, його син Шім'ї.
1CHR|4|27|А в Шім'ї було шістнадцять синів та шість дочок, а брати його не мали багатьох синів, і не помножили ввесь свій рід так, як сини Юдині.
1CHR|4|28|І осілися вони в Беер-Шеві, і в Моладі, і в Хацар-Шуалі,
1CHR|4|29|і в Білзі, і в Ецемі, і в Толаді,
1CHR|4|30|і в Бетуїлі, і в Хормі, і в Ціклаґу,
1CHR|4|31|і в Бет-Маркавоті, і в Хацар-Сусімі, і в Бет-Бір'і, і в Шаараїмі, оце їхні міста аж до зацарювання Давидового.
1CHR|4|32|А їхні осади: Етам, і Аїн, Ріммон, і Тохен, і Ашан, п'ятеро міст.
1CHR|4|33|А всі їхні осади, що навколо тих міст, аж до Баалу; це місця їх оселення та родоводи їх про них.
1CHR|4|34|А Мешовав, і Ямлех, і Йоша, син Амації,
1CHR|4|35|і Йоїл, і Єгу, син Йошів'ї, сина Сераї, сина Асіїлового,
1CHR|4|36|і Елйоенай, і Якова, і Шохая, і Асая, і Адіїл, і Єсіміїл, і Беная,
1CHR|4|37|і Зіза, син Шіф'і, сина Аллона, сина Єдаї, сина Шімрі, сина Шемаї.
1CHR|4|38|Це ті, що входять в імена князів у свої роди, а дім своїх батьків сильно розмножили.
1CHR|4|39|І пішли вони до Мево-Ґедору, аж до східнього боку долини, щоб пошукати пасовиська для своїх отар.
1CHR|4|40|І знайшли вони пасовисько сите та добре, а той край був просторий, і тихий та спокійний, бо від Хама походили ті, що сиділи там колись.
1CHR|4|41|І пішли ці, записані іменами за днів Єзекії, царя Юдиного, і розбили їхні намети там, і побили меінітів, що були знайдені там, що їх учинили закляттям аж до цього дня, й осілися замість них, бо там пасовисько для їхньої дрібної худоби.
1CHR|4|42|А з них, з Симеонових синів, пішли на гору Сеїр п'ять сотень чоловіка, а Пелатія, і Неарія, і Рефая, і Уззіїл, сини Їш'ї, були на чолі їх.
1CHR|4|43|І вони побили останок урятованих Амалика, й осілися там аж до цього дня.
1CHR|5|1|А сини Рувима, Ізраїлевого первородженого, бо він первороджений, та за збезчещення ним ложа свого батька перворідство було дане синам Йосипа, сина Ізраїлевого, та вони не могли приписатися до перворідства.
1CHR|5|2|Бо Юда став найсильнішим серед братів своїх, і князем, сильнішим від нього, а перворідство дісталося Йосипові.
1CHR|5|3|Сини Рувима, Ізраїлевого первородженого: Ханох і Паллу, Хецрон і Кармі.
1CHR|5|4|Йоїлові сини: Шемая син його, його син Ґоґ, син його Шім'ї,
1CHR|5|5|син його Міха, син його Реая, син його Баал,
1CHR|5|6|син його Беера, якого вигнав Тіллеґат-Пілнеесер, цар асирійський. Він був начальником Рувимівців.
1CHR|5|7|А брати його, за його родами, у приписуванні за потомством їх, були: голова Єіїл, і Захарій,
1CHR|5|8|і Бела, син Азаза, сина Шеми, Йоїлового сина, він сидів в Ароері й аж по Нево та Баал-Меон.
1CHR|5|9|А на схід він сидів аж до виходу на пустиню від річки Ефрат, бо їхні череди в ґілеадському краї стали численні.
1CHR|5|10|А за Саулових днів вони провадили війну з агарянами, і ті впали в їхні руки, а вони сиділи в їхніх наметах на всім просторі на схід від Ґілеаду.
1CHR|5|11|А Ґадові сини сиділи навпроти них у башанському краї аж до Салхи.
1CHR|5|12|Йоїл голова, а Шафам другий, і Янай, і Шафат у Башані.
1CHR|5|13|А їхні браття за домами своїх батьків: Михаїл, і Мешуллам, і Шева, і Йорай, і Якан, і Зія, і Евер, семеро.
1CHR|5|14|Оце сини Авіхаїла, сина Хурі, сина Яроаха, сина Ґілеада, сина Михаїла, сина Єшішая, сина Єхдо, сина Буза.
1CHR|5|15|Ахі, син Авдіїла, сина Ґунієвого, голови дому батьків їх.
1CHR|5|16|І сиділи вони в Ґілеаді, в Башані та в залежних від нього містах, та в усіх пасовиськах Шарону, на місцях виходу їх.
1CHR|5|17|Усі вони були переписані в днях Йотама, Юдиного царя, та в днях Єровоама, царя Ізраїлевого.
1CHR|5|18|Синів Рувима, і ґадян, і половини Манасіїного племени, людей військових, що носять щита й меча та натягують лука, та випрактикуваних у війні було сорок і чотири тисячі і сім сотень і шістдесят, що виходили з військом.
1CHR|5|19|І провадили вони війну з агарянами, і з Ітуром, і з Нафішем, і з Нодавом.
1CHR|5|20|І дана була їм поміч на них, і віддані були в їхню руку ті агаряни та всі, що з ними, бо вони кликали до Бога в бою, і Він був ублаганий, бо вони надіялися на Нього.
1CHR|5|21|І вони зайняли їхні череди: їхніх верблюдів п'ятдесят тисяч, і дрібної худоби двісті й п'ятдесят тисяч, і ослів дві тисячі, а людських душ сто тисяч.
1CHR|5|22|Бо трупів попадало багато, бо від Бога була ця війна. І сиділи вони на своєму місці аж до неволі.
1CHR|5|23|А сини половини Манасіїного племени сиділи в краю від Башану аж до Баал-Хермону й Сеніру та гори Гермону. Вони розмножилися.
1CHR|5|24|А оце голови домів їхніх батьків: і Ефер, і Їш'ї, і Еліїл, і Азріїл, і Їрмея, і Годавія, і Яхдіїл, мужі відважні, мужі славні, голови домів їхніх батьків.
1CHR|5|25|Та спроневірилися вони Богові своїх батьків, і блудили за богами народів Краю, яких Бог вигубив перед ними.
1CHR|5|26|І Бог Ізраїлів збудив духа Пула, царя асирійського, і духа Тілленат-Піл'несера, царя асирійського, і він виселив їх, Рувимівців і Ґадівців та половину Манасіїного племени, і запровадив їх у Халах, і Хавор, і Хару, та до річки Ґозан, і вони там аж до цього дня.
1CHR|6|1|(5-27) Левієві сини: Ґершон, Кегат і Мерарі.
1CHR|6|2|(5-28) А сини Кегатові: Амрам, Їцхар, Хеврон, і Уззіїл.
1CHR|6|3|(5-29) А сини Амрамові: Аарон, і Мойсей, і Міріям. А сини Ааронові: Надав і Авігу, Елеазар і Ітамар.
1CHR|6|4|(5-30) Елеазар породив Пінхаса, Пінхас породив Авішую,
1CHR|6|5|(5-31) а Авішуя породив Буккі, а Буккі породив Уззі.
1CHR|6|6|(5-32) А Уззі породив Зерахію, а Зерахія породив Мерайота.
1CHR|6|7|(5-33) Мерайот породив Амарію, а Амарія породив Ахітува.
1CHR|6|8|(5-34) А Ахітув породив Садока, а Садок породив Ахімааца.
1CHR|6|9|(5-35) А Ахімаац породив Азарію, а Азарія породив Йоханана.
1CHR|6|10|(5-36) А Йоханан породив Азарію, це той, що був священиком у Господньому домі, якого вибудував Соломон в Єрусалимі.
1CHR|6|11|(5-37) І Азарія породив Амарію, а Амарія породив Ахітува.
1CHR|6|12|(5-38) А Ахітув породив Садока, а Садок породив Шаллума.
1CHR|6|13|(5-39) А Шаллум породив Хілкійю, а Хілкійя породив Азарію.
1CHR|6|14|(5-40) А Азарія породив Сераю, а Серая породив Єгоцадака.
1CHR|6|15|(5-41) А Єгоцадак пішов до неволі, коли Господь вивів Юду та Єрусалим через Навуходоносора.
1CHR|6|16|(6-1) Сини Левієві: Ґершом, Кегат та Мерарі.
1CHR|6|17|(6-2) А оце ймення Ґершомових синів: Лівні та Шім'ї.
1CHR|6|18|(6-3) А сини Кегатові: Амрам, і Їцхар, і Хеврон, і Уззіїл.
1CHR|6|19|(6-4) Сини Мерарієві: Махлі та Муші. А оце Левієві роди за їхніми батьками:
1CHR|6|20|(6-5) у Ґершома: Лівні його син, син його Яхат, його син Зімма,
1CHR|6|21|(6-6) його син Йоах, його син Іддо, його син Зерах, його син Єатрай.
1CHR|6|22|(6-7) Сини Кегатові: Аммінадав син його, його син Корах, син його Ассір,
1CHR|6|23|(6-8) син його Елкана, син його Ев'ясаф, син його Ассір,
1CHR|6|24|(6-9) син його Тахат, син його Уріїл, син його Уззійя та Саул син його.
1CHR|6|25|(6-10) А сини Елкани: Амасай та Ахімот.
1CHR|6|26|(6-11) Елкана його син, Цофай син його, і Нахат син його,
1CHR|6|27|(6-12) Еліяв син його, Єрохам син його, Елкана син його.
1CHR|6|28|(6-13) А Самуїлові сини: первороджений Йоїл, а другий Авійя.
1CHR|6|29|(6-14) Сини Мерарієві: Махлі, його син Лівні, його син Шім'ї, його син Узза,
1CHR|6|30|(6-15) син його Шім'а, син його Хаґґійя, син його Асая.
1CHR|6|31|(6-16) А оце ті, яких Давид поставив для співання в Господньому домі, від часу миру ковчега.
1CHR|6|32|(6-17) І вони служили перед скинією, скинією заповіту, піснею, аж поки Соломон не збудував Господнього дому в Єрусалимі. І вони ставали, за уставом своїм, на свою службу.
1CHR|6|33|(6-18) А оце ті, що стояли, та їхні сини: співак Геман, син Йоїла, сина Самуїла,
1CHR|6|34|(6-19) сина Елкани, сина Єрохама, сина Еліїла, сина Тоаха,
1CHR|6|35|(6-20) сина Цуфа, сина Елкани, сина Махата, сина Амасая,
1CHR|6|36|(6-21) сина Елкани, сина Йоїла, сина Азарії, сина Цефанії,
1CHR|6|37|(6-22) сина Тахата, сина Ассіра, сина Ев'ясафа, сина Кораха,
1CHR|6|38|(6-23) сина Їцхара, сина Кегата, сина Леві, сина Ізраїля.
1CHR|6|39|(6-24) А брат його Асаф, що стояв на правиці його: Асаф був сином Берехії, сина Шім'ї,
1CHR|6|40|(6-25) сина Михаїла, сина Баасеї, сина Малкійї,
1CHR|6|41|(6-26) сина Етні, сина Зераха, сина Адаї,
1CHR|6|42|(6-27) сина Етана, сина Зіммі, сина Шім'ї,
1CHR|6|43|(6-28) сина Йахата, сина Ґершома, сина Леві.
1CHR|6|44|(6-29) А сини Мерарі, брати їхні на лівиці: Етам, син Кіші, сина Авді, сина Маллуха,
1CHR|6|45|(6-30) сина Хашав'ї, сина Амації, сина Хілкійї,
1CHR|6|46|(6-31) сина Амці, сина Бані, сина Шамері
1CHR|6|47|(6-32) сина Махті, сина Муші, сина Мерарі, сина Леві.
1CHR|6|48|(6-33) А брати їх Левити дані на всяку роботу скинії Божого дому.
1CHR|6|49|(6-34) А Аарон та сини його палили на жертівнику цілопалення та на кадильному жертівнику, і були на всяку роботу Святого Святих, та на очищення Ізраїля, згідно зо всім тим, що наказав був Мойсей, раб Божий.
1CHR|6|50|(6-35) А оце Ааронові сини: Елеазар син його, його син Пінхас, його син Авішуя,
1CHR|6|51|(6-36) його син Буккі, його син Уззі, його син Зерахія,
1CHR|6|52|(6-37) його син Мерайот, його син Амарія, його син Ахітув,
1CHR|6|53|(6-38) його син Садок, його син Ахімаац.
1CHR|6|54|(6-39) А оце місце їхнього сидіння за їхніми осадами, в їхніх границях, синам Аароновим, з роду Кегатівців, бо для них був такий жеребок.
1CHR|6|55|(6-40) І дали їм Хеврон в Юдиному краї, та пасовиська його навколо нього.
1CHR|6|56|(6-41) А міське поле та осади його дали Калеву, синові Ефунне.
1CHR|6|57|(6-42) А Аароновим синам дали міста сховища: Хеврон, і Лівну та її пасовиська, і Яттір, і Ештемоа та пасовиська його,
1CHR|6|58|(6-43) і Хілен та пасовиська його, Девір та пасовиська його,
1CHR|6|59|(6-44) і Ашон та пасовиська його, і Бет-Шемеш та пасовиська його.
1CHR|6|60|(6-45) А з племени Веніяминового: Ґеву та пасовиська її, і Алемет та пасовиська його, і Анатот та пасовиська його, усіх їхніх міст в їхніх родах тринадцять міст.
1CHR|6|61|(6-46) А Кегатовим синам, позосталим із роду племени, дано з половини племени, племени Манасіїного, жеребком десять міст.
1CHR|6|62|(6-47) А Ґершомовим синам, за їхніми родами, з племени Іссахарового, і з племени Асирового, і з племени Нефталимового, і з племени Манасіїного в Башані дано тринадцять міст.
1CHR|6|63|(6-48) Синам Мерарієвим за родами їх із племени Рувимового, і з племени Ґадового, і з племени Завулонового дано за жеребком дванадцять міст.
1CHR|6|64|(6-49) І дали Ізраїлеві сини Левитам ті міста та їхні пасовиська.
1CHR|6|65|(6-50) Вони дали жеребком із племени Юдиних синів, і з племени Симеонових синів, і з племени Веніяминових синів ті міста, що їх вони назвали іменами.
1CHR|6|66|(6-51) А щодо тих, що з родів Кегатових синів, то міста границь їх були від Єфремового племени.
1CHR|6|67|(6-52) І дали їм міста сховища: Сихем та пасовиська його, в Єфремових горах, і Ґезер та пасовиська його,
1CHR|6|68|(6-53) і Йокмеам та пасовиська його, і Бет-Хорон та пасовиська його,
1CHR|6|69|(6-54) і Айялон та пасовиська його, і Ґат-Ріммон та пасовиська його.
1CHR|6|70|(6-55) А з половини Манасіїного племени: Анер та пасовиська його, і Біл'ам та пасовиська його, за родами позосталих Кегатових синів.
1CHR|6|71|(6-56) Ґершомовим синам із роду половини Манасіїного племени: Ґолан у Башані та пасовиська його, і Аштарот та пасовиська його.
1CHR|6|72|(6-57) А з Іссахарового племени: Кедеш та пасовиська його, і Доврат та пасовиська його,
1CHR|6|73|(6-58) і Рамот та пасовиська його, і Анем та пасовиська його.
1CHR|6|74|(6-59) А з Асирового племени: Машал та пасовиська його, і Авдон та пасовиська його,
1CHR|6|75|(6-60) і Хукок та пасовиська його, і Рехов та пасовиська його.
1CHR|6|76|(6-61) А з племени Нефталимового: Кедеш у Ґалілі та пасовиська його, і Хаммон та пасовиська його, і Кір'ятаїм та пасовиська його.
1CHR|6|77|(6-62) А позосталим Мерарієвим синам із Завулонового племени: Ріммон та пасовиська його, Фавор та пасовиська його.
1CHR|6|78|(6-63) А з другого боку Йордану при Єрихоні, на схід від Йордану, з Рувимового племени: Бецер на пустині та пасовиська його, і Ягца та пасовиська її,
1CHR|6|79|(6-64) і Кедемот та пасовиська його, і Мефаат та пасовиська його.
1CHR|6|80|(6-65) А з Ґадового племени: Рамот у Ґілеаді та пасовиська його, і Маханаїм та пасовиська його,
1CHR|6|81|(6-66) і Хешбон та пасовиська його, і Яазір та пасовиська його.
1CHR|7|1|А Іссахарові сини: Тола, і Пуа, Яшув і Шімрон, четверо.
1CHR|7|2|А Толині сини: Уззі, і Рефая, і Єріїл, і Яхмай, і Ївсам, і Самуїл, голови їхніх батьківських домів Толи, хоробрі вояки своїх родів. Число їх за Давидових днів двадцять і дві тисячі і шість сотень.
1CHR|7|3|А сини Уззі: Їзрахія. А сини Їзрахії: Михаїл, і Овадія, і Йоїл, Їшшійя, п'ятеро, вони всі голови.
1CHR|7|4|А в них, за їхніми нащадками, за домом їхніх батьків, були бойові військові ватаги, тридцять і шість тисяч, бо вони мали багато жінок та синів.
1CHR|7|5|А їхніх братів по всіх Іссахарових родах, хоробрих вояків, було вісімдесят і сім тисяч, усі вони переписані.
1CHR|7|6|Веніямин: Бела, і Бекер, і Єдіяїл, троє.
1CHR|7|7|А сини Белині: Ецбон, і Уззі, і Уззіїл, і Єрімот, і Ірі, п'ятеро голів батьківських домів, хоробрі вояки. А в родоводах їх двадцять і дві тисячі тридцять і чотири.
1CHR|7|8|А сини Бехерові: Земіра, і Йоаш, і Еліезер, і Елйоенай, і Омрі, і Єремот, і Авійя, і Анатот, і Алемет, усе це Бехерові сини.
1CHR|7|9|А в родоводах їх, за їхніми нащадками, головами дому їхніх батьків, хоробрих вояків, двадцять тисяч і двісті.
1CHR|7|10|А сини Єдіяїлові: Білган. А сини Білганові: Єуш, і Веніямин, і Егуд, і Кенаана, і Зетан, і Таршіш, і Ахішахар.
1CHR|7|11|Усіх цих Едіяїлових синів, за головами дому батьків, хоробрих вояків, було сімнадцять тисяч і двісті, що виходили з військовим відділом на війну.
1CHR|7|12|І Шуппім, і Хуппім, сини Іра, Хушім син Ахера.
1CHR|7|13|Сини Нефталимові: Яхціїл, і Ґуні, і Єцер, і Шаллум, сини Білги.
1CHR|7|14|Сини Манасіїні: Асріїл, якого породила його наложниця арамітка; вона породила й Махіра, Ґілеадового батька.
1CHR|7|15|А Махір узяв жінку для Хуппіма та Шуппіма, а ім'я його сестрі Мааха, а ім'я другому Целофхад. А в Целофхада були тільки дочки.
1CHR|7|16|І породила Мааха, Махірова жінка, сина, і назвала ім'я йому Переш, а ім'я братові його Шареш. А його сини Улам і Рекем.
1CHR|7|17|А Уламові сини: Бедан. Оце сини Ґілеада, сина Махіра, сина Манасіїного.
1CHR|7|18|А сестра його Молехет породила Ішгода, і Авіезера, і Махлу.
1CHR|7|19|А сини Шеміди були: Ахіян, і Шехем, і Лікхі, і Аніям.
1CHR|7|20|А сини Єфремові: Шутелах, і Веред, син його, і син його Тахат, і син його Ел'ада, і син його Тахат,
1CHR|7|21|і син його Завад, і син його Шутелах, і Езер, і Ел'ад. І повбивали їх люди Ґату, народжені в Краю, бо вони зійшли були забрати їхні череди.
1CHR|7|22|І був у жалобі їх батько Єфрем численні дні, а брати його приходили розважати його.
1CHR|7|23|І ввійшов він до жінки своєї, і зачала вона, і породила сина, а він назвав ім'я йому: Берія, бо зло було в домі його.
1CHR|7|24|А дочка його Шеера. І вона збудувала Бет-Хорон долішній і горішній та Уззен-Шееру.
1CHR|7|25|І син його Рефах, і Решеф, і син його Телах, і син його Тахан,
1CHR|7|26|син його Ладан, син його Аммігуд, син його Елішама,
1CHR|7|27|син його Нон, син його Ісус.
1CHR|7|28|А їхня посілість та місця їхнього оселення Бет-Ел та належні йому міста, а на схід Нааран, а на захід Ґезер та належні йому міста, і Сихем та належні йому міста, аж до Айї та належних йому міст.
1CHR|7|29|А на руки Манасіїних синів: Бет-Шеан та належні йому міста, Танах та належні йому міста, Меґіддо та належні йому міста, Дор та належні йому міста, у них сиділи сини Йосипа, Ізраїлевого сина.
1CHR|7|30|Сини Асирові: Їмна, і Їшва, і Їшві, і Берія, та сестра їх Серах.
1CHR|7|31|А сини Беріїні: Хевер і Малкіїл, він батько Бірзаіта.
1CHR|7|32|А Хевер породив Яфлета, і Шомера, і Хотама, і сестру їх Шую.
1CHR|7|33|А сини Яфлетові: Пасах, і Бімхал, і Ашват, оце сини Яфлетові.
1CHR|7|34|А сини Шемерові: Ахі і Рогаґґа, Яхебба та Арам.
1CHR|7|35|А сини Гелема, його брата: Цофах, і Їмна, і Шелеш, і Амал.
1CHR|7|36|Сини Цофахові: Суах, і Харнефер, і Шуал, і Бері, і Їмра,
1CHR|7|37|Бецер, і Год, і Шамма, і Шілша, і Їтран, і Беера.
1CHR|7|38|А сини Єтерові: Єфунне, і Піспа, і Ара.
1CHR|7|39|А сини Улли: Арах, і Ханніїл, і Ріція.
1CHR|7|40|Усе це Асирові сини, голови батьківських домів, вибрані лицарі вояки, голови начальників. А в родовідних книгах військових записано, число їхніх людей було двадцять і шість тисяч.
1CHR|8|1|А Веніямин породив первородженого свого Белу, другого Ашбелу, і третього Ахраха,
1CHR|8|2|четвертого Наху, і п'ятого Рафу.
1CHR|8|3|А в Бели були сини: Аддар, і Ґера, і Авігуд,
1CHR|8|4|і Авішуя, і Нааман, і Ахоах,
1CHR|8|5|і Ґера, і Шефуфан, і Хурам.
1CHR|8|6|А оце сини Ехудові, вони були голови дому батьків, мешканців Ґеви, та переселено їх до Манахату:
1CHR|8|7|і Нааман, і Ахійя, і Ґера, він їх переселив, і породив Уззу та Ахіхуда.
1CHR|8|8|А Шахараїм породив дітей на моавському полі по тому, як він відіслав своїх жінок Хушім та Баару.
1CHR|8|9|І породив він від Ходеш, своєї жінки: Йовава, і Цівію, і Мешу, і Малкам,
1CHR|8|10|і Єуц, і Сохію, і Мірму, це сини його, голови батьківських домів.
1CHR|8|11|А від Хушім він породив Авітува та Елпаала.
1CHR|8|12|А сини Елпаалові: Евер, і Міш'ам, і Шемер, він збудував Оно й Лод та належні йому міста.
1CHR|8|13|А Берія та Шема вони голови дому батьків, мешканців Айялону; вони вигнали мешканців Ґату.
1CHR|8|14|А Ахйо, Шашак і Єремот,
1CHR|8|15|і Зевадія, і Арад, і Адер,
1CHR|8|16|і Михаїл, і Їшпа, і Йоха сини Берії.
1CHR|8|17|А Зевадія, і Мешуллам, і Хізкі, і Хевер,
1CHR|8|18|і Їшмерай, і Їзлія, і Йовав, сини Елпаалові.
1CHR|8|19|А Яким, і Зіхрі, і Завді,
1CHR|8|20|і Еліенай, і Ціллетай, і Еліїл,
1CHR|8|21|і Адая, і Берая, і Шімрат, сини Шімеієві.
1CHR|8|22|А Їшпан, і Евер, і Еліїл,
1CHR|8|23|і Авдон, і Зіхрі, і Ханан,
1CHR|8|24|і Хананія, і Елам, і Антотійя,
1CHR|8|25|і Їфдея, і Пенуїл, сини Шашакові.
1CHR|8|26|А Шамшерай, і Шехарія, і Аталія,
1CHR|8|27|і Яарешія, і Елійя, і Зіхрі, сини Єрохамові.
1CHR|8|28|Оце голови дому батьків за їхніми нащадками, голови, що вони сиділи в Єрусалимі.
1CHR|8|29|А в Ґів'оні сиділи: батько Ґів'ону, а ім'я його жінці Мааха,
1CHR|8|30|і первороджений син його Авдон, і Цур, і Кіш, і Баал, і Надав,
1CHR|8|31|і Ґедор, і Ахйо, і Зехер.
1CHR|8|32|А Міклот породив Шім'у. І вони теж сиділи в Єрусалимі, при братах своїх, зо своїми братами.
1CHR|8|33|А Нер породив Кіша. А Кіш породив Саула, а Саул породив Йонатана, і Малкі-Шуя, і Авінадава, і Ешбаала.
1CHR|8|34|А син Йонатанів Мерів-Баал, а Мерів-Баал породив Міху.
1CHR|8|35|А сини Міхи: Пітон, і Мелех, і Тареа, і Ахаз.
1CHR|8|36|А Ахаз породив Єгоадду, а Єгоадда породив Алемета, і Азмавета, і Зімрі: а Зімрі породив Моцу.
1CHR|8|37|А Моца породив Бін'ю, його син Рафа, його син Ел'аса, його син Ацел.
1CHR|8|38|А в Ацела було шестеро синів, а оце їхні імена: Азрікам, Бохеру, і Ізмаїл, і Шеар'я, і Овадія, і Ханан, усі вони сини Ацелові.
1CHR|8|39|А сини Ешека, брата його: первороджений його Улам, другий Єуш, третій Еліфелет.
1CHR|8|40|А Уламові сини були мужі хоробрі вояки, що натягували лука й що мали багато синів та онуків, сотню й п'ятдесят. Усі вони з Веніяминових синів.
1CHR|9|1|А ввесь Ізраїль був переписаний, й ось вони були записані в книзі Ізраїлевих царів. А Юда був переселений до Вавилону за своє спроневірення.
1CHR|9|2|А перші мешканці, що сиділи в своїй посілості, по своїх містах, були: Ізраїль, священики, Левити та слуги храму.
1CHR|9|3|А в Єрусалимі сиділи з Юдиних синів, і з Веніяминових синів, і з синів Єфремових та Манасіїних:
1CHR|9|4|Утай, син Аммігуда, сина Омрі, сина Імрі, сина Бані, з синів Переца, Юдиного сина.
1CHR|9|5|А з шілонян: первороджений Асая та сини його.
1CHR|9|6|А з синів Зерахових: Єуїл, та брати їх, шість сотень і дев'ятдесят.
1CHR|9|7|А з синів Веніяминових: Саллу, син Мешуллама, сина Годавії, сина Сенуї,
1CHR|9|8|і Ївнея, син Єрохамів; і Ела, син Уззі, сина Міхрі, і Мешуллам, син Шефатії, сина Реуїла, сина Ївнійї,
1CHR|9|9|і брати їхні за їхніми нащадками, дев'ять сотень і п'ятдесят і шість. Усі ці мужі голови батьків, дому батьків своїх.
1CHR|9|10|А із священиків: Єдая, і Єгоярів, і Яхін.
1CHR|9|11|А Азарія, син Хілкійї, сина Мешуллама, сина Садока, сина Мерайота, сина Ахітава, управитель Божого дому;
1CHR|9|12|і Адая, син Єрохама, сина Пашхура, сина Малкійї; і Масай, син Адіїла, сина Яхзери, сина Мешуллама, сина Мешіллеміта, сина Іммера;
1CHR|9|13|і брати їх, голови дому своїх батьків тисяча й сім сотень і шістдесят, дуже добрі мужі на працю в ділі Божого дому.
1CHR|9|14|А з Левитів: Шемая, син Хассува, сина Азрікама, сина Хашав'ї, з синів Мерарі;
1CHR|9|15|і Бакбаккар, Хереш, і Балал, і Маттанія, син Міхи, сина Зіхрі, сина Асафа;
1CHR|9|16|і Авадія, син Шемаї, сина Ґалала, сина Єдутуна; і Берехія, син Аси, сина Елкани, що сидів в осадах нетоф'ян.
1CHR|9|17|А придверні: Шаллум, і Аккув, і Талмон, і Ахіман, і брати їхні; Шаллум був голова.
1CHR|9|18|І аж дотепер вони в царській брамі на схід, вони придверні таборів Левієвих синів.
1CHR|9|19|А Шаллум, син Коре, сина Ев'ясафа, сина Кораха, і брати його з дому його батька, корахівці, на праці служби, стерегли пороги скинії, а їхні батьки були над Господнім табором, стерегли вхід.
1CHR|9|20|І Пінхас, син Елеазарів, був над ними колись зверхником, і Господь був із ним.
1CHR|9|21|Захарій, син Мешелемії, був придверний при вході скинії заповіту.
1CHR|9|22|Усіх їх, вибраних на придверних при порогах, було двісті й дванадцять. Вони переписані по своїх осадах. Їх поставив Давид та прозорливець Самуїл за їх вірність.
1CHR|9|23|І вони та їхні сини були при брамах Господнього дому, дому скинії, за вартами.
1CHR|9|24|На чотири боки були придверні: на схід, на захід, на північ, на південь.
1CHR|9|25|А брати їхні були по селах, мусіли приходити на сім день, від часу до часу, щоб бути з ними на службі,
1CHR|9|26|бо в службі були чотири перші придверні, вони Левити; вони ж доглядали помешкань та скарбів Божого дому.
1CHR|9|27|І вони всю ніч перебували навколо Божого дому, бо на них був обов'язок варти, і вона щоранку відмикали двері.
1CHR|9|28|І з них були дехто коло службового посуду, бо за числом його приносили, і за числом його виносили.
1CHR|9|29|І з них дехто були призначені до посуду та до всяких святих речей: і над пшеничною мукою, і над вином, і над оливою, і над ладаном, і над пахощами.
1CHR|9|30|А з священичих синів були ті, що мішали запашне на кадило.
1CHR|9|31|А Маттітія з Левитів, він первороджений корахівця Шаллума, був у службі над справою сковорід.
1CHR|9|32|А з синів кегатівців, з їхніх братів, були над хлібом показним, щоб приготовляти щосуботи.
1CHR|9|33|А оце співаки, голови батьківських домів Левитів, по кімнатах, були вільні від іншої праці, бо вдень та вночі були вони при своїй роботі.
1CHR|9|34|Оце голови батьківських домів Левитів за їхніми нащадками, голови, що сиділи в Єрусалимі.
1CHR|9|35|А в Ґів'оні сиділи: батько Ґів'ону Єіїл, а ім'я його жінці Мааха,
1CHR|9|36|і первороджений син його Авдон, і Цур, і Кіш, і Баал, і Нер, і Надав,
1CHR|9|37|і Ґедор, і Ахйо, і Захарій, і Міклот.
1CHR|9|38|А Міклот породив Шім'ама. І вони теж сиділи в Єрусалимі при братах своїх, зо своїми братами.
1CHR|9|39|А Нер породив Кіша, а Кіш породив Саула, а Саул породив Йонатана, і Малкі-Шую, і Авінадава, і Ешбаала.
1CHR|9|40|А син Йонатанів Мерів-Баал, а Мерів-Баал породив Міху.
1CHR|9|41|А сини Міхи: Пітон, і Мелех, і Тахрея.
1CHR|9|42|А Ахаз породив Яру, а Яра породив Алмета, і Азмавета, і Зімрі. А Зімрі породив Моцу.
1CHR|9|43|А Моца породив Бін'ю, його син Рефая, його син Ел'аса, його син Ацел.
1CHR|9|44|А в Ацела було шестеро синів, а оце їхні імена: Азрікам, Бохеру, і Ізмаїл, і Шеар'я, і Овадія, і Ханан, оце сини Ацелові.
1CHR|10|1|А филистимляни воювали з Ізраїлем. І побігли Ізраїлеві мужі перед филистимлянами, і падали трупами на горі Ґілбоа.
1CHR|10|2|І гналися филистимляни за Саулом та за його синами. І повбивали филистимляни Йонатана, і Авінадава, і Малкі-Шуя, Саулових синів...
1CHR|10|3|І став бій тяжкий для Саула, і лучники кинулися на нього, і він злякався тих лучників.
1CHR|10|4|І сказав Саул до свого зброєноші: Витягни меча свого, і пробий мене ним, щоб не прийшли ці необрізані, і не знущалися надо мною! Та не хотів зброєноша, бо дуже боявся. Тоді взяв Саул меча та й упав на нього...
1CHR|10|5|І побачив зброєноша, що помер Саул, і впав і він на меча, та й помер...
1CHR|10|6|І помер Саул і троє синів його, та ввесь його дім померли разом.
1CHR|10|7|І побачили всі ізраїльтяни, що мешкали в долині, що всі втікають, та що помер Саул та сини його, то покидали свої міста й повтікали, а филистимляни поприходили, й осілися в них...
1CHR|10|8|І сталося другого дня, і прийшли филистимляни, щоб пообдирати трупи, та й знайшли Саула та синів його, що лежали на горі Ґілбоа.
1CHR|10|9|І вони пообдирали його, і понесли голову його та зброю його, і послали в филистимські краї навколо, щоб сповістити в домах своїх божків та народові.
1CHR|10|10|І вони поклали зброю його в домі свого бога, а голову його прибили в домі Даґона.
1CHR|10|11|І почув увесь ґілеадський Явеш про все, що филистимляни зробили Саулові,
1CHR|10|12|і встали всі хоробрі, і понесли Саулове тіло та тіла синів його, і принесли до Явешу, та й поховали їхні кості під дубом в Явеші, і постили сім день.
1CHR|10|13|І помер Саул за своє беззаконня, що він ним спроневірився проти Господа через Господнє слово, якого не тримався, а також через те, що питався віщого духа, щоб вивідати,
1CHR|10|14|а не вивідував від Господа. І Він убив його, а царство його передав Давидові, Єссеєвому синові.
1CHR|11|1|І зібрався ввесь Ізраїль до Давида в Хеврон, говорячи: Оце ми кість твоя та тіло твоє!
1CHR|11|2|І давніш, коли Саул був царем, ти водив та приводив Ізраїля на війну. І сказав Господь, Бог твій, тобі: Ти будеш пасти народа Мого, Ізраїля, і ти будеш князем над народом Моїм, Ізраїлем.
1CHR|11|3|І прийшли всі Ізраїлеві старші в Хеврон, а Давид склав із ними умову в Хевроні перед Господнім лицем. І помазали вони Давида царем над Ізраїлем, за Господнім словом через Самуїла.
1CHR|11|4|І пішов Давид та ввесь Ізраїль до Єрусалиму, він Євус, і там були євусеяни, мешканці того краю.
1CHR|11|5|І сказали мешканці Євусу до Давида: Ти не ввійдеш сюди! Та здобув Давид твердиню Сіон, він Місто Давида.
1CHR|11|6|І сказав Давид: Кожен, хто найперше поб'є євусеянина, той стане за голову та за зверхника. І ввійшов найперше Йоав, син Церуїн, і став за голову.
1CHR|11|7|І осівся Давид у твердині, тому назвав ім'я їй: Давидове Місто.
1CHR|11|8|І він збудував місто навколо, від Мілло й аж навколо, а Йоав відновив решту міста.
1CHR|11|9|І Давид ставав усе більшим, а Господь Саваот був із ним.
1CHR|11|10|А оце голови Давидових лицарів, що хоробро трудилися з ним у його царстві, з усім Ізраїлем, щоб настановити його царем, за Господнім словом, над Ізраїлем.
1CHR|11|11|А оце число Давидових лицарів: Яшов'ам, син Гахмоні, голова тридцяти, він махнув своїм списом і побив за один раз три сотні!
1CHR|11|12|А за ним Елеазар, син Додо, ахох'янин, він один із трьох лицарів.
1CHR|11|13|Він був із Давидом у Пас-Дамімі, а филистимляни зібралися там на бій. І була там ділянка поля, повна ячменю, а народ утікав перед филистимлянами.
1CHR|11|14|Та вони стали посеред ділянки, і врятували її та й побили филистимлян. І Господь подав велику перемогу!
1CHR|11|15|І зійшли троє з тих тридцяти на переді на скелю до Давида, до печери Адуллам. А филистимський табір таборував у долині Рефаїм.
1CHR|11|16|Давид же був тоді в твердині, а филистимська залога була тоді в Віфлеємі.
1CHR|11|17|І спрагнув Давид та й сказав: Хто напоїть мене водою з віфлеємської криниці, що в брамі?
1CHR|11|18|І продерлися ці троє до филистимського табору, і зачерпнули води з віфлеємської криниці, що в брамі. І вони винесли й принесли до Давида, та Давид не схотів її пити, і вилив її для Господа,
1CHR|11|19|та й сказав: Борони мене, Боже мій, чинити таке! Чи я буду пити кров цих мужів, що ходили, наражаючи життя своє? Бо життям своїм вони принесли її! І не хотів він пити її. Оце зробили троє цих лицарів.
1CHR|11|20|А Авшай, Йоавів брат, він голова тих трьох. І він махнув своїм списом і побив три сотні! І він мав найславніше ім'я серед трьох.
1CHR|11|21|З тих трьох серед двох він був найшановніший, і став їм за провідника. А до тих трьох не досяг.
1CHR|11|22|Беная, син Єгоядин, син хороброго мужа, великий у ділах, з Кавцеїлу, він побив двох синів Аріїла моавського. І він зійшов і забив лева в середині ями сніжного дня.
1CHR|11|23|І він побив одного єгиптянина, мужа поставного, на п'ять ліктів, а в руці єгиптянина був спис, як ткацький вал. І зійшов він до нього з києм, і вирвав списа з руки того єгиптянина, та й його забив його списом.
1CHR|11|24|Оце зробив Беная, син Єгоядин, і його ім'я було серед тих трьох хоробрих.
1CHR|11|25|З тих тридцяти він був найповажніший, а до тих трьох не досяг. І Давид призначив його до своєї прибічної сторожі.
1CHR|11|26|А хоробрі мужі були ці: Асаїл, Йоавів брат, Елханан, син Додо, із Віфлеєму,
1CHR|11|27|гарор'янин Шаммот, пелонянин Хелес,
1CHR|11|28|Іра, син Іккешів, текоянин, антотянин Авіезер,
1CHR|11|29|хушатянин Сіббехай, ахох'янин Ілай,
1CHR|11|30|нетофатянин Магарай, Хелед, син Баанин, нетофатянин,
1CHR|11|31|Ітай, син Ріваїв, з Ґів'ї Веніяминової, пір'атонянин Беная,
1CHR|11|32|Хурай з Нахале-Ґаашу, арв'янин Авіїл,
1CHR|11|33|бахарум'янин Азмавет, шаалвонянин Ел'яхба,
1CHR|11|34|сини ґізонянина Гашема, Йонатан, син Шаґе, гарар'янин,
1CHR|11|35|Ахійям, син Сахарів, гарар'янин, Еліфал, син Урів,
1CHR|11|36|мехар'янин Хефер, пелонянин Ахійя,
1CHR|11|37|кармелянин Хіцро, Наарай, син Езлаїв,
1CHR|11|38|Йоїл, брат Натанів, Мівхар, син Ґаґрі,
1CHR|11|39|аммонітянин Целек, беротянин Нахрай, зброєноша Йоава, Церуїного сина,
1CHR|11|40|їтрянин Іра, їтрянин Ґарев,
1CHR|11|41|хіттеянин Урійя, Завад, син Ахлая,
1CHR|11|42|Адіна, син Шізин, Рувимівець, голова Рувимівців і над тридцятьма,
1CHR|11|43|Ханан, син Маахин, і мітнянин Йосафат,
1CHR|11|44|аштерянин Уззійя, Шама, і Еуїл, сини ароерянина Хотама,
1CHR|11|45|Єдіаїл, син Шімрі, і Йоха, його брат, тіцянин,
1CHR|11|46|махав'янин Еліїл, і Єрівай, і Йошав'я, сини Ел'наамові, і моавітянин Їтма,
1CHR|11|47|Етіїл, і Овед, і Яасіїл із Цови.
1CHR|12|1|А це ті, що поприходили до Давида в Ціклаґ, коли він ще ховався перед Саулом, сином Кішевим, і вони були серед лицарів, що допомагали в війні,
1CHR|12|2|що були озброєні луком, що кидали правицею та лівицею каміння та стріли з лука, з Саулових братів, від Веніямина:
1CHR|12|3|голова Ахіезер та Йоаш, сини ґів'янина Шемаї, і Єзіїл та Пелет, Азмаветові сини, і Бераха, і аннетотянин Єгу,
1CHR|12|4|і ґів'онянин Їшмая, лицар серед тридцятьох та старший над тридцятьма, і Їрмея, і Яхазіїл, і Йоханан, і ґедерянин Йозавад,
1CHR|12|5|Ел'узай, і Єрімот, і Беал'я, і Шемарія, і гаріф'янин Шефатія,
1CHR|12|6|Елкана, і Їшшійя, і Азареїл, і Йоезер, і Яхов'ам, хорх'яни,
1CHR|12|7|і Йоїла та Зевадія, сини Єрохамові, з Ґедору.
1CHR|12|8|А з ґадян відділилися до Давида до твердині в пустиню лицарі вояки, мужі відважні, на війні, озброєні великим щитом та списом. А їхні обличчя то обличчя лев'ячі, а щодо швидкости вони були, як сарни на горах.
1CHR|12|9|Голова Езер, другий Овадія, третій Еліав,
1CHR|12|10|четвертий Мішманна, п'ятий Їрмея,
1CHR|12|11|шостий Аттай, сьомий Еліїл,
1CHR|12|12|восьмий Йоханан, дев'ятий Елзавад,
1CHR|12|13|десятий Єремія, одинадцятий Махбанай.
1CHR|12|14|Оці були з Ґадових синів, голови військових відділів, малий один на сотню, а великий на тисячу.
1CHR|12|15|Це ті, що перейшли Йордан першого місяця, коли він був переповнений понад усі береги свої, і порозганяли всіх мешканців долин на схід та на захід.
1CHR|12|16|І прийшли з синів Веніяминових та Юдиних аж до твердині до Давида.
1CHR|12|17|А Давид вийшов перед них, і, відповідаючи, сказав їм: Якщо ви прийшли до мене з миром, щоб допомагати мені, буде моє серце з вами за одне, а якщо зрадите мене супроти ворогів моїх, коли нема обмани в руках моїх, то побачить це Бог наших батьків, і покарає!
1CHR|12|18|І зійшов Дух на Амасая, голову тридцяти, і він проказав: Мир, Давиде, тобі, і з тобою, о сину Єссеїв! Мир тобі, і мир тому, хто тобі помагає, бо тобі помагає твій Бог! І прийняв їх Давид, і поставив на чолі війська.
1CHR|12|19|І з Манасії перебігли до Давида, коли він ішов із филистимлянами проти Саула на війну, а він не поміг їм, бо филистимські князі, порадившись, відіслали його, говорячи: За ціну наших голів він хоче перейти до свого пана Саула!
1CHR|12|20|Коли він ішов до Ціклаґу, збігли до нього з Манасії: Аднах, і Йозавад, і Єдіаїл, і Михаїл, і Йозавад, і Елігу, і Ціллетай, голови Манасіїних тисячок.
1CHR|12|21|І вони допомагали Давидові проти юрби, бо вони всі хоробрі вояки, і поставали провідниками військових відділів.
1CHR|12|22|Бо день-у-день приходили вони до Давида помагати йому, аж став табір великий, як табір Божий.
1CHR|12|23|А оце число головних озброєних військових відділів, вони прийшли до Давида в Хеврон, щоб передати Саулове царство йому, за Господнім словом:
1CHR|12|24|Юдиних синів, що носили великого щита та списа, шість тисяч і вісім сотень озброєного війська.
1CHR|12|25|З Симеонових синів хоробрих вояків військового відділу сім тисяч і сто.
1CHR|12|26|З Левієвих синів чотири тисячі й шість сотень.
1CHR|12|27|І Єгояда, проводир синів Ааронових, а з ним три тисячі й сім сотень.
1CHR|12|28|І юнак Садок, хоробрий вояк, та дім його батька, зверхників двадцять і два.
1CHR|12|29|А з Веніяминових синів, Саулових братів, три тисячі, а більша частина їх аж дотепер трималися Саулового дому.
1CHR|12|30|А з Єфремових синів двадцять тисяч і вісім сотень хоробрих вояків, мужів славних дому їхніх батьків.
1CHR|12|31|А з половини Манасіїного племени вісімнадцять тисяч, що були докладно зазначені за іменем, щоб прийти настановити Давида царем.
1CHR|12|32|А з Іссахарових синів, що мали розуміння часу, щоб знати, що буде робити Ізраїль, їх голів було двісті, а всі їхні брати робили за їхнім наказом.
1CHR|12|33|Із Завулона тих, що виходять на війну, що ставляться в бойовому порядку зо всякими військовими речами, п'ятдесят тисяч, щоб допомагати з цілим серцем.
1CHR|12|34|А з Нефталиму тисяча зверхників, а при них зо щитом та списом тридцять і сім тисяч.
1CHR|12|35|А з Данян тих, що ставляться в бойовому порядку двадцять і вісім тисяч і шість сотень.
1CHR|12|36|А з Асира тих, що виходять на війну, щоб ставитися в бойовім порядку, сорок тисяч.
1CHR|12|37|А з того боку Йордану з Рувимівців, і Ґадівців, і з половини Манасії, зо всякими військовими знаряддями для бою сто й двадцять тисяч.
1CHR|12|38|Усі ці люди військові, що ставилися в бойовому порядку, цілим серцем поприходили до Хеврону, щоб настановити Давида царем над усім Ізраїлем. Та й решта Ізраїля були односерді, щоб настановити Давида царем.
1CHR|12|39|І були вони там із Давидом три дні, їли та пили, бо їхні брати наготовили їм.
1CHR|12|40|А також ті, що були близькі до них, аж до Іссахара, і Завулона, і Нефталима, спроваджували хліб ослами, і верблюдами, і мулами, і худобою великою, їжу мучну, спресовані фіґі, і родзинки, і вино, і оливу, і худобу велику, і худобу дрібну, дуже багато, бо радість була в Ізраїлі.
1CHR|13|1|І радився Давид із тисячниками та з сотниками, зо всіма значними.
1CHR|13|2|І сказав Давид до всієї Ізраїлевої громади: Якщо вам це добре, а від Господа, Бога нашого вподобане, пошлімо до наших братів, позосталих по всіх Ізраїлевих краях, а з ними до священиків та Левитів, по містах та по їхніх пасовиськах, і нехай зберуться до нас.
1CHR|13|3|І вернімо ковчега нашого Бога до нас, бо не зверталися ми до нього за Саулових днів.
1CHR|13|4|І сказала вся громада, щоб зробити так, бо слушна була та річ в очах усього народу.
1CHR|13|5|І зібрав Давид усього Ізраїля від єгипетського Шіхору й аж туди, де йдеться до Хамату, щоб спровадити Божого ковчега з Кір'ят-Єаріму.
1CHR|13|6|І пішов Давид та ввесь Ізраїль у Баалу, в Юдин Кір'ят-Єарім, щоб винести звідти ковчега Бога, Господа, що сидить на херувимах, що ім'я Його прикликається.
1CHR|13|7|І повезли Божого ковчега на новому возі з Авінадавового дому, а Узза та Ахйо провадили того воза.
1CHR|13|8|А Давид та ввесь Ізраїль грали перед Божим лицем з усієї сили, і з піснями, і на цитрах, і на арфах, і на бубнах, і на цимбалах, і на сурмах.
1CHR|13|9|І прийшли вони аж до Кідонового току, і простяг Узза свою руку, щоб підхопити ковчега, бо воли нахилили його.
1CHR|13|10|І запалився на Уззу гнів Господній, і Він убив його за те, що простяг руку свою до ковчега. І помер він там перед Господнім лицем...
1CHR|13|11|І зажурився Давид тим, що Господь убив Уззу, і він назвав ім'я тому місцю: Перец-Узза, і так воно зветься аж до цього дня.
1CHR|13|12|І того дня Давид злякався Бога, говорячи: Як я внесу до себе Божого ковчега?
1CHR|13|13|І не повіз Давид ковчега до себе, до Давидового Міста, а направив його до дому ґатянина Овед-Едома.
1CHR|13|14|І пробував Божий ковчег із домом Овед-Едома в його домі три місяці. А Господь поблагословив дім Овед-Едома, та все, що було його.
1CHR|14|1|А Хірам, цар тирський, послав до Давида послів, і кедрового дерева, каменярів та теслярів, щоб збудувати йому дім.
1CHR|14|2|І пізнав Давид, що Господь міцно поставив його царем над Ізраїлем, бо царство його було піднесене високо ради народу його, Ізраїля.
1CHR|14|3|І взяв Давид іще жінок в Єрусалимі, і Давид породив іще синів та дочок.
1CHR|14|4|А оце імена народжених йому в Єрусалимі: Шаммуа і Шовав, Натан і Соломон,
1CHR|14|5|і Ївхар, і Елішуя, і Елпелет,
1CHR|14|6|і Ноґах, і Нефеґ, і Яфія,
1CHR|14|7|і Елішама, і Ел'яда, і Еліфелет.
1CHR|14|8|І почули филистимляни, що Давид був помазаний на царя над усім Ізраїлем, і піднялися всі филистимляни, щоб шукати Давида. А Давид почув про це, і вийшов проти них.
1CHR|14|9|А филистимляни прийшли й стали таборами в долині Рефаїм.
1CHR|14|10|І питався Давид у Бога, говорячи: Чи виходити на филистимлян, і чи даси Ти їх в руку мою? І відказав йому Господь: Вийди, і Я дам їх у руку твою.
1CHR|14|11|І зійшли вони до Баал-Пераціму, і Давид побив їх там. І сказав Давид: Розбив Бог ворогів моїх рукою моєю, як прорив води! Тому назвали ім'я того місця: Баал-Перацім!
1CHR|14|12|А вони позоставили там богів своїх, і Давид наказав, і вони були спалені в огні.
1CHR|14|13|А филистимляни ще отаборилися в долині.
1CHR|14|14|А Давид іще питався Бога, і Бог йому сказав: Не підеш за ними, а поверни від них, і прибудеш до них з-навпроти бальзамового ліска.
1CHR|14|15|І станеться, як ти почуєш шелест ніби кроків на верховіттях бальзамових дерев, тоді вийдеш на бій, бо то вийшов Бог перед тебе, щоб побити филистимський табір.
1CHR|14|16|І зробив Давид так, як наказав йому Бог, і вони побили филистимський табір від Ґів'ону аж до Ґезеру.
1CHR|14|17|І неслося Давидове ім'я по всіх краях, а Господь дав, що всі народи боялись його.
1CHR|15|1|І поробив він собі доми в Давидовому Місті, і приготовив місце на Божого ковчега, і розтягнув для нього скинію.
1CHR|15|2|Тоді Давид сказав, щоб ніхто не носив Божого ковчега, окрім Левитів, бо їх вибрав Господь носити ковчега Господа та служити Йому аж навіки.
1CHR|15|3|І Давид зібрав усього Ізраїля до Єрусалиму, щоб винести Господнього ковчега на його місце, яке приготовив йому він.
1CHR|15|4|І зібрав Давид Ааронових синів та Левитів.
1CHR|15|5|Від Кегатових синів: зверхник Уріїл, а братів його сотня й двадцять.
1CHR|15|6|Від синів Мерарі: зверхник Асая, а братів його двісті й двадцять.
1CHR|15|7|Від Ґершомових синів: зверхник Йоїл, а братів його сотня й тридцять.
1CHR|15|8|Від Еліцафанових синів: зверхник Шемая, а братів його двісті.
1CHR|15|9|Від Хевронових синів: зверхник Еліїл, а братів його вісімдесят.
1CHR|15|10|Від Уззіїлових синів: зверхник Аммінадав, а братів його сотня й дванадцять.
1CHR|15|11|І покликав Давид священиків Садока та Евіятара, та Левитів: Уріїла, Асаю, і Йоїла, Шемаю і Еліїла, і Аммінадава
1CHR|15|12|та й сказав до них: Ви голови родів Левитів. Освятіться ви та ваші брати, і перенесете ковчега Господа, Бога Ізраїлевого, до місця, яке приготовив я йому.
1CHR|15|13|Бо через те, що спочатку не ви це робили, то вдарив нас Господь, Бог наш, бо ми не шукали Його так, як належало.
1CHR|15|14|І освятилися священики та Левити, щоб перенести ковчега Господа, Бога Ізраїлевого.
1CHR|15|15|І понесли сини Левитів Божого ковчега, як наказав був Мойсей за Господнім словом, на плечах своїх, на держаках, на собі.
1CHR|15|16|І сказав Давид зверхникам Левитів, щоб поставили своїх братів співаків на приладдях пісні, на цитрах, арфах, та тих, що грають на цимбалах, щоб піднести голос на радість.
1CHR|15|17|І поставили Левити Гемана, Йоїлового сина, а з братів його Асафа, сина Берехії, а з синів Мерарі, їхніх братів Етана, сина Кушаї.
1CHR|15|18|А з ними їхніх братів других: Захарія, і Яазіїла, і Шемірамота, і Єхіїла, і Унні, Еліава, і Бенаю, і Маасею, і Маттітію, і Еліфлея, і Мікнею, і Овед-Едома, і Єіїла, придверних.
1CHR|15|19|А співаків: Гемана, Асафа та Етана грати на мідяних цимбалах.
1CHR|15|20|А Захарія, і Азіїла, і Шемірамота, і Єхіїла, і Унні, і Еліава, і Маасею, і Бенаю на цитрах, на аламот.
1CHR|15|21|А Маттітію, і Еліфелегу, і Мікнею, і Овед-Едома, і Єїла, і Азазію на арфах, на октаві, щоб починати гру.
1CHR|15|22|А Кенанію, зверхника Левитів, над ношенням; він навчав носити, бо вмів того.
1CHR|15|23|А Берехія та Елкана придверні при ковчезі.
1CHR|15|24|А Шеванія, І Йосафат, і Натанаїл, і Амасай, і Захарій, і Беная, і Еліезер, священики, сурмили в сурми перед Божим ковчегом, а Овед-Едом та Єхійя придверні для ковчега.
1CHR|15|25|І пішов Давид і Ізраїлеві старші та тисячники, щоб перенести ковчега Господнього заповіту з Овед-Едомового дому з радістю.
1CHR|15|26|І сталося, коли Бог допомагав Левитам, що несли ковчега Господнього заповіту, то вони принесли в жертву сім биків та сім баранів.
1CHR|15|27|А Давид був зодягнений в одежу з вісону, як і всі Левити, що несли ковчега, і співаки, і Кенанія, зверхник ношення і співаків, а на Давиді був ще й льняний ефод.
1CHR|15|28|І ввесь Ізраїль ніс ковчега Господнього заповіту з радісним криком, і зо звуком рога, і з сурмами, і з цимбалами, граючи на цитрах та на арфах.
1CHR|15|29|І сталося, коли ковчег Господнього заповіту прийшов аж до Давидового Міста, то Мелхола, Саулова дочка, виглядала через вікно. І побачила вона царя Давида, що танцював та грав, і зневажила його в своєму серці.
1CHR|16|1|І принесли вони Божого ковчега, і поставили його в середині скинії, що розтягнув для нього Давид, і принесли цілопалення та мирні жертви перед Божим лицем.
1CHR|16|2|І покінчив Давид приносити цілопалення та мирні жертви, та й поблагословив народ Ім'ям Господнім.
1CHR|16|3|І він поділив для всякого Ізраїлевого мужа, від чоловіка й аж до жінки, кожному по буханцеві хліба, і по кавалкові м'яса та по виноградному калачеві.
1CHR|16|4|І він попризначував перед Господнім ковчегом із Левитів служачих, щоб вони визнавали, і прославляли, і хвалили Господа, Бога Ізраїлевого:
1CHR|16|5|Асаф був головою, а другий по ньому Захарій, Єіїл, і Шемірамот, і Хіїл, і Маттітія, і Еліяв, і Беная, і Овед-Едом, і Єіїл на знаряддях цитр та на арфах, а Асаф голосно грав на цимбалах.
1CHR|16|6|А священики Беная та Яхазіїл на сурмах, завжди перед ковчегом Божого заповіту.
1CHR|16|7|Того дня, тоді Давид дав уперше псалма на подяку Господеві через Асафа та братів його:
1CHR|16|8|Дякуйте Господу, кличте Ім'я Його, серед народів звіщайте про вчинки Його!
1CHR|16|9|Співайте Йому, грайте Йому, говоріть про всі чуда Його!
1CHR|16|10|Хваліться святим Його Йменням, хай тішиться серце шукаючих Господа!
1CHR|16|11|Пошукуйте Господа й силу Його, лице Його завжди шукайте!
1CHR|16|12|Пам'ятайте про чуда Його, які Він учинив, про ознаки Його та про присуди уст Його
1CHR|16|13|ви, насіння Ізраїля, раба Його, сини Яковові, вибранці Його!
1CHR|16|14|Він Господь, Бог наш, по цілій землі Його присуди!
1CHR|16|15|Пам'ятайте навіки Його заповіта, слово, яке наказав Він на тисячу родів,
1CHR|16|16|що склав Він Його з Авраамом, і присягу Його для Ісака.
1CHR|16|17|І Він поставив його за Закона для Якова, Ізраїлеві заповітом навіки,
1CHR|16|18|говорячи: Дам тобі край ханаанський, як наділ спадщини для вас!
1CHR|16|19|Тоді їх було невелике число, нечисленні були та приходьки на іншій землі,
1CHR|16|20|і від народу ходили вони до народу, і від царства до іншого люду.
1CHR|16|21|Не дозволив нікому Він кривдити їх, і за них Він царям докоряв:
1CHR|16|22|Не доторкуйтеся до Моїх помазанців, а пророкам Моїм не робіте лихого!
1CHR|16|23|Господеві співайте, вся земле, з дня-на-день сповіщайте спасіння Його!
1CHR|16|24|Розповідайте про славу Його між поганами, про чуда Його між усіма народами.
1CHR|16|25|Бо великий Господь і прославлений вельми, і Він найгрізніший над богів усіх!
1CHR|16|26|Бо всі боги народів божки, а Господь небеса сотворив!
1CHR|16|27|Слава та велич перед лицем Його, сила та радість на місці Його.
1CHR|16|28|Дайте Господу, роди народів, дайте Господу славу та силу,
1CHR|16|29|дайте Господу славу Ймення Його, приносьте дарунка й приходьте перед лице Його! Кланяйтеся Господеві в величчі святому!
1CHR|16|30|Перед лицем Його затремти, уся земле, бо міцно поставлений всесвіт, щоб не захитався!
1CHR|16|31|Хай небо радіє, і хай веселиться земля, і хай серед народів говорять: Царює Господь!
1CHR|16|32|Нехай гримить море й його повнота, нехай поле радіє та все, що на ньому!
1CHR|16|33|Тоді перед Господнім лицем дерева лісні заспівають, бо землю судити йде Він.
1CHR|16|34|Дякуйте Господу, добрий бо Він, бо навіки Його милосердя!
1CHR|16|35|І промовте: Спаси нас, о Боже спасіння нашого, і збери нас, і нас урятуй від народів, щоб дякувати Йменню святому Твоєму, щоб Твоєю хвалитися славою!
1CHR|16|36|Благословенний Господь, Бог Ізраїлів, від віку й навіки! А народ увесь сказав: Амінь і Хвала Господеві!
1CHR|16|37|І Давид позоставив там перед ковчегом Господнього заповіту Асафа та братів його, щоб завжди служили перед ковчегом, що в якій день треба було,
1CHR|16|38|і Овед-Едома та братів його, шістдесят і вісьмох; а Овед-Едома, Єдутунового сина, та Хоса за придверних;
1CHR|16|39|а священика Садока та братів його священиків перед Господнім наметом на пагірку, що в Ґів'оні,
1CHR|16|40|щоб приносити цілопалення для Господа на жертівнику цілопалення, завжди ранком та ввечорі, та на все інше, що написане в Законі Господа, що наказав був Ізраїлеві.
1CHR|16|41|А з ними Геман та Єдутун, та решта вибраних, що були докладно зазначені поіменно, щоб Дякувати Господеві, бо навіки Його милосердя!
1CHR|16|42|А з ними сурми та цимбали для тих, що грають, та знаряддя для Божої пісні. А сини Єдутунові сторожі до брами.
1CHR|16|43|І порозходився ввесь народ, кожен до дому свого. А Давид вернувся, щоб поблагословити свій дім.
1CHR|17|1|І сталося, як Давид сидів був у домі своїм, то сказав Давид до пророка Натана: Ось я сиджу в кедровому домі, а ковчег Господнього заповіту під занавісами!...
1CHR|17|2|І сказав Натан до Давида: Зроби все, що в серці твоєму, бо Бог із тобою!
1CHR|17|3|І сталося тієї ночі, і було Боже слово до Натана, говорячи:
1CHR|17|4|Іди, і скажеш Моєму рабові Давидові: Так сказав Господь: Не ти збудуєш Мені цього храма на перебування.
1CHR|17|5|Бо Я не сидів у храмі від дня, коли вивів Ізраїля, аж до дня цього, і ходив від шатра до шатра, і від намету до намету.
1CHR|17|6|Скрізь, де тільки ходив Я між усім Ізраїлем, чи сказав Я хоч слово котрому з Ізраїлевих суддів, яким наказав Я пасти народа Мого: Чому ви не збудували Мені кедрового храма?
1CHR|17|7|А тепер так скажеш рабові Моєму Давидові: Так сказав Господь Саваот: Я взяв тебе з пасовиська від отари, щоб став ти володарем над Моїм народом, Ізраїлем.
1CHR|17|8|І був Я з тобою скрізь, де ти ходив, і винищив Я всіх ворогів Твоїх перед тобою, і зробив Я тобі ім'я, як ім'я тих великих, що на землі.
1CHR|17|9|І дав Я місце Моєму народові Ізраїлеві, і посадив його так, що він перебуватиме на тому самому місці. І він уже не тремтітиме, а кривдники не будуть нищити його, як перше.
1CHR|17|10|А від днів, коли Я настановив суддів над Своїм народом, Ізраїлем, то понизив усіх ворогів твоїх. І звіщаю тобі, що Господь збудує тобі дім.
1CHR|17|11|І станеться, коли виповняться твої дні, щоб піти до батьків своїх, то Я поставлю по тобі твоє насіння, що буде з синів твоїх, і поставлю міцно його царство.
1CHR|17|12|Він збудує Мені храм, а Я поставлю його трона міцно аж навіки.
1CHR|17|13|Я буду йому за батька, а він буде Мені за сина, а милости Своєї Я не відійму від нього, як відняв Я від того, що був перед тобою.
1CHR|17|14|І поставлю його в храмі Своїм та в царстві Своїм аж навіки, і трон його буде міцно стояти навіки.
1CHR|17|15|За всіма цими словами, за всім цим видінням, так говорив Натан до Давида.
1CHR|17|16|І прийшов цар Давид, і сів перед Господнім лицем та й промовив: Хто я, Господи, Боже, і що таке дім мій, що Ти довів мене аж сюди?
1CHR|17|17|Та й це було мале в очах Твоїх, Боже, і Ти говорив про дім Свого раба на майбутнє, і Ти показав мені покоління людське, і підніс мене, Господи Боже!
1CHR|17|18|Що Давид додасть ще до Твого на вшанування Твого раба? А Ти Свого раба знаєш!
1CHR|17|19|Господи, ради Свого раба та за серцем Своїм зробив Ти все це велике, щоб завідомити про всі ті великі речі.
1CHR|17|20|Господи, нема Такого, як Ти, і нема Бога, окрім Тебе, за всім тим, що ми чули своїми ушима.
1CHR|17|21|І який є ще один люд на землі, як Твій народ, Ізраїль, щоб Бог приходив викупити його Собі за народа, і щоб установити Собі ймення великих та страшних речей, щоб вигнати народи перед народом Своїм, якого Ти викупив із Єгипту?
1CHR|17|22|І зробив Ти народ Свій, Ізраїля, Собі за народа аж навіки, і Ти, Господи, став йому за Бога!
1CHR|17|23|А тепер, Господи, нехай стане певним аж навіки те слово, яке говорив Ти про Свого раба, і зроби, як говорив!
1CHR|17|24|А Твоє Ім'я нехай буде міцне, і нехай буде велике аж навіки, щоб казали: Господь Саваот, Бог Ізраїлів Бог для Ізраїля, а дім Твого раба Давида поставлений міцно перед лицем Твоїм.
1CHR|17|25|Бо Ти, Боже мій, об'явив Своєму рабові, що Ти збудуєш йому дім, тому раб Твій знайшов потребу молитися перед лицем Твоїм.
1CHR|17|26|А тепер, Господи, Ти Той Бог, і сказав про Свого раба оце добре.
1CHR|17|27|А тепер був Ти ласкавий поблагословити дім Свого раба, щоб бути навіки перед лицем Твоїм, бо Ти, Господи, поблагословив, і він поблагословлений навіки!
1CHR|18|1|І сталося по тому, і побив Давид филистимлян та поконав їх; і взяв він Ґат та належні йому міста з руки филистимлян.
1CHR|18|2|І побив він Моава, і стали моавітяни Давидовими рабами, що приносили дари.
1CHR|18|3|І побив Давид Гадад'езера, царя цовського, в Хаматі, коли той ішов, щоб поставити владу свою на річці Ефраті.
1CHR|18|4|І здобув Давид від нього тисячі колесниць і сім тисяч верхівців та двадцять тисяч пішого люду. І попідрізував Давид жили коням усіх колесниць, і позоставив із них тільки сотню для колесниць.
1CHR|18|5|І прийшов Арам із Дамаску на поміч Гадад'езерові, цареві цовському, та Давид вибив серед сиріян двадцять і дві тисячі чоловіка.
1CHR|18|6|І поставив Давид у Сирії Дамаській залогу, і сиріяни стали для Давида рабами, що приносили дари. А Господь допомагав Давидові скрізь, де він ходив.
1CHR|18|7|І позабирав Давид золоті щити, що були на Гадад'езерових рабах, і позносив їх до Єрусалиму.
1CHR|18|8|А з Тівхату та з Куну, Гадад'езерових міст, позабирав Давид дуже багато міді, з неї поробив Соломон мідяне море й стовпи, та мідяні речі.
1CHR|18|9|І прочув Тоу, цар хамотський, що Давид побив усе військо Гадад'езера, царя цовського.
1CHR|18|10|І послав він сина свого Гадорама до царя Давида, щоб привітати його, та щоб поблагословити його за те, що воював із Гадад'езером та й побив його, бо Гадад'езер провадив війну з Тоу, а з ним послав всякі речі золоті, і срібні, і мідяні.
1CHR|18|11|І Давид присвятив їх Господеві разом із тим сріблом та золотом, що повиносив від усіх народів з Едому, і з Моаву, і від Аммонових синів та від Амалика.
1CHR|18|12|А Авшай, син Церуїн, побив Едома в Соляній долині, вісімнадцять тисяч.
1CHR|18|13|І поставив він в Едомі залогу, і став увесь Едом Давидовими рабами. А Господь допомагав Давидові скрізь, де він ходив.
1CHR|18|14|І царював Давид над усім Ізраїлем, і чинив суд та справедливість усьому своєму народові.
1CHR|18|15|А Йоав, син Церуїн, був над військом, а Йосафат, син Ахілудів, канцлер.
1CHR|18|16|А Садок, син Ахітувів, та Авімелех, син Ев'ятарів, були священики, а Шавша писар.
1CHR|18|17|А Беная, син Єгоядин, був над керетянином та над пелетянином, а Давидові сини перші при царевій руці.
1CHR|19|1|І сталося по тому, і помер Нахаш, цар аммонітський, а замість нього зацарював син його Ханун.
1CHR|19|2|І сказав Давид: Зроблю я милість Ханунові, Нахашевому синові, як батько його зробив був милість мені. І Давид послав послів, щоб потішити його за його батька. І прибули Давидові раби до аммонітського краю, до Хануна, щоб потішити його.
1CHR|19|3|А начальники аммонітян сказали до Хануна: Чи Давид шанує батька твого в очах твоїх тим, що послав тобі потішителів? Чи ж раби його прийшли до тебе не на те, щоб вивідати, і щоб знищити, і щоб вишпигувати край?
1CHR|19|4|І взяв Ханун Давидових рабів та й оголив їх, й обрізав їхню одежу в половині аж до сидіння, та й відпустив їх...
1CHR|19|5|І пішли й донесли Давидові про тих мужів, а він послав навпроти них, бо ті мужі були дуже осоромлені. І цар їм сказав: Сидіть в Єрихоні, аж поки відросте вам борода, потім повернетесь.
1CHR|19|6|І побачили аммонітяни, що вони зненавиджені в Давида. І послав Ханун та аммонітяни тисячу талантів срібла, щоб винайняти собі колесниці та верхівців з Араму двох річок і з Араму Маахи та з Цови.
1CHR|19|7|І найняли вони собі тридцять і дві тисячі колесниць, і царя Маахи та народ його, і прийшли й таборували перед Медевою. Також аммонітяни зібралися зо своїх міст і прийшли до бою.
1CHR|19|8|А коли Давид прочув про це, то послав Йоава та все військо лицарів.
1CHR|19|9|І повиходили аммонітяни, і вставилися до бою при вході до міста. А царі, що прийшли, вони самі були на полі.
1CHR|19|10|І побачив Йоав, що бойовий фронт став на нього спереду та позаду, то вибрав зо всього вибраного в Ізраїлі, та й установив їх навпроти сиріян.
1CHR|19|11|А решту народу дав під руку свого брата Ав'шая, й їх установили навпроти аммонітян,
1CHR|19|12|і сказав: Якщо сиріяни будуть сильніші від мене, то будеш мені на поміч, а якщо аммонітяни будуть сильніші від тебе, то допоможу тобі.
1CHR|19|13|Будь мужній, і стіймо міцно за народ наш та за міста нашого Бога, а Господь нехай зробить, що добре в очах Його!
1CHR|19|14|А коли Йоав та народ, що був із ним, підійшов перед сиріян до бою, то ті повтікали перед ним.
1CHR|19|15|А аммонітяни побачили, що повтікали сиріяни, то й вони повтікали перед братом його Ав'шаєм, і ввійшли до міста, а Йоав прибув до Єрусалиму.
1CHR|19|16|А коли побачили сиріяни, що вони побиті Ізраїлем, то послали послів, і привели сиріян, що з другого боку Річки, а Шофах, зверхник Гадад'езерового війська, був перед ними.
1CHR|19|17|І було донесено Давидові, і він зібрав усього Ізраїля, і перейшов Йордан та прийшов до них, і вставився проти них. І встановився Давид на бій проти сиріян, і вони воювали з ним.
1CHR|19|18|І побігли сиріяни перед Ізраїлем, а Давид повбивав із сиріян сім тисяч колесниць та сорок тисяч пішого люду. І вбив він Шофаха, зверхника війська...
1CHR|19|19|А коли Гадад'езерові раби побачили, що вони побиті Ізраїлем, то замирилися з Давидом і служили йому. І сиріяни вже не хотіли допомагати аммонітянам.
1CHR|20|1|І сталося по році, того часу, як царі виходили на війну, то Йоав повів військову силу, та й нищив аммонітський край. І прийшов він і обліг Раббу, а Давид сидів в Єрусалимі. І побив Йоав Раббу, і зруйнував її.
1CHR|20|2|І зняв Давид корону їхнього царя з голови його, і знайшов, що вага її талант золота, а на ній каміння дорогоцінне, і була покладена вона на голову Давидову! І він виніс дуже багато здобичі з того міста.
1CHR|20|3|А народ, що був у ньому, повиводив, і перетинав їх пилками, і забивав залізними долотами та сокирами... І так робив Давид усім аммонітським містам. І вернувся Давид та ввесь народ до Єрусалиму.
1CHR|20|4|І сталося по тому, і була війна в Ґезері з филистимлянами. Тоді хушанин Сіббехай убив Сіппая, з Рефаєвих нащадків, і вони були поконані.
1CHR|20|5|І була ще війна з филистимлянами, і Елханан, син Яірів, побив Лахмі, брата ґатянина Ґоліята, а держак списа його був, як ткацький вал!
1CHR|20|6|І була ще війна в Ґаті. А там був чоловік великого зросту, що мав по шість пальців, усього двадцять і чотири. І він також був із нащадків Рефая.
1CHR|20|7|І зневажав він Ізраїля, та забив його Йонатан, син Шім'ї, Давидового брата.
1CHR|20|8|Ці також походили від Рефая в Ґаті, і попадали вони від руки Давида та від руки його слуг.
1CHR|21|1|І повстав сатана на Ізраїля, і намовив Давида перелічити Ізраїля.
1CHR|21|2|І сказав Давид до Йоава та до начальників народу: Ідіть, перелічіть Ізраїля від Беер-Шеви й аж до Дану, і донесіть мені, і я знатиму число їх!
1CHR|21|3|І сказав Йоав: Нехай Господь додасть до народу Свого в сто раз стільки, скільки є! Чи не всі вони, пане мій царю, раби мого пана? Нащо буде шукати цього пан мій, нащо це буде за провину для Ізраїля?
1CHR|21|4|Та цареве слово перемогло Йоава. І вийшов Йоав, і ходив по всьому Ізраїлі, і вернувся до Єрусалиму.
1CHR|21|5|І дав Йоав Давидові число переліку народу. І було всього Ізраїля тисяча тисяч і сто тисяч чоловіка, що витягають меча, а Юди чотири сотні й сімдесят тисяч чоловіка, що витягають меча.
1CHR|21|6|А Левія та Веніямина він не перерахував серед них, бо царське слово було огидою для Йоава...
1CHR|21|7|І було зло в Божих очах на ту річ, і Він ударив Ізраїля!
1CHR|21|8|І сказав Давид до Бога: Я дуже згрішив, що зробив оцю річ! А тепер прости ж гріх Свого раба, бо я зробив дуже нерозумно!...
1CHR|21|9|І сказав Господь до Ґада, Давидового прозорливця, говорячи:
1CHR|21|10|Іди, і будеш говорити Давидові, кажучи: Так говорить Господь: Три карі кладу Я на тебе, вибери собі одну з них, і Я зроблю тобі.
1CHR|21|11|І прийшов Ґад до Давида та й сказав йому: Так сказав Господь: Вибери собі:
1CHR|21|12|чи три роки голоду, чи теж три місяці твого втікання перед ворогами твоїми, а меч ворогів твоїх доганятиме тебе, чи три дні Господнього меча та моровиці в Краю, і Ангол Господній буде нищити по всій Ізраїлевій границі. А тепер розваж, яке слово верну Я Тому, Хто послав мене...
1CHR|21|13|І сказав Давид до Ґада: Тяжко мені дуже! Нехай же впаду я в руку Господа, бо дуже велике Його милосердя, а в руку людську нехай я не впаду!...
1CHR|21|14|І дав Господь моровицю в Ізраїлі, і впало з Ізраїля сімдесят тисяч чоловіка!
1CHR|21|15|І послав Бог Ангола до Єрусалиму, щоб знищити його. А коли він нищив, Господь побачив і пожалував про це лихо. І сказав Він до Ангола, що вигублював: Забагато тепер! Попусти свою руку! А Ангол Господній стояв при тоці євусеянина Орнана.
1CHR|21|16|І підняв Давид очі свої та й побачив Господнього Ангола, що стояв між землею та між небом, а в руці його був витягнений меч, скерований на Єрусалим. І впав Давид та ті старші, покриті веретами, на обличчя свої...
1CHR|21|17|І сказав Давид до Бога: Чи ж не я сказав рахувати в народі? І я той, хто згрішив, і вчинити зло я вчинив зло, а ці вівці що зробили вони, Господи, Боже мій? Нехай же рука Твоя буде на мені та на домі батька мого, а не на народі Твоєму, щоб погубити його...
1CHR|21|18|А Ангол Господній говорив до Ґада, сказати Давидові, щоб Давид пішов поставити жертівника для Господа на току євусеянина Орнана.
1CHR|21|19|І пішов Давид за словом Ґада, що говорив в Господньому Імені.
1CHR|21|20|І обернувся Орнан, і побачив Ангола, а чотири сини його, що були з ним, поховалися. А Орнан молотив пшеницю.
1CHR|21|21|І прийшов Давид до Орнана. І виглянув Орнан, і побачив Давида, і вийшов із току, і поклонився Давидові обличчям до землі.
1CHR|21|22|І сказав Давид до Орнана: Дай же мені місце цього току, й я збудую на ньому жертівника для Господа. Дай мені його за срібло повної ваги, і буде стримана моровиця від народу.
1CHR|21|23|І сказав Орнан до Давида: Візьми собі, і нехай зробить мій пан цар, що добре в очах його. Дивися, я даю цю худобу на цілопалення, а молотарки на дрова, а пшеницю на хлібну жертву. Усе я даю!
1CHR|21|24|І сказав цар Давид до Орнана: Ні, бо купуючи, куплю за срібло повної ваги, бо не піднесу твого в жертві для Господа, і не спалю цілопалення дармо!
1CHR|21|25|І дав Давид Орнанові за місце золота вагою шість сотень шеклів.
1CHR|21|26|І збудував там Давид жертівника для Господа, і приніс цілопалення та мирні жертви. І кликнув він до Господа, і Він відповів йому огнем із небес на жертівник цілопалення.
1CHR|21|27|І сказав Господь до Ангола, і він уклав меча свого до піхов його.
1CHR|21|28|Того часу, як Давид побачив, що Господь відповів йому на току євусеянина Орнана, то приносив там жертву.
1CHR|21|29|А Господня скинія, яку зробив був Мойсей у пустині, та жертівник цілопалення були того часу на пагірку в Ґів'оні.
1CHR|21|30|Та не міг Давид піти перед нього, щоб запитатися в Бога, бо настрашився меча Господнього Ангола.
1CHR|22|1|І Давид сказав: Це той дім Господа Бога, і це жертівник на цілопалення для Ізраїля!
1CHR|22|2|І сказав Давид, щоб зібрати приходьків, що були в Ізраїлевому Краї, і поставив каменярів тесати брили каміння, щоб збудувати Божого дома.
1CHR|22|3|І заготовив Давид силу заліза на цвяхи для брамних дверей та на клямри, і таку силу міді, що їй не було ваги,
1CHR|22|4|і кедрового дерева без числа, бо сидоняни та тиряни спровадили Давидові силу кедрового дерева.
1CHR|22|5|І сказав Давид: Мій син Соломон ще юнак та тендітний, приготую ж йому все на цей храм на збудування для Господа, щоб піднести його високо на славу та на велич для всіх країв. Приготую ж я все для нього! І Давид заготовив безліч усього перед своєю смертю.
1CHR|22|6|І він покликав сина свого Соломона, і наказав йому збудувати храм для Господа, Бога Ізраїля.
1CHR|22|7|І сказав Давид до Соломона: Сину мій, я мав на своєму серці вибудувати храм для Ймення Господа, Бога мого.
1CHR|22|8|Та було про мене Господнє слово, кажучи: Безліч крови пролив ти та війни великі провадив. Не збудуєш ти храма для Мого Ймення, бо багато крови пролив ти на землю перед лицем Моїм!
1CHR|22|9|Ось народиться тобі син, він буде муж мирний, і Я дам йому мир від усіх ворогів його навколо, бо Соломон буде ім'я йому, і Я дам на Ізраїля за його днів мир та тишу.
1CHR|22|10|Він збудує храм для Мого Ймення, і він буде Мені за сина, а Я йому за Батька, і Я міцно поставлю трона царства його над Ізраїлем аж навіки!
1CHR|22|11|Тепер, сину мій, нехай Господь буде з тобою, і буде щастити тобі, і збудуєш ти дім для Господа, Бога свого, як говорив Він про тебе.
1CHR|22|12|Тільки нехай дасть тобі Господь розум та розважність, і нехай поставить тебе над Ізраїлем, і ти будеш стерегти Закон Господа, Бога свого.
1CHR|22|13|Тоді буде щастити тобі, якщо будеш додержувати, щоб чинити устави та права, які наказав був Господь Мойсеєві про Ізраїля. Будь сильний та міцний, не бійся й не страхайся!
1CHR|22|14|І ось я в скудоті своїй заготовив для Господнього дому сто тисяч талантів золота та тисячу тисяч талантів срібла, а для міді та для заліза нема ваги, бо безліч того; і дерева, і каміння заготовив я, а ти до них додаси.
1CHR|22|15|А в тебе безліч робітників для праці, теслярів і каменярів та дереворубів, та всяких здібних на всяку роботу.
1CHR|22|16|Золоту, сріблу, і міді та залізу нема числа. Стань і зроби, і нехай Господь буде з тобою!
1CHR|22|17|І наказав Давид усім Ізраїлевим князям, щоб допомагали синові його Соломонові:
1CHR|22|18|Чи Господь, Бог ваш, не з вами? І Він дав вам мир навколо, бо дав у мою руку мешканців цієї землі, і була здобута ця земля перед лицем Господа та перед народом Його.
1CHR|22|19|Тепер прихиліть серце ваше та душу вашу, щоб шукати Господа, Бога вашого. І встаньте, і збудуйте святиню Господа Бога, щоб перенести ковчега Господнього заповіту та святі Божі речі до храму, збудованого для Господнього Ймення.
1CHR|23|1|А коли Давид постарів і наситився днями, то він поставив царем над Ізраїлем сина свого Соломона.
1CHR|23|2|І зібрав він усіх Ізраїлевих князів, і священиків та Левитів.
1CHR|23|3|І були перелічені Левити від віку тридцяти років і вище, і було число їх, за їхніми головами, за мужчинами тридцять і вісім тисяч.
1CHR|23|4|Із них для керування над роботою Господнього дому двадцять і чотири тисячі, а урядників та суддів шість тисяч,
1CHR|23|5|і чотири тисячі придверних, і чотири тисячі тих, що славлять Господа на музичних знаряддях, які я зробив на славлення.
1CHR|23|6|І поділив їх Давид на черги за синами Левія, для Ґершона, Кегата та Мерарі.
1CHR|23|7|З Ґершонівців Ладан і Шім'ї.
1CHR|23|8|Ладанові сини: голова Єгіїл, і Зетам, і Йоїл, троє.
1CHR|23|9|Сини Шім'ї: Шеломіт, і Хазаїл, і Гаран, троє, вони голови батьківських домів Ладана.
1CHR|23|10|А сини Шім'ї: Яхат, Зіза, і Єуш, і Берія, оце сини Шім'ї, четверо.
1CHR|23|11|І був Яхат головою, а Зіза другий, а Єуш та Берія не мали багато синів, і стали за один батьківський дім при переліченні.
1CHR|23|12|Кегатові сини: Амрам, Іцгар, Хеврон та Уззіїл, четверо.
1CHR|23|13|Амрамові сини: Аарон та Мойсей. І був відділений Аарон, щоб посвятити його до Святого Святих, його та синів його аж навіки, щоб кадити перед лицем Господа, щоб служити Йому та щоб благословляти Ім'ям Його аж навіки.
1CHR|23|14|А Мойсей Божий чоловік, сини його полічені до Левієвого племени.
1CHR|23|15|Сини Мойсеєві: Ґершом та Еліезер.
1CHR|23|16|Сини Ґершомові: Шевуїл, голова.
1CHR|23|17|А сини Еліезерові були: Рехавія, голова; і не було в Еліезера інших синів, а сини Рехавії сильно помножились.
1CHR|23|18|Сини Їцгарові: Шеломіт, голова.
1CHR|23|19|Сини Хевронові: Єрійя голова, Амарія другий, Яхазіїл третій, і Єкам'ам четвертий.
1CHR|23|20|Сини Уззіїлові: Міхал голова, а Їшшійя другий.
1CHR|23|21|Сини Мерарієві: Махлі й Муші. Сини Махлі: Елеазар і Кіш.
1CHR|23|22|І помер Елеазар, і не було в нього синів, бо тільки дочки, і їх побрали собі Кішові сини, їхні брати.
1CHR|23|23|Сини Мушієві: Махлі, і Едер, і Єремот, троє.
1CHR|23|24|Оце сини Левієві за домом батьків їх, голови дому батьків за перегляненням їхнім, числом імен за особами їх, що чинили роботу для будови Господнього дому, від віку двадцяти років і вище.
1CHR|23|25|Бо Давид сказав: Господь, Бог Ізраїля, дав мир Своєму народові, і він осівся в Єрусалимі аж навіки.
1CHR|23|26|І також Левитам не треба носити скинії та всіх речей її для служби їй,
1CHR|23|27|бо за останніми наказами Давида вони становлять число Левієвих синів від віку двадцяти літ і вище.
1CHR|23|28|Бо їхнє становище при руці Ааронових синів для служби Господнього дому над подвір'ями, і над кімнатами, і над чистістю усіх святощів та роботи служби Господнього дому,
1CHR|23|29|і при хлібі виставнім, і при пшеничній муці на хлібну жертву та на прісні коржі, і при сковородах, і при праженні, і при всякій мірі ваги та мірі довжини.
1CHR|23|30|І щоб ставати щоранку на подяку та на хвалу Господа, і так і на вечір.
1CHR|23|31|І при всякому спаленні цілопалень для Господа на суботи, на молодики, і на свята в числі за правом на них, завжди перед лицем Господнім.
1CHR|23|32|І чинили вони охорону скинії заповіту, і сторожу святині, і охорону Ааронових синів, своїх братів, при службі Господнього дому.
1CHR|24|1|А в Ааронових синів такі їхні черги: Ааронові сини: Надав і Авігу, Елеазар і Ітамар.
1CHR|24|2|Та повмирали Надав та Авігу за життя їхнього батька, і не мали вони синів, тому священнодіяли Елеазар та Ітамар.
1CHR|24|3|І поділив їх Давид і Садок, з Елеазарових синів, та Ахімелех, з Ітамарових синів, за їхнім урядом в їхній службі.
1CHR|24|4|І були знайдені Елеазарові сини численнішими, щодо голів чоловіків, від синів Ітамарових. І вони поділили їх: для Елеазарових синів голів дому батьків було шістнадцять, а для Ітамарових синів для дому батьків їх вісім.
1CHR|24|5|І поділили їх жеребками, тих з тими, бо головними в святині та головними перед Богом були з синів Елеазарових та серед синів Ітамарових.
1CHR|24|6|І записав їх Шемая, син Натанаїлів, писар із Левитів, перед царем, і головними, і священиком Садоком, і Ахімелехом, сином Евіятаровим, і головами дому батьків священиків та Левитів. Один батьківський дім був узятий для Елеазара, а один був узятий для Ітамара.
1CHR|24|7|І вийшов перший жеребок для Єгояріва, другий для Єдаї,
1CHR|24|8|третій для Харіма, четвертий для Сеоріма,
1CHR|24|9|п'ятий для Малкійї, шостий для Мійяміна,
1CHR|24|10|сьомий для Гаккоца, восьмий для Авійї,
1CHR|24|11|дев'ятий для Єшуї, десятий для Шеханії,
1CHR|24|12|одинадцятий для Ел'яшіва, дванадцятий для Якіма,
1CHR|24|13|тринадцятий для Хуппи, чотирнадцятий для Єшев'ава,
1CHR|24|14|п'ятнадцятий для Білґи, шістнадцятий для Іммера,
1CHR|24|15|сімнадцятий для Хезіра, вісімнадцятий для Гаппіццеца,
1CHR|24|16|дев'ятнадцятий для Петах'ї, двадцятий для Єхезкела,
1CHR|24|17|двадцять і перший для Яхіна, двадцять і другий для Ґамула,
1CHR|24|18|двадцять і третій для Делаї, двадцять і четвертий для Маазії.
1CHR|24|19|Оце порядок їхньої служби, щоб приходити до Господнього дому за їхньою постановою через Аарона, їхнього батька, як йому наказав був Господь, Бог Ізраїлів.
1CHR|24|20|А від позосталих Левієвих синів: від Амрамових синів Шуваїл, від синів Шуваїлових Єхедія.
1CHR|24|21|Від Рехавії, від синів Рехавії: голова Їшшійя.
1CHR|24|22|Від Їцгарівців: Шеломот, від Шеломотових синів: Яхат.
1CHR|24|23|А сини Хевронові: Єрійя, другий Амарія, третій Яхазіїл, четвертий Єкам'ам.
1CHR|24|24|Сини Уззіїлові: Міха, сини Міхині: Шамір.
1CHR|24|25|Брат Міхи Їшшійя, сини Їшшійїні Захарій.
1CHR|24|26|Сини Мерарієві: Махлі та Муші, сини Яазійї Бено.
1CHR|24|27|Сини Мерарієві, від Яазійї: Бено, і Шогам, і Заккур, і Іврі.
1CHR|24|28|У Махлі: Елеазар, у нього не було синів.
1CHR|24|29|Від Кіша, сини Кішові: Єрахмеїл.
1CHR|24|30|А сини Мушієві: Махлі, і Едер, і Єрімот. Оце сини Левитів, за домом їхніх батьків.
1CHR|24|31|І кидали жеребки і вони відповідно до братів своїх, Ааронових синів, перед царем Давидом, і Садоком, і Ахімелехом, і головами дому батьків священиків та Левитів, голови родин нарівні зо своїм меншим братом.
1CHR|25|1|І відділив Давид та зверхники війська на службу синів Асафа, і Гемана, і Єдутуна, що провіщували на цитрах, і на арфах, і на цимбалах. А число їх, людей праці до служби, було таке:
1CHR|25|2|від Асафових синів: Заккур, і Йосип, і Нетанія, і Асар'їла, Асафові сини, при Асафі, що пророкував при царі.
1CHR|25|3|Від Єдутуна, Єдутунові сини: Ґедалія, і Цері, і Ісая, Хашавія, і Маттітія, шестеро при своєму батькові Єдутуні, що пророкував на цитрі на дяку та на хвалу Господеві.
1CHR|25|4|Від Гемана, Геманові сини: Буккійя, Маттанія, Уззіїл, Шевуїл, і Єрімот, Хананія, Ханані, Еліата, Ґіддалті, і Ромамті, Езер, Йошбекаша, Маллоті, Готір, Махазіот.
1CHR|25|5|Усі ці сини Гемана, царського прозорливця в Божих словах, щоб підвищувати силу. І дав Бог Геманові чотирнадцять синів та три дочки.
1CHR|25|6|Усі вони були при своєму батькові, на співі Господнього дому, на цимбалах, на арфах та цитрах для служби в Божому домі; при царі Асаф, Єдутун та Геман.
1CHR|25|7|І було їхнє число з їхніми братами, вивченими співу для Господа, усіх розуміючих, двісті й вісімдесят і вісім.
1CHR|25|8|І кинули вони жеребки, черга відповідно черзі, як малий, так і великий, учитель з учнем.
1CHR|25|9|І вийшов перший жеребок від Асафа для Йосипа, другий Ґедалія, він і брати його та сини його, дванадцять.
1CHR|25|10|Третій Заккур, сини його та брати його, дванадцять.
1CHR|25|11|Четвертий для Їцрі, сини його та брати його, дванадцять.
1CHR|25|12|П'ятий Нетанія, сини його та брати його, дванадцять.
1CHR|25|13|Шостий Буккійя, сини його та брати його, дванадцять.
1CHR|25|14|Сьомий Єсар'їла, сини його та брати його, дванадцять.
1CHR|25|15|Восьмий Ісая, сини його та брати його, дванадцять.
1CHR|25|16|Дев'ятий Маттанія, сини його та брати його, дванадцять.
1CHR|25|17|Десятий Шім'ї, сини його та брати його, дванадцять.
1CHR|25|18|Одинадцятий Азаріїл, сини його та брати його, дванадцять.
1CHR|25|19|Дванадцятий для Хашав'ї, сини його та брати його, дванадцять.
1CHR|25|20|Тринадцятий для Шуваїла, сини його та брати його, дванадцять.
1CHR|25|21|Чотирнадцятий для Маттітії, сини його та брати його, дванадцять.
1CHR|25|22|П'ятнадцятий для Єремота, сини його та брати його, дванадцять.
1CHR|25|23|Шістнадцятий для Хананії, сини його брати його, дванадцять.
1CHR|25|24|Сімнадцятий для Йошбекаші, сини його та брати його, дванадцять.
1CHR|25|25|Вісімнадцятий для Ханані, сини його та брати його, дванадцять.
1CHR|25|26|Дев'ятнадцятий для Маллоті, сини його та брати його, дванадцять.
1CHR|25|27|Двадцятий для Елійяти, сини його та брати його, дванадцять.
1CHR|25|28|Двадцять і перший для Готіра, сини його та брати його, дванадцять.
1CHR|25|29|Двадцять і другий для Ґіддалті, сини його та брати його, дванадцять.
1CHR|25|30|Двадцять і третій для Махазіота, сини його та брати його, дванадцять.
1CHR|25|31|Двадцять і четвертий для Ромамті-Езера, сини його та брати його, дванадцять.
1CHR|26|1|Черги придверних, від Корахівців: Мешелемія, син Коре, з Асафових синів.
1CHR|26|2|А в Мешелемії сини: первороджений Захарій, другий Єдіаїл, третій Зевадія, четвертий Ятніїл,
1CHR|26|3|п'ятий Елам, шостий Єгоханан, сьомий Ел'єгоенай.
1CHR|26|4|А в Овед-Едома сини: первороджений Шемая, другий Єгозавад, третій Йоах, четвертий Сахар, і п'ятий Натанаїл,
1CHR|26|5|шостий Амміїл, сьомий Іссахар, восьмий Пеуллетай, бо поблагословив його Бог.
1CHR|26|6|У сина його Шемаї народилися сини, що панували над домом їхнього батька, бо вони хоробрі вояки.
1CHR|26|7|Сини Шемаї: Отні, і Рефаїл, і Овед, Елзавад; його брати, мужі хоробрі, Елігу та Шемахія.
1CHR|26|8|Усі ці з Оведових синів; вони й сини та брати їхні кожен хоробрий муж у силі до праці, шістдесят і два для Овед-Едома.
1CHR|26|9|А в Мешелемії було синів та братів, мужів хоробрих, вісімнадцять.
1CHR|26|10|А в Хоси, з синів Мерарі, сини: голова Шімрі, бо хоч не був він первороджений, та батько його настановив його за голову:
1CHR|26|11|другий Хілкійя, третій Тевалія, четвертий Захарій; усіх синів та братів у Хоси тринадцять.
1CHR|26|12|У цих були черги придверних, за головами мужчин, черги відповідно до їхніх братів на служення в Господньому домі.
1CHR|26|13|І кинули вони жеребки, як малий, так і великий, за домом їхніх батьків, для кожної брами.
1CHR|26|14|І впав жеребок на схід для Шелемії. І кинули жеребки для сина його Захарія, мудрого дорадника, і вийшов жеребок його на північ,
1CHR|26|15|для Овед-Едома, на південь, а для синів його комори.
1CHR|26|16|Для Шуппіма та для Хоси на захід, разом із брамою Шаллехет, де підіймається битий шлях, варта навпроти варти.
1CHR|26|17|На схід шість Левитів, на північ четверо на день, на південь четверо на день, а для комори по двоє.
1CHR|26|18|Для Парбару на захід четверо для битого шляху, двоє для Парбару.
1CHR|26|19|Оце черги придверних із синів Корахівців та з синів Мерарі.
1CHR|26|20|А Левити: Ахійя був над скарбами Божого дому та до скарбів святині.
1CHR|26|21|Сини Ладана, сини Ґершонівців, від Ладана, голови дому батьків, від Ладана Ґершонівця: Єхіїлі.
1CHR|26|22|Сини Єхіїлі: Зетам та Йоїл, брат його, над скарбами Господнього дому.
1CHR|26|23|Для Амрамівців, для Їцгарівців, для Хевронівців, для Аззіїлівців:
1CHR|26|24|Шевуїл, син Ґершома, сина Мойсея, володар над скарбами.
1CHR|26|25|А брати його від Еліезера: його син Рехавія, і його син Ісая, і його син Йорам, і його син Зіхрі, і його син Шеломіт.
1CHR|26|26|Цей Шеломіт та брати його були над усіма скарбами святині, які посвятив цар Давид та голови дому батьків, і тисячники, і сотники та зверхники війська,
1CHR|26|27|з воєн та зо здобичі вони присвячували на підтримання Господнього дому,
1CHR|26|28|і все, що посвятив прозорливець Самуїл, і Саул, син Кішів, і Авнер, син Нерів, і Йоав, син Церуїн, усе посвячене було в руці Шеломіта та братів його.
1CHR|26|29|Від Їцгарівців: Кенанія та сини його на зовнішню роботу над Ізраїлем, на писарів та на суддів.
1CHR|26|30|Від Хевронівців: Хашавія та брати його, мужі хоробрі, тисяча й сім сотень, над переглядом Ізраїля з другого боку Йордану на захід, для всякої Господньої праці та для роботи царської.
1CHR|26|31|Від Хевронівців: Єрійя голова для Хевронівця, для його нащадків, за домом батьків. У сороковому році Давидового царювання вони були досліджені, і серед них знайдено хоробрих мужів в гілеадському Язері.
1CHR|26|32|А брати його мужі хоробрі, дві тисячі й сім сотень, голови дому батьків. І цар Давид настановив їх над Рувимівцями і над Ґадівцями та над половиною племени Манасіїного для всякої Божої справи та справи царської.
1CHR|27|1|А Ізраїлеві сини, за їхнім числом, голови батьківських родів і тисячники, і сотники та їхні урядники служили цареві щодо всякої справи відділів, що приходив та відходив місяць у місяць для всіх місяців року; один відділ мав двадцять і чотири тисячі.
1CHR|27|2|Над першим відділом, на перший місяць Яшов'ам, син Завдіїлів, а на відділ його двадцять і чотири тисячі.
1CHR|27|3|Він був з Перецових синів, голова всіх військових зверхників на перший місяць.
1CHR|27|4|А над відділом другого місяця Ахохівець Додай, а володар його відділу Міклот; а на його відділ ішло двадцять і чотири тисячі.
1CHR|27|5|Третій зверхник війська на третій місяць священик Беная, голова, а на його відділ двадцять і чотири тисячі.
1CHR|27|6|Цей Беная лицар із тридцяти й над тридцятьма; а над його відділом був син його Аммізавад.
1CHR|27|7|Четвертий на місяць четвертий Асаїл, брат Йоавів, а по ньому син його Зевадія; а на його відділ двадцять і чотири тисячі.
1CHR|27|8|П'ятий на місяць п'ятий зверхник ізрах'янин Шамут, а на його відділ двадцять і чотири тисячі.
1CHR|27|9|Шостий на місяць шостий Іра, син текоянина Іккеша, а на його відділ двадцять і чотири тисячі.
1CHR|27|10|Сьомий на місяць сьомий пелонянин Хелец з Єфремових синів, а на його відділ двадцять і чотири тисячі.
1CHR|27|11|Восьмий на місяць восьмий хушанин Сіббехай з Зерахівців, а на його відділ двадцять і чотири тисячі.
1CHR|27|12|Дев'ятий на місяць дев'ятий анатонянин Авіезер з Веніяминівців, а на його відділ двадцять і чотири тисячі.
1CHR|27|13|Десятий на місяць десятий нетоф'янин Магарай з Зерахівців, а на його відділ двадцять і чотири тисячі.
1CHR|27|14|Одинадцятий на одинадцятий місяць пір'атонянин Беная з Єфремових синів, а на його відділ двадцять і чотири тисячі.
1CHR|27|15|Дванадцятий на дванадцятий місяць нетоф'янин Хелдай з Отніїла, а на його відділ двадцять і чотири тисячі.
1CHR|27|16|А над Ізраїлевими племенами були: для Рувимівців володар Еліезер, син Зіхрі; для Симеонівців Шефатія, син Маахи.
1CHR|27|17|Для Левія Хашавія, син Кемуїла, для Аарона Садок.
1CHR|27|18|Для Юди Елігу, з Давидових братів, для Іссахара Омрі, син Михаїлів.
1CHR|27|19|Для Завулона Їшмая, син Овадії, для Нефталима Єрімот син Азріїлів.
1CHR|27|20|Для Єфремових синів Осія, син Азазії, для половини Манасіїного племени Йоїл, син Педаї.
1CHR|27|21|Для половини Манасії в Ґілеаді Їддо, син Захарія, для Веніямина Яасіїл, син Авнерів.
1CHR|27|22|Для Дана Азаріїл, син Єрохамів. Оце зверхники Ізраїлевих племен.
1CHR|27|23|А Давид не перелічив їхнього числа від віку двадцяти літ і нижче, бо Господь сказав був, що розмножить Ізраїля, як зорі небесні.
1CHR|27|24|Йоав, син Церуїн, зачав був лічити, та не скінчив. І був за те гнів на Ізраїля, і не ввійшло те число в число хроніки царя Давида.
1CHR|27|25|А над скарбами царськими Азмавет, Адіїлів син, а над скарбами на полі, у містах, і в селах та в баштах Єгонатан, син Уззійї.
1CHR|27|26|А над тими, що робили польову роботу, для праці, на землі Езрі, син Келувів.
1CHR|27|27|А над виноградниками рам'янин Шім'ї, а над тим, що в виноградниках для запасів вина шефам'янин Завді.
1CHR|27|28|А над оливками та над сикоморами, що в Шефелі, ґедерянин Баал-Ханан; а над скарбами оливи Йоаш.
1CHR|27|29|А над великою худобою, що пасеться в Шароні, шаронянин Шітрай, а над великою худобою в долинах Шафат, син Адлаїв.
1CHR|27|30|А над верблюдами їзмаїльтянин Овіл, а над ослицями меронотянин Єхдея.
1CHR|27|31|А над дрібною худобою гаґрянин Язіз. Усі оці зверхники маєтку, що мав цар Давид.
1CHR|27|32|А Йонатан, Давидів дядько, був радник, він чоловік розумний та писар. А Єхіїл, син Нахмоніїв, був із царськими синами.
1CHR|27|33|А Ахітофель радник цареві, а арк'янин Хушай приятель царів.
1CHR|27|34|А по Ахітофелю Єгояда, син Бенаї, та Евіятар, а зверхник царського війська Йоав.
1CHR|28|1|І зібрав Давид усіх Ізраїлевих князів, зверхників племен, і зверхників відділів, що служать цареві, і тисячників, і сотників, і зверхників усякого маєтку та добутку царя та синів його разом з евнухами та лицарями, та всякого хороброго вояка до Єрусалиму.
1CHR|28|2|І встав цар Давид на ноги свої та й сказав: Послухайте мене, брати мої та народе мій! Я серцем своїм був за те, щоб збудувати храм миру для ковчега Господнього заповіту та на підніжок ніг нашого Бога, й я приготовив потрібне на збудування.
1CHR|28|3|А Бог сказав мені: Ти не збудуєш храма для Мого Ймення, бо ти муж воєн і кров проливав.
1CHR|28|4|Та вибрав Господь, Бог Ізраїлів, мене з усього дому батька мого, щоб бути царем над Ізраїлем навіки, бо Юду вибрав Він на володаря, а серед Юдиного дому дім батька мого, а серед синів мого батька мене уподобав Собі, щоб настановити царем над усім Ізраїлем.
1CHR|28|5|А зо всіх моїх синів, бо багатьох синів дав мені Господь то Він вибрав сина мого Соломона, щоб сидів на троні Господнього царства над Ізраїлем.
1CHR|28|6|І Він сказав мені: Соломон, син твій, він збудує храма Мого та двори Мої, бо його Я вибрав Собі за сина, а Я буду йому за Отця.
1CHR|28|7|І міцно поставлю Я царство його аж навіки, якщо він буде сильний, щоб виконувати заповіді Мої та постанови Мої, як цього дня.
1CHR|28|8|А тепер на очах усього Ізраїля, Господнього збору, та в ушах нашого Бога говорю вам: Додержуйте й досліджуйте всі заповіді Господа, Бога вашого, щоб ви посіли цей добрий Край і віддали його в спадщину по собі синам вашим аж навіки.
1CHR|28|9|А тепер, сину мій Соломоне, знай Бога, Отця твого, і служи Йому всім серцем та всією душею, бо Господь вивідує всі серця та знає всякий витвір думок. Якщо будеш шукати Його, то ти знайдеш Його, а якщо залишиш Його, Він залишить тебе назавжди.
1CHR|28|10|Тепер дивися, що Господь вибрав тебе збудувати дім на святиню. Будь міцний та роби!
1CHR|28|11|І Давид дав своєму синові Соломонові взори Господнього дому: притвору, і домів його, і скарбниць його, і горниць його, і кімнат його внутрішніх, і дому для ковчегу,
1CHR|28|12|і взір усього, що було в дусі його для подвір'я Господнього дому, і для всіх кімнат навколо, для скарбів Божого дому та для скарбів святині,
1CHR|28|13|і для відділів священиків та Левитів, і для всякої праці служби Господнього дому, і для всяких речей для служби Господнього дому.
1CHR|28|14|І дав він золота вагою для золота, для всіх речей кожної служби; і срібла для всіх срібних речей вагою, для всіх речей кожної служби;
1CHR|28|15|і вагу для золотих свічників та золотих їхніх лямпадок, вагою кожного свічника та лямпадок його, і для срібних свічників, вагою для свічника та лямпадок його, за роботою кожного свічника.
1CHR|28|16|І дав золота вагою для столів хлібів показних, для кожного столу і срібла для срібних столів,
1CHR|28|17|і видельця, і кропильниці, і чарки чисте золото, і для золотих келіхів вагою для кожного келіха, і для келіхів срібних, вагою для кожного келіха.
1CHR|28|18|А для кадильного жертівника дав очищеного золота вагою, і на подобу воза, для золотих херувимів, що простягають крила свої й покривають над ковчегом Господнього заповіту.
1CHR|28|19|Усе це він зрозумів із письма з Господньої руки, що була над ним, усі роботи взору.
1CHR|28|20|І сказав Давид до сина свого Соломона: Будь сильний і будь відважний, і роби, не бійся та не лякайся, бо Господь Бог, Бог мій, з тобою, Він не покине тебе й не позоставить тебе аж до закінчення всієї праці роботи Господнього дому...
1CHR|28|21|А оце черги священиків та Левитів для всякої служби Божого дому. І будуть з тобою в усякій праці ревні люди, здібні на всяку службу, а начальники та ввесь народ, на всі накази твої.
1CHR|29|1|І сказав цар Давид до всього збору: Син мій Соломон, що його одного Бог вибрав, ще молодий та тендітний, а ця праця велика, бо не для людини ця будова, а для Господа Бога.
1CHR|29|2|А Я всією своєю силою приготовив для храму свого Бога золото на золоті речі, і срібло на срібні, і мідь на мідяні, і залізо на залізні, і дерево на дерев'яні, каміння шогамське та до оправ, каміння нофехське та кольорове, і всякий дорогий камінь та безліч мармурового каміння.
1CHR|29|3|І ще, через моє замилування до дому Бога мого, є в мене скарб власного золота та срібла, і його я віддав для дому свого Бога, понад усе, що я заготовив для святого храму:
1CHR|29|4|три тисячі талантів золота, офірського золота, і сім тисяч очищеного срібла на покриття стін тих домів;
1CHR|29|5|на кожну золоту річ та на кожну срібну, і на всяку працю рукою майстрів. І хто ще жертвує, щоб сьогодні наповнити свою руку пожертвою для Господа?
1CHR|29|6|І стали жертвувати начальники батьківських родів та начальники Ізраїлевих племен, і тисячники та сотники, і начальники праці для царя.
1CHR|29|7|І дали вони на роботу Божого дому золота п'ять тисяч талантів та десять тисяч дарейків, і срібла десять тисяч талантів, і міді десять тисяч і вісім тисяч талантів, а заліза сто тисяч талантів.
1CHR|29|8|А в кого знайшлося при ньому дорогоцінне каміння, ті дали його до скарбниці Господнього дому, до руки Ґершонівця Єхіїла.
1CHR|29|9|І радів народ за їхню жертву, бо вони жертвували Господеві з цілого серця, а також цар Давид радів великою радістю.
1CHR|29|10|І поблагословив Давид Господа на очах усього збору. І сказав Давид: Благословенний Ти, Господи, Боже Ізраїля, нашого батька, від віку й аж до віку!
1CHR|29|11|Твоя, Господи, могутність і сила, і велич, і вічність, і слава, і все на небесах та на землі! Твої, Господи, царства, і Ти піднесений над усім за Голову!
1CHR|29|12|І багатство та слава від Тебе, і Ти пануєш над усім, і в руці Твоїй сила та хоробрість, і в руці Твоїй побільшити та зміцнити все.
1CHR|29|13|А тепер, Боже наш, ми дякуємо Тобі, і славимо Ім'я Твоєї величі.
1CHR|29|14|І хто бо я, і хто народ мій, що маємо силу так жертвувати, як це? Бо все це від Тебе, і з Твоєї руки дали ми Тобі.
1CHR|29|15|Бо ми приходьки перед лицем Твоїм та чужинці, як усі наші батьки! Наші дні на землі мов та тінь, і немає тривалого!
1CHR|29|16|Господи, Боже наш, уся ця безліч, яку ми наготовили на збудування Тобі храму для Ймення Твоєї святости, із Твоєї руки вона, і все це Твоє!
1CHR|29|17|І я знаю, Боже мій, що Ти вивідуєш серце й любиш щирість. У щирості серця свого я пожертвував це все, а тепер бачу я з радістю народ Твій, який знаходиться тут, що жертвує себе Тобі.
1CHR|29|18|Господи, Боже Авраама, Ісака та Якова, наших батьків, збережи ж навіки цей напрямок думок серця народу Твого, і міцно скеруй їхнє серце до Себе!
1CHR|29|19|А моєму синові Соломонові дай серце ціле, щоб виконувати заповіді Твої, свідоцтва Твої та устави Твої, і щоб чинити все, і щоб збудувати цю твердиню, яку я приготовив!
1CHR|29|20|І сказав Давид до всього збору: Поблагословіть же Господа, вашого Бога! І ввесь збір поблагословив Господа, Бога своїх батьків, і нахилилися, і вклонилися всі до землі Господеві й цареві!
1CHR|29|21|І принесли вони для Господа жертви, і спалили цілопалення для Господа другого дня від того дня, тисячу бичків, тисячу баранів, тисячу овечок, і ливні їхні жертви, і безліч жертов за всього Ізраїля.
1CHR|29|22|І вони їли й пили перед Господом того дня з великою радістю, і вдруге настановили Соломона, Давидового сина, і помазали його Господеві на володаря, а Садока на священика.
1CHR|29|23|І сів Соломон на Господньому троні за царя на місці свого батька Давида, і щастило йому, і його слухався ввесь Ізраїль.
1CHR|29|24|І всі князі та лицарі, а також усі сини царя Давида піддалися під Соломона.
1CHR|29|25|І Господь високо звеличив Соломона на очах усього Ізраїля, і дав на нього величність царства, якої не було перед ним ані на жодному цареві над Ізраїлем.
1CHR|29|26|І Давид, син Єссеїв, царював над усім Ізраїлем.
1CHR|29|27|А дні, що він царював над Ізраїлем, були сорок літ: у Хевроні царював він сім років, а в Єрусалимі царював тридцять і три.
1CHR|29|28|І помер він у добрій сивині, ситий днями, багатством та славою, а замість нього зацарював син його Соломон.
1CHR|29|29|А діла царя Давида, перші й останні, ось вони описані в історії провидця Самуїла, і в історії пророка Натана, і в історії прозорливця Ґада,
1CHR|29|30|разом з усім царством його, і лицарськістю його та часами, що перейшли над ним і над Ізраїлем, та над усіма царствами тих країв.
