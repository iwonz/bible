JUDG|1|1|post mortem Iosue consuluerunt filii Israhel Dominum dicentes quis ascendet ante nos contra Chananeum et erit dux belli
JUDG|1|2|dixitque Dominus Iudas ascendet ecce tradidi terram in manus eius
JUDG|1|3|et ait Iudas Symeoni fratri suo ascende mecum in sorte mea et pugna contra Chananeum ut et ego pergam tecum in sorte tua et abiit cum eo Symeon
JUDG|1|4|ascenditque Iudas et tradidit Dominus Chananeum ac Ferezeum in manus eorum et percusserunt in Bezec decem milia virorum
JUDG|1|5|inveneruntque Adonibezec in Bezec et pugnaverunt contra eum ac percusserunt Chananeum et Ferezeum
JUDG|1|6|fugit autem Adonibezec quem secuti conprehenderunt caesis summitatibus manuum eius ac pedum
JUDG|1|7|dixitque Adonibezec septuaginta reges amputatis manuum ac pedum summitatibus colligebant sub mensa mea ciborum reliquias sicut feci ita reddidit mihi Deus adduxeruntque eum in Hierusalem et ibi mortuus est
JUDG|1|8|obpugnantes ergo filii Iuda Hierusalem ceperunt eam et percusserunt in ore gladii tradentes cunctam incendio civitatem
JUDG|1|9|et postea descendentes pugnaverunt contra Chananeum qui habitabat in montanis et ad meridiem et in campestribus
JUDG|1|10|pergensque Iudas contra Chananeum qui habitabat in Hebron cui nomen fuit antiquitus Cariatharbe percussit Sisai et Ahiman et Tholmai
JUDG|1|11|atque inde profectus abiit ad habitatores Dabir cuius nomen vetus erat Cariathsepher id est civitas Litterarum
JUDG|1|12|dixitque Chaleb qui percusserit Cariathsepher et vastaverit eam dabo ei Axam filiam meam uxorem
JUDG|1|13|cumque cepisset eam Othonihel filius Cenez frater Chaleb minor dedit ei filiam suam coniugem
JUDG|1|14|quam pergentem in itinere monuit vir suus ut peteret a patre suo agrum quae cum suspirasset sedens asino dixit ei Chaleb quid habes
JUDG|1|15|at illa respondit da mihi benedictionem quia terram arentem dedisti mihi da et inriguam aquis dedit ergo ei Chaleb inriguum superius et inriguum inferius
JUDG|1|16|filii autem Cinei cognati Mosi ascenderunt de civitate Palmarum cum filiis Iuda in desertum sortis eius quod est ad meridiem Arad et habitaverunt cum eo
JUDG|1|17|abiit autem Iudas cum Symeone fratre suo et percusserunt simul Chananeum qui habitabat in Sephath et interfecerunt eum vocatumque est nomen urbis Horma id est anathema
JUDG|1|18|cepitque Iudas Gazam cum finibus suis et Ascalonem atque Accaron cum terminis suis
JUDG|1|19|fuitque Dominus cum Iuda et montana possedit nec potuit delere habitatores vallis quia falcatis curribus abundabant
JUDG|1|20|dederuntque Chaleb Hebron sicut dixerat Moses qui delevit ex ea tres filios Enach
JUDG|1|21|Iebuseum autem habitatorem Hierusalem non deleverunt filii Beniamin habitavitque Iebuseus cum filiis Beniamin in Hierusalem usque in praesentem diem
JUDG|1|22|domus quoque Ioseph ascendit in Bethel fuitque Dominus cum eis
JUDG|1|23|nam cum obsiderent urbem quae prius Luza vocabatur
JUDG|1|24|viderunt hominem egredientem de civitate dixeruntque ad eum ostende nobis introitum civitatis et faciemus tecum misericordiam
JUDG|1|25|qui cum ostendisset eis percusserunt urbem in ore gladii hominem autem illum et omnem cognationem eius dimiserunt
JUDG|1|26|qui dimissus abiit in terram Etthim et aedificavit ibi civitatem vocavitque eam Luzam quae ita appellatur usque in praesentem diem
JUDG|1|27|Manasses quoque non delevit Bethsan et Thanach cum viculis suis et habitatores Dor et Ieblaam et Mageddo cum viculis suis coepitque Chananeus habitare cum eis
JUDG|1|28|postquam autem confortatus est Israhel fecit eos tributarios et delere noluit
JUDG|1|29|Ephraim etiam non interfecit Chananeum qui habitabat in Gazer sed habitavit cum eo
JUDG|1|30|Zabulon non delevit habitatores Cetron et Naalon sed habitavit Chananeus in medio eius factusque est ei tributarius
JUDG|1|31|Aser quoque non delevit habitatores Achcho et Sidonis Alab et Achazib et Alba et Afec et Roob
JUDG|1|32|habitavitque in medio Chananei habitatoris illius terrae nec interfecit eum
JUDG|1|33|Nepthali non delevit habitatores Bethsemes et Bethanath et habitavit inter Chananeum habitatorem terrae fueruntque ei Bethsemitae et Bethanitae tributarii
JUDG|1|34|artavitque Amorreus filios Dan in monte nec dedit eis locum ut ad planiora descenderent
JUDG|1|35|habitavitque in monte Hares quod interpretatur testaceo in Ahilon et Salabim et adgravata est manus domus Ioseph factusque est ei tributarius
JUDG|1|36|fuit autem terminus Amorrei ab ascensu Scorpionis Petra et superiora loca
JUDG|2|1|ascenditque angelus Domini de Galgal ad locum Flentium et ait eduxi vos de Aegypto et introduxi in terram pro qua iuravi patribus vestris et pollicitus sum ut non facerem irritum pactum meum vobiscum in sempiternum
JUDG|2|2|ita dumtaxat ut non feriretis foedus cum habitatoribus terrae huius et aras eorum subverteretis et noluistis audire vocem meam cur hoc fecistis
JUDG|2|3|quam ob rem nolui delere eos a facie vestra ut habeatis hostes et dii eorum sint vobis in ruinam
JUDG|2|4|cumque loqueretur angelus Domini verba haec ad omnes filios Israhel elevaverunt vocem suam et fleverunt
JUDG|2|5|et vocatum est nomen loci illius Flentium sive Lacrimarum immolaveruntque ibi hostias Domino
JUDG|2|6|dimisit ergo Iosue populum et abierunt filii Israhel unusquisque in possessionem suam ut obtinerent eam
JUDG|2|7|servieruntque Domino cunctis diebus eius et seniorum qui longo post eum vixerunt tempore et noverant omnia opera Domini quae fecerat cum Israhel
JUDG|2|8|mortuus est autem Iosue filius Nun famulus Domini centum et decem annorum
JUDG|2|9|et sepelierunt eum in finibus possessionis suae in Thamnathsare in monte Ephraim a septentrionali plaga montis Gaas
JUDG|2|10|omnisque illa generatio congregata est ad patres suos et surrexerunt alii qui non noverant Dominum et opera quae fecerat cum Israhel
JUDG|2|11|feceruntque filii Israhel malum in conspectu Domini et servierunt Baalim
JUDG|2|12|ac dimiserunt Dominum Deum patrum suorum qui eduxerat eos de terra Aegypti et secuti sunt deos alienos deos quoque populorum qui habitabant in circuitu eorum et adoraverunt eos et ad iracundiam concitaverunt Dominum
JUDG|2|13|dimittentes eum et servientes Baal et Astharoth
JUDG|2|14|iratusque Dominus contra Israhel tradidit eos in manibus diripientium qui ceperunt eos et vendiderunt hostibus qui habitabant per gyrum nec potuerunt resistere adversariis suis
JUDG|2|15|sed quocumque pergere voluissent manus Domini erat super eos sicut locutus est et iuravit eis et vehementer adflicti sunt
JUDG|2|16|suscitavitque Dominus iudices qui liberarent eos de vastantium manibus sed nec illos audire voluerunt
JUDG|2|17|fornicantes cum diis alienis et adorantes eos cito deseruerunt viam per quam ingressi fuerant patres eorum et audientes mandata Domini omnia fecere contraria
JUDG|2|18|cumque Dominus iudices suscitaret in diebus eorum flectebatur misericordia et audiebat adflictorum gemitus et liberabat eos de caede vastantium
JUDG|2|19|postquam autem mortuus esset iudex revertebantur et multo maiora faciebant quam fecerant patres sui sequentes deos alienos et servientes eis et adorantes illos non dimiserunt adinventiones suas et viam durissimam per quam ambulare consueverant
JUDG|2|20|iratusque est furor Domini in Israhel et ait quia irritum fecit gens ista pactum meum quod pepigeram cum patribus eorum et vocem meam audire contempsit
JUDG|2|21|et ego non delebo gentes quas dimisit Iosue et mortuus est
JUDG|2|22|ut in ipsis experiar Israhel utrum custodiant viam Domini et ambulent in ea sicut custodierunt patres eorum an non
JUDG|2|23|dimisit ergo Dominus omnes has nationes et cito subvertere noluit nec tradidit in manibus Iosue
JUDG|3|1|hae sunt gentes quas Dominus dereliquit ut erudiret in eis Israhelem et omnes qui non noverant bella Chananeorum
JUDG|3|2|et postea discerent filii eorum certare cum hostibus et habere consuetudinem proeliandi
JUDG|3|3|quinque satrapas Philisthinorum omnemque Chananeum et Sidonium atque Eveum qui habitabat in monte Libano de monte Baalhermon usque ad introitum Emath
JUDG|3|4|dimisitque eos ut in ipsis experiretur Israhelem utrum audiret mandata Domini quae praeceperat patribus eorum per manum Mosi an non
JUDG|3|5|itaque filii Israhel habitaverunt in medio Chananei et Hetthei et Amorrei et Ferezei et Evei et Iebusei
JUDG|3|6|et duxerunt uxores filias eorum ipsique filias suas eorum filiis tradiderunt et servierunt diis eorum
JUDG|3|7|feceruntque malum in conspectu Domini et obliti sunt Dei sui servientes Baalim et Astharoth
JUDG|3|8|iratusque Dominus contra Israhel tradidit eos in manus Chusanrasathaim regis Mesopotamiae servieruntque ei octo annis
JUDG|3|9|et clamaverunt ad Dominum qui suscitavit eis salvatorem et liberavit eos Othonihel videlicet filium Cenez fratrem Chaleb minorem
JUDG|3|10|fuitque in eo spiritus Domini et iudicavit Israhel egressusque est ad pugnam et tradidit Dominus in manu eius Chusanrasathaim regem Syriae et oppressit eum
JUDG|3|11|quievitque terra quadraginta annis et mortuus est Othonihel filius Cenez
JUDG|3|12|addiderunt autem filii Israhel facere malum in conspectu Domini qui confortavit adversum eos Eglon regem Moab quia fecerunt malum in conspectu eius
JUDG|3|13|et copulavit ei filios Ammon et Amalech abiitque et percussit Israhel atque possedit urbem Palmarum
JUDG|3|14|servieruntque filii Israhel Eglon regi Moab decem et octo annis
JUDG|3|15|et postea clamaverunt ad Dominum qui suscitavit eis salvatorem vocabulo Ahoth filium Gera filii Iemini qui utraque manu utebatur pro dextera miseruntque filii Israhel per illum munera Eglon regi Moab
JUDG|3|16|qui fecit sibi gladium ancipitem habentem in medio capulum longitudinis palmae manus et accinctus est eo subter sagum in dextro femore
JUDG|3|17|obtulitque munera Eglon regi Moab erat autem Eglon crassus nimis
JUDG|3|18|cumque obtulisset ei munera prosecutus est socios qui cum eo venerant
JUDG|3|19|et reversus de Galgalis ubi erant idola dixit ad regem verbum secretum habeo ad te o rex et ille imperavit silentium egressisque omnibus qui circa eum erant
JUDG|3|20|ingressus est Ahoth ad eum sedebat autem in aestivo cenaculo solus dixitque verbum Dei habeo ad te qui statim surrexit de throno
JUDG|3|21|extenditque Ahoth manum sinistram et tulit sicam de dextro femore suo infixitque eam in ventre eius
JUDG|3|22|tam valide ut capulus ferrum sequeretur in vulnere ac pinguissimo adipe stringeretur nec eduxit gladium sed ita ut percusserat reliquit in corpore statimque per secreta naturae alvi stercora proruperunt
JUDG|3|23|Ahoth autem clausis diligentissime ostiis cenaculi et obfirmatis sera
JUDG|3|24|per posticam egressus est servique regis ingressi viderunt clausas fores cenaculi atque dixerunt forsitan purgat alvum in aestivo cubiculo
JUDG|3|25|expectantesque diu donec erubescerent et videntes quod nullus aperiret tulerunt clavem et aperientes invenerunt dominum suum iacentem in terra mortuum
JUDG|3|26|Ahoth autem dum illi turbarentur effugit et pertransiit locum Idolorum unde reversus fuerat venitque in Seirath
JUDG|3|27|et statim insonuit bucina in monte Ephraim descenderuntque cum eo filii Israhel ipso in fronte gradiente
JUDG|3|28|qui dixit ad eos sequimini me tradidit enim Dominus inimicos nostros Moabitas in manus nostras descenderuntque post eum et occupaverunt vada Iordanis quae transmittunt in Moab et non dimiserunt transire quemquam
JUDG|3|29|sed percusserunt Moabitas in tempore illo circiter decem milia omnes robustos et fortes viros nullus eorum evadere potuit
JUDG|3|30|humiliatusque est Moab die illo sub manu Israhel et quievit terra octoginta annis
JUDG|3|31|post hunc fuit Samgar filius Anath qui percussit de Philisthim sescentos viros vomere et ipse quoque defendit Israhel
JUDG|4|1|addideruntque filii Israhel facere malum in conspectu Domini post mortem Ahoth
JUDG|4|2|et tradidit illos Dominus in manu Iabin regis Chanaan qui regnavit in Asor habuitque ducem exercitus sui nomine Sisaram ipse autem habitabat in Aroseth gentium
JUDG|4|3|clamaveruntque filii Israhel ad Dominum nongentos enim habebat falcatos currus et per viginti annos vehementer oppresserat eos
JUDG|4|4|erat autem Debbora prophetis uxor Lapidoth quae iudicabat populum in illo tempore
JUDG|4|5|et sedebat sub palma quae nomine illius vocabatur inter Rama et Bethel in monte Ephraim ascendebantque ad eam filii Israhel in omne iudicium
JUDG|4|6|quae misit et vocavit Barac filium Abinoem de Cedes Nepthalim dixitque ad eum praecepit tibi Dominus Deus Israhel vade et duc exercitum in montem Thabor tollesque tecum decem milia pugnatorum de filiis Nepthalim et de filiis Zabulon
JUDG|4|7|ego autem ducam ad te in loco torrentis Cison Sisaram principem exercitus Iabin et currus eius atque omnem multitudinem et tradam eos in manu tua
JUDG|4|8|dixitque ad eam Barac si venis mecum vadam si nolueris venire non pergam
JUDG|4|9|quae dixit ad eum ibo quidem tecum sed in hac vice tibi victoria non reputabitur quia in manu mulieris tradetur Sisara surrexit itaque Debbora et perrexit cum Barac in Cedes
JUDG|4|10|qui accitis Zabulon et Nepthalim ascendit cum decem milibus pugnatorum habens Debboram in comitatu suo
JUDG|4|11|Aber autem Cineus recesserat quondam a ceteris Cineis fratribus suis filiis Obab cognati Mosi et tetenderat tabernacula usque ad vallem quae vocatur Sennim et erat iuxta Cedes
JUDG|4|12|nuntiatumque est Sisarae quod ascendisset Barac filius Abinoem in montem Thabor
JUDG|4|13|et congregavit nongentos falcatos currus omnemque exercitum de Aroseth gentium ad torrentem Cison
JUDG|4|14|dixitque Debbora ad Barac surge haec est enim dies in qua tradidit Dominus Sisaram in manus tuas en ipse ductor est tuus descendit itaque Barac de monte Thabor et decem milia pugnatorum cum eo
JUDG|4|15|perterruitque Dominus Sisaram et omnes currus eius universamque multitudinem in ore gladii ad conspectum Barac in tantum ut Sisara de curru desiliens pedibus fugeret
JUDG|4|16|et Barac persequeretur fugientes currus et exercitum usque ad Aroseth gentium et omnis hostium multitudo usque ad internicionem caderet
JUDG|4|17|Sisara autem fugiens pervenit ad tentorium Iahel uxoris Aber Cinei erat enim pax inter Iabin regem Asor et domum Aber Cinei
JUDG|4|18|egressa igitur Iahel in occursum Sisarae dixit ad eum intra ad me domine mi intra ne timeas qui ingressus tabernaculum eius et opertus ab ea pallio
JUDG|4|19|dixit ad eam da mihi obsecro paululum aquae quia valde sitio quae aperuit utrem lactis et dedit ei bibere et operuit illum
JUDG|4|20|dixitque Sisara ad eam sta ante ostium tabernaculi et cum venerit aliquis interrogans te et dicens numquid hic est aliquis respondebis nullus est
JUDG|4|21|tulit itaque Iahel uxor Aber clavum tabernaculi adsumens pariter malleum et ingressa abscondite et cum silentio posuit supra tempus capitis eius clavum percussumque malleo defixit in cerebrum usque ad terram qui soporem morti socians defecit et mortuus est
JUDG|4|22|et ecce Barac sequens Sisaram veniebat egressaque Iahel in occursum eius dixit ei veni et ostendam tibi virum quem quaeris qui cum intrasset ad eam vidit Sisaram iacentem mortuum et clavum infixum in tempore eius
JUDG|4|23|humiliavit ergo Deus in die illo Iabin regem Chanaan coram filiis Israhel
JUDG|4|24|qui crescebant cotidie et forti manu opprimebant Iabin regem Chanaan donec delerent eum
JUDG|5|1|cecineruntque Debbora et Barac filius Abinoem in die illo dicentes
JUDG|5|2|qui sponte obtulistis de Israhel animas vestras ad periculum benedicite Domino
JUDG|5|3|audite reges percipite auribus principes ego sum ego sum quae Domino canam psallam Domino Deo Israhel
JUDG|5|4|Domine cum exires de Seir et transires per regiones Edom terra mota est caelique ac nubes stillaverunt aquis
JUDG|5|5|montes fluxerunt a facie Domini et Sinai a facie Domini Dei Israhel
JUDG|5|6|in diebus Samgar filii Anath in diebus Iahel quieverunt semitae et qui ingrediebantur per eas ambulaverunt per calles devios
JUDG|5|7|cessaverunt fortes in Israhel et quieverunt donec surgeret Debbora surgeret mater in Israhel
JUDG|5|8|nova bella elegit Dominus et portas hostium ipse subvertit clypeus et hasta si apparuerint in quadraginta milibus Israhel
JUDG|5|9|cor meum diligit principes Israhel qui propria voluntate obtulistis vos discrimini benedicite Domino
JUDG|5|10|qui ascenditis super nitentes asinos et sedetis in iudicio et ambulatis in via loquimini
JUDG|5|11|ubi conlisi sunt currus et hostium est suffocatus exercitus ibi narrentur iustitiae Domini et clementia in fortes Israhel tunc descendit populus Domini ad portas et obtinuit principatum
JUDG|5|12|surge surge Debbora surge surge et loquere canticum surge Barac et adprehende captivos tuos fili Abinoem
JUDG|5|13|salvatae sunt reliquiae populi Dominus in fortibus dimicavit
JUDG|5|14|ex Ephraim delevit eos in Amalech et post eum ex Beniamin in populos tuos o Amalech de Machir principes descenderunt et de Zabulon qui exercitum ducerent ad bellandum
JUDG|5|15|duces Isachar fuere cum Debbora et Barac vestigia sunt secuti qui quasi in praeceps ac baratrum se discrimini dedit diviso contra se Ruben magnanimorum repperta contentio est
JUDG|5|16|quare habitas inter duos terminos ut audias sibilos gregum diviso contra se Ruben magnanimorum repperta contentio est
JUDG|5|17|Galaad trans Iordanem quiescebat et Dan vacabat navibus Aser habitabat in litore maris et in portibus morabatur
JUDG|5|18|Zabulon vero et Nepthalim obtulerunt animas suas morti in regione Merome
JUDG|5|19|venerunt reges et pugnaverunt pugnaverunt reges Chanaan in Thanach iuxta aquas Mageddo et tamen nihil tulere praedantes
JUDG|5|20|de caelo dimicatum est contra eos stellae manentes in ordine et cursu suo adversum Sisaram pugnaverunt
JUDG|5|21|torrens Cison traxit cadavera eorum torrens Cadumim torrens Cison conculca anima mea robustos
JUDG|5|22|ungulae equorum ceciderunt fugientibus impetu et per praeceps ruentibus fortissimis hostium
JUDG|5|23|maledicite terrae Meroz dixit angelus Domini maledicite habitatoribus eius quia non venerunt ad auxilium Domini in adiutorium fortissimorum eius
JUDG|5|24|benedicta inter mulieres Iahel uxor Aber Cinei benedicatur in tabernaculo suo
JUDG|5|25|aquam petenti lac dedit et in fiala principum obtulit butyrum
JUDG|5|26|sinistram manum misit ad clavum et dexteram ad fabrorum malleos percussitque Sisaram quaerens in capite vulneri locum et tempus valide perforans
JUDG|5|27|inter pedes eius ruit defecit et mortuus est ante pedes illius volvebatur et iacebat exanimis et miserabilis
JUDG|5|28|per fenestram prospiciens ululabat mater eius et de cenaculo loquebatur cur moratur regredi currus eius quare tardaverunt pedes quadrigarum illius
JUDG|5|29|una sapientior ceteris uxoribus eius haec socrui verba respondit
JUDG|5|30|forsitan nunc dividit spolia et pulcherrima feminarum eligitur ei vestes diversorum colorum Sisarae traduntur in praedam et supellex varia ad ornanda colla congeritur
JUDG|5|31|sic pereant omnes inimici tui Domine qui autem diligunt te sicut sol in ortu suo splendet ita rutilent
JUDG|5|32|quievitque terra per quadraginta annos
JUDG|6|1|fecerunt autem filii Israhel malum in conspectu Domini qui tradidit eos in manu Madian septem annis
JUDG|6|2|et oppressi sunt valde ab eis feceruntque sibi antra et speluncas in montibus et munitissima ad repugnandum loca
JUDG|6|3|cumque sevisset Israhel ascendebat Madian et Amalech et ceteri orientalium nationum
JUDG|6|4|et apud eos figentes tentoria sicut erant in herbis cuncta vastabant usque ad introitum Gazae nihilque omnino ad vitam pertinens relinquebant in Israhel non oves non boves non asinos
JUDG|6|5|ipsi enim et universi greges eorum veniebant cum tabernaculis et instar lucustarum universa conplebant innumera multitudo hominum et camelorum quicquid tetigerant devastantes
JUDG|6|6|humiliatusque est Israhel valde in conspectu Madian
JUDG|6|7|et clamavit ad Dominum postulans auxilium contra Madianitas
JUDG|6|8|qui misit ad eos virum prophetam et locutus est haec dicit Dominus Deus Israhel ego vos feci conscendere de Aegypto et eduxi de domo servitutis
JUDG|6|9|et liberavi de manu Aegyptiorum et omnium inimicorum qui adfligebant vos eiecique eos ad introitum vestrum et tradidi vobis terram eorum
JUDG|6|10|et dixi ego Dominus Deus vester ne timeatis deos Amorreorum in quorum terra habitatis et noluistis audire vocem meam
JUDG|6|11|venit autem angelus Domini et sedit sub quercu quae erat in Ephra et pertinebat ad Ioas patrem familiae Ezri cumque Gedeon filius eius excuteret atque purgaret frumenta in torculari ut fugeret Madian
JUDG|6|12|apparuit ei et ait Dominus tecum virorum fortissime
JUDG|6|13|dixitque ei Gedeon obsecro Domine si Dominus nobiscum est cur adprehenderunt nos haec omnia ubi sunt mirabilia eius quae narraverunt patres nostri atque dixerunt de Aegypto eduxit nos Dominus nunc autem dereliquit nos et tradidit in manibus Madian
JUDG|6|14|respexitque ad eum Dominus et ait vade in hac fortitudine tua et liberabis Israhel de manu Madian scito quod miserim te
JUDG|6|15|qui respondens ait obsecro Domine mi in quo liberabo Israhel ecce familia mea infima est in Manasse et ego minimus in domo patris mei
JUDG|6|16|dixitque ei Dominus ego ero tecum et percuties Madian quasi unum virum
JUDG|6|17|et ille si inveni inquit gratiam coram te da mihi signum quod tu sis qui loquaris ad me
JUDG|6|18|ne recedas hinc donec revertar ad te portans sacrificium et offerens tibi qui respondit ego praestolabor adventum tuum
JUDG|6|19|ingressus est itaque Gedeon et coxit hedum et de farinae modio azymos panes carnesque ponens in canistro et ius carnium mittens in ollam tulit omnia sub quercum et obtulit ei
JUDG|6|20|cui dixit angelus Domini tolle carnes et panes azymos et pone super petram illam et ius desuper funde cumque fecisset ita
JUDG|6|21|extendit angelus Domini summitatem virgae quam tenebat in manu et tetigit carnes et azymos panes ascenditque ignis de petra et carnes azymosque consumpsit angelus autem Domini evanuit ex oculis eius
JUDG|6|22|vidensque Gedeon quod esset angelus Domini ait heu mihi Domine Deus quia vidi angelum Domini facie ad faciem
JUDG|6|23|dixitque ei Dominus pax tecum ne timeas non morieris
JUDG|6|24|aedificavit ergo ibi Gedeon altare Domino vocavitque illud Domini pax usque in praesentem diem cum adhuc esset in Ephra quae est familiae Ezri
JUDG|6|25|nocte illa dixit Dominus ad eum tolle taurum patris tui et alterum taurum annorum septem destruesque aram Baal quae est patris tui et nemus quod circa aram est succide
JUDG|6|26|et aedificabis altare Domino Deo tuo in summitate petrae huius super quam sacrificium ante posuisti tollesque taurum secundum et offeres holocaustum super lignorum struem quae de nemore succideris
JUDG|6|27|adsumptis igitur Gedeon decem viris de servis suis fecit sicut praeceperat Dominus timens autem domum patris sui et homines illius civitatis per diem facere noluit sed omnia nocte conplevit
JUDG|6|28|cumque surrexissent viri oppidi eius mane viderunt destructam aram Baal lucumque succisum et taurum alterum inpositum super altare quod tunc aedificatum erat
JUDG|6|29|dixeruntque ad invicem quis hoc fecit cumque perquirerent auctorem facti dictum est Gedeon filius Ioas fecit haec omnia
JUDG|6|30|et dixerunt ad Ioas produc filium tuum ut moriatur quia destruxit aram Baal et succidit nemus
JUDG|6|31|quibus ille respondit numquid ultores estis Baal et pugnatis pro eo qui adversarius eius est moriatur antequam lux crastina veniat si deus est vindicet se de eo qui suffodit aram eius
JUDG|6|32|ex illo die vocatus est Gedeon Hierobbaal eo quod dixisset Ioas ulciscatur se de eo Baal qui suffodit altare eius
JUDG|6|33|igitur omnis Madian et Amalech et orientales populi congregati sunt simul et transeuntes Iordanem castrametati sunt in valle Iezrahel
JUDG|6|34|spiritus autem Domini induit Gedeon qui clangens bucina convocavit domum Abiezer ut sequeretur
JUDG|6|35|misitque nuntios in universum Manassen qui et ipse secutus est eum et alios nuntios in Aser et Zabulon et Nepthalim qui occurrerunt ei
JUDG|6|36|dixitque Gedeon ad Dominum si salvum facis per manum meam Israhel sicut locutus es
JUDG|6|37|ponam vellus hoc lanae in area si ros in solo vellere fuerit et in omni terra siccitas sciam quod per manum meam sicut locutus es liberabis Israhel
JUDG|6|38|factumque est ita et de nocte consurgens expresso vellere concam rore conplevit
JUDG|6|39|dixitque rursus ad Dominum ne irascatur furor tuus contra me si adhuc semel temptavero signum quaerens in vellere oro ut solum vellus siccum sit et omnis terra rore madens
JUDG|6|40|fecitque Dominus nocte illa ut postulaverat et fuit siccitas in solo vellere et ros in omni terra
JUDG|7|1|igitur Hierobbaal qui est et Gedeon de nocte consurgens et omnis populus cum eo venit ad fontem qui vocatur Arad erant autem castra Madian in valle ad septentrionalem plagam collis Excelsi
JUDG|7|2|dixitque Dominus ad Gedeon multus tecum est populus nec tradetur Madian in manus eius ne glorietur contra me Israhel et dicat meis viribus liberatus sum
JUDG|7|3|loquere ad populum et cunctis audientibus praedica qui formidolosus et timidus est revertatur recesseruntque de monte Galaad et reversa sunt ex populo viginti duo milia virorum et tantum decem milia remanserunt
JUDG|7|4|dixitque Dominus ad Gedeon adhuc populus multus est duc eos ad aquas et ibi probabo illos et de quo dixero tibi ut tecum vadat ipse pergat quem ire prohibuero revertatur
JUDG|7|5|cumque descendisset populus ad aquas dixit Dominus ad Gedeon qui lingua lambuerint aquas sicut solent canes lambere separabis eos seorsum qui autem curvatis genibus biberint in altera parte erunt
JUDG|7|6|fuit itaque numerus eorum qui manu ad os proiciente aquas lambuerant trecenti viri omnis autem reliqua multitudo flexo poplite biberat
JUDG|7|7|et ait Dominus ad Gedeon in trecentis viris qui lambuerunt aquas liberabo vos et tradam Madian in manu tua omnis autem reliqua multitudo revertatur in locum suum
JUDG|7|8|sumptis itaque pro numero cibariis et tubis omnem reliquam multitudinem abire praecepit ad tabernacula sua et ipse cum trecentis viris se certamini dedit castra autem Madian erant subter in valle
JUDG|7|9|eadem nocte dixit Dominus ad eum surge et descende in castra quia tradidi eos in manu tua
JUDG|7|10|sin autem solus ire formidas descendat tecum Phara puer tuus
JUDG|7|11|et cum audieris quid loquantur tunc confortabuntur manus tuae et securior ad hostium castra descendes descendit ergo ipse et Phara puer eius in partem castrorum ubi erant armatorum vigiliae
JUDG|7|12|Madian autem et Amalech et omnes orientales populi fusi iacebant in valle ut lucustarum multitudo cameli quoque innumerabiles erant sicut harena quae iacet in litoribus maris
JUDG|7|13|cumque venisset Gedeon narrabat aliquis somnium proximo suo et in hunc modum referebat quod viderat vidi somnium et videbatur mihi quasi subcinericius panis ex hordeo volvi et in Madian castra descendere cumque pervenisset ad tabernaculum percussit illud atque subvertit et terrae funditus coaequavit
JUDG|7|14|respondit is cui loquebatur non est hoc aliud nisi gladius Gedeonis filii Ioas viri Israhelitae tradidit Deus in manu eius Madian et omnia castra eius
JUDG|7|15|cumque audisset Gedeon somnium et interpretationem eius adoravit et reversus ad castra Israhel ait surgite tradidit enim Dominus in manus nostras castra Madian
JUDG|7|16|divisitque trecentos viros in tres partes et dedit tubas in manibus eorum lagoenasque vacuas ac lampadas in medio lagoenarum
JUDG|7|17|et dixit ad eos quod me facere videritis hoc facite ingrediar partem castrorum et quod fecero sectamini
JUDG|7|18|quando personaverit tuba in manu mea vos quoque per castrorum circuitum clangite et conclamate Domino et Gedeoni
JUDG|7|19|ingressusque est Gedeon et trecenti viri qui erant cum eo in parte castrorum incipientibus vigiliis noctis mediae et custodibus suscitatis coeperunt bucinis clangere et conplodere inter se lagoenas
JUDG|7|20|cumque per gyrum castrorum in tribus personarent locis et hydrias confregissent tenuerunt sinistris manibus lampadas et dextris sonantes tubas clamaveruntque gladius Domini et Gedeonis
JUDG|7|21|stantes singuli in loco suo per circuitum castrorum hostilium omnia itaque castra turbata sunt et vociferantes ululantesque fugerunt
JUDG|7|22|et nihilominus insistebant trecenti viri bucinis personantes inmisitque Dominus gladium in omnibus castris et mutua se caede truncabant
JUDG|7|23|fugientes usque Bethseta et crepidinem Abelmeula in Tebbath conclamantes autem viri Israhel de Nepthali et Aser et omni Manasse persequebantur Madian
JUDG|7|24|misitque Gedeon nuntios in omnem montem Ephraim dicens descendite in occursum Madian et occupate aquas usque Bethbera atque Iordanem clamavitque omnis Ephraim et praeoccupavit aquas atque Iordanem usque Bethbera
JUDG|7|25|adprehensosque duos viros Madian Oreb et Zeb interfecit Oreb in petra Oreb Zeb vero in torculari Zeb et persecuti sunt Madian capita Oreb et Zeb portantes ad Gedeon trans fluenta Iordanis
JUDG|8|1|dixeruntque ad eum viri Ephraim quid est hoc quod facere voluisti ut non nos vocares cum ad pugnam pergeres contra Madian iurgantes fortiter et prope vim inferentes
JUDG|8|2|quibus ille respondit quid enim tale facere potui quale vos fecistis nonne melior est racemus Ephraim vindemiis Abiezer
JUDG|8|3|in manus vestras tradidit Dominus principes Madian Oreb et Zeb quid tale facere potui quale vos fecistis quod cum locutus esset requievit spiritus eorum quo tumebant contra eum
JUDG|8|4|cumque venisset Gedeon ad Iordanem transivit eum cum trecentis viris qui secum erant et prae lassitudine fugientes persequi non poterant
JUDG|8|5|dixitque ad viros Soccoth date obsecro panes populo qui mecum est quia valde defecerunt ut possimus persequi Zebee et Salmana reges Madian
JUDG|8|6|responderunt principes Soccoth forsitan palmae manuum Zebee et Salmana in manu tua sunt et idcirco postulas ut demus exercitui tuo panes
JUDG|8|7|quibus ille ait cum ergo tradiderit Dominus Zebee et Salmana in manus meas conteram carnes vestras cum spinis tribulisque deserti
JUDG|8|8|et inde conscendens venit in Phanuhel locutusque est ad viros eius loci similia cui et illi responderunt sicut responderant viri Soccoth
JUDG|8|9|dixit itaque et eis cum reversus fuero victor in pace destruam turrem hanc
JUDG|8|10|Zebee autem et Salmana requiescebant cum omni exercitu suo quindecim milia enim viri remanserant ex omnibus turmis orientalium populorum caesis centum viginti milibus bellatorum et educentium gladium
JUDG|8|11|ascendensque Gedeon per viam eorum qui in tabernaculis morabantur ad orientalem partem Nobee et Iecbaa percussit castra hostium qui securi erant et nihil adversi suspicabantur
JUDG|8|12|fugeruntque Zebee et Salmana quos persequens Gedeon conprehendit turbato omni exercitu eorum
JUDG|8|13|revertensque de bello ante solis ortum
JUDG|8|14|adprehendit puerum de viris Soccoth interrogavitque eum nomina principum et seniorum Soccoth et descripsit septuaginta septem viros
JUDG|8|15|venitque ad Soccoth et dixit eis en Zebee et Salmana super quibus exprobrastis mihi dicentes forsitan manus Zebee et Salmana in manibus tuis sunt et idcirco postulas ut demus viris qui lassi sunt et defecerunt panes
JUDG|8|16|tulit ergo seniores civitatis et spinas deserti ac tribulos et contrivit cum eis atque comminuit viros Soccoth
JUDG|8|17|turrem quoque Phanuhel subvertit occisis habitatoribus civitatis
JUDG|8|18|dixitque ad Zebee et Salmana quales fuerunt viri quos occidistis in Thabor qui responderunt similes tui et unus ex eis quasi filius regis
JUDG|8|19|quibus ille ait fratres mei fuerunt filii matris meae vivit Dominus si servassetis eos non vos occiderem
JUDG|8|20|dixitque Ietther primogenito suo surge et interfice eos qui non eduxit gladium timebat enim quia adhuc puer erat
JUDG|8|21|dixeruntque Zebee et Salmana tu surge et inrue in nos quia iuxta aetatem robur est hominis surrexit Gedeon et interfecit Zebee et Salmana et tulit ornamenta ac bullas quibus colla regalium camelorum decorari solent
JUDG|8|22|dixeruntque omnes viri Israhel ad Gedeon dominare nostri tu et filius tuus et filius filii tui quia liberasti nos de manu Madian
JUDG|8|23|quibus ille ait non dominabor vestri nec dominabitur in vos filius meus sed dominabitur Dominus
JUDG|8|24|dixitque ad eos unam petitionem postulo a vobis date mihi inaures ex praeda vestra inaures enim aureas Ismahelitae habere consuerant
JUDG|8|25|qui responderunt libentissime dabimus expandentesque super terram pallium proiecerunt in eo inaures de praeda
JUDG|8|26|et fuit pondus postulatarum inaurium mille septingenti auri sicli absque ornamentis et monilibus et veste purpurea quibus Madian reges uti soliti erant et praeter torques aureos camelorum
JUDG|8|27|fecitque ex eo Gedeon ephod et posuit illud in civitate sua Ephra fornicatusque est omnis Israhel in eo et factum est Gedeoni et omni domui eius in ruinam
JUDG|8|28|humiliatus est autem Madian coram filiis Israhel nec potuerunt ultra elevare cervices sed quievit terra per quadraginta annos quibus praefuit Gedeon
JUDG|8|29|abiit itaque Hierobbaal filius Ioas et habitavit in domo sua
JUDG|8|30|habuitque septuaginta filios qui egressi sunt de femore eius eo quod plures haberet uxores
JUDG|8|31|concubina autem illius quam habebat in Sychem genuit ei filium nomine Abimelech
JUDG|8|32|mortuusque est Gedeon filius Ioas in senectute bona et sepultus in sepulchro Ioas patris sui in Ephra de familia Ezri
JUDG|8|33|postquam autem mortuus est Gedeon aversi sunt filii Israhel et fornicati cum Baalim percusseruntque cum Baal foedus ut esset eis in deum
JUDG|8|34|nec recordati sunt Domini Dei sui qui eruit eos de manu omnium inimicorum suorum per circuitum
JUDG|8|35|nec fecerunt misericordiam cum domo Hierobbaal Gedeon iuxta omnia bona quae fecerat Israheli
JUDG|9|1|abiit autem Abimelech filius Hierobbaal in Sychem ad fratres matris suae et locutus est ad eos et ad omnem cognationem domus patris matris suae dicens
JUDG|9|2|loquimini ad omnes viros Sychem quid vobis est melius ut dominentur vestri septuaginta viri omnes filii Hierobbaal an ut dominetur vobis unus vir simulque considerate quia os vestrum et caro vestra sum
JUDG|9|3|locutique sunt fratres matris eius de eo ad omnes viros Sychem universos sermones istos et inclinaverunt cor eorum post Abimelech dicentes frater noster est
JUDG|9|4|dederuntque illi septuaginta pondo argenti de fano Baalbrith qui conduxit sibi ex eo viros inopes et vagos secutique sunt eum
JUDG|9|5|et venit in domum patris sui Ephra et occidit fratres suos filios Hierobbaal septuaginta viros super lapidem unum remansitque Ioatham filius Hierobbaal minimus et absconditus est
JUDG|9|6|congregati sunt autem omnes viri Sychem et universae familiae urbis Mello abieruntque et constituerunt regem Abimelech iuxta quercum quae stabat in Sychem
JUDG|9|7|quod cum nuntiatum esset Ioatham ivit et stetit in vertice montis Garizim elevataque voce clamavit et dixit audite me viri Sychem ita audiat vos Deus
JUDG|9|8|ierunt ligna ut unguerent super se regem dixeruntque olivae impera nobis
JUDG|9|9|quae respondit numquid possum deserere pinguedinem meam qua et dii utuntur et homines et venire ut inter ligna promovear
JUDG|9|10|dixeruntque ligna ad arborem ficum veni et super nos regnum accipe
JUDG|9|11|quae respondit eis numquid possum deserere dulcedinem meam fructusque suavissimos et ire ut inter cetera ligna commovear
JUDG|9|12|locuta sunt quoque ligna ad vitem veni et impera nobis
JUDG|9|13|quae respondit numquid possum deserere vinum meum quod laetificat Deum et homines et inter ligna cetera commoveri
JUDG|9|14|dixeruntque omnia ligna ad ramnum veni et impera super nos
JUDG|9|15|quae respondit eis si vere me regem vobis constituitis venite et sub mea umbra requiescite sin autem non vultis egrediatur ignis de ramno et devoret cedros Libani
JUDG|9|16|nunc igitur si recte et absque peccato constituistis super vos regem Abimelech et bene egistis cum Hierobbaal et cum domo eius et reddidistis vicem beneficiis eius qui pugnavit pro vobis
JUDG|9|17|et animam suam dedit periculis ut erueret vos de manu Madian
JUDG|9|18|qui nunc surrexistis contra domum patris mei et interfecistis filios eius septuaginta viros super unum lapidem et constituistis regem Abimelech filium ancillae eius super habitatores Sychem eo quod frater vester sit
JUDG|9|19|si ergo recte et absque vitio egistis cum Hierobbaal et domo eius hodie laetamini in Abimelech et ille laetetur in vobis
JUDG|9|20|sin autem perverse egrediatur ignis ex eo et consumat habitatores Sychem et oppidum Mello egrediaturque ignis de viris Sychem et de oppido Mello et devoret Abimelech
JUDG|9|21|quae cum dixisset fugit et abiit in Bera habitavitque ibi metu Abimelech fratris sui
JUDG|9|22|regnavit itaque Abimelech super Israhel tribus annis
JUDG|9|23|misitque Deus spiritum pessimum inter Abimelech et habitatores Sychem qui coeperunt eum detestari
JUDG|9|24|et scelus interfectionis septuaginta filiorum Hierobbaal et effusionem sanguinis eorum conferre in Abimelech fratrem suum et in ceteros Sycimarum principes qui eum adiuverant
JUDG|9|25|posueruntque insidias adversum eum in montium summitate et dum illius praestolantur adventum exercebant latrocinia agentes praedas de praetereuntibus nuntiatumque est Abimelech
JUDG|9|26|venit autem Gaal filius Obed cum fratribus suis et transivit in Sycimam ad cuius adventum erecti habitatores Sychem
JUDG|9|27|egressi sunt in agros vastantes vineas uvasque calcantes et factis cantantium choris ingressi sunt fanum dei sui et inter epulas et pocula maledicebant Abimelech
JUDG|9|28|clamante Gaal filio Obed quis est Abimelech et quae est Sychem ut serviamus ei numquid non est filius Hierobbaal et constituit principem Zebul servum suum super viros Emmor patris Sychem cur igitur servimus ei
JUDG|9|29|utinam daret aliquis populum istum sub manu mea ut auferrem de medio Abimelech dictumque est Abimelech congrega exercitus multitudinem et veni
JUDG|9|30|Zebul enim princeps civitatis auditis sermonibus Gaal filii Obed iratus est valde
JUDG|9|31|et misit clam ad Abimelech nuntios dicens ecce Gaal filius Obed venit in Sycimam cum fratribus suis et obpugnat adversum te civitatem
JUDG|9|32|surge itaque nocte cum populo qui tecum est et latita in agro
JUDG|9|33|et primo mane oriente sole inrue super civitatem illo autem egrediente adversum te cum populo suo fac ei quod potueris
JUDG|9|34|surrexit itaque Abimelech cum omni exercitu suo nocte et tetendit insidias iuxta Sycimam in quattuor locis
JUDG|9|35|egressusque est Gaal filius Obed et stetit in introitu portae civitatis surrexit autem Abimelech et omnis exercitus cum eo de insidiarum loco
JUDG|9|36|cumque vidisset populum Gaal dixit ad Zebul ecce de montibus multitudo descendit cui ille respondit umbras montium vides quasi hominum capita et hoc errore deciperis
JUDG|9|37|rursumque Gaal ait ecce populus de umbilico terrae descendit et unus cuneus venit per viam quae respicit quercum
JUDG|9|38|cui dixit Zebul ubi est nunc os tuum quo loquebaris quis est Abimelech ut serviamus ei nonne iste est populus quem despiciebas egredere et pugna contra eum
JUDG|9|39|abiit ergo Gaal spectante Sycimarum populo et pugnavit contra Abimelech
JUDG|9|40|qui persecutus est eum fugientem et in urbem conpulit cecideruntque ex parte eius plurimi usque ad portam civitatis
JUDG|9|41|et Abimelech sedit in Ruma Zebul autem Gaal et socios eius expulit de urbe nec in ea passus est commorari
JUDG|9|42|sequenti ergo die egressus est populus in campum quod cum nuntiatum esset Abimelech
JUDG|9|43|tulit exercitum suum et divisit in tres turmas tendens insidias in agris vidensque quod egrederetur populus de civitate surrexit et inruit in eos
JUDG|9|44|cum cuneo suo obpugnans et obsidens civitatem duae autem turmae palantes per campum adversarios sequebantur
JUDG|9|45|porro Abimelech omni illo die obpugnabat urbem quam cepit interfectis habitatoribus eius ipsaque destructa ita ut sal in ea dispergeret
JUDG|9|46|quod cum audissent qui habitabant in turre Sycimorum ingressi sunt fanum dei sui Berith ubi foedus cum eo pepigerant et ex eo locus nomen acceperat qui erat valde munitus
JUDG|9|47|Abimelech quoque audiens viros turris Sycimorum pariter conglobatos
JUDG|9|48|ascendit in montem Selmon cum omni populo suo et arrepta securi praecidit arboris ramum inpositumque ferens umero dixit ad socios quod me vidistis facere cito facite
JUDG|9|49|igitur certatim ramos de arboribus praecidentes sequebantur ducem quos circumdantes praesidio succenderunt atque ita factum est ut fumo et igne mille hominum necarentur viri pariter ac mulieres habitatorum turris Sychem
JUDG|9|50|Abimelech autem inde proficiscens venit ad oppidum Thebes quod circumdans obsidebat exercitu
JUDG|9|51|erat autem turris excelsa in media civitate ad quam confugerant viri simul ac mulieres et omnes principes civitatis clausa firmissime ianua et super turris tectum stantes per propugnacula
JUDG|9|52|accedensque Abimelech iuxta turrem pugnabat fortiter et adpropinquans ostio ignem subponere nitebatur
JUDG|9|53|et ecce una mulier fragmen molae desuper iaciens inlisit capiti Abimelech et confregit cerebrum eius
JUDG|9|54|qui vocavit cito armigerum suum et ait ad eum evagina gladium tuum et percute me ne forte dicatur quod a femina interfectus sim qui iussa perficiens interfecit eum
JUDG|9|55|illoque mortuo omnes qui cum eo erant de Israhel reversi sunt in sedes suas
JUDG|9|56|et reddidit Deus malum quod fecerat Abimelech contra patrem suum interfectis septuaginta fratribus suis
JUDG|9|57|Sycimitis quoque quod operati erant retributum est et venit super eos maledictio Ioatham filii Hierobbaal
JUDG|10|1|post Abimelech surrexit dux in Israhel Thola filius Phoa patrui Abimelech vir de Isachar qui habitavit in Sanir montis Ephraim
JUDG|10|2|et iudicavit Israhel viginti et tribus annis mortuusque ac sepultus est in Sanir
JUDG|10|3|huic successit Iair Galaadites qui iudicavit Israhel per viginti et duos annos
JUDG|10|4|habens triginta filios sedentes super triginta pullos asinarum et principes triginta civitatum quae ex nomine eius appellatae sunt Avothiair id est oppida Iair usque in praesentem diem in terra Galaad
JUDG|10|5|mortuusque est Iair ac sepultus in loco cui est vocabulum Camon
JUDG|10|6|filii autem Israhel peccatis veteribus iungentes nova fecerunt malum in conspectu Domini et servierunt idolis Baalim et Astharoth et diis Syriae ac Sidonis et Moab et filiorum Ammon et Philisthim dimiseruntque Dominum et non colebant eum
JUDG|10|7|contra quos iratus tradidit eos in manu Philisthim et filiorum Ammon
JUDG|10|8|adflictique sunt et vehementer oppressi per annos decem et octo omnes qui habitabant trans Iordanem in terra Amorrei quae est in Galaad
JUDG|10|9|in tantum ut filii Ammon Iordane transmisso vastarent Iudam et Beniamin et Ephraim adflictusque est Israhel nimis
JUDG|10|10|et clamantes ad Dominum dixerunt peccavimus tibi quia dereliquimus Deum nostrum et servivimus Baalim
JUDG|10|11|quibus locutus est Dominus numquid non Aegyptii et Amorrei filiique Ammon et Philisthim
JUDG|10|12|Sidonii quoque et Amalech et Chanaan oppresserunt vos et clamastis ad me et erui vos de manu eorum
JUDG|10|13|et tamen reliquistis me et coluistis deos alienos idcirco non addam ut ultra vos liberem
JUDG|10|14|ite et invocate deos quos elegistis ipsi vos liberent in tempore angustiae
JUDG|10|15|dixeruntque filii Israhel ad Dominum peccavimus redde tu nobis quicquid tibi placet tantum nunc libera nos
JUDG|10|16|quae dicentes omnia de finibus suis alienorum deorum idola proiecerunt et servierunt Deo qui doluit super miseriis eorum
JUDG|10|17|itaque filii Ammon conclamantes in Galaad fixere tentoria contra quos congregati filii Israhel in Maspha castrametati sunt
JUDG|10|18|dixeruntque principes Galaad singuli ad proximos suos qui primus e nobis contra filios Ammon coeperit dimicare erit dux populi Galaad
JUDG|11|1|fuit illo tempore Iepthae Galaadites vir fortissimus atque pugnator filius meretricis mulieris qui natus est de Galaad
JUDG|11|2|habuit autem Galaad uxorem de qua suscepit filios qui postquam creverant eiecerunt Iepthae dicentes heres in domo patris nostri esse non poteris quia de altera matre generatus es
JUDG|11|3|quos ille fugiens atque devitans habitavit in terra Tob congregatique sunt ad eum viri inopes et latrocinantes et quasi principem sequebantur
JUDG|11|4|in illis diebus pugnabant filii Ammon contra Israhel
JUDG|11|5|quibus acriter instantibus perrexerunt maiores natu de Galaad ut tollerent in auxilium sui Iepthae de terra Tob
JUDG|11|6|dixeruntque ad eum veni et esto princeps noster et pugna contra filios Ammon
JUDG|11|7|quibus ille respondit nonne vos estis qui odistis me et eiecistis de domo patris mei et nunc venistis ad me necessitate conpulsi
JUDG|11|8|dixeruntque principes Galaad ad Iepthae ob hanc igitur causam nunc ad te venimus ut proficiscaris nobiscum et pugnes contra filios Ammon sisque dux omnium qui habitant in Galaad
JUDG|11|9|Iepthae quoque dixit eis si vere venistis ad me ut pugnem pro vobis contra filios Ammon tradideritque eos Dominus in manus meas ego ero princeps vester
JUDG|11|10|qui responderunt ei Dominus qui haec audit ipse mediator ac testis est quod nostra promissa faciamus
JUDG|11|11|abiit itaque Iepthae cum principibus Galaad fecitque eum omnis populus principem sui locutusque est Iepthae omnes sermones suos coram Domino in Maspha
JUDG|11|12|et misit nuntios ad regem filiorum Ammon qui ex persona sua dicerent quid mihi et tibi est quia venisti contra me ut vastares terram meam
JUDG|11|13|quibus ille respondit quia tulit Israhel terram meam quando ascendit de Aegypto a finibus Arnon usque Iaboc atque Iordanem nunc igitur cum pace redde mihi eam
JUDG|11|14|per quos rursum mandavit Iepthae et imperavit eis ut dicerent regi Ammon
JUDG|11|15|haec dicit Iepthae non tulit Israhel terram Moab nec terram filiorum Ammon
JUDG|11|16|sed quando de Aegypto conscenderunt ambulavit per solitudinem usque ad mare Rubrum et venit in Cades
JUDG|11|17|misitque nuntios ad regem Edom dicens dimitte ut transeam per terram tuam qui noluit adquiescere precibus eius misit quoque et ad regem Moab qui et ipse transitum praebere contempsit mansit itaque in Cades
JUDG|11|18|et circuivit ex latere terram Edom et terram Moab venitque contra orientalem plagam terrae Moab et castrametatus est trans Arnon nec voluit intrare terminos Moab Arnon quippe confinium est terrae Moab
JUDG|11|19|misit itaque Israhel nuntios ad Seon regem Amorreorum qui habitabat in Esebon et dixerunt ei dimitte ut transeam per terram tuam usque ad fluvium
JUDG|11|20|qui et ipse Israhel verba despiciens non dimisit eum transire per terminos suos sed infinita multitudine congregata egressus est contra eum in Iassa et fortiter resistebat
JUDG|11|21|tradiditque eum Dominus in manu Israhel cum omni exercitu suo qui percussit eum et possedit omnem terram Amorrei habitatoris regionis illius
JUDG|11|22|et universos fines eius de Arnon usque Iaboc et de solitudine usque ad Iordanem
JUDG|11|23|Dominus ergo Deus Israhel subvertit Amorreum pugnante contra illum populo suo Israhel et tu nunc vis possidere terram eius
JUDG|11|24|nonne ea quae possedit Chamos deus tuus tibi iure debentur quae autem Dominus Deus noster victor obtinuit in nostram cedent possessionem
JUDG|11|25|nisi forte melior es Balac filio Sepphor rege Moab aut docere potes quod iurgatus sit contra Israhel et pugnaverit contra eum
JUDG|11|26|quando habitavit in Esebon et viculis eius et in Aroer et villis illius vel in cunctis civitatibus iuxta Iordanem per trecentos annos quare tanto tempore nihil super hac repetitione temptastis
JUDG|11|27|igitur non ego pecco in te sed tu contra me male agis indicens mihi bella non iusta iudicet Dominus arbiter huius diei inter Israhel et inter filios Ammon
JUDG|11|28|noluitque adquiescere rex filiorum Ammon verbis Iepthae quae per nuntios mandaverat
JUDG|11|29|factus est ergo super Iepthae spiritus Domini et circumiens Galaad et Manasse Maspha quoque Galaad et inde transiens ad filios Ammon
JUDG|11|30|votum vovit Domino dicens si tradideris filios Ammon in manus meas
JUDG|11|31|quicumque primus fuerit egressus de foribus domus meae mihique occurrerit revertenti cum pace a filiis Ammon eum holocaustum offeram Domino
JUDG|11|32|transivitque Iepthae ad filios Ammon ut pugnaret contra eos quos tradidit Dominus in manus eius
JUDG|11|33|percussitque ab Aroer usque dum venias in Mennith viginti civitates et usque ad Abel quae est vineis consita plaga magna nimis humiliatique sunt filii Ammon a filiis Israhel
JUDG|11|34|revertenti autem Iepthae in Maspha domum suam occurrit unigenita filia cum tympanis et choris non enim habebat alios liberos
JUDG|11|35|qua visa scidit vestimenta sua et ait heu filia mi decepisti me et ipsa decepta es aperui enim os meum ad Dominum et aliud facere non potero
JUDG|11|36|cui illa respondit pater mi si aperuisti os tuum ad Dominum fac mihi quodcumque pollicitus es concessa tibi ultione atque victoria de hostibus tuis
JUDG|11|37|dixitque ad patrem hoc solum mihi praesta quod deprecor dimitte me ut duobus mensibus circumeam montes et plangam virginitatem meam cum sodalibus meis
JUDG|11|38|cui ille respondit vade et dimisit eam duobus mensibus cumque abisset cum sociis ac sodalibus suis flebat virginitatem suam in montibus
JUDG|11|39|expletisque duobus mensibus reversa est ad patrem suum et fecit ei sicut voverat quae ignorabat virum exinde mos increbuit in Israhel et consuetudo servata est
JUDG|11|40|ut post anni circulum conveniant in unum filiae Israhel et plangant filiam Iepthae Galaaditae diebus quattuor
JUDG|12|1|ecce autem in Ephraim orta seditio est nam transeuntes contra aquilonem dixerunt ad Iepthae quare vadens ad pugnam contra filios Ammon vocare nos noluisti ut pergeremus tecum igitur incendimus domum tuam
JUDG|12|2|quibus ille respondit disceptatio erat mihi et populo meo contra filios Ammon vehemens vocavique vos ut mihi praeberetis auxilium et facere noluistis
JUDG|12|3|quod cernens posui in manibus meis animam meam transivique ad filios Ammon et tradidit eos Dominus in manus meas quid commerui ut adversum me consurgatis in proelium
JUDG|12|4|vocatis itaque ad se cunctis viris Galaad pugnabat contra Ephraim percusseruntque viri Galaad Ephraim quia dixerat fugitivus est Galaad de Ephraim et habitat in medio Ephraim et Manasse
JUDG|12|5|occupaveruntque Galaaditae vada Iordanis per quae Ephraim reversurus erat cumque venisset ad ea de Ephraim numero fugiens atque dixisset obsecro ut me transire permittas dicebant ei Galaaditae numquid Ephrateus es quo dicente non sum
JUDG|12|6|interrogabant eum dic ergo sebboleth quod interpretatur spica qui respondebat tebboleth eadem littera spicam exprimere non valens statimque adprehensum iugulabant in ipso Iordanis transitu et ceciderunt in illo tempore de Ephraim quadraginta duo milia
JUDG|12|7|iudicavitque Iepthae Galaadites Israhel sex annis et mortuus est ac sepultus in civitate sua Galaad
JUDG|12|8|post hunc iudicavit Israhel Abessan de Bethleem
JUDG|12|9|qui habuit triginta filios et totidem filias quas emittens foras maritis dedit et eiusdem numeri filiis suis accepit uxores introducens in domum suam qui septem annis iudicavit Israhel
JUDG|12|10|mortuusque est ac sepultus in Bethleem
JUDG|12|11|cui successit Ahialon Zabulonites et iudicavit Israhelem decem annis
JUDG|12|12|mortuusque est ac sepultus in Zabulon
JUDG|12|13|post hunc iudicavit in Israhel Abdon filius Hellel Farathonites
JUDG|12|14|qui habuit quadraginta filios et triginta ex eis nepotes ascendentes super septuaginta pullos asinarum et iudicavit in Israhel octo annis
JUDG|12|15|mortuusque est ac sepultus in Farathon terrae Ephraim in monte Amalech
JUDG|13|1|rursumque filii Israhel fecerunt malum in conspectu Domini qui tradidit eos in manus Philisthinorum quadraginta annis
JUDG|13|2|erat autem vir quidam de Saraa et de stirpe Dan nomine Manue habens uxorem sterilem
JUDG|13|3|cui apparuit angelus Domini et dixit ad eam sterilis es et absque liberis sed concipies et paries filium
JUDG|13|4|cave ergo ne vinum bibas ac siceram ne inmundum quicquam comedas
JUDG|13|5|quia concipies et paries filium cuius non tanget caput novacula erit enim nazareus Dei ab infantia sua et ex matris utero et ipse incipiet liberare Israhel de manu Philisthinorum
JUDG|13|6|quae cum venisset ad maritum dixit ei vir Dei venit ad me habens vultum angelicum terribilis nimis quem cum interrogassem quis esset et unde venisset et quo nomine vocaretur noluit mihi dicere
JUDG|13|7|sed hoc respondit ecce concipies et paries filium cave ne vinum bibas et siceram et ne aliquo vescaris inmundo erit enim puer nazareus Dei ab infantia sua et ex utero matris usque ad diem mortis suae
JUDG|13|8|oravit itaque Manue Deum et ait obsecro Domine ut vir Dei quem misisti veniat iterum et doceat nos quid debeamus facere de puero qui nasciturus est
JUDG|13|9|exaudivitque Dominus precantem Manue et apparuit rursum angelus Domini uxori eius sedenti in agro Manue autem maritus eius non erat cum ea quae cum vidisset angelum
JUDG|13|10|festinavit et cucurrit ad virum suum nuntiavitque ei dicens ecce apparuit mihi vir quem ante videram
JUDG|13|11|qui surrexit et secutus est uxorem suam veniensque ad virum dixit ei tu es qui locutus es mulieri et ille respondit ego sum
JUDG|13|12|cui Manue quando inquit sermo tuus fuerit expletus quid vis ut faciat puer aut a quo se observare debebit
JUDG|13|13|dixitque angelus Domini ad Manue ab omnibus quae locutus sum uxori tuae abstineat se
JUDG|13|14|et quicquid ex vinea nascitur non comedat vinum et siceram non bibat nullo vescatur inmundo et quod ei praecepi impleat atque custodiat
JUDG|13|15|dixitque Manue ad angelum Domini obsecro te ut adquiescas precibus meis et faciamus tibi hedum de capris
JUDG|13|16|cui respondit angelus si me cogis non comedam panes tuos sin autem vis holocaustum facere offer illud Domino et nesciebat Manue quod angelus Dei esset
JUDG|13|17|dixitque ad eum quod est tibi nomen ut si sermo tuus fuerit expletus honoremus te
JUDG|13|18|cui ille respondit cur quaeris nomen meum quod est mirabile
JUDG|13|19|tulit itaque Manue hedum de capris et libamenta et posuit super petram offerens Domino qui facit mirabilia ipse autem et uxor eius intuebantur
JUDG|13|20|cumque ascenderet flamma altaris in caelum angelus Domini in flamma pariter ascendit quod cum vidisset Manue et uxor eius proni ceciderunt in terram
JUDG|13|21|et ultra non eis apparuit angelus Domini statimque intellexit Manue angelum esse Domini
JUDG|13|22|et dixit ad uxorem suam morte moriemur quia vidimus Deum
JUDG|13|23|cui respondit mulier si Dominus nos vellet occidere de manibus nostris holocaustum et libamenta non suscepisset nec ostendisset nobis haec omnia neque ea quae sunt ventura dixisset
JUDG|13|24|peperit itaque filium et vocavit nomen eius Samson crevitque puer et benedixit ei Dominus
JUDG|13|25|coepitque spiritus Domini esse cum eo in castris Dan inter Saraa et Esthaol
JUDG|14|1|descendit igitur Samson in Thamnatha vidensque ibi mulierem de filiabus Philisthim
JUDG|14|2|ascendit et nuntiavit patri suo et matri dicens vidi mulierem in Thamnatha de filiabus Philisthinorum quam quaeso ut mihi accipiatis uxorem
JUDG|14|3|cui dixerunt pater et mater sua numquid non est mulier in filiabus fratrum tuorum et in omni populo meo quia vis accipere uxorem de Philisthim qui incircumcisi sunt dixitque Samson ad patrem suum hanc mihi accipe quia placuit oculis meis
JUDG|14|4|parentes autem eius nesciebant quod res a Domino fieret et quaereret occasionem contra Philisthim eo enim tempore Philisthim dominabantur Israheli
JUDG|14|5|descendit itaque Samson cum patre suo et matre in Thamnatha cumque venissent ad vineas oppidi apparuit catulus leonis saevus rugiens et occurrit ei
JUDG|14|6|inruit autem spiritus Domini in Samson et dilaceravit leonem quasi hedum in frusta concerperet nihil omnino habens in manu et hoc patri et matri noluit indicare
JUDG|14|7|descenditque et locutus est mulieri quae placuerat oculis eius
JUDG|14|8|et post aliquot dies revertens ut acciperet eam declinavit ut videret cadaver leonis et ecce examen apium in ore leonis erat ac favus mellis
JUDG|14|9|quem cum sumpsisset in manibus comedebat in via veniensque ad patrem suum et matrem dedit eis partem qui et ipsi comederunt nec tamen eis voluit indicare quod mel de corpore leonis adsumpserat
JUDG|14|10|descendit itaque pater eius ad mulierem et fecit filio suo Samson convivium sic enim iuvenes facere consuerant
JUDG|14|11|cum igitur cives loci vidissent eum dederunt ei sodales triginta qui essent cum eo
JUDG|14|12|quibus locutus est Samson proponam vobis problema quod si solveritis mihi intra septem dies convivii dabo vobis triginta sindones et totidem tunicas
JUDG|14|13|sin autem non potueritis solvere vos dabitis mihi triginta sindones et eiusdem numeri tunicas qui responderunt ei propone problema ut audiamus
JUDG|14|14|dixitque eis de comedente exivit cibus et de forte est egressa dulcedo nec potuerunt per tres dies propositionem solvere
JUDG|14|15|cumque adesset dies septimus dixerunt ad uxorem Samson blandire viro tuo et suade ei ut indicet tibi quid significet problema quod si facere nolueris incendimus et te et domum patris tui an idcirco nos vocastis ad nuptias ut spoliaretis
JUDG|14|16|quae fundebat apud Samson lacrimas et querebatur dicens odisti me et non diligis idcirco problema quod proposuisti filiis populi mei non vis mihi exponere at ille respondit patri meo et matri nolui dicere et tibi indicare potero
JUDG|14|17|septem igitur diebus convivii flebat apud eum tandemque die septimo cum ei molesta esset exposuit quae statim indicavit civibus suis
JUDG|14|18|et illi dixerunt ei die septimo ante solis occubitum quid dulcius melle et quid leone fortius qui ait ad eos si non arassetis in vitula mea non invenissetis propositionem meam
JUDG|14|19|inruit itaque in eo spiritus Domini descenditque Ascalonem et percussit ibi triginta viros quorum ablatas vestes dedit his qui problema solverant iratusque nimis ascendit in domum patris sui
JUDG|14|20|uxor autem eius accepit maritum unum de amicis eius et pronubis
JUDG|15|1|post aliquantum autem temporis cum dies triticeae messis instarent venit Samson invisere volens uxorem suam et adtulit ei hedum de capris cumque cubiculum eius solito vellet intrare prohibuit eum pater illius dicens
JUDG|15|2|putavi quod odisses eam et ideo tradidi illam amico tuo sed habet sororem quae iunior et pulchrior illa est sit tibi pro ea uxor
JUDG|15|3|cui respondit Samson ab hac die non erit culpa in me contra Philistheos faciam enim vobis mala
JUDG|15|4|perrexitque et cepit trecentas vulpes caudasque earum iunxit ad caudas et faces ligavit in medio
JUDG|15|5|quas igne succendens dimisit ut huc illucque discurrerent quae statim perrexerunt in segetes Philisthinorum quibus succensis et conportatae iam fruges et adhuc stantes in stipula concrematae sunt in tantum ut vineas quoque et oliveta flamma consumeret
JUDG|15|6|dixeruntque Philisthim quis fecit hanc rem quibus dictum est Samson gener Thamnathei quia tulit uxorem eius et alteri tradidit haec operatus est ascenderuntque Philisthim et conbuserunt tam mulierem quam patrem eius
JUDG|15|7|quibus ait Samson licet haec feceritis tamen adhuc ex vobis expetam ultionem et tunc quiescam
JUDG|15|8|percussitque eos ingenti plaga ita ut stupentes suram femori inponerent et descendens habitavit in spelunca petrae Aetham
JUDG|15|9|igitur ascendentes Philisthim in terra Iuda castrametati sunt et in loco qui postea vocatus est Lehi id est Maxilla eorum est fusus exercitus
JUDG|15|10|dixeruntque ad eos de tribu Iuda cur ascendistis adversum nos qui responderunt ut ligemus Samson venimus et reddamus ei quae in nos operatus est
JUDG|15|11|descenderunt ergo tria milia virorum de Iuda ad specum silicis Aetham dixeruntque ad Samson nescis quod Philisthim imperent nobis quare hoc facere voluisti quibus ille ait sicut fecerunt mihi feci eis
JUDG|15|12|ligare inquiunt te venimus et tradere in manus Philisthinorum iurate respondit mihi quod non me occidatis
JUDG|15|13|dixerunt non te occidimus sed vinctum tradimus ligaveruntque eum duobus novis funibus et tulerunt de petra Aetham
JUDG|15|14|qui cum venisset ad locum Maxillae et Philisthim vociferantes occurrissent ei inruit spiritus Domini in eum et sicut solent ad odorem ignis lina consumi ita vincula quibus ligatus erat dissipata sunt et soluta
JUDG|15|15|inventamque maxillam id est mandibulam asini quae iacebat arripiens interfecit in ea mille viros
JUDG|15|16|et ait in maxilla asini in mandibula pulli asinarum delevi eos et percussi mille viros
JUDG|15|17|cumque haec canens verba conplesset proiecit mandibulam de manu et vocavit nomen loci illius Ramathlehi quod interpretatur elevatio Maxillae
JUDG|15|18|sitiensque valde clamavit ad Dominum et ait tu dedisti in manu servi tui salutem hanc maximam atque victoriam et en siti morior incidamque in manus incircumcisorum
JUDG|15|19|aperuit itaque Dominus molarem dentem in maxilla asini et egressae sunt ex eo aquae quibus haustis refocilavit spiritum et vires recepit idcirco appellatum est nomen loci illius Fons invocantis de maxilla usque in praesentem diem
JUDG|15|20|iudicavitque Israhel in diebus Philisthim viginti annis
JUDG|16|1|abiit quoque in Gazam et vidit ibi meretricem mulierem ingressusque est ad eam
JUDG|16|2|quod cum audissent Philisthim et percrebruisset apud eos intrasse urbem Samson circumdederunt eum positis in porta civitatis custodibus et ibi tota nocte cum silentio praestolantes ut facto mane exeuntem occiderent
JUDG|16|3|dormivit autem Samson usque ad noctis medium et inde consurgens adprehendit ambas portae fores cum postibus suis et sera inpositasque umeris portavit ad verticem montis qui respicit Hebron
JUDG|16|4|post haec amavit mulierem quae habitabat in valle Sorech et vocabatur Dalila
JUDG|16|5|veneruntque ad eam principes Philisthinorum atque dixerunt decipe eum et disce ab illo in quo tantam habeat fortitudinem et quomodo eum superare valeamus et vinctum adfligere quod si feceris dabimus tibi singuli mille centum argenteos
JUDG|16|6|locuta est ergo Dalila ad Samson dic mihi obsecro in quo sit tua maxima fortitudo et quid sit quo ligatus erumpere nequeas
JUDG|16|7|cui respondit Samson si septem nervicis funibus necdum siccis et adhuc humentibus ligatus fuero infirmus ero ut ceteri homines
JUDG|16|8|adtuleruntque ad eam satrapae Philisthinorum septem funes ut dixerat quibus vinxit eum
JUDG|16|9|latentibus apud se insidiis et in cubiculo finem rei expectantibus clamavitque ad eum Philisthim super te Samson qui rupit vincula quomodo si rumpat quis filum de stuppae tortum putamine cum odorem ignis acceperit et non est cognitum in quo esset fortitudo eius
JUDG|16|10|dixitque ad eum Dalila ecce inlusisti mihi et falsum locutus es saltim nunc indica quo ligari debeas
JUDG|16|11|cui ille respondit si ligatus fuero novis funibus qui numquam fuerunt in opere infirmus ero et aliorum hominum similis
JUDG|16|12|quibus rursum Dalila vinxit eum et clamavit Philisthim super te Samson in cubiculo insidiis praeparatis qui ita rupit vincula quasi fila telarum
JUDG|16|13|dixitque Dalila rursum ad eum usquequo decipis me et falsum loqueris ostende quo vinciri debeas si inquit septem crines capitis mei cum licio plexueris et clavum his circumligatum terrae fixeris infirmus ero
JUDG|16|14|quod cum fecisset Dalila dixit ad eum Philisthim super te Samson qui consurgens de somno extraxit clavum cum crinibus et licio
JUDG|16|15|dixitque ad eum Dalila quomodo dicis quod ames me cum animus tuus non sit mecum per tres vices mentitus es mihi et noluisti dicere in quo sit tua maxima fortitudo
JUDG|16|16|cumque molesta ei esset et per multos dies iugiter adhereret spatium ad quietem non tribuens defecit anima eius et ad mortem usque lassata est
JUDG|16|17|tunc aperiens veritatem rei dixit ad eam ferrum numquam ascendit super caput meum quia nazareus id est consecratus Deo sum de utero matris meae si rasum fuerit caput meum recedet a me fortitudo mea et deficiam eroque ut ceteri homines
JUDG|16|18|videns illa quod confessus ei esset omnem animum suum misit ad principes Philisthinorum atque mandavit ascendite adhuc semel quia nunc mihi aperuit cor suum qui ascenderunt adsumpta pecunia quam promiserant
JUDG|16|19|at illa dormire eum fecit super genua sua et in sinu suo reclinare caput vocavitque tonsorem et rasit septem crines eius et coepit abicere eum et a se repellere statim enim ab eo fortitudo discessit
JUDG|16|20|dixitque Philisthim super te Samson qui de somno consurgens dixit in animo suo egrediar sicut ante feci et me excutiam nesciens quod Dominus recessisset ab eo
JUDG|16|21|quem cum adprehendissent Philisthim statim eruerunt oculos eius et duxerunt Gazam vinctum catenis et clausum in carcere molere fecerunt
JUDG|16|22|iamque capilli eius renasci coeperant
JUDG|16|23|et principes Philisthinorum convenerunt in unum ut immolarent hostias magnificas Dagon deo suo et epularentur dicentes tradidit deus noster inimicum nostrum Samson in manus nostras
JUDG|16|24|quod etiam populus videns laudabat deum suum eademque dicebat tradidit deus noster in manus nostras adversarium qui delevit terram nostram et occidit plurimos
JUDG|16|25|laetantesque per convivia sumptis iam epulis praeceperunt ut vocaretur Samson et ante eos luderet qui adductus de carcere ludebat ante eos feceruntque eum stare inter duas columnas
JUDG|16|26|qui dixit puero regenti gressus suos dimitte me ut tangam columnas quibus omnis inminet domus ut recliner super eas et paululum requiescam
JUDG|16|27|domus autem plena erat virorum ac mulierum et erant ibi omnes principes Philisthinorum ac de tecto et solario circiter tria milia utriusque sexus spectabant ludentem Samson
JUDG|16|28|at ille invocato Domino ait Domine Deus memento mei et redde nunc mihi pristinam fortitudinem Deus meus ut ulciscar me de hostibus meis et pro amissione duorum luminum unam ultionem recipiam
JUDG|16|29|et adprehendens ambas columnas quibus innitebatur domus alteramque earum dextera et alteram leva tenens
JUDG|16|30|ait moriatur anima mea cum Philisthim concussisque fortiter columnis cecidit domus super omnes principes et ceteram multitudinem quae ibi erat multoque plures interfecit moriens quam ante vivus occiderat
JUDG|16|31|descendentes autem fratres eius et universa cognatio tulerunt corpus eius et sepelierunt inter Saraa et Esthaol in sepulchro patris Manue iudicavitque Israhel viginti annis
JUDG|17|1|fuit eo tempore vir quidam de monte Ephraim nomine Michas
JUDG|17|2|qui dixit matri suae mille centum argenteos quos separaveras tibi et super quibus me audiente iuraveras ecce ego habeo et apud me sunt cui illa respondit benedictus filius meus Domino
JUDG|17|3|reddidit ergo eos matri suae quae dixerat ei consecravi et vovi argentum hoc Domino ut de manu mea suscipiat filius meus et faciat sculptile atque conflatile et nunc trado illud tibi
JUDG|17|4|reddidit igitur matri suae quae tulit ducentos argenteos et dedit eos argentario ut faceret ex eis sculptile atque conflatile quod fuit in domo Micha
JUDG|17|5|qui aediculam quoque in ea Deo separavit et fecit ephod ac therafin id est vestem sacerdotalem et idola implevitque unius filiorum suorum manum et factus est ei sacerdos
JUDG|17|6|in diebus illis non erat rex in Israhel sed unusquisque quod sibi rectum videbatur hoc faciebat
JUDG|17|7|fuit quoque alter adulescens de Bethleem Iuda et cognatione eius eratque ipse Levites et habitabat ibi
JUDG|17|8|egressusque de civitate Bethleem peregrinari voluit ubicumque sibi commodum repperisset cumque venisset in monte Ephraim iter faciens et declinasset parumper in domum Micha
JUDG|17|9|interrogatus est ab eo unde venis qui respondit Levita sum de Bethleem Iuda et vado ut habitem ubi potuero et utile mihi esse perspexero
JUDG|17|10|mane inquit apud me et esto mihi parens ac sacerdos daboque tibi per annos singulos decem argenteos ac vestem duplicem et quae ad victum necessaria sunt
JUDG|17|11|adquievit et mansit apud hominem fuitque illi quasi unus de filiis
JUDG|17|12|implevitque Micha manum eius et habuit apud se puerum sacerdotem
JUDG|17|13|nunc scio dicens quod bene mihi faciat Deus habenti levitici generis sacerdotem
JUDG|18|1|in diebus illis non erat rex in Israhel et tribus Dan quaerebat possessionem sibi ut habitaret in ea usque ad illum enim diem inter ceteras tribus sortem non acceperat
JUDG|18|2|miserunt igitur filii Dan stirpis et familiae suae quinque viros fortissimos de Saraa et Esthaol ut explorarent terram et diligenter inspicerent dixeruntque eis ite et considerate terram qui cum pergentes venissent in montem Ephraim et intrassent domum Micha requieverunt ibi
JUDG|18|3|et agnoscentes vocem adulescentis Levitae utentesque illius diversorio dixerunt ad eum quis te huc adduxit quid hic agis quam ob causam huc venire voluisti
JUDG|18|4|qui respondit eis haec et haec praestitit mihi Michas et me mercede conduxit ut sim ei sacerdos
JUDG|18|5|rogaveruntque eum ut consuleret Dominum et scire possent an prospero itinere pergerent et res haberet effectum
JUDG|18|6|qui respondit eis ite cum pace Dominus respicit viam vestram et iter quo pergitis
JUDG|18|7|euntes itaque quinque viri venerunt Lais videruntque populum habitantem in ea absque ullo timore iuxta Sidoniorum consuetudinem securum et quietum nullo eis penitus resistente magnarumque opum et procul a Sidone atque a cunctis hominibus separatum
JUDG|18|8|reversique ad fratres suos in Saraa et Esthaol et quid egissent sciscitantibus responderunt
JUDG|18|9|surgite et ascendamus ad eos vidimus enim terram valde opulentam et uberem nolite neglegere nolite cessare eamus et possideamus eam nullus erit labor
JUDG|18|10|intrabimus ad securos in regionem latissimam tradetque nobis Dominus locum in quo nullius rei est penuria eorum quae gignuntur in terra
JUDG|18|11|profecti igitur sunt de cognatione Dan id est de Saraa et Esthaol sescenti viri accincti armis bellicis
JUDG|18|12|ascendentesque manserunt in Cariathiarim Iudae qui locus ex eo tempore castrorum Dan nomen accepit et est post tergum Cariathiarim
JUDG|18|13|inde transierunt in montem Ephraim cumque venissent ad domum Micha
JUDG|18|14|dixerunt quinque viri qui prius missi fuerant ad considerandam terram Lais ceteris fratribus suis nostis quod in domibus istis sit ephod et therafin et sculptile atque conflatile videte quid vobis placeat
JUDG|18|15|et cum paululum declinassent ingressi sunt domum adulescentis Levitae qui erat in domo Micha salutaveruntque eum verbis pacificis
JUDG|18|16|sescenti autem viri ita ut erant armati stabant ante ostium
JUDG|18|17|at illi qui ingressi fuerant domum iuvenis sculptile et ephod et therafin atque conflatile tollere nitebantur et sacerdos stabat ante ostium sescentis viris fortissimis haut procul expectantibus
JUDG|18|18|tulerunt igitur qui intraverant sculptile ephod et idola atque conflatile quibus dixit sacerdos quid facitis
JUDG|18|19|cui responderunt tace et pone digitum super os tuum venique nobiscum ut habeamus te patrem et sacerdotem quid tibi melius est ut sis sacerdos in domo unius viri an in una tribu et familia in Israhel
JUDG|18|20|quod cum audisset adquievit sermonibus eorum et tulit ephod et idola ac sculptile et cum eis profectus est
JUDG|18|21|qui cum pergerent et ante se ire fecissent parvulos et iumenta et omne quod erat pretiosum
JUDG|18|22|iamque a domo Michae essent procul viri qui habitabant in aedibus Michae conclamantes secuti sunt
JUDG|18|23|et post tergum clamare coeperunt qui cum respexissent dixerunt ad Micham quid tibi vis cur clamas
JUDG|18|24|qui respondit deos meos quos mihi feci tulistis et sacerdotem et omnia quae habeo et dicitis quid tibi est
JUDG|18|25|dixeruntque ei filii Dan cave ne ultra loquaris ad nos et veniant ad te viri animo concitati et ipse cum omni domo tua pereas
JUDG|18|26|et sic coepto itinere perrexerunt videns autem Micha quod fortiores se essent reversus est in domum suam
JUDG|18|27|sescenti autem viri tulerunt sacerdotem et quae supra diximus veneruntque in Lais ad populum quiescentem atque securum et percusserunt eos in ore gladii urbemque incendio tradiderunt
JUDG|18|28|nullo penitus ferente praesidium eo quod procul habitarent a Sidone et cum nullo hominum haberent quicquam societatis ac negotii erat autem civitas sita in regione Roob quam rursum extruentes habitaverunt in ea
JUDG|18|29|vocato nomine civitatis Dan iuxta vocabulum patris sui quem genuerat Israhel quae prius Lais dicebatur
JUDG|18|30|posueruntque sibi sculptile et Ionathan filium Gersan filii Mosi ac filios eius sacerdotes in tribu Dan usque ad diem captivitatis suae
JUDG|18|31|mansitque apud eos idolum Michae omni tempore quo fuit domus Dei in Silo in diebus illis non erat rex in Israhel
JUDG|19|1|fuit quidam vir Levites habitans in latere montis Ephraim qui accepit uxorem de Bethleem Iuda
JUDG|19|2|quae reliquit eum et reversa est in domum patris sui Bethleem mansitque apud eum quattuor mensibus
JUDG|19|3|secutusque est eam vir suus volens ei reconciliari atque blandiri et secum reducere habens in comitatu puerum et duos asinos quae suscepit eum et introduxit in domum patris sui quod cum audisset socer eius eumque vidisset occurrit ei laetus
JUDG|19|4|et amplexatus est hominem mansitque gener in domo soceri tribus diebus comedens cum eo et bibens familiariter
JUDG|19|5|die autem quarto de nocte consurgens proficisci voluit quem tenuit socer et ait ad eum gusta prius pauxillum panis et conforta stomachum et sic proficisceris
JUDG|19|6|sederuntque simul et comederunt ac biberunt dixitque pater puellae ad generum suum quaeso te ut hodie hic maneas pariterque laetemur
JUDG|19|7|at ille consurgens coepit velle proficisci et nihilominus obnixe eum socer tenuit et apud se fecit manere
JUDG|19|8|mane facto parabat Levites iter cui rursum socer oro te inquit ut paululum cibi capias et adsumptis viribus donec increscat dies postea proficiscaris comederunt ergo simul
JUDG|19|9|surrexitque adulescens ut pergeret cum uxore sua et puero cui rursum locutus est socer considera quod dies ad occasum declivior sit et propinquet ad vesperum mane apud me etiam hodie et duc laetum diem et cras proficisceris ut vadas in domum tuam
JUDG|19|10|noluit gener adquiescere sermonibus eius sed statim perrexit et venit contra Iebus quae altero nomine vocabatur Hierusalem ducens secum duos asinos onustos et concubinam
JUDG|19|11|iamque aderant iuxta Iebus et dies mutabatur in noctem dixitque puer ad dominum suum veni obsecro declinemus ad urbem Iebuseorum et maneamus in ea
JUDG|19|12|cui respondit dominus non ingrediar oppidum gentis alienae quae non est de filiis Israhel sed transibo usque Gabaa
JUDG|19|13|et cum illuc pervenero manebimus in ea aut certe in urbe Rama
JUDG|19|14|transierunt igitur Iebus et coeptum carpebant iter occubuitque eis sol iuxta Gabaa quae est in tribu Beniamin
JUDG|19|15|deverteruntque ad eam ut manerent ibi quo cum intrassent sedebant in platea civitatis et nullus eos recipere volebat hospitio
JUDG|19|16|et ecce apparuit homo senex revertens de agro et de opere suo vespere qui et ipse erat de monte Ephraim et peregrinus habitabat in Gabaa homines autem regionis illius erant filii Iemini
JUDG|19|17|elevatisque oculis vidit senex sedentem hominem cum sarcinulis suis in platea civitatis et dixit ad eum unde venis et quo vadis
JUDG|19|18|qui respondit ei profecti sumus de Bethleem Iuda et pergimus ad locum nostrum qui est in latere montis Ephraim unde ieramus Bethleem et nunc vadimus ad domum Dei nullusque nos sub tectum suum vult recipere
JUDG|19|19|habentes paleas et faenum in asinorum pabulum et panem ac vinum in meos et ancillae tuae usus et pueri qui mecum est nulla re indigemus nisi hospitio
JUDG|19|20|cui respondit senex pax tecum sit ego praebebo omnia quae necessaria sunt tantum quaeso ne in platea maneas
JUDG|19|21|introduxitque eum in domum suam et pabulum asinis praebuit ac postquam laverunt pedes suos recepit eos in convivium
JUDG|19|22|illis epulantibus et post laborem itineris cibo ac potu reficientibus corpora venerunt viri civitatis illius filii Belial id est absque iugo et circumdantes domum senis fores pulsare coeperunt clamantes ad dominum domus atque dicentes educ virum qui ingressus est domum tuam ut abutamur eo
JUDG|19|23|egressusque est ad eos senex et ait nolite fratres nolite facere malum hoc quia ingressus est homo hospitium meum et cessate ab hac stultitia
JUDG|19|24|habeo filiam virginem et hic homo habet concubinam educam eas ad vos ut humilietis eas et vestram libidinem conpleatis tantum obsecro ne scelus hoc contra naturam operemini in virum
JUDG|19|25|nolebant adquiescere sermonibus eius quod cernens homo eduxit ad eos concubinam suam et eis tradidit inludendam qua cum tota nocte abusi essent dimiserunt eam mane
JUDG|19|26|at mulier recedentibus tenebris venit ad ostium domus ubi manebat dominus suus et ibi corruit
JUDG|19|27|mane facto surrexit homo et aperuit ostium ut coeptam expleret viam et ecce concubina eius iacebat ante ostium sparsis in limine manibus
JUDG|19|28|cui ille putans eam quiescere loquebatur surge ut ambulemus qua nihil respondente intellegens quod erat tulit eam et inposuit asino reversusque est in domum suam
JUDG|19|29|quam cum esset ingressus arripuit gladium et cadaver uxoris cum ossibus suis in duodecim partes ac frusta concidens misit in omnes terminos Israhel
JUDG|19|30|quod cum vidissent singuli conclamabant numquam res talis facta est in Israhel ex eo die quo ascenderunt patres nostri de Aegypto usque in praesens tempus ferte sententiam et in commune decernite quid facto opus sit
JUDG|20|1|egressi sunt itaque omnes filii Israhel et pariter congregati quasi vir unus de Dan usque Bersabee et terra Galaad ad Dominum in Maspha
JUDG|20|2|omnesque anguli populorum et cunctae tribus Israhel in ecclesiam populi Dei convenerunt quadringenta milia peditum pugnatorum
JUDG|20|3|nec latuit filios Beniamin quod ascendissent filii Israhel in Maspha interrogatusque Levita maritus mulieris interfectae quomodo tantum scelus perpetratum esset
JUDG|20|4|respondit veni in Gabaa Beniamin cum uxore mea illucque deverti
JUDG|20|5|et ecce homines civitatis illius circumdederunt nocte domum in qua manebam volentes me occidere et uxorem meam incredibili libidinis furore vexantes denique mortua est
JUDG|20|6|quam arreptam in frusta concidi misique partes in omnes terminos possessionis vestrae quia numquam tantum nefas et tam grande piaculum factum est in Israhel
JUDG|20|7|adestis omnes filii Israhel decernite quid facere debeatis
JUDG|20|8|stansque omnis populus quasi unius hominis sermone respondit non recedemus in tabernacula nostra nec suam quisquam intrabit domum
JUDG|20|9|sed hoc contra Gabaa in commune faciemus
JUDG|20|10|decem viri eligantur e centum ex omnibus tribubus Israhel et centum de mille et mille de decem milibus ut conportent exercitui cibaria et possimus pugnantes contra Gabaa Beniamin reddere ei pro scelere quod meretur
JUDG|20|11|convenitque universus Israhel ad civitatem quasi unus homo eadem mente unoque consilio
JUDG|20|12|et miserunt nuntios ad omnem tribum Beniamin qui dicerent cur tantum nefas in vobis reppertum est
JUDG|20|13|tradite homines de Gabaa qui hoc flagitium perpetrarunt ut moriantur et auferatur malum de Israhel qui noluerunt fratrum suorum filiorum Israhel audire mandatum
JUDG|20|14|sed ex cunctis urbibus quae suae sortis erant convenerunt in Gabaa ut illis ferrent auxilium et contra universum Israhel populum dimicarent
JUDG|20|15|inventique sunt viginti quinque milia de Beniamin educentium gladium praeter habitatores Gabaa
JUDG|20|16|qui septingenti erant viri fortissimi ita sinistra ut dextra proeliantes et sic fundis ad certum iacientes lapides ut capillum quoque possent percutere et nequaquam in alteram partem ictus lapidis deferretur
JUDG|20|17|virorum quoque Israhel absque filiis Beniamin inventa sunt quadringenta milia educentium gladios et paratorum ad pugnam
JUDG|20|18|qui surgentes venerunt in domum Dei hoc est in Silo consulueruntque eum atque dixerunt quis erit in exercitu nostro princeps certaminis contra filios Beniamin quibus respondit Dominus Iudas sit dux vester
JUDG|20|19|statimque filii Israhel surgentes mane castrametati sunt iuxta Gabaa
JUDG|20|20|et inde procedentes ad pugnam contra Beniamin urbem obpugnare coeperunt
JUDG|20|21|egressique filii Beniamin de Gabaa occiderunt de filiis Israhel die illo viginti duo milia viros
JUDG|20|22|rursum filii Israhel et fortitudine et numero confidentes in eodem loco in quo prius certaverant aciem direxerunt
JUDG|20|23|ita tamen ut prius ascenderent et flerent coram Domino usque ad noctem consulerentque eum et dicerent debeo ultra procedere ad dimicandum contra filios Beniamin fratres meos an non quibus ille respondit ascendite ad eum et inite certamen
JUDG|20|24|cumque filii Israhel altero die contra Beniamin ad proelium processissent
JUDG|20|25|eruperunt filii Beniamin de portis Gabaa et occurrentes eis tanta in illos caede baccati sunt ut decem et octo milia virorum educentium gladium prosternerent
JUDG|20|26|quam ob rem omnes filii Israhel venerunt in domum Dei et sedentes flebant coram Domino ieiunaveruntque illo die usque ad vesperam et obtulerunt ei holocausta et pacificas victimas
JUDG|20|27|et super statu suo interrogaverunt eo tempore ibi erat arca foederis Dei
JUDG|20|28|et Finees filius Eleazari filii Aaron praepositus domus consuluerunt igitur Dominum atque dixerunt exire ultra debemus ad pugnam contra filios Beniamin fratres nostros an quiescere quibus ait Dominus ascendite cras enim tradam eos in manus vestras
JUDG|20|29|posueruntque filii Israhel insidias per circuitum urbis Gabaa
JUDG|20|30|et tertia vice sicut semel et bis contra Beniamin exercitum produxerunt
JUDG|20|31|sed et filii Beniamin audacter eruperunt de civitate et fugientes adversarios longius persecuti sunt ita ut vulnerarent ex eis sicut primo et secundo die et caederent per duas semitas terga vertentes quarum una ferebat in Bethel altera in Gabaa atque prosternerent triginta circiter viros
JUDG|20|32|putaverunt enim solito eos more cedere qui fugam arte simulantes iniere consilium ut abstraherent eos de civitate et quasi fugientes ad supradictas semitas perducerent
JUDG|20|33|omnes itaque filii Israhel surgentes de sedibus suis tetenderunt aciem in loco qui vocatur Baalthamar insidiae quoque quae circa urbem erant paulatim se aperire coeperunt
JUDG|20|34|et ab occidentali urbis parte procedere sed et alia decem milia virorum de universo Israhel habitatores urbis ad certamina provocabant ingravatumque est bellum contra filios Beniamin et non intellexerunt quod ex omni parte illis instaret interitus
JUDG|20|35|percussitque eos Dominus in conspectu filiorum Israhel et interfecerunt ex eis in illo die viginti quinque milia et centum viros omnes bellatores et educentes gladium
JUDG|20|36|filii autem Beniamin cum se inferiores esse vidissent coeperunt fugere quod cernentes filii Israhel dederunt eis ad fugiendum locum ut ad praeparatas insidias devenirent quas iuxta urbem posuerant
JUDG|20|37|qui cum repente de latibulis surrexissent et Beniamin terga caedentibus daret ingressi sunt civitatem et percusserunt eam in ore gladii
JUDG|20|38|signum autem dederant filii Israhel his quos in insidiis conlocaverant ut postquam urbem cepissent ignem accenderent et ascendente in altum fumo captam urbem demonstrarent
JUDG|20|39|quod cum cernerent filii Israhel in ipso certamine positi putaverunt enim filii Beniamin eos fugere et instantius sequebantur caesis de exercitu eorum triginta viris
JUDG|20|40|et viderent quasi columnam fumi de civitate conscendere Beniamin quoque retro aspiciens captam cerneret civitatem et flammas in sublime ferri
JUDG|20|41|qui prius simulaverant fugam versa facie fortius resistebant quod cum vidissent filii Beniamin in fugam versi sunt
JUDG|20|42|et ad viam deserti ire coeperunt illuc quoque eos adversariis persequentibus sed et hii qui urbem succenderant occurrerunt eis
JUDG|20|43|atque ita factum est ut ex utraque parte ab hostibus caederentur nec erat ulla morientium requies ceciderunt atque prostrati sunt ad orientalem plagam urbis Gabaa
JUDG|20|44|fuerunt autem qui in eodem loco interfecti sunt decem et octo milia virorum omnes robustissimi pugnatores
JUDG|20|45|quod cum vidissent qui remanserant de Beniamin fugerunt in solitudinem et pergebant ad petram cuius vocabulum est Remmon in illa quoque fuga palantes et in diversa tendentes occiderunt quinque milia viros et cum ultra tenderent persecuti sunt eos et interfecerunt etiam alios duo milia
JUDG|20|46|et sic factum est ut omnes qui ceciderant de Beniamin in diversis locis essent viginti quinque milia pugnatores ad bella promptissimi
JUDG|20|47|remanserunt itaque de omni numero Beniamin qui evadere potuerant et fugere in solitudinem sescenti viri sederuntque in petra Remmon mensibus quattuor
JUDG|20|48|regressi autem filii Israhel omnes reliquias civitatis a viris usque ad iumenta gladio percusserunt cunctasque urbes et viculos Beniamin vorax flamma consumpsit
JUDG|21|1|iuraverunt quoque filii Israhel in Maspha et dixerunt nullus nostrum dabit filiis Beniamin de filiabus suis uxorem
JUDG|21|2|veneruntque omnes ad domum Dei in Silo et in conspectu eius sedentes usque ad vesperam levaverunt vocem et magno ululatu coeperunt flere dicentes
JUDG|21|3|quare Domine Deus Israhel factum est hoc malum in populo tuo ut hodie una tribus auferretur ex nobis
JUDG|21|4|altera autem die diluculo consurgentes extruxerunt altare obtuleruntque ibi holocausta et pacificas victimas et dixerunt
JUDG|21|5|quis non ascendit in exercitu Domini de universis tribubus Israhel grandi enim se iuramento constrinxerant cum essent in Maspha interfici eos qui defuissent
JUDG|21|6|ductique paenitentia filii Israhel super fratre suo Beniamin coeperunt dicere ablata est una tribus de Israhel
JUDG|21|7|unde uxores accipient omnes enim in commune iuravimus non daturos nos his filias nostras
JUDG|21|8|idcirco dixerunt quis est de universis tribubus Israhel qui non ascendit ad Dominum in Maspha et ecce inventi sunt habitatores Iabisgalaad in illo exercitu non fuisse
JUDG|21|9|eo quoque tempore cum essent in Silo nullus ex eis ibi reppertus est
JUDG|21|10|miserunt itaque decem milia viros robustissimos et praeceperunt eis ite et percutite habitatores Iabisgalaad in ore gladii tam uxores quam parvulos eorum
JUDG|21|11|et hoc erit quod observare debetis omne generis masculini et mulieres quae cognoverunt viros interficite
JUDG|21|12|inventaeque sunt de Iabisgalaad quadringentae virgines quae nescierunt viri torum et adduxerunt eas in castra in Silo in terra Chanaan
JUDG|21|13|miseruntque nuntios ad filios Beniamin qui erant in petra Remmon et praeceperunt eis ut eos in pace susciperent
JUDG|21|14|veneruntque filii Beniamin in illo tempore et datae sunt eis uxores de filiabus Iabisgalaad alias autem non reppererunt quas simili modo traderent
JUDG|21|15|universusque Israhel valde doluit et egit paenitudinem super interfectione unius tribus ex Israhel
JUDG|21|16|dixeruntque maiores natu quid faciemus reliquis qui non acceperunt uxores omnes in Beniamin feminae conciderunt
JUDG|21|17|et magna nobis cura ingentique studio providendum est ne una tribus deleatur ex Israhel
JUDG|21|18|filias nostras eis dare non possumus constricti iuramento et maledictione qua diximus maledictus qui dederit de filiabus suis uxorem Beniamin
JUDG|21|19|ceperuntque consilium atque dixerunt ecce sollemnitas Domini est in Silo anniversaria quae sita est ad septentrionem urbis Bethel et ad orientalem plagam viae quae de Bethel tendit ad Sycimam et ad meridiem oppidi Lebona
JUDG|21|20|praeceperuntque filiis Beniamin atque dixerunt ite et latete in vineis
JUDG|21|21|cumque videritis filias Silo ad ducendos choros ex more procedere exite repente de vineis et rapite eas singuli uxores singulas et pergite in terram Beniamin
JUDG|21|22|cumque venerint patres earum ac fratres et adversum vos queri coeperint atque iurgari dicemus eis miseremini eorum non enim rapuerunt eas iure bellantium atque victorum sed rogantibus ut acciperent non dedistis et a vestra parte peccatum est
JUDG|21|23|feceruntque filii Beniamin ut sibi fuerat imperatum et iuxta numerum suum rapuerunt sibi de his quae ducebant choros uxores singulas abieruntque in possessionem suam aedificantes urbes et habitantes in eis
JUDG|21|24|filii quoque Israhel reversi sunt per tribus et familias in tabernacula sua in diebus illis non erat rex in Israhel sed unusquisque quod sibi rectum videbatur hoc faciebat
