JOEL|1|1|The word of the LORD that came to Joel the son of Pethuel.
JOEL|1|2|Hear this, ye old men, and give ear, all ye inhabitants of the land. Hath this been in your days, or even in the days of your fathers?
JOEL|1|3|Tell ye your children of it, and let your children tell their children, and their children another generation.
JOEL|1|4|That which the palmerworm hath left hath the locust eaten; and that which the locust hath left hath the cankerworm eaten; and that which the cankerworm hath left hath the caterpiller eaten.
JOEL|1|5|Awake, ye drunkards, and weep; and howl, all ye drinkers of wine, because of the new wine; for it is cut off from your mouth.
JOEL|1|6|For a nation is come up upon my land, strong, and without number, whose teeth are the teeth of a lion, and he hath the cheek teeth of a great lion.
JOEL|1|7|He hath laid my vine waste, and barked my fig tree: he hath made it clean bare, and cast it away; the branches thereof are made white.
JOEL|1|8|Lament like a virgin girded with sackcloth for the husband of her youth.
JOEL|1|9|The meat offering and the drink offering is cut off from the house of the LORD; the priests, the LORD's ministers, mourn.
JOEL|1|10|The field is wasted, the land mourneth; for the corn is wasted: the new wine is dried up, the oil languisheth.
JOEL|1|11|Be ye ashamed, O ye husbandmen; howl, O ye vinedressers, for the wheat and for the barley; because the harvest of the field is perished.
JOEL|1|12|The vine is dried up, and the fig tree languisheth; the pomegranate tree, the palm tree also, and the apple tree, even all the trees of the field, are withered: because joy is withered away from the sons of men.
JOEL|1|13|Gird yourselves, and lament, ye priests: howl, ye ministers of the altar: come, lie all night in sackcloth, ye ministers of my God: for the meat offering and the drink offering is withholden from the house of your God.
JOEL|1|14|Sanctify ye a fast, call a solemn assembly, gather the elders and all the inhabitants of the land into the house of the LORD your God, and cry unto the LORD,
JOEL|1|15|Alas for the day! for the day of the LORD is at hand, and as a destruction from the Almighty shall it come.
JOEL|1|16|Is not the meat cut off before our eyes, yea, joy and gladness from the house of our God?
JOEL|1|17|The seed is rotten under their clods, the garners are laid desolate, the barns are broken down; for the corn is withered.
JOEL|1|18|How do the beasts groan! the herds of cattle are perplexed, because they have no pasture; yea, the flocks of sheep are made desolate.
JOEL|1|19|O LORD, to thee will I cry: for the fire hath devoured the pastures of the wilderness, and the flame hath burned all the trees of the field.
JOEL|1|20|The beasts of the field cry also unto thee: for the rivers of waters are dried up, and the fire hath devoured the pastures of the wilderness.
JOEL|2|1|Blow ye the trumpet in Zion, and sound an alarm in my holy mountain: let all the inhabitants of the land tremble: for the day of the LORD cometh, for it is nigh at hand;
JOEL|2|2|A day of darkness and of gloominess, a day of clouds and of thick darkness, as the morning spread upon the mountains: a great people and a strong; there hath not been ever the like, neither shall be any more after it, even to the years of many generations.
JOEL|2|3|A fire devoureth before them; and behind them a flame burneth: the land is as the garden of Eden before them, and behind them a desolate wilderness; yea, and nothing shall escape them.
JOEL|2|4|The appearance of them is as the appearance of horses; and as horsemen, so shall they run.
JOEL|2|5|Like the noise of chariots on the tops of mountains shall they leap, like the noise of a flame of fire that devoureth the stubble, as a strong people set in battle array.
JOEL|2|6|Before their face the people shall be much pained: all faces shall gather blackness.
JOEL|2|7|They shall run like mighty men; they shall climb the wall like men of war; and they shall march every one on his ways, and they shall not break their ranks:
JOEL|2|8|Neither shall one thrust another; they shall walk every one in his path: and when they fall upon the sword, they shall not be wounded.
JOEL|2|9|They shall run to and fro in the city; they shall run upon the wall, they shall climb up upon the houses; they shall enter in at the windows like a thief.
JOEL|2|10|The earth shall quake before them; the heavens shall tremble: the sun and the moon shall be dark, and the stars shall withdraw their shining:
JOEL|2|11|And the LORD shall utter his voice before his army: for his camp is very great: for he is strong that executeth his word: for the day of the LORD is great and very terrible; and who can abide it?
JOEL|2|12|Therefore also now, saith the LORD, turn ye even to me with all your heart, and with fasting, and with weeping, and with mourning:
JOEL|2|13|And rend your heart, and not your garments, and turn unto the LORD your God: for he is gracious and merciful, slow to anger, and of great kindness, and repenteth him of the evil.
JOEL|2|14|Who knoweth if he will return and repent, and leave a blessing behind him; even a meat offering and a drink offering unto the LORD your God?
JOEL|2|15|Blow the trumpet in Zion, sanctify a fast, call a solemn assembly:
JOEL|2|16|Gather the people, sanctify the congregation, assemble the elders, gather the children, and those that suck the breasts: let the bridegroom go forth of his chamber, and the bride out of her closet.
JOEL|2|17|Let the priests, the ministers of the LORD, weep between the porch and the altar, and let them say, Spare thy people, O LORD, and give not thine heritage to reproach, that the heathen should rule over them: wherefore should they say among the people, Where is their God?
JOEL|2|18|Then will the LORD be jealous for his land, and pity his people.
JOEL|2|19|Yea, the LORD will answer and say unto his people, Behold, I will send you corn, and wine, and oil, and ye shall be satisfied therewith: and I will no more make you a reproach among the heathen:
JOEL|2|20|But I will remove far off from you the northern army, and will drive him into a land barren and desolate, with his face toward the east sea, and his hinder part toward the utmost sea, and his stink shall come up, and his ill savour shall come up, because he hath done great things.
JOEL|2|21|Fear not, O land; be glad and rejoice: for the LORD will do great things.
JOEL|2|22|Be not afraid, ye beasts of the field: for the pastures of the wilderness do spring, for the tree beareth her fruit, the fig tree and the vine do yield their strength.
JOEL|2|23|Be glad then, ye children of Zion, and rejoice in the LORD your God: for he hath given you the former rain moderately, and he will cause to come down for you the rain, the former rain, and the latter rain in the first month.
JOEL|2|24|And the floors shall be full of wheat, and the vats shall overflow with wine and oil.
JOEL|2|25|And I will restore to you the years that the locust hath eaten, the cankerworm, and the caterpiller, and the palmerworm, my great army which I sent among you.
JOEL|2|26|And ye shall eat in plenty, and be satisfied, and praise the name of the LORD your God, that hath dealt wondrously with you: and my people shall never be ashamed.
JOEL|2|27|And ye shall know that I am in the midst of Israel, and that I am the LORD your God, and none else: and my people shall never be ashamed.
JOEL|2|28|And it shall come to pass afterward, that I will pour out my spirit upon all flesh; and your sons and your daughters shall prophesy, your old men shall dream dreams, your young men shall see visions:
JOEL|2|29|And also upon the servants and upon the handmaids in those days will I pour out my spirit.
JOEL|2|30|And I will shew wonders in the heavens and in the earth, blood, and fire, and pillars of smoke.
JOEL|2|31|The sun shall be turned into darkness, and the moon into blood, before the great and terrible day of the LORD come.
JOEL|2|32|And it shall come to pass, that whosoever shall call on the name of the LORD shall be delivered: for in mount Zion and in Jerusalem shall be deliverance, as the LORD hath said, and in the remnant whom the LORD shall call.
JOEL|3|1|For, behold, in those days, and in that time, when I shall bring again the captivity of Judah and Jerusalem,
JOEL|3|2|I will also gather all nations, and will bring them down into the valley of Jehoshaphat, and will plead with them there for my people and for my heritage Israel, whom they have scattered among the nations, and parted my land.
JOEL|3|3|And they have cast lots for my people; and have given a boy for an harlot, and sold a girl for wine, that they might drink.
JOEL|3|4|Yea, and what have ye to do with me, O Tyre, and Zidon, and all the coasts of Palestine? will ye render me a recompence? and if ye recompense me, swiftly and speedily will I return your recompence upon your own head;
JOEL|3|5|Because ye have taken my silver and my gold, and have carried into your temples my goodly pleasant things:
JOEL|3|6|The children also of Judah and the children of Jerusalem have ye sold unto the Grecians, that ye might remove them far from their border.
JOEL|3|7|Behold, I will raise them out of the place whither ye have sold them, and will return your recompence upon your own head:
JOEL|3|8|And I will sell your sons and your daughters into the hand of the children of Judah, and they shall sell them to the Sabeans, to a people far off: for the LORD hath spoken it.
JOEL|3|9|Proclaim ye this among the Gentiles; Prepare war, wake up the mighty men, let all the men of war draw near; let them come up:
JOEL|3|10|Beat your plowshares into swords and your pruninghooks into spears: let the weak say, I am strong.
JOEL|3|11|Assemble yourselves, and come, all ye heathen, and gather yourselves together round about: thither cause thy mighty ones to come down, O LORD.
JOEL|3|12|Let the heathen be wakened, and come up to the valley of Jehoshaphat: for there will I sit to judge all the heathen round about.
JOEL|3|13|Put ye in the sickle, for the harvest is ripe: come, get you down; for the press is full, the fats overflow; for their wickedness is great.
JOEL|3|14|Multitudes, multitudes in the valley of decision: for the day of the LORD is near in the valley of decision.
JOEL|3|15|The sun and the moon shall be darkened, and the stars shall withdraw their shining.
JOEL|3|16|The LORD also shall roar out of Zion, and utter his voice from Jerusalem; and the heavens and the earth shall shake: but the LORD will be the hope of his people, and the strength of the children of Israel.
JOEL|3|17|So shall ye know that I am the LORD your God dwelling in Zion, my holy mountain: then shall Jerusalem be holy, and there shall no strangers pass through her any more.
JOEL|3|18|And it shall come to pass in that day, that the mountains shall drop down new wine, and the hills shall flow with milk, and all the rivers of Judah shall flow with waters, and a fountain shall come forth out of the house of the LORD, and shall water the valley of Shittim.
JOEL|3|19|Egypt shall be a desolation, and Edom shall be a desolate wilderness, for the violence against the children of Judah, because they have shed innocent blood in their land.
JOEL|3|20|But Judah shall dwell for ever, and Jerusalem from generation to generation.
JOEL|3|21|For I will cleanse their blood that I have not cleansed: for the LORD dwelleth in Zion.
