NUM|1|1|以色列 人出 埃及 地后第二年二月初一，耶和华在 西奈 旷野，在会幕中吩咐 摩西 说：
NUM|1|2|“你要按宗族、父家、人名的数目计算 以色列 全会众，数点所有的男丁。
NUM|1|3|以色列 中凡二十岁以上能出去打仗的，你和 亚伦 要按照他们的队伍数点。
NUM|1|4|每支派要有一个人，就是父家的家长跟你们一起。
NUM|1|5|这是帮助你们的人的名字： 属 吕便 的， 示丢珥 的儿子 以利蓿 ；
NUM|1|6|属 西缅 的， 苏利沙代 的儿子 示路蔑 ；
NUM|1|7|属 犹大 的， 亚米拿达 的儿子 拿顺 ；
NUM|1|8|属 以萨迦 的， 苏押 的儿子 拿坦业 ；
NUM|1|9|属 西布伦 的， 希伦 的儿子 以利押 ；
NUM|1|10|约瑟 子孙、属 以法莲 的， 亚米忽 的儿子 以利沙玛 ；属 玛拿西 的， 比大蓿 的儿子 迦玛列 ；
NUM|1|11|属 便雅悯 的， 基多尼 的儿子 亚比但 ；
NUM|1|12|属 但 的， 亚米沙代 的儿子 亚希以谢 ；
NUM|1|13|属 亚设 的， 俄兰 的儿子 帕结 ；
NUM|1|14|属 迦得 的， 丢珥 的儿子 以利雅萨 ；
NUM|1|15|属 拿弗他利 的， 以南 的儿子 亚希拉 。”
NUM|1|16|这些是从会众中选出来的父系支派的领袖，是 以色列 部队的官长。
NUM|1|17|于是， 摩西 和 亚伦 带着这些按名指定的人，
NUM|1|18|在二月初一召集全会众。会众就照他们的宗族、父家、人名的数目，登记二十岁以上的人口。
NUM|1|19|耶和华怎样吩咐 摩西 ，他就照样在 西奈 的旷野数点他们。
NUM|1|20|以色列 的长子， 吕便 子孙的后代，照着宗族、父家、人名的数目，他们的人口凡二十岁以上能出去打仗的男丁，
NUM|1|21|吕便 支派被数的共有四万六千五百名。
NUM|1|22|西缅 子孙的后代，照着宗族、父家、被数 人名的数目，他们的人口凡二十岁以上能出去打仗的男丁，
NUM|1|23|西缅 支派被数的共有五万九千三百名。
NUM|1|24|迦得 子孙的后代，照着宗族、父家、人名的数目，凡二十岁以上能出去打仗的，
NUM|1|25|迦得 支派被数的共有四万五千六百五十名。
NUM|1|26|犹大 子孙的后代，照着宗族、父家、人名的数目，凡二十岁以上能出去打仗的，
NUM|1|27|犹大 支派被数的共有七万四千六百名。
NUM|1|28|以萨迦 子孙的后代，照着宗族、父家、人名的数目，凡二十岁以上能出去打仗的，
NUM|1|29|以萨迦 支派被数的共有五万四千四百名。
NUM|1|30|西布伦 子孙的后代，照着宗族、父家、人名的数目，凡二十岁以上能出去打仗的，
NUM|1|31|西布伦 支派被数的共有五万七千四百名。
NUM|1|32|约瑟 子孙属 以法莲 子孙的后代，照着宗族、父家、人名的数目，凡二十岁以上能出去打仗的，
NUM|1|33|以法莲 支派被数的共有四万零五百名。
NUM|1|34|玛拿西 子孙的后代，照着宗族、父家、人名的数目，凡二十岁以上能出去打仗的，
NUM|1|35|玛拿西 支派被数的共有三万二千二百名。
NUM|1|36|便雅悯 子孙的后代，照着宗族、父家、人名的数目，凡二十岁以上能出去打仗的，
NUM|1|37|便雅悯 支派被数的共有三万五千四百名。
NUM|1|38|但 子孙的后代，照着宗族、父家、人名的数目，凡二十岁以上能出去打仗的，
NUM|1|39|但 支派被数的共有六万二千七百名。
NUM|1|40|亚设 子孙的后代，照着宗族、父家、人名的数目，凡二十岁以上能出去打仗的，
NUM|1|41|亚设 支派被数的共有四万一千五百名。
NUM|1|42|拿弗他利 子孙的后代，照着宗族、父家、人名的数目，凡二十岁以上能出去打仗的，
NUM|1|43|拿弗他利 支派被数的共有五万三千四百名。
NUM|1|44|这些就是被数点的，是 摩西 、 亚伦 和 以色列 十二个领袖所数点的；每一个领袖代表他们的父家。
NUM|1|45|以色列 人被数点的总数， 以色列 中照着父家，凡二十岁以上能出去打仗的，
NUM|1|46|他们被数点的总数是六十万三千五百五十名。
NUM|1|47|利未 人却没有按照父系支派数在其中。
NUM|1|48|耶和华吩咐 摩西 说：
NUM|1|49|“惟独 利未 支派你不可数点，也不可在 以色列 人中计算他们的人口。
NUM|1|50|你要派 利未 人管理法柜的帐幕和其中一切的器具，以及属帐幕的一切。他们要抬帐幕和其中一切的器具，并要办理帐幕的事务，在帐幕的四围安营。
NUM|1|51|帐幕将往前行的时候， 利未 人要拆卸；将驻扎的时候， 利未 人要支搭帐幕。近前来的外人必被处死。
NUM|1|52|以色列 人要按照各自的队伍安营，各归本营，各归本旗。
NUM|1|53|但 利未 人要在法柜帐幕的四围安营，免得愤怒临到 以色列 会众； 利未 人要负责看守法柜的帐幕。”
NUM|1|54|以色列 人就这样做了。凡耶和华所吩咐 摩西 的，他们都照样做了。
NUM|2|1|耶和华吩咐 摩西 和 亚伦 说：
NUM|2|2|“ 以色列 人各人要在自己的旗帜下，按照自己父家的旗号安营，对着会幕的四围安营。
NUM|2|3|“在东边，向日出的方向， 犹大 营按照他们的队伍，在它的旗帜下安营。 犹大 人的领袖是 亚米拿达 的儿子 拿顺 ，
NUM|2|4|他的军队被数的有七万四千六百名。
NUM|2|5|在他旁边安营的是 以萨迦 支派。 以萨迦 人的领袖是 苏押 的儿子 拿坦业 ，
NUM|2|6|他的军队被数的有五万四千四百名。
NUM|2|7|还有 西布伦 支派， 西布伦 人的领袖是 希伦 的儿子 以利押 ，
NUM|2|8|他的军队被数的有五万七千四百名。
NUM|2|9|凡属 犹大 营，照他们队伍被数的共有十八万六千四百名；他们要作第一队往前行。
NUM|2|10|“在南边，按照他们的队伍是 吕便 营的旗帜。 吕便 人的领袖是 示丢珥 的儿子 以利蓿 ，
NUM|2|11|他的军队被数的有四万六千五百名。
NUM|2|12|在他旁边安营的是 西缅 支派。 西缅 人的领袖是 苏利沙代 的儿子 示路蔑 ，
NUM|2|13|他的军队被数的有五万九千三百名。
NUM|2|14|还有 迦得 支派， 迦得 人的领袖是 丢珥 的儿子 以利雅萨 ，
NUM|2|15|他的军队被数的有四万五千六百五十名。
NUM|2|16|凡属 吕便 营，照他们队伍被数的共有十五万一千四百五十名；他们要作第二队往前行。
NUM|2|17|“会幕与 利未 营在诸营中间往前行。他们怎样安营就怎样往前行，各按本位，各归本旗。
NUM|2|18|“在西边，按照他们的队伍是 以法莲 营的旗帜。 以法莲 人的领袖是 亚米忽 的儿子 以利沙玛 ，
NUM|2|19|他的军队被数的有四万零五百名。
NUM|2|20|在他旁边的是 玛拿西 支派。 玛拿西 人的领袖是 比大蓿 的儿子 迦玛列 ，
NUM|2|21|他的军队被数的有三万二千二百名。
NUM|2|22|还有 便雅悯 支派， 便雅悯 人的领袖是 基多尼 的儿子 亚比但 ，
NUM|2|23|他的军队被数的有三万五千四百名。
NUM|2|24|凡属 以法莲 营，照他们队伍被数的共有十万八千一百名；他们要作第三队往前行。
NUM|2|25|“在北边，按照他们的队伍是 但 营的旗帜。 但 人的领袖是 亚米沙代 的儿子 亚希以谢 ，
NUM|2|26|他的军队被数的有六万二千七百名。
NUM|2|27|在他旁边安营的是 亚设 支派。 亚设 人的领袖是 俄兰 的儿子 帕结 ，
NUM|2|28|他的军队被数的有四万一千五百名。
NUM|2|29|还有 拿弗他利 支派， 拿弗他利 人的领袖是 以南 的儿子 亚希拉 ，
NUM|2|30|他的军队被数的有五万三千四百名。
NUM|2|31|凡属 但 营被数的共有十五万七千六百名；他们随着自己的旗帜行在最后。”
NUM|2|32|以上是 以色列 人按照各自的父家被数的，在诸营中按照各自的队伍被数的，共有六十万三千五百五十名。
NUM|2|33|但 利未 人没有数在 以色列 人中，正如耶和华所吩咐 摩西 的。
NUM|2|34|以色列 人就照着耶和华所吩咐 摩西 的做了，在各自的旗帜下安营，随着各自的宗族、父家起行。
NUM|3|1|耶和华在 西奈山 与 摩西 说话的日子， 亚伦 和 摩西 的后代如下：
NUM|3|2|这些是 亚伦 儿子的名字，长子 拿答 ，及 亚比户 、 以利亚撒 、 以他玛 。
NUM|3|3|这些是 亚伦 儿子的名字，都是受膏的祭司，是 摩西 授圣职使他们担任祭司职分的。
NUM|3|4|拿答 、 亚比户 在 西奈 的旷野向耶和华献上凡火的时候，死在耶和华面前。他们没有儿子。 以利亚撒 和 以他玛 在他们的父亲 亚伦 面前担任祭司的职分。
NUM|3|5|耶和华吩咐 摩西 说：
NUM|3|6|“你要带 利未 支派近前来，站在 亚伦 祭司面前伺候他。
NUM|3|7|他们要替他，又替全会众，在会幕前执行任务，办理帐幕的事。
NUM|3|8|他们要看守会幕一切的器具，为 以色列 人执行任务，办理帐幕的事。
NUM|3|9|你要把 利未 人给 亚伦 和他的儿子；他们是从 以色列 人中选出来完全给他的。
NUM|3|10|你要指派 亚伦 和他的儿子谨守祭司的职分；近前来的外人必被处死。”
NUM|3|11|耶和华吩咐 摩西 说：
NUM|3|12|“看哪，我从 以色列 人中选了 利未 人，代替 以色列 人中所有头胎的长子； 利未 人要归我。
NUM|3|13|因为凡头生的是我的；我在 埃及 地击杀所有头生的那日，就把 以色列 中所有头生的，无论是人或牲畜，都分别为圣归我；他们定要属我。我是耶和华。”
NUM|3|14|耶和华在 西奈 的旷野吩咐 摩西 说：
NUM|3|15|“你要照父家、宗族计算 利未 人。凡一个月以上的男子都要数点。”
NUM|3|16|于是 摩西 遵照耶和华的吩咐，按所指示的数点他们。
NUM|3|17|利未 儿子的名字是 革顺 、 哥辖 、 米拉利 。
NUM|3|18|按照宗族， 革顺 儿子的名字是 立尼 、 示每 。
NUM|3|19|按照宗族， 哥辖 的儿子是 暗兰 、 以斯哈 、 希伯伦 、 乌薛 。
NUM|3|20|按照宗族， 米拉利 的儿子是 抹利 、 母示 。按照父家，这些都是 利未 人的宗族。
NUM|3|21|属 革顺 的有 立尼 族、 示每 族，他们是 革顺 人的宗族。
NUM|3|22|他们被数的，一个月以上所有男子的数目共有七千五百名。
NUM|3|23|这 革顺 人的宗族要在西边，在帐幕后面安营。
NUM|3|24|革顺 人父家的领袖是 拉伊勒 的儿子 以利雅萨 。
NUM|3|25|革顺 的子孙在会幕中要看守的是帐幕、罩棚、罩棚的盖、会幕的门帘、
NUM|3|26|帐幕和祭坛周围院子的帷幔和门帘，以及所有需用的绳子。
NUM|3|27|属 哥辖 的有 暗兰 族、 以斯哈 族、 希伯伦 族、 乌薛 族，他们是 哥辖 人的宗族。
NUM|3|28|一个月以上所有男子的数目共有八千六百 名；他们负责看守圣所。
NUM|3|29|哥辖 子孙的宗族要在帐幕的南边安营。
NUM|3|30|哥辖 人父家宗族的领袖是 乌薛 的儿子 以利撒反 。
NUM|3|31|他们要看守的是约柜、供桌、灯台、祭坛、香坛、祭司在圣所内用的器皿、帘子，与一切相关事奉的物件。
NUM|3|32|亚伦 祭司的儿子 以利亚撒 是 利未 人众领袖的主管，他要监督那些负责看守圣所的人。
NUM|3|33|属 米拉利 的有 抹利 族、 母示 族，他们是 米拉利 的宗族。
NUM|3|34|他们被数的，一个月以上所有男子的数目共有六千二百名。
NUM|3|35|米拉利 宗族的领袖是 亚比亥 的儿子 苏列 ，他们要在帐幕的北边安营。
NUM|3|36|米拉利 子孙的职分是看守帐幕的竖板、横木、柱子、带卯眼的座和一切的器具，就是一切相关事奉的物件，
NUM|3|37|以及院子四围的柱子、其上带卯眼的座、橛子和绳子。
NUM|3|38|在帐幕前东边，向日出的方向，安营的是 摩西 、 亚伦 和 亚伦 的儿子。他们负责看守圣所，是为 以色列 人看守的。近前来的外人必被处死。
NUM|3|39|凡被数的 利未 人，就是 摩西 、 亚伦 照耶和华所指示、按宗族所数的，一个月以上所有的男子共有二万二千名。
NUM|3|40|耶和华对 摩西 说：“你要数点 以色列 人中凡一个月以上头生的男子，登记他们的名字。
NUM|3|41|我是耶和华。你要拣选 利未 人归我，代替所有头生的 以色列 人，也取 利未 人的牲畜代替 以色列 人所有头生的牲畜。”
NUM|3|42|摩西 就遵照耶和华所吩咐的，把所有 以色列 人头生的都数点了。
NUM|3|43|按人名的数目，凡一个月以上头生的男子共有二万二千二百七十三名。
NUM|3|44|耶和华吩咐 摩西 说：
NUM|3|45|“你要拣选 利未 人代替所有头生的 以色列 人，也要取 利未 人的牲畜代替 以色列 人的牲畜。 利未 人要归我，我是耶和华。
NUM|3|46|以色列 人头生的男子比 利未 人多了二百七十三名，必须把他们赎出来；
NUM|3|47|按照人丁，照圣所的舍客勒，每人当付五舍客勒，一舍客勒是二十季拉。
NUM|3|48|你要把这些多出来的人的赎银交给 亚伦 和他的儿子。”
NUM|3|49|于是 摩西 从那被 利未 人所赎以外多出来的人取了赎银。
NUM|3|50|从头生的 以色列 人所取的银子，按照圣所的舍客勒，共计一千三百六十五舍客勒。
NUM|3|51|摩西 遵照耶和华指示的话，把赎银交给 亚伦 和他的儿子，正如耶和华所吩咐的。
NUM|4|1|耶和华吩咐 摩西 和 亚伦 说：
NUM|4|2|“你要照宗族、父家计算 利未 人中 哥辖 子孙的人口，
NUM|4|3|就是从三十岁到五十岁，凡前来任职，在会幕里事奉的人。
NUM|4|4|这是 哥辖 子孙在会幕里有关至圣之物的职责。
NUM|4|5|“拔营的时候， 亚伦 和他儿子要进去，把遮掩的幔子取下，用它来遮盖法柜，
NUM|4|6|又用精美皮料盖在上面，铺上纯蓝色的布，再把杠穿上。
NUM|4|7|他们要用蓝色的布铺在供饼的桌上，将盘、碟，以及浇酒祭的杯和壶摆在上面；经常供的饼也要留在桌上。
NUM|4|8|他们要在这些东西的上面铺上朱红色的布，把精美皮料盖在上面，再把杠穿上。
NUM|4|9|他们要用蓝色的布遮盖供职用的灯台、灯台上的灯盏、灯剪、灯盘，以及所有盛油的器皿；
NUM|4|10|又要用精美皮料把灯台和灯台的一切器具包好，放在抬架上。
NUM|4|11|他们要用蓝色的布铺在金坛上，用精美皮料盖在上面，再把杠穿上。
NUM|4|12|要用蓝色的布把圣所供职用的一切器具包好，再用精美皮料盖在上面，放在抬架上。
NUM|4|13|他们要清理祭坛上的灰，用紫色的布铺在坛上；
NUM|4|14|又要把供职用的一切器具，就是祭坛一切的器具，火盆、肉叉、铲子和盘子，都摆在坛上，铺上精美皮料，再把杠穿上。
NUM|4|15|“拔营的时候， 亚伦 和他儿子把圣所和圣所一切的器具盖好之后， 哥辖 的子孙才好来抬，免得他们摸圣物而死；这是 哥辖 子孙在会幕里所当抬的。
NUM|4|16|“祭司 亚伦 的儿子 以利亚撒 所要照管的是点灯的油和香料，以及常献的素祭和膏油。他要照管整个帐幕和其中所有的，以及圣所和圣所的器具。”
NUM|4|17|耶和华吩咐 摩西 和 亚伦 说：
NUM|4|18|“你们不可使 哥辖 人宗族的这一支从 利未 人中剪除。
NUM|4|19|他们挨近至圣之物的时候，要向他们这样做，使他们存活，不致死亡； 亚伦 和他的儿子要进去，分派各人当做的，当抬的。
NUM|4|20|但是他们不可进去观看圣所的拆卸 ，免得死亡。”
NUM|4|21|耶和华吩咐 摩西 说：
NUM|4|22|“你要照父家、宗族计算 革顺 子孙的人口；
NUM|4|23|从三十岁到五十岁，凡前来任职，在会幕里事奉的，都要数点。
NUM|4|24|这是 革顺 人宗族的职责，要做的事，要抬的东西如下：
NUM|4|25|他们要抬帐幕的幔子、会幕和会幕的盖、外层精美皮料的盖、会幕的门帘、
NUM|4|26|帐幕和祭坛周围院子的帷幔和门帘、绳子，以及所有需用的器具；一切与这些东西相关的事务，他们要尽职。
NUM|4|27|革顺 人的子孙一切的事奉，就是所当抬的，所当做的，都要遵照 亚伦 和他儿子的指示；他们所当抬的，你们要派他们负责。
NUM|4|28|这是 革顺 人子孙的宗族在会幕里的事奉；他们要在 亚伦 祭司的儿子 以他玛 的手下尽职。”
NUM|4|29|“至于 米拉利 的子孙，你要照宗族、父家数点他们；
NUM|4|30|从三十岁到五十岁，凡前来任职，在会幕里事奉的，你都要数点。
NUM|4|31|这是他们在会幕里的事奉，他们负责要抬的是帐幕的竖板、横木、柱子和带卯眼的座，
NUM|4|32|院子四围的柱子和其上带卯眼的座、橛子、绳子和一切的器具，与一切相关事奉的物件。你们要按名指定他们要抬的器具。
NUM|4|33|这是 米拉利 子孙的宗族在会幕里的事奉，都在 亚伦 祭司的儿子 以他玛 的手下。”
NUM|4|34|摩西 、 亚伦 和会众的领袖按照宗族、父家数点 哥辖 人的子孙；
NUM|4|35|从三十岁到五十岁，凡前来任职，在会幕里事奉的，
NUM|4|36|按照宗族被数的共有二千七百五十名。
NUM|4|37|这是所有在会幕里事奉的 哥辖 人宗族中被数的，是 摩西 和 亚伦 遵照耶和华藉 摩西 所指示数点的。
NUM|4|38|革顺 子孙被数的，按照宗族、父家，
NUM|4|39|从三十岁到五十岁，凡前来任职，在会幕里事奉的，
NUM|4|40|按照宗族、父家被数的共有二千六百三十名。
NUM|4|41|这是所有在会幕里事奉的 革顺 子孙宗族中被数的，是 摩西 和 亚伦 遵照耶和华的指示所数点的。
NUM|4|42|米拉利 子孙宗族被数的，按照宗族、父家，
NUM|4|43|从三十岁到五十岁，凡前来任职，在会幕里事奉的，
NUM|4|44|按照宗族被数的共有三千二百名。
NUM|4|45|这是 米拉利 子孙宗族中被数的，是 摩西 和 亚伦 遵照耶和华藉 摩西 所指示数点的。
NUM|4|46|摩西 、 亚伦 和 以色列 领袖按照宗族、父家数点 利未 人，
NUM|4|47|从三十岁到五十岁，凡前来任职，在会幕里事奉，做抬物之工的，
NUM|4|48|他们被数的共有八千五百八十名。
NUM|4|49|按照耶和华藉 摩西 所指示的来分派，各人都有自己所做的事、所抬的物；他们就这样被数点，正如耶和华所吩咐 摩西 的。
NUM|5|1|耶和华吩咐 摩西 说：
NUM|5|2|“你要吩咐 以色列 人，把一切患痲疯 的、患漏症的和因尸体而不洁净的，都送到营外去。
NUM|5|3|无论男女你都要送，把他们送到营外，免得他们玷污了他们的营，这是我住在他们中间的地方。”
NUM|5|4|以色列 人就照样做，把他们送到营外去。耶和华怎样吩咐 摩西 ， 以色列 人就照样做了。
NUM|5|5|耶和华吩咐 摩西 说：
NUM|5|6|“你要吩咐 以色列 人：无论男女，若犯了人所常犯的任何罪 ，以致干犯耶和华，那人就有了罪。
NUM|5|7|他要承认所犯的罪，将所亏负人的如数赔偿，另外再加五分之一，交给所亏负的人。
NUM|5|8|那人若没有至亲可接受所赔偿的，所赔偿的就要归耶和华，交给祭司；另外还要献一只赎罪的公羊为他赎罪。
NUM|5|9|以色列 人一切的圣物中，所奉给祭司的一切礼物都要归给祭司。
NUM|5|10|各人自己的圣物归自己，给祭司的要归给祭司。”
NUM|5|11|耶和华吩咐 摩西 说：
NUM|5|12|“你要吩咐 以色列 人，对他们说：若任何人的妻子背离妇道，对丈夫不贞，
NUM|5|13|有人与她同寝交合，这事瞒过她的丈夫，没有被发现；她玷污自己，没有证人指控她，也没有被捉住；
NUM|5|14|丈夫若生了疑忌的心，对妻子起了疑忌，认为她玷污自己；或是丈夫生了疑忌的心，对妻子起了疑忌，虽然她没有玷污自己，
NUM|5|15|这人要带妻子到祭司那里，同时为她带十分之一伊法大麦面粉作供物。不可浇上油，也不可加乳香，因为这是疑忌的素祭，是纪念的素祭，使人记得罪孽。
NUM|5|16|“祭司要使那妇人近前来，站在耶和华面前。
NUM|5|17|祭司要把圣水盛在瓦器里，从帐幕的地上取些尘土，放在水中。
NUM|5|18|祭司要带那妇人站在耶和华面前，使她蓬头散发，再把纪念的素祭，就是疑忌的素祭，放在她的手掌，祭司手里捧着致诅咒的苦水。
NUM|5|19|祭司要叫妇人起誓，对她说：‘若没有人与你同寝，若你未曾背着丈夫做污秽的事，你就能免去这致诅咒的苦水。
NUM|5|20|但你背着丈夫，玷污自己，跟丈夫以外的人同寝。’
NUM|5|21|祭司叫妇人赌咒起誓，祭司对她说：‘当耶和华使你大腿萎缩，肚腹肿胀时，愿耶和华使你在你百姓中成为诅咒和咒骂；
NUM|5|22|愿这致诅咒的水进入你体内，使你肚腹肿胀，大腿萎缩。’妇人要说：‘阿们，阿们。’
NUM|5|23|“祭司要把这诅咒写在册上，然后用苦水涂去，
NUM|5|24|又叫妇人喝这致诅咒的苦水，这诅咒的水要进入她里面，令她痛苦。
NUM|5|25|祭司要从妇人手中取那疑忌的素祭，把素祭在耶和华面前摇一摇，拿到祭坛前；
NUM|5|26|又要从素祭中取出一把，作为纪念，烧在坛上，然后叫妇人喝这水。
NUM|5|27|祭司叫她喝了以后，她若玷污自己，确实对丈夫不贞，这致诅咒的水必进入她里面，令她痛苦，她的肚腹就要肿胀起来，大腿萎缩；这妇人就在她百姓中成为诅咒。
NUM|5|28|这妇人若没有玷污自己，是贞洁的，就要免受这灾，并且能够生育。
NUM|5|29|“这是疑忌的条例。妻子背离丈夫玷污自己，
NUM|5|30|或是丈夫生了疑忌的心，对妻子起了疑忌，祭司要使那妇人站在耶和华面前，在她身上照这条例而行。
NUM|5|31|男人可免罪责；女人必须担当自己的罪孽。”
NUM|6|1|耶和华吩咐 摩西 说：
NUM|6|2|“你要吩咐 以色列 人，对他们说：无论男女，若许了特别的愿，就是拿细耳人的愿，愿意离俗归耶和华，
NUM|6|3|他就要远离清酒烈酒，也不可喝任何清酒烈酒做的醋；不可喝任何葡萄汁，也不可吃鲜葡萄和干葡萄。
NUM|6|4|在一切离俗的日子，任何葡萄树上所结的，甚至果核和果皮，都不可吃。
NUM|6|5|“在他一切许愿离俗的日子，不可用剃刀剃头。在离俗归耶和华的日子未满之前，他要成为圣，要任由头上的发绺生长。
NUM|6|6|在他一切离俗归耶和华的日子，不可挨近死尸。
NUM|6|7|即使他的父母或兄弟姊妹死了，他也不可因他们使自己不洁净，因为他头上有离俗归上帝的记号 。
NUM|6|8|在他一切离俗的日子，他是归耶和华为圣的。
NUM|6|9|“若在他旁边忽然有人死了，因而玷污了他离俗的头，他要在第七日，得洁净的日子剃头。
NUM|6|10|第八日，他要把两只斑鸠或两只雏鸽带到会幕门口，交给祭司。
NUM|6|11|祭司要献一只作赎罪祭，一只作燔祭，为他赎因尸体而有的罪，并要在当日使他的头分别为圣。
NUM|6|12|他要另选离俗归耶和华的日子，牵一只一岁的小公羊来作赎愆祭。先前的那段日子算为无效，因为他在离俗期间被玷污了。
NUM|6|13|“拿细耳人的条例是这样的：离俗的日子满了，祭司要领他到会幕门口，
NUM|6|14|他要将供物献给耶和华，就是一只没有残疾的一岁小公羊作燔祭，一只没有残疾的一岁小母羊作赎罪祭，和一只没有残疾的公绵羊作平安祭，
NUM|6|15|一篮用油调和的无酵细面饼和抹了油的无酵薄饼，以及同献的素祭和浇酒祭。
NUM|6|16|祭司要来到耶和华面前，献上那人的赎罪祭和燔祭。
NUM|6|17|祭司要把公绵羊和那篮无酵饼献给耶和华作平安祭，又要献上同献的素祭和浇酒祭。
NUM|6|18|拿细耳人要在会幕门口剃离俗的头，把离俗头上的发放在平安祭下的火上。
NUM|6|19|他剃了离俗的头以后，祭司要取那煮好的公绵羊的一条前腿，连同篮子里的一块无酵饼和一块无酵薄饼，放在他手掌上。
NUM|6|20|祭司要拿这些在耶和华面前摇一摇，作为摇祭；这和所摇的胸、所举的腿一样是圣物，是归给祭司的。然后拿细耳人才可以喝酒。
NUM|6|21|“这是拿细耳人许愿的条例，除了他手头财力所及之外，他要为离俗献供物给耶和华。他怎样许愿，就当照离俗的条例做。”
NUM|6|22|耶和华吩咐 摩西 说：
NUM|6|23|“你要吩咐 亚伦 和他儿子说：你们要这样为 以色列 人祝福，对他们说：
NUM|6|24|‘愿耶和华赐福给你，保护你。
NUM|6|25|愿耶和华使他的脸光照你，赐恩给你。
NUM|6|26|愿耶和华向你仰脸，赐你平安。’
NUM|6|27|“他们要如此奉我的名为 以色列 人祝福；我也要赐福给他们。”
NUM|7|1|摩西 竖立帐幕后，就用膏抹了帐幕，使它分别为圣，又用膏抹其中的一切器具，以及祭坛和坛上的一切器具，使它们分别为圣。
NUM|7|2|以色列 的领袖，各父家的家长，都前来奉献。他们是各支派的领袖，管理那些被数的人。
NUM|7|3|他们把自己的供物送到耶和华面前，就是六辆篷车和十二头公牛。每两个领袖奉献一辆车，每个领袖奉献一头牛。他们把这些都带到帐幕前。
NUM|7|4|耶和华对 摩西 说：
NUM|7|5|“你要从他们收下这些，作为会幕事奉的用途，照着 利未 人所事奉的交给他们各人。”
NUM|7|6|于是 摩西 收了车和牛，交给 利未 人。
NUM|7|7|他把两辆车和四头牛，照着 革顺 子孙所事奉的交给他们，
NUM|7|8|又把四辆车和八头牛，照着 米拉利 子孙所事奉的交给他们。他们都在 亚伦 祭司的儿子 以他玛 的手下。
NUM|7|9|但没有交给 哥辖 子孙任何东西，因为他们所事奉的是圣物，必须抬在肩头上。
NUM|7|10|用膏抹祭坛的那一天，众领袖前来为献坛奉献；众领袖都在祭坛前献供物。
NUM|7|11|耶和华对 摩西 说：“众领袖为献坛奉献供物，每天要有一个领袖前来奉献。”
NUM|7|12|第一天献供物的是 犹大 支派的 亚米拿达 的儿子 拿顺 。
NUM|7|13|他的供物是：一个重一百三十舍客勒的银盘，一个重七十舍客勒的银碗，都是按照圣所的舍客勒，里面盛满了调油的细面作素祭；
NUM|7|14|一个重十舍客勒的金碟子，盛满了香；
NUM|7|15|一头公牛犊、一只公绵羊、一只一岁的小公羊作燔祭；
NUM|7|16|一只公山羊作赎罪祭；
NUM|7|17|两头公牛、五只公绵羊、五只公山羊、五只一岁的小公羊作平安祭。这是 亚米拿达 的儿子 拿顺 的供物。
NUM|7|18|第二天来献的是 以萨迦 的领袖， 苏押 的儿子 拿坦业 。
NUM|7|19|他献为供物的是：一个重一百三十舍客勒的银盘，一个重七十舍客勒的银碗，都是按照圣所的舍客勒，里面盛满了调油的细面作素祭；
NUM|7|20|一个重十舍客勒的金碟子，盛满了香；
NUM|7|21|一头公牛犊、一只公绵羊、一只一岁的小公羊作燔祭；
NUM|7|22|一只公山羊作赎罪祭；
NUM|7|23|两头公牛、五只公绵羊、五只公山羊、五只一岁的小公羊作平安祭。这是 苏押 的儿子 拿坦业 的供物。
NUM|7|24|第三天是 西布伦 子孙的领袖， 希伦 的儿子 以利押 。
NUM|7|25|他的供物是：一个重一百三十舍客勒的银盘，一个重七十舍客勒的银碗，都是按照圣所的舍客勒，里面盛满了调油的细面作素祭；
NUM|7|26|一个重十舍客勒的金碟子，盛满了香；
NUM|7|27|一头公牛犊、一只公绵羊、一只一岁的小公羊作燔祭；
NUM|7|28|一只公山羊作赎罪祭；
NUM|7|29|两头公牛、五只公绵羊、五只公山羊、五只一岁的小公羊作平安祭。这是 希伦 的儿子 以利押 的供物。
NUM|7|30|第四天是 吕便 子孙的领袖， 示丢珥 的儿子 以利蓿 。
NUM|7|31|他的供物是：一个重一百三十舍客勒的银盘，一个重七十舍客勒的银碗，都是按照圣所的舍客勒，里面盛满了调油的细面作素祭；
NUM|7|32|一个重十舍客勒的金碟子，盛满了香；
NUM|7|33|一头公牛犊、一只公绵羊、一只一岁的小公羊作燔祭；
NUM|7|34|一只公山羊作赎罪祭；
NUM|7|35|两头公牛、五只公绵羊、五只公山羊、五只一岁的小公羊作平安祭。这是 示丢珥 的儿子 以利蓿 的供物。
NUM|7|36|第五天是 西缅 子孙的领袖， 苏利沙代 的儿子 示路蔑 。
NUM|7|37|他的供物是：一个重一百三十舍客勒的银盘，一个重七十舍客勒的银碗，都是按照圣所的舍客勒，里面盛满了调油的细面作素祭；
NUM|7|38|一个重十舍客勒的金碟子，盛满了香；
NUM|7|39|一头公牛犊、一只公绵羊、一只一岁的小公羊作燔祭；
NUM|7|40|一只公山羊作赎罪祭；
NUM|7|41|两头公牛、五只公绵羊、五只公山羊、五只一岁的小公羊作平安祭。这是 苏利沙代 的儿子 示路蔑 的供物。
NUM|7|42|第六天是 迦得 子孙的领袖， 丢珥 的儿子 以利雅萨 。
NUM|7|43|他的供物是：一个重一百三十舍客勒的银盘，一个重七十舍客勒的银碗，都是按照圣所的舍客勒，里面盛满了调油的细面作素祭；
NUM|7|44|一个重十舍客勒的金碟子，盛满了香；
NUM|7|45|一头公牛犊、一只公绵羊、一只一岁的小公羊作燔祭；
NUM|7|46|一只公山羊作赎罪祭；
NUM|7|47|两头公牛、五只公绵羊、五只公山羊、五只一岁的小公羊作平安祭。这是 丢珥 的儿子 以利雅萨 的供物。
NUM|7|48|第七天是 以法莲 子孙的领袖， 亚米忽 的儿子 以利沙玛 。
NUM|7|49|他的供物是：一个重一百三十舍客勒的银盘，一个重七十舍客勒的银碗，都是按照圣所的舍客勒，里面盛满了调油的细面作素祭；
NUM|7|50|一个重十舍客勒的金碟子，盛满了香；
NUM|7|51|一头公牛犊、一只公绵羊、一只一岁的小公羊作燔祭；
NUM|7|52|一只公山羊作赎罪祭；
NUM|7|53|两头公牛、五只公绵羊、五只公山羊、五只一岁的小公羊作平安祭。这是 亚米忽 的儿子 以利沙玛 的供物。
NUM|7|54|第八天是 玛拿西 子孙的领袖， 比大蓿 的儿子 迦玛列 。
NUM|7|55|他的供物是：一个重一百三十舍客勒的银盘，一个重七十舍客勒的银碗，都是按照圣所的舍客勒，里面盛满了调油的细面作素祭；
NUM|7|56|一个重十舍客勒的金碟子，盛满了香；
NUM|7|57|一头公牛犊、一只公绵羊、一只一岁的小公羊作燔祭；
NUM|7|58|一只公山羊作赎罪祭；
NUM|7|59|两头公牛、五只公绵羊、五只公山羊、五只一岁的小公羊作平安祭。这是 比大蓿 的儿子 迦玛列 的供物。
NUM|7|60|第九天是 便雅悯 子孙的领袖， 基多尼 的儿子 亚比但 。
NUM|7|61|他的供物是：一个重一百三十舍客勒的银盘，一个重七十舍客勒的银碗，都是按照圣所的舍客勒，里面盛满了调油的细面作素祭；
NUM|7|62|一个重十舍客勒的金碟子，盛满了香；
NUM|7|63|一头公牛犊、一只公绵羊、一只一岁的小公羊作燔祭；
NUM|7|64|一只公山羊作赎罪祭；
NUM|7|65|两头公牛、五只公绵羊、五只公山羊、五只一岁的小公羊作平安祭。这是 基多尼 的儿子 亚比但 的供物。
NUM|7|66|第十天是 但 子孙的领袖， 亚米沙代 的儿子 亚希以谢 。
NUM|7|67|他的供物是：一个重一百三十舍客勒的银盘，一个重七十舍客勒的银碗，都是按照圣所的舍客勒，里面盛满了调油的细面作素祭；
NUM|7|68|一个重十舍客勒的金碟子，盛满了香；
NUM|7|69|一头公牛犊、一只公绵羊、一只一岁的小公羊作燔祭；
NUM|7|70|一只公山羊作赎罪祭；
NUM|7|71|两头公牛、五只公绵羊、五只公山羊、五只一岁的小公羊作平安祭。这是 亚米沙代 的儿子 亚希以谢 的供物。
NUM|7|72|第十一天是 亚设 子孙的领袖， 俄兰 的儿子 帕结 。
NUM|7|73|他的供物是：一个重一百三十舍客勒的银盘，一个重七十舍客勒的银碗，都是按照圣所的舍客勒，里面盛满了调油的细面作素祭；
NUM|7|74|一个重十舍客勒的金碟子，盛满了香；
NUM|7|75|一头公牛犊、一只公绵羊、一只一岁的小公羊作燔祭；
NUM|7|76|一只公山羊作赎罪祭；
NUM|7|77|两头公牛、五只公绵羊、五只公山羊、五只一岁的小公羊作平安祭。这是 俄兰 的儿子 帕结 的供物。
NUM|7|78|第十二天是 拿弗他利 子孙的领袖， 以南 儿子 亚希拉 。
NUM|7|79|他的供物是：一个重一百三十舍客勒的银盘，一个重七十舍客勒的银碗，都是按照圣所的舍客勒，里面盛满了调油的细面作素祭；
NUM|7|80|一个重十舍客勒的金碟子，盛满了香；
NUM|7|81|一头公牛犊、一只公绵羊、一只一岁的小公羊作燔祭；
NUM|7|82|一只公山羊作赎罪祭；
NUM|7|83|两头公牛、五只公绵羊、五只公山羊、五只一岁的小公羊作平安祭。这是 以南 的儿子 亚希拉 的供物。
NUM|7|84|用膏抹祭坛的那一天， 以色列 的众领袖为献坛所献的是：银盘十二个、银碗十二个、金碟子十二个；
NUM|7|85|一个银盘重一百三十，一个碗七十。一切器皿的银子，按照圣所的舍客勒共二千四百舍客勒。
NUM|7|86|十二个金碟子盛满了香，按照圣所的舍客勒，一个碟子重十舍客勒，所有碟子的金子共一百二十舍客勒。
NUM|7|87|作燔祭的共有公牛十二头、公羊十二只、一岁的小公羊十二只，和同献的素祭，以及作赎罪祭的公山羊十二只；
NUM|7|88|作平安祭的共有公牛二十四头、公绵羊六十只、公山羊六十只、一岁的小公羊六十只。这就是用膏抹坛之后，为献坛的奉献。
NUM|7|89|摩西 进会幕要与耶和华说话的时候，听见法柜的柜盖以上二基路伯中间有对他说话的声音。耶和华向他说话。
NUM|8|1|耶和华吩咐 摩西 说：
NUM|8|2|“你要吩咐 亚伦 ，对他说：点灯的时候，七盏灯都要照亮灯台前面。”
NUM|8|3|亚伦 就照样做了；他点灯，照亮了灯台前面，正如耶和华所吩咐 摩西 的。
NUM|8|4|灯台是这样造的：灯台是用金子锤出来的，连座带花都是锤出来的。 摩西 照着耶和华所指示的样式造了灯台。
NUM|8|5|耶和华吩咐 摩西 说：
NUM|8|6|“你要从 以色列 人中选出 利未 人来，洁净他们。
NUM|8|7|你要这样做来洁净他们：要用洁净的水弹在他们身上，又叫他们用剃刀剃刮全身，洗净衣服，洁净自己。
NUM|8|8|然后他们要取一头公牛犊，以及同献的素祭，就是调油的细面。你要另取一头公牛犊作赎罪祭。
NUM|8|9|你要带 利未 人到会幕前，并且要召集 以色列 全会众。
NUM|8|10|你要把 利未 人带到耶和华面前， 以色列 人要为 利未 人按手。
NUM|8|11|亚伦 要从 以色列 人中将 利未 人奉献 在耶和华面前，作为摇祭，使他们事奉耶和华。
NUM|8|12|利未 人要按手在那两头牛的头上；你要将一头作赎罪祭，一头作燔祭，献给耶和华，为 利未 人赎罪。
NUM|8|13|你也要使 利未 人站在 亚伦 和他儿子面前，将他们奉献给耶和华，作为摇祭。
NUM|8|14|“你从 以色列 人中将 利未 人分别出来， 利未 人就归我了。
NUM|8|15|你洁净了 利未 人，奉献他们作为摇祭之后，他们就可以进会幕事奉。
NUM|8|16|因为他们是从 以色列 人中全然献给我的；我选他们归我，代替 以色列 人中所有头胎的长子。
NUM|8|17|因为 以色列 人中凡头生的，无论是人或牲畜，都是我的。我在 埃及 地击杀所有头生的那日，已将他们分别为圣归我。
NUM|8|18|我选 利未 人代替 以色列 人中所有头生的。
NUM|8|19|我从 以色列 人中将 利未 人给 亚伦 和他的儿子作为赏赐，在会幕中为 以色列 人事奉，又为 以色列 人赎罪，免得 以色列 人因挨近圣所而遭受灾祸。”
NUM|8|20|摩西 、 亚伦 和 以色列 全会众就向 利未 人这样做。关于 利未 人，凡耶和华怎样吩咐 摩西 ， 以色列 人就向他们照样做了。
NUM|8|21|于是 利未 人从罪中洁净自己，洗净衣服。 亚伦 将他们奉献在耶和华面前，作为摇祭，又为他们赎罪，洁净他们。
NUM|8|22|然后 利未 人进去，在 亚伦 和他儿子面前，在会幕中事奉。关于 利未 人，耶和华怎样吩咐 摩西 ，他们就向 利未 人照样做了。
NUM|8|23|耶和华吩咐 摩西 说：
NUM|8|24|“这是有关 利未 人的：二十五岁以上的人都要前来任职，在会幕里事奉。
NUM|8|25|到了五十岁，他们就要从事奉的工作中退休，不再事奉，
NUM|8|26|只可在会幕里辅助他们的弟兄尽责，他们自己不再事奉了。关于 利未 人的职责，你要向他们这样做。”
NUM|9|1|以色列 人出 埃及 地以后，第二年正月，耶和华在 西奈 的旷野吩咐 摩西 说：
NUM|9|2|“ 以色列 人应当在所定的日期守逾越节。
NUM|9|3|你们要在本月十四日黄昏的时候 ，在所定的日期守这节，按照一切的律例典章守节。”
NUM|9|4|于是 摩西 吩咐 以色列 人守逾越节。
NUM|9|5|正月十四日黄昏的时候，他们就在 西奈 的旷野守逾越节。凡耶和华所吩咐 摩西 的， 以色列 人都照样做了。
NUM|9|6|有几个人因尸体成了不洁净，不能在那日守逾越节。当天他们到 摩西 、 亚伦 面前。
NUM|9|7|那些人对他说：“我们因尸体而不洁净，为何禁止我们，不能和 以色列 人在所定的日期献供物给耶和华呢？”
NUM|9|8|摩西 对他们说：“你们稍等，让我去听耶和华对你们有什么吩咐。”
NUM|9|9|耶和华吩咐 摩西 说：
NUM|9|10|“你要吩咐 以色列 人说：你们和你们后代中，若有人因尸体成了不洁净，或出外远行，仍然要向耶和华守逾越节，
NUM|9|11|他们就要在二月十四日黄昏的时候守节，要吃羔羊，以及无酵饼和苦菜。
NUM|9|12|他们不可留一点食物到早晨；羔羊的骨头一根也不可折断。他们要照逾越节的一切律例守这节。
NUM|9|13|但洁净又不出外远行的人若不守逾越节，那人要从百姓中剪除，因为他没有在所定的日期献供物给耶和华，必须担当自己的罪。
NUM|9|14|若有寄居在你们那里的外人要向耶和华守逾越节，他要照逾越节的律例和典章做。无论是寄居的或是本地人，都用同样的律例。”
NUM|9|15|立起帐幕的那日，有云彩遮盖帐幕，就是法柜的帐幕；从晚上到早晨，云彩在帐幕上，形状如火。
NUM|9|16|经常都是这样：云彩遮盖帐幕，夜间云彩形状如火。
NUM|9|17|云彩几时从帐幕上升， 以色列 人就几时起行；云彩在哪里停住， 以色列 人就在哪里安营。
NUM|9|18|以色列 人遵照耶和华的指示起行，也遵照耶和华的指示安营。云彩在帐幕上停留多久，他们就留在营里多久。
NUM|9|19|云彩在帐幕上停留许多日子， 以色列 人就遵照耶和华的吩咐不起行。
NUM|9|20|有时云彩在帐幕上只停了几天，他们就遵照耶和华的指示留在营里，也遵照耶和华的指示起行。
NUM|9|21|有时云彩从晚上留到早晨；早晨云彩上升，他们就起行。无论是白天是黑夜，当云彩上升的时候，他们就要起行。
NUM|9|22|云彩停留在帐幕上，无论是两天，一个月，或更长的日子， 以色列 人就留在营里不起行；但云彩一上升，他们就起行。
NUM|9|23|他们遵照耶和华的指示安营，也遵照耶和华的指示起行。他们遵守耶和华的吩咐，是耶和华藉 摩西 所指示的话。
NUM|10|1|耶和华吩咐 摩西 说：
NUM|10|2|“你要用银子做两枝号筒，把它们锤出来，给你用来召集会众，拔营起行。
NUM|10|3|吹号的时候，全会众要到你那里，聚集在会幕的门口。
NUM|10|4|若只吹一枝，众领袖，就是 以色列 部队的官长，要到你那里聚集。
NUM|10|5|你们大声吹号的时候，东边安营的要起行。
NUM|10|6|第二次大声吹号的时候，南边安营的要起行。起行的时候，要大声吹号；
NUM|10|7|但召集会众的时候，你们要吹号，却不要吹出大声。
NUM|10|8|亚伦 子孙作祭司的要吹这号筒，作为你们世世代代永远的定例。
NUM|10|9|当你们在自己的土地上，与欺压你们的敌人打仗时，要用号筒吹出大声。你们就在耶和华－你们的上帝面前得蒙记念，也必蒙拯救脱离仇敌。
NUM|10|10|在快乐的日子，节期和初一，献燔祭与平安祭的时候，你们要吹号筒，在你们的上帝面前作为纪念。我是耶和华－你们的上帝。”
NUM|10|11|第二年二月二十日，云彩从法柜的帐幕上升。
NUM|10|12|以色列 人离开 西奈 的旷野，一段一段地往前行，云彩停在 巴兰 的旷野。
NUM|10|13|他们遵照耶和华藉 摩西 所指示的，初次往前行。
NUM|10|14|按照队伍首先起行的是 犹大 营旗帜下的人，带队的是 亚米拿达 的儿子 拿顺 。
NUM|10|15|以萨迦 支派带队的是 苏押 的儿子 拿坦业 。
NUM|10|16|西布伦 支派带队的是 希伦 的儿子 以利押 。
NUM|10|17|帐幕拆卸了， 革顺 的子孙和 米拉利 的子孙就抬着帐幕往前行。
NUM|10|18|按照队伍往前行的是 吕便 营旗帜下的人，带队的是 示丢珥 的儿子 以利蓿 。
NUM|10|19|西缅 支派带队的是 苏利沙代 的儿子 示路蔑 。
NUM|10|20|迦得 支派带队的是 丢珥 的儿子 以利雅萨 。
NUM|10|21|哥辖 人抬着圣物往前行。他们未到以前，帐幕已经立好了。
NUM|10|22|按照队伍往前行的是 以法莲 营旗帜下的人，带队的是 亚米忽 的儿子 以利沙玛 。
NUM|10|23|玛拿西 支派带队的是 比大蓿 的儿子 迦玛列 。
NUM|10|24|便雅悯 支派带队的是 基多尼 的儿子 亚比但 。
NUM|10|25|作全营后卫，按队伍往前行的是 但 营旗帜下的人，带队的是 亚米沙代 的儿子 亚希以谢 。
NUM|10|26|亚设 支派带队的是 俄兰 的儿子 帕结 。
NUM|10|27|拿弗他利 支派带队的是 以南 的儿子 亚希拉 。
NUM|10|28|以色列 人就这样按着队伍往前行。
NUM|10|29|摩西 对他岳父 ， 米甸 人 流珥 的儿子 何巴 说：“我们要往前行，到耶和华所说的地方；他曾说：‘我要将这地赐给你们。’现在请你和我们同去，我们必善待你，因为耶和华已经应许赐福气给 以色列 人。”
NUM|10|30|何巴 对他说：“我不去，我要回本地本族去。”
NUM|10|31|摩西 说：“请你不要离开我们，因为你知道我们要在旷野安营，你可以当我们的眼目。
NUM|10|32|你若和我们同去，将来耶和华以什么福气恩待我们，我们也必这样善待你。”
NUM|10|33|以色列 人离开耶和华的山，往前行了三天的路程。耶和华的约柜在前面行了三天的路程，为他们寻找安歇的地方。
NUM|10|34|他们拔营往前行，日间有耶和华的云彩在他们上面。
NUM|10|35|约柜往前行的时候， 摩西 说： “耶和华啊，求你兴起！ 愿你的仇敌溃散！ 愿恨你的人从你面前逃跑！”
NUM|10|36|约柜停住的时候，他说： “ 以色列 千万人的耶和华啊，求你回来 ！”
NUM|11|1|百姓发怨言，恶言传达到耶和华的耳中。耶和华听见了就怒气发作，耶和华的火在他们中间焚烧，烧毁营的外围。
NUM|11|2|百姓向 摩西 哀求， 摩西 祈求耶和华，火就熄了。
NUM|11|3|那地方就叫做 他备拉 ，因为耶和华的火曾在他们中间焚烧。
NUM|11|4|他们中间的闲杂人动了贪欲的心； 以色列 人又再哭着说：“谁给我们肉吃呢？
NUM|11|5|我们记得在 埃及 的时候，不花钱就可以吃鱼，还有黄瓜、西瓜、韭菜、葱、蒜。
NUM|11|6|现在我们的精力枯干了。除了这吗哪以外，在我们眼前什么都没有。”
NUM|11|7|吗哪好像芫荽子，看上去如同树脂的样子。
NUM|11|8|百姓四处走动捡取吗哪，把它用磨磨碎或用臼捣成粉，在锅中煮了做成饼，滋味好像油烤饼的滋味。
NUM|11|9|夜间露水降在营中，吗哪也随着降下。
NUM|11|10|摩西 听见百姓家家户户在帐棚门口哀哭。因此， 耶和华的怒气大大发作， 摩西 看了也不高兴。
NUM|11|11|摩西 对耶和华说：“你为何苦待仆人？我为何不在你眼前蒙恩，竟把这众百姓的担子加在我身上呢？
NUM|11|12|这众百姓岂是我怀的胎，岂是我生下来的呢？你竟对我说：‘把他们抱在怀里，如养育之父抱着吃奶的婴孩，一直抱到你起誓应许给他们祖宗的土地去。’
NUM|11|13|我从哪里拿肉给这众百姓吃呢？他们都向我哭着说：‘给我们肉吃！’
NUM|11|14|我不能独自带领这众百姓，这对我太沉重了。
NUM|11|15|如果你这样待我，倒不如立刻把我杀了吧！我若在你眼前蒙恩，求你不要让我再受这样的苦。”
NUM|11|16|耶和华对 摩西 说：“你要从 以色列 的长老中为我召集七十个人，就是你所认识，作百姓的长老和官长的，领他们到会幕，使他们和你一同站在那里。
NUM|11|17|我要在那里降临，与你说话，把降给你的灵分给他们。他们就和你分担带领百姓的担子，免得你独自承担。
NUM|11|18|你要对百姓说：‘你们要为了明天使自己分别为圣，你们将有肉吃。因你们哭着说：谁给我们肉吃呢？我们在 埃及 多么好！这声音传到了耶和华的耳中，所以他必给你们肉吃。
NUM|11|19|你们不只吃一天、两天、五天、十天、二十天，
NUM|11|20|而是整整一个月，直到肉从你们的鼻孔喷出来，使你们厌恶。因为你们厌弃那住在你们中间的耶和华，在他面前哭着说：我们为何出 埃及 呢？’”
NUM|11|21|摩西 说：“跟我在一起的百姓，步行的男人就有六十万，你还说：‘我要把肉赐给他们，使他们可以整整吃一个月。’
NUM|11|22|难道宰了羊群牛群，就够给他们吗？或者把海中所有的鱼都捕来，就够给他们吗？”
NUM|11|23|耶和华对 摩西 说：“耶和华的膀臂 岂是缩短了吗？现在你要看我的话向你应验不应验。”
NUM|11|24|摩西 出去，把耶和华的话告诉百姓，并从百姓的长老中召集七十个人来，叫他们站在会幕的四围。
NUM|11|25|耶和华在云中降临，对 摩西 说话，把降给他的灵分给那七十个长老。灵停在他们身上的时候，他们就说预言，以后却没有再说了。
NUM|11|26|但有两个人仍在营里，一个名叫 伊利达 ，一个名叫 米达 。他们本是在那些登记的人中，却没有到会幕那里去。灵停在他们身上，他们就在营里说预言。
NUM|11|27|有一个年轻人跑来告诉 摩西 说：“ 伊利达 和 米达 在营里说预言。”
NUM|11|28|嫩 的儿子 约书亚 ，年轻时就作 摩西 的助手 ，说：“请我主 摩西 禁止他们。”
NUM|11|29|摩西 对他说：“你为我的缘故嫉妒吗？惟愿耶和华的百姓都是先知，愿耶和华把他的灵降在他们身上！”
NUM|11|30|于是， 摩西 回到营里去， 以色列 的长老也回去了。
NUM|11|31|有一阵风从耶和华那里刮起，把鹌鹑从海上刮来，散落在营地和周围；一边约有一天的路程，另一边也约有一天的路程，离地面约有二肘。
NUM|11|32|百姓起来，整天整夜，甚至次日一整天，都在捕捉鹌鹑。每人至少捉到十贺梅珥，各自摆在营的四围。
NUM|11|33|但肉在他们牙间还未咀嚼时，耶和华的怒气向百姓发作，用极重的灾祸击杀百姓。
NUM|11|34|那地方就叫 基博罗．哈他瓦 ，因为他们在那里埋葬了贪欲的百姓。
NUM|11|35|百姓从 基博罗．哈他瓦 起程，到 哈洗录 ，就住在 哈洗录 。
NUM|12|1|摩西 娶了 古实 女子为妻。 米利暗 和 亚伦 因他娶了 古实 女子就批评他，
NUM|12|2|他们说：“难道耶和华只与 摩西 说话吗？他不也与我们说话吗？”耶和华听见了。
NUM|12|3|摩西 为人极其谦和，胜过地面上的任何人。
NUM|12|4|忽然，耶和华对 摩西 、 亚伦 和 米利暗 说：“你们三个人都出来，到会幕这里。”他们三个人就出来了。
NUM|12|5|耶和华在云柱中降临，停在会幕门口，叫 亚伦 和 米利暗 。二人就出来，
NUM|12|6|耶和华说：“你们要听我的话：你们中间若有先知，我－耶和华必在异象中向他显现，在梦中与他说话；
NUM|12|7|但我的仆人 摩西 不是这样，他在我全家是尽忠的。
NUM|12|8|我与他面对面说话，清清楚楚，不用谜语，他甚至看见我的形像。你们为何批评我的仆人 摩西 而不惧怕呢？”
NUM|12|9|耶和华向他们怒气发作，就离开了。
NUM|12|10|当云彩从帐幕上离开时，看哪， 米利暗 长了痲疯，像雪那么白。 亚伦 转向 米利暗 ，看哪，她长了痲疯。
NUM|12|11|亚伦 对 摩西 说：“我主啊，求你不要因我们愚昧，因我们犯罪，就将这罪加在我们身上。
NUM|12|12|求你不要使她像那一出母腹、肉已侵蚀了一半的死胎。”
NUM|12|13|于是 摩西 哀求耶和华说：“上帝啊，求你医治她！”
NUM|12|14|耶和华对 摩西 说：“她父亲若吐唾沫在她脸上，她岂不蒙羞七天吗？现在要把她隔离在营外七天，然后才领她回来。”
NUM|12|15|于是 米利暗 被隔离在营外七天；百姓没有起程，直等到 米利暗 回来。
NUM|12|16|以后百姓从 哈洗录 起行，来到 巴兰 的旷野安营。
NUM|13|1|耶和华吩咐 摩西 说：
NUM|13|2|“你要派人去窥探我所赐给 以色列 人的 迦南 地；每个父系支派要派一个人，是他们中间的族长。”
NUM|13|3|摩西 就遵照耶和华的指示，从 巴兰 旷野差派他们去；他们都是 以色列 人中的领袖。
NUM|13|4|这是他们的名字： 属 吕便 支派的， 撒刻 的儿子 沙母亚 。
NUM|13|5|属 西缅 支派的， 何利 的儿子 沙法 。
NUM|13|6|属 犹大 支派的， 耶孚尼 的儿子 迦勒 。
NUM|13|7|属 以萨迦 支派的， 约色 的儿子 以迦 。
NUM|13|8|属 以法莲 支派的， 嫩 的儿子 何西阿 。
NUM|13|9|属 便雅悯 支派的， 拉孚 的儿子 帕提 。
NUM|13|10|属 西布伦 支派的， 梭底 的儿子 迦叠 。
NUM|13|11|属 约瑟 支派，就是 玛拿西 支派的， 稣西 的儿子 迦底 。
NUM|13|12|属 但 支派的， 基玛利 的儿子 亚米利 。
NUM|13|13|属 亚设 支派的， 米迦勒 的儿子 西帖 。
NUM|13|14|属 拿弗他利 支派的， 缚西 的儿子 拿比 。
NUM|13|15|属 迦得 支派的， 玛基 的儿子 臼利 。
NUM|13|16|这些是 摩西 差派去窥探那地之人的名字。 摩西 叫 嫩 的儿子 何西阿 为 约书亚 。
NUM|13|17|摩西 差派他们去窥探 迦南 地，对他们说：“你们上到 尼革夫 那里，上到山区去，
NUM|13|18|看看那地如何：住那里的百姓是强是弱，是多是少，
NUM|13|19|他们所住的地是好是坏，所住的城镇是营地还是堡垒，
NUM|13|20|那地是肥沃还是贫瘠，当中有树木没有。你们要放胆，把那地的果子带些回来。”那时正是葡萄初熟的季节。
NUM|13|21|他们上去窥探那地，从 寻 的旷野到 利合 ，直到 哈马口 。
NUM|13|22|他们从 尼革夫 上去，到了 希伯仑 。在那里有 亚衲 族的 亚希幔 人、 示筛 人和 挞买 人。 希伯仑 的建造比 埃及 的 琐安 早七年。
NUM|13|23|他们到了 以实各谷 ，从那里砍下葡萄树枝，上面有一挂葡萄，两个人用杠抬着，又带了一些石榴和无花果。
NUM|13|24|以色列 人从那里砍下一挂葡萄，所以那地方就叫 以实各谷 。
NUM|13|25|他们窥探那地四十天之后，就回来了。
NUM|13|26|他们来到 巴兰 旷野的 加低斯 ， 摩西 、 亚伦 ，以及 以色列 全会众那里，向他们和全会众报告，又把那地的果子给他们看。
NUM|13|27|他们告诉 摩西 说：“我们到了你派我们去的那地，果然是流奶与蜜之地；这就是那地的果子。
NUM|13|28|但是住那地的百姓很强悍，城镇又大又坚固，我们也在那里看见了 亚衲 族人。
NUM|13|29|亚玛力 人住在 尼革夫 ； 赫 人、 耶布斯 人和 亚摩利 人住在山区； 迦南 人住在沿海一带和 约旦河 旁。”
NUM|13|30|迦勒 在 摩西 面前安抚百姓，说：“我们立刻上去得那地吧！我们必能征服它。”
NUM|13|31|但那些和他同去的人却说：“我们不能上去攻打那些百姓，因为他们比我们强大。”
NUM|13|32|于是探子中有人向 以色列 人散布有关所窥探之地的谣言，说：“我们所走过、所窥探之地是吞没居民之地，并且我们在那里所看见的百姓都身材高大。
NUM|13|33|我们在那里看见巨人，就是巨人中的 亚衲 族人。我们在自己眼中像蚱蜢一样，而在他们眼中，我们也确是这样。”
NUM|14|1|全会众大声喧嚷，那夜百姓哭号。
NUM|14|2|以色列 众人向 摩西 和 亚伦 发怨言，全会众对他们说：“我们宁愿死在 埃及 地，宁愿死在这旷野！
NUM|14|3|耶和华为什么要把我们领到那地，让我们倒在刀下呢？我们的妻子和孩子必成为掳物。我们回 埃及 去岂不更好吗？”
NUM|14|4|他们彼此说：“我们不如选一个领袖，回 埃及 去吧！”
NUM|14|5|摩西 和 亚伦 在 以色列 全会众面前脸伏于地。
NUM|14|6|窥探那地的人中， 嫩 的儿子 约书亚 和 耶孚尼 的儿子 迦勒 撕裂衣服，
NUM|14|7|对 以色列 全会众说：“我们所走过、所窥探之地是极美之地。
NUM|14|8|耶和华若喜爱我们，就必领我们进入那地，把这流奶与蜜之地赐给我们。
NUM|14|9|但你们不可背叛耶和华，也不要怕那地的百姓，因为他们是我们的食物。保护他们的已经离开他们，耶和华却与我们同在。不要怕他们！”
NUM|14|10|当全会众正说着要拿石头打死他们的时候，耶和华的荣光在会幕中向 以色列 众人显现。
NUM|14|11|耶和华对 摩西 说：“这百姓藐视我要到几时呢？我在他们中间行了这一切神迹，他们还不信我要到几时呢？
NUM|14|12|我要用瘟疫击杀他们，使他们不得承受那地。我要使你成为大国，比他们强大。”
NUM|14|13|摩西 对耶和华说：“ 埃及 人必听见，因你曾施展大能，领这百姓从他们中间出来。
NUM|14|14|埃及 人要告诉这地的居民，他们已经听见你─耶和华是在这百姓中间，因为你─耶和华面对面 显示自己，你的云彩停在他们以上。你日间在云柱中，夜间在火柱中，在他们的前面行。
NUM|14|15|你若把这百姓杀了，好像杀一个人那样，那听见你名声的列国必说：
NUM|14|16|‘耶和华因为不能把这百姓领进他向他们起誓应许之地，所以在旷野把他们杀了。’
NUM|14|17|现在求主显出大能，照你说过的话说：
NUM|14|18|‘耶和华不轻易发怒， 且有丰盛的慈爱。 他赦免罪孽和过犯， 万不以有罪的为无罪， 必惩罚人的罪， 从父到子，直到三、四代。’
NUM|14|19|求你照你的大慈爱赦免这百姓的罪孽，好像你从 埃及 到如今饶恕这百姓一样。”
NUM|14|20|耶和华说：“我照着你的话赦免他们。
NUM|14|21|然而，我指着我的永生与遍地充满了耶和华的荣耀起誓：
NUM|14|22|这些人虽然都看过我的荣耀和我在 埃及 与旷野所行的神迹，仍然这十次试探我，不听从我的话，
NUM|14|23|他们绝不能看见我向他们祖宗所起誓应许之地；凡藐视我的，一个也不得看见。
NUM|14|24|惟独我的仆人 迦勒 ，因他另有一个心志，专心跟从我，我要领他进入他所去过的那地；他的后裔必得那地为业。
NUM|14|25|亚玛力 人和 迦南 人住在谷中，明天你们要转回去，沿着 红海 的路往旷野去。”
NUM|14|26|耶和华对 摩西 和 亚伦 说：
NUM|14|27|“这邪恶的会众向我发怨言要到几时呢？ 以色列 人向我发的怨言，我都听见了。
NUM|14|28|你要告诉他们，耶和华说：‘我指着我的永生起誓，我必照你们在我耳中所说的待你们。
NUM|14|29|你们的尸体必倒在这旷野中。你们中间被数点，凡二十岁以上向我发怨言的，
NUM|14|30|必不得进我所起誓应许给你们居住的那地。惟有 耶孚尼 的儿子 迦勒 和 嫩 的儿子 约书亚 才能进去。
NUM|14|31|你们的孩子，就是你们说要成为掳物的，我必领他们进去，他们就得知你们所厌弃的那地。
NUM|14|32|至于你们，你们的尸体必倒在这旷野中；
NUM|14|33|你们的儿女必在旷野游牧四十年，担当你们不信的罪 ，直到你们的尸体在旷野消灭为止。
NUM|14|34|按你们窥探那地的四十日，一年抵一日，你们要担当你们的罪孽四十年，你们就知道我疏远你们了。’
NUM|14|35|我－耶和华说过，我必这样对待这一切聚集对抗我的邪恶会众。他们必在这旷野中消灭，死在这里。”
NUM|14|36|摩西 所差派去窥探那地的人回来，散布有关那地的谣言，使全会众向 摩西 发怨言，
NUM|14|37|这些散布谣言的人都遭受瘟疫，死在耶和华面前。
NUM|14|38|窥探那地的人中，惟有 嫩 的儿子 约书亚 和 耶孚尼 的儿子 迦勒 得以存活。
NUM|14|39|摩西 把这些话告诉 以色列 众人，他们都极其悲哀。
NUM|14|40|他们清晨起来，上到山顶，说：“看哪，我们要上到耶和华所说的地方；因为我们犯了罪。”
NUM|14|41|摩西 说：“你们为何要这样违背耶和华的指示呢？这事必不能顺利。
NUM|14|42|不要上去，因为耶和华不在你们中间，恐怕你们在仇敌面前被击败。
NUM|14|43|亚玛力 人和 迦南 人都在你们面前，你们必倒在刀下。因为你们背离不跟从耶和华，耶和华必不与你们同在。”
NUM|14|44|他们却擅自上到山顶。但耶和华的约柜和 摩西 都没有离开营地。
NUM|14|45|于是 亚玛力 人和住在那山区的 迦南 人下来，击败他们，追击他们直到 何珥玛 。
NUM|15|1|耶和华吩咐 摩西 说：
NUM|15|2|“你要吩咐 以色列 人，对他们说：你们到了我所赐给你们居住的地，
NUM|15|3|你们要从牛群羊群中取牲畜献给耶和华为火祭，无论是燔祭或祭物，为要还所许特别的愿或甘心祭，或节期的祭，作为献给耶和华的馨香之祭，
NUM|15|4|那献供物的要将十分之一伊法细面和四分之一欣油调和作素祭，献给耶和华。
NUM|15|5|无论是燔祭或祭物，要为每只小绵羊预备四分之一欣酒作浇酒祭。
NUM|15|6|要为每只公绵羊预备十分之二伊法细面，和三分之一欣油调和作素祭，
NUM|15|7|又用三分之一欣酒作浇酒祭，献给耶和华为馨香之祭。
NUM|15|8|你预备公牛献给耶和华作燔祭或祭物，为要还所许特别的愿，或平安祭，
NUM|15|9|就要把十分之三伊法细面和半欣油调和作素祭，和公牛一同献上，
NUM|15|10|又用半欣酒作浇酒祭，献给耶和华为馨香的火祭。
NUM|15|11|“献公牛、或公绵羊、或小绵羊、或小山羊，每只都要这样处理；
NUM|15|12|无论你们所献的数目多少，照着数目每只都要这样处理。
NUM|15|13|凡本地人将馨香的火祭献给耶和华，都要照样处理。
NUM|15|14|若有外人寄居在你们那里，或有人世世代代住在你们中间，愿意将馨香的火祭献给耶和华，你们怎样处理，他也要照样处理。
NUM|15|15|至于会众，无论是你们或寄居的外人都要遵守同一条例；这是你们世世代代永远的定例。在耶和华面前，你们怎样，寄居的也要怎样。
NUM|15|16|你们和寄居在你们那里的外人要遵守同一律法，同一典章。”
NUM|15|17|耶和华吩咐 摩西 说：
NUM|15|18|“你要吩咐 以色列 人，对他们说：你们到了我领你们进去的那地，
NUM|15|19|吃那地的粮食时，要把举祭献给耶和华。
NUM|15|20|你们要用初熟的麦子磨面，做成饼当举祭献上。你们要举上，如同举禾场的举祭。
NUM|15|21|你们世世代代要用初熟的麦子磨面，当举祭献给耶和华。
NUM|15|22|“你们若犯了错，不遵守耶和华所吩咐 摩西 的这一切命令，
NUM|15|23|就是耶和华藉 摩西 一切所命令你们的，从耶和华命令的那日直到你们的世世代代，
NUM|15|24|会众因没有察觉而犯了无心之过，全会众就要将一头公牛犊作燔祭，遵照典章把素祭和浇酒祭一同献给耶和华为馨香的祭，又要献一只公山羊作赎罪祭。
NUM|15|25|祭司要为 以色列 全会众赎罪，他们就必蒙赦免，因为这是无心之过。他们要因自己的无心之过，把供物，就是向耶和华当献的火祭和赎罪祭，带到耶和华面前。
NUM|15|26|以色列 全会众和寄居在他们中间的外人就必蒙赦免，因为这是众百姓的无心之过。
NUM|15|27|“若有一个人无意中犯了罪，他就要献一只一岁的母山羊作赎罪祭。
NUM|15|28|这误犯罪的人因无意中犯了罪，祭司要在耶和华面前为他赎罪，他就必蒙赦免。
NUM|15|29|以色列 中的本地人和寄居在他们中间的外人，若无意中犯了罪，都要遵守同一律法。
NUM|15|30|但那故意犯罪的人，无论是本地人是寄居的，亵渎了耶和华，这人必从百姓中剪除。
NUM|15|31|因为他藐视耶和华的话，违背耶和华的命令，这人一定要剪除；他的罪孽要归到自己身上。”
NUM|15|32|以色列 人还在旷野的时候，发现有一个人在安息日捡柴。
NUM|15|33|发现他捡柴的人把他带到 摩西 、 亚伦 以及全会众那里。
NUM|15|34|他们把他收押在监里，因为还不知道要怎样惩罚他。
NUM|15|35|耶和华吩咐 摩西 说：“这人应当处死；全会众要在营外用石头打死他。”
NUM|15|36|于是全会众把他带到营外，用石头打死他，是照耶和华所吩咐 摩西 的。
NUM|15|37|耶和华对 摩西 说：
NUM|15|38|“你吩咐 以色列 人，对他们说，他们世世代代要在衣服边上缝繸子，并在边上的繸子钉一条蓝色带子。
NUM|15|39|你们要佩带这繸子，好叫你们看见它就记起耶和华一切的命令，并且遵行，不随从自己内心和眼目的情欲而跟着行淫。
NUM|15|40|这样，你们就必记得并遵行我一切的命令，成为圣，归你们的上帝。
NUM|15|41|“我是耶和华－你们的上帝，曾把你们从 埃及 地领出来，要作你们的上帝。我是耶和华－你们的上帝。”
NUM|16|1|利未 的曾孙， 哥辖 的孙子， 以斯哈 的儿子 可拉 ，连同 吕便 子孙中 以利押 的儿子 大坍 和 亚比兰 ，与 比勒 的儿子 安 ，带了
NUM|16|2|以色列 人中的二百五十个领袖，就是有名望、从会众中选出来的人，在 摩西 面前一同起来，
NUM|16|3|聚集攻击 摩西 、 亚伦 ，说：“你们太过分了！全会众人人都成为圣，耶和华也在他们中间。你们为什么抬高自己，在耶和华的会众之上呢？”
NUM|16|4|摩西 听见就脸伏于地，
NUM|16|5|对 可拉 和他所有同伙的人说：“到了早晨，耶和华必指示谁是属他的，谁是成为圣的，就准许谁亲近他。他要叫自己所拣选的人亲近他。
NUM|16|6|可拉 和你所有同伙的人哪，你们要这样做：要拿着香炉，
NUM|16|7|明天在耶和华面前把火盛在炉中，把香放在上面。耶和华拣选谁，谁就成为圣。 利未 的子孙哪，你们太过分了！”
NUM|16|8|摩西 又对 可拉 说：“ 利未 的子孙，听吧！
NUM|16|9|以色列 的上帝将你们从 以色列 会众中分别出来，使你们亲近他，在耶和华的帐幕中事奉，并且站在会众面前替他们供职。这对你们岂是小事吗？
NUM|16|10|耶和华已经准许你和你所有的弟兄，就是 利未 的子孙，一同亲近他，你们还要求祭司的职分吗？
NUM|16|11|所以，你和你所有同伙的人聚集是在攻击耶和华。 亚伦 算什么，你们竟向他发怨言？”
NUM|16|12|摩西 派人去叫 以利押 的儿子 大坍 和 亚比兰 。他们却说：“我们不上去！
NUM|16|13|你把我们从流奶与蜜之地领出来，让我们死在旷野，这岂是小事？你还要自立为王管辖我们吗？
NUM|16|14|你根本没有领我们到流奶与蜜之地，也没有给我们田地和葡萄园作为产业。难道你想要挖这些人的眼睛吗？我们不上去！”
NUM|16|15|摩西 非常生气，就对耶和华说：“求你不要接受他们的供物。我并没有夺过他们一匹驴，也没有害过他们中任何一个人。”
NUM|16|16|摩西 对 可拉 说：“明天，你和你所有同伙的人，以及 亚伦 ，都要站在耶和华面前。
NUM|16|17|你们各人要拿一个香炉，把香放在上面，各人带香炉到耶和华面前，共二百五十个；你和 亚伦 也各拿自己的香炉。”
NUM|16|18|于是他们各人拿一个香炉，盛着火，加上香，和 摩西 、 亚伦 一同站在会幕的门口。
NUM|16|19|可拉 召集全会众到会幕门口攻击 摩西 和 亚伦 。这时，耶和华的荣光向全会众显现。
NUM|16|20|耶和华吩咐 摩西 和 亚伦 说：
NUM|16|21|“你们离开这会众，我好立刻把他们灭绝。”
NUM|16|22|摩西 、 亚伦 脸伏于地，说：“上帝，赐万人气息的上帝啊，一人犯罪，你就要向全会众发怒吗？”
NUM|16|23|耶和华吩咐 摩西 说：
NUM|16|24|“你吩咐会众说：‘你们远离 可拉 、 大坍 和 亚比兰 帐棚的周围。’”
NUM|16|25|摩西 起来，到 大坍 、 亚比兰 那里去； 以色列 的长老也都跟着他去。
NUM|16|26|他吩咐会众说：“你们离开这些恶人的帐棚吧！不可碰他们的任何东西，免得你们因他们一切的罪而消灭。”
NUM|16|27|于是会众远离了 可拉 、 大坍 和 亚比兰 的帐棚。 大坍 和 亚比兰 带着妻子、儿女和小孩子出来，站在自己的帐棚门口。
NUM|16|28|摩西 说：“因这件事，你们就必知道这一切事是耶和华差派我做的，并非出于我的心意。
NUM|16|29|这些人的死若和世人无异，或者他们所遭遇的和其他人相同，那么耶和华就不曾差派我了。
NUM|16|30|但是，倘若耶和华创作一件新事，使地开了裂口，把他们和一切属他们的都吞下去，叫他们活活坠落阴间，你们就知道是这些人藐视了耶和华。”
NUM|16|31|摩西 刚说完这些话，他们脚下的地就裂开，
NUM|16|32|地开了裂口，把他们和他们的家眷，以及一切属 可拉 的人和财物，都吞了下去。
NUM|16|33|他们和一切属他们的，都活活坠落阴间；地在他们上面又合拢起来，他们就从会众中灭亡了。
NUM|16|34|在他们四围的 以色列 众人听见他们的叫声，就都逃跑，说：“恐怕地也要把我们吞下去了！”
NUM|16|35|有火从耶和华那里出来，吞灭了那上香的二百五十人。
NUM|16|36|耶和华吩咐 摩西 说：
NUM|16|37|“你要对 亚伦 祭司的儿子 以利亚撒 说，把香炉从火中移开，再把炭火撒在别处，因为这些香炉是分别为圣的。
NUM|16|38|要把那些犯罪自丧己命之人的香炉锤成薄片，用以包祭坛；因为这些本是他们在耶和华面前献过，分别为圣的，可以给 以色列 人作记号。”
NUM|16|39|于是 以利亚撒 祭司把被烧死的人所献的铜香炉拿来；它们被锤出来，用以包坛，
NUM|16|40|给 以色列 人作纪念，为要叫 亚伦 子孙之外的人不得近前来，在耶和华面前烧香，免得他和 可拉 与同他一伙的人一样，正如耶和华藉 摩西 所吩咐的。
NUM|16|41|第二天， 以色列 全会众都向 摩西 、 亚伦 发怨言说：“你们杀了耶和华的百姓了。”
NUM|16|42|会众聚集攻击 摩西 、 亚伦 的时候， 摩西 和 亚伦 转向会幕，看哪，云彩遮盖会幕，耶和华的荣光显现。
NUM|16|43|摩西 、 亚伦 就来到会幕前。
NUM|16|44|耶和华吩咐 摩西 说：
NUM|16|45|“你们离开这会众，我好立刻把他们灭绝。”他们二人就脸伏于地。
NUM|16|46|摩西 对 亚伦 说：“拿你的香炉，把祭坛的火盛在里面，加上香，赶快带到会众那里，为他们赎罪。因为有愤怒从耶和华面前发出，瘟疫已经开始了。”
NUM|16|47|亚伦 照 摩西 所说的拿了香炉，跑到会众中。看哪，瘟疫已经在百姓中开始了。他就加上香，为百姓赎罪。
NUM|16|48|他站在活人和死人之间，瘟疫就止住了。
NUM|16|49|除了因 可拉 事件死的以外，遭瘟疫死的共有一万四千七百人。
NUM|16|50|亚伦 回到会幕门口 ，到 摩西 那里，瘟疫已经止住了。
NUM|17|1|耶和华吩咐 摩西 说：
NUM|17|2|“你要吩咐 以色列 人，从他们当中取杖，每父家一根；从他们所有的领袖，按着父家，共取十二根。你要把各人的名字写在他的杖上，
NUM|17|3|并要把 亚伦 的名字写在 利未 的杖上，因为各父家的家长都有一根杖。
NUM|17|4|你要把这些杖放在会幕里法柜前，我与你们 相会的地方。
NUM|17|5|我所拣选的人，他的杖必发芽。我就平息了 以色列 人向你们所发的怨言，不再达到我这里。”
NUM|17|6|于是， 摩西 吩咐 以色列 人，他们的众领袖就把杖给他，一个领袖一根杖，按照父家一个领袖一根杖，共有十二根； 亚伦 的杖也在其中。
NUM|17|7|摩西 把这些杖放在耶和华面前，在法柜的帐幕里。
NUM|17|8|第二天， 摩西 进到法柜的帐幕去，看哪， 利未 族 亚伦 的杖已经发芽，长了花苞，开了花，也结出熟的杏子！
NUM|17|9|摩西 把所有的杖从耶和华面前拿出来，给 以色列 众人看。他们都看见了，各领袖就把自己的杖拿去。
NUM|17|10|耶和华吩咐 摩西 说：“把 亚伦 的杖放回法柜前，给这些背叛之子留作记号。你就可以平息他们向我所发的怨言，他们也不会死亡。”
NUM|17|11|摩西 就照样做了；耶和华怎样吩咐他，他就照样做。
NUM|17|12|以色列 人对 摩西 说：“看哪，我们死啦！我们灭亡啦！我们全都灭亡啦！
NUM|17|13|凡挨近耶和华帐幕的，就必死亡。我们都要消灭而死吗？”
NUM|18|1|耶和华对 亚伦 说：“你和你的儿子，以及你父家的人，要一同担当干犯圣所的罪孽；你和你的儿子也要担当干犯祭司职分的罪孽。
NUM|18|2|你也要带你弟兄 利未 人，就是你父系支派的人前来，与你联合，服事你。你和你的儿子要一起在法柜的帐幕前；
NUM|18|3|他们要遵守你的吩咐，负责看守整个帐幕，只是不可挨近圣所的器具和祭坛，免得他们和你们都死亡。
NUM|18|4|他们要与你联合，负责看守会幕和帐幕一切的事；只是外人不可挨近你们。
NUM|18|5|你们要负责看守圣所和祭坛，免得愤怒再临到 以色列 人。
NUM|18|6|看哪，我已从 以色列 人中选了你们的弟兄 利未 人，交给你们为赏赐，归给耶和华，为要在会幕里事奉。
NUM|18|7|你和你的儿子要谨守祭司的职分，负责一切关于祭坛和幔子内的事。我把祭司的职分赐给你们，作为赏赐好事奉我；凡挨近的外人必被处死。”
NUM|18|8|耶和华吩咐 亚伦 说：“看哪，我已将归我的举祭，就是 以色列 人一切分别为圣之物，交给你照管；我把受膏的份赐给你和你的子孙，作为永远当得的份。
NUM|18|9|这是至圣供物中所给你的，一切献给我为至圣的素祭、赎罪祭、赎愆祭，其中所有不被火烧的供物，都要归你和你的子孙。
NUM|18|10|你要把它当作至圣之物吃 ；凡男丁都可以吃。你要以这祭物为圣。
NUM|18|11|这也是你的， 以色列 人所献的举祭和摇祭，我已赐给你和你的儿女，作为永远当得的份；你家中任何洁净的人都可以吃。
NUM|18|12|凡最好的新油、最好的新酒和五谷，就是 以色列 人献给耶和华的初熟之物，我都赐给你。
NUM|18|13|凡他们从地上所带来给耶和华的初熟之物也都要归给你。你家中任何洁净的人都可以吃。
NUM|18|14|以色列 中一切永献的都必归给你。
NUM|18|15|他们所有奉给耶和华的，无论是人是牲畜，凡头胎的，都要归给你；但是人的长子，一定要赎出来。不洁净牲畜中头生的，也要赎出来。
NUM|18|16|其中一个月以上所当赎的，要照你的估价，按圣所的舍客勒，付五舍客勒银子将他赎回，一舍客勒是二十季拉。
NUM|18|17|但是头生的牛，或头生的绵羊，或头生的山羊，却不可赎，因为它们都是圣的。要把它们的血洒在祭坛上，把它们的脂肪焚烧，当作馨香的火祭献给耶和华。
NUM|18|18|它们的肉必归你，像被摇的胸、被举的右腿归你一样。
NUM|18|19|凡 以色列 人所献给耶和华圣物中的举祭，我都赐给你和你的儿女，作为永远当得的份。这要成为你和你的后裔在耶和华面前永远的盐 约。
NUM|18|20|耶和华对 亚伦 说：“你在 以色列 人的境内不可有产业，在他们中间也不可有份。在 以色列 人中，我是你的份，你的产业。
NUM|18|21|“至于 利未 的子孙，看哪，我已赐给他们 以色列 所有出产的十分之一为业，作为他们在会幕中事奉的酬劳。
NUM|18|22|以色列 人不可再挨近会幕，免得他们担当罪而死。
NUM|18|23|惟独 利未 人要在会幕中事奉，他们要担当罪孽，作为你们世世代代永远的定例。他们在 以色列 人中不可有产业；
NUM|18|24|因为 以色列 人出产的十分之一，就是献给耶和华为举祭的，我已赐给 利未 人为业。所以我对他们说，他们不可在 以色列 人中有产业。”
NUM|18|25|耶和华吩咐 摩西 说：
NUM|18|26|“你要吩咐 利未 人，对他们说：你们从 以色列 人中所取的十分之一，就是我给你们为业的，要从这十分之一中取十分之一，作为献给耶和华的举祭。
NUM|18|27|这可算为你们的举祭，如同禾场上的谷，酒池中盛满的酒。
NUM|18|28|这样，从 以色列 人中所收取所有的十分之一，你们要从其中取举祭献给耶和华；你们要把献给耶和华的举祭归给 亚伦 祭司。
NUM|18|29|你们要将给你们一切礼物中最好的，就是分别为圣的，献给耶和华为举祭。
NUM|18|30|你要对 利未 人说：当你们把其中最好的献上为举祭之后，这剩下的就算是你们禾场上的农作物，酒池中的酒。
NUM|18|31|你们和你们的家人可以在任何地方吃；这本是你们的赏赐，是你们在会幕里事奉的酬劳。
NUM|18|32|当你们把其中最好的献上为举祭，就不致于因它担当罪。你们不可玷污 以色列 人的圣物，免得死亡。”
NUM|19|1|耶和华吩咐 摩西 和 亚伦 说：
NUM|19|2|“耶和华所吩咐的律法中，其中一条律例这样说：要吩咐 以色列 人，把一头健康、没有残疾、未曾负轭的红母牛牵到你这里来，
NUM|19|3|交给 以利亚撒 祭司。他要把牛牵到营外，人就在他面前把牛宰了。
NUM|19|4|以利亚撒 祭司要用指头蘸这牛的血，向会幕前面弹七次。
NUM|19|5|人要在他眼前焚烧这母牛，牛的皮、肉、血和粪都要焚烧。
NUM|19|6|祭司要把香柏木、牛膝草和朱红色纱都丢在焚烧牛的火中。
NUM|19|7|祭司要洗衣服，用水洗身，然后才可以进营；祭司必不洁净到晚上。
NUM|19|8|焚烧牛的人也要用水洗衣服，用水洗身，必不洁净到晚上。
NUM|19|9|一个洁净的人要收母牛的灰，存放在营外洁净的地方，为 以色列 会众留作除污秽的水之用。这是为除罪用的。
NUM|19|10|收取母牛灰的人要洗衣服，必不洁净到晚上。这要成为 以色列 人和寄居在他们中间的外人永远的定例。
NUM|19|11|“摸了任何人死尸的，必不洁净七天。
NUM|19|12|那人要在第三天和第七天洁净自己，他就洁净了。若他不在第三天和第七天洁净自己，他就不洁净了。
NUM|19|13|凡摸了死尸，就是死了的人的尸体，又不洁净自己的，就玷污了耶和华的帐幕，这人必从 以色列 中剪除；因为那除污秽的水没有洒在他身上，他就不洁净，污秽还在他身上。
NUM|19|14|“若有人死在帐棚里，条例是这样：凡进那帐棚的，和所有在帐棚里的人，都必不洁净七天。
NUM|19|15|凡敞开的，没有用绳子扎好盖子的器皿，也不洁净。
NUM|19|16|任何人在田野里摸了被刀杀的，或自然死的，或人的骨头，或坟墓，就必不洁净七天。
NUM|19|17|要为这不洁净的人拿一些烧好的除罪灰放在器皿里，倒上清水。
NUM|19|18|一个洁净的人要拿牛膝草蘸在这水中，把水弹在帐棚上，和一切器皿以及帐棚内的人身上，又要弹在那摸了骨头，或摸了被杀的或自然死的，或摸了坟墓的人身上。
NUM|19|19|那洁净的人要在第三天和第七天把水弹在不洁净的人身上，在第七天洁净那人。那人要洗衣服，用水洗澡，到晚上就洁净了。
NUM|19|20|但任何不洁净的人，他若不洁净自己，那人要从会中剪除，因为他玷污了耶和华的圣所，除污秽的水没有洒在他身上，他是不洁净的。
NUM|19|21|这要成为你们永远的定例。此外，那弹除污秽水的人也要洗衣服。凡碰除污秽水的，必不洁净到晚上。
NUM|19|22|不洁净的人所摸的任何东西都不洁净；摸了这东西的人必不洁净到晚上。”
NUM|20|1|正月间， 以色列 全会众到了 寻 的旷野；百姓住在 加低斯 。 米利暗 死在那里，也葬在那里。
NUM|20|2|会众没有水，就聚集反对 摩西 和 亚伦 。
NUM|20|3|百姓与 摩西 争闹，说：“我们恨不得与我们的弟兄一同死在耶和华面前。
NUM|20|4|你们为什么领耶和华的会众到这旷野，使我们和我们的牲畜都死在这里呢？
NUM|20|5|你们为什么领我们从 埃及 上来，把我们带到这坏的地方呢？这地方不能撒种，没有无花果树、葡萄树、石榴树，也没有水喝。”
NUM|20|6|摩西 、 亚伦 离开会众面前，到会幕的门口，脸伏于地；耶和华的荣光向他们显现。
NUM|20|7|耶和华吩咐 摩西 说：
NUM|20|8|“你拿着杖去，和你的哥哥 亚伦 召集会众，在他们眼前吩咐磐石涌出水来，水就会从磐石流出，给会众和他们的牲畜喝。”
NUM|20|9|于是 摩西 遵照耶和华所吩咐他的，从耶和华面前拿了杖去。
NUM|20|10|摩西 和 亚伦 召集会众到磐石前。 摩西 对他们说：“听着，你们这些悖逆的人！我们要叫这磐石流出水来给你们吗？”
NUM|20|11|摩西 举起手来，用杖击打磐石两下，就有许多水流出来，会众和他们的牲畜都喝了。
NUM|20|12|但是耶和华对 摩西 、 亚伦 说：“因为你们不信我，没有在 以色列 人眼前尊我为圣，所以你们必不能领这会众进入我所要赐给他们的地去。”
NUM|20|13|这就是 米利巴 水，因 以色列 人与耶和华争闹，耶和华在他们面前显为圣。
NUM|20|14|摩西 从 加低斯 差遣使者到 以东 王那里，说：“你的弟兄 以色列 这样说：‘你知道我们所遭遇的一切困难。
NUM|20|15|我们的祖先曾下到 埃及 ，我们也在 埃及 住了很多年。然而， 埃及 人却恶待我们和我们的祖先。
NUM|20|16|我们哀求耶和华，他垂听了我们的声音，差遣使者把我们从 埃及 领出来。看哪，我们到了你边界的 加低斯城 。
NUM|20|17|求你让我们穿越你的地。我们不走田间和葡萄园，也不喝井里的水。我们只走王的大路，不偏左右，直到过了你的边界。’”
NUM|20|18|但是， 以东 对他说：“你不可从我这里穿越！否则，我要带刀出去攻击你。”
NUM|20|19|以色列 人对他说：“我们只上大道。如果我和我的牲畜喝了你的水，我必付钱给你。我不求别的事，只求让我步行过去。”
NUM|20|20|以东 说：“你不可经过！”他就率领一大群军队，以强硬的手出来攻击 以色列 。
NUM|20|21|这样， 以东 不肯让 以色列 穿越他的境内， 以色列 就转去，离开他了。
NUM|20|22|以色列 全会众从 加低斯 起行，到了 何珥山 。
NUM|20|23|耶和华在 以东 地边界的 何珥山 对 摩西 、 亚伦 说：
NUM|20|24|“ 亚伦 要归到他祖先 那里。他必不得进入我所赐给 以色列 人的地，因为你们在 米利巴 水的事上违背了我的指示。
NUM|20|25|你要带 亚伦 和他的儿子 以利亚撒 上 何珥山 ，
NUM|20|26|把 亚伦 的圣衣脱下，给他的儿子 以利亚撒 穿上。 亚伦 必归去，死在那里。”
NUM|20|27|摩西 就遵照耶和华的吩咐去做，他们在全会众的眼前上了 何珥山 。
NUM|20|28|摩西 把 亚伦 的圣衣脱下，给他的儿子 以利亚撒 穿上， 亚伦 就死在山顶那里。于是， 摩西 和 以利亚撒 下了山。
NUM|20|29|全会众见 亚伦 死了， 以色列 全家就为 亚伦 举哀三十天。
NUM|21|1|住 尼革夫 的 迦南 人的 亚拉得 王，听说 以色列 从 亚他林 路来，就和 以色列 交战，掳去他们一些人。
NUM|21|2|以色列 向耶和华许愿说：“你若把这百姓真的交在我手中，我就把他们的城镇彻底毁灭。”
NUM|21|3|耶和华垂听了 以色列 的声音，把 迦南 人交出来。 以色列 就把 迦南 人和他们的城镇彻底毁灭。因此，那地方名叫 何珥玛 。
NUM|21|4|他们从 何珥山 起行，绕过 以东 地往 红海 那条路走。在路上，百姓心中烦躁。
NUM|21|5|百姓向上帝和 摩西 发怨言，说：“你们为什么把我们从 埃及 领上来 ，使我们死在旷野呢？这里没有粮食，没有水，我们厌恶这淡而无味的食物。”
NUM|21|6|耶和华派火蛇进入百姓当中去咬他们，于是 以色列 中死了许多百姓。
NUM|21|7|百姓到 摩西 那里，说：“我们有罪了，因为我们向耶和华和你发怨言。求你向耶和华祷告，叫蛇离开我们。”于是 摩西 为百姓祷告。
NUM|21|8|耶和华对 摩西 说：“你要造一条火蛇，挂在杆子上。凡被咬的，一望这蛇就必存活。”
NUM|21|9|摩西 就造了一条铜蛇，挂在杆子上。凡被蛇咬的，一望这铜蛇就活了。
NUM|21|10|以色列 人起行，安营在 阿伯 。
NUM|21|11|又从 阿伯 起行，安营在 以耶．亚巴琳 ，在 摩押 对面的旷野，向日出的方向。
NUM|21|12|又从那里起行，安营在 撒烈谷 。
NUM|21|13|从那里再起行，安营在 亚嫩河 的另一边。这 亚嫩河 在旷野，从 亚摩利 人的境内流出来； 亚嫩河 是 摩押 的边界，在 摩押 和 亚摩利 人之间。
NUM|21|14|所以《耶和华的战记》中提到： “ 苏法 的 哇哈伯 ， 亚嫩河 谷，
NUM|21|15|以及 亚珥 地区众河床的斜坡， 都靠近 摩押 的边境。”
NUM|21|16|以色列 人从那里起行，到了 比珥 。从前耶和华对 摩西 说：“召集百姓，我要给他们水”，说的就是这井。
NUM|21|17|当时， 以色列 人唱这首歌： “井啊，涌出水来！ 你们要向它歌唱！
NUM|21|18|这井是领袖用权杖所挖， 是百姓中的贵族用手杖所掘。” 以色列 人从旷野往 玛他拿 去，
NUM|21|19|从 玛他拿 到 拿哈列 ，从 拿哈列 到 巴末 ，
NUM|21|20|从 巴末 到 摩押 地的谷，又到那可以了望旷野的 毗斯迦山 顶。
NUM|21|21|以色列 差遣使者到 亚摩利 人的王 西宏 那里，说：
NUM|21|22|“求你让我们穿越你的地；我们不岔进田间和葡萄园，也不喝井里的水，只走王的大道，直到过了你的边界。”
NUM|21|23|但 西宏 不让 以色列 人穿越他的境内，就召集他的众百姓出到旷野，要攻击 以色列 ，到了 雅杂 与 以色列 交战。
NUM|21|24|以色列 人用刀杀了他，占领了他的地，从 亚嫩河 到 雅博河 ，直到 亚扪 人的边界，因为 亚扪 人的边防坚固。
NUM|21|25|以色列 人夺取这里所有的城镇，就住在 亚摩利 人的城镇中，包括 希实本 和所属的一切乡镇 。
NUM|21|26|希实本 是 亚摩利 王 西宏 的首都； 西宏 曾与先前的 摩押 王交战，从他手中夺取了他所有的地，直到 亚嫩河 。
NUM|21|27|所以那些作诗歌的说： 你们到 希实本 来吧； 愿 西宏 的城被修造建立。
NUM|21|28|因为有火从 希实本 发出， 有火焰从 西宏 的城冒出， 烧毁了 摩押 的 亚珥 ， 亚嫩河 丘坛的主 。
NUM|21|29|摩押 啊，你有祸了！ 基抹 的百姓啊，你们灭亡了！ 基抹 的男子逃亡， 女子被掳， 交给了 亚摩利 王 西宏 。
NUM|21|30|我们射了他们； 希实本 直到 底本 尽都毁灭 。 我们劫掠，直到 挪法 ； 这 挪法 直延到 米底巴 。
NUM|21|31|这样， 以色列 人就住在 亚摩利 人的地。
NUM|21|32|摩西 差派人去窥探 雅谢 ； 以色列 人占领了 雅谢 附近的乡村，赶出那里的 亚摩利 人。
NUM|21|33|后来， 以色列 人转回，往上 巴珊 的路去。 巴珊 王 噩 率领他的众百姓出来，在 以得来 与他们交战。
NUM|21|34|耶和华对 摩西 说：“不要怕他！因为我已将他和他的众百姓，以及他的地都交在你手中。你要待他如同待住在 希实本 的 亚摩利 王 西宏 一样。”
NUM|21|35|于是他们杀了 巴珊 王和他的众子，以及他的众百姓，没有留下一个幸存者，并且占领了他的地。
NUM|22|1|以色列 人起行，在 摩押 平原， 约旦河 东，对着 耶利哥 安营。
NUM|22|2|西拨 的儿子 巴勒 看见 以色列 向 亚摩利 人所做的一切。
NUM|22|3|摩押 因 以色列 百姓这么多，非常惧怕。 摩押 因 以色列 人的缘故就忧惧。
NUM|22|4|摩押 对 米甸 的长老说：“现在这群人要舔尽我们四围的一切，好像牛舔尽田间的草一样。” 那时， 西拨 的儿子 巴勒 作 摩押 王。
NUM|22|5|他派使者往 大河 附近的 毗夺 去，到 比珥 的儿子 巴兰 的家乡 ，召 巴兰 来，说：“看哪，有一群百姓从 埃及 出来；看哪，他们遮满地面，住在我的对面。
NUM|22|6|现在请你来，为我诅咒这百姓，因为他们比我强大，或许我能打败他们，把他们赶出此地。因为我知道，你为谁祝福，谁就得福；你诅咒谁，谁就受诅咒。”
NUM|22|7|摩押 的长老和 米甸 的长老手里拿着占卜的礼金到 巴兰 那里，将 巴勒 的话告诉他。
NUM|22|8|巴兰 对他们说：“今晚你们在这里过夜，我必照着耶和华向我说的话给你们答覆。” 摩押 的官员就在 巴兰 那里住下。
NUM|22|9|上帝临到 巴兰 那里，说：“你这里的这些人是谁？”
NUM|22|10|巴兰 对上帝说：“ 摩押 王 西拨 的儿子 巴勒 送信给我：
NUM|22|11|‘看哪，从 埃及 出来的百姓遮满了地面，现在请你来，为我诅咒他们，或许我能打败他们，把他们赶走。’”
NUM|22|12|上帝对 巴兰 说：“你不可跟他们去，也不可诅咒这百姓，因为他们是蒙福的。”
NUM|22|13|巴兰 早晨起来，对 巴勒 的官员说：“你们回本地去吧，因为耶和华不允许我和你们一起去。”
NUM|22|14|摩押 的官员就起来，到 巴勒 那里，说：“ 巴兰 不肯和我们一起来。”
NUM|22|15|巴勒 又差遣比这些更多，更尊贵的官员。
NUM|22|16|他们来到 巴兰 那里，对他说：“ 西拨 的儿子 巴勒 这样说：‘请你不要再推辞到我这里来！
NUM|22|17|我必使你得极大的尊荣，无论你向我要什么，我都给你。只求你来为我诅咒这百姓。’”
NUM|22|18|巴兰 回答 巴勒 的臣仆说：“ 巴勒 就是将他满屋的金银给我，我也不能做任何大小的事，违背耶和华－我上帝的指示。
NUM|22|19|现在请你们今晚也在这里住下，我好知道耶和华还要对我说什么。”
NUM|22|20|上帝在夜里临到 巴兰 那里，说：“这些人若来求你，你就起来跟他们去吧，只是你必须照着我对你说的话去做。”
NUM|22|21|巴兰 早晨起来，备了驴，就和 摩押 的官员一同去了。
NUM|22|22|上帝因他去就怒气发作；耶和华的使者站在路中间敌对他。他骑着驴，有两个仆人跟随他。
NUM|22|23|驴看见耶和华的使者站在路中间，手里有拔出来的刀，就离开了路，岔入田间。 巴兰 就打驴，要它回到路上。
NUM|22|24|耶和华的使者站在葡萄园的窄路上，这边有墙，那边也有墙。
NUM|22|25|驴看见耶和华的使者，就往墙挤去，把 巴兰 的脚挤到墙上； 巴兰 再打驴。
NUM|22|26|耶和华的使者又往前去，站在狭窄的地方，那里左右都无路可转。
NUM|22|27|驴看见耶和华的使者，就伏在 巴兰 底下。 巴兰 怒气发作，用杖打驴。
NUM|22|28|耶和华使驴开口，对 巴兰 说：“我向你做了什么，你竟打我这三次呢？”
NUM|22|29|巴兰 对驴说：“因为你戏弄我，我恨不得手中有刀，现在就把你杀了。”
NUM|22|30|驴对 巴兰 说：“我不是你从小直到今天所骑的驴吗？我平时有这样待过你吗？” 巴兰 说：“没有。”
NUM|22|31|耶和华使 巴兰 的眼目明亮，他看见耶和华的使者站在路中间，手里有拔出来的刀； 巴兰 就低头俯伏下拜。
NUM|22|32|耶和华的使者对他说：“你为什么这三次打你的驴呢？看哪，我出来敌对你，因为这路在我面前已经偏离了。
NUM|22|33|驴看见我就从我面前回避了这三次；驴若没有回避我，我早把你杀了，留它存活。”
NUM|22|34|巴兰 对耶和华的使者说：“我有罪了。我不知道你站在路中间阻挡我；现在你若看为不好，我就回去。”
NUM|22|35|耶和华的使者对 巴兰 说：“你和这些人去吧！你只要说我对你说的话。”于是 巴兰 和 巴勒 的官员一同去了。
NUM|22|36|巴勒 听见 巴兰 来了，就到 摩押 的城 去迎接他；这城是在边界的 亚嫩河 旁。
NUM|22|37|巴勒 对 巴兰 说：“我不是急切地派人到你那里去召你吗？你为何不到我这里来呢？我岂不能使你得尊荣吗？”
NUM|22|38|巴兰 对 巴勒 说：“看哪，我已经到你这里来了！现在我岂能擅自说什么呢？上帝将什么话放在我口中，我就说什么。”
NUM|22|39|巴兰 和 巴勒 同去，来到 基列．胡琐 。
NUM|22|40|巴勒 宰了牛羊为祭物，送给 巴兰 和陪伴他的官员。
NUM|22|41|到了早晨， 巴勒 领 巴兰 到 巴末．巴力 ，从那里可以看到一部分 以色列 的百姓。
NUM|23|1|巴兰 对 巴勒 说：“你要在这里为我筑七座坛，又要在这里为我预备七头公牛，七只公羊。”
NUM|23|2|巴勒 照 巴兰 的话做了。 巴勒 和 巴兰 在每座坛上献一头公牛，一只公羊。
NUM|23|3|巴兰 对 巴勒 说：“你站在你的燔祭旁边，我要往前去，或许耶和华会向我显现。他指示我什么事，我必告诉你。”于是 巴兰 上到一个光秃的高地。
NUM|23|4|上帝向 巴兰 显现。 巴兰 对他说：“我预备了七座坛，在每座坛上献了一头公牛，一只公羊。”
NUM|23|5|耶和华把话放在 巴兰 口中，说：“你回到 巴勒 那里，要这样说。”
NUM|23|6|他就回到 巴勒 那里，看哪， 巴勒 和 摩押 的众官员站在燔祭旁边。
NUM|23|7|巴兰 唱起诗歌说： “ 巴勒 领我出 亚兰 ， 摩押 王领我出东方的山脉： ‘来啊，为我诅咒 雅各 ； 来啊，怒骂 以色列 。’
NUM|23|8|上帝没有诅咒的， 我焉能诅咒？ 耶和华没有怒骂的， 我岂能怒骂？
NUM|23|9|我从磐石的巅峰看到他， 我从山丘望见他。 看哪，这是独居的民， 不算在列国中。
NUM|23|10|谁能数点 雅各 的尘土？ 谁能计算 以色列 的尘沙 ？ 我愿如正直人之死而死； 我愿如正直人之终而终。”
NUM|23|11|巴勒 对 巴兰 说：“你向我做的是什么呢？我带你来诅咒我的仇敌，看哪，你竟为他们祝福。”
NUM|23|12|他回答说：“耶和华放在我口中的话，我岂能不谨慎地说呢？”
NUM|23|13|巴勒 对他说：“请你跟我到别的地方，在那里可以看见他们。你只能看见他们的一部分，却不能看见全部。请你在那里为我诅咒他们。”
NUM|23|14|于是 巴勒 领 巴兰 到了 琐腓 的田野，上了 毗斯迦山 顶 ，筑了七座坛，在每座坛上献一头公牛，一只公羊。
NUM|23|15|巴兰 对 巴勒 说：“你站在你的燔祭旁边，我要到那边去看看。”
NUM|23|16|耶和华向 巴兰 显现，把话放在他口中，说：“你回到 巴勒 那里，要这样说。”
NUM|23|17|他回到 巴勒 那里，看哪， 巴勒 站在燔祭旁边， 摩押 的官员也和他在一起。 巴勒 对他说：“耶和华说了什么呢？”
NUM|23|18|巴兰 唱起诗歌说： “ 巴勒 啊，起来，听； 西拨 的儿子啊，侧耳听我。
NUM|23|19|上帝非人，必不致说谎， 也非人子，必不致后悔。 他说了岂不照着做呢？ 他发了言岂不实现呢？
NUM|23|20|看哪，我奉命祝福； 上帝赐福，我不能扭转。
NUM|23|21|他未见 雅各 中有灾难 ， 也未见 以色列 中有祸患 。 耶和华－他的上帝和他同在； 在他中间有欢呼王的声音。
NUM|23|22|上帝领他们出 埃及 ， 为 以色列 有如野牛的角。
NUM|23|23|绝没有法术可以伤 雅各 ， 没有占卜可以害 以色列 。 现在，人论及 雅各 ，论及 以色列 必说： ‘上帝成就了何等的事啊！’
NUM|23|24|看哪，这百姓兴起如母狮， 挺身像公狮， 未曾吃猎物， 未曾喝被杀者的血， 绝不躺卧。”
NUM|23|25|巴勒 对 巴兰 说：“你一点也不要诅咒他们，一点也不要为他们祝福！”
NUM|23|26|巴兰 回答 巴勒 说：“我不是告诉过你：‘凡耶和华所说的，我必须遵行’吗？”
NUM|23|27|巴勒 对 巴兰 说：“来，我领你到别的地方，或许上帝喜欢你在那里为我诅咒他们。”
NUM|23|28|巴勒 就领 巴兰 到那可了望旷野的 毗珥山 顶。
NUM|23|29|巴兰 对 巴勒 说：“你要在这里为我筑七座坛，又要在这里为我预备七头公牛，七只公羊。”
NUM|23|30|巴勒 就照 巴兰 的话做，在每座坛上献一头公牛，一只公羊。
NUM|24|1|巴兰 见耶和华喜欢赐福给 以色列 ，就不像前两次去求法术，却面向旷野。
NUM|24|2|巴兰 举目，看见 以色列 人照着支派扎营。上帝的灵就临到他身上，
NUM|24|3|他唱起诗歌说： “ 比珥 的儿子 巴兰 说， 眼目关闭 的人说，
NUM|24|4|听见上帝的言语， 得见全能者的异象， 俯伏着，眼睛却睁开的人说：
NUM|24|5|雅各 啊，你的帐棚何等华美！ 以色列 啊，你的帐幕何其华丽！
NUM|24|6|如连绵的山谷， 如河畔的园子， 如耶和华栽种的沉香树， 又如水边的香柏木。
NUM|24|7|水要从他的桶里流出， 种子要撒在多水之处。 他的王必超越 亚甲 ， 他的国必要振兴。
NUM|24|8|上帝领他出 埃及 ， 为他有如野牛的角。 他要吞灭那敌对他的国， 压碎他们的骨头， 用箭射透他们。
NUM|24|9|他蹲如公狮， 卧如母狮， 谁敢惹他？ 凡为你祝福的，愿他蒙福； 凡诅咒你的，愿他受诅咒。”
NUM|24|10|巴勒 向 巴兰 怒气发作，就紧握拳头 。 巴勒 对 巴兰 说：“我召你来诅咒我的仇敌，看哪，你竟然这三次为他们祝福。
NUM|24|11|如今你赶快回本地去吧！我想使你大得尊荣，看哪，耶和华却阻止你得尊荣。”
NUM|24|12|巴兰 对 巴勒 说：“我不是对你所差遣到我那里的使者说：
NUM|24|13|‘ 巴勒 就是把他满屋的金银给我，我也不能违背耶和华的指示，随自己的心意做好做歹。耶和华说什么，我就说什么。’
NUM|24|14|现在，看哪，我要回到我的百姓那里。来，让我告诉你这百姓日后要怎样对待你的百姓。”
NUM|24|15|他就唱起诗歌说： “ 比珥 的儿子 巴兰 说， 眼目关闭的人说，
NUM|24|16|听见上帝的言语， 明白至高者的知识， 看见全能者的异象， 俯伏着，眼睛却睁开的人说：
NUM|24|17|我看见他，却不在现时； 我望见他，却不在近处。 有星出于 雅各 ， 有杖从 以色列 兴起， 必打破 摩押 的额头， 必毁坏所有的 塞特 人 。
NUM|24|18|以东 将成为产业， 西珥 将成为它敌人的产业 ； 但 以色列 却要得胜。
NUM|24|19|有一位出于 雅各 的，必掌大权， 他要除灭城中的幸存者。”
NUM|24|20|巴兰 看见 亚玛力 人，就唱起诗歌说： “ 亚玛力 是诸国之首， 但它终必永远沉沦 。”
NUM|24|21|巴兰 看见 基尼 人，就唱起诗歌说： “你的住处坚固； 你的巢窝造在岩石中。
NUM|24|22|然而 基尼 族 必被吞灭， 直到何时 亚述 把你掳去？ ”
NUM|24|23|巴兰 又唱起诗歌说： “哀哉！若上帝做这事， 谁能存活呢？
NUM|24|24|有船只 从 基提 边界来到， 要压制 亚述 ， 要压制 希伯 ； 他也必永远沉沦 。”
NUM|24|25|于是 巴兰 起来，回本地去； 巴勒 也回他的路去了。
NUM|25|1|以色列 人住在 什亭 ，百姓开始与 摩押 女子行淫。
NUM|25|2|这些女子请百姓一同为她们的神明献祭，百姓吃了祭物，跪拜她们的神明。
NUM|25|3|以色列 与 巴力．毗珥 联合，耶和华的怒气就向 以色列 发作。
NUM|25|4|耶和华对 摩西 说：“拿下百姓中所有的领袖，对着太阳把他们悬挂在我面前，使我向 以色列 所发的怒气可以平息。”
NUM|25|5|于是 摩西 对 以色列 的审判官说：“你们的人若有与 巴力．毗珥 联合的，你们各人就要把他们杀了。”
NUM|25|6|摩西 和 以色列 全会众在会幕门口哭泣的时候，看哪，有一个 以色列 人，在他们眼前带着一个 米甸 女子，到他弟兄那里。
NUM|25|7|亚伦 祭司的孙子， 以利亚撒 的儿子 非尼哈 看见了，就从会众中起来，手里拿着枪，
NUM|25|8|跟这 以色列 人进入帐棚，刺穿了二人，就是 以色列 人和那女子的肚腹。这样， 以色列 人遭受的瘟疫就停止了。
NUM|25|9|遭瘟疫死的，有二万四千人。
NUM|25|10|耶和华吩咐 摩西 说：
NUM|25|11|“ 亚伦 祭司的孙子， 以利亚撒 的儿子 非尼哈 ，使我的愤怒转离 以色列 人，因为在他们中间，他以我的妒忌为他的妒忌，使我不在妒忌中毁灭 以色列 人。
NUM|25|12|因此，你要说：‘看哪，我将我平安的约赐给他。
NUM|25|13|这是他和他的后裔永远当祭司职任的约，因他为了上帝而妒忌，他为 以色列 人赎罪。’”
NUM|25|14|那与 米甸 女子一起被杀的 以色列 人，名叫 心利 ，是 撒路 的儿子，是 西缅 一个父家的领袖。
NUM|25|15|那被杀的 米甸 女子，名叫 哥斯比 ，是 苏珥 的女儿； 苏珥 是 米甸 一个父家的领袖。
NUM|25|16|耶和华吩咐 摩西 说：
NUM|25|17|“你要苦害 米甸 人，击杀他们；
NUM|25|18|因为他们用诡计苦害你们，在 毗珥 的事上和他们的姊妹， 米甸 领袖的女儿 哥斯比 的事上，欺骗了你们；在瘟疫的日子，这女子因 毗珥 的事件被杀了。”
NUM|26|1|瘟疫过了之后，耶和华对 摩西 和 亚伦 祭司的儿子 以利亚撒 说：
NUM|26|2|“你们要将 以色列 全会众，按他们的父家，凡二十岁以上能出去为 以色列 打仗的，计算总数。”
NUM|26|3|摩西 和 以利亚撒 祭司在 摩押 平原与 耶利哥 相对的 约旦河 边吩咐他们说：
NUM|26|4|“计算你们中间从二十岁以上的人数。”正如耶和华所吩咐 摩西 的。 从 埃及 地出来的 以色列 人如下：
NUM|26|5|以色列 的长子是 吕便 。 吕便 的众子：属 哈诺 的，有 哈诺 族；属 法路 的，有 法路 族；
NUM|26|6|属 希斯伦 的，有 希斯伦 族；属 迦米 的，有 迦米 族。
NUM|26|7|这就是 吕便 的各族；被数的共有四万三千七百三十名。
NUM|26|8|法路 的儿子是 以利押 。
NUM|26|9|以利押 的儿子是 尼母利 、 大坍 、 亚比兰 。这 大坍 、 亚比兰 ，就是从会中选出来，当 可拉 一伙的人向耶和华争闹的时候，一起向 摩西 、 亚伦 争闹的；
NUM|26|10|地开了裂口，吞了他们和 可拉 ， 可拉 一伙的人也一同死亡。当时火吞灭了二百五十个人；他们就成为鉴戒。
NUM|26|11|然而 可拉 的众子没有死亡。
NUM|26|12|按着宗族， 西缅 的众子：属 尼母利 的，有 尼母利 族；属 雅悯 的，有 雅悯 族；属 雅斤 的，有 雅斤 族；
NUM|26|13|属 谢拉 的，有 谢拉 族；属 扫罗 的，有 扫罗 族。
NUM|26|14|这就是 西缅 的各族，共有二万二千二百名。
NUM|26|15|按着宗族， 迦得 的众子：属 洗分 的，有 洗分 族；属 哈基 的，有 哈基 族；属 书尼 的，有 书尼 族；
NUM|26|16|属 阿斯尼 的，有 阿斯尼 族；属 以利 的，有 以利 族；
NUM|26|17|属 亚律 的，有 亚律 族；属 亚列利 的，有 亚列利 族。
NUM|26|18|这就是 迦得 子孙的各族；他们被数的共有四万零五百名。
NUM|26|19|犹大 的儿子是 珥 和 俄南 。 珥 和 俄南 死在 迦南 地。
NUM|26|20|按着宗族， 犹大 的众子：属 示拉 的，有 示拉 族；属 法勒斯 的，有 法勒斯 族；属 谢拉 的，有 谢拉 族。
NUM|26|21|法勒斯 的众子：属 希斯仑 的，有 希斯仑 族；属 哈母勒 的，有 哈母勒 族。
NUM|26|22|这就是 犹大 的各族；他们被数的共有七万六千五百名。
NUM|26|23|按着宗族， 以萨迦 的众子：属 陀拉 的，有 陀拉 族；属 普瓦 的，有 普瓦 族；
NUM|26|24|属 雅述 的，有 雅述 族；属 伸仑 的，有 伸仑 族。
NUM|26|25|这就是 以萨迦 的各族；他们被数的共有六万四千三百名。
NUM|26|26|按着宗族， 西布伦 的众子：属 西烈 的，有 西烈 族；属 以伦 的，有 以伦 族；属 雅利 的，有 雅利 族。
NUM|26|27|这就是 西布伦 的各族；他们被数的共有六万零五百名。
NUM|26|28|按着宗族， 约瑟 的儿子有 玛拿西 、 以法莲 。
NUM|26|29|玛拿西 的众子：属 玛吉 的，有 玛吉 族； 玛吉 生 基列 ；属 基列 的，有 基列 族。
NUM|26|30|这就是 基列 的众子：属 伊以谢 的，有 伊以谢 族；属 希勒 的，有 希勒 族；
NUM|26|31|属 亚斯烈 的，有 亚斯烈 族；属 示剑 的，有 示剑 族；
NUM|26|32|属 示米大 的，有 示米大 族；属 希弗 的，有 希弗 族。
NUM|26|33|希弗 的儿子 西罗非哈 没有儿子，只有女儿。 西罗非哈 的女儿的名字是 玛拉 、 挪阿 、 曷拉 、 密迦 、 得撒 。
NUM|26|34|这就是 玛拿西 的各族；他们被数的共有五万二千七百名。
NUM|26|35|这就是按着宗族， 以法莲 的众子：属 书提拉 的，有 书提拉 族；属 比结 的，有 比结 族；属 他罕 的，有 他罕 族。
NUM|26|36|这就是 书提拉 的众子：属 以兰 的，有 以兰 族。
NUM|26|37|这就是 以法莲 子孙的各族；他们被数的共有三万二千五百名。按着宗族，以上这些都是 约瑟 的子孙。
NUM|26|38|按着宗族， 便雅悯 的众子：属 比拉 的，有 比拉 族；属 亚实别 的，有 亚实别 族；属 亚希兰 的，有 亚希兰 族；
NUM|26|39|属 书反 的，有 书反 族；属 户反 的，有 户反 族。
NUM|26|40|比拉 的儿子是 亚勒 、 乃幔 ；属 亚勒 的 ，有 亚勒 族；属 乃幔 的，有 乃幔 族。
NUM|26|41|按着宗族，这就是 便雅悯 的子孙；他们被数的共有四万五千六百名。
NUM|26|42|这就是按着宗族， 但 的众子：属 书含 的，有 书含 族。按着宗族，这就是 但 的各族。
NUM|26|43|按照他们被数的， 书含 全宗族共有六万四千四百名。
NUM|26|44|按着宗族， 亚设 的众子：属 音拿 的，有 音拿 族；属 亦施韦 的，有 亦施韦 族；属 比利亚 的，有 比利亚 族。
NUM|26|45|比利亚 的众子：属 希别 的，有 希别 族；属 玛结 的，有 玛结 族。
NUM|26|46|亚设 的女儿名叫 西拉 。
NUM|26|47|这就是 亚设 子孙的各族；他们被数的共有五万三千四百名。
NUM|26|48|按着宗族， 拿弗他利 的众子：属 雅薛 的，有 雅薛 族；属 沽尼 的，有 沽尼 族；
NUM|26|49|属 耶色 的，有 耶色 族；属 示冷 的，有 示冷 族。
NUM|26|50|按着宗族，这就是 拿弗他利 的各族；他们被数的共有四万五千四百名。
NUM|26|51|这就是 以色列 人中被数的，共有六十万零一千七百三十名。
NUM|26|52|耶和华吩咐 摩西 说：
NUM|26|53|“你要按着人名的数目，将地分给这些人为产业。
NUM|26|54|人多的要多给他们产业，人少的要少给他们产业；各照被数的人数分配产业。
NUM|26|55|此外，要以抽签来分地，按着父系各支派的名字承受产业。
NUM|26|56|要根据抽签，看人数的多寡，给他们分配产业。”
NUM|26|57|这就是按着宗族，被数的 利未 人：属 革顺 的，有 革顺 族；属 哥辖 的，有 哥辖 族；属 米拉利 的，有 米拉利 族。
NUM|26|58|这就是 利未 的宗族： 立尼 族、 希伯伦 族、 玛利 族、 母示 族、 可拉 族。 哥辖 生 暗兰 。
NUM|26|59|暗兰 的妻子名叫 约基别 ，是 利未 的女儿，是 利未 在 埃及 所生的。她给 暗兰 生了 亚伦 、 摩西 ，和他们的姊姊 米利暗 。
NUM|26|60|亚伦 生 拿答 、 亚比户 、 以利亚撒 、 以他玛 。
NUM|26|61|拿答 、 亚比户 在耶和华面前献凡火的时候死了。
NUM|26|62|利未 人中，凡一个月以上所有被数的男子，共有二万三千名。他们没有数在 以色列 人中；因为在 以色列 人中，没有分给他们产业。
NUM|26|63|这些是 摩西 和 以利亚撒 祭司所数的；他们在 摩押 平原与 耶利哥 相对的 约旦河 边数点 以色列 人。
NUM|26|64|这些被数的人中，没有一个是 摩西 和 亚伦 祭司先前在 西奈 旷野所数的 以色列 人，
NUM|26|65|因为耶和华论到他们说：“他们必死在旷野。”所以，除了 耶孚尼 的儿子 迦勒 和 嫩 的儿子 约书亚 以外，他们一个也没有存留。
NUM|27|1|约瑟 的儿子 玛拿西 的宗族中，有 玛拿西 的玄孙， 玛吉 的曾孙， 基列 的孙子， 希弗 的儿子 西罗非哈 的女儿，名叫 玛拉 、 挪阿 、 曷拉 、 密迦 、 得撒 。她们前来，
NUM|27|2|站在会幕门口，在 摩西 和 以利亚撒 祭司，以及众领袖与全会众面前，说：
NUM|27|3|“我们的父亲死在旷野。他没有与 可拉 同伙聚集攻击耶和华，是在自己的罪中死的；他没有儿子。
NUM|27|4|为什么因我们的父亲没有儿子就把他的名从他族中除掉呢？求你们在我们父亲的兄弟中分给我们产业。”
NUM|27|5|于是， 摩西 将她们的案件呈到耶和华面前。
NUM|27|6|耶和华对 摩西 说：
NUM|27|7|“ 西罗非哈 的女儿说得有理。你定要在她们父亲的兄弟中，把地分给她们为业，把她们父亲的产业传给她们。
NUM|27|8|你也要吩咐 以色列 人说：‘人死了，若没有儿子，就要把他的产业传给他的女儿。
NUM|27|9|他若没有女儿，就要把他的产业给他的兄弟。
NUM|27|10|他若没有兄弟，就要把他的产业给他父亲的兄弟。
NUM|27|11|他父亲若没有兄弟，就要把他的产业给他族中最近的亲属继承为业。’”这要作 以色列 人的律例典章，是照耶和华所吩咐 摩西 的。
NUM|27|12|耶和华对 摩西 说：“你上这 亚巴琳山脉 ，看我所赐给 以色列 人的地。
NUM|27|13|看了以后，你也必归到你祖先 那里，像你哥哥 亚伦 归去一样。
NUM|27|14|因为你们在 寻 的旷野，当会众争闹的时候，违背了我的命令，在取水之事上没有在会众眼前尊我为圣。”这水就是 寻 的旷野中， 加低斯 的 米利巴 水。
NUM|27|15|摩西 对耶和华说：
NUM|27|16|“愿耶和华，赐万人气息的上帝，立一个人治理会众，
NUM|27|17|可以在他们面前出入，引导他们进出，免得耶和华的会众如同没有牧人的羊群一般。”
NUM|27|18|耶和华对 摩西 说：“ 嫩 的儿子 约书亚 是一个有圣灵的人；你要领他来，为他按手，
NUM|27|19|使他站在 以利亚撒 祭司和全会众面前，在他们眼前委派他，
NUM|27|20|又将你的尊荣给他一些，好使 以色列 全会众都听从他。
NUM|27|21|他要站在 以利亚撒 祭司面前； 以利亚撒 要凭乌陵的判断，在耶和华面前为他求问。他和 以色列 全会众都要照 以利亚撒 的指示出入。”
NUM|27|22|于是 摩西 照耶和华所吩咐他的，将 约书亚 领来，使他站在 以利亚撒 祭司和全会众面前，
NUM|27|23|为他按手，委派他，是照耶和华藉 摩西 所说的。
NUM|28|1|耶和华吩咐 摩西 说：
NUM|28|2|“你要吩咐 以色列 人说：‘你们要按时把我的供物，就是献给我作馨香火祭的食物，献给我。’
NUM|28|3|要对他们说：‘这是当献给耶和华的火祭：每天两只没有残疾一岁的小公羊，作为经常献的燔祭。
NUM|28|4|早晨献第一只小公羊，黄昏献第二只小公羊；
NUM|28|5|又用十分之一伊法细面和四分之一欣捣成的油，调和作为素祭。
NUM|28|6|这是在 西奈山 上规定为经常献的燔祭，是献给耶和华为馨香的火祭。
NUM|28|7|为每只小公羊，要有四分之一欣的浇酒祭；在圣所中，你要将醇酒献给耶和华作浇酒祭。
NUM|28|8|黄昏你献第二只小公羊，要照早晨的素祭和同献的浇酒祭献上，作为馨香的火祭，献给耶和华。’”
NUM|28|9|“在安息日，要献两只没有残疾，一岁的小公羊、十分之二伊法调了油的细面为素祭，和同献的浇酒祭。
NUM|28|10|除了经常献的燔祭和同献的浇酒祭之外，这是每一个安息日当献的燔祭。”
NUM|28|11|“每月初一，要将两头公牛犊、一只公绵羊、七只没有残疾一岁的小公羊，献给耶和华为燔祭。
NUM|28|12|为每头公牛，要用十分之三伊法调了油的细面作为素祭；为那只公绵羊，要用十分之二伊法调了油的细面作为素祭；
NUM|28|13|为每只小公羊，要用十分之一伊法调了油的细面作为素祭。这是馨香的燔祭，是献给耶和华的火祭。
NUM|28|14|每头公牛要有半欣的浇酒祭，每只公绵羊三分之一欣的浇酒祭，每只小公羊四分之一欣的浇酒祭。这是一年之中每月初一当献的燔祭。
NUM|28|15|除了经常献的燔祭和同献的浇酒祭之外，又要将一只公山羊，献给耶和华为赎罪祭。”
NUM|28|16|“正月十四日是向耶和华守的逾越节。
NUM|28|17|这月十五日是节期，要吃无酵饼七日。
NUM|28|18|第一日要有圣会，任何劳动的工都不可做。
NUM|28|19|要把火祭，就是两头公牛犊，一只公绵羊、七只一岁的小公羊，都要没有残疾的，献给耶和华为燔祭。
NUM|28|20|要同时献调了油的细面为素祭：每头公牛要献十分之三伊法；每只公绵羊要献十分之二伊法；
NUM|28|21|为那七只小公羊，每只要献十分之一伊法。
NUM|28|22|此外，要献一只公山羊作赎罪祭，为你们赎罪。
NUM|28|23|除了早晨经常献的燔祭之外，你们也要献这些祭。
NUM|28|24|一连七天，在经常献的燔祭和同献的浇酒祭之外，每天要这样把馨香火祭的食物献给耶和华。
NUM|28|25|第七日要有圣会，任何劳动的工都不可做。”
NUM|28|26|“七七初熟节，就是你们献初熟谷物给耶和华为素祭的那一天，要宣告圣会；任何劳动的工都不可做。
NUM|28|27|要将两头公牛犊，一只公绵羊，七只一岁的小公羊，作为馨香的燔祭献给耶和华。
NUM|28|28|要同时献调了油的细面为素祭：每头公牛要献十分之三伊法；每只公绵羊要献十分之二伊法；
NUM|28|29|为那七只小公羊，每只要献十分之一伊法。
NUM|28|30|此外，要献一只公山羊为你们赎罪。
NUM|28|31|除了经常献的燔祭和同献的素祭，你们也要献上这些没有残疾的，和同献的浇酒祭。”
NUM|29|1|“七月初一，你们当有圣会；任何劳动的工都不可做，是你们当守为吹角的日子。
NUM|29|2|你们要将一头公牛犊、一只公绵羊、七只一岁的小公羊，都是没有残疾的，献给耶和华为馨香的燔祭。
NUM|29|3|要同时献调了油的细面为素祭：每头公牛要献十分之三伊法；每只公绵羊要献十分之二伊法；
NUM|29|4|为那七只小公羊，每只要献十分之一伊法。
NUM|29|5|此外，要献一只公山羊作赎罪祭，为你们赎罪。
NUM|29|6|除了初一的燔祭和同献的素祭、经常献的燔祭与同献的素祭，以及同献的浇酒祭以外，这些都照例作为馨香的火祭献给耶和华。”
NUM|29|7|“七月初十，你们当有圣会；要刻苦己心，任何工都不可做。
NUM|29|8|要将一头公牛犊、一只公绵羊、七只一岁的小公羊，都是没有残疾的，献给耶和华为馨香的燔祭。
NUM|29|9|要同时献调了油的细面为素祭：每头公牛要献十分之三伊法；每只公绵羊要献十分之二伊法；
NUM|29|10|为那七只小公羊，每只要献十分之一伊法。
NUM|29|11|又要献一只公山羊为赎罪祭。这是在赎罪祭和经常献的燔祭，以及同献的素祭和浇酒祭以外所献的。”
NUM|29|12|“七月十五日，你们当有圣会；任何劳动的工都不可做，要向耶和华守节七天。
NUM|29|13|要将十三头公牛犊、两只公绵羊、十四只一岁的小公羊，都是没有残疾的，献上作火祭，是献给耶和华馨香的燔祭。
NUM|29|14|要同时献调了油的细面为素祭：为那十三头公牛犊，每头要献十分之三伊法；为那两只公绵羊，每只要献十分之二伊法；
NUM|29|15|为那十四只小公羊，每只要献十分之一伊法。
NUM|29|16|又要献一只公山羊为赎罪祭。这是在经常献的燔祭、同献的素祭和浇酒祭以外所献的。
NUM|29|17|“第二日要献十二头公牛犊、两只公绵羊、十四只一岁的小公羊，都是没有残疾的，
NUM|29|18|并为公牛、公绵羊和小公羊，按数照例奉献同献的素祭和浇酒祭。
NUM|29|19|又要献一只公山羊为赎罪祭。这是在经常献的燔祭、同献的素祭和浇酒祭以外所献的。
NUM|29|20|“第三日要献十一头公牛、两只公绵羊、十四只一岁的小公羊，都是没有残疾的，
NUM|29|21|并为公牛、公绵羊和小公羊，按数照例奉献同献的素祭和浇酒祭。
NUM|29|22|又要献一只公山羊为赎罪祭。这是在经常献的燔祭、同献的素祭和浇酒祭以外所献的。
NUM|29|23|“第四日要献十头公牛、两只公绵羊、十四只一岁的小公羊，都是没有残疾的，
NUM|29|24|并为公牛、公绵羊和小公羊，按数照例奉献同献的素祭和浇酒祭。
NUM|29|25|又要献一只公山羊为赎罪祭。这是在经常献的燔祭、同献的素祭和浇酒祭以外所献的。
NUM|29|26|“第五日要献九头公牛、两只公绵羊、十四只一岁的小公羊，都是没有残疾的，
NUM|29|27|并为公牛、公绵羊和小公羊，按数照例奉献同献的素祭和浇酒祭。
NUM|29|28|又要献一只公山羊为赎罪祭。这是在经常献的燔祭、同献的素祭和浇酒祭以外所献的。
NUM|29|29|“第六日要献八头公牛、两只公绵羊、十四只一岁的小公羊，都是没有残疾的，
NUM|29|30|并为公牛、公绵羊和小公羊，按数照例奉献同献的素祭和浇酒祭。
NUM|29|31|又要献一只公山羊为赎罪祭。这是在经常献的燔祭、同献的素祭和浇酒祭以外所献的。
NUM|29|32|“第七日要献七头公牛、两只公绵羊、十四只一岁的小公羊，都是没有残疾的，
NUM|29|33|并为公牛、公绵羊和小公羊，按数照例奉献同献的素祭和浇酒祭。
NUM|29|34|又要献一只公山羊为赎罪祭。这是在经常献的燔祭、同献的素祭和浇酒祭以外所献的。
NUM|29|35|“第八日你们当有严肃会；任何劳动的工都不可做；
NUM|29|36|要将一头公牛、一只公绵羊、七只一岁的小公羊，都是没有残疾的，献上作火祭，是献给耶和华馨香的燔祭。
NUM|29|37|要为公牛、公绵羊和小公羊，按数照例奉献同献的素祭和浇酒祭。
NUM|29|38|又要献一只公山羊为赎罪祭。这是在经常献的燔祭、同献的素祭和浇酒祭以外所献的。
NUM|29|39|“这些祭要在你们的节期献给耶和华，都是在所许的愿和甘心献的以外所献的，作为你们的燔祭、素祭、浇酒祭和平安祭。”
NUM|29|40|于是， 摩西 照耶和华所吩咐他的一切话告诉 以色列 人。
NUM|30|1|摩西 对 以色列 各支派的领袖说：“这是耶和华所吩咐的话：
NUM|30|2|人若向耶和华许愿或起誓，要约束自己，就不可食言，必须照口中所出的一切话去做。
NUM|30|3|女子年轻，还在父家的时候，若向耶和华许愿，要约束自己，
NUM|30|4|她父亲听见她所许的愿和约束自己的话，却向她默默不言，她所许的愿和约束自己的话就都有效。
NUM|30|5|但是，若她父亲在听见的日子不允许她一切所许的愿和约束自己的话，这就不算为有效；耶和华也必赦免她，因为她的父亲不允许。
NUM|30|6|她若已出嫁，有愿在身，或口中出了约束自己的冒失话，
NUM|30|7|她丈夫听见了，却在听见的日子向她默默不言，她所许的愿和约束自己的话就都有效。
NUM|30|8|但是，若她丈夫在听见的日子不允许，丈夫就废了她所许的愿和口中所出约束自己的冒失话；耶和华也必赦免她。
NUM|30|9|寡妇或被休的妇人所许的愿，她所有约束自己的话，都是有效的。
NUM|30|10|她若在丈夫家里许了愿或起了誓，要约束自己，
NUM|30|11|丈夫听见了，却向她默默不言，没有不允许，她所许的愿和约束自己的话就都有效。
NUM|30|12|她丈夫听见的日子，若把这些全废了，她口中一切所许的愿或约束自己的话就不算为有效。她丈夫已把这些都废了，耶和华也必赦免她。
NUM|30|13|凡她所许的愿和刻苦约束自己所起的誓，丈夫可以坚立，也可以废去。
NUM|30|14|倘若她丈夫天天向她默默不言，这就算是坚立她一切所许的愿或约束自己的话；因为丈夫在听见的日子向她默默不言，就算是坚立了这些话。
NUM|30|15|但她丈夫听见了，以后若再废了这些话，就要担当妇人的罪孽。”
NUM|30|16|这是关于丈夫待妻子，父亲待女儿，女儿年轻还在父家，耶和华所吩咐 摩西 的条例。
NUM|31|1|耶和华吩咐 摩西 说：
NUM|31|2|“你要为 以色列 人向 米甸 人报仇，然后归到你祖先 那里。”
NUM|31|3|摩西 吩咐百姓说：“要在你们中间叫人带兵器去攻击 米甸 ，为耶和华向 米甸 报仇。
NUM|31|4|从 以色列 众支派中，每支派要派一千人去打仗。”
NUM|31|5|于是从 以色列 千万人中，每支派征召一千人，一共一万二千名，带着兵器预备打仗。
NUM|31|6|摩西 派他们去打仗，每支派一千人；又派 以利亚撒 祭司的儿子 非尼哈 同去； 非尼哈 手里拿着圣所的器皿和吹号的号筒。
NUM|31|7|他们遵照耶和华所吩咐 摩西 的，与 米甸 打仗，杀了所有的男丁。
NUM|31|8|在所杀的人中，他们杀了 米甸 的王，就是 以未 、 利金 、 苏珥 、 户珥 、 利巴 五个 米甸 的王，又用刀杀了 比珥 的儿子 巴兰 。
NUM|31|9|以色列 人掳了 米甸 的妇女和孩童，抢夺他们一切的牲畜、牛羊和所有的财物，
NUM|31|10|又用火焚烧了他们所住的一切城镇和所有的营寨。
NUM|31|11|以色列 人把一切掳物和掠物，连人和牲畜都带走，
NUM|31|12|将俘虏、掠物、掳物带到 摩押 平原，在 约旦河 边与 耶利哥 相对的营地，交给 摩西 和 以利亚撒 祭司，以及 以色列 的会众。
NUM|31|13|摩西 和 以利亚撒 祭司，以及会众中所有的领袖，都出营迎接他们。
NUM|31|14|摩西 向打仗回来的军官，就是千夫长和百夫长发怒。
NUM|31|15|摩西 对他们说：“你们要让这所有的妇女活着吗？
NUM|31|16|看哪，正是这些妇女，因 巴兰 的话，在 毗珥 的事上导致 以色列 人背叛耶和华，以致耶和华的会众遭遇瘟疫。
NUM|31|17|现在，你们要杀所有的男孩，也要把所有曾与男人同房共寝的女子都杀了。
NUM|31|18|但那些未曾与男人同房共寝的女孩，你们可以让她们存活。
NUM|31|19|你们和你们所掳来的人，要住在营外七天；凡杀了人的，和一切摸了尸体的，要在第三日和第七日洁净自己。
NUM|31|20|你们也要洁净一切的衣服，以及用皮革、山羊毛和木头做的任何东西。”
NUM|31|21|以利亚撒 祭司对打仗回来的士兵说：“耶和华所吩咐 摩西 律法中的条例是这样：
NUM|31|22|金、银、铜、铁、锡、铅，
NUM|31|23|凡能耐火的，你们要使它经过火，它就洁净，然而还要用除污秽的水来洁净它；凡不能耐火的，你们要使它经过水。
NUM|31|24|第七日，你们要洗衣服，才为洁净，然后可以进营。”
NUM|31|25|耶和华对 摩西 说：
NUM|31|26|“你和 以利亚撒 祭司，以及会众的各父系家长，要计算所掳掠的人和牲畜的总数。
NUM|31|27|要把所掳掠的分成两半：一半给那出去打仗的精兵，一半给全会众。
NUM|31|28|再从那出去打仗的战士所得的人、牛、驴、羊中，每五百取一，献给耶和华为贡物。
NUM|31|29|要从他们那一半中取出这些，交给 以利亚撒 祭司，作为耶和华的举祭。
NUM|31|30|又要从 以色列 人的那一半中，就是从人、牛、驴、羊，各样牲畜中，每五十取一，交给照管耶和华帐幕的 利未 人。”
NUM|31|31|于是 摩西 和 以利亚撒 祭司遵照耶和华所吩咐 摩西 的做了。
NUM|31|32|除了士兵所夺的财物以外，所掳来的有羊六十七万五千只，
NUM|31|33|牛七万二千头，
NUM|31|34|驴六万一千匹；
NUM|31|35|至于人，就是未曾与男人同房共寝的女子，总共三万二千名。
NUM|31|36|出去打仗之人的那分，就是他们所得的一半，共计羊三十三万七千五百只，
NUM|31|37|其中归耶和华为贡物的羊，六百七十五只；
NUM|31|38|牛三万六千头，其中归耶和华为贡物的七十二头；
NUM|31|39|驴三万零五百匹，其中归耶和华为贡物的六十一匹；
NUM|31|40|人一万六千名，其中归耶和华的三十二名。
NUM|31|41|摩西 把贡物，就是归给耶和华的举祭，交给 以利亚撒 祭司，是照耶和华所吩咐 摩西 的。
NUM|31|42|以色列 人所得的另一半，是 摩西 从打仗的人取来分给他们的。
NUM|31|43|会众的这一半有羊三十三万七千五百只，
NUM|31|44|牛三万六千头，
NUM|31|45|驴三万零五百匹，
NUM|31|46|人一万六千名。
NUM|31|47|无论是人或牲畜， 摩西 都每五十取一，交给照管耶和华帐幕的 利未 人，是照耶和华所吩咐 摩西 的。
NUM|31|48|带领众军队的军官，就是千夫长、百夫长，进到 摩西 那里，
NUM|31|49|对他说：“你的仆人已经计算属下战士的总数，一个也没有少。
NUM|31|50|如今我们把各人所得的金器，就是脚链子、手镯、打印的戒指、耳环、项链，都送给耶和华为供物，好在耶和华面前为我们赎罪。”
NUM|31|51|摩西 和 以利亚撒 祭司就收了他们的金子，就是各样的首饰。
NUM|31|52|千夫长、百夫长所献给耶和华为举祭的金子共有一万六千七百五十舍客勒。
NUM|31|53|打仗的人都把自己所掠夺的各自留下。
NUM|31|54|摩西 和 以利亚撒 祭司收了千夫长、百夫长的金子，就带进会幕，好使 以色列 人在耶和华面前蒙记念。
NUM|32|1|吕便 子孙和 迦得 子孙的牲畜极其众多。他们看到 雅谢 地和 基列 地；看哪，这是可牧放牲畜的地方。
NUM|32|2|吕便 子孙和 迦得 子孙就到 摩西 和 以利亚撒 祭司，以及会众的领袖那里，说：
NUM|32|3|“ 亚他录 、 底本 、 雅谢 、 宁拉 、 希实本 、 以利亚利 、 示班 、 尼波 、 比稳 ，
NUM|32|4|就是耶和华在 以色列 会众面前所攻取之地，是可牧放牲畜之地，而你的仆人也有牲畜。”
NUM|32|5|又说：“我们若在你眼前蒙恩，求你把这地给我们为业；不要领我们过 约旦河 。”
NUM|32|6|摩西 对 迦得 子孙和 吕便 子孙说：“难道你们的弟兄去打仗，你们却留在这里吗？
NUM|32|7|你们为什么使 以色列 人灰心，不渡过去，进入耶和华所赐给他们的那地呢？
NUM|32|8|我从 加低斯．巴尼亚 派你们的父执之辈去窥探那地时，他们就曾这样做过。
NUM|32|9|他们上到 以实各谷 ，窥探了那地之后，竟然使 以色列 人灰心，不愿进入耶和华所赐给他们的地。
NUM|32|10|当日，耶和华的怒气发作，起誓说：
NUM|32|11|‘凡从 埃及 上来二十岁以上的人，断不得看见我对 亚伯拉罕 、 以撒 、 雅各 起誓应许之地，因为他们没有专心跟从我；
NUM|32|12|惟有 基尼洗 族 耶孚尼 的儿子 迦勒 ，还有 嫩 的儿子 约书亚 可以看见，因为他们专心跟从耶和华。’
NUM|32|13|耶和华的怒气向 以色列 发作，使他们在旷野飘流四十年，直到在耶和华眼前作恶的那一代都消灭了。
NUM|32|14|看哪，你们这一伙罪人，竟然接续你们父执之辈，再增加耶和华对 以色列 所发的怒气。
NUM|32|15|你们若转离不跟从他，他要再把 以色列 人撇在旷野；这样，你们就使这众百姓灭亡了。”
NUM|32|16|他们挨近 摩西 ，说：“我们要在这里为牲畜筑圈，为孩童建城。
NUM|32|17|我们自己却要带兵器，急速行在 以色列 人的前面，领他们直到他们的地方。我们的孩童可以留在坚固的城内，躲避当地的居民。
NUM|32|18|我们必不回自己的家，直等到 以色列 人各自承受了自己的产业。
NUM|32|19|我们不和他们在 约旦河 那边分产业，因为我们的产业是在 约旦河 的东边。”
NUM|32|20|摩西 对他们说：“你们若要这么做，若要在耶和华面前带着兵器出去打仗，
NUM|32|21|你们中间所有带兵器的人都要在耶和华面前过 约旦河 ，直到耶和华把仇敌从他面前赶出去。
NUM|32|22|那地在耶和华面前被征服以后，你们方可回来。这样，你们向耶和华和 以色列 才算为无罪，这地也必在耶和华面前归你们为业。
NUM|32|23|倘若你们不这样做，看哪，你们就得罪了耶和华，当知道你们的罪必找上你们。
NUM|32|24|如今你们可以为孩童建城，为羊群筑圈，但你们口所讲出来的话，必须实践。”
NUM|32|25|迦得 子孙和 吕便 子孙对 摩西 说：“你的仆人们必照我主所吩咐的去做。
NUM|32|26|我们的孩子、妻子、牛羊和所有的牲畜都要留在 基列 的各城。
NUM|32|27|但你的仆人，凡能带兵器上战场的，都要照我主所说的话，在耶和华面前渡过去打仗。”
NUM|32|28|于是， 摩西 为他们吩咐 以利亚撒 祭司和 嫩 的儿子 约书亚 ，以及 以色列 人各支派父系的领袖。
NUM|32|29|摩西 对他们说：“ 迦得 子孙和 吕便 子孙，凡带兵器在耶和华面前去打仗的，若与你们一同渡过 约旦河 ，那地被你们征服以后，你们就要把 基列 地给他们为业。
NUM|32|30|倘若他们不带兵器与你们一同渡过去，他们就要在 迦南 地你们中间得产业。”
NUM|32|31|迦得 子孙和 吕便 子孙回答说：“耶和华怎样吩咐仆人，我们就必照样做。
NUM|32|32|我们自己必带着兵器，在耶和华面前渡过去，进入 迦南 地，好使我们在 约旦河 这边得到我们的产业。”
NUM|32|33|摩西 把 亚摩利 王 西宏 的国和 巴珊 王 噩 的国，就是他们的国土和周围的城镇，都给了 迦得 子孙和 吕便 子孙，以及 约瑟 的儿子 玛拿西 半个支派。
NUM|32|34|迦得 子孙建造了 底本 、 亚他录 、 亚罗珥 、
NUM|32|35|亚他录．朔反 、 雅谢 、 约比哈 、
NUM|32|36|伯．宁拉 、 伯．哈兰 ，都是坚固城，并筑有羊圈。
NUM|32|37|吕便 子孙建造了 希实本 、 以利亚利 、 基列亭 、
NUM|32|38|尼波 、 巴力．免 （名字是改了的）、 西比玛 ；他们给建造的城另起别名。
NUM|32|39|玛拿西 的儿子 玛吉 的子孙往 基列 去，占了那地，赶出那里的 亚摩利 人。
NUM|32|40|摩西 把 基列 赐给 玛拿西 的儿子 玛吉 ，他就住在那里。
NUM|32|41|玛拿西 的子孙 睚珥 占了 基列 的城镇，就称这些城镇为 哈倭特．睚珥 。
NUM|32|42|挪巴 占了 基纳 和 基纳 的乡镇，就照自己的名字称 基纳 为 挪巴 。
NUM|33|1|这是 以色列 人按着队伍，在 摩西 、 亚伦 的手下，出 埃及 地的行程。
NUM|33|2|摩西 遵照耶和华的指示记录他们每段行程的起点，这些行程的起点如下：
NUM|33|3|第一个月，就是正月十五日，逾越的第二天，他们从 兰塞 起行，在所有 埃及 人的眼前抬起头 来出去了。
NUM|33|4|那时， 埃及 人正埋葬他们的长子，就是耶和华在他们中间所击杀的；耶和华也惩治了他们的众神明。
NUM|33|5|以色列 人从 兰塞 起行，安营在 疏割 。
NUM|33|6|从 疏割 起行，安营在旷野边上的 以倘 。
NUM|33|7|从 以倘 起行，转向 巴力．洗分 对面的 比．哈希录 ，安营在 密夺 。
NUM|33|8|从 比．哈希录 起行，经过海，进入旷野，在 以倘 的旷野走了三天的路程，就安营在 玛拉 。
NUM|33|9|从 玛拉 起行，来到 以琳 ， 以琳 有十二股水泉，七十棵棕树，就安营在那里。
NUM|33|10|从 以琳 起行，安营在 红海 边。
NUM|33|11|从 红海 边起行，安营在 汛 的旷野。
NUM|33|12|从 汛 的旷野起行，安营在 脱加 。
NUM|33|13|从 脱加 起行，安营在 亚录 。
NUM|33|14|从 亚录 起行，安营在 利非订 ；在那里，百姓没有水喝。
NUM|33|15|从 利非订 起行，安营在 西奈 的旷野。
NUM|33|16|从 西奈 的旷野起行，安营在 基博罗．哈他瓦 。
NUM|33|17|从 基博罗．哈他瓦 起行，安营在 哈洗录 。
NUM|33|18|从 哈洗录 起行，安营在 利提玛 。
NUM|33|19|从 利提玛 起行，安营在 临门．帕烈 。
NUM|33|20|从 临门．帕烈 起行，安营在 立拿 。
NUM|33|21|从 立拿 起行，安营在 勒撒 。
NUM|33|22|从 勒撒 起行，安营在 基希拉他 。
NUM|33|23|从 基希拉他 起行，安营在 沙斐山 。
NUM|33|24|从 沙斐山 起行，安营在 哈拉大 。
NUM|33|25|从 哈拉大 起行，安营在 玛吉希录 。
NUM|33|26|从 玛吉希录 起行，安营在 他哈 。
NUM|33|27|从 他哈 起行，安营在 他拉 。
NUM|33|28|从 他拉 起行，安营在 密加 。
NUM|33|29|从 密加 起行，安营在 哈摩拿 。
NUM|33|30|从 哈摩拿 起行，安营在 摩西录 。
NUM|33|31|从 摩西录 起行，安营在 比尼．亚干 。
NUM|33|32|从 比尼．亚干 起行，安营在 曷．哈及甲 。
NUM|33|33|从 曷．哈及甲 起行，安营在 约巴他 。
NUM|33|34|从 约巴他 起行，安营在 阿博拿 。
NUM|33|35|从 阿博拿 起行，安营在 以旬．迦别 。
NUM|33|36|从 以旬．迦别 起行，安营在 寻 的旷野，就是 加低斯 。
NUM|33|37|从 加低斯 起行，安营在 以东 地边界的 何珥山 。
NUM|33|38|以色列 人出 埃及 地后四十年，五月初一， 亚伦 祭司遵照耶和华的指示，上 何珥山 ，死在那里。
NUM|33|39|亚伦 死在 何珥山 的时候一百二十三岁。
NUM|33|40|住在 迦南 地 尼革夫 的 迦南 人 亚拉得 王听说 以色列 人来了。
NUM|33|41|以色列 人从 何珥山 起行，安营在 撒摩拿 。
NUM|33|42|从 撒摩拿 起行，安营在 普嫩 。
NUM|33|43|从 普嫩 起行，安营在 阿伯 。
NUM|33|44|从 阿伯 起行，安营在 摩押 境内的 以耶．亚巴琳 。
NUM|33|45|从 以耶．亚巴琳 起行，安营在 底本．迦得 。
NUM|33|46|从 底本．迦得 起行，安营在 亚门．低比拉太音 。
NUM|33|47|从 亚门．低比拉太音 起行，安营在 尼波 前面的 亚巴琳山脉 。
NUM|33|48|从 亚巴琳山脉 起行，安营在 约旦河 边， 耶利哥 对面的 摩押 平原。
NUM|33|49|他们在 摩押 平原，沿着 约旦河 安营，从 伯．耶施末 直到 亚伯．什亭 。
NUM|33|50|耶和华在 约旦河 边， 耶利哥 对面的 摩押 平原吩咐 摩西 说：
NUM|33|51|“你要吩咐 以色列 人说：你们过 约旦河 进 迦南 地的时候，
NUM|33|52|要从你们面前赶出那地所有的居民，摧毁他们一切的石像和铸成的偶像，也要拆毁他们一切的丘坛。
NUM|33|53|你们要占领那地，住在那里，因我已把那地赐给你们为业。
NUM|33|54|你们要按照宗族抽签，承受土地：人多的要多给他们产业；人少的要少给他们产业。抽到何地给何人，那地就属于他。你们要按照父系的支派承受产业。
NUM|33|55|倘若你们不把那地的居民从你们面前赶出去，那留下的居民就必成为你们眼中的刺，肋下的荆棘，也必在你们所住的地上扰乱你们；
NUM|33|56|我想要怎样待他们，也必照样待你们。”
NUM|34|1|耶和华吩咐 摩西 说：
NUM|34|2|“你要吩咐 以色列 人，对他们说：你们到了 迦南 地，这就是归你们为业的地， 迦南 地和它四周的边界：
NUM|34|3|你们的南边是从 寻 的旷野起，沿着 以东 的边界；南边的地界从 盐海 东边开始，
NUM|34|4|绕过 亚克拉滨 斜坡的南边，经过 寻 ，直通到 加低斯．巴尼亚 的南边，又通到 哈萨．亚达 ，经过 押们 ，
NUM|34|5|从 押们 转向 埃及 溪谷，直通到海。
NUM|34|6|“你们西边的地界要以 大海 为边界；这就是你们西边的地界。
NUM|34|7|“你们北边的地界要从 大海 开始划界，直到 何珥山 ，
NUM|34|8|从 何珥山 划到 哈马口 ，直通到 西达达 ，
NUM|34|9|又通到 西斐仑 ，直达 哈萨．以难 。这就是你们北边的地界。
NUM|34|10|“东边的地界，你们要从 哈萨．以难 开始划界，直到 示番 ，
NUM|34|11|这地界要从 示番 下到 亚延 东边的 利比拉 ，这地界要下延到 基尼烈海 的东边，
NUM|34|12|这地界又下到 约旦河 ，直通到 盐海 。这就是你们的地和它四围的边界。”
NUM|34|13|摩西 吩咐 以色列 人说：“这就是耶和华吩咐抽签给九个半支派承受为业的地。
NUM|34|14|因为 吕便 子孙的支派按着父家、 迦得 子孙的支派按着父家，和 玛拿西 半个支派已经得到了他们的产业：
NUM|34|15|这两个半支派已经在 耶利哥 对面， 约旦河 东边，向日出的方向承受了产业。”
NUM|34|16|耶和华吩咐 摩西 说：
NUM|34|17|“这是为你们分地为业的人的名字： 以利亚撒 祭司和 嫩 的儿子 约书亚 。
NUM|34|18|你要从每个支派中选一个领袖来分配产业。
NUM|34|19|这些人的名字如下： 犹大 支派， 耶孚尼 的儿子 迦勒 。
NUM|34|20|西缅 子孙的支派， 亚米忽 的儿子 示母利 。
NUM|34|21|便雅悯 支派， 基斯伦 的儿子 以利达 。
NUM|34|22|但 子孙支派的领袖， 约利 的儿子 布基 。
NUM|34|23|约瑟 的子孙， 玛拿西 子孙支派的领袖： 以弗 的儿子 汉尼业 。
NUM|34|24|以法莲 子孙支派的领袖： 拾弗但 的儿子 基摩利 。
NUM|34|25|西布伦 子孙支派的领袖： 帕纳 的儿子 以利撒番 。
NUM|34|26|以萨迦 子孙支派的领袖： 阿散 的儿子 帕铁 。
NUM|34|27|亚设 子孙支派的领袖： 示罗米 的儿子 亚希忽 。
NUM|34|28|拿弗他利 子孙支派的领袖： 亚米忽 的儿子 比大黑 。”
NUM|34|29|这些就是耶和华所吩咐，在 迦南 地为 以色列 人分产业的人。
NUM|35|1|耶和华在 约旦河 边， 耶利哥 对面的 摩押 平原吩咐 摩西 说：
NUM|35|2|“你吩咐 以色列 人，要从所得为业的地中把一些城给 利未 人居住，也要把这些城四围的郊野给 利未 人。
NUM|35|3|这些城镇要归他们居住，郊外可以给他们牧放牛羊、牲畜和所有的动物。
NUM|35|4|你们给 利未 人城的郊外，要从城墙量起，四围往外量一千肘。
NUM|35|5|你们要往东量二千肘，往南量二千肘，往西量二千肘，往北量二千肘为边界，以城为中心；这城镇的郊外要归给他们。”
NUM|35|6|“你们给 利未 人的城镇中，要设立六座逃城，让误杀人的可以逃到那里。此外还要给他们四十二座城。
NUM|35|7|所以，给 利未 人的城一共有四十八座，连同城的郊外都给他们。
NUM|35|8|从 以色列 人所得的产业中给 利未 人的这些城镇，多的要多给，少的要少给；各支派要按照所承受为业之地的多少把城镇给 利未 人。”
NUM|35|9|耶和华吩咐 摩西 说：
NUM|35|10|“你要吩咐 以色列 人，对他们说：你们过了 约旦河 ，进入 迦南 地，
NUM|35|11|要指定几座城，作为你们的逃城，使误杀人的可以逃到那里。
NUM|35|12|这些城要作为逃避报仇者的城，使误杀人的不至于死，等他站在会众面前受审判。
NUM|35|13|“你们指定的城，是要作你们的六座逃城。
NUM|35|14|约旦河 东指定三座， 迦南 地也指定三座，作为逃城。
NUM|35|15|这六座城要给 以色列 人和他们中间的外人，以及寄居者，作为逃城，让误杀人的可以逃到那里。
NUM|35|16|“倘若人用铁器打死人，他是故意杀人的；故意杀人的必被处死。
NUM|35|17|若用手中可以致命的石头打死人，他是故意杀人的；故意杀人的必被处死。
NUM|35|18|若用手中可以致命的木器打死人，他是故意杀人的；故意杀人的必被处死。
NUM|35|19|报血仇者可以亲自杀死那故意杀人的；他一找到凶手，就可以杀死他。
NUM|35|20|人若因怨恨把人推倒，或埋伏等着丢东西砸人，以至于死，
NUM|35|21|或因仇恨用手打死人，打人的必被处死，他是故意杀人的；报血仇者一遇见凶手就可以杀死他。
NUM|35|22|“人若不是出于仇恨，把人推倒，或不是埋伏等着丢东西砸人，
NUM|35|23|或是在不注意的时候，用可以致命的石头扔在人身上，以至于死，彼此没有仇恨，也无意害对方，
NUM|35|24|会众就要照着这些典章，在杀人者和报血仇者中间审判。
NUM|35|25|会众要救这误杀人的脱离报血仇者的手，送他回到他曾逃入的逃城那里。他要住在城中，直到受圣膏的大祭司去世。
NUM|35|26|但误杀人的，无论什么时候，若离开了他所逃入的逃城边界，
NUM|35|27|报血仇者在逃城边界外遇见他，把凶手杀了，报血仇者就没有流人血之罪。
NUM|35|28|因为误杀人的应该住在逃城里，直到大祭司去世。大祭司去世以后，误杀人的才可以回到他所得为业之地。
NUM|35|29|在你们一切的住处，这些都要作为你们世世代代的律例典章。
NUM|35|30|“无论谁杀了人，必须凭几个证人的口，才可把那故意杀人的处死；只凭一个证人，不足以判人死。
NUM|35|31|那犯死罪的杀人犯，你们不可收赎价来代替他的命；他必须被处死。
NUM|35|32|那逃到逃城的人，你们不可向他收赎价，使他在大祭司未死以先回本地居住。
NUM|35|33|这样，你们就不会污秽所住之地，因为血能使地污秽；若有血流在地上，除非流那杀人者的血，否则那地就不得洁净。
NUM|35|34|你们不可玷污所住之地，就是我住在当中的地，因为我－耶和华住在 以色列 人中间。”
NUM|36|1|约瑟 子孙的宗族， 玛拿西 的孙子， 玛吉 的儿子 基列 ，他父系宗族的领袖来到 摩西 和作领袖的 以色列 众父系家长面前，说：
NUM|36|2|“耶和华曾吩咐我主抽签分地给 以色列 人为业，我主也遵照耶和华的吩咐，把我们兄弟 西罗非哈 的产业给他的女儿。
NUM|36|3|她们若嫁给 以色列 别个支派的人，必拿走我们祖宗所遗留的产业，加在她们丈夫支派的产业上。这样，我们抽签所得的产业就要减少了。
NUM|36|4|到了 以色列 人的禧年，她们的产业就必加在她们丈夫支派的产业上。这样，我们祖宗支派的产业就要减少了。”
NUM|36|5|摩西 照耶和华的指示吩咐 以色列 人说：“ 约瑟 子孙支派的人说得有理。
NUM|36|6|关于 西罗非哈 的女儿们，这是耶和华吩咐的话说：‘她们可以随意嫁人，只是必须嫁给同宗，她们父亲支派的人。
NUM|36|7|这样， 以色列 人的产业就不会从这支派转到另一个支派，因为 以色列 人要各自守住祖宗支派的产业。
NUM|36|8|凡在 以色列 支派中得了产业的女儿，必须嫁给同宗，她们父亲支派的人，好使 以色列 人各自承受他们祖宗的产业。
NUM|36|9|产业不可从一个支派转到另一个支派，因为 以色列 支派的人要各自守住自己的产业。’”
NUM|36|10|耶和华怎样吩咐 摩西 ， 西罗非哈 的女儿就照样做。
NUM|36|11|西罗非哈 的女儿 玛拉 、 得撒 、 曷拉 、 密迦 、 挪阿 都嫁给她们叔伯的儿子。
NUM|36|12|她们嫁给了 约瑟 儿子 玛拿西 子孙宗族的人；她们的产业保留在同宗，她们父亲的支派中。
NUM|36|13|这是耶和华在 约旦河 边， 耶利哥 对面的 摩押 平原，藉着 摩西 吩咐 以色列 人的命令和典章。
