1THESS|1|1|Павло й Силуан та Тимофій до Церкви Солунської в Бозі Отці й Господі Ісусі Христі: благодать вам і мир!
1THESS|1|2|Ми дякуємо Богові завжди за всіх вас, згадуючи вас у наших молитвах.
1THESS|1|3|Ми згадуємо безперестанку про ваше діло віри, і про працю любови, і про терпіння надії на Господа нашого Ісуса Христа, перед Богом і Отцем нашим,
1THESS|1|4|знаючи, Богом улюблені браття, про ваше обрання.
1THESS|1|5|Бо наша Євангелія не була для вас тільки у слові, а й у силі, і в Дусі Святім, і з великим упевненням, як знаєте ви, які ми були поміж вами для вас.
1THESS|1|6|І ви стали наслідувачі нам і Господеві, слово прийнявши в великому утискові з радістю Духа Святого,
1THESS|1|7|так що ви стали взірцем для всіх віруючих у Македонії та в Ахаї.
1THESS|1|8|Бо пронеслося Слово Господнє від вас не тільки в Македонії та в Ахаї, а й до кожного міста прийшла ваша віра в Бога, так що вам непотрібно казати чогось.
1THESS|1|9|Вони бо звіщають про нас, який був прихід наш до вас, і як ви навернулись до Бога від ідолів, щоб служити живому й правдивому Богові,
1THESS|1|10|і з неба очікувати Сина Його, що Його воскресив Він із мертвих, Ісуса, що визволює нас від майбутнього гніву.
1THESS|2|1|Самі бо ви знаєте, браття, прихід наш до вас, що не марний він був.
1THESS|2|2|Та хоч ми натерпілися перед тим, і дізнали зневаги в Филипах, як знаєте, проте ми відважилися в нашім Бозі звіщати вам Божу Євангелію з великою боротьбою.
1THESS|2|3|Бо покликання наше було не з обмани, ані з нечистости, ані від лукавства,
1THESS|2|4|але, як Бог визнав нас гідними, щоб нам доручити Євангелію, ми говоримо так, не людям догоджуючи, але Богові, що випробовує наші серця.
1THESS|2|5|Ми слова підлесливого не вживали ніколи, як знаєте, і не винні в зажерливості. Бог свідок тому!
1THESS|2|6|Не шукаємо ми слави в людей, ані в вас, ані в інших.
1THESS|2|7|Хоч могли ми потужними бути, як Христові апостоли, але ми серед вас були тихі, немов годувальниця та, яка доглядає дітей своїх.
1THESS|2|8|Так бувши ласкаві до вас, хотіли ми вам передати не тільки Божу Євангелію, але й душі свої, бо були ви улюблені нам.
1THESS|2|9|Бо ви пам'ятаєте, браття, наше струднення й утому: день і ніч ми робили, щоб жадного з вас не обтяжити, і проповідували вам Божу Євангелію.
1THESS|2|10|Ви свідки та Бог, як свято, і праведно, і бездоганно поводилися ми між вами, віруючими!
1THESS|2|11|Бож знаєте ви, як кожного з вас, немов батько дітей своїх власних,
1THESS|2|12|просили ми вас, і намовлювали та показували, щоб ви гідно поводилися перед Богом, що покликав вас у Своє Царство та в славу.
1THESS|2|13|Тому то й ми дякуємо Богові безперестанку, що, прийнявши почуте від нас Слово Боже, прийняли ви не як слово людське, але як правдиво то є Слово Боже, що й діє в вас, віруючих.
1THESS|2|14|Бо стали ви, браття, наслідувачами Церквам Божим, що в Юдеї в Христі Ісусі, бо те саме і ви були витерпіли від своїх земляків, як і ті від юдеїв,
1THESS|2|15|що вбили вони й Господа Ісуса, і пророків Його, і вигнали нас, і Богові не догоджають, і супротивні всім людям.
1THESS|2|16|Вони забороняють нам говорити поганам, щоб спаслися, щоб тим доповняти їм завжди провини свої. Але Божий гнів їх спіткає вкінці!
1THESS|2|17|А ми, браття, на короткий часок розлучившися з вами лицем, а не серцем, тим із більшим бажанням силкувались побачити ваше лице.
1THESS|2|18|Тим то до вас ми хотіли прийти, я, Павло, раз і двічі, але сатана перешкодив був нам.
1THESS|2|19|Бо хто нам надія, чи радість, чи вінок похвали? Хіба ж то й не ви перед Господом нашим Ісусом в Його приході?
1THESS|2|20|Бо ви наша слава та радість!
1THESS|3|1|Тому то, не стерпівши більше, ми схотіли зостатися в Атенах самі,
1THESS|3|2|і послали Тимофія, нашого брата й служителя Божого в Христовій Євангелії, щоб упевнити вас та потішити в вашій вірі,
1THESS|3|3|щоб ані один не хитався в цім горі. Самі бо ви знаєте, що на те нас призначено.
1THESS|3|4|Бо коли ми були в вас, то казали вам наперед, що маємо страждати, як і сталось, і знаєте ви.
1THESS|3|5|Тому й я, не стерпівши більше, послав довідатись про вашу віру, щоб часом спокусник вас не спокусив, і труд наш не стався б даремний.
1THESS|3|6|А тепер, як вернувся від вас Тимофій і приніс нам радісну звістку про віру та вашу любов, і що завжди ви маєте добру пам'ять про нас, і бажаєте бачити нас, як і ми вас,
1THESS|3|7|через те ми потішились, браття, за вас, у всякому горі та в нашій нужді, ради вашої віри.
1THESS|3|8|Бо тепер ми живемо, якщо в Господі ви стоїте!
1THESS|3|9|Яку бо подяку ми можемо Богові дати за вас, за всю радість, що нею ми тішимося ради вас перед нашим Богом?
1THESS|3|10|Ми вдень та вночі ревно молимося, щоб побачити ваше лице та доповнити те, чого не вистачає вашій вірі.
1THESS|3|11|Сам же Бог і Отець наш, і Господь наш Ісус нехай вирівняє нашу дорогу до вас!
1THESS|3|12|А в вас хай примножить Господь, і нехай збагатить вашу любов один до одного, і до всіх, як і наша є до вас!
1THESS|3|13|Нехай Він зміцнить серця ваші невинними в святості перед Богом і нашим Отцем, при приході Господа нашого Ісуса з усіма святими Його!
1THESS|4|1|А далі, браття, просимо вас та благаємо в Господі Ісусі, щоб, як прийняли ви від нас, як належить поводитись вам та догоджувати Богові, як ви й поводитеся, щоб у тому ще більше зростали!
1THESS|4|2|Бо ви знаєте, які вам накази дали ми Господом Ісусом.
1THESS|4|3|Бо це воля Божа, освячення ваше: щоб ви береглись від розпусти,
1THESS|4|4|щоб кожен із вас умів тримати начиння своє в святості й честі,
1THESS|4|5|а не в пристрасній похоті, як і погани, що Бога не знають.
1THESS|4|6|Щоб ніхто не кривдив і не визискував брата свого в якійбудь справі, бо месник Господь за все це, як і перше казали ми вам та засвідчили.
1THESS|4|7|Бо покликав нас Бог не на нечистість, але на освячення.
1THESS|4|8|Отож, хто оце відкидає, зневажає не людину, а Бога, що нам також дав Свого Духа Святого.
1THESS|4|9|А про братолюбство немає потреби писати до вас, бо самі ви від Бога навчені любити один одного,
1THESS|4|10|бо чините те всім братам у всій Македонії. Благаємо ж, браття, ми вас, щоб у цьому ще більш ви зростали,
1THESS|4|11|і пильно дбали жити спокійно, займатися своїми справами та заробляти своїми руками, як ми вам наказували,
1THESS|4|12|щоб ви перед чужими пристойно поводилися, і щоб ні від кого не залежали!
1THESS|4|13|Не хочу ж я, браття, щоб не відали ви про покійних, щоб ви не сумували, як і інші, що надії не мають.
1THESS|4|14|Коли бо ми віруємо, що Ісус був умер і воскрес, так і покійних через Ісуса приведе Бог із Ним.
1THESS|4|15|Бо це ми вам кажемо словом Господнім, що ми, хто живе, хто полишений до приходу Господнього, ми не попередимо покійних.
1THESS|4|16|Сам бо Господь із наказом, при голосі Архангола та при Божій сурмі зійде з неба, і перше воскреснуть умерлі в Христі,
1THESS|4|17|потім ми, що живемо й зостались, будемо схоплені разом із ними на хмарах на зустріч Господню на повітрі, і так завсіди будемо з Господом.
1THESS|4|18|Отож, потішайте один одного цими словами!
1THESS|5|1|А про часи та про пори, брати, не потрібно писати до вас,
1THESS|5|2|бо самі ви докладно те знаєте, що прийде день Господній так, як злодій вночі.
1THESS|5|3|Бо коли говоритимуть: Мир і безпечність, тоді несподівано прийде загибіль на них, як мука тієї, що носить в утробі, і вони не втечуть!
1THESS|5|4|А ви, браття, не в темряві, щоб той день захопив вас, як злодій.
1THESS|5|5|Бо ви всі сини світла й сини дня. Не належимо ми ночі, ні темряві.
1THESS|5|6|Тож не будемо спати, як інші, а пильнуймо та будьмо тверезі!
1THESS|5|7|Ті бо, що сплять сплять уночі, а ті, що напиваються вночі напиваються.
1THESS|5|8|А ми, що належимо дневі, будьмо тверезі, зодягнувшися в броню віри й любови, та в шолом надії спасіння,
1THESS|5|9|бо Бог нас не призначив на гнів, але щоб спасіння одержали Господом нашим Ісусом Христом,
1THESS|5|10|що помер був за нас, щоб, чи пильнуємо ми чи спимо, укупі з Ним ми жили.
1THESS|5|11|Утішайте тому один одного, і збудовуйте один одного, як і чините ви!
1THESS|5|12|Благаємо ж, браття, ми вас, шануйте тих, що працюють між вами, і в вас старшинують у Господі, і навчають вас вони,
1THESS|5|13|і в великій любові їх майте за їхню працю. Між собою заховуйте мир!
1THESS|5|14|Благаємо ж, браття, ми вас: напоумляйте непорядних, потішайте малодушних, підтримуйте слабих, усім довготерпіть!
1THESS|5|15|Глядіть, щоб ніхто нікому не віддавав злом за зло, але завжди дбайте про добро один для одного й для всіх!
1THESS|5|16|Завжди радійте!
1THESS|5|17|Безперестанку моліться!
1THESS|5|18|Подяку складайте за все, бо така Божа воля про вас у Христі Ісусі.
1THESS|5|19|Духа не вгашайте!
1THESS|5|20|Не гордуйте пророцтвами!
1THESS|5|21|Усе досліджуючи, тримайтеся доброго!
1THESS|5|22|Стережіться лихого в усякому вигляді!
1THESS|5|23|А Сам Бог миру нехай освятить вас цілком досконало, а непорушений дух ваш, і душа, і тіло нехай непорочно збережені будуть на прихід Господа нашого Ісуса Христа!
1THESS|5|24|Вірний Той, Хто вас кличе, Він і вчинить оте!
1THESS|5|25|Браття, моліться за нас!
1THESS|5|26|Привітайте всю браттю святим поцілунком!
1THESS|5|27|Заклинаю вас Господом, цього листа прочитати перед усіма братами!
1THESS|5|28|Благодать Господа нашого Ісуса Христа нехай буде з вами. Амінь!
