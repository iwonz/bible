2JOHN|1|1|The elder unto the elect lady and her children, whom I love in the truth; and not I only, but also all they that have known the truth;
2JOHN|1|2|For the truth's sake, which dwelleth in us, and shall be with us for ever.
2JOHN|1|3|Grace be with you, mercy, and peace, from God the Father, and from the Lord Jesus Christ, the Son of the Father, in truth and love.
2JOHN|1|4|I rejoiced greatly that I found of thy children walking in truth, as we have received a commandment from the Father.
2JOHN|1|5|And now I beseech thee, lady, not as though I wrote a new commandment unto thee, but that which we had from the beginning, that we love one another.
2JOHN|1|6|And this is love, that we walk after his commandments. This is the commandment, That, as ye have heard from the beginning, ye should walk in it.
2JOHN|1|7|For many deceivers are entered into the world, who confess not that Jesus Christ is come in the flesh. This is a deceiver and an antichrist.
2JOHN|1|8|Look to yourselves, that we lose not those things which we have wrought, but that we receive a full reward.
2JOHN|1|9|Whosoever transgresseth, and abideth not in the doctrine of Christ, hath not God. He that abideth in the doctrine of Christ, he hath both the Father and the Son.
2JOHN|1|10|If there come any unto you, and bring not this doctrine, receive him not into your house, neither bid him God speed:
2JOHN|1|11|For he that biddeth him God speed is partaker of his evil deeds.
2JOHN|1|12|Having many things to write unto you, I would not write with paper and ink: but I trust to come unto you, and speak face to face, that our joy may be full.
2JOHN|1|13|The children of thy elect sister greet thee. Amen.
