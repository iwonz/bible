ISA|1|1|Видіння 2377 Ісаї 3470, Амосового 531 сина 1121, яке він був бачив 2372 8804 про Юдею 3063 та про Єрусалим 3389 за днів 3117 Уззії 5818, Йотама 3147, Ахаза 271 та Єзекії 3169, Юдиних 3063 царів 4428.
ISA|1|2|Послухайте ви, небеса, і ти, земле, почуй, бо говорить Господь: Синів Собі виховав й викохав Я, а вони зняли бунт проти Мене!...
ISA|1|3|Віл знає свого власника, а осел ясла пана свого, а Ізраїль не знає Мене, не звертає уваги народ Мій на Мене...
ISA|1|4|О люду ти грішний, народе тяжкої провини, лиходійське насіння, сини-шкідники, ви покинули Господа, ви Святого Ізраїлевого понехтували, обернулись назад!
ISA|1|5|У що будете биті ще, коли неслухняними далі ви будете? Хвора ваша вся голова, і все серце боляще...
ISA|1|6|Від підошви ноги й аж до голови нема цілого місця на ньому: рани й ґудзі, та свіжі порази невичавлені, і не позав'язувані, і оливою не порозм'якшувані...
ISA|1|7|Земля ваша спустошена, огнем спалені ваші міста, поле ваше, на ваших очах поїдають чужинці його, з того всього пустиня, немов з руйнування чужинців!...
ISA|1|8|І позосталась Сіонська дочка, мов курінь в винограднику, мов шатро на ночліг в огірковому полі, як місто обложене...
ISA|1|9|Коли б був Господь Саваот не лишив нам останку малого, ми були б як Содом, до Гоморри ми стали б подібні...
ISA|1|10|Послухайте слова Господнього, содомські князі, почуйте Закон Бога нашого, народе гоморський,
ISA|1|11|нащо Мені многота ваших жертов? говорить Господь. Наситився Я цілопаленнями баранів і жиром ситих телят, а крови биків та овець і козлів не жадаю!
ISA|1|12|Як приходите ви, щоб явитися перед обличчям Моїм, хто жадає того з руки вашої, щоб топтали подвір'я Мої?
ISA|1|13|Не приносьте ви більше марнотного дару, ваше кадило огида для Мене воно; новомісяччя та ті суботи і скликання зборів, не можу знести Я марноти цієї!...
ISA|1|14|Новомісяччя ваші й усі ваші свята ненавидить душа Моя їх: вони стали Мені тягарем, Я змучений зносити їх...
ISA|1|15|Коли ж руки свої простягаєте, Я мружу від вас Свої очі! Навіть коли ви молитву примножуєте, Я не слухаю вас, ваші руки наповнені кров'ю...
ISA|1|16|Умийтесь, очистьте себе! Відкиньте зло ваших учинків із-перед очей Моїх, перестаньте чинити лихе!
ISA|1|17|Навчіться чинити добро, правосуддя жадайте, карайте грабіжника, дайте суд сироті, за вдову заступайтесь!
ISA|1|18|Прийдіть, і будемо правуватися, говорить Господь: коли ваші гріхи будуть як кармазин, стануть білі, мов сніг; якщо будуть червоні, немов багряниця, то стануть мов вовна вони!
ISA|1|19|Як захочете ви та послухаєтесь, то будете добра землі споживати.
ISA|1|20|А коли ви відмовитеся й неслухняними будете, меч пожере вас, бо уста Господні сказали оце!
ISA|1|21|Як стало розпусницею вірне місто: було повне воно правосуддя, справедливість у нім пробувала, тепер же розбійники!
ISA|1|22|Срібло твоє стало жужелицею, твоє питво водою розпущене...
ISA|1|23|Князі твої вперті і друзі злодіям вони, хабара вони люблять усі та женуться за дачкою, не судять вони сироти, удовина справа до них не доходить...
ISA|1|24|Тому то говорить Господь, Господь Саваот, Сильний Ізраїлів: О, буду Я тішитися над Своїми супротивниками, і помщусь на Своїх ворогах!
ISA|1|25|І на тебе Я руку Свою оберну, і твою жужелицю немов лугом витоплю, і все твоє оливо повідкидаю!
ISA|1|26|І верну твоїх суддів, як перше було, і твоїх радників, як напочатку. По цьому тебе будуть звати: місто справедливости, місто вірне!
ISA|1|27|Правосуддям Сіон буде викуплений, а той, хто навернеться в нім, справедливістю.
ISA|1|28|А знищення грішників та винуватців відбудеться разом, і ті, що покинули Господа, будуть понищені.
ISA|1|29|І будете ви посоромлені за ті дуби, що їх пожадали, і застидаєтеся за садки, які вибрали ви.
ISA|1|30|Бо станете ви, як той дуб, що листя всихає йому, і як сад, що не має води.
ISA|1|31|І станеться сильний кострицею, його ж діло за іскру, і вони обоє попаляться разом, і не буде нікого, хто б те погасив!
ISA|2|1|Слово, що його бачив Ісая, син Амосів, про Юдею та про Єрусалим:
ISA|2|2|І станеться на кінці днів, міцно поставлена буде гора дому Господнього на шпилі гір, і піднята буде вона понад згір'я, і полинуть до неї всі люди.
ISA|2|3|І підуть численні народи та й скажуть: Ходіть та зберімось на гору Господню, до дому Бога Якового, і доріг Своїх Він нас навчить, і ми підемо стежками Його! Бо вийде з Сіону Закон, і слово Господнє з Єрусалиму.
ISA|2|4|І Він буде судити між людьми, і буде численні народи розсуджувати. І мечі свої перекують вони на лемеші, а списи свої на серпи. Не підійме меча народ проти народу, і більше не будуть навчатись війни!
ISA|2|5|Доме Яковів, ідіть, і попростуємо в світлі Господньому!
ISA|2|6|Бо Ти був покинув народа Свого, дім Яковів, бо повні безладдя зо сходу вони, та ворожбитів, немов филистимляни, і накладають із дітьми чужинців.
ISA|2|7|І наповнився край його сріблом та золотом, і немає кінця його скарбам. І наповнився край його кіньми, і немає кінця колесницям його.
ISA|2|8|І наповнився край його ідолами, він кланяється ділу рук своїх, тому, що зробили були його пальці,
ISA|2|9|і поклонилась людина, і чоловік упокорився... А Ти їм не даруй!
ISA|2|10|Іди в скелю, і сховайся у порох від страху Господнього, і від пишноти Його величі!
ISA|2|11|Горді очі людини поникнуть, і буде обнижена людська високість, і буде високим Сам тільки Господь того дня!
ISA|2|12|Бо настане день Господа Саваота на все горде й високе, і на все висунене, і понижене буде воно,
ISA|2|13|і на всі кедри ливанські, високі та висунені, і на всілякі башанські дуби,
ISA|2|14|і на всі гори високі, і на всі згір'я піднесені,
ISA|2|15|і на всі башти високі, і на всі мури стрімкі,
ISA|2|16|і на всі кораблі із Таршішу, і на все, на що дивимося пожадливо!
ISA|2|17|І понизиться гордість людини, й обнижена буде високість людей, і буде високим Сам тільки Господь того дня,
ISA|2|18|а божища зовсім минуться!
ISA|2|19|І вони підуть до скельних печер та до пороху в ями від страху Господнього і від пишноти Його величі, коли прийде Він острах збудити на землі!
ISA|2|20|Покине людина того дня божків своїх срібних і божків своїх золотих, що собі наробила була, щоб вклонятись кротам і кажанам,
ISA|2|21|щоб піти у печери й розщілини скельні від страху Господнього і від слави величчя Його, коли прийде Він острах збудити на землі!
ISA|2|22|Відкинься ж собі від людини, що віддих у носі її, бо защо її поважати?
ISA|3|1|Бо Господь ось, Господь Саваот візьме з Єрусалиму й з Юдеї підпору й опору: усяку підпору від хліба, і всяку підпору води,
ISA|3|2|лицаря та вояка, суддю та пророка, і чарівника та старого,
ISA|3|3|п'ятдесятника та родовитого, і радника, і в мистецтві премудрого, і в закляттях умілого,
ISA|3|4|і за правителів дам юнаків, і дітваки запанують над ними!
ISA|3|5|І буде чавити народ один одного, і кожен свого ближнього! Повстане хлопчак на старого, а легковажений на поважаного...
ISA|3|6|Бо схопить брат брата свого в домі батька свого та й скаже: Ти маєш одежу, то будь нашим правителем, і під рукою твоєю хай буде руїна оця!
ISA|3|7|Того дня він підійме свій голос та й скаже: Не буду я рани обв'язувати вам, бо в домі моєму немає ні хліба, ні одягу, не настановляйте мене за правителя люду!
ISA|3|8|Бо рухнув Єрусалим, і впала Юдея, бо їхній язик та їхній чин проти Господа, щоб упертими бути очам Його слави...
ISA|3|9|Проти них свідчить вираз лиця їхнього, а гріх свій вони виявляють, немов той Содом, не перечать. Горе їхній душі, бо вчинили вони собі зло!
ISA|3|10|Скажіте про праведного: Буде добре йому, бо вони споживуть плід учинків своїх.
ISA|3|11|Та горе безбожному, зле, бо йому буде зроблений чин його рук!
ISA|3|12|Народ Мій, дітиська його утискають, а жінки мають гору над ним... Народе ти Мій, твої провідники вчинили блудячим тебе, і дорогу стежок твоїх сплутали!
ISA|3|13|Господь став на прю, і стоїть, щоб судити народи.
ISA|3|14|Господь іде на суд, щоб судитись з старшими народу Свого та з вождями його: Ви виноградника знищили, грабунок з убогого в ваших домах!
ISA|3|15|Що це сталося вам, що народ Мій ви гнобите та утискаєте вбогих? Так говорить Господь, Бог Саваот.
ISA|3|16|І промовив Господь: Зате, що дочки Сіонські загорділи, і ходять витягненошиї, і моргають очима, і все ходять дрібними крочками, і дзвонять спряжками на ногах своїх,
ISA|3|17|тому вчинить Господь тім'я Сіонських дочок паршивим, і їхній сором обнажить Господь!...
ISA|3|18|Того дня поскидає Господь окрасу спряжок на їхніх ногах, і чільця, і місяці,
ISA|3|19|сережки, нараменники, і серпанки,
ISA|3|20|і завої, і ланцюжки на ногах, і пояски, і пляшечки з пахощами, і чарівничі привіски,
ISA|3|21|персні, і сережки носові,
ISA|3|22|чудові убрання, і окриття, і намітки та торби,
ISA|3|23|дзеркала й льняні хитони та турбани, і прозорі покривала.
ISA|3|24|І станеться, замість бальзаму сморід буде, і замість пояса шнур, а замість мистецько укладених кучерів лисина, і замість хитона цінного верета з паском, а замість краси спаленина!
ISA|3|25|Попадають мужі твої від меча, а лицарство твоє на війні,
ISA|3|26|і будуть стогнати та плакати ворота її, і буде спустошена, й сяде на землю Сіонська дочка...
ISA|4|1|І того дня сім жінок схоплять мужа одного, говорячи: Ми будемо їсти свій хліб, і зодягатимем одіж свою, тільки йменням твоїм хай нас кличуть, забери ти наш сором!
ISA|4|2|Того дня буде парость Господня красою та славою, плід же земний величністю та пишнотою для врятованих із Ізраїля.
ISA|4|3|І буде зосталий в Сіоні й полишений в Єрусалимі, святим буде зватися він, кожен, хто жити записаний в Єрусалимі,
ISA|4|4|коли нечистоту Господь змиє з сіонських дочок, а кров Єрусалиму сполоще з-посеред його духом права та духом очищення.
ISA|4|5|І створить Господь над усяким житлом на Сіонській горі та над місцем зібрання удень хмару, вночі ж дим і блиск огню полум'яного, бо над всякою славою буде покрова...
ISA|4|6|І буде шатро удень тінню від спеки, і захистом та укриттям від негоди й дощу!
ISA|5|1|Заспіваю ж я вам про Свойого Улюбленого пісню любовну про Його виноградника! На плодючому версі гори виноградника мав був Мій Приятель.
ISA|5|2|І обкопав Він його, й від каміння очистив його, і виноградом добірним його засадив, і башту поставив посеред його, і витесав у ньому чавило, і чекав, що родитиме він виноград, та він уродив дикі ягоди!
ISA|5|3|Тепер же ти, єрусалимський мешканче та мужу юдейський, розсудіть но між Мною й Моїм виноградником:
ISA|5|4|що ще можна вчинити було для Мого виноградника, але Я не зробив того в ньому? Чому Я чекав, що родитиме він виноград, а він уродив дикі ягоди?
ISA|5|5|А тепер завідомлю Я вас, що зроблю для Свого виноградника: живопліт його викину, і він буде на знищення, горожу його розвалю, і він на потоптання буде,
ISA|5|6|зроблю Я загубу йому, він не буде обтинаний ані підсапуваний, і виросте терня й будяччя на ньому, а хмарам звелю, щоб дощу не давали на нього!
ISA|5|7|Бо виноградник Господа Саваота то Ізраїлів дім, а муж Юди коханий Його саджанець. Сподівавсь правосуддя, та ось кроволиття, сподівавсь справедливости Він, та ось зойк...
ISA|5|8|Горе тим, що долучують дома до дому, а поле до поля приточують, аж місця бракує для інших, так ніби самі сидите серед краю!
ISA|5|9|В мої уші сказав був Господь Саваот: Направду, багато домів попустошені будуть, великі та добрі, і не буде мешканця для них.
ISA|5|10|Бо десять загонів землі виноградника бата одного вродять, а насіння одного хомера породить ефу.
ISA|5|11|Горе тим, що встають рано вранці і женуть за напоєм п'янким, і тривають при нім аж до вечора, щоб вином розпалятись!
ISA|5|12|І сталася цитра та арфа, бубон та сопілка й вино за їхню гулянку, а на діло Господнє не дивляться, не вбачають Його чину рук.
ISA|5|13|Тому піде народ Мій на вигнання непередбачено, і вельможі його голодуватимуть, а натовп його висохне з прагнення...
ISA|5|14|Тому то розширив шеол пожадливість свою і безмірно розкрив свою пащу, і зійде до нього його пишнота, і його натовп, і гуркіт його, й ті, що тішаться в ньому.
ISA|5|15|І людина понижиться, і упокориться муж, а очі високих поникнуть,
ISA|5|16|а Господь Саваот возвеличиться в суді, і Бог Святий виявить святість Свою в справедливості!
ISA|5|17|І пастися будуть овечки, немов би на луці своїй, а зоставлене з ситих чужі поїдять.
ISA|5|18|Горе тим, що вину притягають до себе шнурами марноти, а гріх як мотуззям від воза,
ISA|5|19|та кажуть: Хай квапиться Він, хай принаглить Свій чин, щоб ми бачили, а постанова Святого Ізраїлевого хай наблизиться і нехай прийде і пізнаємо ми!
ISA|5|20|Горе тим, що зло називають добром, а добро злом, що ставлять темноту за світло, а світло за темряву, що ставлять гірке за солодке, а солодке за гірке!
ISA|5|21|Горе мудрим у власних очах та розумним перед собою самим!
ISA|5|22|Горе тим, що хоробрі винце попивати, і силачі на мішання п'янкого напою,
ISA|5|23|що несправедливого чинять в суді за хабар справедливим, а праведність праведного усувають від нього...
ISA|5|24|Тому, як огненний язик пожирає стерню, а від полум'я никне трава, отак спорохнявіє корінь у них, і рознесеться їхній цвіт, немов курява, бо від себе відкинули Закон Господа Саваота, і знехтували вони слово Святого Ізраїлевого!
ISA|5|25|Тому запалився гнів Господа на народ Його, і на нього Він витягнув руку Свою, та й уразив його: і захиталися гори, і сталось їхнього трупу, як сміття серед вулиць!... При цьому всьому не відвернувсь Його гнів, і витягнена ще рука Його!
ISA|5|26|І підійме прапора народу здалека, і засвище йому з кінця краю, і прийде він хутко та легко,
ISA|5|27|немає між ними утомленого та такого, який би спіткнувся! Не дримає ніхто і не спить, а пояс із стегон його не здіймається та не зривається шнур при взутті його.
ISA|5|28|Його стріли погострені, і всі луки його понатягувані. Копита у коней його немов кремінь вважаються, а колеса його немов вихор.
ISA|5|29|Його рик як левиці, і він заричить, немов ті левчуки, і він загарчить, і здобич ухопить, й її понесе, і ніхто не врятує!
ISA|5|30|І на нього ревітиме він того дня, як те море реве... І погляне на землю, а там густа темрява, і світло померкло у хмарах її...
ISA|6|1|Року смерти царя Озії бачив я Господа, що сидів на високому та піднесеному престолі, а кінці одежі Його переповнювали храм.
ISA|6|2|Серафими стояли зверху Його, по шість крил у кожного: двома закривав обличчя своє, і двома закривав ноги свої, а двома літав.
ISA|6|3|І кликав один до одного й говорив: Свят, свят, свят Господь Саваот, уся земля повна слави Його!
ISA|6|4|І захиталися чопи порогів від голосу того, хто кликав, а храм переповнився димом!
ISA|6|5|Тоді я сказав: Горе мені, бо я занапащений! Бо я чоловік нечистоустий, і сиджу посеред народу нечистоустого, а очі мої бачили Царя, Господа Саваота!
ISA|6|6|І прилетів до мене один з Серафимів, а в руці його вугіль розпалений, якого він узяв щипцями з-над жертівника.
ISA|6|7|І він доторкнувся до уст моїх та й сказав: Ось доторкнулося це твоїх уст, і відійшло беззаконня твоє, і гріх твій окуплений.
ISA|6|8|І почув я голос Господа, що говорив: Кого Я пошлю, і хто піде для Нас? А я відказав: Ось я, пошли Ти мене!
ISA|6|9|А Він проказав: Іди, і скажеш народові цьому: Ви будете чути постійно, та не зрозумієте, і будете бачити завжди, але не пізнаєте.
ISA|6|10|Учини затужавілим серце народу цього, і тяжкими зроби його уші, а очі йому позаклеюй, щоб не бачив очима своїми, й ушима своїми не чув, і щоб не зрозумів своїм серцем, і не навернувся, і не був уздоровлений він!
ISA|6|11|І сказав я: Аж доки, о Господи? А Він відказав: Аж доки міста спустіють без мешканця, і доми без людей, а земля спустошена буде зовсім...
ISA|6|12|І віддалить людину Господь, і буде велике опущення серед землі...
ISA|6|13|І коли позостанеться в ній ще десята частина, вона знову спустошена буде... Але мов з теребинту й мов з дубу, зостанеться в них пень по зрубі, насіння бо святости пень їхній!
ISA|7|1|І сталося за днів Ахаза, сина Йотама, Уззіїного сина, царя Юди, вийшов Рецін, цар сирійський, і Пеках, син Ремаліїн, цар Ізраїлів, до Єрусалиму на війну на нього, та не міг звоювати його.
ISA|7|2|І сповіщено Давидів дім, і сказано: Став табором Арам у землі Єфремовій. І захиталося серце його й серце народу його, як хитаються лісові дерева від вітру!
ISA|7|3|І сказав Господь до Ісаї: Вийди навпроти Ахаза, ти та твій син Шеар-Яшув, до кінця водоводу горішнього ставу, на биту дорогу Поля-Валюшників.
ISA|7|4|І скажеш до нього: Стережися й будь спокійний, не бійся, а серце твоє нехай не м'якне через два залишки тих димлячих головешок, від полум'я гніву Реціна й Арама та сина Ремаліїного,
ISA|7|5|за те, що Арам, Єфрем та син Ремаліїн радили проти тебе лихе, говорячи:
ISA|7|6|Ходім на Юдею та її налякаємо, і здобудемо для себе, і настановимо царем серед нього Тавеїлового сина.
ISA|7|7|Так сказав Господь Бог: Цього не станеться й не буде!
ISA|7|8|Бо голова Араму Дамаск, а голова Дамаску Рецін, та ще шістдесят і п'ять літ, і буде зламаний Єфрем, так що перестане бути народом!
ISA|7|9|А голова Єфрему Самарія, а голова Самарії син Ремаліїн. Якщо ви не повірите, то не встоїте.
ISA|7|10|І Господь далі говорив до Ахаза й казав:
ISA|7|11|Зажадай собі знака від Господа, Бога твого, і зійди глибоко до шеолу, або зійди високо догори!
ISA|7|12|А Ахаз відказав: Не пожадаю я, і не буду спокушувати Господа.
ISA|7|13|І він сказав: Послухайте, доме Давидів, чи мало вам трудити людей, що трудите також Бога мого?
ISA|7|14|Тому Господь Сам дасть вам знака: Ось Діва в утробі зачне, і Сина породить, і назвеш ім'я Йому: Еммануїл.
ISA|7|15|Масло та мед буде Він споживати, аж поки не пізнає того, як зло відкидати та добро вибирати.
ISA|7|16|Бо поки пізнає Та Дитина, як зло відкидати та добро вибирати, буде покинена та земля, що ти лякаєшся перед двома царями її.
ISA|7|17|Спровадить Господь на тебе, і на народ твій, і на дім батька твого дні, які не приходили від дня відступлення Єфрема від Юди, спровадить царя асирійського.
ISA|7|18|І станеться в день той, привабить Господь муху, що в кінці рік Єгипту, та бджолу, що в асирійському краї,
ISA|7|19|і вони прилетять, та усядуться всі по проваллях стрімких та по щілинах скельних, і в усіх терновиннях, та на луках усіх...
ISA|7|20|Дня того оголить Господь немов бритвою, найнятою по тім боці ріки, царем асирійським, голову та волосся ніг, забере також бороду.
ISA|7|21|І буде дня того, що хто прогодує корівку та дві штуки худоби дрібної,
ISA|7|22|то станеться, що від многоти молока, що надоїть, споживатиме масло, бо масло та мед буде їсти всякий, хто зостанеться серед землі.
ISA|7|23|І буде дня того: кожне місце, що в нім буде тисяча лоз винограду на тисячу срібла, стане терниною та будяком!
ISA|7|24|Зо стрілами й з луком він буде ходити туди, бо стане терниною та будяком уся земля...
ISA|7|25|А на всі гори, що заступом копано їх, ти не зійдеш туди, бо будеш боятись тернини й будяччя, і стануться місцем вони, куди волів посилатимуть, і топтатимуть вівці його...
ISA|8|1|І промовив до мене Господь: Візьми собі велику таблицю, і напиши на ній людським письмом: Квапиться здобич, скорий грабіж.
ISA|8|2|І взяв я за свідків собі свідків вірних, священика Урію та Захарія, Єверехіїного сина.
ISA|8|3|І зблизився я до пророчиці, і вона зачала, і породила сина. Господь же до мене промовив: Назви ім'я йому: Квапиться здобич, скорий грабіж.
ISA|8|4|Бо поки юнак той умітиме кликати Батьку мій, та: Мамо моя, понесеться багатство Дамаску та здобич Самарії перед обличчя царя асирійського.
ISA|8|5|І Господь ще далі говорив до мене й казав:
ISA|8|6|За те, що народ цей знехтував воду Сілоамську, яка тихо пливе, і має радість з Реціном і з сином Ремаліїним,
ISA|8|7|то тому ось Господь піднесе на них воду ріки, сильну й велику, царя асирійського та всю славу його. І підійметься вона понад усі свої річища, і піде понад усі береги свої.
ISA|8|8|І перейде по Юді вона, заллє та затопить, аж до шиї досягне, і розтягне вона свої крила на всю широчінь твого краю, о Еммануїле!
ISA|8|9|Озлобляйтесь народи, й збентежені будете, почуй, уся земле далека! Озбройтесь, і збентежені будете, озбройтесь, і збентежені будете!
ISA|8|10|Радьте раду і буде вона поруйнована, слово кажіть і не збудеться, бо з нами Бог!
ISA|8|11|Бо так говорив був до мене Господь у силі Своєї руки надо мною, й остерігав мене, щоб не ходити дорогою цього народу, і казав:
ISA|8|12|Не кажіть змова на все, на що каже змова цей народ, і не бійтесь того, чого він боїться, і не лякайтеся!
ISA|8|13|Господа Саваота Його свято шануйте, і Його вам боятись, Його вам лякатись!
ISA|8|14|І буде Він за святиню, і за камінь спотикання, і за скелю спокуси для двох домів Ізраїля, за сітку й за пастку для мешканця Єрусалиму.
ISA|8|15|І спіткнуться об них багатохто, і попадають, і будуть поламані, і заплутаються, і будуть схоплені.
ISA|8|16|Зв'яжи свідоцтво, запечатай Закона між Моїми учнями.
ISA|8|17|І я буду чекати Господа, що ховає лице Своє від Якового дому, і буду надіятись на Нього.
ISA|8|18|Ось я та ті діти, що дав мені Господь, вони на знаки та на чуда в Ізраїлі від Господа Саваота, що пробуває на горі Сіон.
ISA|8|19|А коли вам скажуть: Запитуйте духів померлих та чародіїв, що цвірінькають та муркають, то відповісте: Чи ж народ не звертається до свого Бога? За живих питатися мертвих?
ISA|8|20|До Закону й свідоцтва! Як вони не так кажуть, як це, то немає для них зорі ранньої!
ISA|8|21|І буде блукати утискуваний та голодний. І станеться, коли він зголодніє, то запіниться, і прокляне царя свого та Бога свого, і погляне догори,
ISA|8|22|і подивиться він на землю, аж ось тут горе та темнота, темрява утиску, і він буде пхнутий у темність...
ISA|9|1|(8-23) Бо не буде темноти для того, хто утискуваний. Перша пора злегковажила була край Завулонів та край Нефталимів, а остання прославить дорогу приморську, другий бік Йордану, округу поганів.
ISA|9|2|(9-1) Народ, який в темряві ходить, Світло велике побачить, і над тими, хто сидить у краю тіні смерти, Світло засяє над ними!
ISA|9|3|(9-2) Ти помножиш народ цей, Ти збільшиш йому радість. Вони перед лицем Твоїм будуть радіти, як радіють в жнива, як тішаться в час, коли ділять здобич!
ISA|9|4|(9-3) Бо зламав Ти ярмо тягару його, і кия з рамена його, жезло його пригнобителя, як за днів Мадіяма.
ISA|9|5|(9-4) Усякий бо чобіт військовий, що гупає гучно, та одежа, поплямлена кров'ю, стане все це пожежею, за їжу огню!
ISA|9|6|(9-5) Бо Дитя народилося нам, даний нам Син, і влада на раменах Його, і кликнуть ім'я Йому: Дивний Порадник, Бог сильний, Отець вічности, Князь миру.
ISA|9|7|(9-6) Без кінця буде множитися панування та мир на троні Давида й у царстві його, щоб поставити міцно його й щоб підперти його правосуддям та правдою відтепер й аж навіки, ревність Господа Саваота це зробить!
ISA|9|8|(9-7) Проти Якова слово послав був Господь, а впало воно на Ізраїля,
ISA|9|9|(9-8) і пізнає народ, увесь він, Єфрем та мешканець Самарії, що говорять з пихою й надутістю серця:
ISA|9|10|(9-9) Попадали цегли, а ми побудуємо з каменя тесаного, сікомори позрубувано, та замінимо їх кедрами!
ISA|9|11|(9-10) Та над ним Господь зміцнив противників Реціна, а його ворогів нацькував:
ISA|9|12|(9-11) Арама попереду, а филистимлян позаду, і пожерли Ізраїля цілою пащею... При цьому всьому не відвернувсь Його гнів, і витягнена ще рука Його!
ISA|9|13|(9-12) Та народ не звернувся до Того, Хто вразив його, і не шукали Господа Саваота...
ISA|9|14|(9-13) Тому то Господь відсік від Ізраїля голову й хвіст, пальму й очеретину за одного дня.
ISA|9|15|(9-14) Старий та поважаний це та голова, а пророк, що навчає неправди, це хвіст.
ISA|9|16|(9-15) І сталося, що поводатарі цього народу зробилися звідниками, і гинуть проваджені ними.
ISA|9|17|(9-16) Тому то його юнаками радіти не буде Господь, а до сиріт його й його вдів милосердя не матиме, бо кожен безбожний й злочинець, і злобне всі уста говорять. При цьому всьому не відвернувсь Його гнів, і витягнена ще рука Його!...
ISA|9|18|(9-17) Бо злоба горить, як огонь, пожирає тернину й будяччя, і палає по запустах лісу, і крутяться вверх стовпи диму...
ISA|9|19|(9-18) Від лютости Господа Саваота земля загориться, і стане народ, як пожива огню, і не пощадить жоден брата свого!...
ISA|9|20|(9-19) І різати буде праворуч, та буде голодний, і жертиме зліва, але не насититься, кожен жертиме тіло рамена свого:
ISA|9|21|(9-20) Манасія Єфрема, а Єфрем Манасію, разом обоє на Юду... При цьому всьому не відвернувсь Його гнів, і витягнена ще рука Його!...
ISA|10|1|Горе законодавцям несправедливим, та писарям, які пишуть на лихо,
ISA|10|2|щоб від правосуддя усунути бідних, і щоб відняти права від убогих народу Мого, щоб стали вдовиці здобичею їм, і пограбувати сиріт...
ISA|10|3|А що ви чинитимете в день навіщення, і наглої згуби, що прийде здалека, до кого втечете за поміччю, і де позоставите славу свою?
ISA|10|4|Нічого не лишиться тільки зігнутися між полоненими, і попадати між позабиваними... При цьому всьому не відвернувсь Його гнів, і витягнена ще рука Його!...
ISA|10|5|Біда асирійцеві, жезлові гніву Мого, а кий у руках його це пересердя Моє!
ISA|10|6|На люд нечестивий пошлю Я його, про народ Мого гніву йому накажу, щоб набрати здобичі й вчинити грабунок, і щоб потоптати його, як болото на вулицях.
ISA|10|7|Та не так він собі розуміє, а серце його не так мислить, бо в серці його щоб немало народів понищити та погубити!
ISA|10|8|Бо говорить: Хіба мої провідники разом усі не царі?
ISA|10|9|Чи ж Кално не такий, як Кархеміш? Чи ж Хамат не такий, як Арпад? Хіба ж не така Самарія, як Дамаск?
ISA|10|10|Тому що рука моя царства божків досягла, а в них більші боввани, як в Єрусалимі та в Самарії,
ISA|10|11|то хіба не зроблю я так само для Єрусалиму й бовванів його, як зробив я був для Самарії й божків її?
ISA|10|12|І станеться, як доконає ввесь чин Свій Господь на Сіонській горі та в Єрусалимі, то скаже: Навіщу я плоди гордовитости серця царя асирійського та пишноту чванливих очей його!
ISA|10|13|Бо він каже: Вчинив я це міццю своєї руки й своїм розумом, я бо розумний, і відміняю границі народів, а їхній маєток грабую, й як сильний, скидаю пануючих!
ISA|10|14|І досягла, мов кубло те, багатства народів рука моя, й як збирають покинені яйця, я всю землю зібрав, і ніхто не порушив крилом, і дзюбка не відкрив, і не зацвірінькав...
ISA|10|15|Чи буде сокира пишатися понад свого рубача? Чи понад свого пилувальника буде гордитися пилка? Ніби жезло повищує тих, хто його підіймає, ніби підносить кий того, хто не є дерево!
ISA|10|16|Зате Господь, Бог Саваот пошле сухорлявість на ситих його, і під його славою полум'я буде палати, немов би пожар!
ISA|10|17|І Світло Ізраїля стане огнем, а Святий його полум'ям, і запалить воно, й пожере його терня й будяччя його в один день!
ISA|10|18|І славу лісу його й його саду вигубить Він від душі й аж до тіла, і буде, що знидіє він, мов той хворий,
ISA|10|19|і буде останок дерев його лісу такий нечисленний, що й хлопець їх спише!
ISA|10|20|І станеться в день той, останок Ізраїля і врятовані дому Якова не будуть вже більш опиратись на того, хто б'є їх, й обіпруться у правді на Господа, Святого Ізраїлевого.
ISA|10|21|Рештки навернуться, рештки Якова, до Сильного Бога.
ISA|10|22|Бо коли б був народ твій, Ізраїль, як морський пісок, тільки рештки із нього навернуться! Загибіль призначена є, щоб виповнилась справедливість,
ISA|10|23|бо виконає Господь, Бог Саваот постановлену згубу посеред всієї землі.
ISA|10|24|Тому так промовляє Господь, Бог Саваот: Мій народе, мешканче Сіону, не бійсь асирійця! Він палицею тебе вдарить, і кия свого підійме на тебе, як колись на дорозі єгипетській.
ISA|10|25|Бо мало ще, трохи побуде, та й скінчиться лють, і звернеться гнів Мій на знищення їх!
ISA|10|26|І збудить на нього бича Господь Саваот, як уразив був Він Мадіяма при скелі Орев, і кий Його буде на морі, і його Він простягне, як колись на Єгипет!
ISA|10|27|І станеться в день той, з твого рамена тягар його здійметься, а з-над шиї твоєї ярмо його, і через ситість ярмо буде знищене!
ISA|10|28|Він прийде навпроти Айяту, перейде в Мігрон, свої речі складе до Міхмашу.
ISA|10|29|Перейдуть провалля, Гева ночліг нам, затремтіла Рама, утекла Саулова Гів'а.
ISA|10|30|Заголоси ти, о дочко Галліму, послухай, Лаїше, о бідний Анатоте!
ISA|10|31|Мадмена розбіглась, мешканці Гевіму втікають...
ISA|10|32|Ще сьогодні зостанеться він у Нові; своєю рукою грозить горі дочки Сіону, пагірку Єрусалиму.
ISA|10|33|Ось Господь, Бог Саваот відтинає галузки застрашальною силою, і найвищі поставою будуть постинані, а високі будуть понижені.
ISA|10|34|І буде обтята навколо залізом гущавина лісу, і Ліван упаде від Могутнього!
ISA|11|1|І вийде Пагінчик із пня Єссеєвого, і Галузка дасть плід із коріння його.
ISA|11|2|І спочине на Нім Дух Господній, дух мудрости й розуму, дух поради й лицарства, дух пізнання та страху Господнього.
ISA|11|3|Його уподобання в страху Господньому, і Він не на погляд очей своїх буде судити, і не на послух ушей Своїх буде рішати,
ISA|11|4|але буде судити убогих за правдою, і правосуддя чинитиме слушно сумирним землі. І вдарить Він землю жезлом Своїх уст, а віддихом губ Своїх смерть заподіє безбожному.
ISA|11|5|І станеться поясом клубів Його справедливість, вірність же поясом стегон Його!
ISA|11|6|І замешкає вовк із вівцею, і буде лежати пантера з козлям, і будуть разом телятко й левчук, та теля відгодоване, а дитина мала їх водитиме!
ISA|11|7|А корова й ведмідь будуть пастися разом, разом будуть лежати їхні діти, і лев буде їсти солому, немов та худоба!
ISA|11|8|І буде бавитися немовлятко над діркою гада, і відняте від перс дитинча простягне свою руку над нору гадюки,
ISA|11|9|не вчинять лихого та шкоди не зроблять на всій святій Моїй горі, бо земля буде повна пізнання Господнього так, як море вода покриває!
ISA|11|10|І станеться в день той: до Кореня Єссеєвого, що стане прапором народам, погани звертатися будуть до Нього, і буде славою місце спочинку Його!
ISA|11|11|І станеться в день той, і знову подруге простягне Господь Свою руку, щоб набути останок народу Свого, що полишиться з Ашшуру й з Єгипту, і з Патросу та з Етіопії, і з Еламу й з Шін'ару, і з Хамату, та з морських островів.
ISA|11|12|І поганам підійме Він прапора, і згромадить вигнанців Ізраїля, і розпорошення Юди збере з чотирьох країв світу!
ISA|11|13|І спиниться заздрість Єфрема, і витяті будуть супротивники Юди, не буде вже заздрити Юді Єфрем, а Юда не буде гнобити Єфрема.
ISA|11|14|І вони полетять на плече филистимлян до моря, пограбують гуртом синів сходу, на Едома й Моава вони накладуть свою руку, і діти Аммона їх слухати будуть.
ISA|11|15|І вчинить закляттям Господь затоку моря Єгипетського, і руку Свою простягне на ріку в сильнім вітрі Своїм, і на сім потоків розділить її, й буде можна її у взутті переходити.
ISA|11|16|І буде широка дорога для решти народу Його, що з Ашшуру зостанеться, як була для Ізраїля в день, коли він виходив із краю єгипетського.
ISA|12|1|І ти скажеш дня того: Хвалю Тебе, Господи, бо Ти гнівавсь на мене, та гнів Твій вщухає, й мене Ти порадуєш,
ISA|12|2|оце, Бог спасіння моє! Безпечний я, і не боюсь, бо Господь, Господь сила моя та мій спів, і спасінням для мене Він став!
ISA|12|3|І ви в радості будете черпати воду з спасенних джерел!
ISA|12|4|І скажете ви того дня: Дякуйте Господу, кличте Імення Його, сповістіть між народів про вчинки Його, пригадайте, що Ймення Його превеличне!
ISA|12|5|Співайте для Господа, Він бо величне вчинив, і хай це буде знане по цілій землі!
ISA|12|6|Радій та співай, ти мешканко Сіону, бо серед тебе Великий, Святий Ізраїлів!
ISA|13|1|Пророцтво про Вавилон, що бачив Ісая, син Амосів.
ISA|13|2|Підійміте прапора на лисую гору, кличте їх голосніш, помахайте рукою, щоб ішли у ворота!
ISA|13|3|Я звелів був Своїм посвяченим, теж покликав лицарство Своє на Мій гнів, що зухвало радіють.
ISA|13|4|Чути гамір у горах, як народу численного, чути гомін згромаджених тут царств народів: це переглядає Господь Саваот бойове Своє військо!
ISA|13|5|Приходять з далекого краю, із кінців небес, Господь і знаряддя гніву Його, щоб усю землю понищити!
ISA|13|6|Голосіть, бо близький день Господній, він від Всемогутнього прийде, немов зруйнування...
ISA|13|7|Тому то ослабнуть всі руки, і кожне серце людини зневіриться.
ISA|13|8|І вони налякаються, болі та муки їх схоплять, немов породілля та, будуть тремтіти... Остовпіють один перед одним, полум'яні обличчя то їхні обличчя...
ISA|13|9|Оце день Господній приходить, суворий, і лютість, і полум'я гніву, щоб землю зробити спустошенням, а грішних її повигублювати з неї!
ISA|13|10|Бо зорі небесні та їхні сузір'я не дадуть свого світла, сонце затьмиться при сході своєму, а місяць не буде вже сяяти світлом своїм...
ISA|13|11|І Я покараю всесвіт за зло, а безбожних за їхню провину, бундючність злочинця спиню, а гордість насильників знижу!
ISA|13|12|Я зроблю людину дорожчою від щирого золота, і смертну людину від офірського золота.
ISA|13|13|Тому небеса захитаю, і рухнеться земля з свого місця від лютости Господа Саваота, у День, як палатиме гнів Його...
ISA|13|14|І буде народ, як та сарна сполошена чи як отара, якої зібрати немає кому... До народу свого кожен звернеться, і кожен до краю свого втікатиме.
ISA|13|15|Кожен знайдений буде заколеним, і кожен узятий впаде від меча...
ISA|13|16|А їхні діти на їхніх очах порозбивані будуть, їхні доми пограбовані будуть, а їхніх жінок побезчестять!
ISA|13|17|Оце Я збуджу на них мідян, що срібла не лічать, а золото не чують бажання до нього,
ISA|13|18|і будуть вбивати юнаків їхні луки, і над плодом утроби вони милосердя не матимуть, їхнє око над дітьми не матиме милости...
ISA|13|19|І стане тоді Вавилон, краса царств, пишнота халдейської гордости, таким, як Бог зруйнував був Содом та Гоморру!
ISA|13|20|Не буде назавжди заселений він, нізамешкалий з роду в рід, і араб там не стане наметом, і там пастухи не спочинуть з своєю отарою...
ISA|13|21|Але будуть барложити там звірі пустині, і будуть доми їхні совами повні, і там пробуватимуть струсі, і волохаті демони там танцюватимуть...
ISA|13|22|І завиють шакали в порожніх хоромах його, а гієни в веселих палацах! І близьке вже наступлення часу його, і не забаряться ці його дні!
ISA|14|1|Бо Господь змилосердиться над Яковом, і вибере знову Ізраїля, і на їхній землі їх поселить. І чужинець долучений буде до них, і приєднані будуть до дому Якового.
ISA|14|2|І народи їх візьмуть, і їх попровадять до їхнього місця, а Ізраїлів дім на Господній землі за рабів та за невільниць їх прийме собі на спадщину. І візьмуть вони до неволі тих, хто їх поневолив, і вони над своїми гнобителями запанують!
ISA|14|3|І буде в той день, як Господь дасть тобі відпочинок із терпіння твого та з неспокою твого, та з праці тяжкої, яку ти був мусів робити,
ISA|14|4|то ти заспіваєш оцю пісню глумливу про царя Вавилону та й скажеш: Як гнобитель минувся, минулося гноблення!
ISA|14|5|Господь зламав кия безбожних і жезла пануючих,
ISA|14|6|що народи постійним ударом у лютості бив, що в гніві гнобив був людей переслідуванням безупинним.
ISA|14|7|Спочила була, заспокоїлася вся земля, і виспівує голосно.
ISA|14|8|Кипариси та кедри ливанські тобою втішаються й кажуть: Відколи ти ліг, не приходить на нас дроворуб!
ISA|14|9|Заворушивсь тобою іздолу шеол назустріч твоєму приходу; померлих тобі побудив, усіх проводирів на землі, і підняв з їхніх тронів всіх людських царів.
ISA|14|10|Вони всі зачнуть говорити та й скажуть тобі: І ти ослабів, як і ми, став подібний до нас!
ISA|14|11|Зіпхнута в шеол твоя гордість та гра твоїх арф; вистелено під тобою червою, і червяк накриває тебе...
ISA|14|12|Як спав ти з небес, о сину зірниці досвітньої, ясная зоре, ти розбився об землю, погромнику людів!
ISA|14|13|Ти ж сказав був у серці своєму: Зійду я на небо, повище зір Божих поставлю престола свого, і сяду я на горі збору богів, на кінцях північних,
ISA|14|14|підіймуся понад гори хмар, уподібнюсь Всевишньому!
ISA|14|15|Та скинений ти до шеолу, до найглибшого гробу!
ISA|14|16|Ті, що на тебе дивитися будуть, приглядатися будуть до тебе, звернути увагу на тебе: Чи то той чоловік, що змушував землю тремтіти, що зневолював царства труситись,
ISA|14|17|що він обертав у пустиню вселенну, а міста її бурив, що в'язнів своїх не пускав він додому?
ISA|14|18|Усі царі людів, вони всі у славі лягли, кожен у своїй усипальні,
ISA|14|19|ти ж від гробу свого відкинений геть, мов галузка бридка, оточений вбитими та мечем перешитими, що до гробу між камінь спускаються, як потоптаний труп...
ISA|14|20|Ти не будеш поєднаний з ними у гробі, бо землю свою зруйнував, свій народ повбивав... Насіння злочинців повік не згадається!
ISA|14|21|Його дітям зготуйте різню за вину їхніх батьків, щоб вони не повстали, і землі не вспадкували, і не наповнили світу містами.
ISA|14|22|І на них Я повстану, говорить Господь Саваот, і витну ім'я Вавилону й останок його, і нащадка й онука, говорить Господь!
ISA|14|23|І вчиню Я його їжакові оселею та водним багном, і мітлою вигублення позамітаю його, говорить Господь Саваот!
ISA|14|24|Присягав був Господь Саваот та казав: Поправді, як мислив собі Я, так станеться, й як Я був врадив те сповниться,
ISA|14|25|щоб стовкти асирійця в країні Моїй, і на горах Моїх розтопчу Я його! І ярмо його здійметься з них, і тягар його скинеться з їхніх рамен!
ISA|14|26|Це та рада, яка про всю землю ураджена, і це та рука, що простягнена на всі народи.
ISA|14|27|Бо врадив Господь Саваот, і хто Його раду відмінить? А рука Його витягнена, й хто відверне її?
ISA|14|28|У році смерти царя Ахаза було таке пророцтво:
ISA|14|29|Не тішся, уся филистимськая земле, що зламане жезло, яке тебе вдарило, бо з гадючого кореня виповзе люта змія, і огнистий летючий дракон буде плодом її!
ISA|14|30|І пастися будуть перворідні бідних, і вбогі безпечно лежатимуть, а твій корень Я голодом виморю, і рештки твої він доб'є!
ISA|14|31|Плач же, брамо, ти ж місто, кричи, розпливлася ти, вся филистимськая земле, бо приходить із півночі дим, і не буде нікого, хто відстав би з його вояків!
ISA|14|32|І що відповісться народнім послам? Що Сіона Господь заложив, і сховаються в ньому убогі з народу Його!
ISA|15|1|Пророцтво про Моава. Справді вночі Ар-Моав пограбований був та понищений, справді вночі Кір-Моав пограбований був та понищений.
ISA|15|2|Він пішов до святині, а Дивон на верхів'я, щоб плакати; на Нево й на Медеву голосить Моав. На всіх головах його лисина, обстрижена кожна його борода,
ISA|15|3|на всіх його вулицях підперезались веретою, на дахах його та на площах його всі голосять, з плачу розпливаються...
ISA|15|4|І кричали Ешбон та Ел'але, аж до Ягацу був чутий їхній голос, тому то голосять вояки Моава, і душа його в ньому тремтить.
ISA|15|5|Моє серце кричить про Моава, втікачі його аж до Цоару, до Еглат-Шелішійї, бо з плачем ходять збіччям Лухіту, бо на Хоронаїмській дорозі встає крик загибелі,
ISA|15|6|бо води Німріму спустошенням будуть, бо посохла трава, мурава позникала, немає нічого зеленого...
ISA|15|7|Тому то набутий останок і маєток вони віднесуть за потік степовий.
ISA|15|8|Бо країну Моава той крик оточив, по Еглаїм його голосіння, і по Беер-Елім голосіння його.
ISA|15|9|Бо наповнилась кров'ю димонська вода, бо Я покладу на Димон додаткове: лева для втікачів із Моава, і на останок землі.
ISA|16|1|Овечки пошліть власникові землі, із Сели на пустиню, на гору Сіонської дочки.
ISA|16|2|І станеться, мов те сполошене птаство, з кубла повигонене, будуть дочки Моавські при бродах Арнону:
ISA|16|3|Подай раду, зроби присуд, учини нічну тінь свою повного полудня, сховай вигнаних, біженця не видавай...
ISA|16|4|Нехай мешкають в тебе вигнанці Моаву, стань їм захистом перед грабіжником, бо не стало насильника, скінчився грабунок, загинув топтач із землі...
ISA|16|5|І буде утверджений милістю трон, і сяде на ньому у правді в наметі Давида суддя, що дбатиме за правосуддя та буде в справедливості вправний.
ISA|16|6|Ми чули про гордість Моава, що гордий він дуже, про сваволю його й його гордість, про лютість його, про неслушні його нісенітниці...
ISA|16|7|Буде тому голосити Моав над Моавом, увесь голосити він буде! За паляницями з грон Кір-Харесету плакати будуть насправді побиті,
ISA|16|8|бо посохли хешбонські поля, і виноградник Сівми; володарі народів понищили грозна добірні, які до Язеру сягали й зникали в пустині; галузки ж його розтягалися, і море вони перейшли.
ISA|16|9|Тому то язерським плачем буду плакати за виноградину Сівми. Сльозою своєю тебе орошу, о Хешбоне й Ел'але, бо крик бою напав на твій збір та на жниво твоє.
ISA|16|10|І буде забрана радість та втіха із саду, а по виноградниках пісні не буде й не здійметься окрик. Вина по чавилах не буде топтати чавильник, окрик радости Я припинив!
ISA|16|11|Тому то в жалобі звучать про Моав мої нутрощі, мов би та арфа, а нутро моє про Кір-Херес.
ISA|16|12|І буде, як виявиться, що змучивсь на взгір'ї Моав, і ввійде молитись у святиню свою, та він не осягне нічого.
ISA|16|13|Оце слово, яке говорив був віддавна Господь про Моава.
ISA|16|14|А тепер Господь каже, говорячи: За три роки, однакові з літами наймита, буде зневажена слава Моава з усім велелюддям його, а позосталість мала та дрібна, невелика!
ISA|17|1|Пророцтво про Дамаск. Ось Дамаск вилучається з міст, і стається, як купа руїн.
ISA|17|2|Покинені будуть міста Ароеру, для черід вони будуть, і ті будуть лежати, і не буде кому їх сполошити...
ISA|17|3|Заникне твердиня з Єфрема, і царство з Дамаску, і решта Араму будуть, як слава синів Ізраїля, говорить Господь Саваот!
ISA|17|4|І станеться в день той, слава Якова знидіє, і вихудне товщ його тіла.
ISA|17|5|І буде, немов би жнець збирає збіжжя, а рамено його жне колосся; і буде, немов би збирають колосся в долині Рефаїм.
ISA|17|6|І на ньому зостануться залишки з плодів, як при оббиванні оливки: дві-три ягідки на верховітті, чотири-п'ять на галузках плідної деревини, говорить Господь, Бог Ізраїлів.
ISA|17|7|Того дня зверне людина зір до свого Творця, а очі її на Святого Ізраїлевого дивитися будуть.
ISA|17|8|І не буде звертатись людина до жертівників, чину рук своїх, і не буде дивитись на те, що зробили були її пальці, ні на ашери, ані на стовпи на честь сонця.
ISA|17|9|Того дня її сильні міста будуть, мов ті опустілі місця лісу та верхів'я гір, що їх позоставлено перед синами Ізраїля, і руїною станеться те.
ISA|17|10|Бо забула ти, дочко Ізраїля, Бога спасіння свого, і не пам'ятала про Скелю сили своєї. Тому то садиш розсадника приємного, і пересаджуєш туди чужу виноградину.
ISA|17|11|Того дня, як садила, ти обгородила його, і про посів свій подбала, щоб рано зацвіло. Але жниво минулося в день слабости невигойного болю!...
ISA|17|12|Біда, рев численних народів, гуркочуть, як гуркіт морів, і галас племен, вони галасують, як гуркіт міцної води.
ISA|17|13|Галасують племена, як гуркіт міцної води, та Він їм погрозить, і кожен далеко втече, і буде гнаний, немов та полова на горах за вітром, і мов перед вихром перекотиполе...
ISA|17|14|Як вечір насуне то й жах ось, поки ранок настане не буде його. Це талан наших грабівників, і це доля дерилюдів наших!...
ISA|18|1|Горе тобі, дзвінкокрилий ти краю, що з другого боку річок етіопських,
ISA|18|2|що морем послів посилаєш на човнах папірусових по поверхні води! Ідіть, скороходні посли, до народу високого й блискучезбройного, до народу страшного віддавна й аж досі, до люду пресильного, що топче усе, що річки його землю поперетинали.
ISA|18|3|Усі мешканці всесвіту, що на землі пробуваєте, дивіться, коли піднесеться прапор на горах, слухайте, чи не затрублять у ріг.
ISA|18|4|Бо Господь так промовив до мене: Я буду спокійний, і буду дивитися з місця Свого пробування, як тепло те при світлі ясному, як та хмара роси в спеку жнив!
ISA|18|5|Бо перед жнивами, як скінчиться цвіт, недозріле ж усе стане зрілими грознами, то Він зріже серпами галуззя м'які, а галузки, що стеляться, повідкидає, повідрубує Він.
ISA|18|6|Будуть вони позоставлені разом для хижого птаха гірського й звірини земної, і літо над ним проведе хижий птах, і вся земна звірина над ним перезимує.
ISA|18|7|Того часу принесений буде дарунок для Господа Саваота від народу високого й блискучезбройного, і від народу страшного віддавна й аж досі, від люду пресильного, що топче усе, що річки його землю поперетинали, до місця Ймення Господа Саваота на Сіонській горі.
ISA|19|1|Пророцтво про Єгипет. Ось на хмарі легенькій несеться Господь і прибуде в Єгипет, і затремтять перед лицем Його боввани Єгипту, і серце Єгипту розтане посеред нього.
ISA|19|2|І підбурю єгиптянина на єгиптянина, і будуть точити війну кожен з братом своїм, і кожен із ближнім своїм, місто з містом, а царство із царством.
ISA|19|3|І Єгипет на дусі поникне в своєму нутрі, а раду його Я поплутаю, і вони будуть питати бовванів своїх, і заклиначів духів та духів померлих і своїх ворожбитів.
ISA|19|4|І віддам Я Єгипет у руку жорстокого пана, і цар лютий над ним запанує, говорить Господь, Господь Саваот!
ISA|19|5|І зникне із Моря вода, і висохне Річка, та й стане суха.
ISA|19|6|І засмердяться річки та нужденними стануть, і повисихають притоки Єгипту, пов'яне комиш та очерет.
ISA|19|7|Луги над рікою, над берегом річки, і все, що при річці посіяне, повисихає, розвіється все, і не буде його.
ISA|19|8|І заплачуть рибалки, і будуть ридати всі ті, що гачка закидають до річки, а ті, що розтягують невід на воду, стратять надію.
ISA|19|9|А ті, що працюють при чесанім льоні та тчуть полотно, засоромляться.
ISA|19|10|І будуть основи Єгипту розбиті, всі ж працюючі за плату на дусі впадуть.
ISA|19|11|Дійсно, вельможі Цоану безумні, і нерозумною стала рада мудрих фараонових радників. І як фараонові скажете: Я син мудреців, я син давніх царів?
ISA|19|12|Де ж вони, де твої мудреці? І хай розкажуть тобі й хай пізнають, що порадив Господь Саваот на Єгипет.
ISA|19|13|Стали немудрі вельможі Цоану, вельможі Мемфісу обманені, учинили блудячим Єгипет головніші з племен його.
ISA|19|14|Господь влив у нього дух одуру, і вони вчинили блудячим Єгипет в усякому чині його, як блудить п'яниця в блювоті своїй...
ISA|19|15|І Єгипет не матиме діла, що вміли б вчинити його голова або хвіст, пальмова галузка чи очеретина.
ISA|19|16|Того дня стане Єгипет, немов ті жінки, і тремтітиме, і буде лякатись помаху руки Господа Саваота, що Він нею над ним помахає.
ISA|19|17|І стане юдейська земля для Єгипту за пострах: кожен, кому пригадають про неї, злякається перед задумом Господа Саваота, якого повзяв Він на нього.
ISA|19|18|Того дня буде п'ять міст в єгипетськім краї, що говоритимуть ханаанською мовою й присягатимуть Господом Саваотом. Одне буде зватися Ір-Гахерес.
ISA|19|19|Того дня серед краю єгипетського буде жертівник Господу, і стовп при границі його Господеві.
ISA|19|20|І він буде в єгипетськім краї ознакою й свідком для Господа Саваота, коли будуть взивати до Господа перед гнобителями, то пошле їм спасителя та оборонця, який їх спасе.
ISA|19|21|І стане знаний Господь для Єгипту, і того дня познають єгиптяни Господа, і будуть служити жертвою й жертвою хлібною, і присягнуть обітницю Господеві, і виповнять.
ISA|19|22|І вразить єгиптян Господь, буде бити їх та лікувати, і до Господа звернуться, і Він дасться їм ублагати Себе, і їх вилікує.
ISA|19|23|Того дня буде бита дорога з Єгипту в Асирію, і прийдуть асирійці до єгиптян, а єгиптяни до асирійців, і будуть служити єгиптяни з асирійцями Господеві.
ISA|19|24|Того дня буде Ізраїль третім краєм побіч Єгипту й Асирії, благословенням серед землі,
ISA|19|25|бо Господь Саваот його поблагословив та й сказав: Благословенний народ мій Єгипет, і Ашшур, чин Моїх рук, та Ізраїль, спадщина Моя!
ISA|20|1|Того року, коли Тартан прийшов до Ашдоду, як його послав був Сарґон, цар асирійський, і він воював був з Ашдодом і здобув його,
ISA|20|2|того часу казав був Господь через Ісаю, Амосового сина, говорячи: Іди, і розв'яжеш верету з-над стегон своїх, і здіймеш взуття зо своєї ноги! І він зробив так, ходив нагий та босий.
ISA|20|3|І Господь говорив: Як ходив Мій раб Ісая нагий та босий три роки, це ознака та чудо про Єгипет та про Етіопію,
ISA|20|4|так поведе цар асирійський полонених Єгипту й вигнанців Етіопії, юнаків та старих, нагих та босих, навіть з озадком відкритим. Сором Єгипту!
ISA|20|5|І будуть збентежені та засоромлені за Етіопію, куди звернений зір їхній, та за Єгипет, їхню пишноту.
ISA|20|6|І скаже того дня мешканець того побережжя: Оце таке місце, куди звернений зір наш, куди ми втікали за поміччю, щоб урятуватися перед асирійським царем. І як ми втечемо?
ISA|21|1|Пророцтво про пустиню надморську. Як носяться бурі на півдні, так ворог іде із пустині, із краю страшного.
ISA|21|2|Видіння грізне мені явлене: Грабує грабіжник, пустошник пустошить. Прийди, о Еламе, Мадай обложи, усяким зідханням зробив Я кінець.
ISA|21|3|Тому то наповнилися мої стегна тремтінням, і болі схопили мене, немов породільні ті болі. Я скривився від того, що чув, я від баченого перестрашивсь.
ISA|21|4|Забилося серце моє, тремтіння напало мене несподівано; вечір розкоші моєї змінився мені на страхіття.
ISA|21|5|Поставлений стіл, килимами накрито, їсться та п'ється. Уставайте, правителі, щити намастіть!
ISA|21|6|Бо до мене сказав Господь так: Іди, вартового постав, що побачить, нехай донесе.
ISA|21|7|І коли він похода побачив, по парі їздців, поїзд ослів, поїзд верблюдів, і прислухується він з увагою, із увагою пильною.
ISA|21|8|І він крикнув, як лев: Я завжди стою вдень на варті, о Господи, і стою на сторожі своїй усі ночі!
ISA|21|9|Аж ось іще похід мужів, по двоє їздців. І він відповів та сказав: Упав, упав Вавилон, а всі статуї богів його порозбивані об землю!
ISA|21|10|О мій помолочений ти, сину току мого! Я звістив вам, що чув був від Господа Саваота, Бога Ізраїлевого.
ISA|21|11|Пророцтво про Думу. До мене кричить із Сеїру: Стороже, яка пора ночі? Стороже, яка пора ночі?
ISA|21|12|А сторож сказав: Настав ранок, а все ж іще ніч. Якщо ви питатимете, то питайте та знову прийдіть!
ISA|21|13|Пророцтво про Арабію. У лісі в степу ночувати, ви будете каравани деданів.
ISA|21|14|Мешканці Теманського краю, винесіть воду назустріч для спрагненого, втікача зустрічайте із хлібом!
ISA|21|15|Бо втекли вони перед мечами, перед голим мечем, і перед натягненим луком, і перед тяготою війни.
ISA|21|16|Бо до мене Господь сказав так: Ще за рік, як рік наймита, і вся слава Кедару покінчиться.
ISA|21|17|А понадто полишиться невелике число лучників з лицарів кедарських синів, бо Господь, Бог Ізраїлів, це говорив.
ISA|22|1|Пророцтво про долину Видіння. Що це сталось тобі, що ти висипав увесь на дахи?
ISA|22|2|Місто сповнене галасом, місто гучне, місто веселе! Побиті твої не побиті мечем, і не повмирали в війні.
ISA|22|3|Усі разом утекли твої проводирі, без вистрілу луку пов'язані усі, хто з тобою знайшовся, пов'язані разом, хоч вони повтікали далеко.
ISA|22|4|Тому я сказав: Відверніться від мене, я гірко заплачу! Не силуйтеся потішати мене, що народу мого дочка поруйнована,
ISA|22|5|бо це день збентеження, і стоптання, і заколоту, день Господа, Бога Саваота, у долині Видіння, день розвалення муру та зойку на горах!
ISA|22|6|А Елам узяв сагайдака, у поході мужів з верхівцями, Кір же витяг щита.
ISA|22|7|І сталось, найкращі долини твої понаповнювались колесницями, а при брамі їздці понаставлені.
ISA|22|8|І відкрив він заслону із Юди, і ти поглянув того дня на зброю дому лісу.
ISA|22|9|І побачили в Місті Давидовім щілини, що багато їх стало, і зібрали води з ставу долішнього;
ISA|22|10|і порахували доми в Єрусалимі, і порозбивали доми ті на зміцнення муру;
ISA|22|11|і зробили ви між двома мурами збір для старого ставка, але ви не дивились на Того, Хто це зробив, Хто це віддавна створив, ви не бачили.
ISA|22|12|І Господь, Бог Саваот того дня був покликав на плач, і на голосіння, і на обстригання волосся, і щоб оперезатись веретою.
ISA|22|13|Та ось радість і втіха: забивають худобу велику та ріжуть худобу дрібну, їдять м'ясо й вино попивають, викрикуючи: Будем їсти та пити, бо взавтра помрем!
ISA|22|14|І відкрив Господь Саваот в мої уші: Напевно не проститься вам беззаконство оце, аж поки ви не помрете, промовив Господь, Бог Саваот.
ISA|22|15|Так промовив Господь, Бог Саваот: Іди, увійди до того управителя, до Шевни, що над домом, та й скажеш:
ISA|22|16|Що ти тут маєш, і хто тут у тебе, що гроба для себе тут видовбав? Ти вирубав на висоті свого гроба, ти видовбав в скелі оселю собі,
ISA|22|17|та Господь тебе з силою викине, лицарю, і хапаючи, схопить тебе,
ISA|22|18|звиваючи, звине тебе на клубок, і кине, як кулю, у землю простору, і там ти помреш, і підуть туди й вози славні твої, о ганьбо ти дому свого господаря!
ISA|22|19|І попхну тебе з стану твого, і скину тебе з того місця, на якому стоїш.
ISA|22|20|І станеться в день той, і покличу Свого раба Еліякима, сина Хілкійїного,
ISA|22|21|і на нього хітона твого одягну, і підпережу Я його твоїм поясом, панування твоє дам у руку його, і стане він батьком для мешканця Єрусалиму та для Юдиного дому!
ISA|22|22|І дам ключа дому Давидового на рамено його, і коли він відчинить, не буде кому замикати, коли ж він замкне, то не буде кому відчиняти.
ISA|22|23|І його Я заб'ю, мов кілка, в певне місце, і стане він домові батька свого троном слави.
ISA|22|24|І повісять на ньому всю славу отцівського дому його, нащадки та дикі відростки, увесь посуд малий від мисок й аж до всякого посуду глиняного!
ISA|22|25|Того дня, говорить Господь Саваот, похитнеться кілок, що був в певне місце забитий, і буде відрубаний та й упаде, і знищений буде тягар, що на ньому, бо так каже Господь!...
ISA|23|1|Пророцтво про Тир. Голосіть, кораблі Таршішу, бо Тир поруйнований: без домів і без входу з кіттейського краю... Так було їм відкрито.
ISA|23|2|Замовчіте, мешканці надмор'я! Сидонські купці, які морем пливуть, тебе переповнили.
ISA|23|3|І насіння Шіхору у водах великих, жниво Ріки то набуток його, і народам він став за торговицю.
ISA|23|4|Соромся, Сидоне, сказало бо море, морська твердиня, говорячи: я не терпіла з породу та не породила, і не виховала юнаків, і дівчат я не викохала.
ISA|23|5|Коли до Єгипту ця звістка прибуде, вони затремтять, як на звістку про Тир.
ISA|23|6|Перейдіть до Таршішу, ридайте, мешканці надмор'я!
ISA|23|7|Чи це ваше місто веселе, що початок його з давен-давна? Його ноги несуть його в далечину оселитися.
ISA|23|8|Хто це постановив був про Тир, що корони давав, що князями бували купці його, а його торговці на землі були в шані?
ISA|23|9|Господь Саваот це призначив, щоб збезчестити пиху всякій славі, щоб усіх славних землі злегковажити.
ISA|23|10|Перейди ти свій край, мов Ріка, дочко Таршішу, вже нема перепони
ISA|23|11|Свою руку простяг Він на море, і царства затряс! Господь про Ханаан наказав, щоб твердиню його зруйнувати,
ISA|23|12|і сказав: Не будеш ти більше радіти, збезчещена дівчино, дочко Сидону! Уставай, перейди до Кіттіму, але й там ти спочинку не матимеш.
ISA|23|13|Це земля ханаанська: на ніщо обернувсь цей народ, Ашшур для пустинних звірів влаштував був її. Вони збудували тут башти вартові, і палаци її повалили, у руїну її обернули.
ISA|23|14|Голосіть, кораблі Таршішу, бо спустошена ваша твердиня!
ISA|23|15|І станеться в день той, Тир буде забутий на сімдесят літ, як дні панування одного царя. По семидесяти літах станеться Тирові, як у тій пісні блудниці:
ISA|23|16|Візьми гусла, і пройдися по місті, забута блуднице! Приємно заграй, багато пісень заспівай, щоб тебе пригадали!
ISA|23|17|І буде, як сімдесят літ покінчиться, згадає про Тира Господь, і знову він братиме плату за блудодійство, і чинитиме блуд з усіма царствами світу на поверхні землі.
ISA|23|18|І стане набуток його та прибуток його із торгівлі Господеві присвяченим. Не буде збиратися він і не буде ховатись, бо набуток його буде тим, хто сидітиме перед обличчям Господнім, щоб їсти досита та мати розкішну одежу.
ISA|24|1|Ось Господь нищить землю й пустошить її, й обертає поверхню її, а мешканців її розпорошує.
ISA|24|2|І стане священик як і народ, а пан немов раб, пані, як невільниця її, продавець немов той покупець, боргувальник немов винуватець, віритель як довжник.
ISA|24|3|Земля буде дощенту зруйнована та пограбована вся, бо це слово Господь проказав,
ISA|24|4|засумує, зів'яне земля, ослабіє й зів'яне вселенна, ослабіють вельможі народу землі...
ISA|24|5|Й осквернилась земля під своїми мешканцями, бо переступили закони, постанову порушили, зламали вони заповіта відвічного...
ISA|24|6|Тому землю прокляття поїло, й одержали кару мешканці її, тому то згоріли мешканці землі, і небагато людей позосталося...
ISA|24|7|Сумує вино молоде, виноградина в'яне, усі радісносерді зідхають,
ISA|24|8|спинилися радощі бубнів, галас веселунів перестав, затихла потіха від гусел!
ISA|24|9|При пісні вина вже не п'ють, став гірким п'янкий напій для тих, хто його попиває...
ISA|24|10|Зруйноване місто спустошене, всі доми позамикані, щоб не ввійти...
ISA|24|11|На вулицях крик за вином, усяка радість померкла, веселість землі на вигнання пішла,
ISA|24|12|позосталося в місті спустошення, і розбита на звалище брама...
ISA|24|13|Бо так буде посеред землі, посеред народів, як при оббиванні оливки, немов при визбируванні, коли збір винограду скінчився.
ISA|24|14|Свій голос підіймуть і будуть радіти, через величність Господню викрикувати голосно будуть від моря.
ISA|24|15|Тому Господа славте на сході, на морських островах Ім'я Господа, Бога Ізраїлевого!
ISA|24|16|Ми чуємо співи від краю землі: Слава Праведному! Але я сказав: Гину, гину, ой горе мені: Грабіжники граблять, і грабуючи, граблять грабіжно!
ISA|24|17|Страх і яма та пастка на тебе, мешканче землі!
ISA|24|18|І станеться, той, хто втікатиме від крику жаху, до ями впаде, хто ж із ями виходить, буде схоплений в пастку, бо відкриті розтвори згори, а підстави землі затремтіли...
ISA|24|19|Земля поруйнована зовсім, земля поторощена, вся земля захиталась...
ISA|24|20|Захиталась земля, немов п'яний, і рухається, мов нічліжний курінь, і вчинився над нею тяжким її гріх, і впала вона, й більш не встане!
ISA|24|21|І станеться в день той, Господь навістить військо висоти на висоті, і земних царів на землі,
ISA|24|22|і будуть зібрані разом, мов в'язні до ями, й у в'язницю вони будуть замкнені, а по днях багатьох будуть навіщені!
ISA|24|23|Місяць тоді засоромиться та застидається сонце, бо Господь Саваот зацарював на Сіонській горі та в Єрусалимі, а перед старішими слава Його!
ISA|25|1|Господи, Ти мій Бог! Я буду Тебе величати, хвалитиму Ймення Твоє, бо Ти чудо вчинив, виконав давні приречення, певную правду!
ISA|25|2|Бо Ти купою каменя місто вчинив, укріплене місто руїною, чужинецький палац перестав бути містом, навіки не буде воно відбудоване!
ISA|25|3|Тому буде хвалити Тебе народ сильний, місто людів насильників буде боятись Тебе,
ISA|25|4|бо твердинею став Ти нужденному, твердинею став для убогого в час його утиску, охороною від хуртовини, тінню від спеки, і дух тих насильників був немов хуртовина на стіну!
ISA|25|5|Як спекоту в пустині, Ти крики чужинців приборкав; як тінню від хмари спекоту, спів насильників так Він приглушить.
ISA|25|6|І вчинить Господь Саваот на горі цій гостину з страв ситих, гостину із вин молодих, із шпікового товщу, із очищених вин молодих.
ISA|25|7|І Він на горі цій понищить заслону, заслону над усіма народами, та покриття, що розтягнене над усіма людами.
ISA|25|8|Смерть знищена буде назавжди, і витре сльозу Господь Бог із обличчя усякого, і ганьбу народу Свого він усуне з усієї землі, бо Господь це сказав.
ISA|25|9|І скажуть в той день: Це наш Бог, що на Нього ми мали надію і Він спас нас! Це Господь, що на Нього ми мали надію, тішмося ж ми та радіймо спасінням Його!
ISA|25|10|Бо Господня рука на горі цій спочине, Моав же на місці своєму потоптаний буде, як солома витоптується у гноївці,
ISA|25|11|і простягне він руки свої серед неї, немов той пливак простягає, щоб пливати, і принизить пиху його Він разом з підступами його рук.
ISA|25|12|А високу твердиню цих мурів твоїх Він розвалить, понизить, на землю їх кине, у порох!
ISA|26|1|Того дня заспівають у Юдинім краї пісню таку: У нас сильне місто! Він чинить спасіння за мури й примурки.
ISA|26|2|Відчиняйте ворота, і хай ввійде люд праведний, хто вірність хоронить!
ISA|26|3|Думку, оперту на Тебе, збережеш Ти у повнім спокої, бо на Тебе надію вона покладає.
ISA|26|4|Надійтеся завжди на Господа, бо в Господі, в Господі вічна твердиня!
ISA|26|5|Бо знизив Він тих, хто замешкує на висоті, неприступне те місто понизив його, Він понизив його до землі, повалив аж у порох його!
ISA|26|6|Його топче нога, ноги вбогого, стопи нужденних...
ISA|26|7|Проста дорога для праведного, путь праведного Ти вирівнюєш.
ISA|26|8|І на дорозі судів Твоїх, Господи, маємо надію на Тебе: За Ймення Твоє та за пам'ять Твою пожадання моєї душі,
ISA|26|9|за Тобою душа моя тужить вночі, також дух мій в мені спозаранку шукає Тебе, бо коли на землі Твої суди, то мешканці світу навчаються правди!
ISA|26|10|Хоч буде безбожний помилуваний, то проте справедливости він не навчиться: у краю правоти він чинитиме лихо, а величности Господа він не побачить!
ISA|26|11|Господи, піднялася рука Твоя високо, та не бачать вони! Нехай же побачать горливість Твою до народу, і нехай посоромляться, хай огонь пожере ворогів твоїх!
ISA|26|12|Ти, Господи, вчиниш нам мир, бо й усі чини наші нам Ти доконав!
ISA|26|13|Господи, Боже наш, панували над нами пани окрім Тебе, та тільки Тобою ми згадуємо Ймення Твоє.
ISA|26|14|Померлі вони не оживуть, мертві не встануть вони, тому Ти навідав та вигубив їх, і затер всяку згадку про них.
ISA|26|15|Розмножив Ти, Господи, люд, розмножив Ти люд, і прославив Себе, всі границі землі Ти далеко посунув.
ISA|26|16|Господи, в горі шукали Тебе, шепіт прохання лили, коли Ти їх картав.
ISA|26|17|Як жінка вагітна до породу зближується, в своїх болях тремтить та кричить, так ми стали, о Господи, перед обличчям Твоїм:
ISA|26|18|ми були вагітними та корчилися з болю, немов би родили ми вітер, ми спасіння землі не вчинили, і мешканці всесвіту не народились...
ISA|26|19|Померлі твої оживуть, воскресне й моє мертве тіло. тому пробудіться й співайте, ви мешканці пороху, бо роса Твоя це роса зцілень, і земля викине мертвих!
ISA|26|20|Іди, мій народе, ввійди до покоїв своїх, і свої двері замкни за собою, сховайся на хвилю малу, поки лютість перейде!
ISA|26|21|Бо Господь ось виходить із місця Свого, навідати провини мешканців землі, кожного з них, і відкриє земля свою кров, і вже не закриє забитих своїх!
ISA|27|1|У той день навідає Господь Своїм твердим, і дужим та сильним мечем левіятана, змія прудкого, і левіятана, змія звивкого, і дракона, що в морі, заб'є.
ISA|27|2|У той день заспівайте про нього, про виноградник принадний:
ISA|27|3|Я Господь, його Сторож, щохвилі його Я напоюю; щоб хто не навідав його, стережу його вдень та вночі,
ISA|27|4|Я гніву не маю. Хто Мені дасть тернину й будяччя, на бій Я піду проти них, і спалю їх усіх!...
ISA|27|5|Хіба буде держатися міцно Мого він захисту, щоб мир учинити зо Мною, зо Мною щоб мир учинити!
ISA|27|6|Яків у майбутньому пустить коріння, розцвітеться Ізраїль і пуп'янки пустить, і поверхню вселенної плодом наповнять.
ISA|27|7|Чи Він уразив його, як уразив того, хто бив був його? Чи він був забитий, як забиті були його вбивники?
ISA|27|8|Ти вигнав його, відіслав його й судишся з ним, вигнав його Своїм подувом сильним у день східнього вітру.
ISA|27|9|Тому вина Якова буде окуплена цим, а це плід увесь: усунення з нього гріха, коли він учинить каміння все жертівника побитим, немов грудки крейди, і не стоятимуть більше Астарти, і стовпи на честь сонця.
ISA|27|10|Бо місто укріплене буде самотнє, мешкання покинене та позоставлене, мов би пустиня, там пастися буде теля, і там буде лежати воно, та понищить галузки його.
ISA|27|11|Коли висохнуть віття його, то поламане буде, жінки прийдуть і спалять його... А що це нерозумний народ, тому милосердя до нього Творець його мати не буде, і не буде ласкавий до нього Створитель його...
ISA|27|12|І станеться в день той, плоди помолотить Господь від бігу ріки до потоку єгипетського, а ви по одному позбирані будете, синове Ізраїля!
ISA|27|13|І станеться в день той, і буде засурмлено в велику сурму, і прийдуть, хто гинув у краї асирійському, і вигнанці до краю єгипетського, і будуть вони на святій горі в Єрусалимі вклонятися Господеві.
ISA|28|1|Горе тобі, Самарії, короні пишноти Єфремлян п'яних, квітці зів'ялій краси його гордости, що лежить на верхів'ї долини врожайної, від вина поп'янілих!
ISA|28|2|Ось потужний та сильний у Господа, мов злива із градом, мов буря руїнна, мов повідь сильна, заливна, його кине на землю із силою!
ISA|28|3|Ногами потоптана буде корона пишноти Єфремлян п'яних,
ISA|28|4|і станеться квітка зів'яла краси його гордости, що на верхів'ї долини врожайної, немов передчасно дозріла та смоква, що її як побачить людина, ковтає її, як вона ще в долоні його!
ISA|28|5|Стане Господь Саваот того дня за прекрасну корону, і за пишний вінок для останку народу Його,
ISA|28|6|і духом права тому, хто сидить у суді, і хоробрістю тим, хто до брами повертає бій!
ISA|28|7|І ось ці від вина позбивались з дороги, і від п'янкого напою хитаються: священик і пророк позбивались з дороги напоєм п'янким, від вина збаламутились, від напою п'янкого хитаються, блудять вони у видіннях, у постановах своїх спотикаються...
ISA|28|8|Бо всі столи повні блювотою калу, аж місця нема!...
ISA|28|9|Кого буде навчати пізнання, і кому виясняти об'явлення буде? Відставлених від молока чи від перс повідлучуваних?
ISA|28|10|Бо на заповідь заповідь, заповідь на заповідь, правило на правило, правило на правило, трохи тут, трохи там.
ISA|28|11|Тому незрозумілими устами й іншою мовою буде казати народові цьому
ISA|28|12|Отой, Хто до них говорив: Це спочинок! Дайте змученому відпочити, і це відпочинок, та вони не хотіли послухати.
ISA|28|13|І станеться їм слово Господа: заповідь на заповідь, заповідь на заповідь, правило на правило, правило на правило, трохи тут, трохи там, щоб пішли та попадали навзнак, і щоб були зламані й впали до пастки й зловилися!...
ISA|28|14|Тому то послухайте слова Господнього, ганьбителі, що пануєте над тим народом, що в Єрусалимі!
ISA|28|15|Бо кажете ви: Заповіта ми склали зо смертю і з шеолом зробили умову. Як перейде той бич, мов вода заливна, то не прийде до нас, бо брехню ми зробили притулком своїм, і в брехні ми сховались!
ISA|28|16|Тому Господь Бог сказав так: Оце поклав каменя Я на Сіоні, каменя випробуваного, наріжного, дорогого, міцно закладеного. Хто вірує в нього, не буде той засоромлений!
ISA|28|17|І право за мірило Я покладу, а справедливість вагою; і притулок брехні град понищить, а сховище води заллють!
ISA|28|18|І заповіт ваш із смертю поламаний буде, а ваша умова з шеолом не втримається: як перейде нищівна кара, то вас вона стопче!
ISA|28|19|Коли тільки перейде вона, вона вас забере, бо щоранку вона переходити буде, удень та вночі, і станеться, тільки з тремтінням ви будете слухати звістку про це...
ISA|28|20|Бо буде постеля коротка, щоб на ній розтягнутись, а покривало вузьке, щоб накритися ним...
ISA|28|21|Бо повстане Господь, немов на горі Перацім; затремтить Він у гніві, немов у долині в Гів'оні, щоб Свій чин учинити, предивний Свій чин, щоб зробити роботу Свою, незвичайну роботу Свою!
ISA|28|22|Тож не насміхайтесь тепер, щоб не стали міцнішими ваші кайдани, бо призначене знищення чув я від Господа, Бога Саваота, про всю землю...
ISA|28|23|Візьміть це до ушей і почуйте мій голос, послухайте пильно й почуйте мій голос!
ISA|28|24|Чи кожного дня оре ратай на посів, ралить землю свою й боронує?
ISA|28|25|Чи ж, як рівною зробить поверхню її, він не сіє чорнуху й не кидає кмин, не розсіває пшеницю та просо й ячмінь на означенім місці, а жито в межах її?
ISA|28|26|І за правом напутив його, його Бог його вивчив цього:
ISA|28|27|Бож не бороною чорнуха молотиться, і коло возове не ходить по кмині, а палицею б'ють чорнуху та києм той кмин.
ISA|28|28|Розтирається збіжжя? Ні, бо його не назавжди молотиться конче, і підганяють коло возове та коні на нього, а не розтирають його.
ISA|28|29|І це вийшло від Господа Саваота, чудова порада Його, і велика премудрість Його!
ISA|29|1|Горе Аріїлу, Аріїлу, місту, що Давид у нім таборував! Рік до року додайте, хай свята закінчать свій круг!
ISA|29|2|І притисну Аріїла, і станеться лемент та плач, і він стане на мене, як огнище Боже.
ISA|29|3|І отаборюся проти тебе навколо, і сторожею стисну тебе, і башти поставлю на тебе.
ISA|29|4|І ти будеш понижений, і будеш з землі говорити, і приглушено буде звучати твоє слово. І стане твій голос з землі, мов померлого дух, і шепотітиме з пороху слово твоє.
ISA|29|5|І буде юрба ворогів твоїх, мов тонкий пил, юрба ж насильників мов полова зниклива, і це станеться нагло, раптовно..
ISA|29|6|Господь Саваот тебе громом та трусом навідає, і шумом великим, вихром та бурею, та огняним їдким полум'ям.
ISA|29|7|І буде, як сон, як видіння нічне та юрба всіх народів, що на Аріїла воюють, і всі, хто воює на нього, і проти твердині його, і хто йому докучає.
ISA|29|8|І буде, мов бачить голодний у сні, ніби їсть, а прокинеться він і порожня душа його, і мов спрагнений бачить у сні, ніби п'є, а прокинеться він і ось змучений, а душа його спрагнена! Так буде натовпові всіх народів, що підуть війною на гору Сіон.
ISA|29|9|Одубійте й дивуйтесь, заліпіть собі очі й осліпніть! Вони повпивалися, та не вином, захитались, та не від п'янкого напою,
ISA|29|10|бо вилив Господь на вас духа глибокого сну та закрив ваші очі, затьмарив пророків і ваших голів та провидців!
ISA|29|11|І буде вам кожне видіння, немов би слова запечатаної книжки, що дають її тому, хто вміє читати, та кажуть: Читай но оце, та відказує той: Не можу, вона ж запечатана.
ISA|29|12|І дають оту книжку тому, хто не вміє читати, та кажуть: Читай но оце, та відказує той: Я не вмію читати.
ISA|29|13|І промовив Господь: За те, що народ цей устами своїми наближується, і губами своїми шанує Мене, але серце своє віддалив він від Мене, а страх їхній до Мене заучена заповідь людська,
ISA|29|14|тому Я ось ізнову предивне вчиню з цим народом, вчиню чудо й диво, і загине мудрість премудрих його, а розум розумних його заховається.
ISA|29|15|Горе тим, що глибоко задум ховають від Господа, і чиняться в темряві їхні діла, і що говорять вони: Хто нас бачить, і хто про нас знає?
ISA|29|16|О, ваша фальшивосте! Чи ганчар уважається рівним до глини? Чи зроблене скаже про майстра свого: Він мене не зробив, а твір про свого творця говоритиме: Він не розуміє цього?
ISA|29|17|Хіба за короткого часу Ліван на садка не обернеться, а садок порахований буде за ліс?
ISA|29|18|І в той день слова книжки почують глухі, а очі сліпих із темноти та з темряви бачити будуть,
ISA|29|19|і сумирні побільшать у Господі радість свою, а люди убогі в Святому Ізраїля тішитись будуть!
ISA|29|20|Бо скінчився насильник, і минувся насмішник, і понищені всі ті, хто дбає про кривду,
ISA|29|21|хто судить людину за слово одне, на того ж, хто судить у брамі, вони ставлять пастку, і праведного випихають обманою.
ISA|29|22|Тому то Господь, що викупив Авраама, сказав домові Якова так: Не буде тепер засоромлений Яків, й обличчя його не поблідне тепер,
ISA|29|23|бо як він серед себе побачить дітей своїх, чин Моїх рук, вони будуть святити Моє Ймення, і посвятять Святого Якового, і будуть боятися Бога Ізраїля!
ISA|29|24|Тоді то хто блудить у дусі, ті розум пізнають, а хто ремствує, ті поуки навчаться!
ISA|30|1|Горе синам неслухняним, говорить Господь, що чинять наради, які не від Мене, і складають умови, та без духу Мого, щоб додати гріх на гріх,
ISA|30|2|що йдуть, щоб зійти до Єгипту, але Моїх уст не питали, щоб захисту у фараона шукати, і щоб сховатися в тіні Єгипту!
ISA|30|3|І стане вам соромом захист отой фараонів, а ховання у тіні Єгипту за ганьбу,
ISA|30|4|бо в Цоані були його провідники, і його посланці до Ханесу прийшли.
ISA|30|5|Вони посоромлені будуть усі за народ, що не буде корисний для них, що не буде на поміч і не на пожиток, а на сором та ганьбу...
ISA|30|6|Пророцтво 4853 про Бегемота 929 півдня 5045. В краю 776 утиску 6869 та переслідування 6695, звідки левиця 3833 та лев 3918, гадюка 660 й огнистий 8314 0 летючий 5774 8789 дракон 8314 0, носять 5375 8799 багатство 2428 своє на хребті 3802 молодих 5895 0 ослюків 5895 0, і скарби 214 свої на верблюжім 1581 горбі 1707 до народу 5971, який не поможе 3276 8686.
ISA|30|7|А Єгипет 4714, його поміч 5826 8799 марна 1892 та пуста 7385, тому то я кликнув 7121 8804 на теє 2063: Рагав 7293, сидіти 7674 0 спокійно 7674 0!
ISA|30|8|Тепер увійди, напиши на таблиці для них, і в книжці спиши це, і нехай на пізніші часи воно буде і свідком навіки.
ISA|30|9|Бо це неслухняний народ, це брехливі сини, сини, що не хочуть послухати науки Господньої,
ISA|30|10|що говорять провидцям: Не бачте! а пророкам: Не пророкуйте правдивого нам, говоріть нам гладеньке, передбачте оманливе,
ISA|30|11|уступіться з дороги, збочте з путі, заберіть з-перед нас Святого Ізраїлевого!
ISA|30|12|Тому промовляє Святий Ізраїлів так: За те, що ви нехтуєте оцим словом, і надію кладете на тиск та крутійство, і на це опираєтеся,
ISA|30|13|тому буде для вас ця провина, як вилім, що має впасти, що зяє на мурі високім, що нагло, раптовно приходить руїна його!
ISA|30|14|І Він поруйнує його, як руйнується посуд ганчарський, розбиваючи без милосердя його, і в уламках його не знайдеться ані черепка, щоб із огнища взяти огню чи води зачерпнути з кринички...
ISA|30|15|Бо так промовляє Господь, Бог, Святий Ізраїлів: Коли ви навернетесь та спочинете, то врятовані будете, сила вам буде в утишенні та в сподіванні. Та ви не хотіли,
ISA|30|16|і казали: О ні, бо на конях втечемо, тому то втікати ви будете, На баских ми поїдемо, тому стануть баскими погоничі ваші!...
ISA|30|17|Від крику одного полине одна тисяча, від крику п'ятьох дременете ви всі, аж зостанетеся, немов щогла ота на вершечку гори, і немов прапор на взгір'ї!
ISA|30|18|І проте Господь буде чекати, щоб помилувати вас, і тому Він підійметься, щоб милосердя вчинити над вами. Бо Господи то Бог правосуддя: блаженні всі ті, хто надію на Нього кладе!
ISA|30|19|Бо ти, о народе в Сіоні, що в Єрусалимі сидиш, плакати не будеш ти плакати: милостивим поправді Він буде до тебе на голос благання твого, і як почує його, відповість Він тобі.
ISA|30|20|І дасть вам Господь хліба в утиску і воду в гнобительстві, та твої вчителі вже не будуть ховатись, і очі твої вчителів твоїх бачити будуть.
ISA|30|21|А коли ви відхилитесь праворуч, чи підете ліворуч, то вуха твої будуть чути те слово, яке позад тебе казатиме: Це та дорога, простуйте ви нею!
ISA|30|22|І нечистим учините ви поволоку бовванів своїх із срібла й покриття на божка золотого свого, розпорошиш ти їх, як нечисте, і геть скажеш йому.
ISA|30|23|І Він пошле дощ на насіння твоє, яким будеш обсіювати землю, та хліб урожаю землі, і поживний та ситий він буде. Того дня на широкім пасовиську пастися буде твоя череда,
ISA|30|24|а воли й віслюки, що оброблюють землю, будуть мішанку їсти солону, лопатою й віялкою перечищену.
ISA|30|25|І на кожній високій горі та на кожному взгір'ї високому будуть струмки та потоки води в день великого бою, коли башти попадають.
ISA|30|26|І світло місяця стане, немов світло сонця, світло ж сонця усемеро буде ясніше, як сімох днів, у той день, як Господь перев'яже зламання народу Свого та загоїть поранення вдару Свого!
ISA|30|27|Ось Імення Господнє приходить здалека, палахкотить Його гнів, і здіймається тяжко: Його уста обурення повні, язик же Його, як жерущий огонь,
ISA|30|28|Його ж дух, як потоп заливний, що до шиї сягає, щоб просіяти люди на ситі погибелі... І буде на щелепах людів вуздечка, що тягне до блуду.
ISA|30|29|Буде пісня для вас, як за ночі освячення свята, і радість сердечна, мов у того, хто ходить з сопілкою, щоб вийти на гору Господню до Скелі Ізраїля.
ISA|30|30|І Господь дасть почути велич голосу Свого, опускання ж рамена Свого покаже у гніві бурхливому та в огняному жерущому полум'ї, у бурі й дощі, та в камінному граді!
ISA|30|31|Бо від голосу Господа буде лякатись Ашшур, що жезлом буде битий.
ISA|30|32|І станеться, кожне ударення кия карання Його, що на нього Господь покладе, буде з бубнами й арфою, і Він рухом Своєї руки воюватиме з ним у боях.
ISA|30|33|Бо давно приготовлений Тофет, приготовлений він і для царя, глибоким, широким учинений; на багатті огню його й дров багатенно, запалить його дух Господній, немов би потока сірчаного!
ISA|31|1|Горе тим, що в Єгипет по поміч ідуть, що на коней спираються, і на колесниці надію свою покладають, вони бо численні! та на верхівців, бо вони дуже сильні! але на Святого Ізраїлевого не дивляться, і до Господа не звертаються!
ISA|31|2|Та мудрий і Він, і спровадить лихе, і Своїх слів не відмінить, і підійметься Він проти дому безбожних, і проти помочі несправедливих.
ISA|31|3|А Єгипет не Бог, а людина, а коні їхні тіло, не дух: як простягне Господь Свою руку, то спіткнеться помагач, впаде і підпомаганий, і разом вони всі погинуть!
ISA|31|4|Бо до мене Господь сказав так: Як муркає лев чи левчук над своєю здобиччю, хоч покликана буде на нього юрба пастухів, він голосу їхнього не лякається, та не боїться їхнього крику, так зійде Господь Саваот воювати на Сіонській горі та на взгір'ї її!
ISA|31|5|Як птахи летючі пташат, так Єрусалима Господь Саваот охоронить, охоронить літаючи, та збереже, пощадить та врятує!
ISA|31|6|Верніться до Того, від Кого далеко відпали, синове Ізраїлеві!
ISA|31|7|Бо дня того обридить собі чоловік божків срібних своїх та бовванів своїх золотих, що вам наробили на гріх руки ваші.
ISA|31|8|І Ашшур упаде від меча того нелюда, і його пожере меч нелюдський; і він побіжить не перед мечем, і стануть його юнаки кріпаками...
ISA|31|9|А скеля його проминеться від страху, і владики його затривожаться перед прапором... Так говорить Господь, що має огонь на Сіоні, а в Єрусалимі у Нього горнило.
ISA|32|1|Тож за праведністю царюватиме цар, а князі володітимуть за правосуддям.
ISA|32|2|І станеться кожен, як захист від вітру, і немов та заслона від зливи, як потоки води на пустині, як тінь скелі тяжкої на спраглій землі...
ISA|32|3|І не будуть заплющені очі видющих, і слухатимуть вуха тих, які слухають!
ISA|32|4|І знання розумітиме серце нерозважних, а язик недорікуватих поспішить говорити виразно.
ISA|32|5|Не будуть вже кликати достойним глупця, а на обманця не скажуть шляхетний,
ISA|32|6|бо глупоту говорить безумний, а серце його беззаконня вчиняє, щоб робити лукавство, та щоб говорити до Господа слово облудне, щоб душу голодного випорожнити й напою позбавити спраглого!
ISA|32|7|А лукавий лихі його чини: він лихе замишляє, щоб нищити скромних словами брехливими, як убогий говорить про право,
ISA|32|8|а шляхетний міркує шляхетне, і стоїть при шляхетному.
ISA|32|9|Устаньте, безжурні жінки, почуйте мій голос, дочки безтурботні, послухайте слова мого!
ISA|32|10|Днів багато на рік ви, безтурботні, тремтітимете, бо збір винограду скінчився, а згромадження плоду не прийде!
ISA|32|11|Тремтіть, ви безжурні, дрижіть, безтурботні, роздягніться, себе обнажіть, опережіться по стегнах!
ISA|32|12|За принадні поля будуть битися в груди, за виноградник урожайний...
ISA|32|13|На землі цій народу мого зійде терен й будяччя, по всіх домах радости спаленина, на місті веселому...
ISA|32|14|Бо палац опущений буде, міський гомін замовкне, Офел та башта навік стануть ямами, радістю диких ослів, пасовиськом черід,
ISA|32|15|аж Дух з височини проллється на нас, а пустиня в садок обернеться, а садок порахований буде за ліс!
ISA|32|16|Тоді пробуватиме право в пустині, на ниві ж родючій сидітиме правда.
ISA|32|17|І буде роботою істини мир, а працею правди спокійність й безпека навіки.
ISA|32|18|І осяде народ мій у мешканні спокійнім, і в безпечних місцях, і в спокійних місцях відпочинку.
ISA|32|19|І буде падати град на повалений ліс, і знизиться місто в долину...
ISA|32|20|Блаженні ви, сівачі понад всякими водами, що відпускаєте ногу волові й ослові на волю!
ISA|33|1|Горе тобі, що пустошиш, хоч сам не спустошений, тобі, що грабуєш, хоч тебе й не грабовано! Коли ти пустошити скінчиш, опустошений будеш, коли грабувати скінчиш, тебе пограбують...
ISA|33|2|Господи, змилуйсь над нами, на Тебе надіємось ми! Будь їхнім раменом щоранку та в час утиску нашим спасінням!
ISA|33|3|Від сильного голосу Твого народи втікатимуть, від Твого вивищення розпорошаться люди.
ISA|33|4|І ваша здобич збереться, як збирають тих коників, як літає ота сарана, так кидатись будуть на неї.
ISA|33|5|Величний Господь, бо на височині пробуває; Він наповнив Сіон правосуддям та правдою.
ISA|33|6|І буде безпека за часу твого, щедрота спасіння, мудрости та пізнання. Страх Господній буде він скарбом його.
ISA|33|7|Тож по вулицях їхні хоробрі кричать, гірко плачуть провісники миру.
ISA|33|8|Биті дороги порожніми стали, нема мандрівця на дорозі! Він зламав заповіта, зневажив міста, злегковажив людину...
ISA|33|9|Сумує та слабне земля, засоромився й в'яне Ливан, став Сарон немов пуща, Башан та Кармел своє листя зронили...
ISA|33|10|Нині воскресну, говорить Господь, нині прославлюсь, нині буду вознесений!
ISA|33|11|Заваготієте сіном, стерню ви породите; дух ваш огонь, який вас пожере...
ISA|33|12|І стануть народи за місце паління вапна, за тернину потяту, і будуть огнем вони спалені...
ISA|33|13|Почуйте, далекі, що Я був зробив, і пізнайте, близькі, Мою силу!
ISA|33|14|Затривожились грішні в Сіоні, і трепет безбожних обняв... Хто з нас мешкатиме при жерущім огні? Хто з нас мешкати буде при вічному огнищіу?
ISA|33|15|Хто ходить у правді й говорить правдиве, хто бридиться зиском насилля, хто долоні свої випорожнює, щоб хабара не тримати, хто ухо своє затикає, щоб не чути про кровопролиття, і зажмурює очі свої, щоб не бачити зла,
ISA|33|16|той перебуватиме на високостях, скельні твердині його недоступна оселя, його хліб буде даний йому, вода йому завжди запевнена!
ISA|33|17|Твої очі побачать Царя в Його пишній красі, будуть бачити землю далеку.
ISA|33|18|Твоє серце роздумувати буде про страх: Де Той, Хто рахує? Де Той, Хто все важить? Де Той, Хто обчислює башти?
ISA|33|19|Уже не побачиш народу зухвалого, народу глибокомовного, якого не можна було б розібрати, незрозумілоязикого, якого не можна було б зрозуміти.
ISA|33|20|Подивись на Сіон, на місто наших святкових зібрань, очі твої вгледять Єрусалим, мешкання спокійне, скинію ту незрушиму, кілля її не порушаться ввік, а всі шнури її не порвуться.
ISA|33|21|Бо величний Господь для нас тільки отам, місце потоків й просторих річок, не ходить по ньому весловий байдак, і міцний корабель не перейде його.
ISA|33|22|Бо Господь наш суддя, Господь законодавець для нас, Господь то наш цар, і Він нас спасе!
ISA|33|23|Опустилися шнури твої, не зміцняють підвалини щогли своєї, вітрил не натягують. Тоді будуть ділити награбовану здобич, і навіть криві грабуватимуть.
ISA|33|24|І не скаже мешканець Я хворий! І прощені будуть провини народу, що в ньому живе.
ISA|34|1|Наблизьтеся, люди, щоб чути, народи ж, послухайте! Хай почує земля та все те, що на ній, вселенна й нащадки її!
ISA|34|2|Господній бо гнів на всі люди, а лютість на все їхнє військо: Він їх учинив за закляття, віддав їх на різь!
ISA|34|3|І їхні побиті розкидані будуть, а з трупів їхніх здійметься сморід, розтопляться гори від їхньої крови...
ISA|34|4|І небесні світила усі позникають, а небо, як звій книжковий, буде звинене, і всі його зорі попадають, як спадає оте виноградове листя, й як спадає з фіґовниці плід недозрілий!...
ISA|34|5|Бо на небі напоєний меч Мій, оце він на Едома спускається та на заклятий народ Мій на суд:
ISA|34|6|меч Господній наповнився кров'ю, став ситий від лою, від крови телят та козлів, від лою баранячих нирок, бо Господу жертва в Боцрі й різанина велика в едомській землі...
ISA|34|7|І буйволи зійдуть із ними, і телиці з биками, і напоїться кров'ю їхній край і насититься туком їхній порох,
ISA|34|8|бо це буде день помсти Господньої, рік заплати за заколот проти Сіону!
ISA|34|9|І переміняться в смолу потоки його, його ж порох у сірку, і смолою палючою стане їхній край...
ISA|34|10|Не погасне вночі ані вдень, дим його підійматися буде повік, з роду в рід опустошений буде, на віки віків не перейде по ньому ніхто.
ISA|34|11|І посяде його пелікан та їжак, і перебуватимуть в ньому сова та ворона, і над ним Він розтягне мірильного шнура спустошення та виска знищення...
ISA|34|12|Не буде шляхетних у ньому, щоб царство там проголосити, і стануть нічим усі князі його.
ISA|34|13|І буде тернина рости по палатах його, кропива й будяччя в твердинях його, і він стане мешканням шакалів, подвір'ям для струсів...
ISA|34|14|І будуть стрічатися там дикі звірі пустинні з гієнами, а польовик буде кликати друга свого; Ліліт тільки там заспокоїться і знайде собі відпочинок!
ISA|34|15|Там кублитись буде скакуча гадюка й складатиме яйця, і висиджувати буде та вигріватиме яйця свої... Там теж яструби будуть збиратись один до одного...
ISA|34|16|Пошукайте у книзі Господній й читайте: Із них не забракне ні одного, не будуть шукати один одного, бо уста Його то вони наказали, а Дух Його Він їх зібрав!
ISA|34|17|І Він кинув для них жеребка, а рука Його шнуром мірильним його поділила для них, і посядуть його аж повік, з роду в рід будуть в нім пробувати!
ISA|35|1|Звеселиться пустиня та пуща, і радітиме степ, і зацвіте, мов троянда,
ISA|35|2|розцвітаючи, буде цвісти та радіти, буде втіха також та співання, бо дана йому буде слава Лівану, пишнота Кармелу й Сарону, вони бачитимуть славу Господа, велич нашого Бога!
ISA|35|3|Зміцніть руки охлялі, і підкріпіть спотикливі коліна!
ISA|35|4|Скажіть тим, що вони боязливого серця: Будьте міцні, не лякайтесь! Ось ваш Бог, помста прийде, як Божа відплата, Він прийде й спасе вас!
ISA|35|5|Тоді то розплющаться очі сліпим і відчиняться вуха глухим,
ISA|35|6|Тоді буде скакати кривий, немов олень, і буде співати безмовний язик, бо води в пустині заб'ють джерелом, і потоки в степу!
ISA|35|7|І місце сухе стане ставом, а спрагнений край збірником вод джерельних; леговище шакалів, в якім спочивали, стане місцем тростини й папірусу.
ISA|35|8|І буде там бита дорога та путь, і будуть її називати: дорога свята, не ходитиме нею нечистий, і вона буде належати народові його; не заблудить також нерозумний, як буде тією дорогою йти.
ISA|35|9|Не буде там лева, і дика звірина не піде на неї, не знайдеться там, а будуть ходити лиш викуплені.
ISA|35|10|І Господні викупленці вернуться та до Сіону зо співом увійдуть, і радість довічна на їхній голові! Веселість та радість осягнуть вони, а журба та зідхання втечуть!
ISA|36|1|І сталося, чотирнадцятого року царя Єзекії прийшов Санхерів, цар асирійський, на всі укріплені Юдині міста, та й захопив їх.
ISA|36|2|І послав асирійський цар великого чашника з Лахішу до Єрусалиму, до царя Єзекії, з великим військом, і він став при водоводі горішнього ставу, на битій дорозі поля Валюшників.
ISA|36|3|І вийшов до нього Еліяким, син Хілкійїн, начальник палати, і писар Шевна, та Йоах, син Асафів, канцлер.
ISA|36|4|І сказав їм великий чашник: Скажіть Єзекії: Отак сказав великий цар, цар асирійський: Що це за надія, на яку ти надієшся?
ISA|36|5|Чи думаєш ти, що слово уст, то вже рада та сила до війни? На кого тепер надієшся, що збунтувався проти мене?
ISA|36|6|Ось ти надіявся опертися на оту поламану очеретину, на Єгипет, що коли хто опирається на неї, то вона входить у долоню йому, і продірявлює її. Отакий фараон, цар єгипетський, для всіх, хто надіється на нього!
ISA|36|7|А коли ти скажеш мені: Ми надіємось на Господа, Бога нашого, то чи ж Він не той, що Єзекія повсовував пагірки його та жертівники його, і сказав Юді та Єрусалимові: перед оцим тільки жертівником будете вклонятися?
ISA|36|8|А тепер увійди но в союз з моїм паном, асирійським царем, і я дам тобі дві тисячі коней, якщо ти зможеш собі дати на них верхівців.
ISA|36|9|І як же ти проженеш хоч одного намісника з найменших рабів мого пана? А ти собі надіявся на Єгипет ради колесниць та верхівців!
ISA|36|10|Тепер же, чи без волі Господа прийшов я на цей край, щоб знищити його? Господь сказав був мені: Піди на той край та й знищ його!
ISA|36|11|І сказав Еліяким, і Шевна та Йоах до великого чашника: Говори до своїх рабів по-арамейському, бо ми розуміємо, і не говори до нас по-юдейському в голос при тих людях, що на мурі.
ISA|36|12|І сказав великий чашник: Чи пан мій послав мене говорити ці слова до твого пана та до тебе? Хіба не до цих людей, що сидять на мурі, щоб із вами їсти свій кал та пити свою сечу?
ISA|36|13|І став великий чашник, і кликнув гучним голосом по-юдейському, і сказав: Послухайте слів великого царя, царя асирійського!
ISA|36|14|Так сказав цар: Нехай не дурить вас Єзекія, бо він не зможе врятувати вас!
ISA|36|15|І нехай не запевняє вас Єзекія Господом, говорячи: Рятуючи, врятує вас Господь, і не буде дано цього міста в руку царя асирійського.
ISA|36|16|Не слухайте Єзекії, бо так сказав цар асирійський: Примиріться зо мною, та й вийдіть до мене, та й їжте кожен свій виноград та кожен фіґу свою, і пийте кожен воду зо своєї копанки,
ISA|36|17|аж поки я не прийду й не візьму вас до краю такого ж, як ваш край, до краю збіжжя та виноградного соку, до краю хліба та виноградників.
ISA|36|18|Щоб не намовив вас Єзекія, говорячи: Господь порятує нас! Чи врятували боги тих народів, кожен свій край від руки асирійського царя?
ISA|36|19|Де боги Хамату та Арпаду? Де боги Сефарваїму? І чи врятували вони Самарію від моєї руки?
ISA|36|20|Котрий з-поміж усіх богів цих країв урятував свій край від моєї руки, то невже ж Господь урятує Єрусалим від моєї руки?
ISA|36|21|І мовчали вони, і не відповіли ані слова, бо це був наказ царя, що сказав Не відповідайте йому!
ISA|36|22|І прийшов Еліяким, син Хілкійїн, начальник палати, і писар Шевна, і Йоах, Асафів син, канцлер, з роздертими шатами, до Єзекії, і донесли йому слова великого чашника.
ISA|37|1|І сталося, як почув це цар Єзекія, то роздер свої шати та накрився веретою, і ввійшов до Господнього дому...
ISA|37|2|І послав він Еліякима, керівника палати, і писаря Шевну, та старших із священиків, покритих веретами, до пророка Ісаї, Амосового сина.
ISA|37|3|І сказали вони до нього: Так сказав Єзекія: Цей день це день горя й картання та наруги! Бо підійшли діти аж до виходу утроби, та немає сили породити!
ISA|37|4|Може почує Господь, Бог твій, слова великого чашника, що його послав асирійський цар, пан його, на образу Живого Бога, і Господь, Бог твій, покарає за слова, які чув, а ти принесеш молитву за решту, що ще знаходиться...
ISA|37|5|І прийшли раби царя Єзекії до Ісаї.
ISA|37|6|І сказав їм Ісая Так скажете вашому панові: Так сказав Господь: Не бійся тих слів, що почув ти, якими ображали Мене слуги асирійського царя.
ISA|37|7|Ось Я дам в нього духа, і він почує звістку, і вернеться до свого краю. І Я вражу його мечем у його краї!
ISA|37|8|І вернувся великий чашник, і знайшов асирійського царя, що воював проти Лівни, бо почув, що той рушив із Лахішу.
ISA|37|9|І він почув про Тіргаку, царя етіопського, таке: Він вийшов воювати з тобою! І почув він, і послав послів до Єзекії, говорячи:
ISA|37|10|Так скажете до Єзекії, Юдиного царя, говорячи: Нехай не зводить тебе Бог твій, на Якого ти надієшся, кажучи: Не буде даний Єрусалим у руку асирійського царя.
ISA|37|11|Ось ти чув, що зробили асирійські царі всім краям, щоб учинити їх закляттям, а ти будеш урятований?
ISA|37|12|Чи їх урятували боги тих народів, яких понищили батьки мої: Ґозана, і Харана, і Рецефа, і синів Едена, що в Телассарі?
ISA|37|13|Де він, цар Хамату, і цар Арпаду, і цар міста Сефарваїму, Гени та Івви?
ISA|37|14|І взяв Єзекія ті листи з руки послів, і прочитав їх, і ввійшов у Господній дім. І Єзекія розгорнув одного листа перед Господнім лицем.
ISA|37|15|І Єзекія молився перед Господнім лицем, говорячи:
ISA|37|16|Господи Саваоте, Боже Ізраїлів, що сидиш на Херувимах! Ти Той єдиний Бог для всіх царств землі, Ти створив небеса та землю!
ISA|37|17|Нахили, Господи, ухо Своє та й почуй! Відкрий, Господи, очі Свої та й побач, і почуй всі слова Санхеріва, що прислав ображати Живого Бога.
ISA|37|18|Справді, Господи, асирійські царі попустошили всі народи та їхні краї.
ISA|37|19|І кинули вони їхніх богів на огонь, бо не боги вони, а тільки чин людських рук, дерево та камінь, і понищили їх.
ISA|37|20|А тепер, Господи, Боже наш, спаси нас від руки його, і нехай знають усі царства землі, що Ти Господь, Бог єдиний!
ISA|37|21|І послав Ісая, Амосів син, до Єзекії, говорячи: Так сказав Господь, Бог Ізраїлів: Я почув те, про що ти молився до Мене, про Санхеріва, царя асирійського.
ISA|37|22|Ось те слово, яке Господь говорив про нього: Гордує тобою, сміється із тебе дівиця, сіонська дочка, вслід тобі головою хитає дочка Єрусалиму!
ISA|37|23|Кого лаяв ти та ображав, і на кого повищив ти голос та вгору підніс свої очі? На Святого Ізраїлевого!
ISA|37|24|Через рабів своїх Господа ти ображав та казав: Із безліччю своїх колесниць я вийшов на гори високі, на боки Лівану, і позрубую кедри високі його, добірні його кипариси, і зберусь на вершок його височини, в гущину його саду,
ISA|37|25|я копаю та п'ю чужу воду, і стопою своєї ноги повисушую я всі єгипетські ріки!
ISA|37|26|Хіба ти не чув, що віддавна зробив Я оце, що за днів стародавніх Я це був створив? Тепер же спровадив Я це, що ти нищиш міста поукріплювані, на купу румовищ обертаєш їх.
ISA|37|27|А мешканці їхні безсилі, настрашені та побентежені, вони стали, як зілля оте польове, мов трава зеленіюча, як трава на дахах, як попалене збіжжя, яке не доспіло...
ISA|37|28|І сидіння твоє, і твій вихід та вхід твій Я знаю, і твоє проти Мене обурення.
ISA|37|29|За твоє проти Мене обурення, що гординя твоя надійшла до вух Моїх, то на ніздрі твої Я сережку привішу, а вудило Моє в твої уста, і тебе поверну Я тією дорогою, якою прийшов ти!
ISA|37|30|А оце тобі знак: їжте цього року збіжжя самосійне, а другого року саморосле, а третього року сійте та жніть, і садіть виноградники, та й їжте їхній плід.
ISA|37|31|А врятоване Юдиного дому, що лишилося, пустить коріння додолу, і свого плода дасть угору.
ISA|37|32|Бо з Єрусалиму вийде позостале, а рештки з гори Сіон. Ревність Господа Саваота зробить це.
ISA|37|33|Тому так сказав Господь про асирійського царя: Він не ввійде до міста цього, і туди він не кине стріли, і щитом її не попередить, і вала на нього не висипле.
ISA|37|34|Якою дорогою прийде, то нею й повернеться, у місто ж оце він не ввійде, говорить Господь!
ISA|37|35|І це місто Я обороню на спасіння його ради Себе та ради Давида, Мого раба!
ISA|37|36|І вийшов Ангол Господній, і забив в асирійському таборі сто й вісімдесят і п'ять тисяч. І повставали рано вранці, аж ось усі тіла мертві...
ISA|37|37|А Санхерів, асирійський цар, рушив та й пішов, і вернувся, й осівся в Ніневії.
ISA|37|38|І сталося, коли він молився в домі Нісроха, свого бога, то сини його Адраммелех та Шар'ецер убили його мечем, а самі втекли до краю Арарат... А замість нього зацарював син його Есар-Хаддон.
ISA|38|1|Тими днями смертельно захворів був Єзекія. І прийшов до нього Ісая, Амосів син, пророк, і сказав до нього: Так сказав Господь: Заряди своєму домові, бо ти вмираєш і не будеш жити...
ISA|38|2|І відвернув Єзекія обличчя своє до стіни, і помолився до Господа,
ISA|38|3|та й сказав: О, Господи, згадай же, що я ходив перед обличчям Твоїм правдою та цілим серцем, і робив я добре в очах Твоїх! І заплакав Єзекія ревним плачем!
ISA|38|4|І було Господнє слово до Ісаї, говорячи:
ISA|38|5|Іди й скажеш до Єзекії: Так сказав Господь, Бог батька твого Давида: Почув Я молитву твою, побачив Я сльозу твою! Ось Я додаю до днів твоїх п'ятнадцять літ,
ISA|38|6|і з руки асирійського царя врятую тебе та це місто, й обороню це місто.
ISA|38|7|І оце тобі знак від Господа, що Господь зробить ту річ, про яку говорив:
ISA|38|8|ось я вертаю тінь ступеня, що від сонця зійшла на ступені Ахазові, назад на десять ступенів. І вернулося сонце на десять ступенів тими ступенями, якими зійшло було.
ISA|38|9|Ось писання Єзекії, Юдиного царя, коли він був захворів та видужав з своєї хвороби:
ISA|38|10|Я сказав був: Опівдні днів своїх відійду до шеолових брам, решти років своїх я не матиму...
ISA|38|11|Я сказав: Не побачу я Господа, Господа в краї живих, уже між мешканцями царства померлих не побачу людини...
ISA|38|12|Домівка моя вже розібрана, і від мене відібрана, немов той пастуший намет; я життя своє звинув, мов ткач, від основи мене Він відірве, покінчить мене з дня до ночі...
ISA|38|13|Я кричав аж до ранку... Він, як лев, поторощить всі кості мої, з дня до ночі покінчить зо мною...
ISA|38|14|Пищу я, мов ластівка чи журавель, воркочу, мов той голуб; заниділи очі мої, визираючи до високости... Господи, причавлений я, поручися за мене!
ISA|38|15|Що маю сказати? А що Він сказав був мені, те й вчинив. Тихо змандрую всі літа свої через гіркість моєї душі!
ISA|38|16|Господи, на них, на словах Твоїх, житимуть люди, і в усьому цьому життя моєї душі, уздоров же мене й оживи Ти мене!
ISA|38|17|Ось терпіння це вийшло мені на добро, Ти стримав від гробу гниття мою душу, бо Ти кинув за спину Свою всі гріхи мої,
ISA|38|18|бо не буде ж шеол прославляти Тебе, смерть не буде Тебе вихваляти... Не мають надії на правду Твою ті, хто сходить до гробу.
ISA|38|19|Живий, тільки живий Тебе славити буде, як я ось сьогодні, батько синам розголосить про правду Твою!
ISA|38|20|Господь на спасіння мені, і ми будем співати пісноспіви свої у домі Господнім по всі дні мого життя!
ISA|38|21|А Ісая сказав: Нехай візьмуть грудку фіґ, і нехай розітруть на тому гнояку, і видужає!
ISA|38|22|А Єзекія промовив: Який знак, що я ввійду до Господнього дому?
ISA|39|1|Того часу послав Меродах-Бал'адан, син Бал'аданів, вавилонський цар, листи та дарунка до Єзекії, бо прочув був, що той захворів та видужав.
ISA|39|2|І радів ними Єзекія, і показав їм скарбницю свою, срібло, і золото, і пахощі, і добру оливу, і всю зброївню свою, і все, що знаходилося в його скарбницях. Не було речі, якої не показав би їм Єзекія в домі своїм та в усім володінні своїм.
ISA|39|3|І прийшов пророк Ісая до царя Єзекії та й сказав до нього: Що говорили ці люди? І звідки вони прийшли до тебе? А Єзекія сказав: Вони прийшли до мене з далекого краю, з Вавилону.
ISA|39|4|І той сказав: Що вони бачили в домі твоїм? І Єзекія сказав: Усе, що в домі моїм, вони бачили, не було речі, якої не показав би я їм у скарбницях своїх.
ISA|39|5|І сказав Ісая до Єзекії: Послухай же слова Господа Саваота:
ISA|39|6|Ось приходять дні, і все, що в домі твоєму, і що були зібрали батьки твої аж до цього дня, буде винесене аж до Вавилону. Нічого не позостанеться, говорить Господь...
ISA|39|7|А з синів твоїх, що вийдуть із тебе, яких ти породиш, заберуть, і вони будуть евнухами в палатах вавилонського царя!...
ISA|39|8|І сказав Єзекія до Ісаї: Добре Господнє слово, яке ти сказав! І подумав собі: Так, мир та безпека буде за моїх днів!...
ISA|40|1|Утішайте, втішайте народа Мого, говорить ваш Бог!
ISA|40|2|Промовляйте до серця Єрусалиму, і закличте до нього, що виповнилась його доля тяжка, що вина йому вибачена, що він за свої всі гріхи вдвоє взяв з руки Господа!
ISA|40|3|Голос кличе: На пустині вготуйте дорогу Господню, в степу вирівняйте битий шлях Богу нашому!
ISA|40|4|Хай підійметься всяка долина, і хай знизиться всяка гора та підгірок, і хай стане круте за рівнину, а пасма гірські за долину!
ISA|40|5|І з'явиться слава Господня, і разом побачить її кожне тіло, бо уста Господні оце прорекли!
ISA|40|6|Голос кличе: Звіщай! Я ж спитав: Про що буду звіщати? Всяке тіло трава, всяка ж слава як цвіт польовий:
ISA|40|7|трава засихає, а квітка зів'яне, як подих Господній повіє на неї!... Справді, народ то трава:
ISA|40|8|Трава засихає, а квітка зів'яне, Слово ж нашого Бога повіки стоятиме!
ISA|40|9|На гору високу зберися собі, благовіснику Сіону, свого голоса сильно підвищ, благовіснику Єрусалиму! Підвищ, не лякайся, скажи містам Юди: Ось Бог ваш!
ISA|40|10|Ось прийде Господь, Бог, як сильний, і буде рамено Його панувати для Нього! Ось із Ним нагорода Його, а перед обличчям Його відплата Його.
ISA|40|11|Він отару Свою буде пасти, як Пастир, раменом Своїм позбирає ягнята, і на лоні Своєму носитиме їх, дійняків же провадити буде!
ISA|40|12|Хто води поміряв своєю долонею, а п'ядею виміряв небо, і третиною міри обняв пил землі, і гори ті зважив вагою, а взгір'я шальками?
ISA|40|13|Хто Господнього Духа збагнув, і де та людина, що ради свої подавала Йому?
ISA|40|14|З ким радився Він, і той напоумив Його, та навчав путі права, і пізнання навчив був Його, і Його напоумив дороги розумної?
ISA|40|15|Таж народи як крапля з відра, а важать як порох на шальках! Таж Він острови підіймає, немов ту пилинку!
ISA|40|16|І Ливана не вистачить на запаління жертовне, не стане й звір'я його на цілопалення!
ISA|40|17|Насупроти Нього всі люди немов би ніщо, пораховані в Нього марнотою та порожнечею.
ISA|40|18|І до кого вподобите Бога, і подобу яку ви поставите поруч із Ним?
ISA|40|19|Майстер божка відливає, золотар же його криє золотом, та виливає йому срібляні ланцюжки.
ISA|40|20|Убогий на дара такого бере собі дерево, що не гниє, розшукує вправного майстра, щоб поставив божка, який не захитається.
ISA|40|21|Хіба ви не знаєте, чи ви не чули, чи вам не сповіщено здавна було, чи ви не зрозуміли підвалин землі?
ISA|40|22|Він Той, Хто сидить понад кругом землі, а мешканці її немов та сарана. Він небо простяг, мов тканину тонку, і розтягнув Він його, мов намета на мешкання.
ISA|40|23|Він Той, Хто князів обертає в ніщо, робить суддів землі за марноту:
ISA|40|24|вони не були ще посаджені, і не були ще посіяні, і пень їхній в землі ще не закорінився, та як тільки на них Він дмухнув, вони повсихали, і буря понесла їх, мов ту солому!
ISA|40|25|І до кого Мене прирівняєте, і йому буду рівний? говорить Святий.
ISA|40|26|Підійміть у височину ваші очі й побачте, хто те все створив? Той, Хто зорі виводить за їхнім числом та кличе ім'ям їх усіх! І ніхто не загубиться через всесильність та всемогутність Його.
ISA|40|27|Пощо говориш ти, Якове, і кажеш, Ізраїлю: Закрита дорога моя перед Господом, і від Бога мого відійшло моє право.
ISA|40|28|Хіба ж ти не знаєш, або ти не чув: Бог відвічний Господь, що кінці землі Він створив? Він не змучується та не втомлюється, і не збагненний розум Його.
ISA|40|29|Він змученому дає силу, а безсилому міць.
ISA|40|30|І помучаться хлопці й потомляться, і юнаки спотикнутись спіткнуться,
ISA|40|31|а ті, хто надію складає на Господа, силу відновлять, крила підіймуть, немов ті орли, будуть бігати і не потомляться, будуть ходити і не помучаться!
ISA|41|1|Послухайте мовчки Мене, острови, а народи, чекайте навчання Мого! Хай підійдуть і скажуть: Приступімо всі разом на суд!
ISA|41|2|Хто зо сходу того пробудив, що його супроводить в ході перемога? Він народи дає перед ним та царів на топтання, їхнього меча обертає на порох, його лука в солому розвіяну.
ISA|41|3|Він жене їх, спокійно дорогою йде, якою він не переходив ногами своїми.
ISA|41|4|Хто вчинив та зробив це? Той, хто роди покликав віддавна: Я, Господь, перший, і з останніми Я той же Самий!
ISA|41|5|Бачили це острови та жахалися, кінці землі трипотіли, наближувались та приходили.
ISA|41|6|Один одному допомагає і говорить до брата свого: Будь міцний!
ISA|41|7|І підбадьорує майстер золотаря, а той, хто молотом гладить, того, хто б'є на ковадлі, і каже про споєння: Добре воно! і його зміцнює цвяхами, щоб не хиталось.
ISA|41|8|Та ти, о Ізраїлю, рабе Мій, Якове, що Я тебе вибрав, насіння Авраама, друга Мого,
ISA|41|9|ти, якого Я взяв був із кінців землі та покликав тебе із окраїн її, і сказав був до тебе: Ти раб Мій, Я вибрав тебе й не відкинув тебе,
ISA|41|10|не бійся, з тобою бо Я, і не озирайсь, бо Я Бог твій! Зміцню Я тебе, і тобі поможу, і правицею правди Своєї тебе Я підтримаю.
ISA|41|11|Отож, засоромляться та зніяковіють усі проти тебе запалені, стануть нічим та погинуть твої супротивники.
ISA|41|12|Шукатимеш їх, але їх ти не знайдеш, своїх супротивників; стануть нічим та марнотою ті, хто провадить війну проти тебе.
ISA|41|13|Бо Я Господь, Бог твій, що держить тебе за правицю й говорить до тебе: Не бійся, Я тобі поможу!
ISA|41|14|Не бійся, ти Яковів черве, ти жменько Ізраїлева: Я тобі поможу, говорить Господь, і твій Викупитель Святий Ізраїлів!
ISA|41|15|Ось зроблю Я тебе молотаркою гострою, новою, зубчастою, помолотиш ти гори та їх поторощиш, а підгірки половою вчиниш!
ISA|41|16|Перевієш їх ти, й вітер їх рознесе, і буря їх розпорошить, і ти будеш утішатися Господом, будеш хвалитись Святим Ізраїлевим.
ISA|41|17|Убогі та бідні шукають води, та нема, язик їхній від прагнення висох, Я, Господь, і їх вислухаю, Бог Ізраїлів, не лишу їх!
ISA|41|18|Я ріки відкрию на лисих горах, а джерела посеред долин, оберну Я пустиню на озеро водне, а землю суху на джерела!
ISA|41|19|На пустиню дам кедра, акацію, мирта й маслину, поставлю Я разом в степу кипариса та явора й бука,
ISA|41|20|щоб разом побачили й знали, і пересвідчились та зрозуміли, що Господня рука це зробила, і створив це Святий Ізраїлів!
ISA|41|21|Принесіть свою справу, говорить Господь, припровадьте Мені свої докази, каже Цар Яковів.
ISA|41|22|Хай підійдуть і хай нам розкажуть, що трапиться! Виясніть справи минулі, що вони є, а ми серце наше на те покладемо й пізнаємо їхній кінець, або сповістіть про майбутнє.
ISA|41|23|Розкажіть наперед про майбутнє, і пізнаємо ми, що ви боги. Отож, учиніть ви добро чи зробіть що лихе, щоб ми здивувались і разом побачили.
ISA|41|24|Та ви менш від нічого, і менший ваш чин від марноти, гидота, хто вас вибирає!
ISA|41|25|Я з півночі мужа збудив і прийшов він, зо схід сонця в Ім'я Моє кличе, і він буде чавити князів, мов ту грязюку, й як ганчар глину топче!
ISA|41|26|Хто сказав це віддавна, щоб знали те ми, і щоб наперед ми сказали: Це правда? Та ніхто не сказав, і ніхто не повів, і ніхто не почув ваших слів...
ISA|41|27|Я перший сказав до Сіону: Оце, то вони! А Єрусалимові дам благовісника.
ISA|41|28|І Я дивлюсь, та нікого нема, і немає між ними порадника, щоб відповіли, коли їх запитаю.
ISA|41|29|Тож ніщо всі вони, їхні чини марнота, вітер та порожнеча їхні ідоли!
ISA|42|1|Оце Отрок Мій, що Я підпираю Його, Мій Обранець, що Його полюбила душа Моя. Я злив Свого Духа на Нього, і Він правосуддя народам подасть.
ISA|42|2|Він не буде кричати, і кликати не буде, і на вулицях чути не дасть Свого голосу.
ISA|42|3|Він очеретини надломленої не доломить, і ґнота тліючого не погасить, буде суд видавати за правдою.
ISA|42|4|Не втомиться Він, і не знеможеться, поки присуду не покладе на землі, і будуть чекати Закона Його острови.
ISA|42|5|Говорить отак Бог, Господь, що створив небеса і їх розтягнув, що землю простяг та все те, що із неї виходить, що народові на ній Він дихання дає, і духа всім тим, хто ходить по ній.
ISA|42|6|Я, Господь, покликав Тебе в справедливості, і буду міцно тримати за руки Тебе, і Тебе берегтиму, і дам Я Тебе заповітом народові, за Світло поганам,
ISA|42|7|щоб очі відкрити незрячим, щоб вивести в'язня з в'язниці, а з темниці тих мешканців темряви!
ISA|42|8|Я Господь, оце Ймення Моє, і іншому слави Своєї не дам, ні хвали Своєї божкам.
ISA|42|9|Речі давні прийшли ось, нові ж Я повім, дам почути вам про них, поки виростуть.
ISA|42|10|Заспівайте для Господа пісню нову, від краю землі Йому хвалу! Нехай шумить море, і все, що є в ньому, острови та їхні мешканці!
ISA|42|11|Хай голосно кличуть пустиня й міста її, оселі, що в них проживає Кедар! Хай виспівують мешканці скелі, хай кричать із вершини гірської!
ISA|42|12|Нехай Господу честь віддадуть, і на островах Його славу звіщають!
ISA|42|13|Господь вийде, як лицар, розбудить завзяття Своє, як вояк, підійме Він окрик та буде кричати, переможе Своїх ворогів!
ISA|42|14|Я відвіку мовчав, мовчазний був та стримувався, а тепер Я кричатиму, мов породілля! буду тяжко зідхати й хапати повітря!
ISA|42|15|Спустошу Я гори й підгірки, і всі їхні зілля посушу, і річки оберну в острови, і стави повисушую!
ISA|42|16|І Я попроваджу незрячих дорогою, якої не знають, стежками незнаними їх поведу, оберну перед ними темноту на світло, а нерівне в рівнину. Оце речі, які Я зроблю, і їх не покину!
ISA|42|17|Відступлять назад, посоромляться соромом ті, хто надію складав на божка, хто бовванам казав: Ви наші боги!
ISA|42|18|Почуйте, глухі, а незрячі, прозріте, щоб бачити!
ISA|42|19|Хто сліпий, як не раб Мій, а глухий, як посол Мій, що Я посилаю його? Хто сліпий, як довірений, і сліпий, як раб Господа?
ISA|42|20|Ти бачив багато, але не зберіг, мав вуха відкриті, але не почув.
ISA|42|21|Господь захотів був того ради правди Своєї, збільшив та прославив Закона.
ISA|42|22|Але він народ попустошений та поплюндрований; усі вони по печерах пов'язані та по в'язницях поховані; стали вони за грабіж, і немає визвольника, за здобич, й немає того, хто б сказав: Поверни!
ISA|42|23|Хто з вас візьме оце до вух, на майбутнє почує й послухає?
ISA|42|24|Хто Якова дав на здобич, а Ізраїля грабіжникам? Хіба ж не Господь, що ми проти Нього грішили були і не хотіли ходити путями Його, а Закона Його ми не слухали?
ISA|42|25|І Він вилив на нього жар гніву Свого та насилля війни, що палахкотіло навколо його, та він не пізнав, і в ньому горіло воно, та не брав він до серця цього!
ISA|43|1|А тепер отак каже Господь, що створив тебе, Якове, і тебе вформував, о Ізраїлю: Не бійся, бо Я тебе викупив, Я покликав ім'я твоє, Мій ти!
ISA|43|2|Коли переходитимеш через води, Я буду з тобою, а через річки не затоплять тебе, коли будеш огонь переходити, не попечешся, і не буде палити тебе його полум'я.
ISA|43|3|Бо Я Господь, Бог твій, Святий Ізраїлів, твій Спаситель! Дав Я на викуп за тебе Єгипта, Етіопію й Севу замість тебе.
ISA|43|4|Через те, що ти став дорогий в Моїх очах, шанований став, й Я тебе покохав, то людей замість тебе віддам, а народи за душу твою.
ISA|43|5|Не бійся, бо Я ж із тобою! Зо сходу згромаджу насіння твоє, і з заходу тебе позбираю.
ISA|43|6|Скажу півночі: Дай, а до півдня: Не стримуй! Поприводь ти синів моїх здалека, а дочки мої від окраїн землі,
ISA|43|7|і кожного, хто тільки зветься Іменням Моїм, і кого Я на славу Свою був створив, кого вформував та кого Я вчинив.
ISA|43|8|Приведи ти народа сліпого, хоч очі він має, і глухих, хоч вуха в них є!
ISA|43|9|Нехай разом зберуться всі люди і народи згромадяться: хто поміж ними розкаже про це, і хто розповість про минуле? Нехай дадуть свідків своїх і оправдані будуть, і хай вони чують та скажуть: Це правда!
ISA|43|10|Ви свідки Мої, говорить Господь, та раб Мій, якого Я вибрав, щоб пізнали й Мені ви повірили, та зрозуміли, ще це Я. До Мене не зроблено Бога, і не буде цього по Мені!
ISA|43|11|Я, Я Господь, і крім Мене немає Спасителя!
ISA|43|12|Я розказав, і споміг, і звістив, і Бога чужого немає між вами, ви ж свідки Мої, говорить Господь, а Я Бог!
ISA|43|13|І Я здавна Той Самий, і ніхто не врятує з Моєї руки, як що Я вчиню, то хто це перемінить?
ISA|43|14|Так говорить Господь, ваш Відкупитель, Святий Ізраїлів: Ради вас Я послав у Вавилон, і зганяю усіх втікачів, а халдеїв кораблі їх утіхи.
ISA|43|15|Я Господь, ваш Святий, Творець Ізраїля, Цар ваш!
ISA|43|16|Так говорить Господь, що дорогу на морі дає, а стежку в могутній воді,
ISA|43|17|що випровадив колесницю й коня, військо та силу, що разом лягли і не встали, зотліли, як льон, та погасли...
ISA|43|18|Не згадуйте вже про минуле, і про давнє не думайте!
ISA|43|19|Ось зроблю Я нове, тепер виросте. Чи ж про це ви не знаєте? Теж зроблю Я дорогу в степу, а в пустині річки.
ISA|43|20|Буде славити Мене польова звірина, шакали та струсі, бо воду Я дам на степу, а в пустині річки, щоб напувати народ Мій, вибранця Мого.
ISA|43|21|Цей народ Я Собі вформував, він буде звіщати про славу Мою.
ISA|43|22|Та Мене ти не кликав, о Якове, не змагався за Мене, Ізраїлю.
ISA|43|23|Ти Мені не приводив ягнят цілопалень своїх, і своїми жертвами не шанував ти Мене... Я тебе не силував, щоб приносити жертву хлібну, і кадилом не мучив тебе.
ISA|43|24|Очерету запашного не купував ти за срібло Мені, і не напував ти Мене лоєм жертов своїх, тільки своїми гріхами Мене ти турбував та своїми провинами мучив Мене!...
ISA|43|25|Я, Я є Той, Хто стирає провини твої ради Себе, а гріхів твоїх не пам'ятає!
ISA|43|26|Пригадай ти Мені і судімося разом, розкажи ти Мені, щоб тобі оправдатись!
ISA|43|27|Твій батько був перший згрішив, і відпали від Мене твої посередники,
ISA|43|28|тому Я позбавив священства священиків, і Якова дав на прокляття, і на зневагу Ізраїля!
ISA|44|1|А тепер ось послухай, о Якове, рабе Мій, та Ізраїлю, якого Я вибрав.
ISA|44|2|Так говорить Господь, що тебе учинив і тебе вформував від утроби, і тобі помагає: Не бійся, рабе Мій, Якове, і Єшуруне, якого Я вибрав!
ISA|44|3|Бо виллю Я воду на спрагнене, а текучі потоки на суходіл, виллю Духа Свого на насіння твоє, а благословення Моє на нащадків твоїх,
ISA|44|4|і будуть вони виростати, немов між травою, немов ті тополі при водних потоках!
ISA|44|5|Цей буде казати: Я Господній, а той зватиметься йменням Якова, інший напише своєю рукою: для Господа я, і буде зватися йменням Ізраїля.
ISA|44|6|Так говорить Господь, Цар Ізраїлів та Викупитель його, Господь Саваот: Я перший, і Я останній, і Бога нема, окрім Мене!
ISA|44|7|І хто зветься, як Я? Хай розкаже про те, й хай звістить те Мені з того часу, коли Я заклав у давнині народ, і хай нам розкаже майбутнє й прийдешнє.
ISA|44|8|Не бійтеся та не лякайтесь! Хіба здавна Я не розповів був тобі й не звістив? А ви свідки Мої! Чи є Бог, окрім Мене? І Скелі немає, не знаю ні жодної!
ISA|44|9|Всі, що роблять бовванів, марнота вони, і їхні улюбленці не помагають, а свідками того самі: не бачать вони та не знають, щоб застидатись!
ISA|44|10|Хто бога зробив та ідола вилив, що він не помагає?
ISA|44|11|Тож друзі його посоромлені будуть усі, майстрі ж вони тільки з людей. Хай вони всі зберуться та стануть: вони полякаються та посоромляться разом!
ISA|44|12|Коваль тне з заліза сокиру, і в горючім вугіллі працює, і формує божка молотками та робить його своїм сильним раменом, а при тім той голодний й безсилий, не п'є води й мучиться...
ISA|44|13|А тесля витягує шнура, визначує штифтом його, того ідола, гемблями робить його та окреслює циркулем це, і робить його на подобу людини, як розкішний зразок чоловіка, щоб у домі поставити.
ISA|44|14|Настинає кедрин він собі, і візьме граба й дуба, і міцне собі викохає між лісними деревами, ясен посадить, а дощик вирощує.
ISA|44|15|І стане людині оце все на паливо, і візьме частину із того й зогріється, теж підпалить в печі й спече хліб. Також виробить бога й йому поклоняється, ідолом зробить його, і перед ним на коліна впадає.
ISA|44|16|Половину його він попалить в огні, на половині його варить м'ясо та їсть, печеню пече й насичається, також гріється та приговорює: Як добре, нагрівся, відчув я огонь...
ISA|44|17|А останок його він за бога вчинив, за боввана свого, перед ним на коліна впадає та кланяється, йому молиться й каже: Рятуй же мене, бо ти бог мій!
ISA|44|18|Не знають і не розуміють вони, бо їхні очі зажмурені, щоб не побачити, і стверділи їхні серця, щоб не розуміти!
ISA|44|19|І не покладе він до серця свого, і немає знання ані розуму, щоб проказати: Половину його попалив я в огні, і на вугіллі його я пік хліб, смажив м'ясо та їв. А решту його за огиду вчиню, буду кланятися дерев'яній колоді?
ISA|44|20|Він годується попелом! Звело його серце обманене, і він не врятує своєї душі, та не скаже: Хіба не брехня у правиці моїй?
ISA|44|21|Пам'ятай про це, Якове та Ізраїлю, бо ти раб Мій! Я тебе вформував був для Себе рабом, Мій Ізраїлю, ти не будеш забутий у Мене!
ISA|44|22|Провини твої постирав Я, мов хмару, і немов мряку гріхи твої, навернися ж до Мене, тебе бо Я викупив!
ISA|44|23|Радійте, небеса, бо Господь це зробив; викликуйте радісно, глибини землі; втішайтеся співом, о гори та лісе, та в нім всяке дерево, бо Господь викупив Якова, і прославивсь в Ізраїлі!
ISA|44|24|Так говорить Господь, твій Відкупитель, та Той, що тебе вформував від утроби: Я, Господь, Той, Хто чинить усе: Розтягнув Я Сам небо та землю втвердив, хто при тім був зо Мною?
ISA|44|25|Хто ознаки ламає брехливим, і робить безглуздими чарівників, Хто з нічим мудреців відсилає, і їхні знання обертає в нерозум,
ISA|44|26|Хто сповнює слово Свого раба, і виконує раду Своїх посланців, Хто Єрусалимові каже: Ти будеш заселений! а юдейським містам: Забудовані будете ви, а руїни його відбудую!
ISA|44|27|Хто глибіні проказує: Висохни, а річки твої Я повисушую,
ISA|44|28|Хто до Кіра говорить: Мій пастирю, і всяке Моє пожадання він виконає та Єрусалимові скаже: Збудований будеш! а храмові: Будеш закладений!
ISA|45|1|Так говорить Господь до Свого помазанця Кіра: Я міцно тримаю тебе за правицю, щоб перед обличчям твоїм повалити народи, і з стегон царів розв'яжу пояси, щоб відчинити двері перед тобою, а брами не будуть замикані.
ISA|45|2|Я перед тобою піду й повирівнюю висунене, двері мідні зламаю і порозбиваю залізні засуви.
ISA|45|3|І дам тобі скарби, що в темряві, та багатства заховані, щоб пізнав ти, що Я то Господь, Який кличе тебе за йменням твоїм, Бог Ізраїлів,
ISA|45|4|ради раба Мого Якова й ради вибранця Мого Ізраїля, і кличу тебе твоїм іменням, тебе називаю, хоч ти не знаєш Мене.
ISA|45|5|Я Господь, і нема вже нікого, нема іншого Бога, крім Мене. Я тебе підперізую, хоч ти не знаєш Мене,
ISA|45|6|щоб дізналися зо сходу сонця й з заходу, що крім Мене немає нічого; Я Господь, і нема вже нікого,
ISA|45|7|Я, що світло формую та темність творю, чиню мир і недолю творю, Я Господь, Який робить це все!
ISA|45|8|Спустіть росу згори, небеса, а із хмар хай спливе справедливість! Хай земля відкривається, і хай породить спасіння та правду, хай разом ростуть! Я, Господь, це вчинив!
ISA|45|9|Горе тому, хто з Творцем своїм свариться, черепок із земних черепків! Чи глина повість ганчареві своєму: Що робиш? а діло його: Ти без рук!
ISA|45|10|Горе тому, хто патякає батькові: Пощо ти плодиш? а жінці: Пощо ти родиш?
ISA|45|11|Так говорить Господь, Святий Ізраїлів, і Той, Хто його вформував: Питайте Мене про майбутнє, а долю синів Моїх й чин Моїх рук позоставте Мені!
ISA|45|12|Я землю вчинив і створив людину на ній, небеса Я руками Своїми простяг і про їхні зорі звелів.
ISA|45|13|Я збудив його в правді, і зрівняю йому всі дороги. Він місто Моє побудує і відпустить вигнанців Моїх не за викуп і не за дарунка, говорить Господь Саваот.
ISA|45|14|Так говорить Господь: Праця Єгипту й торгівля Етіопії та високі севаїтяни перейдуть до тебе та будуть твої. Підуть вони за тобою, у кайданах перейдуть, і будуть вклонятись тобі та благати тебе: Тільки в тебе є Бог, і нема більш, нема іншого Бога!
ISA|45|15|Справді Ти Бог таємничий, Бог Ізраїлів, Спаситель!
ISA|45|16|Всі вони засоромляться й зніяковіють, майстрі ідолів підуть у соромі разом,
ISA|45|17|Ізраїль же буде спасений від Господа вічним спасінням: не будете ви засоромлені ані знеславлені аж на вічні віки!
ISA|45|18|Бо так промовляє Господь, Творець неба. Він той Бог, що землю вформував та її вчинив, і міцно поставив її; не як порожнечу її створив, на проживання на ній Він її вформував. Я Господь, і нема більше іншого Бога!
ISA|45|19|Я не говорив в укритті, на темному місці землі. Я не говорив до насіння Якова: Шукаєте дармо Мене! Я Господь, говорю справедливість, звіщаю правдиве!
ISA|45|20|Зберіться й прийдіть, наблизьтеся разом, урятовані всі із поганів! Не знає нічого, хто дерево носить, боввана свого, та що молиться богові, який не поможе.
ISA|45|21|Розкажіть та наблизьте, і хай разом нарадяться: Хто розповів це віддавна, із давніх часів це звістив? Чи ж не Я, ваш Господь? Бож немає вже Бога, крім Мене, окрім Мене нема Бога праведного та Спасителя!
ISA|45|22|Зверніться до Мене й спасетесь, всі кінці землі, бо Я Бог, і нема більше іншого Бога!
ISA|45|23|Я Собою Самим присягав, справедливість із уст Моїх вийшла, те слово, яке не повернеться: усяке коліно вклонятися буде Мені, усякий язик присягне
ISA|45|24|й Мені скаже: Тільки в Господі правда та сила! Прийдуть до Нього та засоромляться всі, що на Нього запалюються.
ISA|45|25|Через Господа усправедливляться, і буде прославлене всяке насіння Ізраїля!
ISA|46|1|Бел упав на коліна, зігнувся Нево, стали ідоли їхні для звірини й худоби. Те, що колись ви носили, накладене, мов той тягар на худобу помучену.
ISA|46|2|Зігнулися й разом упали вони на коліна; не могли врятувати тягара, і самі до полону пішли...
ISA|46|3|Почуйте Мене, доме Яковів, та ввесь залишку дому Ізраїлевого, яких від живота Я підняв, носив від утроби,
ISA|46|4|і Я буду Той Самий до старости вашої, і до сивини вас носитиму, Я вчинив, і Я буду носити, й Я двигатиму й порятую!
ISA|46|5|До кого Мене ви вподобите та прирівняєте, до кого подібним Мене ви учините, щоб схожому бути?
ISA|46|6|Ті, що золото сиплють з киси, срібло ж важать вагою, винаймлюють золотаря, щоб із того їм бога зробив, і перед ним вони падають та поклоняються,
ISA|46|7|носять його на плечі, підіймають його, і ставлять його на місці його. І стоїть, і з місця свого він не рухається; коли ж хто до нього кричить, то він не відповість, і не врятує його від недолі.
ISA|46|8|Пам'ятайте про це та змужнійте, візьміть це на розум, провинники!
ISA|46|9|Пам'ятайте про давнє, відвічне, бо Я Бог, і немає більш Бога, й нікого, як Я,
ISA|46|10|що звіщаю кінець від початку, і наперед що не сталося ще, і що говорю: Мій замір відбудеться, і всяке жадання Своє Я вчиню,
ISA|46|11|що хижого птаха зо сходу прикликую, з краю далекого мужа Своєї поради! Так, Я сказав те й спроваджу, що Я задумав був теє зроблю!
ISA|46|12|Почуйте Мене, твердосерді, далекі від справедливости!
ISA|46|13|Я Свою справедливість наблизив, вона недалеко, а спасіння Моє не припізниться, і дам на Сіоні спасіння, дам Ізраїлеві Свою велич!
ISA|47|1|Зійди й сядь у порох, о діво, дочко Вавилону! Сядь на землю, без трону, о дочко халдеїв! Бо кликати більше не будуть на тебе: тендитна та випещена!
ISA|47|2|Візьми жорна й муки намели, намітку свою відхили, закачай но подолка та стегна відкрий, і бреди через ріки,
ISA|47|3|і буде твій сором відкритий, і стид твій покажеться! Я помсту вчиню, і не буду щадити людини!
ISA|47|4|Наш Відкупитель, Господь Саваот Йому Ймення, Святий Ізраїлів.
ISA|47|5|Сиди мовчки й ввійди до темноти, о дочко халдеїв, бо кликати більше не будуть тебе: Пані царств!
ISA|47|6|Розлютився Я на народ Свій, збезчестив спадщину Своєю, та й віддав їх у руку твою. Ти не виявила милосердя до них: ти над старцем учинила ярмо своє дуже тяжким,
ISA|47|7|та й сказала: Навіки я панею буду! І до серця собі не взяла тих речей, не подумала про свій кінець...
ISA|47|8|А тепер це послухай, розпещена, що безпечно сидиш, що говориш у серці своїм: Я, і більше ніхто! Не буду сидіти вдовою, і не знатиму страти дітей!
ISA|47|9|Та прийдуть на тебе несподівано те й те в один день, страта дітей та вдівство, вони в повній мірі на тебе спадуть при усій многоті твоїх чарів, при силі великій твоїх заклинань!...
ISA|47|10|Ти ж бо надію складала на злобу свою, говорила: Ніхто не побачить мене! Звела тебе мудрість твоя та знання твоє, і сказала ти в серці своїм: Я, і більше ніхто!
ISA|47|11|І прийде на тебе лихе, що відворожити його ти не зможеш, і на тебе нещастя впаде, що не зможеш його окупити, і прийде на тебе раптовно спустошення, про яке ти не знаєш...
ISA|47|12|Ставай же з своїми закляттями та з безліччю чарів своїх, якими ти мучилася від юнацтва свого, може зможеш ти допомогти, може ти настрахаєш!
ISA|47|13|Змучилась ти від великої кількости рад своїх, хай же стануть і хай допоможуть тобі ті, хто небо розрізує, хто до зір придивляється, хто провіщує кожного місяця, що має на тебе прийти!
ISA|47|14|Ось стали вони, мов солома: огонь їх попалить, не врятують своєї душі з руки полум'я, це не жар, щоб погріти себе, ані полум'я, щоб сидіти біля нього...
ISA|47|15|Такими тобі стануть ті, що співпрацювала ти з ними, ворожбити твої від юнацтва твого, кожен буде блудити на свій бік, немає нікого, хто б тебе врятував!
ISA|48|1|Послухайте це, доме Яковів, що зветесь іменням Ізраїлевим, і що вийшли із Юдиних вод, що клянетеся Йменням Господнім та Бога Ізраїля згадуєте, хоч не в правді та не в справедливості!
ISA|48|2|Бо від міста святого вони прозиваються та на Бога Ізраїлевого спираються, Йому Ймення Господь Саваот!
ISA|48|3|Я віддавна звіщав про минуле, із уст Моїх вийшло воно й розповів Я про нього, раптовно зробив, і прийшло.
ISA|48|4|Тому, що Я знав, що впертий ти є, твоя ж шия то м'язи залізні, а чоло твоє мідяне,
ISA|48|5|то звіщав Я віддавна тобі, іще поки прийшло, розповів Я тобі, щоб ти не говорив: Мій божок це зробив, а про це наказав мій бовван та мій ідол.
ISA|48|6|Ти чув, переглянь усе це; і ви хіба не визнаєте цього? Тепер розповів Я тобі новини й таємниці, яких ти не знав.
ISA|48|7|Тепер вони створені, а не віддавна, а перед цим днем ти не чув був про них, щоб не сказати: Оце я їх знав.
ISA|48|8|Та не чув ти й не знав, і віддавна ти не відкривав свого вуха, бо Я знав, що напевно ти зрадиш, і звано тебе від утроби: перевертень.
ISA|48|9|Ради Ймення Свого Я спиняю Свій гнів, і ради слави Своєї Я стримуюся проти тебе, щоб не знищити тебе.
ISA|48|10|Оце перетопив Я тебе, але не як те срібло, у горні недолі тебе дослідив.
ISA|48|11|Ради Себе, ради Себе роблю, бо як буде збезчещене Ймення Моє? А іншому слави Своєї не дам.
ISA|48|12|Почуй Мене, Якове та Ізраїлю, Мій покликаний: Це Я, Я перший, також Я останній!
ISA|48|13|Теж рука Моя землю заклала, і небо напнула правиця Моя, Я закличу до них і вони стануть разом.
ISA|48|14|Зберіться ви всі та й послухайте: Хто серед вас розповів був про те? Кого Господь любить, вчинить волю Його в Вавилоні, рамено ж Його на халдеях.
ISA|48|15|Я, Я говорив і покликав його, спровадив його, і він на дорозі своїй буде мати поводження.
ISA|48|16|Наблизьтесь до Мене, послухайте це: Споконвіку Я не говорив потаємно; від часу, як діялось це, Я був там. А тепер послав Мене Господь Бог та Його Дух.
ISA|48|17|Так говорить Господь, твій Відкупитель, Святий Ізраїлів: Я Господь, Бог твій, що навчає тебе про корисне, що провадить тебе по дорозі, якою ти маєш ходити.
ISA|48|18|О, коли б ти прислухувався до Моїх заповідей, то був би твій спокій, як річка, а твоя справедливість, немов морські хвилі!
ISA|48|19|А насіння твого було б, як піску, а нащадків твого живота немов зернят його, і витяте й вигублене не було б твоє ймення із-перед обличчя Мого!
ISA|48|20|Вирушіть із Вавилону, втечіть від халдеїв, радісним співом звістіть, оце розголосіть, аж до краю землі рознесіть це, скажіть: Господь викупив раба Свого Якова!
ISA|48|21|І спраги не знали вони на пустинях, якими провадив Він їх: воду з скелі пустив їм, Він скелю розбив і вода потекла!
ISA|48|22|Для безбожних спокою немає, говорить Господь.
ISA|49|1|Почуйте Мене, острови, і народи здалека, вважайте: Господь із утроби покликав Мене, Моє Ймення згадав з нутра неньки Моєї.
ISA|49|2|І Мої уста вчинив Він, як той гострий меч, заховав Мене в тіні Своєї руки, і Мене вчинив за добірну стрілу, в Своїм сагайдаці заховав Він Мене.
ISA|49|3|І до Мене прорік: Ти раб Мій, Ізраїлю, Яким Я прославлюсь!
ISA|49|4|І Я відповів: Надаремно трудивсь Я, на порожнечу й марноту зужив Свою силу: Справді ж з Господом право Моє, і нагорода Моя з Моїм Богом.
ISA|49|5|Тепер же промовив Господь, що Мене вформував Собі від живота за раба, щоб навернути Собі Якова, і щоб Ізраїль для Нього був зібраний. І був Я шанований в очах Господніх, а Мій Бог стався міццю Моєю.
ISA|49|6|І Він сказав: Того мало, щоб був Ти Мені за раба, щоб відновити племена Якова, щоб вернути врятованих Ізраїля, але Я вчиню Тебе світлом народів, щоб був Ти спасінням Моїм аж до краю землі!
ISA|49|7|Так говорить Господь, Відкупитель Ізраїлів, Святий його, до погордженого на душі, до обридженого від людей, до раба тих володарів: Побачать царі, і князі повстають, і поклоняться ради Господа, що вірний, ради Святого Ізраїлевого, що вибрав Тебе.
ISA|49|8|Так говорить Господь: За часу вподобання Я відповів Тобі, в день спасіння Тобі допоміг, і стерегтиму Тебе, і дам Я Тебе заповітом народові, щоб край обновити, щоб поділити спадки спустошені,
ISA|49|9|щоб в'язням сказати: Виходьте, а тим, хто в темноті: З'явіться! При дорогах вони будуть пастися, і по всіх лисих горбовинах їхні пасовиська.
ISA|49|10|Не будуть голодні вони, ані спрагнені, і не вдарить їх спека, ні сонце, бо Той, Хто їх милує, їх попровадить і до водних джерел поведе їх.
ISA|49|11|І вчиню Я всі гори Свої за дорогу, і підіймуться биті шляхи Мої.
ISA|49|12|Ось ці здалека прийдуть, а ці ось із півночі й з заходу, а ці з краю Сінім.
ISA|49|13|Радійте, небеса, звеселися ти, земле, ви ж, гори, втішайтеся співом, бо Господь звеселив Свій народ, і змилувався над Своїми убогими!
ISA|49|14|І сказав був Сіон: Господь кинув мене, і Господь мій про мене забув...
ISA|49|15|Чи ж жінка забуде своє немовля, щоб не пожаліти їй сина утроби своєї? Та коли б вони позабували, то Я не забуду про тебе!
ISA|49|16|Отож на долонях Своїх тебе вирізьбив Я, твої мури позавсіди передо Мною.
ISA|49|17|Синове твої поспішаться до тебе, а ті, хто руйнує тебе й ті, хто нищить тебе, повідходять від тебе.
ISA|49|18|Здійми свої очі навколо й побач: всі вони позбиралися й йдуть ось до тебе! Як живий Я, говорить Господь: усіх їх, як оздобу, зодягнеш, та підв'яжешся ними, немов наречена.
ISA|49|19|Бо руїни твої та пустині твої, і зруйнований край твій тепер справді стануть тісними для мешканців, і будуть віддалені ті, хто тебе руйнував.
ISA|49|20|Іще до вух твоїх скажуть синове сирітства твого: Тісне мені місце оце, посунься для мене, й я сяду!
ISA|49|21|І ти скажеш у серці своїм: Хто мені їх зродив, як була осирочена я та самітна, була вигнана та заблудила? І хто виховав їх? Я зосталась сама, а ці, звідки вони?
ISA|49|22|Так сказав Господь Бог: Ось Я підійму Свою руку до людів, і піднесу до народів прапора Свого, і позносять синів твоїх в пазусі, а дочок твоїх поприносять на плечах.
ISA|49|23|І будуть царі за твоїх вихователів, а їхні цариці за няньок твоїх. Лицем до землі вони будуть вклонятись тобі та лизатимуть пил твоїх ніг, і ти пізнаєш, що Я то Господь, що не посоромляться ті, хто на Мене надіється!
ISA|49|24|Чи ж від сильного буде віднята здобич, і чи награбоване гвалтівником урятоване буде?
ISA|49|25|Бо Господь каже так: Полонені відібрані будуть від сильного, і врятована буде здобич насильника, і Я стану на прю із твоїми суперечниками, синів же твоїх Я спасу.
ISA|49|26|І Я змушу твоїх гнобителів їсти тіло своє, і вони повпиваються власною кров'ю, немов би вином молодим... І пізнає тоді кожне тіло, що Я то Господь, твій Спаситель та твій Відкупитель, Потужний Яковів!
ISA|50|1|Так говорить Господь: Де вашої матері лист розводовий, з яким Я її відпустив? Або хто є з Моїх боргувальників, якому Я вас був продав? Тож за ваші провини ви продані, і за ваші гріхи ваша мати відпущена.
ISA|50|2|Чому то нікого немає, коли Я приходжу, і не відповідає ніхто, коли кличу? Чи рука Моя справді короткою стала, щоб викупляти, і хіба рятувати нема в Мені сили? Таж докором Своїм Я висушую море, обертаю ріки в пустиню, їхня риба гниє без води й умирає із прагнення!
ISA|50|3|Небеса зодягаю Я в темряву, і покриттям їхнім верету чиню.
ISA|50|4|Господь Бог Мені дав мову вправну, щоб уміти зміцнити словом змученого, Він щоранку пробуджує, збуджує вухо Мені, щоб слухати, мов учні.
ISA|50|5|Господь Бог відкрив вухо Мені, й Я не став неслухняним, назад не відступив.
ISA|50|6|Підставив Я спину Свою тим, хто б'є, а щоки Свої щипачам, обличчя Свого не сховав від ганьби й плювання.
ISA|50|7|Але Господь Бог допоможе Мені, тому не соромлюся Я, тому Я зробив був обличчя Своє, немов кремінь, і знаю, що не буду застиджений Я.
ISA|50|8|Близько Той, Хто Мене всправедливлює, хто ж стане зо Мною на прю? Станьмо разом, хто Мій супротивник? Хай до Мене підійде!
ISA|50|9|Отож, Господь Бог допоможе Мені, хто ж отой, що признає Мене винуватим?
ISA|50|10|Хто між вами лякається Господа і голос Його Отрока слухає? Хто ходить у темряві, світла ж немає йому, хай надіється він на Господнє Ім'я, і хай на Бога свого опирається!
ISA|50|11|Тож усі, що огонь ви запалюєте, що огненними стрілами ви поузброювані, ходіть у жарі свого огню та в стрілах огненних, які розпалили! З Моєї руки оце станеться вам, і ви будете в муках лежати!
ISA|51|1|Почуйте Мене, хто женеться за правдою, хто пошукує Господа! Погляньте на скелю, з якої ви витесані, і на каменоломню, з якої ви видовбані.
ISA|51|2|Гляньте на Авраама, батька свого, та на Сарру, що вас породила, бо тільки одного його Я покликав, але благословив був його та розмножив його.
ISA|51|3|Бо Сіона Господь потішає, всі руїни його потішає, й обертає пустині його на Еден, його ж степ на Господній садок! Пробуватимуть в ньому утіха та радість, хвала й пісноспіви.
ISA|51|4|Послухай Мене, Мій народе, і візьми до вух, ти племено Моє, бо вийде від Мене Закон, а Своє правосуддя поставлю за світло народам!
ISA|51|5|Близька правда Моя: вийде спасіння Моє, а рамена Мої будуть суд видавати народам. Острови будуть мати надію на Мене і сподівання свої покладуть на рамено Моє.
ISA|51|6|Здійміть свої очі до неба, і погляньте на землю додолу! Бо небо, як дим, продереться, а земля розпадеться, мов одіж, мешканці ж її, як та воша, погинуть, спасіння ж Моє буде вічне, а правда Моя не зламається!
ISA|51|7|Почуйте Мене, знавці правди, народе, що в серці його Мій Закон: Не бійтеся людської ганьби та їхніх образ не лякайтесь,
ISA|51|8|бо поточить їх міль, мов одежу, й як вовну, черва їх зжере, а правда Моя буде вічна, і спасіння моє з роду в рід!
ISA|51|9|Збудися, збудись, зодягнися у силу, рамено Господнє! Збудися, як у давнину, як за покоління віків! Хіба це не ти Рагава зрубало, крокодила здіравило?
ISA|51|10|Хіба це не ти море висушило, води безодні великої, що морську глибину вчинило дорогою, щоб викуплені перейшли?
ISA|51|11|Отак визволенці Господні повернуться та до Сіону зо співом увійдуть, і на їхній голові буде радість відвічна, веселість та втіху осягнуть вони, а журба та зідхання втечуть!
ISA|51|12|Я, Я ваш Той Утішитель! Хто ж то ти, що боїшся людини смертельної й людського сина, що до трави він подібний?
ISA|51|13|І ти забуваєш про Господа, що вчинив був тебе, що напнув небеса Він та землю заклав, і завжди щоденно лякаєшся гніву гнобителя, що готовий тебе погубити. Але де той гнобителів гнів?
ISA|51|14|Закутий в кайдани небавом розв'язаний буде, і не помре він у ямі, і не забракне йому його хліба.
ISA|51|15|Бо Я Господь, Бог твій, що збурює море, й ревуть його хвілі, Господь Саваот Йому Ймення!
ISA|51|16|І кладу Я слова Свої в уста твої та ховаю тебе в тіні рук Своїх, щоб небо напнути та землю закласти, і сказати Сіонові: Ти Мій народ!
ISA|51|17|Збудися, збудися, устань, дочко Єрусалиму, що з руки із Господньої випила ти келіх гніву Його, чашу-келіха одуру випила, вицідила...
ISA|51|18|Зо всіх тих синів, що вона породила, нікого нема, хто б провадив її; зо всіх тих синів, яких виховала, нікого нема, хто б підтримав її...
ISA|51|19|Ці дві речі спіткали тебе, але хто пожаліє тебе? Руїна й недоля, і голод та меч, хто розважить тебе?
ISA|51|20|Синове твої повмлівали, лежали на розі всіх вулиць, мов олень у тенетах, повні гніву Господнього, крику Бога твого...
ISA|51|21|Тому то послухай оцього, убога й сп'яніла, але не з вина:
ISA|51|22|Так говорить Господь твій, Господь і твій Бог, що на прю за народ Свій стає: Ось келіха одуру Я забираю з твоєї руки, чашу-келіха гніву Мого, більше пити його вже не будеш!
ISA|51|23|І дам Я його в руку тих, що гнобили тебе, що вони до твоєї душі говорили: Схились, і по тобі ми перейдемо! І поклала ти спину свою, немов землю, й як вулицю для перехожих...
ISA|52|1|Збудися, збудись, зодягнися, Сіоне, у силу свою, зодягнися у щати пишноти своєї, о Єрусалиме, о місто святе, бо вже необрізаний та занечищений більше не ввійде до тебе!
ISA|52|2|Обтруси з себе порох, устань та сідай, Єрусалиме! Розв'яжи пута шиї своєї, о бранко, о дочко Сіону!
ISA|52|3|Бо Господь каже так: Задармо були ви попродані, тому будете викуплені не за срібло.
ISA|52|4|Бо так Господь Бог промовляє: До Єгипту зійшов був народ Мій впочатку, щоб мешкати там, а Ашшур за ніщо його тиснув.
ISA|52|5|А тепер що Мені тут, говорить Господь, коли взятий даремно народ Мій? Шаліють володарі їхні, говорить Господь, і постійно ввесь день Моє Ймення зневажене...
ISA|52|6|Тому Моє Ймення пізнає народ Мій, тому того дня він пізнає, що Я то Отой, що говорить: Ось Я!
ISA|52|7|Які гарні на горах ноги благовісника, що звіщає про мир, що добро провіщає, що спасіння звіщає, що говорить Сіонові: Царює твій Бог!
ISA|52|8|Слухай, твої сторожі зняли голос, укупі співають, бо бачать вони око-в-око, коли до Сіону Господь повертається.
ISA|52|9|Радійте, співайте сумісно, о єрусалимські руїни, бо народа Свого Господь звеселив, викупив Єрусалима!
ISA|52|10|Господь обнажив на очах усіх народів святеє рамено Своє, і спасіння від нашого Бога побачать всі кінці землі!
ISA|52|11|Уступіться, вступіться та вийдіть ізвідти, нечистого не доторкайтеся, вийдіть з середини його, очистьтеся ви, що носите посуд Господній!
ISA|52|12|Бо не в поспіху вийдете і не навтеки ви підете, бо піде Господь перед вами, за вами ж Ізраїлів Бог.
ISA|52|13|Ось стане розумне робити Мій Отрок, підійметься й буде повищений, і височенним Він стане!
ISA|52|14|Як багато-хто Ним дивувались, такий то був змінений образ Його, що й не був людиною, а вигляд Його, що й не був сином людським!
ISA|52|15|так Він здивує численних народів, царі свої уста замкнуть перед Ним, бо побачать, про що не говорено їм, і зрозуміють, чого не чували вони!...
ISA|53|1|Хто нашій спасенній тій звістці повірив, і над ким відкривалось рамено Господнє?
ISA|53|2|Бо Він виріс перед Ним, мов галузка, і мов корінь з сухої землі, не мав Він принади й не мав пишноти; і ми Його бачили, та краси не було, щоб Його пожадати!
ISA|53|3|Він погорджений був, Його люди покинули, страдник, знайомий з хоробами, і від Якого обличчя ховали, погорджений, і ми не цінували Його...
ISA|53|4|Направду ж Він немочі наші узяв і наші болі поніс, а ми уважали Його за пораненого, ніби Бог Його вдарив поразами й мучив...
ISA|53|5|А Він був ранений за наші гріхи, за наші провини Він мучений був, кара на Ньому була за наш мир, Його ж ранами нас уздоровлено!
ISA|53|6|Усі ми блудили, немов ті овечки, розпорошились кожен на власну дорогу, і на Нього Господь поклав гріх усіх нас!
ISA|53|7|Він гноблений був та понижуваний, але уст Своїх не відкривав. Як ягня був проваджений Він на заколення, й як овечка перед стрижіями своїми мовчить, так і Він не відкривав Своїх уст...
ISA|53|8|Від утиску й суду Він забраний був, і хто збагне Його рід? Бо з краю живих Він відірваний був, за провини Мого народу на смерть Його дано...
ISA|53|9|І з злочинцями визначили Йому гроба Його, та Його поховали в багатого, хоч провини Він не учинив, і не було в Його устах омани...
ISA|53|10|Та зволив Господь, щоб побити Його, щоб муки завдано Йому. Якщо ж душу Свою покладе Він як жертву за гріх, то побачить насіння, і житиме довгії дні, і замір Господній рукою Його буде мати поводження!
ISA|53|11|Він через муки Своєї душі буде бачити плід, та й насититься. Справедливий, Мій Отрок, оправдає пізнанням Своїм багатьох, і їхні гріхи понесе.
ISA|53|12|Тому то дам уділ Йому між великими, і з потужними буде ділити здобич за те, що на смерть віддав душу Свою, і з злочинцями був порахований, хоч гріх багатьох Сам носив і заступавсь за злочинців!
ISA|54|1|Веселися ж, неплідна, яка не родила, співанням утішайся й радій, що мук породільних не мала, бо в покиненої буде більше синів від синів заміжньої, говорить Господь!
ISA|54|2|Пошир місце намету свого, а завіси наметні помешкань твоїх повитягай, не затримуй! Свої шнури продовж, а кілочки свої позміцняй!
ISA|54|3|Бо праворуч і ліворуч поширишся ти, а насіння твоє одідичать народи, і заселять міста опустошені.
ISA|54|4|Не бійся, бо сорому ти не зазнаєш, і не соромся, бо не будеш застиджена, бо про сором свого юнацтва забудеш, а ганьби удівства свого ти не будеш уже пам'ятати!...
ISA|54|5|Бо Муж твій, Творець твій, Господь Саваот йому Ймення, а твій Викупитель Святий Ізраїлів, Він Богом усієї землі буде званий!
ISA|54|6|Бо Господь був покликав тебе, як покинуту жінку й засмучену духом, й як жінку юнацтва Свого, як була ти відкинена, каже твій Бог.
ISA|54|7|На хвильку малу Я тебе був покинув, але з милосердям великим тебе позбираю.
ISA|54|8|У запалі гніву Я сховав був обличчя Своє на хвилину від тебе, та вічною милістю змилуюся над тобою, каже твій Викупитель, Господь.
ISA|54|9|Бо для Мене оце мов ті Ноєві води: як Я присягнув був, що Ноєві води не прийдуть уже над землею, так Я присягнув, щоб на тебе не гніватися й не картати тебе!
ISA|54|10|Бо зрушаться гори й холми захитаються, та милість Моя не відійде від тебе, і заповіт Мого миру не захитається, каже твій милостивець, Господь.
ISA|54|11|Моя дочко убога та бурею гнана, невтішна, ось каміння твої покладу в малахіті, основи ж твої закладу із сапфірів!
ISA|54|12|І пороблю із рубіну карнізи твої, твої ж брами з каміння карбункула, а всю горожу твою з дорогого каміння.
ISA|54|13|Всі сини твої стануть за учнів Господніх, і спокій глибокий настане синам твоїм!
ISA|54|14|Будеш міцно поставлена правдою, стань далеко від утиску, бо не боятимешся, і від страху, бо до тебе не зблизиться він.
ISA|54|15|Коли хто чіплятися буде до тебе, то це не від Мене, хто чіплятися буде до тебе, той перед тобою впаде.
ISA|54|16|Отож, Я створив коваля, який дме на огонь із вугілля, і вироблює зброю свого ремесла; і вигубника теж Я створив, який нищить ту зброю.
ISA|54|17|Жодна зброя, що зроблена буде на тебе, не матиме успіху, і кожнісінького язика, який стане з тобою до суду, осудиш. Це спадщина Господніх рабів, а їхнє оправдання від Мене, говорить Господь!
ISA|55|1|О, всі спрагнені, йдіть до води, а ви, що не маєте срібла, ідіть, купіть живности, й їжте! І йдіть, без срібла купіть живности, і без платні вина й молока!
ISA|55|2|Нащо будете важити срібло за те, що не хліб, і працю вашу за те, що не ситить? Послухайте пильно Мене, й споживайте добро, і нехай розкошує у наситі ваша душа!
ISA|55|3|Нахиліть своє вухо, й до Мене прийдіть, послухайте, й житиме ваша душа! І з Я вами складу заповіта навіки на незмінні Давидові милості.
ISA|55|4|Отож, Його дав Я за свідка народам, за проводиря та владику народам.
ISA|55|5|Тож покличеш народ, що не знаєш його, і той люд, що не знає тебе, і вони поспішаться до тебе, ради Господа, Бога твого, і ради Святого Ізраїлевого, що прославив тебе.
ISA|55|6|Шукайте Господа, доки можна знайти Його, кличте Його, як Він близько!
ISA|55|7|Хай безбожний покине дорогу свою, а крутій свої задуми, і хай до Господа звернеться, і його Він помилує, і до нашого Бога, бо Він пробачає багато!
ISA|55|8|Бо ваші думки не Мої це думки, а дороги Мої то не ваші дороги, говорить Господь.
ISA|55|9|Бо наскільки небо вище за землю, настільки вищі дороги Мої за ваші дороги, а думки Мої за ваші думки.
ISA|55|10|Бо як дощ чи то сніг сходить з неба й туди не вертається, аж поки землі не напоїть і родючою вчинить її, і насіння дає сівачеві, а хліб їдунові,
ISA|55|11|так буде і Слово Моє, що виходить із уст Моїх: порожнім до Мене воно не вертається, але зробить, що Я пожадав, і буде мати поводження в тому, на що Я його посилав!
ISA|55|12|Бо з радістю вийдете ви, і з миром проваджені будете. Гори й холми будуть тішитися перед вами співанням, і всі польові дерева будуть плескати в долоні.
ISA|55|13|На місце тернини зросте кипарис, а замість кропиви появиться мирт. І стане усе Господеві на славу, на вічну ознаку, яка не понищиться!
ISA|56|1|Так говорить Господь: Бережіть правосуддя й чиніть справедливість, незабаром бо прийде спасіння Моє, і появиться правда Моя.
ISA|56|2|Блаженна людина, що робить таке, і син людський, що міцно тримається цього, що хоронить суботу, щоб її не безчестити, та береже свою руку, щоб жодного зла не вчинити!
ISA|56|3|І нехай не повість чужинець, який прилучився до Господа, кажучи: Насправді мене відділив від народу Свого Господь, і скопець хай не скаже: Таж я сухе дерево!
ISA|56|4|Бо так каже Господь про скопців, що суботи Мої бережуть, і вибирають завгодне Мені, і що тримаються міцно Мого заповіту:
ISA|56|5|Я їм дам у Своїм домі та в мурах Своїх місце і ймення, що краще воно за синів та дочок, Я дам йому вічне ім'я, яке не понищиться!
ISA|56|6|А тих чужинців, що пристали до Господа, щоб служити Йому та любити Господнє Ім'я, щоб бути Йому за рабів, усіх, хто хоронить суботу, щоб її не збезчестити, і тих, що тримаються міцно Мого заповіту,
ISA|56|7|їх спроваджу на гору святую Мою та потішу їх в домі молитви Моєї! Цілопалення їхні та їхні жертви будуть Мені до вподоби на Моїм жертівнику, бо Мій дім буде названий домом молитви для всіх народів!
ISA|56|8|Слово Господа Бога, що збирає вигнанців Ізраїля: Я ще позбираю до нього, до його зібраних!
ISA|56|9|Польова вся звірино, прибудьте спожити, також лісова вся звірино!
ISA|56|10|Його вартівники всі сліпі, не знають нічого, всі вони пси німі, які гавкати не можуть, мрійники, лежні, що люблять дрімати!
ISA|56|11|І це пси ненажери, що не знають насичення, і це пастирі ті, що не вміють уважати: усі вони ходять своєю дорогою, кожен з свого кінця до своєї здобичі...
ISA|56|12|Прийдіть но, говорять, візьму я вина, та напою п'янкого нажлуктимось, і буде і цей день, і завтрішній день далеко щедріший!...
ISA|57|1|Праведний умирає, і немає нікого, хто б узяв це до серця, і мужі побожні беруться зо світу, і немає такого, хто б те зрозумів, що від зла забирається праведний з світу!
ISA|57|2|Він відходить із миром; на ложах своїх спочивають, хто ходить прямою дорогою.
ISA|57|3|Та наблизьтесь сюди, ви сини чарівниці, насіння чужоложникове та блудниці,
ISA|57|4|над ким розкошуєте ви, над ким розкриваєте рота, висовуєте язика? Хіба ви не діти переступу, насіння брехні,
ISA|57|5|ви, що палитесь пристрастю серед дубів, під деревом кожним зеленим, що дітей над потоками ріжете, під скельними щілинами?
ISA|57|6|У гладеньких каміннях потоку твій уділ, вони, вони доля твоя! І їм ти лила жертву литу, хлібну жертву приносила! Чи цим Я заспокоєний буду?
ISA|57|7|На горі на високій та висуненій ти поставила ложе своє, і туди ти приходиш приносити жертви.
ISA|57|8|І ти за дверима й одвірком кладеш свого пам'ятника культового, бо ти відступила від Мене, обнажаєшся й входиш, поширюєш ложе своє, і складаєш умову собі з одним з тих, що з ними ти любиш лежати, де місце нагледиш.
ISA|57|9|І ти до Молоха з оливою ходиш, і намножуєш масті свої; і посилаєш далеко своїх посланців, і знижаєшся аж до шеолу.
ISA|57|10|Ти змучувалась на численних дорогах своїх, але не казала: Зрікаюсь! Знайшла ти оживлення сили своєї, тому не ослабла.
ISA|57|11|І за ким побивалася ти та лякалась, що невірною стала й Мене не згадала, не клала на серці своєму? Хіба не тому, що мовчав Я від віку, то ти не боїшся Мене?
ISA|57|12|Я виявлю про справедливість твою та про вчинки твої, та вони не поможуть тобі!
ISA|57|13|Як ти будеш кричати, нехай порятує тебе твоя зграя божків. Але вітер усіх їх розвіє, схопить подих; хто ж на Мене надіється, землю вспадкує й гору святую Мою одідичить!
ISA|57|14|І Він каже: Будуйте дорогу, будуйте дорогу, почистьте дорогу, заберіть перешкоди з дороги народу Мого!
ISA|57|15|Бо так промовляє Високий і Піднесений, повіки Живущий, і Святий Його Ймення: Пробуваю Я на Височині та в святині, і з зламаним та з упокореним, щоб оживляти духа скромних, і щоб оживляти серця згноблених!
ISA|57|16|Бож не вічно Я буду судитись, і не завжди Я гніватись буду, бо дух з-від обличчя Мого зомлів би, та й душі, які Я вчинив.
ISA|57|17|Я гнівався був за гріх користолюбства його, та й уразив його, заховав Я обличчя Своє й лютував, та пішов він, відступний, дорогою серця свого.
ISA|57|18|Я бачив дороги його, і вздоровлю його, і його поведу й дам потіху для нього й для тих, що сумують із ним.
ISA|57|19|Створю Я плід уст: Спокій, спокій далекому та близькому! говорить Господь, і вздоровлю його.
ISA|57|20|А ті несправедливі як море розбурхане, коли бути спокійним не може воно, і коли води його багно й мул викидають.
ISA|57|21|Для безбожних спокою немає, говорить Господь!
ISA|58|1|Кричи на все горло, не стримуйсь, свій голос повищ, мов у сурму, й об'яви ти народові Моєму про їхній переступ, а домові Якова їхні гріхи!
ISA|58|2|Вони бо щоденно шукають Мене та жадають пізнати дороги Мої, мов народ той, що праведне чинить, і права свого Бога не кидає. Питаються в Мене вони про права справедливости, жадають наближення Бога:
ISA|58|3|Нащо ми постимо, коли Ти не бачиш, мучимо душу свою, Ти ж не знаєш того? Отак, у день посту свого ви чините волю свою, і всіх ваших робітників тиснете!
ISA|58|4|Тож на сварку та заколот постите ви, та щоб кулаком бити нахабно... Тепер ви не постите так, щоб ваш голос почутий був на височині!
ISA|58|5|Хіба ж оце піст, що Я вибрав його, той день, коли морить людина душу свою, свою голову гне, як та очеретина, і стелить верету та попіл? Чи ж оце називаєш ти постом та днем уподоби для Господа?
ISA|58|6|Чи ж ось це не той піст, що Я вибрав його: розв'язати кайдани безбожности, пута ярма розв'язати й пустити на волю утиснених, і всяке ярмо розірвати?
ISA|58|7|Чи ж не це, щоб вламати голодному хліба свого, а вбогих бурлаків до дому впровадити? Що як побачиш нагого, щоб вкрити його, і не сховатися від свого рідного?
ISA|58|8|Засяє тоді, мов досвітня зоря, твоє світло, і хутко шкірою рана твоя заросте, і твоя справедливість ходитиме перед тобою, а слава Господня сторожею задньою!
ISA|58|9|Тоді кликати будеш і Господь відповість, будеш кликати і Він скаже: Ось Я! Якщо віддалиш з-поміж себе ярмо, не будеш підносити пальця й казати лихого,
ISA|58|10|і будеш давати голодному хліб свій, і знедолену душу наситиш, тоді то засвітить у темряві світло твоє, і твоя темрява ніби як полудень стане,
ISA|58|11|і буде Господь тебе завжди провадити, і душу твою нагодує в посуху, кості твої позміцняє, і ти станеш, немов той напоєний сад, і мов джерело те, що води його не всихають!
ISA|58|12|І руїни відвічні сини твої позабудовують, поставиш основи довічні, і будуть тебе називати: Замуровник пролому, направник шляхів для поселення!
ISA|58|13|Якщо ради суботи ти стримаєш ногу свою, щоб не чинити своїх забаганок у день Мій святий, і будеш звати суботу приємністю, днем Господнім святим та шанованим, і її пошануєш, не підеш своїми дорогами, діла свого не шукатимеш та не будеш казати даремні слова,
ISA|58|14|тоді в Господі розкошувати ти будеш, і Він посадовить тебе на висотах землі, та зробить, що будеш ти споживати спадщину Якова, батька твого, бо уста Господні сказали оце!
ISA|59|1|Ото ж бо, Господня рука не скоротшала, щоб не помагати, і Його вухо не стало тяжким, щоб не чути,
ISA|59|2|бо то тільки переступи ваші відділювали вас від вашого Бога, і ваші провини ховали обличчя Його від вас, щоб Він не почув,
ISA|59|3|бо ваші долоні заплямлені кров'ю, ваші ж пальці беззаконням, уста ваші говорять неправду, язик ваш белькоче лихе!
ISA|59|4|Немає нікого, хто б кликав на суд, і нікого нема, хто судився б поправді, кожен надію кладе не марноту й говорить неправду, вагітніє бідою й породжує злочин!
ISA|59|5|Висиджують яйця гадючі та тчуть павутиння: хто з'їсть з їхніх яєць, помирає, а з розбитого гадина вийде...
ISA|59|6|Нитки їхні не стануть одежею, і виробами своїми вони не покриються: їхні діла діла кривди, і в їхніх руках чин насильства...
ISA|59|7|Їхні ноги біжать на лихе, і спішать проливати невинну кров, їхні думки думки кривдні, руїна й погибіль на їхніх дорогах!
ISA|59|8|Дороги спокою не знають, і правосуддя немає на їхніх стежках, вони покрутили собі свої стежки, і кожен, хто нею ступає, не знає спокою.
ISA|59|9|Тому віддалилося право від нас, і не сягає до нас справедливість! чекаємо світла, та ось темнота, чекаємо сяйва та й у темнощах ходимо!
ISA|59|10|Ми мацаємо, мов невидющі, за стіну, навпомацки ходимо, мов ті безокі; спотикаємося ми опівдні, немов би смерком, між здоровими ми, як померлі!...
ISA|59|11|Усі ми ревемо, як ведмеді, і мов голуби ті постійно воркочемо, чекаємо права й немає, спасіння й від нас віддалилось воно...
ISA|59|12|Бо помножились наші переступи перед Тобою, і свідкують на нас гріхи наші, бо з нами переступи наші, а наші провини ми знаємо їх!
ISA|59|13|Ми зраджували й говорили неправду на Господа, і повідступали від нашого Бога, казали про утиск та відступ, вагітніли й видумували з свого серця слова неправдиві...
ISA|59|14|І правосуддя назад відступилося, а справедливість здалека стоїть, бо на майдані спіткнулася істина, правда ж не може прийти,
ISA|59|15|і істина зникла, а той, хто від злого відходить, грабований... І це бачить Господь, і лихе в Його очах, що права нема!
ISA|59|16|І Він бачив, що немає нікого, і дивувавсь, що немає заступника... Та рамено Його Йому допомогло, і Його справедливість підперла Його,
ISA|59|17|і Він зодягнув справедливість, як панцер, а шолома спасіння на Свою голову, і зодягнув шати помсти, як одяг, і покрився горливістю, мов би плащем!
ISA|59|18|Надолужить Він гнівом Своїм ворогам згідно з учинками їхніми, Своїм супротивним заплатою, островам надолужить заплату.
ISA|59|19|І будуть боятися Ймення Господнього з заходу, а слави Його зо схід сонця, бо прийде, як річка рвучка, вітер Господній її пожене,
ISA|59|20|і прийде Викупитель Сіонові й тим, хто вернувся із прогріху в Якові, каже Господь.
ISA|59|21|А Я ось із ними умова Моя, говорить Господь: Мій Дух, який на тобі, та слова Мої, що поклав Я до уст твоїх, не уступлять вони з твоїх уст, і з уст нащадків твоїх, і з уст нащадків потомства твого, говорить Господь, відтепер й аж навіки!
ISA|60|1|Уставай, світися, Єрусалиме, бо прийшло твоє світло, а слава Господня над тобою засяла!
ISA|60|2|Бо темрява землю вкриває, а морок народи, та сяє Господь над тобою, і слава Його над тобою з'являється!
ISA|60|3|І підуть народи за світлом твоїм, а царі за ясністю сяйва твого.
ISA|60|4|Здійми свої очі навколо й побач: усі вони зібрані, і до тебе ідуть; сини твої йдуть іздалека, а дочок твоїх на руках он несуть!
ISA|60|5|Побачиш тоді і роз'яснишся ти, сполохнеться й поширшає серце твоє, бо звернеться морське багатство до тебе, і прийде до тебе багатство народів!
ISA|60|6|Безліч верблюдів закриє тебе, молоді ті верблюди з Мідіяну й Ефи, усі вони прийдуть із Шеви, носитимуть золото й ладан та хвали Господні звіщатимуть.
ISA|60|7|Всі отари кедарські зберуться до тебе, барани невайотські послужать тобі, вони підуть усі на Мій вівтар, як жертва приємна, і Я прославлю дім слави Своєї!
ISA|60|8|Хто вони, що летять, як та хмара, і немов голуби до своїх голубників?
ISA|60|9|Бо до Мене збираються мореплавці, і найперше пливуть кораблі із Таршішу, щоб привести синів твоїх здалека, з ними їхнє срібло та їхнє золото для Імені Господа, Бога твого, і для Святого Ізраїля, Він бо прославив тебе.
ISA|60|10|І мури твої побудують чужинці, а їхні царі тобі будуть служити, бо в запалі гніву Свого Я був уразив тебе, а в Своїм уподобанні змилуюся над тобою!
ISA|60|11|І будуть постійно відкритими брами твої, ані вдень, ні вночі не замкнуться вони, щоб приносити до тебе багатство народів, і їхні царі щоб були припроваджені.
ISA|60|12|Бо погинуть народ та те царство, що не схочуть служити тобі, і ці народи понищені будуть зовсім!
ISA|60|13|Слава ліванська прибуде до тебе, кипарис, сосна й бук будуть разом, щоб приоздобити місце святині Моєї, і місце ніг Своїх Я пошаную.
ISA|60|14|І зігнуті прийдуть до тебе сини твоїх кривдників, і кланятись будуть до стіп твоїх ніг усі ненависники, і тебе будуть кликати: Місто Господнє, Сіон Святого Ізраїлевого!
ISA|60|15|За те, що була ти покинута та осоружна, о дочко Сіону, і через тебе ніхто не ходив, то вчиню тебе славою вічною, радістю з роду в рід!
ISA|60|16|І будеш ти ссати молоко із народів, і груди царів будеш ссати, і пізнаєш, що Я то Господь, твій Спаситель, а твій Викупитель Потужний Яковів!
ISA|60|17|Замість міді впроваджу Я золото, і замість заліза впроваджу срібло, і замість дерева мідь, а замість каміння залізо, і дозором твоїм зроблю мир, твоїми ж начальниками справедливість!
ISA|60|18|В твоїм краї не буде вже чуте насилля, руїна й спустошення в межах твоїх, і назвеш свої мури спасінням, а брами свої похвалою!
ISA|60|19|Удень сонце не буде тобі вже за світло, і не буде світити тобі місяць за сяйво, бо буде тобі вічним світлом Господь, а твій Бог за окрасу твою!
ISA|60|20|Не зайде вже сонце твоє, і місяць твій вже не сховається, бо буде тобі вічним світлом Господь, і дні жалоби твоєї покінчаться!
ISA|60|21|А народ твій усі справедливі вони, землю вспадкують навіки, парость Моїх саджанців, чин Моїх рук на прославлення!
ISA|60|22|Цей малий стане тисячею, і наймолодший народом міцним! Я, Господь, цього часу оце приспішу!
ISA|61|1|Дух Господа Бога на мені, бо Господь помазав Мене благовістити сумирним, послав Мене перев'язати зламаних серцем, полоненим звіщати свободу, а в'язням відчинити в'язницю,
ISA|61|2|щоб проголосити рік уподобання Господу, та день помсти для нашого Бога, щоб потішити всіх, хто в жалобі,
ISA|61|3|щоб радість вчинити сіонським жалобникам, щоб замість попелу дати їм оздобу, оливу радости замість жалоби, одежу хвали замість темного духа! І будуть їх звати дубами праведности, саджанцями Господніми, щоб прославивсь Господь!
ISA|61|4|І вони забудують руїни відвічні, відбудують спустошення давні і відновлять міста поруйновані, з роду в рід попустошені.
ISA|61|5|І встануть чужинці та й пастимуть ваші отари, і сини чужинця будуть вам рільниками та вам винарями!
ISA|61|6|І будуть вас кликати: Господні, священики будуть казати на вас: слуги нашого Бога! Ви будете їсти багатство народів, і їхньою славою будете славитись.
ISA|61|7|За ваш сором подвійний і за ганьбу та смуток, ваш уділ, тому то посядуть вони в своїм краї подвійне, радість вічна їм буде!
ISA|61|8|Бо Господь Я, і правосуддя кохаю, і ненавиджу розбій та кривду, і дам їм заплату за чин їхній поправді, і з ними складу заповіта довічного!
ISA|61|9|І буде насіння їхнє знане між людами, і між народами їхні нащадки, усі, хто бачити їх буде, пізнають їх, що вони те насіння, яке благословив був Господь!
ISA|61|10|Я радісно буду втішатися Господом, нехай звеселиться душа моя Богом моїм, бо Він зодягнув мене в шату спасіння, і в одежу праведности мене вбрав, немов молодому, поклав Він на мене вінця, і мов молоду, приоздобив красою мене!
ISA|61|11|Бо так як земля та виводить рослинність свою, й як насіння своє родить сад, так Господь Бог учинить, що виросте правда й хвала перед усіма народами!
ISA|62|1|Не буду мовчати я ради Сіону, і ради Єрусалиму не буду спокійний, аж поки не вийде, як сяйво, його справедливість, а спасіння його як горючий світильник!
ISA|62|2|І побачать народи твою справедливість, а славу твою всі царі, і йменням новим будуть звати тебе, що уста Господні докладно означать його.
ISA|62|3|І ти станеш короною слави в Господній руці й діядемою царства в долоні Бога свого!
ISA|62|4|Вже не скажуть на тебе покинута, а на край твій не будуть казати вже пустиня, бо тебе будуть кликати в ній моя втіха, а край твій заміжня, бо Господь пожадає тебе, і твій край буде взятий за жінку!
ISA|62|5|Як юнак бере панну за жінку, так з тобою одружиться Сам Будівничий, і як тішиться той молодий нареченою, так радітиме Бог твій тобою!
ISA|62|6|На мурах твоїх, Єрусалиме, Я поставив сторожу, ніколи не буде мовчати вона цілий день та всю ніч. Ви, хто пригадує Господа, не замовкніть,
ISA|62|7|і перед Ним не вмовкайте, аж поки не зміцнить, і аж поки не вчинить Він Єрусалима за славу Свою на землі!
ISA|62|8|Господь присягнув був Своєю правицею й потужним раменом Своїм: Направду, не дам уже збіжжя твого ворогам твоїм, і пити не будуть чужинці твого виноградного соку, що ти працював біля нього!
ISA|62|9|Бо ті, хто збирає його, будуть їсти його та й хвалитимуть Господа, і ті, хто громадить його, будуть пити його на подвір'ях святині Моєї!
ISA|62|10|Проходьте, проходьте ви брамами, чистьте дорогу народові! Будуйте дорогу, будуйте дорогу, дорогу ту биту, очистьте від каменя, підійміть над народами прапора!
ISA|62|11|Ось звіщає Господь аж до краю землі: Розкажіте сіонській дочці: Ось приходить Спасіння твоє, ось із Ним нагорода Його, і заплата Його перед Ним!
ISA|62|12|І будуть їх звати народом святим, викупленцями Господа, а на тебе закличуть жадана, незалишене місто!
ISA|63|1|Хто це гряде із Едому, у шатах червоних із Боцри? Хто Той пишний в убранні Своїм, що в величі сили Своєї врочисто гряде? Це Я, що говорить у правді, що владний спасати!
ISA|63|2|Чого то червона одежа Твоя, а шати Твої як у того, хто топче в чавилі?
ISA|63|3|Сам один Я чавило топтав, і не було із народів зо Мною нікого! І Я топтав їх у гніві Своїм, і чавив їх у люті Своїй, і бризкав їх сік на одежу Мою, і Я поплямив всі шати Свої...
ISA|63|4|Бо день помсти у серці Моїм, і надійшов рік Мого викуплення!
ISA|63|5|Я дививсь, але помічника не було, і дивувавсь, бо підпори Мені бракувало, та рамено Моє Мені допомогло, а Мій гнів він підтримав Мене!
ISA|63|6|І топтав Я народи у гніві Своїм, і ламав їх у люті Своїй, і вилив на землю їхню кров!
ISA|63|7|Буду згадувати ласки Господні, Господні хвали за все те, що вчинив нам Господь, за велике добро те для дому Ізраїля, що вчинив Він для них у Своїм милосерді, і в ласці великій Своїй!
ISA|63|8|І сказав: Вони справді народ Мій, сини, що неправди не кажуть, і став Він для них за Спасителя.
ISA|63|9|В усякому утиску їхньому тісно було і Йому, і Ангол обличчя Його їх спасав. Любов'ю Своєю й Своїм милосердям Він викупив їх, і їх підніс і носив їх усі дні в давнину.
ISA|63|10|Та стали вони неслухняними й Духа Святого Його засмутили, і Він обернувся на ворога їм, Він Сам воював проти них...
ISA|63|11|Тоді то народ Його згадає дні давні, Мойсея: Де Той, що їх вивів із моря із пастирем отари Своєї? Де Той, що в нього поклав Свого Духа Святого?
ISA|63|12|Що Він по правиці Мойсея провадив рамено величчя Свого, що Він перед ними розділював воду, щоб зробити Собі вічне Ім'я?
ISA|63|13|Що провадив безоднями їх, як коня на пустині, і вони не спіткнулись?
ISA|63|14|Як сходить у долину худоба, так їх Дух Господній водив до спочинку, так і Ти вів народ Свій, щоб зробити Собі славне Ім'я!
ISA|63|15|Поглянь із небес і побач із мешкання святині Своєї та слави Своєї: Де горливість Твоя та Твої могутні чини? Де велике число милосердя Твого та ласки Твоєї, що супроти мене затрималися?
ISA|63|16|Тільки Ти наш Отець, бо Авраам нас не знає, а Ізраїль нас не пізнає! Ти, Господи, Отець наш, від віку Ім'я Твоє: наш Викупитель!
ISA|63|17|Нащо, Господи, Ти попустив, що ми блудимо з доріг Твоїх, нащо робиш твердим наше серце, щоб ми не боялись Тебе? Вернися ради рабів Своїх, ради племен спадку Свого!
ISA|63|18|Спадщину займав час короткий святий Твій народ, противники наші святиню Твою потоптали!
ISA|63|19|Ми стали такими, немов би відвіку Ти не панував був над нами, немов би не кликалося Твоє Ймення над нами!
ISA|64|1|О, коли б небеса Ти роздер і зійшов, перед обличчям Твоїм розтопилися б гори,
ISA|64|2|як хворост горить від огню, як кипить та вода на огні, отак щоб Ім'я Твоє стало відоме Твоїм ворогам, щоб перед обличчям Твоїм затремтіли народи!
ISA|64|3|Коли Ти чинив страшні речі, ми їх не чекали, коли б Ти зійшов, то перед обличчям Твоїм розтопилися б гори!
ISA|64|4|І відвіку не чули, до ушей не доходило, око не бачило Бога, крім Тебе, Який би зробив так тому, хто надію на Нього кладе!
ISA|64|5|Ти стрічаєш того, хто радіє та праведність чинить, отих, що вони на дорогах Твоїх пам'ятають про Тебе. Та розгнівався Ти, бо ми в тому згрішили навіки та несправедливими стали!
ISA|64|6|І стали всі ми, як нечистий, а вся праведність наша немов поплямована місячним одіж, і в'янемо всі ми, мов листя, а наша провина, як вітер, несе нас...
ISA|64|7|І немає нікого, хто кликав би Ймення Твоє, хто збудився б триматися міцно за Тебе, бо від нас заховав Ти обличчя Своє й через нашу вину Ти покинув нас нидіти...
ISA|64|8|Тепер же, о Господи, Ти наш Отець, ми глина, а Ти наш ганчар, і ми всі чин Твоєї руки!
ISA|64|9|Не гнівайся, Господи, сильно, і не пам'ятай повсякчасно провини! Тож споглянь, ми народ Твій усі!
ISA|64|10|Святі міста Твої стали пустинею, Сіон став пустелею, степом став Єрусалим...
ISA|64|11|Дім святощі нашої й нашої слави, в якім батьки наші хвалили Тебе, погорілищем став, а все наше любе руїною стало...
ISA|64|12|Чи й на це ще Себе будеш стримувати, Господи? Будеш мовчати, й занадто карати нас будеш?
ISA|65|1|Я прихилявся до тих, що Мене не питали, Я знайдений тими, що Мене не шукали. Я казав: Оце Я, оце Я! до народу, що Йменням Моїм не був званий.
ISA|65|2|Я ввесь день простягав Свої руки до люду запеклого, що він, за своїми думками, дорогою ходить недоброю,
ISA|65|3|до народу, що в очі Мене прогнівляє постійно, що жертви приносить в садках та що палить кадило на цеглах,
ISA|65|4|що сидить у гробах та ночує по ямах, їсть свинину, і в їхньому посуді юшка нечиста,
ISA|65|5|що говорить: Спинись, не зближайся до мене, бо святий я для тебе! Оце дим в Моїй ніздрі, огонь, що палає ввесь день!
ISA|65|6|Ось написане перед обличчям Моїм: Я не буду мовчати, але відплачу, і надолужу на їхньому лоні!
ISA|65|7|Укупі переступи ваші й переступи ваших батьків, говорить Господь, що кадили на горах і на взгір'ях Мене зневажали, і заплату їм виміряю Я найперше до їхнього лоня!...
ISA|65|8|Так говорить Господь: Коли в гроні знаходиться сік виноградний, і хтось скаже: Не псуй ти його, бо благословення у ньому, отак Я зроблю ради рабів Своїх, щоб усього не нищити!
ISA|65|9|І насіння Я виведу з Якова, а з Юди спадкоємця гір Моїх, і вибранці Мої одідичать її, і раби Мої житимуть там.
ISA|65|10|І стане Шарон пасовиськом отари, а долина Ахор за ліжницю худоби великої, для народу Мого, що шукали Мене.
ISA|65|11|А ви, що Господа кидаєте, забуваєте гору святу Мою, що ставите Ґаду трапезу, а для Мені виповнюєте жертву литу,
ISA|65|12|то вас відраховую Я для меча, й на коліна впадете ви всі на заріз, бо кликав Я вас, та ви відповіді не дали, говорив був, але ви не чули й робили лихе в Моїх очах, і чого не хотів, вибирали собі!...
ISA|65|13|Тому Господь Бог каже так: Ось будуть раби Мої їсти, а ви будете голодувати, ось будуть раби Мої пити, а ви будете спрагнені, ось будуть раби Мої радіти, а ви посоромлені будете...
ISA|65|14|Ось раби Мої будуть співати від радости серця свого, ви ж кричатимете від сердечного болю, і від скрушення духа заводити будете...
ISA|65|15|І ви своє ймення дасте на прокляття вибранцям Моїм, і Господь Бог тебе вб'є, а рабам Своїм дасть інше ймення,
ISA|65|16|так що хто на землі благословлений буде, буде поблагословлений він вірним Богом, а хто на землі присягає, вірним Богом присягне, бо забудуться утиски давні і заховані будуть вони від очей Моїх!
ISA|65|17|Бо ось Я створю нове небо та землю нову, і не згадаються речі колишні, і не прийдуть на серце!
ISA|65|18|Тож навіки радійте та тіштеся тим, що творю Я, бо ось Я створю Єрусалима на радість, а народа його на веселість!
ISA|65|19|І буду Я Єрусалимом радіти, і втішатися буду народом Своїм, і не почується в ньому вже голос плачу й голос зойку!
ISA|65|20|З цього часу не буде вже юного днями й старого, який своїх днів не поповнить, бо сторокий помре як юнак, а грішник і в віці ста літ буде проклятий!
ISA|65|21|І доми побудують, і мешкати будуть, і засадять вони виноградники, і будуть їхній плід споживати.
ISA|65|22|Не будуть вони будувати, щоб інший сидів, не будуть садити, щоб інший спожив, дні бо народу Мого як дні дерева, і вибранці Мої зуживатимуть чин Своїх рук!
ISA|65|23|Не будуть вони працювати надармо, і не будуть родити на страх, вони бо насіння, благословлене Господом, і нащадки їхні з ними.
ISA|65|24|І станеться, поки покличуть, то Я відповім, вони будуть іще говорити, а Я вже почую!
ISA|65|25|Вовк та вівця будуть пастися разом, і лев буде їсти солому, немов та худоба, а гадові хлібом його буде порох!... Вони не чинитимуть зла й вигубляти не будуть на всій святій Моїй горі, говорить Господь.
ISA|66|1|Так говорить Господь: Небеса Мій престол, а земля то підніжок для ніг Моїх: який же то храм, що для Мене збудуєте ви, і яке ото місце Його відпочинку?
ISA|66|2|Таж усе це створила рука Моя, і так все це сталось, говорить Господь! І при тому дивлюсь Я на вбогого та на розбитого духом, і на тремтячого над Моїм словом.
ISA|66|3|Інакше хто ріже вола одночасно вбиває людину, приносить у жертву ягня переломлює шию собаці, дарунка приносить вживає свинячої крови, складає з кадила частину пригадувальну, одночасно божка благословить... Отак як дороги свої вони повибирали, і до гидот тих своїх уподобання чує душа їхня,
ISA|66|4|так виберу й Я їх на зведення, і предмета їхнього страху на них наведу, за те, що Я кликав і ніхто відповіді не давав, говорив Я й не чули вони, та чинили лихе в Моїх очах, і вибрали те, чого Я не жадав!...
ISA|66|5|Послухайте слова Господнього ті, що на слово Його тремтите: Кажуть ваші брати, що ненавидять вас, що вас ради Ймення Мого виганяють: Хай прославлений буде Господь, і ми вашу радість побачимо! Та будуть вони посоромлені!
ISA|66|6|Голос гомону з міста, голос із храму, це голос Господа, що заплату дає для Своїх ворогів!
ISA|66|7|Поки зазнала дрижання породу, вона породила, і поки прийшов її біль, то сина легенько вона привела...
ISA|66|8|Хто таке коли чув, і хто бачив таке? Чи зроджена буде земля в один день, чи народжений буде народ за одним разом? Бо як тільки зазнала Сіонська дочка породові дрижання, то синів своїх вже породила...
ISA|66|9|Чи Я допроваджу до породу, і не вчиню, щоб вона породила? говорить Господь. Чи Я, що чиню, щоб родила, і стримаю? каже твій Бог.
ISA|66|10|Радійте із Єрусалимом і тіштеся всі ним, хто його покохав! Втішайтесь ним радістю всі, що з-за нього в жалобі були!
ISA|66|11|Щоб ви ссали й наситилися з перс потіхи його, щоб ви ссали та розкошували із перс його слави!
ISA|66|12|Бо Господь каже так: Ось керую до нього Я мир, немов річку, і славу народів, немов той потік заливний: і ви будете ссати, і на руках вас носитимуть, і бавитимуть на колінах!
ISA|66|13|Як когось його ненька втішає, так вас Я потішу, і ви втішені будете Єрусалимом.
ISA|66|14|І побачите це, й серце ваше радітиме, й як трава молода, розцвітуть ваші кості! І в рабах Його пізнана буде Господня рука, і буде Він гніватися на Своїх ворогів.
ISA|66|15|Бо ось прийде Господь ув огні, а Його колесниці мов буря, щоб відплатити жаром гніву Свого, а погрози Свої полум'яним огнем!
ISA|66|16|Бо огнем та мечем Своїм буде судитись Господь з кожним тілом, і буде багато побитих від Господа...
ISA|66|17|А ті, хто освячується й очищає себе у поганських садках, один по одному, всередині, їдять м'ясо свиняче й гидоти та мишу, вони разом загинуть, говорить Господь!...
ISA|66|18|І Я знаю їхні вчинки та їхні думки, і прийду, щоб зібрати всі народи й язики, і прийдуть вони й Мою славу побачать!
ISA|66|19|І знака на них покладу, і пошлю урятованих з них до народів, у Таршіш, Пул, і Лул, в Мешех і Кос, у Тувал та Яван, в острови предалекі, що звістки про Мене не чули й не бачили слави Моєї, і звістять мою славу вони між народами!
ISA|66|20|І вони приведуть усіх ваших братів із народів усіх у дарунок для Господа на конях та на колесницях, і на фурах та мулах, та на верблюдах, на гору святу Мою, до Єрусалиму, говорить Господь, як приносять синове Ізраїлеві дарунка в посудині чистій до дому Господнього.
ISA|66|21|І візьму Я із них за священиків та за Левитів, говорить Господь.
ISA|66|22|Бо як небо нове та нова та земля, що вчиню, стануть перед обличчям Моїм, говорить Господь, так стоятимуть ваші нащадки та ваше ім'я!
ISA|66|23|І станеться, кожного новомісяччя в часі його, і щосуботи за часу її кожне тіло приходитиме, щоб вклонятися перед обличчям Моїм, говорить Господь.
ISA|66|24|І вийдуть вони та й побачать ті трупи людей, що відпали від Мене, бо їхня черва не помре й не погасне огонь їхній, і стануть вони за гидоту для кожного тіла!
