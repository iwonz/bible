DAN|1|1|За третього року царювання Йоякима, Юдиного царя, прийшов Навуходоносор, цар вавилонський, до Єрусалиму, та й обліг його.
DAN|1|2|І дав Господь в його руку Йоякима, Юдиного царя, та частину посуду Божого дому, і він вірправив їх до краю вавилонського, до дому свого бога, а посуд відправив до скарбничного дому свого бога.
DAN|1|3|І сказав цар до Ашпеназа, начальника його евнухів, щоб привести з Ізраїлевих синів, і з царського, і з шляхетського роду,
DAN|1|4|юнаків, що нема в них жодної вади, і вони вродливого вигляду та розумні в усякій мудрості, і здібні до знання, і розуміють науку, і щоб у них була моторність служити в царському палаці, і щоб навчати їх книг та мови халдеїв.
DAN|1|5|І призначив їм цар щоденну поживу, з царської їжі та з вина, що сам його пив, а на їхнє виховання три роки, а по закінченні їх стануть вони перед царським обличчям.
DAN|1|6|І були серед них з Юдиних синів Даниїл, Ананія, Мисаїл та Азарія.
DAN|1|7|А начальник евнухів дав їм інші імена, і дав Даниїлові ім'я Валтасар, а Ананії Шадрах, а Мисаїлові Мешах, а Азарії Авед-Неґо.
DAN|1|8|І поклав Даниїл собі на серце, що він не оскверниться їжею царя та питвом, що той сам його пив, і просив від начальника евнухів, щоб не осквернитися.
DAN|1|9|І дав Бог Даниїлові ласку та милість перед начальником евнухів.
DAN|1|10|І сказав начальник евнухів до Даниїла: Боюсь я свого пана царя, бо він визначив вашу їжу та ваше питво. Бо коли б він побачив ваше обличчя худішим, ніж у тих юнаків, що вашого віку, то ви зробите мою голову винуватою перед царем.
DAN|1|11|І сказав Даниїл до старшого, якого начальник евнухів призначив над Даниїлом, Ананією, Мисаїлом та Азарією:
DAN|1|12|Випробуй но своїх рабів десять день, і нехай дають нам із ярини, і ми будемо їсти, та воду і будемо пити.
DAN|1|13|І нехай з'являться перед тобою наші обличчя та обличчя тих юнаків, що їдять царську їжу, і згідно з тим, що побачиш, зроби зо своїми рабами.
DAN|1|14|І той послухався їх у цьому, і випробовував їх десять день.
DAN|1|15|А по десяти днях їхній вигляд виявився кращим, і вони були здоровіші на тілі, аніж усі ті юнаки, що їли царську їжу.
DAN|1|16|І цей старший відносив їхню їжу та вино їхнього пиття, а давав їм ярину.
DAN|1|17|А ці четверо юнаків, дав їм Бог пізнання та розуміння в кожній книжці та мудрості, а Даниїл розумівся на всякому видінні та снах.
DAN|1|18|А на кінець тих днів, коли цар сказав привести їх, то начальник евнухів привів їх перед обличчя Навуходоносорове.
DAN|1|19|І цар розмовляв з ними, і зо всіх них жоден не був знайдений таким, як Даниїл, Ананія, Мисаїл та Азарія. І вони ставали перед царським обличчям.
DAN|1|20|А всяку справу мудрости та розуму, що шукав від них цар, то він знайшов їх удесятеро мудрішими від усіх чарівників та заклиначів, що були в усьому його царстві.
DAN|1|21|І був Даниїл там аж до першого року царя Кіра.
DAN|2|1|А за другого року Навуходоносорового царювання приснилися Навуходоносорові сни. І занепокоївся дух його, і сон його утік від нього.
DAN|2|2|І сказав цар покликати чарівників та заклиначів, і чаклунів та халдеїв, щоб розповіли цареві його сни. І вони поприходили, і поставали перед царським обличчям.
DAN|2|3|І сказав до них цар: Снився мені сон, і занепокоївся дух мій, щоб пізнати той сон.
DAN|2|4|А халдеї говорили цареві по-арамейському: Царю, живи навіки! Розкажи перше сон своїм рабам, а ми об'явимо розв'язку.
DAN|2|5|Цар відповів та й сказав до халдеїв: Моє слово невідкличне: якщо ви не розповісте мені сна та його розв'язку, будете почетвертовані, а ваші доми обернуться в руїни.
DAN|2|6|А якщо ви розповісте сон та його розв'язку, одержите від мене дари й нагороду та велику честь; тому об'явіть мені сон та його розв'язку.
DAN|2|7|Вони відповіли вдруге та й сказали: Цар перше розкаже сон своїм рабам, а ми об'явимо розв'язку.
DAN|2|8|Цар відповів та й сказав: Я знаю напевно, що ви хочете виграти час, бо бачите, що слово моє невідкличне.
DAN|2|9|Якщо ви не розкажете мені сна, то один у вас задум, бо ви змовилися говорити передо мною лож та неправду, аж поки зміниться час. Тому розкажіть мені сон, і я пізнаю, що ви об'явите мені, і його розв'язку.
DAN|2|10|Халдеї відповіли перед царем та й сказали: Нема на суходолі людини, що могла б об'явити цареву справу, бо жоден великий та панівний цар не питався такої речі від жодного чарівника й заклинача та халдея.
DAN|2|11|А справа, про яку питається цар, тяжка, і немає таких, що об'явили б її перед царем, окрім богів, що не мають своїх мешкань разом із тілом.
DAN|2|12|За це цар розгнівався, та сильно розпінився, і наказав вигубити всіх вавилонських мудреців.
DAN|2|13|І вийшов наказ, і вбивали мудреців, і шукано Даниїла та його товаришів, щоб повбивати.
DAN|2|14|Того часу Даниїл розповів розважно та розумно Арйохові, начальникові царської сторожі, що вийшов був побивати вавилонських мудреців.
DAN|2|15|Він заговорив та й сказав Арйохові, царському владиці: Чому такий жорстокий наказ від царя? Тоді Арйох розповів Даниїлові справу.
DAN|2|16|І Даниїл увійшов, і просив просити від царя, щоб дав йому часу, і він об'явить цареві розв'язку сна.
DAN|2|17|Тоді Даниїл пішов до свого дому, і завідомив про справу товаришів своїх, Ананію, Мисаїла та Азарію,
DAN|2|18|щоб просили милости від Небесного Бога на цю таємницю, щоб не вигубили Даниїла та товаришів його разом з рештою вавилонських мудреців.
DAN|2|19|Тоді Даниїлові відкрита була таємниця в нічному видінні, і Даниїл прославив Небесного Бога.
DAN|2|20|Даниїл заговорив та й сказав: Нехай буде благословенне Боже Ім'я від віку й аж до віку, бо Його мудрість та сила.
DAN|2|21|І Він зміняє часи та пори року, скидає царів і настановляє царів, дає мудрість мудрим, і пізнання розумним.
DAN|2|22|Він відкриває глибоке та сховане, знає те, що в темряві, а світло спочиває з Ним.
DAN|2|23|Тобі, Боже батьків моїх, я дякую та славлю Тебе, що Ти дав мені мудрість та силу, а тепер відкрив мені, що я від Тебе просив, бо Ти відкрив нам справу цареву.
DAN|2|24|Потому Даниїл пішов до Арйоха, якого цар призначив вигубити вавилонських мудреців. Пішов він та й так йому сказав: Не губи вавилонських мудреців! Заведи мене перед царя, і я об'явлю цареві розв'язку сна.
DAN|2|25|Тоді Арйох негайно привів Даниїла перед царя, та й сказав йому так: Знайшов я мужа з синів Юдиного вигнання, що об'явить цареві розв'язку сна.
DAN|2|26|Цар заговорив та й сказав Даниїлові, що йому було ймення Валтасар: Чи ти можеш об'явити мені сон, якого я бачив, та його розв'язку?
DAN|2|27|Даниїл відповів перед царем та й сказав: Таємниці, про яку питається цар, не можуть об'явити цареві ані мудреці, ані заклиначі, ані чарівники, ані віщуни.
DAN|2|28|Але є на небесах Бог, що відкриває таємниці, і Він завідомив царя Навуходоносора про те, що буде в кінці днів. Твій сон та видіння твоєї голови на ложі твоїм оце вони:
DAN|2|29|Тобі царю, приходили на ложе твоє думки твої про те, що буде потім, а Той, Хто відкриває таємницю, показав тобі те, що буде.
DAN|2|30|А мені ця таємниця відкрита не через мудрість, що була б у мені більша від мудрости всіх живих, а тільки на те, щоб об'явити цареві розв'язку, і ти пізнаєш думки свого серця.
DAN|2|31|Ти, царю, бачив, аж ось один великий бовван, бовван цей величезний, а блиск його дуже сильний; він стояв перед тобою, а вигляд його був страшний.
DAN|2|32|Цей бовван такий: голова його з чистого золота, груди його та рамена його зо срібла, нутро його та стегно його з міді,
DAN|2|33|голінки його з заліза, ноги його частинно з заліза, а частинно з глини.
DAN|2|34|Ти бачив, аж ось одірвався камінь сам, не через руки, і вдарив боввана по ногах його, що з заліза та з глини, і розторощив їх.
DAN|2|35|Того часу розторощилося, як одне, залізо, глина, мідь, срібло та золото, і вони стали, немов та полова з току жнив, а вітер їх розвіяв, і не знайшлося по них жодного сліду; а камінь, що вдарив того боввана, став великою горою, і наповнив усю землю.
DAN|2|36|Оце той сон, а його розв'язку зараз скажемо перед царем.
DAN|2|37|Ти, царю, цар над царями, якому Небесний Бог дав царство, владу й міць та славу.
DAN|2|38|І скрізь, де мешкають людські сини, польова звірина та птаство небесне, Він дав їх у твою руку, та вчинив тебе пануючим над усіма ними. Ти голова, що з золота.
DAN|2|39|А по тобі постане інше царство, нижче від тебе, і царство третє, інше, що з міді, яке буде панувати над усією землею.
DAN|2|40|А царство четверте буде сильне, як залізо, бо залізо товче й розбиває все, так і воно стовче й розіб'є, як залізо, що все розбиває.
DAN|2|41|А що ти бачив ноги та пальці частинно з ганчарської глини, частинно з заліза, то це буде поділене царство, і в ньому буде трохи залізної міці, бо ти бачив залізо, змішане з глейкою глиною.
DAN|2|42|А пальці ніг частинно з заліза, а частинно з глини, то й частина царства буде сильна, а частина буде ламлива.
DAN|2|43|А що бачив ти залізо, змішане з глейкою глиною, то вони змішані будуть людським насінням, а не будуть прилягати одне до одного, як залізо не змішується з глиною.
DAN|2|44|А за днів тих царів Небесний Бог поставить царство, що навіки не зруйнується, і те царство не буде віддане іншому народові. Воно потовче й покінчить усі ті царства, а само буде стояти навіки.
DAN|2|45|Бо ти бачив, що з гори відірвався камінь сам, не руками, і потовк залізо, мідь, глину, срібло та золото. Великий Бог об'явив цареві те, що станеться потім. А сон цей певний, і певна його розв'язка!
DAN|2|46|Тоді цар Навуходоносор упав на своє обличчя й поклонився Даниїлові, і наказав приносити йому хлібну жертву та любі пахощі!
DAN|2|47|Цар відповів Даниїлові та й сказав: Направду, що ваш Бог це Бог над богами та Пан над царями, і Він відкриває таємниці, коли міг ти відкрити оцю таємницю!
DAN|2|48|Тоді цар звеличив Даниїла, і дав йому численні дарунки, і вчинив його паном над усім вавилонським краєм, і великим провідником над усіма вавилонськими мудрецями.
DAN|2|49|А Даниїл просив від царя, і він призначив над справами вавилонського краю Шадраха, Мешаха та Авед-Неґо, а Даниїл був при царському дворі.
DAN|3|1|Цар Навуходоносор зробив був золотого боввана, заввишки йому шістдесят ліктів, завширшки йому шість ліктів. Він поставив його в долині Дура в вавилонській окрузі.
DAN|3|2|І цар Навуходоносор послав зібрати сатрапів, заступників, підсатрапів, радників, суддів, вищих урядників та всіх округових володарів, щоб прийшли на посвячення боввана, якого поставив цар Навуходоносор.
DAN|3|3|Того часу зібралися сатрапи, заступники, підсатрапи, радники, скарбники, судді, вищі урядники та всі округові володарі, щоб посвятити боввана, якого поставив цар Навуходоносор, і поставали навпроти боввана, якого поставив Навуходоносор.
DAN|3|4|А оповісник закликав лунким Голосом: До вас говориться, народи, люди та язики!
DAN|3|5|Того часу, коли ви почуєте голос рога, сопілки, гітари, гусел, псалтиря, флейти та всілякого роду музику, падайте й поклоніться золотому бовванові, якого поставив цар Навуходоносор.
DAN|3|6|А той, хто не впаде й не поклониться, тієї хвилі буде вкинений до середини палахкотючої огненної печі.
DAN|3|7|Тому того часу, як усі народи почують голос рога, сопілки, гітари, гусел, псалтиря та всілякого роду музику, попадають всі народи, люди та язики, і поклоняться золотому бовванові, якого поставив цар Навуходоносор.
DAN|3|8|А цього часу наблизилися халдейські мужі, і доносили на юдеїв.
DAN|3|9|Вони заговорили та й сказали цареві Навуходоносорові: Царю, живи навіки!
DAN|3|10|Ти царю, видав наказа, щоб кожен чоловік, хто почує голос рога, сопілки, гітари, гусел, псалтиря й флейти та всілякої музики, упав і поклонився золотому бовванові.
DAN|3|11|А той, хто не впаде й не поклониться, буде вкинений до середини палахкотючої огненної печі.
DAN|3|12|Є юдейські мужі, яких ти призначив над справами вавилонської округи, Шадрах, Мешах та Авед-Неґо, ці мужі не звернули на тебе, царю, уваги: богам твоїм не служать, і золотому бовванові, якого ти поставив, не вклоняються.
DAN|3|13|Тоді Навуходоносор у гніві та в лютості наказав привести Шадраха, Мешаха та Авед-Неґо, і того часу цих людей привели перед царя.
DAN|3|14|Навуходоносор заговорив та й сказав їм: Шадраху, Мешаху та Авед-Неґо, чи це правда, що ви моїм богам не служите, а золотому бовванові, якого я поставив, не вклоняєтеся?
DAN|3|15|Тепер, якщо ви готові, щоб того часу, коли почуєте голос рога, сопілки, гітари, гусел, псалтиря й флейти та всіляких родів музику, попадали й кланялися бовванові, якого я зробив. А якщо ви не поклонитеся, тієї години будете вкинені до середини палахкотючої огненної печі, і хто той Бог, що врятує вас від моїх рук?
DAN|3|16|Шадрах, Мешах та Авед-Неґо відповіли та й сказали цареві Навуходоносорові: Ми не потребуємо відповідати тобі на це слово.
DAN|3|17|Якщо наш Бог, Якому ми служимо, може врятувати нас з палахкотючої огненної печі, то Він урятує й з твоєї руки, о царю!
DAN|3|18|А якщо ні, нехай буде тобі, о царю, знане, що богам твоїм ми не служимо, а золотому бовванові, якого ти поставив, не будемо вклонятися!
DAN|3|19|Тоді Навуходоносор переповнився лютістю, і вигляд його обличчя змінився проти Шадраха, Мешаха та Авед-Неґо. Він відповів, і наказав напалити піч усемеро понад те, як повинно було напалити її.
DAN|3|20|І він наказав хоробрим військовим мужам, що були в його війську, зв'язати Шадраха, Мешаха та Авед-Неґо, щоб укинути до палахкотючої огненної печі.
DAN|3|21|Того часу ці мужі були пов'язані в своїх плащах, у своїх сорочках і в своїх шапках, і в своїх убраннях, і були повкидані до середини палахкотючої огненної печі.
DAN|3|22|А що слово царя було гостре, то піч напалена була надзвичайно сильно, так що тих мужів, що підіймали, щоб укинути Шадраха, Мешаха та Авед-Неґо, забило їх огняне полум'я.
DAN|3|23|А ці три мужі, Шадрах, Мешах та Авед-Неґо, упали до середини палахкотючої огненної печі пов'язані.
DAN|3|24|Тоді цар Навуходоносор здивувався, і поспішно встав, заговорив та й сказав до своїх радників: Чи ж не трьох зв'язаних мужів ми кинули до середини огню? Ті відповіли та й сказали цареві: Певне, царю!
DAN|3|25|Він відповів та й сказав: Таж я бачу чотирьох мужів непов'язаних, що ходять посеред огню, і шкоди їм нема, а вигляд того четвертого подібний до Божого сина!
DAN|3|26|Тоді Навуходоносор наблизився до челюстів палахкотючої огненної печі, заговорив та й сказав: Шадраху, Мешаху та Авед-Неґо, раби Його, Бога Всевишнього, вийдіть і прийдіть! Тоді Шадрах, Мешах та Авед-Неґо вийшли з середини огню.
DAN|3|27|І зібралися сатрапи, заступники, і підсатрапи, і цареві радники, та й побачили тих мужів, що огонь не мав сили над їхнім тілом, і не опалився волос їхньої голови, і їхні плащі не змінилися, і запах огню не ввійшов у них.
DAN|3|28|Навуходоносор заговорив та й сказав: Благословенний Бог Шадраха, Мешаха та Авед-Неґо, що послав Свого Ангола, і врятував Своїх рабів, які надіялися на Нього. І вони не послухалися царського слова, і дали свої тіла на огонь, аби не служити й не кланятися іншому богові, крім Бога свого.
DAN|3|29|А тепер від мене видається наказ, що кожен з народу, люду та язика, який скаже що згірдливе на Бога Шадраха, Мешаха та Авед-Неґо, буде почетвертований, а дім його обернений буде на сміття, бо немає іншого Бога, що міг би так урятувати, як оце.
DAN|3|30|Того часу цар зробив, щоб добре велося Шадрахові, Мешахові та Авед-Неґові в вавилонській окрузі.
DAN|4|1|(3-31) Цар Навуходоносор, до всіх народів, племен та язиків, що мешкають на всій землі: Нехай вам примножиться мир!
DAN|4|2|(3-32) Знаки та чуда, які зробив зо мною Всевишній Бог, уважаю за відповідне об'явити.
DAN|4|3|(3-33) Які великі Його знаки, й які потужні Його чуда! Царство Його царство вічне, а Його панування з покоління в покоління!
DAN|4|4|(4-1) Я, Навуходоносор, був спокійний в своєму домі, і щасливий у палаті своїй.
DAN|4|5|(4-2) Я бачив сон, і він настрашив мене, а думки на моєму ложі та видіння моєї голови налякали мене.
DAN|4|6|(4-3) І був виданий від мене наказ привести перед мене всіх вавилонських мудреців, щоб вони об'явили мені розв'язку сна.
DAN|4|7|(4-4) Того часу поприходили чарівники, заклиначі, халдеї та віщуни, і я розповів перед ними сон, та вони не об'явили мені його розв'язки.
DAN|4|8|(4-5) І аж останній прийшов перед мене Даниїл, якому ім'я Валтасар, як ім'я мого бога, і що в ньому дух Святого Бога. І я розповів йому сон та й сказав:
DAN|4|9|(4-6) Валтасаре, начальнику чарівників, я знаю, що в тобі дух Святого Бога, і всяка таємниця не тяжка тобі. Скажи видіння мого сну, що я бачив, та його розв'язку.
DAN|4|10|(4-7) А видіння моєї голови на моєму ложі такі. Я бачив, аж ось дерево серед землі, а вишина його велика.
DAN|4|11|(4-8) Це дерево стало велике та сильне, і вишина його сягала до Неба, а його обвід до кінця всієї землі.
DAN|4|12|(4-9) Віття його гарне, плід його великий, а в ньому пожива для всіх. Під ним знаходила собі тінь польова звірина, а на його галуззях мешкали птахи небесні, і з нього живилося кожне тіло.
DAN|4|13|(4-10) Бачив я у видіннях своєї голови на моєму ложі, аж ось зійшов з неба Сторож Божий та Святий.
DAN|4|14|(4-11) І він кликнув із силою, і так проказав: Зрубайте це дерево, і повідрубуйте галуззя його, позривайте віття його, і порозсипайте його плід. Нехай розійдеться з-під нього звірина, а птахи з галуззя його!
DAN|4|15|(4-12) Та позоставте в землі пня його кореня, але в путах залізних та мідяних, на зеленій польовій траві. І небесною росою нехай він зрошується, а його частка зо звіриною на польовій траві.
DAN|4|16|(4-13) Його людське серце змінять, і буде дане йому серце звірине, і сім часів перейдуть над ним.
DAN|4|17|(4-14) Через постанову Сторожів Божих це слово, а повідженням Святих ця річ, аж прийде до того, що пізнають живі, що над людським царством панує Всевишній, і кому схоче, дає його, і низького з людей ставить над ним.
DAN|4|18|(4-15) Оцей сон бачив я, цар Навуходоносор, а ти, Валтасаре, скажи його розв'язку, бо всі мудреці мого царства не можуть сказати мені розв'язки, а ти можеш, бо в тобі дух Святого Бога.
DAN|4|19|(4-16) Тоді Даниїл, що ім'я йому Валтасар, остовпів на одну годину, і думки його перестрашили його. Цар заговорив та й сказав: Валтасаре, нехай не страшить тебе цей сон та його розв'язка! Валтасар відповів та й сказав: Мій пане, на ворогів би твоїх цей сон, а його розв'язка на твоїх би неприятелів!
DAN|4|20|(4-17) Дерево, яке ти бачив, що було велике та міцне, і вишина його сягала до неба, а обвід його на всю землю,
DAN|4|21|(4-18) а віття його гарне, і плід його великий, і в ньому пожива для всіх, під ним мешкала польова звірина, а на його галуззях перебували птахи небесні,
DAN|4|22|(4-19) ти, царю, той, що став великий та потужний, і твоя великість побільшилася, і сягнула аж до небес, а панування твоє до кінців землі.
DAN|4|23|(4-20) А що цар бачив Божого Сторожа та Святого, який сходив із небес, і сказав: Зрубайте це дерево, і знищте його, та позоставте в землі пня його кореня, але в путах залізних та мідяних, на зеленій польовій траві; і небесною росою нехай він зрошується, а його частка з польовою звіриною, аж поки перейдуть над ним сім часів,
DAN|4|24|(4-21) то ось розв'язка, царю, і це постанова Всевишнього, що сягає на мого пана царя:
DAN|4|25|(4-22) І тебе виженуть від людей, і з польовою звіриною буде пробування твоє, і дадуть тобі їсти траву, як волам, і з небесної роси тебе зросять, і сім часів перейдуть над тобою, аж поки пізнаєш, що над людським царством панує Всевишній, і дає його тому, кому хоче.
DAN|4|26|(4-23) А що сказали позоставити пня кореня дерева, твоє царство позостанеться тобі, якщо ти пізнаєш, що панує небо.
DAN|4|27|(4-24) Тому, царю, нехай буде до вподоби моя рада тобі, зламай же свої гріхи справедливістю, а свої провини милістю для вбогих, щоб твій мир був довготривалий.
DAN|4|28|(4-25) Усе це сталося над царем Навуходоносором.
DAN|4|29|(4-26) На кінці дванадцяти місяців проходжувався він по царському палацу в Вавилоні.
DAN|4|30|(4-27) Цар заговорив та й сказав: Чи ж це не величний Вавилон, що я збудував його на дім царства міццю потуги своєї та на славу моєї пишноти?
DAN|4|31|(4-28) Ще це слово було в устах царських, коли з неба впав голос: Тобі говорять, царю Навуходоносоре: Оце царство відходить від тебе!
DAN|4|32|(4-29) І від людей тебе відлучать, і з польовою звіриною буде пробування твоє, тобі дадуть на їжу траву, як волам, і сім часів перейдуть над тобою, аж поки не пізнаєш, що над людським царством панує Всевишній, і дає його тому, кому хоче.
DAN|4|33|(4-30) Тієї хвилини виконалося це слово над Навуходоносором, і він був відлучений від людей, і їв траву, як воли, і його тіло зрошувалося з небесної роси, аж його волос став великий, як пір'я орлине, а його пазурі як у птахів.
DAN|4|34|(4-31) А на кінці тих днів я, Навуходоносор, звів свої очі до неба, і мій розум вернувся до мене, й я поблагословив Всевишнього, і вічно Живого хвалив я та славив, що Його панування панування вічне, а царство Його з покоління в покоління.
DAN|4|35|(4-32) А всі мешканці землі пораховані за ніщо, і Він чинить за Своєю Волею серед небесного війська та мешканців землі, і немає нікого, хто спротивився б Його руці та й сказав би Йому: Що Ти робиш?
DAN|4|36|(4-33) Того часу вернувся мій розум до мене, і я вернувся до слави царства свого, і ясність моя вернулася на мене. І шукали мене мої радники та вельможі мої, і над царством своїм я був поставлений знову, і мені була додана дуже велика величність.
DAN|4|37|(4-34) Тепер я, Навуходоносор, хвалю й звеличую та славлю Небесного Царя, що всі чини Його правда, а дорога Його правосуддя, а тих, хто ходить у гордощах, Він може понизити.
DAN|5|1|Цар Валтасар справив велике прийняття для тисячі своїх вельмож, і на очах тієї тисячі пив вино.
DAN|5|2|Коли вино опанувало розум, Валтасар наказав принести золотий та срібний посуд, який виніс був його батько Навуходоносор із храму, що в Єрусалимі, щоб із нього пили цар та вельможі його, його жінки та його наложниці.
DAN|5|3|Тоді принесли золотий посуд, що винесли з храму божого дому, що в Єрусалимі, і пили з них цар та вельможі його, жінки його та його наложниці.
DAN|5|4|Пили вони вино й славили богів золотих та срібних, мідяних, залізних, дерев'яних та камінних.
DAN|5|5|Аж ось тієї хвилини вийшли пальці людської руки, і писали навпроти свічника на вапні стіни царського палацу, і цар бачив зарис руки, що писала.
DAN|5|6|Тоді змінилася ясність царя, і думки його настрашили його, ослабіли суглоби крижів його, і билися коліна його одне об одне.
DAN|5|7|Цар сильно закричав привести заклиначів, халдеїв та віщунів. Цар заговорив та й сказав вавилонським мудрецям: Кожен муж, що прочитає це писання й об'явить мені його розв'язку, той зодягне пурпуру й золотого ланцюга на свою шию, і буде панувати третім у царстві.
DAN|5|8|Тоді поприходили всі царські мудреці, та не могли прочитати писання й об'явити цареві його розв'язку.
DAN|5|9|Тоді цар Валтасар сильно перестрашився, а його ясність змінилася на ньому, і його вельможі були безрадні.
DAN|5|10|На слова царя та вельмож його ввійшла до дому прийняття цариця. Цариця заговорила та й сказала: Царю, живи навіки! Нехай не страшать тебе думки твої, а ясність твоя нехай не міняється!
DAN|5|11|Є в твоєму царстві муж, що в ньому дух святих богів, а за днів твого батька в ньому знаходилась ясність і розум та мудрість, рівна мудрості богів. І цар Навуходоносор, твій батько, настановив його начальником чарівників, заклиначів, халдеїв, віщунів, батько твій цар,
DAN|5|12|бо в ньому, в Даниїлові, якому цар дав ім'я Валтасар, знаходився надмірний дух, і знання та розум розв'язувати сни, і висловлювати загадки та розплутувати вузли. Нехай буде покликаний тепер Даниїл, і нехай він оголосить розв'язку!
DAN|5|13|Того часу Даниїл був приведений перед царя. Цар заговорив та й сказав до Даниїла: Чи ти той Даниїл, що з Юдиних синів вигнання, яких вивів цар, мій батько, з Юдеї?
DAN|5|14|І чув я про тебе, що в тобі дух богів, і що в тобі знаходиться ясність, і розум та надмірна мудрість.
DAN|5|15|А тепер були приведені перед мене мудреці, заклиначі, щоб прочитали оце писання, і розповіли мені його розв'язку, та не могли вони висловити розв'язки цієї речі.
DAN|5|16|А я чув про тебе, що ти можеш розв'язувати недовідоме, і розплутувати вузли. Тож тепер, якщо можеш прочитати це писання, і розповісти мені його розв'язку, то зодягнеш пурпуру, а золотий ланцюг на твою шию, і ти будеш панувати третім у царстві.
DAN|5|17|Тоді Даниїл відповів та й сказав перед царем: Твої дари нехай будуть тобі, а дарунки свої давай іншим. Це писання я прочитаю цареві, і розповім тобі його розв'язку.
DAN|5|18|Ти, царю, Всевишній Бог дав твоєму батькові Навуходоносорові царство, і велич, і славу та пишноту.
DAN|5|19|А через велич, яку Він дав був йому, всі народи, племена та язики тремтіли та лякалися перед ним, бо кого він хотів забивав, а кого хотів лишав при житті, і кого хотів підіймав, а кого хотів понижував.
DAN|5|20|А коли загордилося його серце, а дух його ще більше запишнів, він був скинений з трону свого царства, і його слава була взята від нього.
DAN|5|21|І він був вигнаний з-поміж людських синів, і серце його було зрівняне зо звіриним, а пробування його було з дикими ослами. Годували його травою, як волів, а небесною росою зрошувалося його тіло, аж поки він не пізнав, що в людському царстві панує Всевишній Бог, і Він ставить над ним того, кого хоче.
DAN|5|22|А ти, сину його Валтасаре, не смирив свого серця, хоч усе це знав.
DAN|5|23|І ти піднісся понад Небесного Господа, і посуд храму Його принесли перед тебе, а ти та вельможі твої, жінки твої та наложниці твої пили з них вино, і ти хвалив богів срібних та золотих, мідяних, залізних, дерев'яних та камінних, що не бачать, і не чують та не знають, а Бога, що в руці Його душа твоя й що Його всі дороги твої, ти не прославляв.
DAN|5|24|Того часу від Нього посланий зарис руки, і написане оце писання.
DAN|5|25|А оце писання, що написане: Мене, мене, текел упарсін.
DAN|5|26|Ось розв'язка цієї речі: Мене порахував Бог царство твоє, і покінчив його.
DAN|5|27|Текел ти зважений на вазі, і знайдений легеньким.
DAN|5|28|Перес поділене царство твоє, і віддане мідянам та персам.
DAN|5|29|Тоді наказав Валтасар, і надягли на Даниїла пурпуру, а золотого ланцюга на шию його, і розголосили про нього, що він буде третім пануючим у царстві.
DAN|5|30|Тієї ж ночі був забитий Валтасар, цар халдейський.
DAN|5|31|(6-1) А мідянин Дарій одержав царство в віці шостидесяти й двох років.
DAN|6|1|(6-2) Сподобалося Дарієві, і він поставив над царством сто й двадцять сатрапів, щоб були над усім царством.
DAN|6|2|(6-3) А вище від них три найвищі урядники, що одним із них був Даниїл, яким ці сатрапи здавали звіт, а цар щоб не був пошкодований.
DAN|6|3|(6-4) Тоді цей Даниїл блищав над найвищими урядниками та сатрапами, бо в ньому був високий дух, і цар задумував поставити його над усім царством.
DAN|6|4|(6-5) Тоді найвищі урядники та сатрапи стали шукати причини оскаржити Даниїла в справі царства, але жодної причини чи вади знайти не могли, бо той був вірний, і жодна помилка чи вада не була знайдена на нього.
DAN|6|5|(6-6) Тоді ці люди сказали: Ми не знайдемо на цього Даниїла жодної причини, якщо не знайдемо проти нього в законі його Бога.
DAN|6|6|(6-7) Тоді найвищі урядники та ті сатрапи поспішили до царя, і так йому говорили: Царю Даріє, живи навіки!
DAN|6|7|(6-8) Нарадилися всі найвищі урядники царства, заступники та сатрапи, радники та підсатрапи встановити царську постанову та видати заборону, щоб аж до тридцяти день кожен, хто буде просити яке прохання від якогобудь бога чи людини, крім від тебе, о царю, був укинений до лев'ячої ями.
DAN|6|8|(6-9) Тепер, царю, затверди цю заборону, і напиши це писання, яке не могло б бути змінене за законом мідян та персів, що не міг би бути відмінений.
DAN|6|9|(6-10) Тому цар Дарій написав це писання та заборону.
DAN|6|10|(6-11) А Даниїл, коли довідався, що було написане те писання, пішов до свого дому, а вікна його в його горниці були відчинені навпроти Єрусалиму, і в три усталені порі на день він падав на свої коліна, і молився та славив свого Бога, бо робив так і перед тим.
DAN|6|11|(6-12) Тоді ці мужі поспішили до нього, і знайшли Даниїла, що він просив та благав свого Бога.
DAN|6|12|(6-13) Тоді вони підійшли й розповіли перед царем про царську заборону: Чи ж не написав ти заборони, що кожна людина, яка буде просити аж до тридцяти день від якогобудь бога чи людини, окрім від тебе, царю, буде вкинена до лев'ячої ями? Цар відповів та й сказав: Це слово певне, як право мідян та персів, що не може бути відмінене.
DAN|6|13|(6-14) Тоді вони відповіли та й сказали перед царем: Даниїл, що з вигнання Юдиних синів, не звернув уваги на тебе, о царю, та на заборону, яку написав ти, і в три усталені порі на день приносить свою молитву.
DAN|6|14|(6-15) Тоді цар, як почув це слово, сильно засмутився, і звернув свою думку на Даниїла, щоб його врятувати, і аж до заходу сонця силувався визволити його.
DAN|6|15|(6-16) Того часу ці мужі поспішили до царя, і говорили цареві: Знай, царю, що за правом мідян та персів усяка заборона та постанова, яку цар установить, не може буде змінена.
DAN|6|16|(6-17) Тоді цар звелів, і привели Даниїла, та й кинули до лев'ячої ями. Цар заговорив і сказав Даниїлові: Твій Бог, що ти Йому служиш, Він завжди врятує тебе!
DAN|6|17|(6-18) І принесений був один камінь, і був покладений на отвір ями, а цар запечатав її своєю печаткою та печаткою своїх вельмож, що не буде змінена Даниїлова справа.
DAN|6|18|(6-19) Тоді цар пішов до свого палацу, і провів ніч у пості, і до нього не впроваджено наложниці, а сон його помандрував від нього.
DAN|6|19|(6-20) Того часу цар устав за зірниці на світанку, і в поспіху пішов до лев'ячої ями.
DAN|6|20|(6-21) А як цар наближався до ями, до Даниїла, то кликнув сумним голосом. Цар заговорив та й сказав до Даниїла: Даниїле, рабе Бога Живого, чи твій Бог, Якому ти завжди служиш, міг урятувати тебе від левів?
DAN|6|21|(6-22) Тоді Даниїл заговорив із царем: Царю, навіки живи!
DAN|6|22|(6-23) Мій Бог послав Свого Ангола, і позамикав пащі левів, і вони не пошкодили мені, бо перед Ним знайдено було мене невинним, а також перед тобою, царю, я не зробив шкоди.
DAN|6|23|(6-24) Тоді цар сильно зрадів, і сказав вивести Даниїла з ями. І Даниїл був виведений з ями, і жодної шкоди не знайдено на ньому, бо він вірував у Бога свого.
DAN|6|24|(6-25) І сказав цар, і привели тих мужів, що донесли на Даниїла, і повкидали до лев'ячої ями їх, їхніх дітей та їхніх жінок. І вони не сягнули ще до дна ями, як леви вже похапали їх, і поторощили всі їхні кості.
DAN|6|25|(6-26) Того часу цар Дарій написав до всіх народів, племен та язиків, що мешкали по всій землі: Нехай мир вам примножиться!
DAN|6|26|(6-27) Від мене виданий наказ, щоб у всьому пануванні мого царства тремтіли та боялися перед Даниїловим Богом, бо Він Бог Живий і існує повіки, і царство Його не буде зруйноване, а панування Його аж до кінця.
DAN|6|27|(6-28) Він рятує та визволяє, і чинить знаки та чуда на небі та на землі, Він урятував Даниїла від лев'ячої сили.
DAN|6|28|(6-29) І той Даниїл мав поводження за царювання Дарія та за царювання Кіра перського.
DAN|7|1|За першого року Валтасара, царя вавилонського, бачив Даниїл сон та пророцьке видіння голови своєї на своєму ложі. Того часу записав він сон, сказавши з нього головне.
DAN|7|2|Даниїл заговорив та й сказав: Бачив я в своєму видінні вночі, аж ось чотири небесні вітри вдарили на Велике море.
DAN|7|3|І чотири великі звірі піднялися з моря, різні один від одного.
DAN|7|4|Передній був, як лев, а крила в нього орлині. Я бачив, аж ось були вирвані йому крила, і він був піднятий від землі, і поставлений на ноги, як людина, і серце людське було йому дане.
DAN|7|5|А ось звір інший, другий, подібний до ведмедя, і був поставлений на одному боці, і було три ребрі в його пащі між зубами його. І йому сказали так: Уставай, їж багато м'яса!
DAN|7|6|Потому я бачив, аж ось звір інший, мов пантера, а в нього на спині чотири пташині крилі. Цей звір мав чотири голові, і була йому дана влада.
DAN|7|7|Потому я бачив у видіннях тієї ночі, аж ось четвертий звір, страшний і грізний, та надмірно міцний, і в нього великі залізні зуби. Він жер та торощив, а решту ногами своїми топтав, і він різнився від усіх звірів, що були перед ним, і мав десять рогів.
DAN|7|8|Я приглядався до тих рогів, аж ось поміж ними піднісся ріг інший, малий, а три з тих передніх рогів були вирвані з коренем перед ним. І ось у того рога очі, як очі людські, і уста, що говорили про великі речі.
DAN|7|9|Я бачив, аж ось поставили престоли, і всівся Старий днями. Одежа Його біла, як сніг, а волосся голови Його немов чиста вовна, а престол Його огняне полум'я, колеса Його палахкотючий огонь.
DAN|7|10|Огненна річка пливла й виходила з-перед Нього; тисяча тисяч служили Йому, і десять тисяч десятків тисяч стояли перед Ним; суд усівся, і розгорнулися книги.
DAN|7|11|Я бачив того часу, що від голосу великих слів, які цей ріг говорив, я бачив, аж ось був забитий той звір, і було погублене тіло його, і було віддане на спалення огню.
DAN|7|12|А решті тих звірів відняли їхнє панування, а довгота в житті була їм дана аж до усталеного часу та години.
DAN|7|13|Я бачив у видіннях ночі, аж ось разом з небесними хмарами йшов ніби Син Людський, і прийшов аж до Старого днями, і Його підвели перед Нього.
DAN|7|14|І Йому було дане панування й слава та царство, і всі народи, племена та язики будуть служити Йому. Панування Його панування вічне, яке не спиниться, а царство Його не буде зруйноване.
DAN|7|15|Дух мій, Даниїлів, був засумований через це, і видіння голови моєї стурбували мене.
DAN|7|16|Я наблизився до одного з тих, що стояли, і поспитався від нього про істоту всього того. І він сказав мені, і познайомив мене з розв'язкою цих речей.
DAN|7|17|Ці великі звірі, що їх чотири, це чотири царі встануть з землі.
DAN|7|18|І приймуть царство святі Всевишнього, і будуть міцно держати царювання аж навіки, і аж на віки віків.
DAN|7|19|Тоді хотів я знати певне про четвертого звіра, що різнився від їх усіх, він страшний, надмірний, зуби його залізні, а пазурі його мідяні, він жер та торощив, а решту ногами своїми топтав,
DAN|7|20|і про десять рогів, що на його голові, і про іншого, що піднісся, а три через нього випали, і про цього рога, що мав очі, а уста говорили про великі речі, а вид його більший від його друзів.
DAN|7|21|Я бачив, що цей ріг учинив бій зо святими, і переміг їх.
DAN|7|22|Аж ось прийшов Старий днями, і даний був суд святим Всевишнього, і надійшов умовлений час, і царство взяли святі.
DAN|7|23|Він так сказав: Четвертий звір четверте царство буде на землі, яке буде різнитися від усіх царств, і пожере всю землю, і вимолотить її та розторощить її.
DAN|7|24|А десять рогів визначають, що з того царства встане десять царів, а по них встане інший, що буде різнитися від попередніх, і скине трьох царів.
DAN|7|25|І він буде говорити слова проти Всевишнього, і пригнобить святих Всевишнього, і буде думати позмінювати свята та права, і вони віддані будуть у його руку аж до одного часу, і часів і половини часу.
DAN|7|26|Та засяде суд, і скинуть його панування, щоб його знищити та вигубити аж до кінця.
DAN|7|27|А царство, і панування, і велич царств під усім небом буде дане народові святих Всевишнього. Його царство буде царство вічне, а всі панування Йому будуть служити й будуть слухняні.
DAN|7|28|Аж поти кінець цього слова. Мене, Даниїла, сильно лякали думки мої, і змінилася ясність моя, але це слово я заховав у своїм серці.
DAN|8|1|За третього року царювання царя Валтасара з'явилося мені, Даниїлові, видіння по тому, що з'явилося мені перше.
DAN|8|2|І бачив я в видінні, і сталося в моєму видінні, а я був у твердині Шушані, що в окрузі Еламі, і бачив я в видінні, ніби я був над потоком Улай.
DAN|8|3|І звів я очі свої та й побачив, аж ось один баран стоїть перед потоком, і в нього два роги. А обидва ці роги високі, і один вищий від другого, а той вищий виріс наостанку.
DAN|8|4|Я бачив барана, що колов на захід, і на північ, і на південь, і жоден звір не міг стати проти нього, і не було нікого, хто б урятував від його руки. І він робив за своїм уподобанням, і став величний.
DAN|8|5|І я придивлявся, аж ось козел з кіз приходить із заходу по поверхні всієї землі, і не дотикається до землі. А той козел мав подобу рога між своїми очима.
DAN|8|6|І прийшов він до того барана, що мав ті два роги, якого я бачив, що стояв перед потоком, і помчав на нього в лютості своєї сили.
DAN|8|7|І я бачив його, що він добіг аж до барана, і роз'ярився на нього, та й ударив того барана, і зламав йому ті два роги, а в барана не було сили стати проти нього. І той кинув його на землю, і потоптав його, і не було нікого, хто б вирятував барана від його руки.
DAN|8|8|А козел з кіз став аж надто великий. А коли він зміцнився, то був зламаний той великий ріг, а замість нього виросли чотири подобі рога на чотири вітри неба.
DAN|8|9|А з одного з них вийшов один малий ріг, і з малого став дуже великий до півдня, і до сходу, і до Пишноти.
DAN|8|10|І він побільшився аж до війська небесного, і скинув на землю декого з війська, із зір, і потоптав їх.
DAN|8|11|І він побільшився аж до Вождя того війська, і від Нього була віднята стала жертва, і покинене місце святині Його.
DAN|8|12|І буде віддане йому військо враз із щоденною службою через гріхи, і він кине правду на землю, і зробить, і матиме успіх.
DAN|8|13|І почув я одного святого, що говорив. А інший святий сказав до того, що говорив: Аж доки це видіння про сталу жертву та про нищівний гріх, доки святиня й військо віддані на топтання?
DAN|8|14|І відказав він мені: Аж до двох тисяч і трьох сотень вечорів-ранків, тоді буде визнана очищеною святиня.
DAN|8|15|І сталося, коли я, Даниїл, бачив те видіння, і шукав значення його, ось став передо мною ніби муж.
DAN|8|16|І почув я поміж берегами Улаю людський голос, що кликнув і сказав: Гавриїле, виясни йому це видіння!
DAN|8|17|І він прийшов туди, де я стояв, а коли він прийшов, я настрашився й упав на обличчя своє. І сказав він мені: Зрозумій, сину людський, бо на час кінця це видіння!
DAN|8|18|А коли він говорив зо мною, я зомлів, і припав своїм обличчям до землі, але він діткнувся до мене, і поставив мене на моєму місці,
DAN|8|19|та й сказав: Ось я об'являю тобі, що буде в кінці гніву, бо на кінець призначеного часу це видіння.
DAN|8|20|Той козел, якого ти бачив, що мав ті два роги, це царі мідян та персів.
DAN|8|21|А козел, той волохатий, це цар Греції, а той великий ріг, що між очима його, це перший цар.
DAN|8|22|А той зламаний ріг, і що стали на його місці чотири, це чотири царства постануть із цього народу, але вже не в його силі.
DAN|8|23|А в кінці їхнього царства, коли покінчать своє ті грішники, постане цар нахабний та вправний у підступах.
DAN|8|24|І зміцніє його сила, але не його власною силою, і дивно винищить він, і буде мати успіх, і діятиме. І винищить він сильних і народ святих.
DAN|8|25|А через свою мудрість буде мати успіх, омана буде в його руці, і він звеличиться в своєму серці. І в часі миру він понищить багатьох, і повстане на Владику над владиками, але без руки буде зламаний.
DAN|8|26|А видіння вечора та ранку, про яке було сказано, це правда, та ти сховай це видіння, бо воно відноситься на далекі часи.
DAN|8|27|А я, Даниїл, знемігся й заслаб на кілька днів. І встав я, і робив цареву працю, і остовпів з того видіння, але ніхто того не завважив.
DAN|9|1|За першого року Дарія, Ахашверошового сина, з насіння мідян, що зацарював над халдейським царством,
DAN|9|2|за першого року його царювання я, Даниїл, бачив у книгах число тих років, про які було Господнє слово до пророка Єремії, що сповниться для руїн Єрусалиму сімдесят років.
DAN|9|3|І звернув я своє обличчя до Господа Бога, прохати з молитвою та з благаннями, у пості, у веретищі та в попелі.
DAN|9|4|І молився я Господеві, Богові своєму, і сповідався й казав: О мій Господи, Боже великий і грізний, що стережеш заповіта та милість для тих, хто кохає Тебе, та для тих, хто виконує Твої заповіді!
DAN|9|5|Ми прогрішилися та чинили беззаконня, і були несправедливі, і бунтувалися, і відверталися від Твоїх заповідей та від постанов Твоїх.
DAN|9|6|І не прислухалися ми до Твоїх рабів пророків, що говорили в Твоїм Імені до наших царів, наших начальників та наших батьків, і до всього народу землі.
DAN|9|7|Тобі, Господи, справедливість, а нам сором на обличчя, як цього дня для юдея, і для мешканців Єрусалиму, і для всього Ізраїля, близьких та далеких, по всіх тих краях, куди Ти їх вигнав за їхнє спроневірення, що допустилися його перед Тобою.
DAN|9|8|Господи, сором на обличчя нам, нашим царям, князям нашим та нашим батькам, що згрішили перед Тобою!
DAN|9|9|А Господеві, нашому Богові, милість та прощення, бо ми бунтувалися проти Нього,
DAN|9|10|і не слухалися голосу Господа, нашого Бога, щоб ходити законами Його, які Він дав нам через Своїх рабів пророків.
DAN|9|11|І ввесь Ізраїль переступив Закона Твого, і відвернулися, щоб не слухатися Твого голосу, і було вилите на нас те прокляття й та присяга, що написана в Законі Мойсея, Божого раба, бо ми прогрішилися Йому.
DAN|9|12|І Він сповнив Своє слово, яке говорив на нас та на наших суддів, що судили нас, щоб спровадити на нас велике зло, такого не було вчинено під цілим небом, яке було вчинене в Єрусалимі!
DAN|9|13|Як написано в Мойсеєвому Законі, усе те лихо прийшло на нас, та ми не вблагали Господа, нашого Бога, щоб вернутися нам від свого гріха, і щоб порозумнішати в Твоїй правді.
DAN|9|14|І Господь пильнував того лиха, і спровадив його на нас, бо справедливий Господь, Бог наш, у всіх Своїх чинах, які Він зробив, та ми не слухали Його голосу.
DAN|9|15|А тепер, Господи, Боже наш, що вивів з єгипетського краю Свій народ потужною рукою, і зробив Собі славне Ім'я, як цього дня, згрішили ми, стали несправедливі!
DAN|9|16|Господи, у міру всієї Твоєї справедливости нехай відвернеться гнів Твій та Твоя ревність від Твого міста Єрусалиму, Твоєї святої гори, бо через наші гріхи та через провини наших батьків Єрусалим та народ Твій відданий на ганьбу для всіх наших околиць.
DAN|9|17|І нині прислухайся, Боже наш, до молитви Твого раба та до його благань, і нехай засвітиться Твоє лице над Твоєю спустошеною святинею, ради Господа!
DAN|9|18|Нахили, Боже мій, вухо Своє та й послухай, відкрий Свої очі й побач наші спустошення та те місто, де кликалося Ім'я Твоє в ньому, бо ми кладемо свої благання перед Твоїм лицем не через свої справедливості, але через велику Твою милість.
DAN|9|19|Господи, вислухай! Господи, прости! Господи, прислухайся й зроби! Не опізняйся ради Себе, мій Боже, бо Ім'я Твоє кличеться над Твоїм містом і над Твоїм народом!
DAN|9|20|А ще я говорив і молився, та ісповідував гріх свій та народу мого Ізраїля, і клав свою молитву перед лице Господа, мого Бога, за святу гору мого Бога,
DAN|9|21|і ще я говорив на цій молитві, а той муж Гавриїл, якого я бачив у видінні напочатку, швидко прилетів, і доторкнувся до мене за часу вечірньої хлібної жертви.
DAN|9|22|І він напучував мене, і говорив зо мною та й сказав: Даниїле, я тепер вийшов, щоб умудрити тебе в розумінні.
DAN|9|23|На початку молитов твоїх вийшло слово, і я прийшов об'явити його тобі, бо ти улюблений, і приглянься до цього слова, і придивися до видіння.
DAN|9|24|Сімдесят років-тижнів призначено для твого народу та для міста твоєї святині, аж поки переступ буде докінчений, і міра гріха буде повна, аж поки вина буде спокутувана, і вічна правда приведена, аж поки будуть потверджені видіння й пророк, і щоб помазати Святеє Святих.
DAN|9|25|Та знай і розумій: від виходу наказу, щоб вернути Ізраїля й збудувати Єрусалим, аж до Владики Месії сім тижнів та шістдесят і два тижні. І вернеться народ, і відбудований буде майдан і вулиця, і то буде за тяжкого часу.
DAN|9|26|І по тих шостидесятьох і двох тижнях буде погублений Месія, хоч не буде на Ньому вини. А це місто й святиню знищить народ володаря, що прийде, а кінець його у повідді. І аж до кінця буде війна, гострі спустошення.
DAN|9|27|І Він зміцнить заповіта для багатьох за один тиждень, а за півтижня припинить жертву та жертву хлібну. І на святиню прийде гидота спустошення, поки знищення й рішучий суд кари не виллється на спустошителя.
DAN|10|1|За третього року Кіра, перського царя, було відкрите слово Даниїлові, що звався ім'ям Валтасар, а слово це правда та великий труд; і він зрозумів те слово, і мав зрозуміння того видіння.
DAN|10|2|Тими днями я, Даниїл, був у жалобі три тижні часу.
DAN|10|3|Любої страви я не їв, а м'ясо й вино не входило до моїх уст, і намащуватися не намащувався я аж до виповнення цих трьох тижнів часу.
DAN|10|4|А двадцятого й четвертого дня першого місяця та був я при великій річці, це Хіддекел.
DAN|10|5|І звів я свої очі та й побачив, аж ось один чоловік, одягнений у льняну одіж, а стегна його оперезані золотом з Уфазу.
DAN|10|6|А тіло його як топаз, а обличчя його як вид блискавки, а очі його як огняне полум'я, а рамена його та ноги його ніби блискуча мідь, а звук слів його як гук натовпу.
DAN|10|7|А я, Даниїл, сам бачив це видіння, а люди, що були разом зо мною, не бачили цього видіння, але велике тремтіння спало на них, і вони повтікали в укриття.
DAN|10|8|А я зостався сам, і бачив це велике видіння, і не зосталося в мені сили, а краса обличчя мого змінилася й знищилася, і я не задержав у собі сили...
DAN|10|9|І почув я голос його слів. А як почув я голос його слів, то я зомлів, і припав своїм обличчям до землі.
DAN|10|10|І ось рука доторкнулася до мене, і звела мене на коліна мої та на долоні моїх рук.
DAN|10|11|І сказав він до мене: Даниїле, мужу любий, зрозумій ті слова, що я скажу тобі, і стань на своєму місці, бо тепер я посланий до тебе! А коли він говорив зо мною це слово, устав я й тремтів.
DAN|10|12|А він промовив до мене: Не бійся, Даниїле, бо від першого дня, коли ти дав своє серце, щоб зрозуміти видіння, і щоб упокоритися перед лицем твого Бога, були почуті слова твої, і я прийшов ради твоїх слів.
DAN|10|13|Але князь перського царства стояв проти мене двадцять і один день, і ось Михаїл, один із перших начальників, прийшов допомогти мені, а я позоставив його там при начальниках перських царів.
DAN|10|14|І прийшов я, щоб ти зрозумів, що станеться твоєму народові в кінці днів, бо це видіння ще на наступні дні.
DAN|10|15|А коли він говорив зо мною оці слова, я схилив своє обличчя до землі, і занімів.
DAN|10|16|І ось хтось, як подоба до людських синів, доторкнувся до губ моїх, і я відкрив свої уста, і говорив та й сказав тому, хто стояв передо мною: Мій пане, у цьому видінні обернулися на мене болі мої, і я не задержав сили в собі.
DAN|10|17|І як може цей раб мого пана говорити з оцим моїм паном, коли в мені тепер нема сили, і не залишилося й духу?
DAN|10|18|І знов доторкнувся до мене хтось, як вид людини, і зміцнив мене,
DAN|10|19|та й сказав: Не бійся, любий мужу, мир тобі! Будь міцний і будь сильний! А коли він говорив зо мною, я зміцнився й сказав: Нехай говорить мій пан, бо я зміцнився!
DAN|10|20|І він сказав: Чи ти знаєш, чого я до тебе прийшов? Та тепер я вертаюсь, щоб воювати з перським князем, а коли вийду, то ось прийде грецький князь.
DAN|10|21|Але об'являю тобі записане в книзі правди. І немає нікого, хто зміцняв би мене проти них, окрім вашого князя Михаїла.
DAN|11|1|А я в першому році мідянина Дарія стояв, щоб зміцнити й посилити його.
DAN|11|2|А тепер об'явлю тобі правду. Ось іще три царі повстануть для Персії, а четвертий збагатиться багатством, більшим від усіх, а своєю силою в багатстві своїм підбурить усе проти грецького царства.
DAN|11|3|І повстане хоробрий цар, і запанує великим пануванням, і робитиме за своїм уподобанням.
DAN|11|4|Та коли він повстане, буде зруйноване його царство, і буде розділене на чотири небесні вітри, а не на його нащадків, і не за його пануванням, яким він панував, бо царство його буде вирване й дане іншим, а не їм.
DAN|11|5|І зміцниться південний цар, але один з його князів пересилить його й запанує, його панування панування велике.
DAN|11|6|Але по роках вони поєднаються, і дочка південного царя прийде до царя північного, щоб зробити мир. Але не затримає він сили свого рамена, і не встане потомство його, але буде видана вона й ті, що вели її, і та, що її породила, і той, що міцно тримав її за тих часів.
DAN|11|7|І повстане один із галузки її кореня на його місце, і він вийде проти війська, і ввійде в твердиню північного царя, і буде діяти проти них, і опанує їх.
DAN|11|8|І їхніх богів з їхніми литими бовванами, разом з їхнім улюбленим посудом, золотом та сріблом поведе в неволю до Єгипту, і він роки стоятиме більше від північного царя.
DAN|11|9|І він увійде в царство південного царя, але вернеться до своєї землі.
DAN|11|10|А сини його озброються, і зберуть натовп численних войовників, і один із них конче піде, і все позаливає, і перейде край, і вернеться, і воюватиме аж до його твердині.
DAN|11|11|І розлютиться південний цар, і вийде та й воюватиме з ним, з царем північним, і виставить велике многолюдство, і цей натовп буде відданий у його руку.
DAN|11|12|І буде знищений той натовп, і повищиться його серце, і він кине десятитисячки, та не буде сильний.
DAN|11|13|І вернеться північний цар, і виставить натовп, більший від першого, а на кінець часів та років він конче прийде з великим військом та з численним маєтком.
DAN|11|14|І за того часу багато-хто повстануть на південного царя, а сини насильників твого народу підіймуться, щоб справдилось видіння, і вони спіткнуться.
DAN|11|15|І прийде північний цар, і насипле вала, і здобуде твердинне місто, і не встоять рамена півдня та його добірний народ, і не буде сили встояти.
DAN|11|16|І робитиме той, хто прийде на нього, за своєю вподобою, і не буде того, хто встояв би перед ним. І стане він у Пишному Краї, і буде погибель у його руці.
DAN|11|17|І зверне він своє обличчя, щоб прийти з потугою всього свого царства, і складе договора з ним. І дасть йому молоду дочку за жінку, щоб знищити землю, та це не вдасться, і не станеться йому.
DAN|11|18|І зверне він обличчя своє на острови, і здобуде багато. Але вождь спинить йому наругу його, всемеро заплатить йому за наруги його.
DAN|11|19|І зверне він своє обличчя до твердинь свого краю, і спіткнеться й упаде, і не буде знайдений.
DAN|11|20|А на його місці стане той, що скаже побірникові податків перейти пишноту царства, та за кілька днів від загине, але не від гніву й не від бою.
DAN|11|21|І стане на його місці погорджуваний, та не дадуть йому царської пошани, але він прийде непомітно, й опанує царство лестощами.
DAN|11|22|А війська, що затоплювали, він затопить і знищить, і навіть самого володаря, що з ним поєднався.
DAN|11|23|А від часу поєднання з ним він робитиме оману, і підійметься, і зміцниться малим народом.
DAN|11|24|Він увійде непомітно в ситу округу, і зробить те, чого не робили батьки його та батьки його батьків. Він порозкидає їм награбоване, і здобич, і маєток, і на твердині буде замишляти свої задуми, але до часу.
DAN|11|25|І він збудить свою силу та своє серце на південного царя з великим військом. А південний цар підготовиться до війни з військом великим та дуже міцним, та не встоїть, бо замишляють на нього задуми.
DAN|11|26|А ті, що їдять його поживу, поб'ють його, і його військо позаливає край, і попадають численні забиті.
DAN|11|27|А серце обох цих царів буде на лихе, і при одному столі вони будуть говорити неправду, але не буде успіху, бо кінець буде ще відкладений на означений час.
DAN|11|28|І він вернеться до свого краю з великим маєтком, а його серце буде проти святого заповіту; і він зробить, і вернеться до свого краю.
DAN|11|29|На умовлений час він повернеться, і прийде на південь, але останнє не буде, як перше.
DAN|11|30|І прийдуть на нього кіттейські кораблі, і він налякається, і вернеться, і буде чинити опір святому заповітові, і зробить своє. І він вернеться, і погодиться з тими, хто покинув святий заповіт.
DAN|11|31|І повстануть його війська та й зневажать святиню, твердиню, і спинять сталу жертву, і поставлять гидоту спустошення.
DAN|11|32|А тих, хто чинить несправедливе на заповіт, він прихилить через лестощі. А народ, що знає свого Бога, зміцніє та й діятиме.
DAN|11|33|А розумні з народу навчать багатьох, але спіткнуться об меча та полум'я, об полон та грабіж якийсь час.
DAN|11|34|А коли вони спіткнуться, будуть споможені малою поміччю, хоч до них прилучаться багато-хто лестощами.
DAN|11|35|А дехто з тих розумних спіткнуться, щоб очистити себе, і щоб вибрати, і щоб вибілитися аж до кінцевого часу, бо ще час до умовленого часу.
DAN|11|36|І буде робити той цар за своїм уподобанням, і підійметься, і повищиться понад усякого бога, і на Бога богів говоритиме дивні речі, і матиме успіх, аж поки не довершиться гнів, бо виконається те, що було вирішене.
DAN|11|37|І він не буде придивлятися до богів своїх батьків, і на пожадливість жінок, і на всякого бога не буде дивитися, бо він звеличить себе понад кожного.
DAN|11|38|Але він буде віддавати честь богові твердинь на його місці, та богові, якого не знали батьки його, віддаватиме честь золотом, і сріблом, і дорогоцінним камінням, і речами коштовними.
DAN|11|39|І він посадить у твердині народа чужого бога. Тому, хто пізнає його, примножить славу, і вчинить їх панами над багатьма, і поділить землю на заплату.
DAN|11|40|А в кінцевому часі зудариться з ним південний цар. І кинеться на нього північний цар колесницями, і верхівцями, і численними кораблями, і прийде на краї, і позаливає та перейде їх.
DAN|11|41|І він прийде до Пишного Краю, і багато-хто спіткнуться, та оці втечуть від його руки: Едом, і Моав, і останок Аммонових синів.
DAN|11|42|І він простягне свою руку на краї, і не втече єгипетський край.
DAN|11|43|І він запанує над скарбами золота й срібла, та над усіма коштовними речами Єгипту. А лівійці та етіопляни підуть за ним.
DAN|11|44|Але його налякають вістки зо сходу та з півночі, і він вийде з великою лютістю, щоб багатьох погубити та зробити закляттям.
DAN|11|45|І поставить намети свого палацу між морями та горою пишної святині. Та він прийде до свого кінця, але не буде йому помічника.
DAN|12|1|І повстане того часу Михаїл, великий той князь, що стоїть при синах твого народу, і буде час утиску, якого не було від існування люду аж до цього часу. І того часу буде врятований із народу твого кожен, хто буде знайдений записаним у книзі.
DAN|12|2|І багато-хто з тих, що сплять у земному поросі, збудяться, одні на вічне життя, а одні на наруги, на вічну гидоту.
DAN|12|3|А розумні будуть сяяти, як світила небозводу, а ті, хто привів багатьох до праведности, немов зорі, навіки віків.
DAN|12|4|А ти, Даниїле, заховай ці слова, і запечатай цю книгу аж до часу кінця. Багато-хто дослідять її, і так розмножиться знання.
DAN|12|5|І побачив я, Даниїл, аж ось стоять два інші Анголи, один тут при цьому березі річки, а один там при тому березі річки.
DAN|12|6|І сказав він до мужа, одягненого в льняну одіж, що був над водою річки: Коли буде кінець цим дивним речам?
DAN|12|7|І почув я того мужа, одягненого в льняну одіж, що був над водою річки. І звів він до неба свою правицю та свою лівицю, і присягнув вічно Живим: це буде за час, за часи і за пів часу, і коли скінчиться розбивання сили святого народу, все це сповниться.
DAN|12|8|А я це слухав і не розумів. І сказав я: Мій пане, який цьому кінець?
DAN|12|9|І він сказав: Іди, Даниїле, бо заховані й запечатані ці слова аж до часу кінця.
DAN|12|10|Багато-хто будуть очищені, і вибіляться, і будуть перетоплені; і будуть несправедливі несправедливими, і цього не зрозуміють усі несправедливі, а розумні зрозуміють.
DAN|12|11|А від часу, коли буде припинена стала жертва, щоб була поставлена гидота спустошення, мине тисяча двісті й дев'ятдесят день.
DAN|12|12|Благословенний той, хто чекає, і досягне до тисячі трьох сотень тридцяти й п'яти день!
DAN|12|13|А ти йди до кінця, і відпочинеш, і встанеш на свою долю під кінець тих днів!
