JUDG|1|1|After the death of Joshua, the people of Israel inquired of the LORD, "Who shall go up first for us against the Canaanites, to fight against them?"
JUDG|1|2|The LORD said, "Judah shall go up; behold, I have given the land into his hand."
JUDG|1|3|And Judah said to Simeon his brother, "Come up with me into the territory allotted to me, that we may fight against the Canaanites. And I likewise will go with you into the territory allotted to you." So Simeon went with him.
JUDG|1|4|Then Judah went up and the LORD gave the Canaanites and the Perizzites into their hand, and they defeated 10,000 of them at Bezek.
JUDG|1|5|They found Adoni-bezek at Bezek and fought against him and defeated the Canaanites and the Perizzites.
JUDG|1|6|Adoni-bezek fled, but they pursued him and caught him and cut off his thumbs and his big toes.
JUDG|1|7|And Adoni-bezek said, "Seventy kings with their thumbs and their big toes cut off used to pick up scraps under my table. As I have done, so God has repaid me." And they brought him to Jerusalem, and he died there.
JUDG|1|8|And the men of Judah fought against Jerusalem and captured it and struck it with the edge of the sword and set the city on fire.
JUDG|1|9|And afterward the men of Judah went down to fight against the Canaanites who lived in the hill country, in the Negeb, and in the lowland.
JUDG|1|10|And Judah went against the Canaanites who lived in Hebron (now the name of Hebron was formerly Kiriath-arba), and they defeated Sheshai and Ahiman and Talmai.
JUDG|1|11|From there they went against the inhabitants of Debir. The name of Debir was formerly Kiriath-sepher.
JUDG|1|12|And Caleb said, "He who attacks Kiriath-sepher and captures it, I will give him Achsah my daughter for a wife."
JUDG|1|13|And Othniel the son of Kenaz, Caleb's younger brother, captured it. And he gave him Achsah his daughter for a wife.
JUDG|1|14|When she came to him, she urged him to ask her father for a field. And she dismounted from her donkey, and Caleb said to her, "What do you want?"
JUDG|1|15|She said to him, "Give me a blessing. Since you have set me in the land of the Negeb, give me also springs of water." And Caleb gave her the upper springs and the lower springs.
JUDG|1|16|And the descendants of the Kenite, Moses' father-in-law, went up with the people of Judah from the city of palms into the wilderness of Judah, which lies in the Negeb near Arad, and they went and settled with the people.
JUDG|1|17|And Judah went with Simeon his brother, and they defeated the Canaanites who inhabited Zephath and devoted it to destruction. So the name of the city was called Hormah.
JUDG|1|18|Judah also captured Gaza with its territory, and Ashkelon with its territory, and Ekron with its territory.
JUDG|1|19|And the LORD was with Judah, and he took possession of the hill country, but he could not drive out the inhabitants of the plain because they had chariots of iron.
JUDG|1|20|And Hebron was given to Caleb, as Moses had said. And he drove out from it the three sons of Anak.
JUDG|1|21|But the people of Benjamin did not drive out the Jebusites who lived in Jerusalem, so the Jebusites have lived with the people of Benjamin in Jerusalem to this day.
JUDG|1|22|The house of Joseph also went up against Bethel, and the LORD was with them.
JUDG|1|23|And the house of Joseph scouted out Bethel. (Now the name of the city was formerly Luz.)
JUDG|1|24|And the spies saw a man coming out of the city, and they said to him, "Please show us the way into the city, and we will deal kindly with you."
JUDG|1|25|And he showed them the way into the city. And they struck the city with the edge of the sword, but they let the man and all his family go.
JUDG|1|26|And the man went to the land of the Hittites and built a city and called its name Luz. That is its name to this day.
JUDG|1|27|Manasseh did not drive out the inhabitants of Beth-shean and its villages, or Taanach and its villages, or the inhabitants of Dor and its villages, or the inhabitants of Ibleam and its villages, or the inhabitants of Megiddo and its villages, for the Canaanites persisted in dwelling in that land.
JUDG|1|28|When Israel grew strong, they put the Canaanites to forced labor, but did not drive them out completely.
JUDG|1|29|And Ephraim did not drive out the Canaanites who lived in Gezer, so the Canaanites lived in Gezer among them.
JUDG|1|30|Zebulun did not drive out the inhabitants of Kitron, or the inhabitants of Nahalol, so the Canaanites lived among them, but became subject to forced labor.
JUDG|1|31|Asher did not drive out the inhabitants of Acco, or the inhabitants of Sidon or of Ahlab or of Achzib or of Helbah or of Aphik or of Rehob,
JUDG|1|32|so the Asherites lived among the Canaanites, the inhabitants of the land, for they did not drive them out.
JUDG|1|33|Naphtali did not drive out the inhabitants of Beth-shemesh, or the inhabitants of Beth-anath, so they lived among the Canaanites, the inhabitants of the land. Nevertheless, the inhabitants of Beth-shemesh and of Beth-anath became subject to forced labor for them.
JUDG|1|34|The Amorites pressed the people of Dan back into the hill country, for they did not allow them to come down to the plain.
JUDG|1|35|The Amorites persisted in dwelling in Mount Heres, in Aijalon, and in Shaalbim, but the hand of the house of Joseph rested heavily on them, and they became subject to forced labor.
JUDG|1|36|And the border of the Amorites ran from the ascent of Akrabbim, from Sela and upward.
JUDG|2|1|Now the angel of the LORD went up from Gilgal to Bochim. And he said, "I brought you up from Egypt and brought you into the land that I swore to give to your fathers. I said, 'I will never break my covenant with you,
JUDG|2|2|and you shall make no covenant with the inhabitants of this land; you shall break down their altars.' But you have not obeyed my voice. What is this you have done?
JUDG|2|3|So now I say, I will not drive them out before you, but they shall become thorns in your sides, and their gods shall be a snare to you."
JUDG|2|4|As soon as the angel of the LORD spoke these words to all the people of Israel, the people lifted up their voices and wept.
JUDG|2|5|And they called the name of that place Bochim. And they sacrificed there to the LORD.
JUDG|2|6|When Joshua dismissed the people, the people of Israel went each to his inheritance to take possession of the land.
JUDG|2|7|And the people served the LORD all the days of Joshua, and all the days of the elders who outlived Joshua, who had seen all the great work that the LORD had done for Israel.
JUDG|2|8|And Joshua the son of Nun, the servant of the LORD, died at the age of 110 years.
JUDG|2|9|And they buried him within the boundaries of his inheritance in Timnath-heres, in the hill country of Ephraim, north of the mountain of Gaash.
JUDG|2|10|And all that generation also were gathered to their fathers. And there arose another generation after them who did not know the LORD or the work that he had done for Israel.
JUDG|2|11|And the people of Israel did what was evil in the sight of the LORD and served the Baals.
JUDG|2|12|And they abandoned the LORD, the God of their fathers, who had brought them out of the land of Egypt. They went after other gods, from among the gods of the peoples who were around them, and bowed down to them. And they provoked the LORD to anger.
JUDG|2|13|They abandoned the LORD and served the Baals and the Ashtaroth.
JUDG|2|14|So the anger of the LORD was kindled against Israel, and he gave them over to plunderers, who plundered them. And he sold them into the hand of their surrounding enemies, so that they could no longer withstand their enemies.
JUDG|2|15|Whenever they marched out, the hand of the LORD was against them for harm, as the LORD had warned, and as the LORD had sworn to them. And they were in terrible distress.
JUDG|2|16|Then the LORD raised up judges, who saved them out of the hand of those who plundered them.
JUDG|2|17|Yet they did not listen to their judges, for they whored after other gods and bowed down to them. They soon turned aside from the way in which their fathers had walked, who had obeyed the commandments of the LORD, and they did not do so.
JUDG|2|18|Whenever the LORD raised up judges for them, the LORD was with the judge, and he saved them from the hand of their enemies all the days of the judge. For the LORD was moved to pity by their groaning because of those who afflicted and oppressed them.
JUDG|2|19|But whenever the judge died, they turned back and were more corrupt than their fathers, going after other gods, serving them and bowing down to them. They did not drop any of their practices or their stubborn ways.
JUDG|2|20|So the anger of the LORD was kindled against Israel, and he said, "Because this people have transgressed my covenant that I commanded their fathers and have not obeyed my voice,
JUDG|2|21|I will no longer drive out before them any of the nations that Joshua left when he died,
JUDG|2|22|in order to test Israel by them, whether they will take care to walk in the way of the LORD as their fathers did, or not."
JUDG|2|23|So the LORD left those nations, not driving them out quickly, and he did not give them into the hand of Joshua.
JUDG|3|1|Now these are the nations that the LORD left, to test Israel by them, that is, all in Israel who had not experienced all the wars in Canaan.
JUDG|3|2|It was only in order that the generations of the people of Israel might know war, to teach war to those who had not known it before.
JUDG|3|3|These are the nations: the five lords of the Philistines and all the Canaanites and the Sidonians and the Hivites who lived on Mount Lebanon, from Mount Baal-hermon as far as Lebo-hamath.
JUDG|3|4|They were for the testing of Israel, to know whether Israel would obey the commandments of the LORD, which he commanded their fathers by the hand of Moses.
JUDG|3|5|So the people of Israel lived among the Canaanites, the Hittites, the Amorites, the Perizzites, the Hivites, and the Jebusites.
JUDG|3|6|And their daughters they took to themselves for wives, and their own daughters they gave to their sons, and they served their gods.
JUDG|3|7|And the people of Israel did what was evil in the sight of the LORD. They forgot the LORD their God and served the Baals and the Asheroth.
JUDG|3|8|Therefore the anger of the LORD was kindled against Israel, and he sold them into the hand of Cushan-rishathaim king of Mesopotamia. And the people of Israel served Cushan-rishathaim eight years.
JUDG|3|9|But when the people of Israel cried out to the LORD, the LORD raised up a deliverer for the people of Israel, who saved them, Othniel the son of Kenaz, Caleb's younger brother.
JUDG|3|10|The Spirit of the LORD was upon him, and he judged Israel. He went out to war, and the LORD gave Cushan-rishathaim king of Mesopotamia into his hand. And his hand prevailed over Cushan-rishathaim.
JUDG|3|11|So the land had rest forty years. Then Othniel the son of Kenaz died.
JUDG|3|12|And the people of Israel again did what was evil in the sight of the LORD, and the LORD strengthened Eglon the king of Moab against Israel, because they had done what was evil in the sight of the LORD.
JUDG|3|13|He gathered to himself the Ammonites and the Amalekites, and went and defeated Israel. And they took possession of the city of palms.
JUDG|3|14|And the people of Israel served Eglon the king of Moab eighteen years.
JUDG|3|15|Then the people of Israel cried out to the LORD, and the LORD raised up for them a deliverer, Ehud, the son of Gera, the Benjaminite, a left-handed man. The people of Israel sent tribute by him to Eglon the king of Moab.
JUDG|3|16|And Ehud made for himself a sword with two edges, a cubit in length, and he bound it on his right thigh under his clothes.
JUDG|3|17|And he presented the tribute to Eglon king of Moab. Now Eglon was a very fat man.
JUDG|3|18|And when Ehud had finished presenting the tribute, he sent away the people who carried the tribute.
JUDG|3|19|But he himself turned back at the idols near Gilgal and said, "I have a secret message for you, O king." And he commanded, "Silence." And all his attendants went out from his presence.
JUDG|3|20|And Ehud came to him as he was sitting alone in his cool roof chamber. And Ehud said, "I have a message from God for you." And he arose from his seat.
JUDG|3|21|And Ehud reached with his left hand, took the sword from his right thigh, and thrust it into his belly.
JUDG|3|22|And the hilt also went in after the blade, and the fat closed over the blade, for he did not pull the sword out of his belly; and the dung came out.
JUDG|3|23|Then Ehud went out into the porch and closed the doors of the roof chamber behind him and locked them.
JUDG|3|24|When he had gone, the servants came, and when they saw that the doors of the roof chamber were locked, they thought, "Surely he is relieving himself in the closet of the cool chamber."
JUDG|3|25|And they waited till they were embarrassed. But when he still did not open the doors of the roof chamber, they took the key and opened them, and there lay their lord dead on the floor.
JUDG|3|26|Ehud escaped while they delayed, and he passed beyond the idols and escaped to Seirah.
JUDG|3|27|When he arrived, he sounded the trumpet in the hill country of Ephraim. Then the people of Israel went down with him from the hill country, and he was their leader.
JUDG|3|28|And he said to them, "Follow after me, for the LORD has given your enemies the Moabites into your hand." So they went down after him and seized the fords of the Jordan against the Moabites and did not allow anyone to pass over.
JUDG|3|29|And they killed at that time about 10,000 of the Moabites, all strong, able-bodied men; not a man escaped.
JUDG|3|30|So Moab was subdued that day under the hand of Israel. And the land had rest for eighty years.
JUDG|3|31|After him was Shamgar the son of Anath, who killed 600 of the Philistines with an oxgoad, and he also saved Israel.
JUDG|4|1|And the people of Israel again did what was evil in the sight of the LORD after Ehud died.
JUDG|4|2|And the LORD sold them into the hand of Jabin king of Canaan, who reigned in Hazor. The commander of his army was Sisera, who lived in Harosheth-hagoyim.
JUDG|4|3|Then the people of Israel cried out to the LORD for help, for he had 900 chariots of iron and he oppressed the people of Israel cruelly for twenty years.
JUDG|4|4|Now Deborah, a prophetess, the wife of Lappidoth, was judging Israel at that time.
JUDG|4|5|She used to sit under the palm of Deborah between Ramah and Bethel in the hill country of Ephraim, and the people of Israel came up to her for judgment.
JUDG|4|6|She sent and summoned Barak the son of Abinoam from Kedesh-naphtali and said to him, "Has not the LORD, the God of Israel, commanded you, 'Go, gather your men at Mount Tabor, taking 10,000 from the people of Naphtali and the people of Zebulun.
JUDG|4|7|And I will draw out Sisera, the general of Jabin's army, to meet you by the river Kishon with his chariots and his troops, and I will give him into your hand'?"
JUDG|4|8|Barak said to her, "If you will go with me, I will go, but if you will not go with me, I will not go."
JUDG|4|9|And she said, "I will surely go with you. Nevertheless, the road on which you are going will not lead to your glory, for the LORD will sell Sisera into the hand of a woman." Then Deborah arose and went with Barak to Kedesh.
JUDG|4|10|And Barak called out Zebulun and Naphtali to Kedesh. And 10,000 men went up at his heels, and Deborah went up with him.
JUDG|4|11|Now Heber the Kenite had separated from the Kenites, the descendants of Hobab the father-in-law of Moses, and had pitched his tent as far away as the oak in Zaanannim, which is near Kedesh.
JUDG|4|12|When Sisera was told that Barak the son of Abinoam had gone up to Mount Tabor,
JUDG|4|13|Sisera called out all his chariots, 900 chariots of iron, and all the men who were with him, from Harosheth-hagoyim to the river Kishon.
JUDG|4|14|And Deborah said to Barak, "Up! For this is the day in which the LORD has given Sisera into your hand. Does not the LORD go out before you?" So Barak went down from Mount Tabor with 10,000 men following him.
JUDG|4|15|And the LORD routed Sisera and all his chariots and all his army before Barak by the edge of the sword. And Sisera got down from his chariot and fled away on foot.
JUDG|4|16|And Barak pursued the chariots and the army to Harosheth-hagoyim, and all the army of Sisera fell by the edge of the sword; not a man was left.
JUDG|4|17|But Sisera fled away on foot to the tent of Jael, the wife of Heber the Kenite, for there was peace between Jabin the king of Hazor and the house of Heber the Kenite.
JUDG|4|18|And Jael came out to meet Sisera and said to him, "Turn aside, my lord; turn aside to me; do not be afraid." So he turned aside to her into the tent, and she covered him with a rug.
JUDG|4|19|And he said to her, "Please give me a little water to drink, for I am thirsty." So she opened a skin of milk and gave him a drink and covered him.
JUDG|4|20|And he said to her, "Stand at the opening of the tent, and if any man comes and asks you, 'Is anyone here?' say, 'No.'"
JUDG|4|21|But Jael the wife of Heber took a tent peg, and took a hammer in her hand. Then she went softly to him and drove the peg into his temple until it went down into the ground while he was lying fast asleep from weariness. So he died.
JUDG|4|22|And behold, as Barak was pursuing Sisera, Jael went out to meet him and said to him, "Come, and I will show you the man whom you are seeking." So he went in to her tent, and there lay Sisera dead, with the tent peg in his temple.
JUDG|4|23|So on that day God subdued Jabin the king of Canaan before the people of Israel.
JUDG|4|24|And the hand of the people of Israel pressed harder and harder against Jabin the king of Canaan, until they destroyed Jabin king of Canaan.
JUDG|5|1|Then sang Deborah and Barak the son of Abinoam on that day:
JUDG|5|2|"That the leaders took the lead in Israel, that the people offered themselves willingly, bless the LORD!
JUDG|5|3|"Hear, O kings; give ear, O princes; to the LORD I will sing; I will make melody to the LORD, the God of Israel.
JUDG|5|4|"LORD, when you went out from Seir, when you marched from the region of Edom, the earth trembled and the heavens dropped, yes, the clouds dropped water.
JUDG|5|5|The mountains quaked before the LORD, even Sinai before the LORD, the God of Israel.
JUDG|5|6|"In the days of Shamgar, son of Anath, in the days of Jael, the highways were abandoned, and travelers kept to the byways.
JUDG|5|7|The villagers ceased in Israel; they ceased to be until I arose; I, Deborah, arose as a mother in Israel.
JUDG|5|8|When new gods were chosen, then war was in the gates. Was shield or spear to be seen among forty thousand in Israel?
JUDG|5|9|My heart goes out to the commanders of Israel who offered themselves willingly among the people. Bless the LORD.
JUDG|5|10|"Tell of it, you who ride on white donkeys, you who sit on rich carpets and you who walk by the way.
JUDG|5|11|To the sound of musicians at the watering places, there they repeat the righteous triumphs of the LORD, the righteous triumphs of his villagers in Israel. "Then down to the gates marched the people of the LORD.
JUDG|5|12|"Awake, awake, Deborah! Awake, awake, break out in a song! Arise, Barak, lead away your captives, O son of Abinoam.
JUDG|5|13|Then down marched the remnant of the noble; the people of the LORD marched down for me against the mighty.
JUDG|5|14|From Ephraim their root they marched down into the valley, following you, Benjamin, with your kinsmen; from Machir marched down the commanders, and from Zebulun those who bear the lieutenant's staff;
JUDG|5|15|the princes of Issachar came with Deborah, and Issachar faithful to Barak; into the valley they rushed at his heels. Among the clans of Reuben there were great searchings of heart.
JUDG|5|16|Why did you sit still among the sheepfolds, to hear the whistling for the flocks? Among the clans of Reuben there were great searchings of heart.
JUDG|5|17|Gilead stayed beyond the Jordan; and Dan, why did he stay with the ships? Asher sat still at the coast of the sea, staying by his landings.
JUDG|5|18|Zebulun is a people who risked their lives to the death; Naphtali, too, on the heights of the field.
JUDG|5|19|"The kings came, they fought; then fought the kings of Canaan, at Taanach, by the waters of Megiddo; they got no spoils of silver.
JUDG|5|20|From heaven the stars fought, from their courses they fought against Sisera.
JUDG|5|21|The torrent Kishon swept them away, the ancient torrent, the torrent Kishon. March on, my soul, with might!
JUDG|5|22|"Then loud beat the horses' hoofs with the galloping, galloping of his steeds.
JUDG|5|23|"Curse Meroz, says the angel of the LORD, curse its inhabitants thoroughly, because they did not come to the help of the LORD, to the help of the LORD against the mighty.
JUDG|5|24|"Most blessed of women be Jael, the wife of Heber the Kenite, of tent-dwelling women most blessed.
JUDG|5|25|He asked water and she gave him milk; she brought him curds in a noble's bowl.
JUDG|5|26|She sent her hand to the tent peg and her right hand to the workmen's mallet; she struck Sisera; she crushed his head; she shattered and pierced his temple.
JUDG|5|27|Between her feet he sank, he fell, he lay still; between her feet he sank, he fell; where he sank, there he fell- dead.
JUDG|5|28|"Out of the window she peered, the mother of Sisera wailed through the lattice: 'Why is his chariot so long in coming? Why tarry the hoofbeats of his chariots?'
JUDG|5|29|Her wisest princesses answer, indeed, she answers herself,
JUDG|5|30|'Have they not found and divided the spoil?- A womb or two for every man; spoil of dyed materials for Sisera, spoil of dyed materials embroidered, two pieces of dyed work embroidered for the neck as spoil?'
JUDG|5|31|"So may all your enemies perish, O LORD! But your friends be like the sun as he rises in his might." And the land had rest for forty years.
JUDG|6|1|The people of Israel did what was evil in the sight of the LORD, and the LORD gave them into the hand of Midian seven years.
JUDG|6|2|And the hand of Midian overpowered Israel, and because of Midian the people of Israel made for themselves the dens that are in the mountains and the caves and the strongholds.
JUDG|6|3|For whenever the Israelites planted crops, the Midianites and the Amalekites and the people of the East would come up against them.
JUDG|6|4|They would encamp against them and devour the produce of the land, as far as Gaza, and leave no sustenance in Israel and no sheep or ox or donkey.
JUDG|6|5|For they would come up with their livestock and their tents; they would come like locusts in number- both they and their camels could not be counted- so that they laid waste the land as they came in.
JUDG|6|6|And Israel was brought very low because of Midian. And the people of Israel cried out for help to the LORD.
JUDG|6|7|When the people of Israel cried out to the LORD on account of the Midianites,
JUDG|6|8|the LORD sent a prophet to the people of Israel. And he said to them, "Thus says the LORD, the God of Israel: I led you up from Egypt and brought you out of the house of bondage.
JUDG|6|9|And I delivered you from the hand of the Egyptians and from the hand of all who oppressed you, and drove them out before you and gave you their land.
JUDG|6|10|And I said to you, 'I am the LORD your God; you shall not fear the gods of the Amorites in whose land you dwell.' But you have not obeyed my voice."
JUDG|6|11|Now the angel of the LORD came and sat under the terebinth at Ophrah, which belonged to Joash the Abiezrite, while his son Gideon was beating out wheat in the winepress to hide it from the Midianites.
JUDG|6|12|And the angel of the LORD appeared to him and said to him, "The LORD is with you, O mighty man of valor."
JUDG|6|13|And Gideon said to him, "Please, sir, if the LORD is with us, why then has all this happened to us? And where are all his wonderful deeds that our fathers recounted to us, saying, 'Did not the LORD bring us up from Egypt?' But now the LORD has forsaken us and given us into the hand of Midian."
JUDG|6|14|And the LORD turned to him and said, "Go in this might of yours and save Israel from the hand of Midian; do not I send you?"
JUDG|6|15|And he said to him, "Please, Lord, how can I save Israel? Behold, my clan is the weakest in Manasseh, and I am the least in my father's house."
JUDG|6|16|And the LORD said to him, "But I will be with you, and you shall strike the Midianites as one man."
JUDG|6|17|And he said to him, "If now I have found favor in your eyes, then show me a sign that it is you who speaks with me.
JUDG|6|18|Please do not depart from here until I come to you and bring out my present and set it before you." And he said, "I will stay till you return."
JUDG|6|19|So Gideon went into his house and prepared a young goat and unleavened cakes from an ephah of flour. The meat he put in a basket, and the broth he put in a pot, and brought them to him under the terebinth and presented them.
JUDG|6|20|And the angel of God said to him, "Take the meat and the unleavened cakes, and put them on this rock, and pour the broth over them." And he did so.
JUDG|6|21|Then the angel of the LORD reached out the tip of the staff that was in his hand and touched the meat and the unleavened cakes. And fire sprang up from the rock and consumed the flesh and the unleavened cakes. And the angel of the LORD vanished from his sight.
JUDG|6|22|Then Gideon perceived that he was the angel of the LORD. And Gideon said, "Alas, O Lord GOD! For now I have seen the angel of the LORD face to face."
JUDG|6|23|But the LORD said to him, "Peace be to you. Do not fear; you shall not die."
JUDG|6|24|Then Gideon built an altar there to the LORD and called it, The LORD is Peace. To this day it still stands at Ophrah, which belongs to the Abiezrites.
JUDG|6|25|That night the LORD said to him, "Take your father's bull, and the second bull seven years old, and pull down the altar of Baal that your father has, and cut down the Asherah that is beside it
JUDG|6|26|and build an altar to the LORD your God on the top of the stronghold here, with stones laid in due order. Then take the second bull and offer it as a burnt offering with the wood of the Asherah that you shall cut down."
JUDG|6|27|So Gideon took ten men of his servants and did as the LORD had told him. But because he was too afraid of his family and the men of the town to do it by day, he did it by night.
JUDG|6|28|When the men of the town rose early in the morning, behold, the altar of Baal was broken down, and the Asherah beside it was cut down, and the second bull was offered on the altar that had been built.
JUDG|6|29|And they said to one another, "Who has done this thing?" And after they had searched and inquired, they said, "Gideon the son of Joash has done this thing."
JUDG|6|30|Then the men of the town said to Joash, "Bring out your son, that he may die, for he has broken down the altar of Baal and cut down the Asherah beside it."
JUDG|6|31|But Joash said to all who stood against him, "Will you contend for Baal? Or will you save him? Whoever contends for him shall be put to death by morning. If he is a god, let him contend for himself, because his altar has been broken down."
JUDG|6|32|Therefore on that day Gideon was called Jerubbaal, that is to say, "Let Baal contend against him," because he broke down his altar.
JUDG|6|33|Now all the Midianites and the Amalekites and the people of the East came together, and they crossed the Jordan and encamped in the Valley of Jezreel.
JUDG|6|34|But the Spirit of the LORD clothed Gideon, and he sounded the trumpet, and the Abiezrites were called out to follow him.
JUDG|6|35|And he sent messengers throughout all Manasseh, and they too were called out to follow him. And he sent messengers to Asher, Zebulun, and Naphtali, and they went up to meet them.
JUDG|6|36|Then Gideon said to God, "If you will save Israel by my hand, as you have said,
JUDG|6|37|behold, I am laying a fleece of wool on the threshing floor. If there is dew on the fleece alone, and it is dry on all the ground, then I shall know that you will save Israel by my hand, as you have said."
JUDG|6|38|And it was so. When he rose early next morning and squeezed the fleece, he wrung enough dew from the fleece to fill a bowl with water.
JUDG|6|39|Then Gideon said to God, "Let not your anger burn against me; let me speak just once more. Please let me test just once more with the fleece. Please let it be dry on the fleece only, and on all the ground let there be dew."
JUDG|6|40|And God did so that night; and it was dry on the fleece only, and on all the ground there was dew.
JUDG|7|1|Then Jerubbaal (that is, Gideon) and all the people who were with him rose early and encamped beside the spring of Harod. And the camp of Midian was north of them, by the hill of Moreh, in the valley.
JUDG|7|2|The LORD said to Gideon, "The people with you are too many for me to give the Midianites into their hand, lest Israel boast over me, saying, 'My own hand has saved me.'
JUDG|7|3|Now therefore proclaim in the ears of the people, saying, 'Whoever is fearful and trembling, let him return home and hurry away from Mount Gilead.'"Then 22,000 of the people returned, and 10,000 remained.
JUDG|7|4|And the LORD said to Gideon, "The people are still too many. Take them down to the water, and I will test them for you there, and anyone of whom I say to you, 'This one shall go with you,' shall go with you, and anyone of whom I say to you, 'This one shall not go with you,' shall not go."
JUDG|7|5|So he brought the people down to the water. And the LORD said to Gideon, "Every one who laps the water with his tongue, as a dog laps, you shall set by himself. Likewise, every one who kneels down to drink."
JUDG|7|6|And the number of those who lapped, putting their hands to their mouths, was 300 men, but all the rest of the people knelt down to drink water.
JUDG|7|7|And the LORD said to Gideon, "With the 300 men who lapped I will save you and give the Midianites into your hand, and let all the others go every man to his home."
JUDG|7|8|So the people took provisions in their hands, and their trumpets. And he sent all the rest of Israel every man to his tent, but retained the 300 men. And the camp of Midian was below him in the valley.
JUDG|7|9|That same night the LORD said to him, "Arise, go down against the camp, for I have given it into your hand.
JUDG|7|10|But if you are afraid to go down, go down to the camp with Purah your servant.
JUDG|7|11|And you shall hear what they say, and afterward your hands shall be strengthened to go down against the camp." Then he went down with Purah his servant to the outposts of the armed men who were in the camp.
JUDG|7|12|And the Midianites and the Amalekites and all the people of the East lay along the valley like locusts in abundance, and their camels were without number, as the sand that is on the seashore in abundance.
JUDG|7|13|When Gideon came, behold, a man was telling a dream to his comrade. And he said, "Behold, I dreamed a dream, and behold, a cake of barley bread tumbled into the camp of Midian and came to the tent and struck it so that it fell and turned it upside down, so that the tent lay flat."
JUDG|7|14|And his comrade answered, "This is no other than the sword of Gideon the son of Joash, a man of Israel; God has given into his hand Midian and all the camp."
JUDG|7|15|As soon as Gideon heard the telling of the dream and its interpretation, he worshiped. And he returned to the camp of Israel and said, "Arise, for the LORD has given the host of Midian into your hand."
JUDG|7|16|And he divided the 300 men into three companies and put trumpets into the hands of all of them and empty jars, with torches inside the jars.
JUDG|7|17|And he said to them, "Look at me, and do likewise. When I come to the outskirts of the camp, do as I do.
JUDG|7|18|When I blow the trumpet, I and all who are with me, then blow the trumpets also on every side of all the camp and shout, 'For the LORD and for Gideon.'"
JUDG|7|19|So Gideon and the hundred men who were with him came to the outskirts of the camp at the beginning of the middle watch, when they had just set the watch. And they blew the trumpets and smashed the jars that were in their hands.
JUDG|7|20|Then the three companies blew the trumpets and broke the jars. They held in their left hands the torches, and in their right hands the trumpets to blow. And they cried out, "A sword for the LORD and for Gideon!"
JUDG|7|21|Every man stood in his place around the camp, and all the army ran. They cried out and fled.
JUDG|7|22|When they blew the 300 trumpets, the LORD set every man's sword against his comrade and against all the army. And the army fled as far as Beth-shittah toward Zererah, as far as the border of Abel-meholah, by Tabbath.
JUDG|7|23|And the men of Israel were called out from Naphtali and from Asher and from all Manasseh, and they pursued after Midian.
JUDG|7|24|Gideon sent messengers throughout all the hill country of Ephraim, saying, "Come down against the Midianites and capture the waters against them, as far as Beth-barah, and also the Jordan." So all the men of Ephraim were called out, and they captured the waters as far as Beth-barah, and also the Jordan.
JUDG|7|25|And they captured the two princes of Midian, Oreb and Zeeb. They killed Oreb at the rock of Oreb, and Zeeb they killed at the winepress of Zeeb. Then they pursued Midian, and they brought the heads of Oreb and Zeeb to Gideon across the Jordan.
JUDG|8|1|Then the men of Ephraim said to him, "What is this that you have done to us, not to call us when you went to fight with Midian?" And they accused him fiercely.
JUDG|8|2|And he said to them, "What have I done now in comparison with you? Is not the gleaning of the grapes of Ephraim better than the grape harvest of Abiezer?
JUDG|8|3|God has given into your hands the princes of Midian, Oreb and Zeeb. What have I been able to do in comparison with you?" Then their anger against him subsided when he said this.
JUDG|8|4|And Gideon came to the Jordan and crossed over, he and the 300 men who were with him, exhausted yet pursuing.
JUDG|8|5|So he said to the men of Succoth, "Please give loaves of bread to the people who follow me, for they are exhausted, and I am pursuing after Zebah and Zalmunna, the kings of Midian."
JUDG|8|6|And the officials of Succoth said, "Are the hands of Zebah and Zalmunna already in your hand, that we should give bread to your army?"
JUDG|8|7|So Gideon said, "Well then, when the LORD has given Zebah and Zalmunna into my hand, I will flail your flesh with the thorns of the wilderness and with briers."
JUDG|8|8|And from there he went up to Penuel, and spoke to them in the same way, and the men of Penuel answered him as the men of Succoth had answered.
JUDG|8|9|And he said to the men of Penuel, "When I come again in peace, I will break down this tower."
JUDG|8|10|Now Zebah and Zalmunna were in Karkor with their army, about 15,000 men, all who were left of all the army of the people of the East, for there had fallen 120,000 men who drew the sword.
JUDG|8|11|And Gideon went up by the way of the tent dwellers east of Nobah and Jogbehah and attacked the army, for the army felt secure.
JUDG|8|12|And Zebah and Zalmunna fled, and he pursued them and captured the two kings of Midian, Zebah and Zalmunna, and he threw all the army into a panic.
JUDG|8|13|Then Gideon the son of Joash returned from the battle by the ascent of Heres.
JUDG|8|14|And he captured a young man of Succoth and questioned him. And he wrote down for him the officials and elders of Succoth, seventy-seven men.
JUDG|8|15|And he came to the men of Succoth and said, "Behold Zebah and Zalmunna, about whom you taunted me, saying, 'Are the hands of Zebah and Zalmunna already in your hand, that we should give bread to your men who are exhausted?'"
JUDG|8|16|And he took the elders of the city, and he took thorns of the wilderness and briers and with them taught the men of Succoth a lesson.
JUDG|8|17|And he broke down the tower of Penuel and killed the men of the city.
JUDG|8|18|Then he said to Zebah and Zalmunna, "Where are the men whom you killed at Tabor?" They answered, "As you are, so were they. Every one of them resembled the son of a king."
JUDG|8|19|And he said, "They were my brothers, the sons of my mother. As the LORD lives, if you had saved them alive, I would not kill you."
JUDG|8|20|So he said to Jether his firstborn, "Rise and kill them!" But the young man did not draw his sword, for he was afraid, because he was still a young man.
JUDG|8|21|Then Zebah and Zalmunna said, "Rise yourself and fall upon us, for as the man is, so is his strength." And Gideon arose and killed Zebah and Zalmunna, and he took the crescent ornaments that were on the necks of their camels.
JUDG|8|22|Then the men of Israel said to Gideon, "Rule over us, you and your son and your grandson also, for you have saved us from the hand of Midian."
JUDG|8|23|Gideon said to them, "I will not rule over you, and my son will not rule over you; the LORD will rule over you."
JUDG|8|24|And Gideon said to them, "Let me make a request of you: every one of you give me the earrings from his spoil." (For they had golden earrings, because they were Ishmaelites.)
JUDG|8|25|And they answered, "We will willingly give them." And they spread a cloak, and every man threw in it the earrings of his spoil.
JUDG|8|26|And the weight of the golden earrings that he requested was 1,700 shekels of gold, besides the crescent ornaments and the pendants and the purple garments worn by the kings of Midian, and besides the collars that were around the necks of their camels.
JUDG|8|27|And Gideon made an ephod of it and put it in his city, in Ophrah. And all Israel whored after it there, and it became a snare to Gideon and to his family.
JUDG|8|28|So Midian was subdued before the people of Israel, and they raised their heads no more. And the land had rest forty years in the days of Gideon.
JUDG|8|29|Jerubbaal the son of Joash went and lived in his own house.
JUDG|8|30|Now Gideon had seventy sons, his own offspring, for he had many wives.
JUDG|8|31|And his concubine who was in Shechem also bore him a son, and he called his name Abimelech.
JUDG|8|32|And Gideon the son of Joash died in a good old age and was buried in the tomb of Joash his father, at Ophrah of the Abiezrites.
JUDG|8|33|As soon as Gideon died, the people of Israel turned again and whored after the Baals and made Baal-berith their god.
JUDG|8|34|And the people of Israel did not remember the LORD their God, who had delivered them from the hand of all their enemies on every side,
JUDG|8|35|and they did not show steadfast love to the family of Jerubbaal (that is, Gideon) in return for all the good that he had done to Israel.
JUDG|9|1|Now Abimelech the son of Jerubbaal went to Shechem to his mother's relatives and said to them and to the whole clan of his mother's family,
JUDG|9|2|"Say in the ears of all the leaders of Shechem, 'Which is better for you, that all seventy of the sons of Jerubbaal rule over you, or that one rule over you?' Remember also that I am your bone and your flesh."
JUDG|9|3|And his mother's relatives spoke all these words on his behalf in the ears of all the leaders of Shechem, and their hearts inclined to follow Abimelech, for they said, "He is our brother."
JUDG|9|4|And they gave him seventy pieces of silver out of the house of Baal-berith with which Abimelech hired worthless and reckless fellows, who followed him.
JUDG|9|5|And he went to his father's house at Ophrah and killed his brothers the sons of Jerubbaal, seventy men, on one stone. But Jotham the youngest son of Jerubbaal was left, for he hid himself.
JUDG|9|6|And all the leaders of Shechem came together, and all Beth-millo, and they went and made Abimelech king, by the oak of the pillar at Shechem.
JUDG|9|7|When it was told to Jotham, he went and stood on top of Mount Gerizim and cried aloud and said to them, "Listen to me, you leaders of Shechem, that God may listen to you.
JUDG|9|8|The trees once went out to anoint a king over them, and they said to the olive tree, 'Reign over us.'
JUDG|9|9|But the olive tree said to them, 'Shall I leave my abundance, by which gods and men are honored, and go hold sway over the trees?'
JUDG|9|10|And the trees said to the fig tree, 'You come and reign over us.'
JUDG|9|11|But the fig tree said to them, 'Shall I leave my sweetness and my good fruit and go hold sway over the trees?'
JUDG|9|12|And the trees said to the vine, 'You come and reign over us.'
JUDG|9|13|But the vine said to them, 'Shall I leave my wine that cheers God and men and go hold sway over the trees?'
JUDG|9|14|Then all the trees said to the bramble, 'You come and reign over us.'
JUDG|9|15|And the bramble said to the trees, 'If in good faith you are anointing me king over you, then come and take refuge in my shade, but if not, let fire come out of the bramble and devour the cedars of Lebanon.'
JUDG|9|16|"Now therefore, if you acted in good faith and integrity when you made Abimelech king, and if you have dealt well with Jerubbaal and his house and have done to him as his deeds deserved-
JUDG|9|17|for my father fought for you and risked his life and delivered you from the hand of Midian,
JUDG|9|18|and you have risen up against my father's house this day and have killed his sons, seventy men on one stone, and have made Abimelech, the son of his female servant, king over the leaders of Shechem, because he is your relative-
JUDG|9|19|if you then have acted in good faith and integrity with Jerubbaal and with his house this day, then rejoice in Abimelech, and let him also rejoice in you.
JUDG|9|20|But if not, let fire come out from Abimelech and devour the leaders of Shechem and Beth-millo; and let fire come out from the leaders of Shechem and from Beth-millo and devour Abimelech."
JUDG|9|21|And Jotham ran away and fled and went to Beer and lived there, because of Abimelech his brother.
JUDG|9|22|Abimelech ruled over Israel three years.
JUDG|9|23|And God sent an evil spirit between Abimelech and the leaders of Shechem, and the leaders of Shechem dealt treacherously with Abimelech,
JUDG|9|24|that the violence done to the seventy sons of Jerubbaal might come, and their blood be laid on Abimelech their brother, who killed them, and on the men of Shechem, who strengthened his hands to kill his brothers.
JUDG|9|25|And the leaders of Shechem put men in ambush against him on the mountaintops, and they robbed all who passed by them along that way. And it was told to Abimelech.
JUDG|9|26|And Gaal the son of Ebed moved into Shechem with his relatives, and the leaders of Shechem put confidence in him.
JUDG|9|27|And they went out into the field and gathered the grapes from their vineyards and trod them and held a festival; and they went into the house of their god and ate and drank and reviled Abimelech.
JUDG|9|28|And Gaal the son of Ebed said, "Who is Abimelech, and who are we of Shechem, that we should serve him? Is he not the son of Jerubbaal, and is not Zebul his officer? Serve the men of Hamor the father of Shechem; but why should we serve him?
JUDG|9|29|Would that this people were under my hand! Then I would remove Abimelech. I would say to Abimelech, 'Increase your army, and come out.'"
JUDG|9|30|When Zebul the ruler of the city heard the words of Gaal the son of Ebed, his anger was kindled.
JUDG|9|31|And he sent messengers to Abimelech secretly, saying, "Behold, Gaal the son of Ebed and his relatives have come to Shechem, and they are stirring up the city against you.
JUDG|9|32|Now therefore, go by night, you and the people who are with you, and set an ambush in the field.
JUDG|9|33|Then in the morning, as soon as the sun is up, rise early and rush upon the city. And when he and the people who are with him come out against you, you may do to them as your hand finds to do."
JUDG|9|34|So Abimelech and all the men who were with him rose up by night and set an ambush against Shechem in four companies.
JUDG|9|35|And Gaal the son of Ebed went out and stood in the entrance of the gate of the city, and Abimelech and the people who were with him rose from the ambush.
JUDG|9|36|And when Gaal saw the people, he said to Zebul, "Look, people are coming down from the mountaintops!" And Zebul said to him, "You mistake the shadow of the mountains for men."
JUDG|9|37|Gaal spoke again and said, "Look, people are coming down from the center of the land, and one company is coming from the direction of the Diviners' Oak."
JUDG|9|38|Then Zebul said to him, "Where is your mouth now, you who said, 'Who is Abimelech, that we should serve him?' Are not these the people whom you despised? Go out now and fight with them."
JUDG|9|39|And Gaal went out at the head of the leaders of Shechem and fought with Abimelech.
JUDG|9|40|And Abimelech chased him, and he fled before him. And many fell wounded, up to the entrance of the gate.
JUDG|9|41|And Abimelech lived at Arumah, and Zebul drove out Gaal and his relatives, so that they could not dwell at Shechem.
JUDG|9|42|On the following day, the people went out into the field, and Abimelech was told.
JUDG|9|43|He took his people and divided them into three companies and set an ambush in the fields. And he looked and saw the people coming out of the city. So he rose against them and killed them.
JUDG|9|44|Abimelech and the company that was with him rushed forward and stood at the entrance of the gate of the city, while the two companies rushed upon all who were in the field and killed them.
JUDG|9|45|And Abimelech fought against the city all that day. He captured the city and killed the people who were in it, and he razed the city and sowed it with salt.
JUDG|9|46|When all the leaders of the Tower of Shechem heard of it, they entered the stronghold of the house of El-berith.
JUDG|9|47|Abimelech was told that all the leaders of the Tower of Shechem were gathered together.
JUDG|9|48|And Abimelech went up to Mount Zalmon, he and all the people who were with him. And Abimelech took an axe in his hand and cut down a bundle of brushwood and took it up and laid it on his shoulder. And he said to the men who were with him, "What you have seen me do, hurry and do as I have done."
JUDG|9|49|So every one of the people cut down his bundle and following Abimelech put it against the stronghold, and they set the stronghold on fire over them, so that all the people of the Tower of Shechem also died, about 1,000 men and women.
JUDG|9|50|Then Abimelech went to Thebez and encamped against Thebez and captured it.
JUDG|9|51|But there was a strong tower within the city, and all the men and women and all the leaders of the city fled to it and shut themselves in, and they went up to the roof of the tower.
JUDG|9|52|And Abimelech came to the tower and fought against it and drew near to the door of the tower to burn it with fire.
JUDG|9|53|And a certain woman threw an upper millstone on Abimelech's head and crushed his skull.
JUDG|9|54|Then he called quickly to the young man his armor-bearer and said to him, "Draw your sword and kill me, lest they say of me, 'A woman killed him.'" And his young man thrust him through, and he died.
JUDG|9|55|And when the men of Israel saw that Abimelech was dead, everyone departed to his home.
JUDG|9|56|Thus God returned the evil of Abimelech, which he committed against his father in killing his seventy brothers.
JUDG|9|57|And God also made all the evil of the men of Shechem return on their heads, and upon them came the curse of Jotham the son of Jerubbaal.
JUDG|10|1|After Abimelech there arose to save Israel Tola the son of Puah, son of Dodo, a man of Issachar, and he lived at Shamir in the hill country of Ephraim.
JUDG|10|2|And he judged Israel twenty-three years. Then he died and was buried at Shamir.
JUDG|10|3|After him arose Jair the Gileadite, who judged Israel twenty-two years.
JUDG|10|4|And he had thirty sons who rode on thirty donkeys, and they had thirty cities, called Havvoth-jair to this day, which are in the land of Gilead.
JUDG|10|5|And Jair died and was buried in Kamon.
JUDG|10|6|The people of Israel again did what was evil in the sight of the LORD and served the Baals and the Ashtaroth, the gods of Syria, the gods of Sidon, the gods of Moab, the gods of the Ammonites, and the gods of the Philistines. And they forsook the LORD and did not serve him.
JUDG|10|7|So the anger of the LORD was kindled against Israel, and he sold them into the hand of the Philistines and into the hand of the Ammonites,
JUDG|10|8|and they crushed and oppressed the people of Israel that year. For eighteen years they oppressed all the people of Israel who were beyond the Jordan in the land of the Amorites, which is in Gilead.
JUDG|10|9|And the Ammonites crossed the Jordan to fight also against Judah and against Benjamin and against the house of Ephraim, so that Israel was severely distressed.
JUDG|10|10|And the people of Israel cried out to the LORD, saying, "We have sinned against you, because we have forsaken our God and have served the Baals."
JUDG|10|11|And the LORD said to the people of Israel, "Did I not save you from the Egyptians and from the Amorites, from the Ammonites and from the Philistines?
JUDG|10|12|The Sidonians also, and the Amalekites and the Maonites oppressed you, and you cried out to me, and I saved you out of their hand.
JUDG|10|13|Yet you have forsaken me and served other gods; therefore I will save you no more.
JUDG|10|14|Go and cry out to the gods whom you have chosen; let them save you in the time of your distress."
JUDG|10|15|And the people of Israel said to the LORD, "We have sinned; do to us whatever seems good to you. Only please deliver us this day."
JUDG|10|16|So they put away the foreign gods from among them and served the LORD, and he became impatient over the misery of Israel.
JUDG|10|17|Then the Ammonites were called to arms, and they encamped in Gilead. And the people of Israel came together, and they encamped at Mizpah.
JUDG|10|18|And the people, the leaders of Gilead, said one to another, "Who is the man who will begin to fight against the Ammonites? He shall be head over all the inhabitants of Gilead."
JUDG|11|1|Now Jephthah the Gileadite was a mighty warrior, but he was the son of a prostitute. Gilead was the father of Jephthah.
JUDG|11|2|And Gilead's wife also bore him sons. And when his wife's sons grew up, they drove Jephthah out and said to him, "You shall not have an inheritance in our father's house, for you are the son of another woman."
JUDG|11|3|Then Jephthah fled from his brothers and lived in the land of Tob, and worthless fellows collected around Jephthah and went out with him.
JUDG|11|4|After a time the Ammonites made war against Israel.
JUDG|11|5|And when the Ammonites made war against Israel, the elders of Gilead went to bring Jephthah from the land of Tob.
JUDG|11|6|And they said to Jephthah, "Come and be our leader, that we may fight with the Ammonites."
JUDG|11|7|But Jephthah said to the elders of Gilead, "Did you not hate me and drive me out of my father's house? Why have you come to me now when you are in distress?"
JUDG|11|8|And the elders of Gilead said to Jephthah, "That is why we have turned to you now, that you may go with us and fight with the Ammonites and be our head over all the inhabitants of Gilead."
JUDG|11|9|Jephthah said to the elders of Gilead, "If you bring me home again to fight with the Ammonites, and the LORD gives them over to me, I will be your head."
JUDG|11|10|And the elders of Gilead said to Jephthah, "The LORD will be witness between us, if we do not do as you say."
JUDG|11|11|So Jephthah went with the elders of Gilead, and the people made him head and leader over them. And Jephthah spoke all his words before the LORD at Mizpah.
JUDG|11|12|Then Jephthah sent messengers to the king of the Ammonites and said, "What do you have against me, that you have come to me to fight against my land?"
JUDG|11|13|And the king of the Ammonites answered the messengers of Jephthah, "Because Israel on coming up from Egypt took away my land, from the Arnon to the Jabbok and to the Jordan; now therefore restore it peaceably."
JUDG|11|14|Jephthah again sent messengers to the king of the Ammonites
JUDG|11|15|and said to him, "Thus says Jephthah: Israel did not take away the land of Moab or the land of the Ammonites,
JUDG|11|16|but when they came up from Egypt, Israel went through the wilderness to the Red Sea and came to Kadesh.
JUDG|11|17|Israel then sent messengers to the king of Edom, saying, 'Please let us pass through your land,' but the king of Edom would not listen. And they sent also to the king of Moab, but he would not consent. So Israel remained at Kadesh.
JUDG|11|18|"Then they journeyed through the wilderness and went around the land of Edom and the land of Moab and arrived on the east side of the land of Moab and camped on the other side of the Arnon. But they did not enter the territory of Moab, for the Arnon was the boundary of Moab.
JUDG|11|19|Israel then sent messengers to Sihon king of the Amorites, king of Heshbon, and Israel said to him, 'Please let us pass through your land to our country,'
JUDG|11|20|but Sihon did not trust Israel to pass through his territory, so Sihon gathered all his people together and encamped at Jahaz and fought with Israel.
JUDG|11|21|And the LORD, the God of Israel, gave Sihon and all his people into the hand of Israel, and they defeated them. So Israel took possession of all the land of the Amorites, who inhabited that country.
JUDG|11|22|And they took possession of all the territory of the Amorites from the Arnon to the Jabbok and from the wilderness to the Jordan.
JUDG|11|23|So then the LORD, the God of Israel, dispossessed the Amorites from before his people Israel; and are you to take possession of them?
JUDG|11|24|Will you not possess what Chemosh your god gives you to possess? And all that the LORD our God has dispossessed before us, we will possess.
JUDG|11|25|Now are you any better than Balak the son of Zippor, king of Moab? Did he ever contend against Israel, or did he ever go to war with them?
JUDG|11|26|While Israel lived in Heshbon and its villages, and in Aroer and its villages, and in all the cities that are on the banks of the Arnon, 300 years, why did you not deliver them within that time?
JUDG|11|27|I therefore have not sinned against you, and you do me wrong by making war on me. The LORD, the Judge, decide this day between the people of Israel and the people of Ammon."
JUDG|11|28|But the king of the Ammonites did not listen to the words of Jephthah that he sent to him.
JUDG|11|29|Then the Spirit of the LORD was upon Jephthah, and he passed through Gilead and Manasseh and passed on to Mizpah of Gilead, and from Mizpah of Gilead he passed on to the Ammonites.
JUDG|11|30|And Jephthah made a vow to the LORD and said, "If you will give the Ammonites into my hand,
JUDG|11|31|then whatever comes out from the doors of my house to meet me when I return in peace from the Ammonites shall be the LORD's, and I will offer it up for a burnt offering."
JUDG|11|32|So Jephthah crossed over to the Ammonites to fight against them, and the LORD gave them into his hand.
JUDG|11|33|And he struck them from Aroer to the neighborhood of Minnith, twenty cities, and as far as Abel-keramim, with a great blow. So the Ammonites were subdued before the people of Israel.
JUDG|11|34|Then Jephthah came to his home at Mizpah. And behold, his daughter came out to meet him with tambourines and with dances. She was his only child; beside her he had neither son nor daughter.
JUDG|11|35|And as soon as he saw her, he tore his clothes and said, "Alas, my daughter! You have brought me very low, and you have become the cause of great trouble to me. For I have opened my mouth to the LORD, and I cannot take back my vow."
JUDG|11|36|And she said to him, "My father, you have opened your mouth to the LORD; do to me according to what has gone out of your mouth, now that the LORD has avenged you on your enemies, on the Ammonites."
JUDG|11|37|So she said to her father, "Let this thing be done for me: leave me alone two months, that I may go up and down on the mountains and weep for my virginity, I and my companions."
JUDG|11|38|So he said, "Go." Then he sent her away for two months, and she departed, she and her companions, and wept for her virginity on the mountains.
JUDG|11|39|And at the end of two months, she returned to her father, who did with her according to his vow that he had made. She had never known a man, and it became a custom in Israel
JUDG|11|40|that the daughters of Israel went year by year to lament the daughter of Jephthah the Gileadite four days in the year.
JUDG|12|1|The men of Ephraim were called to arms, and they crossed to Zaphon and said to Jephthah, "Why did you cross over to fight against the Ammonites and did not call us to go with you? We will burn your house over you with fire."
JUDG|12|2|And Jephthah said to them, "I and my people had a great dispute with the Ammonites, and when I called you, you did not save me from their hand.
JUDG|12|3|And when I saw that you would not save me, I took my life in my hand and crossed over against the Ammonites, and the LORD gave them into my hand. Why then have you come up to me this day to fight against me?"
JUDG|12|4|Then Jephthah gathered all the men of Gilead and fought with Ephraim. And the men of Gilead struck Ephraim, because they said, "You are fugitives of Ephraim, you Gileadites, in the midst of Ephraim and Manasseh."
JUDG|12|5|And the Gileadites captured the fords of the Jordan against the Ephraimites. And when any of the fugitives of Ephraim said, "Let me go over," the men of Gilead said to him, "Are you an Ephraimite?" When he said, "No,"
JUDG|12|6|they said to him, "Then say Shibboleth," and he said, "Sibboleth," for he could not pronounce it right. Then they seized him and slaughtered him at the fords of the Jordan. At that time 42,000 of the Ephraimites fell.
JUDG|12|7|Jephthah judged Israel six years. Then Jephthah the Gileadite died and was buried in his city in Gilead.
JUDG|12|8|After him Ibzan of Bethlehem judged Israel.
JUDG|12|9|He had thirty sons, and thirty daughters he gave in marriage outside his clan, and thirty daughters he brought in from outside for his sons. And he judged Israel seven years.
JUDG|12|10|Then Ibzan died and was buried at Bethlehem.
JUDG|12|11|After him Elon the Zebulunite judged Israel, and he judged Israel ten years.
JUDG|12|12|Then Elon the Zebulunite died and was buried at Aijalon in the land of Zebulun.
JUDG|12|13|After him Abdon the son of Hillel the Pirathonite judged Israel.
JUDG|12|14|He had forty sons and thirty grandsons, who rode on seventy donkeys, and he judged Israel eight years.
JUDG|12|15|Then Abdon the son of Hillel the Pirathonite died and was buried at Pirathon in the land of Ephraim, in the hill country of the Amalekites.
JUDG|13|1|And the people of Israel again did what was evil in the sight of the LORD, so the LORD gave them into the hand of the Philistines for forty years.
JUDG|13|2|There was a certain man of Zorah, of the tribe of the Danites, whose name was Manoah. And his wife was barren and had no children.
JUDG|13|3|And the angel of the LORD appeared to the woman and said to her, "Behold, you are barren and have not borne children, but you shall conceive and bear a son.
JUDG|13|4|Therefore be careful and drink no wine or strong drink, and eat nothing unclean,
JUDG|13|5|for behold, you shall conceive and bear a son. No razor shall come upon his head, for the child shall be a Nazirite to God from the womb, and he shall begin to save Israel from the hand of the Philistines."
JUDG|13|6|Then the woman came and told her husband, "A man of God came to me, and his appearance was like the appearance of the angel of God, very awesome. I did not ask him where he was from, and he did not tell me his name,
JUDG|13|7|but he said to me, 'Behold, you shall conceive and bear a son. So then drink no wine or strong drink, and eat nothing unclean, for the child shall be a Nazirite to God from the womb to the day of his death.'"
JUDG|13|8|Then Manoah prayed to the LORD and said, "O Lord, please let the man of God whom you sent come again to us and teach us what we are to do with the child who will be born."
JUDG|13|9|And God listened to the voice of Manoah, and the angel of God came again to the woman as she sat in the field. But Manoah her husband was not with her.
JUDG|13|10|So the woman ran quickly and told her husband, "Behold, the man who came to me the other day has appeared to me."
JUDG|13|11|And Manoah arose and went after his wife and came to the man and said to him, "Are you the man who spoke to this woman?" And he said, "I am."
JUDG|13|12|And Manoah said, "Now when your words come true, what is to be the child's manner of life, and what is his mission?"
JUDG|13|13|And the angel of the LORD said to Manoah, "Of all that I said to the woman let her be careful.
JUDG|13|14|She may not eat of anything that comes from the vine, neither let her drink wine or strong drink, or eat any unclean thing. All that I commanded her let her observe."
JUDG|13|15|Manoah said to the angel of the LORD, "Please let us detain you and prepare a young goat for you."
JUDG|13|16|And the angel of the LORD said to Manoah, "If you detain me, I will not eat of your food. But if you prepare a burnt offering, then offer it to the LORD." (For Manoah did not know that he was the angel of the LORD.)
JUDG|13|17|And Manoah said to the angel of the LORD, "What is your name, so that, when your words come true, we may honor you?"
JUDG|13|18|And the angel of the LORD said to him, "Why do you ask my name, seeing it is wonderful?"
JUDG|13|19|So Manoah took the young goat with the grain offering, and offered it on the rock to the LORD, to the one who works wonders, and Manoah and his wife were watching.
JUDG|13|20|And when the flame went up toward heaven from the altar, the angel of the LORD went up in the flame of the altar. Now Manoah and his wife were watching, and they fell on their faces to the ground.
JUDG|13|21|The angel of the LORD appeared no more to Manoah and to his wife. Then Manoah knew that he was the angel of the LORD.
JUDG|13|22|And Manoah said to his wife, "We shall surely die, for we have seen God."
JUDG|13|23|But his wife said to him, "If the LORD had meant to kill us, he would not have accepted a burnt offering and a grain offering at our hands, or shown us all these things, or now announced to us such things as these."
JUDG|13|24|And the woman bore a son and called his name Samson. And the young man grew, and the LORD blessed him.
JUDG|13|25|And the Spirit of the LORD began to stir him in Mahaneh-dan, between Zorah and Eshtaol.
JUDG|14|1|Samson went down to Timnah, and at Timnah he saw one of the daughters of the Philistines.
JUDG|14|2|Then he came up and told his father and mother, "I saw one of the daughters of the Philistines at Timnah. Now get her for me as my wife."
JUDG|14|3|But his father and mother said to him, "Is there not a woman among the daughters of your relatives, or among all our people, that you must go to take a wife from the uncircumcised Philistines?" But Samson said to his father, "Get her for me, for she is right in my eyes."
JUDG|14|4|His father and mother did not know that it was from the LORD, for he was seeking an opportunity against the Philistines. At that time the Philistines ruled over Israel.
JUDG|14|5|Then Samson went down with his father and mother to Timnah, and they came to the vineyards of Timnah. And behold, a young lion came toward him roaring.
JUDG|14|6|Then the Spirit of the LORD rushed upon him, and although he had nothing in his hand, he tore the lion in pieces as one tears a young goat. But he did not tell his father or his mother what he had done.
JUDG|14|7|Then he went down and talked with the woman, and she was right in Samson's eyes.
JUDG|14|8|After some days he returned to take her. And he turned aside to see the carcass of the lion, and behold, there was a swarm of bees in the body of the lion, and honey.
JUDG|14|9|He scraped it out into his hands and went on, eating as he went. And he came to his father and mother and gave some to them, and they ate. But he did not tell them that he had scraped the honey from the carcass of the lion.
JUDG|14|10|His father went down to the woman, and Samson prepared a feast there, for so the young men used to do.
JUDG|14|11|As soon as the people saw him, they brought thirty companions to be with him.
JUDG|14|12|And Samson said to them, "Let me now put a riddle to you. If you can tell me what it is, within the seven days of the feast, and find it out, then I will give you thirty linen garments and thirty changes of clothes,
JUDG|14|13|but if you cannot tell me what it is, then you shall give me thirty linen garments and thirty changes of clothes." And they said to him, "Put your riddle, that we may hear it."
JUDG|14|14|And he said to them, "Out of the eater came something to eat. Out of the strong came something sweet." And in three days they could not solve the riddle.
JUDG|14|15|On the fourth day they said to Samson's wife, "Entice your husband to tell us what the riddle is, lest we burn you and your father's house with fire. Have you invited us here to impoverish us?"
JUDG|14|16|And Samson's wife wept over him and said, "You only hate me; you do not love me. You have put a riddle to my people, and you have not told me what it is." And he said to her, "Behold, I have not told my father nor my mother, and shall I tell you?"
JUDG|14|17|She wept before him the seven days that their feast lasted, and on the seventh day he told her, because she pressed him hard. Then she told the riddle to her people.
JUDG|14|18|And the men of the city said to him on the seventh day before the sun went down, "What is sweeter than honey? What is stronger than a lion?" And he said to them, "If you had not plowed with my heifer, you would not have found out my riddle."
JUDG|14|19|And the Spirit of the LORD rushed upon him, and he went down to Ashkelon and struck down thirty men of the town and took their spoil and gave the garments to those who had told the riddle. In hot anger he went back to his father's house.
JUDG|14|20|And Samson's wife was given to his companion, who had been his best man.
JUDG|15|1|After some days, at the time of wheat harvest, Samson went to visit his wife with a young goat. And he said, "I will go in to my wife in the chamber." But her father would not allow him to go in.
JUDG|15|2|And her father said, "I really thought that you utterly hated her, so I gave her to your companion. Is not her younger sister more beautiful than she? Please take her instead."
JUDG|15|3|And Samson said to them, "This time I shall be innocent in regard to the Philistines, when I do them harm."
JUDG|15|4|So Samson went and caught 300 foxes and took torches. And he turned them tail to tail and put a torch between each pair of tails.
JUDG|15|5|And when he had set fire to the torches, he let the foxes go into the standing grain of the Philistines and set fire to the stacked grain and the standing grain, as well as the olive orchards.
JUDG|15|6|Then the Philistines said, "Who has done this?" And they said, "Samson, the son-in-law of the Timnite, because he has taken his wife and given her to his companion." And the Philistines came up and burned her and her father with fire.
JUDG|15|7|And Samson said to them, "If this is what you do, I swear I will be avenged on you, and after that I will quit."
JUDG|15|8|And he struck them hip and thigh with a great blow, and he went down and stayed in the cleft of the rock of Etam.
JUDG|15|9|Then the Philistines came up and encamped in Judah and made a raid on Lehi.
JUDG|15|10|And the men of Judah said, "Why have you come up against us?" They said, "We have come up to bind Samson, to do to him as he did to us."
JUDG|15|11|Then 3,000 men of Judah went down to the cleft of the rock of Etam, and said to Samson, "Do you not know that the Philistines are rulers over us? What then is this that you have done to us?" And he said to them, "As they did to me, so have I done to them."
JUDG|15|12|And they said to him, "We have come down to bind you, that we may give you into the hands of the Philistines." And Samson said to them, "Swear to me that you will not attack me yourselves."
JUDG|15|13|They said to him, "No; we will only bind you and give you into their hands. We will surely not kill you." So they bound him with two new ropes and brought him up from the rock.
JUDG|15|14|When he came to Lehi, the Philistines came shouting to meet him. Then the Spirit of the LORD rushed upon him, and the ropes that were on his arms became as flax that has caught fire, and his bonds melted off his hands.
JUDG|15|15|And he found a fresh jawbone of a donkey, and put out his hand and took it, and with it he struck 1,000 men.
JUDG|15|16|And Samson said, "With the jawbone of a donkey, heaps upon heaps, with the jawbone of a donkey have I struck down a thousand men."
JUDG|15|17|As soon as he had finished speaking, he threw away the jawbone out of his hand. And that place was called Ramath-lehi.
JUDG|15|18|And he was very thirsty, and he called upon the LORD and said, "You have granted this great salvation by the hand of your servant, and shall I now die of thirst and fall into the hands of the uncircumcised?"
JUDG|15|19|And God split open the hollow place that is at Lehi, and water came out from it. And when he drank, his spirit returned, and he revived. Therefore the name of it was called En-hakkore; it is at Lehi to this day.
JUDG|15|20|And he judged Israel in the days of the Philistines twenty years.
JUDG|16|1|Samson went to Gaza, and there he saw a prostitute, and he went in to her.
JUDG|16|2|The Gazites were told, "Samson has come here." And they surrounded the place and set an ambush for him all night at the gate of the city. They kept quiet all night, saying, "Let us wait till the light of the morning; then we will kill him."
JUDG|16|3|But Samson lay till midnight, and at midnight he arose and took hold of the doors of the gate of the city and the two posts, and pulled them up, bar and all, and put them on his shoulders and carried them to the top of the hill that is in front of Hebron.
JUDG|16|4|After this he loved a woman in the Valley of Sorek, whose name was Delilah.
JUDG|16|5|And the lords of the Philistines came up to her and said to her, "Seduce him, and see where his great strength lies, and by what means we may overpower him, that we may bind him to humble him. And we will each give you 1,100 pieces of silver."
JUDG|16|6|So Delilah said to Samson, "Please tell me where your great strength lies, and how you might be bound, that one could subdue you."
JUDG|16|7|Samson said to her, "If they bind me with seven fresh bowstrings that have not been dried, then I shall become weak and be like any other man."
JUDG|16|8|Then the lords of the Philistines brought up to her seven fresh bowstrings that had not been dried, and she bound him with them.
JUDG|16|9|Now she had men lying in ambush in an inner chamber. And she said to him, "The Philistines are upon you, Samson!" But he snapped the bowstrings, as a thread of flax snaps when it touches the fire. So the secret of his strength was not known.
JUDG|16|10|Then Delilah said to Samson, "Behold, you have mocked me and told me lies. Please tell me how you might be bound."
JUDG|16|11|And he said to her, "If they bind me with new ropes that have not been used, then I shall become weak and be like any other man."
JUDG|16|12|So Delilah took new ropes and bound him with them and said to him, "The Philistines are upon you, Samson!" And the men lying in ambush were in an inner chamber. But he snapped the ropes off his arms like a thread.
JUDG|16|13|Then Delilah said to Samson, "Until now you have mocked me and told me lies. Tell me how you might be bound." And he said to her, "If you weave the seven locks of my head with the web and fasten it tight with the pin, then I shall become weak and be like any other man."
JUDG|16|14|So while he slept, Delilah took the seven locks of his head and wove them into the web. And she made them tight with the pin and said to him, "The Philistines are upon you, Samson!" But he awoke from his sleep and pulled away the pin, the loom, and the web.
JUDG|16|15|And she said to him, "How can you say, 'I love you,' when your heart is not with me? You have mocked me these three times, and you have not told me where your great strength lies."
JUDG|16|16|And when she pressed him hard with her words day after day, and urged him, his soul was vexed to death.
JUDG|16|17|And he told her all his heart, and said to her, "A razor has never come upon my head, for I have been a Nazirite to God from my mother's womb. If my head is shaved, then my strength will leave me, and I shall become weak and be like any other man."
JUDG|16|18|When Delilah saw that he had told her all his heart, she sent and called the lords of the Philistines, saying, "Come up again, for he has told me all his heart." Then the lords of the Philistines came up to her and brought the money in their hands.
JUDG|16|19|She made him sleep on her knees. And she called a man and had him shave off the seven locks of his head. Then she began to torment him, and his strength left him.
JUDG|16|20|And she said, "The Philistines are upon you, Samson!" And he awoke from his sleep and said, "I will go out as at other times and shake myself free." But he did not know that the LORD had left him.
JUDG|16|21|And the Philistines seized him and gouged out his eyes and brought him down to Gaza and bound him with bronze shackles. And he ground at the mill in the prison.
JUDG|16|22|But the hair of his head began to grow again after it had been shaved.
JUDG|16|23|Now the lords of the Philistines gathered to offer a great sacrifice to Dagon their god and to rejoice, and they said, "Our god has given Samson our enemy into our hand."
JUDG|16|24|And when the people saw him, they praised their god. For they said, "Our god has given our enemy into our hand, the ravager of our country, who has killed many of us."
JUDG|16|25|And when their hearts were merry, they said, "Call Samson, that he may entertain us." So they called Samson out of the prison, and he entertained them. They made him stand between the pillars.
JUDG|16|26|And Samson said to the young man who held him by the hand, "Let me feel the pillars on which the house rests, that I may lean against them."
JUDG|16|27|Now the house was full of men and women. All the lords of the Philistines were there, and on the roof there were about 3,000 men and women, who looked on while Samson entertained.
JUDG|16|28|Then Samson called to the LORD and said, "O Lord GOD, please remember me and please strengthen me only this once, O God, that I may be avenged on the Philistines for my two eyes."
JUDG|16|29|And Samson grasped the two middle pillars on which the house rested, and he leaned his weight against them, his right hand on the one and his left hand on the other.
JUDG|16|30|And Samson said, "Let me die with the Philistines." Then he bowed with all his strength, and the house fell upon the lords and upon all the people who were in it. So the dead whom he killed at his death were more than those whom he had killed during his life.
JUDG|16|31|Then his brothers and all his family came down and took him and brought him up and buried him between Zorah and Eshtaol in the tomb of Manoah his father. He had judged Israel twenty years.
JUDG|17|1|There was a man of the hill country of Ephraim, whose name was Micah.
JUDG|17|2|And he said to his mother, "The 1,100 pieces of silver that were taken from you, about which you uttered a curse, and also spoke it in my ears, behold, the silver is with me; I took it." And his mother said, "Blessed be my son by the LORD."
JUDG|17|3|And he restored the 1,100 pieces of silver to his mother. And his mother said, "I dedicate the silver to the LORD from my hand for my son, to make a carved image and a metal image. Now therefore I will restore it to you."
JUDG|17|4|So when he restored the money to his mother, his mother took 200 pieces of silver and gave it to the silversmith, who made it into a carved image and a metal image. And it was in the house of Micah.
JUDG|17|5|And the man Micah had a shrine, and he made an ephod and household gods, and ordained one of his sons, who became his priest.
JUDG|17|6|In those days there was no king in Israel. Everyone did what was right in his own eyes.
JUDG|17|7|Now there was a young man of Bethlehem in Judah, of the family of Judah, who was a Levite, and he sojourned there.
JUDG|17|8|And the man departed from the town of Bethlehem in Judah to sojourn where he could find a place. And as he journeyed, he came to the hill country of Ephraim to the house of Micah.
JUDG|17|9|And Micah said to him, "Where do you come from?" And he said to him, "I am a Levite of Bethlehem in Judah, and I am going to sojourn where I may find a place."
JUDG|17|10|And Micah said to him, "Stay with me, and be to me a father and a priest, and I will give you ten pieces of silver a year and a suit of clothes and your living." And the Levite went in.
JUDG|17|11|And the Levite was content to dwell with the man, and the young man became to him like one of his sons.
JUDG|17|12|And Micah ordained the Levite, and the young man became his priest, and was in the house of Micah.
JUDG|17|13|Then Micah said, "Now I know that the LORD will prosper me, because I have a Levite as priest."
JUDG|18|1|In those days there was no king in Israel. And in those days the tribe of the people of Dan was seeking for itself an inheritance to dwell in, for until then no inheritance among the tribes of Israel had fallen to them.
JUDG|18|2|So the people of Dan sent five able men from the whole number of their tribe, from Zorah and from Eshtaol, to spy out the land and to explore it. And they said to them, "Go and explore the land." And they came to the hill country of Ephraim, to the house of Micah, and lodged there.
JUDG|18|3|When they were by the house of Micah, they recognized the voice of the young Levite. And they turned aside and said to him, "Who brought you here? What are you doing in this place? What is your business here?"
JUDG|18|4|And he said to them, "This is how Micah dealt with me: he has hired me, and I have become his priest."
JUDG|18|5|And they said to him, "Inquire of God, please, that we may know whether the journey on which we are setting out will succeed."
JUDG|18|6|And the priest said to them, "Go in peace. The journey on which you go is under the eye of the LORD."
JUDG|18|7|Then the five men departed and came to Laish and saw the people who were there, how they lived in security, after the manner of the Sidonians, quiet and unsuspecting, lacking nothing that is in the earth and possessing wealth, and how they were far from the Sidonians and had no dealings with anyone.
JUDG|18|8|And when they came to their brothers at Zorah and Eshtaol, their brothers said to them, "What do you report?"
JUDG|18|9|They said, "Arise, and let us go up against them, for we have seen the land, and behold, it is very good. And will you do nothing? Do not be slow to go, to enter in and possess the land.
JUDG|18|10|As soon as you go, you will come to an unsuspecting people. The land is spacious, for God has given it into your hands, a place where there is no lack of anything that is in the earth."
JUDG|18|11|So 600 men of the tribe of Dan, armed with weapons of war, set out from Zorah and Eshtaol,
JUDG|18|12|and went up and encamped at Kiriath-jearim in Judah. On this account that place is called Mahaneh-dan to this day; behold, it is west of Kiriath-jearim.
JUDG|18|13|And they passed on from there to the hill country of Ephraim, and came to the house of Micah.
JUDG|18|14|Then the five men who had gone to scout out the country of Laish said to their brothers, "Do you know that in these houses there are an ephod, household gods, a carved image, and a metal image? Now therefore consider what you will do."
JUDG|18|15|And they turned aside there and came to the house of the young Levite, at the home of Micah, and asked him about his welfare.
JUDG|18|16|Now the 600 men of the Danites, armed with their weapons of war, stood by the entrance of the gate.
JUDG|18|17|And the five men who had gone to scout out the land went up and entered and took the carved image, the ephod, the household gods, and the metal image, while the priest stood by the entrance of the gate with the 600 men armed with weapons of war.
JUDG|18|18|And when these went into Micah's house and took the carved image, the ephod, the household gods, and the metal image, the priest said to them, "What are you doing?"
JUDG|18|19|And they said to him, "Keep quiet; put your hand on your mouth and come with us and be to us a father and a priest. Is it better for you to be priest to the house of one man, or to be priest to a tribe and clan in Israel?"
JUDG|18|20|And the priest's heart was glad. He took the ephod and the household gods and the carved image and went along with the people.
JUDG|18|21|So they turned and departed, putting the little ones and the livestock and the goods in front of them.
JUDG|18|22|When they had gone a distance from the home of Micah, the men who were in the houses near Micah's house were called out, and they overtook the people of Dan.
JUDG|18|23|And they shouted to the people of Dan, who turned around and said to Micah, "What is the matter with you, that you come with such a company?"
JUDG|18|24|And he said, "You take my gods that I made and the priest, and go away, and what have I left? How then do you ask me, 'What is the matter with you?'"
JUDG|18|25|And the people of Dan said to him, "Do not let your voice be heard among us, lest angry fellows fall upon you, and you lose your life with the lives of your household."
JUDG|18|26|Then the people of Dan went their way. And when Micah saw that they were too strong for him, he turned and went back to his home.
JUDG|18|27|But the people of Dan took what Micah had made, and the priest who belonged to him, and they came to Laish, to a people quiet and unsuspecting, and struck them with the edge of the sword and burned the city with fire.
JUDG|18|28|And there was no deliverer because it was far from Sidon, and they had no dealings with anyone. It was in the valley that belongs to Beth-rehob. Then they rebuilt the city and lived in it.
JUDG|18|29|And they named the city Dan, after the name of Dan their ancestor, who was born to Israel; but the name of the city was Laish at the first.
JUDG|18|30|And the people of Dan set up the carved image for themselves, and Jonathan the son of Gershom, son of Moses, and his sons were priests to the tribe of the Danites until the day of the captivity of the land.
JUDG|18|31|So they set up Micah's carved image that he made, as long as the house of God was at Shiloh.
JUDG|19|1|In those days, when there was no king in Israel, a certain Levite was sojourning in the remote parts of the hill country of Ephraim, who took to himself a concubine from Bethlehem in Judah.
JUDG|19|2|And his concubine was unfaithful to him, and she went away from him to her father's house at Bethlehem in Judah, and was there some four months.
JUDG|19|3|Then her husband arose and went after her, to speak kindly to her and bring her back. He had with him his servant and a couple of donkeys. And she brought him into her father's house. And when the girl's father saw him, he came with joy to meet him.
JUDG|19|4|And his father-in-law, the girl's father, made him stay, and he remained with him three days. So they ate and drank and spent the night there.
JUDG|19|5|And on the fourth day they arose early in the morning, and he prepared to go, but the girl's father said to his son-in-law, "Strengthen your heart with a morsel of bread, and after that you may go."
JUDG|19|6|So the two of them sat and ate and drank together. And the girl's father said to the man, "Be pleased to spend the night, and let your heart be merry."
JUDG|19|7|And when the man rose up to go, his father-in-law pressed him, till he spent the night there again.
JUDG|19|8|And on the fifth day he arose early in the morning to depart. And the girl's father said, "Strengthen your heart and wait until the day declines." So they ate, both of them.
JUDG|19|9|And when the man and his concubine and his servant rose up to depart, his father-in-law, the girl's father, said to him, "Behold, now the day has waned toward evening. Please, spend the night. Behold, the day draws to its close. Lodge here and let your heart be merry, and tomorrow you shall arise early in the morning for your journey, and go home."
JUDG|19|10|But the man would not spend the night. He rose up and departed and arrived opposite Jebus (that is, Jerusalem). He had with him a couple of saddled donkeys, and his concubine was with him.
JUDG|19|11|When they were near Jebus, the day was nearly over, and the servant said to his master, "Come now, let us turn aside to this city of the Jebusites and spend the night in it."
JUDG|19|12|And his master said to him, "We will not turn aside into the city of foreigners, who do not belong to the people of Israel, but we will pass on to Gibeah."
JUDG|19|13|And he said to his young man, "Come and let us draw near to one of these places and spend the night at Gibeah or at Ramah."
JUDG|19|14|So they passed on and went their way. And the sun went down on them near Gibeah, which belongs to Benjamin,
JUDG|19|15|and they turned aside there, to go in and spend the night at Gibeah. And he went in and sat down in the open square of the city, for no one took them into his house to spend the night.
JUDG|19|16|And behold, an old man was coming from his work in the field at evening. The man was from the hill country of Ephraim, and he was sojourning in Gibeah. The men of the place were Benjaminites.
JUDG|19|17|And he lifted up his eyes and saw the traveler in the open square of the city. And the old man said, "Where are you going? and where do you come from?"
JUDG|19|18|And he said to him, "We are passing from Bethlehem in Judah to the remote parts of the hill country of Ephraim, from which I come. I went to Bethlehem in Judah, and I am going to the house of the Lord, but no one has taken me into his house.
JUDG|19|19|We have straw and feed for our donkeys, with bread and wine for me and your female servant and the young man with your servants. There is no lack of anything."
JUDG|19|20|And the old man said, "Peace be to you; I will care for all your wants. Only, do not spend the night in the square."
JUDG|19|21|So he brought him into his house and gave the donkeys feed. And they washed their feet, and ate and drank.
JUDG|19|22|As they were making their hearts merry, behold, the men of the city, worthless fellows, surrounded the house, beating on the door. And they said to the old man, the master of the house, "Bring out the man who came into your house, that we may know him."
JUDG|19|23|And the man, the master of the house, went out to them and said to them, "No, my brothers, do not act so wickedly; since this man has come into my house, do not do this vile thing.
JUDG|19|24|Behold, here are my virgin daughter and his concubine. Let me bring them out now. Violate them and do with them what seems good to you, but against this man do not do this outrageous thing."
JUDG|19|25|But the men would not listen to him. So the man seized his concubine and made her go out to them. And they knew her and abused her all night until the morning. And as the dawn began to break, they let her go.
JUDG|19|26|And as morning appeared, the woman came and fell down at the door of the man's house where her master was, until it was light.
JUDG|19|27|And her master rose up in the morning, and when he opened the doors of the house and went out to go on his way, behold, there was his concubine lying at the door of the house, with her hands on the threshold.
JUDG|19|28|He said to her, "Get up, let us be going." But there was no answer. Then he put her on the donkey, and the man rose up and went away to his home.
JUDG|19|29|And when he entered his house, he took a knife, and taking hold of his concubine he divided her, limb by limb, into twelve pieces, and sent her throughout all the territory of Israel.
JUDG|19|30|And all who saw it said, "Such a thing has never happened or been seen from the day that the people of Israel came up out of the land of Egypt until this day; consider it, take counsel, and speak."
JUDG|20|1|Then all the people of Israel came out, from Dan to Beersheba, including the land of Gilead, and the congregation assembled as one man to the LORD at Mizpah.
JUDG|20|2|And the chiefs of all the people, of all the tribes of Israel, presented themselves in the assembly of the people of God, 400,000 men on foot that drew the sword.
JUDG|20|3|(Now the people of Benjamin heard that the people of Israel had gone up to Mizpah.) And the people of Israel said, "Tell us, how did this evil happen?"
JUDG|20|4|And the Levite, the husband of the woman who was murdered, answered and said, "I came to Gibeah that belongs to Benjamin, I and my concubine, to spend the night.
JUDG|20|5|And the leaders of Gibeah rose against me and surrounded the house against me by night. They meant to kill me, and they violated my concubine, and she is dead.
JUDG|20|6|So I took hold of my concubine and cut her in pieces and sent her throughout all the country of the inheritance of Israel, for they have committed abomination and outrage in Israel.
JUDG|20|7|Behold, you people of Israel, all of you, give your advice and counsel here."
JUDG|20|8|And all the people arose as one man, saying, "None of us will go to his tent, and none of us will return to his house.
JUDG|20|9|But now this is what we will do to Gibeah: we will go up against it by lot,
JUDG|20|10|and we will take ten men of a hundred throughout all the tribes of Israel, and a hundred of a thousand, and a thousand of ten thousand, to bring provisions for the people, that when they come they may repay Gibeah of Benjamin, for all the outrage that they have committed in Israel."
JUDG|20|11|So all the men of Israel gathered against the city, united as one man.
JUDG|20|12|And the tribes of Israel sent men through all the tribe of Benjamin, saying, "What evil is this that has taken place among you?
JUDG|20|13|Now therefore give up the men, the worthless fellows in Gibeah, that we may put them to death and purge evil from Israel." But the Benjaminites would not listen to the voice of their brothers, the people of Israel.
JUDG|20|14|Then the people of Benjamin came together out of the cities to Gibeah to go out to battle against the people of Israel.
JUDG|20|15|And the people of Benjamin mustered out of their cities on that day 26,000 men who drew the sword, besides the inhabitants of Gibeah, who mustered 700 chosen men.
JUDG|20|16|Among all these were 700 chosen men who were left-handed; every one could sling a stone at a hair and not miss.
JUDG|20|17|And the men of Israel, apart from Benjamin, mustered 400,000 men who drew the sword; all these were men of war.
JUDG|20|18|The people of Israel arose and went up to Bethel and inquired of God, "Who shall go up first for us to fight against the people of Benjamin?" And the LORD said, "Judah shall go up first."
JUDG|20|19|Then the people of Israel rose in the morning and encamped against Gibeah.
JUDG|20|20|And the men of Israel went out to fight against Benjamin, and the men of Israel drew up the battle line against them at Gibeah.
JUDG|20|21|The people of Benjamin came out of Gibeah and destroyed on that day 22,000 men of the Israelites.
JUDG|20|22|But the people, the men of Israel, took courage, and again formed the battle line in the same place where they had formed it on the first day.
JUDG|20|23|And the people of Israel went up and wept before the LORD until the evening. And they inquired of the LORD, "Shall we again draw near to fight against our brothers, the people of Benjamin?" And the LORD said, "Go up against them."
JUDG|20|24|So the people of Israel came near against the people of Benjamin the second day.
JUDG|20|25|And Benjamin went against them out of Gibeah the second day, and destroyed 18,000 men of the people of Israel. All these were men who drew the sword.
JUDG|20|26|Then all the people of Israel, the whole army, went up and came to Bethel and wept. They sat there before the LORD and fasted that day until evening, and offered burnt offerings and peace offerings before the LORD.
JUDG|20|27|And the people of Israel inquired of the LORD (for the ark of the covenant of God was there in those days,
JUDG|20|28|and Phinehas the son of Eleazar, son of Aaron, ministered before it in those days), saying, "Shall we go out once more to battle against our brothers, the people of Benjamin, or shall we cease?" And the LORD said, "Go up, for tomorrow I will give them into your hand."
JUDG|20|29|So Israel set men in ambush around Gibeah.
JUDG|20|30|And the people of Israel went up against the people of Benjamin on the third day and set themselves in array against Gibeah, as at other times.
JUDG|20|31|And the people of Benjamin went out against the people and were drawn away from the city. And as at other times they began to strike and kill some of the people in the highways, one of which goes up to Bethel and the other to Gibeah, and in the open country, about thirty men of Israel.
JUDG|20|32|And the people of Benjamin said, "They are routed before us, as at the first." But the people of Israel said, "Let us flee and draw them away from the city to the highways."
JUDG|20|33|And all the men of Israel rose up out of their place and set themselves in array at Baal-tamar, and the men of Israel who were in ambush rushed out of their place from Maareh-geba.
JUDG|20|34|And there came against Gibeah 10,000 chosen men out of all Israel, and the battle was hard, but the Benjaminites did not know that disaster was close upon them.
JUDG|20|35|And the LORD defeated Benjamin before Israel, and the people of Israel destroyed 25,100 men of Benjamin that day. All these were men who drew the sword.
JUDG|20|36|So the people of Benjamin saw that they were defeated. The men of Israel gave ground to Benjamin, because they trusted the men in ambush whom they had set against Gibeah.
JUDG|20|37|Then the men in ambush hurried and rushed against Gibeah; the men in ambush moved out and struck all the city with the edge of the sword.
JUDG|20|38|Now the appointed signal between the men of Israel and the men in the main ambush was that when they made a great cloud of smoke rise up out of the city
JUDG|20|39|the men of Israel should turn in battle. Now Benjamin had begun to strike and kill about thirty men of Israel. They said, "Surely they are defeated before us, as in the first battle."
JUDG|20|40|But when the signal began to rise out of the city in a column of smoke, the Benjaminites looked behind them, and behold, the whole of the city went up in smoke to heaven.
JUDG|20|41|Then the men of Israel turned, and the men of Benjamin were dismayed, for they saw that disaster was close upon them.
JUDG|20|42|Therefore they turned their backs before the men of Israel in the direction of the wilderness, but the battle overtook them. And those who came out of the cities were destroying them in their midst.
JUDG|20|43|Surrounding the Benjaminites, they pursued them and trod them down from Nohah as far as opposite Gibeah on the east.
JUDG|20|44|Eighteen thousand men of Benjamin fell, all of them men of valor.
JUDG|20|45|And they turned and fled toward the wilderness to the rock of Rimmon. Five thousand men of them were cut down in the highways. And they were pursued hard to Gidom, and 2,000 men of them were struck down.
JUDG|20|46|So all who fell that day of Benjamin were 25,000 men who drew the sword, all of them men of valor.
JUDG|20|47|But 600 men turned and fled toward the wilderness to the rock of Rimmon and remained at the rock of Rimmon four months.
JUDG|20|48|And the men of Israel turned back against the people of Benjamin and struck them with the edge of the sword, the city, men and beasts and all that they found. And all the towns that they found they set on fire.
JUDG|21|1|Now the men of Israel had sworn at Mizpah, "No one of us shall give his daughter in marriage to Benjamin."
JUDG|21|2|And the people came to Bethel and sat there till evening before God, and they lifted up their voices and wept bitterly.
JUDG|21|3|And they said, "O LORD, the God of Israel, why has this happened in Israel, that today there should be one tribe lacking in Israel?"
JUDG|21|4|And the next day the people rose early and built there an altar and offered burnt offerings and peace offerings.
JUDG|21|5|And the people of Israel said, "Which of all the tribes of Israel did not come up in the assembly to the LORD?" For they had taken a great oath concerning him who did not come up to the LORD to Mizpah, saying, "He shall surely be put to death."
JUDG|21|6|And the people of Israel had compassion for Benjamin their brother and said, "One tribe is cut off from Israel this day.
JUDG|21|7|What shall we do for wives for those who are left, since we have sworn by the LORD that we will not give them any of our daughters for wives?"
JUDG|21|8|And they said, "What one is there of the tribes of Israel that did not come up to the LORD to Mizpah?" And behold, no one had come to the camp from Jabesh-gilead, to the assembly.
JUDG|21|9|For when the people were mustered, behold, not one of the inhabitants of Jabesh-gilead was there.
JUDG|21|10|So the congregation sent 12,000 of their bravest men there and commanded them, "Go and strike the inhabitants of Jabesh-gilead with the edge of the sword; also the women and the little ones.
JUDG|21|11|This is what you shall do: every male and every woman that has lain with a male you shall devote to destruction."
JUDG|21|12|And they found among the inhabitants of Jabesh-gilead 400 young virgins who had not known a man by lying with him, and they brought them to the camp at Shiloh, which is in the land of Canaan.
JUDG|21|13|Then the whole congregation sent word to the people of Benjamin who were at the rock of Rimmon and proclaimed peace to them.
JUDG|21|14|And Benjamin returned at that time. And they gave them the women whom they had saved alive of the women of Jabesh-gilead, but they were not enough for them.
JUDG|21|15|And the people had compassion on Benjamin because the LORD had made a breach in the tribes of Israel.
JUDG|21|16|Then the elders of the congregation said, "What shall we do for wives for those who are left, since the women are destroyed out of Benjamin?"
JUDG|21|17|And they said, "There must be an inheritance for the survivors of Benjamin, that a tribe not be blotted out from Israel.
JUDG|21|18|Yet we cannot give them wives from our daughters." For the people of Israel had sworn, "Cursed be he who gives a wife to Benjamin."
JUDG|21|19|So they said, "Behold, there is the yearly feast of the LORD at Shiloh, which is north of Bethel, on the east of the highway that goes up from Bethel to Shechem, and south of Lebonah."
JUDG|21|20|And they commanded the people of Benjamin, saying, "Go and lie in ambush in the vineyards
JUDG|21|21|and watch. If the daughters of Shiloh come out to dance in the dances, then come out of the vineyards and snatch each man his wife from the daughters of Shiloh, and go to the land of Benjamin.
JUDG|21|22|And when their fathers or their brothers come to complain to us, we will say to them, 'Grant them graciously to us, because we did not take for each man of them his wife in battle, neither did you give them to them, else you would now be guilty.'"
JUDG|21|23|And the people of Benjamin did so and took their wives, according to their number, from the dancers whom they carried off. Then they went and returned to their inheritance and rebuilt the towns and lived in them.
JUDG|21|24|And the people of Israel departed from there at that time, every man to his tribe and family, and they went out from there every man to his inheritance.
JUDG|21|25|In those days there was no king in Israel. Everyone did what was right in his own eyes.
