AMOS|1|1|The words of Amos, who was among the shepherds of Tekoa, which he saw concerning Israel in the days of Uzziah king of Judah and in the days of Jeroboam the son of Joash, king of Israel, two years before the earthquake.
AMOS|1|2|And he said: "The LORD roars from Zion and utters his voice from Jerusalem; the pastures of the shepherds mourn, and the top of Carmel withers."
AMOS|1|3|Thus says the LORD: "For three transgressions of Damascus, and for four, I will not revoke the punishment, because they have threshed Gilead with threshing sledges of iron.
AMOS|1|4|So I will send a fire upon the house of Hazael, and it shall devour the strongholds of Ben-hadad.
AMOS|1|5|I will break the gate-bar of Damascus, and cut off the inhabitants from the Valley of Aven, and him who holds the scepter from Beth-eden; and the people of Syria shall go into exile to Kir," says the LORD.
AMOS|1|6|Thus says the LORD: "For three transgressions of Gaza, and for four, I will not revoke the punishment, because they carried into exile a whole people to deliver them up to Edom.
AMOS|1|7|So I will send a fire upon the wall of Gaza, and it shall devour her strongholds.
AMOS|1|8|I will cut off the inhabitants from Ashdod, and him who holds the scepter from Ashkelon; I will turn my hand against Ekron, and the remnant of the Philistines shall perish," says the Lord GOD.
AMOS|1|9|Thus says the LORD: "For three transgressions of Tyre, and for four, I will not revoke the punishment, because they delivered up a whole people to Edom, and did not remember the covenant of brotherhood.
AMOS|1|10|So I will send a fire upon the wall of Tyre, and it shall devour her strongholds."
AMOS|1|11|Thus says the LORD: "For three transgressions of Edom, and for four, I will not revoke the punishment, because he pursued his brother with the sword and cast off all pity, and his anger tore perpetually, and he kept his wrath forever.
AMOS|1|12|So I will send a fire upon Teman, and it shall devour the strongholds of Bozrah."
AMOS|1|13|Thus says the LORD: "For three transgressions of the Ammonites, and for four, I will not revoke the punishment, because they have ripped open pregnant women in Gilead, that they might enlarge their border.
AMOS|1|14|So I will kindle a fire in the wall of Rabbah, and it shall devour her strongholds, with shouting on the day of battle, with a tempest in the day of the whirlwind;
AMOS|1|15|and their king shall go into exile, he and his princes together," says the LORD.
AMOS|2|1|Thus says the LORD: "For three transgressions of Moab, and for four, I will not revoke the punishment, because he burned to lime the bones of the king of Edom.
AMOS|2|2|So I will send a fire upon Moab, and it shall devour the strongholds of Kerioth, and Moab shall die amid uproar, amid shouting and the sound of the trumpet;
AMOS|2|3|I will cut off the ruler from its midst, and will kill all its princes with him," says the LORD.
AMOS|2|4|Thus says the LORD: "For three transgressions of Judah, and for four, I will not revoke the punishment, because they have rejected the law of the LORD, and have not kept his statutes, but their lies have led them astray, those after which their fathers walked.
AMOS|2|5|So I will send a fire upon Judah, and it shall devour the strongholds of Jerusalem."
AMOS|2|6|Thus says the LORD: "For three transgressions of Israel, and for four, I will not revoke the punishment, because they sell the righteous for silver, and the needy for a pair of sandals-
AMOS|2|7|those who trample the head of the poor into the dust of the earth and turn aside the way of the afflicted; a man and his father go in to the same girl, so that my holy name is profaned;
AMOS|2|8|they lay themselves down beside every altar on garments taken in pledge, and in the house of their God they drink the wine of those who have been fined.
AMOS|2|9|"Yet it was I who destroyed the Amorite before them, whose height was like the height of the cedars and who was as strong as the oaks; I destroyed his fruit above and his roots beneath.
AMOS|2|10|Also it was I who brought you up out of the land of Egypt and led you forty years in the wilderness, to possess the land of the Amorite.
AMOS|2|11|And I raised up some of your sons for prophets, and some of your young men for Nazirites. Is it not indeed so, O people of Israel?" declares the LORD.
AMOS|2|12|"But you made the Nazirites drink wine, and commanded the prophets, saying, 'You shall not prophesy.'
AMOS|2|13|"Behold, I will press you down in your place, as a cart full of sheaves presses down.
AMOS|2|14|Flight shall perish from the swift, and the strong shall not retain his strength, nor shall the mighty save his life;
AMOS|2|15|he who handles the bow shall not stand, and he who is swift of foot shall not save himself, nor shall he who rides the horse save his life;
AMOS|2|16|and he who is stout of heart among the mighty shall flee away naked in that day," declares the LORD.
AMOS|3|1|Hear this word that the LORD has spoken against you, O people of Israel, against the whole family that I brought up out of the land of Egypt:
AMOS|3|2|"You only have I known of all the families of the earth; therefore I will punish you for all your iniquities.
AMOS|3|3|"Do two walk together, unless they have agreed to meet?
AMOS|3|4|Does a lion roar in the forest, when he has no prey? Does a young lion cry out from his den, if he has taken nothing?
AMOS|3|5|Does a bird fall in a snare on the earth, when there is no trap for it? Does a snare spring up from the ground, when it has taken nothing?
AMOS|3|6|Is a trumpet blown in a city, and the people are not afraid? Does disaster come to a city, unless the LORD has done it?
AMOS|3|7|"For the Lord GOD does nothing without revealing his secret to his servants the prophets.
AMOS|3|8|The lion has roared; who will not fear? The Lord GOD has spoken; who can but prophesy?"
AMOS|3|9|Proclaim to the strongholds in Ashdod and to the strongholds in the land of Egypt, and say, "Assemble yourselves on the mountains of Samaria, and see the great tumults within her, and the oppressed in her midst."
AMOS|3|10|"They do not know how to do right," declares the LORD, "those who store up violence and robbery in their strongholds."
AMOS|3|11|Therefore thus says the Lord GOD: "An adversary shall surround the land and bring down your defenses from you, and your strongholds shall be plundered."
AMOS|3|12|Thus says the LORD: "As the shepherd rescues from the mouth of the lion two legs, or a piece of an ear, so shall the people of Israel who dwell in Samaria be rescued, with the corner of a couch and part of a bed.
AMOS|3|13|"Hear, and testify against the house of Jacob," declares the Lord GOD, the God of hosts,
AMOS|3|14|"that on the day I punish Israel for his transgressions, I will punish the altars of Bethel, and the horns of the altar shall be cut off and fall to the ground.
AMOS|3|15|I will strike the winter house along with the summer house, and the houses of ivory shall perish, and the great houses shall come to an end," declares the LORD.
AMOS|4|1|"Hear this word, you cows of Bashan, who are on the mountain of Samaria, who oppress the poor, who crush the needy, who say to your husbands, 'Bring, that we may drink!'
AMOS|4|2|The Lord GOD has sworn by his holiness that, behold, the days are coming upon you, when they shall take you away with hooks, even the last of you with fishhooks.
AMOS|4|3|And you shall go out through the breaches, each one straight ahead; and you shall be cast out into Harmon," declares the LORD.
AMOS|4|4|"Come to Bethel, and transgress; to Gilgal, and multiply transgression; bring your sacrifices every morning, your tithes every three days;
AMOS|4|5|offer a sacrifice of thanksgiving of that which is leavened, and proclaim freewill offerings, publish them; for so you love to do, O people of Israel!" declares the Lord GOD.
AMOS|4|6|"I gave you cleanness of teeth in all your cities, and lack of bread in all your places, yet you did not return to me," declares the LORD.
AMOS|4|7|"I also withheld the rain from you when there were yet three months to the harvest; I would send rain on one city, and send no rain on another city; one field would have rain, and the field on which it did not rain would wither;
AMOS|4|8|so two or three cities would wander to another city to drink water, and would not be satisfied; yet you did not return to me," declares the LORD.
AMOS|4|9|"I struck you with blight and mildew; your many gardens and your vineyards, your fig trees and your olive trees the locust devoured; yet you did not return to me," declares the LORD.
AMOS|4|10|"I sent among you a pestilence after the manner of Egypt; I killed your young men with the sword, and carried away your horses, and I made the stench of your camp go up into your nostrils; yet you did not return to me," declares the LORD.
AMOS|4|11|"I overthrew some of you, as when God overthrew Sodom and Gomorrah, and you were as a brand plucked out of the burning; yet you did not return to me," declares the LORD.
AMOS|4|12|"Therefore thus I will do to you, O Israel; because I will do this to you, prepare to meet your God, O Israel!"
AMOS|4|13|For behold, he who forms the mountains and creates the wind, and declares to man what is his thought, who makes the morning darkness, and treads on the heights of the earth- the LORD, the God of hosts, is his name!
AMOS|5|1|Hear this word that I take up over you in lamentation, O house of Israel:
AMOS|5|2|"Fallen, no more to rise, is the virgin Israel; forsaken on her land, with none to raise her up."
AMOS|5|3|For thus says the Lord GOD: "The city that went out a thousand shall have a hundred left, and that which went out a hundred shall have ten left to the house of Israel."
AMOS|5|4|For thus says the LORD to the house of Israel: "Seek me and live;
AMOS|5|5|but do not seek Bethel, and do not enter into Gilgal or cross over to Beersheba; for Gilgal shall surely go into exile, and Bethel shall come to nothing."
AMOS|5|6|Seek the LORD and live, lest he break out like fire in the house of Joseph, and it devour, with none to quench it for Bethel,
AMOS|5|7|O you who turn justice to wormwood and cast down righteousness to the earth!
AMOS|5|8|He who made the Pleiades and Orion, and turns deep darkness into the morning and darkens the day into night, who calls for the waters of the sea and pours them out on the surface of the earth, the LORD is his name;
AMOS|5|9|who makes destruction flash forth against the strong, so that destruction comes upon the fortress.
AMOS|5|10|They hate him who reproves in the gate, and they abhor him who speaks the truth.
AMOS|5|11|Therefore because you trample on the poor and you exact taxes of grain from him, you have built houses of hewn stone, but you shall not dwell in them; you have planted pleasant vineyards, but you shall not drink their wine.
AMOS|5|12|For I know how many are your transgressions and how great are your sins- you who afflict the righteous, who take a bribe, and turn aside the needy in the gate.
AMOS|5|13|Therefore he who is prudent will keep silent in such a time, for it is an evil time.
AMOS|5|14|Seek good, and not evil, that you may live; and so the LORD, the God of hosts, will be with you, as you have said.
AMOS|5|15|Hate evil, and love good, and establish justice in the gate; it may be that the LORD, the God of hosts, will be gracious to the remnant of Joseph.
AMOS|5|16|Therefore thus says the LORD, the God of hosts, the Lord: "In all the squares there shall be wailing, and in all the streets they shall say, 'Alas! Alas!' They shall call the farmers to mourning and to wailing those who are skilled in lamentation,
AMOS|5|17|and in all vineyards there shall be wailing, for I will pass through your midst," says the LORD.
AMOS|5|18|Woe to you who desire the day of the LORD! Why would you have the day of the LORD? It is darkness, and not light,
AMOS|5|19|as if a man fled from a lion, and a bear met him, or went into the house and leaned his hand against the wall, and a serpent bit him.
AMOS|5|20|Is not the day of the LORD darkness, and not light, and gloom with no brightness in it?
AMOS|5|21|"I hate, I despise your feasts, and I take no delight in your solemn assemblies.
AMOS|5|22|Even though you offer me your burnt offerings and grain offerings, I will not accept them; and the peace offerings of your fattened animals, I will not look upon them.
AMOS|5|23|Take away from me the noise of your songs; to the melody of your harps I will not listen.
AMOS|5|24|But let justice roll down like waters, and righteousness like an ever-flowing stream.
AMOS|5|25|"Did you bring to me sacrifices and offerings during the forty years in the wilderness, O house of Israel?
AMOS|5|26|You shall take up Sikkuth your king, and Kiyyun your star-god- your images that you made for yourselves,
AMOS|5|27|and I will send you into exile beyond Damascus," says the LORD, whose name is the God of hosts.
AMOS|6|1|"Woe to those who are at ease in Zion, and to those who feel secure on the mountain of Samaria, the notable men of the first of the nations, to whom the house of Israel comes!
AMOS|6|2|Pass over to Calneh, and see, and from there go to Hamath the great; then go down to Gath of the Philistines. Are you better than these kingdoms? Or is their territory greater than your territory,
AMOS|6|3|O you who put far away the day of disaster and bring near the seat of violence?
AMOS|6|4|"Woe to those who lie on beds of ivory and stretch themselves out on their couches, and eat lambs from the flock and calves from the midst of the stall,
AMOS|6|5|who sing idle songs to the sound of the harp and like David invent for themselves instruments of music,
AMOS|6|6|who drink wine in bowls and anoint themselves with the finest oils, but are not grieved over the ruin of Joseph!
AMOS|6|7|Therefore they shall now be the first of those who go into exile, and the revelry of those who stretch themselves out shall pass away."
AMOS|6|8|The Lord GOD has sworn by himself, declares the LORD, the God of hosts: "I abhor the pride of Jacob and hate his strongholds, and I will deliver up the city and all that is in it."
AMOS|6|9|And if ten men remain in one house, they shall die.
AMOS|6|10|And when one's relative, the one who anoints him for burial, shall take him up to bring the bones out of the house, and shall say to him who is in the innermost parts of the house, "Is there still anyone with you?" he shall say, "No"; and he shall say, "Silence! We must not mention the name of the LORD."
AMOS|6|11|For behold, the LORD commands, and the great house shall be struck down into fragments, and the little house into bits.
AMOS|6|12|Do horses run on rocks? Does one plow there with oxen? But you have turned justice into poison and the fruit of righteousness into wormwood-
AMOS|6|13|you who rejoice in Lo-debar, who say, "Have we not by our own strength captured Karnaim for ourselves?"
AMOS|6|14|"For behold, I will raise up against you a nation, O house of Israel," declares the LORD, the God of hosts; "and they shall oppress you from Lebo-hamath to the Brook of the Arabah."
AMOS|7|1|This is what the Lord GOD showed me: behold, he was forming locusts when the latter growth was just beginning to sprout, and behold, it was the latter growth after the king's mowings.
AMOS|7|2|When they had finished eating the grass of the land, I said, "O Lord GOD, please forgive! How can Jacob stand? He is so small!"
AMOS|7|3|The LORD relented concerning this; "It shall not be," said the LORD.
AMOS|7|4|This is what the Lord GOD showed me: behold, the Lord GOD was calling for a judgment by fire, and it devoured the great deep and was eating up the land.
AMOS|7|5|Then I said, "O Lord GOD, please cease! How can Jacob stand? He is so small!"
AMOS|7|6|The LORD relented concerning this; "This also shall not be," said the Lord GOD.
AMOS|7|7|This is what he showed me: behold, the Lord was standing beside a wall built with a plumb line, with a plumb line in his hand.
AMOS|7|8|And the LORD said to me, "Amos, what do you see?" And I said, "A plumb line." Then the Lord said, "Behold, I am setting a plumb line in the midst of my people Israel; I will never again pass by them;
AMOS|7|9|the high places of Isaac shall be made desolate, and the sanctuaries of Israel shall be laid waste, and I will rise against the house of Jeroboam with the sword."
AMOS|7|10|Then Amaziah the priest of Bethel sent to Jeroboam king of Israel, saying, "Amos has conspired against you in the midst of the house of Israel. The land is not able to bear all his words.
AMOS|7|11|For thus Amos has said, "' Jeroboam shall die by the sword, and Israel must go into exile away from his land.'"
AMOS|7|12|And Amaziah said to Amos, "O seer, go, flee away to the land of Judah, and eat bread there, and prophesy there,
AMOS|7|13|but never again prophesy at Bethel, for it is the king's sanctuary, and it is a temple of the kingdom."
AMOS|7|14|Then Amos answered and said to Amaziah, "I was no prophet, nor a prophet's son, but I was a herdsman and a dresser of sycamore figs.
AMOS|7|15|But the LORD took me from following the flock, and the LORD said to me, 'Go, prophesy to my people Israel.'
AMOS|7|16|Now therefore hear the word of the LORD. "You say, 'Do not prophesy against Israel, and do not preach against the house of Isaac.'
AMOS|7|17|Therefore thus says the LORD: "' Your wife shall be a prostitute in the city, and your sons and your daughters shall fall by the sword, and your land shall be divided up with a measuring line; you yourself shall die in an unclean land, and Israel shall surely go into exile away from its land.'"
AMOS|8|1|This is what the Lord GOD showed me: behold, a basket of summer fruit.
AMOS|8|2|And he said, "Amos, what do you see?" And I said, "A basket of summer fruit." Then the LORD said to me, "The end has come upon my people Israel; I will never again pass by them.
AMOS|8|3|The songs of the temple shall become wailings in that day," declares the Lord GOD. "So many dead bodies!" "They are thrown everywhere!" "Silence!"
AMOS|8|4|Hear this, you who trample on the needy and bring the poor of the land to an end,
AMOS|8|5|saying, "When will the new moon be over, that we may sell grain? And the Sabbath, that we may offer wheat for sale, that we may make the ephah small and the shekel great and deal deceitfully with false balances,
AMOS|8|6|that we may buy the poor for silver and the needy for a pair of sandals and sell the chaff of the wheat?"
AMOS|8|7|The LORD has sworn by the pride of Jacob: "Surely I will never forget any of their deeds.
AMOS|8|8|Shall not the land tremble on this account, and everyone mourn who dwells in it, and all of it rise like the Nile, and be tossed about and sink again, like the Nile of Egypt?"
AMOS|8|9|"And on that day," declares the Lord GOD, "I will make the sun go down at noon and darken the earth in broad daylight.
AMOS|8|10|I will turn your feasts into mourning and all your songs into lamentation; I will bring sackcloth on every waist and baldness on every head; I will make it like the mourning for an only son and the end of it like a bitter day.
AMOS|8|11|"Behold, the days are coming," declares the Lord GOD, "when I will send a famine on the land- not a famine of bread, nor a thirst for water, but of hearing the words of the LORD.
AMOS|8|12|They shall wander from sea to sea, and from north to east; they shall run to and fro, to seek the word of the LORD, but they shall not find it.
AMOS|8|13|"In that day the lovely virgins and the young men shall faint for thirst.
AMOS|8|14|Those who swear by the Guilt of Samaria, and say, 'As your god lives, O Dan,' and, 'As the Way of Beersheba lives,' they shall fall, and never rise again."
AMOS|9|1|I saw the LORD standing beside the altar, and he said: "Strike the capitals until the thresholds shake, and shatter them on the heads of all the people; and those who are left of them I will kill with the sword; not one of them shall flee away; not one of them shall escape.
AMOS|9|2|"If they dig into Sheol, from there shall my hand take them; if they climb up to heaven, from there I will bring them down.
AMOS|9|3|If they hide themselves on the top of Carmel, from there I will search them out and take them; and if they hide from my sight at the bottom of the sea, there I will command the serpent, and it shall bite them.
AMOS|9|4|And if they go into captivity before their enemies, there I will command the sword, and it shall kill them; and I will fix my eyes upon them for evil and not for good."
AMOS|9|5|The Lord GOD of hosts, he who touches the earth and it melts, and all who dwell in it mourn, and all of it rises like the Nile, and sinks again, like the Nile of Egypt;
AMOS|9|6|who builds his upper chambers in the heavens and founds his vault upon the earth; who calls for the waters of the sea and pours them out upon the surface of the earth- the LORD is his name.
AMOS|9|7|"Are you not like the Cushites to me, O people of Israel?" declares the LORD. "Did I not bring up Israel from the land of Egypt, and the Philistines from Caphtor and the Syrians from Kir?
AMOS|9|8|Behold, the eyes of the Lord GOD are upon the sinful kingdom, and I will destroy it from the surface of the ground, except that I will not utterly destroy the house of Jacob," declares the LORD.
AMOS|9|9|"For behold, I will command, and shake the house of Israel among all the nations as one shakes with a sieve, but no pebble shall fall to the earth.
AMOS|9|10|All the sinners of my people shall die by the sword, who say, 'Disaster shall not overtake or meet us.'
AMOS|9|11|"In that day I will raise up the booth of David that is fallen and repair its breaches, and raise up its ruins and rebuild it as in the days of old,
AMOS|9|12|that they may possess the remnant of Edom and all the nations who are called by my name," declares the LORD who does this.
AMOS|9|13|"Behold, the days are coming," declares the LORD, "when the plowman shall overtake the reaper and the treader of grapes him who sows the seed; the mountains shall drip sweet wine, and all the hills shall flow with it.
AMOS|9|14|I will restore the fortunes of my people Israel, and they shall rebuild the ruined cities and inhabit them; they shall plant vineyards and drink their wine, and they shall make gardens and eat their fruit.
AMOS|9|15|I will plant them on their land, and they shall never again be uprooted out of the land that I have given them," says the LORD your God.
