1CHR|1|1|Adam, Seth, Enosh;
1CHR|1|2|Kenan, Mahalalel, Jared;
1CHR|1|3|Enoch, Methuselah, Lamech;
1CHR|1|4|Noah, Shem, Ham, and Japheth.
1CHR|1|5|The sons of Japheth: Gomer, Magog, Madai, Javan, Tubal, Meshech, and Tiras.
1CHR|1|6|The sons of Gomer: Ashkenaz, Riphath, and Togarmah.
1CHR|1|7|The sons of Javan: Elishah, Tarshish, Kittim, and Rodanim.
1CHR|1|8|The sons of Ham: Cush, Egypt, Put, and Canaan.
1CHR|1|9|The sons of Cush: Seba, Havilah, Sabta, Raama, and Sabteca. The sons of Raamah: Sheba and Dedan.
1CHR|1|10|Cush fathered Nimrod. He was the first on earth to be a mighty man.
1CHR|1|11|Egypt fathered Ludim, Anamim, Lehabim, Naphtuhim,
1CHR|1|12|Pathrusim, Casluhim (from whom the Philistines came), and Caphtorim.
1CHR|1|13|Canaan fathered Sidon his firstborn and Heth,
1CHR|1|14|and the Jebusites, the Amorites, the Girgashites,
1CHR|1|15|the Hivites, the Arkites, the Sinites,
1CHR|1|16|the Arvadites, the Zemarites, and the Hamathites.
1CHR|1|17|The sons of Shem: Elam, Asshur, Arpachshad, Lud, and Aram. And the sons of Aram: Uz, Hul, Gether, and Meshech.
1CHR|1|18|Arpachshad fathered Shelah, and Shelah fathered Eber.
1CHR|1|19|To Eber were born two sons: the name of the one was Peleg (for in his days the earth was divided), and his brother's name was Joktan.
1CHR|1|20|Joktan fathered Almodad, Sheleph, Hazarmaveth, Jerah,
1CHR|1|21|Hadoram, Uzal, Diklah,
1CHR|1|22|Obal, Abimael, Sheba,
1CHR|1|23|Ophir, Havilah, and Jobab; all these were the sons of Joktan.
1CHR|1|24|Shem, Arpachshad, Shelah;
1CHR|1|25|Eber, Peleg, Reu;
1CHR|1|26|Serug, Nahor, Terah;
1CHR|1|27|Abram, that is, Abraham.
1CHR|1|28|The sons of Abraham: Isaac and Ishmael.
1CHR|1|29|These are their genealogies: the firstborn of Ishmael, Nebaioth, and Kedar, Adbeel, Mibsam,
1CHR|1|30|Mishma, Dumah, Massa, Hadad, Tema,
1CHR|1|31|Jetur, Naphish, and Kedemah. These are the sons of Ishmael.
1CHR|1|32|The sons of Keturah, Abraham's concubine: she bore Zimran, Jokshan, Medan, Midian, Ishbak, and Shuah. The sons of Jokshan: Sheba and Dedan.
1CHR|1|33|The sons of Midian: Ephah, Epher, Hanoch, Abida, and Eldaah. All these were the descendants of Keturah.
1CHR|1|34|Abraham fathered Isaac. The sons of Isaac: Esau and Israel.
1CHR|1|35|The sons of Esau: Eliphaz, Reuel, Jeush, Jalam, and Korah.
1CHR|1|36|The sons of Eliphaz: Teman, Omar, Zepho, Gatam, Kenaz, and of Timna, Amalek.
1CHR|1|37|The sons of Reuel: Nahath, Zerah, Shammah, and Mizzah.
1CHR|1|38|The sons of Seir: Lotan, Shobal, Zibeon, Anah, Dishon, Ezer, and Dishan.
1CHR|1|39|The sons of Lotan: Hori and Hemam; and Lotan's sister was Timna.
1CHR|1|40|The sons of Shobal: Alvan, Manahath, Ebal, Shepho, and Onam. The sons of Zibeon: Aiah and Anah.
1CHR|1|41|The son of Anah: Dishon. The sons of Dishon: Hemdan, Eshban, Ithran, and Cheran.
1CHR|1|42|The sons of Ezer: Bilhan, Zaavan, and Akan. The sons of Dishan: Uz and Aran.
1CHR|1|43|These are the kings who reigned in the land of Edom before any king reigned over the people of Israel: Bela the son of Beor, the name of his city being Dinhabah.
1CHR|1|44|Bela died, and Jobab the son of Zerah of Bozrah reigned in his place.
1CHR|1|45|Jobab died, and Husham of the land of the Temanites reigned in his place.
1CHR|1|46|Husham died, and Hadad the son of Bedad, who defeated Midian in the country of Moab, reigned in his place, the name of his city being Avith.
1CHR|1|47|Hadad died, and Samlah of Masrekah reigned in his place.
1CHR|1|48|Samlah died, and Shaul of Rehoboth on the Euphrates reigned in his place.
1CHR|1|49|Shaul died, and Baal-hanan, the son of Achbor, reigned in his place.
1CHR|1|50|Baal-hanan died, and Hadad reigned in his place, the name of his city being Pai; and his wife's name was Mehetabel, the daughter of Matred, the daughter of Mezahab.
1CHR|1|51|And Hadad died. The chiefs of Edom were: chiefs Timna, Alvah, Jetheth,
1CHR|1|52|Oholibamah, Elah, Pinon,
1CHR|1|53|Kenaz, Teman, Mibzar,
1CHR|1|54|Magdiel, and Iram; these are the chiefs of Edom.
1CHR|2|1|These are the sons of Israel: Reuben, Simeon, Levi, Judah, Issachar, Zebulun,
1CHR|2|2|Dan, Joseph, Benjamin, Naphtali, Gad, and Asher.
1CHR|2|3|The sons of Judah: Er, Onan and Shelah; these three Bath-shua the Canaanite bore to him. Now Er, Judah's firstborn, was evil in the sight of the LORD, and he put him to death.
1CHR|2|4|His daughter-in-law Tamar also bore him Perez and Zerah. Judah had five sons in all.
1CHR|2|5|The sons of Perez: Hezron and Hamul.
1CHR|2|6|The sons of Zerah: Zimri, Ethan, Heman, Calcol, and Dara, five in all.
1CHR|2|7|The son of Carmi: Achan, the troubler of Israel, who broke faith in the matter of the devoted thing;
1CHR|2|8|and Ethan's son was Azariah.
1CHR|2|9|The sons of Hezron that were born to him: Jerahmeel, Ram, and Chelubai.
1CHR|2|10|Ram fathered Amminadab, and Amminadab fathered Nahshon, prince of the sons of Judah.
1CHR|2|11|Nahshon fathered Salmon, Salmon fathered Boaz,
1CHR|2|12|Boaz fathered Obed, Obed fathered Jesse.
1CHR|2|13|Jesse fathered Eliab his firstborn, Abinadab the second, Shimea the third,
1CHR|2|14|Nethanel the fourth, Raddai the fifth,
1CHR|2|15|Ozem the sixth, David the seventh.
1CHR|2|16|And their sisters were Zeruiah and Abigail. The sons of Zeruiah: Abishai, Joab, and Asahel, three.
1CHR|2|17|Abigail bore Amasa, and the father of Amasa was Jether the Ishmaelite.
1CHR|2|18|Caleb the son of Hezron fathered children by his wife Azubah, and by Jerioth; and these were her sons: Jesher, Shobab, and Ardon.
1CHR|2|19|When Azubah died, Caleb married Ephrath, who bore him Hur.
1CHR|2|20|Hur fathered Uri, and Uri fathered Bezalel.
1CHR|2|21|Afterward Hezron went in to the daughter of Machir the father of Gilead, whom he married when he was sixty years old, and she bore him Segub.
1CHR|2|22|And Segub fathered Jair, who had twenty-three cities in the land of Gilead.
1CHR|2|23|But Geshur and Aram took from them Havvoth-jair, Kenath, and its villages, sixty towns. All these were descendants of Machir, the father of Gilead.
1CHR|2|24|After the death of Hezron, Caleb went in to Ephrathah, the wife of Hezron his father, and she bore him Ashhur, the father of Tekoa.
1CHR|2|25|The sons of Jerahmeel, the firstborn of Hezron: Ram, his firstborn, Bunah, Oren, Ozem, and Ahijah.
1CHR|2|26|Jerahmeel also had another wife, whose name was Atarah; she was the mother of Onam.
1CHR|2|27|The sons of Ram, the firstborn of Jerahmeel: Maaz, Jamin, and Eker.
1CHR|2|28|The sons of Onam: Shammai and Jada. The sons of Shammai: Nadab and Abishur.
1CHR|2|29|The name of Abishur's wife was Abihail, and she bore him Ahban and Molid.
1CHR|2|30|The sons of Nadab: Seled and Appaim; and Seled died childless.
1CHR|2|31|The son of Appaim: Ishi. The son of Ishi: Sheshan. The son of Sheshan: Ahlai.
1CHR|2|32|The sons of Jada, Shammai's brother: Jether and Jonathan; and Jether died childless.
1CHR|2|33|The sons of Jonathan: Peleth and Zaza. These were the descendants of Jerahmeel.
1CHR|2|34|Now Sheshan had no sons, only daughters, but Sheshan had an Egyptian slave whose name was Jarha.
1CHR|2|35|So Sheshan gave his daughter in marriage to Jarha his slave, and she bore him Attai.
1CHR|2|36|Attai fathered Nathan, and Nathan fathered Zabad.
1CHR|2|37|Zabad fathered Ephlal, and Ephlal fathered Obed.
1CHR|2|38|Obed fathered Jehu, and Jehu fathered Azariah.
1CHR|2|39|Azariah fathered Helez, and Helez fathered Eleasah.
1CHR|2|40|Eleasah fathered Sismai, and Sismai fathered Shallum.
1CHR|2|41|Shallum fathered Jekamiah, and Jekamiah fathered Elishama.
1CHR|2|42|The sons of Caleb the brother of Jerahmeel: Mareshah his firstborn, who fathered Ziph. The son of Mareshah: Hebron.
1CHR|2|43|The sons of Hebron: Korah, Tappuah, Rekem and Shema.
1CHR|2|44|Shema fathered Raham, the father of Jorkeam; and Rekem fathered Shammai.
1CHR|2|45|The son of Shammai: Maon; and Maon fathered Beth-zur.
1CHR|2|46|Ephah also, Caleb's concubine, bore Haran, Moza, and Gazez; and Haran fathered Gazez.
1CHR|2|47|The sons of Jahdai: Regem, Jotham, Geshan, Pelet, Ephah, and Shaaph.
1CHR|2|48|Maacah, Caleb's concubine, bore Sheber and Tirhanah.
1CHR|2|49|She also bore Shaaph the father of Madmannah, Sheva the father of Machbenah and the father of Gibea; and the daughter of Caleb was Achsah.
1CHR|2|50|These were the descendants of Caleb. The sons of Hur the firstborn of Ephrathah: Shobal the father of Kiriath-jearim,
1CHR|2|51|Salma, the father of Bethlehem, and Hareph the father of Beth-gader.
1CHR|2|52|Shobal the father of Kiriath-jearim had other sons: Haroeh, half of the Menuhoth.
1CHR|2|53|And the clans of Kiriath-jearim: the Ithrites, the Puthites, the Shumathites, and the Mishraites; from these came the Zorathites and the Eshtaolites.
1CHR|2|54|The sons of Salma: Bethlehem, the Netophathites, Atroth-beth-joab and half of the Manahathites, the Zorites.
1CHR|2|55|The clans also of the scribes who lived at Jabez: the Tirathites, the Shimeathites and the Sucathites. These are the Kenites who came from Hammath, the father of the house of Rechab.
1CHR|3|1|These are the sons of David who were born to him in Hebron: the firstborn, Amnon, by Ahinoam the Jezreelite; the second, Daniel, by Abigail the Carmelite,
1CHR|3|2|the third, Absalom, whose mother was Maacah, the daughter of Talmai, king of Geshur; the fourth, Adonijah, whose mother was Haggith;
1CHR|3|3|the fifth, Shephatiah, by Abital; the sixth, Ithream, by his wife Eglah;
1CHR|3|4|six were born to him in Hebron, where he reigned for seven years and six months. And he reigned thirty-three years in Jerusalem.
1CHR|3|5|These were born to him in Jerusalem: Shimea, Shobab, Nathan and Solomon, four by Bath-shua, the daughter of Ammiel;
1CHR|3|6|then Ibhar, Elishama, Eliphelet,
1CHR|3|7|Nogah, Nepheg, Japhia,
1CHR|3|8|Elishama, Eliada, and Eliphelet, nine.
1CHR|3|9|All these were David's sons, besides the sons of the concubines, and Tamar was their sister.
1CHR|3|10|The son of Solomon was Rehoboam, Abijah his son, Asa his son, Jehoshaphat his son,
1CHR|3|11|Joram his son, Ahaziah his son, Joash his son,
1CHR|3|12|Amaziah his son, Azariah his son, Jotham his son,
1CHR|3|13|Ahaz his son, Hezekiah his son, Manasseh his son,
1CHR|3|14|Amon his son, Josiah his son.
1CHR|3|15|The sons of Josiah: Johanan the firstborn, the second Jehoiakim, the third Zedekiah, the fourth Shallum.
1CHR|3|16|The descendants of Jehoiakim: Jeconiah his son, Zedekiah his son;
1CHR|3|17|and the sons of Jeconiah, the captive: Shealtiel his son,
1CHR|3|18|Malchiram, Pedaiah, Shenazzar, Jekamiah, Hosh-ama and Nedabiah;
1CHR|3|19|and the sons of Pedaiah: Zerubbabel and Shimei; and the sons of Zerubbabel: Meshullam and Hananiah, and Shelomith was their sister;
1CHR|3|20|and Hashubah, Ohel, Berechiah, Hasadiah, and Jushab-hesed, five.
1CHR|3|21|The sons of Hananiah: Pelatiah and Jeshaiah, his son Rephaiah, his son Arnan, his son Obadiah, his son Shecaniah.
1CHR|3|22|The son of Shecaniah: Shemaiah. And the sons of Shemaiah: Hattush, Igal, Bariah, Neariah, and Shaphat, six.
1CHR|3|23|The sons of Neariah: Elioenai, Hizkiah, and Azrikam, three.
1CHR|3|24|The sons of Elioenai: Hodaviah, Eliashib, Pelaiah, Akkub, Johanan, Delaiah, and Anani, seven.
1CHR|4|1|The sons of Judah: Perez, Hezron, Carmi, Hur, and Shobal.
1CHR|4|2|Reaiah the son of Shobal fathered Jahath, and Jahath fathered Ahumai and Lahad. These were the clans of the Zorathites.
1CHR|4|3|These were the sons of Etam: Jezreel, Ishma, and Idbash; and the name of their sister was Haz-zelelponi,
1CHR|4|4|and Penuel fathered Gedor, and Ezer fathered Hushah. These were the sons of Hur, the firstborn of Ephrathah, the father of Bethlehem.
1CHR|4|5|Ashhur, the father of Tekoa, had two wives, Helah and Naarah;
1CHR|4|6|Naarah bore him Ahuzzam, Hepher, Temeni, and Haahashtari. These were the sons of Naarah.
1CHR|4|7|The sons of Helah: Zereth, Izhar, and Ethnan.
1CHR|4|8|Koz fathered Anub, Zobebah, and the clans of Aharhel, the son of Harum.
1CHR|4|9|Jabez was more honorable than his brothers; and his mother called his name Jabez, saying, "Because I bore him in pain."
1CHR|4|10|Jabez called upon the God of Israel, saying, "Oh that you would bless me and enlarge my border, and that your hand might be with me, and that you would keep me from harm so that it might not bring me pain!" And God granted what he asked.
1CHR|4|11|Chelub, the brother of Shuhah, fathered Mehir, who fathered Eshton.
1CHR|4|12|Eshton fathered Beth-rapha, Paseah, and Tehinnah, the father of Ir-nahash. These are the men of Recah.
1CHR|4|13|The sons of Kenaz: Othniel and Seraiah; and the sons of Othniel: Hathath and Meonothai.
1CHR|4|14|Meonothai fathered Ophrah; and Seraiah fathered Joab, the father of Ge-harashim, so-called because they were craftsmen.
1CHR|4|15|The sons of Caleb the son of Jephunneh: Iru, Elah, and Naam; and the son of Elah: Kenaz.
1CHR|4|16|The sons of Jehallelel: Ziph, Ziphah, Tiria, and Asarel.
1CHR|4|17|The sons of Ezrah: Jether, Mered, Epher, and Jalon. These are the sons of Bithiah, the daughter of Pharaoh, whom Mered married; and she conceived and bore Miriam, Shammai, and Ishbah, the father of Eshtemoa.
1CHR|4|18|And his Judahite wife bore Jered the father of Gedor, Heber the father of Soco, and Jekuthiel the father of Zanoah.
1CHR|4|19|The sons of the wife of Hodiah, the sister of Naham, were the fathers of Keilah the Garmite and Eshtemoa the Maacathite.
1CHR|4|20|The sons of Shimon: Amnon, Rinnah, Ben-hanan, and Tilon. The sons of Ishi: Zoheth and Ben-zoheth.
1CHR|4|21|The sons of Shelah the son of Judah: Er the father of Lecah, Laadah the father of Mareshah, and the clans of the house of linen workers at Beth-ashbea;
1CHR|4|22|and Jokim, and the men of Cozeba, and Joash, and Saraph, who ruled in Moab and returned to Lehem (now the records are ancient).
1CHR|4|23|These were the potters who were inhabitants of Netaim and Gederah. They lived there in the king's service.
1CHR|4|24|The sons of Simeon: Nemuel, Jamin, Jarib, Zerah, Shaul;
1CHR|4|25|Shallum was his son, Mibsam his son, Mishma his son.
1CHR|4|26|The sons of Mishma: Hammuel his son, Zaccur his son, Shimei his son.
1CHR|4|27|Shimei had sixteen sons and six daughters; but his brothers did not have many children, nor did all their clan multiply like the men of Judah.
1CHR|4|28|They lived in Beersheba, Moladah, Hazar-shual,
1CHR|4|29|Bilhah, Ezem, Tolad,
1CHR|4|30|Bethuel, Hormah, Ziklag,
1CHR|4|31|Beth-marcaboth, Hazar-su-sim, Beth-biri, and Shaaraim. These were their cities until David reigned.
1CHR|4|32|And their villages were Etam, Ain, Rimmon, Tochen, and Ashan, five cities,
1CHR|4|33|along with all their villages that were around these cities as far as Baal. These were their settlements, and they kept a genealogical record.
1CHR|4|34|Meshobab, Jamlech, Joshah the son of Amaziah,
1CHR|4|35|Joel, Jehu the son of Joshibiah, son of Seraiah, son of Asiel,
1CHR|4|36|Elioenai, Jaakobah, Jeshohaiah, Asaiah, Adiel, Jesimiel, Benaiah,
1CHR|4|37|Ziza the son of Shiphi, son of Allon, son of Jedaiah, son of Shimri, son of Shemaiah-
1CHR|4|38|these mentioned by name were princes in their clans, and their fathers' houses increased greatly.
1CHR|4|39|They journeyed to the entrance of Gedor, to the east side of the valley, to seek pasture for their flocks,
1CHR|4|40|where they found rich, good pasture, and the land was very broad, quiet, and peaceful, for the former inhabitants there belonged to Ham.
1CHR|4|41|These, registered by name, came in the days of Hezekiah, king of Judah, and destroyed their tents and the Meunites who were found there, and marked them for destruction to this day, and settled in their place, because there was pasture there for their flocks.
1CHR|4|42|And some of them, five hundred men of the Simeonites, went to Mount Seir, having as their leaders Pelatiah, Neariah, Rephaiah, and Uzziel, the sons of Ishi.
1CHR|4|43|And they defeated the remnant of the Amalekites who had escaped, and they have lived there to this day.
1CHR|5|1|The sons of Reuben the firstborn of Israel (for he was the firstborn, but because he defiled his father's couch, his birthright was given to the sons of Joseph the son of Israel, so that he could not be enrolled as the oldest son;
1CHR|5|2|though Judah became strong among his brothers and a chief came from him, yet the birthright belonged to Joseph),
1CHR|5|3|the sons of Reuben, the firstborn of Israel: Hanoch, Pallu, Hezron, and Carmi.
1CHR|5|4|The sons of Joel: Shemaiah his son, Gog his son, Shimei his son,
1CHR|5|5|Micah his son, Reaiah his son, Baal his son,
1CHR|5|6|Beerah his son, whom Tiglath-pileser king of Assyria carried away into exile; he was a chief of the Reubenites.
1CHR|5|7|And his kinsmen by their clans, when the genealogy of their generations was recorded: the chief, Jeiel, and Zechariah,
1CHR|5|8|and Bela the son of Azaz, son of Shema, son of Joel, who lived in Aroer, as far as Nebo and Baal-meon.
1CHR|5|9|He also lived to the east as far as the entrance of the desert this side of the Euphrates, because their livestock had multiplied in the land of Gilead.
1CHR|5|10|And in the days of Saul they waged war against the Hagrites, who fell into their hand. And they lived in their tents throughout all the region east of Gilead.
1CHR|5|11|The sons of Gad lived over against them in the land of Bashan as far as Salecah:
1CHR|5|12|Joel the chief, Shapham the second, Janai, and Shaphat in Bashan.
1CHR|5|13|And their kinsmen according to their fathers' houses: Michael, Meshullam, Sheba, Jorai, Jacan, Zia and Eber, seven.
1CHR|5|14|These were the sons of Abihail the son of Huri, son of Jaroah, son of Gilead, son of Michael, son of Je-shishai, son of Jahdo, son of Buz.
1CHR|5|15|Ahi the son of Abdiel, son of Guni, was chief in their fathers' houses,
1CHR|5|16|and they lived in Gilead, in Bashan and in its towns, and in all the pasturelands of Sharon to their limits.
1CHR|5|17|All of these were recorded in genealogies in the days of Jotham king of Judah, and in the days of Jeroboam king of Israel.
1CHR|5|18|The Reubenites, the Gadites, and the half-tribe of Manasseh had valiant men who carried shield and sword, and drew the bow, expert in war, 44,760, able to go to war.
1CHR|5|19|They waged war against the Hagrites, Jetur, Naphish, and Nodab.
1CHR|5|20|And when they prevailed over them, the Hagrites and all who were with them were given into their hands, for they cried out to God in the battle, and he granted their urgent plea because they trusted in him.
1CHR|5|21|They carried off their livestock: 50,000 of their camels, 250,000 sheep, 2,000 donkeys, and 100,000 men alive.
1CHR|5|22|For many fell, because the war was of God. And they lived in their place until the exile.
1CHR|5|23|The members of the half-tribe of Manasseh lived in the land. They were very numerous from Bashan to Baal-hermon, Senir, and Mount Hermon.
1CHR|5|24|These were the heads of their fathers' houses: Epher, Ishi, Eliel, Azriel, Jeremiah, Hodaviah, and Jahdiel, mighty warriors, famous men, heads of their fathers' houses.
1CHR|5|25|But they broke faith with the God of their fathers, and whored after the gods of the peoples of the land, whom God had destroyed before them.
1CHR|5|26|So the God of Israel stirred up the spirit of Pul king of Assyria, the spirit of Tiglath-pileser king of Assyria, and he took them into exile, namely, the Reubenites, the Gadites, and the half-tribe of Manasseh, and brought them to Halah, Habor, Hara, and the river Gozan, to this day.
1CHR|6|1|The sons of Levi: Gershon, Kohath, and Merari.
1CHR|6|2|The sons of Kohath: Amram, Izhar, Hebron, and Uzziel.
1CHR|6|3|The children of Amram: Aaron, Moses, and Miriam. The sons of Aaron: Nadab, Abihu, Eleazar, and Ithamar.
1CHR|6|4|Eleazar fathered Phinehas, Phinehas fathered Abishua,
1CHR|6|5|Abishua fathered Bukki, Bukki fathered Uzzi,
1CHR|6|6|Uzzi fathered Zerahiah, Zerahiah fathered Meraioth,
1CHR|6|7|Meraioth fathered Amariah, Amariah fathered Ahitub,
1CHR|6|8|Ahitub fathered Zadok, Zadok fathered Ahimaaz,
1CHR|6|9|Ahimaaz fathered Azariah, Azariah fathered Johanan,
1CHR|6|10|and Johanan fathered Azariah (it was he who served as priest in the house that Solomon built in Jerusalem).
1CHR|6|11|Azariah fathered Amariah, Amariah fathered Ahitub,
1CHR|6|12|Ahitub fathered Zadok, Zadok fathered Shallum,
1CHR|6|13|Shallum fathered Hilkiah, Hilkiah fathered Azariah,
1CHR|6|14|Azariah fathered Seraiah, Seraiah fathered Jehozadak;
1CHR|6|15|and Jehozadak went into exile when the LORD sent Judah and Jerusalem into exile by the hand of Nebuchadnezzar.
1CHR|6|16|The sons of Levi: Gershom, Kohath, and Merari.
1CHR|6|17|And these are the names of the sons of Gershom: Libni and Shimei.
1CHR|6|18|The sons of Kohath: Amram, Izhar, Hebron and Uzziel.
1CHR|6|19|The sons of Merari: Mahli and Mushi. These are the clans of the Levites according to their fathers.
1CHR|6|20|Of Gershom: Libni his son, Jahath his son, Zimmah his son,
1CHR|6|21|Joah his son, Iddo his son, Zerah his son, Jeatherai his son.
1CHR|6|22|The sons of Kohath: Amminadab his son, Korah his son, Assir his son,
1CHR|6|23|Elkanah his son, Ebiasaph his son, Assir his son,
1CHR|6|24|Tahath his son, Uriel his son, Uzziah his son, and Shaul his son.
1CHR|6|25|The sons of Elkanah: Amasai and Ahimoth,
1CHR|6|26|Elkanah his son, Zophai his son, Nahath his son,
1CHR|6|27|Eliab his son, Jeroham his son, Elkanah his son.
1CHR|6|28|The sons of Samuel: Joel his firstborn, the second Abijah.
1CHR|6|29|The sons of Merari: Mahli, Libni his son, Shimei his son, Uzzah his son,
1CHR|6|30|Shimea his son, Haggiah his son, and Asaiah his son.
1CHR|6|31|These are the men whom David put in charge of the service of song in the house of the LORD after the ark rested there.
1CHR|6|32|They ministered with song before the tabernacle of the tent of meeting until Solomon built the house of the LORD in Jerusalem, and they performed their service according to their order.
1CHR|6|33|These are the men who served and their sons. Of the sons of the Kohathites: Heman the singer the son of Joel, son of Samuel,
1CHR|6|34|son of Elkanah, son of Jeroham, son of Eliel, son of Toah,
1CHR|6|35|son of Zuph, son of Elkanah, son of Mahath, son of Amasai,
1CHR|6|36|son of Elkanah, son of Joel, son of Azariah, son of Zephaniah,
1CHR|6|37|son of Tahath, son of Assir, son of Ebiasaph, son of Korah,
1CHR|6|38|son of Izhar, son of Kohath, son of Levi, son of Israel;
1CHR|6|39|and his brother Asaph, who stood on his right hand, namely, Asaph the son of Berechiah, son of Shimea,
1CHR|6|40|son of Michael, son of Baaseiah, son of Malchijah,
1CHR|6|41|son of Ethni, son of Zerah, son of Adaiah,
1CHR|6|42|son of Ethan, son of Zimmah, son of Shimei,
1CHR|6|43|son of Jahath, son of Gershom, son of Levi.
1CHR|6|44|On the left hand were their brothers, the sons of Merari: Ethan the son of Kishi, son of Abdi, son of Malluch,
1CHR|6|45|son of Hashabiah, son of Amaziah, son of Hilkiah,
1CHR|6|46|son of Amzi, son of Bani, son of Shemer,
1CHR|6|47|son of Mahli, son of Mushi, son of Merari, son of Levi.
1CHR|6|48|And their brothers the Levites were appointed for all the service of the tabernacle of the house of God.
1CHR|6|49|But Aaron and his sons made offerings on the altar of burnt offering and on the altar of incense for all the work of the Most Holy Place, and to make atonement for Israel, according to all that Moses the servant of God had commanded.
1CHR|6|50|These are the sons of Aaron: Eleazar his son, Phinehas his son, Abishua his son,
1CHR|6|51|Bukki his son, Uzzi his son, Zerahiah his son,
1CHR|6|52|Meraioth his son, Amariah his son, Ahitub his son,
1CHR|6|53|Zadok his son, Ahimaaz his son.
1CHR|6|54|These are their dwelling places according to their settlements within their borders: to the sons of Aaron of the clans of Kohathites, for theirs was the first lot,
1CHR|6|55|to them they gave Hebron in the land of Judah and its surrounding pasturelands,
1CHR|6|56|but the fields of the city and its villages they gave to Caleb the son of Jephunneh.
1CHR|6|57|To the sons of Aaron they gave the cities of refuge: Hebron, Libnah with its pasturelands, Jattir, Eshtemoa with its pasturelands,
1CHR|6|58|Hilen with its pasturelands, Debir with its pasturelands,
1CHR|6|59|Ashan with its pasturelands, and Beth-shemesh with its pasturelands;
1CHR|6|60|and from the tribe of Benjamin, Gibeon, Geba with its pasturelands, Alemeth with its pasturelands, and Anathoth with its pasturelands. All their cities throughout their clans were thirteen.
1CHR|6|61|To the rest of the Kohathites were given by lot out of the clan of the tribe, out of the half-tribe, the half of Manasseh, ten cities.
1CHR|6|62|To the Gershomites according to their clans were allotted thirteen cities out of the tribes of Issachar, Asher, Naphtali and Manasseh in Bashan.
1CHR|6|63|To the Merarites according to their clans were allotted twelve cities out of the tribes of Reuben, Gad and Zebulun.
1CHR|6|64|So the people of Israel gave the Levites the cities with their pasturelands.
1CHR|6|65|They gave by lot out of the tribes of Judah, Simeon, and Benjamin these cities that are mentioned by name.
1CHR|6|66|And some of the clans of the sons of Kohath had cities of their territory out of the tribe of Ephraim.
1CHR|6|67|They were given the cities of refuge: Shechem with its pasturelands in the hill country of Ephraim, Gezer with its pasturelands,
1CHR|6|68|Jokmeam with its pasturelands, Beth-horon with its pasturelands,
1CHR|6|69|Aijalon with its pasturelands, Gath-rimmon with its pasturelands,
1CHR|6|70|and out of the half-tribe of Manasseh, Aner with its pasturelands, and Bileam with its pasturelands, for the rest of the clans of the Kohathites.
1CHR|6|71|To the Gershomites were given out of the clan of the half-tribe of Manasseh: Golan in Bashan with its pasturelands and Ashtaroth with its pasturelands;
1CHR|6|72|and out of the tribe of Issachar: Kedesh with its pasturelands, Daberath with its pasturelands,
1CHR|6|73|Ramoth with its pasturelands, and Anem with its pasturelands;
1CHR|6|74|out of the tribe of Asher: Mashal with its pasturelands, Abdon with its pasturelands,
1CHR|6|75|Hukok with its pasturelands, and Rehob with its pasturelands;
1CHR|6|76|and out of the tribe of Naphtali: Kedesh in Galilee with its pasturelands, Hammon with its pasturelands, and Kiriathaim with its pasturelands.
1CHR|6|77|To the rest of the Merarites were allotted out of the tribe of Zebulun: Rimmono with its pasturelands, Tabor with its pasturelands,
1CHR|6|78|and beyond the Jordan at Jericho, on the east side of the Jordan, out of the tribe of Reuben: Bezer in the wilderness with its pasturelands, Jahzah with its pasturelands,
1CHR|6|79|Kedemoth with its pasturelands, and Mephaath with its pasturelands;
1CHR|6|80|and out of the tribe of Gad: Ramoth in Gilead with its pasturelands, Mahanaim with its pasturelands,
1CHR|6|81|Heshbon with its pasturelands, and Jazer with its pasturelands.
1CHR|7|1|The sons of Issachar: Tola, Puah, Jashub, and Shimron, four.
1CHR|7|2|The sons of Tola: Uzzi, Rephaiah, Jeriel, Jahmai, Ibsam, and Shemuel, heads of their fathers' houses, namely of Tola, mighty warriors of their generations, their number in the days of David being 22,600.
1CHR|7|3|The son of Uzzi: Izrahiah. And the sons of Izrahiah: Michael, Obadiah, Joel, and Isshiah, all five of them were chief men.
1CHR|7|4|And along with them, by their generations, according to their fathers' houses, were units of the army for war, 36,000, for they had many wives and sons.
1CHR|7|5|Their kinsmen belonging to all the clans of Issachar were in all 87,000 mighty warriors, enrolled by genealogy.
1CHR|7|6|The sons of Benjamin: Bela, Becher, and Jediael, three.
1CHR|7|7|The sons of Bela: Ezbon, Uzzi, Uzziel, Jerimoth, and Iri, five, heads of fathers' houses, mighty warriors. And their enrollment by genealogies was 22,034.
1CHR|7|8|The sons of Becher: Zemirah, Joash, Eliezer, Elioenai, Omri, Jeremoth, Abijah, Anathoth, and Alemeth. All these were the sons of Becher.
1CHR|7|9|And their enrollment by genealogies, according to their generations, as heads of their fathers' houses, mighty warriors, was 22,200.
1CHR|7|10|The son of Jediael: Bilhan. And the sons of Bilhan: Jeush, Benjamin, Ehud, Chenaanah, Zethan, Tarshish, and Ahish-ahar.
1CHR|7|11|All these were the sons of Jediael according to the heads of their fathers' houses, mighty warriors, 17,200, able to go to war.
1CHR|7|12|And Shuppim and Huppim were the sons of Ir, Hushim the son of Aher.
1CHR|7|13|The sons of Naphtali: Jahziel, Guni, Jezer and Shallum, the descendants of Bilhah.
1CHR|7|14|The sons of Manasseh: Asriel, whom his Aramean concubine bore; she bore Machir the father of Gilead.
1CHR|7|15|And Machir took a wife for Huppim and for Shuppim. The name of his sister was Maacah. And the name of the second was Zelophehad, and Zelophehad had daughters.
1CHR|7|16|And Maacah the wife of Machir bore a son, and she called his name Peresh; and the name of his brother was Sheresh; and his sons were Ulam and Rakem.
1CHR|7|17|The son of Ulam: Bedan. These were the sons of Gilead the son of Machir, son of Manasseh.
1CHR|7|18|And his sister Hammolecheth bore Ishhod, Abiezer and Mahlah.
1CHR|7|19|The sons of Shemida were Ahian, Shechem, Likhi, and Aniam.
1CHR|7|20|The sons of Ephraim: Shuthelah, and Bered his son, Tahath his son, Ele-adah his son, Tahath his son,
1CHR|7|21|Zabad his son, Shuthelah his son, and Ezer and Elead, whom the men of Gath who were born in the land killed, because they came down to raid their livestock.
1CHR|7|22|And Ephraim their father mourned many days, and his brothers came to comfort him.
1CHR|7|23|And Ephraim went in to his wife, and she conceived and bore a son. And he called his name Beriah, because disaster had befallen his house.
1CHR|7|24|His daughter was Sheerah, who built both Lower and Upper Beth-horon, and Uzzen-sheerah.
1CHR|7|25|Rephah was his son, Resheph his son, Telah his son, Tahan his son,
1CHR|7|26|Ladan his son, Ammihud his son, Elishama his son,
1CHR|7|27|Nun his son, Joshua his son.
1CHR|7|28|Their possessions and settlements were Bethel and its towns, and to the east Naaran, and to the west Gezer and its towns, Shechem and its towns, and Ayyah and its towns;
1CHR|7|29|also in possession of the Manassites, Beth-shean and its towns, Taanach and its towns, Megiddo and its towns, Dor and its towns. In these lived the sons of Joseph the son of Israel.
1CHR|7|30|The sons of Asher: Imnah, Ishvah, Ishvi, Beriah, and their sister Serah.
1CHR|7|31|The sons of Beriah: Heber, and Malchiel, who fathered Birzaith.
1CHR|7|32|Heber fathered Japhlet, Shomer, Hotham, and their sister Shua.
1CHR|7|33|The sons of Japhlet: Pasach, Bimhal, and Ashvath. These are the sons of Japhlet.
1CHR|7|34|The sons of Shemer his brother: Rohgah, Jehubbah, and Aram.
1CHR|7|35|The sons of Helem his brother: Zophah, Imna, Shelesh, and Amal.
1CHR|7|36|The sons of Zophah: Suah, Harnepher, Shual, Beri, Imrah.
1CHR|7|37|Bezer, Hod, Shamma, Shilshah, Ithran, and Beera.
1CHR|7|38|The sons of Jether: Jephunneh, Pispa, and Ara.
1CHR|7|39|The sons of Ulla: Arah, Hanniel, and Rizia.
1CHR|7|40|All of these were men of Asher, heads of fathers' houses, approved, mighty warriors, chiefs of the princes. Their number enrolled by genealogies, for service in war, was 26,000 men.
1CHR|8|1|Benjamin fathered Bela his firstborn, Ashbel the second, Aharah the third,
1CHR|8|2|Nohah the fourth, and Rapha the fifth.
1CHR|8|3|And Bela had sons: Addar, Gera, Abihud,
1CHR|8|4|Abishua, Naaman, Ahoah,
1CHR|8|5|Gera, Shephu-phan, and Huram.
1CHR|8|6|These are the sons of Ehud (they were heads of fathers' houses of the inhabitants of Geba, and they were carried into exile to Manahath):
1CHR|8|7|Naaman, Ahijah, and Gera, that is, Heglam, who fathered Uzza and Ahihud.
1CHR|8|8|And Shaharaim fathered sons in the country of Moab after he had sent away Hushim and Baara his wives.
1CHR|8|9|He fathered sons by Hodesh his wife: Jobab, Zibia, Mesha, Malcam,
1CHR|8|10|Jeuz, Sachia, and Mirmah. These were his sons, heads of fathers' houses.
1CHR|8|11|He also fathered sons by Hushim: Abitub and Elpaal.
1CHR|8|12|The sons of Elpaal: Eber, Misham, and Shemed, who built Ono and Lod with its towns,
1CHR|8|13|and Beriah and Shema (they were heads of fathers' houses of the inhabitants of Aijalon, who caused the inhabitants of Gath to flee);
1CHR|8|14|and Ahio, Shashak, and Jeremoth.
1CHR|8|15|Zebadiah, Arad, Eder,
1CHR|8|16|Michael, Ishpah, and Joha were sons of Beriah.
1CHR|8|17|Zebadiah, Meshullam, Hizki, Heber,
1CHR|8|18|Ishmerai, Izliah, and Jobab were the sons of Elpaal.
1CHR|8|19|Jakim, Zichri, Zabdi,
1CHR|8|20|Elienai, Zillethai, Eliel,
1CHR|8|21|Adaiah, Beraiah, and Shimrath were the sons of Shimei.
1CHR|8|22|Ishpan, Eber, Eliel,
1CHR|8|23|Abdon, Zichri, Hanan,
1CHR|8|24|Hananiah, Elam, Anthothijah,
1CHR|8|25|Iphdeiah, and Penuel were the sons of Shashak.
1CHR|8|26|Shamsherai, Shehariah, Athaliah,
1CHR|8|27|Jaareshiah, Elijah, and Zichri were the sons of Jeroham.
1CHR|8|28|These were the heads of fathers' houses, according to their generations, chief men. These lived in Jerusalem.
1CHR|8|29|Jeiel the father of Gibeon lived in Gibeon, and the name of his wife was Maacah.
1CHR|8|30|His firstborn son: Abdon, then Zur, Kish, Baal, Nadab,
1CHR|8|31|Gedor, Ahio, Zecher,
1CHR|8|32|and Mikloth (he fathered Shimeah). Now these also lived opposite their kinsmen in Jerusalem, with their kinsmen.
1CHR|8|33|Ner was the father of Kish, Kish of Saul, Saul of Jonathan, Malchi-shua, Abinadab and Eshbaal;
1CHR|8|34|and the son of Jonathan was Merib-baal; and Merib-baal was the father of Micah.
1CHR|8|35|The sons of Micah: Pithon, Melech, Tarea, and Ahaz.
1CHR|8|36|Ahaz fathered Jehoaddah, and Jehoaddah fathered Alemeth, Azmaveth, and Zimri. Zimri fathered Moza.
1CHR|8|37|Moza fathered Binea; Raphah was his son, Eleasah his son, Azel his son.
1CHR|8|38|Azel had six sons, and these are their names: Azrikam, Bocheru, Ishmael, Sheariah, Obadiah, and Hanan. All these were the sons of Azel.
1CHR|8|39|The sons of Eshek his brother: Ulam his firstborn, Jeush the second, and Eliphelet the third.
1CHR|8|40|The sons of Ulam were men who were mighty warriors, bowmen, having many sons and grandsons, 150. All these were Benjaminites.
1CHR|9|1|So all Israel was recorded in genealogies, and these are written in the Book of the Kings of Israel. And Judah was taken into exile in Babylon because of their breach of faith.
1CHR|9|2|Now the first to dwell again in their possessions in their cities were Israel, the priests, the Levites, and the temple servants.
1CHR|9|3|And some of the people of Judah, Benjamin, Ephraim, and Manasseh lived in Jerusalem:
1CHR|9|4|Uthai the son of Ammihud, son of Omri, son of Imri, son of Bani, from the sons of Perez the son of Judah.
1CHR|9|5|And of the Shilonites: Asaiah the firstborn, and his sons.
1CHR|9|6|Of the sons of Zerah: Jeuel and their kinsmen, 690.
1CHR|9|7|Of the Benjaminites: Sallu the son of Meshullam, son of Hodaviah, son of Hassenuah,
1CHR|9|8|Ibneiah the son of Jeroham, Elah the son of Uzzi, son of Michri, and Meshullam the son of Shephatiah, son of Reuel, son of Ibnijah;
1CHR|9|9|and their kinsmen according to their generations, 956. All these were heads of fathers' houses according to their fathers' houses.
1CHR|9|10|Of the priests: Jedaiah, Jehoiarib, Jachin,
1CHR|9|11|and Azariah the son of Hilkiah, son of Meshullam, son of Zadok, son of Meraioth, son of Ahitub, the chief officer of the house of God;
1CHR|9|12|and Adaiah the son of Jeroham, son of Pashhur, son of Malchijah, and Maasai the son of Adiel, son of Jahzerah, son of Meshullam, son of Meshillemith, son of Immer;
1CHR|9|13|besides their kinsmen, heads of their fathers' houses, 1,760, mighty men for the work of the service of the house of God.
1CHR|9|14|Of the Levites: Shemaiah the son of Hasshub, son of Azrikam, son of Hashabiah, of the sons of Merari;
1CHR|9|15|and Bakbakkar, Heresh, Galal and Mattaniah the son of Mica, son of Zichri, son of Asaph;
1CHR|9|16|and Obadiah the son of Shemaiah, son of Galal, son of Jeduthun, and Berechiah the son of Asa, son of Elkanah, who lived in the villages of the Netophathites.
1CHR|9|17|The gatekeepers were Shallum, Akkub, Talmon, Ahiman, and their kinsmen (Shallum was the chief);
1CHR|9|18|until then they were in the king's gate on the east side as the gatekeepers of the camps of the Levites.
1CHR|9|19|Shallum the son of Kore, son of Ebiasaph, son of Korah, and his kinsmen of his fathers' house, the Korahites, were in charge of the work of the service, keepers of the thresholds of the tent, as their fathers had been in charge of the camp of the LORD, keepers of the entrance.
1CHR|9|20|And Phinehas the son of Eleazar was the chief officer over them in time past; the LORD was with him.
1CHR|9|21|Zechariah the son of Meshelemiah was gatekeeper at the entrance of the tent of meeting.
1CHR|9|22|All these, who were chosen as gatekeepers at the thresholds, were 212. They were enrolled by genealogies in their villages. David and Samuel the seer established them in their office of trust.
1CHR|9|23|So they and their sons were in charge of the gates of the house of the LORD, that is, the house of the tent, as guards.
1CHR|9|24|The gatekeepers were on the four sides, east, west, north, and south.
1CHR|9|25|And their kinsmen who were in their villages were obligated to come in every seven days, in turn, to be with these,
1CHR|9|26|for the four chief gatekeepers, who were Levites, were entrusted to be over the chambers and the treasures of the house of God.
1CHR|9|27|And they lodged around the house of God, for on them lay the duty of watching, and they had charge of opening it every morning.
1CHR|9|28|Some of them had charge of the utensils of service, for they were required to count them when they were brought in and taken out.
1CHR|9|29|Others of them were appointed over the furniture and over all the holy utensils, also over the fine flour, the wine, the oil, the incense, and the spices.
1CHR|9|30|Others, of the sons of the priests, prepared the mixing of the spices,
1CHR|9|31|and Mattithiah, one of the Levites, the firstborn of Shallum the Korahite, was entrusted with making the flat cakes.
1CHR|9|32|Also some of their kinsmen of the Kohathites had charge of the showbread, to prepare it every Sabbath.
1CHR|9|33|Now these, the singers, the heads of fathers' houses of the Levites, were in the chambers of the temple free from other service, for they were on duty day and night.
1CHR|9|34|These were heads of fathers' houses of the Levites, according to their generations, leaders. These lived in Jerusalem.
1CHR|9|35|In Gibeon lived the father of Gibeon, Jeiel, and the name of his wife was Maacah,
1CHR|9|36|and his firstborn son Abdon, then Zur, Kish, Baal, Ner, Nadab,
1CHR|9|37|Gedor, Ahio, Zechariah, and Mikloth;
1CHR|9|38|and Mikloth was the father of Shimeam; and these also lived opposite their kinsmen in Jerusalem, with their kinsmen.
1CHR|9|39|Ner fathered Kish, Kish fathered Saul, Saul fathered Jonathan, Malchi-shua, Abinadab, and Eshbaal.
1CHR|9|40|And the son of Jonathan was Merib-baal, and Merib-baal fathered Micah.
1CHR|9|41|The sons of Micah: Pithon, Melech, Tahrea, and Ahaz.
1CHR|9|42|And Ahaz fathered Jarah, and Jarah fathered Alemeth, Azmaveth, and Zimri. And Zimri fathered Moza.
1CHR|9|43|Moza fathered Binea, and Rephaiah was his son, Eleasah his son, Azel his son.
1CHR|9|44|Azel had six sons and these are their names: Azrikam, Bocheru, Ishmael, Sheariah, Obadiah, and Hanan; these were the sons of Azel.
1CHR|10|1|Now the Philistines fought against Israel, and the men of Israel fled before the Philistines and fell slain on Mount Gilboa.
1CHR|10|2|And the Philistines overtook Saul and his sons, and the Philistines struck down Jonathan and Abinadab and Malchi-shua, the sons of Saul.
1CHR|10|3|The battle pressed hard against Saul, and the archers found him, and he was wounded by the archers.
1CHR|10|4|Then Saul said to his armor-bearer, "Draw your sword and thrust me through with it, lest these uncircumcised come and mistreat me." But his armor-bearer would not, for he feared greatly. Therefore Saul took his own sword and fell upon it.
1CHR|10|5|And when his armor-bearer saw that Saul was dead, he also fell upon his sword and died.
1CHR|10|6|Thus Saul died; he and his three sons and all his house died together.
1CHR|10|7|And when all the men of Israel who were in the valley saw that the army had fled and that Saul and his sons were dead, they abandoned their cities and fled, and the Philistines came and lived in them.
1CHR|10|8|The next day, when the Philistines came to strip the slain, they found Saul and his sons fallen on Mount Gilboa.
1CHR|10|9|And they stripped him and took his head and his armor, and sent messengers throughout the land of the Philistines to carry the good news to their idols and to the people.
1CHR|10|10|And they put his armor in the temple of their gods and fastened his head in the temple of Dagon.
1CHR|10|11|But when all Jabesh-gilead heard all that the Philistines had done to Saul,
1CHR|10|12|all the valiant men arose and took away the body of Saul and the bodies of his sons, and brought them to Jabesh. And they buried their bones under the oak in Jabesh and fasted seven days.
1CHR|10|13|So Saul died for his breach of faith. He broke faith with the LORD in that he did not keep the command of the LORD, and also consulted a medium, seeking guidance.
1CHR|10|14|He did not seek guidance from the LORD. Therefore the LORD put him to death and turned the kingdom over to David the son of Jesse.
1CHR|11|1|Then all Israel gathered together to David at Hebron and said, "Behold, we are your bone and flesh.
1CHR|11|2|In times past, even when Saul was king, it was you who led out and brought in Israel. And the LORD your God said to you, 'You shall be shepherd of my people Israel, and you shall be prince over my people Israel.'"
1CHR|11|3|So all the elders of Israel came to the king at Hebron, and David made a covenant with them at Hebron before the LORD. And they anointed David king over Israel, according to the word of the LORD by Samuel.
1CHR|11|4|And David and all Israel went to Jerusalem, that is Jebus, where the Jebusites were, the inhabitants of the land.
1CHR|11|5|The inhabitants of Jebus said to David, "You will not come in here." Nevertheless, David took the stronghold of Zion, that is, the city of David.
1CHR|11|6|David said, "Whoever strikes the Jebusites first shall be chief and commander." And Joab the son of Zeruiah went up first, so he became chief.
1CHR|11|7|And David lived in the stronghold; therefore it was called the city of David.
1CHR|11|8|And he built the city all around from the Millo in complete circuit, and Joab repaired the rest of the city.
1CHR|11|9|And David became greater and greater, for the LORD of hosts was with him.
1CHR|11|10|Now these are the chiefs of David's mighty men, who gave him strong support in his kingdom, together with all Israel, to make him king, according to the word of the LORD concerning Israel.
1CHR|11|11|This is an account of David's mighty men: Jashobeam, a Hachmonite, was chief of the three. He wielded his spear against 300 whom he killed at one time.
1CHR|11|12|And next to him among the three mighty men was Eleazar the son of Dodo, the Ahohite.
1CHR|11|13|He was with David at Pas-dammim when the Philistines were gathered there for battle. There was a plot of ground full of barley, and the men fled from the Philistines.
1CHR|11|14|But he took his stand in the midst of the plot and defended it and killed the Philistines. And the LORD saved them by a great victory.
1CHR|11|15|Three of the thirty chief men went down to the rock to David at the cave of Adullam, when the army of Philistines was encamped in the Valley of Rephaim.
1CHR|11|16|David was then in the stronghold, and the garrison of the Philistines was then at Bethlehem.
1CHR|11|17|And David said longingly, "Oh that someone would give me water to drink from the well of Bethlehem that is by the gate!"
1CHR|11|18|Then the three mighty men broke through the camp of the Philistines and drew water out of the well of Bethlehem that was by the gate and took it and brought it to David. But David would not drink it. He poured it out to the LORD
1CHR|11|19|and said, "Far be it from me before my God that I should do this. Shall I drink the lifeblood of these men? For at the risk of their lives they brought it." Therefore he would not drink it. These things did the three mighty men.
1CHR|11|20|Now Abishai, the brother of Joab, was chief of the thirty. And he wielded his spear against 300 men and killed them and won a name beside the three.
1CHR|11|21|He was the most renowned of the thirty and became their commander, but he did not attain to the three.
1CHR|11|22|And Benaiah the son of Jehoiada was a valiant man of Kabzeel, a doer of great deeds. He struck down two heroes of Moab. He also went down and struck down a lion in a pit on a day when snow had fallen.
1CHR|11|23|And he struck down an Egyptian, a man of great stature, five cubits tall. The Egyptian had in his hand a spear like a weaver's beam, but Benaiah went down to him with a staff and snatched the spear out of the Egyptian's hand and killed him with his own spear.
1CHR|11|24|These things did Benaiah the son of Jehoiada and won a name beside the three mighty men.
1CHR|11|25|He was renowned among the thirty, but he did not attain to the three. And David set him over his bodyguard.
1CHR|11|26|The mighty men were Asahel the brother of Joab, Elhanan the son of Dodo of Bethlehem,
1CHR|11|27|Shammoth of Harod, Helez the Pelonite,
1CHR|11|28|Ira the son of Ikkesh of Tekoa, Abiezer of Anathoth,
1CHR|11|29|Sibbecai the Hushathite, Ilai the Ahohite,
1CHR|11|30|Maharai of Netophah, Heled the son of Baanah of Netophah,
1CHR|11|31|Ithai the son of Ribai of Gibeah of the people of Benjamin, Benaiah of Pirathon,
1CHR|11|32|Hurai of the brooks of Gaash, Abiel the Arbathite,
1CHR|11|33|Azmaveth of Baharum, Eliahba the Shaalbonite,
1CHR|11|34|Hashem the Gizonite, Jonathan the son of Shagee the Hararite,
1CHR|11|35|Ahiam the son of Sachar the Hararite, Eliphal the son of Ur,
1CHR|11|36|Hepher the Mecherathite, Ahijah the Pelonite,
1CHR|11|37|Hezro of Carmel, Naarai the son of Ezbai,
1CHR|11|38|Joel the brother of Nathan, Mibhar the son of Hagri,
1CHR|11|39|Zelek the Ammonite, Naharai of Beeroth, the armor-bearer of Joab the son of Zeruiah,
1CHR|11|40|Ira the Ithrite, Gareb the Ithrite,
1CHR|11|41|Uriah the Hittite, Zabad the son of Ahlai,
1CHR|11|42|Adina the son of Shiza the Reubenite, a leader of the Reubenites, and thirty with him,
1CHR|11|43|Hanan the son of Maacah, and Joshaphat the Mithnite,
1CHR|11|44|Uzzia the Ashterathite, Shama and Jeiel the sons of Hotham the Aroerite,
1CHR|11|45|Jediael the son of Shimri, and Joha his brother, the Tizite,
1CHR|11|46|Eliel the Mahavite, and Jeribai, and Joshaviah, the sons of Elnaam, and Ithmah the Moabite,
1CHR|11|47|Eliel, and Obed, and Jaasiel the Mezobaite.
1CHR|12|1|Now these are the men who came to David at Ziklag, while he could not move about freely because of Saul the son of Kish. And they were among the mighty men who helped him in war.
1CHR|12|2|They were bowmen and could shoot arrows and sling stones with either the right or the left hand; they were Benjaminites, Saul's kinsmen.
1CHR|12|3|The chief was Ahiezer, then Joash, both sons of Shemaah of Gibeah; also Jeziel and Pelet, the sons of Azmaveth; Beracah, Jehu of Anathoth,
1CHR|12|4|Ishmaiah of Gibeon, a mighty man among the thirty and a leader over the thirty; Jeremiah, Jahaziel, Johanan, Jozabad of Gederah,
1CHR|12|5|Eluzai, Jerimoth, Bealiah, Shemariah, Shephatiah the Haruphite;
1CHR|12|6|Elkanah, Isshiah, Azarel, Joezer, and Jashobeam, the Korahites;
1CHR|12|7|And Joelah and Zebadiah, the sons of Jeroham of Gedor.
1CHR|12|8|From the Gadites there went over to David at the stronghold in the wilderness mighty and experienced warriors, expert with shield and spear, whose faces were like the faces of lions and who were swift as gazelles upon the mountains:
1CHR|12|9|Ezer the chief, Obadiah second, Eliab third,
1CHR|12|10|Mishmannah fourth, Jeremiah fifth,
1CHR|12|11|Attai sixth, Eliel seventh,
1CHR|12|12|Johanan eighth, Elzabad ninth,
1CHR|12|13|Jeremiah tenth, Machbannai eleventh.
1CHR|12|14|These Gadites were officers of the army; the least was a match for a hundred men and the greatest for a thousand.
1CHR|12|15|These are the men who crossed the Jordan in the first month, when it was overflowing all its banks, and put to flight all those in the valleys, to the east and to the west.
1CHR|12|16|And some of the men of Benjamin and Judah came to the stronghold to David.
1CHR|12|17|David went out to meet them and said to them, "If you have come to me in friendship to help me, my heart will be joined to you; but if to betray me to my adversaries, although there is no wrong in my hands, then may the God of our fathers see and rebuke you."
1CHR|12|18|Then the Spirit clothed Amasai, chief of the thirty, and he said, "We are yours, O David, and with you, O son of Jesse! Peace, peace to you, and peace to your helpers! For your God helps you." Then David received them and made them officers of his troops.
1CHR|12|19|Some of the men of Manasseh deserted to David when he came with the Philistines for the battle against Saul. (Yet he did not help them, for the rulers of the Philistines took counsel and sent him away, saying, "At peril to our heads he will desert to his master Saul.")
1CHR|12|20|As he went to Ziklag, these men of Manasseh deserted to him: Adnah, Jozabad, Jediael, Michael, Jozabad, Elihu, and Zillethai, chiefs of thousands in Manasseh.
1CHR|12|21|They helped David against the band of raiders, for they were all mighty men of valor and were commanders in the army.
1CHR|12|22|For from day to day men came to David to help him, until there was a great army, like an army of God.
1CHR|12|23|These are the numbers of the divisions of the armed troops who came to David in Hebron to turn the kingdom of Saul over to him, according to the word of the LORD.
1CHR|12|24|The men of Judah bearing shield and spear were 6,800 armed troops.
1CHR|12|25|Of the Simeonites, mighty men of valor for war, 7,100.
1CHR|12|26|Of the Levites 4,600.
1CHR|12|27|The prince Jehoiada, of the house of Aaron, and with him 3,700.
1CHR|12|28|Zadok, a young man mighty in valor, and twenty-two commanders from his own fathers' house.
1CHR|12|29|Of the Benjaminites, the kinsmen of Saul, 3,000, of whom the majority had to that point kept their allegiance to the house of Saul.
1CHR|12|30|Of the Ephraimites 20,800, mighty men of valor, famous men in their fathers' houses.
1CHR|12|31|Of the half-tribe of Manasseh 18,000, who were expressly named to come and make David king.
1CHR|12|32|Of Issachar, men who had understanding of the times, to know what Israel ought to do, 200 chiefs, and all their kinsmen under their command.
1CHR|12|33|Of Zebulun 50,000 seasoned troops, equipped for battle with all the weapons of war, to help David with singleness of purpose.
1CHR|12|34|Of Naphtali 1,000 commanders with whom were 37,000 men armed with shield and spear.
1CHR|12|35|Of the Danites 28,600 men equipped for battle.
1CHR|12|36|Of Asher 40,000 seasoned troops ready for battle.
1CHR|12|37|Of the Reubenites and Gadites and the half-tribe of Manasseh from beyond the Jordan, 120,000 men armed with all the weapons of war.
1CHR|12|38|All these, men of war, arrayed in battle order, came to Hebron with full intent to make David king over all Israel. Likewise, all the rest of Israel were of a single mind to make David king.
1CHR|12|39|And they were there with David for three days, eating and drinking, for their brothers had made preparation for them.
1CHR|12|40|And also their relatives, from as far as Issachar and Zebulun and Naphtali, came bringing food on donkeys and on camels and on mules and on oxen, abundant provisions of flour, cakes of figs, clusters of raisins, and wine and oil, oxen and sheep, for there was joy in Israel.
1CHR|13|1|David consulted with the commanders of thousands and of hundreds, with every leader.
1CHR|13|2|And David said to all the assembly of Israel, "If it seems good to you and from the LORD our God, let us send abroad to our brothers who remain in all the lands of Israel, as well as to the priests and Levites in the cities that have pasturelands, that they may be gathered to us.
1CHR|13|3|Then let us bring again the ark of our God to us, for we did not seek it in the days of Saul."
1CHR|13|4|All the assembly agreed to do so, for the thing was right in the eyes of all the people.
1CHR|13|5|So David assembled all Israel from the Nile of Egypt to Lebo-hamath, to bring the ark of God from Kiriath-jearim.
1CHR|13|6|And David and all Israel went up to Baalah, that is, to Kiriath-jearim that belongs to Judah, to bring up from there the ark of God, which is called by the name of the LORD who sits enthroned above the cherubim.
1CHR|13|7|And they carried the ark of God on a new cart, from the house of Abinadab, and Uzzah and Ahio were driving the cart.
1CHR|13|8|And David and all Israel were rejoicing before God with all their might, with song and lyres and harps and tambourines and cymbals and trumpets.
1CHR|13|9|And when they came to the threshing floor of Chidon, Uzzah put out his hand to take hold of the ark, for the oxen stumbled.
1CHR|13|10|And the anger of the LORD was kindled against Uzzah, and he struck him down because he put out his hand to the ark, and he died there before God.
1CHR|13|11|And David was angry because the LORD had broken out against Uzzah. And that place is called Perez-uzza to this day.
1CHR|13|12|And David was afraid of God that day, and he said, "How can I bring the ark of God home to me?"
1CHR|13|13|So David did not take the ark home into the city of David, but took it aside to the house of Obed-edom the Gittite.
1CHR|13|14|And the ark of God remained with the household of Obed-edom in his house three months. And the LORD blessed the household of Obed-edom and all that he had.
1CHR|14|1|And Hiram king of Tyre sent messengers to David, and cedar trees, also masons and carpenters to build a house for him.
1CHR|14|2|And David knew that the LORD had established him as king over Israel, and that his kingdom was highly exalted for the sake of his people Israel.
1CHR|14|3|And David took more wives in Jerusalem, and David fathered more sons and daughters.
1CHR|14|4|These are the names of the children born to him in Jerusalem: Shammua, Shobab, Nathan, Solomon,
1CHR|14|5|Ibhar, Elishua, Elpelet,
1CHR|14|6|Nogah, Nepheg, Japhia,
1CHR|14|7|Elishama, Beeliada and Eliphelet.
1CHR|14|8|When the Philistines heard that David had been anointed king over all Israel, all the Philistines went up to search for David. But David heard of it and went out against them.
1CHR|14|9|Now the Philistines had come and made a raid in the Valley of Rephaim.
1CHR|14|10|And David inquired of God, "Shall I go up against the Philistines? Will you give them into my hand?" And the LORD said to him, "Go up, and I will give them into your hand."
1CHR|14|11|And he went up to Baal-perazim, and David struck them down there. And David said, "God has broken through my enemies by my hand, like a bursting flood." Therefore the name of that place is called Baal-perazim.
1CHR|14|12|And they left their gods there, and David gave command, and they were burned.
1CHR|14|13|And the Philistines yet again made a raid in the valley.
1CHR|14|14|And when David again inquired of God, God said to him, "You shall not go up after them; go around and come against them opposite the balsam trees.
1CHR|14|15|And when you hear the sound of marching in the tops of the balsam trees, then go out to battle, for God has gone out before you to strike down the army of the Philistines."
1CHR|14|16|And David did as God commanded him, and they struck down the Philistine army from Gibeon to Gezer.
1CHR|14|17|And the fame of David went out into all lands, and the LORD brought the fear of him upon all nations.
1CHR|15|1|David built houses for himself in the city of David. And he prepared a place for the ark of God and pitched a tent for it.
1CHR|15|2|Then David said that no one but the Levites may carry the ark of God, for the LORD had chosen them to carry the ark of the LORD and to minister to him forever.
1CHR|15|3|And David assembled all Israel at Jerusalem to bring up the ark of the LORD to its place, which he had prepared for it.
1CHR|15|4|And David gathered together the sons of Aaron and the Levites:
1CHR|15|5|of the sons of Kohath, Uriel the chief, with 120 of his brothers;
1CHR|15|6|of the sons of Merari, Asaiah the chief, with 220 of his brothers;
1CHR|15|7|of the sons of Gershom, Joel the chief, with 130 of his brothers;
1CHR|15|8|of the sons of Elizaphan, Shemaiah the chief, with 200 of his brothers;
1CHR|15|9|of the sons of Hebron, Eliel the chief, with 80 of his brothers;
1CHR|15|10|of the sons of Uzziel, Amminadab the chief, with 112 of his brothers.
1CHR|15|11|Then David summoned the priests Zadok and Abiathar, and the Levites Uriel, Asaiah, Joel, Shemaiah, Eliel, and Amminadab,
1CHR|15|12|and said to them, "You are the heads of the fathers' houses of the Levites. Consecrate yourselves, you and your brothers, so that you may bring up the ark of the LORD, the God of Israel, to the place that I have prepared for it.
1CHR|15|13|Because you did not carry it the first time, the LORD our God broke out against us, because we did not seek him according to the rule."
1CHR|15|14|So the priests and the Levites consecrated themselves to bring up the ark of the LORD, the God of Israel.
1CHR|15|15|And the Levites carried the ark of God on their shoulders with the poles, as Moses had commanded according to the word of the LORD.
1CHR|15|16|David also commanded the chiefs of the Levites to appoint their brothers as the singers who should play loudly on musical instruments, on harps and lyres and cymbals, to raise sounds of joy.
1CHR|15|17|So the Levites appointed Heman the son of Joel; and of his brothers Asaph the son of Berechiah; and of the sons of Merari, their brothers, Ethan the son of Kushaiah;
1CHR|15|18|and with them their brothers of the second order, Zechariah, Jaaziel, Shemiramoth, Jehiel, Unni, Eliab, Benaiah, Maaseiah, Mattithiah, Eliphelehu, and Mikneiah, and the gatekeepers Obed-edom and Jeiel.
1CHR|15|19|The singers, Heman, Asaph, and Ethan, were to sound bronze cymbals;
1CHR|15|20|Zechariah, Aziel, Shemiramoth, Jehiel, Unni, Eliab, Maaseiah, and Benaiah were to play harps according to Alamoth;
1CHR|15|21|but Mattithiah, Eliphelehu, Mikneiah, Obed-edom, Jeiel, and Azaziah were to lead with lyres according to the Sheminith.
1CHR|15|22|Chenaniah, leader of the Levites in music, should direct the music, for he understood it.
1CHR|15|23|Berechiah and Elkanah were to be gatekeepers for the ark.
1CHR|15|24|Shebaniah, Joshaphat, Nethanel, Amasai, Zechariah, Benaiah, and Eliezer, the priests, should blow the trumpets before the ark of God. Obed-edom and Jehiah were to be gatekeepers for the ark.
1CHR|15|25|So David and the elders of Israel and the commanders of thousands went to bring up the ark of the covenant of the LORD from the house of Obed-edom with rejoicing.
1CHR|15|26|And because God helped the Levites who were carrying the ark of the covenant of the LORD, they sacrificed seven bulls and seven rams.
1CHR|15|27|David was clothed with a robe of fine linen, as also were all the Levites who were carrying the ark, and the singers and Chenaniah the leader of the music of the singers. And David wore a linen ephod.
1CHR|15|28|So all Israel brought up the ark of the covenant of the LORD with shouting, to the sound of the horn, trumpets, and cymbals, and made loud music on harps and lyres.
1CHR|15|29|And as the ark of the covenant of the LORD came to the city of David, Michal the daughter of Saul looked out of the window and saw King David dancing and rejoicing, and she despised him in her heart.
1CHR|16|1|And they brought in the ark of God and set it inside the tent that David had pitched for it, and they offered burnt offerings and peace offerings before God.
1CHR|16|2|And when David had finished offering the burnt offerings and the peace offerings, he blessed the people in the name of the LORD
1CHR|16|3|and distributed to all Israel, both men and women, to each a loaf of bread, a portion of meat, and a cake of raisins.
1CHR|16|4|Then he appointed some of the Levites as ministers before the ark of the LORD, to invoke, to thank, and to praise the LORD, the God of Israel.
1CHR|16|5|Asaph was the chief, and second to him were Zechariah, Jeiel, Shemiramoth, Jehiel, Mattithiah, Eliab, Benaiah, Obed-edom, and Jeiel, who were to play harps and lyres; Asaph was to sound the cymbals,
1CHR|16|6|and Benaiah and Jahaziel the priests were to blow trumpets regularly before the ark of the covenant of God.
1CHR|16|7|Then on that day David first appointed that thanksgiving be sung to the LORD by Asaph and his brothers.
1CHR|16|8|Oh give thanks to the LORD; call upon his name; make known his deeds among the peoples!
1CHR|16|9|Sing to him; sing praises to him; tell of all his wondrous works!
1CHR|16|10|Glory in his holy name; let the hearts of those who seek the LORD rejoice!
1CHR|16|11|Seek the LORD and his strength; seek his presence continually!
1CHR|16|12|Remember the wondrous works that he has done, his miracles and the judgments he uttered,
1CHR|16|13|O offspring of Israel his servant, sons of Jacob, his chosen ones!
1CHR|16|14|He is the LORD our God; his judgments are in all the earth.
1CHR|16|15|Remember his covenant forever, the word that he commanded, for a thousand generations,
1CHR|16|16|the covenant that he made with Abraham, his sworn promise to Isaac,
1CHR|16|17|which he confirmed as a statute to Jacob, as an everlasting covenant to Israel,
1CHR|16|18|saying, "To you I will give the land of Canaan, as your portion for an inheritance."
1CHR|16|19|When you were few in number, and of little account, and sojourners in it,
1CHR|16|20|wandering from nation to nation, from one kingdom to another people,
1CHR|16|21|he allowed no one to oppress them; he rebuked kings on their account,
1CHR|16|22|saying, "Touch not my anointed ones, do my prophets no harm!"
1CHR|16|23|Sing to the LORD, all the earth! Tell of his salvation from day to day.
1CHR|16|24|Declare his glory among the nations, his marvelous works among all the peoples!
1CHR|16|25|For great is the LORD, and greatly to be praised, and he is to be held in awe above all gods.
1CHR|16|26|For all the gods of the peoples are idols, but the LORD made the heavens.
1CHR|16|27|Splendor and majesty are before him; strength and joy are in his place.
1CHR|16|28|Ascribe to the LORD, O clans of the peoples, ascribe to the LORD glory and strength!
1CHR|16|29|Ascribe to the LORD the glory due his name; bring an offering and come before him! Worship the LORD in the splendor of holiness;
1CHR|16|30|tremble before him, all the earth; yes, the world is established; it shall never be moved.
1CHR|16|31|Let the heavens be glad, and let the earth rejoice, and let them say among the nations, "The LORD reigns!"
1CHR|16|32|Let the sea roar, and all that fills it; let the field exult, and everything in it!
1CHR|16|33|Then shall the trees of the forest sing for joy before the LORD, for he comes to judge the earth.
1CHR|16|34|Oh give thanks to the LORD, for he is good; for his steadfast love endures forever!
1CHR|16|35|Say also: "Save us, O God of our salvation, and gather and deliver us from among the nations, that we may give thanks to your holy name, and glory in your praise.
1CHR|16|36|Blessed be the LORD, the God of Israel, from everlasting to everlasting!" Then all the people said, "Amen!" and praised the LORD.
1CHR|16|37|So David left Asaph and his brothers there before the ark of the covenant of the LORD to minister regularly before the ark as each day required,
1CHR|16|38|and also Obed-edom and his sixty-eight brothers, while Obed-edom, the son of Jeduthun, and Hosah were to be gatekeepers.
1CHR|16|39|And he left Zadok the priest and his brothers the priests before the tabernacle of the LORD in the high place that was at Gibeon
1CHR|16|40|to offer burnt offerings to the LORD on the altar of burnt offering regularly morning and evening, to do all that is written in the Law of the LORD that he commanded Israel.
1CHR|16|41|With them were Heman and Jeduthun and the rest of those chosen and expressly named to give thanks to the LORD, for his steadfast love endures forever.
1CHR|16|42|Heman and Jeduthun had trumpets and cymbals for the music and instruments for sacred song. The sons of Jeduthun were appointed to the gate.
1CHR|16|43|Then all the people departed each to his house, and David went home to bless his household.
1CHR|17|1|Now when David lived in his house, David said to Nathan the prophet, "Behold, I dwell in a house of cedar, but the ark of the covenant of the LORD is under a tent."
1CHR|17|2|And Nathan said to David, "Do all that is in your heart, for God is with you."
1CHR|17|3|But that same night the word of the LORD came to Nathan,
1CHR|17|4|"Go and tell my servant David, 'Thus says the LORD: It is not you who will build me a house to dwell in.
1CHR|17|5|For I have not lived in a house since the day I brought up Israel to this day, but I have gone from tent to tent and from dwelling to dwelling.
1CHR|17|6|In all places where I have moved with all Israel, did I speak a word with any of the judges of Israel, whom I commanded to shepherd my people, saying, "Why have you not built me a house of cedar?"'
1CHR|17|7|Now, therefore, thus shall you say to my servant David, 'Thus says the LORD of hosts, I took you from the pasture, from following the sheep, to be prince over my people Israel,
1CHR|17|8|and I have been with you wherever you have gone and have cut off all your enemies from before you. And I will make for you a name, like the name of the great ones of the earth.
1CHR|17|9|And I will appoint a place for my people Israel and will plant them, that they may dwell in their own place and be disturbed no more. And violent men shall waste them no more, as formerly,
1CHR|17|10|from the time that I appointed judges over my people Israel. And I will subdue all your enemies. Moreover, I declare to you that the LORD will build you a house.
1CHR|17|11|When your days are fulfilled to walk with your fathers, I will raise up your offspring after you, one of your own sons, and I will establish his kingdom.
1CHR|17|12|He shall build a house for me, and I will establish his throne forever.
1CHR|17|13|I will be to him a father, and he shall be to me a son. I will not take my steadfast love from him, as I took it from him who was before you,
1CHR|17|14|but I will confirm him in my house and in my kingdom forever, and his throne shall be established forever.'"
1CHR|17|15|In accordance with all these words, and in accordance with all this vision, Nathan spoke to David.
1CHR|17|16|Then King David went in and sat before the LORD and said, "Who am I, O LORD God, and what is my house, that you have brought me thus far?
1CHR|17|17|And this was a small thing in your eyes, O God. You have also spoken of your servant's house for a great while to come, and have shown me future generations, O LORD God!
1CHR|17|18|And what more can David say to you for honoring your servant? For you know your servant.
1CHR|17|19|For your servant's sake, O LORD, and according to your own heart, you have done all this greatness, in making known all these great things.
1CHR|17|20|There is none like you, O LORD, and there is no God besides you, according to all that we have heard with our ears.
1CHR|17|21|And who is like your people Israel, the one nation on earth whom God went to redeem to be his people, making for yourself a name for great and awesome things, in driving out nations before your people whom you redeemed from Egypt?
1CHR|17|22|And you made your people Israel to be your people forever, and you, O LORD, became their God.
1CHR|17|23|And now, O LORD, let the word that you have spoken concerning your servant and concerning his house be established forever, and do as you have spoken,
1CHR|17|24|and your name will be established and magnified forever, saying, 'The LORD of hosts, the God of Israel, is Israel's God,' and the house of your servant David will be established before you.
1CHR|17|25|For you, my God, have revealed to your servant that you will build a house for him. Therefore your servant has found courage to pray before you.
1CHR|17|26|And now, O LORD, you are God, and you have promised this good thing to your servant.
1CHR|17|27|Now you have been pleased to bless the house of your servant, that it may continue forever before you, for it is you, O LORD, who have blessed, and it is blessed forever."
1CHR|18|1|After this David defeated the Philistines and subdued them, and he took Gath and its villages out of the hand of the Philistines.
1CHR|18|2|And he defeated Moab, and the Moabites became servants to David and brought tribute.
1CHR|18|3|David also defeated Hadadezer king of Zobah-Hamath, as he went to set up his monument at the river Euphrates.
1CHR|18|4|And David took from him 1,000 chariots, 7,000 horsemen and 20,000 foot soldiers. And David hamstrung all the chariot horses, but left enough for 100 chariots.
1CHR|18|5|And when the Syrians of Damascus came to help Hadadezer king of Zobah, David struck down 22,000 men of the Syrians.
1CHR|18|6|Then David put garrisons in Syria of Damascus, and the Syrians became servants to David and brought tribute. And the LORD gave victory to David wherever he went.
1CHR|18|7|And David took the shields of gold that were carried by the servants of Hadadezer and brought them to Jerusalem.
1CHR|18|8|And from Tibhath and from Cun, cities of Hadadezer, David took a large amount of bronze. With it Solomon made the bronze sea and the pillars and the vessels of bronze.
1CHR|18|9|When Tou king of Hamath heard that David had defeated the whole army of Hadadezer, king of Zobah,
1CHR|18|10|he sent his son Hadoram to King David, to ask about his health and to bless him because he had fought against Hadadezer and defeated him; for Hadadezer had often been at war with Tou. And he sent all sorts of articles of gold, of silver, and of bronze.
1CHR|18|11|These also King David dedicated to the LORD, together with the silver and gold that he had carried off from all the nations, from Edom, Moab, the Ammonites, the Philistines and Amalek.
1CHR|18|12|And Abishai, the son of Zeruiah, killed 18,000 Edomites in the Valley of Salt.
1CHR|18|13|Then he put garrisons in Edom, and all the Edomites became David's servants. And the LORD gave victory to David wherever he went.
1CHR|18|14|So David reigned over all Israel, and he administered justice and equity to all his people.
1CHR|18|15|And Joab the son of Zeruiah was over the army; and Jehoshaphat the son of Ahilud was recorder;
1CHR|18|16|and Zadok the son of Ahitub and Ahimelech the son of Abiathar were priests; and Shavsha was secretary;
1CHR|18|17|and Benaiah the son of Jehoiada was over the Cherethites and the Pelethites; and David's sons were the chief officials in the service of the king.
1CHR|19|1|Now after this Nahash the king of the Ammonites died, and his son reigned in his place.
1CHR|19|2|And David said, "I will deal kindly with Hanun the son of Nahash, for his father dealt kindly with me." So David sent messengers to console him concerning his father. And David's servants came to the land of the Ammonites to Hanun to console him.
1CHR|19|3|But the princes of the Ammonites said to Hanun, "Do you think, because David has sent comforters to you, that he is honoring your father? Have not his servants come to you to search and to overthrow and to spy out the land?"
1CHR|19|4|So Hanun took David's servants and shaved them and cut off their garments in the middle, at their hips, and sent them away;
1CHR|19|5|and they departed. When David was told concerning the men, he sent messengers to meet them, for the men were greatly ashamed. And the king said, "Remain at Jericho until your beards have grown and then return."
1CHR|19|6|When the Ammonites saw that they had become a stench to David, Hanun and the Ammonites sent 1,000 talents of silver to hire chariots and horsemen from Mesopotamia, from Aram-maacah and from Zobah.
1CHR|19|7|They hired 32,000 chariots and the king of Maacah with his army, who came and encamped before Medeba. And the Ammonites were mustered from their cities and came to battle.
1CHR|19|8|When David heard of it, he sent Joab and all the army of the mighty men.
1CHR|19|9|And the Ammonites came out and drew up in battle array at the entrance of the city, and the kings who had come were by themselves in the open country.
1CHR|19|10|When Joab saw that the battle was set against him both in front and in the rear, he chose some of the best men of Israel and arrayed them against the Syrians.
1CHR|19|11|The rest of his men he put in the charge of Abishai his brother, and they were arrayed against the Ammonites.
1CHR|19|12|And he said, "If the Syrians are too strong for me, then you shall help me, but if the Ammonites are too strong for you, then I will help you.
1CHR|19|13|Be strong, and let us use our strength for our people and for the cities of our God, and may the LORD do what seems good to him."
1CHR|19|14|So Joab and the people who were with him drew near before the Syrians for battle, and they fled before him.
1CHR|19|15|And when the Ammonites saw that the Syrians fled, they likewise fled before Abishai, Joab's brother, and entered the city. Then Joab came to Jerusalem.
1CHR|19|16|But when the Syrians saw that they had been defeated by Israel, they sent messengers and brought out the Syrians who were beyond the Euphrates, with Shophach the commander of the army of Hadadezer at their head.
1CHR|19|17|And when it was told to David, he gathered all Israel together and crossed the Jordan and came to them and drew up his forces against them. And when David set the battle in array against the Syrians, they fought with him.
1CHR|19|18|And the Syrians fled before Israel, and David killed of the Syrians the men of 7,000 chariots and 40,000 foot soldiers, and put to death also Shophach the commander of their army.
1CHR|19|19|And when the servants of Hadadezer saw that they had been defeated by Israel, they made peace with David and became subject to him. So the Syrians were not willing to save the Ammonites any more.
1CHR|20|1|In the spring of the year, the time when kings go out to battle, Joab led out the army and ravaged the country of the Ammonites and came and besieged Rabbah. But David remained at Jerusalem. And Joab struck down Rabbah and overthrew it.
1CHR|20|2|And David took the crown of their king from his head. He found that it weighed a talent of gold, and in it was a precious stone. And it was placed on David's head. And he brought out the spoil of the city, a very great amount.
1CHR|20|3|And he brought out the people who were in it and set them to labor with saws and iron picks and axes. And thus David did to all the cities of the Ammonites. Then David and all the people returned to Jerusalem.
1CHR|20|4|And after this there arose war with the Philistines at Gezer. Then Sibbecai the Hushathite struck down Sippai, who was one of the descendants of the giants, and the Philistines were subdued.
1CHR|20|5|And there was again war with the Philistines, and Elhanan the son of Jair struck down Lahmi the brother of Goliath the Gittite, the shaft of whose spear was like a weaver's beam.
1CHR|20|6|And there was again war at Gath, where there was a man of great stature, who had six fingers on each hand and six toes on each foot, twenty-four in number, and he also was descended from the giants.
1CHR|20|7|And when he taunted Israel, Jonathan the son of Shimea, David's brother, struck him down.
1CHR|20|8|These were descended from the giants in Gath, and they fell by the hand of David and by the hand of his servants.
1CHR|21|1|Then Satan stood against Israel and incited David to number Israel.
1CHR|21|2|So David said to Joab and the commanders of the army, "Go, number Israel, from Beersheba to Dan, and bring me a report, that I may know their number."
1CHR|21|3|But Joab said, "May the LORD add to his people a hundred times as many as they are! Are they not, my lord the king, all of them my lord's servants? Why then should my lord require this? Why should it be a cause of guilt for Israel?"
1CHR|21|4|But the king's word prevailed against Joab. So Joab departed and went throughout all Israel and came back to Jerusalem.
1CHR|21|5|And Joab gave the sum of the numbering of the people to David. In all Israel there were 1,100,000 men who drew the sword, and in Judah 470,000 who drew the sword.
1CHR|21|6|But he did not include Levi and Benjamin in the numbering, for the king's command was abhorrent to Joab.
1CHR|21|7|But God was displeased with this thing, and he struck Israel.
1CHR|21|8|And David said to God, "I have sinned greatly in that I have done this thing. But now, please take away the iniquity of your servant, for I have acted very foolishly."
1CHR|21|9|And the LORD spoke to Gad, David's seer, saying,
1CHR|21|10|"Go and say to David, 'Thus says the LORD, Three things I offer you; choose one of them, that I may do it to you.'"
1CHR|21|11|So Gad came to David and said to him, "Thus says the LORD, 'Choose what you will:
1CHR|21|12|either three years of famine, or three months of devastation by your foes while the sword of your enemies overtakes you, or else three days of the sword of the LORD, pestilence on the land, with the angel of the LORD destroying throughout all the territory of Israel.' Now decide what answer I shall return to him who sent me."
1CHR|21|13|Then David said to Gad, "I am in great distress. Let me fall into the hand of the LORD, for his mercy is very great, but do not let me fall into the hand of man."
1CHR|21|14|So the LORD sent a pestilence on Israel, and 70,000 men of Israel fell.
1CHR|21|15|And God sent the angel to Jerusalem to destroy it, but as he was about to destroy it, the LORD saw, and he relented from the calamity. And he said to the angel who was working destruction, "It is enough; now stay your hand." And the angel of the LORD was standing by the threshing floor of Ornan the Jebusite.
1CHR|21|16|And David lifted his eyes and saw the angel of the LORD standing between earth and heaven, and in his hand a drawn sword stretched out over Jerusalem. Then David and the elders, clothed in sackcloth, fell upon their faces.
1CHR|21|17|And David said to God, "Was it not I who gave command to number the people? It is I who have sinned and done great evil. But these sheep, what have they done? Please let your hand, O LORD my God, be against me and against my father's house. But do not let the plague be on your people."
1CHR|21|18|Now the angel of the LORD had commanded Gad to say to David that David should go up and raise an altar to the LORD on the threshing floor of Ornan the Jebusite.
1CHR|21|19|So David went up at Gad's word, which he had spoken in the name of the LORD.
1CHR|21|20|Now Ornan was threshing wheat. He turned and saw the angel, and his four sons who were with him hid themselves.
1CHR|21|21|As David came to Ornan, Ornan looked and saw David and went out from the threshing floor and paid homage to David with his face to the ground.
1CHR|21|22|And David said to Ornan, "Give me the site of the threshing floor that I may build on it an altar to the LORD- give it to me at its full price- that the plague may be averted from the people."
1CHR|21|23|Then Ornan said to David, "Take it, and let my lord the king do what seems good to him. See, I give the oxen for burnt offerings and the threshing sledges for the wood and the wheat for a grain offering; I give it all."
1CHR|21|24|But King David said to Ornan, "No, but I will buy them for the full price. I will not take for the LORD what is yours, nor offer burnt offerings that cost me nothing."
1CHR|21|25|So David paid Ornan 600 shekels of gold by weight for the site.
1CHR|21|26|And David built there an altar to the LORD and presented burnt offerings and peace offerings and called on the LORD, and the LORD answered him with fire from heaven upon the altar of burnt offering.
1CHR|21|27|Then the LORD commanded the angel, and he put his sword back into its sheath.
1CHR|21|28|At that time, when David saw that the LORD had answered him at the threshing floor of Ornan the Jebusite, he sacrificed there.
1CHR|21|29|For the tabernacle of the LORD, which Moses had made in the wilderness, and the altar of burnt offering were at that time in the high place at Gibeon,
1CHR|21|30|but David could not go before it to inquire of God, for he was afraid of the sword of the angel of the LORD.
1CHR|22|1|Then David said, "Here shall be the house of the LORD God and here the altar of burnt offering for Israel."
1CHR|22|2|David commanded to gather together the resident aliens who were in the land of Israel, and he set stonecutters to prepare dressed stones for building the house of God.
1CHR|22|3|David also provided great quantities of iron for nails for the doors of the gates and for clamps, as well as bronze in quantities beyond weighing,
1CHR|22|4|and cedar timbers without number, for the Sidonians and Tyrians brought great quantities of cedar to David.
1CHR|22|5|For David said, "Solomon my son is young and inexperienced, and the house that is to be built for the LORD must be exceedingly magnificent, of fame and glory throughout all lands. I will therefore make preparation for it." So David provided materials in great quantity before his death.
1CHR|22|6|Then he called for Solomon his son and charged him to build a house for the LORD, the God of Israel.
1CHR|22|7|David said to Solomon, "My son, I had it in my heart to build a house to the name of the LORD my God.
1CHR|22|8|But the word of the LORD came to me, saying, 'You have shed much blood and have waged great wars. You shall not build a house to my name, because you have shed so much blood before me on the earth.
1CHR|22|9|Behold, a son shall be born to you who shall be a man of rest. I will give him rest from all his surrounding enemies. For his name shall be Solomon, and I will give peace and quiet to Israel in his days.
1CHR|22|10|He shall build a house for my name. He shall be my son, and I will be his father, and I will establish his royal throne in Israel forever.'
1CHR|22|11|"Now, my son, the LORD be with you, so that you may succeed in building the house of the LORD your God, as he has spoken concerning you.
1CHR|22|12|Only, may the LORD grant you discretion and understanding, that when he gives you charge over Israel you may keep the law of the LORD your God.
1CHR|22|13|Then you will prosper if you are careful to observe the statutes and the rules that the LORD commanded Moses for Israel. Be strong and courageous. Fear not; do not be dismayed.
1CHR|22|14|With great pains I have provided for the house of the LORD 100,000 talents of gold, a million talents of silver, and bronze and iron beyond weighing, for there is so much of it; timber and stone, too, I have provided. To these you must add.
1CHR|22|15|You have an abundance of workmen: stonecutters, masons, carpenters, and all kinds of craftsmen without number, skilled in working
1CHR|22|16|gold, silver, bronze, and iron. Arise and work! The LORD be with you!"
1CHR|22|17|David also commanded all the leaders of Israel to help Solomon his son, saying,
1CHR|22|18|"Is not the LORD your God with you? And has he not given you peace on every side? For he has delivered the inhabitants of the land into my hand, and the land is subdued before the LORD and his people.
1CHR|22|19|Now set your mind and heart to seek the LORD your God. Arise and build the sanctuary of the LORD God, so that the ark of the covenant of the LORD and the holy vessels of God may be brought into a house built for the name of the LORD."
1CHR|23|1|When David was old and full of days, he made Solomon his son king over Israel.
1CHR|23|2|David assembled all the leaders of Israel and the priests and the Levites.
1CHR|23|3|The Levites, thirty years old and upward, were numbered, and the total was 38,000 men.
1CHR|23|4|"Twenty-four thousand of these," David said, "shall have charge of the work in the house of the LORD, 6,000 shall be officers and judges,
1CHR|23|5|4,000 gatekeepers, and 4,000 shall offer praises to the LORD with the instruments that I have made for praise."
1CHR|23|6|And David organized them in divisions corresponding to the sons of Levi: Gershon, Kohath, and Merari.
1CHR|23|7|The sons of Gershon were Ladan and Shimei.
1CHR|23|8|The sons of Ladan: Jehiel the chief, and Zetham, and Joel, three.
1CHR|23|9|The sons of Shimei: Shelomoth, Haziel, and Haran, three. These were the heads of the fathers' houses of Ladan.
1CHR|23|10|And the sons of Shimei: Jahath, Zina, and Jeush and Beriah. These four were the sons of Shimei.
1CHR|23|11|Jahath was the chief, and Zizah the second; but Jeush and Beriah did not have many sons, therefore they became counted as a single father's house.
1CHR|23|12|The sons of Kohath: Amram, Izhar, Hebron, and Uzziel, four.
1CHR|23|13|The sons of Amram: Aaron and Moses. Aaron was set apart to dedicate the most holy things, that he and his sons forever should make offerings before the LORD and minister to him and pronounce blessings in his name forever.
1CHR|23|14|But the sons of Moses the man of God were named among the tribe of Levi.
1CHR|23|15|The sons of Moses: Gershom and Eliezer.
1CHR|23|16|The sons of Gershom: Shebuel the chief.
1CHR|23|17|The sons of Eliezer: Rehabiah the chief. Eliezer had no other sons, but the sons of Rehabiah were very many.
1CHR|23|18|The sons of Izhar: Shelomith the chief.
1CHR|23|19|The sons of Hebron: Jeriah the chief, Amariah the second, Jahaziel the third, and Jekameam the fourth.
1CHR|23|20|The sons of Uzziel: Micah the chief and Isshiah the second.
1CHR|23|21|The sons of Merari: Mahli and Mushi. The sons of Mahli: Eleazar and Kish.
1CHR|23|22|Eleazar died having no sons, but only daughters; their kinsmen, the sons of Kish, married them.
1CHR|23|23|The sons of Mushi: Mahli, Eder, and Jeremoth, three.
1CHR|23|24|These were the sons of Levi by their fathers' houses, the heads of fathers' houses as they were listed according to the number of the names of the individuals from twenty years old and upward who were to do the work for the service of the house of the LORD.
1CHR|23|25|For David said, "The LORD, the God of Israel, has given rest to his people, and he dwells in Jerusalem forever.
1CHR|23|26|And so the Levites no longer need to carry the tabernacle or any of the things for its service."
1CHR|23|27|For by the last words of David the sons of Levi were numbered from twenty years old and upward.
1CHR|23|28|For their duty was to assist the sons of Aaron for the service of the house of the LORD, having the care of the courts and the chambers, the cleansing of all that is holy, and any work for the service of the house of God.
1CHR|23|29|Their duty was also to assist with the showbread, the flour for the grain offering, the wafers of unleavened bread, the baked offering, the offering mixed with oil, and all measures of quantity or size.
1CHR|23|30|And they were to stand every morning, thanking and praising the LORD, and likewise at evening,
1CHR|23|31|and whenever burnt offerings were offered to the LORD on Sabbaths, new moons and feast days, according to the number required of them, regularly before the LORD.
1CHR|23|32|Thus they were to keep charge of the tent of meeting and the sanctuary, and to attend the sons of Aaron, their brothers, for the service of the house of the LORD.
1CHR|24|1|The divisions of the sons of Aaron were these. The sons of Aaron: Nadab, Abihu, Eleazar, and Ithamar.
1CHR|24|2|But Nadab and Abihu died before their father and had no children, so Eleazar and Ithamar became the priests.
1CHR|24|3|With the help of Zadok of the sons of Eleazar, and Ahimelech of the sons of Ithamar, David organized them according to the appointed duties in their service.
1CHR|24|4|Since more chief men were found among the sons of Eleazar than among the sons of Ithamar, they organized them under sixteen heads of fathers' houses of the sons of Eleazar, and eight of the sons of Ithamar.
1CHR|24|5|They divided them by lot, all alike, for there were sacred officers and officers of God among both the sons of Eleazar and the sons of Ithamar.
1CHR|24|6|And the scribe Shemaiah, the son of Nethanel, a Levite, recorded them in the presence of the king and the princes and Zadok the priest and Ahimelech the son of Abiathar and the heads of the fathers' houses of the priests and of the Levites, one father's house being chosen for Eleazar and one chosen for Ithamar.
1CHR|24|7|The first lot fell to Jehoiarib, the second to Jedaiah,
1CHR|24|8|the third to Harim, the fourth to Seorim,
1CHR|24|9|the fifth to Malchijah, the sixth to Mijamin,
1CHR|24|10|the seventh to Hakkoz, the eighth to Abijah,
1CHR|24|11|the ninth to Jeshua, the tenth to Shecaniah,
1CHR|24|12|the eleventh to Eliashib, the twelfth to Jakim,
1CHR|24|13|the thirteenth to Huppah, the fourteenth to Jeshebeab,
1CHR|24|14|the fifteenth to Bilgah, the sixteenth to Immer,
1CHR|24|15|the seventeenth to Hezir, the eighteenth to Happizzez,
1CHR|24|16|the nineteenth to Pethahiah, the twentieth to Jehezkel,
1CHR|24|17|the twenty-first to Jachin, the twenty-second to Gamul,
1CHR|24|18|the twenty-third to Delaiah, the twenty-fourth to Maaziah.
1CHR|24|19|These had as their appointed duty in their service to come into the house of the LORD according to the procedure established for them by Aaron their father, as the LORD God of Israel had commanded him.
1CHR|24|20|And of the rest of the sons of Levi: of the sons of Amram, Shubael; of the sons of Shubael, Jehdeiah.
1CHR|24|21|Of Rehabiah: of the sons of Rehabiah, Isshiah the chief.
1CHR|24|22|Of the Izharites, Shelomoth; of the sons of Shelomoth, Jahath.
1CHR|24|23|The sons of Hebron: Jeriah the chief, Amariah the second, Jahaziel the third, Jekameam the fourth.
1CHR|24|24|The sons of Uzziel, Micah; of the sons of Micah, Shamir.
1CHR|24|25|The brother of Micah, Isshiah; of the sons of Isshiah, Zechariah.
1CHR|24|26|The sons of Merari: Mahli and Mushi. The sons of Jaaziah: Beno.
1CHR|24|27|The sons of Merari: of Jaaziah, Beno, Shoham, Zaccur and Ibri.
1CHR|24|28|Of Mahli: Eleazar, who had no sons.
1CHR|24|29|Of Kish, the sons of Kish: Jerahmeel.
1CHR|24|30|The sons of Mushi: Mahli, Eder, and Jerimoth. These were the sons of the Levites according to their fathers' houses.
1CHR|24|31|These also, the head of each father's house and his younger brother alike, cast lots, just as their brothers the sons of Aaron, in the presence of King David, Zadok, Ahimelech, and the heads of fathers' houses of the priests and of the Levites.
1CHR|25|1|David and the chiefs of the service also set apart for the service the sons of Asaph, and of Heman, and of Jeduthun, who prophesied with lyres, with harps, and with cymbals. The list of those who did the work and of their duties was:
1CHR|25|2|Of the sons of Asaph: Zaccur, Joseph, Nethaniah, and Asharelah, sons of Asaph, under the direction of Asaph, who prophesied under the direction of the king.
1CHR|25|3|Of Jeduthun, the sons of Jeduthun: Gedaliah, Zeri, Jeshaiah, Shimei, Hashabiah, and Mattithiah, six, under the direction of their father Jeduthun, who prophesied with the lyre in thanksgiving and praise to the LORD.
1CHR|25|4|Of Heman, the sons of Heman: Bukkiah, Mattaniah, Uzziel, Shebuel and Jerimoth, Hananiah, Hanani, Eliathah, Giddalti, and Romamti-ezer, Joshbekashah, Mallothi, Hothir, Mahazioth.
1CHR|25|5|All these were the sons of Heman the king's seer, according to the promise of God to exalt him, for God had given Heman fourteen sons and three daughters.
1CHR|25|6|They were all under the direction of their father in the music in the house of the LORD with cymbals, harps, and lyres for the service of the house of God. Asaph, Jeduthun, and Heman were under the order of the king.
1CHR|25|7|The number of them along with their brothers, who were trained in singing to the LORD, all who were skillful, was 288.
1CHR|25|8|And they cast lots for their duties, small and great, teacher and pupil alike.
1CHR|25|9|The first lot fell for Asaph to Joseph; the second to Gedaliah, to him and his brothers and his sons, twelve;
1CHR|25|10|the third to Zaccur, his sons and his brothers, twelve;
1CHR|25|11|the fourth to Izri, his sons and his brothers, twelve;
1CHR|25|12|the fifth to Nethaniah, his sons and his brothers, twelve;
1CHR|25|13|the sixth to Bukkiah, his sons and his brothers, twelve;
1CHR|25|14|the seventh to Jesharelah, his sons and his brothers, twelve;
1CHR|25|15|the eighth to Jeshaiah, his sons and his brothers, twelve;
1CHR|25|16|the ninth to Mattaniah, his sons and his brothers, twelve;
1CHR|25|17|the tenth to Shimei, his sons and his brothers, twelve;
1CHR|25|18|the eleventh to Azarel, his sons and his brothers, twelve;
1CHR|25|19|the twelfth to Hashabiah, his sons and his brothers, twelve;
1CHR|25|20|to the thirteenth, Shubael, his sons and his brothers, twelve;
1CHR|25|21|to the fourteenth, Mattithiah, his sons and his brothers, twelve;
1CHR|25|22|to the fifteenth, to Jeremoth, his sons and his brothers, twelve;
1CHR|25|23|to the sixteenth, to Hananiah, his sons and his brothers, twelve;
1CHR|25|24|to the seventeenth, to Joshbekashah, his sons and his brothers, twelve;
1CHR|25|25|to the eighteenth, to Hanani, his sons and his brothers, twelve;
1CHR|25|26|to the nineteenth, to Mallothi, his sons and his brothers, twelve;
1CHR|25|27|to the twentieth, to Eliathah, his sons and his brothers, twelve;
1CHR|25|28|to the twenty-first, to Hothir, his sons and his brothers, twelve;
1CHR|25|29|to the twenty-second, to Giddalti, his sons and his brothers, twelve;
1CHR|25|30|to the twenty-third, to Mahazioth, his sons and his brothers, twelve;
1CHR|25|31|to the twenty-fourth, to Romamti-ezer, his sons and his brothers, twelve.
1CHR|26|1|As for the divisions of the gatekeepers: of the Korahites, Meshelemiah the son of Kore, of the sons of Asaph.
1CHR|26|2|And Meshelemiah had sons: Zechariah the firstborn, Jediael the second, Zebadiah the third, Jathniel the fourth,
1CHR|26|3|Elam the fifth, Jehohanan the sixth, Eliehoenai the seventh.
1CHR|26|4|And Obed-edom had sons: Shemaiah the firstborn, Jehozabad the second, Joah the third, Sachar the fourth, Nethanel the fifth,
1CHR|26|5|Ammiel the sixth, Issachar the seventh, Peullethai the eighth, for God blessed him.
1CHR|26|6|Also to his son Shemaiah were sons born who were rulers in their fathers' houses, for they were men of great ability.
1CHR|26|7|The sons of Shemaiah: Othni, Rephael, Obed and Elzabad, whose brothers were able men, Elihu and Semachiah.
1CHR|26|8|All these were of the sons of Obed-edom with their sons and brothers, able men qualified for the service; sixty-two of Obed-edom.
1CHR|26|9|And Meshelemiah had sons and brothers, able men, eighteen.
1CHR|26|10|And Hosah, of the sons of Merari, had sons: Shimri the chief (for though he was not the firstborn, his father made him chief),
1CHR|26|11|Hilkiah the second, Tebaliah the third, Zechariah the fourth: all the sons and brothers of Hosah were thirteen.
1CHR|26|12|These divisions of the gatekeepers, corresponding to their chief men, had duties, just as their brothers did, ministering in the house of the LORD.
1CHR|26|13|And they cast lots by fathers' houses, small and great alike, for their gates.
1CHR|26|14|The lot for the east fell to Shelemiah. They cast lots also for his son Zechariah, a shrewd counselor, and his lot came out for the north.
1CHR|26|15|Obed-edom's came out for the south, and to his sons was allotted the gatehouse.
1CHR|26|16|For Shuppim and Hosah it came out for the west, at the gate of Shallecheth on the road that goes up. Watch corresponded to watch.
1CHR|26|17|On the east there were six each day, on the north four each day, on the south four each day, as well as two and two at the gatehouse.
1CHR|26|18|And for the colonnade on the west there were four at the road and two at the colonnade.
1CHR|26|19|These were the divisions of the gatekeepers among the Korahites and the sons of Merari.
1CHR|26|20|And of the Levites, Ahijah had charge of the treasuries of the house of God and the treasuries of the dedicated gifts.
1CHR|26|21|The sons of Ladan, the sons of the Gershonites belonging to Ladan, the heads of the fathers' houses belonging to Ladan the Gershonite: Jehieli.
1CHR|26|22|The sons of Jehieli, Zetham, and Joel his brother, were in charge of the treasuries of the house of the LORD.
1CHR|26|23|Of the Amramites, the Izharites, the Hebronites, and the Uzzielites-
1CHR|26|24|and Shebuel the son of Gershom, son of Moses, was chief officer in charge of the treasuries.
1CHR|26|25|His brothers: from Eliezer were his son Rehabiah, and his son Jeshaiah, and his son Joram, and his son Zichri, and his son Shelomoth.
1CHR|26|26|This Shelomoth and his brothers were in charge of all the treasuries of the dedicated gifts that David the king and the heads of the fathers' houses and the officers of the thousands and the hundreds and the commanders of the army had dedicated.
1CHR|26|27|From spoil won in battles they dedicated gifts for the maintenance of the house of the LORD.
1CHR|26|28|Also all that Samuel the seer and Saul the son of Kish and Abner the son of Ner and Joab the son of Zeruiah had dedicated- all dedicated gifts were in the care of Shelomoth and his brothers.
1CHR|26|29|Of the Izharites, Chenaniah and his sons were appointed to external duties for Israel, as officers and judges.
1CHR|26|30|Of the Hebronites, Hashabiah and his brothers, 1,700 men of ability, had the oversight of Israel westward of the Jordan for all the work of the LORD and for the service of the king.
1CHR|26|31|Of the Hebronites, Jerijah was chief of the Hebronites of whatever genealogy or fathers' houses. (In the fortieth year of David's reign search was made and men of great ability among them were found at Jazer in Gilead.)
1CHR|26|32|King David appointed him and his brothers, 2,700 men of ability, heads of fathers' houses, to have the oversight of the Reubenites, the Gadites and the half-tribe of the Manassites for everything pertaining to God and for the affairs of the king.
1CHR|27|1|This is the number of the people of Israel, the heads of fathers' houses, the commanders of thousands and hundreds, and their officers who served the king in all matters concerning the divisions that came and went, month after month throughout the year, each division numbering 24,000:
1CHR|27|2|Jashobeam the son of Zabdiel was in charge of the first division in the first month; in his division were 24,000.
1CHR|27|3|He was a descendant of Perez and was chief of all the commanders. He served for the first month.
1CHR|27|4|Dodai the Ahohite was in charge of the division of the second month; in his division were 24,000.
1CHR|27|5|The third commander, for the third month, was Benaiah, the son of Jehoiada the chief priest; in his division were 24,000.
1CHR|27|6|This is the Benaiah who was a mighty man of the thirty and in command of the thirty; Ammizabad his son was in charge of his division.
1CHR|27|7|Asahel the brother of Joab was fourth, for the fourth month, and his son Zebadiah after him; in his division were 24,000.
1CHR|27|8|The fifth commander, for the fifth month, was Shamhuth the Izrahite; in his division were 24,000.
1CHR|27|9|Sixth, for the sixth month, was Ira, the son of Ikkesh the Tekoite; in his division were 24,000.
1CHR|27|10|Seventh, for the seventh month, was Helez the Pelonite, of the sons of Ephraim; in his division were 24,000.
1CHR|27|11|Eighth, for the eighth month, was Sibbecai the Hushathite, of the Zerahites; in his division were 24,000.
1CHR|27|12|Ninth, for the ninth month, was Abiezer of Anathoth, a Benjaminite; in his division were 24,000.
1CHR|27|13|Tenth, for the tenth month, was Maharai of Netophah, of the Zerahites; in his division were 24,000.
1CHR|27|14|Eleventh, for the eleventh month, was Benaiah of Pirathon, of the sons of Ephraim; in his division were 24,000.
1CHR|27|15|Twelfth, for the twelfth month, was Heldai the Netophathite, of Othniel; in his division were 24,000.
1CHR|27|16|Over the tribes of Israel, for the Reubenites, Eliezer the son of Zichri was chief officer; for the Simeonites, Shephatiah the son of Maacah;
1CHR|27|17|for Levi, Hashabiah the son of Kemuel; for Aaron, Zadok;
1CHR|27|18|for Judah, Elihu, one of David's brothers; for Issachar, Omri the son of Michael;
1CHR|27|19|for Zebulun, Ishmaiah the son of Obadiah; for Naphtali, Jeremoth the son of Azriel;
1CHR|27|20|for the Ephraimites, Hoshea the son of Azaziah; for the half-tribe of Manasseh, Joel the son of Pedaiah;
1CHR|27|21|for the half-tribe of Manasseh in Gilead, Iddo the son of Zechariah; for Benjamin, Jaasiel the son of Abner;
1CHR|27|22|for Dan, Azarel the son of Jeroham. These were the leaders of the tribes of Israel.
1CHR|27|23|David did not count those below twenty years of age, for the LORD had promised to make Israel as many as the stars of heaven.
1CHR|27|24|Joab the son of Zeruiah began to count, but did not finish. Yet wrath came upon Israel for this, and the number was not entered in the chronicles of King David.
1CHR|27|25|Over the king's treasuries was Azmaveth the son of Adiel; and over the treasuries in the country, in the cities, in the villages and in the towers, was Jonathan the son of Uzziah;
1CHR|27|26|and over those who did the work of the field for tilling the soil was Ezri the son of Chelub;
1CHR|27|27|and over the vineyards was Shimei the Ramathite; and over the produce of the vineyards for the wine cellars was Zabdi the Shiphmite.
1CHR|27|28|Over the olive and sycamore trees in the Shephelah was Baal-hanan the Gederite; and over the stores of oil was Joash.
1CHR|27|29|Over the herds that pastured in Sharon was Shitrai the Sharonite; over the herds in the valleys was Shaphat the son of Adlai.
1CHR|27|30|Over the camels was Obil the Ishmaelite; and over the donkeys was Jehdeiah the Meronothite. Over the flocks was Jaziz the Hagrite.
1CHR|27|31|All these were stewards of King David's property.
1CHR|27|32|Jonathan, David's uncle, was a counselor, being a man of understanding and a scribe. He and Jehiel the son of Hachmoni attended the king's sons.
1CHR|27|33|Ahithophel was the king's counselor, and Hushai the Archite was the king's friend.
1CHR|27|34|Ahithophel was succeeded by Jehoiada the son of Benaiah, and Abiathar. Joab was commander of the king's army.
1CHR|28|1|David assembled at Jerusalem all the officials of Israel, the officials of the tribes, the officers of the divisions that served the king, the commanders of thousands, the commanders of hundreds, the stewards of all the property and livestock of the king and his sons, together with the palace officials, the mighty men and all the seasoned warriors.
1CHR|28|2|Then King David rose to his feet and said: "Hear me, my brothers and my people. I had it in my heart to build a house of rest for the ark of the covenant of the LORD and for the footstool of our God, and I made preparations for building.
1CHR|28|3|But God said to me, 'You may not build a house for my name, for you are a man of war and have shed blood.'
1CHR|28|4|Yet the LORD God of Israel chose me from all my father's house to be king over Israel forever. For he chose Judah as leader, and in the house of Judah my father's house, and among my father's sons he took pleasure in me to make me king over all Israel.
1CHR|28|5|And of all my sons (for the LORD has given me many sons) he has chosen Solomon my son to sit on the throne of the kingdom of the LORD over Israel.
1CHR|28|6|He said to me, 'It is Solomon your son who shall build my house and my courts, for I have chosen him to be my son, and I will be his father.
1CHR|28|7|I will establish his kingdom forever if he continues strong in keeping my commandments and my rules, as he is today.'
1CHR|28|8|Now therefore in the sight of all Israel, the assembly of the LORD, and in the hearing of our God, observe and seek out all the commandments of the LORD your God, that you may possess this good land and leave it for an inheritance to your children after you forever.
1CHR|28|9|"And you, Solomon my son, know the God of your father and serve him with a whole heart and with a willing mind, for the LORD searches all hearts and understands every plan and thought. If you seek him, he will be found by you, but if you forsake him, he will cast you off forever.
1CHR|28|10|Be careful now, for the LORD has chosen you to build a house for the sanctuary; be strong and do it."
1CHR|28|11|Then David gave Solomon his son the plan of the vestibule of the temple, and of its houses, its treasuries, its upper rooms, and its inner chambers, and of the room for the mercy seat;
1CHR|28|12|and the plan of all that he had in mind for the courts of the house of the LORD, all the surrounding chambers, the treasuries of the house of God, and the treasuries for dedicated gifts;
1CHR|28|13|for the divisions of the priests and of the Levites, and all the work of the service in the house of the LORD; for all the vessels for the service in the house of the LORD,
1CHR|28|14|the weight of gold for all golden vessels for each service, the weight of silver vessels for each service,
1CHR|28|15|the weight of the golden lampstands and their lamps, the weight of gold for each lampstand and its lamps, the weight of silver for a lampstand and its lamps, according to the use of each lampstand in the service,
1CHR|28|16|the weight of gold for each table for the showbread, the silver for the silver tables,
1CHR|28|17|and pure gold for the forks, the basins and the cups; for the golden bowls and the weight of each; for the silver bowls and the weight of each;
1CHR|28|18|for the altar of incense made of refined gold, and its weight; also his plan for the golden chariot of the cherubim that spread their wings and covered the ark of the covenant of the LORD.
1CHR|28|19|All this he made clear to me in writing from the hand of the LORD, all the work to be done according to the plan.
1CHR|28|20|Then David said to Solomon his son, "Be strong and courageous and do it. Do not be afraid and do not be dismayed, for the LORD God, even my God, is with you. He will not leave you or forsake you, until all the work for the service of the house of the LORD is finished.
1CHR|28|21|And behold the divisions of the priests and the Levites for all the service of the house of God; and with you in all the work will be every willing man who has skill for any kind of service; also the officers and all the people will be wholly at your command."
1CHR|29|1|And David the king said to all the assembly, "Solomon my son, whom alone God has chosen, is young and inexperienced, and the work is great, for the palace will not be for man but for the LORD God.
1CHR|29|2|So I have provided for the house of my God, so far as I was able, the gold for the things of gold, the silver for the things of silver, and the bronze for the things of bronze, the iron for the things of iron, and wood for the things of wood, besides great quantities of onyx and stones for setting, antimony, colored stones, all sorts of precious stones and marble.
1CHR|29|3|Moreover, in addition to all that I have provided for the holy house, I have a treasure of my own of gold and silver, and because of my devotion to the house of my God I give it to the house of my God:
1CHR|29|4|3,000 talents of gold, of the gold of Ophir, and 7,000 talents of refined silver, for overlaying the walls of the house,
1CHR|29|5|and for all the work to be done by craftsmen, gold for the things of gold and silver for the things of silver. Who then will offer willingly, consecrating himself today to the LORD?"
1CHR|29|6|Then the leaders of fathers' houses made their freewill offerings, as did also the leaders of the tribes, the commanders of thousands and of hundreds, and the officers over the king's work.
1CHR|29|7|They gave for the service of the house of God 5,000 talents and 10,000 darics of gold, 10,000 talents of silver, 18,000 talents of bronze and 100,000 talents of iron.
1CHR|29|8|And whoever had precious stones gave them to the treasury of the house of the LORD, in the care of Jehiel the Gershonite.
1CHR|29|9|Then the people rejoiced because they had given willingly, for with a whole heart they had offered freely to the LORD. David the king also rejoiced greatly.
1CHR|29|10|Therefore David blessed the LORD in the presence of all the assembly. And David said: "Blessed are you, O LORD, the God of Israel our father, forever and ever.
1CHR|29|11|Yours, O LORD, is the greatness and the power and the glory and the victory and the majesty, for all that is in the heavens and in the earth is yours. Yours is the kingdom, O LORD, and you are exalted as head above all.
1CHR|29|12|Both riches and honor come from you, and you rule over all. In your hand are power and might, and in your hand it is to make great and to give strength to all.
1CHR|29|13|And now we thank you, our God, and praise your glorious name.
1CHR|29|14|"But who am I, and what is my people, that we should be able thus to offer willingly? For all things come from you, and of your own have we given you.
1CHR|29|15|For we are strangers before you and sojourners, as all our fathers were. Our days on the earth are like a shadow, and there is no abiding.
1CHR|29|16|O LORD our God, all this abundance that we have provided for building you a house for your holy name comes from your hand and is all your own.
1CHR|29|17|I know, my God, that you test the heart and have pleasure in uprightness. In the uprightness of my heart I have freely offered all these things, and now I have seen your people, who are present here, offering freely and joyously to you.
1CHR|29|18|O LORD, the God of Abraham, Isaac, and Israel, our fathers, keep forever such purposes and thoughts in the hearts of your people, and direct their hearts toward you.
1CHR|29|19|Grant to Solomon my son a whole heart that he may keep your commandments, your testimonies, and your statutes, performing all, and that he may build the palace for which I have made provision."
1CHR|29|20|Then David said to all the assembly, "Bless the LORD your God." And all the assembly blessed the LORD, the God of their fathers, and bowed their heads and paid homage to the LORD and to the king.
1CHR|29|21|And they offered sacrifices to the LORD, and on the next day offered burnt offerings to the LORD, 1,000 bulls, 1,000 rams, and 1,000 lambs, with their drink offerings, and sacrifices in abundance for all Israel.
1CHR|29|22|And they ate and drank before the LORD on that day with great gladness. And they made Solomon the son of David king the second time, and they anointed him as prince for the LORD, and Zadok as priest.
1CHR|29|23|Then Solomon sat on the throne of the LORD as king in place of David his father. And he prospered, and all Israel obeyed him.
1CHR|29|24|All the leaders and the mighty men, and also all the sons of King David, pledged their allegiance to King Solomon.
1CHR|29|25|And the LORD made Solomon very great in the sight of all Israel and bestowed on him such royal majesty as had not been on any king before him in Israel.
1CHR|29|26|Thus David the son of Jesse reigned over all Israel.
1CHR|29|27|The time that he reigned over Israel was forty years. He reigned seven years in Hebron and thirty-three years in Jerusalem.
1CHR|29|28|Then he died at a good age, full of days, riches, and honor. And Solomon his son reigned in his place.
1CHR|29|29|Now the acts of King David, from first to last, are written in the Chronicles of Samuel the seer, and in the Chronicles of Nathan the prophet, and in the Chronicles of Gad the seer,
1CHR|29|30|with accounts of all his rule and his might and of the circumstances that came upon him and upon Israel and upon all the kingdoms of the countries.
