HEB|1|1|In the past God spoke to our forefathers through the prophets at many times and in various ways,
HEB|1|2|but in these last days he has spoken to us by his Son, whom he appointed heir of all things, and through whom he made the universe.
HEB|1|3|The Son is the radiance of God's glory and the exact representation of his being, sustaining all things by his powerful word. After he had provided purification for sins, he sat down at the right hand of the Majesty in heaven.
HEB|1|4|So he became as much superior to the angels as the name he has inherited is superior to theirs.
HEB|1|5|For to which of the angels did God ever say, "You are my Son; today I have become your Father "? Or again, "I will be his Father, and he will be my Son"?
HEB|1|6|And again, when God brings his firstborn into the world, he says, "Let all God's angels worship him."
HEB|1|7|In speaking of the angels he says, "He makes his angels winds, his servants flames of fire."
HEB|1|8|But about the Son he says, "Your throne, O God, will last for ever and ever, and righteousness will be the scepter of your kingdom.
HEB|1|9|You have loved righteousness and hated wickedness; therefore God, your God, has set you above your companions by anointing you with the oil of joy."
HEB|1|10|He also says, "In the beginning, O Lord, you laid the foundations of the earth, and the heavens are the work of your hands.
HEB|1|11|They will perish, but you remain; they will all wear out like a garment.
HEB|1|12|You will roll them up like a robe; like a garment they will be changed. But you remain the same, and your years will never end."
HEB|1|13|To which of the angels did God ever say, "Sit at my right hand until I make your enemies a footstool for your feet"?
HEB|1|14|Are not all angels ministering spirits sent to serve those who will inherit salvation?
HEB|2|1|We must pay more careful attention, therefore, to what we have heard, so that we do not drift away.
HEB|2|2|For if the message spoken by angels was binding, and every violation and disobedience received its just punishment,
HEB|2|3|how shall we escape if we ignore such a great salvation? This salvation, which was first announced by the Lord, was confirmed to us by those who heard him.
HEB|2|4|God also testified to it by signs, wonders and various miracles, and gifts of the Holy Spirit distributed according to his will.
HEB|2|5|It is not to angels that he has subjected the world to come, about which we are speaking.
HEB|2|6|But there is a place where someone has testified: "What is man that you are mindful of him, the son of man that you care for him?
HEB|2|7|You made him a little lower than the angels; you crowned him with glory and honor
HEB|2|8|and put everything under his feet.? In putting everything under him, God left nothing that is not subject to him. Yet at present we do not see everything subject to him.
HEB|2|9|But we see Jesus, who was made a little lower than the angels, now crowned with glory and honor because he suffered death, so that by the grace of God he might taste death for everyone.
HEB|2|10|In bringing many sons to glory, it was fitting that God, for whom and through whom everything exists, should make the author of their salvation perfect through suffering.
HEB|2|11|Both the one who makes men holy and those who are made holy are of the same family. So Jesus is not ashamed to call them brothers.
HEB|2|12|He says, "I will declare your name to my brothers; in the presence of the congregation I will sing your praises."
HEB|2|13|And again, "I will put my trust in him." And again he says, "Here am I, and the children God has given me."
HEB|2|14|Since the children have flesh and blood, he too shared in their humanity so that by his death he might destroy him who holds the power of death--that is, the devil--
HEB|2|15|and free those who all their lives were held in slavery by their fear of death.
HEB|2|16|For surely it is not angels he helps, but Abraham's descendants.
HEB|2|17|For this reason he had to be made like his brothers in every way, in order that he might become a merciful and faithful high priest in service to God, and that he might make atonement for the sins of the people.
HEB|2|18|Because he himself suffered when he was tempted, he is able to help those who are being tempted.
HEB|3|1|Therefore, holy brothers, who share in the heavenly calling, fix your thoughts on Jesus, the apostle and high priest whom we confess.
HEB|3|2|He was faithful to the one who appointed him, just as Moses was faithful in all God's house.
HEB|3|3|Jesus has been found worthy of greater honor than Moses, just as the builder of a house has greater honor than the house itself.
HEB|3|4|For every house is built by someone, but God is the builder of everything.
HEB|3|5|Moses was faithful as a servant in all God's house, testifying to what would be said in the future.
HEB|3|6|But Christ is faithful as a son over God's house. And we are his house, if we hold on to our courage and the hope of which we boast.
HEB|3|7|So, as the Holy Spirit says: "Today, if you hear his voice,
HEB|3|8|do not harden your hearts as you did in the rebellion, during the time of testing in the desert,
HEB|3|9|where your fathers tested and tried me and for forty years saw what I did.
HEB|3|10|That is why I was angry with that generation, and I said, 'Their hearts are always going astray, and they have not known my ways.'
HEB|3|11|So I declared on oath in my anger, 'They shall never enter my rest.'"
HEB|3|12|See to it, brothers, that none of you has a sinful, unbelieving heart that turns away from the living God.
HEB|3|13|But encourage one another daily, as long as it is called Today, so that none of you may be hardened by sin's deceitfulness.
HEB|3|14|We have come to share in Christ if we hold firmly till the end the confidence we had at first.
HEB|3|15|As has just been said: "Today, if you hear his voice, do not harden your hearts as you did in the rebellion."
HEB|3|16|Who were they who heard and rebelled? Were they not all those Moses led out of Egypt?
HEB|3|17|And with whom was he angry for forty years? Was it not with those who sinned, whose bodies fell in the desert?
HEB|3|18|And to whom did God swear that they would never enter his rest if not to those who disobeyed?
HEB|3|19|So we see that they were not able to enter, because of their unbelief.
HEB|4|1|Therefore, since the promise of entering his rest still stands, let us be careful that none of you be found to have fallen short of it.
HEB|4|2|For we also have had the gospel preached to us, just as they did; but the message they heard was of no value to them, because those who heard did not combine it with faith.
HEB|4|3|Now we who have believed enter that rest, just as God has said, "So I declared on oath in my anger, 'They shall never enter my rest.'"
HEB|4|4|And yet his work has been finished since the creation of the world. For somewhere he has spoken about the seventh day in these words: "And on the seventh day God rested from all his work."
HEB|4|5|And again in the passage above he says, "They shall never enter my rest."
HEB|4|6|It still remains that some will enter that rest, and those who formerly had the gospel preached to them did not go in, because of their disobedience.
HEB|4|7|Therefore God again set a certain day, calling it Today, when a long time later he spoke through David, as was said before: "Today, if you hear his voice, do not harden your hearts."
HEB|4|8|For if Joshua had given them rest, God would not have spoken later about another day.
HEB|4|9|There remains, then, a Sabbath-rest for the people of God;
HEB|4|10|for anyone who enters God's rest also rests from his own work, just as God did from his.
HEB|4|11|Let us, therefore, make every effort to enter that rest, so that no one will fall by following their example of disobedience.
HEB|4|12|For the word of God is living and active. Sharper than any double--edged sword, it penetrates even to dividing soul and spirit, joints and marrow; it judges the thoughts and attitudes of the heart.
HEB|4|13|Nothing in all creation is hidden from God's sight. Everything is uncovered and laid bare before the eyes of him to whom we must give account.
HEB|4|14|Therefore, since we have a great high priest who has gone through the heavens, Jesus the Son of God, let us hold firmly to the faith we profess.
HEB|4|15|For we do not have a high priest who is unable to sympathize with our weaknesses, but we have one who has been tempted in every way, just as we are--yet was without sin.
HEB|4|16|Let us then approach the throne of grace with confidence, so that we may receive mercy and find grace to help us in our time of need.
HEB|5|1|Every high priest is selected from among men and is appointed to represent them in matters related to God, to offer gifts and sacrifices for sins.
HEB|5|2|He is able to deal gently with those who are ignorant and are going astray, since he himself is subject to weakness.
HEB|5|3|This is why he has to offer sacrifices for his own sins, as well as for the sins of the people.
HEB|5|4|No one takes this honor upon himself; he must be called by God, just as Aaron was.
HEB|5|5|So Christ also did not take upon himself the glory of becoming a high priest. But God said to him, "You are my Son; today I have become your Father. "
HEB|5|6|And he says in another place, "You are a priest forever, in the order of Melchizedek."
HEB|5|7|During the days of Jesus' life on earth, he offered up prayers and petitions with loud cries and tears to the one who could save him from death, and he was heard because of his reverent submission.
HEB|5|8|Although he was a son, he learned obedience from what he suffered
HEB|5|9|and, once made perfect, he became the source of eternal salvation for all who obey him
HEB|5|10|and was designated by God to be high priest in the order of Melchizedek.
HEB|5|11|We have much to say about this, but it is hard to explain because you are slow to learn.
HEB|5|12|In fact, though by this time you ought to be teachers, you need someone to teach you the elementary truths of God's word all over again. You need milk, not solid food!
HEB|5|13|Anyone who lives on milk, being still an infant, is not acquainted with the teaching about righteousness.
HEB|5|14|But solid food is for the mature, who by constant use have trained themselves to distinguish good from evil.
HEB|6|1|Therefore let us leave the elementary teachings about Christ and go on to maturity, not laying again the foundation of repentance from acts that lead to death, and of faith in God,
HEB|6|2|instruction about baptisms, the laying on of hands, the resurrection of the dead, and eternal judgment.
HEB|6|3|And God permitting, we will do so.
HEB|6|4|It is impossible for those who have once been enlightened, who have tasted the heavenly gift, who have shared in the Holy Spirit,
HEB|6|5|who have tasted the goodness of the word of God and the powers of the coming age,
HEB|6|6|if they fall away, to be brought back to repentance, because to their loss they are crucifying the Son of God all over again and subjecting him to public disgrace.
HEB|6|7|Land that drinks in the rain often falling on it and that produces a crop useful to those for whom it is farmed receives the blessing of God.
HEB|6|8|But land that produces thorns and thistles is worthless and is in danger of being cursed. In the end it will be burned.
HEB|6|9|Even though we speak like this, dear friends, we are confident of better things in your case--things that accompany salvation.
HEB|6|10|God is not unjust; he will not forget your work and the love you have shown him as you have helped his people and continue to help them.
HEB|6|11|We want each of you to show this same diligence to the very end, in order to make your hope sure.
HEB|6|12|We do not want you to become lazy, but to imitate those who through faith and patience inherit what has been promised.
HEB|6|13|When God made his promise to Abraham, since there was no one greater for him to swear by, he swore by himself,
HEB|6|14|saying, "I will surely bless you and give you many descendants."
HEB|6|15|And so after waiting patiently, Abraham received what was promised.
HEB|6|16|Men swear by someone greater than themselves, and the oath confirms what is said and puts an end to all argument.
HEB|6|17|Because God wanted to make the unchanging nature of his purpose very clear to the heirs of what was promised, he confirmed it with an oath.
HEB|6|18|God did this so that, by two unchangeable things in which it is impossible for God to lie, we who have fled to take hold of the hope offered to us may be greatly encouraged.
HEB|6|19|We have this hope as an anchor for the soul, firm and secure. It enters the inner sanctuary behind the curtain,
HEB|6|20|where Jesus, who went before us, has entered on our behalf. He has become a high priest forever, in the order of Melchizedek.
HEB|7|1|This Melchizedek was king of Salem and priest of God Most High. He met Abraham returning from the defeat of the kings and blessed him,
HEB|7|2|and Abraham gave him a tenth of everything. First, his name means "king of righteousness"; then also, "king of Salem" means "king of peace."
HEB|7|3|Without father or mother, without genealogy, without beginning of days or end of life, like the Son of God he remains a priest forever.
HEB|7|4|Just think how great he was: Even the patriarch Abraham gave him a tenth of the plunder!
HEB|7|5|Now the law requires the descendants of Levi who become priests to collect a tenth from the people--that is, their brothers--even though their brothers are descended from Abraham.
HEB|7|6|This man, however, did not trace his descent from Levi, yet he collected a tenth from Abraham and blessed him who had the promises.
HEB|7|7|And without doubt the lesser person is blessed by the greater.
HEB|7|8|In the one case, the tenth is collected by men who die; but in the other case, by him who is declared to be living.
HEB|7|9|One might even say that Levi, who collects the tenth, paid the tenth through Abraham,
HEB|7|10|because when Melchizedek met Abraham, Levi was still in the body of his ancestor.
HEB|7|11|If perfection could have been attained through the Levitical priesthood (for on the basis of it the law was given to the people), why was there still need for another priest to come--one in the order of Melchizedek, not in the order of Aaron?
HEB|7|12|For when there is a change of the priesthood, there must also be a change of the law.
HEB|7|13|He of whom these things are said belonged to a different tribe, and no one from that tribe has ever served at the altar.
HEB|7|14|For it is clear that our Lord descended from Judah, and in regard to that tribe Moses said nothing about priests.
HEB|7|15|And what we have said is even more clear if another priest like Melchizedek appears,
HEB|7|16|one who has become a priest not on the basis of a regulation as to his ancestry but on the basis of the power of an indestructible life.
HEB|7|17|For it is declared: "You are a priest forever, in the order of Melchizedek."
HEB|7|18|The former regulation is set aside because it was weak and useless
HEB|7|19|(for the law made nothing perfect), and a better hope is introduced, by which we draw near to God.
HEB|7|20|And it was not without an oath! Others became priests without any oath,
HEB|7|21|but he became a priest with an oath when God said to him: "The Lord has sworn and will not change his mind: 'You are a priest forever.'"
HEB|7|22|Because of this oath, Jesus has become the guarantee of a better covenant.
HEB|7|23|Now there have been many of those priests, since death prevented them from continuing in office;
HEB|7|24|but because Jesus lives forever, he has a permanent priesthood.
HEB|7|25|Therefore he is able to save completely those who come to God through him, because he always lives to intercede for them.
HEB|7|26|Such a high priest meets our need--one who is holy, blameless, pure, set apart from sinners, exalted above the heavens.
HEB|7|27|Unlike the other high priests, he does not need to offer sacrifices day after day, first for his own sins, and then for the sins of the people. He sacrificed for their sins once for all when he offered himself.
HEB|7|28|For the law appoints as high priests men who are weak; but the oath, which came after the law, appointed the Son, who has been made perfect forever.
HEB|8|1|The point of what we are saying is this: We do have such a high priest, who sat down at the right hand of the throne of the Majesty in heaven,
HEB|8|2|and who serves in the sanctuary, the true tabernacle set up by the Lord, not by man.
HEB|8|3|Every high priest is appointed to offer both gifts and sacrifices, and so it was necessary for this one also to have something to offer.
HEB|8|4|If he were on earth, he would not be a priest, for there are already men who offer the gifts prescribed by the law.
HEB|8|5|They serve at a sanctuary that is a copy and shadow of what is in heaven. This is why Moses was warned when he was about to build the tabernacle: "See to it that you make everything according to the pattern shown you on the mountain."
HEB|8|6|But the ministry Jesus has received is as superior to theirs as the covenant of which he is mediator is superior to the old one, and it is founded on better promises.
HEB|8|7|For if there had been nothing wrong with that first covenant, no place would have been sought for another.
HEB|8|8|But God found fault with the people and said: "The time is coming, declares the Lord, when I will make a new covenant with the house of Israel and with the house of Judah.
HEB|8|9|It will not be like the covenant I made with their forefathers when I took them by the hand to lead them out of Egypt, because they did not remain faithful to my covenant, and I turned away from them, declares the Lord.
HEB|8|10|This is the covenant I will make with the house of Israel after that time, declares the Lord. I will put my laws in their minds and write them on their hearts. I will be their God, and they will be my people.
HEB|8|11|No longer will a man teach his neighbor, or a man his brother, saying, 'Know the Lord,' because they will all know me, from the least of them to the greatest.
HEB|8|12|For I will forgive their wickedness and will remember their sins no more."
HEB|8|13|By calling this covenant "new," he has made the first one obsolete; and what is obsolete and aging will soon disappear.
HEB|9|1|Now the first covenant had regulations for worship and also an earthly sanctuary.
HEB|9|2|A tabernacle was set up. In its first room were the lampstand, the table and the consecrated bread; this was called the Holy Place.
HEB|9|3|Behind the second curtain was a room called the Most Holy Place,
HEB|9|4|which had the golden altar of incense and the gold-covered ark of the covenant. This ark contained the gold jar of manna, Aaron's staff that had budded, and the stone tablets of the covenant.
HEB|9|5|Above the ark were the cherubim of the Glory, overshadowing the atonement cover. But we cannot discuss these things in detail now.
HEB|9|6|When everything had been arranged like this, the priests entered regularly into the outer room to carry on their ministry.
HEB|9|7|But only the high priest entered the inner room, and that only once a year, and never without blood, which he offered for himself and for the sins the people had committed in ignorance.
HEB|9|8|The Holy Spirit was showing by this that the way into the Most Holy Place had not yet been disclosed as long as the first tabernacle was still standing.
HEB|9|9|This is an illustration for the present time, indicating that the gifts and sacrifices being offered were not able to clear the conscience of the worshiper.
HEB|9|10|They are only a matter of food and drink and various ceremonial washings--external regulations applying until the time of the new order.
HEB|9|11|When Christ came as high priest of the good things that are already here, he went through the greater and more perfect tabernacle that is not man-made, that is to say, not a part of this creation.
HEB|9|12|He did not enter by means of the blood of goats and calves; but he entered the Most Holy Place once for all by his own blood, having obtained eternal redemption.
HEB|9|13|The blood of goats and bulls and the ashes of a heifer sprinkled on those who are ceremonially unclean sanctify them so that they are outwardly clean.
HEB|9|14|How much more, then, will the blood of Christ, who through the eternal Spirit offered himself unblemished to God, cleanse our consciences from acts that lead to death, so that we may serve the living God!
HEB|9|15|For this reason Christ is the mediator of a new covenant, that those who are called may receive the promised eternal inheritance--now that he has died as a ransom to set them free from the sins committed under the first covenant.
HEB|9|16|In the case of a will, it is necessary to prove the death of the one who made it,
HEB|9|17|because a will is in force only when somebody has died; it never takes effect while the one who made it is living.
HEB|9|18|This is why even the first covenant was not put into effect without blood.
HEB|9|19|When Moses had proclaimed every commandment of the law to all the people, he took the blood of calves, together with water, scarlet wool and branches of hyssop, and sprinkled the scroll and all the people.
HEB|9|20|He said, "This is the blood of the covenant, which God has commanded you to keep."
HEB|9|21|In the same way, he sprinkled with the blood both the tabernacle and everything used in its ceremonies.
HEB|9|22|In fact, the law requires that nearly everything be cleansed with blood, and without the shedding of blood there is no forgiveness.
HEB|9|23|It was necessary, then, for the copies of the heavenly things to be purified with these sacrifices, but the heavenly things themselves with better sacrifices than these.
HEB|9|24|For Christ did not enter a man-made sanctuary that was only a copy of the true one; he entered heaven itself, now to appear for us in God's presence.
HEB|9|25|Nor did he enter heaven to offer himself again and again, the way the high priest enters the Most Holy Place every year with blood that is not his own.
HEB|9|26|Then Christ would have had to suffer many times since the creation of the world. But now he has appeared once for all at the end of the ages to do away with sin by the sacrifice of himself.
HEB|9|27|Just as man is destined to die once, and after that to face judgment,
HEB|9|28|so Christ was sacrificed once to take away the sins of many people; and he will appear a second time, not to bear sin, but to bring salvation to those who are waiting for him.
HEB|10|1|The law is only a shadow of the good things that are coming--not the realities themselves. For this reason it can never, by the same sacrifices repeated endlessly year after year, make perfect those who draw near to worship.
HEB|10|2|If it could, would they not have stopped being offered? For the worshipers would have been cleansed once for all, and would no longer have felt guilty for their sins.
HEB|10|3|But those sacrifices are an annual reminder of sins,
HEB|10|4|because it is impossible for the blood of bulls and goats to take away sins.
HEB|10|5|Therefore, when Christ came into the world, he said: "Sacrifice and offering you did not desire, but a body you prepared for me;
HEB|10|6|with burnt offerings and sin offerings you were not pleased.
HEB|10|7|Then I said, 'Here I am--it is written about me in the scroll--I have come to do your will, O God.'"
HEB|10|8|First he said, "Sacrifices and offerings, burnt offerings and sin offerings you did not desire, nor were you pleased with them" (although the law required them to be made).
HEB|10|9|Then he said, "Here I am, I have come to do your will." He sets aside the first to establish the second.
HEB|10|10|And by that will, we have been made holy through the sacrifice of the body of Jesus Christ once for all.
HEB|10|11|Day after day every priest stands and performs his religious duties; again and again he offers the same sacrifices, which can never take away sins.
HEB|10|12|But when this priest had offered for all time one sacrifice for sins, he sat down at the right hand of God.
HEB|10|13|Since that time he waits for his enemies to be made his footstool,
HEB|10|14|because by one sacrifice he has made perfect forever those who are being made holy.
HEB|10|15|The Holy Spirit also testifies to us about this. First he says:
HEB|10|16|"This is the covenant I will make with them after that time, says the Lord. I will put my laws in their hearts, and I will write them on their minds."
HEB|10|17|Then he adds: "Their sins and lawless acts I will remember no more."
HEB|10|18|And where these have been forgiven, there is no longer any sacrifice for sin.
HEB|10|19|Therefore, brothers, since we have confidence to enter the Most Holy Place by the blood of Jesus,
HEB|10|20|by a new and living way opened for us through the curtain, that is, his body,
HEB|10|21|and since we have a great priest over the house of God,
HEB|10|22|let us draw near to God with a sincere heart in full assurance of faith, having our hearts sprinkled to cleanse us from a guilty conscience and having our bodies washed with pure water.
HEB|10|23|Let us hold unswervingly to the hope we profess, for he who promised is faithful.
HEB|10|24|And let us consider how we may spur one another on toward love and good deeds.
HEB|10|25|Let us not give up meeting together, as some are in the habit of doing, but let us encourage one another--and all the more as you see the Day approaching.
HEB|10|26|If we deliberately keep on sinning after we have received the knowledge of the truth, no sacrifice for sins is left,
HEB|10|27|but only a fearful expectation of judgment and of raging fire that will consume the enemies of God.
HEB|10|28|Anyone who rejected the law of Moses died without mercy on the testimony of two or three witnesses.
HEB|10|29|How much more severely do you think a man deserves to be punished who has trampled the Son of God under foot, who has treated as an unholy thing the blood of the covenant that sanctified him, and who has insulted the Spirit of grace?
HEB|10|30|For we know him who said, "It is mine to avenge; I will repay," and again, "The Lord will judge his people."
HEB|10|31|It is a dreadful thing to fall into the hands of the living God.
HEB|10|32|Remember those earlier days after you had received the light, when you stood your ground in a great contest in the face of suffering.
HEB|10|33|Sometimes you were publicly exposed to insult and persecution; at other times you stood side by side with those who were so treated.
HEB|10|34|You sympathized with those in prison and joyfully accepted the confiscation of your property, because you knew that you yourselves had better and lasting possessions.
HEB|10|35|So do not throw away your confidence; it will be richly rewarded.
HEB|10|36|You need to persevere so that when you have done the will of God, you will receive what he has promised.
HEB|10|37|For in just a very little while, "He who is coming will come and will not delay.
HEB|10|38|But my righteous one will live by faith. And if he shrinks back, I will not be pleased with him."
HEB|10|39|But we are not of those who shrink back and are destroyed, but of those who believe and are saved.
HEB|11|1|Now faith is being sure of what we hope for and certain of what we do not see.
HEB|11|2|This is what the ancients were commended for.
HEB|11|3|By faith we understand that the universe was formed at God's command, so that what is seen was not made out of what was visible.
HEB|11|4|By faith Abel offered God a better sacrifice than Cain did. By faith he was commended as a righteous man, when God spoke well of his offerings. And by faith he still speaks, even though he is dead.
HEB|11|5|By faith Enoch was taken from this life, so that he did not experience death; he could not be found, because God had taken him away. For before he was taken, he was commended as one who pleased God.
HEB|11|6|And without faith it is impossible to please God, because anyone who comes to him must believe that he exists and that he rewards those who earnestly seek him.
HEB|11|7|By faith Noah, when warned about things not yet seen, in holy fear built an ark to save his family. By his faith he condemned the world and became heir of the righteousness that comes by faith.
HEB|11|8|By faith Abraham, when called to go to a place he would later receive as his inheritance, obeyed and went, even though he did not know where he was going.
HEB|11|9|By faith he made his home in the promised land like a stranger in a foreign country; he lived in tents, as did Isaac and Jacob, who were heirs with him of the same promise.
HEB|11|10|For he was looking forward to the city with foundations, whose architect and builder is God.
HEB|11|11|By faith Abraham, even though he was past age--and Sarah herself was barren--was enabled to become a father because he considered him faithful who had made the promise.
HEB|11|12|And so from this one man, and he as good as dead, came descendants as numerous as the stars in the sky and as countless as the sand on the seashore.
HEB|11|13|All these people were still living by faith when they died. They did not receive the things promised; they only saw them and welcomed them from a distance. And they admitted that they were aliens and strangers on earth.
HEB|11|14|People who say such things show that they are looking for a country of their own.
HEB|11|15|If they had been thinking of the country they had left, they would have had opportunity to return.
HEB|11|16|Instead, they were longing for a better country--a heavenly one. Therefore God is not ashamed to be called their God, for he has prepared a city for them.
HEB|11|17|By faith Abraham, when God tested him, offered Isaac as a sacrifice. He who had received the promises was about to sacrifice his one and only son,
HEB|11|18|even though God had said to him, "It is through Isaac that your offspring will be reckoned."
HEB|11|19|Abraham reasoned that God could raise the dead, and figuratively speaking, he did receive Isaac back from death.
HEB|11|20|By faith Isaac blessed Jacob and Esau in regard to their future.
HEB|11|21|By faith Jacob, when he was dying, blessed each of Joseph's sons, and worshiped as he leaned on the top of his staff.
HEB|11|22|By faith Joseph, when his end was near, spoke about the exodus of the Israelites from Egypt and gave instructions about his bones.
HEB|11|23|By faith Moses' parents hid him for three months after he was born, because they saw he was no ordinary child, and they were not afraid of the king's edict.
HEB|11|24|By faith Moses, when he had grown up, refused to be known as the son of Pharaoh's daughter.
HEB|11|25|He chose to be mistreated along with the people of God rather than to enjoy the pleasures of sin for a short time.
HEB|11|26|He regarded disgrace for the sake of Christ as of greater value than the treasures of Egypt, because he was looking ahead to his reward.
HEB|11|27|By faith he left Egypt, not fearing the king's anger; he persevered because he saw him who is invisible.
HEB|11|28|By faith he kept the Passover and the sprinkling of blood, so that the destroyer of the firstborn would not touch the firstborn of Israel.
HEB|11|29|By faith the people passed through the Red Sea as on dry land; but when the Egyptians tried to do so, they were drowned.
HEB|11|30|By faith the walls of Jericho fell, after the people had marched around them for seven days.
HEB|11|31|By faith the prostitute Rahab, because she welcomed the spies, was not killed with those who were disobedient.
HEB|11|32|And what more shall I say? I do not have time to tell about Gideon, Barak, Samson, Jephthah, David, Samuel and the prophets,
HEB|11|33|who through faith conquered kingdoms, administered justice, and gained what was promised; who shut the mouths of lions,
HEB|11|34|quenched the fury of the flames, and escaped the edge of the sword; whose weakness was turned to strength; and who became powerful in battle and routed foreign armies.
HEB|11|35|Women received back their dead, raised to life again. Others were tortured and refused to be released, so that they might gain a better resurrection.
HEB|11|36|Some faced jeers and flogging, while still others were chained and put in prison.
HEB|11|37|They were stoned; they were sawed in two; they were put to death by the sword. They went about in sheepskins and goatskins, destitute, persecuted and mistreated--
HEB|11|38|the world was not worthy of them. They wandered in deserts and mountains, and in caves and holes in the ground.
HEB|11|39|These were all commended for their faith, yet none of them received what had been promised.
HEB|11|40|God had planned something better for us so that only together with us would they be made perfect.
HEB|12|1|Therefore, since we are surrounded by such a great cloud of witnesses, let us throw off everything that hinders and the sin that so easily entangles, and let us run with perseverance the race marked out for us.
HEB|12|2|Let us fix our eyes on Jesus, the author and perfecter of our faith, who for the joy set before him endured the cross, scorning its shame, and sat down at the right hand of the throne of God.
HEB|12|3|Consider him who endured such opposition from sinful men, so that you will not grow weary and lose heart.
HEB|12|4|In your struggle against sin, you have not yet resisted to the point of shedding your blood.
HEB|12|5|And you have forgotten that word of encouragement that addresses you as sons: "My son, do not make light of the Lord's discipline, and do not lose heart when he rebukes you,
HEB|12|6|because the Lord disciplines those he loves, and he punishes everyone he accepts as a son."
HEB|12|7|Endure hardship as discipline; God is treating you as sons. For what son is not disciplined by his father?
HEB|12|8|If you are not disciplined (and everyone undergoes discipline), then you are illegitimate children and not true sons.
HEB|12|9|Moreover, we have all had human fathers who disciplined us and we respected them for it. How much more should we submit to the Father of our spirits and live!
HEB|12|10|Our fathers disciplined us for a little while as they thought best; but God disciplines us for our good, that we may share in his holiness.
HEB|12|11|No discipline seems pleasant at the time, but painful. Later on, however, it produces a harvest of righteousness and peace for those who have been trained by it.
HEB|12|12|Therefore, strengthen your feeble arms and weak knees.
HEB|12|13|"Make level paths for your feet," so that the lame may not be disabled, but rather healed.
HEB|12|14|Make every effort to live in peace with all men and to be holy; without holiness no one will see the Lord.
HEB|12|15|See to it that no one misses the grace of God and that no bitter root grows up to cause trouble and defile many.
HEB|12|16|See that no one is sexually immoral, or is godless like Esau, who for a single meal sold his inheritance rights as the oldest son.
HEB|12|17|Afterward, as you know, when he wanted to inherit this blessing, he was rejected. He could bring about no change of mind, though he sought the blessing with tears.
HEB|12|18|You have not come to a mountain that can be touched and that is burning with fire; to darkness, gloom and storm;
HEB|12|19|to a trumpet blast or to such a voice speaking words that those who heard it begged that no further word be spoken to them,
HEB|12|20|because they could not bear what was commanded: "If even an animal touches the mountain, it must be stoned."
HEB|12|21|The sight was so terrifying that Moses said, "I am trembling with fear."
HEB|12|22|But you have come to Mount Zion, to the heavenly Jerusalem, the city of the living God. You have come to thousands upon thousands of angels in joyful assembly,
HEB|12|23|to the church of the firstborn, whose names are written in heaven. You have come to God, the judge of all men, to the spirits of righteous men made perfect,
HEB|12|24|to Jesus the mediator of a new covenant, and to the sprinkled blood that speaks a better word than the blood of Abel.
HEB|12|25|See to it that you do not refuse him who speaks. If they did not escape when they refused him who warned them on earth, how much less will we, if we turn away from him who warns us from heaven?
HEB|12|26|At that time his voice shook the earth, but now he has promised, "Once more I will shake not only the earth but also the heavens."
HEB|12|27|The words "once more" indicate the removing of what can be shaken--that is, created things--so that what cannot be shaken may remain.
HEB|12|28|Therefore, since we are receiving a kingdom that cannot be shaken, let us be thankful, and so worship God acceptably with reverence and awe,
HEB|12|29|for our "God is a consuming fire."
HEB|13|1|Keep on loving each other as brothers.
HEB|13|2|Do not forget to entertain strangers, for by so doing some people have entertained angels without knowing it.
HEB|13|3|Remember those in prison as if you were their fellow prisoners, and those who are mistreated as if you yourselves were suffering.
HEB|13|4|Marriage should be honored by all, and the marriage bed kept pure, for God will judge the adulterer and all the sexually immoral.
HEB|13|5|Keep your lives free from the love of money and be content with what you have, because God has said, "Never will I leave you; never will I forsake you."
HEB|13|6|So we say with confidence, "The Lord is my helper; I will not be afraid. What can man do to me?"
HEB|13|7|Remember your leaders, who spoke the word of God to you. Consider the outcome of their way of life and imitate their faith.
HEB|13|8|Jesus Christ is the same yesterday and today and forever.
HEB|13|9|Do not be carried away by all kinds of strange teachings. It is good for our hearts to be strengthened by grace, not by ceremonial foods, which are of no value to those who eat them.
HEB|13|10|We have an altar from which those who minister at the tabernacle have no right to eat.
HEB|13|11|The high priest carries the blood of animals into the Most Holy Place as a sin offering, but the bodies are burned outside the camp.
HEB|13|12|And so Jesus also suffered outside the city gate to make the people holy through his own blood.
HEB|13|13|Let us, then, go to him outside the camp, bearing the disgrace he bore.
HEB|13|14|For here we do not have an enduring city, but we are looking for the city that is to come.
HEB|13|15|Through Jesus, therefore, let us continually offer to God a sacrifice of praise--the fruit of lips that confess his name.
HEB|13|16|And do not forget to do good and to share with others, for with such sacrifices God is pleased.
HEB|13|17|Obey your leaders and submit to their authority. They keep watch over you as men who must give an account. Obey them so that their work will be a joy, not a burden, for that would be of no advantage to you.
HEB|13|18|Pray for us. We are sure that we have a clear conscience and desire to live honorably in every way.
HEB|13|19|I particularly urge you to pray so that I may be restored to you soon.
HEB|13|20|May the God of peace, who through the blood of the eternal covenant brought back from the dead our Lord Jesus, that great Shepherd of the sheep,
HEB|13|21|equip you with everything good for doing his will, and may he work in us what is pleasing to him, through Jesus Christ, to whom be glory for ever and ever. Amen.
HEB|13|22|Brothers, I urge you to bear with my word of exhortation, for I have written you only a short letter.
HEB|13|23|I want you to know that our brother Timothy has been released. If he arrives soon, I will come with him to see you.
HEB|13|24|Greet all your leaders and all God's people. Those from Italy send you their greetings.
HEB|13|25|Grace be with you all.
