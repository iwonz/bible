JOEL|1|1|The word of the LORD that came to Joel, the son of Pethuel:
JOEL|1|2|Hear this, you elders; give ear, all inhabitants of the land! Has such a thing happened in your days, or in the days of your fathers?
JOEL|1|3|Tell your children of it, and let your children tell their children, and their children to another generation.
JOEL|1|4|What the cutting locust left, the swarming locust has eaten. What the swarming locust left, the hopping locust has eaten, and what the hopping locust left, the destroying locust has eaten.
JOEL|1|5|Awake, you drunkards, and weep, and wail, all you drinkers of wine, because of the sweet wine, for it is cut off from your mouth.
JOEL|1|6|For a nation has come up against my land, powerful and beyond number; its teeth are lions' teeth, and it has the fangs of a lioness.
JOEL|1|7|It has laid waste my vine and splintered my fig tree; it has stripped off their bark and thrown it down; their branches are made white.
JOEL|1|8|Lament like a virgin wearing sackcloth for the bridegroom of her youth.
JOEL|1|9|The grain offering and the drink offering are cut off from the house of the LORD. The priests mourn, the ministers of the LORD.
JOEL|1|10|The fields are destroyed, the ground mourns, because the grain is destroyed, the wine dries up, the oil languishes.
JOEL|1|11|Be ashamed, O tillers of the soil; wail, O vinedressers, for the wheat and the barley, because the harvest of the field has perished.
JOEL|1|12|The vine dries up; the fig tree languishes. Pomegranate, palm, and apple, all the trees of the field are dried up, and gladness dries up from the children of man.
JOEL|1|13|Put on sackcloth and lament, O priests; wail, O ministers of the altar. Go in, pass the night in sackcloth, O ministers of my God! Because grain offering and drink offering are withheld from the house of your God.
JOEL|1|14|Consecrate a fast; call a solemn assembly. Gather the elders and all the inhabitants of the land to the house of the LORD your God, and cry out to the LORD.
JOEL|1|15|Alas for the day! For the day of the LORD is near, and as destruction from the Almighty it comes.
JOEL|1|16|Is not the food cut off before our eyes, joy and gladness from the house of our God?
JOEL|1|17|The seed shrivels under the clods; the storehouses are desolate; the granaries are torn down because the grain has dried up.
JOEL|1|18|How the beasts groan! The herds of cattle are perplexed because there is no pasture for them; even the flocks of sheep suffer.
JOEL|1|19|To you, O LORD, I call. For fire has devoured the pastures of the wilderness, and flame has burned all the trees of the field.
JOEL|1|20|Even the beasts of the field pant for you because the water brooks are dried up, and fire has devoured the pastures of the wilderness.
JOEL|2|1|Blow a trumpet in Zion;sound an alarm on my holy mountain! Let all the inhabitants of the land tremble, for the day of the LORD is coming; it is near,
JOEL|2|2|a day of darkness and gloom, a day of clouds and thick darkness! Like blackness there is spread upon the mountains a great and powerful people; their like has never been before, nor will be again after them through the years of all generations.
JOEL|2|3|Fire devours before them, and behind them a flame burns. The land is like the garden of Eden before them, but behind them a desolate wilderness, and nothing escapes them.
JOEL|2|4|Their appearance is like the appearance of horses, and like war horses they run.
JOEL|2|5|As with the rumbling of chariots, they leap on the tops of the mountains, like the crackling of a flame of fire devouring the stubble, like a powerful army drawn up for battle.
JOEL|2|6|Before them peoples are in anguish; all faces grow pale.
JOEL|2|7|Like warriors they charge; like soldiers they scale the wall. They march each on his way; they do not swerve from their paths.
JOEL|2|8|They do not jostle one another; each marches in his path; they burst through the weapons and are not halted.
JOEL|2|9|They leap upon the city, they run upon the walls, they climb up into the houses, they enter through the windows like a thief.
JOEL|2|10|The earth quakes before them; the heavens tremble. The sun and the moon are darkened, and the stars withdraw their shining.
JOEL|2|11|The LORD utters his voice before his army, for his camp is exceedingly great; he who executes his word is powerful. For the day of the LORD is great and very awesome; who can endure it?
JOEL|2|12|"Yet even now," declares the LORD, "return to me with all your heart, with fasting, with weeping, and with mourning;
JOEL|2|13|and rend your hearts and not your garments." Return to the LORD, your God, for he is gracious and merciful, slow to anger, and abounding in steadfast love; and he relents over disaster.
JOEL|2|14|Who knows whether he will not turn and relent, and leave a blessing behind him, a grain offering and a drink offering for the LORD your God?
JOEL|2|15|Blow the trumpet in Zion; consecrate a fast; call a solemn assembly;
JOEL|2|16|gather the people. Consecrate the congregation; assemble the elders; gather the children, even nursing infants. Let the bridegroom leave his room, and the bride her chamber.
JOEL|2|17|Between the vestibule and the altar let the priests, the ministers of the LORD, weep and say, "Spare your people, O LORD, and make not your heritage a reproach, a byword among the nations. Why should they say among the peoples, 'Where is their God?'"
JOEL|2|18|Then the LORD became jealous for his land and had pity on his people.
JOEL|2|19|The LORD answered and said to his people, "Behold, I am sending to you grain, wine, and oil, and you will be satisfied; and I will no more make you a reproach among the nations.
JOEL|2|20|"I will remove the northerner far from you, and drive him into a parched and desolate land, his vanguard into the eastern sea, and his rear guard into the western sea; the stench and foul smell of him will rise, for he has done great things.
JOEL|2|21|"Fear not, O land; be glad and rejoice, for the LORD has done great things!
JOEL|2|22|Fear not, you beasts of the field, for the pastures of the wilderness are green; the tree bears its fruit; the fig tree and vine give their full yield.
JOEL|2|23|"Be glad, O children of Zion, and rejoice in the LORD your God, for he has given the early rain for your vindication; he has poured down for you abundant rain, the early and the latter rain, as before.
JOEL|2|24|"The threshing floors shall be full of grain; the vats shall overflow with wine and oil.
JOEL|2|25|I will restore to you the years that the swarming locust has eaten, the hopper, the destroyer, and the cutter, my great army, which I sent among you.
JOEL|2|26|"You shall eat in plenty and be satisfied, and praise the name of the LORD your God, who has dealt wondrously with you. And my people shall never again be put to shame.
JOEL|2|27|You shall know that I am in the midst of Israel, and that I am the LORD your God and there is none else. And my people shall never again be put to shame.
JOEL|2|28|"And it shall come to pass afterward, that I will pour out my Spirit on all flesh; your sons and your daughters shall prophesy, your old men shall dream dreams, and your young men shall see visions.
JOEL|2|29|Even on the male and female servants in those days I will pour out my Spirit.
JOEL|2|30|"And I will show wonders in the heavens and on the earth, blood and fire and columns of smoke.
JOEL|2|31|The sun shall be turned to darkness, and the moon to blood, before the great and awesome day of the LORD comes.
JOEL|2|32|And it shall come to pass that everyone who calls on the name of the LORD shall be saved. For in Mount Zion and in Jerusalem there shall be those who escape, as the LORD has said, and among the survivors shall be those whom the LORD calls.
JOEL|3|1|"For behold, in those days and at that time, when I restore the fortunes of Judah and Jerusalem,
JOEL|3|2|I will gather all the nations and bring them down to the Valley of Jehoshaphat. And I will enter into judgment with them there, on behalf of my people and my heritage Israel, because they have scattered them among the nations and have divided up my land,
JOEL|3|3|and have cast lots for my people, and have traded a boy for a prostitute, and have sold a girl for wine and have drunk it.
JOEL|3|4|"What are you to me, O Tyre and Sidon, and all the regions of Philistia? Are you paying me back for something? If you are paying me back, I will return your payment on your own head swiftly and speedily.
JOEL|3|5|For you have taken my silver and my gold, and have carried my rich treasures into your temples.
JOEL|3|6|You have sold the people of Judah and Jerusalem to the Greeks in order to remove them far from their own border.
JOEL|3|7|Behold, I will stir them up from the place to which you have sold them, and I will return your payment on your own head.
JOEL|3|8|I will sell your sons and your daughters into the hand of the people of Judah, and they will sell them to the Sabeans, to a nation far away, for the LORD has spoken."
JOEL|3|9|Proclaim this among the nations: Consecrate for war; stir up the mighty men. Let all the men of war draw near; let them come up.
JOEL|3|10|Beat your plowshares into swords, and your pruning hooks into spears; let the weak say, "I am a warrior."
JOEL|3|11|Hasten and come, all you surrounding nations, and gather yourselves there. Bring down your warriors, O LORD.
JOEL|3|12|Let the nations stir themselves up and come up to the Valley of Jehoshaphat; for there I will sit to judge all the surrounding nations.
JOEL|3|13|Put in the sickle, for the harvest is ripe. Go in, tread, for the winepress is full. The vats overflow, for their evil is great.
JOEL|3|14|Multitudes, multitudes, in the valley of decision! For the day of the LORD is near in the valley of decision.
JOEL|3|15|The sun and the moon are darkened, and the stars withdraw their shining.
JOEL|3|16|The LORD roars from Zion, and utters his voice from Jerusalem, and the heavens and the earth quake. But the LORD is a refuge to his people, a stronghold to the people of Israel.
JOEL|3|17|"So you shall know that I am the LORD your God, who dwell in Zion, my holy mountain. And Jerusalem shall be holy, and strangers shall never again pass through it.
JOEL|3|18|"And in that day the mountains shall drip sweet wine, and the hills shall flow with milk, and all the streambeds of Judah shall flow with water; and a fountain shall come forth from the house of the LORD and water the Valley of Shittim.
JOEL|3|19|"Egypt shall become a desolation and Edom a desolate wilderness, for the violence done to the people of Judah, because they have shed innocent blood in their land.
JOEL|3|20|But Judah shall be inhabited forever, and Jerusalem to all generations.
JOEL|3|21|I will avenge their blood, blood I have not avenged, for the LORD dwells in Zion."
