PROV|1|1|大衛 的兒子， 以色列 王 所羅門 的箴言：
PROV|1|2|要使人懂得智慧和訓誨， 明白通達的言語，
PROV|1|3|使人領受明智的訓誨， 就是公義、公平和正直，
PROV|1|4|使愚蒙人靈巧， 使年輕人有知識，有智謀。
PROV|1|5|智慧人聽見，增長學問， 聰明人得著智謀，
PROV|1|6|明白箴言和譬喻， 懂得智慧人的言詞和謎語。
PROV|1|7|敬畏耶和華是知識的開端； 愚妄人藐視智慧和訓誨。
PROV|1|8|我兒啊，要聽你父親的訓誨， 不可離棄你母親的教誨；
PROV|1|9|因為這要作你頭上恩惠的華冠， 作你頸上的項鏈。
PROV|1|10|我兒啊，罪人若引誘你， 你不可隨從。
PROV|1|11|他們若說：「你與我們同去， 我們要埋伏殺人流血， 無故地潛藏，殺害無辜；
PROV|1|12|我們好像陰間，把他們活活吞下， 囫圇吞下，如吞下那下到地府的人；
PROV|1|13|我們必得各樣寶物， 將所奪來的裝滿房屋；
PROV|1|14|你來與我們同夥， 共用一個錢囊。」
PROV|1|15|我兒啊，不要與他們走同一道路， 禁止你的腳走他們的路徑。
PROV|1|16|因為他們的腳奔跑行惡， 他們急速殺人流血。
PROV|1|17|在飛鳥眼前張設網羅， 一定會徒勞無功；
PROV|1|18|同樣，他們埋伏，是自流己血， 他們潛藏，是自害己命。
PROV|1|19|凡靠暴力歛財的，所行之路都是如此， 這種念頭必奪去自己的生命。
PROV|1|20|智慧 在街市上呼喊， 在廣場上高聲吶喊，
PROV|1|21|在熱鬧街頭呼叫， 在城門口，在城中，發出言語，說：
PROV|1|22|「你們無知的人喜愛無知， 傲慢人喜歡傲慢， 愚昧人恨惡知識， 要到幾時呢？
PROV|1|23|你們當因我的責備回轉， 我要將我的靈澆灌你們， 將我的話指示你們。
PROV|1|24|因為我呼喚，你們不聽， 我招手，無人理會。
PROV|1|25|你們忽視我一切的勸戒， 拒聽我的責備。
PROV|1|26|你們遭難，我就發笑； 驚恐臨到你們， 驚恐如狂風來臨， 災難好像暴風來到， 急難痛苦臨到你們身上， 我必嗤笑。
PROV|1|27|
PROV|1|28|那時，他們就會呼求我，我卻不回答， 懇切尋求我，卻尋不見。
PROV|1|29|因為他們恨惡知識， 選擇不敬畏耶和華，
PROV|1|30|不聽我的勸戒， 藐視我一切的責備，
PROV|1|31|所以他們要自食其果， 飽脹在自己的計謀中。
PROV|1|32|愚蒙人背道，害死自己， 愚昧人安逸，自取滅亡。
PROV|1|33|惟聽從我的，必安然居住， 得享寧靜，不怕災禍。」
PROV|2|1|我兒啊，你若領受我的言語， 珍藏我的命令，
PROV|2|2|留心聽智慧， 專心求聰明；
PROV|2|3|你若呼求明理， 揚聲求聰明，
PROV|2|4|尋找她，如尋找銀子， 搜尋她，如搜尋寶藏，
PROV|2|5|你就懂得敬畏耶和華， 得以認識上帝。
PROV|2|6|因為耶和華賞賜智慧， 知識和聰明都由他口而出。
PROV|2|7|他為正直人珍藏健全的知識， 給行為純正的人作盾牌，
PROV|2|8|為要保護公正的路， 庇護虔誠人的道。
PROV|2|9|那時，你就明白公義、公平、 正直，和一切完善的道路。
PROV|2|10|因為智慧要進入你的心， 知識要使你內心歡愉。
PROV|2|11|智謀要庇護你， 聰明必保護你，
PROV|2|12|救你脫離惡人的道， 脫離言談乖謬的人。
PROV|2|13|他們離棄正直的路， 行走黑暗的道，
PROV|2|14|喜歡作惡， 喜愛惡人的錯謬。
PROV|2|15|他們的路歪曲， 他們偏離中道。
PROV|2|16|智慧要救你遠離陌生女子， 遠離那油嘴滑舌的外邦女子。
PROV|2|17|她離棄年輕時的配偶， 忘了自己神聖的盟約。
PROV|2|18|她的家陷入死亡， 她的路偏向陰魂。
PROV|2|19|凡到她那裏去的，不得回轉， 也得不到生命的路。
PROV|2|20|智慧使你行善人的道， 守義人的路。
PROV|2|21|正直人必在地上居住， 完全人必在其上存留；
PROV|2|22|惟惡人要從地上剪除， 奸詐人要被拔出。
PROV|3|1|我兒啊，不要忘記我的教誨， 你的心要謹守我的命令，
PROV|3|2|因為它們 必加給你長久的日子， 生命的年數與平安。
PROV|3|3|不可使慈愛和誠信離開你， 要繫在你頸項上，刻在你心版上。
PROV|3|4|這樣，你必在上帝和世人眼前 蒙恩惠，有美好的見識。
PROV|3|5|你要專心仰賴耶和華， 不可倚靠自己的聰明，
PROV|3|6|在你一切所行的路上都要認定他， 他必使你的道路平直。
PROV|3|7|不要自以為有智慧； 要敬畏耶和華，遠離惡事。
PROV|3|8|這便醫治你的肉體 ， 滋潤你的百骨。
PROV|3|9|你要以財物 和一切初熟的土產尊崇耶和華，
PROV|3|10|這樣，你的倉庫必充滿有餘， 你的酒池有新酒盈溢。
PROV|3|11|我兒啊，不可輕看耶和華的管教， 也不可厭煩他的責備，
PROV|3|12|因為耶和華所愛的，他必責備， 正如父親責備所喜愛的兒子。
PROV|3|13|得智慧，得聰明的， 這人有福了。
PROV|3|14|因為智慧的獲利勝過銀子， 所得的盈餘強如金子，
PROV|3|15|比寶石 更寶貴， 你一切所喜愛的，都不足與其比較。
PROV|3|16|她的右手有長壽， 左手有富貴。
PROV|3|17|她的道是安樂， 她的路全是平安。
PROV|3|18|她給持守她的人作生命樹， 謹守她的必定蒙福。
PROV|3|19|耶和華以智慧奠立地基， 以聰明鋪設諸天，
PROV|3|20|以知識使深淵裂開， 使天空滴下甘露。
PROV|3|21|我兒啊，要謹守健全的知識和智謀， 不可使它們偏離你的眼目。
PROV|3|22|這樣，它們必使你的生命有活力， 又作你頸項的美飾。
PROV|3|23|那時，你就坦然行路， 不致跌倒。
PROV|3|24|你躺下，必不懼怕； 你躺臥，睡得香甜。
PROV|3|25|忽然來的驚恐，你不要害怕； 惡人遭毀滅，也不要恐懼，
PROV|3|26|因為耶和華是你的倚靠， 他必保護你的腳不陷入羅網。
PROV|3|27|你的手若有行善的力量， 不可推辭，要施與那應得的人。
PROV|3|28|你若手頭方便， 不可對鄰舍說： 「去吧，明天再來，我必給你。」
PROV|3|29|你的鄰舍既在你附近安居， 不可設計害他。
PROV|3|30|人若未曾加害你， 不可無故與他相爭。
PROV|3|31|不可嫉妒殘暴的人， 不可選擇他的任何道路。
PROV|3|32|因為走偏方向的人是耶和華所憎惡的； 正直人為他所親密。
PROV|3|33|耶和華詛咒惡人的家； 義人的居所他卻賜福。
PROV|3|34|他譏誚那愛譏誚的人； 但賜恩給謙卑的人。
PROV|3|35|智慧人必承受尊榮； 愚昧人高升卻是羞辱。
PROV|4|1|孩子們，要聽父親的訓誨， 留心明白道理。
PROV|4|2|因我給你們好的教導， 不可離棄我的教誨。
PROV|4|3|當我在父親面前還是小孩， 是母親獨一嬌兒的時候，
PROV|4|4|他教導我說：「你的心要持守我的話， 遵守我的命令，你就會存活。
PROV|4|5|要獲得智慧，要獲得聰明， 不可忘記， 也不可偏離我口中的言語。
PROV|4|6|不可離棄智慧，智慧就庇護你， 要愛她，她就保護你。
PROV|4|7|智慧為首，所以要獲得智慧， 要用你一切所有的換取聰明。
PROV|4|8|高舉智慧，她就使你升高， 擁抱智慧，她就使你尊榮。
PROV|4|9|她必將恩惠的華冠加在你頭上， 把榮冕賜給你。」
PROV|4|10|我兒啊，要聽，要領受我的言語， 你就必延年益壽。
PROV|4|11|我已指教你走智慧的道， 引導你行正直的路。
PROV|4|12|你行走，腳步沒有阻礙； 你奔跑，也不致跌倒。
PROV|4|13|要持定訓誨，不可放鬆； 要謹守它，因為它是你的生命。
PROV|4|14|不可行惡人的路， 不要走壞人的道；
PROV|4|15|要躲避，不可經過， 要轉離而去。
PROV|4|16|他們若不行惡，難以成眠， 不使人跌倒，就睡臥不安；
PROV|4|17|因為他們以邪惡當餅吃， 以暴力當酒喝。
PROV|4|18|但義人的路好像黎明的光， 越照越明，直到正午。
PROV|4|19|惡人的道幽暗， 自己不知因何跌倒。
PROV|4|20|我兒啊，要留心聽我的話， 側耳聽我的言語，
PROV|4|21|不可使它們偏離你的眼目， 要存記在你心中。
PROV|4|22|因為找到它們的，就找到生命， 得到全身的醫治。
PROV|4|23|你要保守你心，勝過保守一切， 因為生命的泉源由心發出。
PROV|4|24|要離開歪曲的口， 轉離偏邪的嘴唇。
PROV|4|25|你的兩眼要向前看， 你的雙目 直視前方。
PROV|4|26|要修平 你腳下的路， 你一切的道就必穩固。
PROV|4|27|不可偏左偏右， 你的腳要離開邪惡。
PROV|5|1|我兒啊，要留心聽我的智慧， 側耳聽我的聰明，
PROV|5|2|為要使你謹守智謀， 嘴唇保護知識。
PROV|5|3|因為陌生女子的嘴唇滴下蜂蜜， 她的口比油更滑，
PROV|5|4|後來卻苦似茵蔯， 銳利如兩刃的劍。
PROV|5|5|她的腳墜落死亡， 她的腳步踏入陰間，
PROV|5|6|她無法找到生命的道路， 她的路變遷不定，自己卻不知道。
PROV|5|7|孩子們，現在要聽從我， 不可離棄我口中的言語。
PROV|5|8|你所行的道要遠離她， 不可靠近她家的門口，
PROV|5|9|免得將你的尊榮給別人， 將你的歲月給殘忍的人；
PROV|5|10|免得陌生人滿得你的財富， 你勞苦所得的歸入外邦人的家。
PROV|5|11|在你人生終結，你皮肉和身體衰殘時， 你必唉聲嘆氣，
PROV|5|12|說：「我為何恨惡管教， 心裏輕看責備呢？
PROV|5|13|我不聽從教師的話， 也沒有側耳聽那教導我的。
PROV|5|14|在聚集的會眾中， 我幾乎墜入深淵。」
PROV|5|15|你要喝自己池中的水， 飲自己井裏的活水。
PROV|5|16|你的泉源豈可溢流在外？ 你的河水豈可流到街上？
PROV|5|17|讓它們惟獨歸你， 不可與陌生人同享。
PROV|5|18|要使你的泉源蒙福， 要喜愛你年輕時的妻子。
PROV|5|19|她如可愛的母鹿，如優美的母羊， 願她的胸懷使你時時滿足， 願你常常迷戀她的愛情。
PROV|5|20|我兒啊，你為何迷戀陌生女子？ 為何擁抱外邦女子的胸懷？
PROV|5|21|因為人所行的道都在耶和華眼前， 他察驗 人一切的路。
PROV|5|22|惡人被自己的罪孽抓住， 被自己罪惡的繩索纏繞。
PROV|5|23|他因不受管教而死亡， 因極度愚昧而走迷。
PROV|6|1|我兒啊，你若為朋友擔保， 替陌生人擊掌，
PROV|6|2|你就被口中的言語套住， 被嘴裏的言語抓住。
PROV|6|3|我兒啊，你既落在朋友手中，當這樣行才可救自己： 你要謙卑自己，去懇求你的朋友。
PROV|6|4|不要讓你的眼睛睡覺， 不可容你的眼皮打盹。
PROV|6|5|要救自己，如羚羊脫離獵人的手， 如鳥脫離捕鳥人的手。
PROV|6|6|懶惰人哪， 你去察看螞蟻的動作，就可得智慧。
PROV|6|7|螞蟻沒有領袖， 沒有官長，沒有君王，
PROV|6|8|尚且在夏天預備食物， 在收割時儲存糧食。
PROV|6|9|懶惰人哪，你要睡到幾時呢？ 你甚麼時候才睡醒呢？
PROV|6|10|再睡片時，打盹片時， 抱著雙臂躺臥片時，
PROV|6|11|你的貧窮就如盜賊來到， 你的貧乏彷彿拿盾牌的人來臨。
PROV|6|12|無賴的惡徒 行事全憑歪曲的口，
PROV|6|13|他眨眼傳神， 以腳示意，用指點劃，
PROV|6|14|存心乖謬， 常設惡謀，散播紛爭。
PROV|6|15|所以，災難必突然臨到他， 他必頃刻被毀，無從醫治。
PROV|6|16|耶和華所恨惡的有六樣， 他心所憎惡的共有七樣：
PROV|6|17|就是高傲的眼，撒謊的舌， 殺害無辜的手，
PROV|6|18|圖謀惡計的心， 飛奔行惡的腳，
PROV|6|19|口吐謊言的假證人， 並在弟兄間散播紛爭的人。
PROV|6|20|我兒啊，要遵守你父親的命令， 不可離棄你母親的教誨。
PROV|6|21|要常掛在你心上， 繫在你頸項上。
PROV|6|22|你行走，她必引導你， 你躺臥，她必保護你， 你睡醒，她必與你談論。
PROV|6|23|因為誡命是燈，教誨是光， 管教的責備是生命的道，
PROV|6|24|要保護你遠離邪惡的婦女， 遠離外邦女子諂媚的舌頭。
PROV|6|25|你不要因她的美色而動心， 也不要被她的眼皮勾引。
PROV|6|26|因為連最後一塊餅都會被妓女拿走 ； 有夫之婦會獵取寶貴的生命。
PROV|6|27|人若兜火在懷中， 他的衣服豈能不燒著呢？
PROV|6|28|人若走在火炭上， 他的腳豈能不燙傷呢？
PROV|6|29|與鄰舍之妻同寢的，也是如此， 凡親近她的，難免受罰。
PROV|6|30|賊因飢餓偷竊充飢， 人不藐視他，
PROV|6|31|但若被抓到，要賠償七倍， 他必賠上家中一切財物。
PROV|6|32|與婦人行姦淫的，便是無知， 做這事的，必毀了自己。
PROV|6|33|他必受損傷和羞辱， 他的羞恥不得消除。
PROV|6|34|丈夫因嫉恨發怒， 報仇的時候絕不留情。
PROV|6|35|他不接受任何賠償， 你送許多禮物，他也不肯和解。
PROV|7|1|我兒啊，要遵守我的言語， 存記我的命令。
PROV|7|2|遵守我的命令就得存活， 謹守我的教誨，好像保護眼中的瞳人。
PROV|7|3|要繫在你指頭上， 刻在你心版上。
PROV|7|4|對智慧說「你是我的姊妹」， 稱呼聰明為親人，
PROV|7|5|她就保護你遠離陌生女子， 遠離油嘴滑舌的外邦女子。
PROV|7|6|我曾在我房屋的窗戶內， 透過窗格子往外觀看，
PROV|7|7|看見在愚蒙人中， 注意到孩兒中有一個無知的青年，
PROV|7|8|從街上經過，靠近她的巷口， 直往她家的路去，
PROV|7|9|在黃昏，在傍晚， 在半夜，黑暗之中。
PROV|7|10|看哪，有一個女子來迎接他， 是妓女的打扮，有詭詐的心思。
PROV|7|11|她喧嚷，不守約束， 她的腳在家裏留不住，
PROV|7|12|有時在街市，有時在廣場， 或在各巷口等候。
PROV|7|13|她拉住那青年吻他， 厚著臉皮對他說：
PROV|7|14|「我已獻了平安祭， 今日我還了所許的願。
PROV|7|15|因此，我出來迎接你， 渴望見你的面，我總算找到你了！
PROV|7|16|我已在床上鋪好被單， 是 埃及 麻織的花紋布，
PROV|7|17|又用沒藥、沉香、桂皮 薰了我的床。
PROV|7|18|你來，讓我們飽享愛情，直到早晨， 讓我們彼此親愛歡樂。
PROV|7|19|因為我丈夫不在家， 出門遠行，
PROV|7|20|他手帶錢囊， 要到月圓才回家。」
PROV|7|21|這女子用許多巧言引誘他， 用諂媚的嘴唇催逼他。
PROV|7|22|青年立刻跟隨她，好像牛去被宰殺， 又像愚妄人帶著腳鐐去受刑，
PROV|7|23|直到箭穿進他的肝，如同雀鳥急投羅網， 卻不知會賠上自己的生命。
PROV|7|24|孩子們，現在要聽從我， 要留心聽我口中的言語。
PROV|7|25|你的心不可偏向她的道， 不要誤入她的迷途。
PROV|7|26|因為她擊倒許多人， 無數的人被她殺戮 。
PROV|7|27|她的家是在陰間之路， 下到死亡之宮。
PROV|8|1|智慧豈不呼喚？ 聰明豈不揚聲？
PROV|8|2|她站立在十字路口， 在道路旁高處的頂上，
PROV|8|3|在城門旁，城門口， 入口處，她呼喊：
PROV|8|4|「人哪，我呼喚你們， 我向世人揚聲。
PROV|8|5|愚蒙人哪，你們要學習靈巧， 愚昧人哪，你們的心要明辨。
PROV|8|6|你們當聽，因我要說尊貴的事， 我要張開嘴唇講正直的事。
PROV|8|7|我的口要發出真理， 我的嘴唇憎惡邪惡。
PROV|8|8|我口中的言語都是公義， 並無奸詐和歪曲。
PROV|8|9|聰明人看為正確， 有知識的，都以為正直。
PROV|8|10|你們當領受我的訓誨，勝過領受銀子， 寧得知識，強如得上選的金子。
PROV|8|11|「因為智慧比寶石更美， 一切可喜愛的都不足與其比較。
PROV|8|12|我－智慧以靈巧為居所， 又尋得知識和智謀。
PROV|8|13|敬畏耶和華就是恨惡邪惡； 我恨惡驕傲、狂妄、惡道，和乖謬的口。
PROV|8|14|我有策略和健全的知識， 我聰明，又有能力。
PROV|8|15|君王藉我治國， 王子藉我定公平，
PROV|8|16|王公貴族，所有公義的審判官， 都藉我掌權 。
PROV|8|17|愛我的，我也愛他， 懇切尋求我的，必尋見。
PROV|8|18|財富和尊榮在我， 恆久的財寶和繁榮 也在我。
PROV|8|19|我的果實勝過金子，強如純金， 我的出產超乎上選的銀子。
PROV|8|20|我在公義的道上走， 在公平的路中行，
PROV|8|21|使愛我的承受財產， 充滿他們的庫房。
PROV|8|22|「耶和華在造化的起頭， 在太初創造萬物之先，就有 了我。
PROV|8|23|從亙古，從太初， 未有大地以前，我已被立。
PROV|8|24|沒有深淵， 沒有大水的泉源，我已出生。
PROV|8|25|大山未曾奠定， 小山未有之先，我已出生。
PROV|8|26|那時，他還沒有創造大地和田野， 並世上頭一撮塵土。
PROV|8|27|他立高天，我在那裏， 他在淵面的周圍劃出圓圈，
PROV|8|28|上使穹蒼堅硬， 下使淵源穩固，
PROV|8|29|為滄海定出範圍，使水不越過界限， 奠定大地的根基。
PROV|8|30|那時，我在他旁邊為工程師， 天天充滿喜樂，時時在他面前歡笑，
PROV|8|31|在他的全地歡笑， 喜愛住在人世間。
PROV|8|32|「孩子們，現在要聽從我， 謹守我道的有福了。
PROV|8|33|要聽訓誨，得智慧， 不可棄絕。
PROV|8|34|聽從我，天天在我門口守望， 在我門框旁等候的，那人有福了。
PROV|8|35|因為尋得我的，就尋得生命， 他必蒙耶和華的恩惠。
PROV|8|36|得罪我的，害了自己的生命， 凡恨惡我的，喜愛死亡。」
PROV|9|1|智慧建造房屋， 鑿成七根柱子，
PROV|9|2|宰殺牲畜，調好美酒， 又擺設筵席，
PROV|9|3|派遣女僕出去， 自己在城中至高處呼喚：
PROV|9|4|「誰是愚蒙的人，讓他轉到這裏來！」 又對那無知的人說：
PROV|9|5|「你們來，吃我的餅， 喝我調的酒。
PROV|9|6|你們要離棄愚蒙，就得存活， 並要走明智的道路。」
PROV|9|7|糾正傲慢人的，必招羞辱， 責備惡人的，必被侮辱。
PROV|9|8|不要責備傲慢人，免得他恨你； 要責備智慧人，他必愛你。
PROV|9|9|教導智慧人，他就越有智慧， 指示義人，他就增長學問。
PROV|9|10|敬畏耶和華是智慧的開端， 認識至聖者便是聰明。
PROV|9|11|藉著我，你的日子必增多， 你生命的年數也必加添。
PROV|9|12|你若有智慧，是自己有智慧； 你若傲慢，就自己承擔。
PROV|9|13|愚昧的女子喧嚷， 她是愚蒙，一無所知。
PROV|9|14|她坐在自己家門口， 在城中高處的座位上，
PROV|9|15|呼喚過路的， 向那些在路上直走的人說：
PROV|9|16|「誰是愚蒙的人，讓他轉到這裏來！」 又對那無知的人說：
PROV|9|17|「偷來的水是甜的， 暗藏的餅是美的。」
PROV|9|18|人卻不知有陰魂在她那裏， 她召喚的人是在陰間的深處。
PROV|10|1|所羅門的箴言： 智慧之子使父親喜樂； 愚昧之子使母親擔憂。
PROV|10|2|不義之財毫無益處； 惟有公義能救人脫離死亡。
PROV|10|3|耶和華不使義人捱餓； 惡人所欲的，耶和華必拒絕。
PROV|10|4|手懶的，必致窮乏； 手勤的，卻要富足。
PROV|10|5|夏天儲存的，是智慧之子； 收割時沉睡的，是蒙羞之子。
PROV|10|6|福祉臨到義人頭上； 惡人的口藏匿殘暴。
PROV|10|7|義人的稱號帶來祝福； 惡人的名字必然敗壞。
PROV|10|8|智慧的心，領受誡命； 愚妄的嘴唇，必致傾倒。
PROV|10|9|行正直路的，步步安穩； 走彎曲道的，必致敗露。
PROV|10|10|擠眉弄眼的，使人憂患； 愚妄的嘴唇，必致傾倒。
PROV|10|11|義人的口是生命的泉源； 惡人的口藏匿殘暴。
PROV|10|12|恨能挑啟爭端； 愛能遮掩一切過錯。
PROV|10|13|聰明人嘴裏有智慧； 無知的人背上受刑杖。
PROV|10|14|智慧人積存知識； 愚妄人的口速致敗壞。
PROV|10|15|有錢人的財物是他堅固的城； 貧寒人的貧乏使他敗壞。
PROV|10|16|義人的報酬帶來生命； 惡人的所得用來犯罪。
PROV|10|17|遵守訓誨的，行在生命道上； 離棄責備的，走迷了路。
PROV|10|18|隱藏怨恨的，有說謊的嘴唇； 口出毀謗的，是愚昧人。
PROV|10|19|多言多語難免有過； 節制嘴唇是有智慧。
PROV|10|20|義人的舌如上選的銀子； 惡人的心所值無幾。
PROV|10|21|義人的嘴唇牧養多人； 愚妄人因無知而死亡。
PROV|10|22|耶和華所賜的福使人富足， 並不加上憂慮。
PROV|10|23|愚昧人以行惡為樂； 聰明人以智慧為樂。
PROV|10|24|惡人所怕的，必臨到他； 義人的心願，必蒙應允。
PROV|10|25|暴風一過，惡人歸於無有； 義人卻有永久的根基。
PROV|10|26|懶惰人使那差他的人， 如醋倒牙，如煙薰目。
PROV|10|27|敬畏耶和華使人長壽； 惡人的年歲必減少。
PROV|10|28|義人的盼望帶來喜樂； 惡人的指望必致滅沒。
PROV|10|29|耶和華的道是正直人的保障； 卻成了作惡人的敗壞。
PROV|10|30|義人永不動搖； 惡人不得住在地上。
PROV|10|31|義人的口結出智慧； 乖謬的舌必被割斷。
PROV|10|32|義人的嘴唇懂得令人喜悅； 惡人的口只知乖謬。
PROV|11|1|詭詐的天平為耶和華所憎惡； 公平的法碼為他所喜悅。
PROV|11|2|驕傲來，羞恥也來； 謙遜人卻有智慧。
PROV|11|3|正直人的純正必引導自己； 奸詐人的邪惡必毀滅自己。
PROV|11|4|遭怒的日子錢財無益； 惟有公義能救人脫離死亡。
PROV|11|5|完全人的義修平自己的路； 但惡人必因自己的惡跌倒。
PROV|11|6|正直人的義必拯救自己； 奸詐人必被自己的慾望纏住。
PROV|11|7|惡人一死，他的指望就滅絕； 罪人的盼望也必滅絕。
PROV|11|8|義人得脫離患難， 有惡人來代替他。
PROV|11|9|不虔敬的人用口敗壞鄰舍； 義人卻因知識得救。
PROV|11|10|義人享福，全城喜樂； 惡人滅亡，人人歡呼。
PROV|11|11|因正直人的祝福，城必升高； 因邪惡人的口，它必傾覆。
PROV|11|12|藐視鄰舍的，便是無知； 聰明人卻靜默不言。
PROV|11|13|到處傳話的，洩漏機密； 內心老實的，保守祕密。
PROV|11|14|無智謀，民就敗落； 謀士多，就必得勝。
PROV|11|15|為陌生人擔保的，必受虧損； 恨惡擊掌的，卻得安穩。
PROV|11|16|恩慈的婦女得尊榮； 強壯的男子得財富。
PROV|11|17|仁慈的人善待自己； 殘忍的人擾害己身。
PROV|11|18|惡人做事，得虛幻的報酬； 撒公義種子的，得實在的報償。
PROV|11|19|真正行義的，必得生命； 追求邪惡的，必致死亡。
PROV|11|20|心中歪曲的，為耶和華所憎惡； 行為正直的，為他所喜悅。
PROV|11|21|擊掌保證，惡人難免受罰； 義人的後裔必得拯救。
PROV|11|22|婦女美貌而無見識， 如同金環戴在豬鼻上。
PROV|11|23|義人的心願盡是好的； 惡人的指望卻帶來憤怒。
PROV|11|24|有施捨的，錢財增添； 吝惜過度，反致窮乏。
PROV|11|25|慷慨待人，必然豐裕； 滋潤人的，連自己也得滋潤。
PROV|11|26|屯糧不賣的，百姓必詛咒他； 願意出售的，祝福臨到頭上。
PROV|11|27|懇切求善的，就求得恩寵； 但那求惡的，惡必臨到他。
PROV|11|28|倚靠財富的，自己必跌倒； 義人必興旺如綠葉。
PROV|11|29|擾害己家的，必承受虛空 ； 愚妄人作心中有智慧者的僕人。
PROV|11|30|義人的果實是生命樹； 智慧人必能得人。
PROV|11|31|看哪，義人在地上尚且受報， 何況惡人和罪人呢？
PROV|12|1|喜愛管教的，就是喜愛知識； 恨惡責備的，卻像畜牲。
PROV|12|2|善人蒙耶和華的恩寵； 設詭計的，耶和華必定罪。
PROV|12|3|人靠惡行不能堅立； 義人的根必不動搖。
PROV|12|4|才德的妻子是丈夫的冠冕； 蒙羞的婦人使丈夫骨頭朽爛。
PROV|12|5|義人的思念是公平； 惡人的計謀是詭詐。
PROV|12|6|惡人的言論埋伏流人的血； 正直人的口卻拯救人。
PROV|12|7|惡人傾覆，歸於無有； 義人的家卻屹立不倒。
PROV|12|8|人按自己的智慧得稱讚； 心中偏邪的，必被藐視。
PROV|12|9|被人藐視，但有自己僕人 的， 勝過妄自尊大，卻缺乏食物。
PROV|12|10|義人顧惜他牲畜的命； 惡人的憐憫也是殘忍。
PROV|12|11|耕種自己田地的，必得飽食； 追求虛浮的，卻是無知。
PROV|12|12|惡人想得壞人的獵物； 義人的根結出果實。
PROV|12|13|嘴唇的過錯是惡人的圈套； 但義人必脫離患難。
PROV|12|14|人因口所結的果實，必飽得美福； 人手所做的，必歸到自己身上。
PROV|12|15|愚妄人所行的，在自己眼中看為正直； 惟智慧人從善如流。
PROV|12|16|愚妄人的惱怒立時顯露； 通達人卻能忍辱。
PROV|12|17|說出真話的，顯明公義； 作假見證的，顯出詭詐。
PROV|12|18|說話浮躁，猶如刺刀； 智慧人的舌頭卻能醫治。
PROV|12|19|誠實的嘴唇永遠堅立； 說謊的舌頭只存片時。
PROV|12|20|圖謀惡事的，心存詭詐； 勸人和睦的，便得喜樂。
PROV|12|21|義人不遭災害； 惡人滿受禍患。
PROV|12|22|說謊的嘴唇，為耶和華所憎惡； 行事誠實，為他所喜悅。
PROV|12|23|通達人隱藏知識； 愚昧人的心彰顯愚昧。
PROV|12|24|殷勤人的手必掌權； 懶惰的人必服苦役。
PROV|12|25|人心憂慮，就必沉重； 一句良言，使心歡樂。
PROV|12|26|義人引導他的鄰舍 ； 惡人的道叫人迷失。
PROV|12|27|懶惰的人不烤獵物； 殷勤的人卻得寶貴的財物。
PROV|12|28|在公義的路上有生命； 在其道上並無死亡。
PROV|13|1|智慧之子聽父親的訓誨； 傲慢人不聽責備。
PROV|13|2|人因口所結的果實，必享美福； 奸詐人卻意圖殘暴。
PROV|13|3|謹慎守口的，得保生命； 大張嘴唇的，必致敗亡。
PROV|13|4|懶惰的人奢求，卻無所得； 殷勤的人必然豐裕。
PROV|13|5|義人恨惡謊言； 惡人可憎可恥。
PROV|13|6|行為純正的，有公義保護； 犯罪的，被罪惡傾覆。
PROV|13|7|假冒富足的，一無所有； 裝作窮乏的，多有財物。
PROV|13|8|財富可作人的生命贖價； 窮乏人卻聽不見威嚇的話。
PROV|13|9|義人的光使人歡喜 ； 惡人的燈要熄滅。
PROV|13|10|驕傲挑啟紛爭； 聽勸言卻有智慧。
PROV|13|11|不勞而獲之財 必減少； 逐漸積蓄的必增多。
PROV|13|12|盼望遲延，令人心憂； 願望實現，就是得到生命樹。
PROV|13|13|藐視訓言的，自取滅亡； 敬畏誡命的，必得善報。
PROV|13|14|智慧人的教誨是生命的泉源， 使人避開死亡的圈套。
PROV|13|15|美好的見識使人得寵； 奸詐人的道路恆久奸詐 。
PROV|13|16|通達人都憑知識行事； 愚昧人張揚自己的愚昧。
PROV|13|17|邪惡的使者必陷入禍患； 忠信的使臣帶來醫治。
PROV|13|18|棄絕管教的，必貧窮受辱； 領受責備的，必享尊榮。
PROV|13|19|願望實現，心覺甘甜； 遠離惡事，為愚昧人所憎惡。
PROV|13|20|與智慧人同行的，必得智慧； 和愚昧人作伴的，必受虧損。
PROV|13|21|禍患追趕罪人； 義人卻得善報。
PROV|13|22|善人給子孫遺留產業； 罪人積財卻歸義人。
PROV|13|23|窮乏人開墾的地雖多產糧食， 卻因不公而被奪走。
PROV|13|24|不忍用杖打兒子的，是恨惡他； 疼愛兒子的，勤加管教。
PROV|13|25|義人吃喝食慾滿足； 惡人肚腹卻是缺乏。
PROV|14|1|婦人的智慧建立家室； 愚昧卻親手拆毀它 。
PROV|14|2|行事正直的，敬畏耶和華； 偏離正路的，卻藐視他。
PROV|14|3|在愚妄人的口中有驕傲的杖； 智慧人的嘴唇必保護自己。
PROV|14|4|沒有牛，槽就空空； 土產豐盛卻憑牛的力氣。
PROV|14|5|誠實的證人不說謊； 虛假的證人口吐謊言。
PROV|14|6|傲慢人枉尋智慧； 聰明人易得知識。
PROV|14|7|不要到愚昧人面前， 你無法從他嘴唇裏知道知識。
PROV|14|8|通達人的智慧使他認清自己的道路； 愚昧人的愚昧卻是自欺。
PROV|14|9|愚妄人嘲笑贖愆祭 ； 但正直人蒙悅納。
PROV|14|10|心中的苦楚，只有自己知道； 心裏的喜樂，陌生人無法分享。
PROV|14|11|惡人的房屋必倒塌； 正直人的帳棚必興旺。
PROV|14|12|有一條路，人以為正， 至終成為死亡之路。
PROV|14|13|人在喜笑中，心也會憂愁； 快樂的終點就是愁苦。
PROV|14|14|心中背道的，必滿嘗其果； 善人必從自己的行為得到回報。
PROV|14|15|無知的人甚麼話都信； 通達人謹慎自己的腳步。
PROV|14|16|智慧人有所懼怕，就遠離惡事； 愚昧人卻狂傲自恃。
PROV|14|17|輕易發怒的，行事愚昧； 擅長詭計的，被人恨惡。
PROV|14|18|愚蒙人承受愚昧為產業； 通達人得知識為冠冕。
PROV|14|19|壞人在善人面前俯伏； 惡人在義人門口也是如此。
PROV|14|20|窮乏人，連鄰舍也恨他； 有錢人，愛他的人眾多。
PROV|14|21|藐視鄰舍的，這人有罪； 施恩給困苦人的，這人有福。
PROV|14|22|謀惡的，豈非走入迷途？ 謀善的，有慈愛和誠實。
PROV|14|23|任何勤勞總有收穫； 僅耍嘴皮必致窮乏。
PROV|14|24|智慧人的冠冕是富有智慧； 愚昧人的愚昧終究是愚昧。
PROV|14|25|誠實作證，救人性命； 口吐謊言是詭詐。
PROV|14|26|敬畏耶和華的，大有倚靠； 他的兒女也有避難所。
PROV|14|27|敬畏耶和華是生命的泉源， 使人離開死亡的圈套。
PROV|14|28|君王的榮耀在乎民多； 沒有百姓，王就衰敗。
PROV|14|29|不輕易發怒的，大有聰明； 性情暴躁的，大顯愚昧。
PROV|14|30|平靜的心使肉體有生氣； 嫉妒使骨頭朽爛。
PROV|14|31|欺壓貧寒人的，是蔑視造他的主； 憐憫貧窮人的，是尊敬主。
PROV|14|32|惡人因所行的惡必被推倒； 義人臨死 ，有所投靠。
PROV|14|33|智慧安居在聰明人的心中， 在愚昧人的心中卻不認識 。
PROV|14|34|公義使邦國高舉； 罪惡是百姓的羞辱。
PROV|14|35|君王的恩寵臨到智慧的臣僕； 但其憤怒臨到蒙羞的臣僕。
PROV|15|1|回答柔和，使怒消退； 言語粗暴，觸動怒氣。
PROV|15|2|智慧人的舌善發知識； 愚昧人的口吐出愚昧。
PROV|15|3|耶和華的眼目無處不在， 惡人善人，他都鑒察。
PROV|15|4|溫良的舌是生命樹； 邪惡的舌使人心碎。
PROV|15|5|愚妄人藐視父親的管教； 領受責備，使人精明。
PROV|15|6|義人家中多有財富； 惡人獲利反受擾害。
PROV|15|7|智慧人的嘴傳揚知識； 愚昧人的心並非如此。
PROV|15|8|惡人獻祭，為耶和華所憎惡； 正直人祈禱，為他所喜悅。
PROV|15|9|惡人的道路，為耶和華所憎惡； 追求公義的，為他所喜愛。
PROV|15|10|背棄正路的，必受嚴刑； 恨惡責備的，必致死亡。
PROV|15|11|陰間和冥府 尚且在耶和華面前， 何況世人的心呢？
PROV|15|12|傲慢人不愛受責備， 也不去接近智慧人。
PROV|15|13|心中喜樂，面有喜色； 心裏憂愁，靈就憂傷。
PROV|15|14|聰明人的心追求知識； 愚昧人的口吞吃愚昧。
PROV|15|15|困苦人的日子都是愁苦； 心中歡暢的，常享宴席。
PROV|15|16|財寶稀少，敬畏耶和華， 強如財寶眾多，煩亂不安。
PROV|15|17|有愛，吃素菜， 強如相恨，吃肥牛。
PROV|15|18|暴怒的人挑啟爭端； 忍怒的人止息紛爭。
PROV|15|19|懶惰人的道像荊棘的籬笆； 正直人的路是平坦大道。
PROV|15|20|智慧之子使父親喜樂； 愚昧的人藐視母親。
PROV|15|21|無知的人以愚昧為樂； 聰明的人按正直而行。
PROV|15|22|不先商議，所謀無效； 謀士眾多，所謀得成。
PROV|15|23|口善應對，自覺喜樂； 話合其時，何等美好。
PROV|15|24|生命之道使智慧人上升， 使他遠離底下的陰間。
PROV|15|25|耶和華必拆毀驕傲人的家， 卻要立定寡婦的地界。
PROV|15|26|惡謀為耶和華所憎惡； 良言卻是純淨的。
PROV|15|27|暴力歛財的，擾害己家； 恨惡賄賂的，必得存活。
PROV|15|28|義人的心思量應答； 惡人的口吐出惡言。
PROV|15|29|耶和華遠離惡人， 卻聽義人的祈禱。
PROV|15|30|眼睛發光，使心喜樂； 好的信息，滋潤骨頭。
PROV|15|31|耳聽使人得生命的責備， 必居住在智慧人之中。
PROV|15|32|棄絕管教的，輕看自己的生命； 領受責備的，卻得智慧的心。
PROV|15|33|敬畏耶和華是智慧的訓誨； 要得尊榮，先有謙卑。
PROV|16|1|心中的籌謀在乎人， 舌頭的應對出於耶和華。
PROV|16|2|人一切所行的，在自己眼中看為純潔， 惟有耶和華衡量人的內心。
PROV|16|3|你所做的，要交託耶和華， 你所謀的，就必堅立。
PROV|16|4|耶和華造萬物各適其用， 就是惡人也為禍患的日子所造。
PROV|16|5|凡心裏驕傲的，為耶和華所憎惡； 擊掌保證，他難免受罰。
PROV|16|6|因慈愛和信實，罪孽得贖； 敬畏耶和華的，遠離惡事。
PROV|16|7|人所行的若蒙耶和華喜悅， 耶和華也使仇敵與他和好。
PROV|16|8|少獲利，行事公義， 強如多獲利，行事不義。
PROV|16|9|人心籌算自己的道路； 惟耶和華指引他的腳步。
PROV|16|10|王的嘴唇有聖言， 審判之時，他的口必不差錯。
PROV|16|11|公道的秤和天平屬耶和華， 囊中一切的法碼是他所定。
PROV|16|12|作惡，為王所憎惡， 因國位是靠公義堅立。
PROV|16|13|公義的嘴唇，王喜悅， 說正直話的，他喜愛。
PROV|16|14|王的震怒是死亡的使者， 但智慧人能平息王怒。
PROV|16|15|王臉上的光使人有生命， 他的恩惠好像雲帶來的春雨。
PROV|16|16|得智慧勝過得金子， 選聰明強如選銀子。
PROV|16|17|正直人的道遠離惡事， 謹守己路的，保全性命。
PROV|16|18|驕傲在敗壞以先， 內心高傲在跌倒之前。
PROV|16|19|心裏謙卑與困苦人來往， 強如與驕傲人同分戰利品。
PROV|16|20|留心訓言的 ，必得福樂； 倚靠耶和華的，這人有福。
PROV|16|21|心中有智慧的，必稱為聰明人； 嘴唇的甜言，增長人的學問。
PROV|16|22|人有智慧就有生命的泉源； 愚妄人必受愚妄的懲戒。
PROV|16|23|智慧人的心使他的口謹慎， 又使他的嘴唇增長學問。
PROV|16|24|良言如同蜂巢， 使心甘甜，使骨得醫治。
PROV|16|25|有一條路，人以為正， 至終卻成為死亡之路。
PROV|16|26|勞力的人為自己勞力， 因為他的口腹催逼他。
PROV|16|27|匪徒圖謀奸惡， 嘴唇上的言語彷彿燒焦的火。
PROV|16|28|乖謬的人散播紛爭， 造謠的離間密友。
PROV|16|29|殘暴的人引誘鄰舍， 領他走不好的道路。
PROV|16|30|緊閉雙目的，圖謀乖謬； 緊咬嘴唇的，成就惡事。
PROV|16|31|白髮是榮耀的冠冕， 行在公義道上的，必能得著。
PROV|16|32|不輕易發怒的，勝過勇士； 控制自己脾氣的，強如取城。
PROV|16|33|人雖可擲籤在膝上， 定事卻由耶和華。
PROV|17|1|一塊乾餅，大家相安； 勝過宴席滿屋，大家相爭。
PROV|17|2|明智的僕人必管轄蒙羞的兒子， 並在兄弟中同分產業。
PROV|17|3|鼎為煉銀，爐為煉金， 惟有耶和華熬煉人心。
PROV|17|4|行惡的，留心聽惡毒的嘴唇； 說謊的，側耳聽邪惡的舌頭。
PROV|17|5|譏笑窮乏人的，是蔑視造他的主； 幸災樂禍的，難免受罰。
PROV|17|6|子孫為老人的冠冕； 父母是兒女的榮耀。
PROV|17|7|愚頑人說美言並不相宜， 君子說謊言也不合宜。
PROV|17|8|賄賂在餽贈者的眼中看為玉石， 隨處運轉都得順利。
PROV|17|9|包容過錯的，尋求友愛； 喋喋不休的，離間密友。
PROV|17|10|一句責備的話深入聰明人的心， 強如打愚昧人一百下。
PROV|17|11|惡人只尋求背叛， 殘忍的使者必奉差攻擊他。
PROV|17|12|寧可遇見失喪小熊的母熊， 也不願遇見正行愚昧的愚昧人。
PROV|17|13|以惡報善的， 禍患必不離他的家。
PROV|17|14|紛爭掀起，如同缺口的水； 因此，爭端尚未爆發就當制止。
PROV|17|15|定惡人為義的，定義人為有罪的， 都為耶和華所憎惡。
PROV|17|16|愚昧人既無知， 為何手拿銀錢去買智慧呢？
PROV|17|17|朋友時常親愛， 弟兄為患難而生。
PROV|17|18|在鄰舍面前擊掌擔保的， 是無知的人。
PROV|17|19|喜愛爭吵的，是喜愛過犯； 門蓋得高的，自取敗壞。
PROV|17|20|心中歪曲的，得不著福樂； 舌頭顛倒是非的，陷在禍患中。
PROV|17|21|生愚昧之子的，自己必愁苦； 愚頑人的父親毫無喜樂。
PROV|17|22|喜樂的心能治好疾病； 憂傷的靈使骨頭枯乾。
PROV|17|23|惡人暗中受賄賂， 以致彎曲公正的路。
PROV|17|24|聰明人面前有智慧； 愚昧人眼望地的盡頭。
PROV|17|25|愚昧的兒子使父親愁煩， 使那生他的母親憂苦。
PROV|17|26|刑罰義人實為不善， 責打正直的君子也不宜。
PROV|17|27|節制言語的，有見識； 性情溫良的人，有聰明。
PROV|17|28|愚妄人若靜默不言，可算為智慧， 閉上嘴唇也可算為聰明。
PROV|18|1|孤僻的人只顧自己的心願 ， 他鄙視一切健全的知識。
PROV|18|2|愚昧人不喜愛聰明， 只喜愛表達自己的心意。
PROV|18|3|邪惡來，藐視跟著來； 羞恥到，辱罵同時到。
PROV|18|4|人的口所講的話如同深水， 智慧之泉如湧流的河水。
PROV|18|5|偏袒惡人的情面，是不好的。 審判時使義人受屈，也是不善。
PROV|18|6|愚昧人的嘴唇挑起爭端， 一開口就招鞭打。
PROV|18|7|愚昧人的口自取敗壞， 他的嘴唇是自己生命的圈套。
PROV|18|8|造謠者的話如同美食， 深入人的肚腹。
PROV|18|9|做工懈怠的， 是破壞者的兄弟。
PROV|18|10|耶和華的名是堅固臺， 義人奔入就得安穩。
PROV|18|11|有錢人的財物是他堅固的城， 在他幻想中，猶如高牆。
PROV|18|12|敗壞之先，人心驕傲； 要得尊榮，先有謙卑。
PROV|18|13|未聽完就回話的， 就是他的愚昧和羞辱。
PROV|18|14|人的心靈忍耐疾病； 心靈憂傷，誰能承當呢？
PROV|18|15|聰明人的心得知識； 智慧人的耳求知識。
PROV|18|16|人的禮物為他開路， 引他到高位的人面前。
PROV|18|17|先訴情由的，似乎有理； 另一人來到，就察出實情。
PROV|18|18|掣籤能止息紛爭， 也能化解雙方激烈的爭辯。
PROV|18|19|被冒犯的弟兄 強如難以攻下的堅城； 紛爭如同城堡的門閂。
PROV|18|20|人的肚腹必因口所結的果實飽足； 他必因嘴唇所出的感到滿足。
PROV|18|21|生死在舌頭的掌握之下， 喜愛弄舌的，必吃它所結的果實。
PROV|18|22|得著妻子的，得著好處， 他是蒙了耶和華的恩惠。
PROV|18|23|窮乏人說哀求的話； 有錢人卻用威嚇的話回答。
PROV|18|24|朋友太多的人，必受損害 ； 但有一知己比兄弟更親密。
PROV|19|1|行為純正的窮乏人 勝過嘴唇歪曲的愚昧人。
PROV|19|2|熱心而無見識，實為不善； 腳步急快的，易入歧途。
PROV|19|3|人因愚昧自毀前途， 他的心卻埋怨耶和華。
PROV|19|4|財富使朋友增多； 貧寒人連僅有的朋友也離棄他。
PROV|19|5|作假見證的，難免受罰； 口吐謊言的，不能逃脫。
PROV|19|6|有權貴的，許多人求他賞臉； 愛送禮的，人都作他的朋友。
PROV|19|7|窮乏人連兄弟都恨他， 何況朋友，更是遠離他！ 他用言語追隨，他們卻不在。
PROV|19|8|得著智慧的，愛惜生命； 持守聰明的，尋得好處。
PROV|19|9|作假見證的，難免受罰； 口吐謊言的，必定滅亡。
PROV|19|10|愚昧人奢華度日並不相宜， 僕人管轄王子，也不應該。
PROV|19|11|人有見識就不輕易發怒， 寬恕人的過失便是自己的榮耀。
PROV|19|12|王的憤怒好像獅子吼叫； 他的恩惠卻如草上的甘露。
PROV|19|13|愚昧的兒子是父親的禍患， 妻子的爭吵如雨連連滴漏。
PROV|19|14|房屋錢財是祖宗所遺留的； 惟有賢慧的妻是耶和華所賜的。
PROV|19|15|懶惰使人沉睡， 懈怠的人必捱餓。
PROV|19|16|遵守誡命的，保全生命； 輕忽己路的，必致死亡。
PROV|19|17|憐憫貧寒人的，就是借給耶和華， 他的報償，耶和華必歸還他。
PROV|19|18|趁還有指望，管教你的兒子， 不可執意摧毀他。
PROV|19|19|暴怒的人必受懲罰， 你若救他，必須再救。
PROV|19|20|要聽勸言，接受訓誨， 使你終久有智慧。
PROV|19|21|人心多有計謀； 惟有耶和華的籌算才能成就。
PROV|19|22|仁慈的人令人喜愛 ， 窮乏人強如說謊言的。
PROV|19|23|敬畏耶和華的，得著生命， 他必飽足安居，不遭禍患。
PROV|19|24|懶惰人把手埋入盤裏， 連縮回送進口中也不肯。
PROV|19|25|責打傲慢人，能使無知的人變精明； 責備聰明人，他就明白知識。
PROV|19|26|虐待父親、驅逐母親的， 是蒙羞致辱之子。
PROV|19|27|我兒啊，停止聽 那叫你偏離知識言語的教導 。
PROV|19|28|卑劣的見證嘲笑公平， 惡人的口吞下罪孽。
PROV|19|29|刑罰是為傲慢人預備的， 鞭打則是為愚昧人的背預備的。
PROV|20|1|酒能使人傲慢，烈酒使人喧嚷， 凡沉溺其中的，都無智慧。
PROV|20|2|王的威嚇如獅子吼叫， 激怒他的是自害己命。
PROV|20|3|止息紛爭是人的尊榮， 愚妄人爭鬧不休。
PROV|20|4|懶惰人因冬寒不去耕種， 到收割時，他去尋找，一無所得。
PROV|20|5|人心中的籌算如同深水， 惟聰明人才能汲引出來。
PROV|20|6|很多人聲稱自己忠信， 但誠信的人誰能遇著呢？
PROV|20|7|義人行為純正， 他後代的子孫有福了！
PROV|20|8|王坐在審判的位上， 以眼目驅散一切邪惡。
PROV|20|9|誰能說：「我已經潔淨了我的心， 脫淨了我的罪？」
PROV|20|10|兩樣的法碼和兩樣的伊法 ， 都為耶和華所憎惡。
PROV|20|11|孩童的行動或純潔，或正直， 都以行為顯明自己。
PROV|20|12|能聽的耳，能看的眼， 二者都為耶和華所造。
PROV|20|13|不要貪睡，免致貧窮； 眼要睜開，就可吃飽。
PROV|20|14|買東西的說：「不好，不好！」 及至離去，他卻自誇。
PROV|20|15|有金子和許多寶石， 惟知識的嘴唇是貴重的珍寶。
PROV|20|16|誰為陌生人擔保，就拿誰的衣服； 誰為外邦人作保，誰就要承當。
PROV|20|17|靠謊言而得的食物，令人愉悅； 到後來，他的口必充滿碎石。
PROV|20|18|計謀憑籌算立定， 打仗要憑智謀。
PROV|20|19|到處傳話的，洩漏機密； 口無遮攔的，不可與他結交。
PROV|20|20|咒罵父母的， 他的燈必熄滅，在漆黑中。
PROV|20|21|起初很快得來的產業， 終久卻不是福。
PROV|20|22|你不要說：「我要以惡報惡」； 要等候耶和華，他必拯救你。
PROV|20|23|兩樣的法碼為耶和華所憎惡， 詭詐的天平也為不善。
PROV|20|24|人的腳步為耶和華所定， 人豈能明白自己的道路呢？
PROV|20|25|人冒失地聲稱：「這是神聖的！」 許願之後才細想，就是自陷圈套。
PROV|20|26|智慧的王驅散惡人， 用輪子滾過他們。
PROV|20|27|人的靈是耶和華的燈， 鑒察人的內心深處。
PROV|20|28|慈愛和誠實庇護君王， 他的王位因慈愛而立穩。
PROV|20|29|強壯是青年的榮耀； 白髮為老人的尊榮。
PROV|20|30|鞭傷除淨邪惡， 責打可潔淨人心深處。
PROV|21|1|王的心在耶和華手中像河水， 他能使它隨意流轉。
PROV|21|2|人一切所行的，在自己眼中看為正直， 惟有耶和華衡量人心。
PROV|21|3|行公義和公平 比獻祭更蒙耶和華悅納。
PROV|21|4|眼高心傲，就是惡人的燈， 都是罪。
PROV|21|5|殷勤籌劃的，足致豐裕； 行事急躁的，必致缺乏。
PROV|21|6|用詭詐之舌所得的財富 如被吹散的霧氣，趨向滅亡 。
PROV|21|7|惡人的殘暴必掃去自己， 因他們不肯按公平行事。
PROV|21|8|有罪的人其路彎曲； 純潔的人行為正直。
PROV|21|9|寧可住在房頂的一角， 也不與好爭吵的婦人同住。
PROV|21|10|惡人的心渴想邪惡， 他的眼並不憐憫鄰舍。
PROV|21|11|傲慢人受懲罰，愚蒙人可得智慧； 智慧人受訓誨，便得知識。
PROV|21|12|公義的上帝 鑒察惡人的家， 他傾覆惡人，以致滅亡。
PROV|21|13|塞耳不聽貧寒人哀求的， 他自己呼求，也不蒙應允。
PROV|21|14|暗中送的禮物挽回怒氣， 懷裏的賄賂能止息暴怒。
PROV|21|15|秉公行義使義人喜樂， 卻使作惡的人敗壞。
PROV|21|16|人偏離智慧的路， 必與陰魂為伍 。
PROV|21|17|愛宴樂的，必致窮乏； 貪愛酒和油的，必不富足。
PROV|21|18|惡人作義人的贖價， 奸詐人代替正直人。
PROV|21|19|寧可住在曠野之地， 也不與爭吵易怒的婦人同住。
PROV|21|20|智慧人的居所積蓄寶物與膏油 ； 愚昧人卻揮霍一空。
PROV|21|21|追求公義慈愛的， 就尋得生命、公義 和尊榮。
PROV|21|22|智慧人爬上勇士的城牆， 摧毀他所倚靠的堡壘。
PROV|21|23|謹守口和舌的， 就保護自己免受災難。
PROV|21|24|心驕氣傲的人名叫傲慢， 他行事出於狂妄驕傲。
PROV|21|25|懶惰人的慾望害死自己， 因為他的手不肯做工；
PROV|21|26|有人終日貪得無饜， 義人卻施捨而不吝惜。
PROV|21|27|惡人獻的祭是可憎的， 何況他存惡意來獻呢？
PROV|21|28|不實的見證必消滅； 惟聆聽真情的，他的證詞有力。
PROV|21|29|惡人臉無羞恥； 正直人行事堅定 。
PROV|21|30|沒有人能以智慧、聰明、 謀略抵擋耶和華。
PROV|21|31|馬是為打仗之日預備的； 得勝卻在於耶和華。
PROV|22|1|美名勝過大財， 宏恩強如金銀。
PROV|22|2|有錢人與窮乏人相遇 ， 他們都為耶和華所造。
PROV|22|3|通達人見禍就藏躲； 愚蒙人卻前往受害。
PROV|22|4|敬畏耶和華心存謙卑， 就得財富、尊榮、生命為賞賜。
PROV|22|5|歪曲的人路上有荊棘和羅網， 保護自己生命的，必要遠離。
PROV|22|6|教養孩童走當行的道， 就是到老他也不偏離。
PROV|22|7|有錢人管轄窮乏人， 欠債的是債主的僕人。
PROV|22|8|撒不義種子的必收割災禍， 他逞怒的杖也必廢掉。
PROV|22|9|眼目仁慈的必蒙福， 因他將食物分給貧寒人。
PROV|22|10|趕出傲慢人，爭端就消除， 紛爭和羞辱也必止息。
PROV|22|11|喜愛清心，嘴唇有恩言的， 王必與他為友。
PROV|22|12|耶和華的眼目保護知識， 卻毀壞奸詐人的言語。
PROV|22|13|懶惰人說：「外面有獅子， 我在街上必被殺害。」
PROV|22|14|陌生女子的口是深坑， 耶和華所憎惡的，必陷在其中。
PROV|22|15|愚昧迷住孩童的心， 用管教的杖可以遠遠趕除。
PROV|22|16|欺壓貧寒人為要利己的， 並送禮給有錢人的，都必缺乏。
PROV|22|17|你要側耳聽智慧人的言語 ， 留心領會我的知識。
PROV|22|18|你若心中存記， 嘴唇也準備就緒，這是美的。
PROV|22|19|我今日特地指教你， 為要使你倚靠耶和華。
PROV|22|20|謀略和知識的美事 ， 我豈沒有寫給你嗎？
PROV|22|21|要使你明白真情實理， 好將實情回覆那差你來的人。
PROV|22|22|不可因人貧寒就搶奪他， 也不可在城門口欺壓困苦人，
PROV|22|23|因耶和華必為他們辯護， 也必奪取那搶奪者的命。
PROV|22|24|不可結交好生氣的人， 也不可與暴怒的人來往，
PROV|22|25|恐怕你效法他的行為， 自己就陷在圈套裏。
PROV|22|26|不要為人擊掌擔保， 也不要為債務作保。
PROV|22|27|你若沒有甚麼可償還， 何必使人奪去你睡臥的床呢？
PROV|22|28|祖先所立的地界， 你不可挪移。
PROV|22|29|你看見辦事殷勤的人嗎？ 他必侍立在君王面前， 不在平庸的人面前。
PROV|23|1|你若與長官坐席， 要留意在你面前的是誰。
PROV|23|2|你若是胃口大的人， 就當拿刀放在喉嚨上。
PROV|23|3|不可貪戀長官的美食， 因為那是欺哄人的食物。
PROV|23|4|不要勞碌求富， 要有聰明來節制。
PROV|23|5|你定睛在財富，它就消失， 因為它必長翅膀，如鷹向天飛去。
PROV|23|6|守財奴 的飯，你不要吃， 也不要貪戀他的美味；
PROV|23|7|因為他的心怎樣算計 ， 他為人就是這樣。 他雖對你說：請吃，請喝， 他的心卻與你相背。
PROV|23|8|你所吃的那點食物必吐出來， 你恭維的話語也必落空。
PROV|23|9|不要說話給愚昧人聽， 因他必藐視你智慧的言語。
PROV|23|10|不可挪移古時的地界， 也不可侵佔孤兒的田地，
PROV|23|11|因他們的救贖者 大有能力， 他必向你為他們辯護。
PROV|23|12|你要留心領受訓誨， 側耳聽從知識的言語。
PROV|23|13|不可不管教孩童， 因為你用杖打他，他不會死。
PROV|23|14|你用杖打他， 就可以救他的性命免下陰間。
PROV|23|15|我兒啊，你若心存智慧， 我的心就甚歡喜。
PROV|23|16|你的嘴唇若說正直話， 我的心腸也必快樂。
PROV|23|17|你的心不要羨慕罪人， 卻要羨慕常常敬畏耶和華的人，
PROV|23|18|因為你必有前途， 你的指望也不致斷絕。
PROV|23|19|我兒啊，你當聽，當存智慧， 好在正道上引導你的心。
PROV|23|20|不可與好飲酒的人在一起， 也不要跟貪吃肉的人來往，
PROV|23|21|因為貪食好酒的，必致貧窮， 愛睡覺的，必穿破爛衣服。
PROV|23|22|你要聽從生你的父親； 不可因母親年老而輕看她。
PROV|23|23|你當獲得真理，不可出賣， 智慧、訓誨和聰明也是一樣。
PROV|23|24|義人的父親必大大快樂， 生智慧兒子的，必因他歡喜。
PROV|23|25|願你的父母歡喜， 願那生你的母親快樂。
PROV|23|26|我兒啊，要將你的心歸我， 你的眼目也要喜愛 我的道路。
PROV|23|27|妓女是深坑， 外邦女子是窄井。
PROV|23|28|她像強盜埋伏， 她使奸詐的人增多。
PROV|23|29|誰有禍患？誰有災難？ 誰有紛爭？誰有焦慮？ 誰無故受傷？誰的眼目紅赤？
PROV|23|30|就是那流連飲酒的人， 常去尋找調和的酒。
PROV|23|31|酒發紅，在杯中閃爍時， 你不可觀看； 雖下咽舒暢， 終究它必咬你如蛇，刺你如毒蛇。
PROV|23|32|
PROV|23|33|你的眼睛必看見怪異的事， 你的心必發出乖謬的話。
PROV|23|34|你必像躺在深海中， 或臥在桅杆頂上，
PROV|23|35|說：「人擊打我，但我未受傷， 重擊我，我不覺得。 我幾時清醒， 還要再去尋酒。」
PROV|24|1|你不要嫉妒惡人， 也不要渴望與他們相處，
PROV|24|2|因為他們的心圖謀暴行， 他們的嘴唇談論奸惡。
PROV|24|3|房屋因智慧建造， 因聰明立穩；
PROV|24|4|又因知識， 屋內充滿各樣美好寶貴的財物。
PROV|24|5|有智慧的勇士大有能力， 有知識的人力上加力。
PROV|24|6|你去打仗，要憑智謀； 謀士眾多，就必得勝。
PROV|24|7|對愚妄人，智慧高不可及， 所以他在城門不敢開口。
PROV|24|8|圖謀行惡的， 必稱為奸詐人。
PROV|24|9|愚妄人的籌劃盡是罪惡， 傲慢者為人所憎惡。
PROV|24|10|在患難時你若灰心， 你的力量就微小。
PROV|24|11|人被拉到死亡，你要解救； 人將被殺，你須攔阻。
PROV|24|12|你若說：「看哪，這事我們不知道」， 那衡量人心的豈不明白嗎？ 保護你性命的豈不知道嗎？ 他豈不按各人所做的報應各人嗎？
PROV|24|13|我兒啊，你要吃蜜，因為它是美好的， 要讓甘甜的蜜滴入你的口。
PROV|24|14|你要知道，智慧對你的生命正像如此。 你若找著，必有前途， 你的指望也不致斷絕。
PROV|24|15|你這惡人，不可埋伏攻擊義人的家， 也不可毀壞他安居之所。
PROV|24|16|因為義人雖七次跌倒，仍必興起； 惡人卻被禍患傾倒。
PROV|24|17|你的仇敵跌倒，你不要歡喜， 他傾倒，你的心不要快樂；
PROV|24|18|恐怕耶和華看見就不喜悅， 將怒氣從仇敵身上轉過來。
PROV|24|19|不要為作惡的心懷不平， 也不要嫉妒惡人，
PROV|24|20|因為壞人沒有前途， 惡人的燈也必熄滅。
PROV|24|21|我兒啊，你要敬畏耶和華與君王， 不可結交反覆無常的人，
PROV|24|22|因為他們的災難必忽然興起。 誰能知道耶和華與君王所施行的毀滅呢？
PROV|24|23|以下也是智慧人的箴言： 審判時看人情面是不好的。
PROV|24|24|對惡人說「你是義人」的， 萬民必詛咒，萬族必惱恨。
PROV|24|25|責備惡人的，必得喜悅， 美好的福分也必臨到他。
PROV|24|26|應對合宜的， 猶如與人親吻。
PROV|24|27|你要在外面預備材料， 在田間為自己準備齊全， 然後才建造你的房屋。
PROV|24|28|不可無故作證反對鄰舍， 也不可用嘴唇欺騙人。
PROV|24|29|不可說：「人怎樣待我，我也怎樣待他， 我必照他所做的報復他。」
PROV|24|30|我經過懶惰人的田地， 走過無知人的葡萄園，
PROV|24|31|看哪，它長滿了荊棘， 蕁麻蓋地面， 石牆也坍塌了。
PROV|24|32|我看見就留心思想， 我看著就領受訓誨。
PROV|24|33|再睡片時，打盹片時， 抱著雙臂躺臥片時，
PROV|24|34|你的貧窮就如盜賊來到， 你的貧乏彷彿拿盾牌的人來臨。
PROV|25|1|以下也是 所羅門 的箴言，是 猶大 王 希西家 的人所謄錄的。
PROV|25|2|隱藏事情是上帝的榮耀； 查明事情乃君王的榮耀。
PROV|25|3|天之高，地之深， 君王之心測不透。
PROV|25|4|除去銀子的渣滓， 銀匠就做出器皿來。
PROV|25|5|除去王面前的惡人， 國位就靠公義堅立。
PROV|25|6|不可在君王面前妄自尊大， 也不要站在大人的位上。
PROV|25|7|寧可讓人家說「請你上到這裏來」， 強如在你覲見的貴人面前令你退下。
PROV|25|8|不要冒失出去與人爭訟 ， 免得你的鄰舍羞辱你， 最後你就不知怎麼做。
PROV|25|9|要與鄰舍爭辯你的案情， 不可洩漏他人的隱密，
PROV|25|10|恐怕聽見的人責罵你， 你就難以擺脫臭名。
PROV|25|11|一句話說得合宜， 就如金蘋果在銀網子裏
PROV|25|12|智慧人的勸戒在順從的人耳中， 好像金環和金首飾。
PROV|25|13|忠信的使者對那差他的人， 就如收割時有冰雪的涼氣， 使主人的心舒暢。
PROV|25|14|人空誇禮物而不肯贈送， 就好像有風有雲卻無雨。
PROV|25|15|恆常的忍耐可以勸服君王， 柔和的舌頭能折斷骨頭。
PROV|25|16|你得了蜜，吃夠就好， 免得過飽就吐出來。
PROV|25|17|你的腳要少進鄰舍的家， 免得他厭煩你，恨惡你。
PROV|25|18|作假見證陷害鄰舍的， 就是大錘，是利刀，是快箭。
PROV|25|19|患難時倚靠奸詐的人， 好像牙齒斷裂，又如腳脫臼。
PROV|25|20|對傷心的人唱歌， 就如冷天脫他的衣服， 又如在鹼上倒醋 。
PROV|25|21|你的仇敵若餓了，就給他飯吃， 若渴了，就給他水喝；
PROV|25|22|因為你這樣做，就是把炭火堆在他的頭上， 耶和華必回報你。
PROV|25|23|正如北風生雨， 毀謗的舌頭也生怒容。
PROV|25|24|寧可住在房頂的一角， 也不與好爭吵的婦人同住。
PROV|25|25|有好消息從遙遠的地方來， 就如涼水滋潤口渴的人。
PROV|25|26|義人在惡人面前退縮， 好像攪渾之泉，污染之井。
PROV|25|27|吃蜜過多是不好的， 自求榮耀也是一樣。
PROV|25|28|人不克制自己的心， 就像毀壞的城沒有牆。
PROV|26|1|愚昧人得尊榮不相宜， 正如夏天落雪，收割時下雨。
PROV|26|2|詛咒不會無故臨到 ， 正如麻雀掠過，燕子翻飛。
PROV|26|3|鞭子是為打馬，轡頭是為勒驢， 刑杖正是為打愚昧人的背。
PROV|26|4|不要照愚昧人的愚昧話回答他， 免得你與他一樣。
PROV|26|5|要照愚昧人的愚昧話回答他， 免得他自以為有智慧。
PROV|26|6|藉愚昧人的手寄信的， 就像砍斷雙腳，喝下殘暴。
PROV|26|7|箴言在愚昧人的口中， 正如瘸子的腳懸空無用。
PROV|26|8|將尊榮給愚昧人的， 就像石頭綁在彈弓上。
PROV|26|9|箴言在愚昧人的口中， 好像荊棘刺入醉漢的手。
PROV|26|10|雇愚昧人的，與雇過路人的， 就像弓箭手射傷任何人。
PROV|26|11|愚昧人重複做愚昧之事， 就如狗轉過來吃自己所吐的。
PROV|26|12|你看見自以為有智慧的人嗎？ 愚昧人比他更有指望。
PROV|26|13|懶惰人說：「道路有猛獅， 街上有壯獅。」
PROV|26|14|懶惰人在床上， 就像門在軸心上轉動一樣。
PROV|26|15|懶惰人把手埋入盤裏， 就是送進口中也覺得累。
PROV|26|16|懶惰人眼看自己 比七個善於應對的人更有智慧。
PROV|26|17|過路時捲入與己無關的紛爭， 好像人揪住狗耳一般。
PROV|26|18|人欺騙鄰舍，卻說 「我只是開玩笑而已」， 他就像瘋狂的人拋擲致死的火把和利箭。
PROV|26|19|
PROV|26|20|火缺了柴就必熄滅； 無人造謠，紛爭就止息。
PROV|26|21|好爭吵的人煽動爭端， 就如餘火加炭，火上加柴一樣。
PROV|26|22|造謠者的話如同美食， 深入人的肚腹。
PROV|26|23|火熱的 嘴唇，邪惡的心， 好像銀渣包在瓦器上。
PROV|26|24|仇敵用嘴唇掩飾， 心裏卻藏著詭詐；
PROV|26|25|他用甜言蜜語，你不能相信他， 因為他心中有七樣可憎惡的事。
PROV|26|26|他雖用詭詐掩飾怨恨， 他的邪惡必在集會中顯露。
PROV|26|27|挖陷坑的，自己必陷在其中； 滾石頭的，石頭反滾在他身上。
PROV|26|28|虛謊的舌憎恨他所壓傷的人； 諂媚的口敗壞人的事。
PROV|27|1|不要為明天自誇， 因為你不知道每天會發生何事。
PROV|27|2|要讓陌生人誇獎你，不可用口自誇； 讓外邦人稱讚你，不可用嘴唇稱讚自己。
PROV|27|3|石頭沉，沙土重， 愚妄人的惱怒比這兩樣更沉重。
PROV|27|4|憤怒為殘忍，怒氣像狂瀾， 惟有嫉妒，誰能擋得住呢？
PROV|27|5|當面的責備 勝過隱藏的愛情。
PROV|27|6|朋友加的傷痕出於忠誠； 敵人的親吻卻是多餘。
PROV|27|7|人吃飽了，厭惡蜂房的蜜； 人飢餓了，一切苦物都覺甘甜。
PROV|27|8|人離故鄉漂泊， 就像雀鳥離窩四處飛翔。
PROV|27|9|膏油與香料使人心喜悅， 朋友誠心的勸勉也是如此甘美。
PROV|27|10|你的朋友和父親的朋友， 你都不可離棄。 你遭難時，不要上兄弟的家去； 相近的鄰舍強如遠方的兄弟。
PROV|27|11|我兒啊，你要做智慧人，好叫我的心歡喜， 使我可以回答那辱罵我的人。
PROV|27|12|通達人見禍就藏躲； 愚蒙人卻前往受害。
PROV|27|13|誰為陌生人擔保，就拿誰的衣服； 誰為外邦女子作保，誰就要承當。
PROV|27|14|清晨起來大聲給朋友祝福的， 就算是詛咒他。
PROV|27|15|下雨天連連滴漏， 好爭吵的婦人就像這樣；
PROV|27|16|攔阻她的，就是攔阻風， 又像用右手抓油。
PROV|27|17|以鐵磨鐵，越磨越利， 朋友當面琢磨，也是如此。
PROV|27|18|看守無花果樹的，必吃樹上的果子； 敬奉主人的，必得尊榮。
PROV|27|19|水中照臉，彼此相符； 人心相映，也是如此。
PROV|27|20|陰間和冥府 永不滿足， 人的眼目也是如此。
PROV|27|21|鼎為煉銀，爐為煉金， 口中的稱讚也試煉人。
PROV|27|22|用杵把愚妄人與穀粒一同搗在臼中， 他的愚昧還是離不了他。
PROV|27|23|你要詳細知道你羊群的景況， 留心照顧你的牛群，
PROV|27|24|因為財富不能永留， 冠冕豈能存到萬代？
PROV|27|25|青草除去，嫩草長出， 山上的菜蔬也被採收。
PROV|27|26|綿羊可以做衣服， 公山羊可作田地的價值，
PROV|27|27|並有母山羊奶夠你吃， 夠你養家和女僕的生活。
PROV|28|1|惡人雖無人追趕也逃跑； 義人卻膽壯像獅子。
PROV|28|2|地上因有罪過，君王就多更換； 因聰明和有見識的人，國必長存。
PROV|28|3|窮乏人欺壓貧寒人， 好像暴雨掃過，不留糧食。
PROV|28|4|離棄律法的，誇獎惡人； 遵守律法的，卻與惡人相爭。
PROV|28|5|惡人不明白公義； 惟有尋求耶和華的，無不明白。
PROV|28|6|行為純正的窮乏人 勝過行事歪曲的有錢人。
PROV|28|7|謹守教誨的，是聰明之子； 與貪食者為伍的，卻羞辱其父。
PROV|28|8|人以厚利增加財富， 是給那憐憫貧寒人的積財。
PROV|28|9|轉耳不聽教誨的， 他的祈禱也可憎。
PROV|28|10|誘惑正直人行惡道的，必掉在自己的坑裏； 惟有完全人必承受福分。
PROV|28|11|有錢人自以為有智慧， 但聰明的貧寒人能看穿他。
PROV|28|12|義人高升，有大榮耀； 惡人興起，人就躲藏。
PROV|28|13|遮掩自己過犯的，必不順利； 承認且離棄過犯的，必蒙憐憫。
PROV|28|14|常存敬畏的，這人有福了； 心裏剛硬的，必陷在禍患裏。
PROV|28|15|邪惡的君王壓制貧民， 好像吼叫的獅子，又如覓食的熊。
PROV|28|16|無知的君王多行暴虐； 恨惡非分之財的，必年長日久。
PROV|28|17|背負流人血之罪的，必逃跑直到地府； 願無人幫助他！
PROV|28|18|行為正直的，必蒙拯救； 行事彎曲的，立時跌倒。
PROV|28|19|耕種自己田地的，糧食充足； 追求虛浮的，窮困潦倒。
PROV|28|20|誠實人必多得福； 想要急速發財的，難免受罰。
PROV|28|21|看人情面是不好的； 卻有人因一塊餅而犯法。
PROV|28|22|守財奴 想要急速發財， 卻不知窮乏必臨到他身上。
PROV|28|23|責備人的，後來蒙人喜悅， 多於那用舌頭諂媚人的。
PROV|28|24|搶奪父母竟說「這不是罪過」， 此人與毀滅者同類。
PROV|28|25|心中貪婪的，挑起爭端； 倚靠耶和華的，必得豐裕。
PROV|28|26|心中自以為是的，就是愚昧人； 憑智慧行事的，必蒙拯救。
PROV|28|27|賙濟窮乏人的，不致缺乏； 遮眼不看的，多受詛咒。
PROV|28|28|惡人興起，人就躲藏； 惡人敗亡，義人必增多。
PROV|29|1|人屢次受責罰，仍然硬著頸項， 他必頃刻被毀，無從醫治。
PROV|29|2|義人增多，民就喜樂； 惡人掌權，民就嘆息。
PROV|29|3|愛慕智慧的，使父親喜樂； 結交妓女的，卻浪費錢財。
PROV|29|4|王藉公平，使國堅定； 強索貢物的，使它毀壞。
PROV|29|5|諂媚鄰舍的， 就是設網羅絆他的腳。
PROV|29|6|惡人犯罪，自陷圈套； 惟獨義人歡呼喜樂。
PROV|29|7|義人關注貧寒人的案情； 惡人不明瞭這種知識。
PROV|29|8|傲慢人煽動全城； 智慧人止息眾怒。
PROV|29|9|智慧人與愚妄人有爭訟， 或怒或笑，總不得安寧。
PROV|29|10|好流人血的，恨惡完全人， 正直人卻顧惜 他的性命。
PROV|29|11|愚昧人怒氣全發； 智慧人自我平息。
PROV|29|12|君王若聽謊言， 他一切臣僕都是奸惡。
PROV|29|13|窮乏人和欺壓者相遇 ， 耶和華使他們的眼目明亮。
PROV|29|14|君王憑誠信判斷貧寒人， 他的國位必永遠堅立。
PROV|29|15|杖打和責備能增加智慧； 任性的少年使母親羞愧。
PROV|29|16|惡人多，過犯也加多， 義人必看見他們敗亡。
PROV|29|17|管教你的兒子，他就使你得安寧， 也使你心裏喜樂。
PROV|29|18|沒有異象 ，民就放肆； 惟遵守律法的，便為有福。
PROV|29|19|僕人不能靠言語受教； 他即使明白，也不回應。
PROV|29|20|你見過言語急躁的人嗎？ 愚昧人比他更有指望。
PROV|29|21|人將僕人從小嬌養， 至終必帶來憂傷 。
PROV|29|22|好生氣的人挑起爭端， 暴怒的人多多犯錯。
PROV|29|23|人的高傲使自己蒙羞； 心裏謙遜的，必得尊榮。
PROV|29|24|與盜賊分贓的，是恨惡自己的性命； 他雖聽見發誓的聲音，也不告訴人。
PROV|29|25|懼怕人的，陷入圈套； 惟有倚靠耶和華的，必得安穩。
PROV|29|26|求王恩的人多； 人獲公正來自耶和華。
PROV|29|27|不義之人，義人憎惡； 行事正直的，惡人憎惡。
PROV|30|1|雅基 的兒子、 瑪撒 人 亞古珥 的言語 ，是這人對 以鐵 和 烏甲 說的。
PROV|30|2|我比眾人更像畜牲， 也沒有人的聰明。
PROV|30|3|我沒有學好智慧， 也不認識至聖者。
PROV|30|4|誰升天又降下來？ 誰聚風在手掌中？ 誰包水在衣服裏？ 誰立定地的四極？ 他名叫甚麼？ 他兒子名叫甚麼？ 你知道嗎？
PROV|30|5|上帝的言語句句都是煉淨的， 投靠他的，他便作他們的盾牌。
PROV|30|6|你不可加添他的言語， 恐怕他責備你，你就顯為說謊的。
PROV|30|7|我求你兩件事， 在我未死之先，不要拒絕我：
PROV|30|8|求你使虛假和謊言遠離我， 使我不貧窮也不富足， 賜給我需用的飲食。
PROV|30|9|免得我飽足了，就不認你，說： 「耶和華是誰呢？」 又恐怕我貧窮就偷竊， 以致褻瀆我上帝的名。
PROV|30|10|不要向主人讒害他的僕人， 恐怕他詛咒你，你便算為有罪。
PROV|30|11|有一類人，詛咒父親， 不給母親祝福。
PROV|30|12|有一類人，自以為純潔， 卻沒有洗淨自己的污穢。
PROV|30|13|有一類人，眼目何其高傲， 眼皮也是高舉。
PROV|30|14|有一類人，牙如劍，齒如刀， 要吞滅地上的困苦人和世間的貧窮人。
PROV|30|15|水蛭有兩個女兒： 「給呀，給呀。」 有三樣不知足的， 不說「夠了」的有四樣：
PROV|30|16|陰間和不生育的子宮， 吸水不足的地，還有不說「夠了」的火。
PROV|30|17|嘲笑父親、藐視而不聽從母親的， 谷中的烏鴉必啄他的眼睛，小鷹也必吃它。
PROV|30|18|我所測不透的奇妙有三樣， 我所不知道的有四樣：
PROV|30|19|就是鷹在空中飛的道， 蛇在磐石上爬的道， 船在海中行的道， 男與女交合的道。
PROV|30|20|淫婦的道是這樣， 她吃了，把嘴一擦就說： 「我沒有行惡。」
PROV|30|21|使地震動的有三樣， 地承擔不起的有四樣：
PROV|30|22|就是僕人作王， 愚頑人吃得飽足，
PROV|30|23|令人憎惡的女子出嫁， 婢女取代她的女主人。
PROV|30|24|地上有四樣東西雖小，卻甚聰明：
PROV|30|25|螞蟻是無力之類， 卻在夏天預備糧食。
PROV|30|26|石獾並非強壯之類， 卻在巖石中造房子。
PROV|30|27|蝗蟲沒有君王， 卻分隊而出。
PROV|30|28|壁虎你用手就可抓住， 牠卻住在王宮。
PROV|30|29|腳步威武的有三樣， 行走威武的有四樣：
PROV|30|30|獅子－百獸中最勇猛的、 無論遇見甚麼絕不退縮，
PROV|30|31|獵狗，公山羊， 和有整排士兵的君王。
PROV|30|32|你若行事愚頑，自高自傲， 或是設計惡謀，就當用手摀口。
PROV|30|33|攪動牛奶必成乳酪， 扭鼻子必出血， 照樣，激發烈怒必挑起爭端。
PROV|31|1|瑪撒 王 利慕伊勒 的言語，就是他母親教導他的 。
PROV|31|2|我兒，怎麼了？ 我腹中生的兒，怎麼了？ 我許願而得的兒，怎麼了？
PROV|31|3|不要將你的精力給婦女， 也不要有敗壞君王的行為。
PROV|31|4|利慕伊勒 啊，君王不宜，君王不宜喝酒， 王子尋找烈酒也不相宜；
PROV|31|5|恐怕喝了就忘記所頒的法令， 顛倒所有困苦人的是非。
PROV|31|6|可以把烈酒給將亡的人喝， 把酒給心裏愁苦的人喝，
PROV|31|7|讓他喝了，就忘記他的貧窮， 不再記得他的苦楚。
PROV|31|8|你當為不能自辯的人 開口， 為所有孤獨無助者伸冤。
PROV|31|9|你當開口按公義判斷， 當為困苦和貧窮的人辯護。
PROV|31|10|才德的婦人誰能得著呢？ 她的價值遠勝過寶石。
PROV|31|11|她丈夫心裏信賴她， 必不缺少利益；
PROV|31|12|她終其一生， 使丈夫有益無損。
PROV|31|13|她尋找羊毛和麻， 歡喜用手做工。
PROV|31|14|她好像商船， 從遠方運來糧食，
PROV|31|15|未到黎明她就起來， 把食物分給家中的人， 將當做的工分派女僕。
PROV|31|16|她想得田地，就去買來， 用手中的成果栽葡萄園。
PROV|31|17|她以能力束腰， 使膀臂有力。
PROV|31|18|她覺得自己獲利不錯， 她的燈終夜不滅。
PROV|31|19|她伸手拿捲線桿， 她的手掌把住紡車。
PROV|31|20|她張手賙濟困苦人， 伸手幫助貧窮人。
PROV|31|21|她不因下雪為家裏的人擔心， 因為全家都穿上朱紅衣服。
PROV|31|22|她為自己製作被單， 她的衣服是細麻和紫色布做的。
PROV|31|23|她丈夫在城門口與本地的長老同坐， 為人所認識。
PROV|31|24|她做細麻布衣裳來賣， 又將腰帶賣給商家。
PROV|31|25|能力和威儀是她的衣服， 她想到日後的景況就喜笑。
PROV|31|26|她開口就發智慧， 她舌上有仁慈的教誨。
PROV|31|27|她管理家務， 並不吃閒飯。
PROV|31|28|她的兒女起來稱她有福， 她的丈夫也稱讚她：
PROV|31|29|「才德的女子很多， 惟獨你超過一切。」
PROV|31|30|魅力是虛假的，美貌是虛浮的； 惟敬畏耶和華的婦女必得稱讚。
PROV|31|31|她手中的成果你們要賞給她， 願她的工作在城門口榮耀她。
