2TIM|1|1|Paulus apostolus Christi Iesu per voluntatem Dei secundum promissionem vitae quae est in Christo Iesu
2TIM|1|2|Timotheo carissimo filio gratia misericordia pax a Deo Patre et Christo Iesu Domino nostro
2TIM|1|3|gratias ago Deo cui servio a progenitoribus in conscientia pura quam sine intermissione habeam tui memoriam in orationibus meis nocte ac die
2TIM|1|4|desiderans te videre memor lacrimarum tuarum ut gaudio implear
2TIM|1|5|recordationem accipiens eius fidei quae est in te non ficta quae et habitavit primum in avia tua Loide et matre tua Eunice certus sum autem quod et in te
2TIM|1|6|propter quam causam admoneo te ut resuscites gratiam Dei quae est in te per inpositionem manuum mearum
2TIM|1|7|non enim dedit nobis Deus spiritum timoris sed virtutis et dilectionis et sobrietatis
2TIM|1|8|noli itaque erubescere testimonium Domini nostri neque me vinctum eius sed conlabora evangelio secundum virtutem Dei
2TIM|1|9|qui nos liberavit et vocavit vocatione sancta non secundum opera nostra sed secundum propositum suum et gratiam quae data est nobis in Christo Iesu ante tempora saecularia
2TIM|1|10|manifestata est autem nunc per inluminationem salvatoris nostri Iesu Christi qui destruxit quidem mortem inluminavit autem vitam et incorruptionem per evangelium
2TIM|1|11|in quo positus sum ego praedicator et apostolus et magister gentium
2TIM|1|12|ob quam causam etiam haec patior sed non confundor scio enim cui credidi et certus sum quia potens est depositum meum servare in illum diem
2TIM|1|13|formam habe sanorum verborum quae a me audisti in fide et dilectione in Christo Iesu
2TIM|1|14|bonum depositum custodi per Spiritum Sanctum qui habitat in nobis
2TIM|1|15|scis hoc quod aversi sunt a me omnes qui in Asia sunt ex quibus est Phygelus et Hermogenes
2TIM|1|16|det misericordiam Dominus Onesifori domui quia saepe me refrigeravit et catenam meam non erubuit
2TIM|1|17|sed cum Romam venisset sollicite me quaesivit et invenit
2TIM|1|18|det illi Dominus invenire misericordiam a Domino in illa die et quanta Ephesi ministravit melius tu nosti
2TIM|2|1|tu ergo fili mi confortare in gratia quae est in Christo Iesu
2TIM|2|2|et quae audisti a me per multos testes haec commenda fidelibus hominibus qui idonei erunt et alios docere
2TIM|2|3|labora sicut bonus miles Christi Iesu
2TIM|2|4|nemo militans inplicat se negotiis saecularibus ut ei placeat cui se probavit
2TIM|2|5|nam et qui certat in agone non coronatur nisi legitime certaverit
2TIM|2|6|laborantem agricolam oportet primum de fructibus accipere
2TIM|2|7|intellege quae dico dabit enim tibi Dominus in omnibus intellectum
2TIM|2|8|memor esto Iesum Christum resurrexisse a mortuis ex semine David secundum evangelium meum
2TIM|2|9|in quo laboro usque ad vincula quasi male operans sed verbum Dei non est alligatum
2TIM|2|10|ideo omnia sustineo propter electos ut et ipsi salutem consequantur quae est in Christo Iesu cum gloria caelesti
2TIM|2|11|fidelis sermo nam si conmortui sumus et convivemus
2TIM|2|12|si sustinemus et conregnabimus si negabimus et ille negabit nos
2TIM|2|13|si non credimus ille fidelis manet negare se ipsum non potest
2TIM|2|14|haec commone testificans coram Domino noli verbis contendere in nihil utile ad subversionem audientium
2TIM|2|15|sollicite cura te ipsum probabilem exhibere Deo operarium inconfusibilem recte tractantem verbum veritatis
2TIM|2|16|profana autem inaniloquia devita multum enim proficient ad impietatem
2TIM|2|17|et sermo eorum ut cancer serpit ex quibus est Hymeneus et Philetus
2TIM|2|18|qui a veritate exciderunt dicentes resurrectionem iam factam et subvertunt quorundam fidem
2TIM|2|19|sed firmum fundamentum Dei stetit habens signaculum hoc cognovit Dominus qui sunt eius et discedat ab iniquitate omnis qui nominat nomen Domini
2TIM|2|20|in magna autem domo non solum sunt vasa aurea et argentea sed et lignea et fictilia et quaedam quidem in honorem quaedam autem in contumeliam
2TIM|2|21|si quis ergo emundaverit se ab istis erit vas in honorem sanctificatum et utile Domino ad omne opus bonum paratum
2TIM|2|22|iuvenilia autem desideria fuge sectare vero iustitiam fidem caritatem pacem cum his qui invocant Dominum de corde puro
2TIM|2|23|stultas autem et sine disciplina quaestiones devita sciens quia generant lites
2TIM|2|24|servum autem Domini non oportet litigare sed mansuetum esse ad omnes docibilem patientem
2TIM|2|25|cum modestia corripientem eos qui resistunt nequando det illis Deus paenitentiam ad cognoscendam veritatem
2TIM|2|26|et resipiscant a diaboli laqueis a quo capti tenentur ad ipsius voluntatem
2TIM|3|1|hoc autem scito quod in novissimis diebus instabunt tempora periculosa
2TIM|3|2|et erunt homines se ipsos amantes cupidi elati superbi blasphemi parentibus inoboedientes ingrati scelesti
2TIM|3|3|sine affectione sine pace criminatores incontinentes inmites sine benignitate
2TIM|3|4|proditores protervi tumidi voluptatium amatores magis quam Dei
2TIM|3|5|habentes speciem quidem pietatis virtutem autem eius abnegantes et hos devita
2TIM|3|6|ex his enim sunt qui penetrant domos et captivas ducunt mulierculas oneratas peccatis quae ducuntur variis desideriis
2TIM|3|7|semper discentes et numquam ad scientiam veritatis pervenientes
2TIM|3|8|quemadmodum autem Iannes et Mambres restiterunt Mosi ita et hii resistunt veritati homines corrupti mente reprobi circa fidem
2TIM|3|9|sed ultra non proficient insipientia enim eorum manifesta erit omnibus sicut et illorum fuit
2TIM|3|10|tu autem adsecutus es meam doctrinam institutionem propositum fidem longanimitatem dilectionem patientiam
2TIM|3|11|persecutiones passiones qualia mihi facta sunt Antiochiae Iconii Lystris quales persecutiones sustinui et ex omnibus me eripuit Dominus
2TIM|3|12|et omnes qui volunt pie vivere in Christo Iesu persecutionem patientur
2TIM|3|13|mali autem homines et seductores proficient in peius errantes et in errorem mittentes
2TIM|3|14|tu vero permane in his quae didicisti et credita sunt tibi sciens a quo didiceris
2TIM|3|15|et quia ab infantia sacras litteras nosti quae te possint instruere ad salutem per fidem quae est in Christo Iesu
2TIM|3|16|omnis scriptura divinitus inspirata et utilis ad docendum ad arguendum ad corrigendum ad erudiendum in iustitia
2TIM|3|17|ut perfectus sit homo Dei ad omne opus bonum instructus
2TIM|4|1|testificor coram Deo et Christo Iesu qui iudicaturus est vivos ac mortuos et adventum ipsius et regnum eius
2TIM|4|2|praedica verbum insta oportune inportune argue obsecra increpa in omni patientia et doctrina
2TIM|4|3|erit enim tempus cum sanam doctrinam non sustinebunt sed ad sua desideria coacervabunt sibi magistros prurientes auribus
2TIM|4|4|et a veritate quidem auditum avertent ad fabulas autem convertentur
2TIM|4|5|tu vero vigila in omnibus labora opus fac evangelistae ministerium tuum imple
2TIM|4|6|ego enim iam delibor et tempus meae resolutionis instat
2TIM|4|7|bonum certamen certavi cursum consummavi fidem servavi
2TIM|4|8|in reliquo reposita est mihi iustitiae corona quam reddet mihi Dominus in illa die iustus iudex non solum autem mihi sed et his qui diligunt adventum eius
2TIM|4|9|festina venire ad me cito
2TIM|4|10|Demas enim me dereliquit diligens hoc saeculum et abiit Thessalonicam Crescens in Galliam Titus in Dalmatiam
2TIM|4|11|Lucas est mecum solus Marcum adsume et adduc tecum est enim mihi utilis in ministerium
2TIM|4|12|Tychicum autem misi Ephesum
2TIM|4|13|paenulam quam reliqui Troade apud Carpum veniens adfers et libros maxime autem membranas
2TIM|4|14|Alexander aerarius multa mala mihi ostendit reddat ei Dominus secundum opera eius
2TIM|4|15|quem et tu devita valde enim restitit verbis nostris
2TIM|4|16|in prima mea defensione nemo mihi adfuit sed omnes me dereliquerunt non illis reputetur
2TIM|4|17|Dominus autem mihi adstitit et confortavit me ut per me praedicatio impleatur et audiant omnes gentes et liberatus sum de ore leonis
2TIM|4|18|liberabit me Dominus ab omni opere malo et salvum faciet in regnum suum caeleste cui gloria in saecula saeculorum amen
2TIM|4|19|saluta Priscam et Aquilam et Onesifori domum
2TIM|4|20|Erastus remansit Corinthi Trophimum autem reliqui infirmum Mileti
2TIM|4|21|festina ante hiemem venire salutat te Eubulus et Pudens et Linus et Claudia et fratres omnes
2TIM|4|22|Dominus Iesus cum spiritu tuo gratia nobiscum amen
