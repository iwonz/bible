EZRA|1|1|В первый год Кира, царя Персидского, во исполнение слова Господня из уст Иеремии, возбудил Господь дух Кира, царя Персидского, и он повелел объявить по всему царству своему, словесно и письменно:
EZRA|1|2|так говорит Кир, царь Персидский: все царства земли дал мне Господь Бог небесный, и Он повелел мне построить Ему дом в Иерусалиме, что в Иудее.
EZRA|1|3|Кто есть из вас, из всего народа Его, – да будет Бог его с ним, – и пусть он идет в Иерусалим, что в Иудее, и строит дом Господа Бога Израилева, Того Бога, Который в Иерусалиме.
EZRA|1|4|А все оставшиеся во всех местах, где бы тот ни жил, пусть помогут ему жители места того серебром и золотом и [иным] имуществом, и скотом, с доброхотным даянием для дома Божия, что в Иерусалиме.
EZRA|1|5|И поднялись главы поколений Иудиных и Вениаминовых, и священники и левиты, всякий, [в ком] возбудил Бог дух его, чтобы пойти строить дом Господень, который в Иерусалиме.
EZRA|1|6|И все соседи их вспомоществовали им серебряными сосудами, золотом, [иным] имуществом, и скотом, и дорогими вещами, сверх всякого доброхотного даяния [для храма].
EZRA|1|7|И царь Кир вынес сосуды дома Господня, которые Навуходоносор взял из Иерусалима и положил в доме бога своего, –
EZRA|1|8|и вынес их Кир, царь Персидский, рукою Мифредата сокровищехранителя, а он счетом сдал их Шешбацару князю Иудину.
EZRA|1|9|И вот число их: блюд золотых тридцать, блюд серебряных тысяча, ножей двадцать девять,
EZRA|1|10|чаш золотых тридцать, чаш серебряных двойных четыреста десять, других сосудов тысяча:
EZRA|1|11|всех сосудов, золотых и серебряных, пять тысяч четыреста. Все [это] взял [с собою] Шешбацар, при отправлении переселенцев из Вавилона в Иерусалим.
EZRA|2|1|Вот сыны страны из пленников переселения, которых Навуходоносор, царь Вавилонский, отвел в Вавилон, возвратившиеся в Иерусалим и Иудею, каждый в свой город, –
EZRA|2|2|пришедшие с Зоровавелем, Иисусом, Неемиею, Сараием, Реелаем, Мардохеем, Билшаном, Мисфаром, Бигваем, Рехумом, Вааном. Число людей народа Израилева:
EZRA|2|3|сыновей Пароша две тысячи сто семьдесят два;
EZRA|2|4|сыновей Сафатии триста семьдесят два;
EZRA|2|5|сыновей Араха семьсот семьдесят пять;
EZRA|2|6|сыновей Пахаф–Моава, из сыновей Иисуса [и] Иоава, две тысячи восемьсот двенадцать;
EZRA|2|7|сыновей Елама тысяча двести пятьдесят четыре;
EZRA|2|8|сыновей Заттуя девятьсот сорок пять;
EZRA|2|9|сыновей Закхая семьсот шестьдесят;
EZRA|2|10|сыновей Вания шестьсот сорок два;
EZRA|2|11|сыновей Бебая шестьсот двадцать три;
EZRA|2|12|сыновей Азгада тысяча двести двадцать два;
EZRA|2|13|сыновей Адоникама шестьсот шестьдесят шесть;
EZRA|2|14|сыновей Бигвая две тысячи пятьдесят шесть;
EZRA|2|15|сыновей Адина четыреста пятьдесят четыре;
EZRA|2|16|сыновей Атера, из [дома] Езекии, девяносто восемь;
EZRA|2|17|сыновей Бецая триста двадцать три;
EZRA|2|18|сыновей Иоры сто двенадцать;
EZRA|2|19|сыновей Хашума двести двадцать три;
EZRA|2|20|сыновей Гиббара девяносто пять;
EZRA|2|21|уроженцев Вифлеема сто двадцать три;
EZRA|2|22|жителей Нетофы пятьдесят шесть;
EZRA|2|23|жителей Анафофа сто двадцать восемь;
EZRA|2|24|уроженцев Азмавефа сорок два;
EZRA|2|25|уроженцев Кириаф–Иарима, Кефиры и Беерофа семьсот сорок три;
EZRA|2|26|уроженцев Рамы и Гевы шестьсот двадцать один;
EZRA|2|27|жителей Михмаса сто двадцать два;
EZRA|2|28|жителей Вефиля и Гая двести двадцать три;
EZRA|2|29|уроженцев Нево пятьдесят два;
EZRA|2|30|уроженцев Магбиша сто пятьдесят шесть;
EZRA|2|31|сыновей другого Елама тысяча двести пятьдесят четыре;
EZRA|2|32|сыновей Харима триста двадцать;
EZRA|2|33|уроженцев Лидды, Хадида и Оно семьсот двадцать пять;
EZRA|2|34|уроженцев Иерихона триста сорок пять;
EZRA|2|35|уроженцев Сенаи три тысячи шестьсот тридцать.
EZRA|2|36|Священников: сыновей Иедаии, из дома Иисусова, девятьсот семьдесят три;
EZRA|2|37|сыновей Иммера тысяча пятьдесят два;
EZRA|2|38|сыновей Пашхура тысяча двести сорок семь;
EZRA|2|39|сыновей Харима тысяча семнадцать.
EZRA|2|40|Левитов: сыновей Иисуса и Кадмиила, из сыновей Годавии, семьдесят четыре;
EZRA|2|41|певцов: сыновей Асафа сто двадцать восемь;
EZRA|2|42|сыновей привратников: сыновья Шаллума, сыновья Атера, сыновья Талмона, сыновья Аккува, сыновья Хатиты, сыновья Шовая, – всего сто тридцать девять.
EZRA|2|43|Нефинеев: сыновья Цихи, сыновья Хасуфы, сыновья Таббаофа,
EZRA|2|44|сыновья Кероса, сыновья Сиаги, сыновья Фадона,
EZRA|2|45|сыновья Лебаны, сыновья Хагабы, сыновья Аккува,
EZRA|2|46|сыновья Хагава, сыновья Шамлая, сыновья Ханана,
EZRA|2|47|сыновья Гиддела, сыновья Гахара, сыновья Реаии,
EZRA|2|48|сыновья Рецина, сыновья Некоды, сыновья Газзама,
EZRA|2|49|сыновья Уззы, сыновья Пасеаха, сыновья Бесая,
EZRA|2|50|сыновья Асны, сыновья Меунима, сыновья Нефисима,
EZRA|2|51|сыновья Бакбука, сыновья Хакуфы, сыновья Хархура,
EZRA|2|52|сыновья Бацлуфа, сыновья Мехиды, сыновья Харши,
EZRA|2|53|сыновья Баркоса, сыновья Сисры, сыновья Фамаха,
EZRA|2|54|сыновья Нециаха, сыновья Хатифы;
EZRA|2|55|сыновья рабов Соломоновых: сыновья Сотая, сыновья Гассоферефа, сыновья Феруды,
EZRA|2|56|сыновья Иаалы, сыновья Даркона, сыновья Гиддела,
EZRA|2|57|сыновья Сефатии, сыновья Хаттила, сыновья Похереф–Гаццебайима, сыновья Амия, –
EZRA|2|58|всего – нефинеев и сыновей рабов Соломоновых триста девяносто два.
EZRA|2|59|И вот вышедшие из Тел–Мелаха, Тел–Харши, Херуб–Аддан–Иммера, которые не могли показать о поколении своем и о племени своем – от Израиля ли они:
EZRA|2|60|сыновья Делайи, сыновья Товии, сыновья Некоды, шестьсот пятьдесят два.
EZRA|2|61|И из сыновей священнических: сыновья Хабайи, сыновья Гаккоца, сыновья Верзеллия, который взял жену из дочерей Верзеллия Галаадитянина и стал называться именем их.
EZRA|2|62|Они искали своей записи родословной, и не нашлось ее, а [потому] исключены из священства.
EZRA|2|63|И Тиршафа сказал им, чтоб они не ели великой святыни, доколе не восстанет священник с уримом и туммимом.
EZRA|2|64|Все общество вместе [состояло] из сорока двух тысяч трехсот шестидесяти [человек],
EZRA|2|65|кроме рабов их и рабынь их, которых [было] семь тысяч триста тридцать семь; и при них певцов и певиц двести.
EZRA|2|66|Коней у них семьсот тридцать шесть, лошаков у них двести сорок пять;
EZRA|2|67|верблюдов у них четыреста тридцать пять, ослов шесть тысяч семьсот двадцать.
EZRA|2|68|Из глав поколений [некоторые], придя к дому Господню, что в Иерусалиме, доброхотно жертвовали на дом Божий, чтобы восстановить его на основании его.
EZRA|2|69|По достатку своему, они дали в сокровищницу на [производство] работ шестьдесят одну тысячу драхм золота и пять тысяч мин серебра и сто священнических одежд.
EZRA|2|70|И стали жить священники и левиты, и народ и певцы, и привратники и нефинеи в городах своих, и весь Израиль в городах своих.
EZRA|3|1|Когда наступил седьмой месяц, и сыны Израилевы [уже были] в городах, тогда собрался народ, как один человек, в Иерусалиме.
EZRA|3|2|И встал Иисус, сын Иоседеков, и братья его священники, и Зоровавель, сын Салафиилов, и братья его, и соорудили они жертвенник Богу Израилеву, чтобы возносить на нем всесожжения, как написано в законе Моисея, человека Божия.
EZRA|3|3|И поставили жертвенник на основании его, так как они [были] в страхе от иноземных народов; и стали возносить на нем всесожжения Господу, всесожжения утренние и вечерние.
EZRA|3|4|И совершили праздник кущей, как предписано, с ежедневным всесожжением в определенном числе, по уставу [каждого] дня.
EZRA|3|5|И после того [совершали] всесожжение постоянное, и в новомесячия, и во все праздники, посвященные Господу, и добровольное приношение Господу от всякого усердствующего.
EZRA|3|6|С первого же дня седьмого месяца начали возносить всесожжения Господу. А храму Господню [еще] не было положено основание.
EZRA|3|7|И стали выдавать серебро каменотесам и плотникам, и пищу и питье и масло Сидонянам и Тирянам, чтоб они доставляли кедровый лес с Ливана по морю в Яфу, с дозволения им Кира, царя Персидского.
EZRA|3|8|Во второй год по приходе своем к дому Божию в Иерусалим, во второй месяц Зоровавель, сын Салафиилов, и Иисус, сын Иоседеков, и прочие братья их, священники и левиты, и все пришедшие из плена в Иерусалим положили начало и поставили левитов от двадцати лет и выше для надзора за работами дома Господня.
EZRA|3|9|И стали Иисус, сыновья его и братья его, Кадмиил и сыновья его, сыновья Иуды, как один [человек], для надзора за производителями работ в доме Божием, [а также и] сыновья Хенадада, сыновья их и братья их левиты.
EZRA|3|10|Когда строители положили основание храму Господню, тогда поставили священников в облачении их с трубами и левитов, сыновей Асафовых, с кимвалами, чтобы славить Господа по уставу Давида, царя Израилева.
EZRA|3|11|И начали они попеременно петь: "хвалите" и: "славьте Господа", "ибо – благ, ибо вовек милость Его к Израилю". И весь народ восклицал громогласно, славя Господа за то, что положено основание дома Господня.
EZRA|3|12|Впрочем многие из священников и левитов и глав поколений, старики, которые видели прежний храм, при основании этого храма пред глазами их, плакали громко, но многие и восклицали от радости громогласно.
EZRA|3|13|И не мог народ распознать восклицаний радости от воплей плача народного, потому что народ восклицал громко, и голос слышен был далеко.
EZRA|4|1|И услышали враги Иуды и Вениамина, что возвратившиеся из плена строят храм Господу Богу Израилеву;
EZRA|4|2|и пришли они к Зоровавелю и к главам поколений, и сказали им: будем и мы строить с вами, потому что мы, как и вы, прибегаем к Богу вашему, и Ему приносим жертвы от дней Асардана, царя Сирийского, который перевел нас сюда.
EZRA|4|3|И сказал им Зоровавель и Иисус и прочие главы поколений Израильских: не строить вам вместе с нами дом нашему Богу; мы одни будем строить [дом] Господу, Богу Израилеву, как повелел нам царь Кир, царь Персидский.
EZRA|4|4|И стал народ земли той ослаблять руки народа Иудейского и препятствовать ему в строении;
EZRA|4|5|и подкупали против них советников, чтобы разрушить предприятие их, во все дни Кира, царя Персидского, и до царствования Дария, царя Персидского.
EZRA|4|6|А в царствование Ахашвероша, в начале царствования его, написали обвинение на жителей Иудеи и Иерусалима.
EZRA|4|7|И во дни Артаксеркса писали Бишлам, Мифредат, Табеел и прочие товарищи их к Артаксерксу, царю Персидскому. Письмо же написано [было] буквами Сирийскими и на Сирийском языке.
EZRA|4|8|Рехум советник и Шимшай писец писали одно письмо против Иерусалима к царю Артаксерксу такое:
EZRA|4|9|Тогда–то. Рехум советник и Шимшай писец и прочие товарищи их, – Динеи и Афарсафхеи, Тарпелеи, Апарсы, Арехьяне, Вавилоняне, Сусанцы, Даги, Еламитяне,
EZRA|4|10|и прочие народы, которых переселил Аснафар, великий и славный и поселил в городах Самарийских и в прочих [городах] за рекою, и прочее.
EZRA|4|11|И вот список с письма, которое послали к нему: Царю Артаксерксу – рабы твои, люди, [живущие] за рекою, и прочее.
EZRA|4|12|Да будет известно царю, что Иудеи, которые вышли от тебя, пришли к нам в Иерусалим, строят [этот] мятежный и негодный город, и стены делают, и основания [их уже] исправили.
EZRA|4|13|Да будет же известно царю, что если этот город будет построен и стены восстановлены, то [ни] подати, [ни] налога, ни пошлины не будут давать, и царской казне сделан будет ущерб.
EZRA|4|14|Так как мы едим соль от дворца царского, и ущерб для царя не можем видеть, поэтому мы посылаем донесение к царю:
EZRA|4|15|пусть поищут в памятной книге отцов твоих, – и найдешь в книге памятной, и узнаешь, что город сей – город мятежный и вредный для царей и областей, и [что] отпадения бывали в нем издавна, за что город сей и опустошен.
EZRA|4|16|Посему мы уведомляем царя, что если город сей будет достроен и стены его доделаны, то после этого не будет у тебя владения за рекою.
EZRA|4|17|Царь послал ответ Рехуму советнику и Шимшаю писцу и прочим товарищам их, которые живут в Самарии и [в] прочих [городах] заречных: Мир... и прочее.
EZRA|4|18|Письмо, которое вы прислали нам, внятно прочитано предо мною;
EZRA|4|19|и от меня дано повеление, – и разыскивали, и нашли, что город этот издавна восставал против царей, и производились в нем мятежи и волнения,
EZRA|4|20|и [что были] в Иерусалиме цари могущественные и владевшие всем заречьем, и им давали подать, налоги и пошлины.
EZRA|4|21|Итак дайте приказание, чтобы люди сии перестали работать, и [чтобы] город сей не строился, доколе от меня не будет дано повеление.
EZRA|4|22|И будьте осторожны, чтобы не сделать в этом недосмотра. К чему допускать размножение вредного в ущерб царям?
EZRA|4|23|Как скоро это письмо царя Артаксеркса было прочитано пред Рехумом и Шимшаем писцом и товарищами их, они немедленно пошли в Иерусалим к Иудеям, и сильною вооруженною рукою остановили работу их.
EZRA|4|24|Тогда остановилась работа при доме Божием, который в Иерусалиме, и остановка сия продолжалась до второго года царствования Дария, царя Персидского.
EZRA|5|1|Но пророк Аггей и пророк Захария, сын Адды, говорили Иудеям, которые в Иудее и Иерусалиме, пророческие речи во имя Бога Израилева.
EZRA|5|2|Тогда встали Зоровавель, сын Салафиилов, и Иисус, сын Иоседеков, и начали строить дом Божий в Иерусалиме, и с ними пророки Божии, подкреплявшие их.
EZRA|5|3|В то время пришел к ним Фафнай, заречный областеначальник, и Шефар–Бознай и товарищи их, и так сказали им: кто дал вам разрешение строить дом сей и доделывать стены сии?
EZRA|5|4|Тогда мы сказали им имена тех людей, которые строят это здание.
EZRA|5|5|Но око Бога их было над старейшинами Иудейскими, и те не возбраняли им, доколе дело не отправили к Дарию, и доколе не пришло решение по этому делу.
EZRA|5|6|Вот содержание письма, которое послал Фафнай, заречный областеначальник, и Шефар–Бознай с товарищами своими Афарсахеями, которые за рекою, к царю Дарию.
EZRA|5|7|В донесении, которое они послали к нему, вот что написано: Дарию царю – всякий мир!
EZRA|5|8|Да будет известно царю, что мы ходили в Иудейскую область, к дому Бога великого; и строится он из больших камней, и дерево вкладывается в стены; и работа сия производится быстро и с успехом идет в руках их.
EZRA|5|9|Тогда мы спросили у старейшин тех и так сказали им: кто дал вам разрешение строить дом сей и стены сии доделывать?
EZRA|5|10|И сверх того об именах их мы спросили их, чтобы дать знать тебе и написать имена тех людей, которые главными у них.
EZRA|5|11|И они ответили нам такими словами: мы рабы Бога неба и земли и строим дом, который был построен за много лет прежде сего, – и великий царь у Израиля строил его и довершил его.
EZRA|5|12|Когда же отцы наши прогневали Бога небесного, Он предал их в руку Навуходоносора, царя Вавилонского, Халдеянина; и дом сей он разрушил, и народ переселил в Вавилон.
EZRA|5|13|Но в первый год Кира, царя Вавилонского, царь Кир дал разрешение построить сей дом Божий;
EZRA|5|14|да и сосуды дома Божия, золотые и серебряные, которые Навуходоносор вынес из храма Иерусалимского и отнес в храм Вавилонский, – вынес Кир царь из храма Вавилонского; и отдали [их] по имени Шешбацару, которого он назначил областеначальником,
EZRA|5|15|и сказал ему: возьми сии сосуды, пойди и отнеси их в храм Иерусалимский, и пусть дом Божий строится на своем месте.
EZRA|5|16|Тогда Шешбацар тот пришел, положил основания дома Божия в Иерусалиме; и с тех пор доселе он строится, и еще не кончен.
EZRA|5|17|Итак, если царю благоугодно, пусть поищут в доме царских сокровищ, там в Вавилоне, точно ли царем Киром дано разрешение строить сей дом Божий в Иерусалиме, и царскую волю о сем пусть пришлют к нам.
EZRA|6|1|Тогда царь Дарий дал повеление, и разыскивали в Вавилоне в книгохранилище, куда полагали сокровища.
EZRA|6|2|И найден в Екбатане во дворце, который в области Мидии, один свиток, и в нем написано так: "Для памяти:
EZRA|6|3|в первый год царя Кира, царь Кир дал повеление о доме Божием в Иерусалиме: пусть строится дом на том месте, где приносят жертвы, и пусть будут положены прочные основания для него; вышина его в шестьдесят локтей, ширина его в шестьдесят локтей;
EZRA|6|4|рядов из камней больших три, и ряд из дерева один; издержки же пусть выдаются из царского дома.
EZRA|6|5|Да и сосуды дома Божия, золотые и серебряные, которые Навуходоносор вынес из храма Иерусалимского и отнес в Вавилон, пусть возвратятся и пойдут в храм Иерусалимский, [каждый] на место свое, и помещены будут в доме Божием.
EZRA|6|6|Итак, Фафнай, заречный областеначальник, и Шефар–Бознай, с товарищами вашими Афарсахеями, которые за рекою, – удалитесь оттуда.
EZRA|6|7|Не останавливайте работы при сем доме Божием; пусть Иудейский областеначальник и Иудейские старейшины строят сей дом Божий на месте его.
EZRA|6|8|И от меня дается повеление о том, чем вы должны содействовать старейшинам тем Иудейским в построении того дома Божия, и [именно]: из имущества царского – [из] заречной подати – немедленно берите и давайте тем людям, чтобы работа не останавливалась;
EZRA|6|9|и сколько нужно – тельцов ли, или овнов и агнцев, на всесожжения Богу небесному, также пшеницы, соли, вина и масла, как скажут священники Иерусалимские, пусть будет выдаваемо им изо дня в день без задержки,
EZRA|6|10|чтоб они приносили жертву приятную Богу небесному и молились о жизни царя и сыновей его.
EZRA|6|11|Мною же дается повеление, что [если] какой человек изменит это определение, то будет вынуто бревно из дома его, и будет поднят он и пригвожден к нему, а дом его за то будет обращен в развалины.
EZRA|6|12|И Бог, Которого имя там обитает, да низложит всякого царя и народ, который простер бы руку свою, чтобы изменить [сие] ко вреду этого дома Божия в Иерусалиме. Я, Дарий, дал это повеление; да будет оно в точности исполняемо".
EZRA|6|13|Тогда Фафнай, заречный областеначальник, Шефар–Бознай и товарищи их, – как повелел царь Дарий, так в точности и делали.
EZRA|6|14|И старейшины Иудейские строили и преуспевали, по пророчеству Аггея пророка и Захарии, сына Адды. И построили и окончили, по воле Бога Израилева и по воле Кира и Дария и Артаксеркса, царей Персидских.
EZRA|6|15|И окончен дом сей к третьему дню месяца Адара, в шестой год царствования царя Дария.
EZRA|6|16|И совершили сыны Израилевы, священники и левиты и прочие, возвратившиеся из плена, освящение сего дома Божия с радостью.
EZRA|6|17|И принесли при освящении сего дома Божия: сто волов, двести овнов, четыреста агнцев и двенадцать козлов в жертву за грех за всего Израиля, по числу колен Израилевых.
EZRA|6|18|И поставили священников по отделениям их, и левитов по чередам их на службу Божию в Иерусалиме, как предписано в книге Моисея.
EZRA|6|19|И совершили возвратившиеся из плена пасху в четырнадцатый день первого месяца,
EZRA|6|20|потому что очистились священники и левиты, – все они, как один, [были] чисты; и закололи агнцев пасхальных для всех, возвратившихся из плена, для братьев своих священников и для себя.
EZRA|6|21|И ели сыны Израилевы, возвратившиеся из переселения, и все отделившиеся к ним от нечистоты народов земли, чтобы прибегать к Господу Богу Израилеву.
EZRA|6|22|И праздновали праздник опресноков семь дней в радости, потому что обрадовал их Господь и обратил к ним сердце царя Ассирийского, чтобы подкреплять руки их при строении дома Господа Бога Израилева.
EZRA|7|1|После сих происшествий, в царствование Артаксеркса, царя Персидского, Ездра, сын Сераии, сын Азарии, сын Хелкии,
EZRA|7|2|сын Шаллума, сын Садока, сын Ахитува,
EZRA|7|3|сын Амарии, сын Азарии, сын Марайофа,
EZRA|7|4|сын Захарии, сын Уззия, сын Буккия,
EZRA|7|5|сын Авишуя, сын Финееса, сын Елеазара, сын Аарона первосвященника, –
EZRA|7|6|сей Ездра вышел из Вавилона. Он был книжник, сведущий в законе Моисеевом, который дал Господь Бог Израилев. И дал ему царь все по желанию его, так как рука Господа Бога его [была] над ним.
EZRA|7|7|[С ним] пошли в Иерусалим и [некоторые] из сынов Израилевых, и из священников и левитов, и певцов и привратников и нефинеев в седьмой год царя Артаксеркса.
EZRA|7|8|И пришел он в Иерусалим в пятый месяц, – в седьмой же год царя.
EZRA|7|9|Ибо в первый день первого месяца [было] начало выхода из Вавилона, и в первый день пятого месяца он пришел в Иерусалим, так как благодеющая рука Бога его была над ним,
EZRA|7|10|потому что Ездра расположил сердце свое к тому, чтобы изучать закон Господень и исполнять [его], и учить в Израиле закону и правде.
EZRA|7|11|И вот содержание письма, которое дал царь Артаксеркс Ездре священнику, книжнику, учившему словам заповедей Господа и законов Его в Израиле:
EZRA|7|12|Артаксеркс, царь царей, Ездре священнику, учителю закона Бога небесного совершенному, и прочее.
EZRA|7|13|От меня дано повеление, чтобы в царстве моем всякий из народа Израилева и из священников его и левитов, желающий идти в Иерусалим, шел с тобою.
EZRA|7|14|Так как ты посылаешься от царя и семи советников его, чтобы обозреть Иудею и Иерусалим по закону Бога твоего, находящемуся в руке твоей,
EZRA|7|15|и чтобы доставить серебро и золото, которое царь и советники его пожертвовали Богу Израилеву, Которого жилище в Иерусалиме,
EZRA|7|16|и все серебро и золото, которое ты соберешь во всей области Вавилонской, вместе с доброхотными даяниями от народа и священников, которые пожертвуют они для дома Бога своего, что в Иерусалиме;
EZRA|7|17|поэтому немедленно купи на эти деньги волов, овнов, агнцев и хлебных приношений к ним и возлияний для них, и принеси их на жертвенник дома Бога вашего в Иерусалиме.
EZRA|7|18|И что тебе и братьям твоим заблагорассудится сделать из остального серебра и золота, то по воле Бога вашего делайте.
EZRA|7|19|И сосуды, которые даны тебе для служб [в] доме Бога твоего, поставь пред Богом Иерусалимским.
EZRA|7|20|И прочее потребное для дома Бога твоего, что ты признаешь нужным, давай из дома царских сокровищ.
EZRA|7|21|И от меня царя Артаксеркса дается повеление всем сокровищехранителям, которые за рекою: все, чего потребует у вас Ездра священник, учитель закона Бога небесного, немедленно давайте:
EZRA|7|22|серебра до ста талантов, и пшеницы до ста коров, и вина до ста батов, и до ста же батов масла, а соли без обозначения [количества].
EZRA|7|23|Все, что повелено Богом небесным, должно делаться со тщанием для дома Бога небесного; дабы не [было] гнева [Его] на царство, царя и сыновей его.
EZRA|7|24|И даем вам знать, чтобы [ни] на кого [из] священников или левитов, певцов, привратников, нефинеев и служащих при этом доме Божием, не налагать [ни] подати, [ни] налога, ни пошлины.
EZRA|7|25|Ты же, Ездра, по премудрости Бога твоего, которая в руке твоей, поставь правителей и судей, чтоб они судили весь народ за рекою, – всех знающих законы Бога твоего, а кто не знает, тех учите.
EZRA|7|26|Кто же не будет исполнять закон Бога твоего и закон царя, над тем немедленно пусть производят суд, на смерть ли, или на изгнание, или на денежную пеню, или на заключение в темницу.
EZRA|7|27|Благословен Господь, Бог отцов наших, вложивший в сердце царя – украсить дом Господень, который в Иерусалиме,
EZRA|7|28|и склонивший на меня милость царя и советников его, и всех могущественных князей царя! И я ободрился, ибо рука Господа Бога моего [была] надо мною, и собрал я глав Израиля, чтоб они пошли со мною.
EZRA|8|1|И вот главы поколений и родословие тех, которые вышли со мною из Вавилона, в царствование царя Артаксеркса:
EZRA|8|2|из сыновей Финееса Гирсон; из сыновей Ифамара Даниил; из сыновей Давида Хаттуш;
EZRA|8|3|из сыновей Шехании, из сыновей Пароша Захария, и с ним по списку родословному сто пятьдесят [человек] мужеского пола;
EZRA|8|4|из сыновей Пахаф–Моава Эльегоенай, сын Зерахии, и с ним двести [человек] мужеского пола;
EZRA|8|5|из сыновей Шехания, сын Яхазиила, и с ним триста [человек] мужеского пола;
EZRA|8|6|из сыновей Адина Евед, сын Ионафана, и с ним пятьдесят [человек] мужеского пола;
EZRA|8|7|из сыновей Елама Иешаия, сын Афалии, и с ним семьдесят [человек] мужеского пола;
EZRA|8|8|из сыновей Сафатии Зевадия, сын Михаилов, и с ним восемьдесят [человек] мужеского пола;
EZRA|8|9|из сыновей Иоава Овадия, сын Иехиелов, и с ним двести восемнадцать [человек] мужеского пола;
EZRA|8|10|из сыновей Шеломиф, сын Иосифии, и с ним сто шестьдесят [человек] мужеского пола;
EZRA|8|11|из сыновей Бевая Захария, сын Бевая, и с ним двадцать восемь [человек] мужеского пола;
EZRA|8|12|из сыновей Азгада Иоханан, сын Гаккатана, и с ним сто десять [человек] мужеского пола;
EZRA|8|13|из сыновей Адоникама последние, и вот имена их: Елифелет, Иеиел и Шемаия, и с ними шестьдесят [человек] мужеского пола;
EZRA|8|14|из сыновей Бигвая, Уфай и Заббуд, и с ними семьдесят [человек] мужеского пола.
EZRA|8|15|Я собрал их у реки, втекающей в Агаву, и мы простояли там три дня, и когда я осмотрел народ и священников, то из сынов Левия [никого] там не нашел.
EZRA|8|16|И послал я позвать Елиезера, Ариэла, Шемаию, и Элнафана, и Иарива, и Элнафана, и Нафана, и Захарию, и Мешуллама – главных, и Иоярива и Элнафана – ученых;
EZRA|8|17|и дал им поручение к Иддо, главному в местности Касифье, и вложил им в уста, что говорить к Иддо и братьям его, нефинеям в местности Касифье, чтобы они привели к нам служителей для дома Бога нашего.
EZRA|8|18|И привели они к нам, так как благодеющая рука Бога нашего была над нами, человека умного из сыновей Махлия, сына Левиина, сына Израилева, именно Шеревию, и сыновей его и братьев его, восемнадцать [человек];
EZRA|8|19|и Хашавию и с ним Иешаию из сыновей Мерариных, братьев его и сыновей их двадцать;
EZRA|8|20|и из нефинеев, которых дал Давид и князья [его] на прислугу левитам, двести двадцать нефинеев; все они названы поименно.
EZRA|8|21|И провозгласил я там пост у реки Агавы, чтобы смириться нам пред лицем Бога нашего, просить у Него благополучного пути для себя и для детей наших и для всего имущества нашего,
EZRA|8|22|так как мне стыдно было просить у царя войска и всадников для охранения нашего от врага на пути, ибо мы, говоря с царем, сказали: рука Бога нашего для всех прибегающих к Нему [есть] благодеющая, а на всех оставляющих Его – могущество Его и гнев Его!
EZRA|8|23|Итак мы постились и просили Бога нашего о сем, и Он услышал нас.
EZRA|8|24|И я отделил из начальствующих над священниками двенадцать [человек]: Шеревию, Хашавию и с ними десять из братьев их;
EZRA|8|25|и отдал им весом серебро, и золото, и сосуды, – все, пожертвованное [для] дома Бога нашего, что пожертвовали царь, и советники его, и князья его, и все Израильтяне, [там] находившиеся.
EZRA|8|26|И отдал на руки им весом: серебра – шестьсот пятьдесят талантов, и серебряных сосудов на сто талантов, золота – сто талантов;
EZRA|8|27|и чаш золотых – двадцать, в тысячу драхм, и два сосуда из лучшей блестящей меди, ценимой как золото.
EZRA|8|28|И сказал я им: вы – святыня Господу, и сосуды – святыня, и серебро и золото – доброхотное даяние Господу Богу отцов ваших.
EZRA|8|29|Будьте же бдительны и сберегите [это], доколе весом не сдадите начальствующим над священниками и левитами и главам поколений Израилевых в Иерусалиме, в хранилище при доме Господнем.
EZRA|8|30|И приняли священники и левиты взвешенное серебро, и золото, и сосуды, чтоб отнести в Иерусалим в дом Бога нашего.
EZRA|8|31|И отправились мы от реки Агавы в двенадцатый день первого месяца, чтобы идти в Иерусалим; и рука Бога нашего была над нами, и спасала нас от руки врага и от подстерегающих нас на пути.
EZRA|8|32|И пришли мы в Иерусалим, и пробыли там три дня.
EZRA|8|33|В четвертый день мы сдали весом серебро, и золото, и сосуды в дом Бога нашего, на руки Меремофу, сыну Урии, священнику, и с ним Елеазару, сыну Финеесову, и с ними Иозаваду, сыну Иисусову, и Ноадии, сыну Виннуя, левитам,
EZRA|8|34|все счетом и весом. И все взвешенное записано в то же время.
EZRA|8|35|Пришедшие из плена переселенцы принесли во всесожжение Богу Израилеву двенадцать тельцов из всего Израиля, девяносто шесть овнов, семьдесят семь агнцев и двенадцать козлов в жертву за грех: все это во всесожжение Господу.
EZRA|8|36|И отдали царские повеления царским сатрапам и заречным областеначальникам, и они почтили народ и дом Божий.
EZRA|9|1|По окончании сего, подошли ко мне начальствующие и сказали: народ Израилев и священники и левиты не отделились от народов иноплеменных с мерзостями их, от Хананеев, Хеттеев, Ферезеев, Иевусеев, Аммонитян, Моавитян, Египтян и Аморреев,
EZRA|9|2|потому что взяли дочерей их за себя и за сыновей своих, и смешалось семя святое с народами иноплеменными, и притом рука знатнейших и главнейших была в сем беззаконии первою.
EZRA|9|3|Услышав это слово, я разодрал нижнюю и верхнюю одежду мою и рвал волосы на голове моей и на бороде моей, и сидел печальный.
EZRA|9|4|Тогда собрались ко мне все, убоявшиеся слов Бога Израилева по причине преступления переселенцев, и я сидел в печали до вечерней жертвы.
EZRA|9|5|А во время вечерней жертвы я встал с места сетования моего, и в разодранной нижней и верхней одежде пал на колени мои и простер руки мои к Господу Богу моему
EZRA|9|6|и сказал: Боже мой! стыжусь и боюсь поднять лице мое к Тебе, Боже мой, потому что беззакония наши стали выше головы, и вина наша возросла до небес.
EZRA|9|7|Со дней отцов наших мы в великой вине до сего дня, и за беззакония наши преданы были мы, цари наши, священники наши, в руки царей иноземных, под меч, в плен и на разграбление и на посрамление, как это и ныне.
EZRA|9|8|И вот, по малом времени, даровано нам помилование от Господа Бога нашего, и Он оставил у нас [несколько] уцелевших и дал нам утвердиться на месте святыни Его, и просветил глаза наши Бог наш, и дал нам ожить немного в рабстве нашем.
EZRA|9|9|Мы – рабы, но и в рабстве нашем не оставил нас Бог наш. И склонил Он к нам милость царей Персидских, чтоб они дали нам ожить, воздвигнуть дом Бога нашего и восстановить [его] из развалин его, и дали нам ограждение в Иудее и в Иерусалиме.
EZRA|9|10|И ныне, что скажем мы, Боже наш, после этого? Ибо мы отступили от заповедей Твоих,
EZRA|9|11|которые заповедал Ты чрез рабов Твоих пророков, говоря: земля, в которую идете вы, чтоб овладеть ею, земля нечистая, она осквернена нечистотою иноплеменных народов, их мерзостями, которыми они наполнили ее от края до края в осквернениях своих.
EZRA|9|12|Итак дочерей ваших не выдавайте за сыновей их, и дочерей их не берите за сыновей ваших, и не ищите мира их и блага их во веки, чтобы укрепиться вам и питаться благами земли той и передать ее в наследие сыновьям вашим на веки.
EZRA|9|13|И после всего, постигшего нас за худые дела наши и за великую вину нашу, – ибо Ты, Боже наш, пощадил нас не по мере беззакония нашего и дал нам такое избавление, –
EZRA|9|14|неужели мы опять будем нарушать заповеди Твои и вступать в родство с этими отвратительными народами? Не прогневаешься ли Ты на нас даже до истребления [нас], так что не будет уцелевших и не будет спасения?
EZRA|9|15|Господи Боже Израилев! праведен Ты. Ибо мы остались уцелевшими до сего дня; и вот мы в беззакониях наших пред лицем Твоим, хотя после этого не надлежало бы нам стоять пред лицем Твоим.
EZRA|10|1|Когда [так] молился Ездра и исповедывался, плача и повергаясь пред домом Божиим, стеклось к нему весьма большое собрание Израильтян, мужчин и женщин и детей, потому что и народ много плакал.
EZRA|10|2|И отвечал Шехания, сын Иехиила из сыновей Еламовых, и сказал Ездре: мы сделали преступление пред Богом нашим, что взяли [себе] жен иноплеменных из народов земли, но есть еще надежда для Израиля в этом деле;
EZRA|10|3|заключим теперь завет с Богом нашим, что, по совету господина моего и благоговеющих пред заповедями Бога нашего, мы отпустим [от себя] всех жен и [детей], рожденных ими, – и да будет по закону!
EZRA|10|4|Встань, потому что это твое дело, и мы с тобою: ободрись и действуй!
EZRA|10|5|И встал Ездра, и велел начальствующим над священниками, левитами и всем Израилем дать клятву, что они сделают так. И они дали клятву.
EZRA|10|6|И встал Ездра и пошел от дома Божия в жилище Иоханана, сына Елияшивова, и пришел туда. Хлеба он не ел и воды не пил, потому что плакал о преступлении переселенцев.
EZRA|10|7|И объявили в Иудее и в Иерусалиме всем [бывшим] в плену, чтоб они собрались в Иерусалим;
EZRA|10|8|а кто не придет чрез три дня, на все имение того, по определению начальствующих и старейшин, будет положено заклятие, и сам он будет отлучен от общества переселенцев.
EZRA|10|9|И собрались все жители Иудеи и земли Вениаминовой в Иерусалим в три дня. Это [было] в девятом месяце, в двадцатый день месяца. И сидел весь народ на площади у дома Божия, дрожа как по этому делу, так и от дождей.
EZRA|10|10|И встал Ездра священник и сказал им: вы сделали преступление, взяв себе жен иноплеменных, и тем увеличили вину Израиля.
EZRA|10|11|Итак покайтесь [в сем] пред Господом Богом отцов ваших, и исполните волю Его, и отлучите себя от народов земли и от жен иноплеменных.
EZRA|10|12|И отвечало все собрание, и сказало громким голосом: как ты сказал, так и сделаем.
EZRA|10|13|Однако же народ многочислен и время [теперь] дождливое, и нет возможности стоять на улице. Да и это дело не одного дня и не двух, потому что мы много в этом деле погрешили.
EZRA|10|14|Пусть наши начальствующие заступят место всего общества, и все в городах наших, которые взяли жен иноплеменных, пусть приходят сюда в назначенные времена и с ними старейшины каждого города и судьи его, доколе не отвратится от нас пылающий гнев Бога нашего за это дело.
EZRA|10|15|Тогда Ионафан, сын Асаила, и Яхзеия, сын Фиквы, стали над этим делом, и Мешуллам и Шавфай левит были помощниками им.
EZRA|10|16|И сделали так вышедшие из плена. И отделены [на это] Ездра священник, главы поколений, от каждого поколения их, и все они [названы] поименно. И сделали они заседание в первый день десятого месяца, для исследования сего дела;
EZRA|10|17|и окончили [исследование] о всех, которые взяли жен иноплеменных, к первому дню первого месяца.
EZRA|10|18|И нашлись из сыновей священнических, которые взяли жен иноплеменных, – из сыновей Иисуса, сына Иоседекова, и братьев его: Маасея, Елиезер, Иарив и Гедалия;
EZRA|10|19|и они дали руки свои [во уверение], что отпустят жен своих, и [что они] повинны [принести] в жертву овна за свою вину;
EZRA|10|20|и из сыновей Иммера: Хананий и Зевадия;
EZRA|10|21|и из сыновей Харима: Маасея, Елия, Шемаия, Иехиил и Уззия;
EZRA|10|22|и из сыновей Пашхура: Елиоенай, Маасея, Исмаил, Нафанаил, Иозавад и Эласа;
EZRA|10|23|и из левитов: Иозавад, Шимей и Келаия, он же Клита, Пафахия, Иуда и Елиезер;
EZRA|10|24|и из певцов: Елияшив; и из привратников: Шаллум, Телем и Урий;
EZRA|10|25|а из Израильтян, – из сыновей Пароша: Рамаия, Иззия, Малхия, Миямин, Елеазар, Малхия и Венаия;
EZRA|10|26|и из сыновей Елама: Матфания, Захария, Иехиел, Авдий, Иремоф и Елия;
EZRA|10|27|и из сыновей Заффу: Елиоенай, Елияшив, Матфания, Иремоф, Завад и Азиса;
EZRA|10|28|и из сыновей Бевая: Иоханан, Ханания, Забвай и Афлай;
EZRA|10|29|и из сыновей Вания: Мешуллам, Маллух, Адая, Иашув, Шеал и Иерамоф;
EZRA|10|30|и из сыновей Пахаф–Моава: Адна, Хелал, Венаия, Маасея, Матфания, Веселеил, Биннуй и Манассия;
EZRA|10|31|и из сыновей Харима: Елиезер, Ишшия, Малхия, Шемаия, Симеон,
EZRA|10|32|Вениамин, Маллух, Шемария;
EZRA|10|33|и из сыновей Хашума: Мафнай, Мафафа, Завад, Елифелет, Иеремай, Манассия и Шимей;
EZRA|10|34|и из сыновей Вания: Маадай, Амрам и Уел,
EZRA|10|35|Бенаия, Бидья, Келуги,
EZRA|10|36|Ванея, Меремоф, Елиашив,
EZRA|10|37|Матфания, Мафнай, Иаасай,
EZRA|10|38|Ваний, Биннуй, Шимей,
EZRA|10|39|Шелемия, Нафан, Адаия,
EZRA|10|40|Махнадбай, Шашай, Шарай,
EZRA|10|41|Азариел, Шелемиягу, Шемария,
EZRA|10|42|Шаллум, Амария и Иосиф;
EZRA|10|43|и из сыновей Нево: Иеиел, Матфифия, Завад, Зевина, Иаддай, Иоель и Бенаия.
EZRA|10|44|Все сии взяли [за себя] жен иноплеменных, и некоторые из сих жен родили им детей.
