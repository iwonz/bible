1COR|1|1|Paulus vocatus apostolus Christi Iesu per voluntatem Dei et Sosthenes frater
1COR|1|2|ecclesiae Dei quae est Corinthi sanctificatis in Christo Iesu vocatis sanctis cum omnibus qui invocant nomen Domini nostri Iesu Christi in omni loco ipsorum et nostro
1COR|1|3|gratia vobis et pax a Deo Patre nostro et Domino Iesu Christo
1COR|1|4|gratias ago Deo meo semper pro vobis in gratia Dei quae data est vobis in Christo Iesu
1COR|1|5|quia in omnibus divites facti estis in illo in omni verbo et in omni scientia
1COR|1|6|sicut testimonium Christi confirmatum est in vobis
1COR|1|7|ita ut nihil vobis desit in ulla gratia expectantibus revelationem Domini nostri Iesu Christi
1COR|1|8|qui et confirmabit vos usque ad finem sine crimine in die adventus Domini nostri Iesu Christi
1COR|1|9|fidelis Deus per quem vocati estis in societatem Filii eius Iesu Christi Domini nostri
1COR|1|10|obsecro autem vos fratres per nomen Domini nostri Iesu Christi ut id ipsum dicatis omnes et non sint in vobis scismata sitis autem perfecti in eodem sensu et in eadem sententia
1COR|1|11|significatum est enim mihi de vobis fratres mei ab his qui sunt Chloes quia contentiones inter vos sunt
1COR|1|12|hoc autem dico quod unusquisque vestrum dicit ego quidem sum Pauli ego autem Apollo ego vero Cephae ego autem Christi
1COR|1|13|divisus est Christus numquid Paulus crucifixus est pro vobis aut in nomine Pauli baptizati estis
1COR|1|14|gratias ago Deo quod neminem vestrum baptizavi nisi Crispum et Gaium
1COR|1|15|ne quis dicat quod in nomine meo baptizati sitis
1COR|1|16|baptizavi autem et Stephanae domum ceterum nescio si quem alium baptizaverim
1COR|1|17|non enim misit me Christus baptizare sed evangelizare non in sapientia verbi ut non evacuetur crux Christi
1COR|1|18|verbum enim crucis pereuntibus quidem stultitia est his autem qui salvi fiunt id est nobis virtus Dei est
1COR|1|19|scriptum est enim perdam sapientiam sapientium et prudentiam prudentium reprobabo
1COR|1|20|ubi sapiens ubi scriba ubi conquisitor huius saeculi nonne stultam fecit Deus sapientiam huius mundi
1COR|1|21|nam quia in Dei sapientia non cognovit mundus per sapientiam Deum placuit Deo per stultitiam praedicationis salvos facere credentes
1COR|1|22|quoniam et Iudaei signa petunt et Graeci sapientiam quaerunt
1COR|1|23|nos autem praedicamus Christum crucifixum Iudaeis quidem scandalum gentibus autem stultitiam
1COR|1|24|ipsis autem vocatis Iudaeis atque Graecis Christum Dei virtutem et Dei sapientiam
1COR|1|25|quia quod stultum est Dei sapientius est hominibus et quod infirmum est Dei fortius est hominibus
1COR|1|26|videte enim vocationem vestram fratres quia non multi sapientes secundum carnem non multi potentes non multi nobiles
1COR|1|27|sed quae stulta sunt mundi elegit Deus ut confundat sapientes et infirma mundi elegit Deus ut confundat fortia
1COR|1|28|et ignobilia mundi et contemptibilia elegit Deus et quae non sunt ut ea quae sunt destrueret
1COR|1|29|ut non glorietur omnis caro in conspectu eius
1COR|1|30|ex ipso autem vos estis in Christo Iesu qui factus est sapientia nobis a Deo et iustitia et sanctificatio et redemptio
1COR|1|31|ut quemadmodum scriptum est qui gloriatur in Domino glorietur
1COR|2|1|et ego cum venissem ad vos fratres veni non per sublimitatem sermonis aut sapientiae adnuntians vobis testimonium Christi
1COR|2|2|non enim iudicavi scire me aliquid inter vos nisi Iesum Christum et hunc crucifixum
1COR|2|3|et ego in infirmitate et timore et tremore multo fui apud vos
1COR|2|4|et sermo meus et praedicatio mea non in persuasibilibus sapientiae verbis sed in ostensione Spiritus et virtutis
1COR|2|5|ut fides vestra non sit in sapientia hominum sed in virtute Dei
1COR|2|6|sapientiam autem loquimur inter perfectos sapientiam vero non huius saeculi neque principum huius saeculi qui destruuntur
1COR|2|7|sed loquimur Dei sapientiam in mysterio quae abscondita est quam praedestinavit Deus ante saecula in gloriam nostram
1COR|2|8|quam nemo principum huius saeculi cognovit si enim cognovissent numquam Dominum gloriae crucifixissent
1COR|2|9|sed sicut scriptum est quod oculus non vidit nec auris audivit nec in cor hominis ascendit quae praeparavit Deus his qui diligunt illum
1COR|2|10|nobis autem revelavit Deus per Spiritum suum Spiritus enim omnia scrutatur etiam profunda Dei
1COR|2|11|quis enim scit hominum quae sint hominis nisi spiritus hominis qui in ipso est ita et quae Dei sunt nemo cognovit nisi Spiritus Dei
1COR|2|12|nos autem non spiritum mundi accepimus sed Spiritum qui ex Deo est ut sciamus quae a Deo donata sunt nobis
1COR|2|13|quae et loquimur non in doctis humanae sapientiae verbis sed in doctrina Spiritus spiritalibus spiritalia conparantes
1COR|2|14|animalis autem homo non percipit ea quae sunt Spiritus Dei stultitia est enim illi et non potest intellegere quia spiritaliter examinatur
1COR|2|15|spiritalis autem iudicat omnia et ipse a nemine iudicatur
1COR|2|16|quis enim cognovit sensum Domini qui instruat eum nos autem sensum Christi habemus
1COR|3|1|et ego fratres non potui vobis loqui quasi spiritalibus sed quasi carnalibus tamquam parvulis in Christo
1COR|3|2|lac vobis potum dedi non escam nondum enim poteratis sed ne nunc quidem potestis adhuc enim estis carnales
1COR|3|3|cum enim sit inter vos zelus et contentio nonne carnales estis et secundum hominem ambulatis
1COR|3|4|cum enim quis dicit ego quidem sum Pauli alius autem ego Apollo nonne homines estis quid igitur est Apollo quid vero Paulus
1COR|3|5|ministri eius cui credidistis et unicuique sicut Dominus dedit
1COR|3|6|ego plantavi Apollo rigavit sed Deus incrementum dedit
1COR|3|7|itaque neque qui plantat est aliquid neque qui rigat sed qui incrementum dat Deus
1COR|3|8|qui plantat autem et qui rigat unum sunt unusquisque autem propriam mercedem accipiet secundum suum laborem
1COR|3|9|Dei enim sumus adiutores Dei agricultura estis Dei aedificatio estis
1COR|3|10|secundum gratiam Dei quae data est mihi ut sapiens architectus fundamentum posui alius autem superaedificat unusquisque autem videat quomodo superaedificet
1COR|3|11|fundamentum enim aliud nemo potest ponere praeter id quod positum est qui est Christus Iesus
1COR|3|12|si quis autem superaedificat supra fundamentum hoc aurum argentum lapides pretiosos ligna faenum stipulam
1COR|3|13|uniuscuiusque opus manifestum erit dies enim declarabit quia in igne revelabitur et uniuscuiusque opus quale sit ignis probabit
1COR|3|14|si cuius opus manserit quod superaedificavit mercedem accipiet
1COR|3|15|si cuius opus arserit detrimentum patietur ipse autem salvus erit sic tamen quasi per ignem
1COR|3|16|nescitis quia templum Dei estis et Spiritus Dei habitat in vobis
1COR|3|17|si quis autem templum Dei violaverit disperdet illum Deus templum enim Dei sanctum est quod estis vos
1COR|3|18|nemo se seducat si quis videtur inter vos sapiens esse in hoc saeculo stultus fiat ut sit sapiens
1COR|3|19|sapientia enim huius mundi stultitia est apud Deum scriptum est enim conprehendam sapientes in astutia eorum
1COR|3|20|et iterum Dominus novit cogitationes sapientium quoniam vanae sunt
1COR|3|21|itaque nemo glorietur in hominibus omnia enim vestra sunt
1COR|3|22|sive Paulus sive Apollo sive Cephas sive mundus sive vita sive mors sive praesentia sive futura omnia enim vestra sunt
1COR|3|23|vos autem Christi Christus autem Dei
1COR|4|1|sic nos existimet homo ut ministros Christi et dispensatores mysteriorum Dei
1COR|4|2|hic iam quaeritur inter dispensatores ut fidelis quis inveniatur
1COR|4|3|mihi autem pro minimo est ut a vobis iudicer aut ab humano die sed neque me ipsum iudico
1COR|4|4|nihil enim mihi conscius sum sed non in hoc iustificatus sum qui autem iudicat me Dominus est
1COR|4|5|itaque nolite ante tempus iudicare quoadusque veniat Dominus qui et inluminabit abscondita tenebrarum et manifestabit consilia cordium et tunc laus erit unicuique a Deo
1COR|4|6|haec autem fratres transfiguravi in me et Apollo propter vos ut in nobis discatis ne supra quam scriptum est unus adversus alterum infletur pro alio
1COR|4|7|quis enim te discernit quid autem habes quod non accepisti si autem accepisti quid gloriaris quasi non acceperis
1COR|4|8|iam saturati estis iam divites facti estis sine nobis regnastis et utinam regnaretis ut et nos vobiscum regnaremus
1COR|4|9|puto enim Deus nos apostolos novissimos ostendit tamquam morti destinatos quia spectaculum facti sumus mundo et angelis et hominibus
1COR|4|10|nos stulti propter Christum vos autem prudentes in Christo nos infirmi vos autem fortes vos nobiles nos autem ignobiles
1COR|4|11|usque in hanc horam et esurimus et sitimus et nudi sumus et colaphis caedimur et instabiles sumus
1COR|4|12|et laboramus operantes manibus nostris maledicimur et benedicimus persecutionem patimur et sustinemus
1COR|4|13|blasphemamur et obsecramus tamquam purgamenta huius mundi facti sumus omnium peripsima usque adhuc
1COR|4|14|non ut confundam vos haec scribo sed ut filios meos carissimos moneo
1COR|4|15|nam si decem milia pedagogorum habeatis in Christo sed non multos patres nam in Christo Iesu per evangelium ego vos genui
1COR|4|16|rogo ergo vos imitatores mei estote
1COR|4|17|ideo misi ad vos Timotheum qui est filius meus carissimus et fidelis in Domino qui vos commonefaciat vias meas quae sunt in Christo sicut ubique in omni ecclesia doceo
1COR|4|18|tamquam non venturus sim ad vos sic inflati sunt quidam
1COR|4|19|veniam autem cito ad vos si Dominus voluerit et cognoscam non sermonem eorum qui inflati sunt sed virtutem
1COR|4|20|non enim in sermone est regnum Dei sed in virtute
1COR|4|21|quid vultis in virga veniam ad vos an in caritate et spiritu mansuetudinis
1COR|5|1|omnino auditur inter vos fornicatio et talis fornicatio qualis nec inter gentes ita ut uxorem patris aliquis habeat
1COR|5|2|et vos inflati estis et non magis luctum habuistis ut tollatur de medio vestrum qui hoc opus fecit
1COR|5|3|ego quidem absens corpore praesens autem spiritu iam iudicavi ut praesens eum qui sic operatus est
1COR|5|4|in nomine Domini nostri Iesu Christi congregatis vobis et meo spiritu cum virtute Domini Iesu
1COR|5|5|tradere huiusmodi Satanae in interitum carnis ut spiritus salvus sit in die Domini Iesu
1COR|5|6|non bona gloriatio vestra nescitis quia modicum fermentum totam massam corrumpit
1COR|5|7|expurgate vetus fermentum ut sitis nova consparsio sicut estis azymi etenim pascha nostrum immolatus est Christus
1COR|5|8|itaque epulemur non in fermento veteri neque in fermento malitiae et nequitiae sed in azymis sinceritatis et veritatis
1COR|5|9|scripsi vobis in epistula ne commisceamini fornicariis
1COR|5|10|non utique fornicariis huius mundi aut avaris aut rapacibus aut idolis servientibus alioquin debueratis de hoc mundo exisse
1COR|5|11|nunc autem scripsi vobis non commisceri si is qui frater nominatur est fornicator aut avarus aut idolis serviens aut maledicus aut ebriosus aut rapax cum eiusmodi nec cibum sumere
1COR|5|12|quid enim mihi de his qui foris sunt iudicare nonne de his qui intus sunt vos iudicatis
1COR|5|13|nam eos qui foris sunt Deus iudicabit auferte malum ex vobis ipsis
1COR|6|1|audet aliquis vestrum habens negotium adversus alterum iudicari apud iniquos et non apud sanctos
1COR|6|2|an nescitis quoniam sancti de mundo iudicabunt et si in vobis iudicabitur mundus indigni estis qui de minimis iudicetis
1COR|6|3|nescitis quoniam angelos iudicabimus quanto magis saecularia
1COR|6|4|saecularia igitur iudicia si habueritis contemptibiles qui sunt in ecclesia illos constituite ad iudicandum
1COR|6|5|ad verecundiam vestram dico sic non est inter vos sapiens quisquam qui possit iudicare inter fratrem suum
1COR|6|6|sed frater cum fratre iudicio contendit et hoc apud infideles
1COR|6|7|iam quidem omnino delictum est in vobis quod iudicia habetis inter vos quare non magis iniuriam accipitis quare non magis fraudem patimini
1COR|6|8|sed vos iniuriam facitis et fraudatis et hoc fratribus
1COR|6|9|an nescitis quia iniqui regnum Dei non possidebunt nolite errare neque fornicarii neque idolis servientes neque adulteri
1COR|6|10|neque molles neque masculorum concubitores neque fures neque avari neque ebriosi neque maledici neque rapaces regnum Dei possidebunt
1COR|6|11|et haec quidam fuistis sed abluti estis sed sanctificati estis sed iustificati estis in nomine Domini nostri Iesu Christi et in Spiritu Dei nostri
1COR|6|12|omnia mihi licent sed non omnia expediunt omnia mihi licent sed ego sub nullius redigar potestate
1COR|6|13|esca ventri et venter escis Deus autem et hunc et haec destruet corpus autem non fornicationi sed Domino et Dominus corpori
1COR|6|14|Deus vero et Dominum suscitavit et nos suscitabit per virtutem suam
1COR|6|15|nescitis quoniam corpora vestra membra Christi sunt tollens ergo membra Christi faciam membra meretricis absit
1COR|6|16|an nescitis quoniam qui adheret meretrici unum corpus efficitur erunt enim inquit duo in carne una
1COR|6|17|qui autem adheret Domino unus spiritus est
1COR|6|18|fugite fornicationem omne peccatum quodcumque fecerit homo extra corpus est qui autem fornicatur in corpus suum peccat
1COR|6|19|an nescitis quoniam membra vestra templum est Spiritus Sancti qui in vobis est quem habetis a Deo et non estis vestri
1COR|6|20|empti enim estis pretio magno glorificate et portate Deum in corpore vestro
1COR|7|1|de quibus autem scripsistis bonum est homini mulierem non tangere
1COR|7|2|propter fornicationes autem unusquisque suam uxorem habeat et unaquaeque suum virum habeat
1COR|7|3|uxori vir debitum reddat similiter autem et uxor viro
1COR|7|4|mulier sui corporis potestatem non habet sed vir similiter autem et vir sui corporis potestatem non habet sed mulier
1COR|7|5|nolite fraudare invicem nisi forte ex consensu ad tempus ut vacetis orationi et iterum revertimini in id ipsum ne temptet vos Satanas propter incontinentiam vestram
1COR|7|6|hoc autem dico secundum indulgentiam non secundum imperium
1COR|7|7|volo autem omnes homines esse sicut me ipsum sed unusquisque proprium habet donum ex Deo alius quidem sic alius vero sic
1COR|7|8|dico autem non nuptis et viduis bonum est illis si sic maneant sicut et ego
1COR|7|9|quod si non se continent nubant melius est enim nubere quam uri
1COR|7|10|his autem qui matrimonio iuncti sunt praecipio non ego sed Dominus uxorem a viro non discedere
1COR|7|11|quod si discesserit manere innuptam aut viro suo reconciliari et vir uxorem ne dimittat
1COR|7|12|nam ceteris ego dico non Dominus si quis frater uxorem habet infidelem et haec consentit habitare cum illo non dimittat illam
1COR|7|13|et si qua mulier habet virum infidelem et hic consentit habitare cum illa non dimittat virum
1COR|7|14|sanctificatus est enim vir infidelis in muliere fideli et sanctificata est mulier infidelis per virum fidelem alioquin filii vestri inmundi essent nunc autem sancti sunt
1COR|7|15|quod si infidelis discedit discedat non est enim servituti subiectus frater aut soror in eiusmodi in pace autem vocavit nos Deus
1COR|7|16|unde enim scis mulier si virum salvum facies aut unde scis vir si mulierem salvam facies
1COR|7|17|nisi unicuique sicut divisit Dominus unumquemque sicut vocavit Deus ita ambulet et sic in omnibus ecclesiis doceo
1COR|7|18|circumcisus aliquis vocatus est non adducat praeputium in praeputio aliquis vocatus est non circumcidatur
1COR|7|19|circumcisio nihil est et praeputium nihil est sed observatio mandatorum Dei
1COR|7|20|unusquisque in qua vocatione vocatus est in ea permaneat
1COR|7|21|servus vocatus es non sit tibi curae sed et si potes liber fieri magis utere
1COR|7|22|qui enim in Domino vocatus est servus libertus est Domini similiter qui liber vocatus est servus est Christi
1COR|7|23|pretio empti estis nolite fieri servi hominum
1COR|7|24|unusquisque in quo vocatus est fratres in hoc maneat apud Deum
1COR|7|25|de virginibus autem praeceptum Domini non habeo consilium autem do tamquam misericordiam consecutus a Domino ut sim fidelis
1COR|7|26|existimo ergo hoc bonum esse propter instantem necessitatem quoniam bonum est homini sic esse
1COR|7|27|alligatus es uxori noli quaerere solutionem solutus es ab uxore noli quaerere uxorem
1COR|7|28|si autem acceperis uxorem non peccasti et si nupserit virgo non peccavit tribulationem tamen carnis habebunt huiusmodi ego autem vobis parco
1COR|7|29|hoc itaque dico fratres tempus breve est reliquum est ut qui habent uxores tamquam non habentes sint
1COR|7|30|et qui flent tamquam non flentes et qui gaudent tamquam non gaudentes et qui emunt tamquam non possidentes
1COR|7|31|et qui utuntur hoc mundo tamquam non utantur praeterit enim figura huius mundi
1COR|7|32|volo autem vos sine sollicitudine esse qui sine uxore est sollicitus est quae Domini sunt quomodo placeat Deo
1COR|7|33|qui autem cum uxore est sollicitus est quae sunt mundi quomodo placeat uxori et divisus est
1COR|7|34|et mulier innupta et virgo cogitat quae Domini sunt ut sit sancta et corpore et spiritu quae autem nupta est cogitat quae sunt mundi quomodo placeat viro
1COR|7|35|porro hoc ad utilitatem vestram dico non ut laqueum vobis iniciam sed ad id quod honestum est et quod facultatem praebeat sine inpedimento Dominum observandi
1COR|7|36|si quis autem turpem se videri existimat super virgine sua quod sit superadulta et ita oportet fieri quod vult faciat non peccat nubat
1COR|7|37|nam qui statuit in corde suo firmus non habens necessitatem potestatem autem habet suae voluntatis et hoc iudicavit in corde suo servare virginem suam bene facit
1COR|7|38|igitur et qui matrimonio iungit virginem suam bene facit et qui non iungit melius facit
1COR|7|39|mulier alligata est quanto tempore vir eius vivit quod si dormierit vir eius liberata est cui vult nubat tantum in Domino
1COR|7|40|beatior autem erit si sic permanserit secundum meum consilium puto autem quod et ego Spiritum Dei habeo
1COR|8|1|de his autem quae idolis sacrificantur scimus quia omnes scientiam habemus scientia inflat caritas vero aedificat
1COR|8|2|si quis se existimat scire aliquid nondum cognovit quemadmodum oporteat eum scire
1COR|8|3|si quis autem diligit Deum hic cognitus est ab eo
1COR|8|4|de escis autem quae idolis immolantur scimus quia nihil est idolum in mundo et quod nullus Deus nisi unus
1COR|8|5|nam et si sunt qui dicantur dii sive in caelo sive in terra siquidem sunt dii multi et domini multi
1COR|8|6|nobis tamen unus Deus Pater ex quo omnia et nos in illum et unus Dominus Iesus Christus per quem omnia et nos per ipsum
1COR|8|7|sed non in omnibus est scientia quidam autem conscientia usque nunc idoli quasi idolothytum manducant et conscientia ipsorum cum sit infirma polluitur
1COR|8|8|esca autem nos non commendat Deo neque si non manducaverimus deficiemus neque si manducaverimus abundabimus
1COR|8|9|videte autem ne forte haec licentia vestra offendiculum fiat infirmibus
1COR|8|10|si enim quis viderit eum qui habet scientiam in idolio recumbentem nonne conscientia eius cum sit infirma aedificabitur ad manducandum idolothyta
1COR|8|11|et peribit infirmus in tua scientia frater propter quem Christus mortuus est
1COR|8|12|sic autem peccantes in fratres et percutientes conscientiam eorum infirmam in Christo peccatis
1COR|8|13|quapropter si esca scandalizat fratrem meum non manducabo carnem in aeternum ne fratrem meum scandalizem
1COR|9|1|non sum liber non sum apostolus nonne Iesum Dominum nostrum vidi non opus meum vos estis in Domino
1COR|9|2|si aliis non sum apostolus sed tamen vobis sum nam signaculum apostolatus mei vos estis in Domino
1COR|9|3|mea defensio apud eos qui me interrogant haec est
1COR|9|4|numquid non habemus potestatem manducandi et bibendi
1COR|9|5|numquid non habemus potestatem sororem mulierem circumducendi sicut et ceteri apostoli et fratres Domini et Cephas
1COR|9|6|aut solus ego et Barnabas non habemus potestatem hoc operandi
1COR|9|7|quis militat suis stipendiis umquam quis plantat vineam et fructum eius non edit quis pascit gregem et de lacte gregis non manducat
1COR|9|8|numquid secundum hominem haec dico an et lex haec non dicit
1COR|9|9|scriptum est enim in lege Mosi non alligabis os bovi trituranti numquid de bubus cura est Deo
1COR|9|10|an propter nos utique dicit nam propter nos scripta sunt quoniam debet in spe qui arat arare et qui triturat in spe fructus percipiendi
1COR|9|11|si nos vobis spiritalia seminavimus magnum est si nos carnalia vestra metamus
1COR|9|12|si alii potestatis vestrae participes sunt non potius nos sed non usi sumus hac potestate sed omnia sustinemus ne quod offendiculum demus evangelio Christi
1COR|9|13|nescitis quoniam qui in sacrario operantur quae de sacrario sunt edunt qui altario deserviunt cum altario participantur
1COR|9|14|ita et Dominus ordinavit his qui evangelium adnuntiant de evangelio vivere
1COR|9|15|ego autem nullo horum usus sum non scripsi autem haec ut ita fiant in me bonum est enim mihi magis mori quam ut gloriam meam quis evacuet
1COR|9|16|nam si evangelizavero non est mihi gloria necessitas enim mihi incumbit vae enim mihi est si non evangelizavero
1COR|9|17|si enim volens hoc ago mercedem habeo si autem invitus dispensatio mihi credita est
1COR|9|18|quae est ergo merces mea ut evangelium praedicans sine sumptu ponam evangelium ut non abutar potestate mea in evangelio
1COR|9|19|nam cum liber essem ex omnibus omnium me servum feci ut plures lucri facerem
1COR|9|20|et factus sum Iudaeis tamquam Iudaeus ut Iudaeos lucrarer
1COR|9|21|his qui sub lege sunt quasi sub lege essem cum ipse non essem sub lege ut eos qui sub lege erant lucri facerem his qui sine lege erant tamquam sine lege essem cum sine lege Dei non essem sed in lege essem Christi ut lucri facerem eos qui sine lege erant
1COR|9|22|factus sum infirmis infirmus ut infirmos lucri facerem omnibus omnia factus sum ut omnes facerem salvos
1COR|9|23|omnia autem facio propter evangelium ut particeps eius efficiar
1COR|9|24|nescitis quod hii qui in stadio currunt omnes quidem currunt sed unus accipit bravium sic currite ut conprehendatis
1COR|9|25|omnis autem qui in agone contendit ab omnibus se abstinet et illi quidem ut corruptibilem coronam accipiant nos autem incorruptam
1COR|9|26|ego igitur sic curro non quasi in incertum sic pugno non quasi aerem verberans
1COR|9|27|sed castigo corpus meum et in servitutem redigo ne forte cum aliis praedicaverim ipse reprobus efficiar
1COR|10|1|nolo enim vos ignorare fratres quoniam patres nostri omnes sub nube fuerunt et omnes mare transierunt
1COR|10|2|et omnes in Mose baptizati sunt in nube et in mari
1COR|10|3|et omnes eandem escam spiritalem manducaverunt
1COR|10|4|et omnes eundem potum spiritalem biberunt bibebant autem de spiritali consequenti eos petra petra autem erat Christus
1COR|10|5|sed non in pluribus eorum beneplacitum est Deo nam prostrati sunt in deserto
1COR|10|6|haec autem in figura facta sunt nostri ut non simus concupiscentes malorum sicut et illi concupierunt
1COR|10|7|neque idolorum cultores efficiamini sicut quidam ex ipsis quemadmodum scriptum est sedit populus manducare et bibere et surrexerunt ludere
1COR|10|8|neque fornicemur sicut quidam ex ipsis fornicati sunt et ceciderunt una die viginti tria milia
1COR|10|9|neque temptemus Christum sicut quidam eorum temptaverunt et a serpentibus perierunt
1COR|10|10|neque murmuraveritis sicut quidam eorum murmuraverunt et perierunt ab exterminatore
1COR|10|11|haec autem omnia in figura contingebant illis scripta sunt autem ad correptionem nostram in quos fines saeculorum devenerunt
1COR|10|12|itaque qui se existimat stare videat ne cadat
1COR|10|13|temptatio vos non adprehendat nisi humana fidelis autem Deus qui non patietur vos temptari super id quod potestis sed faciet cum temptatione etiam proventum ut possitis sustinere
1COR|10|14|propter quod carissimi mihi fugite ab idolorum cultura
1COR|10|15|ut prudentibus loquor vos iudicate quod dico
1COR|10|16|calicem benedictionis cui benedicimus nonne communicatio sanguinis Christi est et panis quem frangimus nonne participatio corporis Domini est
1COR|10|17|quoniam unus panis unum corpus multi sumus omnes quidem de uno pane participamur
1COR|10|18|videte Israhel secundum carnem nonne qui edunt hostias participes sunt altaris
1COR|10|19|quid ergo dico quod idolis immolatum sit aliquid aut quod idolum sit aliquid
1COR|10|20|sed quae immolant gentes daemoniis immolant et non Deo nolo autem vos socios fieri daemoniorum non potestis calicem Domini bibere et calicem daemoniorum
1COR|10|21|non potestis mensae Domini participes esse et mensae daemoniorum
1COR|10|22|an aemulamur Dominum numquid fortiores illo sumus omnia licent sed non omnia expediunt
1COR|10|23|omnia licent sed non omnia aedificant
1COR|10|24|nemo quod suum est quaerat sed quod alterius
1COR|10|25|omne quod in macello venit manducate nihil interrogantes propter conscientiam
1COR|10|26|Domini est terra et plenitudo eius
1COR|10|27|si quis vocat vos infidelium et vultis ire omne quod vobis adponitur manducate nihil interrogantes propter conscientiam
1COR|10|28|si quis autem dixerit hoc immolaticium est idolis nolite manducare propter illum qui indicavit et propter conscientiam
1COR|10|29|conscientiam autem dico non tuam sed alterius ut quid enim libertas mea iudicatur ab alia conscientia
1COR|10|30|si ego cum gratia participo quid blasphemor pro eo quod gratias ago
1COR|10|31|sive ergo manducatis sive bibitis vel aliud quid facitis omnia in gloriam Dei facite
1COR|10|32|sine offensione estote Iudaeis et gentilibus et ecclesiae Dei
1COR|10|33|sicut et ego per omnia omnibus placeo non quaerens quod mihi utile est sed quod multis ut salvi fiant
1COR|11|1|imitatores mei estote sicut et ego Christi
1COR|11|2|laudo autem vos fratres quod omnia mei memores estis et sicut tradidi vobis praecepta mea tenetis
1COR|11|3|volo autem vos scire quod omnis viri caput Christus est caput autem mulieris vir caput vero Christi Deus
1COR|11|4|omnis vir orans aut prophetans velato capite deturpat caput suum
1COR|11|5|omnis autem mulier orans aut prophetans non velato capite deturpat caput suum unum est enim atque si decalvetur
1COR|11|6|nam si non velatur mulier et tondeatur si vero turpe est mulieri tonderi aut decalvari velet caput suum
1COR|11|7|vir quidem non debet velare caput quoniam imago et gloria est Dei mulier autem gloria viri est
1COR|11|8|non enim vir ex muliere est sed mulier ex viro
1COR|11|9|etenim non est creatus vir propter mulierem sed mulier propter virum
1COR|11|10|ideo debet mulier potestatem habere supra caput propter angelos
1COR|11|11|verumtamen neque vir sine muliere neque mulier sine viro in Domino
1COR|11|12|nam sicut mulier de viro ita et vir per mulierem omnia autem ex Deo
1COR|11|13|vos ipsi iudicate decet mulierem non velatam orare Deum
1COR|11|14|nec ipsa natura docet vos quod vir quidem si comam nutriat ignominia est illi
1COR|11|15|mulier vero si comam nutriat gloria est illi quoniam capilli pro velamine ei dati sunt
1COR|11|16|si quis autem videtur contentiosus esse nos talem consuetudinem non habemus neque ecclesiae Dei
1COR|11|17|hoc autem praecipio non laudans quod non in melius sed in deterius convenitis
1COR|11|18|primum quidem convenientibus vobis in ecclesia audio scissuras esse et ex parte credo
1COR|11|19|nam oportet et hereses esse ut et qui probati sunt manifesti fiant in vobis
1COR|11|20|convenientibus ergo vobis in unum iam non est dominicam cenam manducare
1COR|11|21|unusquisque enim suam cenam praesumit ad manducandum et alius quidem esurit alius autem ebrius est
1COR|11|22|numquid domos non habetis ad manducandum et bibendum aut ecclesiam Dei contemnitis et confunditis eos qui non habent quid dicam vobis laudo vos in hoc non laudo
1COR|11|23|ego enim accepi a Domino quod et tradidi vobis quoniam Dominus Iesus in qua nocte tradebatur accepit panem
1COR|11|24|et gratias agens fregit et dixit hoc est corpus meum pro vobis hoc facite in meam commemorationem
1COR|11|25|similiter et calicem postquam cenavit dicens hic calix novum testamentum est in meo sanguine hoc facite quotienscumque bibetis in meam commemorationem
1COR|11|26|quotienscumque enim manducabitis panem hunc et calicem bibetis mortem Domini adnuntiatis donec veniat
1COR|11|27|itaque quicumque manducaverit panem vel biberit calicem Domini indigne reus erit corporis et sanguinis Domini
1COR|11|28|probet autem se ipsum homo et sic de pane illo edat et de calice bibat
1COR|11|29|qui enim manducat et bibit indigne iudicium sibi manducat et bibit non diiudicans corpus
1COR|11|30|ideo inter vos multi infirmes et inbecilles et dormiunt multi
1COR|11|31|quod si nosmet ipsos diiudicaremus non utique iudicaremur
1COR|11|32|dum iudicamur autem a Domino corripimur ut non cum hoc mundo damnemur
1COR|11|33|itaque fratres mei cum convenitis ad manducandum invicem expectate
1COR|11|34|si quis esurit domi manducet ut non in iudicium conveniatis cetera autem cum venero disponam
1COR|12|1|de spiritalibus autem nolo vos ignorare fratres
1COR|12|2|scitis quoniam cum gentes essetis ad simulacra muta prout ducebamini euntes
1COR|12|3|ideo notum vobis facio quod nemo in Spiritu Dei loquens dicit anathema Iesu et nemo potest dicere Dominus Iesus nisi in Spiritu Sancto
1COR|12|4|divisiones vero gratiarum sunt idem autem Spiritus
1COR|12|5|et divisiones ministrationum sunt idem autem Dominus
1COR|12|6|et divisiones operationum sunt idem vero Deus qui operatur omnia in omnibus
1COR|12|7|unicuique autem datur manifestatio Spiritus ad utilitatem
1COR|12|8|alii quidem per Spiritum datur sermo sapientiae alii autem sermo scientiae secundum eundem Spiritum
1COR|12|9|alteri fides in eodem Spiritu alii gratia sanitatum in uno Spiritu
1COR|12|10|alii operatio virtutum alii prophetatio alii discretio spirituum alii genera linguarum alii interpretatio sermonum
1COR|12|11|haec autem omnia operatur unus atque idem Spiritus dividens singulis prout vult
1COR|12|12|sicut enim corpus unum est et membra habet multa omnia autem membra corporis cum sint multa unum corpus sunt ita et Christus
1COR|12|13|etenim in uno Spiritu omnes nos in unum corpus baptizati sumus sive Iudaei sive gentiles sive servi sive liberi et omnes unum Spiritum potati sumus
1COR|12|14|nam et corpus non est unum membrum sed multa
1COR|12|15|si dixerit pes quoniam non sum manus non sum de corpore non ideo non est de corpore
1COR|12|16|et si dixerit auris quia non sum oculus non sum de corpore non ideo non est de corpore
1COR|12|17|si totum corpus oculus ubi auditus si totum auditus ubi odoratus
1COR|12|18|nunc autem posuit Deus membra unumquodque eorum in corpore sicut voluit
1COR|12|19|quod si essent omnia unum membrum ubi corpus
1COR|12|20|nunc autem multa quidem membra unum autem corpus
1COR|12|21|non potest dicere oculus manui opera tua non indigeo aut iterum caput pedibus non estis mihi necessarii
1COR|12|22|sed multo magis quae videntur membra corporis infirmiora esse necessariora sunt
1COR|12|23|et quae putamus ignobiliora membra esse corporis his honorem abundantiorem circumdamus et quae inhonesta sunt nostra abundantiorem honestatem habent
1COR|12|24|honesta autem nostra nullius egent sed Deus temperavit corpus ei cui deerat abundantiorem tribuendo honorem
1COR|12|25|ut non sit scisma in corpore sed id ipsum pro invicem sollicita sint membra
1COR|12|26|et si quid patitur unum membrum conpatiuntur omnia membra sive gloriatur unum membrum congaudent omnia membra
1COR|12|27|vos autem estis corpus Christi et membra de membro
1COR|12|28|et quosdam quidem posuit Deus in ecclesia primum apostolos secundo prophetas tertio doctores deinde virtutes exin gratias curationum opitulationes gubernationes genera linguarum
1COR|12|29|numquid omnes apostoli numquid omnes prophetae numquid omnes doctores
1COR|12|30|numquid omnes virtutes numquid omnes gratiam habent curationum numquid omnes linguis loquuntur numquid omnes interpretantur
1COR|12|31|aemulamini autem charismata maiora et adhuc excellentiorem viam vobis demonstro
1COR|13|1|si linguis hominum loquar et angelorum caritatem autem non habeam factus sum velut aes sonans aut cymbalum tinniens
1COR|13|2|et si habuero prophetiam et noverim mysteria omnia et omnem scientiam et habuero omnem fidem ita ut montes transferam caritatem autem non habuero nihil sum
1COR|13|3|et si distribuero in cibos pauperum omnes facultates meas et si tradidero corpus meum ut ardeam caritatem autem non habuero nihil mihi prodest
1COR|13|4|caritas patiens est benigna est caritas non aemulatur non agit perperam non inflatur
1COR|13|5|non est ambitiosa non quaerit quae sua sunt non inritatur non cogitat malum
1COR|13|6|non gaudet super iniquitatem congaudet autem veritati
1COR|13|7|omnia suffert omnia credit omnia sperat omnia sustinet
1COR|13|8|caritas numquam excidit sive prophetiae evacuabuntur sive linguae cessabunt sive scientia destruetur
1COR|13|9|ex parte enim cognoscimus et ex parte prophetamus
1COR|13|10|cum autem venerit quod perfectum est evacuabitur quod ex parte est
1COR|13|11|cum essem parvulus loquebar ut parvulus sapiebam ut parvulus cogitabam ut parvulus quando factus sum vir evacuavi quae erant parvuli
1COR|13|12|videmus nunc per speculum in enigmate tunc autem facie ad faciem nunc cognosco ex parte tunc autem cognoscam sicut et cognitus sum
1COR|13|13|nunc autem manet fides spes caritas tria haec maior autem his est caritas
1COR|14|1|sectamini caritatem aemulamini spiritalia magis autem ut prophetetis
1COR|14|2|qui enim loquitur lingua non hominibus loquitur sed Deo nemo enim audit Spiritu autem loquitur mysteria
1COR|14|3|nam qui prophetat hominibus loquitur aedificationem et exhortationem et consolationes
1COR|14|4|qui loquitur lingua semet ipsum aedificat qui autem prophetat ecclesiam aedificat
1COR|14|5|volo autem omnes vos loqui linguis magis autem prophetare nam maior est qui prophetat quam qui loquitur linguis nisi si forte ut interpretetur ut ecclesia aedificationem accipiat
1COR|14|6|nunc autem fratres si venero ad vos linguis loquens quid vobis prodero nisi si vobis loquar aut in revelatione aut scientia aut prophetia aut in doctrina
1COR|14|7|tamen quae sine anima sunt vocem dantia sive tibia sive cithara nisi distinctionem sonituum dederint quomodo scietur quod canitur aut quod citharizatur
1COR|14|8|etenim si incertam vocem det tuba quis parabit se ad bellum
1COR|14|9|ita et vos per linguam nisi manifestum sermonem dederitis quomodo scietur id quod dicitur eritis enim in aera loquentes
1COR|14|10|tam multa ut puta genera linguarum sunt in mundo et nihil sine voce est
1COR|14|11|si ergo nesciero virtutem vocis ero ei cui loquor barbarus et qui loquitur mihi barbarus
1COR|14|12|sic et vos quoniam aemulatores estis spirituum ad aedificationem ecclesiae quaerite ut abundetis
1COR|14|13|et ideo qui loquitur lingua oret ut interpretetur
1COR|14|14|nam si orem lingua spiritus meus orat mens autem mea sine fructu est
1COR|14|15|quid ergo est orabo spiritu orabo et mente psallam spiritu psallam et mente
1COR|14|16|ceterum si benedixeris spiritu qui supplet locum idiotae quomodo dicet amen super tuam benedictionem quoniam quid dicas nescit
1COR|14|17|nam tu quidem bene gratias agis sed alter non aedificatur
1COR|14|18|gratias ago Deo quod omnium vestrum lingua loquor
1COR|14|19|sed in ecclesia volo quinque verba sensu meo loqui ut et alios instruam quam decem milia verborum in lingua
1COR|14|20|fratres nolite pueri effici sensibus sed malitia parvuli estote sensibus autem perfecti estote
1COR|14|21|in lege scriptum est quoniam in aliis linguis et labiis aliis loquar populo huic et nec sic exaudient me dicit Dominus
1COR|14|22|itaque linguae in signum sunt non fidelibus sed infidelibus prophetia autem non infidelibus sed fidelibus
1COR|14|23|si ergo conveniat universa ecclesia in unum et omnes linguis loquantur intrent autem idiotae aut infideles nonne dicent quod insanitis
1COR|14|24|si autem omnes prophetent intret autem quis infidelis vel idiota convincitur ab omnibus diiudicatur ab omnibus
1COR|14|25|occulta cordis eius manifesta fiunt et ita cadens in faciem adorabit Deum pronuntians quod vere Deus in vobis est
1COR|14|26|quid ergo est fratres cum convenitis unusquisque vestrum psalmum habet doctrinam habet apocalypsin habet linguam habet interpretationem habet omnia ad aedificationem fiant
1COR|14|27|sive lingua quis loquitur secundum duos aut ut multum tres et per partes et unus interpretetur
1COR|14|28|si autem non fuerit interpres taceat in ecclesia sibi autem loquatur et Deo
1COR|14|29|prophetae duo aut tres dicant et ceteri diiudicent
1COR|14|30|quod si alii revelatum fuerit sedenti prior taceat
1COR|14|31|potestis enim omnes per singulos prophetare ut omnes discant et omnes exhortentur
1COR|14|32|et spiritus prophetarum prophetis subiecti sunt
1COR|14|33|non enim est dissensionis Deus sed pacis sicut in omnibus ecclesiis sanctorum
1COR|14|34|mulieres in ecclesiis taceant non enim permittitur eis loqui sed subditas esse sicut et lex dicit
1COR|14|35|si quid autem volunt discere domi viros suos interrogent turpe est enim mulieri loqui in ecclesia
1COR|14|36|an a vobis verbum Dei processit aut in vos solos pervenit
1COR|14|37|si quis videtur propheta esse aut spiritalis cognoscat quae scribo vobis quia Domini sunt mandata
1COR|14|38|si quis autem ignorat ignorabitur
1COR|14|39|itaque fratres aemulamini prophetare et loqui linguis nolite prohibere
1COR|14|40|omnia autem honeste et secundum ordinem fiant
1COR|15|1|notum autem vobis facio fratres evangelium quod praedicavi vobis quod et accepistis in quo et statis
1COR|15|2|per quod et salvamini qua ratione praedicaverim vobis si tenetis nisi si frustra credidistis
1COR|15|3|tradidi enim vobis in primis quod et accepi quoniam Christus mortuus est pro peccatis nostris secundum scripturas
1COR|15|4|et quia sepultus est et quia resurrexit tertia die secundum scripturas
1COR|15|5|et quia visus est Cephae et post haec undecim
1COR|15|6|deinde visus est plus quam quingentis fratribus simul ex quibus multi manent usque adhuc quidam autem dormierunt
1COR|15|7|deinde visus est Iacobo deinde apostolis omnibus
1COR|15|8|novissime autem omnium tamquam abortivo visus est et mihi
1COR|15|9|ego enim sum minimus apostolorum qui non sum dignus vocari apostolus quoniam persecutus sum ecclesiam Dei
1COR|15|10|gratia autem Dei sum id quod sum et gratia eius in me vacua non fuit sed abundantius illis omnibus laboravi non ego autem sed gratia Dei mecum
1COR|15|11|sive enim ego sive illi sic praedicamus et sic credidistis
1COR|15|12|si autem Christus praedicatur quod resurrexit a mortuis quomodo quidam dicunt in vobis quoniam resurrectio mortuorum non est
1COR|15|13|si autem resurrectio mortuorum non est neque Christus resurrexit
1COR|15|14|si autem Christus non resurrexit inanis est ergo praedicatio nostra inanis est et fides vestra
1COR|15|15|invenimur autem et falsi testes Dei quoniam testimonium diximus adversus Deum quod suscitaverit Christum quem non suscitavit si mortui non resurgunt
1COR|15|16|nam si mortui non resurgunt neque Christus resurrexit
1COR|15|17|quod si Christus non resurrexit vana est fides vestra adhuc enim estis in peccatis vestris
1COR|15|18|ergo et qui dormierunt in Christo perierunt
1COR|15|19|si in hac vita tantum in Christo sperantes sumus miserabiliores sumus omnibus hominibus
1COR|15|20|nunc autem Christus resurrexit a mortuis primitiae dormientium
1COR|15|21|quoniam enim per hominem mors et per hominem resurrectio mortuorum
1COR|15|22|et sicut in Adam omnes moriuntur ita et in Christo omnes vivificabuntur
1COR|15|23|unusquisque autem in suo ordine primitiae Christus deinde hii qui sunt Christi in adventu eius
1COR|15|24|deinde finis cum tradiderit regnum Deo et Patri cum evacuaverit omnem principatum et potestatem et virtutem
1COR|15|25|oportet autem illum regnare donec ponat omnes inimicos sub pedibus eius
1COR|15|26|novissima autem inimica destruetur mors omnia enim subiecit sub pedibus eius cum autem dicat
1COR|15|27|omnia subiecta sunt sine dubio praeter eum qui subiecit ei omnia
1COR|15|28|cum autem subiecta fuerint illi omnia tunc ipse Filius subiectus erit illi qui sibi subiecit omnia ut sit Deus omnia in omnibus
1COR|15|29|alioquin quid facient qui baptizantur pro mortuis si omnino mortui non resurgunt ut quid et baptizantur pro illis
1COR|15|30|ut quid et nos periclitamur omni hora
1COR|15|31|cotidie morior per vestram gloriam fratres quam habeo in Christo Iesu Domino nostro
1COR|15|32|si secundum hominem ad bestias pugnavi Ephesi quid mihi prodest si mortui non resurgunt manducemus et bibamus cras enim moriemur
1COR|15|33|nolite seduci corrumpunt mores bonos conloquia mala
1COR|15|34|evigilate iuste et nolite peccare ignorantiam enim Dei quidam habent ad reverentiam vobis loquor
1COR|15|35|sed dicet aliquis quomodo resurgunt mortui quali autem corpore veniunt
1COR|15|36|insipiens tu quod seminas non vivificatur nisi prius moriatur
1COR|15|37|et quod seminas non corpus quod futurum est seminas sed nudum granum ut puta tritici aut alicuius ceterorum
1COR|15|38|Deus autem dat illi corpus sicut voluit et unicuique seminum proprium corpus
1COR|15|39|non omnis caro eadem caro sed alia hominum alia pecorum alia caro volucrum alia autem piscium
1COR|15|40|et corpora caelestia et corpora terrestria sed alia quidem caelestium gloria alia autem terrestrium
1COR|15|41|alia claritas solis alia claritas lunae et alia claritas stellarum stella enim ab stella differt in claritate
1COR|15|42|sic et resurrectio mortuorum seminatur in corruptione surgit in incorruptione
1COR|15|43|seminatur in ignobilitate surgit in gloria seminatur in infirmitate surgit in virtute
1COR|15|44|seminatur corpus animale surgit corpus spiritale si est corpus animale est et spiritale sic et scriptum est
1COR|15|45|factus est primus homo Adam in animam viventem novissimus Adam in spiritum vivificantem
1COR|15|46|sed non prius quod spiritale est sed quod animale est deinde quod spiritale
1COR|15|47|primus homo de terra terrenus secundus homo de caelo caelestis
1COR|15|48|qualis terrenus tales et terreni et qualis caelestis tales et caelestes
1COR|15|49|igitur sicut portavimus imaginem terreni portemus et imaginem caelestis
1COR|15|50|hoc autem dico fratres quoniam caro et sanguis regnum Dei possidere non possunt neque corruptio incorruptelam possidebit
1COR|15|51|ecce mysterium vobis dico omnes quidem resurgemus sed non omnes inmutabimur
1COR|15|52|in momento in ictu oculi in novissima tuba canet enim et mortui resurgent incorrupti et nos inmutabimur
1COR|15|53|oportet enim corruptibile hoc induere incorruptelam et mortale hoc induere inmortalitatem
1COR|15|54|cum autem mortale hoc induerit inmortalitatem tunc fiet sermo qui scriptus est absorta est mors in victoria
1COR|15|55|ubi est mors victoria tua ubi est mors stimulus tuus
1COR|15|56|stimulus autem mortis peccatum est virtus vero peccati lex
1COR|15|57|Deo autem gratias qui dedit nobis victoriam per Dominum nostrum Iesum Christum
1COR|15|58|itaque fratres mei dilecti stabiles estote et inmobiles abundantes in opere Domini semper scientes quod labor vester non est inanis in Domino
1COR|16|1|de collectis autem quae fiunt in sanctos sicut ordinavi ecclesiis Galatiae ita et vos facite
1COR|16|2|per unam sabbati unusquisque vestrum apud se ponat recondens quod ei beneplacuerit ut non cum venero tunc collectae fiant
1COR|16|3|cum autem praesens fuero quos probaveritis per epistulas hos mittam perferre gratiam vestram in Hierusalem
1COR|16|4|quod si dignum fuerit ut et ego eam mecum ibunt
1COR|16|5|veniam autem ad vos cum Macedoniam pertransiero nam Macedoniam pertransibo
1COR|16|6|apud vos autem forsitan manebo vel etiam hiemabo ut vos me deducatis quocumque iero
1COR|16|7|nolo enim vos modo in transitu videre spero enim me aliquantum temporis manere apud vos si Dominus permiserit
1COR|16|8|permanebo autem Ephesi usque ad pentecosten
1COR|16|9|ostium enim mihi apertum est magnum et evidens et adversarii multi
1COR|16|10|si autem venerit Timotheus videte ut sine timore sit apud vos opus enim Domini operatur sicut et ego
1COR|16|11|ne quis ergo illum spernat deducite autem illum in pace ut veniat ad me expecto enim illum cum fratribus
1COR|16|12|de Apollo autem fratre multum rogavi eum ut veniret ad vos cum fratribus et utique non fuit voluntas ut nunc veniret veniet autem cum ei vacuum fuerit
1COR|16|13|vigilate state in fide viriliter agite et confortamini
1COR|16|14|omnia vestra in caritate fiant
1COR|16|15|obsecro autem vos fratres nostis domum Stephanae et Fortunati quoniam sunt primitiae Achaiae et in ministerium sanctorum ordinaverunt se ipsos
1COR|16|16|ut et vos subditi sitis eiusmodi et omni cooperanti et laboranti
1COR|16|17|gaudeo autem in praesentia Stephanae et Fortunati et Achaici quoniam id quod vobis deerat ipsi suppleverunt
1COR|16|18|refecerunt enim et meum spiritum et vestrum cognoscite ergo qui eiusmodi sunt
1COR|16|19|salutant vos ecclesiae Asiae salutant vos in Domino multum Aquila et Prisca cum domestica sua ecclesia
1COR|16|20|salutant vos fratres omnes salutate invicem in osculo sancto
1COR|16|21|salutatio mea manu Pauli
1COR|16|22|si quis non amat Dominum Iesum Christum sit anathema maranatha
1COR|16|23|gratia Domini Iesu vobiscum
1COR|16|24|caritas mea cum omnibus vobis in Christo Iesu amen
