LUKE|1|1|Forasmuch as many have taken in hand to set forth in order a declaration of those things which are most surely believed among us,
LUKE|1|2|Even as they delivered them unto us, which from the beginning were eyewitnesses, and ministers of the word;
LUKE|1|3|It seemed good to me also, having had perfect understanding of all things from the very first, to write unto thee in order, most excellent Theophilus,
LUKE|1|4|That thou mightest know the certainty of those things, wherein thou hast been instructed.
LUKE|1|5|THERE was in the days of Herod, the king of Judaea, a certain priest named Zacharias, of the course of Abia: and his wife was of the daughters of Aaron, and her name was Elisabeth.
LUKE|1|6|And they were both righteous before God, walking in all the commandments and ordinances of the Lord blameless.
LUKE|1|7|And they had no child, because that Elisabeth was barren, and they both were now well stricken in years.
LUKE|1|8|And it came to pass, that while he executed the priest's office before God in the order of his course,
LUKE|1|9|According to the custom of the priest's office, his lot was to burn incense when he went into the temple of the Lord.
LUKE|1|10|And the whole multitude of the people were praying without at the time of incense.
LUKE|1|11|And there appeared unto him an angel of the Lord standing on the right side of the altar of incense.
LUKE|1|12|And when Zacharias saw him, he was troubled, and fear fell upon him.
LUKE|1|13|But the angel said unto him, Fear not, Zacharias: for thy prayer is heard; and thy wife Elisabeth shall bear thee a son, and thou shalt call his name John.
LUKE|1|14|And thou shalt have joy and gladness; and many shall rejoice at his birth.
LUKE|1|15|For he shall be great in the sight of the Lord, and shall drink neither wine nor strong drink; and he shall be filled with the Holy Ghost, even from his mother's womb.
LUKE|1|16|And many of the children of Israel shall he turn to the Lord their God.
LUKE|1|17|And he shall go before him in the spirit and power of Elias, to turn the hearts of the fathers to the children, and the disobedient to the wisdom of the just; to make ready a people prepared for the Lord.
LUKE|1|18|And Zacharias said unto the angel, Whereby shall I know this? for I am an old man, and my wife well stricken in years.
LUKE|1|19|And the angel answering said unto him, I am Gabriel, that stand in the presence of God; and am sent to speak unto thee, and to shew thee these glad tidings.
LUKE|1|20|And, behold, thou shalt be dumb, and not able to speak, until the day that these things shall be performed, because thou believest not my words, which shall be fulfilled in their season.
LUKE|1|21|And the people waited for Zacharias, and marvelled that he tarried so long in the temple.
LUKE|1|22|And when he came out, he could not speak unto them: and they perceived that he had seen a vision in the temple: for he beckoned unto them, and remained speechless.
LUKE|1|23|And it came to pass, that, as soon as the days of his ministration were accomplished, he departed to his own house.
LUKE|1|24|And after those days his wife Elisabeth conceived, and hid herself five months, saying,
LUKE|1|25|Thus hath the Lord dealt with me in the days wherein he looked on me, to take away my reproach among men.
LUKE|1|26|And in the sixth month the angel Gabriel was sent from God unto a city of Galilee, named Nazareth,
LUKE|1|27|To a virgin espoused to a man whose name was Joseph, of the house of David; and the virgin's name was Mary.
LUKE|1|28|And the angel came in unto her, and said, Hail, thou that art highly favoured, the Lord is with thee: blessed art thou among women.
LUKE|1|29|And when she saw him, she was troubled at his saying, and cast in her mind what manner of salutation this should be.
LUKE|1|30|And the angel said unto her, Fear not, Mary: for thou hast found favour with God.
LUKE|1|31|And, behold, thou shalt conceive in thy womb, and bring forth a son, and shalt call his name JESUS.
LUKE|1|32|He shall be great, and shall be called the Son of the Highest: and the Lord God shall give unto him the throne of his father David:
LUKE|1|33|And he shall reign over the house of Jacob for ever; and of his kingdom there shall be no end.
LUKE|1|34|Then said Mary unto the angel, How shall this be, seeing I know not a man?
LUKE|1|35|And the angel answered and said unto her, The Holy Ghost shall come upon thee, and the power of the Highest shall overshadow thee: therefore also that holy thing which shall be born of thee shall be called the Son of God.
LUKE|1|36|And, behold, thy cousin Elisabeth, she hath also conceived a son in her old age: and this is the sixth month with her, who was called barren.
LUKE|1|37|For with God nothing shall be impossible.
LUKE|1|38|And Mary said, Behold the handmaid of the Lord; be it unto me according to thy word. And the angel departed from her.
LUKE|1|39|And Mary arose in those days, and went into the hill country with haste, into a city of Juda;
LUKE|1|40|And entered into the house of Zacharias, and saluted Elisabeth.
LUKE|1|41|And it came to pass, that, when Elisabeth heard the salutation of Mary, the babe leaped in her womb; and Elisabeth was filled with the Holy Ghost:
LUKE|1|42|And she spake out with a loud voice, and said, Blessed art thou among women, and blessed is the fruit of thy womb.
LUKE|1|43|And whence is this to me, that the mother of my Lord should come to me?
LUKE|1|44|For, lo, as soon as the voice of thy salutation sounded in mine ears, the babe leaped in my womb for joy.
LUKE|1|45|And blessed is she that believed: for there shall be a performance of those things which were told her from the Lord.
LUKE|1|46|And Mary said, My soul doth magnify the Lord,
LUKE|1|47|And my spirit hath rejoiced in God my Saviour.
LUKE|1|48|For he hath regarded the low estate of his handmaiden: for, behold, from henceforth all generations shall call me blessed.
LUKE|1|49|For he that is mighty hath done to me great things; and holy is his name.
LUKE|1|50|And his mercy is on them that fear him from generation to generation.
LUKE|1|51|He hath shewed strength with his arm; he hath scattered the proud in the imagination of their hearts.
LUKE|1|52|He hath put down the mighty from their seats, and exalted them of low degree.
LUKE|1|53|He hath filled the hungry with good things; and the rich he hath sent empty away.
LUKE|1|54|He hath holpen his servant Israel, in remembrance of his mercy;
LUKE|1|55|As he spake to our fathers, to Abraham, and to his seed for ever.
LUKE|1|56|And Mary abode with her about three months, and returned to her own house.
LUKE|1|57|Now Elisabeth's full time came that she should be delivered; and she brought forth a son.
LUKE|1|58|And her neighbours and her cousins heard how the Lord had shewed great mercy upon her; and they rejoiced with her.
LUKE|1|59|And it came to pass, that on the eighth day they came to circumcise the child; and they called him Zacharias, after the name of his father.
LUKE|1|60|And his mother answered and said, Not so; but he shall be called John.
LUKE|1|61|And they said unto her, There is none of thy kindred that is called by this name.
LUKE|1|62|And they made signs to his father, how he would have him called.
LUKE|1|63|And he asked for a writing table, and wrote, saying, His name is John. And they marvelled all.
LUKE|1|64|And his mouth was opened immediately, and his tongue loosed, and he spake, and praised God.
LUKE|1|65|And fear came on all that dwelt round about them: and all these sayings were noised abroad throughout all the hill country of Judaea.
LUKE|1|66|And all they that heard them laid them up in their hearts, saying, What manner of child shall this be! And the hand of the Lord was with him.
LUKE|1|67|And his father Zacharias was filled with the Holy Ghost, and prophesied, saying,
LUKE|1|68|Blessed be the Lord God of Israel; for he hath visited and redeemed his people,
LUKE|1|69|And hath raised up an horn of salvation for us in the house of his servant David;
LUKE|1|70|As he spake by the mouth of his holy prophets, which have been since the world began:
LUKE|1|71|That we should be saved from our enemies, and from the hand of all that hate us;
LUKE|1|72|To perform the mercy promised to our fathers, and to remember his holy covenant;
LUKE|1|73|The oath which he sware to our father Abraham,
LUKE|1|74|That he would grant unto us, that we being delivered out of the hand of our enemies might serve him without fear,
LUKE|1|75|In holiness and righteousness before him, all the days of our life.
LUKE|1|76|And thou, child, shalt be called the prophet of the Highest: for thou shalt go before the face of the Lord to prepare his ways;
LUKE|1|77|To give knowledge of salvation unto his people by the remission of their sins,
LUKE|1|78|Through the tender mercy of our God; whereby the dayspring from on high hath visited us,
LUKE|1|79|To give light to them that sit in darkness and in the shadow of death, to guide our feet into the way of peace.
LUKE|1|80|And the child grew, and waxed strong in spirit, and was in the deserts till the day of his shewing unto Israel.
LUKE|2|1|And it came to pass in those days, that there went out a decree from Caesar Augustus that all the world should be taxed.
LUKE|2|2|(And this taxing was first made when Cyrenius was governor of Syria.)
LUKE|2|3|And all went to be taxed, every one into his own city.
LUKE|2|4|And Joseph also went up from Galilee, out of the city of Nazareth, into Judaea, unto the city of David, which is called Bethlehem; (because he was of the house and lineage of David:)
LUKE|2|5|To be taxed with Mary his espoused wife, being great with child.
LUKE|2|6|And so it was, that, while they were there, the days were accomplished that she should be delivered.
LUKE|2|7|And she brought forth her firstborn son, and wrapped him in swaddling clothes, and laid him in a manger; because there was no room for them in the inn.
LUKE|2|8|And there were in the same country shepherds abiding in the field, keeping watch over their flock by night.
LUKE|2|9|And, lo, the angel of the Lord came upon them, and the glory of the Lord shone round about them: and they were sore afraid.
LUKE|2|10|And the angel said unto them, Fear not: for, behold, I bring you good tidings of great joy, which shall be to all people.
LUKE|2|11|For unto you is born this day in the city of David a Saviour, which is Christ the Lord.
LUKE|2|12|And this shall be a sign unto you; Ye shall find the babe wrapped in swaddling clothes, lying in a manger.
LUKE|2|13|And suddenly there was with the angel a multitude of the heavenly host praising God, and saying,
LUKE|2|14|Glory to God in the highest, and on earth peace, good will toward men.
LUKE|2|15|And it came to pass, as the angels were gone away from them into heaven, the shepherds said one to another, Let us now go even unto Bethlehem, and see this thing which is come to pass, which the Lord hath made known unto us.
LUKE|2|16|And they came with haste, and found Mary, and Joseph, and the babe lying in a manger.
LUKE|2|17|And when they had seen it, they made known abroad the saying which was told them concerning this child.
LUKE|2|18|And all they that heard it wondered at those things which were told them by the shepherds.
LUKE|2|19|But Mary kept all these things, and pondered them in her heart.
LUKE|2|20|And the shepherds returned, glorifying and praising God for all the things that they had heard and seen, as it was told unto them.
LUKE|2|21|And when eight days were accomplished for the circumcising of the child, his name was called JESUS, which was so named of the angel before he was conceived in the womb.
LUKE|2|22|And when the days of her purification according to the law of Moses were accomplished, they brought him to Jerusalem, to present him to the Lord;
LUKE|2|23|(As it is written in the law of the LORD, Every male that openeth the womb shall be called holy to the Lord;)
LUKE|2|24|And to offer a sacrifice according to that which is said in the law of the Lord, A pair of turtledoves, or two young pigeons.
LUKE|2|25|And, behold, there was a man in Jerusalem, whose name was Simeon; and the same man was just and devout, waiting for the consolation of Israel: and the Holy Ghost was upon him.
LUKE|2|26|And it was revealed unto him by the Holy Ghost, that he should not see death, before he had seen the Lord's Christ.
LUKE|2|27|And he came by the Spirit into the temple: and when the parents brought in the child Jesus, to do for him after the custom of the law,
LUKE|2|28|Then took he him up in his arms, and blessed God, and said,
LUKE|2|29|Lord, now lettest thou thy servant depart in peace, according to thy word:
LUKE|2|30|For mine eyes have seen thy salvation,
LUKE|2|31|Which thou hast prepared before the face of all people;
LUKE|2|32|A light to lighten the Gentiles, and the glory of thy people Israel.
LUKE|2|33|And Joseph and his mother marvelled at those things which were spoken of him.
LUKE|2|34|And Simeon blessed them, and said unto Mary his mother, Behold, this child is set for the fall and rising again of many in Israel; and for a sign which shall be spoken against;
LUKE|2|35|(Yea, a sword shall pierce through thy own soul also,) that the thoughts of many hearts may be revealed.
LUKE|2|36|And there was one Anna, a prophetess, the daughter of Phanuel, of the tribe of Aser: she was of a great age, and had lived with an husband seven years from her virginity;
LUKE|2|37|And she was a widow of about fourscore and four years, which departed not from the temple, but served God with fastings and prayers night and day.
LUKE|2|38|And she coming in that instant gave thanks likewise unto the Lord, and spake of him to all them that looked for redemption in Jerusalem.
LUKE|2|39|And when they had performed all things according to the law of the Lord, they returned into Galilee, to their own city Nazareth.
LUKE|2|40|And the child grew, and waxed strong in spirit, filled with wisdom: and the grace of God was upon him.
LUKE|2|41|Now his parents went to Jerusalem every year at the feast of the passover.
LUKE|2|42|And when he was twelve years old, they went up to Jerusalem after the custom of the feast.
LUKE|2|43|And when they had fulfilled the days, as they returned, the child Jesus tarried behind in Jerusalem; and Joseph and his mother knew not of it.
LUKE|2|44|But they, supposing him to have been in the company, went a day's journey; and they sought him among their kinsfolk and acquaintance.
LUKE|2|45|And when they found him not, they turned back again to Jerusalem, seeking him.
LUKE|2|46|And it came to pass, that after three days they found him in the temple, sitting in the midst of the doctors, both hearing them, and asking them questions.
LUKE|2|47|And all that heard him were astonished at his understanding and answers.
LUKE|2|48|And when they saw him, they were amazed: and his mother said unto him, Son, why hast thou thus dealt with us? behold, thy father and I have sought thee sorrowing.
LUKE|2|49|And he said unto them, How is it that ye sought me? wist ye not that I must be about my Father's business?
LUKE|2|50|And they understood not the saying which he spake unto them.
LUKE|2|51|And he went down with them, and came to Nazareth, and was subject unto them: but his mother kept all these sayings in her heart.
LUKE|2|52|And Jesus increased in wisdom and stature, and in favour with God and man.
LUKE|3|1|Now in the fifteenth year of the reign of Tiberius Caesar, Pontius Pilate being governor of Judaea, and Herod being tetrarch of Galilee, and his brother Philip tetrarch of Ituraea and of the region of Trachonitis, and Lysanias the tetrarch of Abilene,
LUKE|3|2|Annas and Caiaphas being the high priests, the word of God came unto John the son of Zacharias in the wilderness.
LUKE|3|3|And he came into all the country about Jordan, preaching the baptism of repentance for the remission of sins;
LUKE|3|4|As it is written in the book of the words of Esaias the prophet, saying, The voice of one crying in the wilderness, Prepare ye the way of the Lord, make his paths straight.
LUKE|3|5|Every valley shall be filled, and every mountain and hill shall be brought low; and the crooked shall be made straight, and the rough ways shall be made smooth;
LUKE|3|6|And all flesh shall see the salvation of God.
LUKE|3|7|Then said he to the multitude that came forth to be baptized of him, O generation of vipers, who hath warned you to flee from the wrath to come?
LUKE|3|8|Bring forth therefore fruits worthy of repentance, and begin not to say within yourselves, We have Abraham to our father: for I say unto you, That God is able of these stones to raise up children unto Abraham.
LUKE|3|9|And now also the axe is laid unto the root of the trees: every tree therefore which bringeth not forth good fruit is hewn down, and cast into the fire.
LUKE|3|10|And the people asked him, saying, What shall we do then?
LUKE|3|11|He answereth and saith unto them, He that hath two coats, let him impart to him that hath none; and he that hath meat, let him do likewise.
LUKE|3|12|Then came also publicans to be baptized, and said unto him, Master, what shall we do?
LUKE|3|13|And he said unto them, Exact no more than that which is appointed you.
LUKE|3|14|And the soldiers likewise demanded of him, saying, And what shall we do? And he said unto them, Do violence to no man, neither accuse any falsely; and be content with your wages.
LUKE|3|15|And as the people were in expectation, and all men mused in their hearts of John, whether he were the Christ, or not;
LUKE|3|16|John answered, saying unto them all, I indeed baptize you with water; but one mightier than I cometh, the latchet of whose shoes I am not worthy to unloose: he shall baptize you with the Holy Ghost and with fire:
LUKE|3|17|Whose fan is in his hand, and he will throughly purge his floor, and will gather the wheat into his garner; but the chaff he will burn with fire unquenchable.
LUKE|3|18|And many other things in his exhortation preached he unto the people.
LUKE|3|19|But Herod the tetrarch, being reproved by him for Herodias his brother Philip's wife, and for all the evils which Herod had done,
LUKE|3|20|Added yet this above all, that he shut up John in prison.
LUKE|3|21|Now when all the people were baptized, it came to pass, that Jesus also being baptized, and praying, the heaven was opened,
LUKE|3|22|And the Holy Ghost descended in a bodily shape like a dove upon him, and a voice came from heaven, which said, Thou art my beloved Son; in thee I am well pleased.
LUKE|3|23|And Jesus himself began to be about thirty years of age, being (as was supposed) the son of Joseph, which was the son of Heli,
LUKE|3|24|Which was the son of Matthat, which was the son of Levi, which was the son of Melchi, which was the son of Janna, which was the son of Joseph,
LUKE|3|25|Which was the son of Mattathias, which was the son of Amos, which was the son of Naum, which was the son of Esli, which was the son of Nagge,
LUKE|3|26|Which was the son of Maath, which was the son of Mattathias, which was the son of Semei, which was the son of Joseph, which was the son of Juda,
LUKE|3|27|Which was the son of Joanna, which was the son of Rhesa, which was the son of Zorobabel, which was the son of Salathiel, which was the son of Neri,
LUKE|3|28|Which was the son of Melchi, which was the son of Addi, which was the son of Cosam, which was the son of Elmodam, which was the son of Er,
LUKE|3|29|Which was the son of Jose, which was the son of Eliezer, which was the son of Jorim, which was the son of Matthat, which was the son of Levi,
LUKE|3|30|Which was the son of Simeon, which was the son of Juda, which was the son of Joseph, which was the son of Jonan, which was the son of Eliakim,
LUKE|3|31|Which was the son of Melea, which was the son of Menan, which was the son of Mattatha, which was the son of Nathan, which was the son of David,
LUKE|3|32|Which was the son of Jesse, which was the son of Obed, which was the son of Booz, which was the son of Salmon, which was the son of Naasson,
LUKE|3|33|Which was the son of Aminadab, which was the son of Aram, which was the son of Esrom, which was the son of Phares, which was the son of Juda,
LUKE|3|34|Which was the son of Jacob, which was the son of Isaac, which was the son of Abraham, which was the son of Thara, which was the son of Nachor,
LUKE|3|35|Which was the son of Saruch, which was the son of Ragau, which was the son of Phalec, which was the son of Heber, which was the son of Sala,
LUKE|3|36|Which was the son of Cainan, which was the son of Arphaxad, which was the son of Sem, which was the son of Noe, which was the son of Lamech,
LUKE|3|37|Which was the son of Mathusala, which was the son of Enoch, which was the son of Jared, which was the son of Maleleel, which was the son of Cainan,
LUKE|3|38|Which was the son of Enos, which was the son of Seth, which was the son of Adam, which was the son of God.
LUKE|4|1|And Jesus being full of the Holy Ghost returned from Jordan, and was led by the Spirit into the wilderness,
LUKE|4|2|Being forty days tempted of the devil. And in those days he did eat nothing: and when they were ended, he afterward hungered.
LUKE|4|3|And the devil said unto him, If thou be the Son of God, command this stone that it be made bread.
LUKE|4|4|And Jesus answered him, saying, It is written, That man shall not live by bread alone, but by every word of God.
LUKE|4|5|And the devil, taking him up into an high mountain, shewed unto him all the kingdoms of the world in a moment of time.
LUKE|4|6|And the devil said unto him, All this power will I give thee, and the glory of them: for that is delivered unto me; and to whomsoever I will I give it.
LUKE|4|7|If thou therefore wilt worship me, all shall be thine.
LUKE|4|8|And Jesus answered and said unto him, Get thee behind me, Satan: for it is written, Thou shalt worship the Lord thy God, and him only shalt thou serve.
LUKE|4|9|And he brought him to Jerusalem, and set him on a pinnacle of the temple, and said unto him, If thou be the Son of God, cast thyself down from hence:
LUKE|4|10|For it is written, He shall give his angels charge over thee, to keep thee:
LUKE|4|11|And in their hands they shall bear thee up, lest at any time thou dash thy foot against a stone.
LUKE|4|12|And Jesus answering said unto him, It is said, Thou shalt not tempt the Lord thy God.
LUKE|4|13|And when the devil had ended all the temptation, he departed from him for a season.
LUKE|4|14|And Jesus returned in the power of the Spirit into Galilee: and there went out a fame of him through all the region round about.
LUKE|4|15|And he taught in their synagogues, being glorified of all.
LUKE|4|16|And he came to Nazareth, where he had been brought up: and, as his custom was, he went into the synagogue on the sabbath day, and stood up for to read.
LUKE|4|17|And there was delivered unto him the book of the prophet Esaias. And when he had opened the book, he found the place where it was written,
LUKE|4|18|The Spirit of the Lord is upon me, because he hath anointed me to preach the gospel to the poor; he hath sent me to heal the brokenhearted, to preach deliverance to the captives, and recovering of sight to the blind, to set at liberty them that are bruised,
LUKE|4|19|To preach the acceptable year of the Lord.
LUKE|4|20|And he closed the book, and he gave it again to the minister, and sat down. And the eyes of all them that were in the synagogue were fastened on him.
LUKE|4|21|And he began to say unto them, This day is this scripture fulfilled in your ears.
LUKE|4|22|And all bare him witness, and wondered at the gracious words which proceeded out of his mouth. And they said, Is not this Joseph's son?
LUKE|4|23|And he said unto them, Ye will surely say unto me this proverb, Physician, heal thyself: whatsoever we have heard done in Capernaum, do also here in thy country.
LUKE|4|24|And he said, Verily I say unto you, No prophet is accepted in his own country.
LUKE|4|25|But I tell you of a truth, many widows were in Israel in the days of Elias, when the heaven was shut up three years and six months, when great famine was throughout all the land;
LUKE|4|26|But unto none of them was Elias sent, save unto Sarepta, a city of Sidon, unto a woman that was a widow.
LUKE|4|27|And many lepers were in Israel in the time of Eliseus the prophet; and none of them was cleansed, saving Naaman the Syrian.
LUKE|4|28|And all they in the synagogue, when they heard these things, were filled with wrath,
LUKE|4|29|And rose up, and thrust him out of the city, and led him unto the brow of the hill whereon their city was built, that they might cast him down headlong.
LUKE|4|30|But he passing through the midst of them went his way,
LUKE|4|31|And came down to Capernaum, a city of Galilee, and taught them on the sabbath days.
LUKE|4|32|And they were astonished at his doctrine: for his word was with power.
LUKE|4|33|And in the synagogue there was a man, which had a spirit of an unclean devil, and cried out with a loud voice,
LUKE|4|34|Saying, Let us alone; what have we to do with thee, thou Jesus of Nazareth? art thou come to destroy us? I know thee who thou art; the Holy One of God.
LUKE|4|35|And Jesus rebuked him, saying, Hold thy peace, and come out of him. And when the devil had thrown him in the midst, he came out of him, and hurt him not.
LUKE|4|36|And they were all amazed, and spake among themselves, saying, What a word is this! for with authority and power he commandeth the unclean spirits, and they come out.
LUKE|4|37|And the fame of him went out into every place of the country round about.
LUKE|4|38|And he arose out of the synagogue, and entered into Simon's house. And Simon's wife's mother was taken with a great fever; and they besought him for her.
LUKE|4|39|And he stood over her, and rebuked the fever; and it left her: and immediately she arose and ministered unto them.
LUKE|4|40|Now when the sun was setting, all they that had any sick with divers diseases brought them unto him; and he laid his hands on every one of them, and healed them.
LUKE|4|41|And devils also came out of many, crying out, and saying, Thou art Christ the Son of God. And he rebuking them suffered them not to speak: for they knew that he was Christ.
LUKE|4|42|And when it was day, he departed and went into a desert place: and the people sought him, and came unto him, and stayed him, that he should not depart from them.
LUKE|4|43|And he said unto them, I must preach the kingdom of God to other cities also: for therefore am I sent.
LUKE|4|44|And he preached in the synagogues of Galilee.
LUKE|5|1|And it came to pass, that, as the people pressed upon him to hear the word of God, he stood by the lake of Gennesaret,
LUKE|5|2|And saw two ships standing by the lake: but the fishermen were gone out of them, and were washing their nets.
LUKE|5|3|And he entered into one of the ships, which was Simon's, and prayed him that he would thrust out a little from the land. And he sat down, and taught the people out of the ship.
LUKE|5|4|Now when he had left speaking, he said unto Simon, Launch out into the deep, and let down your nets for a draught.
LUKE|5|5|And Simon answering said unto him, Master, we have toiled all the night, and have taken nothing: nevertheless at thy word I will let down the net.
LUKE|5|6|And when they had this done, they inclosed a great multitude of fishes: and their net brake.
LUKE|5|7|And they beckoned unto their partners, which were in the other ship, that they should come and help them. And they came, and filled both the ships, so that they began to sink.
LUKE|5|8|When Simon Peter saw it, he fell down at Jesus' knees, saying, Depart from me; for I am a sinful man, O Lord.
LUKE|5|9|For he was astonished, and all that were with him, at the draught of the fishes which they had taken:
LUKE|5|10|And so was also James, and John, the sons of Zebedee, which were partners with Simon. And Jesus said unto Simon, Fear not; from henceforth thou shalt catch men.
LUKE|5|11|And when they had brought their ships to land, they forsook all, and followed him.
LUKE|5|12|And it came to pass, when he was in a certain city, behold a man full of leprosy: who seeing Jesus fell on his face, and besought him, saying, Lord, if thou wilt, thou canst make me clean.
LUKE|5|13|And he put forth his hand, and touched him, saying, I will: be thou clean. And immediately the leprosy departed from him.
LUKE|5|14|And he charged him to tell no man: but go, and shew thyself to the priest, and offer for thy cleansing, according as Moses commanded, for a testimony unto them.
LUKE|5|15|But so much the more went there a fame abroad of him: and great multitudes came together to hear, and to be healed by him of their infirmities.
LUKE|5|16|And he withdrew himself into the wilderness, and prayed.
LUKE|5|17|And it came to pass on a certain day, as he was teaching, that there were Pharisees and doctors of the law sitting by, which were come out of every town of Galilee, and Judaea, and Jerusalem: and the power of the Lord was present to heal them.
LUKE|5|18|And, behold, men brought in a bed a man which was taken with a palsy: and they sought means to bring him in, and to lay him before him.
LUKE|5|19|And when they could not find by what way they might bring him in because of the multitude, they went upon the housetop, and let him down through the tiling with his couch into the midst before Jesus.
LUKE|5|20|And when he saw their faith, he said unto him, Man, thy sins are forgiven thee.
LUKE|5|21|And the scribes and the Pharisees began to reason, saying, Who is this which speaketh blasphemies? Who can forgive sins, but God alone?
LUKE|5|22|But when Jesus perceived their thoughts, he answering said unto them, What reason ye in your hearts?
LUKE|5|23|Whether is easier, to say, Thy sins be forgiven thee; or to say, Rise up and walk?
LUKE|5|24|But that ye may know that the Son of man hath power upon earth to forgive sins, (he said unto the sick of the palsy,) I say unto thee, Arise, and take up thy couch, and go into thine house.
LUKE|5|25|And immediately he rose up before them, and took up that whereon he lay, and departed to his own house, glorifying God.
LUKE|5|26|And they were all amazed, and they glorified God, and were filled with fear, saying, We have seen strange things to day.
LUKE|5|27|And after these things he went forth, and saw a publican, named Levi, sitting at the receipt of custom: and he said unto him, Follow me.
LUKE|5|28|And he left all, rose up, and followed him.
LUKE|5|29|And Levi made him a great feast in his own house: and there was a great company of publicans and of others that sat down with them.
LUKE|5|30|But their scribes and Pharisees murmured against his disciples, saying, Why do ye eat and drink with publicans and sinners?
LUKE|5|31|And Jesus answering said unto them, They that are whole need not a physician; but they that are sick.
LUKE|5|32|I came not to call the righteous, but sinners to repentance.
LUKE|5|33|And they said unto him, Why do the disciples of John fast often, and make prayers, and likewise the disciples of the Pharisees; but thine eat and drink?
LUKE|5|34|And he said unto them, Can ye make the children of the bridechamber fast, while the bridegroom is with them?
LUKE|5|35|But the days will come, when the bridegroom shall be taken away from them, and then shall they fast in those days.
LUKE|5|36|And he spake also a parable unto them; No man putteth a piece of a new garment upon an old; if otherwise, then both the new maketh a rent, and the piece that was taken out of the new agreeth not with the old.
LUKE|5|37|And no man putteth new wine into old bottles; else the new wine will burst the bottles, and be spilled, and the bottles shall perish.
LUKE|5|38|But new wine must be put into new bottles; and both are preserved.
LUKE|5|39|No man also having drunk old wine straightway desireth new: for he saith, The old is better.
LUKE|6|1|And it came to pass on the second sabbath after the first, that he went through the corn fields; and his disciples plucked the ears of corn, and did eat, rubbing them in their hands.
LUKE|6|2|And certain of the Pharisees said unto them, Why do ye that which is not lawful to do on the sabbath days?
LUKE|6|3|And Jesus answering them said, Have ye not read so much as this, what David did, when himself was an hungred, and they which were with him;
LUKE|6|4|How he went into the house of God, and did take and eat the shewbread, and gave also to them that were with him; which it is not lawful to eat but for the priests alone?
LUKE|6|5|And he said unto them, That the Son of man is Lord also of the sabbath.
LUKE|6|6|And it came to pass also on another sabbath, that he entered into the synagogue and taught: and there was a man whose right hand was withered.
LUKE|6|7|And the scribes and Pharisees watched him, whether he would heal on the sabbath day; that they might find an accusation against him.
LUKE|6|8|But he knew their thoughts, and said to the man which had the withered hand, Rise up, and stand forth in the midst. And he arose and stood forth.
LUKE|6|9|Then said Jesus unto them, I will ask you one thing; Is it lawful on the sabbath days to do good, or to do evil? to save life, or to destroy it?
LUKE|6|10|And looking round about upon them all, he said unto the man, Stretch forth thy hand. And he did so: and his hand was restored whole as the other.
LUKE|6|11|And they were filled with madness; and communed one with another what they might do to Jesus.
LUKE|6|12|And it came to pass in those days, that he went out into a mountain to pray, and continued all night in prayer to God.
LUKE|6|13|And when it was day, he called unto him his disciples: and of them he chose twelve, whom also he named apostles;
LUKE|6|14|Simon, (whom he also named Peter,) and Andrew his brother, James and John, Philip and Bartholomew,
LUKE|6|15|Matthew and Thomas, James the son of Alphaeus, and Simon called Zelotes,
LUKE|6|16|And Judas the brother of James, and Judas Iscariot, which also was the traitor.
LUKE|6|17|And he came down with them, and stood in the plain, and the company of his disciples, and a great multitude of people out of all Judaea and Jerusalem, and from the sea coast of Tyre and Sidon, which came to hear him, and to be healed of their diseases;
LUKE|6|18|And they that were vexed with unclean spirits: and they were healed.
LUKE|6|19|And the whole multitude sought to touch him: for there went virtue out of him, and healed them all.
LUKE|6|20|And he lifted up his eyes on his disciples, and said, Blessed be ye poor: for yours is the kingdom of God.
LUKE|6|21|Blessed are ye that hunger now: for ye shall be filled. Blessed are ye that weep now: for ye shall laugh.
LUKE|6|22|Blessed are ye, when men shall hate you, and when they shall separate you from their company, and shall reproach you, and cast out your name as evil, for the Son of man's sake.
LUKE|6|23|Rejoice ye in that day, and leap for joy: for, behold, your reward is great in heaven: for in the like manner did their fathers unto the prophets.
LUKE|6|24|But woe unto you that are rich! for ye have received your consolation.
LUKE|6|25|Woe unto you that are full! for ye shall hunger. Woe unto you that laugh now! for ye shall mourn and weep.
LUKE|6|26|Woe unto you, when all men shall speak well of you! for so did their fathers to the false prophets.
LUKE|6|27|But I say unto you which hear, Love your enemies, do good to them which hate you,
LUKE|6|28|Bless them that curse you, and pray for them which despitefully use you.
LUKE|6|29|And unto him that smiteth thee on the one cheek offer also the other; and him that taketh away thy cloak forbid not to take thy coat also.
LUKE|6|30|Give to every man that asketh of thee; and of him that taketh away thy goods ask them not again.
LUKE|6|31|And as ye would that men should do to you, do ye also to them likewise.
LUKE|6|32|For if ye love them which love you, what thank have ye? for sinners also love those that love them.
LUKE|6|33|And if ye do good to them which do good to you, what thank have ye? for sinners also do even the same.
LUKE|6|34|And if ye lend to them of whom ye hope to receive, what thank have ye? for sinners also lend to sinners, to receive as much again.
LUKE|6|35|But love ye your enemies, and do good, and lend, hoping for nothing again; and your reward shall be great, and ye shall be the children of the Highest: for he is kind unto the unthankful and to the evil.
LUKE|6|36|Be ye therefore merciful, as your Father also is merciful.
LUKE|6|37|Judge not, and ye shall not be judged: condemn not, and ye shall not be condemned: forgive, and ye shall be forgiven:
LUKE|6|38|Give, and it shall be given unto you; good measure, pressed down, and shaken together, and running over, shall men give into your bosom. For with the same measure that ye mete withal it shall be measured to you again.
LUKE|6|39|And he spake a parable unto them, Can the blind lead the blind? shall they not both fall into the ditch?
LUKE|6|40|The disciple is not above his master: but every one that is perfect shall be as his master.
LUKE|6|41|And why beholdest thou the mote that is in thy brother's eye, but perceivest not the beam that is in thine own eye?
LUKE|6|42|Either how canst thou say to thy brother, Brother, let me pull out the mote that is in thine eye, when thou thyself beholdest not the beam that is in thine own eye? Thou hypocrite, cast out first the beam out of thine own eye, and then shalt thou see clearly to pull out the mote that is in thy brother's eye.
LUKE|6|43|For a good tree bringeth not forth corrupt fruit; neither doth a corrupt tree bring forth good fruit.
LUKE|6|44|For every tree is known by his own fruit. For of thorns men do not gather figs, nor of a bramble bush gather they grapes.
LUKE|6|45|A good man out of the good treasure of his heart bringeth forth that which is good; and an evil man out of the evil treasure of his heart bringeth forth that which is evil: for of the abundance of the heart his mouth speaketh.
LUKE|6|46|And why call ye me, Lord, Lord, and do not the things which I say?
LUKE|6|47|Whosoever cometh to me, and heareth my sayings, and doeth them, I will shew you to whom he is like:
LUKE|6|48|He is like a man which built an house, and digged deep, and laid the foundation on a rock: and when the flood arose, the stream beat vehemently upon that house, and could not shake it: for it was founded upon a rock.
LUKE|6|49|But he that heareth, and doeth not, is like a man that without a foundation built an house upon the earth; against which the stream did beat vehemently, and immediately it fell; and the ruin of that house was great.
LUKE|7|1|Now when he had ended all his sayings in the audience of the people, he entered into Capernaum.
LUKE|7|2|And a certain centurion's servant, who was dear unto him, was sick, and ready to die.
LUKE|7|3|And when he heard of Jesus, he sent unto him the elders of the Jews, beseeching him that he would come and heal his servant.
LUKE|7|4|And when they came to Jesus, they besought him instantly, saying, That he was worthy for whom he should do this:
LUKE|7|5|For he loveth our nation, and he hath built us a synagogue.
LUKE|7|6|Then Jesus went with them. And when he was now not far from the house, the centurion sent friends to him, saying unto him, Lord, trouble not thyself: for I am not worthy that thou shouldest enter under my roof:
LUKE|7|7|Wherefore neither thought I myself worthy to come unto thee: but say in a word, and my servant shall be healed.
LUKE|7|8|For I also am a man set under authority, having under me soldiers, and I say unto one, Go, and he goeth; and to another, Come, and he cometh; and to my servant, Do this, and he doeth it.
LUKE|7|9|When Jesus heard these things, he marvelled at him, and turned him about, and said unto the people that followed him, I say unto you, I have not found so great faith, no, not in Israel.
LUKE|7|10|And they that were sent, returning to the house, found the servant whole that had been sick.
LUKE|7|11|And it came to pass the day after, that he went into a city called Nain; and many of his disciples went with him, and much people.
LUKE|7|12|Now when he came nigh to the gate of the city, behold, there was a dead man carried out, the only son of his mother, and she was a widow: and much people of the city was with her.
LUKE|7|13|And when the Lord saw her, he had compassion on her, and said unto her, Weep not.
LUKE|7|14|And he came and touched the bier: and they that bare him stood still. And he said, Young man, I say unto thee, Arise.
LUKE|7|15|And he that was dead sat up, and began to speak. And he delivered him to his mother.
LUKE|7|16|And there came a fear on all: and they glorified God, saying, That a great prophet is risen up among us; and, That God hath visited his people.
LUKE|7|17|And this rumour of him went forth throughout all Judaea, and throughout all the region round about.
LUKE|7|18|And the disciples of John shewed him of all these things.
LUKE|7|19|And John calling unto him two of his disciples sent them to Jesus, saying, Art thou he that should come? or look we for another?
LUKE|7|20|When the men were come unto him, they said, John Baptist hath sent us unto thee, saying, Art thou he that should come? or look we for another?
LUKE|7|21|And in that same hour he cured many of their infirmities and plagues, and of evil spirits; and unto many that were blind he gave sight.
LUKE|7|22|Then Jesus answering said unto them, Go your way, and tell John what things ye have seen and heard; how that the blind see, the lame walk, the lepers are cleansed, the deaf hear, the dead are raised, to the poor the gospel is preached.
LUKE|7|23|And blessed is he, whosoever shall not be offended in me.
LUKE|7|24|And when the messengers of John were departed, he began to speak unto the people concerning John, What went ye out into the wilderness for to see? A reed shaken with the wind?
LUKE|7|25|But what went ye out for to see? A man clothed in soft raiment? Behold, they which are gorgeously apparelled, and live delicately, are in kings' courts.
LUKE|7|26|But what went ye out for to see? A prophet? Yea, I say unto you, and much more than a prophet.
LUKE|7|27|This is he, of whom it is written, Behold, I send my messenger before thy face, which shall prepare thy way before thee.
LUKE|7|28|For I say unto you, Among those that are born of women there is not a greater prophet than John the Baptist: but he that is least in the kingdom of God is greater than he.
LUKE|7|29|And all the people that heard him, and the publicans, justified God, being baptized with the baptism of John.
LUKE|7|30|But the Pharisees and lawyers rejected the counsel of God against themselves, being not baptized of him.
LUKE|7|31|And the Lord said, Whereunto then shall I liken the men of this generation? and to what are they like?
LUKE|7|32|They are like unto children sitting in the marketplace, and calling one to another, and saying, We have piped unto you, and ye have not danced; we have mourned to you, and ye have not wept.
LUKE|7|33|For John the Baptist came neither eating bread nor drinking wine; and ye say, He hath a devil.
LUKE|7|34|The Son of man is come eating and drinking; and ye say, Behold a gluttonous man, and a winebibber, a friend of publicans and sinners!
LUKE|7|35|But wisdom is justified of all her children.
LUKE|7|36|And one of the Pharisees desired him that he would eat with him. And he went into the Pharisee's house, and sat down to meat.
LUKE|7|37|And, behold, a woman in the city, which was a sinner, when she knew that Jesus sat at meat in the Pharisee's house, brought an alabaster box of ointment,
LUKE|7|38|And stood at his feet behind him weeping, and began to wash his feet with tears, and did wipe them with the hairs of her head, and kissed his feet, and anointed them with the ointment.
LUKE|7|39|Now when the Pharisee which had bidden him saw it, he spake within himself, saying, This man, if he were a prophet, would have known who and what manner of woman this is that toucheth him: for she is a sinner.
LUKE|7|40|And Jesus answering said unto him, Simon, I have somewhat to say unto thee. And he saith, Master, say on.
LUKE|7|41|There was a certain creditor which had two debtors: the one owed five hundred pence, and the other fifty.
LUKE|7|42|And when they had nothing to pay, he frankly forgave them both. Tell me therefore, which of them will love him most?
LUKE|7|43|Simon answered and said, I suppose that he, to whom he forgave most. And he said unto him, Thou hast rightly judged.
LUKE|7|44|And he turned to the woman, and said unto Simon, Seest thou this woman? I entered into thine house, thou gavest me no water for my feet: but she hath washed my feet with tears, and wiped them with the hairs of her head.
LUKE|7|45|Thou gavest me no kiss: but this woman since the time I came in hath not ceased to kiss my feet.
LUKE|7|46|My head with oil thou didst not anoint: but this woman hath anointed my feet with ointment.
LUKE|7|47|Wherefore I say unto thee, Her sins, which are many, are forgiven; for she loved much: but to whom little is forgiven, the same loveth little.
LUKE|7|48|And he said unto her, Thy sins are forgiven.
LUKE|7|49|And they that sat at meat with him began to say within themselves, Who is this that forgiveth sins also?
LUKE|7|50|And he said to the woman, Thy faith hath saved thee; go in peace.
LUKE|8|1|And it came to pass afterward, that he went throughout every city and village, preaching and shewing the glad tidings of the kingdom of God: and the twelve were with him,
LUKE|8|2|And certain women, which had been healed of evil spirits and infirmities, Mary called Magdalene, out of whom went seven devils,
LUKE|8|3|And Joanna the wife of Chuza Herod's steward, and Susanna, and many others, which ministered unto him of their substance.
LUKE|8|4|And when much people were gathered together, and were come to him out of every city, he spake by a parable:
LUKE|8|5|A sower went out to sow his seed: and as he sowed, some fell by the way side; and it was trodden down, and the fowls of the air devoured it.
LUKE|8|6|And some fell upon a rock; and as soon as it was sprung up, it withered away, because it lacked moisture.
LUKE|8|7|And some fell among thorns; and the thorns sprang up with it, and choked it.
LUKE|8|8|And other fell on good ground, and sprang up, and bare fruit an hundredfold. And when he had said these things, he cried, He that hath ears to hear, let him hear.
LUKE|8|9|And his disciples asked him, saying, What might this parable be?
LUKE|8|10|And he said, Unto you it is given to know the mysteries of the kingdom of God: but to others in parables; that seeing they might not see, and hearing they might not understand.
LUKE|8|11|Now the parable is this: The seed is the word of God.
LUKE|8|12|Those by the way side are they that hear; then cometh the devil, and taketh away the word out of their hearts, lest they should believe and be saved.
LUKE|8|13|They on the rock are they, which, when they hear, receive the word with joy; and these have no root, which for a while believe, and in time of temptation fall away.
LUKE|8|14|And that which fell among thorns are they, which, when they have heard, go forth, and are choked with cares and riches and pleasures of this life, and bring no fruit to perfection.
LUKE|8|15|But that on the good ground are they, which in an honest and good heart, having heard the word, keep it, and bring forth fruit with patience.
LUKE|8|16|No man, when he hath lighted a candle, covereth it with a vessel, or putteth it under a bed; but setteth it on a candlestick, that they which enter in may see the light.
LUKE|8|17|For nothing is secret, that shall not be made manifest; neither any thing hid, that shall not be known and come abroad.
LUKE|8|18|Take heed therefore how ye hear: for whosoever hath, to him shall be given; and whosoever hath not, from him shall be taken even that which he seemeth to have.
LUKE|8|19|Then came to him his mother and his brethren, and could not come at him for the press.
LUKE|8|20|And it was told him by certain which said, Thy mother and thy brethren stand without, desiring to see thee.
LUKE|8|21|And he answered and said unto them, My mother and my brethren are these which hear the word of God, and do it.
LUKE|8|22|Now it came to pass on a certain day, that he went into a ship with his disciples: and he said unto them, Let us go over unto the other side of the lake. And they launched forth.
LUKE|8|23|But as they sailed he fell asleep: and there came down a storm of wind on the lake; and they were filled with water, and were in jeopardy.
LUKE|8|24|And they came to him, and awoke him, saying, Master, master, we perish. Then he arose, and rebuked the wind and the raging of the water: and they ceased, and there was a calm.
LUKE|8|25|And he said unto them, Where is your faith? And they being afraid wondered, saying one to another, What manner of man is this! for he commandeth even the winds and water, and they obey him.
LUKE|8|26|And they arrived at the country of the Gadarenes, which is over against Galilee.
LUKE|8|27|And when he went forth to land, there met him out of the city a certain man, which had devils long time, and ware no clothes, neither abode in any house, but in the tombs.
LUKE|8|28|When he saw Jesus, he cried out, and fell down before him, and with a loud voice said, What have I to do with thee, Jesus, thou Son of God most high? I beseech thee, torment me not.
LUKE|8|29|(For he had commanded the unclean spirit to come out of the man. For oftentimes it had caught him: and he was kept bound with chains and in fetters; and he brake the bands, and was driven of the devil into the wilderness.)
LUKE|8|30|And Jesus asked him, saying, What is thy name? And he said, Legion: because many devils were entered into him.
LUKE|8|31|And they besought him that he would not command them to go out into the deep.
LUKE|8|32|And there was there an herd of many swine feeding on the mountain: and they besought him that he would suffer them to enter into them. And he suffered them.
LUKE|8|33|Then went the devils out of the man, and entered into the swine: and the herd ran violently down a steep place into the lake, and were choked.
LUKE|8|34|When they that fed them saw what was done, they fled, and went and told it in the city and in the country.
LUKE|8|35|Then they went out to see what was done; and came to Jesus, and found the man, out of whom the devils were departed, sitting at the feet of Jesus, clothed, and in his right mind: and they were afraid.
LUKE|8|36|They also which saw it told them by what means he that was possessed of the devils was healed.
LUKE|8|37|Then the whole multitude of the country of the Gadarenes round about besought him to depart from them; for they were taken with great fear: and he went up into the ship, and returned back again.
LUKE|8|38|Now the man out of whom the devils were departed besought him that he might be with him: but Jesus sent him away, saying,
LUKE|8|39|Return to thine own house, and shew how great things God hath done unto thee. And he went his way, and published throughout the whole city how great things Jesus had done unto him.
LUKE|8|40|And it came to pass, that, when Jesus was returned, the people gladly received him: for they were all waiting for him.
LUKE|8|41|And, behold, there came a man named Jairus, and he was a ruler of the synagogue: and he fell down at Jesus' feet, and besought him that he would come into his house:
LUKE|8|42|For he had one only daughter, about twelve years of age, and she lay a dying. But as he went the people thronged him.
LUKE|8|43|And a woman having an issue of blood twelve years, which had spent all her living upon physicians, neither could be healed of any,
LUKE|8|44|Came behind him, and touched the border of his garment: and immediately her issue of blood stanched.
LUKE|8|45|And Jesus said, Who touched me? When all denied, Peter and they that were with him said, Master, the multitude throng thee and press thee, and sayest thou, Who touched me?
LUKE|8|46|And Jesus said, Somebody hath touched me: for I perceive that virtue is gone out of me.
LUKE|8|47|And when the woman saw that she was not hid, she came trembling, and falling down before him, she declared unto him before all the people for what cause she had touched him, and how she was healed immediately.
LUKE|8|48|And he said unto her, Daughter, be of good comfort: thy faith hath made thee whole; go in peace.
LUKE|8|49|While he yet spake, there cometh one from the ruler of the synagogue's house, saying to him, Thy daughter is dead; trouble not the Master.
LUKE|8|50|But when Jesus heard it, he answered him, saying, Fear not: believe only, and she shall be made whole.
LUKE|8|51|And when he came into the house, he suffered no man to go in, save Peter, and James, and John, and the father and the mother of the maiden.
LUKE|8|52|And all wept, and bewailed her: but he said, Weep not; she is not dead, but sleepeth.
LUKE|8|53|And they laughed him to scorn, knowing that she was dead.
LUKE|8|54|And he put them all out, and took her by the hand, and called, saying, Maid, arise.
LUKE|8|55|And her spirit came again, and she arose straightway: and he commanded to give her meat.
LUKE|8|56|And her parents were astonished: but he charged them that they should tell no man what was done.
LUKE|9|1|Then he called his twelve disciples together, and gave them power and authority over all devils, and to cure diseases.
LUKE|9|2|And he sent them to preach the kingdom of God, and to heal the sick.
LUKE|9|3|And he said unto them, Take nothing for your journey, neither staves, nor scrip, neither bread, neither money; neither have two coats apiece.
LUKE|9|4|And whatsoever house ye enter into, there abide, and thence depart.
LUKE|9|5|And whosoever will not receive you, when ye go out of that city, shake off the very dust from your feet for a testimony against them.
LUKE|9|6|And they departed, and went through the towns, preaching the gospel, and healing every where.
LUKE|9|7|Now Herod the tetrarch heard of all that was done by him: and he was perplexed, because that it was said of some, that John was risen from the dead;
LUKE|9|8|And of some, that Elias had appeared; and of others, that one of the old prophets was risen again.
LUKE|9|9|And Herod said, John have I beheaded: but who is this, of whom I hear such things? And he desired to see him.
LUKE|9|10|And the apostles, when they were returned, told him all that they had done. And he took them, and went aside privately into a desert place belonging to the city called Bethsaida.
LUKE|9|11|And the people, when they knew it, followed him: and he received them, and spake unto them of the kingdom of God, and healed them that had need of healing.
LUKE|9|12|And when the day began to wear away, then came the twelve, and said unto him, Send the multitude away, that they may go into the towns and country round about, and lodge, and get victuals: for we are here in a desert place.
LUKE|9|13|But he said unto them, Give ye them to eat. And they said, We have no more but five loaves and two fishes; except we should go and buy meat for all this people.
LUKE|9|14|For they were about five thousand men. And he said to his disciples, Make them sit down by fifties in a company.
LUKE|9|15|And they did so, and made them all sit down.
LUKE|9|16|Then he took the five loaves and the two fishes, and looking up to heaven, he blessed them, and brake, and gave to the disciples to set before the multitude.
LUKE|9|17|And they did eat, and were all filled: and there was taken up of fragments that remained to them twelve baskets.
LUKE|9|18|And it came to pass, as he was alone praying, his disciples were with him: and he asked them, saying, Whom say the people that I am?
LUKE|9|19|They answering said, John the Baptist; but some say, Elias; and others say, that one of the old prophets is risen again.
LUKE|9|20|He said unto them, But whom say ye that I am? Peter answering said, The Christ of God.
LUKE|9|21|And he straitly charged them, and commanded them to tell no man that thing;
LUKE|9|22|Saying, The Son of man must suffer many things, and be rejected of the elders and chief priests and scribes, and be slain, and be raised the third day.
LUKE|9|23|And he said to them all, If any man will come after me, let him deny himself, and take up his cross daily, and follow me.
LUKE|9|24|For whosoever will save his life shall lose it: but whosoever will lose his life for my sake, the same shall save it.
LUKE|9|25|For what is a man advantaged, if he gain the whole world, and lose himself, or be cast away?
LUKE|9|26|For whosoever shall be ashamed of me and of my words, of him shall the Son of man be ashamed, when he shall come in his own glory, and in his Father's, and of the holy angels.
LUKE|9|27|But I tell you of a truth, there be some standing here, which shall not taste of death, till they see the kingdom of God.
LUKE|9|28|And it came to pass about an eight days after these sayings, he took Peter and John and James, and went up into a mountain to pray.
LUKE|9|29|And as he prayed, the fashion of his countenance was altered, and his raiment was white and glistering.
LUKE|9|30|And, behold, there talked with him two men, which were Moses and Elias:
LUKE|9|31|Who appeared in glory, and spake of his decease which he should accomplish at Jerusalem.
LUKE|9|32|But Peter and they that were with him were heavy with sleep: and when they were awake, they saw his glory, and the two men that stood with him.
LUKE|9|33|And it came to pass, as they departed from him, Peter said unto Jesus, Master, it is good for us to be here: and let us make three tabernacles; one for thee, and one for Moses, and one for Elias: not knowing what he said.
LUKE|9|34|While he thus spake, there came a cloud, and overshadowed them: and they feared as they entered into the cloud.
LUKE|9|35|And there came a voice out of the cloud, saying, This is my beloved Son: hear him.
LUKE|9|36|And when the voice was past, Jesus was found alone. And they kept it close, and told no man in those days any of those things which they had seen.
LUKE|9|37|And it came to pass, that on the next day, when they were come down from the hill, much people met him.
LUKE|9|38|And, behold, a man of the company cried out, saying, Master, I beseech thee, look upon my son: for he is mine only child.
LUKE|9|39|And, lo, a spirit taketh him, and he suddenly crieth out; and it teareth him that he foameth again, and bruising him hardly departeth from him.
LUKE|9|40|And I besought thy disciples to cast him out; and they could not.
LUKE|9|41|And Jesus answering said, O faithless and perverse generation, how long shall I be with you, and suffer you? Bring thy son hither.
LUKE|9|42|And as he was yet a coming, the devil threw him down, and tare him. And Jesus rebuked the unclean spirit, and healed the child, and delivered him again to his father.
LUKE|9|43|And they were all amazed at the mighty power of God. But while they wondered every one at all things which Jesus did, he said unto his disciples,
LUKE|9|44|Let these sayings sink down into your ears: for the Son of man shall be delivered into the hands of men.
LUKE|9|45|But they understood not this saying, and it was hid from them, that they perceived it not: and they feared to ask him of that saying.
LUKE|9|46|Then there arose a reasoning among them, which of them should be greatest.
LUKE|9|47|And Jesus, perceiving the thought of their heart, took a child, and set him by him,
LUKE|9|48|And said unto them, Whosoever shall receive this child in my name receiveth me: and whosoever shall receive me receiveth him that sent me: for he that is least among you all, the same shall be great.
LUKE|9|49|And John answered and said, Master, we saw one casting out devils in thy name; and we forbad him, because he followeth not with us.
LUKE|9|50|And Jesus said unto him, Forbid him not: for he that is not against us is for us.
LUKE|9|51|And it came to pass, when the time was come that he should be received up, he stedfastly set his face to go to Jerusalem,
LUKE|9|52|And sent messengers before his face: and they went, and entered into a village of the Samaritans, to make ready for him.
LUKE|9|53|And they did not receive him, because his face was as though he would go to Jerusalem.
LUKE|9|54|And when his disciples James and John saw this, they said, Lord, wilt thou that we command fire to come down from heaven, and consume them, even as Elias did?
LUKE|9|55|But he turned, and rebuked them, and said, Ye know not what manner of spirit ye are of.
LUKE|9|56|For the Son of man is not come to destroy men's lives, but to save them. And they went to another village.
LUKE|9|57|And it came to pass, that, as they went in the way, a certain man said unto him, Lord, I will follow thee whithersoever thou goest.
LUKE|9|58|And Jesus said unto him, Foxes have holes, and birds of the air have nests; but the Son of man hath not where to lay his head.
LUKE|9|59|And he said unto another, Follow me. But he said, Lord, suffer me first to go and bury my father.
LUKE|9|60|Jesus said unto him, Let the dead bury their dead: but go thou and preach the kingdom of God.
LUKE|9|61|And another also said, Lord, I will follow thee; but let me first go bid them farewell, which are at home at my house.
LUKE|9|62|And Jesus said unto him, No man, having put his hand to the plough, and looking back, is fit for the kingdom of God.
LUKE|10|1|After these things the LORD appointed other seventy also, and sent them two and two before his face into every city and place, whither he himself would come.
LUKE|10|2|Therefore said he unto them, The harvest truly is great, but the labourers are few: pray ye therefore the Lord of the harvest, that he would send forth labourers into his harvest.
LUKE|10|3|Go your ways: behold, I send you forth as lambs among wolves.
LUKE|10|4|Carry neither purse, nor scrip, nor shoes: and salute no man by the way.
LUKE|10|5|And into whatsoever house ye enter, first say, Peace be to this house.
LUKE|10|6|And if the son of peace be there, your peace shall rest upon it: if not, it shall turn to you again.
LUKE|10|7|And in the same house remain, eating and drinking such things as they give: for the labourer is worthy of his hire. Go not from house to house.
LUKE|10|8|And into whatsoever city ye enter, and they receive you, eat such things as are set before you:
LUKE|10|9|And heal the sick that are therein, and say unto them, The kingdom of God is come nigh unto you.
LUKE|10|10|But into whatsoever city ye enter, and they receive you not, go your ways out into the streets of the same, and say,
LUKE|10|11|Even the very dust of your city, which cleaveth on us, we do wipe off against you: notwithstanding be ye sure of this, that the kingdom of God is come nigh unto you.
LUKE|10|12|But I say unto you, that it shall be more tolerable in that day for Sodom, than for that city.
LUKE|10|13|Woe unto thee, Chorazin! woe unto thee, Bethsaida! for if the mighty works had been done in Tyre and Sidon, which have been done in you, they had a great while ago repented, sitting in sackcloth and ashes.
LUKE|10|14|But it shall be more tolerable for Tyre and Sidon at the judgment, than for you.
LUKE|10|15|And thou, Capernaum, which art exalted to heaven, shalt be thrust down to hell.
LUKE|10|16|He that heareth you heareth me; and he that despiseth you despiseth me; and he that despiseth me despiseth him that sent me.
LUKE|10|17|And the seventy returned again with joy, saying, Lord, even the devils are subject unto us through thy name.
LUKE|10|18|And he said unto them, I beheld Satan as lightning fall from heaven.
LUKE|10|19|Behold, I give unto you power to tread on serpents and scorpions, and over all the power of the enemy: and nothing shall by any means hurt you.
LUKE|10|20|Notwithstanding in this rejoice not, that the spirits are subject unto you; but rather rejoice, because your names are written in heaven.
LUKE|10|21|In that hour Jesus rejoiced in spirit, and said, I thank thee, O Father, Lord of heaven and earth, that thou hast hid these things from the wise and prudent, and hast revealed them unto babes: even so, Father; for so it seemed good in thy sight.
LUKE|10|22|All things are delivered to me of my Father: and no man knoweth who the Son is, but the Father; and who the Father is, but the Son, and he to whom the Son will reveal him.
LUKE|10|23|And he turned him unto his disciples, and said privately, Blessed are the eyes which see the things that ye see:
LUKE|10|24|For I tell you, that many prophets and kings have desired to see those things which ye see, and have not seen them; and to hear those things which ye hear, and have not heard them.
LUKE|10|25|And, behold, a certain lawyer stood up, and tempted him, saying, Master, what shall I do to inherit eternal life?
LUKE|10|26|He said unto him, What is written in the law? how readest thou?
LUKE|10|27|And he answering said, Thou shalt love the Lord thy God with all thy heart, and with all thy soul, and with all thy strength, and with all thy mind; and thy neighbour as thyself.
LUKE|10|28|And he said unto him, Thou hast answered right: this do, and thou shalt live.
LUKE|10|29|But he, willing to justify himself, said unto Jesus, And who is my neighbour?
LUKE|10|30|And Jesus answering said, A certain man went down from Jerusalem to Jericho, and fell among thieves, which stripped him of his raiment, and wounded him, and departed, leaving him half dead.
LUKE|10|31|And by chance there came down a certain priest that way: and when he saw him, he passed by on the other side.
LUKE|10|32|And likewise a Levite, when he was at the place, came and looked on him, and passed by on the other side.
LUKE|10|33|But a certain Samaritan, as he journeyed, came where he was: and when he saw him, he had compassion on him,
LUKE|10|34|And went to him, and bound up his wounds, pouring in oil and wine, and set him on his own beast, and brought him to an inn, and took care of him.
LUKE|10|35|And on the morrow when he departed, he took out two pence, and gave them to the host, and said unto him, Take care of him; and whatsoever thou spendest more, when I come again, I will repay thee.
LUKE|10|36|Which now of these three, thinkest thou, was neighbour unto him that fell among the thieves?
LUKE|10|37|And he said, He that shewed mercy on him. Then said Jesus unto him, Go, and do thou likewise.
LUKE|10|38|Now it came to pass, as they went, that he entered into a certain village: and a certain woman named Martha received him into her house.
LUKE|10|39|And she had a sister called Mary, which also sat at Jesus' feet, and heard his word.
LUKE|10|40|But Martha was cumbered about much serving, and came to him, and said, Lord, dost thou not care that my sister hath left me to serve alone? bid her therefore that she help me.
LUKE|10|41|And Jesus answered and said unto her, Martha, Martha, thou art careful and troubled about many things:
LUKE|10|42|But one thing is needful: and Mary hath chosen that good part, which shall not be taken away from her.
LUKE|11|1|And it came to pass, that, as he was praying in a certain place, when he ceased, one of his disciples said unto him, Lord, teach us to pray, as John also taught his disciples.
LUKE|11|2|And he said unto them, When ye pray, say, Our Father which art in heaven, Hallowed be thy name. Thy kingdom come. Thy will be done, as in heaven, so in earth.
LUKE|11|3|Give us day by day our daily bread.
LUKE|11|4|And forgive us our sins; for we also forgive every one that is indebted to us. And lead us not into temptation; but deliver us from evil.
LUKE|11|5|And he said unto them, Which of you shall have a friend, and shall go unto him at midnight, and say unto him, Friend, lend me three loaves;
LUKE|11|6|For a friend of mine in his journey is come to me, and I have nothing to set before him?
LUKE|11|7|And he from within shall answer and say, Trouble me not: the door is now shut, and my children are with me in bed; I cannot rise and give thee.
LUKE|11|8|I say unto you, Though he will not rise and give him, because he is his friend, yet because of his importunity he will rise and give him as many as he needeth.
LUKE|11|9|And I say unto you, Ask, and it shall be given you; seek, and ye shall find; knock, and it shall be opened unto you.
LUKE|11|10|For every one that asketh receiveth; and he that seeketh findeth; and to him that knocketh it shall be opened.
LUKE|11|11|If a son shall ask bread of any of you that is a father, will he give him a stone? or if he ask a fish, will he for a fish give him a serpent?
LUKE|11|12|Or if he shall ask an egg, will he offer him a scorpion?
LUKE|11|13|If ye then, being evil, know how to give good gifts unto your children: how much more shall your heavenly Father give the Holy Spirit to them that ask him?
LUKE|11|14|And he was casting out a devil, and it was dumb. And it came to pass, when the devil was gone out, the dumb spake; and the people wondered.
LUKE|11|15|But some of them said, He casteth out devils through Beelzebub the chief of the devils.
LUKE|11|16|And others, tempting him, sought of him a sign from heaven.
LUKE|11|17|But he, knowing their thoughts, said unto them, Every kingdom divided against itself is brought to desolation; and a house divided against a house falleth.
LUKE|11|18|If Satan also be divided against himself, how shall his kingdom stand? because ye say that I cast out devils through Beelzebub.
LUKE|11|19|And if I by Beelzebub cast out devils, by whom do your sons cast them out? therefore shall they be your judges.
LUKE|11|20|But if I with the finger of God cast out devils, no doubt the kingdom of God is come upon you.
LUKE|11|21|When a strong man armed keepeth his palace, his goods are in peace:
LUKE|11|22|But when a stronger than he shall come upon him, and overcome him, he taketh from him all his armour wherein he trusted, and divideth his spoils.
LUKE|11|23|He that is not with me is against me: and he that gathereth not with me scattereth.
LUKE|11|24|When the unclean spirit is gone out of a man, he walketh through dry places, seeking rest; and finding none, he saith, I will return unto my house whence I came out.
LUKE|11|25|And when he cometh, he findeth it swept and garnished.
LUKE|11|26|Then goeth he, and taketh to him seven other spirits more wicked than himself; and they enter in, and dwell there: and the last state of that man is worse than the first.
LUKE|11|27|And it came to pass, as he spake these things, a certain woman of the company lifted up her voice, and said unto him, Blessed is the womb that bare thee, and the paps which thou hast sucked.
LUKE|11|28|But he said, Yea rather, blessed are they that hear the word of God, and keep it.
LUKE|11|29|And when the people were gathered thick together, he began to say, This is an evil generation: they seek a sign; and there shall no sign be given it, but the sign of Jonas the prophet.
LUKE|11|30|For as Jonas was a sign unto the Ninevites, so shall also the Son of man be to this generation.
LUKE|11|31|The queen of the south shall rise up in the judgment with the men of this generation, and condemn them: for she came from the utmost parts of the earth to hear the wisdom of Solomon; and, behold, a greater than Solomon is here.
LUKE|11|32|The men of Nineve shall rise up in the judgment with this generation, and shall condemn it: for they repented at the preaching of Jonas; and, behold, a greater than Jonas is here.
LUKE|11|33|No man, when he hath lighted a candle, putteth it in a secret place, neither under a bushel, but on a candlestick, that they which come in may see the light.
LUKE|11|34|The light of the body is the eye: therefore when thine eye is single, thy whole body also is full of light; but when thine eye is evil, thy body also is full of darkness.
LUKE|11|35|Take heed therefore that the light which is in thee be not darkness.
LUKE|11|36|If thy whole body therefore be full of light, having no part dark, the whole shall be full of light, as when the bright shining of a candle doth give thee light.
LUKE|11|37|And as he spake, a certain Pharisee besought him to dine with him: and he went in, and sat down to meat.
LUKE|11|38|And when the Pharisee saw it, he marvelled that he had not first washed before dinner.
LUKE|11|39|And the Lord said unto him, Now do ye Pharisees make clean the outside of the cup and the platter; but your inward part is full of ravening and wickedness.
LUKE|11|40|Ye fools, did not he that made that which is without make that which is within also?
LUKE|11|41|But rather give alms of such things as ye have; and, behold, all things are clean unto you.
LUKE|11|42|But woe unto you, Pharisees! for ye tithe mint and rue and all manner of herbs, and pass over judgment and the love of God: these ought ye to have done, and not to leave the other undone.
LUKE|11|43|Woe unto you, Pharisees! for ye love the uppermost seats in the synagogues, and greetings in the markets.
LUKE|11|44|Woe unto you, scribes and Pharisees, hypocrites! for ye are as graves which appear not, and the men that walk over them are not aware of them.
LUKE|11|45|Then answered one of the lawyers, and said unto him, Master, thus saying thou reproachest us also.
LUKE|11|46|And he said, Woe unto you also, ye lawyers! for ye lade men with burdens grievous to be borne, and ye yourselves touch not the burdens with one of your fingers.
LUKE|11|47|Woe unto you! for ye build the sepulchres of the prophets, and your fathers killed them.
LUKE|11|48|Truly ye bear witness that ye allow the deeds of your fathers: for they indeed killed them, and ye build their sepulchres.
LUKE|11|49|Therefore also said the wisdom of God, I will send them prophets and apostles, and some of them they shall slay and persecute:
LUKE|11|50|That the blood of all the prophets, which was shed from the foundation of the world, may be required of this generation;
LUKE|11|51|From the blood of Abel unto the blood of Zacharias which perished between the altar and the temple: verily I say unto you, It shall be required of this generation.
LUKE|11|52|Woe unto you, lawyers! for ye have taken away the key of knowledge: ye entered not in yourselves, and them that were entering in ye hindered.
LUKE|11|53|And as he said these things unto them, the scribes and the Pharisees began to urge him vehemently, and to provoke him to speak of many things:
LUKE|11|54|Laying wait for him, and seeking to catch something out of his mouth, that they might accuse him.
LUKE|12|1|In the mean time, when there were gathered together an innumerable multitude of people, insomuch that they trode one upon another, he began to say unto his disciples first of all, Beware ye of the leaven of the Pharisees, which is hypocrisy.
LUKE|12|2|For there is nothing covered, that shall not be revealed; neither hid, that shall not be known.
LUKE|12|3|Therefore whatsoever ye have spoken in darkness shall be heard in the light; and that which ye have spoken in the ear in closets shall be proclaimed upon the housetops.
LUKE|12|4|And I say unto you my friends, Be not afraid of them that kill the body, and after that have no more that they can do.
LUKE|12|5|But I will forewarn you whom ye shall fear: Fear him, which after he hath killed hath power to cast into hell; yea, I say unto you, Fear him.
LUKE|12|6|Are not five sparrows sold for two farthings, and not one of them is forgotten before God?
LUKE|12|7|But even the very hairs of your head are all numbered. Fear not therefore: ye are of more value than many sparrows.
LUKE|12|8|Also I say unto you, Whosoever shall confess me before men, him shall the Son of man also confess before the angels of God:
LUKE|12|9|But he that denieth me before men shall be denied before the angels of God.
LUKE|12|10|And whosoever shall speak a word against the Son of man, it shall be forgiven him: but unto him that blasphemeth against the Holy Ghost it shall not be forgiven.
LUKE|12|11|And when they bring you unto the synagogues, and unto magistrates, and powers, take ye no thought how or what thing ye shall answer, or what ye shall say:
LUKE|12|12|For the Holy Ghost shall teach you in the same hour what ye ought to say.
LUKE|12|13|And one of the company said unto him, Master, speak to my brother, that he divide the inheritance with me.
LUKE|12|14|And he said unto him, Man, who made me a judge or a divider over you?
LUKE|12|15|And he said unto them, Take heed, and beware of covetousness: for a man's life consisteth not in the abundance of the things which he possesseth.
LUKE|12|16|And he spake a parable unto them, saying, The ground of a certain rich man brought forth plentifully:
LUKE|12|17|And he thought within himself, saying, What shall I do, because I have no room where to bestow my fruits?
LUKE|12|18|And he said, This will I do: I will pull down my barns, and build greater; and there will I bestow all my fruits and my goods.
LUKE|12|19|And I will say to my soul, Soul, thou hast much goods laid up for many years; take thine ease, eat, drink, and be merry.
LUKE|12|20|But God said unto him, Thou fool, this night thy soul shall be required of thee: then whose shall those things be, which thou hast provided?
LUKE|12|21|So is he that layeth up treasure for himself, and is not rich toward God.
LUKE|12|22|And he said unto his disciples, Therefore I say unto you, Take no thought for your life, what ye shall eat; neither for the body, what ye shall put on.
LUKE|12|23|The life is more than meat, and the body is more than raiment.
LUKE|12|24|Consider the ravens: for they neither sow nor reap; which neither have storehouse nor barn; and God feedeth them: how much more are ye better than the fowls?
LUKE|12|25|And which of you with taking thought can add to his stature one cubit?
LUKE|12|26|If ye then be not able to do that thing which is least, why take ye thought for the rest?
LUKE|12|27|Consider the lilies how they grow: they toil not, they spin not; and yet I say unto you, that Solomon in all his glory was not arrayed like one of these.
LUKE|12|28|If then God so clothe the grass, which is to day in the field, and to morrow is cast into the oven; how much more will he clothe you, O ye of little faith?
LUKE|12|29|And seek not ye what ye shall eat, or what ye shall drink, neither be ye of doubtful mind.
LUKE|12|30|For all these things do the nations of the world seek after: and your Father knoweth that ye have need of these things.
LUKE|12|31|But rather seek ye the kingdom of God; and all these things shall be added unto you.
LUKE|12|32|Fear not, little flock; for it is your Father's good pleasure to give you the kingdom.
LUKE|12|33|Sell that ye have, and give alms; provide yourselves bags which wax not old, a treasure in the heavens that faileth not, where no thief approacheth, neither moth corrupteth.
LUKE|12|34|For where your treasure is, there will your heart be also.
LUKE|12|35|Let your loins be girded about, and your lights burning;
LUKE|12|36|And ye yourselves like unto men that wait for their lord, when he will return from the wedding; that when he cometh and knocketh, they may open unto him immediately.
LUKE|12|37|Blessed are those servants, whom the lord when he cometh shall find watching: verily I say unto you, that he shall gird himself, and make them to sit down to meat, and will come forth and serve them.
LUKE|12|38|And if he shall come in the second watch, or come in the third watch, and find them so, blessed are those servants.
LUKE|12|39|And this know, that if the goodman of the house had known what hour the thief would come, he would have watched, and not have suffered his house to be broken through.
LUKE|12|40|Be ye therefore ready also: for the Son of man cometh at an hour when ye think not.
LUKE|12|41|Then Peter said unto him, Lord, speakest thou this parable unto us, or even to all?
LUKE|12|42|And the Lord said, Who then is that faithful and wise steward, whom his lord shall make ruler over his household, to give them their portion of meat in due season?
LUKE|12|43|Blessed is that servant, whom his lord when he cometh shall find so doing.
LUKE|12|44|Of a truth I say unto you, that he will make him ruler over all that he hath.
LUKE|12|45|But and if that servant say in his heart, My lord delayeth his coming; and shall begin to beat the menservants and maidens, and to eat and drink, and to be drunken;
LUKE|12|46|The lord of that servant will come in a day when he looketh not for him, and at an hour when he is not aware, and will cut him in sunder, and will appoint him his portion with the unbelievers.
LUKE|12|47|And that servant, which knew his lord's will, and prepared not himself, neither did according to his will, shall be beaten with many stripes.
LUKE|12|48|But he that knew not, and did commit things worthy of stripes, shall be beaten with few stripes. For unto whomsoever much is given, of him shall be much required: and to whom men have committed much, of him they will ask the more.
LUKE|12|49|I am come to send fire on the earth; and what will I, if it be already kindled?
LUKE|12|50|But I have a baptism to be baptized with; and how am I straitened till it be accomplished!
LUKE|12|51|Suppose ye that I am come to give peace on earth? I tell you, Nay; but rather division:
LUKE|12|52|For from henceforth there shall be five in one house divided, three against two, and two against three.
LUKE|12|53|The father shall be divided against the son, and the son against the father; the mother against the daughter, and the daughter against the mother; the mother in law against her daughter in law, and the daughter in law against her mother in law.
LUKE|12|54|And he said also to the people, When ye see a cloud rise out of the west, straightway ye say, There cometh a shower; and so it is.
LUKE|12|55|And when ye see the south wind blow, ye say, There will be heat; and it cometh to pass.
LUKE|12|56|Ye hypocrites, ye can discern the face of the sky and of the earth; but how is it that ye do not discern this time?
LUKE|12|57|Yea, and why even of yourselves judge ye not what is right?
LUKE|12|58|When thou goest with thine adversary to the magistrate, as thou art in the way, give diligence that thou mayest be delivered from him; lest he hale thee to the judge, and the judge deliver thee to the officer, and the officer cast thee into prison.
LUKE|12|59|I tell thee, thou shalt not depart thence, till thou hast paid the very last mite.
LUKE|13|1|There were present at that season some that told him of the Galilaeans, whose blood Pilate had mingled with their sacrifices.
LUKE|13|2|And Jesus answering said unto them, Suppose ye that these Galilaeans were sinners above all the Galilaeans, because they suffered such things?
LUKE|13|3|I tell you, Nay: but, except ye repent, ye shall all likewise perish.
LUKE|13|4|Or those eighteen, upon whom the tower in Siloam fell, and slew them, think ye that they were sinners above all men that dwelt in Jerusalem?
LUKE|13|5|I tell you, Nay: but, except ye repent, ye shall all likewise perish.
LUKE|13|6|He spake also this parable; A certain man had a fig tree planted in his vineyard; and he came and sought fruit thereon, and found none.
LUKE|13|7|Then said he unto the dresser of his vineyard, Behold, these three years I come seeking fruit on this fig tree, and find none: cut it down; why cumbereth it the ground?
LUKE|13|8|And he answering said unto him, Lord, let it alone this year also, till I shall dig about it, and dung it:
LUKE|13|9|And if it bear fruit, well: and if not, then after that thou shalt cut it down.
LUKE|13|10|And he was teaching in one of the synagogues on the sabbath.
LUKE|13|11|And, behold, there was a woman which had a spirit of infirmity eighteen years, and was bowed together, and could in no wise lift up herself.
LUKE|13|12|And when Jesus saw her, he called her to him, and said unto her, Woman, thou art loosed from thine infirmity.
LUKE|13|13|And he laid his hands on her: and immediately she was made straight, and glorified God.
LUKE|13|14|And the ruler of the synagogue answered with indignation, because that Jesus had healed on the sabbath day, and said unto the people, There are six days in which men ought to work: in them therefore come and be healed, and not on the sabbath day.
LUKE|13|15|The Lord then answered him, and said, Thou hypocrite, doth not each one of you on the sabbath loose his ox or his ass from the stall, and lead him away to watering?
LUKE|13|16|And ought not this woman, being a daughter of Abraham, whom Satan hath bound, lo, these eighteen years, be loosed from this bond on the sabbath day?
LUKE|13|17|And when he had said these things, all his adversaries were ashamed: and all the people rejoiced for all the glorious things that were done by him.
LUKE|13|18|Then said he, Unto what is the kingdom of God like? and whereunto shall I resemble it?
LUKE|13|19|It is like a grain of mustard seed, which a man took, and cast into his garden; and it grew, and waxed a great tree; and the fowls of the air lodged in the branches of it.
LUKE|13|20|And again he said, Whereunto shall I liken the kingdom of God?
LUKE|13|21|It is like leaven, which a woman took and hid in three measures of meal, till the whole was leavened.
LUKE|13|22|And he went through the cities and villages, teaching, and journeying toward Jerusalem.
LUKE|13|23|Then said one unto him, Lord, are there few that be saved? And he said unto them,
LUKE|13|24|Strive to enter in at the strait gate: for many, I say unto you, will seek to enter in, and shall not be able.
LUKE|13|25|When once the master of the house is risen up, and hath shut to the door, and ye begin to stand without, and to knock at the door, saying, Lord, Lord, open unto us; and he shall answer and say unto you, I know you not whence ye are:
LUKE|13|26|Then shall ye begin to say, We have eaten and drunk in thy presence, and thou hast taught in our streets.
LUKE|13|27|But he shall say, I tell you, I know you not whence ye are; depart from me, all ye workers of iniquity.
LUKE|13|28|There shall be weeping and gnashing of teeth, when ye shall see Abraham, and Isaac, and Jacob, and all the prophets, in the kingdom of God, and you yourselves thrust out.
LUKE|13|29|And they shall come from the east, and from the west, and from the north, and from the south, and shall sit down in the kingdom of God.
LUKE|13|30|And, behold, there are last which shall be first, and there are first which shall be last.
LUKE|13|31|The same day there came certain of the Pharisees, saying unto him, Get thee out, and depart hence: for Herod will kill thee.
LUKE|13|32|And he said unto them, Go ye, and tell that fox, Behold, I cast out devils, and I do cures to day and to morrow, and the third day I shall be perfected.
LUKE|13|33|Nevertheless I must walk to day, and to morrow, and the day following: for it cannot be that a prophet perish out of Jerusalem.
LUKE|13|34|O Jerusalem, Jerusalem, which killest the prophets, and stonest them that are sent unto thee; how often would I have gathered thy children together, as a hen doth gather her brood under her wings, and ye would not!
LUKE|13|35|Behold, your house is left unto you desolate: and verily I say unto you, Ye shall not see me, until the time come when ye shall say, Blessed is he that cometh in the name of the Lord.
LUKE|14|1|And it came to pass, as he went into the house of one of the chief Pharisees to eat bread on the sabbath day, that they watched him.
LUKE|14|2|And, behold, there was a certain man before him which had the dropsy.
LUKE|14|3|And Jesus answering spake unto the lawyers and Pharisees, saying, Is it lawful to heal on the sabbath day?
LUKE|14|4|And they held their peace. And he took him, and healed him, and let him go;
LUKE|14|5|And answered them, saying, Which of you shall have an ass or an ox fallen into a pit, and will not straightway pull him out on the sabbath day?
LUKE|14|6|And they could not answer him again to these things.
LUKE|14|7|And he put forth a parable to those which were bidden, when he marked how they chose out the chief rooms; saying unto them.
LUKE|14|8|When thou art bidden of any man to a wedding, sit not down in the highest room; lest a more honourable man than thou be bidden of him;
LUKE|14|9|And he that bade thee and him come and say to thee, Give this man place; and thou begin with shame to take the lowest room.
LUKE|14|10|But when thou art bidden, go and sit down in the lowest room; that when he that bade thee cometh, he may say unto thee, Friend, go up higher: then shalt thou have worship in the presence of them that sit at meat with thee.
LUKE|14|11|For whosoever exalteth himself shall be abased; and he that humbleth himself shall be exalted.
LUKE|14|12|Then said he also to him that bade him, When thou makest a dinner or a supper, call not thy friends, nor thy brethren, neither thy kinsmen, nor thy rich neighbours; lest they also bid thee again, and a recompence be made thee.
LUKE|14|13|But when thou makest a feast, call the poor, the maimed, the lame, the blind:
LUKE|14|14|And thou shalt be blessed; for they cannot recompense thee: for thou shalt be recompensed at the resurrection of the just.
LUKE|14|15|And when one of them that sat at meat with him heard these things, he said unto him, Blessed is he that shall eat bread in the kingdom of God.
LUKE|14|16|Then said he unto him, A certain man made a great supper, and bade many:
LUKE|14|17|And sent his servant at supper time to say to them that were bidden, Come; for all things are now ready.
LUKE|14|18|And they all with one consent began to make excuse. The first said unto him, I have bought a piece of ground, and I must needs go and see it: I pray thee have me excused.
LUKE|14|19|And another said, I have bought five yoke of oxen, and I go to prove them: I pray thee have me excused.
LUKE|14|20|And another said, I have married a wife, and therefore I cannot come.
LUKE|14|21|So that servant came, and shewed his lord these things. Then the master of the house being angry said to his servant, Go out quickly into the streets and lanes of the city, and bring in hither the poor, and the maimed, and the halt, and the blind.
LUKE|14|22|And the servant said, Lord, it is done as thou hast commanded, and yet there is room.
LUKE|14|23|And the lord said unto the servant, Go out into the highways and hedges, and compel them to come in, that my house may be filled.
LUKE|14|24|For I say unto you, That none of those men which were bidden shall taste of my supper.
LUKE|14|25|And there went great multitudes with him: and he turned, and said unto them,
LUKE|14|26|If any man come to me, and hate not his father, and mother, and wife, and children, and brethren, and sisters, yea, and his own life also, he cannot be my disciple.
LUKE|14|27|And whosoever doth not bear his cross, and come after me, cannot be my disciple.
LUKE|14|28|For which of you, intending to build a tower, sitteth not down first, and counteth the cost, whether he have sufficient to finish it?
LUKE|14|29|Lest haply, after he hath laid the foundation, and is not able to finish it, all that behold it begin to mock him,
LUKE|14|30|Saying, This man began to build, and was not able to finish.
LUKE|14|31|Or what king, going to make war against another king, sitteth not down first, and consulteth whether he be able with ten thousand to meet him that cometh against him with twenty thousand?
LUKE|14|32|Or else, while the other is yet a great way off, he sendeth an ambassage, and desireth conditions of peace.
LUKE|14|33|So likewise, whosoever he be of you that forsaketh not all that he hath, he cannot be my disciple.
LUKE|14|34|Salt is good: but if the salt have lost his savour, wherewith shall it be seasoned?
LUKE|14|35|It is neither fit for the land, nor yet for the dunghill; but men cast it out. He that hath ears to hear, let him hear.
LUKE|15|1|Then drew near unto him all the publicans and sinners for to hear him.
LUKE|15|2|And the Pharisees and scribes murmured, saying, This man receiveth sinners, and eateth with them.
LUKE|15|3|And he spake this parable unto them, saying,
LUKE|15|4|What man of you, having an hundred sheep, if he lose one of them, doth not leave the ninety and nine in the wilderness, and go after that which is lost, until he find it?
LUKE|15|5|And when he hath found it, he layeth it on his shoulders, rejoicing.
LUKE|15|6|And when he cometh home, he calleth together his friends and neighbours, saying unto them, Rejoice with me; for I have found my sheep which was lost.
LUKE|15|7|I say unto you, that likewise joy shall be in heaven over one sinner that repenteth, more than over ninety and nine just persons, which need no repentance.
LUKE|15|8|Either what woman having ten pieces of silver, if she lose one piece, doth not light a candle, and sweep the house, and seek diligently till she find it?
LUKE|15|9|And when she hath found it, she calleth her friends and her neighbours together, saying, Rejoice with me; for I have found the piece which I had lost.
LUKE|15|10|Likewise, I say unto you, there is joy in the presence of the angels of God over one sinner that repenteth.
LUKE|15|11|And he said, A certain man had two sons:
LUKE|15|12|And the younger of them said to his father, Father, give me the portion of goods that falleth to me. And he divided unto them his living.
LUKE|15|13|And not many days after the younger son gathered all together, and took his journey into a far country, and there wasted his substance with riotous living.
LUKE|15|14|And when he had spent all, there arose a mighty famine in that land; and he began to be in want.
LUKE|15|15|And he went and joined himself to a citizen of that country; and he sent him into his fields to feed swine.
LUKE|15|16|And he would fain have filled his belly with the husks that the swine did eat: and no man gave unto him.
LUKE|15|17|And when he came to himself, he said, How many hired servants of my father's have bread enough and to spare, and I perish with hunger!
LUKE|15|18|I will arise and go to my father, and will say unto him, Father, I have sinned against heaven, and before thee,
LUKE|15|19|And am no more worthy to be called thy son: make me as one of thy hired servants.
LUKE|15|20|And he arose, and came to his father. But when he was yet a great way off, his father saw him, and had compassion, and ran, and fell on his neck, and kissed him.
LUKE|15|21|And the son said unto him, Father, I have sinned against heaven, and in thy sight, and am no more worthy to be called thy son.
LUKE|15|22|But the father said to his servants, Bring forth the best robe, and put it on him; and put a ring on his hand, and shoes on his feet:
LUKE|15|23|And bring hither the fatted calf, and kill it; and let us eat, and be merry:
LUKE|15|24|For this my son was dead, and is alive again; he was lost, and is found. And they began to be merry.
LUKE|15|25|Now his elder son was in the field: and as he came and drew nigh to the house, he heard musick and dancing.
LUKE|15|26|And he called one of the servants, and asked what these things meant.
LUKE|15|27|And he said unto him, Thy brother is come; and thy father hath killed the fatted calf, because he hath received him safe and sound.
LUKE|15|28|And he was angry, and would not go in: therefore came his father out, and intreated him.
LUKE|15|29|And he answering said to his father, Lo, these many years do I serve thee, neither transgressed I at any time thy commandment: and yet thou never gavest me a kid, that I might make merry with my friends:
LUKE|15|30|But as soon as this thy son was come, which hath devoured thy living with harlots, thou hast killed for him the fatted calf.
LUKE|15|31|And he said unto him, Son, thou art ever with me, and all that I have is thine.
LUKE|15|32|It was meet that we should make merry, and be glad: for this thy brother was dead, and is alive again; and was lost, and is found.
LUKE|16|1|And he said also unto his disciples, There was a certain rich man, which had a steward; and the same was accused unto him that he had wasted his goods.
LUKE|16|2|And he called him, and said unto him, How is it that I hear this of thee? give an account of thy stewardship; for thou mayest be no longer steward.
LUKE|16|3|Then the steward said within himself, What shall I do? for my lord taketh away from me the stewardship: I cannot dig; to beg I am ashamed.
LUKE|16|4|I am resolved what to do, that, when I am put out of the stewardship, they may receive me into their houses.
LUKE|16|5|So he called every one of his lord's debtors unto him, and said unto the first, How much owest thou unto my lord?
LUKE|16|6|And he said, An hundred measures of oil. And he said unto him, Take thy bill, and sit down quickly, and write fifty.
LUKE|16|7|Then said he to another, And how much owest thou? And he said, An hundred measures of wheat. And he said unto him, Take thy bill, and write fourscore.
LUKE|16|8|And the lord commended the unjust steward, because he had done wisely: for the children of this world are in their generation wiser than the children of light.
LUKE|16|9|And I say unto you, Make to yourselves friends of the mammon of unrighteousness; that, when ye fail, they may receive you into everlasting habitations.
LUKE|16|10|He that is faithful in that which is least is faithful also in much: and he that is unjust in the least is unjust also in much.
LUKE|16|11|If therefore ye have not been faithful in the unrighteous mammon, who will commit to your trust the true riches?
LUKE|16|12|And if ye have not been faithful in that which is another man's, who shall give you that which is your own?
LUKE|16|13|No servant can serve two masters: for either he will hate the one, and love the other; or else he will hold to the one, and despise the other. Ye cannot serve God and mammon.
LUKE|16|14|And the Pharisees also, who were covetous, heard all these things: and they derided him.
LUKE|16|15|And he said unto them, Ye are they which justify yourselves before men; but God knoweth your hearts: for that which is highly esteemed among men is abomination in the sight of God.
LUKE|16|16|The law and the prophets were until John: since that time the kingdom of God is preached, and every man presseth into it.
LUKE|16|17|And it is easier for heaven and earth to pass, than one tittle of the law to fail.
LUKE|16|18|Whosoever putteth away his wife, and marrieth another, committeth adultery: and whosoever marrieth her that is put away from her husband committeth adultery.
LUKE|16|19|There was a certain rich man, which was clothed in purple and fine linen, and fared sumptuously every day:
LUKE|16|20|And there was a certain beggar named Lazarus, which was laid at his gate, full of sores,
LUKE|16|21|And desiring to be fed with the crumbs which fell from the rich man's table: moreover the dogs came and licked his sores.
LUKE|16|22|And it came to pass, that the beggar died, and was carried by the angels into Abraham's bosom: the rich man also died, and was buried;
LUKE|16|23|And in hell he lift up his eyes, being in torments, and seeth Abraham afar off, and Lazarus in his bosom.
LUKE|16|24|And he cried and said, Father Abraham, have mercy on me, and send Lazarus, that he may dip the tip of his finger in water, and cool my tongue; for I am tormented in this flame.
LUKE|16|25|But Abraham said, Son, remember that thou in thy lifetime receivedst thy good things, and likewise Lazarus evil things: but now he is comforted, and thou art tormented.
LUKE|16|26|And beside all this, between us and you there is a great gulf fixed: so that they which would pass from hence to you cannot; neither can they pass to us, that would come from thence.
LUKE|16|27|Then he said, I pray thee therefore, father, that thou wouldest send him to my father's house:
LUKE|16|28|For I have five brethren; that he may testify unto them, lest they also come into this place of torment.
LUKE|16|29|Abraham saith unto him, They have Moses and the prophets; let them hear them.
LUKE|16|30|And he said, Nay, father Abraham: but if one went unto them from the dead, they will repent.
LUKE|16|31|And he said unto him, If they hear not Moses and the prophets, neither will they be persuaded, though one rose from the dead.
LUKE|17|1|Then said he unto the disciples, It is impossible but that offences will come: but woe unto him, through whom they come!
LUKE|17|2|It were better for him that a millstone were hanged about his neck, and he cast into the sea, than that he should offend one of these little ones.
LUKE|17|3|Take heed to yourselves: If thy brother trespass against thee, rebuke him; and if he repent, forgive him.
LUKE|17|4|And if he trespass against thee seven times in a day, and seven times in a day turn again to thee, saying, I repent; thou shalt forgive him.
LUKE|17|5|And the apostles said unto the Lord, Increase our faith.
LUKE|17|6|And the Lord said, If ye had faith as a grain of mustard seed, ye might say unto this sycamine tree, Be thou plucked up by the root, and be thou planted in the sea; and it should obey you.
LUKE|17|7|But which of you, having a servant plowing or feeding cattle, will say unto him by and by, when he is come from the field, Go and sit down to meat?
LUKE|17|8|And will not rather say unto him, Make ready wherewith I may sup, and gird thyself, and serve me, till I have eaten and drunken; and afterward thou shalt eat and drink?
LUKE|17|9|Doth he thank that servant because he did the things that were commanded him? I trow not.
LUKE|17|10|So likewise ye, when ye shall have done all those things which are commanded you, say, We are unprofitable servants: we have done that which was our duty to do.
LUKE|17|11|And it came to pass, as he went to Jerusalem, that he passed through the midst of Samaria and Galilee.
LUKE|17|12|And as he entered into a certain village, there met him ten men that were lepers, which stood afar off:
LUKE|17|13|And they lifted up their voices, and said, Jesus, Master, have mercy on us.
LUKE|17|14|And when he saw them, he said unto them, Go shew yourselves unto the priests. And it came to pass, that, as they went, they were cleansed.
LUKE|17|15|And one of them, when he saw that he was healed, turned back, and with a loud voice glorified God,
LUKE|17|16|And fell down on his face at his feet, giving him thanks: and he was a Samaritan.
LUKE|17|17|And Jesus answering said, Were there not ten cleansed? but where are the nine?
LUKE|17|18|There are not found that returned to give glory to God, save this stranger.
LUKE|17|19|And he said unto him, Arise, go thy way: thy faith hath made thee whole.
LUKE|17|20|And when he was demanded of the Pharisees, when the kingdom of God should come, he answered them and said, The kingdom of God cometh not with observation:
LUKE|17|21|Neither shall they say, Lo here! or, lo there! for, behold, the kingdom of God is within you.
LUKE|17|22|And he said unto the disciples, The days will come, when ye shall desire to see one of the days of the Son of man, and ye shall not see it.
LUKE|17|23|And they shall say to you, See here; or, see there: go not after them, nor follow them.
LUKE|17|24|For as the lightning, that lighteneth out of the one part under heaven, shineth unto the other part under heaven; so shall also the Son of man be in his day.
LUKE|17|25|But first must he suffer many things, and be rejected of this generation.
LUKE|17|26|And as it was in the days of Noe, so shall it be also in the days of the Son of man.
LUKE|17|27|They did eat, they drank, they married wives, they were given in marriage, until the day that Noe entered into the ark, and the flood came, and destroyed them all.
LUKE|17|28|Likewise also as it was in the days of Lot; they did eat, they drank, they bought, they sold, they planted, they builded;
LUKE|17|29|But the same day that Lot went out of Sodom it rained fire and brimstone from heaven, and destroyed them all.
LUKE|17|30|Even thus shall it be in the day when the Son of man is revealed.
LUKE|17|31|In that day, he which shall be upon the housetop, and his stuff in the house, let him not come down to take it away: and he that is in the field, let him likewise not return back.
LUKE|17|32|Remember Lot's wife.
LUKE|17|33|Whosoever shall seek to save his life shall lose it; and whosoever shall lose his life shall preserve it.
LUKE|17|34|I tell you, in that night there shall be two men in one bed; the one shall be taken, and the other shall be left.
LUKE|17|35|Two women shall be grinding together; the one shall be taken, and the other left.
LUKE|17|36|Two men shall be in the field; the one shall be taken, and the other left.
LUKE|17|37|And they answered and said unto him, Where, Lord? And he said unto them, Wheresoever the body is, thither will the eagles be gathered together.
LUKE|18|1|And he spake a parable unto them to this end, that men ought always to pray, and not to faint;
LUKE|18|2|Saying, There was in a city a judge, which feared not God, neither regarded man:
LUKE|18|3|And there was a widow in that city; and she came unto him, saying, Avenge me of mine adversary.
LUKE|18|4|And he would not for a while: but afterward he said within himself, Though I fear not God, nor regard man;
LUKE|18|5|Yet because this widow troubleth me, I will avenge her, lest by her continual coming she weary me.
LUKE|18|6|And the Lord said, Hear what the unjust judge saith.
LUKE|18|7|And shall not God avenge his own elect, which cry day and night unto him, though he bear long with them?
LUKE|18|8|I tell you that he will avenge them speedily. Nevertheless when the Son of man cometh, shall he find faith on the earth?
LUKE|18|9|And he spake this parable unto certain which trusted in themselves that they were righteous, and despised others:
LUKE|18|10|Two men went up into the temple to pray; the one a Pharisee, and the other a publican.
LUKE|18|11|The Pharisee stood and prayed thus with himself, God, I thank thee, that I am not as other men are, extortioners, unjust, adulterers, or even as this publican.
LUKE|18|12|I fast twice in the week, I give tithes of all that I possess.
LUKE|18|13|And the publican, standing afar off, would not lift up so much as his eyes unto heaven, but smote upon his breast, saying, God be merciful to me a sinner.
LUKE|18|14|I tell you, this man went down to his house justified rather than the other: for every one that exalteth himself shall be abased; and he that humbleth himself shall be exalted.
LUKE|18|15|And they brought unto him also infants, that he would touch them: but when his disciples saw it, they rebuked them.
LUKE|18|16|But Jesus called them unto him, and said, Suffer little children to come unto me, and forbid them not: for of such is the kingdom of God.
LUKE|18|17|Verily I say unto you, Whosoever shall not receive the kingdom of God as a little child shall in no wise enter therein.
LUKE|18|18|And a certain ruler asked him, saying, Good Master, what shall I do to inherit eternal life?
LUKE|18|19|And Jesus said unto him, Why callest thou me good? none is good, save one, that is, God.
LUKE|18|20|Thou knowest the commandments, Do not commit adultery, Do not kill, Do not steal, Do not bear false witness, Honour thy father and thy mother.
LUKE|18|21|And he said, All these have I kept from my youth up.
LUKE|18|22|Now when Jesus heard these things, he said unto him, Yet lackest thou one thing: sell all that thou hast, and distribute unto the poor, and thou shalt have treasure in heaven: and come, follow me.
LUKE|18|23|And when he heard this, he was very sorrowful: for he was very rich.
LUKE|18|24|And when Jesus saw that he was very sorrowful, he said, How hardly shall they that have riches enter into the kingdom of God!
LUKE|18|25|For it is easier for a camel to go through a needle's eye, than for a rich man to enter into the kingdom of God.
LUKE|18|26|And they that heard it said, Who then can be saved?
LUKE|18|27|And he said, The things which are impossible with men are possible with God.
LUKE|18|28|Then Peter said, Lo, we have left all, and followed thee.
LUKE|18|29|And he said unto them, Verily I say unto you, There is no man that hath left house, or parents, or brethren, or wife, or children, for the kingdom of God's sake,
LUKE|18|30|Who shall not receive manifold more in this present time, and in the world to come life everlasting.
LUKE|18|31|Then he took unto him the twelve, and said unto them, Behold, we go up to Jerusalem, and all things that are written by the prophets concerning the Son of man shall be accomplished.
LUKE|18|32|For he shall be delivered unto the Gentiles, and shall be mocked, and spitefully entreated, and spitted on:
LUKE|18|33|And they shall scourge him, and put him to death: and the third day he shall rise again.
LUKE|18|34|And they understood none of these things: and this saying was hid from them, neither knew they the things which were spoken.
LUKE|18|35|And it came to pass, that as he was come nigh unto Jericho, a certain blind man sat by the way side begging:
LUKE|18|36|And hearing the multitude pass by, he asked what it meant.
LUKE|18|37|And they told him, that Jesus of Nazareth passeth by.
LUKE|18|38|And he cried, saying, Jesus, thou son of David, have mercy on me.
LUKE|18|39|And they which went before rebuked him, that he should hold his peace: but he cried so much the more, Thou son of David, have mercy on me.
LUKE|18|40|And Jesus stood, and commanded him to be brought unto him: and when he was come near, he asked him,
LUKE|18|41|Saying, What wilt thou that I shall do unto thee? And he said, Lord, that I may receive my sight.
LUKE|18|42|And Jesus said unto him, Receive thy sight: thy faith hath saved thee.
LUKE|18|43|And immediately he received his sight, and followed him, glorifying God: and all the people, when they saw it, gave praise unto God.
LUKE|19|1|And Jesus entered and passed through Jericho.
LUKE|19|2|And, behold, there was a man named Zacchaeus, which was the chief among the publicans, and he was rich.
LUKE|19|3|And he sought to see Jesus who he was; and could not for the press, because he was little of stature.
LUKE|19|4|And he ran before, and climbed up into a sycomore tree to see him: for he was to pass that way.
LUKE|19|5|And when Jesus came to the place, he looked up, and saw him, and said unto him, Zacchaeus, make haste, and come down; for to day I must abide at thy house.
LUKE|19|6|And he made haste, and came down, and received him joyfully.
LUKE|19|7|And when they saw it, they all murmured, saying, That he was gone to be guest with a man that is a sinner.
LUKE|19|8|And Zacchaeus stood, and said unto the Lord: Behold, Lord, the half of my goods I give to the poor; and if I have taken any thing from any man by false accusation, I restore him fourfold.
LUKE|19|9|And Jesus said unto him, This day is salvation come to this house, forsomuch as he also is a son of Abraham.
LUKE|19|10|For the Son of man is come to seek and to save that which was lost.
LUKE|19|11|And as they heard these things, he added and spake a parable, because he was nigh to Jerusalem, and because they thought that the kingdom of God should immediately appear.
LUKE|19|12|He said therefore, A certain nobleman went into a far country to receive for himself a kingdom, and to return.
LUKE|19|13|And he called his ten servants, and delivered them ten pounds, and said unto them, Occupy till I come.
LUKE|19|14|But his citizens hated him, and sent a message after him, saying, We will not have this man to reign over us.
LUKE|19|15|And it came to pass, that when he was returned, having received the kingdom, then he commanded these servants to be called unto him, to whom he had given the money, that he might know how much every man had gained by trading.
LUKE|19|16|Then came the first, saying, Lord, thy pound hath gained ten pounds.
LUKE|19|17|And he said unto him, Well, thou good servant: because thou hast been faithful in a very little, have thou authority over ten cities.
LUKE|19|18|And the second came, saying, Lord, thy pound hath gained five pounds.
LUKE|19|19|And he said likewise to him, Be thou also over five cities.
LUKE|19|20|And another came, saying, Lord, behold, here is thy pound, which I have kept laid up in a napkin:
LUKE|19|21|For I feared thee, because thou art an austere man: thou takest up that thou layedst not down, and reapest that thou didst not sow.
LUKE|19|22|And he saith unto him, Out of thine own mouth will I judge thee, thou wicked servant. Thou knewest that I was an austere man, taking up that I laid not down, and reaping that I did not sow:
LUKE|19|23|Wherefore then gavest not thou my money into the bank, that at my coming I might have required mine own with usury?
LUKE|19|24|And he said unto them that stood by, Take from him the pound, and give it to him that hath ten pounds.
LUKE|19|25|(And they said unto him, Lord, he hath ten pounds.)
LUKE|19|26|For I say unto you, That unto every one which hath shall be given; and from him that hath not, even that he hath shall be taken away from him.
LUKE|19|27|But those mine enemies, which would not that I should reign over them, bring hither, and slay them before me.
LUKE|19|28|And when he had thus spoken, he went before, ascending up to Jerusalem.
LUKE|19|29|And it came to pass, when he was come nigh to Bethphage and Bethany, at the mount called the mount of Olives, he sent two of his disciples,
LUKE|19|30|Saying, Go ye into the village over against you; in the which at your entering ye shall find a colt tied, whereon yet never man sat: loose him, and bring him hither.
LUKE|19|31|And if any man ask you, Why do ye loose him? thus shall ye say unto him, Because the Lord hath need of him.
LUKE|19|32|And they that were sent went their way, and found even as he had said unto them.
LUKE|19|33|And as they were loosing the colt, the owners thereof said unto them, Why loose ye the colt?
LUKE|19|34|And they said, The Lord hath need of him.
LUKE|19|35|And they brought him to Jesus: and they cast their garments upon the colt, and they set Jesus thereon.
LUKE|19|36|And as he went, they spread their clothes in the way.
LUKE|19|37|And when he was come nigh, even now at the descent of the mount of Olives, the whole multitude of the disciples began to rejoice and praise God with a loud voice for all the mighty works that they had seen;
LUKE|19|38|Saying, Blessed be the King that cometh in the name of the Lord: peace in heaven, and glory in the highest.
LUKE|19|39|And some of the Pharisees from among the multitude said unto him, Master, rebuke thy disciples.
LUKE|19|40|And he answered and said unto them, I tell you that, if these should hold their peace, the stones would immediately cry out.
LUKE|19|41|And when he was come near, he beheld the city, and wept over it,
LUKE|19|42|Saying, If thou hadst known, even thou, at least in this thy day, the things which belong unto thy peace! but now they are hid from thine eyes.
LUKE|19|43|For the days shall come upon thee, that thine enemies shall cast a trench about thee, and compass thee round, and keep thee in on every side,
LUKE|19|44|And shall lay thee even with the ground, and thy children within thee; and they shall not leave in thee one stone upon another; because thou knewest not the time of thy visitation.
LUKE|19|45|And he went into the temple, and began to cast out them that sold therein, and them that bought;
LUKE|19|46|Saying unto them, It is written, My house is the house of prayer: but ye have made it a den of thieves.
LUKE|19|47|And he taught daily in the temple. But the chief priests and the scribes and the chief of the people sought to destroy him,
LUKE|19|48|And could not find what they might do: for all the people were very attentive to hear him.
LUKE|20|1|And it came to pass, that on one of those days, as he taught the people in the temple, and preached the gospel, the chief priests and the scribes came upon him with the elders,
LUKE|20|2|And spake unto him, saying, Tell us, by what authority doest thou these things? or who is he that gave thee this authority?
LUKE|20|3|And he answered and said unto them, I will also ask you one thing; and answer me:
LUKE|20|4|The baptism of John, was it from heaven, or of men?
LUKE|20|5|And they reasoned with themselves, saying, If we shall say, From heaven; he will say, Why then believed ye him not?
LUKE|20|6|But and if we say, Of men; all the people will stone us: for they be persuaded that John was a prophet.
LUKE|20|7|And they answered, that they could not tell whence it was.
LUKE|20|8|And Jesus said unto them, Neither tell I you by what authority I do these things.
LUKE|20|9|Then began he to speak to the people this parable; A certain man planted a vineyard, and let it forth to husbandmen, and went into a far country for a long time.
LUKE|20|10|And at the season he sent a servant to the husbandmen, that they should give him of the fruit of the vineyard: but the husbandmen beat him, and sent him away empty.
LUKE|20|11|And again he sent another servant: and they beat him also, and entreated him shamefully, and sent him away empty.
LUKE|20|12|And again he sent a third: and they wounded him also, and cast him out.
LUKE|20|13|Then said the lord of the vineyard, What shall I do? I will send my beloved son: it may be they will reverence him when they see him.
LUKE|20|14|But when the husbandmen saw him, they reasoned among themselves, saying, This is the heir: come, let us kill him, that the inheritance may be ours.
LUKE|20|15|So they cast him out of the vineyard, and killed him. What therefore shall the lord of the vineyard do unto them?
LUKE|20|16|He shall come and destroy these husbandmen, and shall give the vineyard to others. And when they heard it, they said, God forbid.
LUKE|20|17|And he beheld them, and said, What is this then that is written, The stone which the builders rejected, the same is become the head of the corner?
LUKE|20|18|Whosoever shall fall upon that stone shall be broken; but on whomsoever it shall fall, it will grind him to powder.
LUKE|20|19|And the chief priests and the scribes the same hour sought to lay hands on him; and they feared the people: for they perceived that he had spoken this parable against them.
LUKE|20|20|And they watched him, and sent forth spies, which should feign themselves just men, that they might take hold of his words, that so they might deliver him unto the power and authority of the governor.
LUKE|20|21|And they asked him, saying, Master, we know that thou sayest and teachest rightly, neither acceptest thou the person of any, but teachest the way of God truly:
LUKE|20|22|Is it lawful for us to give tribute unto Caesar, or no?
LUKE|20|23|But he perceived their craftiness, and said unto them, Why tempt ye me?
LUKE|20|24|Shew me a penny. Whose image and superscription hath it? They answered and said, Caesar's.
LUKE|20|25|And he said unto them, Render therefore unto Caesar the things which be Caesar's, and unto God the things which be God's.
LUKE|20|26|And they could not take hold of his words before the people: and they marvelled at his answer, and held their peace.
LUKE|20|27|Then came to him certain of the Sadducees, which deny that there is any resurrection; and they asked him,
LUKE|20|28|Saying, Master, Moses wrote unto us, If any man's brother die, having a wife, and he die without children, that his brother should take his wife, and raise up seed unto his brother.
LUKE|20|29|There were therefore seven brethren: and the first took a wife, and died without children.
LUKE|20|30|And the second took her to wife, and he died childless.
LUKE|20|31|And the third took her; and in like manner the seven also: and they left no children, and died.
LUKE|20|32|Last of all the woman died also.
LUKE|20|33|Therefore in the resurrection whose wife of them is she? for seven had her to wife.
LUKE|20|34|And Jesus answering said unto them, The children of this world marry, and are given in marriage:
LUKE|20|35|But they which shall be accounted worthy to obtain that world, and the resurrection from the dead, neither marry, nor are given in marriage:
LUKE|20|36|Neither can they die any more: for they are equal unto the angels; and are the children of God, being the children of the resurrection.
LUKE|20|37|Now that the dead are raised, even Moses shewed at the bush, when he calleth the Lord the God of Abraham, and the God of Isaac, and the God of Jacob.
LUKE|20|38|For he is not a God of the dead, but of the living: for all live unto him.
LUKE|20|39|Then certain of the scribes answering said, Master, thou hast well said.
LUKE|20|40|And after that they durst not ask him any question at all.
LUKE|20|41|And he said unto them, How say they that Christ is David's son?
LUKE|20|42|And David himself saith in the book of Psalms, The LORD said unto my Lord, Sit thou on my right hand,
LUKE|20|43|Till I make thine enemies thy footstool.
LUKE|20|44|David therefore calleth him Lord, how is he then his son?
LUKE|20|45|Then in the audience of all the people he said unto his disciples,
LUKE|20|46|Beware of the scribes, which desire to walk in long robes, and love greetings in the markets, and the highest seats in the synagogues, and the chief rooms at feasts;
LUKE|20|47|Which devour widows' houses, and for a shew make long prayers: the same shall receive greater damnation.
LUKE|21|1|And he looked up, and saw the rich men casting their gifts into the treasury.
LUKE|21|2|And he saw also a certain poor widow casting in thither two mites.
LUKE|21|3|And he said, Of a truth I say unto you, that this poor widow hath cast in more than they all:
LUKE|21|4|For all these have of their abundance cast in unto the offerings of God: but she of her penury hath cast in all the living that she had.
LUKE|21|5|And as some spake of the temple, how it was adorned with goodly stones and gifts, he said,
LUKE|21|6|As for these things which ye behold, the days will come, in the which there shall not be left one stone upon another, that shall not be thrown down.
LUKE|21|7|And they asked him, saying, Master, but when shall these things be? and what sign will there be when these things shall come to pass?
LUKE|21|8|And he said, Take heed that ye be not deceived: for many shall come in my name, saying, I am Christ; and the time draweth near: go ye not therefore after them.
LUKE|21|9|But when ye shall hear of wars and commotions, be not terrified: for these things must first come to pass; but the end is not by and by.
LUKE|21|10|Then said he unto them, Nation shall rise against nation, and kingdom against kingdom:
LUKE|21|11|And great earthquakes shall be in divers places, and famines, and pestilences; and fearful sights and great signs shall there be from heaven.
LUKE|21|12|But before all these, they shall lay their hands on you, and persecute you, delivering you up to the synagogues, and into prisons, being brought before kings and rulers for my name's sake.
LUKE|21|13|And it shall turn to you for a testimony.
LUKE|21|14|Settle it therefore in your hearts, not to meditate before what ye shall answer:
LUKE|21|15|For I will give you a mouth and wisdom, which all your adversaries shall not be able to gainsay nor resist.
LUKE|21|16|And ye shall be betrayed both by parents, and brethren, and kinsfolks, and friends; and some of you shall they cause to be put to death.
LUKE|21|17|And ye shall be hated of all men for my name's sake.
LUKE|21|18|But there shall not an hair of your head perish.
LUKE|21|19|In your patience possess ye your souls.
LUKE|21|20|And when ye shall see Jerusalem compassed with armies, then know that the desolation thereof is nigh.
LUKE|21|21|Then let them which are in Judaea flee to the mountains; and let them which are in the midst of it depart out; and let not them that are in the countries enter thereinto.
LUKE|21|22|For these be the days of vengeance, that all things which are written may be fulfilled.
LUKE|21|23|But woe unto them that are with child, and to them that give suck, in those days! for there shall be great distress in the land, and wrath upon this people.
LUKE|21|24|And they shall fall by the edge of the sword, and shall be led away captive into all nations: and Jerusalem shall be trodden down of the Gentiles, until the times of the Gentiles be fulfilled.
LUKE|21|25|And there shall be signs in the sun, and in the moon, and in the stars; and upon the earth distress of nations, with perplexity; the sea and the waves roaring;
LUKE|21|26|Men's hearts failing them for fear, and for looking after those things which are coming on the earth: for the powers of heaven shall be shaken.
LUKE|21|27|And then shall they see the Son of man coming in a cloud with power and great glory.
LUKE|21|28|And when these things begin to come to pass, then look up, and lift up your heads; for your redemption draweth nigh.
LUKE|21|29|And he spake to them a parable; Behold the fig tree, and all the trees;
LUKE|21|30|When they now shoot forth, ye see and know of your own selves that summer is now nigh at hand.
LUKE|21|31|So likewise ye, when ye see these things come to pass, know ye that the kingdom of God is nigh at hand.
LUKE|21|32|Verily I say unto you, This generation shall not pass away, till all be fulfilled.
LUKE|21|33|Heaven and earth shall pass away: but my words shall not pass away.
LUKE|21|34|And take heed to yourselves, lest at any time your hearts be overcharged with surfeiting, and drunkenness, and cares of this life, and so that day come upon you unawares.
LUKE|21|35|For as a snare shall it come on all them that dwell on the face of the whole earth.
LUKE|21|36|Watch ye therefore, and pray always, that ye may be accounted worthy to escape all these things that shall come to pass, and to stand before the Son of man.
LUKE|21|37|And in the day time he was teaching in the temple; and at night he went out, and abode in the mount that is called the mount of Olives.
LUKE|21|38|And all the people came early in the morning to him in the temple, for to hear him.
LUKE|22|1|Now the feast of unleavened bread drew nigh, which is called the Passover.
LUKE|22|2|And the chief priests and scribes sought how they might kill him; for they feared the people.
LUKE|22|3|Then entered Satan into Judas surnamed Iscariot, being of the number of the twelve.
LUKE|22|4|And he went his way, and communed with the chief priests and captains, how he might betray him unto them.
LUKE|22|5|And they were glad, and covenanted to give him money.
LUKE|22|6|And he promised, and sought opportunity to betray him unto them in the absence of the multitude.
LUKE|22|7|Then came the day of unleavened bread, when the passover must be killed.
LUKE|22|8|And he sent Peter and John, saying, Go and prepare us the passover, that we may eat.
LUKE|22|9|And they said unto him, Where wilt thou that we prepare?
LUKE|22|10|And he said unto them, Behold, when ye are entered into the city, there shall a man meet you, bearing a pitcher of water; follow him into the house where he entereth in.
LUKE|22|11|And ye shall say unto the goodman of the house, The Master saith unto thee, Where is the guestchamber, where I shall eat the passover with my disciples?
LUKE|22|12|And he shall shew you a large upper room furnished: there make ready.
LUKE|22|13|And they went, and found as he had said unto them: and they made ready the passover.
LUKE|22|14|And when the hour was come, he sat down, and the twelve apostles with him.
LUKE|22|15|And he said unto them, With desire I have desired to eat this passover with you before I suffer:
LUKE|22|16|For I say unto you, I will not any more eat thereof, until it be fulfilled in the kingdom of God.
LUKE|22|17|And he took the cup, and gave thanks, and said, Take this, and divide it among yourselves:
LUKE|22|18|For I say unto you, I will not drink of the fruit of the vine, until the kingdom of God shall come.
LUKE|22|19|And he took bread, and gave thanks, and brake it, and gave unto them, saying, This is my body which is given for you: this do in remembrance of me.
LUKE|22|20|Likewise also the cup after supper, saying, This cup is the new testament in my blood, which is shed for you.
LUKE|22|21|But, behold, the hand of him that betrayeth me is with me on the table.
LUKE|22|22|And truly the Son of man goeth, as it was determined: but woe unto that man by whom he is betrayed!
LUKE|22|23|And they began to enquire among themselves, which of them it was that should do this thing.
LUKE|22|24|And there was also a strife among them, which of them should be accounted the greatest.
LUKE|22|25|And he said unto them, The kings of the Gentiles exercise lordship over them; and they that exercise authority upon them are called benefactors.
LUKE|22|26|But ye shall not be so: but he that is greatest among you, let him be as the younger; and he that is chief, as he that doth serve.
LUKE|22|27|For whether is greater, he that sitteth at meat, or he that serveth? is not he that sitteth at meat? but I am among you as he that serveth.
LUKE|22|28|Ye are they which have continued with me in my temptations.
LUKE|22|29|And I appoint unto you a kingdom, as my Father hath appointed unto me;
LUKE|22|30|That ye may eat and drink at my table in my kingdom, and sit on thrones judging the twelve tribes of Israel.
LUKE|22|31|And the Lord said, Simon, Simon, behold, Satan hath desired to have you, that he may sift you as wheat:
LUKE|22|32|But I have prayed for thee, that thy faith fail not: and when thou art converted, strengthen thy brethren.
LUKE|22|33|And he said unto him, Lord, I am ready to go with thee, both into prison, and to death.
LUKE|22|34|And he said, I tell thee, Peter, the cock shall not crow this day, before that thou shalt thrice deny that thou knowest me.
LUKE|22|35|And he said unto them, When I sent you without purse, and scrip, and shoes, lacked ye any thing? And they said, Nothing.
LUKE|22|36|Then said he unto them, But now, he that hath a purse, let him take it, and likewise his scrip: and he that hath no sword, let him sell his garment, and buy one.
LUKE|22|37|For I say unto you, that this that is written must yet be accomplished in me, And he was reckoned among the transgressors: for the things concerning me have an end.
LUKE|22|38|And they said, Lord, behold, here are two swords. And he said unto them, It is enough.
LUKE|22|39|And he came out, and went, as he was wont, to the mount of Olives; and his disciples also followed him.
LUKE|22|40|And when he was at the place, he said unto them, Pray that ye enter not into temptation.
LUKE|22|41|And he was withdrawn from them about a stone's cast, and kneeled down, and prayed,
LUKE|22|42|Saying, Father, if thou be willing, remove this cup from me: nevertheless not my will, but thine, be done.
LUKE|22|43|And there appeared an angel unto him from heaven, strengthening him.
LUKE|22|44|And being in an agony he prayed more earnestly: and his sweat was as it were great drops of blood falling down to the ground.
LUKE|22|45|And when he rose up from prayer, and was come to his disciples, he found them sleeping for sorrow,
LUKE|22|46|And said unto them, Why sleep ye? rise and pray, lest ye enter into temptation.
LUKE|22|47|And while he yet spake, behold a multitude, and he that was called Judas, one of the twelve, went before them, and drew near unto Jesus to kiss him.
LUKE|22|48|But Jesus said unto him, Judas, betrayest thou the Son of man with a kiss?
LUKE|22|49|When they which were about him saw what would follow, they said unto him, Lord, shall we smite with the sword?
LUKE|22|50|And one of them smote the servant of the high priest, and cut off his right ear.
LUKE|22|51|And Jesus answered and said, Suffer ye thus far. And he touched his ear, and healed him.
LUKE|22|52|Then Jesus said unto the chief priests, and captains of the temple, and the elders, which were come to him, Be ye come out, as against a thief, with swords and staves?
LUKE|22|53|When I was daily with you in the temple, ye stretched forth no hands against me: but this is your hour, and the power of darkness.
LUKE|22|54|Then took they him, and led him, and brought him into the high priest's house. And Peter followed afar off.
LUKE|22|55|And when they had kindled a fire in the midst of the hall, and were set down together, Peter sat down among them.
LUKE|22|56|But a certain maid beheld him as he sat by the fire, and earnestly looked upon him, and said, This man was also with him.
LUKE|22|57|And he denied him, saying, Woman, I know him not.
LUKE|22|58|And after a little while another saw him, and said, Thou art also of them. And Peter said, Man, I am not.
LUKE|22|59|And about the space of one hour after another confidently affirmed, saying, Of a truth this fellow also was with him: for he is a Galilaean.
LUKE|22|60|And Peter said, Man, I know not what thou sayest. And immediately, while he yet spake, the cock crew.
LUKE|22|61|And the Lord turned, and looked upon Peter. And Peter remembered the word of the Lord, how he had said unto him, Before the cock crow, thou shalt deny me thrice.
LUKE|22|62|And Peter went out, and wept bitterly.
LUKE|22|63|And the men that held Jesus mocked him, and smote him.
LUKE|22|64|And when they had blindfolded him, they struck him on the face, and asked him, saying, Prophesy, who is it that smote thee?
LUKE|22|65|And many other things blasphemously spake they against him.
LUKE|22|66|And as soon as it was day, the elders of the people and the chief priests and the scribes came together, and led him into their council, saying,
LUKE|22|67|Art thou the Christ? tell us. And he said unto them, If I tell you, ye will not believe:
LUKE|22|68|And if I also ask you, ye will not answer me, nor let me go.
LUKE|22|69|Hereafter shall the Son of man sit on the right hand of the power of God.
LUKE|22|70|Then said they all, Art thou then the Son of God? And he said unto them, Ye say that I am.
LUKE|22|71|And they said, What need we any further witness? for we ourselves have heard of his own mouth.
LUKE|23|1|And the whole multitude of them arose, and led him unto Pilate.
LUKE|23|2|And they began to accuse him, saying, We found this fellow perverting the nation, and forbidding to give tribute to Caesar, saying that he himself is Christ a King.
LUKE|23|3|And Pilate asked him, saying, Art thou the King of the Jews? And he answered him and said, Thou sayest it.
LUKE|23|4|Then said Pilate to the chief priests and to the people, I find no fault in this man.
LUKE|23|5|And they were the more fierce, saying, He stirreth up the people, teaching throughout all Jewry, beginning from Galilee to this place.
LUKE|23|6|When Pilate heard of Galilee, he asked whether the man were a Galilaean.
LUKE|23|7|And as soon as he knew that he belonged unto Herod's jurisdiction, he sent him to Herod, who himself also was at Jerusalem at that time.
LUKE|23|8|And when Herod saw Jesus, he was exceeding glad: for he was desirous to see him of a long season, because he had heard many things of him; and he hoped to have seen some miracle done by him.
LUKE|23|9|Then he questioned with him in many words; but he answered him nothing.
LUKE|23|10|And the chief priests and scribes stood and vehemently accused him.
LUKE|23|11|And Herod with his men of war set him at nought, and mocked him, and arrayed him in a gorgeous robe, and sent him again to Pilate.
LUKE|23|12|And the same day Pilate and Herod were made friends together: for before they were at enmity between themselves.
LUKE|23|13|And Pilate, when he had called together the chief priests and the rulers and the people,
LUKE|23|14|Said unto them, Ye have brought this man unto me, as one that perverteth the people: and, behold, I, having examined him before you, have found no fault in this man touching those things whereof ye accuse him:
LUKE|23|15|No, nor yet Herod: for I sent you to him; and, lo, nothing worthy of death is done unto him.
LUKE|23|16|I will therefore chastise him, and release him.
LUKE|23|17|(For of necessity he must release one unto them at the feast.)
LUKE|23|18|And they cried out all at once, saying, Away with this man, and release unto us Barabbas:
LUKE|23|19|(Who for a certain sedition made in the city, and for murder, was cast into prison.)
LUKE|23|20|Pilate therefore, willing to release Jesus, spake again to them.
LUKE|23|21|But they cried, saying, Crucify him, crucify him.
LUKE|23|22|And he said unto them the third time, Why, what evil hath he done? I have found no cause of death in him: I will therefore chastise him, and let him go.
LUKE|23|23|And they were instant with loud voices, requiring that he might be crucified. And the voices of them and of the chief priests prevailed.
LUKE|23|24|And Pilate gave sentence that it should be as they required.
LUKE|23|25|And he released unto them him that for sedition and murder was cast into prison, whom they had desired; but he delivered Jesus to their will.
LUKE|23|26|And as they led him away, they laid hold upon one Simon, a Cyrenian, coming out of the country, and on him they laid the cross, that he might bear it after Jesus.
LUKE|23|27|And there followed him a great company of people, and of women, which also bewailed and lamented him.
LUKE|23|28|But Jesus turning unto them said, Daughters of Jerusalem, weep not for me, but weep for yourselves, and for your children.
LUKE|23|29|For, behold, the days are coming, in the which they shall say, Blessed are the barren, and the wombs that never bare, and the paps which never gave suck.
LUKE|23|30|Then shall they begin to say to the mountains, Fall on us; and to the hills, Cover us.
LUKE|23|31|For if they do these things in a green tree, what shall be done in the dry?
LUKE|23|32|And there were also two other, malefactors, led with him to be put to death.
LUKE|23|33|And when they were come to the place, which is called Calvary, there they crucified him, and the malefactors, one on the right hand, and the other on the left.
LUKE|23|34|Then said Jesus, Father, forgive them; for they know not what they do. And they parted his raiment, and cast lots.
LUKE|23|35|And the people stood beholding. And the rulers also with them derided him, saying, He saved others; let him save himself, if he be Christ, the chosen of God.
LUKE|23|36|And the soldiers also mocked him, coming to him, and offering him vinegar,
LUKE|23|37|And saying, If thou be the king of the Jews, save thyself.
LUKE|23|38|And a superscription also was written over him in letters of Greek, and Latin, and Hebrew, THIS IS THE KING OF THE JEWS.
LUKE|23|39|And one of the malefactors which were hanged railed on him, saying, If thou be Christ, save thyself and us.
LUKE|23|40|But the other answering rebuked him, saying, Dost not thou fear God, seeing thou art in the same condemnation?
LUKE|23|41|And we indeed justly; for we receive the due reward of our deeds: but this man hath done nothing amiss.
LUKE|23|42|And he said unto Jesus, Lord, remember me when thou comest into thy kingdom.
LUKE|23|43|And Jesus said unto him, Verily I say unto thee, To day shalt thou be with me in paradise.
LUKE|23|44|And it was about the sixth hour, and there was a darkness over all the earth until the ninth hour.
LUKE|23|45|And the sun was darkened, and the veil of the temple was rent in the midst.
LUKE|23|46|And when Jesus had cried with a loud voice, he said, Father, into thy hands I commend my spirit: and having said thus, he gave up the ghost.
LUKE|23|47|Now when the centurion saw what was done, he glorified God, saying, Certainly this was a righteous man.
LUKE|23|48|And all the people that came together to that sight, beholding the things which were done, smote their breasts, and returned.
LUKE|23|49|And all his acquaintance, and the women that followed him from Galilee, stood afar off, beholding these things.
LUKE|23|50|And, behold, there was a man named Joseph, a counsellor; and he was a good man, and a just:
LUKE|23|51|(The same had not consented to the counsel and deed of them;) he was of Arimathaea, a city of the Jews: who also himself waited for the kingdom of God.
LUKE|23|52|This man went unto Pilate, and begged the body of Jesus.
LUKE|23|53|And he took it down, and wrapped it in linen, and laid it in a sepulchre that was hewn in stone, wherein never man before was laid.
LUKE|23|54|And that day was the preparation, and the sabbath drew on.
LUKE|23|55|And the women also, which came with him from Galilee, followed after, and beheld the sepulchre, and how his body was laid.
LUKE|23|56|And they returned, and prepared spices and ointments; and rested the sabbath day according to the commandment.
LUKE|24|1|Now upon the first day of the week, very early in the morning, they came unto the sepulchre, bringing the spices which they had prepared, and certain others with them.
LUKE|24|2|And they found the stone rolled away from the sepulchre.
LUKE|24|3|And they entered in, and found not the body of the Lord Jesus.
LUKE|24|4|And it came to pass, as they were much perplexed thereabout, behold, two men stood by them in shining garments:
LUKE|24|5|And as they were afraid, and bowed down their faces to the earth, they said unto them, Why seek ye the living among the dead?
LUKE|24|6|He is not here, but is risen: remember how he spake unto you when he was yet in Galilee,
LUKE|24|7|Saying, The Son of man must be delivered into the hands of sinful men, and be crucified, and the third day rise again.
LUKE|24|8|And they remembered his words,
LUKE|24|9|And returned from the sepulchre, and told all these things unto the eleven, and to all the rest.
LUKE|24|10|It was Mary Magdalene and Joanna, and Mary the mother of James, and other women that were with them, which told these things unto the apostles.
LUKE|24|11|And their words seemed to them as idle tales, and they believed them not.
LUKE|24|12|Then arose Peter, and ran unto the sepulchre; and stooping down, he beheld the linen clothes laid by themselves, and departed, wondering in himself at that which was come to pass.
LUKE|24|13|And, behold, two of them went that same day to a village called Emmaus, which was from Jerusalem about threescore furlongs.
LUKE|24|14|And they talked together of all these things which had happened.
LUKE|24|15|And it came to pass, that, while they communed together and reasoned, Jesus himself drew near, and went with them.
LUKE|24|16|But their eyes were holden that they should not know him.
LUKE|24|17|And he said unto them, What manner of communications are these that ye have one to another, as ye walk, and are sad?
LUKE|24|18|And the one of them, whose name was Cleopas, answering said unto him, Art thou only a stranger in Jerusalem, and hast not known the things which are come to pass there in these days?
LUKE|24|19|And he said unto them, What things? And they said unto him, Concerning Jesus of Nazareth, which was a prophet mighty in deed and word before God and all the people:
LUKE|24|20|And how the chief priests and our rulers delivered him to be condemned to death, and have crucified him.
LUKE|24|21|But we trusted that it had been he which should have redeemed Israel: and beside all this, to day is the third day since these things were done.
LUKE|24|22|Yea, and certain women also of our company made us astonished, which were early at the sepulchre;
LUKE|24|23|And when they found not his body, they came, saying, that they had also seen a vision of angels, which said that he was alive.
LUKE|24|24|And certain of them which were with us went to the sepulchre, and found it even so as the women had said: but him they saw not.
LUKE|24|25|Then he said unto them, O fools, and slow of heart to believe all that the prophets have spoken:
LUKE|24|26|Ought not Christ to have suffered these things, and to enter into his glory?
LUKE|24|27|And beginning at Moses and all the prophets, he expounded unto them in all the scriptures the things concerning himself.
LUKE|24|28|And they drew nigh unto the village, whither they went: and he made as though he would have gone further.
LUKE|24|29|But they constrained him, saying, Abide with us: for it is toward evening, and the day is far spent. And he went in to tarry with them.
LUKE|24|30|And it came to pass, as he sat at meat with them, he took bread, and blessed it, and brake, and gave to them.
LUKE|24|31|And their eyes were opened, and they knew him; and he vanished out of their sight.
LUKE|24|32|And they said one to another, Did not our heart burn within us, while he talked with us by the way, and while he opened to us the scriptures?
LUKE|24|33|And they rose up the same hour, and returned to Jerusalem, and found the eleven gathered together, and them that were with them,
LUKE|24|34|Saying, The Lord is risen indeed, and hath appeared to Simon.
LUKE|24|35|And they told what things were done in the way, and how he was known of them in breaking of bread.
LUKE|24|36|And as they thus spake, Jesus himself stood in the midst of them, and saith unto them, Peace be unto you.
LUKE|24|37|But they were terrified and affrighted, and supposed that they had seen a spirit.
LUKE|24|38|And he said unto them, Why are ye troubled? and why do thoughts arise in your hearts?
LUKE|24|39|Behold my hands and my feet, that it is I myself: handle me, and see; for a spirit hath not flesh and bones, as ye see me have.
LUKE|24|40|And when he had thus spoken, he shewed them his hands and his feet.
LUKE|24|41|And while they yet believed not for joy, and wondered, he said unto them, Have ye here any meat?
LUKE|24|42|And they gave him a piece of a broiled fish, and of an honeycomb.
LUKE|24|43|And he took it, and did eat before them.
LUKE|24|44|And he said unto them, These are the words which I spake unto you, while I was yet with you, that all things must be fulfilled, which were written in the law of Moses, and in the prophets, and in the psalms, concerning me.
LUKE|24|45|Then opened he their understanding, that they might understand the scriptures,
LUKE|24|46|And said unto them, Thus it is written, and thus it behoved Christ to suffer, and to rise from the dead the third day:
LUKE|24|47|And that repentance and remission of sins should be preached in his name among all nations, beginning at Jerusalem.
LUKE|24|48|And ye are witnesses of these things.
LUKE|24|49|And, behold, I send the promise of my Father upon you: but tarry ye in the city of Jerusalem, until ye be endued with power from on high.
LUKE|24|50|And he led them out as far as to Bethany, and he lifted up his hands, and blessed them.
LUKE|24|51|And it came to pass, while he blessed them, he was parted from them, and carried up into heaven.
LUKE|24|52|And they worshipped him, and returned to Jerusalem with great joy:
LUKE|24|53|And were continually in the temple, praising and blessing God. Amen.
