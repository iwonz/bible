PS|1|1|beatus vir qui non abiit in consilio impiorum et in via peccatorum non stetit et in cathedra pestilentiae non sedit
PS|1|2|sed in lege Domini voluntas eius et in lege eius meditabitur die ac nocte
PS|1|3|et erit tamquam lignum quod plantatum est secus decursus aquarum quod fructum suum dabit in tempore suo et folium eius non defluet et omnia quaecumque faciet prosperabuntur
PS|1|4|non sic impii non sic; sed tamquam pulvis quem proicit ventus a facie terrae;
PS|1|5|ideo non resurgent impii in iudicio neque peccatores in consilio iustorum
PS|1|6|quoniam novit Dominus viam iustorum et iter impiorum peribit
PS|2|1|psalmus David quare fremuerunt gentes et populi meditati sunt inania
PS|2|2|adstiterunt reges terrae et principes convenerunt in unum adversus Dominum et adversus christum eius diapsalma
PS|2|3|disrumpamus vincula eorum et proiciamus a nobis iugum ipsorum
PS|2|4|qui habitat in caelis inridebit eos et Dominus subsannabit eos
PS|2|5|tunc loquetur ad eos in ira sua et in furore suo conturbabit eos
PS|2|6|ego autem constitutus sum rex ab eo super Sion montem sanctum eius praedicans praeceptum eius
PS|2|7|Dominus dixit ad me filius meus es tu ego hodie genui te
PS|2|8|postula a me et dabo tibi gentes hereditatem tuam et possessionem tuam terminos terrae
PS|2|9|reges eos in virga ferrea tamquam vas figuli confringes eos
PS|2|10|et nunc reges intellegite erudimini qui iudicatis terram
PS|2|11|servite Domino in timore et exultate ei in tremore
PS|2|12|adprehendite disciplinam nequando irascatur Dominus et pereatis de via iusta
PS|2|13|cum exarserit in brevi ira eius beati omnes qui confidunt in eo
PS|3|1|psalmus David cum fugeret a facie Abessalon filii sui
PS|3|2|Domine quid multiplicati sunt qui tribulant me multi insurgunt adversum me
PS|3|3|multi dicunt animae meae non est salus ipsi in Deo eius; diapsalma
PS|3|4|tu autem Domine susceptor meus es gloria mea et exaltans caput meum
PS|3|5|voce mea ad Dominum clamavi et exaudivit me de monte sancto suo diapsalma
PS|3|6|ego dormivi et soporatus sum exsurrexi quia Dominus suscipiet me
PS|3|7|non timebo milia populi circumdantis me exsurge Domine salvum me fac Deus meus
PS|3|8|quoniam tu percussisti omnes adversantes mihi sine causa dentes peccatorum contrivisti
PS|3|9|Domini est salus et super populum tuum benedictio tua
PS|4|1|in finem in carminibus psalmus David
PS|4|2|cum invocarem exaudivit me Deus iustitiae meae in tribulatione dilatasti mihi miserere mei et exaudi orationem meam
PS|4|3|filii hominum usquequo gravi corde ut quid diligitis vanitatem et quaeritis mendacium diapsalma
PS|4|4|et scitote quoniam mirificavit Dominus sanctum suum Dominus exaudiet me cum clamavero ad eum
PS|4|5|irascimini et nolite peccare quae dicitis in cordibus vestris in cubilibus vestris conpungimini diapsalma
PS|4|6|sacrificate sacrificium iustitiae et sperate in Domino multi dicunt quis ostendet nobis bona
PS|4|7|signatum est super nos lumen vultus tui Domine dedisti laetitiam in corde meo
PS|4|8|a fructu frumenti et vini et olei sui multiplicati sunt
PS|4|9|in pace in id ipsum dormiam et requiescam
PS|4|10|quoniam tu Domine singulariter in spe constituisti me
PS|5|1|in finem pro ea quae hereditatem consequitur psalmus David
PS|5|2|verba mea auribus percipe Domine intellege clamorem meum
PS|5|3|intende voci orationis meae rex meus et Deus meus
PS|5|4|quoniam ad te orabo Domine mane exaudies vocem meam
PS|5|5|mane adstabo tibi et videbo quoniam non deus volens iniquitatem tu es
PS|5|6|neque habitabit iuxta te malignus neque permanebunt iniusti ante oculos tuos
PS|5|7|odisti omnes qui operantur iniquitatem perdes %omnes; qui loquuntur mendacium virum sanguinum et dolosum abominabitur Dominus
PS|5|8|ego autem in multitudine misericordiae tuae introibo in domum tuam adorabo ad templum sanctum tuum in timore tuo
PS|5|9|Domine deduc me in iustitia tua propter inimicos meos dirige in conspectu meo viam tuam
PS|5|10|quoniam non est in ore eorum veritas cor eorum vanum est
PS|5|11|sepulchrum patens est guttur eorum linguis suis dolose agebant iudica illos Deus decidant a cogitationibus suis secundum multitudinem impietatum eorum expelle eos quoniam inritaverunt te Domine
PS|5|12|et laetentur omnes qui sperant in te in aeternum exultabunt et habitabis in eis et gloriabuntur in te omnes qui diligunt nomen tuum
PS|5|13|quoniam tu benedices iusto Domine ut scuto bonae voluntatis coronasti nos
PS|6|1|in finem in carminibus pro octava psalmus David
PS|6|2|Domine ne in furore tuo arguas me neque in ira tua corripias me
PS|6|3|miserere mei Domine quoniam infirmus sum sana me Domine quoniam conturbata sunt ossa mea
PS|6|4|et anima mea turbata est valde et tu Domine usquequo
PS|6|5|convertere Domine eripe animam meam salvum me fac propter misericordiam tuam
PS|6|6|quoniam non est in morte qui memor sit tui in inferno autem quis confitebitur tibi
PS|6|7|laboravi in gemitu meo lavabo per singulas noctes lectum meum in lacrimis meis stratum meum rigabo
PS|6|8|turbatus est a furore oculus meus inveteravi inter omnes inimicos meos
PS|6|9|discedite a me omnes qui operamini iniquitatem quoniam exaudivit Dominus vocem fletus mei
PS|6|10|exaudivit Dominus deprecationem meam Dominus orationem meam suscepit
PS|6|11|erubescant et conturbentur vehementer omnes inimici mei convertantur et erubescant valde velociter
PS|7|1|psalmus David quem cantavit Domino pro verbis Chusi filii Iemini
PS|7|2|Domine Deus meus in te speravi salvum me fac ex omnibus persequentibus me et libera me
PS|7|3|nequando rapiat ut leo animam meam dum non est qui redimat neque qui salvum faciat
PS|7|4|Domine Deus meus si feci istud si est iniquitas in manibus meis
PS|7|5|si reddidi retribuentibus mihi mala decidam merito ab inimicis meis inanis
PS|7|6|persequatur inimicus animam meam et conprehendat et conculcet in terra vitam meam et gloriam meam in pulverem deducat diapsalma
PS|7|7|exsurge Domine in ira tua exaltare in finibus inimicorum meorum et exsurge Domine Deus meus in praecepto quod mandasti
PS|7|8|et synagoga populorum circumdabit te et propter hanc in altum regredere
PS|7|9|Dominus iudicat populos iudica me Domine secundum iustitiam meam et secundum innocentiam meam super me
PS|7|10|consummetur nequitia peccatorum et diriges iustum et scrutans corda et renes Deus
PS|7|11|iustum adiutorium meum a Deo qui salvos facit rectos corde
PS|7|12|Deus iudex iustus et fortis et patiens numquid irascitur per singulos dies
PS|7|13|nisi conversi fueritis gladium suum vibrabit arcum suum tetendit et paravit illum
PS|7|14|et in eo paravit vasa mortis sagittas suas ardentibus effecit
PS|7|15|ecce parturiit iniustitiam et; concepit dolorem et peperit iniquitatem
PS|7|16|lacum aperuit et effodit eum et incidet in foveam quam fecit
PS|7|17|convertetur dolor eius in caput eius et in verticem ipsius iniquitas eius descendet
PS|7|18|confitebor Domino secundum iustitiam eius et psallam nomini Domini altissimi
PS|8|1|in finem pro torcularibus psalmus David
PS|8|2|Domine Dominus noster quam admirabile est nomen tuum in universa terra quoniam elevata est magnificentia tua super caelos
PS|8|3|ex ore infantium et lactantium perfecisti laudem propter inimicos tuos ut destruas inimicum et ultorem
PS|8|4|quoniam videbo caelos tuos; opera digitorum tuorum lunam et stellas quae tu fundasti
PS|8|5|quid est homo quod memor es eius aut filius hominis quoniam visitas eum
PS|8|6|minuisti eum paulo minus ab angelis gloria et honore coronasti eum
PS|8|7|et constituisti eum super opera manuum tuarum
PS|8|8|omnia subiecisti sub pedibus eius oves et boves universas insuper et pecora campi
PS|8|9|volucres caeli et pisces maris qui perambulant semitas maris
PS|8|10|Domine Dominus noster quam admirabile est nomen tuum in universa terra
PS|9|1|in finem pro occultis filii psalmus David
PS|9|2|confitebor tibi Domine in toto corde meo narrabo omnia mirabilia tua
PS|9|3|laetabor et exultabo in te psallam nomini tuo Altissime
PS|9|4|in convertendo inimicum meum retrorsum infirmabuntur et peribunt a facie tua
PS|9|5|quoniam fecisti iudicium meum et causam meam sedisti super thronum qui iudicas iustitiam
PS|9|6|increpasti gentes %et; periit impius nomen eorum delisti in aeternum et in saeculum %saeculi;
PS|9|7|inimici defecerunt frameae in finem et civitates destruxisti periit memoria eorum cum sonitu
PS|9|8|et Dominus in aeternum permanet paravit in iudicio thronum suum
PS|9|9|et ipse iudicabit orbem terrae in aequitate iudicabit populos in iustitia
PS|9|10|et factus est Dominus refugium pauperi adiutor in oportunitatibus in tribulatione
PS|9|11|et sperent in te qui noverunt nomen tuum quoniam non dereliquisti quaerentes te Domine
PS|9|12|psallite Domino qui habitat in Sion adnuntiate inter gentes studia eius
PS|9|13|quoniam requirens sanguinem eorum recordatus est non est oblitus clamorem pauperum
PS|9|14|miserere mei Domine vide humilitatem meam de inimicis meis
PS|9|15|qui exaltas me de portis mortis ut adnuntiem omnes laudationes tuas in portis filiae Sion
PS|9|16|exultabo in salutari tuo infixae sunt gentes in interitu quem fecerunt in laqueo isto quem absconderunt conprehensus est pes eorum
PS|9|17|cognoscitur Dominus iudicia faciens in operibus manuum suarum conprehensus est peccator canticum diapsalmatis
PS|9|18|convertantur peccatores in infernum omnes gentes quae obliviscuntur Deum
PS|9|19|quoniam non in finem oblivio erit pauperis patientia pauperum non peribit in finem
PS|9|20|exsurge Domine non confortetur homo iudicentur gentes in conspectu tuo
PS|9|21|constitue Domine legislatorem super eos sciant gentes quoniam homines sunt diapsalma
PS|9|22|ut quid Domine recessisti longe dispicis in oportunitatibus in tribulatione
PS|9|23|dum superbit impius incenditur pauper conprehenduntur in consiliis quibus cogitant
PS|9|24|quoniam laudatur peccator in desideriis animae suae et iniquus benedicitur
PS|9|25|exacerbavit Dominum peccator secundum multitudinem irae suae non quaeret
PS|9|26|non est Deus in conspectu eius inquinatae sunt viae illius in omni tempore auferuntur iudicia tua a facie eius omnium inimicorum suorum dominabitur
PS|9|27|dixit enim in corde suo non movebor a generatione in generationem sine malo
PS|9|28|cuius maledictione os plenum est et amaritudine et dolo sub lingua eius labor et dolor
PS|9|29|sedet in insidiis cum divitibus in occultis ut interficiat innocentem
PS|9|30|oculi eius in pauperem respiciunt insidiatur in abscondito quasi leo in spelunca sua insidiatur ut rapiat pauperem rapere pauperem dum adtrahit eum
PS|9|31|in laqueo suo humiliabit eum inclinabit se et cadet cum dominatus fuerit pauperum
PS|9|32|dixit enim in corde suo oblitus est Deus avertit faciem suam ne videat in finem
PS|9|33|exsurge Domine Deus exaltetur manus tua ne obliviscaris pauperum
PS|9|34|propter quid inritavit impius Deum dixit enim in corde suo non requiret
PS|9|35|vides quoniam tu laborem et dolorem consideras ut tradas eos in manus tuas tibi derelictus est pauper orfano tu eras adiutor
PS|9|36|contere brachium peccatoris et maligni quaeretur peccatum illius et non invenietur
PS|9|37|Dominus regnabit in aeternum et in saeculum %saeculi; peribitis gentes de terra illius
PS|9|38|desiderium pauperum exaudivit Dominus praeparationem cordis eorum audivit auris tua
PS|9|39|iudicare pupillo et humili ut non adponat ultra magnificare se homo super terram
PS|10|1|in finem psalmus David
PS|10|2|in Domino confido quomodo dicitis animae meae transmigra in montes sicut passer
PS|10|3|quoniam ecce peccatores intenderunt arcum paraverunt sagittas suas in faretra ut sagittent in obscuro rectos corde
PS|10|4|quoniam quae perfecisti destruxerunt iustus %autem; quid fecit
PS|10|5|Dominus in templo sancto suo Dominus in caelo sedis eius oculi eius %in pauperem; respiciunt palpebrae eius interrogant filios hominum
PS|10|6|Dominus interrogat iustum et impium qui autem diligit iniquitatem odit animam suam
PS|10|7|pluet super peccatores laqueos ignis et sulphur et spiritus procellarum pars calicis eorum
PS|10|8|quoniam iustus Dominus %et; iustitias dilexit aequitatem vidit vultus eius
PS|11|1|in finem pro octava psalmus David
PS|11|2|salvum me fac Domine quoniam defecit sanctus quoniam deminutae sunt veritates a filiis hominum
PS|11|3|vana locuti sunt unusquisque ad proximum suum labia dolosa in corde et corde locuti sunt
PS|11|4|disperdat Dominus universa labia dolosa linguam magniloquam
PS|11|5|qui dixerunt linguam nostram magnificabimus labia nostra a nobis sunt quis noster dominus est
PS|11|6|propter miseriam inopum et gemitum pauperum nunc exsurgam dicit Dominus ponam in salutari fiducialiter agam in eo
PS|11|7|eloquia Domini eloquia casta argentum igne examinatum probatum terrae purgatum septuplum
PS|11|8|tu Domine servabis nos et custodies nos a generatione hac et in aeternum
PS|11|9|in circuitu impii ambulant secundum altitudinem tuam multiplicasti filios hominum
PS|12|1|in finem psalmus David usquequo Domine oblivisceris me in finem usquequo avertis faciem tuam a me
PS|12|2|quamdiu ponam consilia in anima mea dolorem in corde meo per diem
PS|12|3|usquequo exaltabitur inimicus meus super me
PS|12|4|respice exaudi me Domine Deus meus inlumina oculos meos ne umquam obdormiam in mortem
PS|12|5|nequando dicat inimicus meus praevalui adversus eum qui tribulant me exultabunt si motus fuero
PS|12|6|ego autem in misericordia tua speravi exultabit cor meum in salutari tuo cantabo Domino qui bona tribuit mihi et psallam nomini Domini altissimi
PS|13|1|in finem psalmus David dixit insipiens in corde suo non est Deus corrupti sunt et abominabiles facti sunt in studiis %suis; non est qui faciat bonum %non est usque ad unum;
PS|13|2|Dominus de caelo prospexit super filios hominum ut videat si est intellegens %aut; requirens Deum
PS|13|3|omnes declinaverunt simul inutiles facti sunt non est qui faciat bonum non est usque ad unum = sepulchrum patens est guttur eorum = linguis suis dolose agebant = venenum aspidum sub labiis eorum = quorum os maledictione et amaritudine plenum est = veloces pedes eorum ad effundendum sanguinem = contritio et infelicitas in viis eorum = et viam pacis non cognoverunt % non est timor Dei ante oculos eorum;
PS|13|4|nonne cognoscent omnes qui operantur iniquitatem qui devorant plebem meam sicut escam panis
PS|13|5|Dominum non invocaverunt illic trepidaverunt timore %ubi non erat timor;
PS|13|6|quoniam Deus in generatione iusta consilium inopis confudistis quoniam Dominus spes eius est
PS|13|7|quis dabit ex Sion salutare Israhel cum averterit Dominus captivitatem plebis suae exultabit Iacob et laetabitur Israhel
PS|14|1|psalmus David Domine quis habitabit in tabernaculo tuo aut quis requiescet in monte sancto tuo
PS|14|2|qui ingreditur sine macula et operatur iustitiam
PS|14|3|qui loquitur veritatem in corde suo qui non egit dolum in lingua sua nec fecit proximo suo malum et obprobrium non accepit adversus proximos suos
PS|14|4|ad nihilum deductus est in conspectu eius malignus timentes autem Dominum glorificat qui iurat proximo suo et non decipit
PS|14|5|qui pecuniam suam non dedit ad usuram et munera super innocentes non accepit qui facit haec non movebitur in aeternum
PS|15|1|tituli inscriptio ipsi David conserva me Domine quoniam in te speravi
PS|15|2|dixi Domino Dominus meus es tu quoniam bonorum meorum non eges
PS|15|3|sanctis qui sunt in terra eius mirificavit mihi; omnes voluntates meas in eis
PS|15|4|multiplicatae sunt infirmitates eorum postea adceleraverunt non congregabo conventicula eorum de sanguinibus nec memor ero nominum eorum per labia mea
PS|15|5|Dominus pars hereditatis meae et calicis mei tu es qui restitues hereditatem meam mihi
PS|15|6|funes ceciderunt mihi in praeclaris etenim hereditas mea praeclara est mihi
PS|15|7|benedicam Domino qui tribuit mihi intellectum insuper et usque ad noctem increpaverunt me renes mei
PS|15|8|providebam Dominum in conspectu meo semper quoniam a dextris est mihi ne commovear
PS|15|9|propter hoc laetatum est cor meum et exultavit lingua mea insuper et caro mea requiescet in spe
PS|15|10|quoniam non derelinques animam meam in inferno non dabis sanctum tuum videre corruptionem notas mihi fecisti vias vitae adimplebis me laetitia cum vultu tuo delectatio in dextera tua usque in finem
PS|16|1|oratio David exaudi Domine iustitiam meam intende deprecationem meam auribus percipe orationem meam non in labiis dolosis
PS|16|2|de vultu tuo iudicium meum prodeat oculi tui videant aequitates
PS|16|3|probasti cor meum visitasti nocte igne me examinasti et non est inventa in me iniquitas
PS|16|4|ut non loquatur os meum opera hominum propter verba labiorum tuorum ego custodivi vias duras
PS|16|5|perfice gressus meos in semitis tuis ut non moveantur vestigia mea
PS|16|6|ego clamavi quoniam exaudisti me Deus inclina aurem tuam mihi et exaudi verba mea
PS|16|7|mirifica misericordias tuas qui salvos facis sperantes in te
PS|16|8|a resistentibus dexterae tuae custodi me ut pupillam oculi sub umbra alarum tuarum proteges me
PS|16|9|a facie impiorum qui me adflixerunt inimici mei animam meam circumdederunt super me;
PS|16|10|adipem suum concluserunt os eorum locutum est superbia
PS|16|11|proicientes me nunc circumdederunt me oculos suos statuerunt declinare in terram
PS|16|12|susceperunt me sicut leo paratus ad praedam et sicut catulus leonis habitans in abditis
PS|16|13|exsurge Domine praeveni eum et subplanta eum eripe animam meam ab impio frameam tuam
PS|16|14|ab inimicis manus tuae Domine a paucis de terra divide eos in vita eorum de absconditis tuis adimpletus est venter eorum saturati sunt filiis et dimiserunt reliquias suas parvulis suis
PS|16|15|ego autem in iustitia apparebo conspectui tuo satiabor cum apparuerit gloria tua
PS|17|1|in finem puero Domini David quae locutus est Domino verba cantici huius in die qua eripuit eum Dominus de manu omnium inimicorum eius et de manu Saul et dixit
PS|17|2|diligam te Domine fortitudo mea
PS|17|3|Dominus firmamentum meum et refugium meum et liberator meus Deus meus adiutor meus et sperabo in eum protector meus et cornu salutis meae et susceptor meus
PS|17|4|laudans invocabo Dominum et ab inimicis meis salvus ero
PS|17|5|circumdederunt me dolores mortis et torrentes iniquitatis conturbaverunt me
PS|17|6|dolores inferni circumdederunt me praeoccupaverunt me laquei mortis
PS|17|7|cum tribularer invocavi Dominum et ad Deum meum clamavi exaudivit de templo %sancto; suo vocem meam et clamor meus in conspectu eius introibit in aures eius
PS|17|8|et commota est et contremuit terra et fundamenta montium conturbata sunt et commota sunt quoniam iratus est eis
PS|17|9|ascendit fumus in ira eius et ignis a facie eius exarsit carbones succensi sunt ab eo
PS|17|10|inclinavit caelos et descendit et caligo sub pedibus eius
PS|17|11|et ascendit super cherubin et volavit volavit super pinnas ventorum
PS|17|12|et posuit tenebras latibulum suum in circuitu eius tabernaculum eius tenebrosa aqua in nubibus aeris
PS|17|13|prae fulgore in conspectu eius nubes eius; transierunt grando et carbones ignis
PS|17|14|et intonuit de caelo Dominus et Altissimus dedit vocem suam grando et carbones ignis;
PS|17|15|et misit sagittas et dissipavit eos et fulgora multiplicavit et conturbavit eos
PS|17|16|et apparuerunt fontes aquarum et revelata sunt fundamenta orbis terrarum ab increpatione tua Domine ab inspiratione spiritus irae tuae
PS|17|17|misit de summo et accepit me adsumpsit me de aquis multis
PS|17|18|eripiet me de inimicis meis fortissimis et ab his qui oderunt me quoniam confirmati sunt super me
PS|17|19|praevenerunt me in die adflictionis meae et factus est Dominus protector meus
PS|17|20|et eduxit me in latitudinem salvum me faciet quoniam voluit me
PS|17|21|%et; retribuet mihi Dominus secundum iustitiam meam %et; secundum puritatem manuum mearum retribuet mihi
PS|17|22|quia custodivi vias Domini nec impie gessi a Deo meo
PS|17|23|quoniam omnia iudicia eius in conspectu meo sunt et iustitias eius non reppuli a me
PS|17|24|et ero inmaculatus cum eo et observabo ab iniquitate mea
PS|17|25|et retribuet mihi Dominus secundum iustitiam meam et secundum puritatem manuum mearum in conspectu oculorum eius
PS|17|26|cum sancto sanctus eris et cum viro innocente innocens eris
PS|17|27|et cum electo electus eris et cum perverso perverteris
PS|17|28|quoniam tu populum humilem salvum facies et oculos superborum humiliabis
PS|17|29|quoniam tu inluminas lucernam meam Domine Deus meus inluminas tenebras meas
PS|17|30|quoniam in te eripiar a temptatione et in Deo meo transgrediar murum
PS|17|31|Deus meus inpolluta via eius eloquia Domini igne examinata protector est omnium sperantium in eum
PS|17|32|quoniam quis deus praeter Dominum et quis deus praeter Deum nostrum
PS|17|33|Deus qui praecingit me virtute et posuit inmaculatam viam meam
PS|17|34|qui perfecit pedes meos tamquam cervorum et super excelsa statuens me
PS|17|35|qui doces manus meas in proelium et posuisti arcum aereum brachia mea
PS|17|36|et dedisti mihi protectionem salutis tuae et dextera tua suscepit me et disciplina tua correxit me in finem et disciplina tua ipsa me docebit
PS|17|37|dilatasti gressus meos subtus me et non sunt infirmata vestigia mea
PS|17|38|persequar inimicos meos et conprehendam illos et non convertar donec deficiant
PS|17|39|confringam illos nec poterunt stare cadent subtus pedes meos
PS|17|40|et praecinxisti me virtute ad bellum subplantasti insurgentes in me subtus me
PS|17|41|et inimicos meos dedisti mihi dorsum et odientes me disperdisti
PS|17|42|clamaverunt nec erat qui salvos faceret ad Dominum nec exaudivit eos
PS|17|43|et comminuam illos ut pulverem ante faciem venti ut lutum platearum delebo eos
PS|17|44|eripe me de contradictionibus populi constitues me in caput gentium
PS|17|45|populus quem non cognovi servivit mihi in auditu auris oboedivit mihi
PS|17|46|filii alieni mentiti sunt mihi filii alieni inveterati sunt et claudicaverunt a semitis suis
PS|17|47|vivit Dominus et benedictus Deus meus et exaltetur Deus salutis meae
PS|17|48|Deus qui dat vindictas mihi et subdidit populos sub me liberator meus de gentibus iracundis
PS|17|49|et ab insurgentibus in me exaltabis me a viro iniquo eripies me
PS|17|50|propterea confitebor tibi in nationibus Domine et psalmum dicam nomini tuo
PS|17|51|magnificans salutes regis eius et faciens misericordiam christo suo David et semini eius usque in saeculum
PS|18|1|in finem psalmus David
PS|18|2|caeli enarrant gloriam Dei et opera manuum eius adnuntiat firmamentum
PS|18|3|dies diei eructat verbum et nox nocti indicat scientiam
PS|18|4|non sunt loquellae neque sermones quorum non audiantur voces eorum
PS|18|5|in omnem terram exivit sonus eorum et in fines orbis terrae verba eorum
PS|18|6|in sole posuit tabernaculum suum et ipse tamquam sponsus procedens de thalamo suo exultavit ut gigans ad currendam viam %suam;
PS|18|7|a summo caeli egressio eius et occursus eius usque ad summum eius nec est qui se abscondat a calore eius
PS|18|8|lex Domini inmaculata convertens animas testimonium Domini fidele sapientiam praestans parvulis
PS|18|9|iustitiae Domini rectae laetificantes corda praeceptum Domini lucidum inluminans oculos
PS|18|10|timor Domini sanctus permanens in saeculum saeculi iudicia Domini vera iustificata in semet ipsa
PS|18|11|desiderabilia super aurum et lapidem pretiosum multum et dulciora super mel et favum
PS|18|12|etenim servus tuus custodit ea in custodiendis illis retributio multa
PS|18|13|delicta quis intellegit ab occultis meis munda me
PS|18|14|et ab alienis parce servo tuo si mei non fuerint dominati tunc inmaculatus ero et emundabor a delicto maximo
PS|18|15|et erunt ut conplaceant eloquia oris mei et meditatio cordis mei in conspectu tuo semper Domine adiutor meus et redemptor meus
PS|19|1|in finem psalmus David
PS|19|2|exaudiat te Dominus in die tribulationis protegat te nomen Dei Iacob
PS|19|3|mittat tibi auxilium de sancto et de Sion tueatur te
PS|19|4|memor sit omnis sacrificii tui et holocaustum tuum pingue fiat diapsalma
PS|19|5|tribuat tibi secundum cor tuum et omne consilium tuum confirmet
PS|19|6|laetabimur in salutari tuo et in nomine Dei nostri magnificabimur
PS|19|7|impleat Dominus omnes petitiones tuas nunc cognovi quoniam salvum fecit Dominus christum suum exaudiet illum de caelo sancto suo in potentatibus salus dexterae eius
PS|19|8|hii in curribus et hii in equis nos autem in nomine Domini Dei nostri invocabimus
PS|19|9|ipsi obligati sunt et ceciderunt nos vero surreximus et erecti sumus
PS|19|10|Domine salvum fac regem et exaudi nos in die qua invocaverimus te
PS|20|1|in finem psalmus David
PS|20|2|Domine in virtute tua laetabitur rex et super salutare tuum exultabit vehementer
PS|20|3|desiderium animae eius tribuisti ei et voluntate labiorum eius non fraudasti eum diapsalma
PS|20|4|quoniam praevenisti eum in benedictionibus dulcedinis posuisti in capite eius coronam de lapide pretioso
PS|20|5|vitam petiit a te et tribuisti ei longitudinem dierum in saeculum et in saeculum saeculi
PS|20|6|magna gloria eius in salutari tuo gloriam et magnum decorem inpones super eum
PS|20|7|quoniam dabis eum benedictionem in saeculum saeculi laetificabis eum in gaudio cum vultu tuo
PS|20|8|quoniam rex sperat in Domino et in misericordia Altissimi non commovebitur
PS|20|9|inveniatur manus tua omnibus inimicis tuis dextera tua inveniat %omnes; qui te oderunt
PS|20|10|pones eos ut clibanum ignis in tempore vultus tui Dominus in ira sua conturbabit eos et devorabit eos ignis
PS|20|11|fructum eorum de terra perdes et semen eorum a filiis hominum
PS|20|12|quoniam declinaverunt in te mala cogitaverunt consilia quae non potuerunt %stabilire;
PS|20|13|quoniam pones eos dorsum in reliquis tuis praeparabis vultum eorum
PS|20|14|exaltare Domine in virtute tua cantabimus et psallemus virtutes tuas
PS|21|1|in finem pro adsumptione matutina psalmus David
PS|21|2|Deus Deus meus respice me; quare me dereliquisti longe a salute mea verba delictorum meorum
PS|21|3|Deus meus clamabo per diem et non exaudies et nocte et non ad insipientiam mihi
PS|21|4|tu autem in sancto habitas Laus Israhel
PS|21|5|in te speraverunt patres nostri speraverunt et liberasti eos
PS|21|6|ad te clamaverunt et salvi facti sunt in te speraverunt et non sunt confusi
PS|21|7|ego autem sum vermis et non homo obprobrium hominum et abiectio plebis
PS|21|8|omnes videntes me deriserunt me locuti sunt labiis moverunt caput
PS|21|9|speravit in Domino eripiat eum salvum faciat eum quoniam vult eum
PS|21|10|quoniam tu es qui extraxisti me de ventre spes mea ab uberibus matris meae
PS|21|11|in te proiectus sum ex utero de ventre matris meae Deus meus es tu
PS|21|12|ne discesseris a me quoniam tribulatio proxima est quoniam non est qui adiuvet
PS|21|13|circumdederunt me vituli multi tauri pingues obsederunt me
PS|21|14|aperuerunt super me os suum sicut leo rapiens et rugiens
PS|21|15|sicut aqua effusus sum et dispersa sunt universa ossa mea factum est cor meum tamquam cera liquescens in medio ventris mei
PS|21|16|aruit tamquam testa virtus mea et lingua mea adhesit faucibus meis et in limum mortis deduxisti me
PS|21|17|quoniam circumdederunt me canes multi concilium malignantium obsedit me foderunt manus meas et pedes meos
PS|21|18|dinumeraverunt omnia ossa mea ipsi vero consideraverunt et inspexerunt me
PS|21|19|diviserunt sibi vestimenta mea et super vestem meam miserunt sortem
PS|21|20|tu autem Domine ne elongaveris auxilium tuum ad defensionem meam conspice
PS|21|21|erue a framea animam meam et de manu canis unicam meam
PS|21|22|salva me ex ore leonis et a cornibus unicornium humilitatem meam
PS|21|23|narrabo nomen tuum fratribus meis in media ecclesia laudabo te
PS|21|24|qui timetis Dominum laudate eum universum semen Iacob magnificate eum
PS|21|25|timeat eum omne semen Israhel quoniam non sprevit neque dispexit deprecationem pauperis nec avertit faciem suam a me et cum clamarem ad eum exaudivit %me;
PS|21|26|apud te laus mea in ecclesia magna vota mea reddam in conspectu timentium eum
PS|21|27|edent pauperes et saturabuntur et laudabunt Dominum qui requirunt eum vivent corda eorum in saeculum saeculi
PS|21|28|reminiscentur et convertentur ad Dominum universi fines terrae et adorabunt in conspectu eius universae familiae gentium
PS|21|29|quoniam Dei est regnum et %ipse; dominabitur gentium
PS|21|30|manducaverunt et adoraverunt omnes pingues terrae in conspectu eius cadent omnes qui descendunt in terram
PS|21|31|et anima mea illi vivet et semen meum serviet ipsi
PS|21|32|adnuntiabitur Domino generatio ventura et adnuntiabunt iustitiam eius populo qui nascetur quem fecit %Dominus;
PS|22|1|psalmus David Dominus reget me et nihil mihi deerit
PS|22|2|in loco pascuae %ibi; me conlocavit super aquam refectionis educavit me
PS|22|3|animam meam convertit deduxit me super semitas iustitiae propter nomen suum
PS|22|4|nam et si ambulavero in medio umbrae mortis non timebo mala quoniam tu mecum es virga tua et baculus tuus ipsa me consolata sunt
PS|22|5|parasti in conspectu meo mensam adversus eos qui tribulant me inpinguasti in oleo caput meum et calix meus inebrians quam praeclarus est
PS|22|6|et misericordia tua subsequitur me omnibus diebus vitae meae et ut inhabitem in domo Domini in longitudinem dierum
PS|23|1|psalmus David prima sabbati Domini est terra et plenitudo eius orbis terrarum et %universi; qui habitant in eo
PS|23|2|quia; ipse super maria fundavit eum et super flumina praeparavit eum
PS|23|3|quis ascendit in montem Domini aut quis stabit in loco sancto eius
PS|23|4|innocens manibus et mundo corde qui non accepit in vano animam suam nec iuravit in dolo proximo suo
PS|23|5|hic accipiet benedictionem a Domino et misericordiam a Deo salvatore suo
PS|23|6|haec est generatio quaerentium eum quaerentium faciem Dei Iacob diapsalma
PS|23|7|adtollite portas principes vestras et elevamini portae aeternales et introibit rex gloriae
PS|23|8|quis est iste rex gloriae Dominus fortis et potens Dominus potens in proelio
PS|23|9|adtollite portas principes vestras et elevamini portae aeternales et introibit rex gloriae
PS|23|10|quis est iste rex gloriae Dominus virtutum ipse est rex gloriae diapsalma
PS|24|1|psalmus David ad te Domine levavi animam meam
PS|24|2|Deus meus in te confido non erubescam
PS|24|3|neque inrideant me inimici mei etenim universi qui sustinent te non confundentur
PS|24|4|confundantur %omnes; iniqua agentes supervacue vias tuas Domine demonstra mihi %et; semitas tuas doce me
PS|24|5|dirige me in veritatem tuam et doce me quoniam tu es Deus salvator meus et te sustinui tota die
PS|24|6|reminiscere miserationum tuarum Domine et misericordiarum tuarum quia a saeculo sunt
PS|24|7|delicta iuventutis meae et ignorantias meas ne memineris secundum misericordiam tuam memento mei tu; propter bonitatem tuam Domine
PS|24|8|dulcis et rectus Dominus propter hoc legem dabit delinquentibus in via
PS|24|9|diriget mansuetos in iudicio docebit mites vias suas
PS|24|10|universae viae Domini misericordia et veritas requirentibus testamentum eius et testimonia eius
PS|24|11|propter nomen tuum Domine et propitiaberis peccato meo multum est enim
PS|24|12|quis est homo qui timet Dominum legem statuet ei in via quam elegit
PS|24|13|anima eius in bonis demorabitur et semen ipsius hereditabit terram
PS|24|14|firmamentum est Dominus timentibus eum et testamentum ipsius ut manifestetur illis
PS|24|15|oculi mei semper ad Dominum quoniam ipse evellet de laqueo pedes meos
PS|24|16|respice in me et miserere mei quia unicus et pauper sum ego
PS|24|17|tribulationes cordis mei multiplicatae sunt de necessitatibus meis erue me
PS|24|18|vide humilitatem meam et laborem meum et dimitte universa delicta mea
PS|24|19|respice inimicos meos quoniam multiplicati sunt et odio iniquo oderunt me
PS|24|20|custodi animam meam et erue me non erubescam quoniam speravi in te
PS|24|21|innocentes et recti adheserunt mihi quia sustinui te
PS|24|22|libera Deus Israhel ex omnibus tribulationibus suis
PS|25|1|psalmus David iudica me Domine quoniam ego in innocentia mea ingressus sum et in Domino sperans non infirmabor
PS|25|2|proba me Domine et tempta me ure renes meos et cor meum
PS|25|3|quoniam misericordia tua ante oculos meos est et conplacui in veritate tua
PS|25|4|non sedi cum concilio vanitatis et cum iniqua gerentibus non introibo
PS|25|5|odivi ecclesiam malignantium et cum impiis non sedebo
PS|25|6|lavabo inter innocentes manus meas et circumdabo altare tuum Domine
PS|25|7|ut audiam vocem laudis et enarrem universa mirabilia tua
PS|25|8|Domine dilexi decorem domus tuae et locum habitationis gloriae tuae
PS|25|9|ne perdas cum impiis animam meam et cum viris sanguinum vitam meam
PS|25|10|in quorum manibus iniquitates sunt dextera eorum repleta est muneribus
PS|25|11|ego autem in innocentia mea ingressus sum redime me et miserere mei
PS|25|12|pes meus stetit in directo in ecclesiis benedicam %te; Domine
PS|26|1|David priusquam liniretur Dominus inluminatio mea et salus mea quem timebo Dominus protector vitae meae a quo trepidabo
PS|26|2|dum adpropiant super me nocentes ut edant carnes meas qui tribulant me et inimici mei ipsi infirmati sunt et ceciderunt
PS|26|3|si consistant adversus me castra non timebit cor meum si exsurgat adversus me proelium in hoc ego sperabo
PS|26|4|unam petii a Domino hanc requiram ut inhabitem in domo Domini omnes dies vitae meae ut videam voluntatem Domini et visitem templum eius
PS|26|5|quoniam abscondit me in tabernaculo in die malorum protexit me in abscondito tabernaculi sui
PS|26|6|in petra exaltavit me et nunc exaltavit caput meum super inimicos meos circuivi et immolavi in tabernaculo eius hostiam vociferationis cantabo et psalmum dicam Domino
PS|26|7|exaudi Domine vocem meam qua clamavi miserere mei et exaudi me
PS|26|8|tibi dixit cor meum exquisivit facies mea faciem tuam Domine requiram
PS|26|9|ne avertas faciem tuam a me ne declines in ira a servo tuo adiutor meus esto ne derelinquas me neque dispicias me Deus salvator meus
PS|26|10|quoniam pater meus et mater mea dereliquerunt me Dominus autem adsumpsit me
PS|26|11|legem pone mihi Domine in via tua et dirige me in semita recta propter inimicos meos
PS|26|12|ne tradideris me in animas tribulantium me quoniam insurrexerunt in me testes iniqui et mentita est iniquitas sibi
PS|26|13|credo videre bona Domini in terra viventium
PS|26|14|expecta Dominum viriliter age et confortetur cor tuum et sustine Dominum
PS|27|1|huic David ad te Domine clamabo Deus meus ne sileas a me nequando taceas a me et adsimilabor descendentibus in lacum
PS|27|2|exaudi vocem deprecationis meae dum oro ad te dum extollo manus meas ad templum sanctum tuum
PS|27|3|ne simul tradas me cum peccatoribus et cum operantibus iniquitatem %ne perdideris me; qui loquuntur pacem cum proximo suo mala autem sunt in cordibus eorum
PS|27|4|da illis secundum opera ipsorum et secundum nequitiam adinventionum ipsorum secundum opera manuum eorum tribue illis redde retributionem eorum ipsis
PS|27|5|quoniam non intellexerunt opera Domini et in opera manuum eius destrues illos et non aedificabis eos
PS|27|6|benedictus Dominus quoniam exaudivit vocem deprecationis meae
PS|27|7|Dominus adiutor meus et protector meus in ipso speravit cor meum et adiutus sum et refloruit caro mea et ex voluntate mea confitebor ei
PS|27|8|Dominus fortitudo plebis suae et protector salvationum christi sui est
PS|27|9|salvam fac plebem tuam et benedic hereditati tuae et rege eos et extolle eos usque in aeternum
PS|28|1|psalmus David in consummatione tabernaculi adferte Domino filii Dei adferte Domino filios arietum
PS|28|2|adferte Domino gloriam et honorem adferte Domino gloriam nomini eius adorate Dominum in atrio sancto eius
PS|28|3|vox Domini super aquas Deus maiestatis intonuit Dominus super aquas multas
PS|28|4|vox Domini in virtute vox Domini in magnificentia
PS|28|5|vox Domini confringentis cedros et confringet Dominus cedros Libani
PS|28|6|et comminuet eas tamquam vitulum Libani et dilectus quemadmodum filius unicornium
PS|28|7|vox Domini intercidentis flammam ignis
PS|28|8|vox Domini concutientis desertum et commovebit Dominus desertum Cades
PS|28|9|vox Domini praeparantis cervos et revelabit condensa et in templo eius omnis dicet gloriam
PS|28|10|Dominus diluvium inhabitare facit et sedebit Dominus rex in aeternum
PS|28|11|Dominus virtutem populo suo dabit Dominus benedicet populo suo in pace
PS|29|1|psalmus cantici in dedicatione domus David
PS|29|2|exaltabo te Domine quoniam suscepisti me nec delectasti inimicos meos super me
PS|29|3|Domine Deus meus clamavi ad te et sanasti me
PS|29|4|Domine eduxisti ab inferno animam meam salvasti me a descendentibus in lacum
PS|29|5|psallite Domino sancti eius et confitemini memoriae sanctitatis eius
PS|29|6|quoniam ira in indignatione eius et vita in voluntate eius ad vesperum demorabitur fletus et ad matutinum laetitia
PS|29|7|ego autem dixi in abundantia mea non movebor in aeternum
PS|29|8|Domine in voluntate tua praestitisti decori meo virtutem avertisti faciem tuam et factus sum conturbatus
PS|29|9|ad te Domine clamabo et ad Deum meum deprecabor
PS|29|10|quae utilitas in sanguine meo dum descendo in corruptionem numquid confitebitur tibi pulvis aut adnuntiabit veritatem tuam
PS|29|11|audivit Dominus et misertus est mei Dominus factus est adiutor meus
PS|29|12|convertisti planctum meum in gaudium mihi conscidisti saccum meum et circumdedisti me laetitia
PS|29|13|ut cantet tibi gloria mea et non conpungar Domine Deus meus in aeternum confitebor tibi
PS|30|1|in finem psalmus David
PS|30|2|in te Domine speravi non confundar in aeternum in iustitia tua libera me
PS|30|3|inclina ad me aurem tuam adcelera ut eruas me esto mihi in Deum protectorem et in domum refugii ut salvum me facias
PS|30|4|quoniam fortitudo mea et refugium meum es tu et propter nomen tuum deduces me et enutries me
PS|30|5|educes me de laqueo hoc quem absconderunt mihi quoniam tu es protector meus
PS|30|6|in manus tuas commendabo spiritum meum redemisti me Domine Deus veritatis
PS|30|7|odisti observantes vanitates supervacue ego autem in Domino speravi
PS|30|8|exultabo et laetabor in misericordia tua quoniam respexisti humilitatem meam salvasti de necessitatibus animam meam
PS|30|9|nec conclusisti me in manibus inimici statuisti in loco spatioso pedes meos
PS|30|10|miserere mei Domine quoniam tribulor conturbatus est in ira oculus meus anima mea et venter meus
PS|30|11|quoniam defecit in dolore vita mea et anni mei in gemitibus infirmata est in paupertate virtus mea et ossa mea conturbata sunt
PS|30|12|super omnes inimicos meos factus sum obprobrium et vicinis meis valde et timor notis meis qui videbant me foras fugerunt a me
PS|30|13|oblivioni datus sum tamquam mortuus a corde factus sum tamquam vas perditum
PS|30|14|quoniam audivi vituperationem multorum commorantium in circuitu in eo dum convenirent simul adversus me accipere animam meam consiliati sunt
PS|30|15|ego autem in te speravi Domine dixi Deus meus es tu
PS|30|16|in manibus tuis sortes meae eripe me de manu inimicorum meorum et a persequentibus me
PS|30|17|inlustra faciem tuam super servum tuum salvum me fac in misericordia tua
PS|30|18|Domine ne confundar quoniam invocavi te erubescant impii et deducantur in infernum
PS|30|19|muta fiant labia dolosa quae loquuntur adversus iustum iniquitatem in superbia et in abusione
PS|30|20|quam magna multitudo dulcedinis tuae %Domine; quam abscondisti timentibus te perfecisti eis qui sperant in te in conspectu filiorum hominum
PS|30|21|abscondes eos in abdito faciei tuae a conturbatione hominum proteges eos in tabernaculo a contradictione linguarum
PS|30|22|benedictus Dominus quoniam mirificavit misericordiam suam mihi in civitate munita
PS|30|23|ego autem dixi in excessu mentis meae proiectus sum a facie oculorum tuorum ideo exaudisti vocem orationis meae dum clamarem ad te
PS|30|24|diligite Dominum omnes sancti eius %quoniam; veritates requirit Dominus et retribuit abundanter facientibus superbiam
PS|30|25|viriliter agite et confortetur cor vestrum omnes qui speratis in Domino
PS|31|1|huic David intellectus beati quorum remissae sunt iniquitates et quorum tecta sunt peccata
PS|31|2|beatus vir cui non inputabit Dominus peccatum nec est in spiritu eius dolus
PS|31|3|quoniam tacui inveteraverunt ossa mea dum clamarem tota die
PS|31|4|quoniam die ac nocte gravata est super me manus tua conversus sum in aerumna mea; dum configitur %mihi; spina diapsalma
PS|31|5|delictum meum cognitum tibi; feci et iniustitiam meam non abscondi dixi confitebor adversus me iniustitiam meam Domino et tu remisisti impietatem peccati mei diapsalma
PS|31|6|pro hac orabit ad te omnis sanctus in tempore oportuno verumtamen in diluvio aquarum multarum ad eum non adproximabunt
PS|31|7|tu es refugium meum a tribulatione quae circumdedit me exultatio mea erue me a circumdantibus me diapsalma
PS|31|8|intellectum tibi dabo et instruam te in via hac qua gradieris firmabo super te oculos meos
PS|31|9|nolite fieri sicut equus et mulus quibus non est intellectus in camo et freno maxillas eorum constringe qui non adproximant ad te
PS|31|10|multa flagella peccatoris sperantem autem in Domino misericordia circumdabit
PS|31|11|laetamini in Domino et exultate iusti et gloriamini omnes recti corde
PS|32|1|psalmus David exultate iusti in Domino rectos decet laudatio
PS|32|2|confitemini Domino in cithara in psalterio decem cordarum psallite illi
PS|32|3|cantate ei canticum novum bene psallite in vociferatione
PS|32|4|quia rectum est verbum Domini et omnia opera eius in fide
PS|32|5|diligit misericordiam et iudicium misericordia Domini plena est terra
PS|32|6|verbo Domini caeli firmati sunt et spiritu oris eius omnis virtus eorum
PS|32|7|congregans sicut in utre aquas maris ponens in thesauris abyssos
PS|32|8|timeat Dominum omnis terra ab eo autem commoveantur omnes inhabitantes orbem
PS|32|9|quoniam ipse dixit et facta sunt ipse mandavit et creata sunt
PS|32|10|Dominus dissipat consilia gentium reprobat autem cogitationes populorum %et reprobat consilia principum;
PS|32|11|consilium autem Domini in aeternum manet cogitationes cordis eius in generatione et generationem
PS|32|12|beata gens cuius est Dominus Deus eius populus quem elegit in hereditatem sibi
PS|32|13|de caelo respexit Dominus vidit omnes filios hominum
PS|32|14|de praeparato habitaculo suo respexit super omnes qui habitant terram
PS|32|15|qui finxit singillatim corda eorum qui intellegit omnia opera illorum
PS|32|16|non salvatur rex per multam virtutem et gigans non salvabitur in multitudine virtutis suae
PS|32|17|fallax equus ad salutem in abundantia autem virtutis suae non salvabitur
PS|32|18|ecce oculi Domini super metuentes eum qui sperant super misericordia eius
PS|32|19|ut eruat a morte animas eorum et alat eos in fame
PS|32|20|anima nostra sustinet Dominum quoniam adiutor et protector noster est
PS|32|21|quia in eo laetabitur cor nostrum et in nomine sancto eius speravimus
PS|32|22|fiat misericordia tua Domine super nos quemadmodum speravimus in te
PS|33|1|David cum inmutavit vultum suum coram Abimelech et dimisit eum et abiit
PS|33|2|benedicam Dominum in omni tempore semper laus eius in ore meo
PS|33|3|in Domino laudabitur anima mea audiant mansueti et laetentur
PS|33|4|magnificate Dominum mecum et exaltemus nomen eius in id ipsum
PS|33|5|exquisivi Dominum et exaudivit me et ex omnibus tribulationibus meis eripuit me
PS|33|6|accedite ad eum et inluminamini et facies vestrae non confundentur
PS|33|7|iste pauper clamavit et Dominus exaudivit %eum; et de omnibus tribulationibus eius salvavit eum
PS|33|8|vallabit angelus Domini in circuitu timentium eum et eripiet eos
PS|33|9|gustate et videte quoniam suavis est Dominus beatus vir qui sperat in eo
PS|33|10|timete Dominum %omnes; sancti eius quoniam non est inopia timentibus eum
PS|33|11|divites eguerunt et esurierunt inquirentes autem Dominum non minuentur omni bono diapsalma
PS|33|12|venite filii audite me timorem Domini docebo vos
PS|33|13|quis est homo qui vult vitam cupit videre dies bonos
PS|33|14|prohibe linguam tuam a malo et labia tua ne loquantur dolum
PS|33|15|deverte a malo et fac bonum inquire pacem et persequere eam
PS|33|16|oculi Domini super iustos et aures eius in precem eorum
PS|33|17|facies Domini super facientes mala ut perdat de terra memoriam eorum
PS|33|18|clamaverunt iusti et Dominus exaudivit et ex omnibus tribulationibus eorum liberavit eos
PS|33|19|iuxta est Dominus his qui tribulato sunt corde et humiles spiritu salvabit
PS|33|20|multae tribulationes iustorum et de omnibus his liberavit eos
PS|33|21|Dominus custodit omnia ossa eorum unum ex his non conteretur
PS|33|22|mors peccatorum pessima et qui oderunt iustum delinquent
PS|33|23|redimet Dominus animas servorum suorum et non delinquent omnes qui sperant in eum
PS|34|1|huic David iudica Domine nocentes me expugna expugnantes me
PS|34|2|adprehende arma et scutum et exsurge in adiutorium mihi
PS|34|3|effunde frameam et conclude adversus eos qui persequuntur me dic animae meae salus tua ego sum
PS|34|4|confundantur et revereantur quaerentes animam meam avertantur retrorsum et confundantur cogitantes mihi mala
PS|34|5|fiant tamquam pulvis ante faciem venti et angelus Domini coartans eos
PS|34|6|fiat via illorum tenebrae et lubricum et angelus Domini persequens eos
PS|34|7|quoniam gratis absconderunt mihi interitum laquei sui supervacue exprobraverunt animam meam
PS|34|8|veniat illi laqueus quem ignorat et captio quam abscondit conprehendat eum et in laqueo cadat in ipso
PS|34|9|anima autem mea exultabit in Domino delectabitur super salutari suo
PS|34|10|omnia ossa mea dicent Domine quis similis tui eripiens inopem de manu fortiorum eius egenum et pauperem a diripientibus eum
PS|34|11|surgentes testes iniqui quae ignorabam interrogabant me
PS|34|12|retribuebant mihi mala pro bonis sterilitatem animae meae
PS|34|13|ego autem cum mihi molesti essent induebar cilicio humiliabam in ieiunio animam meam et oratio mea in sinum meum convertetur
PS|34|14|quasi proximum quasi fratrem nostrum sic conplacebam quasi lugens et contristatus sic humiliabar
PS|34|15|et adversum me laetati sunt et convenerunt congregata sunt super me flagella et ignoravi
PS|34|16|dissipati sunt nec conpuncti temptaverunt me subsannaverunt me subsannatione frenduerunt super me dentibus suis
PS|34|17|Domine quando respicies restitue animam meam a malignitate eorum a leonibus unicam meam
PS|34|18|confitebor tibi in ecclesia magna in populo gravi laudabo te
PS|34|19|non supergaudeant mihi qui adversantur mihi inique qui oderunt me gratis et annuunt oculis
PS|34|20|quoniam mihi quidem pacifice loquebantur et in iracundia terrae loquentes; dolos cogitabant
PS|34|21|et dilataverunt super me os suum dixerunt euge euge viderunt oculi nostri
PS|34|22|vidisti Domine ne sileas Domine ne discedas a me
PS|34|23|exsurge et intende iudicio meo Deus meus et Dominus meus in causam meam
PS|34|24|iudica me secundum iustitiam tuam Domine Deus meus et non supergaudeant mihi
PS|34|25|non dicant in cordibus suis euge euge animae nostrae nec dicant devoravimus eum
PS|34|26|erubescant et revereantur simul qui gratulantur malis meis induantur confusione et reverentia qui magna loquuntur super me
PS|34|27|exultent et laetentur qui volunt iustitiam meam et dicant semper magnificetur Dominus qui volunt pacem servi eius
PS|34|28|et lingua mea meditabitur iustitiam tuam tota die laudem tuam
PS|35|1|in finem servo Domini David
PS|35|2|dixit iniustus ut delinquat in semet ipso non est timor Dei ante oculos eius
PS|35|3|quoniam dolose egit in conspectu eius ut inveniatur iniquitas eius ad odium
PS|35|4|verba oris eius iniquitas et dolus noluit intellegere ut bene ageret
PS|35|5|iniquitatem meditatus est in cubili suo adstetit omni viae non bonae malitiam autem non odivit
PS|35|6|Domine in caelo misericordia tua et veritas tua usque ad nubes
PS|35|7|iustitia tua sicut montes Dei iudicia tua abyssus multa homines et iumenta salvabis Domine
PS|35|8|quemadmodum multiplicasti misericordiam tuam Deus filii autem hominum in tegmine alarum tuarum sperabunt
PS|35|9|inebriabuntur ab ubertate domus tuae et torrente voluntatis tuae potabis eos
PS|35|10|quoniam apud te fons vitae in lumine tuo videbimus lumen
PS|35|11|praetende misericordiam tuam scientibus te et iustitiam tuam his qui recto sunt corde
PS|35|12|non veniat mihi pes superbiae et manus peccatoris non moveat me
PS|35|13|ibi ceciderunt qui operantur iniquitatem expulsi sunt nec potuerunt stare
PS|36|1|ipsi David noli aemulari in malignantibus neque zelaveris facientes iniquitatem
PS|36|2|quoniam tamquam faenum velociter arescent et quemadmodum holera herbarum cito decident
PS|36|3|spera in Domino et fac bonitatem et inhabita terram et pasceris in divitiis eius
PS|36|4|delectare in Domino et dabit tibi petitiones cordis tui
PS|36|5|revela Domino viam tuam et spera in eum et ipse faciet
PS|36|6|et educet quasi lumen iustitiam tuam et iudicium tuum tamquam meridiem
PS|36|7|subditus esto Domino et ora eum noli aemulari in eo qui prosperatur in via sua in homine faciente iniustitias
PS|36|8|desine ab ira et derelinque furorem noli aemulari ut maligneris
PS|36|9|quoniam qui malignantur exterminabuntur sustinentes autem Dominum ipsi hereditabunt terram
PS|36|10|et adhuc pusillum et non erit peccator et quaeres locum eius et non invenies
PS|36|11|mansueti autem hereditabunt terram et delectabuntur in multitudine pacis
PS|36|12|observabit peccator iustum et stridebit super eum dentibus suis
PS|36|13|Dominus autem inridebit eum quia prospicit quoniam veniet dies eius
PS|36|14|gladium evaginaverunt peccatores intenderunt arcum suum ut decipiant pauperem et inopem ut trucident rectos corde
PS|36|15|gladius eorum intret in corda ipsorum et arcus ipsorum confringatur
PS|36|16|melius est modicum iusto super divitias peccatorum multas
PS|36|17|quoniam brachia peccatorum conterentur confirmat autem iustos Dominus
PS|36|18|novit Dominus dies inmaculatorum et hereditas eorum in aeternum erit
PS|36|19|non confundentur in tempore malo et in diebus famis saturabuntur
PS|36|20|quia peccatores peribunt inimici vero Domini mox honorificati fuerint et exaltati deficientes quemadmodum fumus defecerunt
PS|36|21|mutuabitur peccator et non solvet iustus autem miseretur et tribuet
PS|36|22|quia benedicentes ei hereditabunt terram maledicentes autem ei disperibunt
PS|36|23|apud Dominum gressus hominis dirigentur et viam eius volet
PS|36|24|cum ceciderit non conlidetur quia Dominus subponit manum suam
PS|36|25|iunior fui et senui et non vidi iustum derelictum nec semen eius quaerens panes
PS|36|26|tota die miseretur et commodat et semen illius in benedictione erit
PS|36|27|declina a malo et fac bonum et inhabita in saeculum saeculi
PS|36|28|quia Dominus amat iudicium et non derelinquet sanctos suos in aeternum conservabuntur iniusti punientur et semen impiorum peribit
PS|36|29|iusti autem hereditabunt terram et inhabitabunt in saeculum %saeculi; super eam
PS|36|30|os iusti meditabitur sapientiam et lingua eius loquetur iudicium
PS|36|31|lex Dei eius in corde ipsius et non subplantabuntur gressus eius
PS|36|32|considerat peccator iustum et quaerit mortificare eum
PS|36|33|Dominus autem non derelinquet eum in manus eius nec damnabit eum cum iudicabitur illi
PS|36|34|expecta Dominum et custodi viam eius et exaltabit te ut hereditate capias terram cum perierint peccatores videbis
PS|36|35|vidi impium superexaltatum et elevatum sicut cedros Libani
PS|36|36|et transivi et ecce non erat et quaesivi eum et non est inventus locus eius
PS|36|37|custodi innocentiam et vide aequitatem quoniam sunt reliquiae homini pacifico
PS|36|38|iniusti autem disperibunt simul reliquiae impiorum peribunt
PS|36|39|salus autem iustorum a Domino et protector eorum in tempore tribulationis
PS|36|40|et adiuvabit eos Dominus et liberabit eos et eruet eos a peccatoribus et salvabit eos quia speraverunt in eo
PS|37|1|psalmus David in rememorationem de sabbato
PS|37|2|Domine ne in furore tuo arguas me neque in ira tua corripias me
PS|37|3|quoniam sagittae tuae infixae sunt mihi et confirmasti super me manum tuam
PS|37|4|non est sanitas carni meae a facie irae tuae non est pax ossibus meis a facie peccatorum meorum
PS|37|5|quoniam iniquitates meae supergressae sunt caput meum sicut onus grave gravatae sunt super me
PS|37|6|putruerunt et corruptae sunt cicatrices meae a facie insipientiae meae
PS|37|7|miser factus sum et curvatus sum usque ad finem tota die contristatus ingrediebar
PS|37|8|quoniam lumbi mei impleti sunt inlusionibus et non est sanitas in carne mea
PS|37|9|adflictus sum et humiliatus sum nimis rugiebam a gemitu cordis mei
PS|37|10|Domine ante te omne desiderium meum et gemitus meus a te non est absconditus
PS|37|11|cor meum conturbatum est dereliquit me virtus mea et lumen oculorum meorum et ipsum non est mecum
PS|37|12|amici mei et proximi mei adversus me adpropinquaverunt et steterunt et qui iuxta me erant de longe steterunt
PS|37|13|et vim faciebant qui quaerebant animam meam et qui inquirebant mala mihi locuti sunt vanitates et dolos tota die meditabantur
PS|37|14|ego autem tamquam surdus non audiebam et sicut mutus non aperiens os suum
PS|37|15|et factus sum sicut homo non audiens et non habens in ore suo redargutiones
PS|37|16|quoniam in te Domine speravi tu exaudies Domine Deus meus
PS|37|17|quia dixi nequando supergaudeant mihi inimici mei et dum commoventur pedes mei super me magna locuti sunt
PS|37|18|quoniam ego in flagella paratus et dolor meus in conspectu meo semper
PS|37|19|quoniam iniquitatem meam adnuntiabo %et; cogitabo pro peccato meo
PS|37|20|inimici autem mei vivent et firmati sunt super me et multiplicati sunt qui oderunt me inique
PS|37|21|qui retribuunt mala pro bonis detrahebant mihi quoniam sequebar bonitatem
PS|37|22|non derelinquas me Domine Deus meus ne discesseris a me
PS|37|23|intende in adiutorium meum Domine salutis meae
PS|38|1|in finem Idithun canticum David
PS|38|2|dixi custodiam vias meas ut non delinquam in lingua mea posui ori meo custodiam cum consisteret peccator adversum me
PS|38|3|obmutui et humiliatus sum et silui a bonis et dolor meus renovatus est
PS|38|4|concaluit cor meum intra me et in meditatione mea exardescet ignis
PS|38|5|locutus sum in lingua mea notum fac mihi Domine finem meum et numerum dierum meorum quis est ut sciam quid desit mihi
PS|38|6|ecce mensurabiles posuisti dies meos et substantia mea tamquam nihilum ante te verumtamen universa vanitas omnis homo vivens diapsalma
PS|38|7|verumtamen in imagine pertransit homo sed et frustra conturbatur thesaurizat et ignorat cui congregabit ea
PS|38|8|et nunc quae est expectatio mea nonne Dominus et substantia mea apud te est
PS|38|9|ab omnibus iniquitatibus meis erue me obprobrium insipienti dedisti me
PS|38|10|obmutui %et; non aperui os meum quoniam tu fecisti
PS|38|11|amove a me plagas tuas
PS|38|12|a fortitudine manus tuae ego defeci in increpationibus propter iniquitatem corripuisti hominem et tabescere fecisti sicut araneam animam eius verumtamen vane %conturbatur; omnis homo diapsalma
PS|38|13|exaudi orationem meam Domine et deprecationem meam auribus percipe lacrimas meas ne sileas quoniam advena sum apud te et peregrinus sicut omnes patres mei
PS|38|14|remitte mihi ut refrigerer priusquam abeam et amplius non ero
PS|39|1|in finem David psalmus
PS|39|2|expectans expectavi Dominum et intendit mihi
PS|39|3|et exaudivit preces meas et eduxit me de lacu miseriae et de luto fecis et statuit super petram pedes meos et direxit gressus meos
PS|39|4|et inmisit in os meum canticum novum carmen Deo nostro videbunt multi et timebunt et sperabunt in Domino
PS|39|5|beatus vir cuius est nomen Domini spes ipsius et non respexit in vanitates et insanias falsas
PS|39|6|multa fecisti tu Domine Deus meus mirabilia tua et cogitationibus tuis non est qui similis sit tibi adnuntiavi et locutus sum multiplicati sunt super numerum
PS|39|7|sacrificium et oblationem noluisti aures autem perfecisti mihi holocaustum et pro peccato non postulasti
PS|39|8|tunc dixi ecce venio in capite libri scriptum est de me
PS|39|9|ut facerem voluntatem tuam Deus meus volui et legem tuam in medio cordis mei
PS|39|10|adnuntiavi iustitiam in ecclesia magna ecce labia mea non prohibebo Domine tu scisti
PS|39|11|iustitiam tuam non abscondi in corde meo veritatem tuam et salutare tuum dixi non abscondi misericordiam tuam et veritatem tuam a concilio multo
PS|39|12|tu autem Domine ne longe facias miserationes tuas a me misericordia tua et veritas tua semper susceperunt me
PS|39|13|quoniam circumdederunt me mala quorum non est numerus conprehenderunt me iniquitates meae et non potui ut viderem multiplicatae sunt super capillos capitis mei et cor meum dereliquit me
PS|39|14|conplaceat tibi Domine ut eruas me Domine ad adiuvandum me respice
PS|39|15|confundantur et revereantur simul qui quaerunt animam meam ut auferant eam convertantur retrorsum et revereantur qui volunt mihi mala
PS|39|16|ferant confestim confusionem suam qui dicunt mihi euge euge
PS|39|17|exultent et laetentur super te omnes quaerentes te et dicant semper magnificetur Dominus qui diligunt salutare tuum
PS|39|18|ego autem mendicus sum et pauper Dominus sollicitus est mei adiutor meus et protector meus tu es Deus meus ne tardaveris
PS|40|1|in finem psalmus David
PS|40|2|beatus qui intellegit super egenum et pauperem in die mala liberabit eum Dominus
PS|40|3|Dominus conservet eum et vivificet eum et beatum faciat eum in terra et non tradat eum in animam inimicorum eius
PS|40|4|Dominus opem ferat illi super lectum doloris eius universum stratum eius versasti in infirmitate eius
PS|40|5|ego dixi Domine miserere mei sana animam meam quoniam peccavi tibi
PS|40|6|inimici mei dixerunt mala mihi quando morietur et peribit nomen eius
PS|40|7|et si ingrediebatur ut videret vane loquebatur cor eius congregavit iniquitatem sibi egrediebatur foras et loquebatur
PS|40|8|in id ipsum adversum me susurrabant omnes inimici mei adversus me cogitabant mala mihi
PS|40|9|verbum iniquum constituerunt adversus me numquid qui dormit non adiciet ut resurgat
PS|40|10|etenim homo pacis meae in quo speravi qui edebat panes meos magnificavit super me subplantationem
PS|40|11|tu autem Domine miserere mei et resuscita me et retribuam eis
PS|40|12|in hoc cognovi quoniam voluisti me quoniam non gaudebit inimicus meus super me
PS|40|13|me autem propter innocentiam suscepisti et confirmasti me in conspectu tuo in aeternum
PS|40|14|benedictus Dominus Deus Israhel a saeculo et in saeculum fiat fiat
PS|41|1|in finem in intellectum filiis Core
PS|41|2|quemadmodum desiderat cervus ad fontes aquarum ita desiderat anima mea ad te Deus
PS|41|3|sitivit anima mea ad Deum fortem; vivum quando veniam et parebo ante faciem Dei
PS|41|4|fuerunt mihi lacrimae meae panis die ac nocte dum dicitur mihi cotidie ubi est Deus tuus
PS|41|5|haec recordatus sum et effudi in me animam meam quoniam transibo in loco tabernaculi admirabilis usque ad domum Dei in voce exultationis et confessionis sonus epulantis
PS|41|6|quare tristis es anima mea et quare conturbas me spera in Deo quoniam confitebor illi salutare vultus mei
PS|41|7|Deus meus ad me ipsum anima mea conturbata est propterea memor ero tui de terra Iordanis et Hermoniim a monte modico
PS|41|8|abyssus ad; abyssum invocat in voce cataractarum tuarum omnia excelsa tua et fluctus tui super me transierunt
PS|41|9|in die mandavit Dominus misericordiam suam et nocte canticum eius apud me oratio Deo vitae meae
PS|41|10|dicam Deo susceptor meus es quare oblitus es mei quare contristatus incedo dum adfligit me inimicus
PS|41|11|dum confringuntur ossa mea exprobraverunt mihi qui tribulant me dum dicunt mihi per singulos dies ubi est Deus tuus
PS|41|12|quare tristis es anima mea et quare conturbas me spera in Deum quoniam adhuc; confitebor illi salutare vultus mei et; Deus meus
PS|42|1|psalmus David iudica me Deus et discerne causam meam de gente non sancta ab homine iniquo et doloso erue me
PS|42|2|quia tu es Deus fortitudo mea quare me reppulisti quare tristis incedo dum adfligit me inimicus
PS|42|3|emitte lucem tuam et veritatem tuam ipsa me deduxerunt et adduxerunt in montem sanctum tuum et in tabernacula tua
PS|42|4|et introibo ad altare Dei ad Deum qui laetificat iuventutem meam confitebor tibi in cithara Deus Deus meus
PS|42|5|quare tristis es anima mea et quare conturbas me spera in Deum quoniam adhuc; confitebor illi salutare vultus mei et; Deus meus
PS|43|1|in finem filiis Core ad intellectum
PS|43|2|Deus auribus nostris audivimus patres nostri adnuntiaverunt nobis opus quod operatus es in diebus eorum in diebus antiquis
PS|43|3|manus tua gentes disperdit et plantasti eos adflixisti populos et expulisti eos
PS|43|4|nec enim in gladio suo possederunt terram et brachium eorum non salvavit eos sed dextera tua et brachium tuum et inluminatio faciei tuae quoniam conplacuisti in eis
PS|43|5|tu es ipse rex meus et Deus meus qui mandas salutes Iacob
PS|43|6|in te inimicos nostros ventilabimus cornu et in nomine tuo spernemus insurgentes in nobis
PS|43|7|non enim in arcu meo sperabo et gladius meus non salvabit me
PS|43|8|salvasti enim nos de adfligentibus nos et odientes nos confudisti
PS|43|9|in Deo laudabimur tota die et in nomine tuo confitebimur in saeculum diapsalma
PS|43|10|nunc autem reppulisti et confudisti nos et non egredieris in virtutibus nostris
PS|43|11|avertisti nos retrorsum post inimicos nostros et qui oderunt nos diripiebant sibi
PS|43|12|dedisti nos tamquam oves escarum et in gentibus dispersisti nos
PS|43|13|vendidisti populum tuum sine pretio et non fuit multitudo in commutationibus nostris
PS|43|14|posuisti nos obprobrium vicinis nostris subsannationem et derisum his qui in circuitu nostro
PS|43|15|posuisti nos in similitudinem gentibus commotionem capitis in populis
PS|43|16|tota die verecundia mea contra me est et confusio faciei meae cooperuit me
PS|43|17|a voce exprobrantis et obloquentis a facie inimici et persequentis
PS|43|18|haec omnia venerunt super nos nec obliti sumus te et inique non egimus in testamento tuo
PS|43|19|et non recessit retrorsum cor nostrum et declinasti semitas nostras a via tua
PS|43|20|quoniam humiliasti nos in loco adflictionis et cooperuit nos umbra mortis
PS|43|21|si obliti sumus nomen Dei nostri et %si; expandimus manus nostras ad deum alienum
PS|43|22|nonne Deus requiret ista ipse enim novit abscondita cordis quoniam propter te mortificamur omni die aestimati sumus sicut oves occisionis
PS|43|23|exsurge quare dormis Domine exsurge %et; ne repellas in finem
PS|43|24|quare faciem tuam avertis oblivisceris inopiae nostrae et tribulationis nostrae
PS|43|25|quoniam humiliata est in pulvere anima nostra conglutinatus est in terra venter noster
PS|43|26|exsurge adiuva nos et redime nos propter nomen tuum
PS|44|1|in finem pro his qui commutabuntur filiis Core ad intellectum canticum pro dilecto
PS|44|2|eructavit cor meum verbum bonum dico ego opera mea regi lingua mea calamus scribae velociter scribentis
PS|44|3|speciosus forma prae filiis hominum diffusa est gratia in labiis tuis propterea benedixit te Deus in aeternum
PS|44|4|accingere gladio tuo super femur tuum potentissime
PS|44|5|specie tua et pulchritudine tua et intende prospere procede et regna propter veritatem et mansuetudinem et iustitiam et deducet te mirabiliter dextera tua
PS|44|6|sagittae tuae acutae populi sub te cadent in corde inimicorum regis
PS|44|7|sedis tua Deus in saeculum saeculi virga directionis virga regni tui
PS|44|8|dilexisti iustitiam et odisti iniquitatem propterea unxit te Deus Deus tuus oleo laetitiae prae consortibus tuis
PS|44|9|murra et gutta et cassia a vestimentis tuis a domibus eburneis ex quibus delectaverunt te
PS|44|10|filiae regum in honore tuo adstetit regina a dextris tuis in vestitu deaurato circumdata varietate
PS|44|11|audi filia et vide et inclina aurem tuam et obliviscere populum tuum et domum patris tui
PS|44|12|et concupiscet rex decorem tuum quoniam ipse est dominus tuus et adorabunt eum
PS|44|13|et; filiae Tyri in muneribus vultum tuum deprecabuntur divites plebis
PS|44|14|omnis gloria eius filiae regis ab intus in fimbriis aureis
PS|44|15|circumamicta varietatibus adducentur regi virgines post eam proximae eius adferentur tibi
PS|44|16|adferentur in laetitia et exultatione adducentur in templum regis
PS|44|17|pro patribus tuis nati sunt tibi filii constitues eos principes super omnem terram
PS|44|18|memor ero nominis tui in omni generatione et generatione propterea populi confitebuntur tibi in aeternum et in saeculum saeculi
PS|45|1|in finem pro filiis Core pro arcanis psalmus
PS|45|2|Deus noster refugium et virtus adiutor in tribulationibus quae invenerunt nos nimis
PS|45|3|propterea non timebimus dum turbabitur terra et transferentur montes in cor maris
PS|45|4|sonaverunt et turbatae sunt aquae eorum conturbati sunt montes in fortitudine eius diapsalma
PS|45|5|fluminis impetus laetificat civitatem Dei sanctificavit tabernaculum suum Altissimus
PS|45|6|Deus in medio eius non commovebitur adiuvabit eam Deus mane diluculo
PS|45|7|conturbatae sunt gentes inclinata sunt regna dedit vocem suam mota est terra
PS|45|8|Dominus virtutum nobiscum susceptor noster Deus Iacob diapsalma
PS|45|9|venite et videte opera Domini quae posuit prodigia super terram
PS|45|10|auferens bella usque ad finem terrae arcum conteret et confringet arma et scuta conburet in igne
PS|45|11|vacate et videte quoniam ego sum Deus exaltabor in gentibus exaltabor in terra
PS|45|12|Dominus virtutum nobiscum susceptor noster Deus Iacob
PS|46|1|in finem pro filiis Core psalmus
PS|46|2|omnes gentes plaudite manibus iubilate Deo in voce exultationis
PS|46|3|quoniam Dominus excelsus terribilis rex magnus super omnem terram
PS|46|4|subiecit populos nobis et gentes sub pedibus nostris
PS|46|5|elegit nobis hereditatem suam speciem Iacob quam dilexit diapsalma
PS|46|6|ascendit Deus in iubilo Dominus in voce tubae
PS|46|7|psallite Deo nostro psallite psallite regi nostro psallite
PS|46|8|quoniam rex omnis terrae Deus psallite sapienter
PS|46|9|regnavit Deus super gentes Deus sedit super sedem sanctam suam
PS|46|10|principes populorum congregati sunt cum Deo Abraham quoniam Dei fortes terrae vehementer elevati sunt
PS|47|1|canticum psalmi filiis Core secunda sabbati
PS|47|2|magnus Dominus et laudabilis nimis in civitate Dei nostri in monte sancto eius
PS|47|3|fundatur exultatione universae terrae montes Sion latera aquilonis civitas regis magni
PS|47|4|Deus in domibus eius cognoscitur cum suscipiet eam
PS|47|5|quoniam ecce reges congregati sunt convenerunt in unum
PS|47|6|ipsi videntes sic admirati sunt conturbati sunt commoti sunt
PS|47|7|tremor adprehendit eos ibi dolores ut parturientis
PS|47|8|in spiritu vehementi conteres naves Tharsis
PS|47|9|sicut audivimus sic vidimus in civitate Domini virtutum in civitate Dei nostri Deus fundavit eam in aeternum diapsalma
PS|47|10|suscepimus Deus misericordiam tuam in medio templi tui
PS|47|11|secundum nomen tuum Deus sic et laus tua in fines terrae iustitia plena est dextera tua
PS|47|12|laetetur mons Sion exultent filiae Iudaeae propter iudicia tua %Domine;
PS|47|13|circumdate Sion et conplectimini eam narrate in turribus eius
PS|47|14|ponite corda vestra in virtute eius et distribuite domus eius ut enarretis in progeniem alteram
PS|47|15|quoniam hic est Deus Deus noster in aeternum et in saeculum saeculi ipse reget nos in saecula
PS|48|1|in finem filiis Core psalmus
PS|48|2|audite haec omnes gentes auribus percipite omnes qui habitatis orbem
PS|48|3|quique terriginae et filii hominum in unum dives et pauper
PS|48|4|os meum loquetur sapientiam et meditatio cordis mei prudentiam
PS|48|5|inclinabo in parabolam aurem meam aperiam in psalterio propositionem meam
PS|48|6|cur timebo in die malo iniquitas calcanei mei circumdabit me
PS|48|7|qui confidunt in virtute sua et in multitudine divitiarum suarum gloriantur
PS|48|8|frater non redimit redimet homo non dabit Deo placationem suam
PS|48|9|et pretium redemptionis animae suae et laboravit in aeternum
PS|48|10|et vivet adhuc; in finem
PS|48|11|non videbit interitum cum viderit sapientes morientes simul insipiens et stultus peribunt et relinquent alienis divitias suas
PS|48|12|%et; sepulchra eorum domus illorum in aeternum tabernacula eorum in progeniem et progeniem vocaverunt nomina sua in terris suis
PS|48|13|et homo cum in honore esset non intellexit conparatus est iumentis insipientibus et similis factus est illis
PS|48|14|haec via illorum scandalum ipsis et postea in ore suo conplacebunt diapsalma
PS|48|15|sicut oves in inferno positi sunt mors depascet eos et dominabuntur eorum iusti in matutino et auxilium eorum veterescet in inferno a gloria eorum
PS|48|16|verumtamen Deus redimet animam meam de manu inferi cum acceperit me diapsalma
PS|48|17|ne timueris cum dives factus fuerit homo et cum multiplicata fuerit gloria domus eius
PS|48|18|quoniam cum interierit non sumet omnia neque descendet cum eo pone; gloria eius
PS|48|19|quia anima eius in vita ipsius benedicetur confitebitur tibi cum benefeceris ei
PS|48|20|introibit usque in progenies patrum suorum usque in aeternum non videbit lumen
PS|48|21|homo in honore cum esset non intellexit conparatus est iumentis %insipientibus; et similis factus est illis
PS|49|1|psalmus Asaph Deus deorum Dominus locutus est et vocavit terram a solis ortu usque ad occasum
PS|49|2|ex Sion species decoris eius
PS|49|3|Deus manifeste veniet Deus noster et non silebit ignis in conspectu eius exardescet et in circuitu eius tempestas valida
PS|49|4|advocabit caelum desursum et terram discernere populum suum
PS|49|5|congregate illi sanctos eius qui ordinant testamentum eius super sacrificia
PS|49|6|et adnuntiabunt caeli iustitiam eius quoniam Deus iudex est diapsalma
PS|49|7|audi populus meus et loquar tibi Israhel et testificabor tibi Deus Deus tuus ego sum
PS|49|8|non in sacrificiis tuis arguam te holocausta autem tua in conspectu meo sunt semper
PS|49|9|non accipiam de domo tua vitulos neque de gregibus tuis hircos
PS|49|10|quoniam meae sunt omnes ferae silvarum iumenta in montibus et boves
PS|49|11|cognovi omnia volatilia caeli et pulchritudo agri mecum est
PS|49|12|si esuriero non dicam tibi meus est enim orbis terrae et plenitudo eius
PS|49|13|numquid manducabo carnes taurorum aut sanguinem hircorum potabo
PS|49|14|immola Deo sacrificium laudis et redde Altissimo vota tua
PS|49|15|et invoca me in die tribulationis et eruam te et honorificabis me diapsalma
PS|49|16|peccatori autem dixit Deus quare tu enarras iustitias meas et adsumis testamentum meum per os tuum
PS|49|17|tu vero odisti disciplinam et proiecisti sermones meos retrorsum
PS|49|18|si videbas furem currebas cum eo et cum adulteris portionem tuam ponebas
PS|49|19|os tuum abundavit malitia et lingua tua concinnabat dolos
PS|49|20|sedens adversus fratrem tuum loquebaris et adversus filium matris tuae ponebas scandalum
PS|49|21|haec fecisti et tacui existimasti inique quod ero tui similis arguam te et statuam contra faciem tuam
PS|49|22|intellegite nunc haec qui obliviscimini Deum nequando rapiat et non sit qui eripiat
PS|49|23|sacrificium laudis honorificabit me et illic iter quod ostendam illi salutare Dei
PS|50|1|in finem psalmus David
PS|50|2|cum venit ad eum Nathan propheta quando intravit ad Bethsabee
PS|50|3|miserere mei Deus secundum %magnam; misericordiam tuam %et; secundum multitudinem miserationum tuarum dele iniquitatem meam
PS|50|4|amplius lava me ab iniquitate mea et a peccato meo munda me
PS|50|5|quoniam iniquitatem meam ego cognosco et peccatum meum contra me est semper
PS|50|6|tibi soli peccavi et malum coram te feci ut iustificeris in sermonibus tuis et vincas cum iudicaris
PS|50|7|ecce enim in iniquitatibus conceptus sum et in peccatis concepit me mater mea
PS|50|8|ecce enim veritatem dilexisti incerta et occulta sapientiae tuae manifestasti mihi
PS|50|9|asparges me hysopo et mundabor lavabis me et super nivem dealbabor
PS|50|10|auditui meo dabis gaudium et laetitiam exultabunt ossa humiliata
PS|50|11|averte faciem tuam a peccatis meis et omnes iniquitates meas dele
PS|50|12|cor mundum crea in me Deus et spiritum rectum innova in visceribus meis
PS|50|13|ne proicias me a facie tua et spiritum sanctum tuum ne auferas a me
PS|50|14|redde mihi laetitiam salutaris tui et spiritu principali confirma me
PS|50|15|docebo iniquos vias tuas et impii ad te convertentur
PS|50|16|libera me de sanguinibus Deus Deus salutis meae exultabit lingua mea iustitiam tuam
PS|50|17|Domine labia mea aperies et os meum adnuntiabit laudem tuam
PS|50|18|quoniam si voluisses sacrificium dedissem utique holocaustis non delectaberis
PS|50|19|sacrificium Deo spiritus contribulatus cor contritum et humiliatum Deus non spernet
PS|50|20|benigne fac Domine in bona voluntate tua Sion et aedificentur muri Hierusalem
PS|50|21|tunc acceptabis sacrificium iustitiae oblationes et holocausta tunc inponent super altare tuum vitulos
PS|51|1|in finem intellectus David
PS|51|2|cum venit Doec Idumeus et adnuntiavit Saul et dixit venit David in domo Achimelech
PS|51|3|quid gloriatur in malitia qui potens est iniquitate
PS|51|4|tota die iniustitiam cogitavit lingua tua sicut novacula acuta fecisti dolum
PS|51|5|dilexisti malitiam super benignitatem iniquitatem magis quam loqui aequitatem diapsalma
PS|51|6|dilexisti omnia verba praecipitationis linguam dolosam
PS|51|7|propterea Deus destruet te in finem evellet te et emigrabit te de tabernaculo et radicem tuam de terra viventium diapsalma
PS|51|8|videbunt iusti et timebunt et super eum ridebunt et dicent
PS|51|9|ecce homo qui non posuit Deum adiutorem suum sed speravit in multitudine divitiarum suarum et praevaluit in vanitate sua
PS|51|10|ego autem sicut oliva fructifera in domo Dei speravi in misericordia Dei in aeternum et in saeculum saeculi
PS|51|11|confitebor tibi in saeculum quia fecisti et expectabo nomen tuum quoniam bonum in conspectu sanctorum tuorum
PS|52|1|in finem pro Melech intellegentiae David dixit insipiens in corde suo non est Deus
PS|52|2|corrupti sunt et abominabiles facti sunt in iniquitatibus non est qui faciat bonum
PS|52|3|Deus de caelo prospexit in filios hominum ut videat si est intellegens %aut; requirens Deum
PS|52|4|omnes declinaverunt simul inutiles facti sunt non est qui faciat bonum non est usque ad unum
PS|52|5|nonne scient %omnes; qui operantur iniquitatem qui devorant plebem meam ut cibum panis
PS|52|6|Deum non invocaverunt illic trepidabunt timore ubi non fuit timor quoniam Deus dissipavit ossa eorum qui hominibus placent confusi sunt quoniam Deus sprevit eos
PS|52|7|quis dabit ex Sion salutare Israhel dum convertit Deus captivitatem plebis suae exultabit Iacob et laetabitur Israhel
PS|53|1|in finem in carminibus intellectus David
PS|53|2|cum venissent Ziphei et dixissent ad Saul nonne David absconditus est apud nos
PS|53|3|Deus in nomine tuo salvum me fac et in virtute tua iudica me
PS|53|4|Deus exaudi orationem meam auribus percipe verba oris mei
PS|53|5|quoniam alieni insurrexerunt adversum me et fortes quaesierunt animam meam non proposuerunt Deum ante conspectum suum diapsalma
PS|53|6|ecce enim Deus adiuvat me Dominus susceptor animae meae
PS|53|7|avertet mala inimicis meis in veritate tua disperde illos
PS|53|8|voluntarie sacrificabo tibi confitebor nomini tuo Domine quoniam bonum
PS|53|9|quoniam ex omni tribulatione eripuisti me et super inimicos meos despexit oculus meus
PS|54|1|in finem in carminibus intellectus David
PS|54|2|exaudi Deus orationem meam et ne despexeris deprecationem meam
PS|54|3|intende mihi et exaudi me contristatus sum in exercitatione mea et conturbatus sum
PS|54|4|a voce inimici et a tribulatione peccatoris quoniam declinaverunt in me iniquitatem et in ira molesti erant mihi
PS|54|5|cor meum conturbatum est in me et formido mortis cecidit super me
PS|54|6|timor et tremor venit super me et contexit me tenebra
PS|54|7|et dixi quis dabit mihi pinnas sicut columbae et volabo et requiescam
PS|54|8|ecce elongavi fugiens et mansi in solitudine diapsalma
PS|54|9|expectabam eum qui salvum me fecit a pusillanimitate spiritus et a tempestate
PS|54|10|praecipita Domine divide linguas eorum quoniam vidi iniquitatem et contradictionem in civitate
PS|54|11|die et nocte circumdabit eam super muros eius et iniquitas et labor in medio eius
PS|54|12|et iniustitia et non defecit de plateis eius usura et dolus
PS|54|13|quoniam si inimicus maledixisset mihi sustinuissem utique et si is qui oderat me super me magna locutus fuisset abscondissem me forsitan ab eo
PS|54|14|tu vero homo unianimis dux meus et notus meus
PS|54|15|qui simul mecum dulces capiebas cibos in domo Dei ambulavimus cum consensu
PS|54|16|veniat mors super illos et descendant in infernum viventes quoniam nequitiae in habitaculis eorum in medio eorum
PS|54|17|ego %autem; ad Deum clamavi et Dominus salvabit me
PS|54|18|vespere et mane et meridie narrabo et adnuntiabo et exaudiet vocem meam
PS|54|19|redimet in pace animam meam ab his qui adpropinquant mihi quoniam inter multos erant mecum
PS|54|20|exaudiet Deus et humiliabit illos qui est ante saecula diapsalma non enim est illis commutatio et non timuerunt Deum
PS|54|21|extendit manum suam in retribuendo contaminaverunt testamentum eius
PS|54|22|divisi sunt ab ira vultus eius et adpropinquavit cor illius molliti sunt sermones eius super oleum et ipsi sunt iacula
PS|54|23|iacta super Dominum curam tuam et ipse te enutriet non dabit in aeternum fluctuationem iusto
PS|54|24|tu vero Deus deduces eos in puteum interitus viri sanguinum et doli non dimidiabunt dies suos ego autem sperabo in te Domine
PS|55|1|in finem pro populo qui a sanctis longe factus est David in tituli inscriptione cum tenuerunt eum Allophili in Geth
PS|55|2|miserere mei Deus quoniam conculcavit me homo tota die inpugnans tribulavit me
PS|55|3|conculcaverunt me inimici mei tota die quoniam multi bellantes adversum me
PS|55|4|ab altitudine diei timebo ego vero in te sperabo
PS|55|5|in Deo laudabo sermones meos in Deo speravi non timebo quid faciat mihi caro
PS|55|6|tota die verba mea execrabantur adversum me omnia consilia eorum in malum
PS|55|7|inhabitabunt et abscondent ipsi calcaneum meum observabunt sicut sustinuerunt animam meam
PS|55|8|pro nihilo salvos facies illos in ira populos confringes Deus
PS|55|9|vitam meam adnuntiavi tibi posuisti lacrimas meas in conspectu tuo sicut et in promissione tua
PS|55|10|tunc convertentur inimici mei retrorsum in quacumque die invocavero te ecce cognovi quoniam Deus meus es
PS|55|11|in Deo laudabo verbum in Domino laudabo sermonem in Deo speravi non timebo quid faciat mihi homo
PS|55|12|in me sunt Deus vota tua; % quae; reddam laudationes tibi
PS|55|13|quoniam eripuisti animam meam de morte et pedes meos de lapsu ut placeam coram Deo in lumine viventium
PS|56|1|in finem ne disperdas David in tituli inscriptione cum fugeret a facie Saul in spelunca
PS|56|2|miserere mei Deus miserere mei quoniam in te confidit anima mea et in umbra alarum tuarum sperabo donec transeat iniquitas
PS|56|3|clamabo ad Deum altissimum Deum qui benefecit mihi
PS|56|4|misit de caelo et liberavit me dedit in obprobrium conculcantes me diapsalma misit Deus misericordiam suam et veritatem suam
PS|56|5|et eripuit animam meam de medio catulorum leonum dormivi conturbatus filii hominum dentes eorum arma et sagittae et lingua eorum gladius acutus
PS|56|6|exaltare super caelos Deus et in omnem terram gloria tua
PS|56|7|laqueum paraverunt pedibus meis et incurvaverunt animam meam foderunt ante faciem meam foveam et inciderunt in eam diapsalma
PS|56|8|paratum cor meum Deus paratum cor meum cantabo et psalmum dicam
PS|56|9|exsurge gloria mea exsurge psalterium et cithara exsurgam diluculo
PS|56|10|confitebor tibi in populis Domine psalmum dicam tibi in gentibus
PS|56|11|quoniam magnificata est usque ad caelos misericordia tua et usque ad nubes veritas tua
PS|56|12|exaltare super caelos Deus et super omnem terram gloria tua
PS|57|1|in finem ne disperdas David in tituli inscriptione
PS|57|2|si vere utique iustitiam loquimini recta iudicate filii hominum
PS|57|3|etenim in corde iniquitates operamini in terra iniustitiam manus vestrae concinnant
PS|57|4|alienati sunt peccatores a vulva erraverunt ab utero locuti sunt falsa
PS|57|5|furor illis secundum similitudinem serpentis sicut aspidis surdae et obturantis aures suas
PS|57|6|quae non exaudiet vocem incantantium et venefici incantantis sapienter
PS|57|7|Deus conteret dentes eorum in ore ipsorum molas leonum confringet Dominus
PS|57|8|ad nihilum devenient tamquam aqua decurrens intendit arcum suum donec infirmentur
PS|57|9|sicut cera quae fluit auferentur supercecidit ignis et non viderunt solem
PS|57|10|priusquam intellegerent spinae vestrae ramnum sicut viventes sicut in ira absorbet vos
PS|57|11|laetabitur iustus cum viderit vindictam manus suas lavabit in sanguine peccatoris
PS|57|12|et dicet homo si utique est fructus iusto utique est Deus iudicans eos in terra
PS|58|1|in finem ne disperdas David in tituli inscriptione quando misit Saul et custodivit domum eius ut interficeret eum
PS|58|2|eripe me de inimicis meis Deus et ab insurgentibus in me libera me
PS|58|3|eripe me de operantibus iniquitatem et de viris sanguinum salva me
PS|58|4|quia ecce ceperunt animam meam inruerunt in me fortes
PS|58|5|neque iniquitas mea neque peccatum meum Domine sine iniquitate cucurri et direxi
PS|58|6|exsurge in occursum meum et vide et tu Domine Deus virtutum Deus Israhel intende ad visitandas omnes gentes non miserearis omnibus qui operantur iniquitatem diapsalma
PS|58|7|convertentur ad vesperam et famem patientur ut canes et circuibunt civitatem
PS|58|8|ecce loquentur in ore suo et gladius in labiis eorum quoniam quis audivit
PS|58|9|et tu Domine deridebis eos ad nihilum deduces omnes gentes
PS|58|10|fortitudinem meam ad te custodiam quia Deus susceptor meus
PS|58|11|Deus meus voluntas eius praeveniet me
PS|58|12|Deus ostendet mihi super inimicos meos ne occidas eos nequando obliviscantur populi mei disperge illos in virtute tua et depone eos protector meus Domine
PS|58|13|delictum oris eorum sermonem labiorum ipsorum et conprehendantur in superbia sua et de execratione et mendacio adnuntiabuntur
PS|58|14|in consummatione in ira consummationis et non erunt et scient quia Deus dominatur Iacob finium terrae diapsalma
PS|58|15|convertentur ad vesperam et famem patientur ut canes et circuibunt civitatem
PS|58|16|ipsi dispergentur ad manducandum si vero non fuerint saturati et murmurabunt
PS|58|17|ego autem cantabo fortitudinem tuam et exultabo mane misericordiam tuam quia factus es susceptor meus et refugium meum in die tribulationis meae
PS|58|18|adiutor meus tibi psallam quia Deus susceptor meus es Deus meus misericordia mea
PS|59|1|in finem his qui inmutabuntur in tituli inscriptione David in doctrina
PS|59|2|cum succendit Syriam Mesopotamiam et Syriam Soba et convertit Ioab et percussit vallem Salinarum duodecim milia
PS|59|3|Deus reppulisti nos et destruxisti nos iratus es et misertus es nobis
PS|59|4|commovisti terram et turbasti eam sana contritiones eius quia commota est
PS|59|5|ostendisti populo tuo dura potasti nos vino conpunctionis
PS|59|6|dedisti metuentibus te significationem ut fugiant a facie arcus diapsalma ut liberentur dilecti tui
PS|59|7|salvum fac dextera tua et exaudi me
PS|59|8|Deus locutus est in sancto suo laetabor et partibor Sicima et convallem tabernaculorum metibor
PS|59|9|meus est Galaad et meus %est; Manasses et Effraim fortitudo capitis mei Iuda rex meus
PS|59|10|Moab olla spei meae in Idumeam extendam calciamentum meum mihi alienigenae subditi sunt
PS|59|11|quis deducet me in civitatem munitam quis deducet me usque in Idumeam
PS|59|12|nonne tu Deus qui reppulisti nos et non egredieris Deus in virtutibus nostris
PS|59|13|da nobis auxilium de tribulatione et vana salus hominis
PS|59|14|in Deo faciemus virtutem et ipse ad nihilum deducet tribulantes nos
PS|60|1|in finem in hymnis David
PS|60|2|exaudi Deus deprecationem meam intende orationi meae
PS|60|3|a finibus terrae ad te clamavi dum anxiaretur cor meum in petra exaltasti me deduxisti me
PS|60|4|quia factus es spes mea turris fortitudinis a facie inimici
PS|60|5|inhabitabo in tabernaculo tuo in saecula protegar in velamento alarum tuarum diapsalma
PS|60|6|quoniam tu Deus meus exaudisti orationem meam dedisti hereditatem timentibus nomen tuum
PS|60|7|dies super dies regis adicies annos eius usque in diem generationis et generationis
PS|60|8|permanet in aeternum in conspectu Dei misericordiam et veritatem quis requiret eius
PS|60|9|sic psalmum dicam nomini tuo in saeculum saeculi ut reddam vota mea de die in diem
PS|61|1|in finem pro Idithun psalmus David
PS|61|2|nonne Deo subiecta erit anima mea ab ipso enim salutare meum
PS|61|3|nam et ipse Deus meus et salutaris meus susceptor meus non movebor amplius
PS|61|4|quousque inruitis in hominem interficitis universi vos tamquam parieti inclinato et maceriae depulsae
PS|61|5|verumtamen pretium meum cogitaverunt repellere cucurri in siti ore suo benedicebant et corde suo maledicebant diapsalma
PS|61|6|verumtamen Deo subiecta esto anima mea quoniam ab ipso patientia mea
PS|61|7|quia ipse Deus meus et salvator meus adiutor meus non emigrabo
PS|61|8|in Deo salutare meum et gloria mea Deus auxilii mei et spes mea in Deo est
PS|61|9|sperate in eo omnis congregatio populi effundite coram illo corda vestra Deus adiutor noster in aeternum
PS|61|10|verumtamen vani filii hominum mendaces filii hominum in stateris ut decipiant ipsi de vanitate in id ipsum
PS|61|11|nolite sperare in iniquitate et rapinas nolite concupiscere divitiae si affluant nolite cor adponere
PS|61|12|semel locutus est Deus duo haec audivi quia potestas Dei
PS|61|13|et tibi Domine misericordia quia tu reddes unicuique iuxta opera sua
PS|62|1|psalmus David cum esset in deserto Iudaeae
PS|62|2|Deus Deus meus ad te de luce vigilo sitivit in te anima mea quam multipliciter tibi caro mea
PS|62|3|in terra deserta et invia et inaquosa sic in sancto apparui tibi ut viderem virtutem tuam et gloriam tuam
PS|62|4|quoniam melior est misericordia tua super vitas labia mea laudabunt te
PS|62|5|sic benedicam te in vita mea in nomine tuo levabo manus meas
PS|62|6|sicut adipe et pinguidine repleatur anima mea et labia exultationis laudabit os meum
PS|62|7|si memor fui tui super stratum meum in matutinis meditabar in te
PS|62|8|quia fuisti adiutor meus et in velamento alarum tuarum exultabo
PS|62|9|adhesit anima mea post te me suscepit dextera tua
PS|62|10|ipsi vero in vanum quaesierunt animam meam introibunt in inferiora terrae
PS|62|11|tradentur in manus gladii partes vulpium erunt
PS|62|12|rex vero laetabitur in Deo laudabitur omnis qui iurat in eo quia obstructum est os loquentium iniqua
PS|63|1|in finem psalmus David
PS|63|2|exaudi Deus orationem meam cum deprecor a timore inimici eripe animam meam
PS|63|3|protexisti me a conventu malignantium a multitudine operantium iniquitatem
PS|63|4|quia exacuerunt ut gladium linguas suas intenderunt arcum rem amaram
PS|63|5|ut sagittent in occultis inmaculatum
PS|63|6|subito sagittabunt eum et non timebunt firmaverunt sibi sermonem nequam narraverunt ut absconderent laqueos dixerunt quis videbit eos
PS|63|7|scrutati sunt iniquitates defecerunt scrutantes scrutinio accedet homo et cor altum
PS|63|8|et exaltabitur Deus sagittae parvulorum factae sunt plagae eorum
PS|63|9|et infirmatae sunt contra eos linguae eorum conturbati sunt omnes qui videbant eos
PS|63|10|et timuit omnis homo et adnuntiaverunt opera Dei et facta eius intellexerunt
PS|63|11|laetabitur iustus in Domino et sperabit in eo et laudabuntur omnes recti corde
PS|64|1|in finem psalmus David canticum; Hieremiae et Aggei de verbo peregrinationis quando incipiebant proficisci
PS|64|2|te decet hymnus Deus in Sion et tibi reddetur votum in Hierusalem
PS|64|3|exaudi orationem ad te omnis caro veniet
PS|64|4|verba iniquorum praevaluerunt super nos et impietatibus nostris tu propitiaberis
PS|64|5|beatus quem elegisti et adsumpsisti inhabitabit in atriis tuis replebimur in bonis domus tuae sanctum est templum tuum
PS|64|6|mirabile in aequitate exaudi nos Deus salutaris noster spes omnium finium terrae et in mari longe
PS|64|7|praeparans montes in virtute tua accinctus potentia
PS|64|8|qui conturbas profundum maris sonum fluctuum eius turbabuntur gentes
PS|64|9|et timebunt qui inhabitant terminos a signis tuis exitus matutini et vespere delectabis
PS|64|10|visitasti terram et inebriasti eam multiplicasti locupletare eam flumen Dei repletum est aquis parasti cibum illorum quoniam ita est praeparatio eius
PS|64|11|rivos eius inebria multiplica genimina eius in stillicidiis eius laetabitur germinans
PS|64|12|benedices coronae anni benignitatis tuae et campi tui replebuntur ubertate
PS|64|13|pinguescent speciosa deserti et exultatione colles accingentur
PS|64|14|induti sunt arietes ovium et valles abundabunt frumento clamabunt etenim hymnum dicent
PS|65|1|in finem canticum psalmi resurrectionis iubilate Deo omnis terra
PS|65|2|psalmum dicite nomini eius date gloriam laudi eius
PS|65|3|dicite Deo quam terribilia sunt opera tua Domine in multitudine virtutis tuae mentientur tibi inimici tui
PS|65|4|omnis terra adorent te et psallant tibi psalmum dicant nomini tuo diapsalma
PS|65|5|venite et videte opera Dei terribilis in consiliis super filios hominum
PS|65|6|qui convertit mare in aridam in flumine pertransibunt pede ibi laetabimur in ipso
PS|65|7|qui dominatur in virtute sua in aeternum oculi eius super gentes respiciunt qui exasperant non exaltentur in semet ipsis diapsalma
PS|65|8|benedicite gentes Deum nostrum et auditam facite vocem laudis eius
PS|65|9|qui posuit animam meam ad vitam et non dedit in commotionem pedes meos
PS|65|10|quoniam probasti nos Deus igne nos examinasti sicut examinatur argentum
PS|65|11|induxisti nos in laqueum posuisti tribulationes in dorso nostro
PS|65|12|inposuisti homines super capita nostra transivimus per ignem et aquam et eduxisti nos in refrigerium
PS|65|13|introibo in domum tuam in holocaustis reddam tibi vota mea
PS|65|14|quae distinxerunt labia mea et locutum est os meum in tribulatione mea
PS|65|15|holocausta medullata offeram tibi cum incensu arietum offeram tibi boves cum hircis diapsalma
PS|65|16|venite audite et narrabo omnes qui timetis Deum quanta fecit animae meae
PS|65|17|ad ipsum ore meo clamavi et exaltavi sub lingua mea
PS|65|18|iniquitatem si aspexi in corde meo non exaudiat Dominus
PS|65|19|propterea exaudivit Deus adtendit voci deprecationis meae
PS|65|20|benedictus Deus qui non amovit orationem meam et misericordiam suam a me
PS|66|1|in finem in hymnis psalmus cantici
PS|66|2|Deus misereatur nostri et benedicat nobis inluminet vultum suum super nos et misereatur nostri diapsalma
PS|66|3|ut cognoscamus in terra viam tuam in omnibus gentibus salutare tuum
PS|66|4|confiteantur tibi populi Deus confiteantur tibi populi omnes
PS|66|5|laetentur et exultent gentes quoniam iudicas populos in aequitate et gentes in terra diriges diapsalma
PS|66|6|confiteantur tibi populi Deus confiteantur tibi populi omnes
PS|66|7|terra dedit fructum suum benedicat nos Deus Deus noster
PS|66|8|benedicat nos Deus et metuant eum omnes fines terrae
PS|67|1|in finem David psalmus cantici
PS|67|2|exsurgat Deus et dissipentur inimici eius et fugiant qui oderunt eum a facie eius
PS|67|3|sicut deficit fumus deficiant sicut fluit cera a facie ignis sic pereant peccatores a facie Dei
PS|67|4|et iusti epulentur exultent in conspectu Dei delectentur in laetitia
PS|67|5|cantate Deo psalmum dicite nomini eius iter facite ei qui ascendit super occasum Dominus nomen illi et exultate in conspectu eius turbabuntur a facie eius
PS|67|6|patris orfanorum et iudicis viduarum Deus in loco sancto suo
PS|67|7|Deus inhabitare facit unius moris in domo qui educit vinctos in fortitudine similiter eos qui exasperant qui habitant in sepulchris
PS|67|8|Deus cum egredereris in conspectu populi tui cum pertransieris in deserto diapsalma
PS|67|9|terra mota est etenim caeli distillaverunt a facie Dei Sinai a facie Dei Israhel
PS|67|10|pluviam voluntariam segregabis Deus hereditati tuae et infirmata est tu vero perfecisti eam
PS|67|11|animalia tua habitant in ea parasti in dulcedine tua pauperi Deus
PS|67|12|Dominus dabit verbum evangelizantibus virtute multa
PS|67|13|rex virtutum dilecti dilecti; et speciei domus dividere spolia
PS|67|14|si dormiatis inter medios cleros pinnae columbae deargentatae et posteriora dorsi eius in pallore auri
PS|67|15|dum discernit Caelestis reges super eam nive dealbabuntur in Selmon
PS|67|16|mons Dei mons pinguis mons coagulatus mons pinguis
PS|67|17|ut quid suspicamini montes coagulatos mons in quo beneplacitum est Deo habitare in eo etenim Dominus habitabit in finem
PS|67|18|currus Dei decem milibus multiplex milia laetantium Dominus in eis in Sina in sancto
PS|67|19|ascendisti in altum cepisti captivitatem accepisti dona in hominibus etenim non credentes inhabitare Dominum Deus
PS|67|20|benedictus Dominus die cotidie prosperum iter faciet nobis Deus salutarium nostrorum diapsalma
PS|67|21|Deus noster Deus salvos faciendi et Domini Domini exitus mortis
PS|67|22|verumtamen Deus confringet capita inimicorum suorum verticem capilli perambulantium in delictis suis
PS|67|23|dixit Dominus ex Basan convertam convertam in profundis maris
PS|67|24|ut intinguatur pes tuus in sanguine lingua canum tuorum ex inimicis ab ipso
PS|67|25|viderunt ingressus tui Deus ingressus Dei mei regis mei qui est in sancto
PS|67|26|praevenerunt principes coniuncti psallentibus in medio iuvencularum tympanistriarum
PS|67|27|in ecclesiis benedicite Deum Dominum de fontibus Israhel
PS|67|28|ibi Beniamin adulescentulus in mentis excessu principes Iuda duces eorum principes Zabulon principes Nepthali
PS|67|29|manda Deus virtutem tuam confirma Deus hoc quod operatus es nobis
PS|67|30|a templo tuo in Hierusalem tibi adferent reges munera
PS|67|31|increpa feras harundinis congregatio taurorum in vaccis populorum ut excludant eos qui probati sunt argento dissipa gentes quae bella volunt
PS|67|32|venient legati ex Aegypto Aethiopia praeveniet manus eius Deo
PS|67|33|regna terrae cantate Deo psallite Domino diapsalma %psallite Deo;
PS|67|34|qui ascendit super caelum caeli ad orientem ecce dabit voci suae vocem virtutis
PS|67|35|date gloriam Deo super Israhel magnificentia eius et virtus eius in nubibus
PS|67|36|mirabilis Deus in sanctis suis Deus Israhel ipse dabit virtutem et fortitudinem plebi suae benedictus Deus
PS|68|1|in finem pro his qui commutabuntur David
PS|68|2|salvum me fac Deus quoniam intraverunt aquae usque ad animam meam
PS|68|3|infixus sum in limum profundi et non est substantia veni in altitudines maris et tempestas demersit me
PS|68|4|laboravi clamans raucae factae sunt fauces meae defecerunt oculi mei dum spero in Deum meum
PS|68|5|multiplicati sunt super capillos capitis mei qui oderunt me gratis confortati sunt qui persecuti sunt me inimici mei iniuste quae non rapui tunc exsolvebam
PS|68|6|Deus tu scis insipientiam meam et delicta mea a te non sunt abscondita
PS|68|7|non erubescant in me qui expectant te Domine Domine virtutum non confundantur super me qui quaerunt te Deus Israhel
PS|68|8|quoniam propter te sustinui obprobrium operuit confusio faciem meam
PS|68|9|extraneus factus sum fratribus meis et peregrinus filiis matris meae
PS|68|10|quoniam zelus domus tuae comedit me et obprobria exprobrantium tibi ceciderunt super me
PS|68|11|et operui in ieiunio animam meam et factum est in obprobrium mihi
PS|68|12|et posui vestimentum meum cilicium et factus sum illis in parabolam
PS|68|13|adversum me exercebantur qui sedebant in porta et in me psallebant qui bibebant vinum
PS|68|14|ego vero orationem meam ad te Domine tempus beneplaciti Deus in multitudine misericordiae tuae exaudi me in veritate salutis tuae
PS|68|15|eripe me de luto ut non infigar liberer ab his qui oderunt me et de profundis aquarum
PS|68|16|non me demergat tempestas aquae neque absorbeat me profundum neque urgeat super me puteus os suum
PS|68|17|exaudi me Domine quoniam benigna est misericordia tua secundum multitudinem miserationum tuarum respice me
PS|68|18|et ne avertas faciem tuam a puero tuo quoniam tribulor velociter exaudi me
PS|68|19|intende animae meae et libera eam propter inimicos meos eripe me
PS|68|20|tu scis inproperium meum et confusionem et reverentiam meam
PS|68|21|in conspectu tuo sunt omnes qui tribulant me inproperium expectavit cor meum et miseriam et sustinui qui simul contristaretur et non fuit et qui consolaretur et non inveni
PS|68|22|et dederunt in escam meam fel et in siti mea potaverunt me aceto
PS|68|23|fiat mensa eorum coram ipsis in laqueum et in retributiones et in scandalum
PS|68|24|obscurentur oculi eorum ne videant et dorsum eorum semper incurva
PS|68|25|effunde super eos iram tuam et furor irae tuae conprehendat eos
PS|68|26|fiat habitatio eorum deserta et in tabernaculis eorum non sit qui inhabitet
PS|68|27|quoniam quem tu percussisti persecuti sunt et super dolorem vulnerum meorum addiderunt
PS|68|28|adpone iniquitatem super iniquitatem eorum et non intrent in iustitia tua
PS|68|29|deleantur de libro viventium et cum iustis non scribantur
PS|68|30|ego sum pauper et dolens salus tua Deus suscepit me
PS|68|31|laudabo nomen Dei cum cantico magnificabo eum in laude
PS|68|32|et placebit Deo super vitulum novellum cornua producentem et ungulas
PS|68|33|videant pauperes et laetentur quaerite Deum et vivet anima vestra
PS|68|34|quoniam exaudivit pauperes Dominus et vinctos suos non despexit
PS|68|35|laudent illum caeli et terra mare et omnia reptilia in eis
PS|68|36|quoniam Deus salvam faciet Sion et aedificabuntur civitates Iudaeae et inhabitabunt ibi et hereditate adquirent eam
PS|68|37|et semen servorum eius possidebunt eam et qui diligunt nomen eius habitabunt in ea
PS|69|1|in finem David in rememoratione eo quod salvum me fecit Dominus
PS|69|2|Deus in adiutorium meum intende Domine ad adiuvandum me festina;
PS|69|3|confundantur et revereantur qui quaerunt animam meam
PS|69|4|avertantur retrorsum et erubescant qui volunt mihi mala avertantur statim erubescentes qui dicunt %mihi; euge euge
PS|69|5|exultent et laetentur in te omnes qui quaerunt te et dicant semper magnificetur Deus qui diligunt salutare tuum
PS|69|6|ego vero egenus et pauper Deus adiuva me adiutor meus et liberator meus es tu Domine ne moreris
PS|69|7|
PS|69|8|
PS|69|9|
PS|70|1|David psalmus filiorum Ionadab et priorum captivorum in te Domine speravi non confundar in aeternum
PS|70|2|in iustitia tua libera me et eripe me inclina ad me aurem tuam et salva me
PS|70|3|esto mihi in Deum protectorem et in locum munitum ut salvum me facias quoniam firmamentum meum et refugium meum es tu
PS|70|4|Deus meus eripe me de manu peccatoris de manu contra legem agentis et iniqui
PS|70|5|quoniam tu es patientia mea Domine Domine spes mea a iuventute mea
PS|70|6|in te confirmatus sum ex utero de ventre matris meae tu es protector meus in te cantatio mea semper
PS|70|7|tamquam prodigium factus sum multis et tu adiutor fortis
PS|70|8|repleatur os meum laude ut cantem gloriam tuam tota die magnitudinem tuam
PS|70|9|non proicias me in tempore senectutis cum deficiet virtus mea ne derelinquas me
PS|70|10|quia dixerunt inimici mei mihi et qui custodiebant animam meam consilium fecerunt in unum
PS|70|11|dicentes Deus dereliquit eum persequimini et conprehendite eum quia non est qui eripiat
PS|70|12|Deus ne elongeris a me Deus meus in adiutorium meum respice
PS|70|13|confundantur et deficiant detrahentes animae meae operiantur confusione et pudore qui quaerunt mala mihi
PS|70|14|ego autem semper sperabo et adiciam super omnem laudem tuam
PS|70|15|os meum adnuntiabit iustitiam tuam tota die salutem tuam quoniam non cognovi litteraturam
PS|70|16|introibo in potentiam Domini Domine memorabor iustitiae tuae solius
PS|70|17|Deus docuisti me ex iuventute mea et usque nunc pronuntiabo mirabilia tua
PS|70|18|et usque in senectam et senium Deus ne derelinquas me donec adnuntiem brachium tuum generationi omni quae ventura est potentiam tuam
PS|70|19|et iustitiam tuam Deus usque in altissima quae fecisti magnalia Deus quis similis tibi
PS|70|20|quantas ostendisti mihi tribulationes multas et malas et conversus vivificasti me et de abyssis terrae iterum reduxisti me
PS|70|21|multiplicasti magnificentiam tuam et conversus consolatus es me
PS|70|22|nam et ego confitebor tibi in vasis psalmi veritatem tuam Deus psallam tibi in cithara Sanctus Israhel
PS|70|23|exultabunt labia mea cum cantavero tibi et anima mea quam redemisti
PS|70|24|sed et lingua mea tota die meditabitur iustitiam tuam cum confusi et reveriti fuerint qui quaerunt mala mihi
PS|71|1|in Salomonem
PS|71|2|Deus iudicium tuum regi da et iustitiam tuam filio regis iudicare populum tuum in iustitia et pauperes tuos in iudicio
PS|71|3|suscipiant montes pacem populo et colles iustitiam
PS|71|4|iudicabit pauperes populi et salvos faciet filios pauperum et humiliabit calumniatorem
PS|71|5|et permanebit cum sole et ante lunam generationes generationum
PS|71|6|descendet sicut pluvia in vellus et sicut stillicidia stillantia super terram
PS|71|7|orietur in diebus eius iustitia et abundantia pacis donec auferatur luna
PS|71|8|et dominabitur a mari usque ad mare et a flumine usque ad terminos orbis terrarum
PS|71|9|coram illo procident Aethiopes et inimici eius terram lingent
PS|71|10|reges Tharsis et insulae munera offerent reges Arabum et Saba dona adducent
PS|71|11|et adorabunt eum omnes reges omnes gentes servient ei
PS|71|12|quia liberavit pauperem a potente et pauperem cui non erat adiutor
PS|71|13|parcet pauperi et inopi et animas pauperum salvas faciet
PS|71|14|ex usuris et iniquitate redimet animas eorum et honorabile nomen eorum coram illo
PS|71|15|et vivet et dabitur ei de auro Arabiae et orabunt de ipso semper tota die benedicent ei
PS|71|16|erit firmamentum in terra in summis montium superextolletur super Libanum fructus eius et florebunt de civitate sicut faenum terrae
PS|71|17|sit nomen eius benedictum in saecula ante solem permanet nomen eius et benedicentur in ipso omnes tribus terrae omnes gentes beatificabunt eum
PS|71|18|benedictus Dominus Deus Deus Israhel qui facit mirabilia solus
PS|71|19|et benedictum nomen maiestatis eius in aeternum et replebitur maiestate eius omnis terra fiat fiat
PS|71|20|defecerunt laudes David filii Iesse
PS|72|1|psalmus Asaph quam bonus Israhel Deus his qui recto sunt corde
PS|72|2|mei autem paene moti sunt pedes paene effusi sunt gressus mei
PS|72|3|quia zelavi super iniquis pacem peccatorum videns
PS|72|4|quia non est respectus morti eorum et firmamentum in plaga eorum
PS|72|5|in labore hominum non sunt et cum hominibus non flagellabuntur
PS|72|6|ideo tenuit eos superbia operti sunt iniquitate et impietate sua
PS|72|7|prodiet quasi ex adipe iniquitas eorum transierunt in affectum cordis
PS|72|8|cogitaverunt et locuti sunt in nequitia iniquitatem in excelso locuti sunt
PS|72|9|posuerunt in caelum os suum et lingua eorum transivit in terra
PS|72|10|ideo convertetur populus meus hic et dies pleni invenientur in eis
PS|72|11|et dixerunt quomodo scit Deus et si est scientia in Excelso
PS|72|12|ecce ipsi peccatores et abundantes in saeculo obtinuerunt divitias
PS|72|13|%et dixi; ergo sine causa iustificavi cor meum et lavi inter innocentes manus meas
PS|72|14|et fui flagellatus tota die et castigatio mea in matutino
PS|72|15|si dicebam narrabo sic ecce nationem filiorum tuorum reprobavi
PS|72|16|et existimabam cognoscere hoc labor est ante me
PS|72|17|donec intrem in sanctuarium Dei intellegam in novissimis eorum
PS|72|18|verumtamen propter dolos posuisti eis deiecisti eos dum adlevarentur
PS|72|19|quomodo facti sunt in desolationem subito defecerunt perierunt propter iniquitatem suam
PS|72|20|velut somnium surgentium Domine in civitate tua imaginem ipsorum ad nihilum rediges
PS|72|21|quia inflammatum est cor meum et renes mei commutati sunt
PS|72|22|et ego ad nihilum redactus sum et nescivi
PS|72|23|ut iumentum factus sum apud te et ego semper tecum
PS|72|24|tenuisti manum dexteram meam et in voluntate tua deduxisti me et cum gloria suscepisti me
PS|72|25|quid enim mihi est in caelo et a te quid volui super terram
PS|72|26|defecit caro mea et cor meum Deus cordis mei et pars mea Deus in aeternum
PS|72|27|quia ecce qui elongant se a te peribunt perdidisti omnem qui fornicatur abs te
PS|72|28|mihi autem adherere Deo bonum est ponere in Domino Deo spem meam ut adnuntiem omnes praedicationes tuas % in portis filiae Sion;
PS|73|1|intellectus Asaph ut quid Deus reppulisti in finem iratus est furor tuus super oves pascuae tuae
PS|73|2|memor esto congregationis tuae quam possedisti ab initio redemisti virgam hereditatis tuae mons Sion in quo habitasti in eo
PS|73|3|leva manus tuas in superbias eorum in finem quanta malignatus est inimicus in sancto
PS|73|4|et gloriati sunt qui oderunt te in medio sollemnitatis tuae posuerunt signa sua signa
PS|73|5|et non cognoverunt sicut in exitu super summum quasi in silva lignorum securibus
PS|73|6|exciderunt ianuas eius in id ipsum in securi et ascia deiecerunt %eam;
PS|73|7|incenderunt igni sanctuarium tuum in terra polluerunt tabernaculum nominis tui
PS|73|8|dixerunt in corde suo cognatio eorum simul quiescere faciamus omnes dies festos Dei a terra
PS|73|9|signa nostra non vidimus iam non est propheta et nos non cognoscet amplius
PS|73|10|usquequo Deus inproperabit inimicus inritat adversarius nomen tuum in finem
PS|73|11|ut quid avertis manum tuam et dexteram tuam de medio sinu tuo in finem
PS|73|12|Deus autem rex noster ante saeculum operatus est salutes in medio terrae
PS|73|13|tu confirmasti in virtute tua mare contribulasti capita draconum in aquis
PS|73|14|tu confregisti capita draconis dedisti eum escam populis Aethiopum
PS|73|15|tu disrupisti fontem et torrentes tu siccasti fluvios Aetham;
PS|73|16|tuus est dies et tua est nox tu fabricatus es auroram et solem
PS|73|17|tu fecisti omnes terminos terrae aestatem et ver tu plasmasti ea
PS|73|18|memor esto huius inimicus inproperavit Dominum et populus insipiens incitavit nomen tuum
PS|73|19|ne tradas bestiis animam confitentem tibi animas pauperum tuorum ne obliviscaris in finem
PS|73|20|respice in testamentum tuum quia repleti sunt qui obscurati sunt terrae domibus iniquitatum
PS|73|21|ne avertatur humilis factus confusus pauper et inops laudabunt nomen tuum
PS|73|22|exsurge Deus iudica causam tuam memor esto inproperiorum tuorum eorum qui ab insipiente sunt tota die
PS|73|23|ne obliviscaris voces inimicorum tuorum superbia eorum qui te oderunt ascendit semper
PS|74|1|in finem ne corrumpas psalmus Asaph cantici
PS|74|2|confitebimur tibi Deus confitebimur et invocabimus nomen tuum narrabimus mirabilia tua
PS|74|3|cum accepero tempus ego iustitias iudicabo
PS|74|4|liquefacta est terra et omnes qui habitant in ea ego confirmavi columnas eius diapsalma
PS|74|5|dixi iniquis nolite inique facere et delinquentibus nolite exaltare cornu
PS|74|6|nolite extollere in altum cornu vestrum nolite loqui adversus Deum iniquitatem
PS|74|7|quia neque ab oriente neque ab occidente neque a desertis montibus
PS|74|8|quoniam Deus iudex est hunc humiliat et hunc exaltat
PS|74|9|quia calix in manu Domini vini meri plenus mixto et inclinavit ex hoc in hoc verum fex eius non est exinanita bibent omnes peccatores terrae
PS|74|10|ego autem adnuntiabo in saeculum cantabo Deo Iacob
PS|74|11|et omnia cornua peccatorum confringam et exaltabuntur cornua iusti
PS|75|1|in finem in laudibus psalmus Asaph canticum ad Assyrium
PS|75|2|notus in Iudaea Deus in Israhel magnum nomen eius
PS|75|3|et factus est in pace locus eius et habitatio eius in Sion
PS|75|4|ibi confregit potentias arcuum scutum et gladium et bellum diapsalma
PS|75|5|inluminas tu mirabiliter de montibus aeternis
PS|75|6|turbati sunt omnes insipientes corde dormierunt somnum suum et nihil invenerunt omnes viri divitiarum manibus suis
PS|75|7|ab increpatione tua Deus Iacob dormitaverunt qui ascenderunt equos
PS|75|8|tu terribilis es et quis resistet tibi ex tunc ira tua
PS|75|9|de caelo auditum fecisti iudicium terra timuit et quievit
PS|75|10|cum exsurgeret in iudicium Deus ut salvos faceret omnes mansuetos terrae diapsalma
PS|75|11|quoniam cogitatio hominis confitebitur tibi et reliquiae cogitationis diem festum agent tibi
PS|75|12|vovete et reddite Domino Deo vestro omnes qui in circuitu eius adferent munera terribili
PS|75|13|et ei qui aufert spiritus principum terribili apud reges terrae
PS|76|1|in finem pro Idithun psalmus Asaph
PS|76|2|voce mea ad Dominum clamavi voce mea ad Deum et intendit me
PS|76|3|in die tribulationis meae Deum exquisivi manibus meis nocte contra eum et non sum deceptus rennuit consolari anima mea
PS|76|4|memor fui Dei et delectatus sum exercitatus sum et defecit spiritus meus diapsalma
PS|76|5|anticipaverunt vigilias oculi mei turbatus sum et non sum locutus
PS|76|6|cogitavi dies antiquos et annos aeternos in mente habui
PS|76|7|et meditatus sum nocte cum corde meo exercitabar et scobebam spiritum meum
PS|76|8|numquid in aeternum proiciet Deus et non adponet ut conplacitior sit adhuc
PS|76|9|aut in finem misericordiam suam abscidet a generatione in generationem
PS|76|10|aut obliviscetur misereri Deus aut continebit in ira sua misericordias suas diapsalma
PS|76|11|et dixi nunc coepi haec mutatio dexterae Excelsi
PS|76|12|memor fui operum Domini quia memor ero ab initio mirabilium tuorum
PS|76|13|et meditabor in omnibus operibus tuis et in adinventionibus tuis exercebor
PS|76|14|Deus in sancto via tua quis deus magnus sicut Deus noster
PS|76|15|tu es Deus qui facis mirabilia notam fecisti in populis virtutem tuam
PS|76|16|redemisti in brachio tuo populum tuum filios Iacob et Ioseph diapsalma
PS|76|17|viderunt te aquae Deus viderunt te aquae et timuerunt et turbatae sunt abyssi
PS|76|18|multitudo sonitus aquarum vocem dederunt nubes etenim sagittae tuae transeunt
PS|76|19|vox tonitrui tui in rota inluxerunt coruscationes tuae orbi terrae commota est et contremuit terra
PS|76|20|in mari via tua et semitae tuae in aquis multis et vestigia tua non cognoscentur
PS|76|21|deduxisti sicut oves populum tuum in manu Mosi et Aaron
PS|77|1|intellectus Asaph adtendite populus meus legem meam inclinate aurem vestram in verba oris mei
PS|77|2|aperiam in parabola os meum eloquar propositiones ab initio
PS|77|3|quanta audivimus et cognovimus ea et patres nostri narraverunt nobis
PS|77|4|non sunt occultata a filiis eorum in generationem alteram narrantes laudes Domini et virtutes eius et mirabilia eius quae fecit
PS|77|5|et suscitavit testimonium in Iacob et legem posuit in Israhel quanta mandavit patribus nostris nota facere ea filiis suis
PS|77|6|ut cognoscat generatio altera filii qui nascentur et exsurgent et narrabunt filiis suis
PS|77|7|ut ponant in Deo spem suam et non obliviscantur opera Dei et mandata eius exquirant
PS|77|8|ne fiant sicut patres eorum generatio prava et exasperans generatio quae non direxit cor suum et non est creditus cum Deo spiritus eius
PS|77|9|filii Effrem intendentes et mittentes arcus conversi sunt in die belli
PS|77|10|non custodierunt testamentum Dei et in lege eius noluerunt ambulare
PS|77|11|et obliti sunt benefactorum eius et mirabilium eius quae ostendit eis
PS|77|12|coram patribus eorum quae fecit mirabilia in terra Aegypti in campo Taneos
PS|77|13|interrupit mare et perduxit eos statuit aquas quasi utrem
PS|77|14|et deduxit eos in nube diei et tota nocte in inluminatione ignis
PS|77|15|interrupit petram in heremo et adaquavit eos velut in abysso multa
PS|77|16|et eduxit aquam de petra et deduxit tamquam flumina aquas
PS|77|17|et adposuerunt adhuc peccare ei in ira excitaverunt Excelsum in inaquoso
PS|77|18|et temptaverunt Deum in cordibus suis ut peterent escas animabus suis
PS|77|19|et male locuti sunt de Deo dixerunt numquid poterit Deus parare mensam in deserto
PS|77|20|quoniam percussit petram et fluxerunt aquae et torrentes inundaverunt numquid et panem potest dare aut parare mensam populo suo
PS|77|21|ideo audivit Dominus et distulit et ignis accensus est in Iacob et ira ascendit in Israhel
PS|77|22|quia non crediderunt in Deo nec speraverunt in salutare eius
PS|77|23|et mandavit nubibus desuper et ianuas caeli aperuit
PS|77|24|et pluit illis manna ad manducandum et panem caeli dedit eis
PS|77|25|panem angelorum manducavit homo cibaria misit eis in abundantiam
PS|77|26|transtulit austrum de caelo et induxit in virtute sua africum
PS|77|27|et pluit super eos sicut pulverem carnes et sicut harenam maris volatilia pinnata
PS|77|28|et ceciderunt in medio castrorum eorum circa tabernacula eorum
PS|77|29|et manducaverunt et saturati sunt nimis et desiderium eorum adtulit eis
PS|77|30|non sunt fraudati a desiderio suo adhuc escae eorum erant in ore ipsorum
PS|77|31|et ira Dei ascendit in eos et occidit pingues eorum et electos Israhel inpedivit
PS|77|32|in omnibus his peccaverunt adhuc et non crediderunt mirabilibus eius
PS|77|33|et defecerunt in vanitate dies eorum et anni eorum cum festinatione
PS|77|34|cum occideret eos quaerebant eum et revertebantur et diluculo veniebant ad Deum
PS|77|35|et rememorati sunt quia Deus adiutor est eorum et Deus excelsus redemptor eorum est
PS|77|36|et dilexerunt eum in ore suo et lingua sua mentiti sunt ei
PS|77|37|cor autem ipsorum non erat rectum cum eo nec fideles habiti sunt in testamento eius
PS|77|38|ipse autem est misericors et propitius fiet peccatis eorum et non perdet eos et abundabit ut avertat iram suam et non accendet omnem iram suam
PS|77|39|et recordatus est quia caro sunt spiritus vadens et non rediens
PS|77|40|quotiens exacerbaverunt eum in deserto in ira concitaverunt eum in inaquoso
PS|77|41|et conversi sunt et temptaverunt Deum et Sanctum Israhel exacerbaverunt
PS|77|42|non sunt recordati manus eius die qua redemit eos de manu tribulantis
PS|77|43|sicut posuit in Aegypto signa sua et prodigia sua in campo Taneos
PS|77|44|et convertit in sanguine flumina eorum et imbres eorum ne biberent
PS|77|45|misit in eos cynomiam et comedit eos et ranam et disperdit eos
PS|77|46|et dedit erugini fructus eorum et labores eorum lucustae
PS|77|47|et occidit in grandine vineam eorum et moros eorum in pruina
PS|77|48|et tradidit grandini iumenta eorum et possessionem eorum igni
PS|77|49|misit in eos iram indignationis suae indignationem et iram et tribulationem inmissionem per angelos malos
PS|77|50|viam fecit semitae irae suae non pepercit a morte animarum eorum et iumenta eorum in morte conclusit
PS|77|51|et percussit omne primitivum in terra Aegypti primitias laborum eorum in tabernaculis Cham
PS|77|52|et abstulit sicut oves populum suum et perduxit eos tamquam gregem in deserto
PS|77|53|et deduxit eos in spe et non timuerunt et inimicos eorum operuit mare
PS|77|54|et induxit eos in montem sanctificationis suae montem quem adquisivit dextera eius et eiecit a facie eorum gentes et sorte divisit eis terram in funiculo distributionis
PS|77|55|et habitare fecit in tabernaculis eorum tribus Israhel
PS|77|56|et temptaverunt et exacerbaverunt Deum excelsum et testimonia eius non custodierunt
PS|77|57|et averterunt se et non servaverunt pactum quemadmodum patres eorum conversi sunt in arcum pravum
PS|77|58|et in ira concitaverunt eum in collibus suis et in sculptilibus suis ad aemulationem eum provocaverunt
PS|77|59|audivit Deus et sprevit et ad nihilum redegit valde Israhel
PS|77|60|et reppulit tabernaculum Selo tabernaculum suum ubi habitavit in hominibus
PS|77|61|et tradidit in captivitatem virtutem eorum et pulchritudinem eorum in manus inimici
PS|77|62|et conclusit in gladio populum suum et hereditatem suam sprevit
PS|77|63|iuvenes eorum comedit ignis et virgines eorum non sunt lamentatae
PS|77|64|sacerdotes eorum in gladio ceciderunt et viduae eorum non plorabuntur
PS|77|65|et excitatus est tamquam dormiens Dominus tamquam potens crapulatus a vino
PS|77|66|et percussit inimicos suos in posteriora obprobrium sempiternum dedit illis
PS|77|67|et reppulit tabernaculum Ioseph et tribum Effrem non elegit
PS|77|68|et elegit tribum Iuda montem Sion quem dilexit
PS|77|69|et aedificavit sicut unicornium sanctificium suum in terra quam fundavit in saecula
PS|77|70|et elegit David servum suum et sustulit eum de gregibus ovium de post fetantes accepit eum
PS|77|71|pascere Iacob servum suum et Israhel hereditatem suam
PS|77|72|et pavit eos in innocentia cordis sui et in intellectibus manuum suarum deduxit eos
PS|78|1|psalmus Asaph Deus venerunt gentes in hereditatem tuam polluerunt templum sanctum tuum posuerunt Hierusalem in pomorum custodiam
PS|78|2|posuerunt morticina servorum tuorum escas volatilibus caeli carnes sanctorum tuorum bestiis terrae
PS|78|3|effuderunt sanguinem ipsorum tamquam aquam in circuitu Hierusalem et non erat qui sepeliret
PS|78|4|facti sumus obprobrium vicinis nostris subsannatio et inlusio his qui circum nos sunt
PS|78|5|usquequo Domine irasceris in finem accendetur velut ignis zelus tuus
PS|78|6|effunde iram tuam in gentes quae te non noverunt et in regna quae nomen tuum non invocaverunt
PS|78|7|quia comederunt Iacob et locum eius desolaverunt
PS|78|8|ne memineris iniquitatum nostrarum antiquarum cito anticipent nos misericordiae tuae quia pauperes facti sumus nimis
PS|78|9|adiuva nos Deus salutaris noster propter gloriam nominis tui Domine libera nos et propitius esto peccatis nostris propter nomen tuum
PS|78|10|ne forte dicant in gentibus ubi est Deus eorum et innotescat in nationibus coram oculis nostris ultio sanguinis servorum tuorum qui effusus est
PS|78|11|introeat in conspectu tuo gemitus conpeditorum secundum magnitudinem brachii tui posside filios mortificatorum
PS|78|12|et redde vicinis nostris septuplum in sinu eorum inproperium ipsorum quod exprobraverunt tibi Domine
PS|78|13|nos autem populus tuus et oves pascuae tuae confitebimur tibi in saeculum in generationem et generationem adnuntiabimus laudem tuam
PS|79|1|in finem pro his qui commutabuntur testimonium Asaph psalmus
PS|79|2|qui regis Israhel intende qui deducis tamquam oves Ioseph qui sedes super cherubin manifestare
PS|79|3|coram Effraim et Beniamin et Manasse excita potentiam tuam et veni ut salvos facias nos
PS|79|4|Deus converte nos et ostende faciem tuam et salvi erimus
PS|79|5|Domine Deus virtutum quousque irasceris super orationem servi tui
PS|79|6|cibabis nos pane lacrimarum et potum dabis nobis in lacrimis in mensura
PS|79|7|posuisti nos in contradictionem vicinis nostris et inimici nostri subsannaverunt nos
PS|79|8|Deus virtutum converte nos et ostende faciem tuam et salvi erimus
PS|79|9|vineam de Aegypto transtulisti eiecisti gentes et plantasti eam
PS|79|10|dux itineris fuisti in conspectu eius et plantasti radices eius et implevit terram
PS|79|11|operuit montes umbra eius et arbusta eius cedros Dei
PS|79|12|extendit palmites suos usque ad mare et usque ad Flumen propagines eius
PS|79|13|ut quid destruxisti maceriam eius et vindemiant eam omnes qui praetergrediuntur viam
PS|79|14|exterminavit eam aper de silva et singularis ferus depastus est eam
PS|79|15|Deus virtutum convertere respice de caelo et vide et visita vineam istam
PS|79|16|et perfice eam quam plantavit dextera tua et super filium quem confirmasti tibi
PS|79|17|incensa igni et suffossa ab increpatione vultus tui peribunt
PS|79|18|fiat manus tua super virum dexterae tuae et super filium hominis quem confirmasti tibi
PS|79|19|et non discedimus a te vivificabis nos et nomen tuum invocabimus
PS|79|20|Domine Deus virtutum converte nos et ostende faciem tuam et salvi erimus
PS|80|1|in finem pro torcularibus Asaph
PS|80|2|exultate Deo adiutori nostro iubilate Deo Iacob
PS|80|3|sumite psalmum et date tympanum psalterium iucundum cum cithara
PS|80|4|bucinate in neomenia tuba in insigni die sollemnitatis nostrae
PS|80|5|quia praeceptum Israhel est et iudicium Dei Iacob
PS|80|6|testimonium in Ioseph posuit illud cum exiret de terra Aegypti linguam quam non noverat audivit
PS|80|7|devertit ab oneribus dorsum eius manus eius in cofino servierunt
PS|80|8|in tribulatione invocasti me et liberavi te exaudivi te in abscondito tempestatis probavi te apud aquam Contradictionis diapsalma
PS|80|9|audi populus meus et contestabor te Israhel si audias me
PS|80|10|non erit in te deus recens nec adorabis deum alienum
PS|80|11|ego enim sum Dominus Deus tuus qui eduxi te de terra Aegypti dilata os tuum et implebo illud
PS|80|12|et non audivit populus meus vocem meam et Israhel non intendit mihi
PS|80|13|et dimisi illos secundum desideria cordis eorum ibunt in adinventionibus suis
PS|80|14|si populus meus audisset me Israhel si in viis meis ambulasset
PS|80|15|pro nihilo forsitan inimicos eorum humiliassem et super tribulantes eos misissem manum meam
PS|80|16|inimici Domini mentiti sunt ei et erit tempus eorum in saeculo
PS|80|17|et cibavit illos ex adipe frumenti et de petra melle saturavit illos
PS|81|1|psalmus Asaph Deus stetit in synagoga deorum in medio autem Deus deiudicat
PS|81|2|usquequo iudicatis iniquitatem et facies peccatorum sumitis diapsalma
PS|81|3|iudicate egenum et pupillum humilem et pauperem iustificate
PS|81|4|eripite pauperem et egenum de manu peccatoris liberate
PS|81|5|nescierunt neque intellexerunt in tenebris ambulant movebuntur omnia fundamenta terrae
PS|81|6|ego dixi dii estis et filii Excelsi omnes
PS|81|7|vos autem sicut homines moriemini et sicut unus de principibus cadetis
PS|81|8|surge Deus iudica terram quoniam tu hereditabis in omnibus gentibus
PS|82|1|canticum psalmi Asaph
PS|82|2|Deus quis similis erit tibi ne taceas neque conpescaris Deus
PS|82|3|quoniam ecce inimici tui sonaverunt et qui oderunt te extulerunt caput
PS|82|4|super populum tuum malignaverunt consilium et cogitaverunt adversus sanctos tuos
PS|82|5|dixerunt venite et disperdamus eos de gente et non memoretur nomen Israhel ultra
PS|82|6|quoniam cogitaverunt unianimiter simul adversum te testamentum disposuerunt
PS|82|7|tabernacula Idumeorum et Ismahelitae Moab et Aggareni
PS|82|8|Gebal et Ammon et Amalech alienigenae cum habitantibus Tyrum
PS|82|9|etenim Assur venit cum illis facti sunt in adiutorium filiis Loth diapsalma
PS|82|10|fac illis sicut Madiam et Sisarae sicut Iabin in torrente Cison
PS|82|11|disperierunt in Endor facti sunt ut stercus terrae
PS|82|12|pone principes eorum sicut Oreb et Zeb et Zebee et Salmana omnes principes eorum
PS|82|13|qui dixerunt hereditate possideamus sanctuarium Dei
PS|82|14|Deus meus pone illos ut rotam sicut stipulam ante faciem venti
PS|82|15|sicut ignis qui conburit silvam sicut flamma conburens montes
PS|82|16|ita persequeris illos in tempestate tua et in ira tua turbabis eos
PS|82|17|imple facies illorum ignominia et quaerent nomen tuum Domine
PS|82|18|erubescant et conturbentur in saeculum saeculi et confundantur et pereant
PS|82|19|et cognoscant quia nomen tibi Dominus tu solus Altissimus in omni terra
PS|83|1|in finem pro torcularibus filiis Core psalmus
PS|83|2|quam dilecta tabernacula tua Domine virtutum
PS|83|3|concupiscit et defecit anima mea in atria Domini cor meum et caro mea exultavit in Deum vivum
PS|83|4|etenim passer invenit %sibi; domum et turtur nidum sibi ubi ponat pullos suos altaria tua Domine virtutum rex meus et Deus meus
PS|83|5|beati qui habitant in domo tua in saecula saeculorum laudabunt te diapsalma
PS|83|6|beatus vir cui est auxilium abs te ascensiones in corde suo disposuit
PS|83|7|in valle lacrimarum in loco quem posuit
PS|83|8|etenim benedictiones dabit legis dator ibunt de virtute in virtutem videbitur Deus deorum in Sion
PS|83|9|Domine Deus virtutum exaudi orationem meam auribus percipe Deus Iacob diapsalma
PS|83|10|protector noster aspice Deus et respice in faciem christi tui
PS|83|11|quia melior est dies una in atriis tuis super milia elegi abiectus esse in domo Dei mei magis quam habitare in tabernaculis peccatorum
PS|83|12|quia misericordiam et veritatem %diligit; Deus gratiam et gloriam dabit Dominus
PS|83|13|non privabit bonis eos qui ambulant in innocentia Domine virtutum beatus vir qui sperat in te
PS|84|1|in finem filiis Core psalmus
PS|84|2|benedixisti Domine terram tuam avertisti captivitatem Iacob
PS|84|3|remisisti iniquitates plebis tuae operuisti omnia peccata eorum diapsalma
PS|84|4|mitigasti omnem iram tuam avertisti ab ira indignationis tuae
PS|84|5|converte nos Deus salutum nostrarum et averte iram tuam a nobis
PS|84|6|numquid in aeternum irasceris nobis aut extendes iram tuam a generatione in generationem
PS|84|7|Deus tu conversus vivificabis nos et plebs tua laetabitur in te
PS|84|8|ostende nobis Domine misericordiam tuam et salutare tuum da nobis
PS|84|9|audiam quid loquatur % in me; Dominus Deus quoniam loquetur pacem in plebem suam et super sanctos suos et in eos qui convertuntur ad cor
PS|84|10|verumtamen prope timentes eum salutare ipsius ut inhabitet gloria in terra nostra
PS|84|11|misericordia et veritas obviaverunt % sibi; iustitia et pax osculatae sunt
PS|84|12|veritas de terra orta est et iustitia de caelo prospexit
PS|84|13|etenim Dominus dabit benignitatem et terra nostra dabit fructum suum
PS|84|14|iustitia ante eum ambulabit et ponet in via gressus suos
PS|85|1|oratio ipsi David inclina Domine aurem tuam %et; exaudi me quoniam inops et pauper sum ego
PS|85|2|custodi animam meam quoniam sanctus sum salvum fac servum tuum Deus meus sperantem in te
PS|85|3|miserere mei Domine quoniam ad te clamabo tota die
PS|85|4|laetifica animam servi tui quoniam ad te Domine animam meam levavi
PS|85|5|quoniam tu Domine suavis et mitis et multae misericordiae omnibus invocantibus te
PS|85|6|auribus percipe Domine orationem meam et intende voci orationis meae
PS|85|7|in die tribulationis meae clamavi ad te quia exaudisti me
PS|85|8|non est similis tui in diis Domine et non est secundum opera tua
PS|85|9|omnes gentes quascumque fecisti venient et adorabunt coram te Domine et glorificabunt nomen tuum
PS|85|10|quoniam magnus es tu et faciens mirabilia tu es Deus solus
PS|85|11|deduc me Domine in via tua et ingrediar in veritate tua laetetur cor meum ut timeat nomen tuum
PS|85|12|confitebor tibi Domine Deus meus in toto corde meo et glorificabo nomen tuum in aeternum
PS|85|13|quia misericordia tua magna est super me et eruisti animam meam ex inferno inferiori
PS|85|14|Deus iniqui insurrexerunt super me et synagoga potentium quaesierunt animam meam et non proposuerunt te in conspectu suo
PS|85|15|et tu Domine Deus miserator et misericors patiens et multae misericordiae et verax
PS|85|16|respice in me et miserere mei da imperium tuum puero tuo et salvum fac filium ancillae tuae
PS|85|17|fac mecum signum in bono et videant qui oderunt me et confundantur quoniam tu Domine adiuvasti me et consolatus es me
PS|86|1|filiis Core psalmus cantici fundamenta eius in montibus sanctis
PS|86|2|diligit Dominus portas Sion super omnia tabernacula Iacob
PS|86|3|gloriosa dicta sunt de te civitas Dei diapsalma
PS|86|4|memor ero Raab et Babylonis scientibus me ecce alienigenae et Tyrus et populus Aethiopum hii fuerunt illic
PS|86|5|numquid Sion dicet homo et homo natus est in ea et ipse fundavit eam Altissimus
PS|86|6|Dominus narrabit in scriptura populorum et principum horum qui fuerunt in ea diapsalma
PS|86|7|sicut laetantium omnium habitatio in te
PS|87|1|canticum psalmi filiis Core in finem pro Maeleth ad respondendum intellectus Eman Ezraitae
PS|87|2|Domine Deus salutis meae die clamavi et nocte coram te
PS|87|3|intret in conspectu tuo oratio mea inclina aurem tuam ad precem meam
PS|87|4|quia repleta est malis anima mea et vita mea in inferno adpropinquavit
PS|87|5|aestimatus sum cum descendentibus in lacum factus sum sicut homo sine adiutorio
PS|87|6|inter mortuos liber sicut vulnerati dormientes in sepulchris quorum non es memor amplius et ipsi de manu tua repulsi sunt
PS|87|7|posuerunt me in lacu inferiori in tenebrosis et in umbra mortis
PS|87|8|super me confirmatus est furor tuus et omnes fluctus tuos induxisti super me diapsalma
PS|87|9|longe fecisti notos meos a me posuerunt me abominationem sibi traditus sum et non egrediebar
PS|87|10|oculi mei languerunt prae inopia clamavi ad te Domine tota die expandi ad te manus meas
PS|87|11|numquid mortuis facies mirabilia aut medici suscitabunt et confitebuntur tibi diapsalma
PS|87|12|numquid narrabit aliquis in sepulchro misericordiam tuam et veritatem tuam in perditione
PS|87|13|numquid cognoscentur in tenebris mirabilia tua et iustitia tua in terra oblivionis
PS|87|14|et ego ad te Domine clamavi et mane oratio mea praeveniet te
PS|87|15|ut quid Domine repellis orationem meam avertis faciem tuam a me
PS|87|16|pauper sum ego et in laboribus a iuventute mea exaltatus autem humiliatus sum et conturbatus
PS|87|17|in me transierunt irae tuae et terrores tui conturbaverunt me
PS|87|18|circuierunt me sicut aqua tota die circumdederunt me simul
PS|87|19|elongasti a me amicum et proximum et notos meos a miseria
PS|88|1|intellectus Aethan Ezraitae
PS|88|2|misericordias Domini in aeternum cantabo in generationem et generationem adnuntiabo veritatem tuam in ore meo
PS|88|3|quoniam dixisti in aeternum misericordia aedificabitur in caelis praeparabitur veritas tua in eis;
PS|88|4|disposui testamentum electis meis iuravi David servo meo
PS|88|5|usque in aeternum praeparabo semen tuum et aedificabo in generationem et generationem sedem tuam diapsalma
PS|88|6|confitebuntur caeli mirabilia tua Domine etenim veritatem tuam in ecclesia sanctorum
PS|88|7|quoniam quis in nubibus aequabitur Domino similis erit Domino in filiis Dei
PS|88|8|Deus qui glorificatur in consilio sanctorum magnus et horrendus super omnes qui in circuitu eius sunt
PS|88|9|Domine Deus virtutum quis similis tibi potens es Domine et veritas tua in circuitu tuo
PS|88|10|tu dominaris potestatis maris motum autem fluctuum eius tu mitigas
PS|88|11|tu humiliasti sicut vulneratum superbum in brachio virtutis tuae dispersisti inimicos tuos
PS|88|12|tui sunt caeli et tua est terra orbem terrae et plenitudinem eius tu fundasti
PS|88|13|aquilonem et mare tu creasti Thabor et Hermon in nomine tuo exultabunt
PS|88|14|tuum brachium cum potentia firmetur manus tua et exaltetur dextera tua
PS|88|15|iustitia et iudicium praeparatio sedis tuae misericordia et veritas praecedent faciem tuam
PS|88|16|beatus populus qui scit iubilationem Domine in lumine vultus tui ambulabunt
PS|88|17|et in nomine tuo exultabunt tota die et in iustitia tua exaltabuntur
PS|88|18|quoniam gloria virtutis eorum tu es et in beneplacito tuo exaltabitur cornu nostrum
PS|88|19|quia Domini est adsumptio nostra; et Sancti Israhel regis nostri
PS|88|20|tunc locutus es in visione sanctis tuis et dixisti posui adiutorium in potentem exaltavi electum de plebe mea
PS|88|21|inveni David servum meum in oleo sancto meo linui eum
PS|88|22|manus enim mea auxiliabitur ei et brachium meum confirmabit eum
PS|88|23|nihil proficiet inimicus in eo et filius iniquitatis non adponet nocere eum
PS|88|24|et concidam a facie ipsius inimicos eius et odientes eum in fugam convertam
PS|88|25|et veritas mea et misericordia mea cum ipso et in nomine meo exaltabitur cornu eius
PS|88|26|et ponam in mari manum eius et in fluminibus dexteram eius
PS|88|27|ipse invocabit me pater meus es tu Deus meus et susceptor salutis meae
PS|88|28|et ego primogenitum ponam illum excelsum prae regibus terrae
PS|88|29|in aeternum servabo illi misericordiam meam et testamentum meum fidele ipsi
PS|88|30|et ponam in saeculum saeculi semen eius et thronum eius sicut dies caeli
PS|88|31|si dereliquerint filii eius legem meam et in iudiciis meis non ambulaverint
PS|88|32|si iustitias meas profanaverint et mandata mea non custodierint
PS|88|33|visitabo in virga iniquitates eorum et in verberibus peccata eorum
PS|88|34|misericordiam autem meam non dispergam ab eo neque nocebo in veritate mea
PS|88|35|neque profanabo testamentum meum et quae procedunt de labiis meis non faciam irrita
PS|88|36|semel iuravi in sancto meo si David mentiar
PS|88|37|semen eius in aeternum manebit
PS|88|38|et thronus eius sicut sol in conspectu meo et sicut luna perfecta in aeternum et testis in caelo fidelis diapsalma
PS|88|39|tu vero reppulisti et despexisti distulisti christum tuum
PS|88|40|evertisti testamentum servi tui profanasti in terram sanctuarium eius
PS|88|41|destruxisti omnes sepes eius posuisti firmamenta eius formidinem
PS|88|42|diripuerunt eum omnes transeuntes viam factus est obprobrium vicinis suis
PS|88|43|exaltasti dexteram deprimentium eum laetificasti omnes inimicos eius
PS|88|44|avertisti adiutorium gladii eius et non es auxiliatus ei in bello
PS|88|45|destruxisti eum a mundatione sedem eius in terram conlisisti
PS|88|46|minorasti dies temporis eius perfudisti eum confusione diapsalma
PS|88|47|usquequo Domine avertis in finem exardescet sicut ignis ira tua
PS|88|48|memorare quae mea substantia numquid enim vane constituisti omnes filios hominum
PS|88|49|quis est homo qui vivet et non videbit mortem eruet animam suam de manu inferi diapsalma
PS|88|50|ubi sunt misericordiae tuae antiquae Domine sicut iurasti David in veritate tua
PS|88|51|memor esto Domine obprobrii servorum tuorum quod continui in sinu meo multarum gentium
PS|88|52|quod exprobraverunt inimici tui Domine quod exprobraverunt commutationem christi tui
PS|88|53|benedictus Dominus in aeternum fiat fiat
PS|89|1|oratio Mosi hominis Dei Domine refugium tu factus es nobis in generatione et generatione
PS|89|2|priusquam montes fierent et formaretur terra et orbis a saeculo usque in saeculum tu es Deus
PS|89|3|ne avertas hominem in humilitatem et dixisti convertimini filii hominum
PS|89|4|quoniam mille anni ante oculos tuos tamquam dies hesterna quae praeteriit et custodia in nocte
PS|89|5|quae pro nihilo habentur eorum anni erunt
PS|89|6|mane sicut herba transeat mane floreat et transeat vespere decidat induret et arescat
PS|89|7|quia defecimus in ira tua et in furore tuo turbati sumus
PS|89|8|posuisti iniquitates nostras in conspectu tuo saeculum nostrum in inluminatione vultus tui
PS|89|9|quoniam omnes dies nostri defecerunt in ira tua defecimus anni nostri sicut aranea meditabantur
PS|89|10|dies annorum nostrorum in ipsis septuaginta anni si autem in potentatibus octoginta anni et amplius eorum labor et dolor quoniam supervenit mansuetudo et corripiemur
PS|89|11|quis novit potestatem irae tuae et prae timore tuo iram tuam
PS|89|12|dinumerare dexteram tuam sic notam fac et conpeditos corde in sapientia
PS|89|13|convertere Domine usquequo et deprecabilis esto super servos tuos
PS|89|14|repleti sumus mane misericordia tua et exultavimus et delectati sumus in omnibus diebus nostris
PS|89|15|laetati sumus pro diebus quibus nos humiliasti annis quibus vidimus mala
PS|89|16|et respice in servos tuos et in opera tua et dirige filios eorum
PS|89|17|et sit splendor Domini Dei nostri super nos et opera manuum nostrarum dirige super nos et opus manuum nostrarum dirige;
PS|90|1|laus cantici David qui habitat in adiutorio Altissimi in protectione Dei caeli commorabitur
PS|90|2|dicet Domino susceptor meus es tu et refugium meum Deus meus sperabo in eum
PS|90|3|quoniam ipse liberabit me de laqueo venantium et a verbo aspero
PS|90|4|in scapulis suis obumbrabit te et sub pinnis eius sperabis
PS|90|5|scuto circumdabit te veritas eius non timebis a timore nocturno
PS|90|6|a sagitta volante in die a negotio perambulante in tenebris ab incursu et daemonio meridiano
PS|90|7|cadent a latere tuo mille et decem milia a dextris tuis ad te autem non adpropinquabit
PS|90|8|verumtamen oculis tuis considerabis et retributionem peccatorum videbis
PS|90|9|quoniam tu Domine spes mea Altissimum posuisti refugium tuum
PS|90|10|non accedent ad te mala et flagellum non adpropinquabit tabernaculo tuo
PS|90|11|quoniam angelis suis mandabit de te ut custodiant te in omnibus viis tuis
PS|90|12|in manibus portabunt te ne forte offendas ad lapidem pedem tuum
PS|90|13|super aspidem et basiliscum ambulabis %et; conculcabis leonem et draconem
PS|90|14|quoniam in me speravit et liberabo eum protegam eum quia cognovit nomen meum
PS|90|15|clamabit ad me et exaudiam eum cum ipso sum in tribulatione eripiam eum et clarificabo eum
PS|90|16|longitudine dierum replebo eum et ostendam illi salutare meum
PS|91|1|psalmus cantici in die sabbati
PS|91|2|bonum est confiteri Domino et psallere nomini tuo Altissime
PS|91|3|ad adnuntiandum mane misericordiam tuam et veritatem tuam per noctem
PS|91|4|in decacordo psalterio cum cantico in cithara
PS|91|5|quia delectasti me Domine in factura tua et in operibus manuum tuarum exultabo
PS|91|6|quam magnificata sunt opera tua Domine nimis profundae factae sunt cogitationes tuae
PS|91|7|vir insipiens non cognoscet et stultus non intelleget haec
PS|91|8|cum exorti fuerint peccatores sicut faenum et apparuerint omnes qui operantur iniquitatem ut intereant in saeculum %saeculi;
PS|91|9|tu autem Altissimus in aeternum Domine
PS|91|10|quoniam ecce inimici tui Domine; quoniam ecce inimici tui peribunt et dispergentur omnes qui operantur iniquitatem
PS|91|11|et exaltabitur sicut unicornis cornu meum et senectus mea in misericordia uberi
PS|91|12|et despexit oculus meus inimicis meis et insurgentibus in me malignantibus audiet auris mea
PS|91|13|iustus ut palma florebit ut cedrus Libani multiplicabitur
PS|91|14|plantati in domo Domini in atriis Dei nostri florebunt
PS|91|15|adhuc multiplicabuntur in senecta uberi et bene patientes erunt
PS|91|16|ut adnuntient quoniam rectus Dominus Deus noster et non est iniquitas in eo
PS|92|1|laus cantici David in die ante sabbatum quando inhabitata est terra Dominus regnavit decore indutus est indutus est Dominus fortitudine et praecinxit se etenim firmavit orbem terrae qui non commovebitur
PS|92|2|parata sedis tua ex tunc a saeculo tu es
PS|92|3|elevaverunt flumina Domine elevaverunt flumina vocem suam elevabunt flumina fluctus suos;
PS|92|4|a vocibus aquarum multarum mirabiles elationes maris mirabilis in altis Dominus
PS|92|5|testimonia tua credibilia facta sunt nimis domum tuam decet sanctitudo Domine in longitudine dierum
PS|93|1|psalmus David quarta sabbati Deus ultionum Dominus Deus ultionum libere egit
PS|93|2|exaltare qui iudicas terram redde retributionem superbis
PS|93|3|usquequo peccatores Domine usquequo peccatores gloriabuntur
PS|93|4|effabuntur et loquentur iniquitatem loquentur omnes qui operantur iniustitiam
PS|93|5|populum tuum Domine humiliaverunt et hereditatem tuam vexaverunt
PS|93|6|viduam et advenam interfecerunt et pupillos occiderunt
PS|93|7|et dixerunt non videbit Dominus nec intelleget Deus Iacob
PS|93|8|intellegite qui insipientes estis in populo et stulti aliquando sapite
PS|93|9|qui plantavit aurem non audiet aut qui finxit oculum non considerat
PS|93|10|qui corripit gentes non arguet qui docet hominem scientiam
PS|93|11|Dominus scit cogitationes hominum quoniam vanae sunt
PS|93|12|beatus homo quem tu erudieris Domine et de lege tua docueris eum
PS|93|13|ut mitiges ei a diebus malis donec fodiatur peccatori fovea
PS|93|14|quia non repellet Dominus plebem suam et hereditatem suam non derelinquet
PS|93|15|quoadusque iustitia convertatur in iudicium et qui iuxta illam omnes qui recto sunt corde diapsalma
PS|93|16|quis consurget mihi adversus malignantes aut quis stabit mecum adversus operantes iniquitatem
PS|93|17|nisi quia Dominus adiuvit me paulo minus habitavit in inferno anima mea
PS|93|18|si dicebam motus est pes meus misericordia tua Domine adiuvabat me
PS|93|19|secundum multitudinem dolorum meorum in corde meo consolationes tuae laetificaverunt animam meam
PS|93|20|numquid aderit tibi sedis iniquitatis qui fingis dolorem in praecepto
PS|93|21|captabunt in animam iusti et sanguinem innocentem condemnabunt
PS|93|22|et factus est Dominus mihi in refugium et Deus meus in adiutorem spei meae
PS|93|23|et reddet illis iniquitatem ipsorum et in malitia eorum disperdet eos disperdet illos Dominus Deus noster
PS|94|1|laus cantici David venite exultemus Domino iubilemus Deo salutari nostro
PS|94|2|praeoccupemus faciem eius in confessione et in psalmis iubilemus ei
PS|94|3|quoniam Deus magnus Dominus et rex magnus super omnes deos
PS|94|4|quia in manu eius fines terrae et altitudines montium ipsius sunt
PS|94|5|quoniam ipsius est mare et ipse fecit illud et siccam manus eius formaverunt
PS|94|6|venite adoremus et procidamus et ploremus ante Dominum qui fecit nos
PS|94|7|quia ipse est Deus noster et nos populus pascuae eius et oves manus eius
PS|94|8|hodie si vocem eius audieritis nolite obdurare corda vestra
PS|94|9|sicut in inritatione secundum diem temptationis in deserto ubi temptaverunt me patres vestri probaverunt me; et viderunt opera mea
PS|94|10|quadraginta annis offensus fui generationi illi et dixi semper errant corde
PS|94|11|et isti non cognoverunt vias meas ut iuravi in ira mea si intrabunt in requiem meam
PS|95|1|quando domus aedificabatur post captivitatem canticum huic David cantate Domino canticum novum cantate Domino omnis terra
PS|95|2|cantate Domino benedicite nomini eius adnuntiate diem de die salutare eius
PS|95|3|adnuntiate inter gentes gloriam eius in omnibus populis mirabilia eius
PS|95|4|quoniam magnus Dominus et laudabilis valde terribilis est super omnes deos
PS|95|5|quoniam omnes dii gentium daemonia at vero Dominus caelos fecit
PS|95|6|confessio et pulchritudo in conspectu eius sanctimonia et magnificentia in sanctificatione eius
PS|95|7|adferte Domino patriae gentium adferte Domino gloriam et honorem
PS|95|8|adferte Domino gloriam nomini eius tollite hostias et introite in atria eius
PS|95|9|adorate Dominum in atrio sancto eius commoveatur a facie eius universa terra
PS|95|10|dicite in gentibus quia Dominus regnavit etenim correxit orbem qui non movebitur iudicabit populos in aequitate
PS|95|11|laetentur caeli et exultet terra commoveatur mare et plenitudo eius
PS|95|12|gaudebunt campi et omnia quae in eis sunt tunc exultabunt omnia ligna silvarum
PS|95|13|a facie Domini quia venit quoniam venit iudicare terram iudicabit orbem terrae in aequitate et populos in veritate sua
PS|96|1|huic David quando terra eius restituta est Dominus regnavit exultet terra laetentur insulae multae
PS|96|2|nubes et caligo in circuitu eius iustitia et iudicium correctio sedis eius
PS|96|3|ignis ante ipsum praecedet et inflammabit in circuitu inimicos eius
PS|96|4|adluxerunt fulgora eius orbi terrae vidit et commota est terra
PS|96|5|montes sicut cera fluxerunt a facie Domini; a facie Domini omnis terrae
PS|96|6|adnuntiaverunt caeli iustitiam eius et viderunt omnes populi gloriam eius
PS|96|7|confundantur omnes qui adorant sculptilia qui gloriantur in simulacris suis adorate eum omnes angeli eius
PS|96|8|audivit et laetata est Sion et exultaverunt filiae Iudaeae propter iudicia tua Domine
PS|96|9|quoniam tu Dominus Altissimus super omnem terram nimis superexaltatus es super omnes deos
PS|96|10|qui diligitis Dominum odite malum custodit animas sanctorum suorum de manu peccatoris liberabit eos
PS|96|11|lux orta est iusto et rectis corde laetitia
PS|96|12|laetamini iusti in Domino et confitemini memoriae sanctificationis eius
PS|97|1|psalmus David cantate Domino canticum novum quoniam mirabilia fecit salvavit sibi dextera eius et brachium sanctum eius
PS|97|2|notum fecit Dominus salutare suum in conspectu gentium revelavit iustitiam suam
PS|97|3|recordatus est misericordiae suae et veritatem suam domui Israhel viderunt omnes termini terrae salutare Dei nostri
PS|97|4|iubilate Domino omnis terra cantate et exultate et psallite
PS|97|5|psallite Domino in cithara in cithara et voce psalmi
PS|97|6|in tubis ductilibus et voce tubae corneae iubilate in conspectu regis Domini
PS|97|7|moveatur mare et plenitudo eius orbis terrarum et qui habitant in eo
PS|97|8|flumina plaudent manu simul montes exultabunt
PS|97|9|a conspectu Domini quoniam venit iudicare terram iudicabit orbem terrarum in iustitia et populos in aequitate
PS|98|1|psalmus David Dominus regnavit irascantur populi qui sedet super cherubin moveatur terra
PS|98|2|Dominus in Sion magnus et excelsus est super omnes populos
PS|98|3|confiteantur nomini tuo magno quoniam terribile et sanctum est
PS|98|4|et honor regis iudicium diligit tu parasti directiones iudicium et iustitiam in Iacob tu fecisti
PS|98|5|exaltate Dominum Deum nostrum et adorate scabillum pedum eius quoniam sanctum est
PS|98|6|Moses et Aaron in sacerdotibus eius et Samuhel inter eos qui invocant nomen eius invocabant Dominum et ipse exaudiebat illos
PS|98|7|in columna nubis loquebatur ad eos custodiebant testimonia eius et praeceptum quod dedit illis
PS|98|8|Domine Deus noster tu exaudiebas illos Deus tu propitius fuisti eis et ulciscens in omnes adinventiones eorum
PS|98|9|exaltate Dominum Deum nostrum et adorate in monte sancto eius quoniam sanctus Dominus Deus noster
PS|99|1|psalmus in confessione
PS|99|2|iubilate Domino omnis terra servite Domino in laetitia introite in conspectu eius in exultatione
PS|99|3|scitote quoniam Dominus ipse est Deus ipse fecit nos et non ipsi nos populus eius et oves pascuae eius
PS|99|4|introite portas eius in confessione atria eius in hymnis confitemini illi laudate nomen eius
PS|99|5|quoniam suavis Dominus in aeternum misericordia eius et usque in generationem et generationem veritas eius
PS|100|1|David psalmus misericordiam et iudicium cantabo tibi Domine psallam
PS|100|2|et intellegam in via inmaculata quando venies ad me perambulabam in innocentia cordis mei in medio domus meae
PS|100|3|non proponebam ante oculos meos rem iniustam facientes praevaricationes odivi non adhesit mihi
PS|100|4|cor pravum declinante a me maligno non cognoscebam
PS|100|5|detrahentem secreto proximo suo hunc persequebar superbo oculo et insatiabili corde cum hoc non edebam
PS|100|6|oculi mei ad fideles terrae ut sederent mecum ambulans in via inmaculata hic mihi ministrabat
PS|100|7|non habitabat in medio domus meae qui facit superbiam qui loquitur iniqua non direxit in conspectu oculorum meorum
PS|100|8|in matutino interficiebam omnes peccatores terrae ut disperderem de civitate Domini omnes operantes iniquitatem
PS|101|1|oratio pauperis cum anxius fuerit et coram Domino effuderit precem suam
PS|101|2|Domine exaudi orationem meam et clamor meus ad te veniat
PS|101|3|non avertas faciem tuam a me in quacumque die tribulor inclina ad me aurem tuam in quacumque die invocavero te velociter exaudi me
PS|101|4|quia defecerunt sicut fumus dies mei et ossa mea sicut gremium aruerunt
PS|101|5|percussum est ut faenum et aruit cor meum quia oblitus sum comedere panem meum
PS|101|6|a voce gemitus mei adhesit os meum carni meae
PS|101|7|similis factus sum pelicano solitudinis factus sum sicut nycticorax in domicilio
PS|101|8|vigilavi et factus sum sicut passer solitarius in tecto
PS|101|9|tota die exprobrabant mihi inimici mei et qui laudabant me adversus me iurabant
PS|101|10|quia cinerem tamquam panem manducavi et poculum meum cum fletu miscebam
PS|101|11|a facie irae et indignationis tuae quia elevans adlisisti me
PS|101|12|dies mei sicut umbra declinaverunt et ego sicut faenum arui
PS|101|13|tu autem Domine in aeternum permanes et memoriale tuum in generationem et generationem
PS|101|14|tu exsurgens misereberis Sion quia tempus miserendi eius quia venit tempus
PS|101|15|quoniam placuerunt servis tuis lapides eius et terrae eius miserebuntur
PS|101|16|et timebunt gentes nomen Domini et omnes reges terrae gloriam tuam
PS|101|17|quia aedificabit Dominus Sion et videbitur in gloria sua
PS|101|18|respexit in orationem humilium et non sprevit precem eorum
PS|101|19|scribantur haec in generationem alteram et populus qui creabitur laudabit Dominum
PS|101|20|quia prospexit de excelso sancto suo Dominus de caelo in terram aspexit
PS|101|21|ut audiret gemitum conpeditorum ut solvat filios interemptorum
PS|101|22|ut adnuntiet in Sion nomen Domini et laudem suam in Hierusalem
PS|101|23|in conveniendo populos in unum et reges ut serviant Domino
PS|101|24|respondit ei in via virtutis suae paucitatem dierum meorum nuntia mihi
PS|101|25|ne revoces me in dimidio dierum meorum in generationem et generationem anni tui
PS|101|26|initio tu Domine terram fundasti et opera manuum tuarum sunt caeli
PS|101|27|ipsi peribunt tu autem permanes et omnes sicut vestimentum veterescent et sicut opertorium mutabis eos et mutabuntur
PS|101|28|tu autem idem ipse es et anni tui non deficient
PS|101|29|filii servorum tuorum habitabunt et semen eorum in saeculum dirigetur
PS|102|1|ipsi David benedic anima mea Domino et omnia quae intra me sunt nomini sancto eius
PS|102|2|benedic anima mea Domino et noli oblivisci omnes retributiones eius
PS|102|3|qui propitiatur omnibus iniquitatibus tuis qui sanat omnes infirmitates tuas
PS|102|4|qui redimit de interitu vitam tuam qui coronat te in misericordia et miserationibus
PS|102|5|qui replet in bonis desiderium tuum renovabitur ut aquilae iuventus tua
PS|102|6|faciens misericordias Dominus et iudicium omnibus iniuriam patientibus
PS|102|7|notas fecit vias suas Mosi filiis Israhel voluntates suas
PS|102|8|miserator et misericors Dominus longanimis et multum misericors
PS|102|9|non in perpetuum irascetur neque in aeternum comminabitur
PS|102|10|non secundum peccata nostra fecit nobis nec secundum iniustitias nostras retribuit nobis
PS|102|11|quoniam secundum altitudinem caeli a terra corroboravit misericordiam suam super timentes se
PS|102|12|quantum distat ortus ab occidente longe fecit a nobis iniquitates nostras
PS|102|13|quomodo miseretur pater filiorum misertus est Dominus timentibus se
PS|102|14|quoniam ipse cognovit figmentum nostrum recordatus est quoniam pulvis sumus
PS|102|15|homo sicut faenum dies eius tamquam flos agri sic efflorebit
PS|102|16|quoniam spiritus pertransivit in illo et non subsistet et non cognoscet amplius locum suum
PS|102|17|misericordia autem Domini ab aeterno et usque in aeternum super timentes eum et iustitia illius in filios filiorum
PS|102|18|his qui servant testamentum eius et memores sunt mandatorum ipsius ad faciendum ea
PS|102|19|Dominus in caelo paravit sedem suam et regnum ipsius omnibus dominabitur
PS|102|20|benedicite Domino angeli eius potentes virtute facientes verbum illius ad audiendam vocem sermonum eius
PS|102|21|benedicite Domino omnes virtutes eius ministri eius qui facitis voluntatem eius
PS|102|22|benedicite Domino omnia opera eius in omni loco dominationis ipsius benedic anima mea Domino
PS|103|1|ipsi David benedic anima mea Domino Domine Deus meus magnificatus es vehementer confessionem et decorem induisti
PS|103|2|amictus lumine sicut vestimento extendens caelum sicut pellem
PS|103|3|qui tegis in aquis superiora eius qui ponis nubem ascensum tuum qui ambulas super pinnas ventorum
PS|103|4|qui facis angelos tuos spiritus et ministros tuos ignem urentem
PS|103|5|qui fundasti terram super stabilitatem suam non inclinabitur in saeculum saeculi
PS|103|6|abyssus sicut vestimentum amictus eius super montes stabunt aquae
PS|103|7|ab increpatione tua fugient a voce tonitrui tui formidabunt
PS|103|8|ascendunt montes et descendunt campi in locum quem fundasti eis
PS|103|9|terminum posuisti quem non transgredientur neque convertentur operire terram
PS|103|10|qui emittis fontes in convallibus inter medium montium pertransibunt aquae
PS|103|11|potabunt omnes bestiae agri expectabunt onagri in siti sua
PS|103|12|super ea volucres caeli habitabunt de medio petrarum dabunt vocem
PS|103|13|rigans montes de superioribus suis de fructu operum tuorum satiabitur terra
PS|103|14|producens faenum iumentis et herbam servituti hominum ut educas panem de terra
PS|103|15|et vinum laetificat cor hominis ut exhilaret faciem in oleo et panis cor hominis confirmat
PS|103|16|saturabuntur ligna campi et cedri Libani quas plantavit
PS|103|17|illic passeres nidificabunt erodii domus dux est eorum
PS|103|18|montes excelsi cervis petra refugium erinaciis
PS|103|19|fecit lunam in tempora sol cognovit occasum suum
PS|103|20|posuisti tenebras et facta est nox in ipsa pertransibunt omnes bestiae silvae
PS|103|21|catuli leonum rugientes ut rapiant et quaerant a Deo escam sibi
PS|103|22|ortus est sol et congregati sunt et in cubilibus suis conlocabuntur
PS|103|23|exibit homo ad opus suum et ad operationem suam usque ad vesperum
PS|103|24|quam magnificata sunt opera tua Domine omnia in sapientia fecisti impleta est terra possessione tua
PS|103|25|hoc mare magnum et spatiosum manibus; illic reptilia quorum non est numerus animalia pusilla cum magnis
PS|103|26|illic naves pertransibunt draco iste quem formasti ad inludendum ei
PS|103|27|omnia a te expectant ut des illis escam in tempore
PS|103|28|dante te illis colligent aperiente te manum tuam omnia implebuntur bonitate
PS|103|29|avertente autem te faciem turbabuntur auferes spiritum eorum et deficient et in pulverem suum revertentur
PS|103|30|emittes spiritum tuum et creabuntur et renovabis faciem terrae
PS|103|31|sit gloria Domini in saeculum laetabitur Dominus in operibus suis
PS|103|32|qui respicit terram et facit eam tremere qui tangit montes et fumigant
PS|103|33|cantabo Domino in vita mea psallam Deo meo quamdiu sum
PS|103|34|iucundum sit ei eloquium meum ego vero delectabor in Domino
PS|103|35|deficiant peccatores a terra et iniqui ita ut non sint benedic anima mea Domino
PS|104|1|alleluia confitemini Domino et invocate nomen eius adnuntiate inter gentes opera eius
PS|104|2|cantate ei et psallite ei narrate omnia mirabilia eius
PS|104|3|laudamini in nomine sancto eius laetetur cor quaerentium Dominum
PS|104|4|quaerite Dominum et confirmamini quaerite faciem eius semper
PS|104|5|mementote mirabilium eius quae fecit prodigia eius et iudicia oris eius
PS|104|6|semen Abraham servi eius filii Iacob electi eius
PS|104|7|ipse Dominus Deus noster in universa terra iudicia eius
PS|104|8|memor fuit in saeculum testamenti sui verbi quod mandavit in mille generationes
PS|104|9|quod disposuit ad Abraham et iuramenti sui ad Isaac
PS|104|10|et statuit illud Iacob in praeceptum et Israhel in testamentum aeternum
PS|104|11|dicens tibi dabo terram Chanaan funiculum hereditatis vestrae
PS|104|12|cum essent numero breves paucissimos et incolas eius
PS|104|13|et pertransierunt de gente in gentem et de regno ad populum alterum
PS|104|14|non reliquit hominem nocere eis et corripuit pro eis reges
PS|104|15|nolite tangere christos meos et in prophetis meis nolite malignari
PS|104|16|et vocavit famem super terram omne firmamentum panis contrivit
PS|104|17|misit ante eos virum in servum venundatus est Ioseph
PS|104|18|humiliaverunt in conpedibus pedes eius ferrum pertransiit anima eius
PS|104|19|donec veniret verbum eius eloquium Domini inflammavit eum
PS|104|20|misit rex et solvit eum princeps populorum et dimisit eum
PS|104|21|constituit eum dominum domus suae et principem omnis possessionis suae
PS|104|22|ut erudiret principes eius sicut semet ipsum et senes eius prudentiam doceret
PS|104|23|et intravit Israhel in Aegyptum et Iacob accola fuit in terra Cham
PS|104|24|et auxit populum eius vehementer et firmavit eum super inimicos eius
PS|104|25|convertit cor eorum ut odirent populum eius ut dolum facerent in servos eius
PS|104|26|misit Mosen servum suum Aaron quem elegit ipsum
PS|104|27|posuit in eis verba signorum suorum et prodigiorum in terra Cham
PS|104|28|misit tenebras et obscuravit et non exacerbavit sermones suos
PS|104|29|convertit aquas eorum in sanguinem et occidit pisces eorum
PS|104|30|dedit terra eorum ranas in penetrabilibus regum ipsorum
PS|104|31|dixit et venit cynomia et scinifes in omnibus finibus eorum
PS|104|32|posuit pluvias eorum grandinem ignem conburentem in terra ipsorum
PS|104|33|et percussit vineas eorum et ficulneas eorum et contrivit lignum finium eorum
PS|104|34|dixit et venit lucusta et bruchus cuius non erat numerus
PS|104|35|et comedit omne faenum in terra eorum et comedit omnem fructum terrae eorum
PS|104|36|et percussit omne primogenitum in terra eorum primitias omnis laboris eorum
PS|104|37|et eduxit eos in argento et auro et non erat in tribubus eorum infirmus
PS|104|38|laetata est Aegyptus in profectione eorum quia incubuit timor eorum super eos
PS|104|39|expandit nubem in protectionem eorum et ignem ut luceret eis per noctem
PS|104|40|petierunt et venit coturnix et panem caeli saturavit eos
PS|104|41|disrupit petram et fluxerunt aquae abierunt in sicco flumina
PS|104|42|quoniam memor fuit verbi sancti sui quod habuit ad Abraham puerum suum
PS|104|43|et eduxit populum suum in exultatione %et; electos suos in laetitia
PS|104|44|et dedit illis regiones gentium et labores populorum possederunt
PS|104|45|ut custodiant iustificationes eius et legem eius requirant
PS|105|1|alleluia confitemini Domino quoniam bonus quoniam in saeculum misericordia eius
PS|105|2|quis loquetur potentias Domini auditas faciet omnes laudes eius
PS|105|3|beati qui custodiunt iudicium et faciunt iustitiam in omni tempore
PS|105|4|memento nostri Domine in beneplacito populi tui visita nos in salutari tuo
PS|105|5|ad videndum in bonitate electorum tuorum ad laetandum in laetitia gentis tuae et lauderis cum hereditate tua
PS|105|6|peccavimus cum patribus nostris iniuste egimus iniquitatem fecimus
PS|105|7|patres nostri in Aegypto non intellexerunt mirabilia tua non fuerunt memores multitudinis misericordiae tuae et inritaverunt ascendentes in mare mare; Rubrum
PS|105|8|et salvavit eos propter nomen suum ut notam faceret potentiam suam
PS|105|9|et increpuit mare Rubrum et exsiccatum est et deduxit eos in abyssis sicut in deserto
PS|105|10|et salvavit eos de manu odientium et redemit eos de manu inimici
PS|105|11|et operuit aqua tribulantes eos unus ex eis non remansit
PS|105|12|et crediderunt in verbis eius et laudaverunt laudem eius
PS|105|13|cito fecerunt obliti sunt operum eius non sustinuerunt consilium eius
PS|105|14|et concupierunt concupiscentiam in deserto et temptaverunt Deum in inaquoso
PS|105|15|et dedit eis petitionem ipsorum et misit saturitatem in anima eorum
PS|105|16|et inritaverunt Mosen in castris Aaron sanctum Domini
PS|105|17|aperta est terra et degluttivit Dathan et operuit super congregationem Abiron
PS|105|18|et exarsit ignis in synagoga eorum flamma conbusit peccatores
PS|105|19|et fecerunt vitulum in Choreb et adoraverunt sculptile
PS|105|20|et mutaverunt gloriam suam in similitudine vituli comedentis faenum
PS|105|21|obliti sunt Deum qui salvavit eos qui fecit magnalia in Aegypto
PS|105|22|mirabilia in terra Cham terribilia in mari Rubro
PS|105|23|et dixit ut disperderet eos si non Moses electus eius stetisset in confractione in conspectu eius ut averteret iram eius ne disperderet eos
PS|105|24|et pro nihilo habuerunt terram desiderabilem non crediderunt verbo eius
PS|105|25|et murmurabant in tabernaculis suis non exaudierunt vocem Domini
PS|105|26|et elevavit manum suam super eos ut prosterneret eos in deserto
PS|105|27|et ut deiceret semen eorum in nationibus et dispergeret eos in regionibus
PS|105|28|et initiati sunt Beelphegor et comederunt sacrificia mortuorum
PS|105|29|et inritaverunt eum in adinventionibus suis et multiplicata est in eis ruina
PS|105|30|et stetit Finees et placavit et cessavit quassatio
PS|105|31|et reputatum est ei in iustitiam in generatione et generationem usque in sempiternum
PS|105|32|et inritaverunt ad aquam Contradictionis et vexatus est Moses propter eos
PS|105|33|quia exacerbaverunt spiritum eius et distinxit in labiis suis
PS|105|34|non disperdiderunt gentes quas dixit Dominus illis
PS|105|35|et commixti sunt inter gentes et didicerunt opera eorum
PS|105|36|et servierunt sculptilibus eorum et factum est illis in scandalum
PS|105|37|et immolaverunt filios suos et filias suas daemoniis
PS|105|38|et effuderunt sanguinem innocentem sanguinem filiorum suorum et filiarum suarum; quas sacrificaverunt sculptilibus Chanaan et interfecta est terra in sanguinibus
PS|105|39|et contaminata est in operibus eorum et fornicati sunt in adinventionibus suis
PS|105|40|et iratus est furore Dominus in populo suo et abominatus est hereditatem suam
PS|105|41|et tradidit eos in manus gentium et dominati sunt eorum qui oderant eos
PS|105|42|et tribulaverunt eos inimici eorum et humiliati sunt sub manibus eorum
PS|105|43|saepe liberavit eos ipsi autem exacerbaverunt eum in consilio suo et humiliati sunt in iniquitatibus suis
PS|105|44|et vidit cum tribularentur et audiret orationem eorum
PS|105|45|et memor fuit testamenti sui et paenituit eum secundum multitudinem misericordiae suae
PS|105|46|et dedit eos in misericordias in conspectu omnium qui ceperant eos
PS|105|47|salvos fac nos Domine Deus noster et congrega nos de nationibus ut confiteamur nomini tuo sancto et gloriemur in laude tua
PS|105|48|benedictus Dominus Deus Israhel a saeculo et usque in saeculum et dicet omnis populus fiat fiat
PS|106|1|alleluia confitemini Domino quoniam bonus quoniam in saeculum misericordia eius
PS|106|2|dicant qui redempti sunt a Domino quos redemit de manu inimici de regionibus congregavit eos
PS|106|3|a solis ortu et occasu et ab aquilone et mari
PS|106|4|erraverunt in solitudine in inaquoso viam civitatis habitaculi non invenerunt
PS|106|5|esurientes et sitientes anima eorum in ipsis defecit
PS|106|6|et clamaverunt ad Dominum cum tribularentur et de necessitatibus eorum eripuit eos
PS|106|7|et deduxit eos in viam rectam ut irent in civitatem habitationis
PS|106|8|confiteantur Domino misericordiae eius et mirabilia eius filiis hominum
PS|106|9|quia satiavit animam inanem et animam esurientem satiavit bonis
PS|106|10|sedentes in tenebris et umbra mortis vinctos in mendicitate et ferro
PS|106|11|quia exacerbaverunt eloquia Dei et consilium Altissimi inritaverunt
PS|106|12|et humiliatum est in laboribus cor eorum infirmati sunt nec fuit qui adiuvaret
PS|106|13|et clamaverunt ad Dominum cum tribularentur et de necessitatibus eorum liberavit eos
PS|106|14|et eduxit eos de tenebris et umbra mortis et vincula eorum disrupit
PS|106|15|confiteantur Domino misericordiae eius et mirabilia eius filiis hominum
PS|106|16|quia contrivit portas aereas et vectes ferreos confregit
PS|106|17|suscepit eos de via iniquitatis eorum propter iniustitias enim suas humiliati sunt
PS|106|18|omnem escam abominata est anima eorum et adpropinquaverunt usque ad portas mortis
PS|106|19|et clamaverunt ad Dominum cum tribularentur et de necessitatibus eorum liberavit eos
PS|106|20|misit verbum suum et sanavit eos et eripuit eos de interitionibus eorum
PS|106|21|confiteantur Domino misericordiae eius et mirabilia eius filiis hominum
PS|106|22|et sacrificent sacrificium laudis et adnuntient opera eius in exultatione
PS|106|23|qui descendunt mare in navibus facientes operationem in aquis multis
PS|106|24|ipsi viderunt opera Domini et mirabilia eius in profundo
PS|106|25|dixit et stetit spiritus procellae et exaltati sunt fluctus eius
PS|106|26|ascendunt usque ad caelos et descendunt usque ad abyssos anima eorum in malis tabescebat
PS|106|27|turbati sunt et moti sunt sicut ebrius et omnis sapientia eorum devorata est
PS|106|28|et clamaverunt ad Dominum cum tribularentur et de necessitatibus eorum eduxit eos
PS|106|29|et statuit procellam %eius; in auram et siluerunt fluctus eius
PS|106|30|et laetati sunt quia siluerunt et deduxit eos in portum voluntatis eorum
PS|106|31|confiteantur Domino misericordiae eius et mirabilia eius filiis hominum
PS|106|32|exaltent eum in ecclesia plebis et in cathedra seniorum laudent eum
PS|106|33|posuit flumina in desertum et exitus aquarum in sitim
PS|106|34|terram fructiferam in salsuginem a malitia inhabitantium in ea
PS|106|35|posuit desertum in stagna aquarum et terram sine aqua in exitus aquarum
PS|106|36|et conlocavit illic esurientes et constituerunt civitatem habitationis
PS|106|37|et seminaverunt agros et plantaverunt vineas et fecerunt fructum nativitatis
PS|106|38|et benedixit eis et multiplicati sunt nimis et iumenta eorum non minoravit
PS|106|39|et pauci facti sunt et vexati sunt a tribulatione malorum et dolore
PS|106|40|effusa est contemptio super principes et errare fecit eos in invio et non in via
PS|106|41|et adiuvit pauperem de inopia et posuit sicut oves familias
PS|106|42|videbunt recti et laetabuntur et omnis iniquitas oppilabit os suum
PS|106|43|quis sapiens et custodiet haec et intellegent misericordias Domini
PS|107|1|canticum psalmi David
PS|107|2|paratum cor meum Deus paratum cor meum cantabo et psallam in gloria mea
PS|107|3|exsurge psalterium et cithara exsurgam diluculo
PS|107|4|confitebor tibi in populis Domine et psallam tibi in nationibus
PS|107|5|quia magna super caelos misericordia tua et usque ad nubes veritas tua
PS|107|6|exaltare super caelos Deus et super omnem terram gloria tua
PS|107|7|ut liberentur dilecti tui salvum fac dextera tua et exaudi me
PS|107|8|Deus locutus est in sancto suo exaltabor et dividam Sicima et convallem tabernaculorum dimetiar
PS|107|9|meus est Galaad et meus est Manasse et Effraim susceptio capitis mei Iuda rex meus
PS|107|10|Moab lebes spei meae in Idumeam extendam calciamentum meum mihi alienigenae amici facti sunt
PS|107|11|quis deducet me in civitatem munitam quis deducet me usque in Idumeam
PS|107|12|nonne tu Deus qui reppulisti nos et non exibis Deus in virtutibus nostris
PS|107|13|da nobis auxilium de tribulatione quia vana salus hominis
PS|107|14|in Deo faciemus virtutem et ipse ad nihilum deducet inimicos nostros
PS|108|1|in finem David psalmus
PS|108|2|Deus laudem meam ne tacueris quia os peccatoris et os dolosi super me apertum est
PS|108|3|locuti sunt adversum me lingua dolosa et sermonibus odii circuierunt me et expugnaverunt me gratis
PS|108|4|pro eo ut me diligerent detrahebant mihi ego autem orabam
PS|108|5|et posuerunt adversus me mala pro bonis et odium pro dilectione mea
PS|108|6|constitue super eum peccatorem et diabulus stet a dextris eius
PS|108|7|cum iudicatur exeat condemnatus et oratio eius fiat in peccatum
PS|108|8|fiant dies eius pauci et episcopatum eius accipiat alter
PS|108|9|fiant filii eius orfani et uxor eius vidua
PS|108|10|nutantes transferantur filii eius et mendicent eiciantur de habitationibus suis
PS|108|11|scrutetur fenerator omnem substantiam eius et diripiant alieni labores eius
PS|108|12|non sit illi adiutor nec sit qui misereatur pupillis eius
PS|108|13|fiant nati eius in interitum in generatione una deleatur nomen eius
PS|108|14|in memoriam redeat iniquitas patrum eius in conspectu Domini et peccatum matris eius non deleatur
PS|108|15|fiant contra Dominum semper et dispereat de terra memoria eorum
PS|108|16|pro eo quod non est recordatus facere misericordiam
PS|108|17|et persecutus est hominem inopem et mendicum et conpunctum corde mortificare
PS|108|18|et dilexit maledictionem et veniet ei et noluit benedictionem et elongabitur ab eo et induit maledictionem sicut vestimentum et intravit sicut aqua in interiora eius et sicut oleum in ossibus eius
PS|108|19|fiat ei sicut vestimentum quo operitur et sicut zona qua semper praecingitur
PS|108|20|hoc opus eorum qui detrahunt mihi apud Dominum et qui loquuntur mala adversus animam meam
PS|108|21|et tu Domine Domine fac mecum propter nomen tuum quia suavis misericordia tua libera me
PS|108|22|quia egenus et pauper ego sum et cor meum turbatum est intra me
PS|108|23|sicut umbra cum declinat ablatus sum excussus sum sicut lucustae
PS|108|24|genua mea infirmata sunt a ieiunio et caro mea inmutata est propter oleum
PS|108|25|et ego factus sum obprobrium illis viderunt me moverunt capita sua
PS|108|26|adiuva me Domine Deus meus salvum fac me secundum misericordiam tuam
PS|108|27|et sciant quia manus tua haec tu Domine fecisti eam
PS|108|28|maledicent illi et tu benedices qui insurgunt in me confundantur servus autem tuus laetabitur
PS|108|29|induantur qui detrahunt mihi pudore et operiantur sicut deploide confusione sua
PS|108|30|confitebor Domino nimis in ore meo et in medio multorum laudabo eum
PS|108|31|quia adstetit a dextris pauperis ut salvam faceret a persequentibus animam meam
PS|109|1|David psalmus dixit Dominus Domino meo sede a dextris meis donec ponam inimicos tuos scabillum pedum tuorum
PS|109|2|virgam virtutis tuae emittet Dominus ex Sion dominare in medio inimicorum tuorum
PS|109|3|tecum principium in die virtutis tuae in splendoribus sanctorum ex utero ante luciferum genui te
PS|109|4|iuravit Dominus et non paenitebit eum tu es sacerdos in aeternum secundum ordinem Melchisedech
PS|109|5|Dominus a dextris tuis confregit in die irae suae reges
PS|109|6|iudicabit in nationibus implebit cadavera conquassabit capita in terra multorum
PS|109|7|de torrente in via bibet propterea exaltabit caput
PS|110|1|alleluia reversionis Aggei et Zacchariae confitebor tibi Domine in toto corde meo in consilio iustorum et congregatione
PS|110|2|magna opera Domini exquisita in omnes voluntates eius
PS|110|3|confessio et magnificentia opus eius et iustitia eius manet in saeculum saeculi
PS|110|4|memoriam fecit mirabilium suorum misericors et miserator Dominus
PS|110|5|escam dedit timentibus se memor erit in saeculum testamenti sui
PS|110|6|virtutem operum suorum adnuntiabit populo suo
PS|110|7|ut det illis hereditatem gentium opera manuum eius veritas et iudicium
PS|110|8|fidelia omnia mandata eius confirmata in saeculum saeculi facta in veritate et aequitate
PS|110|9|redemptionem misit populo suo mandavit in aeternum testamentum suum sanctum et terribile nomen eius
PS|110|10|initium sapientiae timor Domini intellectus bonus omnibus facientibus eum laudatio eius manet in saeculum %saeculi;
PS|111|1|alleluia reversionis Aggei et Zacchariae beatus vir qui timet Dominum in mandatis eius volet nimis
PS|111|2|potens in terra erit semen eius generatio rectorum benedicetur
PS|111|3|gloria et divitiae in domo eius et iustitia eius manet in saeculum saeculi
PS|111|4|exortum est in tenebris lumen rectis misericors et miserator et iustus
PS|111|5|iucundus homo qui miseretur et commodat disponet sermones suos in iudicio
PS|111|6|quia in aeternum non commovebitur
PS|111|7|in memoria aeterna erit iustus ab auditione mala non timebit paratum cor eius sperare in Domino
PS|111|8|confirmatum est cor eius non commovebitur donec dispiciat inimicos suos
PS|111|9|dispersit dedit pauperibus iustitia eius manet in saeculum saeculi cornu eius exaltabitur in gloria
PS|111|10|peccator videbit et irascetur dentibus suis fremet et tabescet desiderium peccatorum peribit
PS|112|1|alleluia laudate pueri Dominum laudate nomen Domini
PS|112|2|sit nomen Domini benedictum ex hoc nunc et usque in saeculum
PS|112|3|a solis ortu usque ad occasum laudabile nomen Domini
PS|112|4|excelsus super omnes gentes Dominus super caelos gloria eius
PS|112|5|quis sicut Dominus Deus noster qui in altis habitat
PS|112|6|et humilia respicit in caelo et in terra
PS|112|7|suscitans a terra inopem et de stercore erigens pauperem
PS|112|8|ut conlocet eum cum principibus cum principibus populi sui
PS|112|9|qui habitare facit sterilem in domo matrem filiorum laetantem
PS|113|1|alleluia in exitu Israhel de Aegypto domus Iacob de populo barbaro
PS|113|2|facta est Iudaea sanctificatio eius Israhel potestas eius
PS|113|3|mare vidit et fugit Iordanis conversus est retrorsum
PS|113|4|montes exultaverunt ut arietes colles sicut agni ovium
PS|113|5|quid est tibi mare quod fugisti et tu Iordanis quia conversus es retrorsum
PS|113|6|montes exultastis sicut arietes et colles sicut agni ovium
PS|113|7|a facie Domini mota est terra a facie Dei Iacob
PS|113|8|qui convertit petram in stagna aquarum et rupem in fontes aquarum
PS|113|9|non nobis Domine non nobis sed nomini tuo da gloriam
PS|113|10|super misericordia tua et veritate tua nequando dicant gentes ubi est Deus eorum
PS|113|11|Deus autem noster in caelo omnia quaecumque voluit fecit
PS|113|12|simulacra gentium argentum et aurum opera manuum hominum
PS|113|13|os habent et non loquentur oculos habent et non videbunt
PS|113|14|aures habent et non audient nares habent et non odorabuntur
PS|113|15|manus habent et non palpabunt pedes habent et non ambulabunt non clamabunt in gutture suo
PS|113|16|similes illis fiant qui faciunt ea et omnes qui confidunt in eis
PS|113|17|domus Israhel speravit in Domino adiutor eorum et protector eorum est
PS|113|18|domus Aaron speravit in Domino adiutor eorum et protector eorum est
PS|113|19|qui timent Dominum speraverunt in Domino adiutor eorum et protector eorum est
PS|113|20|Dominus memor fuit nostri et benedixit nobis benedixit domui Israhel benedixit domui Aaron
PS|113|21|benedixit omnibus qui timent Dominum pusillis cum maioribus
PS|113|22|adiciat Dominus super vos super vos et super filios vestros
PS|113|23|benedicti vos Domino qui fecit caelum et terram
PS|113|24|caelum caeli Domino terram autem dedit filiis hominum
PS|113|25|non mortui laudabunt te Domine neque omnes qui descendunt in infernum
PS|113|26|sed nos qui vivimus benedicimus Domino ex hoc nunc et usque in saeculum
PS|114|1|alleluia dilexi quoniam exaudiet Dominus vocem orationis meae
PS|114|2|quia inclinavit aurem suam mihi et in diebus meis invocabo te
PS|114|3|circumdederunt me dolores mortis pericula inferni invenerunt me tribulationem et dolorem inveni
PS|114|4|et nomen Domini invocavi o Domine libera animam meam
PS|114|5|misericors Dominus et iustus et Deus noster miseretur
PS|114|6|custodiens parvulos Dominus humiliatus sum et liberavit me
PS|114|7|convertere anima mea in requiem tuam quia Dominus benefecit tibi
PS|114|8|quia eripuit animam meam de morte oculos meos a lacrimis pedes meos a lapsu
PS|114|9|placebo Domino in regione vivorum
PS|115|1|alleluia credidi propter quod locutus sum ego autem humiliatus sum nimis
PS|115|2|ego dixi in excessu meo omnis homo mendax
PS|115|3|quid retribuam Domino pro omnibus quae retribuit mihi
PS|115|4|calicem salutaris accipiam et nomen Domini invocabo
PS|115|5|vota mea Domino reddam coram omni populo eius
PS|115|6|pretiosa in conspectu Domini mors sanctorum eius
PS|115|7|o Domine quia ego servus tuus ego servus tuus et filius ancillae tuae disrupisti vincula mea
PS|115|8|tibi sacrificabo hostiam laudis et in nomine Domini invocabo
PS|115|9|vota mea Domino reddam in conspectu omnis populi eius
PS|115|10|in atriis domus Domini in medio tui Hierusalem
PS|116|1|alleluia laudate Dominum omnes gentes laudate eum omnes populi
PS|116|2|quoniam confirmata est super nos misericordia eius et veritas Domini manet in saeculum
PS|117|1|alleluia confitemini Domino quoniam bonus quoniam in saeculum misericordia eius
PS|117|2|dicat nunc Israhel quoniam bonus quoniam in saeculum misericordia eius
PS|117|3|dicat nunc domus Aaron quoniam in saeculum misericordia eius
PS|117|4|dicant nunc qui timent Dominum quoniam in saeculum misericordia eius
PS|117|5|de tribulatione invocavi Dominum et exaudivit me in latitudinem Dominus
PS|117|6|Dominus mihi adiutor non timebo quid faciat mihi homo
PS|117|7|Dominus mihi adiutor et ego despiciam inimicos meos
PS|117|8|bonum est confidere in Domino quam confidere in homine
PS|117|9|bonum est sperare in Domino quam sperare in principibus
PS|117|10|omnes gentes circumierunt me et in nomine Domini quia; ultus sum in eos
PS|117|11|circumdantes circumdederunt me in nomine autem Domini quia; ultus sum in eos
PS|117|12|circumdederunt me sicut apes et exarserunt sicut ignis in spinis et in nomine Domini quia; ultus sum in eos
PS|117|13|inpulsus eversus sum ut caderem et Dominus suscepit me
PS|117|14|fortitudo mea et laudatio mea Dominus et factus est mihi in salutem
PS|117|15|vox exultationis et salutis in tabernaculis iustorum
PS|117|16|dextera Domini fecit virtutem dextera Domini exaltavit me dextera Domini fecit virtutem
PS|117|17|non moriar sed vivam et narrabo opera Domini
PS|117|18|castigans castigavit me Dominus et morti non tradidit me
PS|117|19|aperite mihi portas iustitiae ingressus in eas confitebor Domino
PS|117|20|haec porta Domini iusti intrabunt in eam
PS|117|21|confitebor tibi quoniam exaudisti me et factus es mihi in salutem
PS|117|22|lapidem quem reprobaverunt aedificantes hic factus est in caput anguli
PS|117|23|a Domino factum est istud hoc est mirabile in oculis nostris
PS|117|24|haec est dies quam fecit Dominus exultemus et laetemur in ea
PS|117|25|o Domine salvum fac o Domine prosperare
PS|117|26|benedictus qui venturus est in nomine Domini benediximus vobis de domo Domini
PS|117|27|Deus Dominus et inluxit nobis constituite diem sollemnem in condensis usque ad cornua altaris
PS|117|28|Deus meus es tu et confitebor tibi Deus meus % es tu; et exaltabo te confitebor tibi quoniam exaudisti me et factus es mihi in salutem
PS|117|29|confitemini Domino quoniam bonus quoniam in saeculum misericordia eius
PS|118|1|alleluia aleph beati inmaculati in via qui ambulant in lege Domini
PS|118|2|beati qui scrutantur testimonia eius in toto corde exquirent eum
PS|118|3|non enim qui operantur iniquitatem in viis eius ambulaverunt
PS|118|4|tu mandasti mandata tua custodire nimis
PS|118|5|utinam dirigantur viae meae ad custodiendas iustificationes tuas
PS|118|6|tunc non confundar cum perspexero in omnibus mandatis tuis
PS|118|7|confitebor tibi in directione cordis in eo quod didici iudicia iustitiae tuae
PS|118|8|iustificationes tuas custodiam non me derelinquas usquequaque
PS|118|9|beth in quo corriget adulescentior viam suam in custodiendo sermones tuos
PS|118|10|in toto corde meo exquisivi te non repellas me a mandatis tuis
PS|118|11|in corde meo abscondi eloquia tua ut non peccem tibi
PS|118|12|benedictus es Domine doce me iustificationes tuas
PS|118|13|in labiis meis pronuntiavi omnia iudicia oris tui
PS|118|14|in via testimoniorum tuorum delectatus sum sicut in omnibus divitiis
PS|118|15|in mandatis tuis exercebor et considerabo vias tuas
PS|118|16|in iustificationibus tuis meditabor non obliviscar sermones tuos
PS|118|17|gimel retribue servo tuo vivifica me et custodiam sermones tuos
PS|118|18|revela oculos meos et considerabo mirabilia de lege tua
PS|118|19|incola ego sum in terra non abscondas a me mandata tua
PS|118|20|concupivit anima mea desiderare iustificationes tuas in omni tempore
PS|118|21|increpasti superbos maledicti qui declinant a mandatis tuis
PS|118|22|aufer a me obprobrium et contemptum quia testimonia tua exquisivi
PS|118|23|etenim sederunt principes et adversum me loquebantur servus autem tuus exercebatur in iustificationibus tuis
PS|118|24|nam et testimonia tua meditatio mea et consilium meum iustificationes tuae
PS|118|25|deleth adhesit pavimento anima mea vivifica me secundum verbum tuum
PS|118|26|vias meas enuntiavi et exaudisti me doce me iustificationes tuas
PS|118|27|viam iustificationum tuarum instrue me et exercebor in mirabilibus tuis
PS|118|28|dormitavit anima mea prae taedio confirma me in verbis tuis
PS|118|29|viam iniquitatis amove a me et lege tua miserere mei
PS|118|30|viam veritatis elegi iudicia tua non sum oblitus
PS|118|31|adhesi testimoniis tuis Domine noli me confundere
PS|118|32|viam mandatorum tuorum cucurri cum dilatasti cor meum
PS|118|33|he legem pone mihi Domine viam iustificationum tuarum et exquiram eam semper
PS|118|34|da mihi intellectum et scrutabor legem tuam et custodiam illam in toto corde meo
PS|118|35|deduc me in semita mandatorum tuorum quia ipsam volui
PS|118|36|inclina cor meum in testimonia tua et non in avaritiam
PS|118|37|averte oculos meos ne videant vanitatem in via tua vivifica me
PS|118|38|statue servo tuo eloquium tuum in timore tuo
PS|118|39|amputa obprobrium meum quod suspicatus sum quia iudicia tua iucunda
PS|118|40|ecce concupivi mandata tua in aequitate tua vivifica me
PS|118|41|vav et veniat super me misericordia tua Domine salutare tuum secundum eloquium tuum
PS|118|42|et respondebo exprobrantibus mihi verbum quia speravi in sermonibus tuis
PS|118|43|et ne auferas de ore meo verbum veritatis usquequaque quia in iudiciis tuis supersperavi
PS|118|44|et custodiam legem tuam semper in saeculum et in saeculum saeculi
PS|118|45|et ambulabam in latitudine quia mandata tua exquisivi
PS|118|46|et loquebar in testimoniis tuis in conspectu regum et non confundebar
PS|118|47|et meditabar in mandatis tuis quae dilexi
PS|118|48|et levavi manus meas ad mandata quae dilexi et exercebar in iustificationibus tuis
PS|118|49|zai memor esto verbi tui servo tuo in quo mihi spem dedisti
PS|118|50|haec me consolata est in humilitate mea quia eloquium tuum vivificavit me
PS|118|51|superbi inique agebant usquequaque a lege autem tua non declinavi
PS|118|52|memor fui iudiciorum tuorum a saeculo Domine et consolatus sum
PS|118|53|defectio tenuit me prae peccatoribus derelinquentibus legem tuam
PS|118|54|cantabiles mihi erant iustificationes tuae in loco peregrinationis meae
PS|118|55|memor fui in nocte nominis tui Domine et custodivi legem tuam
PS|118|56|haec facta est mihi quia iustificationes tuas exquisivi
PS|118|57|heth portio mea Dominus dixi custodire legem tuam
PS|118|58|deprecatus sum faciem tuam in toto corde meo miserere mei secundum eloquium tuum
PS|118|59|cogitavi vias meas et avertisti pedes meos in testimonia tua
PS|118|60|paratus sum et non sum turbatus ut custodiam mandata tua
PS|118|61|funes peccatorum circumplexi sunt me et legem tuam non sum oblitus
PS|118|62|media nocte surgebam ad confitendum tibi super iudicia iustificationis tuae
PS|118|63|particeps ego sum omnium timentium te et custodientium mandata tua
PS|118|64|misericordia Domini plena est terra iustificationes tuas doce me
PS|118|65|teth bonitatem fecisti cum servo tuo Domine secundum verbum tuum
PS|118|66|bonitatem et disciplinam et scientiam doce me quia mandatis tuis credidi
PS|118|67|priusquam humiliarer ego deliqui propterea eloquium tuum custodivi
PS|118|68|bonus es tu et in bonitate tua doce me iustificationes tuas
PS|118|69|multiplicata est super me iniquitas superborum ego autem in toto corde scrutabor mandata tua
PS|118|70|coagulatum est sicut lac cor eorum ego vero legem tuam meditatus sum
PS|118|71|bonum mihi quia humiliasti me ut discam iustificationes tuas
PS|118|72|bonum mihi lex oris tui super milia auri et argenti
PS|118|73|ioth manus tuae fecerunt me et plasmaverunt me da mihi intellectum et discam mandata tua
PS|118|74|qui timent te videbunt me et laetabuntur quia in verba tua supersperavi
PS|118|75|cognovi Domine quia aequitas iudicia tua et veritate humiliasti me
PS|118|76|fiat misericordia tua ut consoletur me secundum eloquium tuum servo tuo
PS|118|77|veniant mihi miserationes tuae et vivam quia lex tua meditatio mea est
PS|118|78|confundantur superbi quia iniuste iniquitatem fecerunt in me ego autem exercebor in mandatis tuis
PS|118|79|convertantur mihi timentes te et qui noverunt testimonia tua
PS|118|80|fiat cor meum inmaculatum in iustificationibus tuis ut non confundar
PS|118|81|caf defecit in salutare tuum anima mea in verbum tuum supersperavi
PS|118|82|defecerunt oculi mei in eloquium tuum dicentes quando consolaberis me
PS|118|83|quia factus sum sicut uter in pruina iustificationes tuas non sum oblitus
PS|118|84|quot sunt dies servo tuo quando facies de persequentibus me iudicium
PS|118|85|narraverunt mihi iniqui fabulationes sed non ut lex tua
PS|118|86|omnia mandata tua veritas inique persecuti sunt me adiuva me
PS|118|87|paulo minus consummaverunt me in terra ego autem non dereliqui mandata tua
PS|118|88|secundum misericordiam tuam vivifica me et custodiam testimonia oris tui
PS|118|89|lamed in aeternum Domine verbum tuum permanet in caelo
PS|118|90|in generationem et generationem veritas tua fundasti terram et permanet
PS|118|91|ordinatione tua perseverat dies quoniam omnia serviunt tibi
PS|118|92|nisi quod lex tua meditatio mea est tunc forte perissem in humilitate mea
PS|118|93|in aeternum non obliviscar iustificationes tuas quia in ipsis vivificasti me
PS|118|94|tuus sum ego salvum me fac quoniam iustificationes tuas exquisivi
PS|118|95|me expectaverunt peccatores ut perderent me testimonia tua intellexi
PS|118|96|omni consummationi vidi finem latum mandatum tuum nimis
PS|118|97|mem quomodo dilexi legem tuam tota die meditatio mea est
PS|118|98|super inimicos meos prudentem me fecisti mandato tuo quia in aeternum mihi est
PS|118|99|super omnes docentes me intellexi quia testimonia tua meditatio mea est
PS|118|100|super senes intellexi quia mandata tua quaesivi
PS|118|101|ab omni via mala prohibui pedes meos ut custodiam verba tua
PS|118|102|a iudiciis tuis non declinavi quia tu legem posuisti mihi
PS|118|103|quam dulcia faucibus meis eloquia tua super mel ori meo
PS|118|104|a mandatis tuis intellexi propterea odivi omnem viam iniquitatis
PS|118|105|nun lucerna pedibus meis verbum tuum et lumen semitis meis
PS|118|106|iuravi et statui custodire iudicia iustitiae tuae
PS|118|107|humiliatus sum usquequaque Domine vivifica me secundum verbum tuum
PS|118|108|voluntaria oris mei beneplacita fac Domine et iudicia tua doce me
PS|118|109|anima mea in manibus meis semper et legem tuam non sum oblitus
PS|118|110|posuerunt peccatores laqueum mihi et de mandatis tuis non erravi
PS|118|111|hereditate adquisivi testimonia tua in aeternum quia exultatio cordis mei sunt
PS|118|112|inclinavi cor meum ad faciendas iustificationes tuas in aeternum propter retributionem
PS|118|113|samech iniquos odio habui et legem tuam dilexi
PS|118|114|adiutor meus et susceptor meus es tu in verbum tuum supersperavi
PS|118|115|declinate a me maligni et scrutabor mandata Dei mei
PS|118|116|suscipe me secundum eloquium tuum et vivam et non confundas me ab expectatione mea
PS|118|117|adiuva me et salvus ero et meditabor in iustificationibus tuis semper
PS|118|118|sprevisti omnes discedentes a iustitiis tuis quia iniusta cogitatio eorum
PS|118|119|praevaricantes reputavi omnes peccatores terrae ideo dilexi testimonia tua
PS|118|120|confige timore tuo carnes meas a iudiciis %enim; tuis timui
PS|118|121|ain feci iudicium et iustitiam non tradas me calumniantibus me
PS|118|122|suscipe servum tuum in bonum non calumnientur me superbi
PS|118|123|oculi mei defecerunt in salutare tuum et in eloquium iustitiae tuae
PS|118|124|fac cum servo tuo secundum misericordiam tuam et iustificationes tuas doce me
PS|118|125|servus tuus sum ego da mihi intellectum et sciam testimonia tua
PS|118|126|tempus faciendi Domino dissipaverunt legem tuam
PS|118|127|ideo dilexi mandata tua super aurum et topazion
PS|118|128|propterea ad omnia mandata tua dirigebar omnem viam iniquam odio habui
PS|118|129|fe mirabilia testimonia tua ideo scrutata est ea anima mea
PS|118|130|declaratio sermonum tuorum inluminat et intellectum dat parvulis
PS|118|131|os meum aperui et adtraxi spiritum quia mandata tua desiderabam
PS|118|132|aspice in me et miserere mei secundum iudicium diligentium nomen tuum
PS|118|133|gressus meos dirige secundum eloquium tuum et non dominetur mei omnis iniustitia
PS|118|134|redime me a calumniis hominum et custodiam mandata tua
PS|118|135|faciem tuam inlumina super servum tuum et doce me iustificationes tuas
PS|118|136|exitus aquarum deduxerunt oculi mei quia non custodierunt legem tuam
PS|118|137|sade iustus es Domine et rectum iudicium tuum
PS|118|138|mandasti iustitiam testimonia tua et veritatem tuam nimis
PS|118|139|tabescere me fecit zelus meus quia obliti sunt verba tua inimici mei
PS|118|140|ignitum eloquium tuum vehementer et servus tuus dilexit illud
PS|118|141|adulescentulus sum ego et contemptus iustificationes tuas non sum oblitus
PS|118|142|iustitia tua iustitia in aeternum et lex tua veritas
PS|118|143|tribulatio et angustia invenerunt me mandata tua meditatio mea
PS|118|144|aequitas testimonia tua in aeternum intellectum da mihi et vivam
PS|118|145|cof clamavi in toto corde exaudi me Domine iustificationes tuas requiram
PS|118|146|clamavi te salvum me fac et custodiam mandata tua
PS|118|147|praeveni in maturitate et clamavi in verba tua supersperavi
PS|118|148|praevenerunt oculi mei ad diluculum ut meditarer eloquia tua
PS|118|149|vocem meam audi secundum misericordiam tuam Domine secundum iudicium tuum vivifica me
PS|118|150|adpropinquaverunt persequentes me iniquitate a lege autem tua longe facti sunt
PS|118|151|prope es tu Domine et omnes viae tuae veritas
PS|118|152|initio cognovi de testimoniis tuis quia in aeternum fundasti ea
PS|118|153|res vide humilitatem meam et eripe me quia legem tuam non sum oblitus
PS|118|154|iudica iudicium meum et redime me propter eloquium tuum vivifica me
PS|118|155|longe a peccatoribus salus quia iustificationes tuas non exquisierunt
PS|118|156|misericordiae tuae multae Domine secundum iudicia tua vivifica me
PS|118|157|multi qui persequuntur me et tribulant me a testimoniis tuis non declinavi
PS|118|158|vidi praevaricantes et tabescebam quia eloquia tua non custodierunt
PS|118|159|vide quoniam mandata tua dilexi Domine in misericordia tua vivifica me
PS|118|160|principium verborum tuorum veritas et in aeternum omnia iudicia iustitiae tuae
PS|118|161|sen principes persecuti sunt me gratis et a verbis tuis formidavit cor meum
PS|118|162|laetabor ego super eloquia tua sicut qui invenit spolia multa
PS|118|163|iniquitatem odio habui et abominatus sum legem autem tuam dilexi
PS|118|164|septies in die laudem dixi tibi super iudicia iustitiae tuae
PS|118|165|pax multa diligentibus legem tuam et non est illis scandalum
PS|118|166|expectabam salutare tuum Domine et mandata tua dilexi
PS|118|167|custodivit anima mea testimonia tua et dilexi ea vehementer
PS|118|168|servavi mandata tua et testimonia tua quia omnes viae meae in conspectu tuo
PS|118|169|thau adpropinquet deprecatio mea in conspectu tuo Domine iuxta eloquium tuum da mihi intellectum
PS|118|170|intret postulatio mea in conspectu tuo secundum eloquium tuum eripe me
PS|118|171|eructabunt labia mea hymnum cum docueris me iustificationes tuas
PS|118|172|pronuntiabit lingua mea eloquium tuum quia omnia mandata tua aequitas
PS|118|173|fiat manus tua ut salvet me quoniam mandata tua elegi
PS|118|174|concupivi salutare tuum Domine et lex tua meditatio mea
PS|118|175|vivet anima mea et laudabit te et iudicia tua adiuvabunt me
PS|118|176|erravi sicut ovis quae periit quaere servum tuum quia mandata tua non sum oblitus
PS|119|1|canticum graduum ad Dominum cum tribularer clamavi et exaudivit me
PS|119|2|Domine libera animam meam a labiis iniquis a lingua dolosa
PS|119|3|quid detur tibi et quid adponatur tibi ad linguam dolosam
PS|119|4|sagittae potentis acutae cum carbonibus desolatoriis
PS|119|5|heu mihi quia incolatus meus prolongatus est habitavi cum habitationibus Cedar
PS|119|6|multum incola fuit anima mea
PS|119|7|cum his qui oderant pacem eram pacificus cum loquebar illis inpugnabant me gratis
PS|120|1|canticum graduum levavi oculos meos in montes unde veniet auxilium mihi
PS|120|2|auxilium meum a Domino qui fecit caelum et terram
PS|120|3|non det in commotionem pedem tuum neque dormitet qui custodit te
PS|120|4|ecce non dormitabit neque dormiet qui custodit Israhel
PS|120|5|Dominus custodit te Dominus protectio tua super manum dexteram tuam
PS|120|6|per diem sol non uret te neque luna per noctem
PS|120|7|Dominus custodit te ab omni malo custodiat animam tuam Dominus
PS|120|8|Dominus custodiat introitum tuum et exitum tuum ex hoc nunc et usque in saeculum
PS|121|1|canticum graduum huic David laetatus sum in his quae dicta sunt mihi in domum Domini ibimus
PS|121|2|stantes erant pedes nostri in atriis tuis Hierusalem
PS|121|3|Hierusalem quae aedificatur ut civitas cuius participatio eius in id ipsum
PS|121|4|illic enim ascenderunt tribus tribus Domini testimonium Israhel ad confitendum nomini Domini
PS|121|5|quia illic sederunt sedes in iudicium sedes super domum David
PS|121|6|rogate quae ad pacem sunt Hierusalem et abundantia diligentibus te
PS|121|7|fiat pax in virtute tua et abundantia in turribus tuis
PS|121|8|propter fratres meos et proximos meos loquebar pacem de te
PS|121|9|propter domum Domini Dei nostri quaesivi bona tibi
PS|122|1|canticum graduum ad te levavi oculos meos qui habitas in caelo
PS|122|2|ecce sicut oculi servorum in manibus dominorum suorum sicut oculi ancillae in manibus dominae eius ita oculi nostri ad Dominum Deum nostrum donec misereatur nostri
PS|122|3|miserere nostri Domine miserere nostri quia multum repleti sumus despectione
PS|122|4|quia multum repleta est anima nostra obprobrium abundantibus et despectio superbis
PS|123|1|canticum graduum huic David nisi quia Dominus erat in nobis dicat nunc Israhel
PS|123|2|nisi quia Dominus erat in nobis cum exsurgerent in nos homines
PS|123|3|forte vivos degluttissent nos cum irasceretur furor eorum in nos
PS|123|4|forsitan aqua absorbuisset nos
PS|123|5|torrentem pertransivit anima nostra forsitan pertransisset anima nostra aquam intolerabilem
PS|123|6|benedictus Dominus qui non dedit nos in captionem dentibus eorum
PS|123|7|anima nostra sicut passer erepta est de laqueo venantium laqueus contritus est et nos liberati sumus
PS|123|8|adiutorium nostrum in nomine Domini qui fecit caelum et terram
PS|124|1|canticum graduum qui confidunt in Domino sicut mons Sion non commovebitur in aeternum qui habitat
PS|124|2|in Hierusalem montes in circuitu eius et Dominus in circuitu populi sui ex hoc nunc et usque in saeculum
PS|124|3|quia non relinquet virgam peccatorum super sortem iustorum ut non extendant iusti ad iniquitatem manus suas
PS|124|4|benefac Domine bonis et rectis corde
PS|124|5|declinantes autem in obligationes adducet Dominus cum operantibus iniquitatem pax super Israhel
PS|125|1|canticum graduum in convertendo Dominum captivitatem Sion facti sumus sicut consolati
PS|125|2|tunc repletum est gaudio os nostrum et lingua nostra exultatione tunc dicent inter gentes magnificavit Dominus facere cum eis
PS|125|3|magnificavit Dominus facere nobiscum facti sumus laetantes
PS|125|4|converte Domine captivitatem nostram sicut torrens in austro
PS|125|5|qui seminant in lacrimis in exultatione metent
PS|125|6|euntes ibant et flebant portantes semina sua venientes autem venient in exultatione portantes manipulos suos
PS|126|1|canticum graduum Salomonis nisi Dominus aedificaverit domum in vanum laboraverunt qui aedificant eam nisi Dominus custodierit civitatem frustra vigilavit qui custodit
PS|126|2|vanum est vobis ante lucem surgere surgere postquam sederitis qui manducatis panem doloris cum dederit dilectis suis somnum
PS|126|3|ecce hereditas Domini filii mercis fructus ventris
PS|126|4|sicut sagittae in manu potentis ita filii excussorum
PS|126|5|beatus vir qui implebit desiderium suum ex ipsis non confundentur cum loquentur inimicis suis in porta
PS|127|1|canticum graduum beati omnes qui timent Dominum qui ambulant in viis eius
PS|127|2|labores manuum tuarum quia; manducabis beatus es et bene tibi erit
PS|127|3|uxor tua sicut vitis abundans in lateribus domus tuae filii tui sicut novella olivarum in circuitu mensae tuae
PS|127|4|ecce sic benedicetur homo qui timet Dominum
PS|127|5|benedicat te Dominus ex Sion et videas bona Hierusalem omnibus diebus vitae tuae
PS|127|6|et videas filios filiorum tuorum pax super Israhel
PS|128|1|canticum graduum saepe expugnaverunt me a iuventute mea dicat nunc Israhel
PS|128|2|saepe expugnaverunt me a iuventute mea etenim non potuerunt mihi
PS|128|3|supra dorsum meum fabricabantur peccatores prolongaverunt iniquitatem suam
PS|128|4|Dominus iustus concidet cervices peccatorum
PS|128|5|confundantur et convertantur retrorsum omnes qui oderunt Sion
PS|128|6|fiant sicut faenum tectorum quod priusquam evellatur exaruit
PS|128|7|de quo non implevit manum suam qui metit et sinum suum qui manipulos colligit
PS|128|8|et non dixerunt qui praeteribant benedictio Domini super vos benediximus vobis in nomine Domini
PS|129|1|canticum graduum de profundis clamavi ad te Domine
PS|129|2|Domine exaudi vocem meam fiant aures tuae intendentes in vocem deprecationis meae
PS|129|3|si iniquitates observabis Domine Domine quis sustinebit
PS|129|4|quia apud te propitiatio est propter legem tuam sustinui te Domine sustinuit anima mea in verbum eius
PS|129|5|speravit anima mea in Domino
PS|129|6|a custodia matutina usque ad noctem speret Israhel in Domino
PS|129|7|quia apud Dominum misericordia et copiosa apud eum redemptio
PS|129|8|et ipse redimet Israhel ex omnibus iniquitatibus eius
PS|130|1|canticum graduum David Domine non est exaltatum cor meum neque elati sunt oculi mei neque ambulavi in magnis neque in mirabilibus super me
PS|130|2|si non humiliter sentiebam sed exaltavi animam meam sicut ablactatum super matrem suam ita retributio in anima mea
PS|130|3|speret Israhel in Domino ex hoc nunc et usque in saeculum
PS|131|1|canticum graduum memento Domine David et omnis mansuetudinis eius
PS|131|2|sicut iuravit Domino votum vovit Deo Iacob
PS|131|3|si introiero in tabernaculum domus meae si ascendero in lectum strati mei
PS|131|4|si dedero somnum oculis meis et palpebris meis dormitationem
PS|131|5|et requiem temporibus meis donec inveniam locum Domino tabernaculum Deo Iacob
PS|131|6|ecce audivimus eam in Efrata invenimus eam in campis silvae
PS|131|7|introibimus in tabernacula eius adorabimus in loco ubi steterunt pedes eius
PS|131|8|surge Domine in requiem tuam tu et arca sanctificationis tuae
PS|131|9|sacerdotes tui induentur iustitia et sancti tui exultabunt
PS|131|10|propter David servum tuum non avertas faciem christi tui
PS|131|11|iuravit Dominus David veritatem et non frustrabit eum de fructu ventris tui ponam super sedem tuam
PS|131|12|si custodierint filii tui testamentum meum et testimonia mea haec quae docebo eos et filii eorum usque in saeculum sedebunt super sedem tuam
PS|131|13|quoniam elegit Dominus Sion elegit eam in habitationem sibi
PS|131|14|haec requies mea in saeculum saeculi hic habitabo quoniam elegi eam
PS|131|15|viduam eius benedicens benedicam pauperes eius saturabo panibus
PS|131|16|sacerdotes eius induam salutari et sancti eius exultatione exultabunt
PS|131|17|illic producam cornu David paravi lucernam christo meo
PS|131|18|inimicos eius induam confusione super ipsum autem efflorebit sanctificatio mea
PS|132|1|canticum graduum David ecce quam bonum et quam iucundum habitare fratres in unum
PS|132|2|sicut unguentum in capite quod descendit in barbam barbam Aaron quod descendit in ora vestimenti eius
PS|132|3|sicut ros Hermon qui descendit in montes Sion quoniam illic mandavit Dominus benedictionem et vitam usque in saeculum
PS|133|1|canticum graduum ecce nunc benedicite Dominum omnes servi Domini qui statis in domo Domini %in atriis domus Dei nostri;
PS|133|2|in noctibus extollite manus vestras in sancta et benedicite Domino
PS|133|3|benedicat te Dominus ex Sion qui fecit caelum et terram
PS|134|1|alleluia laudate nomen Domini laudate servi Dominum
PS|134|2|qui statis in domo Domini in atriis domus Dei nostri
PS|134|3|laudate Dominum quia bonus Dominus psallite nomini eius quoniam suave
PS|134|4|quoniam Iacob elegit sibi Dominus Israhel in possessionem sibi
PS|134|5|quia ego cognovi quod magnus est Dominus et Deus noster prae omnibus diis
PS|134|6|omnia quae voluit Dominus fecit in caelo et in terra in mare et in omnibus abyssis
PS|134|7|educens nubes ab extremo terrae fulgora in pluviam fecit qui producit ventos de thesauris suis
PS|134|8|qui percussit primogenita Aegypti ab homine usque ad pecus
PS|134|9|emisit signa et prodigia in medio tui Aegypte in Pharaonem et in omnes servos eius
PS|134|10|qui percussit gentes multas et occidit reges fortes
PS|134|11|Seon regem Amorreorum et Og regem Basan et omnia regna Chanaan
PS|134|12|et dedit terram eorum hereditatem hereditatem Israhel populo suo
PS|134|13|Domine nomen tuum in aeternum Domine memoriale tuum in generationem et generationem
PS|134|14|quia iudicabit Dominus populum suum et in servis suis deprecabitur
PS|134|15|simulacra gentium argentum et aurum opera manuum hominum
PS|134|16|os habent et non loquentur oculos habent et non videbunt
PS|134|17|aures habent et non audient neque enim est spiritus in ore eorum
PS|134|18|similes illis fiant qui faciunt ea et omnes qui sperant in eis
PS|134|19|domus Israhel benedicite Domino domus Aaron benedicite Domino
PS|134|20|domus Levi benedicite Domino qui timetis Dominum benedicite Domino
PS|134|21|benedictus Dominus ex Sion qui habitat in Hierusalem
PS|135|1|alleluia confitemini Domino quoniam bonus quoniam in aeternum misericordia eius
PS|135|2|confitemini Deo deorum quoniam in aeternum misericordia eius
PS|135|3|confitemini Domino dominorum quoniam in aeternum misericordia eius
PS|135|4|qui facit mirabilia magna solus quoniam in aeternum misericordia eius
PS|135|5|qui fecit caelos in intellectu quoniam in aeternum misericordia eius
PS|135|6|qui firmavit terram super aquas quoniam in aeternum misericordia eius
PS|135|7|qui fecit luminaria magna quoniam in aeternum misericordia eius
PS|135|8|solem in potestatem diei quoniam in aeternum misericordia eius
PS|135|9|lunam et stellas in potestatem noctis quoniam in aeternum misericordia eius
PS|135|10|qui percussit Aegyptum cum primogenitis eorum quoniam in aeternum misericordia eius
PS|135|11|qui eduxit Israhel de medio eorum quoniam in aeternum misericordia eius
PS|135|12|in manu potenti et brachio excelso quoniam in aeternum misericordia eius
PS|135|13|qui divisit Rubrum mare in divisiones quoniam in aeternum misericordia eius
PS|135|14|et duxit Israhel per medium eius quoniam in aeternum misericordia eius
PS|135|15|et excussit Pharaonem et virtutem eius in mari Rubro quoniam in aeternum misericordia eius
PS|135|16|qui transduxit populum suum in deserto quoniam in aeternum misericordia eius
PS|135|17|qui percussit reges magnos quoniam in aeternum misericordia eius
PS|135|18|et occidit reges fortes quoniam in aeternum misericordia eius
PS|135|19|Seon regem Amorreorum quoniam in aeternum misericordia eius
PS|135|20|et Og regem Basan quoniam in aeternum misericordia eius
PS|135|21|et dedit terram eorum hereditatem quoniam in aeternum misericordia eius
PS|135|22|hereditatem Israhel servo suo quoniam in aeternum misericordia eius
PS|135|23|quia in humilitate nostra memor fuit nostri quoniam in aeternum misericordia eius
PS|135|24|et redemit nos ab inimicis nostris quoniam in aeternum misericordia eius
PS|135|25|qui dat escam omni carni quoniam in aeternum misericordia eius
PS|135|26|confitemini Deo caeli quoniam in aeternum misericordia eius confitemini Domino dominorum quoniam in aeternum misericordia eius
PS|136|1|David Hieremiae super flumina Babylonis illic sedimus et flevimus cum recordaremur Sion
PS|136|2|in salicibus in medio eius suspendimus organa nostra
PS|136|3|quia illic interrogaverunt nos qui captivos duxerunt nos verba cantionum et qui abduxerunt nos hymnum cantate nobis de canticis Sion
PS|136|4|quomodo cantabimus canticum Domini in terra aliena
PS|136|5|si oblitus fuero tui Hierusalem oblivioni detur dextera mea
PS|136|6|adhereat lingua mea faucibus meis si non meminero tui si non praeposuero Hierusalem in principio laetitiae meae
PS|136|7|memor esto Domine filiorum Edom diem Hierusalem qui dicunt exinanite exinanite usque ad fundamentum in ea
PS|136|8|filia Babylonis misera beatus qui retribuet tibi retributionem tuam quam retribuisti nobis
PS|136|9|beatus qui tenebit et adlidet parvulos tuos ad petram
PS|137|1|ipsi David confitebor tibi Domine in toto corde meo quoniam audisti verba oris mei in conspectu angelorum psallam tibi
PS|137|2|adorabo ad templum sanctum tuum et confitebor nomini tuo super misericordia tua et veritate tua quoniam magnificasti super omne nomen sanctum tuum
PS|137|3|in quacumque die invocavero te exaudi me multiplicabis me in anima mea virtute
PS|137|4|confiteantur tibi Domine omnes reges terrae quia audierunt omnia verba oris tui
PS|137|5|et cantent in viis Domini quoniam magna gloria Domini
PS|137|6|quoniam excelsus Dominus et humilia respicit et alta a longe cognoscit
PS|137|7|si ambulavero in medio tribulationis vivificabis me super iram inimicorum meorum extendisti manum tuam et salvum me fecit dextera tua
PS|137|8|Dominus retribuet propter me Domine misericordia tua in saeculum opera manuum tuarum ne dispicias
PS|138|1|in finem David psalmus
PS|138|2|Domine probasti me et cognovisti me tu cognovisti sessionem meam et surrectionem meam
PS|138|3|intellexisti cogitationes meas de longe semitam meam et funiculum meum investigasti
PS|138|4|et omnes vias meas praevidisti quia non est sermo in lingua mea
PS|138|5|ecce Domine tu cognovisti omnia novissima et antiqua tu formasti me et posuisti super me manum tuam
PS|138|6|mirabilis facta est scientia tua ex me confortata est non potero ad eam
PS|138|7|quo ibo ab spiritu tuo et quo a facie tua fugiam
PS|138|8|si ascendero in caelum tu illic es si descendero ad infernum ades
PS|138|9|si sumpsero pinnas meas diluculo et habitavero in extremis maris
PS|138|10|etenim illuc manus tua deducet me et tenebit me dextera tua
PS|138|11|et dixi forsitan tenebrae conculcabunt me et nox inluminatio in deliciis meis
PS|138|12|quia tenebrae non obscurabuntur a te et nox sicut dies inluminabitur sicut tenebrae eius ita et lumen eius
PS|138|13|quia tu possedisti renes meos suscepisti me de utero matris meae
PS|138|14|confitebor tibi quia terribiliter magnificatus es mirabilia opera tua et anima mea cognoscit nimis
PS|138|15|non est occultatum os meum a te quod fecisti in occulto et substantia mea in inferioribus terrae
PS|138|16|inperfectum meum viderunt oculi tui et in libro tuo omnes scribentur die formabuntur et nemo in eis
PS|138|17|mihi autem nimis honorificati sunt amici tui Deus nimis confirmati sunt principatus eorum
PS|138|18|dinumerabo eos et super harenam multiplicabuntur exsurrexi et adhuc sum tecum
PS|138|19|si occideris Deus peccatores et viri sanguinum declinate a me
PS|138|20|quia dices in cogitatione accipient in vanitate civitates tuas
PS|138|21|nonne qui oderunt te Domine oderam et super inimicos tuos tabescebam
PS|138|22|perfecto odio oderam illos inimici facti sunt mihi
PS|138|23|proba me Deus et scito cor meum interroga me et cognosce semitas meas
PS|138|24|et vide si via iniquitatis in me est et deduc me in via aeterna
PS|139|1|in finem psalmus David
PS|139|2|eripe me Domine ab homine malo a viro iniquo eripe me
PS|139|3|qui cogitaverunt iniquitates in corde tota die constituebant proelia
PS|139|4|acuerunt linguam suam sicut serpentis venenum aspidum sub labiis eorum diapsalma
PS|139|5|custodi me Domine de manu peccatoris ab hominibus iniquis eripe me qui cogitaverunt subplantare gressus meos
PS|139|6|absconderunt superbi laqueum mihi et funes extenderunt in laqueum iuxta iter scandalum posuerunt mihi diapsalma
PS|139|7|dixi Domino Deus meus es tu exaudi Domine vocem deprecationis meae
PS|139|8|Domine Domine virtus salutis meae obumbrasti super caput meum in die belli
PS|139|9|non tradas Domine desiderio meo peccatori cogitaverunt contra me ne derelinquas me ne forte exaltentur diapsalma
PS|139|10|caput circuitus eorum labor labiorum ipsorum operiet eos
PS|139|11|cadent super eos carbones in igne deicies eos in miseriis non subsistent
PS|139|12|vir linguosus non dirigetur in terra virum iniustum mala capient in interitu
PS|139|13|cognovi quia faciet Dominus iudicium inopis et vindictam pauperum
PS|139|14|verumtamen iusti confitebuntur nomini tuo habitabunt recti cum vultu tuo
PS|140|1|psalmus David Domine clamavi ad te exaudi me intende voci meae cum clamavero ad te
PS|140|2|dirigatur oratio mea sicut incensum in conspectu tuo elevatio manuum mearum sacrificium vespertinum
PS|140|3|pone Domine custodiam ori meo et ostium circumstantiae labiis meis
PS|140|4|non declines cor meum in verba malitiae ad excusandas excusationes in peccatis cum hominibus operantibus iniquitatem et non communicabo cum electis eorum
PS|140|5|corripiet me iustus in misericordia et increpabit me oleum %autem; peccatoris non inpinguet caput meum quoniam adhuc et oratio mea in beneplacitis eorum
PS|140|6|absorti sunt iuncti petrae iudices eorum audient verba mea quoniam potuerunt
PS|140|7|sicut crassitudo terrae erupta est super terram dissipata sunt ossa nostra secus infernum
PS|140|8|quia ad te Domine Domine oculi mei in te speravi non auferas animam meam
PS|140|9|custodi me a laqueo quem statuerunt mihi et ab scandalis operantium iniquitatem
PS|140|10|cadent in retiaculo eius peccatores singulariter sum ego donec transeam
PS|141|1|intellectus David cum esset in spelunca oratio
PS|141|2|voce mea ad Dominum clamavi voce mea ad Dominum deprecatus sum
PS|141|3|effundo in conspectu eius deprecationem meam tribulationem meam ante ipsum pronuntio
PS|141|4|in deficiendo ex me spiritum meum et tu cognovisti semitas meas in via hac qua ambulabam absconderunt laqueum mihi
PS|141|5|considerabam ad dexteram et videbam et non erat qui cognosceret me periit fuga a me et non est qui requirit animam meam
PS|141|6|clamavi ad te Domine dixi tu es spes mea portio mea in terra viventium
PS|141|7|intende ad deprecationem meam quia humiliatus sum nimis libera me a persequentibus me quia confortati sunt super me
PS|141|8|educ de custodia animam meam ad confitendum nomini tuo me expectant iusti donec retribuas mihi
PS|142|1|psalmus David quando filius eum persequebatur Domine exaudi orationem meam auribus percipe obsecrationem meam in veritate tua exaudi me in tua iustitia
PS|142|2|et non intres in iudicio cum servo tuo quia non iustificabitur in conspectu tuo omnis vivens
PS|142|3|quia persecutus est inimicus animam meam humiliavit in terra vitam meam conlocavit me in obscuris sicut mortuos saeculi
PS|142|4|et anxiatus est super me spiritus meus in me turbatum est cor meum
PS|142|5|memor fui dierum antiquorum meditatus sum in omnibus operibus tuis in factis manuum tuarum meditabar
PS|142|6|expandi manus meas ad te anima mea sicut terra sine aqua tibi diapsalma
PS|142|7|velociter exaudi me Domine defecit spiritus meus non avertas faciem tuam a me et similis ero descendentibus in lacum
PS|142|8|auditam mihi fac mane misericordiam tuam quia in te speravi notam fac mihi viam in qua ambulem quia ad te levavi animam meam
PS|142|9|eripe me de inimicis meis Domine ad te confugi
PS|142|10|doce me facere voluntatem tuam quia Deus meus es tu spiritus tuus bonus deducet me in terra recta
PS|142|11|propter nomen tuum Domine vivificabis me in aequitate tua educes de tribulatione animam meam
PS|142|12|et in misericordia tua disperdes inimicos meos et perdes omnes qui tribulant animam meam quoniam ego servus tuus sum
PS|143|1|David adversus Goliad benedictus Dominus Deus meus qui docet manus meas ad proelium digitos meos ad bellum
PS|143|2|misericordia mea et refugium meum susceptor meus et liberator meus protector meus et in eo speravi qui subdis populum meum sub me
PS|143|3|Domine quid est homo quia innotuisti ei aut filius hominis quia reputas eum
PS|143|4|homo vanitati similis factus est dies eius sicut umbra praetereunt
PS|143|5|Domine inclina caelos tuos et descende tange montes et fumigabunt
PS|143|6|fulgora coruscationem et dissipabis eos emitte sagittas tuas et conturbabis eos
PS|143|7|emitte manum tuam de alto eripe me et libera me de aquis multis de manu filiorum alienorum
PS|143|8|quorum os locutum est vanitatem et dextera eorum dextera iniquitatis
PS|143|9|Deus canticum novum cantabo tibi in psalterio decacordo psallam tibi
PS|143|10|qui das salutem regibus qui redimit David servum suum de gladio maligno
PS|143|11|eripe me et eripe me de manu filiorum alienigenarum quorum os locutum est vanitatem et dextera eorum dextera iniquitatis
PS|143|12|quorum filii sicut novella plantationis in iuventute sua filiae eorum conpositae circumornatae ut similitudo templi
PS|143|13|promptuaria eorum plena eructantia ex hoc in illud oves eorum fetosae abundantes in egressibus suis
PS|143|14|boves eorum crassi non est ruina maceriae neque transitus neque clamor in plateis eorum
PS|143|15|beatum dixerunt populum cui haec sunt beatus populus cuius Dominus Deus eius
PS|144|1|laudatio David exaltabo te Deus meus rex et benedicam nomini tuo in saeculum et in saeculum saeculi
PS|144|2|per singulos dies benedicam tibi et laudabo nomen tuum in saeculum et in saeculum saeculi
PS|144|3|magnus Dominus et laudabilis nimis et magnitudinis eius non est finis
PS|144|4|generatio et generatio laudabit opera tua et potentiam tuam pronuntiabunt
PS|144|5|magnificentiam gloriae sanctitatis tuae loquentur et mirabilia tua narrabunt
PS|144|6|et virtutem terribilium tuorum dicent et magnitudinem tuam narrabunt
PS|144|7|memoriam abundantiae suavitatis tuae eructabunt et iustitia tua exultabunt
PS|144|8|miserator et misericors Dominus patiens et multum misericors
PS|144|9|suavis Dominus universis et miserationes eius super omnia opera eius
PS|144|10|confiteantur tibi Domine omnia opera tua et sancti tui confiteantur tibi
PS|144|11|gloriam regni tui dicent et potentiam tuam loquentur
PS|144|12|ut notam faciant filiis hominum potentiam tuam et gloriam magnificentiae regni tui
PS|144|13|regnum tuum regnum omnium saeculorum et dominatio tua in omni generatione et progenie fidelis Dominus in omnibus verbis suis et sanctus in omnibus operibus suis
PS|144|14|adlevat Dominus omnes qui corruunt et erigit omnes elisos
PS|144|15|oculi omnium in te sperant et tu das escam illorum in tempore oportuno
PS|144|16|aperis tu manum tuam et imples omne animal benedictione
PS|144|17|iustus Dominus in omnibus viis suis et sanctus in omnibus operibus suis
PS|144|18|prope est Dominus omnibus invocantibus eum omnibus invocantibus eum in veritate
PS|144|19|voluntatem timentium se faciet et deprecationem eorum exaudiet et salvos faciet eos
PS|144|20|custodit Dominus omnes diligentes se et omnes peccatores disperdet
PS|144|21|laudationem Domini loquetur os meum et benedicat omnis caro nomini sancto eius in saeculum et in saeculum saeculi
PS|145|1|alleluia Aggei et Zacchariae
PS|145|2|lauda anima mea Dominum laudabo Dominum in vita mea psallam Deo meo quamdiu fuero nolite confidere in principibus
PS|145|3|in filiis hominum quibus non est salus
PS|145|4|exibit spiritus eius et revertetur in terram suam in illa die peribunt omnes cogitationes eorum
PS|145|5|beatus cuius Deus Iacob adiutor eius spes eius in Domino Deo ipsius
PS|145|6|qui fecit caelum et terram mare et omnia quae in eis
PS|145|7|qui custodit veritatem in saeculum facit iudicium iniuriam patientibus dat escam esurientibus Dominus solvit conpeditos
PS|145|8|Dominus inluminat caecos Dominus erigit adlisos Dominus diligit iustos
PS|145|9|Dominus custodit advenas pupillum et viduam suscipiet et viam peccatorum disperdet
PS|145|10|regnabit Dominus in saecula Deus tuus Sion in generationem et generationem
PS|146|1|alleluia Aggei et Zacchariae laudate Dominum quoniam bonum psalmus Deo nostro sit iucunda decoraque; laudatio
PS|146|2|aedificans Hierusalem Dominus dispersiones Israhel congregabit
PS|146|3|qui sanat contritos corde et alligat contritiones illorum
PS|146|4|qui numerat multitudinem stellarum et omnibus eis nomina vocans
PS|146|5|magnus Dominus noster et magna virtus eius et sapientiae eius non est numerus
PS|146|6|suscipiens mansuetos Dominus humilians autem peccatores usque ad terram
PS|146|7|praecinite Domino in confessione psallite Deo nostro in cithara
PS|146|8|qui operit caelum nubibus et parat terrae pluviam qui producit in montibus faenum et herbam servituti hominum
PS|146|9|et dat iumentis escam ipsorum et pullis corvorum invocantibus eum
PS|146|10|non in fortitudine equi voluntatem habebit nec in tibiis viri beneplacitum erit ei
PS|146|11|beneplacitum est Domino super timentes eum et in eis qui sperant super misericordia eius
PS|147|1|alleluia lauda Hierusalem Dominum lauda Deum tuum Sion
PS|147|2|quoniam confortavit seras portarum tuarum benedixit filiis tuis in te
PS|147|3|qui posuit fines tuos pacem et adipe frumenti satiat te
PS|147|4|qui emittit eloquium suum terrae velociter currit sermo eius
PS|147|5|qui dat nivem sicut lanam nebulam sicut cinerem spargit
PS|147|6|mittit cristallum suum sicut buccellas ante faciem frigoris eius quis sustinebit
PS|147|7|emittet verbum suum et liquefaciet ea flabit spiritus eius et fluent aquae
PS|147|8|qui adnuntiat verbum suum Iacob iustitias et iudicia sua Israhel
PS|147|9|non fecit taliter omni nationi et iudicia sua non manifestavit eis
PS|148|1|alleluia laudate Dominum de caelis laudate eum in excelsis
PS|148|2|laudate eum omnes angeli eius laudate eum omnes virtutes eius
PS|148|3|laudate eum sol et luna laudate eum omnes stellae et lumen
PS|148|4|laudate eum caeli caelorum et aqua quae super caelum est
PS|148|5|laudent nomen Domini quia ipse dixit et facta sunt ipse mandavit et creata sunt
PS|148|6|statuit ea in saeculum et in saeculum saeculi praeceptum posuit et non praeteribit
PS|148|7|laudate Dominum de terra dracones et omnes abyssi
PS|148|8|ignis grando nix glacies spiritus procellarum quae faciunt verbum eius
PS|148|9|montes et omnes colles ligna fructifera et omnes cedri
PS|148|10|bestiae et universa pecora serpentes et volucres pinnatae
PS|148|11|reges terrae et omnes populi principes et omnes iudices terrae
PS|148|12|iuvenes et virgines senes cum iunioribus laudent nomen Domini
PS|148|13|quia exaltatum est nomen eius solius
PS|148|14|confessio eius super caelum et terram et exaltabit cornu populi sui hymnus omnibus sanctis eius filiis Israhel populo adpropinquanti sibi
PS|149|1|alleluia cantate Domino canticum novum laus eius in ecclesia sanctorum
PS|149|2|laetetur Israhel in eo qui fecit eum et filii Sion exultent in rege suo
PS|149|3|laudent nomen eius in choro in tympano et psalterio psallant ei
PS|149|4|quia beneplacitum est Domino in populo suo et exaltabit mansuetos in salute
PS|149|5|exultabunt sancti in gloria laetabuntur in cubilibus suis
PS|149|6|exaltationes Dei in gutture eorum et gladii ancipites in manibus eorum
PS|149|7|ad faciendam vindictam in nationibus increpationes in populis
PS|149|8|ad alligandos reges eorum in conpedibus et nobiles eorum in manicis ferreis
PS|149|9|ut faciant in eis iudicium conscriptum gloria haec est omnibus sanctis eius
PS|150|1|alleluia laudate Dominum in sanctis eius laudate eum in firmamento virtutis eius
PS|150|2|laudate eum in virtutibus eius laudate eum secundum multitudinem magnitudinis eius
PS|150|3|laudate eum in sono tubae laudate eum in psalterio et cithara
PS|150|4|laudate eum in tympano et choro laudate eum in cordis et organo
PS|150|5|laudate eum in cymbalis bene sonantibus laudate eum in cymbalis iubilationis
PS|150|6|omnis spiritus laudet Dominum
