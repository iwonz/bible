MAL|1|1|Пророцтво Господнього слова до Ізраїля через Малахію.
MAL|1|2|Я вас покохав, говорить Господь, а ви кажете: Як Ти нас покохав? Чи ж не брат Ісав Якову? каже Господь, а Я Якова був покохав,
MAL|1|3|а Ісава зненавидів, і зробив його гори спустошенням, а спадок його для шакалів пустині.
MAL|1|4|Коли скаже Едом: Ми зруйновані, та знову збудуємо руїни, то так промовляє Господь Саваот: Вони побудують, а Я розвалю! І звати їх будуть: Країна безбожности, і народ, на якого навіки розгнівавсь Господь!
MAL|1|5|І ваші очі побачать оце, і ви скажете: Стане великий Господь понад границю Ізраїлеву!
MAL|1|6|Шанує син батька, а раб свого пана; та якщо Я вам батько, де пошана Моя? А якщо Я вам пан, де страх передо Мною? говорить Господь Саваот вам, священики, що погорджуєте Моїм Іменням та й кажете: Чим ми погордили Йменням Твоїм?
MAL|1|7|На жертівник Мій ви приносите хліб занечищений і кажете: Чим Тебе ми зневажили? Тим, що кажете ви: Трапеза Господня вона погорджена!
MAL|1|8|І коли ви проносите в жертву сліпе, це не зле? І як кульгаве та хворе приносите, чи ж це не зле? Принеси но подібне своєму намісникові, чи тебе він вподобає, чи підійме обличчя твоє? промовляє Господь Саваот.
MAL|1|9|А тепер ублагайте ви Боже лице, і хай стане для нас милостивим. З ваших рук це було, то хіба кому з вас Він обличчя підійме? говорить Господь Саваот.
MAL|1|10|Нехай хто серед вас замкне двері святині, і не буде надармо освічувати Мого жертівника! Я не маю вподоби до вас, говорить Господь Саваот, і з ваших рук не вподобаю дару!
MAL|1|11|Бо від сходу сонця й аж по захід його звеличиться Ймення Моє між народами, і кадиться в кожному місці для Ймення Мого дар чистий, бо звеличиться Ймення Моє між народами, каже Господь Саваот.
MAL|1|12|Ви ж Його зневажаєте, кажучи: Трапеза Господня вона занечищена, й дохід її, обриджена страва її.
MAL|1|13|І до того говорите: Ось стільки праці! і ним нехтуєте, говорить Господь Саваот, і приносите крадене, і кульгаве та хворе, і таку жертву хлібну приносите. Чи буде воно Мені миле з рук ваших? говорить Господь.
MAL|1|14|І проклятий обманець, що в стаді його є самець, а він обіцяє та в жертву дає Господеві зіпсуте, а Я Цар великий, говорить Господь, і серед народів грізне Моє Ймення!
MAL|2|1|А тепер до вас заповідь цяя, священики!
MAL|2|2|Якщо ви не послухаєтесь, і не покладете на серце собі, щоб Іменню Моєму давати хвалу, говорить Господь Саваот, то пошлю Я прокляття на вас, і прокляну благословення ваші, і вже проклинаю, бо ви не берете до серця цього!
MAL|2|3|Ось Я обітну вам рамено, і розпорошу нечистість на ваших обличчях, нечистість свят ваших, і до неї вас винесуть.
MAL|2|4|І пізнаєте ви, що Я заповідь вам цю послав, щоб був заповіт Мій з Левієм, каже Господь Саваот.
MAL|2|5|Заповіт Мій з ним був для життя та для миру, і Я дав йому страх, і він налякався Мене, та боявсь перед Іменням Моїм.
MAL|2|6|Закон правди в устах його був, і не знайшлась на губах його кривда, у мирі й простоті ходив він зо Мною, і багато-кого відвернув від вини.
MAL|2|7|Бо уста священикові знання стережуть та Закона шукають із уст його, бо він Ангол Господа Саваота.
MAL|2|8|А ви відхилились з дороги, вчинили таке, що багато спіткнулись в Законі, Левієвого заповіта понищили, говорить Господь Саваот.
MAL|2|9|Тому то і Я вас зробив погорджуваними й низькими для всього народу, бо не стережете доріг Моїх ви, та не безсторонні в Законі.
MAL|2|10|Чи Отець нам усім не один? Хіба Бог не один нас створив? Чому ж один одного зраджуємо ми, щоб нам зневажати заповіт батьків наших?
MAL|2|11|Зраджує Юда, і робиться нечисть серед Ізраїля та в Єрусалимі, бо Юда зневажив святиню Господню, яку покохав був, і дочку бога чужого за жінку узяв.
MAL|2|12|Нехай Господь вигубить кожного, хто таке робить, того, хто чуває та відповідає з наметів Якова, і хто дар приносить Господу Саваоту.
MAL|2|13|І робите й друге таке: Господнього жертівника ви слізьми покриваєте, плачем та стогнанням, бо до дарів уже Він не звернеться більше, і милої жертви з рук ваших не візьме.
MAL|2|14|А ви ще й говорите: Защо? За те, що засвідчив Господь між тобою й жоною юнацтва твого, якій ти невірність вчинив, а вона ж твоя подруга, і дружина умови твоєї!
MAL|2|15|Хіба Бог не один нас учинив? І залишок духу Його. А що цей один? Насіння від Бога шукав. Тому свого духа пильнуйте, і дружину юнацтва свойого не зраджуйте!
MAL|2|16|Бо ненавиджу розвід, говорить Господь, Бог Ізраїлів, і того, хто вкриває насильством одежу свою, промовляє Господь Саваот. Тому свого духа пильнуйте, і не зраджуйте!
MAL|2|17|Словами своїми ви мучите Господа, та й питаєте ще: Чим ми мучимо? Говоренням вашим: Кожен, хто чинить лихе, той добрий у Господніх очах, і Він у них уподобання має, або: Де Бог правосуддя?
MAL|3|1|Ось Я посилаю Свого Ангола, і він перед обличчям Моїм приготує дорогу. І нагло прибуде до храму Свого Господь, Якого шукаєте ви, і Ангол заповіту, Якого жадаєте. Ось іде Він, говорить Господь Саваот!
MAL|3|2|І хто витерпить день Його прибуття, і хто встоїть, коли Він з'явиться? Бо Він, як огонь той у золотаря, і як у пральників луг.
MAL|3|3|І Він сяде топити та чистити срібло, і очистить синів Левія, і їх перечистить, як золото й срібло, і будуть для Господа жертву приносити в правді.
MAL|3|4|Тоді буде дар Юди та Єрусалиму приємний для Господа, як за днів віковічних і за років стародавніх.
MAL|3|5|І прибуду до вас Я на суд, і буду свідком швидким проти чарівників, і на перелюбників, і проти тих, хто присягу складає на лжу, і проти тих, хто заплатою наймита тисне, вдову й сироту, хто відхилює право чужинця, Мене ж не боїться, говорить Господь Саваот.
MAL|3|6|Бо Я, Господь, не змінююся, тому ви, сини Яковові, не будете знищені.
MAL|3|7|Від устав Моїх ви відступили з днів ваших батьків, і їх не стерегли. Верніться ж до Мене, і вернусь Я до вас! промовляє Господь Саваот. Та говорите ви: У чому повернемось?
MAL|3|8|Чи Бога людина обманить? Мене ж ви обманюєте, ще й говорите: Чим ми Тебе обманили? Десятиною та приносами!
MAL|3|9|Прокляттям ви прокляті, а Мене обманили, о люду ти ввесь!
MAL|3|10|Принесіть же ви всю десятину до дому скарбниці, щоб страва була в Моїм храмі, і тим Мене випробуйте, промовляє Господь Саваот: чи небесних отворів вам не відчиню, та не виллю вам благословення аж надмір?
MAL|3|11|І ради вас насварю Я все те, що жере, і воно не понищить вам земного плоду, і не заб'є винограду вам на полі, говорить Господь Саваот.
MAL|3|12|І будуть всі люди вважати вас блаженними, бо будете ви любим Краєм, говорить Господь Саваот.
MAL|3|13|Жорсткі ваші слова проти Мене, говорить Господь, а ви кажете: Що ми на Тебе сказали?
MAL|3|14|Ви кажете: Марність служити для Бога! І що за користь, що ми стережемо Його службу, та ходимо в жалобі перед лицем Господа Саваота?
MAL|3|15|А тепер ми вважаємо пишних щасливими, і ті, хто вчиняє безбожне, будуються та випробовують Бога, і втікають...
MAL|3|16|Змовлялись тоді один з одним і ті, хто страх перед Господом має, і прислухавсь Господь, і почув, і перед обличчям Його була писана пам'ятна книга про тих, хто страх перед Господом має, і хто поважає Ймення Його.
MAL|3|17|І будуть Мені вони власністю, каже Господь Саваот, на той день, що вчиню, і змилосерджусь над ними, як змилосерджується чоловік над синами своїми, що служать йому.
MAL|3|18|І ви знову побачите різне між праведним та нечестивим, між тим, хто Богові служить, та тим, хто не служить Йому.
MAL|4|1|Бо ось наступає той день, що палає, як піч, і стануть всі пишні та кожен, хто чинить безбожне, соломою, і спалить їх день той, який наступає, говорить Господь Саваот, Який не позоставить їм кореня, ані галузки.
MAL|4|2|А для вас, хто Ймення Мойого боїться, зійде Сонце Правди та лікування в промінях Його, і ви вийдете та поскакаєте, мов ті ситі телята!
MAL|4|3|І безбожних топтати ви будете, бо стануть за попіл вони під п'ятами ніг ваших у той день, що його Я вчиню, промовляє Господь Саваот.
MAL|4|4|Згадайте Закона Мойсея, Мого раба, що йому наказав на Хориві устави й права щодо всього Ізраїля.
MAL|4|5|Ось Я пошлю вам пророка Іллю, перше ніж день Господній настане, великий й страшний!
MAL|4|6|І приверне він серце батьків до синів, і серце синівське до їхніх батьків, щоб Я не прийшов, і не вразив цей Край прокляттям!
