GEN|1|1|起初，上帝創造天地。
GEN|1|2|地是空虛混沌，深淵上面一片黑暗；上帝的靈 運行在水面上。
GEN|1|3|上帝說：「要有光」，就有了光。
GEN|1|4|上帝看光是好的，於是上帝就把光和暗分開。
GEN|1|5|上帝稱光為「晝」，稱暗為「夜」。有晚上，有早晨，這是第一日。
GEN|1|6|上帝說：「眾水之間要有穹蒼，把水和水分開。」
GEN|1|7|上帝就造了穹蒼，把穹蒼以下的水和穹蒼以上的水分開。事就這樣成了。
GEN|1|8|上帝稱穹蒼為「天」。有晚上，有早晨，這是第二日。
GEN|1|9|上帝說：「天下面的水要聚集在一處，使乾地露出來。」事就這樣成了。
GEN|1|10|上帝稱乾地為「地」，稱聚集在一起的水為「海」。上帝看為好的。
GEN|1|11|上帝說：「地要長出植物，就是含種子的五穀菜蔬，和會結果子、果子裏有種子的樹，在地上各從其類。」事就這樣成了。
GEN|1|12|於是地長出了植物：含種子的五穀菜蔬，各從其類；會結果子、果子裏有種子的樹，各從其類。上帝看為好的。
GEN|1|13|有晚上，有早晨，這是第三日。
GEN|1|14|上帝說：「天上要有光體來分晝夜，讓它們作記號，定季節、日子、年份，
GEN|1|15|它們要在天空發光，照在地上。」事就這樣成了。
GEN|1|16|於是上帝造了兩個大光體，大的管晝，小的管夜，又造了星辰。
GEN|1|17|上帝把這些光體擺列在天空，照在地上，
GEN|1|18|管理晝夜，分別光暗。上帝看為好的。
GEN|1|19|有晚上，有早晨，這是第四日。
GEN|1|20|上帝說：「水要滋生眾多有生命之物；要有鳥飛在地面以上，天空之中。」
GEN|1|21|上帝就創造了大魚和在水裏滋生的各樣活動的生物，各從其類，以及各樣有翅膀的鳥，各從其類。上帝看為好的。
GEN|1|22|上帝就賜福給這一切，說：「要繁殖增多，充滿在海的水裏；飛鳥也要在地上增多。」
GEN|1|23|有晚上，有早晨，這是第五日。
GEN|1|24|上帝說：「地要生出有生命之物，各從其類，就是牲畜、爬行動物、地上的走獸，各從其類。」事就這樣成了。
GEN|1|25|於是上帝造了地上的走獸，各從其類；牲畜，各從其類；和地上一切的爬行動物，各從其類。上帝看為好的。
GEN|1|26|上帝說：「我們要照著我們的形像，按著我們的樣式造人，使他們管理海裏的魚、天空的鳥、地上的牲畜和全地，以及地上爬的一切爬行動物。」
GEN|1|27|上帝就照著他的形像創造人，照著上帝的形像創造他們 ；他創造了他們，有男有女。
GEN|1|28|上帝賜福給他們，上帝對他們說：「要生養眾多，遍滿這地，治理它；要管理海裏的魚、天空的鳥和地上各樣活動的生物。」
GEN|1|29|上帝說：「看哪，我把全地一切含種子的五穀菜蔬和一切會結果子、果子裏有種子的樹，都賜給你們；這些都可作食物。
GEN|1|30|至於地上一切的走獸、天空一切的飛鳥，並一切在地上爬行的，有生命的動物，我把綠色植物賜給牠們作食物。」事就這樣成了。
GEN|1|31|上帝看一切所造的，看哪，都非常好。有晚上，有早晨，這是第六日。
GEN|2|1|天和地，以及萬象都完成了。
GEN|2|2|到第七日，上帝已經完成了造物之工，就在第七日安息了，歇了他所做一切的工。
GEN|2|3|上帝賜福給第七日，將它分別為聖，因為在這日，上帝安息了，歇了他所做一切創造的工。
GEN|2|4|這就是天地創造的來歷。 在耶和華上帝造地和天的時候，
GEN|2|5|地上還沒有田野的草木，田間的菜蔬還沒有長出來，因為耶和華上帝還沒有降雨在地上，也沒有人耕種土地。
GEN|2|6|但是，有霧氣從地上騰，滋潤整個土地的表面。
GEN|2|7|耶和華上帝用地上的塵土造人，將生命之氣吹進他的鼻孔，這人就成了有靈的活人 。
GEN|2|8|耶和華上帝在東方的 伊甸 栽了一個園子，把所造的人安置在那裏。
GEN|2|9|耶和華上帝使各樣的樹從土地裏長出來，可以悅人的眼目，好作食物。園子當中有生命樹和知善惡的樹 。
GEN|2|10|有一條河從 伊甸 流出來，滋潤那園子，從那裏分成四個源頭：
GEN|2|11|第一條名叫 比遜 ，它環繞 哈腓拉 全地，在那裏有金子。
GEN|2|12|那地的金子很好，在那裏也有珍珠 和紅瑪瑙。
GEN|2|13|第二條河名叫 基訓 ，它環繞 古實 全地。
GEN|2|14|第三條河名叫 底格里斯 ，它流到 亞述 的東邊。第四條河就是 幼發拉底 。
GEN|2|15|耶和華上帝把那人安置在 伊甸園 ，讓他耕耘看管。
GEN|2|16|耶和華上帝吩咐那人說：「園中各樣樹上所出的，你可以隨意吃，
GEN|2|17|只是知善惡的樹所出的，你不可吃，因為你吃它的日子必定死！」
GEN|2|18|耶和華上帝說：「那人單獨一個不好，我要為他造一個配偶幫助他。」
GEN|2|19|耶和華上帝用泥土造了野地各樣的走獸和天空各樣的飛鳥，都帶到那人面前，看他叫甚麼。那人怎樣叫各樣的動物，那就是牠的名字。
GEN|2|20|那人就給一切牲畜、天空的飛鳥和野地各樣的走獸都起了名。只是 亞當 沒有找到配偶幫助他。
GEN|2|21|耶和華上帝使他沉睡，他就睡了；於是取下他的一根肋骨，又在原處把肉合起來。
GEN|2|22|耶和華上帝就用那人身上所取的肋骨造了一個女人，帶她到那人面前。
GEN|2|23|那人說： 「這正是我骨中的骨， 肉中的肉， 可以稱她為女人， 因為她是從男人身上取出來的。」
GEN|2|24|因此，人要離開父母，與妻子結合，二人成為一體。
GEN|2|25|當時夫妻二人赤身露體，並不覺得羞恥。
GEN|3|1|耶和華上帝所造的，惟有蛇比田野一切的走獸更狡猾。蛇對女人說：「上帝豈是真說，你們不可吃園中任何樹上所出的嗎？」
GEN|3|2|女人對蛇說：「園中樹上的果子，我們都可以吃；
GEN|3|3|只是園子中間那棵樹的果子，上帝曾說：『你們不可吃，也不可摸，免得你們死。』」
GEN|3|4|蛇對女人說：「你們不一定死；
GEN|3|5|因為上帝知道，你們吃的日子眼睛就開了，你們就像上帝一樣知道善惡。」
GEN|3|6|於是女人見那棵樹好作食物，又悅人的眼目，那樹令人喜愛，能使人有智慧，她就摘下果子吃了，又給了與她一起的丈夫，他也吃了。
GEN|3|7|他們二人的眼睛就開了，知道自己赤身露體，就編織無花果樹的葉子，為自己做成裙子。
GEN|3|8|天起了涼風，那人和他妻子聽見耶和華上帝在園中來回行走的聲音，就藏在園裏的樹木中，躲避耶和華上帝的面。
GEN|3|9|耶和華上帝呼喚那人，對他說：「你在哪裏？」
GEN|3|10|他說：「我在園中聽見你的聲音，我就害怕；因為我赤身露體，我就藏了起來。」
GEN|3|11|耶和華上帝說：「誰告訴你，你是赤身露體呢？莫非你吃了那樹上所出的，就是我吩咐你不可吃的嗎？」
GEN|3|12|那人說：「你賜給我、與我一起的女人，是她把那樹上所出的給我，我就吃了。」
GEN|3|13|耶和華上帝對女人說：「你怎麼會做這種事呢？」女人說：「那蛇引誘我，我就吃了。」
GEN|3|14|耶和華上帝對蛇說： 「你既做了這事，就必受詛咒， 比一切的牲畜和野獸更重。 你必用肚子行走， 終生吃土。
GEN|3|15|我要使你和女人彼此為仇， 你的後裔和女人的後裔也彼此為仇。 他要傷你的頭， 你要傷他的腳跟。 」
GEN|3|16|又對女人說： 「我必多多加增你懷胎的痛苦， 你生兒女時必多受痛苦。 你必戀慕你丈夫， 他必管轄你。」
GEN|3|17|又對 亞當 說： 「你既聽從你妻子的話， 吃了那樹上所出的， 就是我吩咐你不可吃的， 土地必因你的緣故受詛咒； 你必終生勞苦才能從土地得吃的。
GEN|3|18|土地必給你長出荊棘和蒺藜來； 你也要吃田間的五穀菜蔬。
GEN|3|19|你必汗流滿面才有食物可吃， 直到你歸了土地， 因為你是從土地而出的。 你本是塵土，仍要歸回塵土。」
GEN|3|20|那人給他妻子起名叫 夏娃 ，因為她是眾生之母 。
GEN|3|21|耶和華上帝用獸皮做衣服給 亞當 和他的妻子穿。
GEN|3|22|耶和華上帝說：「看哪，那人已經像我們中間的一個，知道善惡，現在恐怕他又伸手摘生命樹所出的來吃，就永遠活著。」
GEN|3|23|耶和華上帝就驅逐他出 伊甸園 ，使他耕種土地，他原是從土地裏被取出來的。
GEN|3|24|耶和華上帝把那人趕出去，就在 伊甸園 東邊安設基路伯和發出火焰轉動的劍，把守生命樹的道路。
GEN|4|1|那人和他妻子 夏娃 同房， 夏娃 就懷孕，生了 該隱 ，她說：「我靠耶和華得了一個男的。」
GEN|4|2|她又生了 該隱 的弟弟 亞伯 。 亞伯 是牧羊的； 該隱 是耕地的。
GEN|4|3|過了一些日子， 該隱 拿地裏的出產為供物獻給耶和華；
GEN|4|4|亞伯 也把他羊群中頭生的和羊的脂肪獻上。耶和華看中了 亞伯 和他的供物，
GEN|4|5|卻看不中 該隱 和他的供物。 該隱 就非常生氣，沉下臉來。
GEN|4|6|耶和華對 該隱 說：「你為甚麼生氣呢？你為甚麼沉下臉來呢？
GEN|4|7|你若做得對，豈不仰起頭來嗎？你若做得不對，罪就伏在門前。它想要控制你，你卻要制伏它。」
GEN|4|8|該隱 與他弟弟 亞伯 說話 。 二人正在田間時， 該隱 起來攻擊他弟弟 亞伯 ，把他殺了。
GEN|4|9|耶和華對 該隱 說：「你弟弟 亞伯 在哪裏？」他說：「我不知道！我豈是看守我弟弟的嗎？」
GEN|4|10|耶和華說：「你做了甚麼事呢？你弟弟血的聲音從地裏向我哀號。
GEN|4|11|現在你必從這地受詛咒，這地開了口，從你手裏接受你弟弟的血。
GEN|4|12|你耕種土地，它不再給你效力；你必流離飄蕩在地上。」
GEN|4|13|該隱 對耶和華說：「我的懲罰太重，過於我所能承當的。
GEN|4|14|看哪，今日你趕我離開這塊土地，不能見你的面；我必流離飄蕩在地上，凡遇見我的必殺我。」
GEN|4|15|耶和華對他說：「既然如此 ，凡殺 該隱 的，必遭報七倍。」耶和華就給 該隱 立一個記號，免得人遇見他就殺他。
GEN|4|16|於是 該隱 離開了耶和華的面，去住在 伊甸 東邊 挪得 之地。
GEN|4|17|該隱 與妻子同房，她就懷孕，生了 以諾 。 該隱 建造一座城，就照他兒子的名字稱那城為 以諾 。
GEN|4|18|以諾 生 以拿 ， 以拿 生 米戶雅利 ， 米戶雅利 生 瑪土撒利 ， 瑪土撒利 生 拉麥 。
GEN|4|19|拉麥 娶了兩個妻子：一個名叫 亞大 ，一個名叫 洗拉 。
GEN|4|20|亞大 生 雅八 ； 雅八 是住帳棚、牧養牲畜之人的祖師。
GEN|4|21|雅八 的兄弟名叫 猶八 ；他是所有彈琴吹簫之人的祖師。
GEN|4|22|洗拉 又生了 土八‧該隱 ；他是打造各樣銅器鐵器的工匠。 土八‧該隱 的妹妹是 拿瑪 。
GEN|4|23|拉麥 對他兩個妻子說： 亞大 、 洗拉 啊，聽我的聲音； 拉麥 的妻子啊，側耳聽我的言語： 大人傷我，我把他殺了； 小孩損我，我把他害了 。
GEN|4|24|若殺 該隱 ，遭報七倍， 殺 拉麥 的，必遭報七十七倍。
GEN|4|25|亞當 又與妻子同房，她就生了一個兒子，給他起名叫 塞特 ，說：「上帝給我立了另一個子嗣代替 亞伯 ，因為 該隱 殺了他。」
GEN|4|26|塞特 也生了一個兒子，起名叫 以挪士 。那時候，人開始求告耶和華的名。
GEN|5|1|這是 亞當 後代的家譜。當上帝造人的日子，他照著自己的樣式造人。
GEN|5|2|他造男造女。在他們被造的日子，上帝賜福給他們，稱他們為人。
GEN|5|3|亞當 活到一百三十歲，生了一個兒子，形像樣式和自己相似，就給他起名叫 塞特 。
GEN|5|4|亞當 生 塞特 之後，又活了八百年，並且生兒育女。
GEN|5|5|亞當 共活了九百三十年，就死了。
GEN|5|6|塞特 活到一百零五歲，生了 以挪士 。
GEN|5|7|塞特 生 以挪士 之後，又活了八百零七年，並且生兒育女。
GEN|5|8|塞特 共活了九百一十二年，就死了。
GEN|5|9|以挪士 活到九十歲，生了 該南 。
GEN|5|10|以挪士 生 該南 之後，又活了八百一十五年，並且生兒育女。
GEN|5|11|以挪士 共活了九百零五年，就死了。
GEN|5|12|該南 活到七十歲，生了 瑪勒列 。
GEN|5|13|該南 生 瑪勒列 之後，又活了八百四十年，並且生兒育女。
GEN|5|14|該南 共活了九百一十年，就死了。
GEN|5|15|瑪勒列 活到六十五歲，生了 雅列 。
GEN|5|16|瑪勒列 生 雅列 之後，又活了八百三十年，並且生兒育女。
GEN|5|17|瑪勒列 共活了八百九十五年，就死了。
GEN|5|18|雅列 活到一百六十二歲，生了 以諾 。
GEN|5|19|雅列 生 以諾 之後，又活了八百年，並且生兒育女。
GEN|5|20|雅列 共活了九百六十二年，就死了。
GEN|5|21|以諾 活到六十五歲，生了 瑪土撒拉 。
GEN|5|22|以諾 生 瑪土撒拉 之後，與上帝同行三百年，並且生兒育女。
GEN|5|23|以諾 共活了三百六十五年。
GEN|5|24|以諾 與上帝同行，上帝把他接去，他就不在了。
GEN|5|25|瑪土撒拉 活到一百八十七歲，生了 拉麥 。
GEN|5|26|瑪土撒拉 生 拉麥 之後，又活了七百八十二年，並且生兒育女。
GEN|5|27|瑪土撒拉 共活了九百六十九年，就死了。
GEN|5|28|拉麥 活到一百八十二歲，生了一個兒子，
GEN|5|29|給他起名叫 挪亞 ，說：「在耶和華所詛咒的地上，這個兒子必使我們從工作和手中的勞苦得到安慰。」
GEN|5|30|拉麥 生 挪亞 之後，又活了五百九十五年，並且生兒育女。
GEN|5|31|拉麥 共活了七百七十七年，就死了。
GEN|5|32|挪亞 活到五百歲，生了 閃 、 含 和 雅弗 。
GEN|6|1|當人開始在地面上增多、又生女兒的時候，
GEN|6|2|上帝的兒子們看見人的女子美貌，就隨意挑選，娶來為妻。
GEN|6|3|耶和華說：「人既屬乎血氣，我的靈就不永遠住在他裏面；然而他的年歲還可到一百二十年。」
GEN|6|4|那時候有巨人在地上，後來也有；上帝的兒子們和人的女子們交合，生了孩子。那些人就是古代的勇士，有名的人物。
GEN|6|5|耶和華見人在地上罪大惡極，終日心裏所想的盡都是惡事，
GEN|6|6|耶和華就因造人在地上感到遺憾，心中憂傷。
GEN|6|7|耶和華說：「我要把所造的人和走獸，爬行動物，以及天空的飛鳥，都從地面上除滅，因為我造了他們感到遺憾。」
GEN|6|8|只有 挪亞 在耶和華眼前蒙恩。
GEN|6|9|這是 挪亞 的後代。 挪亞 是個義人，在他的世代中是個完全人。 挪亞 與上帝同行。
GEN|6|10|挪亞 生了三個兒子，就是 閃 、 含 和 雅弗 。
GEN|6|11|這地在上帝面前敗壞了，地上充滿了暴力。
GEN|6|12|上帝觀看這地，看哪，它敗壞了，因為凡血肉之軀在地上的行為都敗壞了。
GEN|6|13|上帝對 挪亞 說：「在我面前，凡血肉之軀的結局已經臨到，因著他們，地上充滿了暴力。看哪，我要把他們和這地一起毀滅。
GEN|6|14|你要為自己用歌斐木造一艘方舟，並在方舟內造房間，內外都要抹上瀝青。
GEN|6|15|方舟的造法是這樣：要長三百肘，寬五十肘，高三十肘。
GEN|6|16|方舟上面要造天窗，向上一肘。方舟的門要開在旁邊。方舟要分上、中、下三層。
GEN|6|17|看哪，我要使洪水氾濫在地上，毀滅天下凡有生命氣息的血肉之軀，地上的一切都要滅亡。
GEN|6|18|但我要與你立約；你同你的兒子、妻子和媳婦都要進入方舟。
GEN|6|19|凡有血肉的動物，每樣一對，一公一母，你要帶進方舟，好跟你一起保全生命。
GEN|6|20|飛鳥各從其類，牲畜各從其類，地上的爬行動物各從其類，每樣一對，都要到你那裏，好保全生命。
GEN|6|21|你要拿各樣可吃的食物，儲存在你那裏，作你和牠們的糧食。」
GEN|6|22|挪亞 就去做了；凡上帝吩咐他的，他都照樣去做。
GEN|7|1|耶和華對 挪亞 說：「你和你的全家都要進入方舟，因為在這世代中，我看你在我面前是個義人。
GEN|7|2|凡潔淨的牲畜，你要各取七公七母；不潔淨的牲畜，你要各取一公一母；
GEN|7|3|天空的飛鳥也要各取七公七母，為了要留種，活在全地面上。
GEN|7|4|因為再過七天，我要降雨在地上四十晝夜，把我所造的一切生物從地面上除滅。」
GEN|7|5|挪亞 就遵照耶和華吩咐他的去做。
GEN|7|6|當洪水 在地上氾濫的時候， 挪亞 已六百歲。
GEN|7|7|挪亞 同他的兒子、妻子和媳婦都進入方舟，躲避洪水。
GEN|7|8|潔淨的牲畜和不潔淨的牲畜，飛鳥及所有爬行在土地上的，
GEN|7|9|都一對一對，有公有母，到 挪亞 那裏，進入方舟，正如上帝所吩咐 挪亞 的。
GEN|7|10|過了七天，洪水氾濫在地上。
GEN|7|11|挪亞 六百歲那一年的二月十七日，就在那一天，大深淵的泉源都裂開，天上的窗戶也敞開了，
GEN|7|12|四十晝夜有大雨降在地上。
GEN|7|13|正在那日， 挪亞 和他的兒子 閃 、 含 、 雅弗 ，以及 挪亞 的妻子和三個媳婦，都一同進入方舟。
GEN|7|14|他們和一切走獸，各從其類；一切牲畜，各從其類；地上爬的一切爬行動物，各從其類；一切的鳥，就是一切有翅膀的飛禽，各從其類；
GEN|7|15|凡有生命氣息的血肉之軀，都一對一對到 挪亞 那裏，進入方舟。
GEN|7|16|凡有血肉的，都一公一母進入方舟，正如上帝所吩咐 挪亞 的。耶和華就把他關在方舟裏。
GEN|7|17|洪水在地上氾濫四十天，水往上漲，使方舟浮起，方舟就從地上漂起來。
GEN|7|18|水勢洶湧，在地上大大上漲，方舟在水面上漂蕩。
GEN|7|19|水勢在地上極其浩大，普天下所有的高山都淹沒了。
GEN|7|20|水勢洶湧，比山高出十五肘 ，山嶺都淹沒了。
GEN|7|21|凡有血肉在地上行動的，就是飛鳥、牲畜、走獸和地上成群的群聚動物，以及所有的人，都死了。
GEN|7|22|在乾地上凡鼻孔裏有生命氣息的都死了。
GEN|7|23|耶和華除滅了地面上各類的生物，包括人和牲畜、爬行動物，以及天空的飛鳥；他們就都從地上除滅了，只剩下 挪亞 和那些與他同在方舟裏的。
GEN|7|24|水勢洶湧，在地上共一百五十天。
GEN|8|1|上帝記念 挪亞 和 挪亞 方舟裏的一切走獸牲畜。上帝使風吹地，水勢漸落。
GEN|8|2|深淵的泉源和天上的窗戶都關閉了，雨不再從天降下。
GEN|8|3|水從地上逐漸消退。過了一百五十天，水就退了。
GEN|8|4|七月十七日，方舟停在 亞拉臘山 上。
GEN|8|5|水繼續退去，直到十月；十月初一，山頂都露出來了。
GEN|8|6|過了四十天， 挪亞 打開他所造的方舟的窗戶，
GEN|8|7|放出一隻烏鴉。那烏鴉飛來飛去，直到地上的水都乾了。
GEN|8|8|他又從他那裏放出一隻鴿子，要看水從地面上退了沒有。
GEN|8|9|但全地面都是水，鴿子找不到落腳之地，就回到方舟 挪亞 那裏。 挪亞 伸手接了鴿子，把牠帶進方舟。
GEN|8|10|挪亞 又另外等了七天，再把鴿子從方舟放出去。
GEN|8|11|到了晚上，鴿子回到他那裏，看哪，嘴裏有一片剛啄下來的橄欖葉， 挪亞 就知道水已經從地上退了。
GEN|8|12|他又另外等了七天，再放出鴿子，這次鴿子不再回到他那裏了。
GEN|8|13|當 挪亞 六百零一歲，正月初一的時候，地上的水都乾了。 挪亞 打開方舟的蓋觀看，看哪，地面乾了。
GEN|8|14|到了二月二十七日，地就都乾了。
GEN|8|15|上帝對 挪亞 說：
GEN|8|16|「你同你的妻子、兒子、媳婦都要出方舟。
GEN|8|17|凡與你一起有血肉的生物，就是飛鳥、牲畜和地上爬的一切爬行動物，都要帶出來。 牠們要在地上滋生，繁殖增多。」
GEN|8|18|於是 挪亞 同他的兒子、妻子、媳婦都出來了。
GEN|8|19|一切走獸、爬行動物和飛鳥，地上所有的動物，各從其類，也都出了方舟。
GEN|8|20|挪亞 為耶和華築了一座壇，拿各種潔淨的牲畜和各種潔淨的飛鳥，獻在壇上為燔祭。
GEN|8|21|耶和華聞了那馨香之氣，耶和華心裏說：「我不再因人的緣故詛咒土地，因為人從幼年就心裏懷著惡念；我也不再照我曾做的毀滅一切生物了。
GEN|8|22|地還存在的時候，撒種、收割、寒暑、冬夏、晝夜都永不止息。」
GEN|9|1|上帝賜福給 挪亞 和他的兒子，對他們說：「你們要生養眾多，遍滿這地。
GEN|9|2|地上一切的走獸、天空一切的飛鳥、所有爬行在土地上的和海裏一切的魚都必怕你們，畏懼你們，牠們都要交在你們手裏。
GEN|9|3|凡活的動物都可作你們的食物。這一切我都賜給你們，如同綠色的菜蔬一樣。
GEN|9|4|只是帶著生命的肉，就是帶著血的，你們不可吃。
GEN|9|5|流你們血、害你們命的，我必向他追討；我要向一切走獸追討，向人和向人的弟兄追討人命。
GEN|9|6|凡流人血的，他的血也必被人所流，因為上帝造人，是照自己的形像造的。
GEN|9|7|你們要生養眾多，在地上繁衍昌盛。」
GEN|9|8|上帝對 挪亞 和同他一起的兒子說：
GEN|9|9|「看哪，我要與你們和你們後裔立我的約，
GEN|9|10|包括和你們一起所有的生物，就是飛鳥、牲畜、地上一切的走獸，凡從方舟裏出來地上一切的生物。
GEN|9|11|我與你們立我的約：凡有血肉的，不再被洪水滅絕，也不再有洪水毀壞這地了。」
GEN|9|12|上帝說：「這是我與你們，以及和你們一起的一切生物所立之約的記號，直到萬代：
GEN|9|13|我把彩虹放在雲中，這就是我與地立約的記號了。
GEN|9|14|我使雲遮地的時候，會有彩虹出現在雲中，
GEN|9|15|我就記念我與你們，以及各樣有血肉的生物所立的約：不再有洪水氾濫去毀滅一切有血肉的了。
GEN|9|16|彩虹出現在雲中，我看見了，就要記念上帝與地上一切有血肉的生物所立的永約。」
GEN|9|17|上帝對 挪亞 說：「這就是我與地上一切有血肉的立約的記號。」
GEN|9|18|挪亞 的兒子，從方舟出來的，有 閃 、 含 和 雅弗 。 含 是 迦南 的父親。
GEN|9|19|這是 挪亞 的三個兒子，他們的後裔散佈全地。
GEN|9|20|挪亞 是農夫，是他開始栽葡萄園的。
GEN|9|21|他喝了一些酒就醉了，在他的帳棚裏赤著身子。
GEN|9|22|迦南 的父親 含 看見他父親赤身，就到外面告訴他的兩個兄弟。
GEN|9|23|於是 閃 和 雅弗 拿了外衣搭在二人肩上，倒退著進去，遮蓋父親的赤身；他們背著臉，看不見父親的赤身。
GEN|9|24|挪亞 酒醒以後，知道小兒子向他所做的事，
GEN|9|25|就說： 「 迦南 當受詛咒， 必給他弟兄作奴僕的奴僕。」
GEN|9|26|又說： 「耶和華— 閃 的上帝是應當稱頌的！ 願 迦南 作 閃 的奴僕。
GEN|9|27|願上帝使 雅弗 擴張， 願他住在 閃 的帳棚裏； 願 迦南 作他的奴僕。」
GEN|9|28|洪水以後， 挪亞 又活了三百五十年。
GEN|9|29|挪亞 共活了九百五十年，就死了。
GEN|10|1|這是 挪亞 的兒子 閃 、 含 、 雅弗 的後代。洪水以後，他們都生了兒子。
GEN|10|2|雅弗 的兒子是 歌篾 、 瑪各 、 瑪代 、 雅完 、 土巴 、 米設 、 提拉 。
GEN|10|3|歌篾 的兒子是 亞實基拿 、 利法 、 陀迦瑪 。
GEN|10|4|雅完 的兒子是 以利沙 、 他施 、 基提 、 羅單 人 。
GEN|10|5|從這些人中有沿海國家的人散居各處，有自己的土地，各有各的語言、宗族、國家。
GEN|10|6|含 的兒子是 古實 、 麥西 、 弗 、 迦南 。
GEN|10|7|古實 的兒子是 西巴 、 哈腓拉 、 撒弗他 、 拉瑪 、 撒弗提迦 。 拉瑪 的兒子是 示巴 、 底但 。
GEN|10|8|古實 又生 寧錄 ，他是地上第一個勇士。
GEN|10|9|他在耶和華面前是個英勇的獵人，所以有話說：「像 寧錄 在耶和華面前是個英勇的獵人。」
GEN|10|10|他王國的開始是在 巴別 、 以力 、 亞甲 、 甲尼 ，都在 示拿 地。
GEN|10|11|他從那地出來往 亞述 去，建造了 尼尼微 、 利河伯 、 迦拉 ，
GEN|10|12|以及 尼尼微 和 迦拉 之間的 利鮮 ，那是座大城。
GEN|10|13|麥西 生 路低 人、 亞拿米 人、 利哈比 人、 拿弗土希 人、
GEN|10|14|帕斯魯細 人、 迦斯路希 人、 迦斐託 人； 非利士 人是從 迦斐託 人 出來的。
GEN|10|15|迦南 生了長子 西頓 ，又生 赫
GEN|10|16|和 耶布斯 人、 亞摩利 人、 革迦撒 人、
GEN|10|17|希未 人、 亞基 人、 西尼 人、
GEN|10|18|亞瓦底 人、 洗瑪利 人、 哈馬 人，後來 迦南 的家族散開了。
GEN|10|19|迦南 的疆界是從 西頓 到 基拉耳 ，直到 迦薩 ，又到 所多瑪 、 蛾摩拉 、 押瑪 、 洗扁 ，直到 拉沙 。
GEN|10|20|這就是 含 的後裔，各有自己的宗族、語言、土地和國家。
GEN|10|21|閃 也生了兒子，他是 雅弗 的哥哥 ，是 希伯 人的祖先。
GEN|10|22|閃 的兒子是 以攔 、 亞述 、 亞法撒 、 路德 、 亞蘭 。
GEN|10|23|亞蘭 的兒子是 烏斯 、 戶勒 、 基帖 、 瑪施 。
GEN|10|24|亞法撒 生 沙拉 ， 沙拉 生 希伯 。
GEN|10|25|希伯 生了兩個兒子，一個名叫 法勒 ，因為那時人分地居住； 法勒 的兄弟名叫 約坍 。
GEN|10|26|約坍 生 亞摩答 、 沙列 、 哈薩瑪非 、 耶拉 、
GEN|10|27|哈多蘭 、 烏薩 、 德拉 、
GEN|10|28|俄巴路 、 亞比瑪利 、 示巴 、
GEN|10|29|阿斐 、 哈腓拉 、 約巴 ，這些都是 約坍 的兒子。
GEN|10|30|他們所住的地方是從 米沙 直到 西發 ，到東邊的山。
GEN|10|31|這就是 閃 的後裔，各有自己的宗族、語言、土地和國家。
GEN|10|32|這些是 挪亞 兒子的宗族，按著他們的後代立國。洪水以後，邦國就從他們散佈在地上。
GEN|11|1|那時，全地只有一種語言，都說一樣的話。
GEN|11|2|他們向東遷移的時候，在 示拿 地找到一片平原，就住在那裏。
GEN|11|3|他們彼此商量說：「來，讓我們來做磚，把磚燒透了。」他們就拿磚當石頭，又拿柏油當泥漿。
GEN|11|4|他們說：「來，讓我們建造一座城和一座塔，塔頂通天。我們要為自己立名，免得我們分散在全地面上。」
GEN|11|5|耶和華降臨，要看世人所建造的城和塔。
GEN|11|6|耶和華說：「看哪，他們成了同一個民族，都有一樣的語言。這只是他們開始做的事，現在他們想要做的任何事，就沒有甚麼可攔阻他們了。
GEN|11|7|來，我們下去，在那裏變亂他們的語言，使他們彼此語言不通。」
GEN|11|8|於是耶和華使他們從那裏分散在全地面上；他們就停止建造那城了。
GEN|11|9|因為耶和華在那裏變亂了全地的語言，把人從那裏分散在全地面上，所以那城名叫 巴別 。
GEN|11|10|這是 閃 的後代。洪水以後二年， 閃 一百歲生了 亞法撒 。
GEN|11|11|閃 生 亞法撒 之後又活了五百年，並且生兒育女。
GEN|11|12|亞法撒 活到三十五歲，生了 沙拉 。
GEN|11|13|亞法撒 生 沙拉 之後又活了四百零三年，並且生兒育女。
GEN|11|14|沙拉 活到三十歲，生了 希伯 。
GEN|11|15|沙拉 生 希伯 之後又活了四百零三年，並且生兒育女。
GEN|11|16|希伯 活到三十四歲，生了 法勒 。
GEN|11|17|希伯 生 法勒 之後又活了四百三十年，並且生兒育女。
GEN|11|18|法勒 活到三十歲，生了 拉吳 。
GEN|11|19|法勒 生 拉吳 之後又活了二百零九年，並且生兒育女。
GEN|11|20|拉吳 活到三十二歲，生了 西鹿 。
GEN|11|21|拉吳 生 西鹿 之後又活了二百零七年，並且生兒育女。
GEN|11|22|西鹿 活到三十歲，生了 拿鶴 。
GEN|11|23|西鹿 生 拿鶴 之後又活了二百年，並且生兒育女。
GEN|11|24|拿鶴 活到二十九歲，生了 他拉 。
GEN|11|25|拿鶴 生 他拉 之後又活了一百一十九年，並且生兒育女。
GEN|11|26|他拉 活到七十歲，生了 亞伯蘭 、 拿鶴 和 哈蘭 。
GEN|11|27|這是 他拉 的後代。 他拉 生 亞伯蘭 、 拿鶴 和 哈蘭 ； 哈蘭 生 羅得 。
GEN|11|28|哈蘭 死在他父親 他拉 的面前，死在他的出生地 迦勒底 的 吾珥 。
GEN|11|29|亞伯蘭 、 拿鶴 各娶了妻。 亞伯蘭 的妻子名叫 撒萊 ， 拿鶴 的妻子名叫 密迦 ，是 哈蘭 的女兒。 哈蘭 是 密迦 和 亦迦 的父親。
GEN|11|30|撒萊 不生育，沒有孩子。
GEN|11|31|他拉 帶著他兒子 亞伯蘭 和他孫子， 哈蘭 的兒子 羅得 ，以及他的媳婦， 亞伯蘭 的妻子 撒萊 ，一同出了 迦勒底 的 吾珥 ，要往 迦南 地去；他們來到 哈蘭 ，就住在那裏。
GEN|11|32|他拉 共活了二百零五年，就死在 哈蘭 。
GEN|12|1|耶和華對 亞伯蘭 說：「你要離開本地、本族、父家，往我所要指示你的地去。
GEN|12|2|我必使你成為大國，我必賜福給你，使你的名為大；你要使別人得福 。
GEN|12|3|為你祝福的，我必賜福給他；詛咒你的，我必詛咒他。地上的萬族都必因你得福。」
GEN|12|4|亞伯蘭 就遵照耶和華的吩咐去了； 羅得 也和他同去。 亞伯蘭 離開 哈蘭 的時候年七十五歲。
GEN|12|5|亞伯蘭 帶著他妻子 撒萊 和姪兒 羅得 ，以及他們在 哈蘭 積蓄的財物、獲得的人口，往 迦南 地去。他們就來到了 迦南 地。
GEN|12|6|亞伯蘭 經過那地，直到 示劍 地方， 摩利 橡樹那裏；當時 迦南 人住在那地。
GEN|12|7|耶和華向 亞伯蘭 顯現，說：「我要把這地賜給你的後裔。」 亞伯蘭 就在那裏為向他顯現的耶和華築了一座壇。
GEN|12|8|從那裏他又遷到 伯特利 東邊的山，支搭帳棚；西邊是 伯特利 ，東邊是 艾 。他在那裏又為耶和華築了一座壇，求告耶和華的名。
GEN|12|9|後來 亞伯蘭 漸漸遷往 尼革夫 去。
GEN|12|10|那地遭遇饑荒。 亞伯蘭 因那地的饑荒嚴重，就下到 埃及 ，要在那裏寄居。
GEN|12|11|將近 埃及 ，他對妻子 撒萊 說：「看哪，我知道你是美貌的女人。
GEN|12|12|埃及 人看見你會說：『這是他的妻子』，他們就會殺我，卻讓你活著。
GEN|12|13|所以，請你說你是我的妹妹，使我可以因你得平安，我的性命也因你存活。」
GEN|12|14|亞伯蘭 到達 埃及 時， 埃及 人看見那女人極其美貌。
GEN|12|15|法老的臣僕看見了她，就在法老面前稱讚她。那女人就被帶進法老的宮中。
GEN|12|16|法老就因她厚待 亞伯蘭 ，給了 亞伯蘭 許多牛、羊、公驢、奴僕、婢女、母驢、駱駝。
GEN|12|17|耶和華因 亞伯蘭 妻子 撒萊 的緣故，降大災擊打法老和他的全家。
GEN|12|18|法老召了 亞伯蘭 來，說：「你向我做的是甚麼事呢？為甚麼沒有告訴我她是你的妻子？
GEN|12|19|為甚麼說『她是我的妹妹』，以致我把她接來要作我的妻子呢？現在 ，看哪，你的妻子在這裏，帶她走吧！」
GEN|12|20|於是法老吩咐人把 亞伯蘭 和他妻子，以及他一切所有的都送走了。
GEN|13|1|亞伯蘭 帶著他的妻子與 羅得 ，以及一切所有的，從 埃及 上 尼革夫 去。
GEN|13|2|亞伯蘭 的牲畜和金銀極多。
GEN|13|3|他從 尼革夫 漸漸往 伯特利 去，到了 伯特利 和 艾 的中間，當初他支搭帳棚的地方，
GEN|13|4|也是他起先築壇的地方。 亞伯蘭 在那裏求告耶和華的名。
GEN|13|5|與 亞伯蘭 同行的 羅得 也有牛群、羊群、帳棚。
GEN|13|6|那地容不下他們住在一起；因為他們的財物非常多，使他們不能同住一起。
GEN|13|7|當時， 迦南 人與 比利洗 人在那地居住。 亞伯蘭 的牧人和 羅得 的牧人之間起了爭端。
GEN|13|8|亞伯蘭 就對 羅得 說：「你我不可以相爭，你的牧人和我的牧人也不可以相爭，因為我們是一家人。
GEN|13|9|遍地不都在你眼前嗎？請你離開我吧！你向左，我就向右；你向右，我就向左。」
GEN|13|10|羅得 舉目，看見 約旦河 整個平原，直到 瑣珥 ，都是水源充足之地。在耶和華未毀滅 所多瑪 、 蛾摩拉 以前，那地好像耶和華的園子，又像 埃及 地。
GEN|13|11|於是 羅得 選擇了 約旦河 整個平原。 羅得 往東遷移，他們就彼此分開了。
GEN|13|12|亞伯蘭 住在 迦南 地； 羅得 住在平原的城鎮，他漸漸遷移帳棚，直到 所多瑪 。
GEN|13|13|所多瑪 人在耶和華面前罪大惡極。
GEN|13|14|羅得 離開 亞伯蘭 以後，耶和華對 亞伯蘭 說：「你要從你所在的地方，舉目向東西南北觀看；
GEN|13|15|你所看見一切的地，我都要把它賜給你和你的後裔，直到永遠。
GEN|13|16|我要使你的後裔好像地上的塵沙，人若能數地上的塵沙，才能數你的後裔。
GEN|13|17|你起來，縱橫走遍這地，因為我必把這地賜給你。」
GEN|13|18|亞伯蘭 就遷移帳棚，來到 希伯崙 ， 幔利 的橡樹那裏居住，在那裏為耶和華築了一座壇。
GEN|14|1|當 暗拉非 作 示拿 王， 亞略 作 以拉撒 王， 基大老瑪 作 以攔 王， 提達 作 戈印 王的時候，
GEN|14|2|他們攻打 所多瑪 王 比拉 、 蛾摩拉 王 比沙 、 押瑪 王 示納 、 洗扁 王 善以別 和 比拉 王， 比拉 就是 瑣珥 。
GEN|14|3|這些王都會合在 西訂谷 ， 西訂谷 就是 鹽海 。
GEN|14|4|他們已經服事 基大老瑪 十二年，第十三年就背叛了。
GEN|14|5|第十四年， 基大老瑪 和與他結盟的王都來了，在 亞特律‧加寧 擊敗 利乏音 人，在 哈麥 擊敗 蘇西 人，在 沙微‧基列亭 擊敗 以米 人，
GEN|14|6|在 何利 人的 西珥山 擊敗 何利 人，一直到靠近曠野的 伊勒‧巴蘭 。
GEN|14|7|他們轉回，來到 安‧密巴 ，就是 加低斯 ，擊敗了 亞瑪力 全地的人，以及住在 哈洗遜‧他瑪 的 亞摩利 人。
GEN|14|8|於是 所多瑪 王、 蛾摩拉 王、 押瑪 王、 洗扁 王和 比拉 王， 比拉 就是 瑣珥 ，都出來，在 西訂谷 擺陣，與他們交戰，
GEN|14|9|就是與 以攔 王 基大老瑪 、 戈印 王 提達 、 示拿 王 暗拉非 、 以拉撒 王 亞略 交戰；這就是四王對五王之戰。
GEN|14|10|西訂谷 有許多柏油坑。 所多瑪 王和 蛾摩拉 王逃跑，掉在坑裏，其餘的人都往山上逃跑。
GEN|14|11|四王就把 所多瑪 和 蛾摩拉 所有的財物和所有的糧食都擄掠去了；
GEN|14|12|他們也把 亞伯蘭 的姪兒 羅得 和 羅得 的財物都擄掠去了。當時 羅得 住在 所多瑪 。
GEN|14|13|有一個逃脫的人來告訴 希伯來 人 亞伯蘭 ； 亞伯蘭 正住在 亞摩利 人 幔利 的橡樹那裏。 幔利 、 以實各 和 亞乃 都是弟兄，曾與 亞伯蘭 結盟。
GEN|14|14|亞伯蘭 聽見他姪兒 被擄去，就把三百一十八個生在他家中、受過訓練的壯丁全都出動 去追，一直到 但 。
GEN|14|15|在夜間，他和他的僕人分隊擊敗了敵人，並且追殺他們，直到 大馬士革 北邊的 何把 。
GEN|14|16|他把一切被擄掠的財物奪回，也把他姪兒 羅得 和他的財物，以及人和婦女都奪回來。
GEN|14|17|亞伯蘭 擊敗 基大老瑪 和與他結盟的王回來的時候， 所多瑪 王出來，在 沙微谷 迎接他， 沙微谷 就是 王的谷 。
GEN|14|18|又有 撒冷 王 麥基洗德 帶著餅和酒出來；他是至高上帝的祭司。
GEN|14|19|他為 亞伯蘭 祝福，說： 「願至高的上帝、 天地的主賜福給 亞伯蘭 ！
GEN|14|20|至高的上帝把敵人交在你手裏， 他是應當稱頌的！」 亞伯蘭 就把所有的拿出十分之一給他。
GEN|14|21|所多瑪 王對 亞伯蘭 說：「你把人還給我，財物你自己拿去吧！」
GEN|14|22|亞伯蘭 對 所多瑪 王說：「我指著耶和華—至高的上帝、天地的主起誓：
GEN|14|23|凡是你的東西，就是一根線、一條鞋帶，我都不拿，免得你說：『是我使 亞伯蘭 富足！』
GEN|14|24|我甚麼都不要，只是僕人所吃的，以及與我同去的 亞乃 、 以實各 、 幔利 所應得的份，讓他們拿去吧！」
GEN|15|1|這些事以後，耶和華的話在異象中臨到 亞伯蘭 ，說：「 亞伯蘭 哪，不要懼怕！我是你的盾牌，你必得豐富的賞賜。」
GEN|15|2|亞伯蘭 說：「主耶和華啊，我還沒有兒子，你能賜我甚麼呢？承受我家業的是 大馬士革 人 以利以謝 。」
GEN|15|3|亞伯蘭 又說：「看哪，你沒有給我後嗣。你看，那生在我家中的人要繼承我。」
GEN|15|4|看哪，耶和華的話又臨到他，說：「這人不會繼承你，你本身所生的才會繼承你。」
GEN|15|5|於是耶和華帶他到外面，說：「你向天觀看，去數星星，你能數得清嗎？」又對他說：「你的後裔將要如此。」
GEN|15|6|亞伯蘭 信耶和華，耶和華就以此算他為義。
GEN|15|7|耶和華又對他說：「我是耶和華，曾領你出 迦勒底 的 吾珥 ，為要把這地賜你為業。」
GEN|15|8|亞伯蘭 說：「主耶和華啊，我怎能知道我必得這地為業呢？」
GEN|15|9|耶和華對他說：「你為我取一頭三歲的母牛犢，一隻三歲的母山羊，一隻三歲的公綿羊，一隻斑鳩和一隻雛鴿。」
GEN|15|10|亞伯蘭 就把這些都取來，每樣從中間劈成兩半，一半對著另一半排列，只有鳥沒有劈開。
GEN|15|11|當鷙鳥下來，落在這些屍體上時， 亞伯蘭 就把牠們趕走了。
GEN|15|12|日落的時候， 亞伯蘭 沉睡了。看哪，有大而可怕的黑暗落在他身上。
GEN|15|13|耶和華對 亞伯蘭 說：「你要確實知道，你的後裔必寄居在別人的地，服事那地的人；那地的人要虐待他們四百年。
GEN|15|14|但我要懲罰他們所服事的那國，以後他們必帶著許多財物從那裏出來。
GEN|15|15|至於你，你要平平安安歸到你祖先那裏，必享長壽，被人埋葬。
GEN|15|16|到了第四代，他們必回到這裏，因為 亞摩利 人的罪惡到現在還沒有滿盈。」
GEN|15|17|日落天黑的時候，看哪，有冒煙的爐和燒著的火把從那些肉塊中經過。
GEN|15|18|在那日，耶和華與 亞伯蘭 立約，說：「我已賜給你的後裔這一片地，從 埃及河 直到 大河 ， 幼發拉底河 ，
GEN|15|19|就是 基尼 人、 基尼洗 人、 甲摩尼 人、
GEN|15|20|赫 人、 比利洗 人、 利乏音 人、
GEN|15|21|亞摩利 人、 迦南 人、 革迦撒 人、 耶布斯 人的地。」
GEN|16|1|亞伯蘭 的妻子 撒萊 沒有為他生孩子。 撒萊 有一個婢女，是 埃及 人，名叫 夏甲 。
GEN|16|2|撒萊 對 亞伯蘭 說：「看哪，耶和華使我不能生育。你來和我的婢女同房，也許我可以從她得孩子 。」 亞伯蘭 聽從了 撒萊 的話。
GEN|16|3|於是 亞伯蘭 的妻子 撒萊 把她的婢女， 埃及 人 夏甲 ，給了丈夫為妾；那時 亞伯蘭 在 迦南 已經住了十年。
GEN|16|4|亞伯蘭 與 夏甲 同房， 夏甲 就懷了孕。她看見自己有孕，就輕視她的女主人。
GEN|16|5|撒萊 對 亞伯蘭 說：「我因你受了委屈。我把我的婢女放在你懷中，她見自己懷了孕，就輕視我。願耶和華在你我之間判斷。」
GEN|16|6|亞伯蘭 對 撒萊 說：「看哪，婢女在你手裏，你可以照你看為好的對待她。」於是， 撒萊 虐待她，她就從 撒萊 面前逃走了。
GEN|16|7|耶和華的使者在曠野的水泉旁，在 書珥 路上的水泉旁遇見 夏甲 ，
GEN|16|8|對她說：「 撒萊 的婢女 夏甲 ，你從哪裏來？要到哪裏去？」她說：「我從我的女主人 撒萊 面前逃出來。」
GEN|16|9|耶和華的使者對她說：「你要回到你的女主人那裏，屈服在她手下。」
GEN|16|10|耶和華的使者對她說： 「我必使你的後裔極其繁多， 多到不可勝數。」
GEN|16|11|耶和華的使者又對她說： 「看哪，你已懷孕， 要生一個兒子。 你要給他起名叫 以實瑪利 ， 因為耶和華聽見了你的苦楚。
GEN|16|12|他為人必像野驢。 他的手要攻打人， 人的手也要攻打他； 他必常與他的眾弟兄作對 。」
GEN|16|13|夏甲 就稱那向她說話的耶和華為「你是看見 的上帝」，因為她說：「他看見了我之後，我還能在這裏看見他嗎？」
GEN|16|14|所以這井名叫 庇耳‧拉海‧萊 ，看哪，它位於 加低斯 和 巴列 的中間。
GEN|16|15|後來 夏甲 為 亞伯蘭 生了一個兒子； 亞伯蘭 給 夏甲 生的兒子起名叫 以實瑪利 。
GEN|16|16|夏甲 為 亞伯蘭 生 以實瑪利 的時候， 亞伯蘭 年八十六歲。
GEN|17|1|亞伯蘭 九十九歲時，耶和華向他顯現，對他說：「我是全能的上帝。你當在我面前行走，作完全的人，
GEN|17|2|我要與你立約，使你的後裔極其繁多。」
GEN|17|3|亞伯蘭 臉伏於地；上帝又對他說：
GEN|17|4|「看哪，這就是我與你立的約，你要成為多國的父。
GEN|17|5|從今以後，你的名字不再叫 亞伯蘭 ，要叫 亞伯拉罕 ，因為我已經立你作多國之父。
GEN|17|6|我必使你生養極其繁多；國度要從你而立，君王要從你而出。
GEN|17|7|我要與你，以及你世世代代的後裔堅立我的約，成為永遠的約，是要作你和你後裔的上帝。
GEN|17|8|我要把你現在寄居的地，就是 迦南 全地，賜給你和你的後裔永遠為業；我也必作他們的上帝。」
GEN|17|9|上帝又對 亞伯拉罕 說：「你和你的後裔一定要世世代代遵守我的約。
GEN|17|10|這就是我與你，以及你的後裔所立的約，是你們所當遵守的，你們所有的男子都要受割禮。
GEN|17|11|你們要割去肉體的包皮，這是我與你們立約的記號。
GEN|17|12|你們世世代代的男子，無論是在家裏生的，或是用銀子從外人買來而不是你後裔生的，都要在生下來的第八日受割禮。
GEN|17|13|你家裏生的和你用銀子買的，都必須受割禮。這樣，我的約就在你們肉體上成為永遠的約。
GEN|17|14|不受割禮的男子都必從民中剪除，因他違背了我的約。」
GEN|17|15|上帝又對 亞伯拉罕 說：「至於你的妻子 撒萊 ，不可再叫她 撒萊 ，她的名要叫 撒拉 。
GEN|17|16|我必賜福給她，也要從她賜一個兒子給你。我必賜福給 撒拉 ，她要興起多國；必有百姓的君王從她而出。」
GEN|17|17|亞伯拉罕 就臉伏於地竊笑，心裏想：「一百歲的人還能有孩子嗎？ 撒拉 已經九十歲了，還能生育嗎？」
GEN|17|18|亞伯拉罕 對上帝說：「但願 以實瑪利 活在你面前。」
GEN|17|19|上帝說：「不！你妻子 撒拉 必為你生一個兒子，你要給他起名叫 以撒 。我要與他堅立我的約，成為他後裔永遠的約。
GEN|17|20|至於 以實瑪利 ，我已聽見你了：看哪，我必賜福給他，使他興旺，極其繁多。他必生十二個族長，我要使他成為大國。
GEN|17|21|到明年所定的時候， 撒拉 必為你生 以撒 ，我要與他堅立我的約。」
GEN|17|22|上帝和 亞伯拉罕 說完了話，就離開他上升去了。
GEN|17|23|在那一天， 亞伯拉罕 遵照上帝所說的，給他的兒子 以實瑪利 和家裏所有的男丁，無論是在家裏生的，或是用銀子買來的，都行了割禮 。
GEN|17|24|亞伯拉罕 受割禮時，年九十九歲。
GEN|17|25|他兒子 以實瑪利 受割禮時，年十三歲。
GEN|17|26|在那一天， 亞伯拉罕 和他兒子 以實瑪利 一同受了割禮。
GEN|17|27|家裏所有的男人，無論是在家裏生的，或是用銀子從外人買來的，也都一同受了割禮。
GEN|18|1|耶和華在 幔利 橡樹那裏向 亞伯拉罕 顯現。天正熱的時候， 亞伯拉罕 坐在帳棚門口。
GEN|18|2|他舉目觀看，看哪，有三個人站在他附近。他一看見，就從帳棚門口跑去迎接他們，俯伏在地，
GEN|18|3|說：「我主，我若在你眼前蒙恩，請不要離開你的僕人走過去。
GEN|18|4|容我拿點水來，請你們洗腳，在樹下休息。
GEN|18|5|既然你們來到僕人這裏了，我再拿點餅來，讓你們恢復心力，然後再走。」他們說：「就照你說的去做吧。」
GEN|18|6|亞伯拉罕 急忙進帳棚到 撒拉 那裏，說：「你趕快拿三細亞細麵，揉麵做餅。」
GEN|18|7|亞伯拉罕 又跑到牛群裏，牽了一頭又嫩又好的牛犢來，交給僕人，僕人就急忙去預備。
GEN|18|8|亞伯拉罕 取了乳酪和奶，以及預備好了的牛犢來，擺在他們面前，自己在樹下站在旁邊，他們就吃了。
GEN|18|9|他們對 亞伯拉罕 說：「你妻子 撒拉 在哪裏？」他說：「看哪，在帳棚裏。」
GEN|18|10|有一位說：「明年這時候 ，我一定會回到你這裏。看哪，你的妻子 撒拉 會生一個兒子。」 撒拉 在那人後面的帳棚門口也聽見了。
GEN|18|11|亞伯拉罕 和 撒拉 都年紀老邁， 撒拉 的月經已停了。
GEN|18|12|撒拉 心裏竊笑，說：「我已衰老，我的主也老了，怎能有這喜事呢？」
GEN|18|13|耶和華對 亞伯拉罕 說：「 撒拉 為甚麼竊笑，說：『我已年老，果真能生育嗎？』
GEN|18|14|耶和華豈有難成的事嗎？到了所定的時候，我必回到你這裏。明年這時候， 撒拉 會生一個兒子。」
GEN|18|15|撒拉 因為害怕，就不承認，說：「我沒有笑。」那人說：「不，你的確笑了。」
GEN|18|16|三人從那裏起程，面向 所多瑪 觀望， 亞伯拉罕 與他們同行，要送他們一程。
GEN|18|17|耶和華說：「我所要做的事豈可瞞著 亞伯拉罕 呢？
GEN|18|18|亞伯拉罕 必要成為強大的國；地上的萬國都必因他得福。
GEN|18|19|我揀選他 ，為要叫他命令他的子孫和後代家屬遵行耶和華的道，秉公行義，使耶和華所應許 亞伯拉罕 的話都實現了。」
GEN|18|20|耶和華說：「 所多瑪 和 蛾摩拉 罪惡極其嚴重，控告他們的聲音很大。
GEN|18|21|我要下去察看他們所做的，是否真的像那達到我這裏的聲音一樣；如果不是，我也要知道。」
GEN|18|22|二人轉身離開那裏，往 所多瑪 去；但 亞伯拉罕 仍然站在耶和華面前。
GEN|18|23|亞伯拉罕 近前來，說：「你真的要把義人和惡人一同剿滅嗎？
GEN|18|24|假若那城裏有五十個義人，你真的還要剿滅，不因城裏這五十個義人饒了那地方嗎？
GEN|18|25|你絕不會做這樣的事，把義人與惡人一同殺了，使義人與惡人一樣。你絕不會這樣！審判全地的主豈不做公平的事嗎？」
GEN|18|26|耶和華說：「我若在 所多瑪城 裏找到五十個義人，我就為他們的緣故饒恕那整個地方。」
GEN|18|27|亞伯拉罕 回答說：「看哪，我雖只是塵土灰燼，還敢向主說話。
GEN|18|28|假若這五十個義人少了五個，你就因為少了五個而毀滅全城嗎？」他說：「我在那裏若找到四十五個，就不毀滅。」
GEN|18|29|亞伯拉罕 又對他說：「假若在那裏找到四十個呢？」他說：「為這四十個的緣故，我也不做。」
GEN|18|30|亞伯拉罕 說：「求主不要生氣，容我說，假若在那裏找到三十個呢？」他說：「我在那裏若找到三十個，我也不做。」
GEN|18|31|亞伯拉罕 說：「看哪，我還敢向主說，假若在那裏找到二十個呢？」他說：「為這二十個的緣故，我也不毀滅。」
GEN|18|32|亞伯拉罕 說：「求主不要生氣，我再說一次，假若在那裏找到十個呢？」他說：「為這十個的緣故，我也不毀滅。」
GEN|18|33|耶和華與 亞伯拉罕 說完了話就走了； 亞伯拉罕 也回到自己的地方去了。
GEN|19|1|兩個天使在傍晚到了 所多瑪 ， 羅得 正坐在 所多瑪 的城門口。 羅得 一看見，就起身迎接他們，臉伏於地下拜，
GEN|19|2|說：「看哪，我主，請你們轉到僕人家裏過夜，洗你們的腳，清早起來再上路。」他們說：「不！我們要在廣場上過夜。」
GEN|19|3|羅得 懇切地請他們，他們就轉向他，進到他屋裏。 羅得 為他們預備宴席，烤無酵餅，他們就吃了。
GEN|19|4|他們還沒有躺下， 所多瑪城 的人，連老帶少所有的人，個個都來圍住那屋子。
GEN|19|5|他們呼叫 羅得 ，對他說：「今天晚上到你這裏來的人在哪裏？把他們帶出來，讓我們親近他們。」
GEN|19|6|羅得 出了門，把身後的門關上，到眾人那裏，
GEN|19|7|說：「我的弟兄們，請你們不要做這惡事。
GEN|19|8|看哪，我有兩個女兒，還沒有親近過男人，讓我領她們出來給你們，就照你們看為好的對待她們吧！只是這兩個人既然到我舍下，請不要向他們做這事。」
GEN|19|9|眾人說：「站到一邊去吧！」又說：「這個人來寄居，還想扮審判官呢！現在我們要害你比害他們更厲害。」眾人就往前衝向 羅得 ，要攻破大門。
GEN|19|10|那兩個人伸出手來，把 羅得 拉進屋子他們那裏，就關上門。
GEN|19|11|他們擊打門外的人，無論老少，都眼睛迷糊，找門找得很煩躁。
GEN|19|12|那兩個人對 羅得 說：「你這裏還有甚麼人嗎？無論是女婿，是兒女，這城中所有屬你的人，你都要把他們從這地方帶出去。
GEN|19|13|我們要毀滅這地方，因為控告城內百姓的聲音在耶和華面前非常大，耶和華派我們來毀滅這城。」
GEN|19|14|羅得 出去，告訴娶了 他女兒的女婿們說：「起來，離開這地方，因為耶和華要毀滅這城。」他的女婿們卻以為他說的是笑話。
GEN|19|15|天亮了，天使催逼 羅得 說：「起來！帶著你的妻子和你這裏的兩個女兒出去，免得你因這城的罪孽同被剿滅。」
GEN|19|16|但 羅得 遲延不走。二人因為耶和華憐憫 羅得 ，就拉著他的手和他妻子的手，以及他兩個女兒的手，把他們領出來，安置在城外；
GEN|19|17|領他們出來以後，就說：「逃命吧！不可回頭看，也不可在平原站住。要往山上逃跑，免得你被剿滅。」
GEN|19|18|羅得 對他們說：「我主啊，不要這樣！
GEN|19|19|看哪，你僕人已經在你眼前蒙恩，你又向我大施慈愛，救我的性命。但是我不能逃到山上去，恐怕這災禍追上我，我就死了。
GEN|19|20|看哪，這城又近又小，比較容易逃到那裏。這不是一座小城嗎？求你容我逃到那裏，使我的性命可以存活。」
GEN|19|21|天使對他說：「看哪，這事我也應允你，不傾覆你所說的這城。
GEN|19|22|你要趕快逃到那城，因為你還沒有到那裏，我不能做甚麼。」因此那城名叫 瑣珥 。
GEN|19|23|羅得 到了 瑣珥 ，太陽已經升出地面。
GEN|19|24|當時，耶和華把硫磺與火，從天上耶和華那裏降與 所多瑪 和 蛾摩拉 ，
GEN|19|25|把那些城和全平原，城裏所有的居民和土地上生長的，都毀滅了。
GEN|19|26|羅得 的妻子在他後邊回頭一看，就變成了一根鹽柱。
GEN|19|27|亞伯拉罕 清早起來，到了他先前站在耶和華面前的地方，
GEN|19|28|面向 所多瑪 和 蛾摩拉 ，以及平原全地觀望。他觀看，看哪，那地有濃煙上騰，好像燒窯的濃煙。
GEN|19|29|當上帝毀滅平原諸城的時候，他記念 亞伯拉罕 ；在傾覆 羅得 所住之城的時候，就把 羅得 從傾覆中帶出來。
GEN|19|30|羅得 因為怕住在 瑣珥 ，就同他兩個女兒從 瑣珥 上去，住在山上。他和兩個女兒住在一個洞裏。
GEN|19|31|大女兒對小女兒說：「我們的父親老了，這地又沒有男人可以照世上的禮俗來與我們結合。
GEN|19|32|來！我們叫父親喝酒，然後與他同寢。這樣，我們可以從我們的父親存留後裔。」
GEN|19|33|於是，那晚她們叫父親喝酒，大女兒就進去和她父親同寢；她幾時躺下，幾時起來，父親都不知道。
GEN|19|34|第二天，大女兒對小女兒說：「看哪，我昨夜與父親同寢。今晚我們再叫他喝酒，你進去與他同寢。這樣，我們可以從父親存留後裔。」
GEN|19|35|於是，那晚她們又叫父親喝酒，小女兒起來與她父親同寢；她幾時躺下，幾時起來，父親都不知道。
GEN|19|36|這樣， 羅得 的兩個女兒都從她們的父親懷了孕。
GEN|19|37|大女兒生了兒子，給他起名叫 摩押 ，就是現今 摩押 人的始祖。
GEN|19|38|小女兒也生了兒子，給他起名叫 便‧亞米 ，就是現今 亞捫 人的始祖。
GEN|20|1|亞伯拉罕 從那裏往 尼革夫 遷移，寄居在 加低斯 和 書珥 之間的 基拉耳 。
GEN|20|2|亞伯拉罕 稱他的妻子 撒拉 為妹妹。 基拉耳 王 亞比米勒 派人把 撒拉 帶走。
GEN|20|3|夜間，上帝在夢中來到 亞比米勒 那裏，對他說：「看哪，你要死了，因為你帶來的女人，她是有丈夫的女子！」
GEN|20|4|亞比米勒 還未親近 撒拉 ；他說：「主啊，連公義的國，你也要毀滅嗎？
GEN|20|5|那人豈不是自己對我說『她是我妹妹』嗎？連這女人自己也說：『他是我哥哥。』我做這事是心正手潔的。」
GEN|20|6|上帝在夢中對他說：「我也知道你做這事是心中正直的；是我攔阻了你，免得你得罪我。所以我不讓你侵犯她。
GEN|20|7|現在你當把這人的妻子歸還給他；因為他是先知，他要為你禱告，使你存活。你若不歸還，你當知道，你和你所有的人都必定死。」
GEN|20|8|亞比米勒 清早起來，叫了他的眾臣僕來，把這一切事說給他們聽，他們就很害怕。
GEN|20|9|亞比米勒 召了 亞伯拉罕 來，對他說：「你怎麼向我這樣做呢？我甚麼事得罪你，你竟使我和我的國陷在大罪中呢？你對我做了不該做的事了！」
GEN|20|10|亞比米勒 對 亞伯拉罕 說：「你看見甚麼才做這事呢？」
GEN|20|11|亞伯拉罕 說：「我以為這地方的人根本不敬畏上帝，必為我妻子的緣故殺我。
GEN|20|12|況且她也真是我的妹妹；她與我是同父異母的，後來作了我的妻子。
GEN|20|13|當上帝叫我離開父家、飄流在外的時候，我對她說：我們無論走到甚麼地方，你要對人說：『他是我哥哥』，這就是你以慈愛待我了。」
GEN|20|14|亞比米勒 把牛、羊、奴僕、婢女送給 亞伯拉罕 ，也把他的妻子 撒拉 歸還給他。
GEN|20|15|亞比米勒 說：「看哪，我的地都在你面前，你看為好的地方就居住吧。」
GEN|20|16|他對 撒拉 說：「看哪，我給你哥哥一千銀子。看哪，這要在你全家人面前遮羞 ，向眾人證實你是清白的。」
GEN|20|17|亞伯拉罕 向上帝禱告，上帝就醫好 亞比米勒 和他的妻子，以及他的使女們，他們就能生育。
GEN|20|18|因耶和華為 亞伯拉罕 的妻子 撒拉 的緣故，已經使 亞比米勒 家中的婦人不能懷孕。
GEN|21|1|耶和華照著他所說的眷顧 撒拉 ，耶和華實現了他對 撒拉 的應許。
GEN|21|2|亞伯拉罕 年老，到上帝對他說的那所定的時候， 撒拉 懷了孕，給他生了一個兒子。
GEN|21|3|亞伯拉罕 給 撒拉 所生的兒子起名叫 以撒 。
GEN|21|4|以撒 出生後第八日， 亞伯拉罕 遵照上帝所吩咐的，為 以撒 行割禮。
GEN|21|5|他兒子 以撒 出生的時候， 亞伯拉罕 年一百歲。
GEN|21|6|撒拉 說：「上帝使我歡笑，凡聽見的人必與我一同歡笑」，
GEN|21|7|又說：「誰能預先對 亞伯拉罕 說， 撒拉 要乳養孩子呢？因為在他年老的時候，我為他生了一個兒子。」
GEN|21|8|孩子漸漸長大，就斷了奶。 以撒 斷奶的那一天， 亞伯拉罕 擺設豐盛的宴席。
GEN|21|9|那時， 撒拉 看見 埃及 人 夏甲 為 亞伯拉罕 所生的兒子戲笑，
GEN|21|10|就對 亞伯拉罕 說：「你把這使女和她兒子趕出去！因為這使女的兒子不可與我的兒子 以撒 一同承受產業。」
GEN|21|11|亞伯拉罕 為這事非常憂愁，因為關乎他的兒子。
GEN|21|12|上帝對 亞伯拉罕 說：「你不必為這孩子和你的使女憂愁。 撒拉 對你說的話，你都要聽從；因為從 以撒 生的，才要稱為你的後裔。
GEN|21|13|至於使女的兒子，我也必使他成為一國，因為他是你的後裔。」
GEN|21|14|亞伯拉罕 清早起來，拿餅和一皮袋水，給了 夏甲 ，搭在她肩上，把她和孩子一起送走。 夏甲 就走了，但她卻在 別是巴 的曠野流浪。
GEN|21|15|皮袋的水用完了， 夏甲 就把孩子放在一棵小樹下，
GEN|21|16|自己走開約有一箭之遠，相對而坐，說：「我不忍心看見孩子死」。她就坐在對面，放聲大哭。
GEN|21|17|上帝聽見孩子的聲音，上帝的使者就從天上呼叫 夏甲 說：「 夏甲 ，你為何這樣呢？不要害怕，上帝已經聽見孩子在那裏的聲音了。
GEN|21|18|起來！把孩子扶起來，用你的手握住他，因我必使他成為大國。」
GEN|21|19|上帝開了 夏甲 的眼睛，她就看見一口水井。她就去，把皮袋裝滿了水，給孩子喝。
GEN|21|20|上帝與這孩子同在，他就漸漸長大，住在曠野，成了一個弓箭手。
GEN|21|21|他住在 巴蘭 的曠野；他母親從 埃及 地為他娶了一個妻子。
GEN|21|22|那時候， 亞比米勒 和他的將軍 非各 對 亞伯拉罕 說：「凡你所做的事，上帝都與你同在。
GEN|21|23|我願你如今在這裏指著上帝對我起誓，不要虧待我和我的兒子，以及我的子孫。我怎樣忠誠待你，你也要照樣忠誠待我和你所寄居的這地。」
GEN|21|24|亞伯拉罕 說：「我願意起誓。」
GEN|21|25|先前， 亞比米勒 的僕人霸佔了一口水井， 亞伯拉罕 為這事責備 亞比米勒 。
GEN|21|26|亞比米勒 說：「我不知道誰做了這事，你也沒有告訴我，我到今日才聽到。」
GEN|21|27|亞伯拉罕 把羊和牛給了 亞比米勒 ，二人就彼此立約。
GEN|21|28|亞伯拉罕 把七隻小母羊另放在一處。
GEN|21|29|亞比米勒 對 亞伯拉罕 說：「你把這七隻小母羊另放一處是甚麼意思呢？」
GEN|21|30|他說：「你要從我手裏接受這七隻小母羊，作我挖了這口井的證據。」
GEN|21|31|所以他給那地方起名叫 別是巴 ，因為他們二人在那裏起了誓。
GEN|21|32|他們在 別是巴 立了約， 亞比米勒 就和他的將軍 非各 起身回 非利士 人的地去了。
GEN|21|33|亞伯拉罕 就在 別是巴 種了一棵柳樹，在那裏求告耶和華—永恆上帝的名。
GEN|21|34|亞伯拉罕 在 非利士 人的地寄居了許多日子。
GEN|22|1|這些事以後，上帝考驗 亞伯拉罕 ，對他說：「 亞伯拉罕 ！」他說：「我在這裏。」
GEN|22|2|上帝說：「你要帶你的兒子，就是你所愛的獨子 以撒 ，往 摩利亞 地去，在我指示你的一座山上，把他獻為燔祭。」
GEN|22|3|亞伯拉罕 清早起來，預備了驢，帶著跟他一起的兩個僕人和他兒子 以撒 ，劈好了燔祭的柴，就起身往上帝指示他的地方去了。
GEN|22|4|到了第三日， 亞伯拉罕 舉目遙望那地方。
GEN|22|5|亞伯拉罕 對他的僕人說：「你們和驢留在這裏，我和孩子要去那裏敬拜，然後回到你們這裏來。」
GEN|22|6|亞伯拉罕 把燔祭的柴放在他兒子 以撒 身上，自己手裏拿著火與刀；於是二人同行。
GEN|22|7|以撒 對他父親 亞伯拉罕 說：「我父啊！」 亞伯拉罕 說：「我兒，我在這裏。」 以撒 說：「看哪，火與柴都有了，但燔祭的羔羊在哪裏呢？」
GEN|22|8|亞伯拉罕 說：「我兒，上帝必自己預備燔祭的羔羊。」於是二人同行。
GEN|22|9|他們到了上帝指示他的地方， 亞伯拉罕 在那裏築壇，把柴擺好，綁了他兒子 以撒 ，放在壇的柴上。
GEN|22|10|亞伯拉罕 就伸手拿刀，要殺他的兒子。
GEN|22|11|耶和華的使者從天上呼喚他說：「 亞伯拉罕 ！ 亞伯拉罕 ！」他說：「我在這裏。」
GEN|22|12|天使說：「不可在這孩子身上下手！一點也不可傷害他！現在我知道你是敬畏上帝的人了，因為你沒有把你的兒子，就是你的獨子，留下不給我。」
GEN|22|13|亞伯拉罕 舉目觀看，看哪，一隻公綿羊兩角纏在灌木叢中。 亞伯拉罕 就去牽了那隻公綿羊，獻為燔祭，代替他的兒子。
GEN|22|14|亞伯拉罕 給那地方起名叫「耶和華以勒」 。直到今日人還說：「在耶和華的山上必有預備。」
GEN|22|15|耶和華的使者第二次從天上呼喚 亞伯拉罕 ，
GEN|22|16|說：「耶和華說：『你既行了這事，沒有留下你的兒子，就是你的獨子，我指著自己起誓：
GEN|22|17|我必多多賜福給你，我必使你的後裔大大增多，如同天上的星、海邊的沙。你的後裔必得仇敵的城門，
GEN|22|18|並且地上的萬國都必因你的後裔得福，因為你聽從了我的話。』」
GEN|22|19|於是 亞伯拉罕 回到他僕人那裏。他們一同起身，往 別是巴 去， 亞伯拉罕 就住在 別是巴 。
GEN|22|20|這些事以後，有人告訴 亞伯拉罕 說：「看哪， 密迦 也為你兄弟 拿鶴 生了幾個兒子：
GEN|22|21|長子 烏斯 、他的兄弟 布斯 、 亞蘭 的父親 基摩利 、
GEN|22|22|基薛 、 哈瑣 、 必達 、 益拉 和 彼土利 。」
GEN|22|23|彼土利 生 利百加 。這八個人都是 密迦 為 亞伯拉罕 的兄弟 拿鶴 生的。
GEN|22|24|拿鶴 的妾名叫 流瑪 ，她也生了 提八 、 迦含 、 他轄 和 瑪迦 。
GEN|23|1|撒拉 享壽一百二十七歲，這是 撒拉 一生的歲數 。
GEN|23|2|撒拉 死在 迦南 地的 基列‧亞巴 ，就是 希伯崙 。 亞伯拉罕 來哀悼 撒拉 ，為她哭泣。
GEN|23|3|然後， 亞伯拉罕 起來，離開死人面前，對 赫 人說：
GEN|23|4|「我在你們中間是外人，是寄居的。請給我你們那裏的一塊墳地，我好埋葬我的亡妻，使她不在我的面前。」
GEN|23|5|赫 人回答 亞伯拉罕 說：
GEN|23|6|「我主請聽。你在我們中間是一位尊貴的王子，只管在我們最好的墳地裏埋葬你的死人；我們沒有一人會拒絕你在他的墳地裏埋葬你的死人。」
GEN|23|7|於是， 亞伯拉罕 起來，向當地的百姓 赫 人下拜，
GEN|23|8|對他們說：「你們若願意讓我埋葬我的亡妻，使她不在我面前，就請聽我，為我求 瑣轄 的兒子 以弗崙 ，
GEN|23|9|把他田地盡頭的 麥比拉洞 賣給我。他可以按照足價賣給我，作為我在你們中間的墳地。」
GEN|23|10|那時， 以弗崙 正坐在 赫 人中間。 赫 人 以弗崙 就回答 亞伯拉罕 ，說給所有出入城門的 赫 人聽：
GEN|23|11|「不，我主請聽。我要把這塊田送給你，連田間的洞也送給你，在我同族的人眼前都給你，讓你埋葬你的死人。」
GEN|23|12|亞伯拉罕 就在當地的百姓面前下拜，
GEN|23|13|對 以弗崙 說，也給當地百姓聽：「你若應允，請你聽我。我要把田的價錢給你，請你收下，我就在那裏埋葬我的死人。」
GEN|23|14|以弗崙 回答 亞伯拉罕 說：
GEN|23|15|「我主請聽。四百舍客勒銀子的地，在你我中間算甚麼呢？只管埋葬你的死人吧！」
GEN|23|16|亞伯拉罕 聽從了 以弗崙 。 亞伯拉罕 就照著他說給 赫 人聽的，把買賣通用的銀子，秤了四百舍客勒銀子給 以弗崙 。
GEN|23|17|於是， 以弗崙 把那塊位於 幔利 對面的 麥比拉 田，和其中的洞，以及田間周圍的樹木都成交了，
GEN|23|18|在所有出入城門的 赫 人眼前，賣給 亞伯拉罕 作為他的產業。
GEN|23|19|後來， 亞伯拉罕 把他妻子 撒拉 安葬在 迦南 地 幔利 對面的 麥比拉 田間的洞裏， 幔利 就是 希伯崙 。
GEN|23|20|從此，那塊田和田間的洞就從 赫 人移交給 亞伯拉罕 作墳地的產業。
GEN|24|1|亞伯拉罕 年紀老邁，耶和華在一切事上都賜福給他。
GEN|24|2|亞伯拉罕 對他家中管理他一切產業最老的僕人說：「把你的手放在我大腿底下。
GEN|24|3|我要叫你指著耶和華—天和地的上帝起誓，不要為我兒子娶我所居住的 迦南 地的女子為妻。
GEN|24|4|你要往我的本地本族去，為我的兒子 以撒 娶妻。」
GEN|24|5|僕人對他說：「如果那女子不肯跟我來到這地，我必須把你的兒子帶回到你出來的地方嗎？」
GEN|24|6|亞伯拉罕 對他說：「你要謹慎，不可帶我兒子回那裏去。
GEN|24|7|耶和華—天上的上帝曾帶領我離開父家和本族的地，對我說話，向我起誓說：『我要將這地賜給你的後裔。』他要差遣使者在你面前，你就可以從那裏為我兒子娶妻。
GEN|24|8|倘若那女子不肯跟你來，我叫你起的誓就與你無關了，只是你不可帶我的兒子回到那裏去。」
GEN|24|9|僕人就把手放在他主人 亞伯拉罕 的大腿底下，為這事向他起誓。
GEN|24|10|那僕人從他主人的駱駝中取了十匹駱駝，他手中也帶著他主人各樣的貴重物品離開 ，起身往 美索不達米亞 去，到了 拿鶴 的城。
GEN|24|11|傍晚時，眾女子出來打水，他就讓駱駝跪在城外的水井旁。
GEN|24|12|他說：「耶和華—我主人 亞伯拉罕 的上帝啊，求你施恩給我的主人 亞伯拉罕 ，讓我今日就遇見吧！
GEN|24|13|看哪，我站在井旁，城內居民的女子們正出來打水。
GEN|24|14|我向哪一個少女說：『請你放下水瓶來，給我水喝』，她若說：『請喝！我也給你的駱駝喝』，願她作你所選定給你僕人 以撒 的妻。這樣，我就知道你施恩給我的主人了。」
GEN|24|15|話還沒說完，看哪， 利百加 肩頭上扛著水瓶出來。 利百加 是 彼土利 所生的； 彼土利 是 亞伯拉罕 的兄弟 拿鶴 妻子 密迦 的兒子。
GEN|24|16|那少女容貌極其美麗，是未曾與人親近的童女。她下到井旁，打滿了瓶子的水，就上來。
GEN|24|17|僕人跑上前去迎著她，說：「請你讓我喝你瓶子裏的一點水。」
GEN|24|18|少女說：「我主請喝！」就急忙拿下瓶子托在手上，給他喝水。
GEN|24|19|那少女給他喝足了，又說：「我也為你的駱駝打水，直到駱駝喝足了。」
GEN|24|20|她就急忙把瓶子裏的水倒在槽裏，又跑到井旁打水，為所有的駱駝打了水。
GEN|24|21|那人定睛看著少女，一句話也不說，要知道耶和華是否使他的道路亨通。
GEN|24|22|駱駝喝足了，那人就拿出一個比加 重的金環，一對十舍客勒重的金手鐲，
GEN|24|23|說：「請告訴我，你是誰的女兒？你父親家裏有沒有地方可以讓我們過夜？」
GEN|24|24|少女說：「我是 密迦 為 拿鶴 生的兒子 彼土利 的女兒。」
GEN|24|25|又說：「我們家裏有充足的乾草和飼料，也有住宿的地方。」
GEN|24|26|那人就低頭向耶和華敬拜，
GEN|24|27|說：「耶和華—我主人 亞伯拉罕 的上帝是應當稱頌的，因他不斷以慈愛信實待我主人。至於我，耶和華一路引領我，直到我主人的兄弟家裏。」
GEN|24|28|那少女跑去，把這些話告訴她母親家裏的人。
GEN|24|29|利百加 有一個哥哥，名叫 拉班 ， 拉班 就跑到外面井旁那人那裏。
GEN|24|30|當他看見金環和戴在他妹妹手上的金鐲，又聽見他妹妹 利百加 說的話：「那人如此對我說」，他就來到那人面前，看哪，他還站在井旁的駱駝旁邊，
GEN|24|31|就對他說：「你這蒙耶和華賜福的人，請進來吧！為甚麼站在外面？我已經收拾了房屋，也為駱駝預備了地方。」
GEN|24|32|那人就進了 拉班 的家。 拉班 卸了駱駝，用飼料餵牠們，拿水給那人和隨從他的人洗腳，
GEN|24|33|把食物擺在他面前，請他吃。他卻說：「我不吃，等我把我的事情說完了再吃。」 拉班 說：「請說。」
GEN|24|34|他說：「我是 亞伯拉罕 的僕人。
GEN|24|35|耶和華大大地賜福給我主人，使他發達，賜給他羊群、牛群、金銀、奴僕、婢女、駱駝和驢。
GEN|24|36|我主人的妻子 撒拉 年老的時候為我主人生了一個兒子；我主人把他一切所有的都給了他。
GEN|24|37|我主人叫我起誓說：『不要為我兒子娶我所居住的 迦南 地的女子為妻。
GEN|24|38|你要往我父家、我本族那裏去，為我的兒子娶妻。』
GEN|24|39|我對我主人說：『恐怕那女子不肯跟我來。』
GEN|24|40|他就說：『我所事奉的耶和華必要差遣他的使者與你同去，使你的道路亨通，你就可以在我父家、我本族那裏，為我的兒子娶妻。
GEN|24|41|只要你到了我本族那裏，我叫你起的誓就與你無關。他們若不把女子交給你，我叫你起的誓也與你無關。』
GEN|24|42|「我今日到了井旁，就說：『耶和華—我主人 亞伯拉罕 的上帝啊，願你使我所行的道路亨通。
GEN|24|43|看哪，我站在井旁，對哪一個出來打水的女子說：請你讓我喝你瓶子裏的一點水，
GEN|24|44|她若說：你只管喝，我也為你的駱駝打水；願那女子作耶和華給我主人兒子所選定的妻子。』
GEN|24|45|「我心裏的話還沒有說完，看哪， 利百加 肩頭上扛著水瓶出來，下到井旁打水。我對她說：『請你給我水喝。』
GEN|24|46|她就急忙從肩頭上拿下瓶子來，說：『請喝！我也給你的駱駝喝。』我就喝了；她也給我的駱駝喝了。
GEN|24|47|我問她說：『你是誰的女兒？』她說：『我是 彼土利 的女兒， 彼土利 是 密迦 和 拿鶴 生的兒子。』我就把環子戴在她鼻子上，把鐲子戴在她雙手上。
GEN|24|48|然後我低頭向耶和華敬拜，稱頌耶和華—我主人 亞伯拉罕 的上帝，因為他引導我走合適的道路，使我得著我主人兄弟的孫女，給我主人的兒子為妻。
GEN|24|49|現在你們若願以慈愛誠信待我主人，就告訴我；若不然，也告訴我，使我可以或向左，或向右。」
GEN|24|50|拉班 和 彼土利 回答說：「這事既然出於耶和華，我們不能向你說好說歹。
GEN|24|51|看哪， 利百加 就在你面前，可以將她帶去，遵照耶和華所說的，給你主人的兒子為妻。」
GEN|24|52|亞伯拉罕 的僕人聽見他們這些話，就向耶和華俯伏在地。
GEN|24|53|僕人拿出金器、銀器和衣服送給 利百加 ，又將貴重的物品送給她哥哥和她母親。
GEN|24|54|然後，僕人和隨從的人才吃喝，並且住了一夜。早晨起來，僕人說：「請讓我回我主人那裏去吧。」
GEN|24|55|利百加 的哥哥和母親說：「讓她同我們再住幾天，也許十天，然後她可以去。」
GEN|24|56|僕人對他們說：「耶和華既然使我道路亨通，你們就不要耽誤我，請讓我走，回我主人那裏去吧！」
GEN|24|57|他們說：「我們把她叫來問問她 。」
GEN|24|58|他們就叫了 利百加 來，對她說：「你和這人同去嗎？」她說：「我去。」
GEN|24|59|於是他們送他們的妹妹 利百加 和她的奶媽，同 亞伯拉罕 的僕人，以及隨從他的人走了。
GEN|24|60|他們就為 利百加 祝福，對她說： 「我們的妹妹啊， 願你作千萬人的母親！ 願你的後裔得著仇敵的城門！」
GEN|24|61|利百加 和她的女僕們起來，騎上駱駝，跟著那人去。僕人就帶著 利百加 走了。
GEN|24|62|那時， 以撒 住在 尼革夫 。他剛從 庇耳‧拉海‧萊 回來。
GEN|24|63|傍晚時， 以撒 出來，到田間默想。他舉目一看，看哪，來了一隊駱駝。
GEN|24|64|利百加 舉目看見 以撒 ，就急忙下了駱駝，
GEN|24|65|對那僕人說：「這從田間走來迎接我們的人是誰？」僕人說：「他是我的主人。」 利百加 就拿面紗蓋住自己。
GEN|24|66|僕人把他所做的一切事都告訴 以撒 。
GEN|24|67|以撒 就領 利百加 進了母親 撒拉 的帳棚，娶了她為妻，並且愛她。 以撒 自從母親離世以後，這才得了安慰。
GEN|25|1|亞伯拉罕 再娶了一個妻子，名叫 基土拉 。
GEN|25|2|她為他生了 心蘭 、 約珊 、 米但 、 米甸 、 伊施巴 和 書亞 。
GEN|25|3|約珊 生了 示巴 和 底但 。 底但 的子孫是 亞書利 族、 利都是 族和 利烏米 族。
GEN|25|4|米甸 的兒子是 以法 、 以弗 、 哈諾 、 亞比大 和 以勒大 。這些都是 基土拉 的子孫。
GEN|25|5|亞伯拉罕 把他一切所有的都給了 以撒 。
GEN|25|6|至於 亞伯拉罕 妾的兒子， 亞伯拉罕 趁著自己還活著的時候把財物分給他們，打發他們離開他的兒子 以撒 ，往東方去，直到東方之地。
GEN|25|7|這是 亞伯拉罕 一生的年日，他活了一百七十五年。
GEN|25|8|亞伯拉罕 壽高年邁，安享天年，息勞而終，歸到他祖先 那裏。
GEN|25|9|他兩個兒子 以撒 、 以實瑪利 把他安葬在 麥比拉 洞裏。這洞在 幔利 的對面、 赫 人 瑣轄 的兒子 以弗崙 的田中，
GEN|25|10|就是 亞伯拉罕 向 赫 人買的那塊田。 亞伯拉罕 和他妻子 撒拉 都葬在那裏。
GEN|25|11|亞伯拉罕 死了以後，上帝賜福給他的兒子 以撒 。 以撒 住在 庇耳‧拉海‧萊 附近。
GEN|25|12|這是 撒拉 的婢女、 埃及 人 夏甲 為 亞伯拉罕 生的兒子 以實瑪利 的後代。
GEN|25|13|以實瑪利 兒子們的名字，按著他們後代的名字如下： 以實瑪利 的長子 尼拜約 ，又有 基達 、 亞德別 、 米比衫 、
GEN|25|14|米施瑪 、 度瑪 、 瑪撒 、
GEN|25|15|哈大 、 提瑪 、 伊突 、 拿非施 ，和 基底瑪 。
GEN|25|16|這些都是 以實瑪利 的兒子們。他們的村莊和營寨按著他們命名；他們作了十二族的族長。
GEN|25|17|以實瑪利 一生的歲數是一百三十七歲，斷氣而死，歸到他祖先那裏。
GEN|25|18|他的子孫住在 哈腓拉 ，直到 埃及 東邊的 書珥 ，向著 亞述 ，在他眾弟兄的對面安頓下來 。
GEN|25|19|這是 亞伯拉罕 的兒子 以撒 的後代。 亞伯拉罕 生 以撒 。
GEN|25|20|以撒 四十歲時娶 利百加 為妻。 利百加 是 巴旦‧亞蘭 地的 亞蘭 人 彼土利 的女兒，是 亞蘭 人 拉班 的妹妹。
GEN|25|21|以撒 因他妻子不生育，就為她祈求耶和華。耶和華應允他的祈求，他的妻子 利百加 就懷了孕。
GEN|25|22|胎兒們在她腹中彼此相爭，她就說：「若是如此，我為甚麼會這樣呢 ？」她就去求問耶和華。
GEN|25|23|耶和華對她說： 兩國在你腹中； 兩族要從你身上分立。 這族必強於那族； 將來大的要服侍小的。
GEN|25|24|到了生產的日期，看哪，腹中是對雙胞胎。
GEN|25|25|先出生的身體帶紅，渾身有毛，好像皮衣；他們就給他起名叫 以掃 。
GEN|25|26|隨後， 以掃 的弟弟也出生，他的手抓住 以掃 的腳跟，因此給他起名叫 雅各 。兩個兒子出生時， 以撒 六十歲。
GEN|25|27|兩個孩子漸漸長大， 以掃 善於打獵，常在田野； 雅各 為人安靜，常住在帳棚裏。
GEN|25|28|以撒 愛 以掃 ，因為常吃他的野味； 利百加 卻愛 雅各 。
GEN|25|29|有一天， 雅各 熬了湯， 以掃 從田野回來，疲憊不堪。
GEN|25|30|以掃 對 雅各 說：「我累死了，請你讓我吃這紅的，這紅的湯吧！」因此 以掃 又叫 以東 。
GEN|25|31|雅各 說：「你今日把長子的名分賣給我吧。」
GEN|25|32|以掃 說：「看哪，我快要死了，這長子的名分對我有甚麼用呢？」
GEN|25|33|雅各 說：「你今日對我起誓吧。」 以掃 就向他起誓，把長子的名分賣給了 雅各 。
GEN|25|34|於是 雅各 把餅和豆湯給了 以掃 ， 以掃 吃喝以後，起來走了。這樣， 以掃 輕看他長子的名分。
GEN|26|1|那地有了饑荒，不是 亞伯拉罕 的時候曾有過的那次饑荒， 以撒 就到 基拉耳 ， 非利士 人的王 亞比米勒 那裏去。
GEN|26|2|耶和華向 以撒 顯現，說：「你不要下 埃及 去，要住在我所指示你的地。
GEN|26|3|你要寄居在這地，我必與你同在，賜福給你，因為我要將這一切的地都賜給你和你的後裔。我必堅定我向你父親 亞伯拉罕 所起的誓。
GEN|26|4|我要使你的後裔增多，好像天上的星，又要將這一切的地賜給你的後裔，並且地上的萬國都必因你的後裔得福，
GEN|26|5|因為 亞伯拉罕 聽從我的話，遵守我的吩咐、誡令、律例和教導。」
GEN|26|6|於是， 以撒 住在 基拉耳 。
GEN|26|7|那地方的人問起他的妻子，他就說：「她是我的妹妹。」原來他害怕說「我的妻子」。他想：「或許這地方的人會因 利百加 殺我，因為她容貌美麗。」
GEN|26|8|他在那裏住了一段很長的日子。有一天， 非利士 人的王 亞比米勒 從窗戶往外觀看，看哪， 以撒 在撫愛他的妻子 利百加 。
GEN|26|9|亞比米勒 召 以撒 來，說：「看哪，她實在是你的妻子，你怎麼說『她是我的妹妹』呢？」 以撒 對他說：「因為我想，恐怕我會因她而死。」
GEN|26|10|亞比米勒 說：「你向我們做的是甚麼事呢？百姓中有一個人幾乎要和你的妻子同寢，你就把我們陷在罪中了。」
GEN|26|11|於是 亞比米勒 命令眾百姓說：「凡侵犯這個人，或他妻子的，必要把他處死。」
GEN|26|12|以撒 在那地耕種，那一年有百倍的收成。耶和華賜福給他，
GEN|26|13|他就發達，日漸昌盛，成了大富翁。
GEN|26|14|他有羊群牛群，又有許多僕人， 非利士 人就嫉妒他。
GEN|26|15|他父親 亞伯拉罕 在世的時候，他父親的僕人所挖的井， 非利士 人全都塞住，填滿了土。
GEN|26|16|亞比米勒 對 以撒 說：「你離開我們去吧，因為你比我們強盛得多。」
GEN|26|17|以撒 就離開那裏，在 基拉耳谷 支搭帳棚，住在那裏。
GEN|26|18|他父親 亞伯拉罕 在世的時候所挖的水井，在 亞伯拉罕 死後，都被 非利士 人塞住了， 以撒 就重新把井挖出來，仍照他父親所取的名為它們命名。
GEN|26|19|以撒 的僕人在谷中挖井，就在那裏得了一口活水井。
GEN|26|20|基拉耳 的牧人與 以撒 的牧人相爭，說：「這水是我們的。」 以撒 就給那井起名叫 埃色 ，因為他們和他相爭。
GEN|26|21|以撒 的僕人又挖了一口井，他們又為這井相爭， 以撒 就給這井起名叫 西提拿 。
GEN|26|22|以撒 離開那裏，又挖了一口井，他們不再為這井相爭了，他就給那井起名叫 利河伯 。他說：「耶和華現在給我們寬闊之地，我們必在這地興旺。」
GEN|26|23|以撒 從那裏上 別是巴 去。
GEN|26|24|當夜耶和華向他顯現，說：「我是你父親 亞伯拉罕 的上帝。不要懼怕，因為我與你同在，要賜福給你，也要為我僕人 亞伯拉罕 的緣故，使你的後裔增多。」
GEN|26|25|以撒 就在那裏築了一座壇，求告耶和華的名，並且在那裏支搭帳棚；他的僕人就在那裏挖了一口井。
GEN|26|26|亞比米勒 同他的顧問 亞戶撒 和他軍隊的元帥 非各 ，從 基拉耳 來到 以撒 那裏。
GEN|26|27|以撒 對他們說：「你們既然恨我，趕我離開你們，為甚麼又到我這裏來呢？」
GEN|26|28|他們說：「我們明明看見耶和華與你同在；因此就說，讓我們雙方彼此起誓，我們跟你立約，
GEN|26|29|使你不加害我們，正如我們未曾侵犯你，素來善待你，並且送你平平安安地走。你是蒙耶和華賜福的！」
GEN|26|30|以撒 為他們擺設宴席，他們就一起吃喝。
GEN|26|31|他們清早起來，彼此起誓。 以撒 送他們走，他們就平平安安地離開他去了。
GEN|26|32|那一天， 以撒 的僕人來，把挖井的消息告訴他，說：「我們得到水了。」
GEN|26|33|他就給那井起名叫 示巴 ，因此那城名叫 別是巴 ，直到今日。
GEN|26|34|以掃 四十歲的時候娶了 赫 人 比利 的女兒 猶滴 ，和 赫 人 以倫 的女兒 巴實抹 為妻。
GEN|26|35|她們使 以撒 和 利百加 心裏愁煩。
GEN|27|1|以撒 年老，眼睛昏花，不能看見，就叫他大兒子 以掃 來，對他說：「我兒。」 以掃 對他說：「我在這裏。」
GEN|27|2|他說：「看哪，我老了，不知道哪一天死。
GEN|27|3|現在拿你打獵的工具，就是箭囊和弓，到田野去為我打獵，
GEN|27|4|照我所愛的做成美味，拿來給我吃，好讓我在未死之前為你祝福。」
GEN|27|5|以撒 對他兒子 以掃 說話的時候， 利百加 聽見了。 以掃 往田野去打獵，要把獵物帶回來。
GEN|27|6|利百加 就對她兒子 雅各 說：「看哪，我聽見你父親對你哥哥 以掃 說：
GEN|27|7|『你去把獵物帶回來，做成美味給我吃，讓我在未死之前，在耶和華面前為你祝福。』
GEN|27|8|現在，我兒，你要聽我的話，照我所吩咐你的，
GEN|27|9|到羊群裏去，從那裏牽兩隻肥美的小山羊來給我，我就照你父親所愛的，把牠們做成美味給他。
GEN|27|10|然後，你拿到你父親那裏給他吃，好讓他在未死之前為你祝福。」
GEN|27|11|雅各 對他母親 利百加 說：「看哪，我哥哥 以掃 渾身都有毛，我身上卻是光滑的；
GEN|27|12|倘若父親摸著我，我在他眼中就是騙子了。這樣，我就自招詛咒，而不是祝福。」
GEN|27|13|他母親對他說：「我兒，你所受的詛咒臨到我身上吧！你只管聽我的話，去牽小山羊來給我。」
GEN|27|14|他就去牽來，交給他母親。他母親就照他父親所愛的，做成美味。
GEN|27|15|利百加 把大兒子 以掃 在家裏最好的衣服給她小兒子 雅各 穿，
GEN|27|16|又用小山羊的皮包在 雅各 的手上和頸項光滑的地方，
GEN|27|17|就把所做的美味和餅交在她兒子 雅各 的手裏。
GEN|27|18|雅各 來到他父親那裏，說：「我的父親！」他說：「我在這裏。我兒，你是誰？」
GEN|27|19|雅各 對他父親說：「我是你的長子 以掃 。我已照你吩咐我的做了。請起來坐著，吃我的野味，你好為我祝福。」
GEN|27|20|以撒 對他兒子說：「我兒，你怎麼這樣快就找到了呢？」他說：「因為這是耶和華—你的上帝使我遇見的。」
GEN|27|21|以撒 對 雅各 說：「我兒，靠近一點，讓我摸摸你，你真的是我的兒子 以掃 嗎？」
GEN|27|22|雅各 就靠近他父親 以撒 。 以撒 摸著他，說：「聲音是 雅各 的聲音，手卻是 以掃 的手。」
GEN|27|23|以撒 認不出他來，因為他手上有毛，像他哥哥 以掃 的手一樣。於是， 以撒 就為他祝福。
GEN|27|24|以撒 說：「你真的是我兒子 以掃 嗎？」他說：「我是。」
GEN|27|25|以撒 說：「拿給我，讓我吃我兒子的野味，我好為你祝福。」 雅各 拿給他，他就吃了，又拿酒給他，他也喝了。
GEN|27|26|他父親 以撒 對他說：「我兒，靠近一點來親我！」
GEN|27|27|他就近前親吻父親。他父親一聞他衣服上的香氣，就為他祝福，說： 「看，我兒的香氣 好像耶和華賜福之田地的香氣。
GEN|27|28|願上帝賜你天上的甘露， 地上的肥土， 和豐富的五穀新酒。
GEN|27|29|願萬民事奉你， 萬族向你下拜。 願你作你弟兄的主， 你母親的兒子向你下拜。 詛咒你的，願他受詛咒； 祝福你的，願他蒙祝福。」
GEN|27|30|以撒 為 雅各 祝福完畢， 雅各 才從他父親那裏出來，他哥哥 以掃 正打獵回來。
GEN|27|31|以掃 也做了美味，拿來給他父親，對他父親說：「父親，請起來，吃你兒子的野味，你好為我祝福。」
GEN|27|32|他父親 以撒 對他說：「你是誰？」他說：「我是你的兒子，你的長子 以掃 。」
GEN|27|33|以撒 就大大戰兢，說：「那麼，是誰打了獵物拿來給我呢？你未來之前我已經吃了，也為他祝福了，他將來就必蒙福。」
GEN|27|34|以掃 聽了他父親的話，就大聲痛哭，對他父親說：「我父啊，求你也為我祝福！」
GEN|27|35|以撒 說：「你弟弟已經用詭計來把你的福分奪去了。」
GEN|27|36|以掃 說：「他名叫 雅各 ，豈不是這樣嗎？他欺騙了我兩次：他先前奪了我長子的名分，看哪，他現在又奪了我的福分。」 以掃 又說：「你沒有留下給我的祝福嗎？」
GEN|27|37|以撒 回答 以掃 說：「看哪，我已立他作你的主，使他的弟兄都給他作僕人，並賜他五穀新酒可以養生。我兒，那麼，現在我還能為你做甚麼呢？」
GEN|27|38|以掃 對他父親說：「我父啊，你只有一個祝福嗎？我父啊，求你也為我祝福！」 以掃 就放聲而哭。
GEN|27|39|他父親 以撒 回答說： 「看哪，你所住的地方必缺乏肥沃的土地， 缺乏天上的甘露 。
GEN|27|40|你必倚靠刀劍度日， 又必服侍你的兄弟； 到你強盛的時候， 必從你頸項上掙開他的軛。
GEN|27|41|以掃 因他父親給 雅各 的祝福，就怨恨 雅各 ，心裏說：「為我父親居喪的時候近了，到那時候，我要殺我的弟弟 雅各 。」
GEN|27|42|有人把 利百加 大兒子 以掃 的話告訴 利百加 ，她就派人去，叫了她小兒子 雅各 來，對他說：「看哪，你哥哥 以掃 想要殺你來洩恨。
GEN|27|43|現在，我兒，聽我的話，起來，逃往 哈蘭 ，到我哥哥 拉班 那裏去，
GEN|27|44|同他住一段日子，直等到你哥哥的怒氣消了。
GEN|27|45|等到你哥哥向你消了怒氣，忘了你向他所做的事，我就派人去，把你從那裏帶回來。我何必在一天之內喪失你們二人呢？」
GEN|27|46|利百加 對 以撒 說：「我因這 赫 人的女子活得不耐煩了；倘若 雅各 也從本地女子中娶像這樣的 赫 人女子為妻，我為甚麼要活著呢？」
GEN|28|1|以撒 叫了 雅各 來，為他祝福，並吩咐他說：「你不要娶 迦南 的女子為妻。
GEN|28|2|你起身往 巴旦‧亞蘭 去，到你外祖父 彼土利 的家，從你舅父 拉班 的女兒中娶一位作你的妻子。
GEN|28|3|願全能的上帝賜福給你，使你生養眾多，成為許多民族，
GEN|28|4|將應許 亞伯拉罕 的福賜給你和你的後裔，使你承受你所寄居的地為業，就是上帝賜給 亞伯拉罕 的地。」
GEN|28|5|以撒 送 雅各 走了， 雅各 就往 巴旦‧亞蘭 去，到 亞蘭 人 彼土利 的兒子 拉班 那裏， 拉班 是 利百加 的哥哥， 利百加 是 雅各 和 以掃 的母親。
GEN|28|6|以掃 見 以撒 已經為 雅各 祝福，而且送他往 巴旦‧亞蘭 去，在那裏娶妻，並且見 以撒 祝福 雅各 的時候吩咐他說：「不要娶 迦南 的女子為妻」，
GEN|28|7|又見 雅各 聽從父母的話往 巴旦‧亞蘭 去了，
GEN|28|8|以掃 就看出他父親 以撒 看 迦南 女子不順眼。
GEN|28|9|於是他往 以實瑪利 那裏去，在兩個妻子之外， 又娶了 瑪哈拉 為妻，她是 亞伯拉罕 兒子 以實瑪利 的女兒，是 尼拜約 的妹妹。
GEN|28|10|雅各 離開 別是巴 ，往 哈蘭 去。
GEN|28|11|到了一個地方，因為已經日落，就在那裏過夜。他拾起那地方的一塊石頭枕在頭下，就躺在那地方。
GEN|28|12|他做夢，看哪，一個梯子立在地上，梯子的頂端直伸到天；看哪，上帝的使者在梯子上，上去下來。
GEN|28|13|看哪，耶和華站在梯子上面 ，說：「我是耶和華—你祖父 亞伯拉罕 的上帝， 以撒 的上帝。你現在躺臥之地，我要將它賜給你和你的後裔。
GEN|28|14|你的後裔必像地上的塵沙，必向東西南北開展；地上萬族必因你和你的後裔得福。
GEN|28|15|看哪，我必與你同在，無論你往哪裏去，我必保佑你，領你歸回這地。我總不離棄你，直到我實現了對你所說的話。」
GEN|28|16|雅各 睡醒了，說：「耶和華真的在這裏，我竟不知道！」
GEN|28|17|他就懼怕，說：「這地方何等可畏！這不是別的，是上帝的殿，是天的門。」
GEN|28|18|雅各 清早起來，拿起枕在頭下的石頭，立作柱子，澆油在上面。
GEN|28|19|他給那地方起名叫 伯特利 ；那地方原先名叫 路斯 。
GEN|28|20|雅各 許願說：「上帝若與我同在，在我所行的路上保佑我，給我食物吃，衣服穿，
GEN|28|21|使我平平安安回到我父親的家，我就必以耶和華為我的上帝。
GEN|28|22|我所立為柱子的這塊石頭必作上帝的殿；凡你所賜給我的，我必將十分之一獻給你。」
GEN|29|1|雅各 起行，到了東方人之地。
GEN|29|2|他觀看，看哪，田間有一口井，看哪，有三群羊臥在井旁；因為人都取那井裏的水給羊喝。井口上的那塊石頭很大。
GEN|29|3|羊群都在那裏聚集，人就把石頭移開井口，取水給羊喝，然後又把石頭放回井口原處。
GEN|29|4|雅各 對他們說：「弟兄們，你們從哪裏來？」他們說：「我們是從 哈蘭 來的。」
GEN|29|5|他對他們說：「你們認識 拿鶴 的孫子 拉班 嗎？」他們說：「我們認識。」
GEN|29|6|雅各 對他們說：「他平安嗎？」他們說：「平安。看哪，他女兒 拉結 和羊一起來了。」
GEN|29|7|雅各 說：「看哪，日正當中，不是牲畜聚集的時候。你們取水給羊喝，再去牧放吧！」
GEN|29|8|他們說：「我們不能這樣，必須等所有的羊群聚集，人把石頭移開井口，我們才可以取水給羊喝。」
GEN|29|9|雅各 正和他們說話的時候， 拉結 和她父親的羊來了，因為她是牧羊的。
GEN|29|10|雅各 看見他舅父 拉班 的女兒 拉結 和舅父 拉班 的羊群，就上前把石頭移開井口，取水給舅父 拉班 的羊喝。
GEN|29|11|雅各 親了 拉結 ，就放聲大哭。
GEN|29|12|雅各 告訴 拉結 ，自己是她父親的親戚 ，是 利百加 的兒子。 拉結 就跑去告訴她父親。
GEN|29|13|拉班 聽見外甥 雅各 的消息，就跑去迎接他，抱著他，親他，帶他到自己的家。 雅各 把這一切的事告訴 拉班 。
GEN|29|14|拉班 對他說：「你實在是我的骨肉。」 雅各 就和他同住了一個月。
GEN|29|15|拉班 對 雅各 說：「雖然你是我的親戚，怎麼可以讓你白白服事我呢？告訴我，你要甚麼作工資呢？」
GEN|29|16|拉班 有兩個女兒，大的名叫 利亞 ，小的名叫 拉結 。
GEN|29|17|利亞 的雙眼無神， 拉結 卻長得美貌秀麗。
GEN|29|18|雅各 愛 拉結 ，就說：「我願為你的小女兒 拉結 服事你七年。」
GEN|29|19|拉班 說：「我把她給你，勝過給別人，你與我同住吧！」
GEN|29|20|雅各 就為 拉結 服事了七年；他因為愛 拉結 ，就看這七年如同幾天。
GEN|29|21|雅各 對 拉班 說：「日期已經滿了，請把我的妻子給我，我好與她同房。」
GEN|29|22|拉班 就擺設宴席，請了當地所有的人。
GEN|29|23|到了晚上， 拉班 帶女兒 利亞 來送給 雅各 ， 雅各 就與她同房。
GEN|29|24|拉班 也把自己的婢女 悉帕 給女兒 利亞 作婢女。
GEN|29|25|到了早晨，看哪，她是 利亞 ， 雅各 對 拉班 說：「你向我做的是甚麼事呢？我服事你，不是為 拉結 嗎？你為甚麼欺騙我呢？」
GEN|29|26|拉班 說：「大女兒還沒有給人就先把小女兒給人，我們這地方沒有這樣的規矩。
GEN|29|27|你先為這個滿了七日，我們就把那個也給你，不過你要另外再服事我七年。」
GEN|29|28|雅各 就這樣做了。滿了 利亞 的七日， 拉班 就把女兒 拉結 給 雅各 為妻。
GEN|29|29|拉班 又把自己的婢女 辟拉 給女兒 拉結 作婢女。
GEN|29|30|雅各 也與 拉結 同房，並且愛 拉結 勝過愛 利亞 ，於是他又服事了 拉班 七年。
GEN|29|31|耶和華見 利亞 失寵 ，就使她生育， 拉結 卻不生育。
GEN|29|32|利亞 懷孕生子，給他起名叫 呂便 ，因為她說：「耶和華看見我的苦情，如今我的丈夫必愛我。」
GEN|29|33|她又懷孕生子，給他起名叫 西緬 ，說：「耶和華因為聽見我失寵，所以又賜給我這個兒子。」
GEN|29|34|她又懷孕生子，說：「我給丈夫生了三個兒子，現在，這次他必親近我了。」因此， 雅各 給他起名叫 利未 。
GEN|29|35|她又懷孕生子，說：「這次我要讚美耶和華。」因此給他起名叫 猶大 。於是她停了生育。
GEN|30|1|拉結 見自己不給 雅各 生孩子，就嫉妒她姊姊，對 雅各 說：「你給我孩子，不然，讓我死了吧。」
GEN|30|2|雅各 對 拉結 生氣，說：「是我代替上帝使你生不出孩子的嗎？」
GEN|30|3|拉結 說：「看哪，我的使女 辟拉 在這裏，你可以與她同房，使她生子歸在我膝下，我也可以藉著她得孩子 。」
GEN|30|4|拉結 就把她的婢女 辟拉 給丈夫為妾， 雅各 與她同房。
GEN|30|5|辟拉 懷孕，為 雅各 生了一個兒子。
GEN|30|6|拉結 給他起名叫 但 ，說：「上帝為我伸冤，也聽了我的聲音，賜給我一個兒子。」
GEN|30|7|拉結 的婢女 辟拉 又懷孕，為 雅各 生了第二個兒子。
GEN|30|8|拉結 給他起名叫 拿弗他利 ，說：「我與我姊姊大大較力，並且得勝了。」
GEN|30|9|利亞 見自己停了生育，就把她的婢女 悉帕 給 雅各 為妾。
GEN|30|10|利亞 的婢女 悉帕 為 雅各 生了一個兒子。
GEN|30|11|利亞 給他起名叫 迦得 ，說：「真是幸運！」
GEN|30|12|利亞 的婢女 悉帕 又為 雅各 生了第二個兒子。
GEN|30|13|利亞 給他起名叫 亞設 ，說：「我真有福啊，眾女子都要稱我有福。」
GEN|30|14|收割麥子的時候， 呂便 到田裏去，找到曼陀羅草 ，就拿給他的母親 利亞 。 拉結 對 利亞 說：「請你給我一些你兒子的曼陀羅草吧。」
GEN|30|15|利亞 對她說：「你奪走了我的丈夫還是小事嗎？你還要奪取我兒子的曼陀羅草嗎？」 拉結 說：「今夜他可以與你同寢，來交換你兒子的曼陀羅草。」
GEN|30|16|到了晚上， 雅各 從田裏回來， 利亞 出來迎接他，說：「你要與我同寢，因為我真的用我兒子的曼陀羅草把你雇下了。」那一夜， 雅各 就與她同寢。
GEN|30|17|上帝應允了 利亞 ，她就懷孕，為 雅各 生了第五個兒子。
GEN|30|18|利亞 給他起名叫 以薩迦 ，說：「上帝給了我工價，因為我把婢女給了我的丈夫。」
GEN|30|19|利亞 又懷孕，為 雅各 生了第六個兒子。
GEN|30|20|利亞 給他起名叫 西布倫 ，說：「上帝賜給我厚禮了；這次，我丈夫必看重我，因為我為他生了六個兒子。」
GEN|30|21|後來她又生了一個女兒，給她起名叫 底拿 。
GEN|30|22|上帝顧念 拉結 ，應允她，使她能生育。
GEN|30|23|拉結 懷孕生子，說：「上帝除去了我的羞恥。」
GEN|30|24|拉結 就給他起名叫 約瑟 ，說：「願耶和華再增添一個兒子給我。」
GEN|30|25|拉結 生 約瑟 之後， 雅各 對 拉班 說：「請讓我走，回到我的本鄉本土去。
GEN|30|26|請你把我服事你所得的妻子和孩子給我，讓我走吧！我怎樣服事你，你都知道。」
GEN|30|27|拉班 對他說：「願你看得起我，因我占卜得知，耶和華賜福給我是因你的緣故。」
GEN|30|28|又說：「請為我定你的工資，我就給你。」
GEN|30|29|雅各 對他說：「我怎樣服事你，你的牲畜在我這裏變得怎樣，你都知道。
GEN|30|30|我未來以前，你擁有的很少，現在卻已大量增加，因為耶和華隨著我的腳步賜福給你。現在，我到甚麼時候才可以成家立業呢？」
GEN|30|31|拉班 說：「我該給你甚麼呢？」 雅各 說：「你甚麼也不必給我，只要你為我做這件事，我就繼續牧放你的羊群。
GEN|30|32|今天我要走遍你的羊群，把綿羊中凡有點的、有斑的，和小綿羊中凡是黑色的羊；以及山羊中凡有斑的、有點的，都從那裏挑出來，作為我的工資。
GEN|30|33|以後你來當面查看我的工資，任何我這裏的山羊不是有點有斑的，小綿羊不是黑色的，就算是我偷的。這就可以證明我是正直的。」
GEN|30|34|拉班 說：「看哪，就照你所說的做吧。」
GEN|30|35|當日， 拉班 把有紋的、有斑的公山羊，一切有點的、有斑的、有少許白色 的母山羊，以及小綿羊中所有黑色的 ，都挑出來，交在他兒子們的手裏，
GEN|30|36|又使自己和 雅各 相隔三天的路程。 雅各 就牧放 拉班 其餘的羊。
GEN|30|37|雅各 拿楊樹、杏樹、楓樹的嫩枝，把皮剝出白色的條紋，使枝子露出白色來。
GEN|30|38|他把剝了皮的枝子對著羊群，插在羊喝水的水溝和水槽裏。羊來喝水的時候，牠們彼此交配。
GEN|30|39|羊對著枝子交配，就生下有紋的、有點的、有斑的來。
GEN|30|40|雅各 把小綿羊分出來，讓羊對著 拉班 羊群中有紋的和所有黑色的。於是他把自己的羊群分開，不叫牠們和 拉班 的羊混在一起。
GEN|30|41|當肥壯的羊交配的時候， 雅各 就把枝子插在水溝裏，使羊對著枝子交配。
GEN|30|42|可是當瘦弱的羊交配的時候，他就不插枝子。這樣，瘦弱的就歸 拉班 ，肥壯的就歸 雅各 。
GEN|30|43|於是這人極其發達，擁有許多的羊群、奴僕、婢女、駱駝和驢。
GEN|31|1|雅各 聽見 拉班 兒子們的話，說：「 雅各 把我們父親所有的都奪去了！他從我們父親所擁有的獲得這一切的財富。」
GEN|31|2|雅各 見 拉班 的臉色，看哪，待他不如從前了。
GEN|31|3|耶和華對 雅各 說：「你要回你祖先之地，到你本族那裏去，我必與你同在。」
GEN|31|4|雅各 就派人叫 拉結 和 利亞 到田野他的羊群那裏去，
GEN|31|5|對她們說：「我看你們父親待我的臉色不如從前了，但我父親的上帝向來與我同在。
GEN|31|6|你們也知道，我盡了全力服事你們的父親。
GEN|31|7|可是你們的父親欺騙我，十次更改我的工資，但上帝不容許他害我。
GEN|31|8|他若說：『有點的歸給你作工資』，羊群所生的都是有點的；他若說：『有紋的歸給你作工資』，羊群所生的都是有紋的。
GEN|31|9|這樣，上帝把你們父親的牲畜拿來賜給我了。
GEN|31|10|「羊群交配的時候，我在夢中舉目一看，看哪，跳母羊的公羊都是有紋的、有點的、有花斑的。
GEN|31|11|上帝的使者在夢中呼叫我說：『 雅各 。』我說：『我在這裏。』
GEN|31|12|他說：『你舉目觀看，跳母羊的公羊都是有紋的、有點的、有花斑的。 拉班 向你所做的一切，我都看見了。
GEN|31|13|我是 伯特利 的上帝；你曾在那裏用油膏過柱子，向我許過願。現在你起來，離開這地，回你本族之地去吧！』」
GEN|31|14|拉結 和 利亞 回答 雅各 說：「在我們父親家裏還有我們可分得的產業嗎？
GEN|31|15|我們不是被他看作外人嗎？因為他賣了我們，還吞吃了我們的銀錢。
GEN|31|16|上帝從我們父親所拿走的一切財物，都是我們和我們孩子的。現在，凡上帝所吩咐你的，你只管去做吧！」
GEN|31|17|雅各 起來，叫他的孩子和妻子都騎上駱駝，
GEN|31|18|又趕著他一切的牲畜和他所得的一切財物，就是他在 巴旦‧亞蘭 所得的，他擁有的牲畜 ，往 迦南 地他父親 以撒 那裏去了。
GEN|31|19|當時 拉班 去剪羊毛， 拉結 偷了他父親家中的神像。
GEN|31|20|雅各 瞞住 亞蘭 人 拉班 ，不通知他就逃走了。
GEN|31|21|雅各 帶著他所有的逃走了；他起程，渡過 大河 ，面向著 基列山 。
GEN|31|22|到第三天，有人告訴 拉班 ， 雅各 逃跑了。
GEN|31|23|拉班 帶著他的弟兄們去追他，追了七天，就在 基列山 追上了。
GEN|31|24|夜間，上帝來到 亞蘭 人 拉班 那裏，在夢中對他說：「你要小心，不可對 雅各 說好說歹。」
GEN|31|25|拉班 追上 雅各 。 雅各 在山上支搭帳棚； 拉班 和他的弟兄們也在 基列山 上支搭帳棚。
GEN|31|26|拉班 對 雅各 說：「你做的是甚麼事呢？你瞞著我把我的女兒們帶走，好像用刀劍擄去一般。
GEN|31|27|你為甚麼暗暗地逃跑，瞞著我，不通知我一聲，叫我可以歡樂、唱歌、擊鼓、彈琴送你回去呢？
GEN|31|28|為甚麼不容許我與外孫和女兒吻別呢？你現在所做的真是愚蠢！
GEN|31|29|我的手本有能力害你，只是你父親的上帝昨夜對我說：『你要小心，不可對 雅各 說好說歹。』
GEN|31|30|現在你既然這麼想念你的父家，不得不去，為甚麼又偷了我的神明呢？」
GEN|31|31|雅各 回答 拉班 說：「因為我害怕，我想，恐怕你把你的女兒從我這裏奪走。
GEN|31|32|至於你的神明，你若在誰那裏搜出來，就不讓誰活。當著我們弟兄面前，你認一認在我這裏有甚麼東西是你的，你就拿去吧。」原來 雅各 並不知道 拉結 偷了神明。
GEN|31|33|拉班 進了 雅各 、 利亞 ，以及兩個使女的帳棚，卻沒有找到，就從 利亞 的帳棚出來，進入 拉結 的帳棚。
GEN|31|34|拉結 拿了神像，藏在駱駝的鞍子裏，自己坐在上面。 拉班 搜遍了那帳棚，並沒有找到。
GEN|31|35|拉結 對她父親說：「請我主不要生氣，因為我恰有月事，不能在你面前起來。」 拉班 搜尋，卻找不到神像。
GEN|31|36|於是 雅各 發怒，斥責 拉班 。 雅各 對 拉班 說：「我有甚麼過犯，有甚麼罪惡，你竟這樣火速地追我？
GEN|31|37|你搜遍了我一切的物件，你找到甚麼呢？可以放在你我弟兄面前，叫他們在我們兩個之間評評理。
GEN|31|38|我在你那裏這二十年，你的母綿羊、母山羊沒有掉過胎。你羊群中的公綿羊，我沒有吃過；
GEN|31|39|被野獸撕裂的，我沒有帶來給你，是我自己賠償的。無論是白日被偷的，或是黑夜被偷的，你都從我手中索取。
GEN|31|40|我常常白日受盡炎熱，黑夜受盡寒霜，不得合眼入睡。
GEN|31|41|我這二十年在你家裏，為你兩個女兒服事了你十四年，為你的羊群服事了你六年，你卻十次更改我的工資。
GEN|31|42|若不是我父親 以撒 所敬畏的上帝，就是 亞伯拉罕 的上帝與我同在，你如今必定打發我空手而去。上帝看見我的苦情和我手的辛勞，就在昨夜責備了你。」
GEN|31|43|拉班 回答 雅各 說：「這兩個女兒是我的女兒，這些孩子是我的孩子，這些羊群也都是我的羊群；凡你所看見的都是我的。我的女兒和她們所生的孩子，我今日還能對他們做甚麼呢？
GEN|31|44|現在，來吧！讓我和你立約，作你我之間的證據。」
GEN|31|45|雅各 就拿一塊石頭立作柱子，
GEN|31|46|對弟兄們說：「大家來堆積石頭。」他們拿石頭堆成一堆，於是在那裏，在石堆旁邊吃喝。
GEN|31|47|拉班 稱那石堆為 伊迦爾‧撒哈杜他 ， 雅各 卻稱那石堆為 迦累得 。
GEN|31|48|拉班 說：「今日這石堆成為你我之間的證據。」因此這地方名叫 迦累得 ，
GEN|31|49|又叫 米斯巴 ，因為他說：「我們彼此離別以後，願耶和華在你我中間鑒察 。
GEN|31|50|你若苦待我的女兒，或在我的女兒以外另娶妻，雖沒有人在場，你看，有上帝在你我中間作證。」
GEN|31|51|拉班 又對 雅各 說：「看哪，這石堆，看哪，這柱子，是我在你我中間所立的。
GEN|31|52|這石堆是證據，這柱子也是證據。我必不越過這石堆去害你；你也不可越過這石堆和柱子來害我。
GEN|31|53|願 亞伯拉罕 的上帝和 拿鶴 的上帝，就是他們父親的上帝 ，在你我中間判斷。」 雅各 就指著他父親 以撒 所敬畏的上帝起誓，
GEN|31|54|又在山上獻祭，請弟兄們來吃飯。他們吃了飯，就在山上過夜。
GEN|31|55|拉班 清早起來，與他外孫和女兒親吻，為他們祝福，就回到自己的地方去了。
GEN|32|1|雅各 繼續行路，上帝的使者遇見他。
GEN|32|2|雅各 看見他們就說：「這是上帝的軍營。」於是給那地方起名叫 瑪哈念 。
GEN|32|3|雅各 派使者在他前面到 西珥 地，就是 以東 地他哥哥 以掃 那裏。
GEN|32|4|他吩咐他們說：「你們要對我主 以掃 說：『你的僕人 雅各 這樣說：我在 拉班 那裏寄居，延遲到如今。
GEN|32|5|我有牛、驢、羊群、奴僕、婢女，現在派人來報告我主，為了要在你眼前蒙恩。』」
GEN|32|6|使者回到 雅各 那裏，說：「我們到了你哥哥 以掃 那裏。他正迎著你來，並且有四百人和他一起。」
GEN|32|7|雅各 就很懼怕，而且愁煩。他把跟他同行的人和羊群、牛群、駱駝分成兩隊，
GEN|32|8|說：「 以掃 若來擊殺其中一隊，剩下的另一隊還可以逃脫。」
GEN|32|9|雅各 說：「耶和華—我祖父 亞伯拉罕 的上帝，我父親 以撒 的上帝啊，你曾對我說：『回你本地本族去，我要厚待你。』
GEN|32|10|你向僕人所施的一切慈愛和信實，我一點也不配得。我先前只用我的一根杖過這 約旦河 ，如今我卻成了兩隊。
GEN|32|11|求你救我脫離我哥哥的手，脫離 以掃 的手，因為我怕他來殺我，連母親和兒女都不放過。
GEN|32|12|你曾說：『我必定厚待你，使你的後裔如同海邊的沙，多得不可勝數。』」
GEN|32|13|當夜， 雅各 在那裏住宿，就從他手中所擁有的拿禮物要送給他哥哥 以掃 ，
GEN|32|14|就是二百隻母山羊、二十隻公山羊、二百隻母綿羊、二十隻公綿羊、
GEN|32|15|三十匹哺乳的母駱駝和牠們的小駱駝、四十頭母牛、十頭公牛、二十匹母驢和十匹公驢。
GEN|32|16|他把每種牲畜各分一群，交在僕人手中，對僕人說：「你們要在我的前頭過去，使群和群之間保持一段距離」。
GEN|32|17|他又吩咐領頭的人說：「我哥哥 以掃 遇見你的時候，問你說：『你是誰的人？要往哪裏去？你前面這些是誰的？』
GEN|32|18|你就說：『是你僕人 雅各 的，是送給我主 以掃 的禮物。看哪，他自己也在我們後面。』」
GEN|32|19|他又吩咐第二、第三和所有趕畜群的人說：「你們遇見 以掃 的時候要照這樣的話對他說，
GEN|32|20|你們還要說：『看哪，你僕人 雅各 在我們後面。』」因 雅各 說：「我藉著在我前面送去的禮物給他面子，然後再見他的面，或許他會寬容我。」
GEN|32|21|於是禮物在他前面過去了；那夜， 雅各 在營中住宿。
GEN|32|22|他夜間起來，帶著兩個妻子，兩個婢女和十一個孩子，過了 雅博 渡口。
GEN|32|23|他帶著他們，送他們過河，他所有的一切也都過去，
GEN|32|24|只剩下 雅各 一人。有一個人來和他摔跤，直到黎明。
GEN|32|25|那人見自己勝不過他，就摸了他的大腿窩一下。 雅各 的大腿窩就在和那人摔跤的時候扭了。
GEN|32|26|那人說：「天快亮了，讓我走吧！」 雅各 說：「你不給我祝福，我就不讓你走。」
GEN|32|27|那人說：「你叫甚麼名字？」他說：「 雅各 。」
GEN|32|28|那人說：「你的名字不要再叫 雅各 ，要叫 以色列 ，因為你與上帝和人較力，都得勝了。」
GEN|32|29|雅各 問他說：「請告訴我你的名字。」那人說：「何必問我的名字呢？」於是他在那裏為 雅各 祝福。
GEN|32|30|雅各 就給那地方起名叫 毗努伊勒 ，說：「我面對面見了上帝，我的性命仍得保全。」
GEN|32|31|太陽剛出來的時候， 雅各 經過 毗努伊勒 ，他的大腿就瘸了。
GEN|32|32|因此， 以色列 人不吃大腿窩的筋，直到今日，因為那人摸了 雅各 大腿窩的筋。
GEN|33|1|雅各 舉目觀看，看哪， 以掃 來了，有四百人和他一起。 雅各 就把孩子們分開交給 利亞 、 拉結 和兩個婢女。
GEN|33|2|他叫兩個婢女和她們的孩子走在前頭， 利亞 和她的孩子跟在後面，而 拉結 和 約瑟 在最後。
GEN|33|3|他自己卻走到他們前面，一連七次俯伏在地才挨近他哥哥。
GEN|33|4|以掃 跑來迎接他，將他抱住，伏在他的頸項上親他，他們都哭了。
GEN|33|5|以掃 舉目看見婦人和孩子，就說：「這些和你一起的是誰呢？」 雅各 說：「這些孩子是上帝施恩給你僕人的。」
GEN|33|6|於是兩個婢女和她們的孩子前來下拜，
GEN|33|7|利亞 和她的孩子也前來下拜，隨後 約瑟 和 拉結 也前來下拜。
GEN|33|8|以掃 說：「我所遇見的這些畜群是甚麼意思呢？」 雅各 說：「是為了要在我主眼前蒙恩。」
GEN|33|9|以掃 說：「弟弟啊，我的已經夠了，你的你自己留著吧！」
GEN|33|10|雅各 說：「不，我若在你眼前蒙恩，就請你從我手裏收下這禮物；因為我見了你的面，如同見了上帝的面，並且你也寬容了我。
GEN|33|11|請你收下我帶來給你的禮物，因為上帝恩待我，使我一切都充足。」 雅各 再三求他，他才收下。
GEN|33|12|以掃 說：「讓我們起身前行，我和你一起走吧。」
GEN|33|13|雅各 對他說：「我主知道孩子們還年幼嬌嫩，我的牛羊也正在哺乳中，只要催趕一天，群羊都會死了。
GEN|33|14|請我主在僕人前面先走，我要按著在我面前的牲畜和孩子的步伐慢慢前進，直走到 西珥 我主那裏。」
GEN|33|15|以掃 說：「讓我把跟隨我的人留幾個在你這裏。」 雅各 說：「何必這樣呢？只要能在我主眼前蒙恩就夠了。」
GEN|33|16|於是， 以掃 當日起行，回 西珥 去了。
GEN|33|17|雅各 就往 疏割 去，在那裏為自己蓋房屋，又為牲畜搭棚，因此那地方叫 疏割 。
GEN|33|18|雅各 從 巴旦‧亞蘭 平安地回到 迦南 地的 示劍城 ，他在城的前面支搭帳棚。
GEN|33|19|他用一百可錫塔 從 示劍 的父親 哈抹 的眾子手中買了搭帳棚的那塊地。
GEN|33|20|雅各 在那裏築了一座壇，起名叫 伊利‧伊羅伊‧以色列 。
GEN|34|1|利亞 給 雅各 所生的女兒 底拿 出去，要探望那地的女子們。
GEN|34|2|那地的族長 希未 人 哈抹 的兒子 示劍 看見她，就拉住她，與她同寢，玷辱了她。
GEN|34|3|示劍 的心喜歡 雅各 的女兒 底拿 ，愛上這少女，甜言蜜語地安慰她。
GEN|34|4|示劍 對他父親 哈抹 說：「求你為我聘這女孩為妻。」
GEN|34|5|雅各 聽見 示劍 污辱了他的女兒 底拿 。那時他的兒子們正和牲畜在田野， 雅各 就沉默，等他們回來。
GEN|34|6|示劍 的父親 哈抹 出來，到 雅各 那裏，要和他講話。
GEN|34|7|雅各 的兒子們聽見這事，就從田野回來，人人悲憤，十分惱怒，因 示劍 在 以色列 中做了醜事，與 雅各 的女兒同寢，這本是不該做的事。
GEN|34|8|哈抹 和他們談話，說：「我兒子 示劍 的心喜歡你們家的女兒，請你們把她嫁給我的兒子。
GEN|34|9|你們與我們彼此結親；你們可以把你們家的女兒嫁給我們，也可以娶我們家的女兒。
GEN|34|10|你們與我們同住吧！這地都在你們面前，只管在這裏居住，做買賣，置產業。」
GEN|34|11|示劍 對女子的父親和兄弟們說：「願你們看得起我，你們向我要甚麼，我必給你們，
GEN|34|12|無論向我要多貴重的聘金和禮物，我必照你們所說的給你們，只要你們將這少女嫁給我。」
GEN|34|13|雅各 的兒子們因 示劍 污辱了他們的妹妹 底拿 ，就用詭詐的話回答 示劍 和他父親 哈抹 ，
GEN|34|14|對他們說：「我們不能做這樣的事，把我們的妹妹嫁給沒有受割禮的人為妻，因為那是我們的羞恥。
GEN|34|15|惟有一個條件，我們才答應你們，就是你們所有的男丁都要受割禮，和我們一樣，
GEN|34|16|我們就把我們家的女兒嫁給你們，也娶你們家的女兒；我們就與你們同住，大家成為一族人。
GEN|34|17|倘若你們不聽從我們受割禮，我們就帶我們家的女兒走了。」
GEN|34|18|這些話在 哈抹 和他兒子 示劍 的眼中看為美。
GEN|34|19|那年輕人毫不遲延做這事，因為他愛上了 雅各 的女兒；他在他父親家中也是最受人尊重的。
GEN|34|20|哈抹 和他兒子 示劍 到他們的城門口，對城裏的人講說：
GEN|34|21|「這些人對我們友善，不如允許他們在這地居住，做買賣；看哪，這地寬闊，足以容納他們。我們可以娶他們家的女兒，也可以把我們家的女兒嫁給他們。
GEN|34|22|惟有一個條件，這些人才答應和我們同住，成為一族人，就是我們中間所有的男丁都要受割禮，和他們一樣。
GEN|34|23|他們的牲畜、財物和一切的牲口豈不都歸給我們嗎？只要答應他們，他們就與我們同住。」
GEN|34|24|凡從城門出入的人都聽從了 哈抹 和他兒子 示劍 的話。於是，凡從城門出入的男丁都受了割禮。
GEN|34|25|到第三天，他們正疼痛的時候， 雅各 的兩個兒子，就是 底拿 的哥哥 西緬 和 利未 ，各拿刀劍，不動聲色地來到城中，把所有的男丁都殺了，
GEN|34|26|又用刀殺了 哈抹 和他兒子 示劍 ，把 底拿 從 示劍 家裏帶走，就離開了。
GEN|34|27|雅各 的兒子們因為他們的妹妹受污辱，就來到被殺的人那裏，洗劫那城，
GEN|34|28|奪走了他們的羊群、牛群和驢，以及城裏和田間所有的；
GEN|34|29|又俘擄搶劫他們一切的財物、孩童、婦女，以及房屋中所有的。
GEN|34|30|雅各 對 西緬 和 利未 說：「你們連累了我，使我在這地的居民中，就是在 迦南 人和 比利洗 人中壞了名聲。我的人丁稀少，他們必聚集來擊殺我，我和全家的人都要被滅絕。」
GEN|34|31|他們卻說：「他豈可待我們的妹妹如同妓女呢？」
GEN|35|1|上帝對 雅各 說：「起來！上 伯特利 去，住在那裏。在那裏築一座壇給上帝，就是你逃避你哥哥 以掃 的時候向你顯現的上帝。」
GEN|35|2|雅各 就對他家中的人，以及所有和他一起的人說：「除掉你們中間外邦的神明，要自潔，更換衣服。
GEN|35|3|我們要起來，上 伯特利 去，在那裏我要築一座壇給上帝，就是在我遭難的日子應允我，在我行走的路上與我同在的上帝。」
GEN|35|4|他們就把手中所有外邦的神明和自己耳朵上的環子交給 雅各 ； 雅各 把它們埋在 示劍 那裏的橡樹下。
GEN|35|5|他們起行。上帝使周圍城鎮的人都驚恐，就不追趕 雅各 的兒子們了。
GEN|35|6|於是 雅各 和所有與他一起的人到了 迦南 地的 路斯 ，就是 伯特利 。
GEN|35|7|他在那裏築了一座壇，給那地方起名叫 伊勒‧伯特利 ，因為他逃避他哥哥的時候，上帝曾在那裏向他顯現。
GEN|35|8|利百加 的奶媽 底波拉 死了，葬在 伯特利 下邊的橡樹下；那棵樹名叫 亞倫‧巴古 。
GEN|35|9|雅各 從 巴旦‧亞蘭 回來，上帝又向他顯現，賜福給他。
GEN|35|10|上帝對他說：「你的名原是 雅各 ，從今以後不要再叫 雅各 ，你的名要叫 以色列 。」於是，上帝就叫他的名為 以色列 。
GEN|35|11|上帝又對他說：「我是全能的上帝；你要生養眾多，將來有一國和許多的國從你而來，又有許多君王從你生出 。
GEN|35|12|至於我賜給 亞伯拉罕 和 以撒 的地，我必賜給你；我必賜這地給你的後裔。」
GEN|35|13|上帝就從與 雅各 說話的那地方升上去了。
GEN|35|14|雅各 就在上帝與他說話的地方立了一根柱子，就是石柱，在它上面獻澆酒祭，又澆油。
GEN|35|15|雅各 就給上帝與他說話的那地方起名叫 伯特利 。
GEN|35|16|他們從 伯特利 起行，到 以法他 還有一段路程， 拉結 生產，生得十分艱難。
GEN|35|17|她生得十分艱難的時候，接生婆對她說：「不要怕，你又要有一個兒子了。」
GEN|35|18|她快要死，還有一口氣的時候，就給她兒子起名叫 便‧俄尼 ；他父親卻給他起名叫 便雅憫 。
GEN|35|19|拉結 死了，葬在往 以法他 的路旁； 以法他 就是 伯利恆 。
GEN|35|20|雅各 在她的墳上立了一塊碑，就是 拉結 的墓碑，到今日還在。
GEN|35|21|以色列 起行，在 以得臺 的那一邊支搭帳棚。
GEN|35|22|以色列 住在那地的時候， 呂便 去與他父親的妾 辟拉 同寢， 以色列 也聽見了這件事 。 雅各 共有十二個兒子。
GEN|35|23|利亞 的兒子是 雅各 的長子 呂便 ，還有 西緬 、 利未 、 猶大 、 以薩迦 、 西布倫 。
GEN|35|24|拉結 的兒子是 約瑟 、 便雅憫 。
GEN|35|25|拉結 的婢女 辟拉 的兒子是 但 、 拿弗他利 。
GEN|35|26|利亞 的婢女 悉帕 的兒子是 迦得 、 亞設 。這是 雅各 在 巴旦‧亞蘭 所生的兒子。
GEN|35|27|雅各 來到他父親 以撒 那裏，到了 幔利 ， 基列‧亞巴 ，就是 希伯崙 ，是 亞伯拉罕 和 以撒 寄居的地方。
GEN|35|28|以撒 共活了一百八十年。
GEN|35|29|以撒 年紀老邁，安享天年，息勞而終，歸到他祖先 那裏。他兩個兒子 以掃 和 雅各 把他安葬了。
GEN|36|1|這是 以掃 的後代， 以掃 就是 以東 。
GEN|36|2|以掃 娶 迦南 的女子為妻，就是 赫 人 以倫 的女兒 亞大 和 希未 人 祭便 的孫女， 亞拿 的女兒 阿何利巴瑪 ，
GEN|36|3|又娶了 以實瑪利 的女兒， 尼拜約 的妹妹 巴實抹 。
GEN|36|4|亞大 為 以掃 生了 以利法 ； 巴實抹 生了 流珥 ；
GEN|36|5|阿何利巴瑪 生了 耶烏施 、 雅蘭 、 可拉 。這些都是 以掃 的兒子，是在 迦南 地生的。
GEN|36|6|以掃 帶著他的妻子、兒女和家中所有的人，以及他的牛羊、牲畜和一切財物，就是他在 迦南 地所得的，往別處去，離開了他的兄弟 雅各 。
GEN|36|7|因為他們擁有的很多，不能住在一起。因為牲畜的緣故，寄居的地方容不下他們。
GEN|36|8|於是 以掃 住在 西珥山 ； 以掃 就是 以東 。
GEN|36|9|這是 以掃 的後代，他是 西珥山 裏 以東 人的始祖。
GEN|36|10|以掃 子孫的名字如下： 以掃 的妻子 亞大 生 以利法 ； 以掃 的妻子 巴實抹 生 流珥 。
GEN|36|11|以利法 的兒子是 提幔 、 阿抹 、 洗玻 、 迦坦 、 基納斯 。
GEN|36|12|亭納 是 以掃 兒子 以利法 的妾，她為 以利法 生了 亞瑪力 。這是 以掃 的妻子 亞大 的子孫。
GEN|36|13|流珥 的兒子是 拿哈 、 謝拉 、 沙瑪 、 米撒 。這是 以掃 妻子 巴實抹 的子孫。
GEN|36|14|以掃 的妻子 阿何利巴瑪 是 祭便 的孫女， 亞拿 的女兒。她為 以掃 生了 耶烏施 、 雅蘭 、 可拉 。
GEN|36|15|這是 以掃 子孫中作族長的： 以掃 的長子 以利法 的子孫中，有 提幔 族長、 阿抹 族長、 洗玻 族長、 基納斯 族長、
GEN|36|16|可拉 族長、 迦坦 族長、 亞瑪力 族長。這是在 以東 地，從 以利法 所出的族長，是 亞大 的子孫。
GEN|36|17|以掃 的兒子 流珥 的子孫中，有 拿哈 族長、 謝拉 族長、 沙瑪 族長、 米撒 族長。這是在 以東 地，從 流珥 所出的族長，是 以掃 妻子 巴實抹 的子孫。
GEN|36|18|以掃 的妻子 阿何利巴瑪 的子孫中，有 耶烏施 族長、 雅蘭 族長、 可拉 族長。這是從 以掃 的妻子， 亞拿 的女兒 阿何利巴瑪 的子孫中所出的族長。
GEN|36|19|以上的族長都是 以掃 的子孫； 以掃 就是 以東 。
GEN|36|20|這是那地原來的居民， 何利 人 西珥 的子孫： 羅坍 、 朔巴 、 祭便 、 亞拿 、
GEN|36|21|底順 、 以察 、 底珊 。這是在 以東 地，從 何利 人 西珥 子孫中所出的族長。
GEN|36|22|羅坍 的兒子是 何利 、 希幔 ， 羅坍 的妹妹是 亭納 。
GEN|36|23|朔巴 的兒子是 亞勒文 、 瑪拿轄 、 以巴錄 、 示玻 、 阿南 。
GEN|36|24|祭便 的兒子是 愛亞 、 亞拿 ，當時在曠野牧放他父親 祭便 的驢，發現溫泉的就是這 亞拿 。
GEN|36|25|亞拿 的兒子是 底順 ， 亞拿 的女兒是 阿何利巴瑪 。
GEN|36|26|底順 的兒子是 欣但 、 伊是班 、 益蘭 、 基蘭 。
GEN|36|27|以察 的兒子是 辟罕 、 撒番 、 亞干 。
GEN|36|28|底珊 的兒子是 烏斯 、 亞蘭 。
GEN|36|29|這是從 何利 人所出的族長： 羅坍 族長、 朔巴 族長、 祭便 族長、 亞拿 族長、
GEN|36|30|底順 族長、 以察 族長、 底珊 族長。這是從 何利 人所出的族長，都在 西珥 地，按著族長 來分。
GEN|36|31|以色列 未有君王治理之前，這些是在 以東 地作王的。
GEN|36|32|比珥 的兒子 比拉 在 以東 作王，他的城名叫 亭哈巴 。
GEN|36|33|比拉 死了， 波斯拉 人 謝拉 的兒子 約巴 接續他作王。
GEN|36|34|約巴 死了， 提幔 人之地的 戶珊 接續他作王。
GEN|36|35|戶珊 死了， 比達 的兒子 哈達 接續他作王， 哈達 曾在 摩押 地擊敗 米甸 人，他的城名叫 亞未得 。
GEN|36|36|哈達 死了， 瑪士利加 人 桑拉 接續他作王。
GEN|36|37|桑拉 死了， 大河 邊的 利河伯 人 掃羅 接續他作王。
GEN|36|38|掃羅 死了， 亞革波 的兒子 巴勒‧哈南 接續他作王。
GEN|36|39|亞革波 的兒子 巴勒‧哈南 死了， 哈達爾 接續他作王，他的城名叫 巴烏 。他的妻子名叫 米希她別 ，是 米‧薩合 的孫女， 瑪特列 的女兒。
GEN|36|40|這些是 以掃 的族長，按著他們的宗族、住處和名字： 亭納 族長、 亞勒瓦 族長、 耶帖 族長、
GEN|36|41|阿何利巴瑪 族長、 以拉 族長、 比嫩 族長、
GEN|36|42|基納斯 族長、 提幔 族長、 米比薩 族長、
GEN|36|43|瑪基疊 族長、 以蘭 族長。這些是 以東 人在所得為業的地上，按著他們住處的族長。 以掃 是 以東 人的始祖。
GEN|37|1|雅各 住在 迦南 地，就是他父親寄居的地。
GEN|37|2|這是 雅各 的事蹟。 約瑟 十七歲與他哥哥們一同牧羊。他是個少年，與他父親的妾 辟拉 和 悉帕 的兒子們常在一起。 約瑟 把他們的惡行報給父親。
GEN|37|3|以色列 愛 約瑟 過於其他的兒子，因為 約瑟 是他年老生的；他給 約瑟 做了一件長袍 。
GEN|37|4|哥哥們見父親愛 約瑟 過於他們，就恨 約瑟 ，不與他說友善的話。
GEN|37|5|約瑟 做了一個夢，告訴他哥哥們，他們就更加恨他。
GEN|37|6|約瑟 對他們說：「請聽我做的這個夢：
GEN|37|7|看哪，我們在田裏捆禾稼；看哪，我的捆起來站著；看哪，你們的捆圍著我的捆下拜。」
GEN|37|8|他的哥哥們對他說：「難道你真的要作我們的王嗎？難道你真的要統治我們嗎？」他們就因他的夢和他的話更加恨他。
GEN|37|9|後來他又做了另一個夢，告訴他哥哥們說：「看哪，我又做了一個夢；看哪，太陽、月亮和十一顆星都向我下拜。」
GEN|37|10|約瑟 告訴他父親和哥哥們，他父親就責備他說：「你做的這是甚麼夢！難道我和你母親、你的兄弟真的要俯伏在地，來向你下拜嗎？」
GEN|37|11|他的哥哥們都嫉妒他，他父親卻把這事存在心裏。
GEN|37|12|約瑟 的哥哥們到 示劍 去放他們父親的羊。
GEN|37|13|以色列 對 約瑟 說：「你哥哥們不是在 示劍 放羊嗎？來，我派你到他們那裏去。」 約瑟 對他說：「我在這裏。」
GEN|37|14|以色列 對他說：「你去看看你哥哥們是否平安，羊群是否平安，再回來告訴我。」於是他派 約瑟 出 希伯崙谷 ， 約瑟 就往 示劍 去了。
GEN|37|15|有人遇見他，看哪，他在田野走迷了路。那人問他說：「你找甚麼？」
GEN|37|16|他說：「我找我的哥哥們，請告訴我，他們在哪裏放羊。」
GEN|37|17|那人說：「他們已經離開這裏走了，我聽見他們說：『我們往 多坍 去。』」 約瑟 就去追哥哥們，在 多坍 找到了他們。
GEN|37|18|他們遠遠看見他，趁他還沒有走近他們，就圖謀要殺死他。
GEN|37|19|他們彼此說：「看哪！那做夢的來了。
GEN|37|20|現在，來吧！我們把他殺了，丟在一個坑裏，就說有惡獸把他吃了。我們且看他的夢將來怎麼樣。」
GEN|37|21|呂便 聽見了，要救 約瑟 脫離他們的手，說：「我們不可害他的性命」；
GEN|37|22|呂便 又對他們說：「不可流他的血，可以把他丟在這曠野的坑裏，不可下手害他。」 呂便 要救他脫離他們的手，把他還給他父親。
GEN|37|23|約瑟 到了他哥哥們那裏，他們就剝去他的外衣，就是他身上那件長袍。
GEN|37|24|他們抓住他，把他丟在坑裏。那坑是空的，裏頭沒有水。
GEN|37|25|他們坐下吃飯，舉目觀看，看哪，有一群 以實瑪利 人從 基列 來，用駱駝馱著香料、乳香、沒藥，要帶下 埃及 去。
GEN|37|26|猶大 對他的兄弟們說：「我們殺我們的弟弟，遮掩他的血有甚麼好處呢？
GEN|37|27|來，我們把他賣給 以實瑪利 人，不要下手害他，因為他是我們的弟弟，我們的骨肉。」他的兄弟們就聽從了他。
GEN|37|28|那時，有些 米甸 的商人從那裏經過，就把 約瑟 從坑裏拉上來。他們以二十塊銀子把 約瑟 賣給 以實瑪利 人，他們就把 約瑟 帶到 埃及 去了。
GEN|37|29|呂便 回到坑旁，看哪， 約瑟 不在坑裏，就撕裂自己的衣服，
GEN|37|30|回到他兄弟們那裏，說：「孩子不在了。我往哪裏去才好呢？」
GEN|37|31|於是，他們宰了一隻公山羊，拿了 約瑟 的那件外衣染上了血，
GEN|37|32|派人把長袍送到他們的父親那裏，說：「我們發現這個， 請認一認，是不是你兒子的外衣？」
GEN|37|33|他認出來，就說：「這是我兒子的外衣，惡獸把他吃了， 約瑟 一定被撕碎了！」
GEN|37|34|雅各 就撕裂衣服，腰間圍上麻布，為他兒子哀傷了多日。
GEN|37|35|他的兒女都起來安慰他，他卻不肯受安慰，說：「我必哀傷著下陰間，到我兒子那裏。」 約瑟 的父親就為他哀哭。
GEN|37|36|米甸 人把 約瑟 賣到 埃及 ，給法老的官員，就是護衛長 波提乏 。
GEN|38|1|那時， 猶大 離開他兄弟們下去，到一個名叫 希拉 的 亞杜蘭 人的家附近支搭帳棚。
GEN|38|2|猶大 在那裏看見一個名叫 拔．書亞 的 迦南 女子，就娶她為妻，與她同房，
GEN|38|3|她就懷孕生了兒子， 猶大 給他起名叫 珥 。
GEN|38|4|她又懷孕生了兒子，給他起名叫 俄南 。
GEN|38|5|她又再生了兒子，給他起名叫 示拉 。她生 示拉 的時候， 猶大 正在 基悉 。
GEN|38|6|猶大 為長子 珥 娶妻，名叫 她瑪 。
GEN|38|7|猶大 的長子 珥 在耶和華眼中看為惡，耶和華就殺死了他。
GEN|38|8|猶大 對 俄南 說：「你當與你哥哥的妻子同房，向她盡你的本分，為你哥哥生子立後。」
GEN|38|9|俄南 知道如果與嫂嫂同房，所生的孩子不屬於自己，就洩在地上，不為哥哥生子立後。
GEN|38|10|俄南 所做的在耶和華眼中看為惡，耶和華也殺死了他。
GEN|38|11|猶大 對他媳婦 她瑪 說：「你去住在你父親家裏守寡，等我兒子 示拉 長大。」因為他說：「恐怕 示拉 也像兩個哥哥一樣死去。」 她瑪 就去，住在她父親家裏。
GEN|38|12|過了一段很長的日子， 猶大 的妻子， 書亞 的女兒死了。 猶大 受到了安慰，就和他朋友 亞杜蘭 人 希拉 上 亭拿 去，到他的剪羊毛的人那裏。
GEN|38|13|有人告訴 她瑪 說：「看哪，你的公公上 亭拿 剪羊毛去了。」
GEN|38|14|她瑪 見 示拉 已經長大，卻還沒有娶她為妻，就脫去她寡婦的衣裳，用面紗蒙著，蓋住自己，坐在往 亭拿 的路上， 伊拿印 城門口。
GEN|38|15|猶大 看見她，以為是妓女，因為她蒙著臉。
GEN|38|16|猶大 就轉到路邊她那裏，說：「來吧！讓我與你同寢。」他並不知道她就是他的媳婦。 她瑪 說：「你要與我同寢，把甚麼給我呢？」
GEN|38|17|猶大 說：「我從羊群裏取一隻小山羊，派人送來給你。」 她瑪 說：「在未送之前，你能給我一個信物嗎？」
GEN|38|18|他說：「我給你甚麼信物呢？」 她瑪 說：「你的印、你的帶子 和你手裏的杖。」於是 猶大 給了她，與她同寢，她就從 猶大 懷了孕。
GEN|38|19|她瑪 起來走了，除去面紗，照常穿上寡婦的衣裳。
GEN|38|20|猶大 託他朋友 亞杜蘭 人送一隻小山羊去，要從那女人手裏取回信物，卻找不到她。
GEN|38|21|他問那地方的人說：「 伊拿印 路旁的神廟娼妓在哪裏？」他們說：「這裏沒有神廟娼妓。」
GEN|38|22|他回到 猶大 那裏說：「我找不到她，並且那地方的人說：『這裏沒有神廟娼妓。』」
GEN|38|23|猶大 說：「讓她拿去吧，免得我們被人譏笑。看哪，我把這小山羊送去了，可是你找不到她。」
GEN|38|24|大約過了三個月，有人告訴 猶大 說：「你的媳婦 她瑪 行淫，並且，看哪，她因行淫而懷了孕。」 猶大 說：「拉她出來，把她燒了！」
GEN|38|25|她瑪 被拉出來的時候，就派人到她公公那裏，對他說：「這些東西是誰的，我就是從誰懷了孕。」她又說：「請你認一認，這印、這帶子和這杖是誰的？」
GEN|38|26|猶大 承認說：「她比我更有理，因為我沒有把她給我的兒子 示拉 。」 猶大 再也不跟她同寢。
GEN|38|27|她瑪 生產的時候到了，看哪，腹裏懷的是雙胞胎。
GEN|38|28|生產的時候，一個孩子伸出手來；接生婆拿紅線綁在他手上，說：「這是頭生的。」
GEN|38|29|這孩子把手收回去，看哪，他哥哥生出來了；接生婆說：「你竟然為自己衝出一個裂縫！」於是，他的名字叫 法勒斯 。
GEN|38|30|後來，那手上有紅線的兄弟也生出來，他的名字叫 謝拉 。
GEN|39|1|約瑟 被帶下 埃及 去。有一個 埃及 人 波提乏 ，是法老的官員，是護衛長，他從那些帶 約瑟 下來的 以實瑪利 人手中把 約瑟 買了去。
GEN|39|2|約瑟 在他 埃及 主人的家中，耶和華與他同在，他是一個通達的人。
GEN|39|3|他主人見耶和華與他同在，又見耶和華使他手裏所辦的事都順利，
GEN|39|4|約瑟 就在主人眼前蒙恩，伺候他主人，主人派他管理家務，把一切所有的都交在他手裏。
GEN|39|5|自從主人派 約瑟 管理家務和他一切所有的，耶和華就因 約瑟 的緣故賜福給那 埃及 人的家；凡家裏和田間一切所有的，都蒙耶和華賜福。
GEN|39|6|波提乏 把他一切所有的都交在 約瑟 手中，除了自己所吃的食物，其他的事一概不知。 約瑟 英俊健美。
GEN|39|7|這些事以後， 約瑟 主人的妻子以目送情給 約瑟 ，說：「你與我同寢吧！」
GEN|39|8|約瑟 拒絕，對他主人的妻子說：「看哪，一切家務我主人一概不知，他把所有的都交在我手裏。
GEN|39|9|在這家裏沒有人比我更大，除你以外，他也沒有留下一樣不交給我，因為你是他的妻子。我怎能行這麼大的惡，得罪上帝呢？」
GEN|39|10|她天天這樣對 約瑟 說， 約瑟 卻不聽從她，不與她同寢，也不和她在一起。
GEN|39|11|有一天， 約瑟 進屋裏去辦事，家裏沒有一個人在那屋子裏，
GEN|39|12|婦人就拉住他的衣服，說：「你與我同寢吧！」 約瑟 把衣服留在她手裏，逃出外面去了。
GEN|39|13|婦人看見 約瑟 把衣服留在她手裏逃到外面，
GEN|39|14|就叫了家裏的人來，對他們說：「看，他帶了一個 希伯來 人到我們這裏戲弄我們。他到我這裏來，要與我同寢，我就大聲喊叫。
GEN|39|15|他聽見我放聲大喊，就把他的衣服留在我這裏，逃出外面去了。」
GEN|39|16|婦人把 約瑟 的衣服放在身邊，直到他主人回家，
GEN|39|17|就用這樣的話對他說：「你帶到我們這裏來的那 希伯來 僕人進來要調戲我，
GEN|39|18|我放聲大喊，他就把衣服留在我身邊，逃到外面。」
GEN|39|19|主人聽見他妻子對他說的話，說：「你的僕人就是這樣對待我」，就非常生氣。
GEN|39|20|約瑟 的主人把他抓起來，關在監獄裏，就是王的囚犯被關的地方。於是 約瑟 在那裏坐牢。
GEN|39|21|但耶和華與 約瑟 同在，向他施恩，使他在監獄長的眼前蒙恩。
GEN|39|22|監獄長就把監獄裏所有的囚犯都交在 約瑟 手下；在那裏的一切事都由他處理。
GEN|39|23|任何交在 約瑟 手中的事，監獄長一概不察，因為耶和華與 約瑟 同在，耶和華使他所做的都順利。
GEN|40|1|這些事以後， 埃及 王的司酒長和司膳長得罪了他們的主 埃及 王。
GEN|40|2|法老就對司酒長和司膳長兩個官員發怒，
GEN|40|3|把他們關在護衛長府內的監獄裏，就是 約瑟 被囚的地方。
GEN|40|4|護衛長把他們交給 約瑟 ， 約瑟 就伺候他們。他們被關了一段日子。
GEN|40|5|關在監獄裏的這兩個人，就是 埃及 王的司酒長和司膳長，在同一個晚上各自做了一個夢，每個夢都有自己的解釋。
GEN|40|6|到了早晨， 約瑟 來到他們那裏看他們，看哪，他們很憂愁。
GEN|40|7|他就問一同關在他主人府內法老的官員，說：「你們今日為甚麼面帶愁容呢？」
GEN|40|8|他們對他說：「我們各自做了一個夢，卻沒有人能講解。」 約瑟 對他們說：「解夢不是出於上帝嗎？請你們把夢告訴我。」
GEN|40|9|司酒長就把夢告訴 約瑟 ，對他說：「在我的夢中，看哪，有一棵葡萄樹在我面前，
GEN|40|10|樹上有三根枝子。枝子發了芽，開了花，結出串串成熟的葡萄。
GEN|40|11|法老的杯在我手中，我就拿葡萄擠在法老的杯裏，把杯遞到他手中。」
GEN|40|12|約瑟 對他說：「夢的解釋是這樣：三根枝子就是三天；
GEN|40|13|三天之內，法老要讓你抬起頭來，叫你官復原職。你仍要遞杯在法老的手中，像先前作他的司酒長一樣。
GEN|40|14|但你得福的時候，請你記得我，向我施慈愛，在法老面前提起我，救我出這監牢。
GEN|40|15|我實在是從 希伯來 人之地被拐來的，我在這裏也沒有做過甚麼，好叫他們把我關在牢裏。」
GEN|40|16|司膳長見夢解得好，就對 約瑟 說：「在我夢中，看哪，我頭上頂著三個裝餅的籃子；
GEN|40|17|最上面的籃子裏有為法老烤的各樣食物，有飛鳥來吃我頭上籃子裏的食物。」
GEN|40|18|約瑟 說：「夢的解釋是這樣：三個籃子就是三天；
GEN|40|19|三天之內，法老要讓你抬起頭來，身首異處，把你掛在木架上，必有飛鳥來吃你身上的肉。」
GEN|40|20|到了第三天，正是法老的生日，他為眾臣僕擺設宴席，使司酒長和司膳長從眾臣僕中抬起頭來，
GEN|40|21|讓司酒長官復原職，仍舊遞杯在法老手中，
GEN|40|22|卻把司膳長掛起來，正如 約瑟 向他們所講解的。
GEN|40|23|然而，司酒長不記得 約瑟 ，竟忘了他。
GEN|41|1|過了兩年，法老做夢，看哪，自己站在 尼羅河 邊，
GEN|41|2|看哪，有七頭母牛從 尼羅河 裏上來，長相俊美，肌肉肥壯，在蘆葦中吃草。
GEN|41|3|看哪，隨後又有七頭母牛從 尼羅河 裏上來，長相醜陋，肌肉乾瘦，與那七頭母牛一同站在河邊。
GEN|41|4|這長相醜陋，肌肉乾瘦的七頭母牛吃了那長相俊美又肥壯的七頭母牛。法老就醒了。
GEN|41|5|他又睡著，第二次做夢，看哪，一株麥桿長了七個穗子，又肥大又佳美，
GEN|41|6|看哪，隨後又長出七個穗子，又細弱又被東風吹焦了。
GEN|41|7|這細弱的穗子吞了那七個又肥大又飽滿的穗子。法老醒了，看哪，是個夢。
GEN|41|8|到了早晨，法老心裏不安，就派人把 埃及 所有的術士和智慧人都召來。法老把所做的夢告訴他們，但是沒有人能為法老解夢。
GEN|41|9|那時司酒長對法老說：「我今日想起我的罪來。
GEN|41|10|從前法老對臣僕發怒，把我和司膳長關在護衛長府內的監牢裏。
GEN|41|11|我們兩人在同一晚上各做一夢，每個夢都有各自的解釋。
GEN|41|12|同我們在一起有一個 希伯來 的年輕人，是護衛長的僕人。我們告訴他，他就為我們解夢，照著各人的夢講解。
GEN|41|13|後來事情正如他給我們講解的實現了，我官復原職，司膳長被掛起來了。」
GEN|41|14|於是法老派人去召 約瑟 ，他們就急忙把他從牢裏提出來。他就剃頭刮臉，換衣服，進到法老面前。
GEN|41|15|法老對 約瑟 說：「我做了一個夢，沒有人能講解。我聽人說，你聽了夢就能講解。」
GEN|41|16|約瑟 回答法老說：「這不在乎我。上帝必應允法老平安。」
GEN|41|17|法老對 約瑟 說：「在我的夢中，看哪，我站在 尼羅河 邊，
GEN|41|18|看哪，有七頭母牛從 尼羅河 裏上來，肌肉肥壯，外形俊美，在蘆葦中吃草。
GEN|41|19|看哪，隨後又有七頭母牛上來，虛弱，外形很醜陋，肌肉又乾瘦，在 埃及 全地，我沒有見過這樣醜陋的牛。
GEN|41|20|這乾瘦又醜陋的母牛吃了那先前的七頭肥母牛，
GEN|41|21|進了肚子以後卻看不出已經進了肚子，那醜陋的長相仍舊和先前一樣。我就醒了。
GEN|41|22|我又在夢中觀看，看哪，一株麥桿長了七個穗子，又飽滿又佳美，
GEN|41|23|看哪，隨後又長出七個穗子，枯槁，細弱，又被東風吹焦了。
GEN|41|24|這些細弱的穗子吞了那七個佳美的穗子。我告訴術士，卻沒有人能為我講解。」
GEN|41|25|約瑟 對法老說：「法老的夢是同一個。上帝已把要做的事指示法老了。
GEN|41|26|七頭好母牛是七年，七個佳美的穗子也是七年，這是同一個夢。
GEN|41|27|那隨後上來的七頭乾瘦又醜陋的母牛是七年；那七個空心，被東風吹焦的穗子也一樣，都是七個荒年。
GEN|41|28|這就是我對法老所說，上帝已把要做的事顯明給法老了。
GEN|41|29|看哪，必有七個大豐年來到 埃及 全地，
GEN|41|30|隨後又有七個荒年，甚至 埃及 地的人都忘了先前的豐收，這地必被饑荒所滅。
GEN|41|31|因為那後來的饑荒非常嚴重，就不覺得這地先前有豐收。
GEN|41|32|至於法老兩次做夢，是因為上帝已經確定這事，上帝必速速成就。
GEN|41|33|現在，請法老選一個聰明又有智慧的人，委派他治理 埃及 地。
GEN|41|34|請法老這樣做，委派官員治理這地，在七個豐年的期間，徵收 埃及 地出產的五分之一，
GEN|41|35|叫他們聚集未來豐年一切的糧食，積存五穀歸在法老的手下作糧食，儲藏在各城裏。
GEN|41|36|這糧食可以為這地作儲備，為了 埃及 地要來的七個荒年，免得這地被饑荒所滅。」
GEN|41|37|這事在法老和他眾臣僕眼中都覺得好。
GEN|41|38|法老對臣僕說：「像這樣的人，有上帝的靈在他裏面，我們豈能找得著呢？」
GEN|41|39|法老對 約瑟 說：「上帝既指示你這一切事，就沒有人像你這樣聰明又有智慧。
GEN|41|40|你可以治理我的家；我的百姓都必服從你口中的命令。惟獨在寶座上，我比你大。」
GEN|41|41|法老又對 約瑟 說：「看，我委派你治理 埃及 全地。」
GEN|41|42|法老就脫下手上帶印的戒指，戴在 約瑟 的手上，給他穿上細麻衣，把金鏈戴在他的頸項上，
GEN|41|43|又給 約瑟 坐他的副座車，在他前面有人呼叫說：「跪下 。」於是，法老委派他治理 埃及 全地。
GEN|41|44|法老對 約瑟 說：「我是法老，若沒有你的命令， 埃及 全地的人都不可擅自辦事 。」
GEN|41|45|法老給 約瑟 起名叫 撒發那特‧巴內亞 ，又將 安城 的祭司 波提‧非拉 的女兒 亞西納 給他為妻。 約瑟 就出去治理 埃及 地。
GEN|41|46|約瑟 在 埃及 王法老面前侍立的時候年三十歲。 約瑟 從法老面前出去，巡行 埃及 全地。
GEN|41|47|七個豐年之內，地的出產極其豐盛 ，
GEN|41|48|約瑟 聚集 埃及 地七年一切的糧食，把糧食積存在各城裏，就是把各城周圍田地的糧食都積存在該城裏。
GEN|41|49|約瑟 積存的五穀很多，如同海邊的沙，無法計算，數也數不清。
GEN|41|50|荒年未到以前， 安城 的祭司 波提‧非拉 的女兒 亞西納 為 約瑟 生了兩個兒子。
GEN|41|51|約瑟 給長子起名叫 瑪拿西 ，因為他說：「上帝使我忘了一切的困苦和我父的全家。」
GEN|41|52|他給次子起名叫 以法蓮 ，因為他說：「上帝使我在受苦的地方興盛。」
GEN|41|53|埃及 地的七個豐年一過，
GEN|41|54|七個荒年就來了，正如 約瑟 所說的。各地都有饑荒，惟獨 埃及 全地有糧食。
GEN|41|55|等到 埃及 全地也有了饑荒，眾百姓就向法老哀求糧食。法老對所有的 埃及 人說：「你們到 約瑟 那裏去，凡他所說的，你們都要做。」
GEN|41|56|當時饑荒遍滿了全地， 約瑟 就開了各處的糧倉 ，賣糧食給 埃及 人。 埃及 地的饑荒非常嚴重。
GEN|41|57|各地的人都去 埃及 ，到 約瑟 那裏買糧食，因為全地的饑荒非常嚴重。
GEN|42|1|雅各 見 埃及 有糧，就對兒子們說：「你們為甚麼彼此對看呢？」
GEN|42|2|他又說：「看哪，我聽見 埃及 有糧，你們可以下到那裏，從那裏為我們買些糧來，我們就可以存活，不至於死。」
GEN|42|3|於是， 約瑟 的十個哥哥都下去，到 埃及 買糧食。
GEN|42|4|至於 約瑟 的弟弟 便雅憫 ， 雅各 沒有派他和哥哥們同去，因為 雅各 說：「恐怕他遭難。」
GEN|42|5|以色列 的兒子們來了，在前來的人當中，為要買糧食，因為 迦南 地也有饑荒。
GEN|42|6|當時在 埃及 地掌權的人是 約瑟 ，賣糧給各地眾百姓的就是他。 約瑟 的哥哥們來了，臉伏於地，向他下拜。
GEN|42|7|約瑟 看見他哥哥們，就認出他們，卻對他們裝作陌生人，向他們說嚴厲的話，對他們說：「你們從哪裏來？」他們說：「我們從 迦南 地來買糧。」
GEN|42|8|約瑟 認得他哥哥們，他們卻不認得他。
GEN|42|9|約瑟 想起從前所做的那兩個夢，就對他們說：「你們是奸細，你們來是要窺探這地的虛實。」
GEN|42|10|他們對他說：「我主啊，不是的，僕人們是來買糧的。
GEN|42|11|我們都是同一個人的兒子，我們是誠實的人。僕人們並不是奸細。」
GEN|42|12|約瑟 對他們說：「不，你們一定是窺探這地的虛實來的。」
GEN|42|13|他們說：「僕人們本是兄弟十二人，我們都是 迦南 地同一個人的兒子。看哪，最小的今日在我們父親那裏，有一個不在了。」
GEN|42|14|約瑟 對他們說：「我剛才對你們說過了，你們是奸細！
GEN|42|15|我指著法老的性命起誓，若是你們最小的弟弟不到這裏來，你們就不可以離開這裏；這樣你們就可以證實自己了。
GEN|42|16|要派你們當中的一個人去，把你們的弟弟帶來。至於你們，都要關在這裏，好證實你們的話是不是真的。若不是，我指著法老的性命起誓，你們一定是奸細。」
GEN|42|17|於是 約瑟 把他們一起都關在監裏三天。
GEN|42|18|第三天， 約瑟 對他們說：「我是敬畏上帝的，你們這麼做就可以活。
GEN|42|19|如果你們是誠實的人，留你們兄弟中的一個關在監牢裏，你們帶糧食回去，救你們家的饑荒，
GEN|42|20|再把你們最小的弟弟帶到我這裏來。如此，你們的話就是真的了，你們也不至於死。」他們就照樣做了。
GEN|42|21|他們彼此說：「我們在弟弟身上實在犯了罪。他哀求我們的時候，我們看見他的痛苦，卻不肯聽，所以這場苦難臨到我們。」
GEN|42|22|呂便 回答他們說：「我不是對你們說過，不可傷害那孩子嗎？只是你們不肯聽，看哪，他的血在追討了。」
GEN|42|23|他們不知道 約瑟 在聽，因為在他們之間有傳譯官。
GEN|42|24|約瑟 轉身離開他們，哭了一場，又回來對他們說話，就從他們中間抓了 西緬 ，在他們眼前捆綁他。
GEN|42|25|約瑟 吩咐人把他們的器皿裝滿糧食，把各人的銀子退還在各人的袋裏，又給他們路上需用的食物。人就為他們這樣做了。
GEN|42|26|他們把糧食馱在驢上，離開那裏去了。
GEN|42|27|到了住宿的地方，有一個人打開袋子，要拿飼料餵驢，就看見自己的銀子，看哪，仍在袋口上。
GEN|42|28|他對兄弟們說：「我的銀子退回來了，看哪，還在我袋子裏！」他們戰戰兢兢，心都快跳出來了，彼此說：「上帝向我們做的是甚麼呢？」
GEN|42|29|他們來到 迦南 地他們的父親 雅各 那裏，把所遭遇的事都告訴他，說：
GEN|42|30|「那地的主對我們說嚴厲的話，把我們當作窺探那地的奸細。
GEN|42|31|我們對他說：『我們是誠實的人，並不是奸細。
GEN|42|32|我們本是兄弟十二人，都是同一個父親的兒子，有一個不在了，最小的今日和我們父親在 迦南 地。』
GEN|42|33|那地的主對我們說：『只有這樣我才知道你們是誠實的人：留你們兄弟中的一個在我這裏，你們帶糧食回去，救你們家的饑荒，
GEN|42|34|再把你們最小的弟弟帶到我這裏來，我就知道你們不是奸細，是誠實的人。然後，我就把你們的兄弟交還你們，你們也可以在此地做買賣。』」
GEN|42|35|後來他們倒空袋子，看哪，各人的銀囊都在袋子裏。他們和父親看見銀囊就都害怕。
GEN|42|36|他們的父親 雅各 對他們說：「你們害我喪失了我的兒子： 約瑟 不在了， 西緬 也不在了，你們還要帶走 便雅憫 ！這些事都臨到我身上了。」
GEN|42|37|呂便 對他父親說：「我若不帶他回來給你，你可以殺我的兩個兒子。只管把他交在我手裏，我必帶他回來給你。」
GEN|42|38|雅各 說：「我的兒子不可與你們一同下去。他哥哥死了，只剩下他。他若在你們行走的路上遭難，你們就害我白髮蒼蒼、悲悲慘慘下陰間去了。」
GEN|43|1|那地的饑荒非常嚴重。
GEN|43|2|他們從 埃及 帶來的糧食吃完了，父親對他們說：「你們再去給我們買些糧來。」
GEN|43|3|猶大 對他說：「那人嚴厲地警告我們說：『你們的弟弟若不和你們同來，你們就不要來見我的面。』
GEN|43|4|你若派我們的弟弟跟我們同去，我們就下去給你買糧；
GEN|43|5|你若不派他去，我們就不下去，因為那人對我們說：『你們的弟弟若不和你們同來，你們就不要來見我的面。』」
GEN|43|6|以色列 說：「你們為甚麼這樣害我，告訴那人你們還有弟弟呢？」
GEN|43|7|他們說：「那人詳細問到我們和我們的家人，說：『你們的父親還在嗎？你們還有兄弟嗎？』我們就按著他的這些話告訴他，我們怎麼知道他會說：『把你們的弟弟帶下來』呢？」
GEN|43|8|猶大 又對他父親 以色列 說：「請派這年輕人和我同去，我們就動身前去，好叫我們和你，以及我們的孩子都得存活，不至於死。
GEN|43|9|我為他擔保，你可以從我手中要人，我若不帶他回來交在你面前，我就對你永遠擔當這罪。
GEN|43|10|我們若沒有耽擱，現在第二趟都回來了。」
GEN|43|11|父親 以色列 對他們說：「如果必須如此，你們要這樣做：把本地土產中最好的乳香、蜂蜜、香料、沒藥、堅果、杏仁各取一點，放在器皿裏，帶下去送給那人作禮物。
GEN|43|12|手裏要帶雙倍的銀子，把退還在你們袋口的銀子親手帶回去；或許那是個失誤。
GEN|43|13|帶著你們的弟弟，動身再去見那人。
GEN|43|14|願全能的上帝使你們在那人面前蒙憐憫，放你們另一個兄弟和 便雅憫 回來。我若要失喪兒子，就喪了吧！」
GEN|43|15|於是，他們拿著那些禮物，手裏也帶雙倍的銀子，並且帶著 便雅憫 ，動身下到 埃及 ，站在 約瑟 面前。
GEN|43|16|約瑟 見 便雅憫 和他們同來，就對管家說：「把這些人領到屋裏。要宰殺牲畜，預備宴席，因為中午這些人要跟我吃飯。」
GEN|43|17|那人就照 約瑟 所說的去做，領他們進 約瑟 的屋裏。
GEN|43|18|這些人因為被領到 約瑟 的屋裏，就害怕，說：「領我們到這裏來，必是因為當初退還在我們袋裏的銀子，要設計害我們，抓我們去當奴隸，搶奪我們的驢。」
GEN|43|19|他們就挨近 約瑟 的管家，在屋子門口和他說話，
GEN|43|20|說：「我主啊，求求你，我們當初下來，真的是要買糧食。
GEN|43|21|後來到了住宿的地方，我們打開袋子，看哪，各人的銀子還在自己的袋口上，銀子的分量一點不少。現在我們親手把它帶回來，
GEN|43|22|我們手裏又帶了另外的銀子來買糧食。我們不知道是誰把銀子放在我們袋裏的。」
GEN|43|23|他說：「你們平安！不要害怕，是你們的上帝和你們父親的上帝把財寶放在你們的袋裏。你們的銀子，我已經收了。」他就把 西緬 帶出來，交給他們。
GEN|43|24|那人領這些人進 約瑟 的屋裏，給他們水洗腳，又給他們飼料餵驢。
GEN|43|25|他們預備好禮物，等候 約瑟 中午來，因為他們聽說他們要在那裏吃飯。
GEN|43|26|約瑟 來到家裏，他們就把手中的禮物拿進屋裏給他，俯伏在地，向他下拜。
GEN|43|27|約瑟 問他們安，又說：「你們的父親，就是你們所說的那位老人家平安嗎？他還在嗎？」
GEN|43|28|他們說：「你僕人，我們的父親平安，他還在。」於是他們低頭下拜。
GEN|43|29|約瑟 舉目看見他同母的弟弟 便雅憫 ，就說：「你們向我所說那最小的弟弟就是這位嗎？」又說：「我兒啊，願上帝賜恩給你！」
GEN|43|30|約瑟 愛弟之情激動，就急忙找個地方去哭。他進入自己的房間，哭了一場。
GEN|43|31|他洗了臉出來，勉強忍住，就說：「開飯吧！」
GEN|43|32|他們為 約瑟 單獨擺了一席，為那些人又擺了一席，也為和 約瑟 同吃飯的 埃及 人另擺了一席，因為 埃及 人不和 希伯來 人一同吃飯；那是 埃及 人所厭惡的。
GEN|43|33|兄弟們被安排在 約瑟 面前坐席，都按著長幼的次序，這些人彼此感到詫異。
GEN|43|34|約瑟 把他面前的食物分給他們，但 便雅憫 所得的比別人多五倍。他們就喝酒，和 約瑟 一同暢飲。
GEN|44|1|約瑟 吩咐管家說：「按照他們的驢子所能馱的，把這些人的袋子裝滿糧食，再把各人的銀子放在各人的袋口上，
GEN|44|2|我的杯，就是那個銀杯，要和買糧的銀子一同放在最年輕的那個人的袋口上。」管家就照 約瑟 所說的話去做了。
GEN|44|3|天一亮，這些人和他們的驢子就被送走了。
GEN|44|4|他們出城走了不遠， 約瑟 對管家說：「起來，去追那些人，追上了就對他們說：『你們為甚麼以惡報善呢？
GEN|44|5|這不是我主人用來飲酒，確實用它來占卜的嗎？你們這麼做是不對的！』」
GEN|44|6|管家追上他們，把這些話對他們說了。
GEN|44|7|他們對他說：「我主為甚麼說這樣的話呢？你僕人們絕不會做這樣的事。
GEN|44|8|看哪，我們從前在袋口上發現的銀子，尚且從 迦南 地帶來還你，我們又怎麼會從你主人家裏偷竊金銀呢？
GEN|44|9|你僕人中無論在誰那裏找到杯子，就叫他死，我們也要作我主的奴隸。」
GEN|44|10|管家說：「現在就照你們的話做吧！在誰那裏找到杯子，誰就作我的奴隸，其餘的人都沒有罪。」
GEN|44|11|於是他們各人急忙把袋子卸在地上，各人打開自己的袋子。
GEN|44|12|管家就搜查，從年長的開始到年幼的為止，那杯竟在 便雅憫 的袋子裏找到了。
GEN|44|13|他們就撕裂衣服，各人把馱子抬在驢上，回城去了。
GEN|44|14|猶大 和他兄弟們來到 約瑟 的屋裏， 約瑟 還在那裏，他們就在他面前俯伏於地。
GEN|44|15|約瑟 對他們說：「你們做的是甚麼事呢？你們豈不知像我這樣的人必懂得占卜嗎？」
GEN|44|16|猶大 說：「我們對我主能說甚麼呢？還有甚麼話可說呢？我們還能為自己表白嗎？上帝已經查出你僕人的罪孽了。看哪，我們與那在他手中找到杯子的人都是我主的奴隸。」
GEN|44|17|約瑟 說：「我絕不能做這樣的事！誰的手中找到杯子，誰就作我的奴隸。至於你們，可以平平安安上到你們父親那裏去。」
GEN|44|18|猶大 挨近他，說：「我主啊，求求你，讓僕人說一句話給我主聽，不要向僕人發烈怒，因為你如同法老一樣。
GEN|44|19|我主曾問僕人們說：『你們有父親、兄弟沒有？』
GEN|44|20|我們對我主說：『我們有父親，他已經年老，還有他老年所生的一個小兒子。他哥哥死了，他的母親只剩下他一個孩子，父親也疼愛他。』
GEN|44|21|你對僕人說：『把他帶下到我這裏來，讓我親眼看看他。』
GEN|44|22|我們對我主說：『這年輕人不能離開他父親，若是離開，父親就會死。』
GEN|44|23|你對僕人說：『你們最小的弟弟若不和你們一同下來，你們就不要來見我的面。』
GEN|44|24|我們上到你僕人，我們父親那裏，就把我主的話告訴了他。
GEN|44|25|後來，我們的父親說：『你們再去給我買些糧來。』
GEN|44|26|我們說：『我們不能下去。最小的弟弟若和我們同去，我們就可以下去。因為，最小的弟弟若不和我們同去，我們必不能見那人的面。』
GEN|44|27|你僕人，我父親對我們說：『你們知道我的妻子給我生了兩個兒子。
GEN|44|28|一個離開我走了，我說他必是被野獸撕碎了，直到如今我再沒有見過他；
GEN|44|29|現在你們又要把這個從我面前帶走。倘若他遭難，那麼你們就害我白髮蒼蒼、悲悲慘慘下陰間去了。』
GEN|44|30|如今我回到你僕人，我父親那裏，若沒有這年輕人和我們同去，我父親的命是與這年輕人的命相連的，
GEN|44|31|當我們的父親看見沒有了這年輕人，他就會死。這樣，我們就害你僕人，我們的父親白髮蒼蒼、悲悲慘慘下陰間去了。
GEN|44|32|僕人曾向我父親為這年輕人擔保，說：『我若不帶他回來交給父親，我就在父親面前永遠擔當這罪。』
GEN|44|33|現在，求你把僕人留下，代替這年輕人作我主的奴隸，讓這年輕人和他哥哥們一同上去。
GEN|44|34|若這年輕人不和我一起，我怎能上到我父親那裏呢？恐怕我要看到災禍臨到我父親了。」
GEN|45|1|約瑟 在所有侍立在他旁邊的人面前情不自禁，就喊叫說：「每一個人都離開我，出去吧！」 約瑟 和兄弟相認的時候沒有一人站在他那裏。
GEN|45|2|他放聲大哭， 埃及 人聽見了，法老家中的人也聽見了。
GEN|45|3|約瑟 對他兄弟們說：「我就是 約瑟 。我的父親還在嗎？」他兄弟們不敢回答他，因為他們在他面前都很驚惶。
GEN|45|4|約瑟 又對他兄弟們說：「靠近我一點。」他們就近前來。他說：「我是被你們賣到 埃及 的兄弟 約瑟 。
GEN|45|5|現在，不要因為把我賣到這裏而憂傷，對自己生氣，因為上帝差我在你們以先來，為要保全性命。
GEN|45|6|現在這地的饑荒已經二年了，還有五年不能耕種，沒有收成。
GEN|45|7|上帝差我在你們以先來，為要給你們在世上存留餘種，大施拯救，保全你們的性命。
GEN|45|8|這樣看來，差我到這裏來的不是你們，而是上帝。他又使我如同法老之父，作他全家之主，和 埃及 全地掌權的人。
GEN|45|9|你們要趕緊上到我父親那裏，對他說：『你兒子 約瑟 這樣說：上帝已立我作全 埃及 之主，請你下到我這裏來，不要耽擱。
GEN|45|10|你和你的兒子孫子，羊群牛群，以及一切所有的，都可以住在 歌珊 地，與我相近。
GEN|45|11|我要在那裏奉養你，因為還有五年的饑荒，免得你和你的家屬，以及一切所有的，都陷入窮困中。』
GEN|45|12|看哪，你們的眼睛和我弟弟 便雅憫 的眼睛都看見，是我親口對你們說話。
GEN|45|13|你們要把我在 埃及 一切的尊榮和你們所有看見的事情都告訴我父親，也要趕緊請我父親下到這裏來。」
GEN|45|14|於是 約瑟 伏在他弟弟 便雅憫 的頸項上哭， 便雅憫 也在他的頸項上哭。
GEN|45|15|他又親眾兄弟，伏著他們哭。過後，他的兄弟就和他說話。
GEN|45|16|這消息傳到法老的宮裏，說：「 約瑟 的兄弟們來了。」法老和他的臣僕眼中都看為好。
GEN|45|17|法老對 約瑟 說：「你要吩咐你的兄弟們說：『你們要這樣做：把馱子抬在牲口上，動身到 迦南 地去，
GEN|45|18|請你們的父親和你們的家屬都到我這裏來，我要把 埃及 地的美物賜給你們，你們也要吃這地肥美的出產。』
GEN|45|19|你要吩咐他們：『要這樣做：從 埃及 地帶著車輛去，把你們的孩子和妻子，以及你們的父親都接來。
GEN|45|20|你們的眼不要顧惜你們的家具，因為 埃及 全地的美物都是你們的。』」
GEN|45|21|以色列 的兒子們就照樣做了。 約瑟 遵照法老的吩咐，給他們車輛和路上需用的食物。
GEN|45|22|他又給所有哥哥每人一套衣服， 卻給 便雅憫 三百銀子，五套衣服。
GEN|45|23|他也送給父親十匹公驢，馱著 埃及 的美物，以及十匹母驢，馱著給他父親在路上需用的穀物、餅和糧食。
GEN|45|24|於是 約瑟 送他的兄弟們回去，對他們說：「你們不要在路上爭吵。」
GEN|45|25|他們從 埃及 上去，來到 迦南 地他們的父親 雅各 那裏，
GEN|45|26|告訴他說：「 約瑟 還活著，並且作了 埃及 全地掌權的人。」 雅各 心裏冰涼，因為不信他們。
GEN|45|27|他們就把 約瑟 對他們所說一切的話都告訴了他。他看見 約瑟 派來接他的車輛，他們父親 雅各 的靈就甦醒了。
GEN|45|28|以色列 說：「夠了！我的兒子 約瑟 還活著，我要趁我未死之前去見他。」
GEN|46|1|以色列 帶著一切所有的，起程到 別是巴 去，獻祭給他父親 以撒 的上帝。
GEN|46|2|夜間，上帝在異象中對 以色列 說：「 雅各 ！ 雅各 ！」他說：「我在這裏。」
GEN|46|3|上帝說：「我是上帝，你父親的上帝。不要害怕下 埃及 去，因為我必使你在那裏成為大國。
GEN|46|4|我要和你同下 埃及 去，也必定帶你上來； 約瑟 要親手合上你的眼睛。」
GEN|46|5|雅各 就從 別是巴 起行。 以色列 的兒子讓他們的父親 雅各 和他們的孩子、妻子都坐在法老為 雅各 派來的車上。
GEN|46|6|他們也帶著 迦南 地所得的牲畜和財物來到 埃及 。 雅各 和他所有的子孫都一同來了。
GEN|46|7|他把他的兒子、孫子、女兒、孫女，他所有的子孫一同帶到 埃及 。
GEN|46|8|這些是來到 埃及 的 以色列 人， 雅各 和他子孫的名字： 雅各 的長子是 呂便 。
GEN|46|9|呂便 的兒子是 哈諾 、 法路 、 希斯倫 、 迦米 。
GEN|46|10|西緬 的兒子是 耶母利 、 雅憫 、 阿轄 、 雅斤 、 瑣轄 ，還有 迦南 女子生的兒子 掃羅 。
GEN|46|11|利未 的兒子是 革順 、 哥轄 、 米拉利 。
GEN|46|12|猶大 的兒子是 珥 、 俄南 、 示拉 、 法勒斯 、 謝拉 ； 珥 與 俄南 死在 迦南 地。 法勒斯 的兒子是 希斯崙 、 哈母勒 。
GEN|46|13|以薩迦 的兒子是 陀拉 、 普瓦 、 約伯 、 伸崙 。
GEN|46|14|西布倫 的兒子是 西烈 、 以倫 、 雅利 。
GEN|46|15|這是 利亞 在 巴旦‧亞蘭 為 雅各 所生的兒孫，還有女兒 底拿 ，兒孫共三十三人。
GEN|46|16|迦得 的兒子是 洗非芸 、 哈基 、 書尼 、 以斯本 、 以利 、 亞羅底 、 亞列利 。
GEN|46|17|亞設 的兒子是 音拿 、 亦施瓦 、 亦施韋 、 比利亞 ，還有他們的妹妹 西拉 。 比利亞 的兒子是 希別 、 瑪結 。
GEN|46|18|這是 拉班 給他女兒 利亞 的婢女 悉帕 的兒孫，她為 雅各 所生的共有十六人。
GEN|46|19|雅各 之妻 拉結 的兒子是 約瑟 和 便雅憫 。
GEN|46|20|約瑟 在 埃及 地生了 瑪拿西 和 以法蓮 ，是 安城 的祭司 波提非拉 的女兒 亞西納 為 約瑟 生的。
GEN|46|21|便雅憫 的兒子是 比拉 、 比結 、 亞實別 、 基拉 、 乃幔 、 以希 、 羅實 、 母平 、 戶平 、 亞勒 。
GEN|46|22|這是 拉結 為 雅各 所生的兒孫，共有十四人。
GEN|46|23|但 的兒子是 戶伸 。
GEN|46|24|拿弗他利 的兒子是 雅薛 、 沽尼 、 耶色 、 示冷 。
GEN|46|25|這是 拉班 給他女兒 拉結 的婢女 辟拉 的兒孫，她為 雅各 所生的共有七人。
GEN|46|26|那與 雅各 同到 埃及 的，除了他媳婦之外，凡從他生的共有六十六人。
GEN|46|27|還有 約瑟 在 埃及 所生的兩個兒子。到 埃及 的 雅各 全家共有七十人。
GEN|46|28|雅各 派 猶大 先到 約瑟 那裏，請他先指示到 歌珊 去的路；於是他們來到了 歌珊 地。
GEN|46|29|約瑟 備好座車，上 歌珊 去迎接他的父親 以色列 。他見到父親，就伏在父親的頸項上，在父親的頸項上哭了許久。
GEN|46|30|以色列 對 約瑟 說：「我見了你的面，知道你還活著，現在我可以死了。」
GEN|46|31|約瑟 對他兄弟和他父親的全家說：「我要上去告訴法老，對他說：『我在 迦南 地的兄弟和我父親的全家，都到我這裏來了。
GEN|46|32|他們是牧羊人，是牧放牲畜的人；他們把羊群牛群和一切所有的都帶來了。』
GEN|46|33|等到法老召見你們，說：『你們是做甚麼的？』
GEN|46|34|你們就說：『你的僕人，從幼年直到現在，都是牧放牲畜的人，我們和我們的祖宗都是這樣。』如此，你們就可以住在 歌珊 地，因為凡牧羊的都被 埃及 人厭惡。」
GEN|47|1|約瑟 進去告訴法老說：「我的父親和我的兄弟帶著羊群牛群，以及他們一切所有的，從 迦南 地來了。看哪，他們正在 歌珊 地。」
GEN|47|2|約瑟 從他所有兄弟中挑選五個人，引他們到法老面前。
GEN|47|3|法老對 約瑟 的兄弟說：「你們是做甚麼的？」他們對法老說：「你僕人是牧羊的，我們和我們的祖宗都是這樣。」
GEN|47|4|他們又對法老說：「 迦南 地的饑荒非常嚴重，僕人的羊群沒有牧草，所以我們來到這地寄居。現在求你准許僕人住在 歌珊 地。」
GEN|47|5|法老對 約瑟 說：「你的父親和你的兄弟到你這裏來了，
GEN|47|6|埃及 地都在你面前，只管讓你父親和你兄弟住在最好的地，他們可以住在 歌珊 地。你若知道他們中間有能幹的人，就派他們看管我的牲畜。」
GEN|47|7|約瑟 帶他父親 雅各 來，站在法老面前， 雅各 就為法老祝福。
GEN|47|8|法老對 雅各 說：「你平生的年日是多少呢？」
GEN|47|9|雅各 對法老說：「我在世寄居的年日是一百三十年，我一生的歲月又短又苦，比不上我祖先在世寄居的年日。」
GEN|47|10|雅各 又為法老祝福，就從法老面前退出去了。
GEN|47|11|約瑟 安頓他的父親和兄弟，遵照法老的命令，把 埃及 境內最好的地，就是 蘭塞 地，給他們作為產業。
GEN|47|12|約瑟 用糧食供給他父親和兄弟們，以及他父親全家的人，照扶養親屬的人口供給。
GEN|47|13|饑荒非常嚴重，全地都絕了糧， 埃及 地和 迦南 地都因饑荒耗損了。
GEN|47|14|約瑟 收集了 埃及 地和 迦南 地所有的銀子，就是眾人買糧的銀子， 約瑟 就把那些銀子都帶到法老的宮裏。
GEN|47|15|埃及 地和 迦南 地的銀子都花光了， 埃及 眾人到 約瑟 那裏，說：「我們的銀子都用完了，求你給我們糧食吧！我們為甚麼要死在你面前呢？」
GEN|47|16|約瑟 說：「銀子若是用完了，可以把你們的牲畜賣給我，我就以你們的牲畜換糧食給你們。」
GEN|47|17|於是他們把牲畜帶到 約瑟 那裏， 約瑟 就拿糧食換了他們的馬、羊、牛、驢；那一年他因換他們一切的牲畜，用糧食養活他們。
GEN|47|18|那一年過去，第二年他們又來到 約瑟 那裏，對他說：「不瞞我主，我們的銀子都花光了，牲畜也都歸於我主了。我們在我主面前，除了自己的身體和土地以外，一無所剩。
GEN|47|19|你為甚麼要眼看著我們人死地荒呢？求你用糧食買我們和我們的地，我們和我們的地就要為法老效力。求你給我們種子，使我們可以存活，不致死亡，土地也不致荒蕪。」
GEN|47|20|於是， 約瑟 為法老買了 埃及 所有的土地， 埃及 人因饑荒所迫，都賣了自己的田地；那些地都歸給法老了。
GEN|47|21|至於百姓，從 埃及 邊界的一端到另一端， 約瑟 使他們作奴隸。
GEN|47|22|只有祭司的土地， 約瑟 沒有買，因為祭司從法老領取薪俸，靠法老的薪俸過活，所以沒有賣自己的土地。
GEN|47|23|約瑟 對百姓說：「看哪，我今日為法老買了你們和你們的土地。看，這些種子是給你們的，你們可以耕種土地。
GEN|47|24|將來收割的時候，你們要把五分之一納給法老，另外四分可以給你們作田地的種子，作你們和你們全家大小的食物。」
GEN|47|25|他們說：「你救了我們的性命，願我們在我主眼前蒙恩，我們情願作法老的奴隸。」
GEN|47|26|於是 約瑟 為 埃及 的土地立下定例，直到今日，就是收成的五分之一要歸法老。惟獨祭司的土地例外，不歸於法老。
GEN|47|27|以色列 人住在 埃及 境內的 歌珊 地。他們在那裏得了產業，並且生養眾多。
GEN|47|28|雅各 住在 埃及 地十七年。 雅各 一生的年日是一百四十七年。
GEN|47|29|以色列 的死期快到了，就叫了他兒子 約瑟 來，對他說：「我若在你眼前蒙恩，把你的手放在我大腿底下，以慈愛和誠實向我承諾，必不將我葬在 埃及 。
GEN|47|30|我與我祖先同睡的時候，你要將我帶出 埃及 ，把我葬在他們所葬的地方。」 約瑟 說：「我必遵照你的吩咐去做。」
GEN|47|31|雅各 說：「你向我起誓吧！」 約瑟 就向他起了誓。於是 以色列 在床頭 敬拜。
GEN|48|1|這些事以後，有人告訴 約瑟 說：「看哪，你的父親病了。」他就帶著兩個兒子 瑪拿西 和 以法蓮 同去。
GEN|48|2|有人告訴 雅各 說：「看哪，你的兒子 約瑟 到你這裏來了。」 以色列 就勉強在床上坐起來。
GEN|48|3|雅各 對 約瑟 說：「全能的上帝曾在 迦南 地的 路斯 向我顯現，賜福給我，
GEN|48|4|對我說：『看哪，我必使你生養眾多，成為許多民族，又要將這地賜給你的後裔，永遠為業。』
GEN|48|5|我未到 埃及 你那裏之前，你在 埃及 地所生的 以法蓮 和 瑪拿西 這兩個兒子，現在他們是我的，正如 呂便 和 西緬 是我的一樣。
GEN|48|6|你在他們以後所生的後裔就是你的，這些後裔可以在自己兄弟的名下得產業。
GEN|48|7|至於我，我從 巴旦 回來的時候， 拉結 在我身旁死了，就是在往 迦南 地的路上，離 以法他 還有一段路程。我就把她葬在往 以法他 的路旁； 以法他 就是 伯利恆 。」
GEN|48|8|以色列 看見 約瑟 的兒子，就說：「這些是誰？」
GEN|48|9|約瑟 對他父親說：「這是上帝在這裏賜給我的兒子。」 以色列 說：「領他們到我跟前，我要為他們祝福。」
GEN|48|10|以色列 年紀老邁，眼睛昏花，不能看見。 約瑟 領他們到他跟前，他就和他們親吻，抱著他們。
GEN|48|11|以色列 對 約瑟 說：「我沒有想到能夠見你的面。看哪，上帝還讓我看見你的兒子。」
GEN|48|12|約瑟 把他們從 以色列 兩膝中間領出來，自己臉伏於地下拜。
GEN|48|13|然後， 約瑟 牽著他們兩個，帶到父親跟前，右手牽 以法蓮 到 以色列 的左邊，左手牽 瑪拿西 到 以色列 的右邊。
GEN|48|14|以色列 卻伸出右手來，按在次子 以法蓮 的頭上，又交叉伸出左手來，按在長子 瑪拿西 的頭上。
GEN|48|15|他就為 約瑟 祝福說： 「願我祖父 亞伯拉罕 和我父親 以撒 所事奉的上帝， 就是一生牧養我直到今日的上帝，
GEN|48|16|救贖我脫離一切患難的那位使者，賜福給這兩個孩子。 願我的名，我祖父 亞伯拉罕 和我父親 以撒 的名藉著他們得以流傳。 又願他們在全地上多多繁衍。」
GEN|48|17|約瑟 見父親把右手按在 以法蓮 的頭上，他看為不好，就提起他父親的手，要從 以法蓮 的頭上移到 瑪拿西 的頭上。
GEN|48|18|約瑟 對父親說：「我父，不是這樣。這個才是長子，請你把右手按在他頭上。」
GEN|48|19|他父親卻不肯，說：「我知道，我兒，我知道。他也要成為一族，也要強大。可是他的弟弟將來比他還要強大；他弟弟的後裔要成為許多國家。」
GEN|48|20|以色列 就在當日為他們祝福，說：「 以色列 人要指著你們祝福，說：『願上帝使你如 以法蓮 、 瑪拿西 一樣。』」於是他立 以法蓮 在 瑪拿西 之上。
GEN|48|21|以色列 又對 約瑟 說：「看哪，我快要死了，但上帝必與你們同在，領你們回到你們祖先之地。
GEN|48|22|從前我用刀用弓從 亞摩利 人手下奪取的那一份，我要把它賜給你，使你比你的兄弟多得一份 。」
GEN|49|1|雅各 叫了他的兒子來，說：「你們都來聚集，讓我把你們日後要遇到的事告訴你們。
GEN|49|2|雅各 的兒子們，你們要聚集，要聆聽， 聽你們父親 以色列 的話。
GEN|49|3|呂便 啊，你是我的長子，我的力量， 我壯年頭生之子， 極有尊榮，權力超群。
GEN|49|4|你卻放縱如水，必不得居首位； 因為你上了你父親的床， 你 上了我的榻，污辱了它！
GEN|49|5|西緬 和 利未 是兄弟； 他們的刀劍是殘暴的兵器。
GEN|49|6|願我的心不與他們同謀， 願我的靈 不與他們合夥； 因為他們在烈怒中殺人， 任意割斷牛腿的筋。
GEN|49|7|他們火爆的烈怒可詛， 他們兇殘的憤恨可咒！ 我要把他們分散在 雅各 中， 使他們散居在 以色列 。
GEN|49|8|猶大 啊，你的兄弟必讚美你， 你的手必掐住仇敵的頸項， 你父親的兒子要向你下拜。
GEN|49|9|猶大 是隻小獅子； 我兒啊，你捕獲了獵物就上去。 他蹲伏，他躺臥，如公獅， 又如母獅，誰敢惹他呢？
GEN|49|10|權杖必不離 猶大 ， 統治者的杖必不離他兩腳之間， 直等細羅 來到， 萬民都要歸順他。
GEN|49|11|猶大 把小驢拴在葡萄樹上， 把驢駒拴在佳美的葡萄樹上。 他在葡萄酒中洗衣服， 在葡萄汁 中洗長袍。
GEN|49|12|他的眼睛比 酒紅潤， 他的牙齒比奶潔白。
GEN|49|13|西布倫 必住在海邊， 必成為停船的港口； 他的疆界必延到 西頓 。
GEN|49|14|以薩迦 是匹強壯的驢， 臥在羊圈之中。
GEN|49|15|他看見居所安舒， 土地肥美， 就屈肩負重， 成為服勞役的僕人。
GEN|49|16|但 必為他的百姓伸冤 ， 作為 以色列 支派之一。
GEN|49|17|但 必作道旁的蛇， 路邊的毒蛇， 咬傷馬蹄， 使騎馬的人向後墜落。
GEN|49|18|耶和華啊，我等候你的救恩。
GEN|49|19|迦得 必被襲擊者襲擊 ， 他卻要襲擊他們的腳跟。
GEN|49|20|亞設 必出豐盛的糧食， 要供應君王的佳肴。
GEN|49|21|拿弗他利 是被釋放的母鹿， 他要生出可愛的小鹿 。
GEN|49|22|約瑟 是多結果子的樹枝， 是泉旁多結果的枝子； 他的枝條伸出牆外。
GEN|49|23|弓箭手惡意攻擊他， 敵對他，向他射箭。
GEN|49|24|但他的弓仍舊堅硬， 他的手臂靈活敏捷， 這是因 雅各 的大能者的手， 從那裏，他是 以色列 的牧者， 以色列 的磐石 。
GEN|49|25|你父親的上帝必幫助你； 全能者必賜福給你： 天上的福， 深淵下面蘊藏的福， 以及生育哺養的福。
GEN|49|26|你父親的福 勝過我祖先的福， 直到永世山嶺的極限。 這些福必降在 約瑟 的頭上， 臨到那與兄弟有分別之人的頭頂上。
GEN|49|27|便雅憫 是隻抓撕掠物的狼， 早晨要吃他的獵物， 晚上要分他的擄物。」
GEN|49|28|這一切是 以色列 的十二個支派。這是他們的父親對他們所說的話，他按照各人的福分為他們祝福。
GEN|49|29|他又吩咐他們說：「我快要歸到我祖先 那裏。你們要將我葬在 赫 人 以弗崙 田間的洞裏，與我的祖先在一處，
GEN|49|30|就是在 迦南 地 幔利 對面的 麥比拉 田間的洞裏，那田是 亞伯拉罕 向 赫 人 以弗崙 買來作墳地的產業。
GEN|49|31|亞伯拉罕 和他的妻子 撒拉 葬在那裏； 以撒 和他的妻子 利百加 也葬在那裏。我也在那裏葬了 利亞 。
GEN|49|32|那塊田和田間的洞是向 赫 人買的。」
GEN|49|33|雅各 囑咐眾子完畢後，就把腳收在床上斷了氣，歸到他祖先 那裏去了。
GEN|50|1|約瑟 伏在他父親的臉上，在他臉上哭，又親他。
GEN|50|2|約瑟 吩咐伺候他的醫生們用香料塗他父親，醫生就用香料塗了 以色列 。
GEN|50|3|四十天滿了，就是塗香料所規定的日子滿了。 埃及 人為他哀哭了七十天。
GEN|50|4|過了哀悼的日子， 約瑟 對法老家中的人說：「我若在你們眼前蒙恩，請你們對法老說：
GEN|50|5|『我父親曾叫我起誓說：看哪，我快要死了，你要將我葬在 迦南 地，在我為自己所掘的墳墓裏。』現在求你准我上去葬我父親，然後我必回來。」
GEN|50|6|法老說：「你可以上去，照你父親叫你起的誓，將他安葬。」
GEN|50|7|於是 約瑟 上去葬他父親。與他一同上去的有法老的眾臣僕和法老家中的長老，以及 埃及 地所有的長老，
GEN|50|8|還有 約瑟 的全家和他的兄弟們，以及他父親的家屬；只留下他們的孩子和羊群牛群在 歌珊 地。
GEN|50|9|又有車輛和駕駛兵和他一同上去，隊伍非常龐大。
GEN|50|10|他們到了 約旦河 東 亞達 的禾場，就在那裏大大地號咷痛哭。 約瑟 為他父親哀哭了七天。
GEN|50|11|迦南 的居民看見 亞達 禾場上的哀哭，就說：「這是 埃及 人一場極大的哀哭。」因此那地方名叫 亞伯‧麥西 ，是在 約旦河 東。
GEN|50|12|雅各 的兒子們遵照父親的吩咐去辦了，
GEN|50|13|他們把他送到 迦南 地，葬在 幔利 對面的 麥比拉 田間的洞裏；那田是 亞伯拉罕 向 赫 人 以弗崙 買來作墳地的產業。
GEN|50|14|約瑟 葬了他父親以後，就和他的兄弟，以及所有同他上去葬他父親的人，都回 埃及 去了。
GEN|50|15|約瑟 的哥哥們見父親死了，就說：「也許 約瑟 仍然懷恨我們，會照我們從前待他一切的惡，重重報復我們。」
GEN|50|16|他們就傳口信給 約瑟 說：「你父親未死之前曾吩咐說：
GEN|50|17|『你們要對 約瑟 這樣說：從前你哥哥們惡待你，你要饒恕他們的過犯和罪惡。』現在求你饒恕你父親的上帝之僕人們的過犯。」他們對 約瑟 說了這話， 約瑟 就哭了。
GEN|50|18|他的哥哥們又來俯伏在他面前，說：「看哪，我們是你的奴隸。」
GEN|50|19|約瑟 對他們說：「不要怕，我豈能代替上帝呢？
GEN|50|20|從前你們的意思是要害我，但上帝的意思原是好的，要使許多百姓得以存活，成就今日的光景。
GEN|50|21|現在你們不要害怕，我必養活你們和你們的孩子。」於是 約瑟 安慰他們，講了使他們安心的話。
GEN|50|22|約瑟 和他父親的家屬都住在 埃及 。 約瑟 活了一百一十年。
GEN|50|23|約瑟 看到 以法蓮 第三代的子孫。 瑪拿西 的孫子， 瑪吉 的兒子，出生時都放在 約瑟 的膝上。
GEN|50|24|約瑟 對他的兄弟說：「我快要死了，但上帝必定看顧你們，領你們從這地上去，到他起誓應許給 亞伯拉罕 、 以撒 、 雅各 之地。」
GEN|50|25|約瑟 叫 以色列 的子孫起誓：「上帝必定眷顧你們，你們要把我的骸骨從這裏帶上去。」
GEN|50|26|約瑟 死了，那時他一百一十歲。人用香料塗了他，把他收殮在棺材裏，停放在 埃及 。
EXOD|1|1|以色列 的眾兒子各帶著家眷，和 雅各 一同來到 埃及 ，他們的名字如下：
EXOD|1|2|呂便 、 西緬 、 利未 、 猶大 、
EXOD|1|3|以薩迦 、 西布倫 、 便雅憫 、
EXOD|1|4|但 、 拿弗他利 、 迦得 、 亞設 。
EXOD|1|5|凡從 雅各 生的，共有七十人。那時， 約瑟 已經在 埃及 。
EXOD|1|6|約瑟 和他所有的兄弟，以及那一代的人都死了。
EXOD|1|7|然而， 以色列 人生養眾多，繁衍昌盛，極其強盛，遍滿了那地。
EXOD|1|8|有一位不認識 約瑟 的新王興起，統治 埃及 。
EXOD|1|9|他對自己的百姓說：「看哪， 以色列 人的百姓比我們還多，又比我們強盛。
EXOD|1|10|來吧，讓我們機巧地待他們，恐怕他們增多起來，將來若有戰爭，他們就聯合我們的仇敵來攻擊我們，然後離開這地去了。」
EXOD|1|11|於是 埃及 人派監工管轄他們，用勞役苦待他們。他們為法老建造儲貨城，就是 比東 和 蘭塞 。
EXOD|1|12|可是越苦待他們，他們就越發增多，更加繁衍， 埃及 人就因 以色列 人愁煩。
EXOD|1|13|埃及 人嚴厲地強迫 以色列 人做工，
EXOD|1|14|使他們因苦工而生活痛苦；無論是和泥，是做磚，是做田間各樣的工，一切的工 埃及 人都嚴厲地對待他們。
EXOD|1|15|埃及 王又對 希伯來 的接生婆，一個名叫 施弗拉 ，另一個名叫 普阿 的說：
EXOD|1|16|「你們為 希伯來 婦人接生，臨盆的時候要注意 ，若是男的，就把他殺了，若是女的，就讓她活。」
EXOD|1|17|但是接生婆敬畏上帝，不照 埃及 王的吩咐去做，卻讓男孩活著。
EXOD|1|18|埃及 王召了接生婆來，對她們說：「你們為甚麼做這事，讓男孩活著呢？」
EXOD|1|19|接生婆對法老說：「因為 希伯來 婦人與 埃及 婦人不同； 希伯來 婦人健壯，接生婆還沒有到，她們已經生產了。」
EXOD|1|20|上帝恩待接生婆； 以色列 人增多起來，極其強盛。
EXOD|1|21|接生婆因為敬畏上帝，上帝就叫她們成立家室。
EXOD|1|22|法老吩咐他的眾百姓說：「把所生的 每一個男孩都丟到 尼羅河 裏去，讓所有的女孩存活。」
EXOD|2|1|有一個 利未 家的人娶了一個 利未 女子為妻。
EXOD|2|2|那女人懷孕，生了一個兒子，見他俊美，就把他藏了三個月，
EXOD|2|3|後來不能再藏，就取了一個蒲草箱，抹上柏油和樹脂，將孩子放在裏面，把箱子擱在 尼羅河 邊的蘆葦中。
EXOD|2|4|孩子的姊姊遠遠站著，要知道他究竟會怎樣。
EXOD|2|5|法老的女兒來到 尼羅河 邊洗澡，她的女僕們在河邊行走。她看見在蘆葦中的箱子，就派一個使女把它拿來。
EXOD|2|6|她打開箱子，看見那孩子。看哪，男孩在哭，她就可憐他，說：「這是 希伯來 人的一個孩子。」
EXOD|2|7|孩子的姊姊對法老的女兒說：「我去叫一個 希伯來 婦人來作奶媽，替你乳養這孩子，好嗎？」
EXOD|2|8|法老的女兒對她說：「去吧！」那女孩就去叫了孩子的母親來。
EXOD|2|9|法老的女兒對她說：「你把這孩子抱去，替我乳養這孩子，我必給你工錢。」那婦人就把孩子接過來，乳養他。
EXOD|2|10|孩子長大了，婦人把他帶到法老的女兒那裏，就作了她的兒子。她給孩子起名叫 摩西 ，說：「因我把他從水裏拉出來。」
EXOD|2|11|過了一段日子， 摩西 長大了，他出去到他同胞那裏，看見他們的勞役。他看見一個 埃及 人打他的同胞，一個 希伯來 人。
EXOD|2|12|他左右觀看，見沒有人，就把 埃及 人打死了，藏在沙土裏。
EXOD|2|13|第二天他出去，看哪，有兩個 希伯來 人在打架，他就對那兇惡的人說：「你為甚麼打你同族的人呢？」
EXOD|2|14|那人說：「誰立你作我們的領袖和審判官呢？難道你要殺我，像殺那 埃及 人一樣嗎？」 摩西 就懼怕，說：「這事一定是讓人知道了。」
EXOD|2|15|法老聽見這事，就設法要殺 摩西 。於是 摩西 逃走，躲避法老，到了 米甸 地，坐在井旁。
EXOD|2|16|米甸 的祭司有七個女兒；她們來打水，打滿了槽，要給父親的羊群喝水。
EXOD|2|17|有一些牧羊人來，把她們趕走， 摩西 卻起來幫助她們，取水給她們的羊群喝。
EXOD|2|18|她們回到父親 流珥 那裏；他說：「今日你們為何這麼快就回來了呢？」
EXOD|2|19|她們說：「有一個 埃及 人來救我們脫離牧羊人的手，他甚至打水給我們的羊群喝。」
EXOD|2|20|他對女兒們說：「那人在哪裏？你們為甚麼撇下他呢？去請他來吃飯吧！」
EXOD|2|21|摩西 願意和那人同住， 那人就把女兒 西坡拉 給 摩西 為妻。
EXOD|2|22|西坡拉 生了一個兒子， 摩西 給他起名叫 革舜 ，因他說：「我在外地作了寄居者。」
EXOD|2|23|過了許多年， 埃及 王死了。 以色列 人因做苦工，就嘆息哀求；他們因苦工所發出的哀聲達於上帝。
EXOD|2|24|上帝聽見他們的哀聲，就記念他與 亞伯拉罕 、 以撒 、 雅各 所立的約。
EXOD|2|25|上帝看顧 以色列 人，上帝是知道的 。
EXOD|3|1|摩西 牧放他岳父 米甸 祭司 葉特羅 的羊群，他領羊群往曠野的那一邊去，到了上帝的山，就是 何烈山 。
EXOD|3|2|耶和華的使者在荊棘的火焰中向他顯現。 摩西 觀看，看哪，荊棘在火中焚燒，卻沒有燒燬。
EXOD|3|3|摩西 說：「我要轉過去看這大異象，這荊棘為何沒有燒燬呢？」
EXOD|3|4|耶和華見 摩西 轉過去看，上帝就從荊棘裏呼叫他說：「 摩西 ！ 摩西 ！」他說：「我在這裏。」
EXOD|3|5|上帝說：「不要靠近這裏。把你腳上的鞋脫下來，因為你所站的地方是聖地」。
EXOD|3|6|他又說：「我是你父親的上帝，是 亞伯拉罕 的上帝， 以撒 的上帝， 雅各 的上帝。」 摩西 蒙上臉，因為怕看上帝。
EXOD|3|7|耶和華說：「我確實看見了我百姓在 埃及 所受的困苦，我也聽見了他們因受監工苦待所發的哀聲；我確實知道他們的痛苦。
EXOD|3|8|我下來是要救他們脫離 埃及 人的手，領他們從那地上來，到美好與寬闊之地，到流奶與蜜之地，就是 迦南 人、 赫 人、 亞摩利 人、 比利洗 人、 希未 人、 耶布斯 人之地。
EXOD|3|9|現在，看哪， 以色列 人的哀聲達到我這裏，我也看見 埃及 人怎樣欺壓他們。
EXOD|3|10|現在，你去，我要差派你到法老那裏，把我的百姓 以色列 人從 埃及 領出來。」
EXOD|3|11|摩西 對上帝說：「我是甚麼人，竟能去見法老，把 以色列 人從 埃及 領出來呢？」
EXOD|3|12|上帝說：「我必與你同在。這就是我差派你去，給你的憑據：你把百姓從 埃及 領出來之後，你們必在這山上事奉上帝。」
EXOD|3|13|摩西 對上帝說：「看哪，我到 以色列 人那裏，對他們說：『你們祖宗的上帝差派我到你們這裏來。』他們若對我說：『他叫甚麼名字？』我要對他們說甚麼呢？」
EXOD|3|14|上帝對 摩西 說：「我是自有永有的」；又說：「你要對 以色列 人這樣說：『那自有永有的差派我到你們這裏來。』」
EXOD|3|15|上帝又對 摩西 說：「你要對 以色列 人這樣說：『耶和華－你們祖宗的上帝，就是 亞伯拉罕 的上帝， 以撒 的上帝， 雅各 的上帝差派我到你們這裏來。』這是我的名，直到永遠；這也是我的稱號 ，直到萬代。
EXOD|3|16|你去召集 以色列 的長老，對他們說：『耶和華－你們祖宗的上帝，就是 亞伯拉罕 的上帝， 以撒 的上帝， 雅各 的上帝向我顯現，說：我實在眷顧了你們，眷顧你們在 埃及 的遭遇。
EXOD|3|17|我也曾說：要把你們從 埃及 的困苦中領出來，往 迦南 人、 赫 人、 亞摩利 人、 比利洗 人、 希未 人、 耶布斯 人的地去，就是到流奶與蜜之地。』
EXOD|3|18|他們必聽你的話。你和 以色列 的長老要到 埃及 王那裏，對他說：『耶和華－ 希伯來 人的上帝向我們顯現，現在求你讓我們往曠野去，走三天的路程，為要向耶和華我們的上帝獻祭。』
EXOD|3|19|我知道若不用大能的手， 埃及 王不會放你們走。
EXOD|3|20|因此，我必伸出我的手，在 埃及 施行我一切的神蹟，擊打這地，然後，他才放你們走。
EXOD|3|21|我必使 埃及 人看得起你們，你們離開的時候就不至於空手而去。
EXOD|3|22|每一個婦女必向她的鄰舍，以及寄居在她家裏的女人，索取金器、銀器和衣裳，給你們的兒女穿戴。這樣你們就掠奪了 埃及 人。」
EXOD|4|1|摩西 回答說：「看哪！他們不會信我，也不會聽我的話，因為他們必說：『耶和華並沒有向你顯現。』」
EXOD|4|2|耶和華對 摩西 說：「你手裏的是甚麼？」他說：「是杖。」
EXOD|4|3|耶和華說：「把它丟在地上！」他一丟在地上，杖就變成一條蛇； 摩西 逃走避開牠。
EXOD|4|4|耶和華對 摩西 說：「伸出手來，拿住牠的尾巴─ 摩西 就伸出手，抓住牠，牠就在 摩西 的手掌中變為杖─
EXOD|4|5|為了要使他們信耶和華他們祖宗的上帝，就是 亞伯拉罕 的上帝， 以撒 的上帝， 雅各 的上帝，曾向你顯現了。」
EXOD|4|6|耶和華又對他說：「把手放進懷裏。」他就把手放進懷裏。當他把手抽出來，看哪，手竟然長了痲瘋 ，像雪一樣白。
EXOD|4|7|耶和華說：「把手放回懷裏─他就把手放回懷裏。當他把手從懷裏再抽出來，看哪，手復原了，與全身的肉一樣─
EXOD|4|8|倘若他們不信你，也不聽第一個神蹟的聲音，他們會信第二個神蹟的聲音。
EXOD|4|9|倘若他們不信這兩個神蹟，不聽你的話，你就從 尼羅河 裏取些水，倒在乾的地上。你從 尼羅河 裏所取的水必在乾地上變成血。」
EXOD|4|10|摩西 對耶和華說：「主啊，求求你，我並不是一個能言善道的人，以前這樣，就是你對僕人說話以後也是這樣，因為我是拙口笨舌的。」
EXOD|4|11|耶和華對他說：「誰造人的口呢？誰使人口啞、耳聾、目明、眼瞎呢？豈不是我－耶和華嗎？
EXOD|4|12|現在，去吧，我必賜你口才，指教你應當說的。」
EXOD|4|13|摩西 說：「主啊，求求你，你要藉著誰的手，就差派誰去吧！」
EXOD|4|14|耶和華的怒氣向 摩西 發作，說：「你不是有一個哥哥 利未 人 亞倫 嗎？我知道他是個能言善道的人。看哪，他正出來迎接你。他一見到你，心裏就歡喜。
EXOD|4|15|你要跟他說話，把話放在他的口裏，我要賜你口才，也要賜他口才，又要教你們做當做的事。
EXOD|4|16|他要替你向百姓說話；他要當你的口，你要當他的上帝。
EXOD|4|17|你手裏要拿這杖，用它來行神蹟。」
EXOD|4|18|於是， 摩西 回到他岳父 葉特羅 那裏，對他說：「請你讓我回 埃及 我同胞那裏，看他們還在不在。」 葉特羅 對 摩西 說：「平平安安地去吧！」
EXOD|4|19|耶和華在 米甸 對 摩西 說：「你要回 埃及 去，因為那些尋索你命的人都死了。」
EXOD|4|20|摩西 就帶著妻子和兩個兒子，讓他們騎上驢，回 埃及 地去。 摩西 手裏拿著上帝的杖。
EXOD|4|21|耶和華對 摩西 說：「你回到 埃及 去的時候，要留意將我交在你手中的一切奇事行在法老面前。但我要任憑他的心剛硬，他必不放百姓走。
EXOD|4|22|你要對法老說：『耶和華如此說： 以色列 是我的兒子，我的長子。
EXOD|4|23|我對你說過：放我的兒子走，好事奉我。你還是不肯放他走。看哪，我要殺你頭生的兒子。』」
EXOD|4|24|在路上住宿的地方，耶和華遇見 摩西 ，想要殺他。
EXOD|4|25|西坡拉 就拿一塊火石，割下她兒子的包皮，碰觸 摩西 的腳，說：「你真是我血的新郎了。」
EXOD|4|26|這樣，耶和華才放了他。那時， 西坡拉 說：「你因割禮就是血的新郎 了」。
EXOD|4|27|耶和華對 亞倫 說：「你往曠野去迎接 摩西 。」他就去，在上帝的山遇見 摩西 ，就親他。
EXOD|4|28|摩西 將耶和華差派他所說的話和吩咐他所行的神蹟都告訴了 亞倫 。
EXOD|4|29|摩西 和 亞倫 就去召集 以色列 的眾長老。
EXOD|4|30|亞倫 將耶和華對 摩西 所說的一切話述說了一遍，又在百姓眼前行了那些神蹟，
EXOD|4|31|百姓就信了。他們聽見耶和華眷顧 以色列 人，鑒察他們的困苦，就低頭敬拜。
EXOD|5|1|後來， 摩西 和 亞倫 去對法老說：「耶和華－ 以色列 的上帝這樣說：『放我的百姓走，好讓他們在曠野向我守節。』」
EXOD|5|2|法老說：「耶和華是誰，要我聽他的話，讓 以色列 人去？我不認識耶和華，也不放 以色列 人走！」
EXOD|5|3|他們說：「 希伯來 人的上帝已向我們顯現了。求你讓我們往曠野去，走三天的路程，向耶和華我們的上帝獻祭，免得他用瘟疫、刀劍攻擊我們。」
EXOD|5|4|埃及 王對他們說：「 摩西 、 亞倫 ！你們為甚麼叫百姓不做工呢？去，服你們的勞役吧！」
EXOD|5|5|他又說：「看哪，這地的 以色列 人如今這麼多，你們竟然叫他們歇下勞役！」
EXOD|5|6|當天，法老吩咐監工和工頭說：
EXOD|5|7|「你們不可照以前一樣提供草給百姓做磚，要叫他們自己去撿草。
EXOD|5|8|他們平時做磚的數目，你們仍舊向他們要，一點不可減少，因為他們是懶惰的，所以才呼求說：『讓我們去向我們的上帝獻祭。』
EXOD|5|9|你們要把更重的工作加在這些人身上，使他們在其中勞碌，不去理會謊言。」
EXOD|5|10|監工和工頭出來對百姓說：「法老這樣說：『我不給你們草，
EXOD|5|11|你們自己在哪裏能找到草，就往哪裏去找吧！但你們的工作一點也不可減少。』」
EXOD|5|12|於是，百姓分散在 埃及 全地，撿碎秸當草用。
EXOD|5|13|監工催逼他們，說：「你們每天要做完一天的工，與先前有草一樣。」
EXOD|5|14|法老的監工擊打他們所派的 以色列 工頭，說：「為甚麼昨天和今天你們沒有按照以前做磚的數目，完成你們的工作呢？」
EXOD|5|15|以色列 人的工頭來哀求法老說：「為甚麼這樣待你的僕人呢？
EXOD|5|16|監工不把草給僕人，並且對我們說：『做磚吧！』看哪，你僕人挨了打，其實是你百姓的錯。」
EXOD|5|17|法老卻說：「懶惰，你們真是懶惰！所以你們說：『讓我們去向耶和華獻祭吧。』
EXOD|5|18|現在，去做工吧！草是不會給你們，磚卻要如數交納。」
EXOD|5|19|以色列 人的工頭聽見「你們每天做磚的工作一點也不可減少」，就知道惹上禍了。
EXOD|5|20|他們離開法老出來，正遇見 摩西 和 亞倫 站在那裏等候他們，
EXOD|5|21|就向他們說：「願耶和華鑒察你們，施行判斷，因為你們使我們在法老和他臣僕面前有了臭名，把刀遞在他們手中來殺我們。」
EXOD|5|22|摩西 回到耶和華那裏，說：「主啊，你為甚麼苦待這百姓呢？為甚麼差派我呢？
EXOD|5|23|自從我到法老那裏，奉你的名說話，他就苦待這百姓，你卻一點也沒有拯救你的百姓。」
EXOD|6|1|耶和華對 摩西 說：「現在你必看見我向法老所行的事，使他因我大能的手放 以色列 人走，因我大能的手把他們趕出他的地。」
EXOD|6|2|上帝吩咐 摩西 ，對他說：「我是耶和華。
EXOD|6|3|我從前向 亞伯拉罕 、 以撒 、 雅各 顯現為全能的上帝；至於我的名耶和華，我未曾讓他們知道。
EXOD|6|4|我要與他們堅立我的約，要把 迦南 地，他們寄居的地賜給他們。
EXOD|6|5|我聽見 以色列 人被 埃及 人奴役的哀聲，我就記念我的約。
EXOD|6|6|所以你要對 以色列 人說：『我是耶和華；我要除去 埃及 人加給你們的勞役，救你們脫離他們的奴役。我要用伸出來的膀臂，藉嚴厲的懲罰救贖你們。
EXOD|6|7|我要以你們為我的百姓，我也要作你們的上帝。我除去 埃及 人加給你們的勞役，你們就知道我是耶和華你們的上帝。
EXOD|6|8|我起誓應許給 亞伯拉罕 、 以撒 、 雅各 的地，我要領你們進去，將那地賜給你們為業。我是耶和華。』」
EXOD|6|9|摩西 把這話告訴 以色列 人，但是他們因心裏愁煩，又因苦工，就不肯聽 摩西 的話。
EXOD|6|10|耶和華吩咐 摩西 說：
EXOD|6|11|「你去對 埃及 王法老說，讓 以色列 人離開他的地。」
EXOD|6|12|摩西 在耶和華面前說：「看哪， 以色列 人尚且不聽我，法老怎麼會聽我這不會講話的人呢？」
EXOD|6|13|耶和華吩咐 摩西 和 亞倫 ，命令他們到 以色列 人和 埃及 王法老那裏，把 以色列 人從 埃及 地領出來。
EXOD|6|14|以色列 人族長的名字如下： 以色列 長子 呂便 的兒子是 哈諾 、 法路 、 希斯倫 、 迦米 ；這是 呂便 的家族。
EXOD|6|15|西緬 的兒子是 耶母利 、 雅憫 、 阿轄 、 雅斤 、 瑣轄 ，和 迦南 女子生的兒子 掃羅 ；這是 西緬 的家族。
EXOD|6|16|以下是 利未 的兒子按著家譜的名字： 革順 、 哥轄 、 米拉利 。 利未 一生的歲數是一百三十七歲。
EXOD|6|17|革順 的兒子按著家族是 立尼 、 示每 。
EXOD|6|18|哥轄 的兒子是 暗蘭 、 以斯哈 、 希伯倫 、 烏薛 。 哥轄 一生的歲數是一百三十三歲。
EXOD|6|19|米拉利 的兒子是 抹利 和 母示 ；這是 利未 按著家譜的家族。
EXOD|6|20|暗蘭 娶了他父親的妹妹 約基別 為妻，她為他生了 亞倫 和 摩西 。 暗蘭 一生的歲數是一百三十七歲。
EXOD|6|21|以斯哈 的兒子是 可拉 、 尼斐 、 細基利 。
EXOD|6|22|烏薛 的兒子是 米沙利 、 以利撒反 、 西提利 。
EXOD|6|23|亞倫 娶了 亞米拿達 的女兒， 拿順 的妹妹， 以利沙巴 為妻，她為他生了 拿答 、 亞比戶 、 以利亞撒 、 以他瑪 。
EXOD|6|24|可拉 的兒子是 亞惜 、 以利加拿 、 亞比亞撒 ；這是 可拉 的家族。
EXOD|6|25|亞倫 的兒子 以利亞撒 娶了 普鐵 的一個女兒為妻，她為他生了 非尼哈 。這是 利未 人按著家族的族長。
EXOD|6|26|這就是曾聽見耶和華說「把 以色列 人按著隊伍從 埃及 地領出來」的 亞倫 和 摩西 ，
EXOD|6|27|對 埃及 王法老說要將 以色列 人從 埃及 領出來的，也是這 摩西 和 亞倫 。
EXOD|6|28|當耶和華在 埃及 地對 摩西 說話的時候，
EXOD|6|29|耶和華對 摩西 說：「我是耶和華；我對你所說的一切話，你都要告訴 埃及 王法老。」
EXOD|6|30|摩西 在耶和華面前說：「看哪，我是不會講話的人，法老怎麼會聽我呢？」
EXOD|7|1|耶和華對 摩西 說：「我使你在法老面前像上帝一樣，你的哥哥 亞倫 是你的代言人 。
EXOD|7|2|凡我所吩咐你的，你都要說。你的哥哥 亞倫 要對法老說，讓 以色列 人離開他的地。
EXOD|7|3|我要使法老的心固執，我也要在 埃及 地多行神蹟奇事。
EXOD|7|4|法老必不聽從你們，因此我要伸手嚴厲地懲罰 埃及 ，把我的軍隊，就是我的百姓 以色列 人從 埃及 地領出來。
EXOD|7|5|我伸手攻擊 埃及 ，把 以色列 人從他們中間領出來的時候， 埃及 人就知道我是耶和華。」
EXOD|7|6|摩西 和 亞倫 就去做；他們照耶和華吩咐的去做了。
EXOD|7|7|摩西 和 亞倫 與法老說話的時候， 摩西 八十歲， 亞倫 八十三歲。
EXOD|7|8|耶和華對 摩西 和 亞倫 說：
EXOD|7|9|「法老若吩咐你們說：『你們行一件奇事吧！』你就對 亞倫 說：『把杖丟在法老面前！杖會變成蛇。』」
EXOD|7|10|摩西 和 亞倫 到法老那裏去，照耶和華所吩咐的去做。 亞倫 把杖丟在法老和他臣僕面前，杖就變成蛇。
EXOD|7|11|法老也召了智慧人和行邪術的人來，這些 埃及 術士也用邪術照樣做。
EXOD|7|12|他們各人丟下自己的杖，杖就變成蛇；但 亞倫 的杖吞了他們的杖。
EXOD|7|13|法老心裏剛硬，不聽 摩西 和 亞倫 ，正如耶和華所說的。
EXOD|7|14|耶和華對 摩西 說：「法老心硬，不肯放百姓走。
EXOD|7|15|明天早晨你要到法老那裏去，看哪，他出來往水邊去，你要到 尼羅河 邊去迎見他，手裏拿著那根變過蛇的杖。
EXOD|7|16|你要對他說：『耶和華－ 希伯來 人的上帝差派我到你這裏，說：放我的百姓走，到曠野事奉我。看哪，到如今你還是不聽。
EXOD|7|17|耶和華如此說：看哪，我要用我手裏的杖擊打 尼羅河 中的水，水就變成血；這樣，你就知道我是耶和華。
EXOD|7|18|河裏的魚必死，河也要發臭， 埃及 人就厭惡喝這河裏的水。』」
EXOD|7|19|耶和華對 摩西 說：「你要對 亞倫 說：『拿你的杖，伸出你的手在 埃及 所有的水上，在他們的江、河、池塘，所有水聚集的地方上，叫水變成血。在 埃及 全地，無論在木器中，石器中，都必有血。』」
EXOD|7|20|摩西 和 亞倫 就照耶和華所吩咐的去做。 亞倫 在法老和他臣僕眼前舉杖擊打 尼羅河 裏的水，河裏的水都變成血了。
EXOD|7|21|河裏的魚死了，河也臭了， 埃及 人就不能喝這河裏的水； 埃及 遍地都有了血。
EXOD|7|22|但是， 埃及 的術士也用邪術照樣做了；法老心裏剛硬，不聽 摩西 和 亞倫 ，正如耶和華所說的。
EXOD|7|23|法老轉身回宮去，並不把這事放在心上。
EXOD|7|24|所有的 埃及 人都沿著 尼羅河 邊挖掘，要找水喝，因為他們不能喝河裏的水。
EXOD|7|25|耶和華擊打 尼羅河 後，過了七天。
EXOD|8|1|耶和華對 摩西 說：「你要到法老那裏，對他說：『耶和華如此說：放我的百姓走，好事奉我。
EXOD|8|2|你若不肯放他們走，看哪，我必以青蛙之災擊打你的疆土。
EXOD|8|3|尼羅河 要滋生青蛙；這青蛙要上來進你的宮殿和你的臥房，上你的床榻，進你臣僕的房屋，上你百姓的身上，進你的爐灶和你的揉麵盆。
EXOD|8|4|這些青蛙要跳上你、你百姓和你眾臣僕的身上。』」
EXOD|8|5|耶和華對 摩西 說：「你要對 亞倫 說：『伸出你手裏的杖在江、河、池塘上，把青蛙帶上 埃及 地來。』」
EXOD|8|6|亞倫 伸手在 埃及 的眾水上，青蛙就上來，遮滿了 埃及 地。
EXOD|8|7|術士也用他們的邪術照樣去做，把青蛙帶上 埃及 地。
EXOD|8|8|法老召 摩西 和 亞倫 來，說：「請你們祈求耶和華使這些青蛙離開我和我的百姓，我就讓這百姓去向耶和華獻祭。」
EXOD|8|9|摩西 對法老說：「悉聽尊便，告訴我何時為你、你臣僕和你的百姓祈求，使青蛙被剪除，離開你和你的宮殿，只留在 尼羅河 裏。」
EXOD|8|10|他說：「明天。」 摩西 說：「就照你的話吧，為要叫你知道沒有像耶和華我們上帝的，
EXOD|8|11|青蛙必會離開你、你宮殿、你臣僕和你的百姓，只留在 尼羅河 裏。」
EXOD|8|12|於是 摩西 和 亞倫 離開法老出去。 摩西 為了青蛙的事呼求耶和華，因為他帶來青蛙攪擾法老。
EXOD|8|13|耶和華就照 摩西 的請求去做；在屋裏、院中、田間的青蛙都死了。
EXOD|8|14|眾人把青蛙聚攏成堆，地就發出臭氣。
EXOD|8|15|但法老見災禍舒緩了，就硬著心，不聽從他們，正如耶和華所說的。
EXOD|8|16|耶和華對 摩西 說：「你要對 亞倫 說：『伸出你的杖擊打地上的塵土，使塵土在 埃及 全地變成蚊子 。』」
EXOD|8|17|他們就照樣做了。 亞倫 伸出他手裏的杖，擊打地上的塵土，人和牲畜身上就有了蚊子； 埃及 全地的塵土都變成蚊子了。
EXOD|8|18|術士也用邪術要照樣產生蚊子，卻做不成。於是人和牲畜的身上都有了蚊子。
EXOD|8|19|術士對法老說：「這是上帝的手指。」法老心裏剛硬，不聽 摩西 和 亞倫 ，正如耶和華所說的。
EXOD|8|20|耶和華對 摩西 說：「你要清早起來，站在法老面前。看哪，法老來到水邊，你就對他說：『耶和華如此說：放我的百姓走，好事奉我。
EXOD|8|21|你若不放我的百姓走，看哪，我要派成群的蒼蠅到你、你臣僕和你百姓身上，進你的宮殿； 埃及 人的房屋和他們所住的地都要滿了成群的蒼蠅。
EXOD|8|22|那一日，我必把我百姓所住的 歌珊 地分別出來，使那裏沒有成群的蒼蠅，好叫你知道我─耶和華是在全地之中。
EXOD|8|23|我要施行救贖，區隔我的百姓和你的百姓。明天必有這神蹟。』」
EXOD|8|24|耶和華就這樣做了。大群的蒼蠅進入法老的宮殿和他臣僕的房屋；在 埃及 全地，地就因這成群的蒼蠅毀壞了。
EXOD|8|25|法老召了 摩西 和 亞倫 來，說：「去，在此地向你們的上帝獻祭。」
EXOD|8|26|摩西 說：「這樣做是不妥的，因為我們要獻給耶和華－我們上帝的祭物是 埃及 人所厭惡的；看哪，我們在 埃及 人眼前獻他們所厭惡的，他們豈不拿石頭打死我們嗎？
EXOD|8|27|我們要遵照耶和華－我們上帝所吩咐我們的，往曠野去，走三天路程，向他獻祭。」
EXOD|8|28|法老說：「我可以放你們走，在曠野向耶和華－你們的上帝獻祭，只是不可走得太遠。你們要為我祈禱。」
EXOD|8|29|摩西 說：「看哪，我要從你這裏出去祈求耶和華，使成群的蒼蠅明天離開法老、法老的臣僕和法老的百姓；法老卻不可再欺騙，不讓百姓去向耶和華獻祭。」
EXOD|8|30|於是 摩西 離開法老，去祈求耶和華。
EXOD|8|31|耶和華就照 摩西 的請求去做，使成群的蒼蠅離開法老、他的臣僕和他的百姓，一隻也沒有留下。
EXOD|8|32|但這一次法老又硬著心，不放百姓走。
EXOD|9|1|耶和華對 摩西 說：「你要到法老那裏，對他說：『耶和華－ 希伯來 人的上帝如此說：放我的百姓走，好事奉我。
EXOD|9|2|你若不肯放他們走，仍要強留他們，
EXOD|9|3|看哪，耶和華的手必以嚴重的瘟疫加在你田間的牲畜上，就是在馬、驢、駱駝、牛群和羊群的身上。
EXOD|9|4|耶和華卻要分別 以色列 的牲畜和 埃及 的牲畜，凡屬 以色列 人的，一隻都不死。』」
EXOD|9|5|耶和華就設定時間，說：「明天耶和華必在此地行這事。」
EXOD|9|6|第二天，耶和華行了這事。 埃及 的牲畜全都死了，只是 以色列 人的牲畜，一隻都沒有死。
EXOD|9|7|法老派人去，看哪， 以色列 人的牲畜連一隻都沒有死。可是法老硬著心，不放百姓走。
EXOD|9|8|耶和華對 摩西 和 亞倫 說：「你們從爐裏滿滿捧出爐灰， 摩西 要在法老眼前把它撒在空中。
EXOD|9|9|這灰要在 埃及 全地變成塵土，使 埃及 全地的人和牲畜身上起泡生瘡。」
EXOD|9|10|摩西 和 亞倫 取了爐灰，站在法老面前。 摩西 把它撒在空中，人和牲畜的身上就起泡生瘡了。
EXOD|9|11|因為這瘡，術士在 摩西 面前站立不住，術士和所有 埃及 人的身上都生了瘡。
EXOD|9|12|但耶和華任憑法老的心剛硬，不聽 摩西 和 亞倫 ，正如耶和華對 摩西 所說的。
EXOD|9|13|耶和華對 摩西 說：「你要清早起來，站在法老面前，對他說：『耶和華－ 希伯來 人的上帝如此說：放我的百姓走，好事奉我。
EXOD|9|14|因為這一次我要使一切的災禍臨到你自己，你臣僕和你百姓的身上，為要叫你知道在全地沒有像我的。
EXOD|9|15|現在，我若伸手用瘟疫攻擊你和你的百姓，你就會從地上除滅了。
EXOD|9|16|然而，我讓你存活，是為了要使你看見我的大能，並要使我的名傳遍全地。
EXOD|9|17|可是你仍然向我的百姓自高自大，不放他們走。
EXOD|9|18|看哪，明天大約這時候，我必使大量的冰雹降下，這是從 埃及 立國直到如今沒有出現過的。
EXOD|9|19|現在，你要派人把你的牲畜和你田間一切所有的帶去躲避；任何在田間，無論是人是牲畜沒有回到屋內的，冰雹必降在他們身上，他們就必死。』」
EXOD|9|20|法老的臣僕中，懼怕耶和華這話的，就讓他的奴僕和牲畜逃進屋裏。
EXOD|9|21|但那不把耶和華這話放在心上的，就把他的奴僕和牲畜留在田裏。
EXOD|9|22|耶和華對 摩西 說：「你向天伸出你的手，使冰雹降在 埃及 全地，降在 埃及 地的人和牲畜身上，以及田間各樣菜蔬上。」
EXOD|9|23|摩西 向天伸杖，耶和華就打雷下雹，有火降到地上；耶和華下雹在 埃及 地上。
EXOD|9|24|那時，有雹，也有火在雹中閃爍，極其嚴重；自從 埃及 立國以來，全地沒有像這樣的。
EXOD|9|25|在 埃及 全地，冰雹擊打田間所有的人和牲畜，擊打一切的菜蔬，也打壞了田間一切的樹木。
EXOD|9|26|惟獨 以色列 人所住的 歌珊 地沒有冰雹。
EXOD|9|27|法老差派人去召 摩西 和 亞倫 來，對他們說：「這一次我犯罪了。耶和華是公義的；我和我的百姓是邪惡的。
EXOD|9|28|請你們祈求耶和華，因上帝的雷轟和冰雹已經夠了。我要放你們走，你們不用再留下來了。」
EXOD|9|29|摩西 對他說：「我一出城就向耶和華舉起雙手；雷必止住，也不再有冰雹，叫你知道地是屬於耶和華的。
EXOD|9|30|至於你和你的臣僕，我知道你們仍然不敬畏耶和華上帝。」
EXOD|9|31|那時，亞麻和大麥被摧毀了，因為大麥已經吐穗，亞麻也開了花。
EXOD|9|32|只是小麥和粗麥沒有被摧毀，因為它們還沒有長成。
EXOD|9|33|摩西 離開法老出了城，向耶和華舉起雙手，雷和雹就止住，雨也不再下在地上了。
EXOD|9|34|法老見雨、雹、雷止住，又再犯罪；他和他的臣僕都硬著心。
EXOD|9|35|法老的心剛硬，不放 以色列 人走，正如耶和華藉著 摩西 所說的。
EXOD|10|1|耶和華對 摩西 說：「你要到法老那裏，因我使他硬著心，也使他臣僕硬著心，為要在他們中間 顯出我的這些神蹟來，
EXOD|10|2|並要叫你將我嚴厲對付 埃及 的事，和在他們中間所行的神蹟，傳於兒子和孫子的耳中，好叫你們知道我是耶和華。」
EXOD|10|3|摩西 和 亞倫 就到法老那裏，對他說：「耶和華－ 希伯來 人的上帝這樣說：『你在我面前不肯謙卑要到幾時呢？放我的百姓走，好事奉我。
EXOD|10|4|你若不肯放我的百姓走，看哪，明天我要使蝗蟲進入你的境內，
EXOD|10|5|遮滿地面 ，甚至地也看不見了。牠們要吃那冰雹後所剩，就是留給你們的；並且要吃那生長在田間的一切樹木。
EXOD|10|6|你的宮殿和你眾臣僕的房屋，以及一切 埃及 人的房屋，都要被蝗蟲佔滿；你祖宗和你祖宗的祖宗在世以來，直到今日都沒有見過。』」 摩西 就轉身離開法老出去。
EXOD|10|7|法老的臣僕對法老說：「這傢伙成為我們的羅網要到幾時呢？讓這些人去事奉耶和華－他們的上帝吧！ 埃及 快要滅亡了，你還不知道嗎？」
EXOD|10|8|於是 摩西 和 亞倫 被召回來見法老。法老對他們說：「去，事奉耶和華－你們的上帝吧！但要去的是哪些人呢？」
EXOD|10|9|摩西 說：「我們要帶著年老的和年少的同去，要帶著我們的兒子和女兒，以及我們的羊群牛群一起去，因為我們要向耶和華守節。」
EXOD|10|10|法老對他們說：「願耶和華與你們同在吧！我若讓你們帶著你們的孩子同去，看，災禍就在你們面前 ！
EXOD|10|11|不可都去！你們壯年人去事奉耶和華吧，因為這是你們所求的。」於是法老把他們從自己面前趕出去。
EXOD|10|12|耶和華對 摩西 說：「你向 埃及 地伸出你的手，使蝗蟲上到 埃及 地，吃地上冰雹後所剩一切的植物。」
EXOD|10|13|摩西 就向 埃及 地伸杖；整整一晝一夜，耶和華使東風颳在 埃及 地上，到了早晨，東風把蝗蟲颳了來。
EXOD|10|14|蝗蟲上到 埃及 全地，落在 埃及 全境，非常厲害；蝗蟲這麼多，是空前絕後的。
EXOD|10|15|蝗蟲遮滿地面，地上一片黑暗。牠們吃盡了地上一切的植物和冰雹過後所剩樹上的果子。 埃及 全地，無論是樹木，是田間的植物，連一點綠的也沒有留下。
EXOD|10|16|於是法老急忙召了 摩西 和 亞倫 來，說：「我得罪了耶和華－你們的上帝，又得罪了你們。
EXOD|10|17|現在求你，就這一次，饒恕我的罪，祈求耶和華－你們的上帝救我脫離這次的死亡。」
EXOD|10|18|摩西 就離開法老，去祈求耶和華。
EXOD|10|19|耶和華轉變風向，使強勁的西風吹來，把蝗蟲颳起，吹入 紅海 ；在 埃及 全境連一隻也沒有留下。
EXOD|10|20|但耶和華任憑法老的心剛硬，不放 以色列 人走。
EXOD|10|21|耶和華對 摩西 說：「你向天伸出你的手，使黑暗籠罩 埃及 地；這黑暗甚至可以摸得到。」
EXOD|10|22|摩西 向天伸出他的手，濃密的黑暗就籠罩了 埃及 全地三天之久。
EXOD|10|23|三天內，人人彼此看不見，誰也不敢起身離開原地；但所有 以色列 人住的地方卻有光。
EXOD|10|24|法老就召 摩西 來，說：「去，事奉耶和華吧！只是你們的羊群牛群要留下來。你們的孩子可以和你們同去。」
EXOD|10|25|摩西 說：「你必須把祭物和燔祭牲交在我們手中，讓我們可以向耶和華我們的上帝獻祭。
EXOD|10|26|我們的牲畜也要與我們同去，連一蹄也不留下，因為我們要從牲畜中挑選來事奉耶和華－我們的上帝。未到那裏之前，我們還不知道要用甚麼來事奉耶和華。」
EXOD|10|27|但耶和華任憑法老的心剛硬，法老不肯放他們走。
EXOD|10|28|法老對 摩西 說：「離開我去吧！你要小心，不要再見我的面，因為再見我面的那日，你就必死！」
EXOD|10|29|摩西 說：「就照你說的，我也不要再見你的面了！」
EXOD|11|1|耶和華對 摩西 說：「我要再降一個災禍給法老和 埃及 ，然後他必讓你們離開這裏。他放你們走的時候，一定會趕你們全都離開這裏。
EXOD|11|2|你要傳於百姓耳中，叫他們男的女的各向鄰舍索取金器銀器。」
EXOD|11|3|耶和華使 埃及 人看得起他的百姓 ，並且 摩西 在 埃及 地，在法老臣僕和百姓眼中看為偉大。
EXOD|11|4|摩西 說：「耶和華如此說：『約到半夜，我必出去走遍 埃及 。
EXOD|11|5|凡在 埃及 地，從坐寶座的法老到推磨 的婢女所生的長子，以及一切頭生的牲畜，都必死。
EXOD|11|6|埃及 全地必有大大的哀號，這將是空前絕後的。
EXOD|11|7|至於 以色列 人中，無論是人是牲畜，連狗也不敢向他們吠叫，使你們知道耶和華區別 埃及 和 以色列 。』
EXOD|11|8|你所有的這些臣僕都要下到我這裏，向我下拜說：『請你和跟從你的百姓都離開吧！』然後我才離開。」於是， 摩西 氣憤憤地離開法老出去了。
EXOD|11|9|耶和華對 摩西 說：「法老必不聽你們，為了要使我在 埃及 地多行奇事。」
EXOD|11|10|摩西 和 亞倫 在法老面前行了這一切奇事，但耶和華任憑法老的心剛硬，不讓 以色列 人離開他的地。
EXOD|12|1|耶和華在 埃及 地對 摩西 和 亞倫 說：
EXOD|12|2|「你們要以本月為正月，為一年之首。
EXOD|12|3|你們要吩咐 以色列 全會眾說：本月初十，各人要按著家庭 取羔羊，一家一隻羔羊。
EXOD|12|4|若一家的人太少，吃不了一隻羔羊，就要按照人數和隔壁的鄰舍共取一隻；你們要按每人的食量來估算羔羊。
EXOD|12|5|你們要從綿羊或山羊中取一隻無殘疾、一歲的公羔羊，
EXOD|12|6|要把牠留到本月十四日；那日黃昏的時候， 以色列 全會眾要把羔羊宰了。
EXOD|12|7|他們要取一些血，塗在他們吃羔羊的房屋兩邊的門框上和門楣上。
EXOD|12|8|當晚要吃羔羊的肉；要用火烤了，與無酵餅和苦菜一起吃。
EXOD|12|9|不可吃生的，或用水煮的，要把羔羊連頭帶腿和內臟用火烤了吃。
EXOD|12|10|一點也不可留到早晨；若有留到早晨的，要用火燒了。
EXOD|12|11|你們要這樣吃羔羊：腰間束帶，腳上穿鞋，手中拿杖，快快地吃。這是耶和華的逾越。
EXOD|12|12|因為那夜我要走遍 埃及 地，把 埃及 地一切頭生的，無論是人是牲畜，都擊殺了；我要對 埃及 所有的神明施行審判。我是耶和華。
EXOD|12|13|這血要在你們所住的房屋上作記號；我一見這血，就逾越你們。我擊打 埃及 地的時候，災殃必不臨到你們身上施行毀滅。」
EXOD|12|14|「你們要記念這日，世世代代守這日為耶和華的節日，作為你們永遠的定例。
EXOD|12|15|你們要吃無酵餅七日。第一日要把酵從你們各家中除去，因為從第一日到第七日，任何吃有酵之物的，必從 以色列 中剪除。
EXOD|12|16|第一日當有聖會，第七日也當有聖會。在這兩日，任何工作都不可做，只能預備各人的食物，這是惟一可做的工作。
EXOD|12|17|你們要守除酵節，因為我在這一日把你們的軍隊從 埃及 地領出來。所以，你們要世世代代守這日，立為永遠的定例。
EXOD|12|18|從正月十四日晚上，直到二十一日晚上，你們要吃無酵餅。
EXOD|12|19|在你們各家中，七日之內不可有酵，因為凡吃有酵之物的，無論是寄居的，是本地的，必從 以色列 的會中剪除。
EXOD|12|20|任何有酵的物，你們都不可吃；在你們一切的住處要吃無酵餅。」
EXOD|12|21|於是， 摩西 召了 以色列 的眾長老來，對他們說：「你們要為家人取羔羊，把逾越的羔羊宰了。
EXOD|12|22|要拿一把牛膝草，蘸盆裏的血，把盆裏的血塗在門楣上和兩邊的門框上。直到早晨你們誰也不可出自己家裏的門。
EXOD|12|23|因為耶和華要走遍 埃及 ，施行擊殺，他看見血在門楣上和兩邊的門框上，耶和華就必逾越那門，不讓滅命者進你們的家，施行擊殺。
EXOD|12|24|你們要守這命令，作為你們和你們子孫永遠的定例。
EXOD|12|25|日後，你們到了耶和華所應許賜給你們的那地，就要守這禮儀。
EXOD|12|26|你們的兒女對你們說：『這禮儀是甚麼意思呢？』
EXOD|12|27|你們就說：『這是獻給耶和華逾越節的祭物。當耶和華擊殺 埃及 人的時候，他逾越了 以色列 人在 埃及 的房屋，救了我們各家。』」於是百姓低頭敬拜。
EXOD|12|28|以色列 人就去做；他們照耶和華吩咐 摩西 和 亞倫 的去做了。
EXOD|12|29|到了半夜，耶和華把 埃及 地所有頭生的，就是從坐寶座的法老，到關在牢裏的人的長子，以及一切頭生的牲畜，盡都殺了。
EXOD|12|30|法老和他眾臣僕，以及所有的 埃及 人，都在夜間起來了。在 埃及 有大大的哀號，因為沒有一家不死人的。
EXOD|12|31|夜間，法老召了 摩西 和 亞倫 來，說：「起來！你們和 以色列 人，都離開我的百姓出去，照你們所說的，去事奉耶和華吧！
EXOD|12|32|照你們所說的，連羊群牛群也帶走，也為我祝福吧！」
EXOD|12|33|埃及 人催促百姓趕快離開那地，因為 埃及 人說：「我們都快死了。」
EXOD|12|34|百姓就拿著沒有發酵的生麵，把揉麵盆包在衣服中，扛在肩上。
EXOD|12|35|以色列 人照 摩西 的話去做，向 埃及 人索取金器、銀器和衣裳。
EXOD|12|36|耶和華使 埃及 人看得起他的百姓， 埃及 人就給了他們所要的。他們就掠奪了 埃及 人。
EXOD|12|37|以色列 人從 蘭塞 起程，往 疏割 去。除了小孩，步行的男人約有六十萬。
EXOD|12|38|又有許多不同族群的人，以及眾多的羊群牛群，和他們一同上去。
EXOD|12|39|他們用 埃及 帶出來的生麵烤成無酵餅。這生麵是沒有發酵的；因為他們被催促離開 埃及 ，不能耽延，就沒有為自己預備食物。
EXOD|12|40|以色列 人住在 埃及 共四百三十年。
EXOD|12|41|正滿四百三十年的那一天，耶和華的全軍從 埃及 地出來了。
EXOD|12|42|這是向耶和華守的夜，他領他們出 埃及 地；這是 以色列 眾人世世代代要向耶和華守的夜。
EXOD|12|43|耶和華對 摩西 和 亞倫 說：「逾越節的條例是這樣：外邦人不可吃這羔羊。
EXOD|12|44|但是你們用銀子買來，又受過割禮的奴僕可以吃。
EXOD|12|45|寄居的和雇工都不可吃。
EXOD|12|46|應當在一個屋子裏吃，不可把肉帶到屋外，骨頭一根也不可折斷。
EXOD|12|47|以色列 全會眾都要守這禮儀。
EXOD|12|48|若有外人寄居在你那裏，要向耶和華守逾越節，他所有的男子務要先受割禮，然後才可以當他是本地人，容許他守這禮儀。但未受割禮的都不可吃這羔羊。
EXOD|12|49|本地人和寄居在你們中間的外人當守同一個條例。」
EXOD|12|50|以色列 眾人就去做，他們照耶和華吩咐 摩西 和 亞倫 的去做了。
EXOD|12|51|正當那日，耶和華將 以色列 人按著他們的隊伍從 埃及 地領了出來。
EXOD|13|1|耶和華吩咐 摩西 說：
EXOD|13|2|「頭生的要分別為聖歸我； 以色列 中凡頭生的，無論是人是牲畜，都是我的。」
EXOD|13|3|摩西 對百姓說：「你們要記念從 埃及 為奴之家出來的這日，因為耶和華用大能的手將你們從這地領出來。有酵之物都不可吃。
EXOD|13|4|亞筆月的這一日你們走出來了。
EXOD|13|5|將來耶和華領你進 迦南 人、 赫 人、 亞摩利 人、 希未 人、 耶布斯 人之地，就是他向你祖宗起誓應許給你的那流奶與蜜之地，那時你要在這一個月守這禮儀。
EXOD|13|6|你要吃無酵餅七日，在第七日要向耶和華守節。
EXOD|13|7|這七日之內，要吃無酵餅；在你的全境內不可見有酵之物，也不可見酵母。
EXOD|13|8|當那日，你要告訴你的兒子說：『這樣做是因為耶和華在我出 埃及 的時候為我所做的事。』
EXOD|13|9|這要在你手上作記號，在你額上 作紀念，使耶和華的教導常在你口中，因為耶和華用大能的手將你從 埃及 領出來。
EXOD|13|10|所以你每年要按著日期守這條例。」
EXOD|13|11|「當耶和華照他向你和你祖宗所起的誓將你領進 迦南 人之地，把那地賜給你的時候，
EXOD|13|12|你要將一切頭生的獻給耶和華；你牲畜中頭生的，公的都歸耶和華。
EXOD|13|13|然而，凡頭生的驢，你要用羔羊贖回；若不贖牠，就要打斷牠的頸項。你兒子中的長子都要贖出來。
EXOD|13|14|日後，你的兒子問你說：『這是甚麼意思？』你就說：『耶和華用大能的手將我們從 埃及 為奴之家領出來。
EXOD|13|15|那時法老固執，不肯放我們走，耶和華就把 埃及 地所有頭生的，無論是人是牲畜，都殺了。因此，我把一切頭生的公的牲畜獻給耶和華為祭，卻將所有頭生的兒子贖出來。
EXOD|13|16|這要在你手上作記號，在你額上作經匣 ，因為耶和華用大能的手將我們從 埃及 領出來。』」
EXOD|13|17|法老放百姓走的時候， 非利士 人之地的路雖近，上帝卻不領他們從那裏走，因為上帝說：「恐怕百姓遇見戰爭就後悔，轉回 埃及 去。」
EXOD|13|18|上帝領百姓繞道而行，走曠野的路到 紅海 。 以色列 人出 埃及 地，都帶著兵器上去 。
EXOD|13|19|摩西 把 約瑟 的骸骨一起帶走；因為 約瑟 曾叫 以色列 人鄭重地起誓，對他們說：「上帝必定眷顧你們，你們要把我的骸骨從這裏一起帶上去。」
EXOD|13|20|他們從 疏割 起程，在曠野邊上的 以倘 安營。
EXOD|13|21|耶和華走在他們前面，日間用雲柱引領他們的路，夜間用火柱照亮他們，使他們日夜都可以行走。
EXOD|13|22|日間的雲柱，夜間的火柱，總不離開百姓的面前。
EXOD|14|1|耶和華吩咐 摩西 說：
EXOD|14|2|「你吩咐 以色列 人轉回，要在 比‧哈希錄 前面， 密奪 和海的中間， 巴力‧洗分 的前面安營。你們要在對面，靠近海邊安營。
EXOD|14|3|以色列 人這樣做，法老必說：『他們在此地迷了路，曠野把他們困住了。』
EXOD|14|4|我要任憑法老的心剛硬，他要追趕他們。我必在法老和他全軍身上得榮耀， 埃及 人就知道我是耶和華。」於是 以色列 人照樣做了。
EXOD|14|5|有人報告 埃及 王說：「百姓逃跑了！」法老和他的臣僕對百姓改變了心意，說：「我們放 以色列 人走，不再服事我們，我們怎麼會做這種事呢？」
EXOD|14|6|法老就預備戰車，帶領他的軍兵同去，
EXOD|14|7|他帶了六百輛特選的戰車和 埃及 所有的戰車，每輛都有軍官。
EXOD|14|8|耶和華任憑 埃及 王法老的心剛硬，他就追趕 以色列 人； 以色列 人卻抬起頭 來出去了。
EXOD|14|9|埃及 人追趕他們，法老一切的馬匹、戰車、戰車長，與軍兵就在海邊上，靠近 比‧哈希錄 ，在 巴力‧洗分 的前面，在他們安營的地方追上了。
EXOD|14|10|法老逼近的時候， 以色列 人舉目，看哪， 埃及 人追來了，就非常懼怕， 以色列 人向耶和華哀求。
EXOD|14|11|他們對 摩西 說：「難道 埃及 沒有墳地，你要把我們帶來死在曠野嗎？你為甚麼這樣待我們，將我們從 埃及 領出來呢？
EXOD|14|12|我們在 埃及 豈沒有對你說過，不要攪擾我們，讓我們服事 埃及 人嗎？因為服事 埃及 人總比死在曠野好。」
EXOD|14|13|摩西 對百姓說：「不要怕，要站穩，看耶和華今天向你們所要施行的拯救，因為你們今天所看見的 埃及 人必永遠不再看見了。
EXOD|14|14|耶和華必為你們爭戰，你們要安靜！」
EXOD|14|15|耶和華對 摩西 說：「你為甚麼向我哀求呢？你吩咐 以色列 人往前走。
EXOD|14|16|你舉手向海伸杖，把水分開。 以色列 人要下到海中，走在乾地上。
EXOD|14|17|看哪，我要任憑 埃及 人的心剛硬，他們就跟著下去。我要在法老和他的全軍、戰車、戰車長身上得榮耀。
EXOD|14|18|我在法老和他的戰車、戰車長身上得榮耀的時候， 埃及 人就知道我是耶和華。」
EXOD|14|19|在 以色列 營前行走的上帝的使者移動，走到他們後面；雲也從他們的前面移動，站在他們後面。
EXOD|14|20|它來到 埃及 營和 以色列 營的中間：一邊有雲和黑暗，另一邊它照亮夜晚，整夜彼此不得接近。
EXOD|14|21|摩西 向海伸手，耶和華就用強勁的東風，使海水在一夜間退去，海就成了乾地；水分開了。
EXOD|14|22|以色列 人下到海中，走在乾地上，水在他們左右成了牆壁。
EXOD|14|23|埃及 人追趕他們，法老一切的馬匹、戰車和戰車長都跟著下到海中。
EXOD|14|24|破曉時分，耶和華從雲柱、火柱中瞭望 埃及 的軍兵，使 埃及 的軍兵混亂。
EXOD|14|25|他使他們的車輪脫落 ，難以前行， 埃及 人說：「我們從 以色列 人面前逃跑吧！因耶和華為他們作戰，攻擊 埃及 了。」
EXOD|14|26|耶和華對 摩西 說：「你要向海伸手，使水回流到 埃及 人，他們的戰車和戰車長身上。」
EXOD|14|27|摩西 就向海伸手，到了天亮的時候，海恢復原狀。 埃及 人逃避水的時候，耶和華把他們推入海中。
EXOD|14|28|海水回流，淹沒了戰車和戰車長，以及那些跟著 以色列 人下到海中的法老全軍，連一個也沒有剩下。
EXOD|14|29|以色列 人卻在海中走乾地，水在他們的左右成了牆壁。
EXOD|14|30|那一日，耶和華拯救 以色列 脫離 埃及 人的手。 以色列 人看見 埃及 人死在海邊。
EXOD|14|31|以色列 人看見耶和華向 埃及 人所施展的大能，百姓就敬畏耶和華，並且信服耶和華和他的僕人 摩西 。
EXOD|15|1|那時， 摩西 和 以色列 人向耶和華唱這歌，說： 「我要向耶和華歌唱，因他大大得勝， 將馬和騎馬的投在海中。
EXOD|15|2|耶和華是我的力量，是我的詩歌， 他也成了我的拯救。 這是我的上帝，我要讚美他； 我父親的上帝，我要尊崇他。
EXOD|15|3|耶和華是戰士； 耶和華是他的名。
EXOD|15|4|「法老的戰車、軍兵，他已拋在海中； 法老精選的軍官都沉於 紅海 。
EXOD|15|5|深水淹沒他們； 他們好像石頭墜到深處。
EXOD|15|6|耶和華啊，你的右手施展能力，大顯榮耀； 耶和華啊，你的右手摔碎仇敵。
EXOD|15|7|你大發威嚴，摧毀了你的敵人； 你發出烈怒，吞滅他們如同碎秸。
EXOD|15|8|因你鼻中的氣，水就聚成堆， 大水豎立如壘， 海的中心深水凝結。
EXOD|15|9|仇敵說：『我要追趕，我要追上， 我要分擄物，在他們身上滿足我的心願， 我要拔刀，親手毀滅他們。』
EXOD|15|10|你用風一吹，海水就淹沒他們； 他們像鉛沉在大水之中。
EXOD|15|11|「耶和華啊，眾神明中，誰能像你？ 誰能像你，至聖至榮， 可頌可畏，施行奇事！
EXOD|15|12|你伸出右手， 地就吞滅他們。
EXOD|15|13|「你以慈愛引領你所救贖的百姓； 你以能力引導他們到你的聖所。
EXOD|15|14|萬民聽見就戰抖； 疼痛抓住 非利士 的居民。
EXOD|15|15|那時， 以東 的族長驚惶， 摩押 的英雄被戰兢抓住， 迦南 所有的居民都融化。
EXOD|15|16|驚駭恐懼臨到他們； 耶和華啊，因你膀臂的大能， 他們如石頭寂靜不動， 等候你百姓過去， 等候你所贖的百姓過去。
EXOD|15|17|你要將他們領進去，栽在你產業的山上， 耶和華啊，就是你為自己所造的住處， 主啊，就是你手所建立的聖所。
EXOD|15|18|耶和華必作王，直到永永遠遠！」
EXOD|15|19|法老的馬匹、戰車和戰車長下到海中，耶和華使海水回流到他們身上； 以色列 人卻走在海中的乾地上。
EXOD|15|20|那時， 米利暗 女先知， 亞倫 的姊姊，手裏拿著鈴鼓；眾婦女也跟她出去打鼓跳舞。
EXOD|15|21|米利暗 回應他們： 「你們要歌頌耶和華，因他大大得勝， 將馬和騎馬的投在海中。」
EXOD|15|22|摩西 領 以色列 人從 紅海 起程，到了 書珥 的曠野，在曠野走了三天，找不到水。
EXOD|15|23|到了 瑪拉 ，他們不能喝 瑪拉 的水，因為水是苦的；所以那地名叫 瑪拉 。
EXOD|15|24|百姓就向 摩西 發怨言，說：「我們喝甚麼呢？」
EXOD|15|25|摩西 呼求耶和華，耶和華指示他一棵樹 。他把樹丟在水裏，水就變甜了。 耶和華在那裏為他們定了律例、典章，在那裏考驗他們。
EXOD|15|26|他說：「你若留心聽從耶和華－你上帝的話，行我眼中看為正的事，側耳聽我的誡令，遵守我一切的律例，我就不將所加於 埃及 人的疾病加在你身上，因為我是醫治你的耶和華。」
EXOD|15|27|他們到了 以琳 ，在那裏有十二股水泉，七十棵棕樹；他們就在那裏的水邊安營。
EXOD|16|1|以色列 全會眾從 以琳 起程，在出 埃及 之後第二個月十五日到了 以琳 和 西奈 中間， 汛 的曠野。
EXOD|16|2|以色列 全會眾在曠野向 摩西 和 亞倫 發怨言。
EXOD|16|3|以色列 人對他們說：「我們寧願在 埃及 地死在耶和華手中！那時我們坐在肉鍋旁，吃餅得飽。你們卻將我們領出來，到這曠野，要叫這全會眾都餓死啊！」
EXOD|16|4|耶和華對 摩西 說：「看哪，我要從天降食物給你們。百姓可以出去，每天收集當天的分量。這樣，我就可以考驗他們是否遵行我的指示。
EXOD|16|5|到第六天，他們預備食物，所收集的分量要比每天所收的多一倍。」
EXOD|16|6|摩西 和 亞倫 對 以色列 眾人說：「到了晚上，你們就知道是耶和華將你們從 埃及 地領出來的。
EXOD|16|7|早晨，你們要看見耶和華的榮耀，因為耶和華聽見你們向他所發的怨言了。我們算甚麼，你們竟然向我們發怨言呢？」
EXOD|16|8|摩西 又說：「耶和華晚上必給你們肉吃，早晨必給你們食物得飽，因為耶和華已經聽見你們向他所發的怨言。我們算甚麼呢？你們的怨言不是向我們發的，而是向耶和華發的。」
EXOD|16|9|摩西 對 亞倫 說：「你對 以色列 全會眾說：『你們來到耶和華面前，因為他已經聽見你們的怨言了。』」
EXOD|16|10|亞倫 正對 以色列 全會眾說話的時候，他們轉向曠野，看哪，耶和華的榮光在雲中顯現。
EXOD|16|11|耶和華吩咐 摩西 說：
EXOD|16|12|「我已經聽見 以色列 人的怨言了。你要對他們說：『到黃昏的時候 ，你們要吃肉，早晨也必有食物得飽。你們就知道我是耶和華－你們的上帝。』」
EXOD|16|13|到了晚上，有鵪鶉上來，遮滿營地；早晨，營地周圍有一層露水。
EXOD|16|14|那一層露水蒸發之後，看哪，曠野的表面出現了小圓物，好像地上的薄霜一樣。
EXOD|16|15|以色列 人看見了，不知道是甚麼，就彼此說：「這是甚麼？ 」 摩西 對他們說：「這是耶和華給你們吃的食物。
EXOD|16|16|耶和華所吩咐的是這樣：『你們每個人要按自己的食量收集，各人要為帳棚裏的人收集，按照人口數每個人一俄梅珥。』」
EXOD|16|17|以色列 人就照樣去做；有的收多，有的收少。
EXOD|16|18|用俄梅珥量一量，多收的沒有餘，少收的也沒有缺；各人都按著自己的食量收集。
EXOD|16|19|摩西 對他們說：「任何人都不可以把所收的留到早晨。」
EXOD|16|20|然而他們不聽從 摩西 ，當中有人把食物留到早晨，食物就生蟲發臭了。 摩西 就向他們發怒。
EXOD|16|21|他們每日早晨按著各人的食量收集；太陽一發熱，食物就融化了。
EXOD|16|22|到第六天，他們收集了雙倍的食物，每個人二俄梅珥。會眾的官長來告訴 摩西 ，
EXOD|16|23|摩西 對他們說：「耶和華吩咐：『明天是安息日，是向耶和華守的聖安息日。你們要烤的就烤，要煮的就煮，所剩下的都留到早晨。』」
EXOD|16|24|他們就照 摩西 的吩咐把剩下的留到早晨，這些食物既不發臭，裏頭也沒有生蟲。
EXOD|16|25|摩西 說：「你們今天就吃這些吧！因為今天是向耶和華守的安息日，你們在野外必找不著食物了。
EXOD|16|26|六天可以收集，第七天是安息日，這一天甚麼也沒有了。」
EXOD|16|27|第七天，百姓中有人出去收，甚麼也找不著。
EXOD|16|28|耶和華對 摩西 說：「你們不肯遵守我的誡令和教導，要到幾時呢？
EXOD|16|29|你們看，耶和華既然將安息日賜給你們，所以第六天他就賜給你們兩天的食物，第七天各人都要留在自己的地方，不許任何人從這裏出去。」
EXOD|16|30|於是百姓在第七天安息了。
EXOD|16|31|以色列 家給這食物取名叫嗎哪，它的樣子像芫荽子，顏色是白的，吃起來像和蜜的薄餅。
EXOD|16|32|摩西 說：「耶和華所吩咐的是這樣：『要裝滿一俄梅珥的嗎哪留給你們的後代，使他們可以看見我領你們出 埃及 地的時候，在曠野所給你們吃的食物。』」
EXOD|16|33|摩西 對 亞倫 說：「你拿一個罐子，裝滿一俄梅珥的嗎哪，存在耶和華面前，留給你們的後代。」
EXOD|16|34|耶和華怎麼吩咐 摩西 ， 亞倫 就照樣做，把嗎哪存留作見證 。
EXOD|16|35|以色列 人吃嗎哪共四十年，直到進入有人居住的地方；他們吃嗎哪，直到 迦南 地的邊境。
EXOD|16|36|一俄梅珥是一伊法的十分之一。
EXOD|17|1|以色列 全會眾遵照耶和華的吩咐，從 汛 的曠野一段一段地往前行。他們在 利非訂 安營，但百姓沒有水喝。
EXOD|17|2|百姓就與 摩西 爭鬧，說：「給我們水喝吧！」 摩西 對他們說：「你們為甚麼與我爭鬧呢？你們為甚麼試探耶和華呢？」
EXOD|17|3|百姓在那裏口渴要喝水，就向 摩西 發怨言，說：「你為甚麼把我們從 埃及 領出來，使我們和我們的兒女，以及牲畜都渴死呢？」
EXOD|17|4|摩西 就呼求耶和華說：「我要怎樣對待這百姓呢？他們差一點就要拿石頭打死我了。」
EXOD|17|5|耶和華對 摩西 說：「你帶著 以色列 的幾個長老，走在百姓前面，手裏拿著你先前擊打 尼羅河 的杖，去吧！
EXOD|17|6|看哪，我要在 何烈 的磐石那裏，站在你面前。你要擊打磐石，水就會從磐石流出來，給百姓喝。」 摩西 就在 以色列 的長老眼前這樣做了。
EXOD|17|7|他給那地方起名叫 瑪撒 ，又叫 米利巴 ，因為 以色列 人在那裏爭鬧，並且試探耶和華，說：「耶和華是否在我們中間呢？」
EXOD|17|8|那時， 亞瑪力 來到 利非訂 ，和 以色列 爭戰。
EXOD|17|9|摩西 對 約書亞 說：「你為我們選出人來，出去和 亞瑪力 爭戰。明天我要站在山頂上，手裏拿著上帝的杖。」
EXOD|17|10|於是， 約書亞 照著 摩西 對他所說的話去做，和 亞瑪力 爭戰。 摩西 、 亞倫 和 戶珥 都上了山頂。
EXOD|17|11|摩西 何時舉手， 以色列 就得勝；何時垂手， 亞瑪力 就得勝。
EXOD|17|12|但 摩西 的雙手沉重，他們就搬一塊石頭來放在他下面，他就坐在上面。 亞倫 與 戶珥 扶著他的手，一個在這邊，一個在那邊，他的手就穩住，直到日落。
EXOD|17|13|約書亞 用刀打敗了 亞瑪力 和他的百姓。
EXOD|17|14|耶和華對 摩西 說：「你要把這事記錄在書上作紀念，又念給 約書亞 聽：我要把 亞瑪力 的名字從天下全然塗去。」
EXOD|17|15|摩西 築了一座壇，起名叫「耶和華尼西 」。
EXOD|17|16|他說：「我指著耶和華的寶座發誓 ，耶和華必世世代代和 亞瑪力 爭戰。」
EXOD|18|1|摩西 的岳父， 米甸 祭司 葉特羅 ，聽見上帝為 摩西 和為他百姓 以色列 所行的一切事，就是耶和華將 以色列 從 埃及 領了出來。
EXOD|18|2|摩西 的岳父 葉特羅 帶著 西坡拉 ，就是 摩西 先前送回家的妻子，
EXOD|18|3|又帶著她的兩個兒子：一個名叫 革舜 ，因為 摩西 說：「我在外地作了寄居者」；
EXOD|18|4|另一個名叫 以利以謝 ，因為他說：「我父親的上帝幫助我，救我脫離法老的刀。」
EXOD|18|5|摩西 的岳父 葉特羅 帶著 摩西 的妻子和兩個兒子來到上帝的山，就是 摩西 在曠野安營的地方。
EXOD|18|6|他對 摩西 說：「我是 你岳父 葉特羅 ，帶著你的妻子和兩個兒子來到你這裏。」
EXOD|18|7|摩西 迎接他的岳父，向他下拜，親他，彼此問安，然後進入帳棚。
EXOD|18|8|摩西 將耶和華為 以色列 的緣故向法老和 埃及 人所行的一切事，他們在路上遭遇的一切艱難，以及耶和華怎樣搭救他們，都述說給他的岳父聽。
EXOD|18|9|葉特羅 因耶和華待 以色列 的一切恩惠，就是拯救他們脫離 埃及 人的手，就非常喜樂。
EXOD|18|10|葉特羅 說：「耶和華是應當稱頌的，他救了你們脫離 埃及 人和法老的手，將這百姓從 埃及 人的手裏救出來 。
EXOD|18|11|現在，從 埃及 人狂傲地對待 以色列 人這件事上，我知道耶和華比萬神更大。」
EXOD|18|12|摩西 的岳父 葉特羅 把燔祭和祭物獻給上帝。 亞倫 和 以色列 的眾長老都來了，與 摩西 的岳父在上帝面前吃飯。
EXOD|18|13|第二天， 摩西 坐著審判百姓，百姓從早到晚站在 摩西 的旁邊。
EXOD|18|14|摩西 的岳父看見他為百姓所做的一切事，就說：「你為百姓所做的，這是甚麼事呢？你為甚麼獨自一人坐著，而眾百姓從早到晚都站在你旁邊呢？」
EXOD|18|15|摩西 對岳父說：「這是因為百姓到我這裏來求問上帝。
EXOD|18|16|他們有事的時候，就到我這裏來，我就在雙方之間作判決；我又叫他們知道上帝的律例和法度。」
EXOD|18|17|摩西 的岳父對他說：「你這樣做不好。
EXOD|18|18|你和這些與你在一起的百姓都必疲憊，因為這事太重，你獨自一人做不了。
EXOD|18|19|現在，聽我的話，我給你出個主意，願上帝與你同在。你要代替百姓到上帝面前，將事件帶到上帝那裏，
EXOD|18|20|又要用律例和法度警戒他們，指示他們當行的道，當做的事。
EXOD|18|21|你也要從百姓中選出有才能的人，敬畏上帝、誠實可靠、恨惡不義之財的人，派他們作千夫長、百夫長、五十夫長、十夫長來管理百姓。
EXOD|18|22|他們要隨時審判百姓；重大的事要送到你這裏，小事就由他們自行判決。這樣，你就可以輕省一些，他們可以與你分擔。
EXOD|18|23|你若這樣做，上帝也這樣吩咐你，你就能承受得住，眾百姓也可以和睦地回到自己的地方。」
EXOD|18|24|摩西 聽了他岳父的話，照著他所說的一切去做。
EXOD|18|25|摩西 從 以色列 人中選出有才能的人，立他們為百姓的領袖，作千夫長、百夫長、五十夫長、十夫長。
EXOD|18|26|他們隨時審判百姓：難斷的事就送到 摩西 那裏，各樣小事就由他們自行判決。
EXOD|18|27|於是， 摩西 給他的岳父送行，他就回到本地去了。
EXOD|19|1|以色列 人出 埃及 地以後，第三個月的初一，就在那一天他們來到了 西奈 的曠野。
EXOD|19|2|他們從 利非訂 起程，來到 西奈 的曠野，在那裏的山下安營。
EXOD|19|3|摩西 到上帝那裏，耶和華從山上呼喚他說：「你要這樣告訴 雅各 家，對 以色列 人說：
EXOD|19|4|『我向 埃及 人所行的事，你們都看見了， 我如鷹將你們背在翅膀上，帶你們來歸我。
EXOD|19|5|如今你們若真的聽從我的話，遵守我的約，就要在萬民中作屬我的子民 ，因為全地都是我的。
EXOD|19|6|你們要歸我作祭司的國度，為神聖的國民。』這些話你要告訴 以色列 人。」
EXOD|19|7|摩西 去召了百姓中的長老來，將耶和華吩咐他的話當面告訴他們。
EXOD|19|8|百姓都同聲回答：「凡耶和華所說的，我們一定遵行。」 摩西 就將百姓的話回覆耶和華。
EXOD|19|9|耶和華對 摩西 說：「看哪，我要在密雲中臨到你那裏，叫百姓在我與你說話的時候可以聽見，就可以永遠相信你了。」於是， 摩西 將百姓的話稟告耶和華。
EXOD|19|10|耶和華對 摩西 說：「你往百姓那裏去，使他們今天明天分別為聖，又叫他們洗衣服。
EXOD|19|11|第三天要預備好，因為第三天耶和華要在眾百姓眼前降臨在 西奈山 。
EXOD|19|12|你要在山的周圍給百姓劃定界限，說：『你們當謹慎，不可上山去，也不可摸山的邊界。凡摸這山的，必被處死。
EXOD|19|13|不可用手碰他，要用石頭打死，或射死；無論是人是牲畜，都不可活。』到角聲拉長的時候，他們才可到山腳來。」
EXOD|19|14|摩西 下山到百姓那裏去，使他們分別為聖，他們就洗衣服。
EXOD|19|15|他對百姓說：「第三天要預備好；不可親近女人。」
EXOD|19|16|到了第三天早晨，山上有雷轟、閃電和密雲，並且角聲非常響亮，營中的百姓盡都戰抖。
EXOD|19|17|摩西 率領百姓出營迎見上帝，都站在山下。
EXOD|19|18|西奈山 全山冒煙，因為耶和華在火中降臨山上。山的煙霧上騰，彷彿燒窯，整座山劇烈震動。
EXOD|19|19|角聲越來越響， 摩西 說話，上帝以聲音回答他。
EXOD|19|20|耶和華降臨在 西奈山 頂上，耶和華召 摩西 上山頂， 摩西 就上去了。
EXOD|19|21|耶和華對 摩西 說：「你下去警告百姓，免得他們闖過來看耶和華，就會有許多人死亡。
EXOD|19|22|那些親近耶和華的祭司也要把自己分別為聖，免得耶和華忽然出來擊殺他們。」
EXOD|19|23|摩西 對耶和華說：「百姓不能上 西奈山 ，因為你已經警告我們說：『要在山的周圍劃定界限，使山成聖。』」
EXOD|19|24|耶和華對他說：「下去吧，你要和 亞倫 一起上來；只是祭司和百姓不可闖上來到耶和華這裏，免得耶和華忽然出來擊殺他們。」
EXOD|19|25|於是， 摩西 下到百姓那裏告訴他們。
EXOD|20|1|上帝吩咐這一切的話，說：
EXOD|20|2|「我是耶和華－你的上帝，曾將你從 埃及 地為奴之家領出來。
EXOD|20|3|「除了我以外，你不可有別的神。
EXOD|20|4|「不可為自己雕刻偶像，也不可做甚麼形像，彷彿上天、下地和地底下水中的百物。
EXOD|20|5|不可跪拜那些像，也不可事奉它們，因為我耶和華─你的上帝是忌邪 的上帝。恨我的，我必懲罰他們的罪，自父及子，直到三、四代；
EXOD|20|6|愛我，守我誡命的，我必向他們施慈愛，直到千代。
EXOD|20|7|「不可妄稱耶和華－你上帝的名，因為妄稱耶和華名的，耶和華必不以他為無罪。
EXOD|20|8|「當記念安息日，守為聖日。
EXOD|20|9|六日要勞碌做你一切的工，
EXOD|20|10|但第七日是向耶和華─你的上帝當守的安息日。這一日你和你的兒女、奴僕、婢女、牲畜，以及你城裏寄居的客旅，都不可做任何的工。
EXOD|20|11|因為六日之內，耶和華造天、地、海和其中的萬物，第七日就安息了；所以耶和華賜福與安息日，定為聖日。
EXOD|20|12|「當孝敬父母，使你的日子在耶和華－你上帝所賜你的地上得以長久。
EXOD|20|13|「不可殺人。
EXOD|20|14|「不可姦淫。
EXOD|20|15|「不可偷盜。
EXOD|20|16|「不可做假見證陷害你的鄰舍。
EXOD|20|17|「不可貪戀你鄰舍的房屋；不可貪戀你鄰舍的妻子、奴僕、婢女、牛驢，以及他一切所有的。」
EXOD|20|18|眾百姓見雷轟、閃電、角聲、山上冒煙，百姓看見 就都戰抖，遠遠站著。
EXOD|20|19|他們對 摩西 說：「請你向我們說話，我們必聽；不要讓上帝向我們說話，免得我們死亡。」
EXOD|20|20|摩西 對百姓說：「不要害怕；因為上帝降臨是要考驗你們，要你們敬畏他，不致犯罪。」
EXOD|20|21|於是百姓遠遠站著，但 摩西 卻挨近上帝所在的幽暗中。
EXOD|20|22|耶和華對 摩西 說：「你要向 以色列 人這樣說：『你們親自看見我從天上向你們說話了。
EXOD|20|23|你們不可為我製造偶像，不可為自己造任何金銀的神像。
EXOD|20|24|你要為我築一座土壇，在上面獻牛羊為燔祭和平安祭。凡在我叫你記念我名的地方，我必到那裏賜福給你。
EXOD|20|25|你若為我築一座石壇，不可用鑿過的石頭，因為你在石頭上動了工具，就使壇污穢了。
EXOD|20|26|你不可用臺階上我的壇，免得露出你的下體來。』」
EXOD|21|1|「你在百姓面前所要立的典章是這樣：
EXOD|21|2|「你若買 希伯來 人作奴僕，他服事你六年，第七年他可以自由，白白地離去。
EXOD|21|3|他若單身來就可以單身去；他若是有妻子的，他的妻子可以同他離去。
EXOD|21|4|若他主人給他娶了妻，妻子為他生了兒子或女兒，妻子和兒女要歸主人，他要獨自離去。
EXOD|21|5|倘若奴僕聲明：『我愛我的主人和我的妻子兒女，不願意自由離去。』
EXOD|21|6|他的主人就要帶他到審判官 前，再帶他到門或門框那裏，用錐子穿他的耳朵，他就要永遠服事主人。
EXOD|21|7|「人若賣女兒作婢女，婢女不可像男的奴僕那樣離去。
EXOD|21|8|主人若選定她歸自己，後來看不順眼，就要允許她贖身；主人既然對她失信，就沒有權柄把她賣給外邦人。
EXOD|21|9|主人若選定她給自己的兒子，就當照女兒的規矩對待她。
EXOD|21|10|若另娶一個，她的飲食、衣服和房事不可減少。
EXOD|21|11|若不向她行這三樣，她就可以白白離去，不必付贖金。」
EXOD|21|12|「打人致死的，必被處死。
EXOD|21|13|他若不是出於預謀 ，而是上帝交在他手中，我就設立一個地方，讓他可以逃到那裏。
EXOD|21|14|人若蓄意用詭計殺了他的鄰舍，就是逃到我的壇那裏，也當把他捉去處死。
EXOD|21|15|「打父母的，必被處死。
EXOD|21|16|「誘拐人口的，無論是把人賣了，或是扣留在他手中，必被處死。
EXOD|21|17|「咒罵父母的，必被處死。
EXOD|21|18|「人若彼此爭吵，一個用石頭或拳頭打另一個，被打的人沒有死去，卻要躺臥在床，
EXOD|21|19|若他還能起來扶杖行走，那打他的可免處刑，卻要賠償他不能工作的損失，並要把他完全醫好。
EXOD|21|20|「人若用棍子打奴僕或婢女，當場死在他的手下，他必受報應。
EXOD|21|21|若能撐過一兩天，主人就不必受懲罰，因為那是他的財產。
EXOD|21|22|「人若彼此打鬥，傷害有孕的婦人，以致胎兒掉了出來，隨後卻無別的傷害，那傷害她的人，總要按婦人的丈夫所提出的，照審判官所裁定的賠償。
EXOD|21|23|若有別的傷害，就要以命抵命，
EXOD|21|24|以眼還眼，以牙還牙，以手還手，以腳還腳，
EXOD|21|25|以灼傷還灼傷，以損傷還損傷，以鞭打還鞭打。
EXOD|21|26|「人若打奴僕或婢女的眼睛，毀了一隻，就要因他的眼讓他自由離去。
EXOD|21|27|若打掉了奴僕或婢女的一顆牙，就要因他的牙讓他自由離去。」
EXOD|21|28|「牛若牴死男人或女人，總要用石頭打死那牛，卻不可吃牠的肉；牛的主人可免處刑。
EXOD|21|29|倘若那牛向來是牴人的，牛的主人雖然受過警告，仍不把牠拴好，以致把男人或女人牴死，牛要用石頭打死，主人也要被處死。
EXOD|21|30|若罰他付贖命的賠款，他就要照所罰的數目贖他的命。
EXOD|21|31|牛若牴了男孩或女孩，也要照這條例處理。
EXOD|21|32|牛若牴了奴僕或婢女，就要把三十舍客勒銀子給他的主人，牛要用石頭打死。
EXOD|21|33|「人若敞開井口，或挖井不蓋住它，有牛或驢掉進井裏，
EXOD|21|34|井的主人要拿錢賠償牲畜的主人，死牲畜要歸自己。
EXOD|21|35|「人的牛若牴死鄰舍的牛，他們就要賣了那活牛，平分價錢；也要平分死牛。
EXOD|21|36|若這牛向來是以好牴人出名的，主人竟不把牛拴好，他必要以牛賠牛，死牛卻歸自己。」
EXOD|22|1|「人若偷牛或羊，無論是宰了或賣了，他就要以五牛賠一牛， 四羊賠一羊。
EXOD|22|2|賊挖洞，若被發現而被打死，打的人沒有流血的罪。
EXOD|22|3|若太陽已經出來，打的人就有流血的罪。賊總要賠償，若他一無所有，就要被賣來還他所偷的東西。
EXOD|22|4|若發現他所偷的，無論是牛、驢，或羊，在他手中還活著，他就要加倍賠償。
EXOD|22|5|「人若在田間或葡萄園裏牧放牲畜，任憑牲畜上別人田裏去吃 ，他就要拿自己田間和葡萄園裏上好的賠償。
EXOD|22|6|「若火冒出，延燒到荊棘，以致將堆積的禾捆，直立的莊稼，或田地，都燒盡了，那點火的必要賠償。
EXOD|22|7|「人若將銀錢或物件託鄰舍保管，東西從這人的家中被偷去，若找到了賊，賊要加倍賠償；
EXOD|22|8|若找不到賊，這家的主人就要到審判官 那裏，聲明 自己沒有伸手拿鄰舍的物件。
EXOD|22|9|「關於任何侵害的案件，無論是為牛、驢、羊、衣服，或任何失物，有一人說：『這是我的』，雙方就要將案件帶到審判官面前，審判官定誰有罪，誰就要加倍賠償給他的鄰舍。
EXOD|22|10|「人將驢、牛、羊，或別的牲畜託鄰舍看管，若牲畜死亡，受了傷，或被搶走，無人看見，
EXOD|22|11|雙方要在耶和華前起誓，受託人要表明自己沒有伸手拿鄰舍的東西，原主要接受誓言，受託人不必賠償。
EXOD|22|12|牲畜若從受託人那裏被偷去，他就要賠償原主；
EXOD|22|13|若被野獸撕碎，受託人要帶回來作證據，被撕碎的就不必賠償。
EXOD|22|14|「人若向鄰舍借牲畜 ，所借的或傷或死，原主沒有在場，借的人總要賠償。
EXOD|22|15|若原主在場，借的人不必賠償；若是租用的，只要付租金 。」
EXOD|22|16|「人若引誘沒有訂婚的處女，與她同寢，他就必須交出聘禮，娶她為妻。
EXOD|22|17|若女子的父親堅決不將女子給他，他就要按著處女的聘禮交出錢來。
EXOD|22|18|「行邪術的女人，不可讓她存活。
EXOD|22|19|「凡與獸交合的，必被處死。
EXOD|22|20|「向別神獻祭，不單單獻給耶和華的，那人必要滅絕。
EXOD|22|21|「不可虧待寄居的，也不可欺壓他，因為你們在 埃及 地也作過寄居的。
EXOD|22|22|不可苛待寡婦和孤兒；
EXOD|22|23|若你確實苛待他，他向我苦苦哀求，我一定會聽他的呼求，
EXOD|22|24|並要發烈怒，用刀殺你們，使你們的妻子成為寡婦，兒女成為孤兒。
EXOD|22|25|「我的子民中有困苦人在你那裏，你若借錢給他，不可如放債的向他取利息。
EXOD|22|26|你果真拿了鄰舍的外衣作抵押，也要在日落前還給他；
EXOD|22|27|因為他只有這一件用來作被子，是他蔽體的衣服。他還可以拿甚麼睡覺呢？當他哀求我，我就應允，因為我是有恩惠的。
EXOD|22|28|「不可毀謗上帝；也不可詛咒你百姓的領袖。
EXOD|22|29|「不可遲延獻你的莊稼、酒和油 。 「要將你頭生的兒子歸給我。
EXOD|22|30|你的牛羊也要照樣做：七天當跟著牠母親，第八天你要把牠歸給我。
EXOD|22|31|「你們要分別為聖歸給我。因此，田間被野獸撕裂的肉，你們不可吃，要把它丟給狗。」
EXOD|23|1|「不可散佈謠言；不可與惡人連手作惡意的見證。
EXOD|23|2|不可附和群眾作惡；不可在訴訟中附和群眾歪曲公正，作歪曲的見證；
EXOD|23|3|也不可在訴訟中偏袒貧寒人。
EXOD|23|4|「若遇見你仇敵的牛或驢迷了路，務必牽回來交給他。
EXOD|23|5|若看見恨你的人的驢被壓在重馱之下，不可走開，務要和他一同卸下驢的重馱。
EXOD|23|6|「不可在貧窮人的訴訟中屈枉正直。
EXOD|23|7|當遠離誣告的事。不可殺害無辜和義人，因我必不以惡人為義。
EXOD|23|8|不可接受賄賂，因為賄賂能使明眼人變瞎，又能曲解義人的證詞。
EXOD|23|9|「不可欺壓寄居的，因為你們在 埃及 地作過寄居的，知道寄居者的心情。」
EXOD|23|10|「六年你要耕種田地，收集地的出產。
EXOD|23|11|只是第七年你要讓地歇息，不耕不種，使你百姓中的貧窮人有吃的；他們吃剩的，野獸可以吃。你的葡萄園和橄欖園也要照樣辦理。
EXOD|23|12|「六日你要做工，第七日要安息，使牛、驢可以歇息，也讓你使女的兒子和寄居的可以恢復精力。
EXOD|23|13|「凡我對你們說的話，你們都要謹守。別神的名，你不可提，也不可用口說給人聽。」
EXOD|23|14|「一年三次，你要向我守節。
EXOD|23|15|你要守除酵節，照我所吩咐你的，在亞筆月內所定的日期吃無酵餅七天，因為你是在這月離開了 埃及 。誰也不可空手來朝見我。
EXOD|23|16|你要守收割節，收田間所種、勞碌所得初熟之物。你年底收藏田間勞碌所得時，要守收藏節。
EXOD|23|17|所有的男丁都要一年三次朝見主耶和華。
EXOD|23|18|「不可將我祭牲的血和有酵之物一同獻上，也不可將我節期中祭牲的脂肪留到早晨。
EXOD|23|19|「要把地裏最好的初熟之物帶到耶和華－你上帝的殿中。 「不可用母山羊的奶來煮牠的小山羊。」
EXOD|23|20|「看哪，我要差遣使者在你前面，在路上保護你，領你到我所預備的地方。
EXOD|23|21|你們要在他面前謹慎，聽從他的話。不可抗拒 他，否則他必不赦免你們的過犯，因為我的名在他身上。
EXOD|23|22|「你若真的聽從他的話，照我一切所說的去做，我就以你的仇敵為仇敵，以你的敵人為敵人。
EXOD|23|23|「我的使者要走在你前面，領你到 亞摩利 人、 赫 人、 比利洗 人、 迦南 人、 希未 人、 耶布斯 人那裏，我必將他們除滅。
EXOD|23|24|你不可跪拜事奉他們的神明，也不可隨從他們的習俗，卻要徹底廢除，完全打碎他們的柱像。
EXOD|23|25|你們要事奉耶和華－你們的上帝，他必賜福給你的糧食和水，也必從你中間除去疾病。
EXOD|23|26|你境內必沒有流產的、不生育的。我要使你享滿你年日的數目。
EXOD|23|27|凡你所到的地方，我要使那裏的眾百姓在你面前驚慌失措，又要使你所有的仇敵轉身逃跑。
EXOD|23|28|我要派瘟疫 在你的前面，把 希未 人、 迦南 人、 赫 人從你面前趕出去。
EXOD|23|29|我不在一年之內把他們從你面前趕出去，恐怕地會荒廢，野地的走獸增多危害你。
EXOD|23|30|我要逐漸把他們從你面前趕出去，直到你的人數增多，承受那地為業。
EXOD|23|31|我要定你的疆界，從 紅海 直到 非利士海 ，從曠野直到 大河 。我要把那地的居民交在你手中，你要把他們從你面前趕出去。
EXOD|23|32|不可跟他們和他們的神明立約。
EXOD|23|33|他們不可住在你的地上，免得他們使你得罪我。你若事奉他們的神明，必成為你的圈套。」
EXOD|24|1|耶和華對 摩西 說：「你和 亞倫 、 拿答 、 亞比戶 ，以及 以色列 長老中的七十人，都要上到耶和華這裏來，遠遠地下拜。
EXOD|24|2|只有 摩西 可以接近耶和華，其他的人卻不可接近；百姓也不可和他一同上來。」
EXOD|24|3|摩西 下山，向百姓陳述耶和華一切的命令和典章。眾百姓齊聲說：「耶和華所吩咐的一切，我們都必遵行。」
EXOD|24|4|摩西 將耶和華一切的命令都寫下來。 他清早起來，在山腳築了一座壇，按著 以色列 十二支派立了十二根石柱。
EXOD|24|5|他差派 以色列 的年輕人去獻燔祭，又宰牛獻給耶和華為平安祭。
EXOD|24|6|摩西 將血的一半盛在盆中，另一半灑在壇上。
EXOD|24|7|然後，他拿起約書來，念給百姓聽。他們說：「耶和華所吩咐的一切，我們都必遵行，也必聽從。」
EXOD|24|8|摩西 把血灑在百姓身上，說：「看哪！這是立約的血，是耶和華按照這一切的命令和你們立約的憑據。」
EXOD|24|9|摩西 、 亞倫 、 拿答 、 亞比戶 ，以及 以色列 長老中的七十人都上去，
EXOD|24|10|看見了 以色列 的上帝。在他的腳下，彷彿有藍寶石鋪道，明淨如天。
EXOD|24|11|他不把手伸在 以色列 領袖的身上。他們瞻仰上帝，又吃又喝。
EXOD|24|12|耶和華對 摩西 說：「你上山到我這裏來，就在那裏，我要將石版，就是我所寫的律法和誡命賜給你，使你可以教導他們。」
EXOD|24|13|摩西 和他的助手 約書亞 站起來； 摩西 上了上帝的山。
EXOD|24|14|摩西 對長老們說：「你們在這裏等我們，直到我們再回到你們這裏。看哪， 亞倫 和 戶珥 與你們同在。誰有訴訟，可以去找他們。」
EXOD|24|15|摩西 上山，有雲彩把山遮蓋。
EXOD|24|16|耶和華的榮耀駐在 西奈山 ，雲彩遮蓋了山六天，第七天他從雲中呼叫 摩西 。
EXOD|24|17|耶和華的榮耀在山頂上，在 以色列 人眼前，形狀如吞噬的火。
EXOD|24|18|摩西 進入雲中，登上了山。 摩西 在山上四十晝夜。
EXOD|25|1|耶和華吩咐 摩西 說：
EXOD|25|2|「你要吩咐 以色列 人獻禮物給我。凡甘心樂意獻給我的禮物，你們都可以收下。
EXOD|25|3|要從他們收的禮物是：金、銀、銅，
EXOD|25|4|藍色、紫色、朱紅色紗 ，細麻，山羊毛，
EXOD|25|5|染紅的公羊皮、精美的皮料，金合歡木，
EXOD|25|6|點燈的油，做膏油的香料、做香的香料，
EXOD|25|7|紅瑪瑙與寶石，可以鑲嵌在以弗得和胸袋上。
EXOD|25|8|他們要為我造聖所，使我住在他們中間。
EXOD|25|9|你們要按照我指示你的，帳幕和其中一切器具的樣式，照樣去做。」
EXOD|25|10|「他們要用金合歡木做一個櫃子，長二肘半，寬一肘半，高一肘半。
EXOD|25|11|你要把它裏裏外外包上純金，四圍要鑲上金邊。
EXOD|25|12|要鑄造四個金環，安在櫃子的四腳上；這邊兩個環，那邊兩個環。
EXOD|25|13|要用金合歡木做兩根槓，包上金子。
EXOD|25|14|要把槓穿過櫃旁的環，以便抬櫃。
EXOD|25|15|這槓要留在櫃的環內，不可抽出來。
EXOD|25|16|要把我所要賜給你的法版 放在櫃裏。
EXOD|25|17|要用純金做一個櫃蓋 ，長二肘半，寬一肘半。
EXOD|25|18|要造兩個用金子錘出的基路伯，從櫃蓋的兩端錘出它們。
EXOD|25|19|這端錘出一個基路伯，那端錘出一個基路伯；從櫃蓋的兩端錘出兩個基路伯。
EXOD|25|20|二基路伯的翅膀要向上張開，用翅膀遮住櫃蓋，臉要彼此相對；基路伯的臉要朝向櫃蓋。
EXOD|25|21|要把櫃蓋安在櫃的上邊，又要把我所要賜給你的法版放在櫃裏。
EXOD|25|22|我要在那裏與你相會，並要從法版之櫃的櫃蓋上，兩個基路伯的中間，將我要吩咐 以色列 人的一切事告訴你。」
EXOD|25|23|「你要用金合歡木做一張供桌，長二肘，寬一肘，高一肘半，
EXOD|25|24|把它包上純金，四圍鑲上金邊。
EXOD|25|25|供桌的四圍各做一掌寬的邊緣，邊緣周圍要鑲上金邊。
EXOD|25|26|要為供桌做四個金環，把環安在四個桌腳的四角上。
EXOD|25|27|環要靠近邊緣，以便穿槓抬供桌。
EXOD|25|28|要用金合歡木做兩根槓，包上金子，用來抬供桌。
EXOD|25|29|要用純金做桌上的盤、碟，以及澆酒祭的壺和杯。
EXOD|25|30|要把供餅擺在桌上，常在我面前。」
EXOD|25|31|「要造一座用純金錘出的燈臺。燈臺的座、幹、杯、花萼和花瓣，都要和燈臺接連一塊。
EXOD|25|32|燈臺兩旁要伸出六根枝子：這邊三根，那邊三根。
EXOD|25|33|這邊枝子上有三個杯，形狀像杏花，有花萼有花瓣；那邊枝子上也有三個杯，形狀像杏花，有花萼有花瓣。從燈臺伸出來的六根枝子都是如此。
EXOD|25|34|燈臺本身要有四個杯，形狀像杏花，有花萼有花瓣。
EXOD|25|35|燈臺的第一對枝子下面有花萼，燈臺的第二對枝子下面有花萼，燈臺的第三對枝子下面也有花萼；燈臺伸出的六根枝子都是如此。
EXOD|25|36|花萼和枝子都要和燈臺接連一塊，全是從一塊純金錘出來的。
EXOD|25|37|要做燈臺的七盞燈，燈要點燃，照亮前面。
EXOD|25|38|要用純金做燈剪和燈盤。
EXOD|25|39|做燈臺和這一切的器具要用一他連得純金。
EXOD|25|40|要謹慎，照著在山上指示你的樣式去做。」
EXOD|26|1|「你要用十幅幔子做帳幕。這些幔子要用搓的細麻和藍色、紫色、朱紅色紗織成，並且以刺繡的手藝繡上基路伯。
EXOD|26|2|每幅幔子要長二十八肘，每幅幔子寬四肘，全部的幔子尺寸都要一樣。
EXOD|26|3|這五幅幔子要彼此相連；那五幅也彼此相連。
EXOD|26|4|在這一組相連幔子的末幅邊上要縫藍色的鈕環；在另一組相連幔子的末幅邊上也要照樣做。
EXOD|26|5|這幅幔子上要縫五十個鈕環，另一組相連幔子的末幅上也縫五十個鈕環，環環相對。
EXOD|26|6|要做五十個金鉤，用鉤子使幔子彼此相連，成為一個帳幕。
EXOD|26|7|「你要用山羊毛織十一幅幔子來作帳幕的罩棚。
EXOD|26|8|每幅幔子要長三十肘，每幅幔子寬四肘；十一幅幔子的尺寸都要一樣。
EXOD|26|9|要把五幅幔子連成一幅，又把六幅幔子連成一幅，這第六幅幔子要在罩棚的前面摺上去。
EXOD|26|10|在這一組相連幔子的末幅邊上要縫五十個鈕環；在另一組相連幔子的末幅邊上也縫五十個鈕環。
EXOD|26|11|要做五十個銅鉤，鉤在鈕環中，使罩棚相連成為一個。
EXOD|26|12|罩棚幔子餘下垂著的，那餘下的半幅要垂在帳幕的背面。
EXOD|26|13|罩棚的幔子兩旁所餘下的，這邊一肘，那邊一肘，要垂在帳幕的兩邊，蓋住帳幕。
EXOD|26|14|要用染紅的公羊皮做罩棚的蓋，再用精美皮料做外層的蓋。
EXOD|26|15|「你要用金合歡木做豎立帳幕的木板，
EXOD|26|16|木板要長十肘，每塊板寬一肘半，
EXOD|26|17|每塊板有兩個榫頭可以彼此銜接。帳幕一切的板都要這樣做。
EXOD|26|18|你要做帳幕的木板：南面，就是面向南方的那一邊，要做二十塊板。
EXOD|26|19|在這二十塊板底下要做四十個帶卯眼的銀座；兩個卯眼接連這塊板上的兩個榫頭，另外兩個卯眼接連那塊板上的兩個榫頭。
EXOD|26|20|帳幕的第二邊，就是北面，也要做二十塊板，
EXOD|26|21|和四十個帶卯眼的銀座；這塊板底下有兩個卯眼，那塊板底下也有兩個卯眼。
EXOD|26|22|帳幕的後面，就是西面，要做六塊板。
EXOD|26|23|帳幕後面的角落要做兩塊板。
EXOD|26|24|下端的板是成雙的，上端要連在一起，直到頂端的第一個環子；兩塊板都要這樣，做成兩個角落。
EXOD|26|25|一共有八塊板和十六個帶卯眼的銀座；這塊板底下有兩個卯眼，那塊板底下也有兩個卯眼。
EXOD|26|26|「你要用金合歡木做橫木：為帳幕這面的板做五根橫木，
EXOD|26|27|為帳幕那面的板做五根橫木，又為帳幕後面，就是朝西的板做五根橫木。
EXOD|26|28|板腰間的橫木，要從一頭通到另一頭。
EXOD|26|29|板要包上金子，又要做板上的金環來套橫木；橫木也要包上金子。
EXOD|26|30|要照著在山上所指示你的樣式，把帳幕豎立起來。
EXOD|26|31|「你要用藍色、紫色、朱紅色紗，和搓的細麻織幔子，以刺繡的手藝繡上基路伯。
EXOD|26|32|要把幔子掛在四根包金的金合歡木柱子上，柱子有金鉤，並且安在四個帶卯眼的銀座上。
EXOD|26|33|要把幔子垂掛在鉤子上，把法櫃抬進幔子內；這幔子要將聖所和至聖所隔開。
EXOD|26|34|又要把櫃蓋安在至聖所內的法櫃上，
EXOD|26|35|把供桌安在幔子的外面，供桌在北面，燈臺在帳幕的南面，和供桌相對。
EXOD|26|36|「你要用藍色、紫色、朱紅色紗，和搓的細麻，以刺繡的手藝為帳幕織門簾。
EXOD|26|37|要用金合歡木為簾子做五根柱子，包上金子。柱子有金鉤，又為柱子鑄造五個帶卯眼的銅座。」
EXOD|27|1|「你要用金合歡木做祭壇，長五肘，寬五肘，這壇是正方形的，高三肘。
EXOD|27|2|要在壇的四角做四個翹角，與壇接連一塊；要把壇包上銅。
EXOD|27|3|要做桶子來盛壇上的灰，又要做鏟子、盤子、肉叉和火盆；壇上一切的器具都要用銅做。
EXOD|27|4|要為壇做一個銅網，在網的四角做四個銅環，
EXOD|27|5|把網安在壇四圍的邊的下面，使網垂到壇的半腰。
EXOD|27|6|又要用金合歡木為壇做槓，包上銅。
EXOD|27|7|這槓要穿過壇兩旁的環子，用來抬壇。
EXOD|27|8|要用板做壇，壇的中心是空的，都照著在山上所指示你的樣式做。」
EXOD|27|9|「你要做帳幕的院子。南面，就是面向南方的那一邊，要用搓的細麻做院子的帷幔，長一百肘，
EXOD|27|10|院子要有二十根柱子，二十個帶卯眼的銅座。要用銀做柱子的鉤和箍。
EXOD|27|11|北面的長度也一樣，帷幔長一百肘，要有二十根柱子，二十個帶卯眼的銅座。要用銀做柱子的鉤和箍。
EXOD|27|12|院子的西面有帷幔，寬五十肘，帷幔要有十根柱子，十個帶卯眼的座。
EXOD|27|13|院子的東面，就是面向東方的那一邊，寬五十肘。
EXOD|27|14|一邊的帷幔有十五肘，要有三根柱子，三個帶卯眼的座。
EXOD|27|15|另一邊的帷幔也有十五肘，要有三根柱子，三個帶卯眼的座。
EXOD|27|16|院子的門要有二十肘長的簾子，用藍色、紫色、朱紅色紗，和搓的細麻，以刺繡的手藝織成；要有四根柱子，四個帶卯眼的座。
EXOD|27|17|院子四圍一切的柱子都要用銀子箍著，要用銀做柱子的鉤子，用銅做帶卯眼的座。
EXOD|27|18|院子要長一百肘，寬五十肘 ，高五肘。要用搓的細麻做帷幔，用銅做帶卯眼的座。
EXOD|27|19|帳幕中各樣用途的器具，以及帳幕一切的橛子和院子裏一切的橛子，都要用銅做。」
EXOD|27|20|「你要吩咐 以色列 人，把搗成的純橄欖油拿來給你，用以點燈，使燈經常點著；
EXOD|27|21|在會幕中法櫃前的幔子外， 亞倫 和他的兒子要從晚上到早晨，在耶和華面前照管這燈。這要成為 以色列 人世世代代永遠的定例。」
EXOD|28|1|「你要從 以色列 人中，叫你的哥哥 亞倫 和他的兒子 拿答 、 亞比戶 、 以利亞撒 、 以他瑪 一同親近你，作事奉我的祭司。
EXOD|28|2|你要為你哥哥 亞倫 做聖衣，以示尊嚴和華美。
EXOD|28|3|要吩咐一切心中有智慧的，就是我用智慧的靈所充滿的人，為 亞倫 做衣服，使他分別為聖，作事奉我的祭司。
EXOD|28|4|所要做的是胸袋、以弗得、外袍、織成的內袍、禮冠和腰帶。他們要為你哥哥 亞倫 和他的兒子做聖衣，使他們作祭司事奉我。
EXOD|28|5|要用金色、藍色、紫色、朱紅色紗，和細麻去縫製。
EXOD|28|6|「他們要用金色、藍色、紫色、朱紅色紗，和搓的細麻，以刺繡的手藝做以弗得。
EXOD|28|7|以弗得當有兩條肩帶，接上兩端，使它相連。
EXOD|28|8|以弗得的精緻帶子，要以一樣的手藝，用金色、藍色、紫色、朱紅色紗，和搓的細麻縫製，與以弗得接連在一起。
EXOD|28|9|要取兩塊紅瑪瑙，在上面刻 以色列 兒子的名字：
EXOD|28|10|六個名字在一塊寶石上，六個名字在另一塊寶石上，都按照他們出生的次序。
EXOD|28|11|要以雕刻寶石的手藝，如同刻印章，把 以色列 兒子的名字刻在這兩塊寶石上，並把寶石鑲在金槽裏。
EXOD|28|12|要把這兩塊寶石安在以弗得的兩條肩帶上，為 以色列 人作紀念石。 亞倫 要在耶和華面前把他們的名字帶在兩肩上，作為紀念。
EXOD|28|13|要用金子做兩個槽，
EXOD|28|14|再用純金打兩條鏈子，像編成的繩子一樣，把這編成的金鏈扣在槽上。」
EXOD|28|15|「你要以刺繡的手藝做一個決斷的胸袋，和做以弗得的方法一樣，用金色、藍色、紫色、朱紅色紗，和搓的細麻縫製。
EXOD|28|16|胸袋是正方形的，疊成兩層，長一虎口，寬一虎口。
EXOD|28|17|要在上面鑲四行寶石：第一行是紅寶石、紅璧璽、紅玉；
EXOD|28|18|第二行是綠寶石、藍寶石、金剛石；
EXOD|28|19|第三行是紫瑪瑙、白瑪瑙、紫晶；
EXOD|28|20|第四行是水蒼玉、紅瑪瑙、碧玉。這些都要鑲在金槽中。
EXOD|28|21|這些寶石要有 以色列 十二個兒子的名字，如同刻印章，每一顆有自己的名字，代表十二個支派。
EXOD|28|22|要在胸袋上用純金打鏈子，像編成的繩子一樣。
EXOD|28|23|要為胸袋做兩個金環，把這兩個環安在胸袋的兩端。
EXOD|28|24|要把那兩條編成的金鏈繫在胸袋兩端的兩個環上。
EXOD|28|25|又要把鏈子的另外兩端扣在兩個槽上，安在以弗得前面的肩帶上。
EXOD|28|26|要做兩個金環，安在胸袋的兩端，在以弗得裏面的邊上。
EXOD|28|27|再做兩個金環，安在以弗得前面兩條肩帶的下邊，靠近接縫處，在以弗得精緻帶子的上面。
EXOD|28|28|要用藍色的帶子把胸袋的環與以弗得的環繫住，使胸袋綁在以弗得的精緻帶子上，不致鬆脫。
EXOD|28|29|亞倫 進聖所的時候，要把刻著 以色列 兒子名字的決斷胸袋帶著，放在心上，在耶和華面前常作紀念。
EXOD|28|30|又要將烏陵和土明 放在決斷胸袋裏； 亞倫 進到耶和華面前的時候，要放在心上。這樣， 亞倫 在耶和華面前要把 以色列 人的決斷胸袋常常帶著，放在心上。」
EXOD|28|31|「你要做以弗得的外袍，顏色全是藍的。
EXOD|28|32|袍上方的中間要留一個領口，領口周圍的領邊要以手藝編織而成，好像鎧甲的領口，免得破裂。
EXOD|28|33|袍子下襬，就是下襬的周圍要用藍色、紫色、朱紅色紗做石榴，周圍的石榴中間要有金鈴鐺：
EXOD|28|34|一個金鈴鐺一個石榴，一個金鈴鐺一個石榴，在袍子下襬的周圍。
EXOD|28|35|亞倫 供職的時候要穿這袍。他進入聖所到耶和華面前，以及出來的時候，袍上的鈴聲必被聽見，使他不至於死。
EXOD|28|36|「你要用純金做一面牌，如同刻印章，在上面刻『歸耶和華為聖』。
EXOD|28|37|要用藍色的帶子把牌繫在禮冠上，在禮冠的正前面。
EXOD|28|38|這牌必在 亞倫 的額上， 亞倫 要擔當干犯聖物的罪孽；這聖物是 以色列 人在一切聖禮物上所分別為聖的。這牌要常在他的額上，使他們可以在耶和華面前蒙悅納。
EXOD|28|39|要用細麻編織內袍，用細麻做禮冠，又以刺繡的手藝做腰帶。
EXOD|28|40|「你要為 亞倫 的兒子做內袍、腰帶、頭巾，以示尊嚴和華美。
EXOD|28|41|要把這些給你哥哥 亞倫 和他的兒子穿戴，又要膏他們，授予聖職，使他們分別為聖，作事奉我的祭司。
EXOD|28|42|要用細麻布給他們做褲子來遮掩下體，從腰間直到大腿。
EXOD|28|43|亞倫 和他兒子進入會幕，或接近祭壇，在聖所供職的時候要穿上褲子，免得擔當罪孽而死。這要成為 亞倫 和他後裔永遠的定例。」
EXOD|29|1|「這是你使他們分別為聖，作事奉我的祭司時要做的事：取一頭公牛犢，兩隻無殘疾的公綿羊，
EXOD|29|2|無酵餅、用油調和的無酵餅，和抹油的無酵薄餅；這些餅都要用細麥麵做成。
EXOD|29|3|這些餅要裝在一個籃子裏，用籃子帶來，又把公牛和兩隻公綿羊牽來。
EXOD|29|4|要帶 亞倫 和他兒子到會幕的門口，用水洗他們。
EXOD|29|5|要拿服裝，給 亞倫 穿上內袍和以弗得的外袍，以及以弗得，又帶上胸袋，束上以弗得精緻的帶子。
EXOD|29|6|要把禮冠戴在他頭上，將聖冕加在禮冠上，
EXOD|29|7|把膏油倒在他頭上膏他。
EXOD|29|8|要帶他的兒子來，給他們穿上內袍。
EXOD|29|9|要給 亞倫 和他的兒子束上腰帶，裹上頭巾，他們就憑永遠的定例得祭司的職分。又要授聖職給 亞倫 和他的兒子。
EXOD|29|10|「你要把公牛牽到會幕前， 亞倫 和他的兒子要按手在公牛的頭上。
EXOD|29|11|你要在耶和華面前，在會幕的門口宰這公牛。
EXOD|29|12|要取些公牛的血，用指頭抹在祭壇的四個翹角上，把其餘的血全倒在壇的底座上。
EXOD|29|13|要把所有包著內臟的脂肪、肝上的網油、兩個腎和腎上的脂肪，都燒在壇上。
EXOD|29|14|只是公牛的肉、皮、糞都要在營外用火焚燒；這牛是贖罪祭。
EXOD|29|15|「你要牽一隻公綿羊來， 亞倫 和他兒子要按手在這羊的頭上。
EXOD|29|16|你要宰這羊，把血灑在祭壇的周圍。
EXOD|29|17|再把羊切成肉塊，洗淨內臟和腿，連肉塊和頭放在一處。
EXOD|29|18|要把全羊燒在壇上。這是獻給耶和華的燔祭，是獻給耶和華馨香的火祭。」
EXOD|29|19|「你要把第二隻公綿羊牽來， 亞倫 和他兒子要按手在這羊的頭上。
EXOD|29|20|你要宰這羊，取些血抹在 亞倫 的右耳垂和他兒子的右耳垂上，又抹在他們右手的大拇指和右腳的大腳趾上，然後把其餘的血灑在壇的周圍。
EXOD|29|21|你要取些膏油和壇上的血，彈在 亞倫 和他的衣服上，以及他兒子和他們的衣服上； 亞倫 和他的衣服，他兒子和他們的衣服都成為聖了。
EXOD|29|22|「你要取這羊的脂肪，肥尾巴、包著內臟的脂肪、肝上的網油、兩個腎、腎上的脂肪和右腿，這是聖職禮所獻的公綿羊；
EXOD|29|23|再從耶和華面前那裝無酵餅的籃子中取一個餅、一個油餅和一個薄餅，
EXOD|29|24|把它們都放在 亞倫 的手和他兒子的手上，在耶和華面前搖一搖，作為搖祭。
EXOD|29|25|然後，你要從他們手中接過來，放在燔祭上，一起燒在壇上，作為耶和華面前馨香之氣；這是獻給耶和華的火祭。
EXOD|29|26|「你要取 亞倫 聖職禮所獻公綿羊的胸，在耶和華面前搖一搖，作為搖祭；這份就是你的。
EXOD|29|27|那搖祭的胸和舉祭的腿，就是聖職禮獻公綿羊時所搖的、所舉的，你要使它們分別為聖，是歸給 亞倫 和他兒子的。
EXOD|29|28|這是 亞倫 和他子孫憑永遠的定例從 以色列 人中所應得的；因為這是舉祭，是從 以色列 人的平安祭中取出，作為獻給耶和華的舉祭。
EXOD|29|29|「 亞倫 的聖衣要傳給他的子孫，使他們在受膏和承接聖職的時候穿上。
EXOD|29|30|他的子孫接續他當祭司的，每逢進入會幕在聖所供職的時候，要穿這聖衣七天。
EXOD|29|31|「你要拿聖職禮所獻的公綿羊，在聖處煮牠的肉。
EXOD|29|32|亞倫 和他兒子要在會幕的門口吃這羊的肉和籃子裏的餅。
EXOD|29|33|他們要吃那些用來贖罪之物，好承接聖職，使他們分別為聖。外人不可吃，因為這是聖物。
EXOD|29|34|那聖職禮所獻的肉或餅，若有剩餘留到早晨，就要把剩下的用火燒了，不可再吃，因為這是聖物。
EXOD|29|35|「你要這樣照我一切所吩咐的，向 亞倫 和他兒子行授聖職禮七天。
EXOD|29|36|為了贖罪，每天要獻一頭公牛為贖罪祭。你要為祭壇贖罪，使壇潔淨，並要用膏抹壇，使壇成為聖。
EXOD|29|37|要為壇贖罪七天，使壇成為聖，壇就成為至聖。凡觸摸壇的都成為聖。」
EXOD|29|38|「這是你要獻在壇上的：每天不可間斷地獻兩隻一歲的羔羊；
EXOD|29|39|早晨獻第一隻羔羊，黃昏獻第二隻羔羊。
EXOD|29|40|獻第一隻羔羊時，要同時獻上十分之一伊法細麵，調和四分之一欣搗成的油，再獻四分之一欣酒作澆酒祭。
EXOD|29|41|黃昏你獻第二隻羔羊，要照早晨的素祭和同獻的澆酒祭獻上，作為獻給耶和華馨香的火祭。
EXOD|29|42|這要在耶和華面前，在會幕的門口，作為你們世世代代經常獻的燔祭。我要在那裏與你們 相會，和你說話。
EXOD|29|43|我要在那裏與 以色列 人相會，會幕就要因我的榮耀成為聖。
EXOD|29|44|我要使會幕和祭壇分別為聖，也要使 亞倫 和他的兒子分別為聖，作事奉我的祭司。
EXOD|29|45|我要住在 以色列 人中，作他們的上帝。
EXOD|29|46|他們必知道我是耶和華－他們的上帝，是將他們從 埃及 地領出來的，為要住在他們中間。我是耶和華－他們的上帝 。」
EXOD|30|1|「你要用金合歡木做一座燒香的壇，
EXOD|30|2|長一肘，寬一肘，這壇是正方形的，高二肘。壇的四個翹角與壇接連一塊。
EXOD|30|3|要把壇的上面與壇的四圍，以及壇的四個翹角包上純金；又要在壇的四圍鑲上金邊。
EXOD|30|4|要在壇的兩個對側，金邊下面做兩個金環，用來穿槓抬壇。
EXOD|30|5|要用金合歡木做槓，包上金子。
EXOD|30|6|要把壇放在法櫃前的幔子外，對著法櫃上的櫃蓋，就是我與你相會的地方。
EXOD|30|7|亞倫 要在壇上燒芬芳的香；每早晨整理燈的時候，他都要燒這香。
EXOD|30|8|黃昏點燈的時候， 亞倫 也要燒這香。這是你們世世代代在耶和華面前常燒的香。
EXOD|30|9|在這壇上不可燒別樣的香，不可獻燔祭、素祭，也不可獻澆酒祭。
EXOD|30|10|亞倫 每年一次要為壇的四個翹角贖罪。他每年一次要用贖罪祭的血為壇贖罪，作為世世代代的定例。這壇在耶和華面前是至聖的。」
EXOD|30|11|耶和華吩咐 摩西 說：
EXOD|30|12|「你數點 以色列 人，計算人頭時，被數的每一個人要把他生命的贖價獻給耶和華，免得災殃在數點中臨到他們。
EXOD|30|13|每一個被數的人要按照聖所的舍客勒，付半舍客勒，一舍客勒是二十季拉；這半舍客勒是獻給耶和華的禮物。
EXOD|30|14|每一個被數的人，就是二十歲以上的，要將這禮物獻給耶和華。
EXOD|30|15|富有的不必多付，貧窮的也不可少出，各人都要獻半舍客勒給耶和華，作你們生命的贖價。
EXOD|30|16|你要向 以色列 人收這贖罪的銀子，用在會幕的事工。這要在耶和華面前為 以色列 人作紀念，作你們生命的贖價。」
EXOD|30|17|耶和華吩咐 摩西 說：
EXOD|30|18|「你要用銅做洗濯盆和盆座，用來洗濯。要將盆放在會幕和祭壇的中間，盆裏盛水。
EXOD|30|19|亞倫 和他的兒子要用這盆洗手洗腳。
EXOD|30|20|他們進會幕，或是走近壇前供職，獻火祭給耶和華的時候，必須用水洗濯，免得死亡；
EXOD|30|21|他們要洗手洗腳，免得死亡。這是 亞倫 和他的後裔世世代代永遠的定例。」
EXOD|30|22|耶和華吩咐 摩西 說：
EXOD|30|23|「你要取上等的香料，就是五百舍客勒流質的沒藥、二百五十香肉桂、二百五十香菖蒲，
EXOD|30|24|和五百桂皮，都按照聖所的舍客勒；再取一欣橄欖油，
EXOD|30|25|以做香的方法調和製成聖膏油，它就成為聖膏油。
EXOD|30|26|要用這膏油抹會幕和法櫃，
EXOD|30|27|供桌和供桌的一切器具，燈臺和燈臺的器具 ，以及香壇、
EXOD|30|28|燔祭壇和壇的一切器具，洗濯盆和盆座。
EXOD|30|29|你要使這些分別為聖，成為至聖；凡觸摸它們的都成為聖。
EXOD|30|30|要膏 亞倫 和他的兒子，使他們分別為聖，作事奉我的祭司。
EXOD|30|31|你要吩咐 以色列 人說：『你們要世世代代以這油為我的聖膏油。
EXOD|30|32|不可把這油倒在別人身上，也不可用配製這膏油的方法製成同樣的膏油。這膏油是聖的，你們要以它為聖。
EXOD|30|33|凡調和與此類似的膏油，或將它膏在別人身上的，這人要從百姓中剪除。』」
EXOD|30|34|耶和華吩咐 摩西 說：「你要取香料，就是拿他弗、施喜列、喜利比拿，這些香料再加純乳香，每樣都要相同的分量。
EXOD|30|35|你要用這些加上鹽，以配製香料的方法，製成純淨又神聖的香。
EXOD|30|36|要取一點這香，搗成細的粉，放在會幕中的法櫃前，就是我和你相會的地方。你們要以這香為至聖。
EXOD|30|37|你們不可用這配製的方法為自己做香；要以這香為聖，歸於耶和華。
EXOD|30|38|為要聞香味而配製同樣的香的，這人要從百姓中剪除。」
EXOD|31|1|耶和華吩咐 摩西 說：
EXOD|31|2|「你看，我已經題名召 猶大 支派中 戶珥 的孫子， 烏利 的兒子 比撒列 。
EXOD|31|3|我以上帝的靈充滿他，使他有智慧，有聰明，有知識，能做各樣的工，
EXOD|31|4|能設計圖案，用金、銀、銅製造各物，
EXOD|31|5|又能雕刻鑲嵌用的寶石，雕刻木頭，做各樣的工。
EXOD|31|6|看哪，我委派 但 支派中 亞希撒抹 的兒子 亞何利亞伯 與他同工。凡心裏有智慧的，我更要賜給他們智慧的心，能做我所吩咐你的一切，
EXOD|31|7|就是會幕、法櫃和其上的櫃蓋、會幕中一切的器具、
EXOD|31|8|供桌和供桌的器具、純金的燈臺和燈臺的一切器具、香壇、
EXOD|31|9|燔祭壇和壇的一切器具、洗濯盆與盆座、
EXOD|31|10|供祭司職分用的精緻禮服， 亞倫 祭司的聖衣和他兒子的衣服，
EXOD|31|11|以及膏油和聖所用的芬芳的香。他們都要照我所吩咐的一切去做。」
EXOD|31|12|耶和華對 摩西 說：
EXOD|31|13|「你要吩咐 以色列 人說：『你們務要守我的安息日，因為這是你我之間世世代代的記號，叫你們知道我是耶和華，是使你們分別為聖的。
EXOD|31|14|你們要守安息日，以它為聖日。凡干犯這日的，必被處死；凡在這日做工的，那人必從百姓中剪除。
EXOD|31|15|六日要做工，但第七日是向耶和華守完全安息的安息聖日。凡在安息日做工的，必被處死。』
EXOD|31|16|以色列 人要守安息日，世世代代守安息日為永遠的約。
EXOD|31|17|這是我和 以色列 人之間永遠的記號，因為六日之內耶和華造天地，第七日就安息舒暢。」
EXOD|31|18|耶和華在 西奈山 和 摩西 說完了話，就把兩塊法版交給他，是上帝用指頭寫的石版。
EXOD|32|1|百姓見 摩西 遲遲不下山，就聚集到 亞倫 那裏，對他說：「起來！為我們造神明，在我們前面引路，因為領我們出 埃及 地的那個 摩西 ，我們不知道他遭遇了甚麼事。」
EXOD|32|2|亞倫 對他們說：「你們去摘下你們妻子、兒女耳上的金環，拿來給我。」
EXOD|32|3|眾百姓就摘下他們耳上的金環，拿來給 亞倫 。
EXOD|32|4|亞倫 從他們手裏接過來，用模子塑造它，把它鑄成一頭牛犢。他們就說：「 以色列 啊，這是領你出 埃及 地的神明！」
EXOD|32|5|亞倫 看見，就在牛犢面前築壇。 亞倫 宣告說：「明日要向耶和華守節。」
EXOD|32|6|次日清早，百姓起來獻燔祭和平安祭，就坐下吃喝，起來玩樂。
EXOD|32|7|耶和華吩咐 摩西 ：「下去吧，因為你從 埃及 領上來的百姓已經敗壞了。
EXOD|32|8|他們這麼快偏離了我所吩咐的道，為自己鑄了一頭牛犢，向它跪拜，向它獻祭，說：『 以色列 啊，這就是領你出 埃及 地的神明。』」
EXOD|32|9|耶和華對 摩西 說：「我看這百姓，看哪，他們真是硬著頸項的百姓。
EXOD|32|10|現在，你且由著我，我要向他們發烈怒，滅絕他們，但我要使你成為大國。」
EXOD|32|11|摩西 就懇求耶和華－他的上帝，說：「耶和華啊，你為甚麼向你的百姓發烈怒呢？這百姓是你用大能大力的手從 埃及 地領出來的！
EXOD|32|12|為甚麼讓 埃及 人說：『他領他們出去，是要降災禍給他們，在山中把他們殺了，將他們從地上除滅』呢？求你回心轉意，不發你的烈怒，不降災禍給你的百姓。
EXOD|32|13|求你記念你的僕人 亞伯拉罕 、 以撒 、 以色列 。你曾向他們指著自己起誓說：『我必使你們的後裔像天上的星那樣多，並且我要將所應許的這全地賜給你們的後裔，讓他們永遠承受為業。』」
EXOD|32|14|於是耶和華改變心意，不把所說的災禍降給他的百姓。
EXOD|32|15|摩西 轉身下山，手裏拿著兩塊法版。這版的兩面都寫著字，正面背面都有字。
EXOD|32|16|版是上帝的工作，字是上帝寫的字，刻在版上。
EXOD|32|17|約書亞 一聽見百姓呼喊的聲音，就對 摩西 說：「在營裏有戰爭的聲音。」
EXOD|32|18|摩西 說：「這不是打勝仗的聲音，也不是打敗仗的聲音，我聽見的是歌唱的聲音。」
EXOD|32|19|摩西 走近營前，看見牛犢，又看見人在跳舞，就發烈怒，把兩塊版從手中扔到山下摔碎了。
EXOD|32|20|他將他們所鑄的牛犢用火焚燒，磨得粉碎，撒在水面上，叫 以色列 人喝。
EXOD|32|21|摩西 對 亞倫 說：「這百姓向你做了甚麼呢？你竟使他們陷入大罪中！」
EXOD|32|22|亞倫 說：「求我主不要發烈怒。你知道這百姓，他們是向惡的。
EXOD|32|23|他們對我說：『你為我們造神明，在我們前面引路，因為領我們出 埃及 地的那個 摩西 ，我們不知道他遭遇了甚麼事。』
EXOD|32|24|我對他們說：『凡有金環的可以摘下來』，他們就給了我。我把金環扔在火中，這牛犢就出來了。」
EXOD|32|25|摩西 見百姓放肆，因 亞倫 縱容他們，使這事成了敵人的笑柄，
EXOD|32|26|就站在營門前，說：「凡屬耶和華的人，都到我這裏來！」於是 利未 人都聚集到他那裏。
EXOD|32|27|他對他們說：「耶和華－ 以色列 的上帝這樣說：『你們各人把刀佩在腰間，從這門到那門，來回走遍全營，各人要殺自己的弟兄、鄰舍和親人。』」
EXOD|32|28|利未 人遵照 摩西 的話做了。那一天百姓中倒下的約有三千人。
EXOD|32|29|摩西 說：「今天你們要奉獻自己 來事奉耶和華，因為各人犧牲自己的兒子和弟兄，使耶和華今天賜福給你們。」
EXOD|32|30|第二天， 摩西 對百姓說：「你們犯了大罪。我如今要上耶和華那裏去，或許可以為你們贖罪。」
EXOD|32|31|摩西 回到耶和華那裏，說：「唉！這百姓犯了大罪，為自己造了金的神明。
EXOD|32|32|現在，求你赦免他們的罪；不然，就把我從你所寫的冊上除名。」
EXOD|32|33|耶和華對 摩西 說：「誰得罪我，我就把他從我的冊上除去。
EXOD|32|34|現在你去，領這百姓往我所告訴你的地方去，看哪，我的使者必在你的前面引路。到了該懲罰的時候，我必懲罰他們的罪。」
EXOD|32|35|耶和華降災與百姓，因為他們和 亞倫 一起造了牛犢。
EXOD|33|1|耶和華吩咐 摩西 說：「去，離開這裏，你和你從 埃及 地領出來的百姓要上到我起誓應許給 亞伯拉罕 、 以撒 和 雅各 之地去；我曾對他們說：『我要將這地賜給你的後裔』。
EXOD|33|2|我要差遣使者在你前面，把 迦南 人、 亞摩利 人、 赫 人、 比利洗 人、 希未 人、 耶布斯 人趕出
EXOD|33|3|那流奶與蜜之地。但我不與你們上去，因為你們是硬著頸項的百姓，免得我在路上把你們滅絕。」
EXOD|33|4|百姓一聽見這壞的信息，他們就悲哀，沒有人佩戴首飾。
EXOD|33|5|耶和華對 摩西 說：「你對 以色列 人說：『你們是硬著頸項的百姓，我若在你們中間一起上去，只一瞬間，就必把你們滅絕。現在把你們身上的首飾摘下來，我好知道該怎樣處置你們。』」
EXOD|33|6|以色列 人離開 何烈山 以後，就把身上的首飾全都摘下來。
EXOD|33|7|摩西 拿一個帳棚支搭在營外，離營有一段距離，他稱這帳棚為會幕。凡求問耶和華的，就到營外的會幕那裏去。
EXOD|33|8|當 摩西 出營到會幕去的時候，百姓就都起來，各人站在自己帳棚的門口，望著 摩西 ，直到他進了會幕。
EXOD|33|9|摩西 進會幕的時候，雲柱就降下來，停在會幕的門前，耶和華就與 摩西 說話。
EXOD|33|10|眾百姓看見雲柱停在會幕的門前，就都起來，各人在自己帳棚的門口下拜。
EXOD|33|11|耶和華與 摩西 面對面說話，好像人與朋友說話。 摩西 回到營裏去，他的年輕助手 嫩 的兒子 約書亞 卻沒有離開會幕。
EXOD|33|12|摩西 對耶和華說：「看，你曾對我說：『將這百姓領上去』；卻沒有讓我知道你要差派誰與我同去。你還說：『我按你的名認識你，你也在我眼前蒙了恩。』
EXOD|33|13|我如今若在你眼前蒙恩，求你將你的道指示我，使我可以認識你，並在你眼前蒙恩。求你顧念這國是你的子民。」
EXOD|33|14|耶和華說：「我必親自去，讓你安心。」
EXOD|33|15|摩西 說：「你若不親自去，就不要把我們從這裏領上去。
EXOD|33|16|現在，人如何得知我和你的百姓在你眼前蒙恩呢？豈不是因為你與我們同去，使我和你的百姓與地面上的萬民有分別嗎？」
EXOD|33|17|耶和華對 摩西 說：「你所說的這件事，我也會去做，因為你在我眼前蒙了恩，並且我按你的名認識你。」
EXOD|33|18|摩西 說：「求你顯出你的榮耀給我看。」
EXOD|33|19|耶和華說：「我要顯示我一切的美善，在你面前經過，並要在你面前宣告耶和華的名。我要恩待誰就恩待誰，要憐憫誰就憐憫誰。」
EXOD|33|20|他又說：「只是你不能看見我的面，因為沒有人看見我還可以存活。」
EXOD|33|21|耶和華說：「看哪，靠近我這裏有個地方，你可以站在這磐石上。
EXOD|33|22|當我的榮耀經過的時候，我必將你放在磐石縫裏，用我的手掌遮掩你，等我過去，
EXOD|33|23|然後我要將我的手掌收回，你就可以看見我的背，卻看不到我的面。」
EXOD|34|1|耶和華對 摩西 說：「你要鑿出兩塊石版，和先前的一樣；我要把你摔碎的那版上先前所寫的字，寫在這版上。
EXOD|34|2|明日早晨，你要預備好了，上 西奈山 ，在山頂那裏站在我面前。
EXOD|34|3|誰也不可和你上去，整座山都不可見到人，也不可有羊群牛群在山下吃草。」
EXOD|34|4|摩西 就鑿出兩塊石版，和先前的一樣。他清晨起來，遵照耶和華吩咐他的，上 西奈山 去，手裏拿著兩塊石版。
EXOD|34|5|耶和華在雲中降臨，與 摩西 一同站在那裏，宣告耶和華的名。
EXOD|34|6|耶和華在他面前經過，宣告： 「耶和華，耶和華， 有憐憫，有恩惠的上帝， 不輕易發怒， 且有豐盛的慈愛和信實，
EXOD|34|7|為千代的人存留慈愛， 赦免罪孽、過犯和罪惡， 萬不以有罪的為無罪， 必懲罰人的罪， 自父及子，直到三、四代。」
EXOD|34|8|摩西 急忙俯伏在地敬拜，
EXOD|34|9|說：「主啊，我若在你眼前蒙恩，求主在我們中間同行。雖然這是硬著頸項的百姓，求你赦免我們的罪孽和罪惡，接納我們為你的產業。」
EXOD|34|10|耶和華說：「看哪，我要立約，要在你眾百姓面前行奇妙的事，是在全地萬國中未曾做過的。你周圍的萬民要看見我藉著你所行，耶和華可畏懼的作為。
EXOD|34|11|「我今天所吩咐你的，你要謹守。看哪，我要從你面前趕出 亞摩利 人、 迦南 人、 赫 人、 比利洗 人、 希未 人、 耶布斯 人。
EXOD|34|12|你要謹慎，不可與你所要去那地的居民立約，免得他們成為你中間的圈套。
EXOD|34|13|你要拆毀他們的祭壇，打碎他們的柱像，砍斷他們的 亞舍拉 。
EXOD|34|14|不可敬拜別神，因為耶和華是忌邪 的上帝，他的名是忌邪者。
EXOD|34|15|你不可與那地的居民立約，因為他們隨從自己的神明行淫；祭他們神明的時候，有人邀請你參加，你就會吃他的祭物。
EXOD|34|16|你為你兒子娶他們的女兒為妻，他們的女兒因著隨從她們的神明行淫，就引誘你的兒子也隨從她們的神明行淫。
EXOD|34|17|「不可為自己鑄造神像。
EXOD|34|18|「你要守除酵節，照我所吩咐你的，在亞筆月內所定的日期吃無酵餅七天，因為你是在亞筆月內出了 埃及 。
EXOD|34|19|「凡頭生的都是我的；無論是牛是羊，一切頭生的公的牲畜都要分別出來 。
EXOD|34|20|頭生的驢可以用羔羊代贖。若不贖牠，就要打斷牠的頸項。凡頭生的兒子都要贖出來。沒有人可以空手來朝見我。
EXOD|34|21|「六日你要做工，第七日要安息，即使在耕種或收割的時候也要安息。
EXOD|34|22|在收割初熟麥子的時候要守七七節，又要在年底守收藏節。
EXOD|34|23|你所有的男丁要一年三次朝見主耶和華－ 以色列 的上帝。
EXOD|34|24|我要從你面前趕走列國，擴張你的疆界。你一年三次上去朝見耶和華－你上帝的時候，必沒有人貪圖你的地。
EXOD|34|25|「不可將我祭牲的血和有酵之物一同獻上。逾越節的祭牲也不可留到早晨。
EXOD|34|26|土地裏上好的初熟之物要奉到耶和華－你上帝的殿。不可用母山羊的奶來煮牠的小山羊。」
EXOD|34|27|耶和華對 摩西 說：「你要將這些話寫上，因為我按這話與你和 以色列 人立約。」
EXOD|34|28|摩西 在耶和華那裏四十晝夜，不吃飯不喝水。他把這約的話，那十條誡命 ，寫在版上。
EXOD|34|29|摩西 下 西奈山 。 摩西 從山上下來的時候，手裏拿著兩塊法版。 摩西 不知道自己臉上的皮膚因耶和華和他說話而發光。
EXOD|34|30|亞倫 和 以色列 眾人看見 摩西 ，看哪，他臉上的皮膚發光，他們就怕靠近他。
EXOD|34|31|摩西 叫他們來， 亞倫 和會眾的官長回到他那裏， 摩西 就跟他們說話。
EXOD|34|32|隨後 以色列 眾人都近前來，他就把耶和華在 西奈山 與他所說的一切話都吩咐他們。
EXOD|34|33|摩西 跟他們說完了話，就用面紗蒙上臉。
EXOD|34|34|但 摩西 進到耶和華面前與他說話的時候，就把面紗揭下，直到出來。 摩西 出來，將所吩咐他的話告訴 以色列 人。
EXOD|34|35|以色列 人看見 摩西 的臉，他臉上的皮膚發光。 摩西 就用面紗蒙上臉，直到他進去與耶和華說話才揭下。
EXOD|35|1|摩西 召集 以色列 全會眾，對他們說：「這是耶和華吩咐你們遵行的事：
EXOD|35|2|六日要做工，第七日你們要奉為向耶和華守完全安息的安息聖日。凡在這日做工的，要被處死。
EXOD|35|3|在安息日這一天，不可在你們一切的住處生火。」
EXOD|35|4|摩西 對 以色列 全會眾說：「這是耶和華所吩咐的話，說：
EXOD|35|5|要從你們當中拿禮物獻給耶和華；凡甘心樂意的，可以把耶和華的禮物拿來，就是金、銀、銅，
EXOD|35|6|藍色、紫色、朱紅色紗，細麻，山羊毛，
EXOD|35|7|染紅的公羊皮，精美的皮料，金合歡木，
EXOD|35|8|點燈的油，做膏油的香料、做香的香料，
EXOD|35|9|紅瑪瑙與寶石，可以鑲嵌在以弗得和胸袋上。」
EXOD|35|10|「你們當中凡心裏有智慧的都要來，製造一切耶和華所吩咐的，
EXOD|35|11|就是帳幕、帳幕的罩棚、帳幕的蓋、鉤子、豎板、橫木、柱子和帶卯眼的座，
EXOD|35|12|櫃子、櫃子的槓、櫃蓋和遮掩的幔子，
EXOD|35|13|供桌、供桌的槓、供桌一切的器具和供餅，
EXOD|35|14|燈臺、燈臺的器具、燈和點燈的油，
EXOD|35|15|香壇、壇的槓、膏油和芬芳的香，帳幕門口的門簾，
EXOD|35|16|燔祭壇、壇的銅網、壇的槓和壇的一切器具，洗濯盆和盆座，
EXOD|35|17|院子的帷幔、柱子、帶卯眼的座和院子的門簾，
EXOD|35|18|帳幕的橛子、院子的橛子和繩子，
EXOD|35|19|以及聖所事奉用的精緻禮服， 亞倫 祭司的聖衣和他兒子的衣服，供祭司職分用。」
EXOD|35|20|以色列 全會眾從 摩西 的面前出去。
EXOD|35|21|凡心受感動，靈被驅策的，都帶耶和華的禮物來，為要造會幕和其中一切的器具，以及縫製聖衣。
EXOD|35|22|凡甘心樂意的，連男帶女都來了，各將金器，就是胸針、耳環、打印的戒指，和項鏈帶來，搖著金器的搖祭獻給耶和華。
EXOD|35|23|凡有藍色、紫色、朱紅色紗、細麻、山羊毛、染紅的公羊皮、精美皮料的，都拿了來；
EXOD|35|24|凡願意獻銀和銅作禮物的，都拿禮物來獻給耶和華；凡有金合歡木可做各種用途的也都拿了來。
EXOD|35|25|凡心中有智慧，可以親手紡織的婦女，也把所紡的藍色、紫色、朱紅色紗，和細麻都拿了來。
EXOD|35|26|凡有智慧，心裏受感動的婦女都來紡山羊毛。
EXOD|35|27|眾官長把紅瑪瑙和寶石，可以鑲嵌在以弗得與胸袋上的，都拿了來，
EXOD|35|28|又拿做香，做膏油，和點燈所需的香料和油來。
EXOD|35|29|以色列 人，無論男女，凡心裏受感動的，都帶甘心祭來獻給耶和華，為要做耶和華藉 摩西 所吩咐的一切工。
EXOD|35|30|摩西 對 以色列 人說：「看， 猶大 支派中 戶珥 的孫子， 烏利 的兒子 比撒列 ，耶和華已經題名召他，
EXOD|35|31|又以上帝的靈充滿他，使他有智慧、聰明、知識，能做各樣的工，
EXOD|35|32|能設計圖案，用金、銀、銅製造各物，
EXOD|35|33|又能雕刻鑲嵌用的寶石，雕刻木頭，做各樣精巧的工。
EXOD|35|34|耶和華又賜給他和 但 支派中， 亞希撒抹 的兒子 亞何利亞伯 能教導人的心。
EXOD|35|35|耶和華使他們的心滿有智慧，能做各樣的工，無論是雕刻的工，圖案設計的工，用藍色、紫色、朱紅色紗，和細麻作刺繡的工，以及編織的工，他們都能勝任，也能設計圖案。」
EXOD|36|1|比撒列 和 亞何利亞伯 ，以及一切心裏有智慧，蒙耶和華賜智慧和聰明，懂得做聖所各樣用途之工的人，都照耶和華所吩咐的去做。
EXOD|36|2|摩西 把 比撒列 和 亞何利亞伯 ，以及那些蒙耶和華賜他心裏有智慧，心受感動願意前來做工的人都召來。
EXOD|36|3|這些人就從 摩西 收了 以色列 人為建造聖所，以及聖所各用途之工而奉獻的禮物。每天早晨，百姓繼續把甘心祭拿來。
EXOD|36|4|凡有智慧能做聖所一切工的人，都各自離開他們原本的工作前來，
EXOD|36|5|對 摩西 說：「百姓送來的禮物很多，已經超過耶和華吩咐建造之工所需要的了。」
EXOD|36|6|摩西 吩咐，他們就在營中傳令說：「無論男女，不必再為聖所的禮物做任何的工。」這樣才使百姓停止，不再拿禮物來，
EXOD|36|7|他們所有的材料已經足夠整個工程之用，而且有餘。
EXOD|36|8|做工的人當中，凡心裏有智慧的，用十幅幔子做帳幕，幔子是用搓的細麻和藍色、紫色、朱紅色紗織成的，並且以刺繡的手藝繡上基路伯。
EXOD|36|9|每幅幔子長二十八肘，每幅幔子寬四肘，全部的幔子都是一樣的尺寸。
EXOD|36|10|他使這五幅幔子彼此相連，又使那五幅幔子彼此相連。
EXOD|36|11|他在這一組相連幔子的末幅邊上縫了藍色的鈕環；在另一組相連幔子的末幅邊上也照樣做。
EXOD|36|12|他在這幅幔子上縫五十個鈕環，在另一組相連幔子的末幅上也縫五十個鈕環，環環相對。
EXOD|36|13|他又做了五十個金鉤，用鉤子使幔子彼此相連，成為一個帳幕。
EXOD|36|14|他用山羊毛織十一幅幔子，作為帳幕上的罩棚。
EXOD|36|15|每幅幔子長三十肘，每幅幔子寬四肘；十一幅幔子都是一樣的尺寸。
EXOD|36|16|他把五幅幔子連成一幅，又把六幅幔子連成一幅。
EXOD|36|17|他在這一組相連幔子的末幅邊上縫了五十個鈕環；在另一組相連幔子的末幅邊上也縫了五十個鈕環。
EXOD|36|18|他又做五十個銅鉤，使罩棚相連成為一個。
EXOD|36|19|他用染紅的公羊皮做罩棚的蓋，再用精美皮料做外層的蓋。
EXOD|36|20|他用金合歡木做豎立帳幕的木板，
EXOD|36|21|木板長十肘，每塊板寬一肘半，
EXOD|36|22|每塊板有兩個榫頭可以彼此銜接。帳幕一切的板都是這樣做。
EXOD|36|23|他做帳幕的木板：南面，就是面向南方的那一邊，做二十塊板，
EXOD|36|24|在這二十塊板底下做了四十個帶卯眼的銀座：兩個卯眼接連這塊板上的兩個榫頭，另外兩個卯眼接連那塊板上的兩個榫頭。
EXOD|36|25|他在帳幕的第二邊，就是北面，也做二十塊板，
EXOD|36|26|和四十個帶卯眼的銀座；這塊板底下有兩個卯眼，那塊板底下也有兩個卯眼。
EXOD|36|27|他在帳幕的後面，就是西面，做六塊板，
EXOD|36|28|在帳幕後面的角落做兩塊板。
EXOD|36|29|下端的板是成雙的，上端連在一起，直到頂端的第一個環子；兩塊板都是這樣，做成兩個角落。
EXOD|36|30|一共有八塊板和十六個帶卯眼的銀座，每塊板底下有兩個卯眼。
EXOD|36|31|他用金合歡木做橫木：為帳幕這面的板做五根橫木，
EXOD|36|32|為帳幕那面的板做五根橫木，又為帳幕後面，就是朝西的板做五根橫木，
EXOD|36|33|他做了板腰間的橫木，從一頭通到另一頭。
EXOD|36|34|他將板包上金子，又做板上的金環來套橫木；橫木也包上金子。
EXOD|36|35|他用藍色、紫色、朱紅色紗，和搓的細麻織幔子，以刺繡的手藝繡上基路伯。
EXOD|36|36|他又用金合歡木為幔子做四根柱子，包上金子，柱子有金鉤，又為柱子鑄了四個帶卯眼的銀座。
EXOD|36|37|他用藍色、紫色、朱紅色紗，和搓的細麻，以刺繡的手藝為帳幕織門簾，
EXOD|36|38|又為簾子做五根柱子和柱子的鉤子，把柱頂和柱子的箍包上金子。柱子有五個帶卯眼的銅座。
EXOD|37|1|比撒列 用金合歡木做一個櫃子，長二肘半，寬一肘半，高一肘半。
EXOD|37|2|裏裏外外包上金子，四圍鑲上金邊。
EXOD|37|3|他又鑄了四個金環，安在櫃子的四腳上；這邊兩個環，那邊兩個環。
EXOD|37|4|他用金合歡木做了兩根槓，包上金子，
EXOD|37|5|又把槓穿過櫃旁的環，以便抬櫃。
EXOD|37|6|他用純金做了一個櫃蓋，長二肘半，寬一肘半，
EXOD|37|7|他造兩個用金子錘出的基路伯，從櫃蓋的兩端錘出它們。
EXOD|37|8|這端一個基路伯，那端一個基路伯；從櫃蓋的兩端錘出兩個基路伯。
EXOD|37|9|二基路伯的翅膀向上張開，用翅膀遮住櫃蓋，臉彼此相對；基路伯的臉朝向櫃蓋。
EXOD|37|10|他用金合歡木做了一張供桌，長二肘，寬一肘，高一肘半，
EXOD|37|11|把它包上純金，四圍鑲上金邊。
EXOD|37|12|供桌的四圍各做了一掌寬的邊緣，邊緣鑲上金邊。
EXOD|37|13|他又鑄了四個金環，把環安在四個桌腳的四角上。
EXOD|37|14|環靠近邊緣，以便穿槓抬供桌。
EXOD|37|15|他用金合歡木做了兩根槓，包上金子，用來抬供桌。
EXOD|37|16|他又用純金做了桌上的器具，就是盤、碟，以及澆酒祭的杯和壺。
EXOD|37|17|他造一座用純金錘出的燈臺；燈臺的座、幹、杯、花萼和花瓣，都和燈臺接連一塊。
EXOD|37|18|燈臺兩旁伸出六根枝子：這邊三根，那邊三根。
EXOD|37|19|這邊的枝子上有三個杯，形狀像杏花，有花萼有花瓣；那邊的枝子上也有三個杯，形狀像杏花，有花萼有花瓣。從燈臺伸出來的六根枝子都是如此。
EXOD|37|20|燈臺本身有四個杯，形狀像杏花，有花萼有花瓣。
EXOD|37|21|燈臺的第一對枝子下面有花萼，燈臺的第二對枝子下面有花萼，燈臺的第三對枝子下面也有花萼；燈臺伸出的六根枝子都是如此。
EXOD|37|22|花萼和枝子都和燈臺接連一塊，全是從一塊純金錘出來的。
EXOD|37|23|他用純金做燈臺的七盞燈，以及燈剪和燈盤。
EXOD|37|24|他用一他連得的純金做燈臺和燈臺的一切器具。
EXOD|37|25|他用金合歡木做香壇，長一肘，寬一肘，這壇是正方形的，高二肘。壇的四個翹角與壇接連一塊。
EXOD|37|26|他把壇的上面與壇的四圍，以及壇的四個翹角包上純金，又在壇的四圍鑲上金邊。
EXOD|37|27|他在壇的兩個對側，金邊下面做了兩個金環，用來穿槓抬壇。
EXOD|37|28|他又用金合歡木做槓，包上金子。
EXOD|37|29|他按配製香料的方法製成聖膏油和芬芳的純香。
EXOD|38|1|他用金合歡木做燔祭壇，長五肘，寬五肘，是正方形的，高三肘。
EXOD|38|2|在壇的四角做四個翹角，與壇接連一塊，把壇包上銅。
EXOD|38|3|他做壇的一切器具，就是桶子、鏟子、盤子、肉叉和火盆；這一切器具都是用銅做的。
EXOD|38|4|他又為壇做一個銅網，安在壇四圍的邊的下面，垂到壇的半腰。
EXOD|38|5|他在銅網的四角上鑄了四個環，用來穿槓。
EXOD|38|6|他用金合歡木做槓，包上銅，
EXOD|38|7|把槓穿過壇兩旁的環子，用來抬壇。他用板做壇，壇的中心是空的。
EXOD|38|8|他用銅做洗濯盆和盆座，是用會幕門前事奉之婦人的銅鏡做的。
EXOD|38|9|他又做院子，在南面，就是面向南方的那一邊，用搓的細麻做院子的帷幔，一百肘。
EXOD|38|10|帷幔有二十根柱子，二十個帶卯眼的銅座；柱子的鉤和箍都是銀的。
EXOD|38|11|北面的帷幔一百肘。帷幔有二十根柱子，二十個帶卯眼的銅座；柱子的鉤和箍都是銀的。
EXOD|38|12|西面的帷幔五十肘。帷幔有十根柱子，十個帶卯眼的座；柱子的鉤和箍都是銀的。
EXOD|38|13|院子的東面，就是面向東方的那一邊，五十肘。
EXOD|38|14|一邊的帷幔有十五肘，有三根柱子，三個帶卯眼的座。
EXOD|38|15|另一邊也一樣，院子門口左右的帷幔也有十五肘，有三根柱子，三個帶卯眼的座。
EXOD|38|16|院子四面的帷幔都是用搓的細麻做的。
EXOD|38|17|柱子帶卯眼的座是銅的，柱子的鉤和箍是銀的，柱頂是用銀包的。院子一切的柱子都是用銀子箍著的。
EXOD|38|18|院子的門簾是以刺繡的手藝，用藍色、紫色、朱紅色紗，和搓的細麻織的，長二十肘，寬也就是高五肘，與院子帷幔的高度相同。
EXOD|38|19|門簾有四根柱子，四個帶卯眼的銅座；柱子上的鉤和箍是銀的，柱頂是用銀包的。
EXOD|38|20|帳幕一切的橛子和院子四圍的橛子都是銅的。
EXOD|38|21|這是帳幕，就是法櫃帳幕中物件的總數，是照 摩西 的吩咐， 亞倫 祭司的兒子 以他瑪 經手， 利未 人數點的。
EXOD|38|22|凡耶和華吩咐 摩西 的，都是由 猶大 支派中 戶珥 的孫子， 烏利 的兒子 比撒列 去做的；
EXOD|38|23|與他同工的有 但 支派中 亞希撒抹 的兒子 亞何利亞伯 ；他是雕刻師，也是設計師，又是用藍色、紫色、朱紅色紗，和細麻的刺繡師。
EXOD|38|24|為聖所一切工作用的金子，就是所奉獻的金子，按聖所的舍客勒，一共是二十九他連得，七百三十舍客勒。
EXOD|38|25|會中被數的人所獻的銀子，按聖所的舍客勒，一共是一百他連得，一千七百七十五舍客勒。
EXOD|38|26|凡曾被數的，就是二十歲以上的人，共有六十萬三千五百五十人。按聖所的舍客勒，每人半舍客勒，就是一比加。
EXOD|38|27|一百他連得銀子是用來鑄造聖所帶卯眼的座和幔子下帶卯眼的座；用一百他連得鑄造一百個帶卯眼的座，每個帶卯眼的座一他連得。
EXOD|38|28|一千七百七十五舍客勒是用來鑄造柱子的鉤，包柱頂，以及箍著柱子。
EXOD|38|29|所奉獻的銅共有七十他連得，二千四百舍客勒。
EXOD|38|30|這些銅是用來做會幕門口帶卯眼的座，銅壇、壇的銅網和壇的一切器具，
EXOD|38|31|院子四圍帶卯眼的座和院子門口帶卯眼的座，以及帳幕一切的橛子和院子四圍所有的橛子。
EXOD|39|1|他們用藍色、紫色、朱紅色紗縫製精緻的禮服，在聖所用以供職；他們為 亞倫 做聖衣，是照耶和華所吩咐 摩西 的。
EXOD|39|2|以弗得是用金色、藍色、紫色、朱紅色紗，和搓的細麻做的。
EXOD|39|3|他們把金子錘成薄片，剪成細線，與藍色、紫色、朱紅色紗，以刺繡的手藝織在一起。
EXOD|39|4|他們又為以弗得做兩條相連的肩帶，接連在以弗得的兩端。
EXOD|39|5|以弗得的精緻帶子以一樣的手藝，用金色、藍色、紫色、朱紅色紗，和搓的細麻縫製，與以弗得接連在一起，是照耶和華所吩咐 摩西 的。
EXOD|39|6|他們琢出兩塊紅瑪瑙，鑲在金槽裏，如同刻印章，刻上 以色列 眾子的名字。
EXOD|39|7|他把這兩塊寶石安在以弗得的兩條肩帶上，為 以色列 人作紀念石，是照耶和華所吩咐 摩西 的。
EXOD|39|8|胸袋是以刺繡的手藝，如同以弗得的做法，用金色、藍色、紫色、朱紅色紗，和搓的細麻縫製。
EXOD|39|9|胸袋是正方形的，他們把它做成兩層，這兩層各長一虎口，寬一虎口。
EXOD|39|10|他們在上面鑲四行寶石：第一行是紅寶石、紅璧璽、紅玉；
EXOD|39|11|第二行是綠寶石、藍寶石、金剛石；
EXOD|39|12|第三行是紫瑪瑙、白瑪瑙、紫晶；
EXOD|39|13|第四行是水蒼玉、紅瑪瑙、碧玉。這些都鑲在金槽中。
EXOD|39|14|這些寶石有 以色列 十二個兒子的名字，如同刻印章，每一顆有自己的名字，代表十二個支派。
EXOD|39|15|他們在胸袋上用純金打鏈子，像編成的繩子一樣。
EXOD|39|16|他們又做了兩個金槽和兩個金環，把這兩個環安在胸袋的兩端。
EXOD|39|17|他們把那兩條編成的金鏈繫在胸袋兩端的兩個環上，
EXOD|39|18|又把鏈子的另外兩端扣在兩個槽上，安在以弗得前面的肩帶上。
EXOD|39|19|他們做了兩個金環，安在胸袋的兩端，在以弗得裏面的邊上，
EXOD|39|20|又做兩個金環，安在以弗得前面兩條肩帶的下邊，靠近接縫處，在精緻帶子的上面。
EXOD|39|21|他們用藍色的帶子把胸袋的環與以弗得的環繫住，使胸袋綁在以弗得精緻的帶子上，不致鬆脫，是照耶和華所吩咐 摩西 的。
EXOD|39|22|以弗得的外袍是以編織的手藝做的，顏色全是藍的。
EXOD|39|23|袍上方的中間留了一個領口，領口的周圍織出領邊，好像鎧甲的領口，免得破裂。
EXOD|39|24|他們在袍子下襬用藍色、紫色、朱紅色紗，和搓的細麻 做石榴，
EXOD|39|25|又用純金鑄了鈴鐺，把鈴鐺釘在石榴中間，袍子下襬周圍的石榴中間：
EXOD|39|26|一個鈴鐺一個石榴，一個鈴鐺一個石榴，在袍子下襬的周圍，用以供職，是照耶和華所吩咐 摩西 的。
EXOD|39|27|他們用編織的工為 亞倫 和他的兒子做細麻布內袍、
EXOD|39|28|細麻布禮冠、細麻布精緻頭巾，和搓的細麻布褲子，
EXOD|39|29|又用藍色、紫色、朱紅色紗，和搓的細麻，以刺繡的手藝做腰帶，是照耶和華所吩咐 摩西 的。
EXOD|39|30|他們用純金做一面聖冠上的牌，如同刻印章，在上面寫著「歸耶和華為聖」，
EXOD|39|31|又用藍色的帶子把牌繫在禮冠上，是照耶和華所吩咐 摩西 的。
EXOD|39|32|會幕的帳幕一切的工程就這樣做完了。凡耶和華所吩咐 摩西 的， 以色列 人都照樣做了。
EXOD|39|33|他們把帳幕運到 摩西 那裏，帳幕和帳幕的一切器具，就是鉤、板、橫木、柱子、帶卯眼的座，
EXOD|39|34|染紅公羊皮的蓋、精美皮料的蓋、遮掩的幔子，
EXOD|39|35|法櫃、櫃的槓、櫃蓋，
EXOD|39|36|供桌、供桌的一切器具、供餅，
EXOD|39|37|純金的燈臺、擺列的燈、燈臺的一切器具、點燈的油，
EXOD|39|38|金壇、膏油、芬芳的香、帳幕的門簾，
EXOD|39|39|銅壇、壇的銅網、壇的槓、壇的一切器具，洗濯盆和盆座，
EXOD|39|40|院子的帷幔、柱子、帶卯眼的座、院子的門簾、繩子、橛子，帳幕，就是會幕使用的一切器具，
EXOD|39|41|以及聖所事奉用的精緻禮服， 亞倫 祭司的聖衣和他兒子的衣服，供祭司職分用。
EXOD|39|42|這一切工作都是 以色列 人照耶和華所吩咐 摩西 做的。
EXOD|39|43|摩西 看見這一切的工，看哪，耶和華怎樣吩咐，他們就照樣做了， 摩西 就為他們祝福。
EXOD|40|1|耶和華吩咐 摩西 說：
EXOD|40|2|「正月初一，你要立起會幕的帳幕，
EXOD|40|3|把法櫃安放在裏面，用幔子將櫃遮掩。
EXOD|40|4|把供桌搬進去，擺設桌上的器具。又把燈臺搬進去，點上燈。
EXOD|40|5|把金香壇安在法櫃前，掛上帳幕的門簾。
EXOD|40|6|把燔祭壇安在會幕的帳幕門前。
EXOD|40|7|把洗濯盆安在會幕和壇的中間，在盆裏盛水。
EXOD|40|8|又要在院子周圍支起帷幔，把院子的門簾掛上。
EXOD|40|9|你要用膏油抹帳幕和其中所有的，使帳幕和一切器具分別為聖，就都成為聖。
EXOD|40|10|又要抹燔祭壇和壇的一切器具，使壇分別為聖，壇就成為至聖。
EXOD|40|11|要抹洗濯盆和盆座，使盆分別為聖。
EXOD|40|12|你要帶 亞倫 和他兒子到會幕門口，用水洗身。
EXOD|40|13|要給 亞倫 穿上聖衣，又膏他，使他分別為聖，作事奉我的祭司。
EXOD|40|14|又要帶他的兒子來，給他們穿上內袍。
EXOD|40|15|你怎樣膏他們的父親，也要照樣膏他們，使他們成為事奉我的祭司。他們受了膏，就必世世代代永遠得祭司的職分。」
EXOD|40|16|摩西 這樣做了；耶和華怎樣吩咐 摩西 ，他就照樣做了。
EXOD|40|17|第二年正月初一，帳幕就立起來。
EXOD|40|18|摩西 支起帳幕，安上帶卯眼的座，安上板，穿上橫木，立起柱子。
EXOD|40|19|他在帳幕的上面搭上罩棚，把罩棚外層的蓋子蓋在其上，是照著耶和華所吩咐他的。
EXOD|40|20|他把法版放在櫃裏，把槓穿在櫃的兩旁，把櫃蓋安在櫃上。
EXOD|40|21|把櫃抬進帳幕，掛上遮掩櫃的幔子，把法櫃遮蓋了，是照耶和華所吩咐 摩西 的。
EXOD|40|22|他把供桌安在會幕內，在帳幕的北邊，幔子的外面。
EXOD|40|23|把餅擺設在供桌上，在耶和華面前，是照耶和華所吩咐 摩西 的。
EXOD|40|24|他把燈臺安在會幕內，在帳幕的南邊，供桌的對面，
EXOD|40|25|並在耶和華面前點燈，是照耶和華所吩咐 摩西 的。
EXOD|40|26|他把金壇安在會幕內，幔子的前面，
EXOD|40|27|又在壇上燒芬芳的香，是照耶和華所吩咐 摩西 的。
EXOD|40|28|他又掛上帳幕的門簾。
EXOD|40|29|在會幕的帳幕門口安設燔祭壇，把燔祭和素祭獻在壇上，是照耶和華所吩咐 摩西 的。
EXOD|40|30|他又把洗濯盆安在會幕和祭壇的中間，盆裏盛水，以便洗濯。
EXOD|40|31|摩西 和 亞倫 ，以及 亞倫 的兒子用這盆洗手洗腳。
EXOD|40|32|他們進會幕或走近壇的時候，就都洗濯，是照耶和華所吩咐 摩西 的。
EXOD|40|33|他在帳幕和祭壇的四圍支起院子的帷幔，把院子的門簾掛上。這樣， 摩西 就做完了工。
EXOD|40|34|那時，雲彩遮蓋會幕，耶和華的榮光充滿了帳幕。
EXOD|40|35|摩西 不能進會幕，因為雲彩停在其上，耶和華的榮光充滿了帳幕。
EXOD|40|36|每逢雲彩從帳幕升上去， 以色列 人就起程前行；
EXOD|40|37|雲彩若不升上去，他們就不起程，直等到雲彩升上去。
EXOD|40|38|在他們所行的路上，在 以色列 全家的眼前，白天，耶和華的雲彩在帳幕上，黑夜，有火在雲彩中。
LEV|1|1|耶和華從會幕中呼叫 摩西 ，吩咐他說：
LEV|1|2|「你要吩咐 以色列 人，對他們說：你們中間若有人要獻供物給耶和華，可以從牛群羊群中獻牲畜為供物。
LEV|1|3|「他的供物若以牛為燔祭，要獻一頭沒有殘疾的公牛，獻在會幕的門口，他就可以在耶和華面前蒙悅納。
LEV|1|4|他要按手在燔祭牲的頭上，為自己贖罪，就蒙悅納。
LEV|1|5|他要在耶和華面前宰公牛犢； 亞倫 子孫作祭司的要獻上血，把血灑在會幕門口壇的周圍。
LEV|1|6|他要剝去燔祭牲的皮，把燔祭牲切成塊。
LEV|1|7|亞倫 祭司的子孫要在壇上生火，把柴擺在火上。
LEV|1|8|亞倫 子孫作祭司的要把肉塊連頭和脂肪，擺在壇上燒著火的柴上。
LEV|1|9|燔祭牲的內臟與小腿要用水洗淨，祭司要把整隻全燒在壇上，當作燔祭，是獻給耶和華為馨香的火祭。
LEV|1|10|「人的供物若以綿羊或山羊為燔祭，要獻一隻沒有殘疾的公羊。
LEV|1|11|他要在壇的北邊，在耶和華面前宰羊； 亞倫 子孫作祭司的要把血灑在壇的周圍。
LEV|1|12|他要把燔祭牲切成塊，祭司就要把肉塊連頭和脂肪，擺在壇上燒著火的柴上。
LEV|1|13|內臟與小腿要用水洗淨，祭司要把整隻獻上，全燒在壇上。這是燔祭，是獻給耶和華為馨香的火祭。
LEV|1|14|「人獻給耶和華的供物若以鳥為燔祭，就要獻斑鳩或雛鴿為他的供物。
LEV|1|15|祭司要把鳥拿到壇前，扭斷牠的頭，把鳥燒在壇上，鳥的血要流在壇的旁邊；
LEV|1|16|又要把鳥的嗉囊和裏面的髒物 除掉，丟在壇東邊倒灰的地方。
LEV|1|17|他要拿著鳥的兩個翅膀，把鳥撕開，卻不可撕斷；祭司要把牠擺在壇上燒著火的柴上焚燒。這是燔祭，是獻給耶和華為馨香的火祭。」
LEV|2|1|「若有人獻素祭為供物給耶和華，就要獻細麵為供物，把油澆在上面，加上乳香，
LEV|2|2|帶到 亞倫 子孫作祭司的那裏。祭司要從細麵中取出滿滿的一把，又取些油和所有的乳香，把這些作為紀念的燒在壇上，是獻給耶和華為馨香的火祭。
LEV|2|3|素祭所剩的要歸給 亞倫 和他的子孫；在獻給耶和華的火祭中，這是至聖的。
LEV|2|4|「若獻爐中烤的素祭為供物，要用調了油的無酵細麵餅，或抹了油的無酵薄餅。
LEV|2|5|若以鐵盤上的素祭為供物，就要用調了油的無酵細麵，
LEV|2|6|分成小塊，澆上油；這是素祭。
LEV|2|7|若以煎鍋煎的素祭為供物，就要用油與細麵做成。
LEV|2|8|要把這樣做成的素祭帶到耶和華面前，拿給祭司，祭司要帶到壇前。
LEV|2|9|祭司要從素祭中取出作為紀念的燒在壇上，是獻給耶和華為馨香的火祭。
LEV|2|10|素祭所剩的要歸給 亞倫 和他的子孫；在獻給耶和華的火祭中，這是至聖的。
LEV|2|11|「凡獻給耶和華的素祭都不可以有酵，因為你們不可把任何的酵或蜜燒了，當作火祭獻給耶和華。
LEV|2|12|你們可以把這些獻給耶和華當作初熟的供物，但是不可獻在壇上作為馨香的祭。
LEV|2|13|凡獻為素祭的供物都要用鹽調和；在素祭中，不可缺少你與上帝立約的鹽。一切的供物都要加鹽獻上。
LEV|2|14|「你若獻初熟之物給耶和華為素祭，就要獻在火中烘過的新麥穗，就是磨碎的新穀物，當作初熟之物的素祭。
LEV|2|15|你要加上油和乳香；這是素祭。
LEV|2|16|祭司要把供物中作為紀念的，就是一些磨碎的新穀物和一些油，以及所有的乳香，都焚燒，是獻給耶和華的火祭。」
LEV|3|1|「人獻平安祭為供物，若是從牛群中獻，無論是公的母的，要用沒有殘疾的，獻在耶和華面前。
LEV|3|2|他要按手在供物的頭上，在會幕的門口宰了牠。 亞倫 子孫作祭司的，要把血灑在壇的周圍。
LEV|3|3|從平安祭中，他要把火祭獻給耶和華，就是包著內臟的脂肪和內臟上所有的脂肪，
LEV|3|4|兩個腎和腎上的脂肪，即靠近腎兩旁的脂肪，以及肝上的網油，連同腎一起取下。
LEV|3|5|亞倫 的子孫要把這些擺在燒著火的柴上，燒在壇的燔祭上，是獻給耶和華為馨香的火祭。
LEV|3|6|「人向耶和華獻平安祭為供物，若是從羊群中獻，無論是公的母的，要用沒有殘疾的。
LEV|3|7|若他獻一隻綿羊為供物，就要把牠獻在耶和華面前。
LEV|3|8|要按手在供物的頭上，在會幕前宰了牠。 亞倫 的子孫要把血灑在壇的周圍。
LEV|3|9|從平安祭中，他要取脂肪當作火祭獻給耶和華，就是靠近脊骨處取下的整條肥尾巴，包著內臟的脂肪和內臟上所有的脂肪，
LEV|3|10|兩個腎和腎上的脂肪，即靠近腎兩旁的脂肪，以及肝上的網油，連同腎一起取下。
LEV|3|11|祭司要把這些燒在壇上，是獻給耶和華為食物的火祭。
LEV|3|12|「人的供物若是山羊，就要把牠獻在耶和華面前。
LEV|3|13|要按手在牠的頭上，在會幕前宰了牠。 亞倫 的子孫要把血灑在壇的周圍，
LEV|3|14|又要從供物中把火祭獻給耶和華，就是包著內臟的脂肪和內臟上所有的脂肪，
LEV|3|15|兩個腎和腎上的脂肪，即靠近腎兩旁的脂肪，以及肝上的網油，連同腎一起取下。
LEV|3|16|祭司要把這些燒在壇上，作為馨香火祭的食物；所有的脂肪都是耶和華的。
LEV|3|17|在你們一切的住處，脂肪和血都不可吃，這要成為你們世世代代永遠的定例。」
LEV|4|1|耶和華吩咐 摩西 說：
LEV|4|2|「你要吩咐 以色列 人說：若有人無意中犯罪，在任何事上犯了一條耶和華所吩咐的禁令，
LEV|4|3|或是受膏的祭司犯了罪，使百姓陷在罪裏，他就當為自己所犯的罪，把沒有殘疾的公牛犢獻給耶和華為贖罪祭。
LEV|4|4|他要把公牛牽到會幕的門口，在耶和華面前按手在牛的頭上，把牛宰於耶和華面前。
LEV|4|5|受膏的祭司要取些公牛的血，帶到會幕那裏。
LEV|4|6|祭司要把手指蘸在血中，在耶和華面前對著聖所的幔子彈血七次，
LEV|4|7|又要把一些血抹在會幕內，耶和華面前香壇的四個翹角上，再把公牛其餘的血全倒在會幕門口燔祭壇的底座上；
LEV|4|8|又要取出這頭贖罪祭公牛所有的脂肪，就是包著內臟的脂肪和內臟上所有的脂肪，
LEV|4|9|兩個腎和腎上的脂肪，即靠近腎兩旁的脂肪，以及肝上的網油，連同腎一起取下，
LEV|4|10|正如從平安祭的牛身上所取的，祭司要把這些燒在燔祭壇上。
LEV|4|11|但公牛的皮和所有的肉，以及頭、腿、內臟、糞，
LEV|4|12|就是全公牛，要搬到營外清潔的地方倒灰之處，放在柴上用火焚燒。
LEV|4|13|「 以色列 全會眾若犯了錯，在任何事上犯了一條耶和華所吩咐的禁令，而有了罪，會眾看不出這隱藏的事；
LEV|4|14|他們一知道犯了罪，就要獻一頭公牛犢為贖罪祭，牽牠到會幕前。
LEV|4|15|會眾的長老要在耶和華面前按手在公牛的頭上，把牛宰於耶和華面前。
LEV|4|16|受膏的祭司要取些公牛的血，帶到會幕那裏。
LEV|4|17|祭司要用手指蘸一些血，在耶和華面前對著幔子彈七次，
LEV|4|18|又要把一些血抹在會幕內，耶和華面前壇的四個翹角上，再把其餘的血全倒在會幕門口燔祭壇的底座上。
LEV|4|19|他要取出公牛所有的脂肪，燒在壇上。
LEV|4|20|他要處理這牛，正如處理那頭贖罪祭的公牛一樣，他要如此去做。祭司要為他們贖罪，他們就蒙赦免。
LEV|4|21|他要把牛搬到營外燒了，像燒前一頭公牛一樣；這是會眾的贖罪祭。
LEV|4|22|「官長若犯罪，在任何事上無意中犯了一條耶和華－他的上帝所吩咐的禁令，而有了罪，
LEV|4|23|他一知道自己犯了罪，就要牽一隻沒有殘疾的公山羊為供物。
LEV|4|24|他要按手在羊的頭上，在耶和華面前宰燔祭牲的地方把牠宰了；這是贖罪祭。
LEV|4|25|祭司要用手指蘸一些贖罪祭牲的血，抹在燔祭壇的四個翹角上，再把其餘的血倒在燔祭壇的底座上。
LEV|4|26|祭牲所有的脂肪都要燒在壇上，正如平安祭的脂肪一樣。祭司要為他的罪贖了他，他就蒙赦免。
LEV|4|27|「這地的百姓若有人無意中犯罪，在任何事上犯了一條耶和華所吩咐的禁令，而有了罪，
LEV|4|28|他一知道自己犯了罪，就要為所犯的罪牽一隻沒有殘疾的母山羊為供物。
LEV|4|29|他要按手在贖罪祭牲的頭上，在燔祭牲的地方把牠宰了。
LEV|4|30|祭司要用手指蘸一些祭牲的血，抹在燔祭壇的四個翹角上，再把其餘的血全倒在壇的底座上；
LEV|4|31|又要把祭牲所有的脂肪都取下，正如取平安祭牲的脂肪一樣。祭司要把脂肪燒在壇上，在耶和華面前作為馨香的祭。祭司要為他贖罪，他就蒙赦免。
LEV|4|32|「人若牽一隻綿羊為贖罪祭作供物，就要牽一隻沒有殘疾的母羊。
LEV|4|33|他要按手在贖罪祭牲的頭上，在宰燔祭牲的地方宰了牠，作為贖罪祭。
LEV|4|34|祭司要用手指蘸一些贖罪祭牲的血，抹在燔祭壇的四個翹角上，再把其餘的血全倒在壇的底座上；
LEV|4|35|又要把祭牲所有的脂肪都取下，正如取平安祭的羊的脂肪一樣。祭司要按獻給耶和華火祭的條例，把脂肪燒在壇上。祭司要為他所犯的罪贖了他，他就蒙赦免。」
LEV|5|1|「若有人犯了罪，就是聽見了誓言，他本來可以作證，卻不把所看見、所知道的說出來，必須擔當他的罪孽。
LEV|5|2|若有人摸了任何不潔之物，無論是野獸的不潔屍體，家畜的不潔屍體，或是群聚動物的不潔屍體，他雖不察覺，也是不潔淨，就有罪了。
LEV|5|3|或是他摸了人的不潔之物，就是任何使人成為不潔的不潔之物，他雖不察覺，但一知道，就有罪了。
LEV|5|4|若有人隨口發誓，或出於惡意，或出於善意，這人無論在甚麼事上隨意發誓，雖不察覺，但一知道，就在這其中的一件事上有罪了。
LEV|5|5|當他在這其中的一件事上有罪的時候，就要承認所犯的罪，
LEV|5|6|並要為所犯的罪，把他的贖愆祭牲，就是羊群中的一隻母綿羊或母山羊，獻給耶和華為贖罪祭，祭司要為他的罪贖了他。
LEV|5|7|「若他的力量不夠獻一隻綿羊，就要為所犯的罪，把兩隻斑鳩或是兩隻雛鴿獻給耶和華為贖愆祭：一隻作贖罪祭，一隻作燔祭。
LEV|5|8|他要把這些帶到祭司那裏，祭司就先把贖罪祭獻上，從鳥的頸項上扭斷牠的頭，但不把鳥撕斷。
LEV|5|9|祭司要把一些贖罪祭牲的血彈在祭壇的邊上，其餘的血要倒在壇的底座上；這是贖罪祭。
LEV|5|10|他要依照條例獻第二隻鳥為燔祭。祭司要為他所犯的罪贖了他，他就蒙赦免。
LEV|5|11|「他的力量若不夠獻兩隻斑鳩或兩隻雛鴿，就要為所犯的罪把供物，就是十分之一伊法細麵，獻上為贖罪祭；不可加上油，也不可加上乳香，因為這是贖罪祭。
LEV|5|12|他要把細麵帶到祭司那裏，祭司要取出滿滿的一把，作為紀念，按照獻火祭給耶和華的條例把它燒在壇上；這是贖罪祭。
LEV|5|13|至於他在這幾件事中所犯的任何罪，祭司要為他贖了，他就蒙赦免。剩下的都歸給祭司，和素祭一樣。」
LEV|5|14|耶和華吩咐 摩西 說：
LEV|5|15|「若有人在耶和華的聖物上無意中犯了罪，有了過犯，就要獻羊群中一隻沒有殘疾的公綿羊給耶和華為贖愆祭，或依聖所的舍客勒所估定的銀子，作為贖愆祭。
LEV|5|16|他要為在聖物上的疏忽賠償，另外加五分之一，把這些都交給祭司。祭司要用贖愆祭的公綿羊為他贖罪，他就蒙赦免。
LEV|5|17|「若有人犯罪，在任何事上犯了一條耶和華所吩咐的禁令，他雖不察覺，仍算有罪，必須擔當自己的罪孽。
LEV|5|18|他要牽羊群中一隻沒有殘疾的公綿羊，或照你所估定的價值，給祭司作贖愆祭。祭司要為他贖他因不知道而無意中所犯的罪，他就蒙赦免。
LEV|5|19|這是贖愆祭；因他確實得罪了耶和華。」
LEV|6|1|耶和華吩咐 摩西 說：
LEV|6|2|「若有人犯罪，得罪了耶和華，就是在鄰舍寄託他的東西或抵押品上行詭詐，或搶奪，或欺壓鄰舍，
LEV|6|3|或是撿了失物行了詭詐，起了假誓，在人所做的任何事上犯了罪；
LEV|6|4|他既犯了罪，有了過犯，就要歸還他所搶奪的，或是因欺壓所得的，或是別人寄託他的，或是他所撿到的失物，
LEV|6|5|或是起假誓得來的任何東西，就要全數歸還，另外再加五分之一。在查出他有罪的日子，就要立刻賠還給原主。
LEV|6|6|他要獻羊群中一隻沒有殘疾的公綿羊，給耶和華為贖愆祭，或照你所估定的價值，給祭司 作贖愆祭。
LEV|6|7|祭司要在耶和華面前為他贖罪；他無論做了甚麼事，以致有了罪，都必蒙赦免。」
LEV|6|8|耶和華吩咐 摩西 說：
LEV|6|9|「你要吩咐 亞倫 和他的子孫說，燔祭的條例是這樣：燔祭要放在壇的底盤上，從晚上到天亮，壇上的火要不斷地燒著。
LEV|6|10|祭司要穿上細麻布衣服，又要把細麻布褲子穿在身上，把在壇上燒剩的燔祭灰收起來，放在壇的旁邊。
LEV|6|11|然後，他要脫去這衣服，穿上別的衣服，把灰拿到營外潔淨之處。
LEV|6|12|壇上的火要不斷地燒著，不可熄滅。每日早晨，祭司要在壇上燒柴，把燔祭擺在壇上，並燒平安祭牲的脂肪。
LEV|6|13|壇上的火要不斷地燒著，不可熄滅。」
LEV|6|14|「素祭的條例是這樣： 亞倫 的子孫要在壇前把這祭獻在耶和華面前。
LEV|6|15|祭司要從素祭中的細麵取出一把，再取些油和素祭上所有的乳香，把這些作為紀念的燒在壇上，是獻給耶和華為馨香的祭。
LEV|6|16|亞倫 和他子孫要吃素祭剩下的；要在聖處吃這無酵餅，在會幕的院子裏吃。
LEV|6|17|烤餅不可加酵。這是從獻給我的火祭中歸給他們的一份；如贖罪祭和贖愆祭一樣，這份是至聖的。
LEV|6|18|亞倫 子孫中的男丁都要吃，因為這是你們世世代代從獻給耶和華的火祭中，他們永遠應得的份。凡摸這些祭物的都要成為聖。」
LEV|6|19|耶和華吩咐 摩西 說：
LEV|6|20|「這是 亞倫 受膏的日子，他和他的子孫所要獻給耶和華的供物：十分之一伊法細麵，如他們經常獻的素祭，早晨一半，晚上一半。
LEV|6|21|要在鐵盤上用油調和，調勻後，就拿去烤。素祭烤熟了要分成小塊，作為獻給耶和華馨香的祭。
LEV|6|22|亞倫 子孫中接續他受膏為祭司的，要把這素祭獻上，全燒給耶和華。這是永遠的定例。
LEV|6|23|祭司一切的素祭要全部燒了，不可以吃。」
LEV|6|24|耶和華吩咐 摩西 說：
LEV|6|25|「你要吩咐 亞倫 和他的子孫說，贖罪祭的條例是這樣：要在耶和華面前宰燔祭牲的地方宰贖罪祭牲；這是至聖的。
LEV|6|26|獻贖罪祭的祭司要吃這祭物；要在聖處，就是在會幕的院子裏吃。
LEV|6|27|凡摸這祭肉的都要成為聖；這祭牲的血若濺在衣服上，你要在聖處洗淨那濺到血的衣服 。
LEV|6|28|煮這祭物的瓦器要打碎；若祭物是在銅器裏煮，要把這銅器擦淨，用水沖洗。
LEV|6|29|祭司中所有的男丁都可以吃；這是至聖的。
LEV|6|30|若將任何贖罪祭的血帶進會幕，為要在聖所贖罪，那肉就不可吃，要用火焚燒。」
LEV|7|1|「贖愆祭的條例是這樣：這祭是至聖的。
LEV|7|2|人在哪裏宰燔祭牲，也要在哪裏宰贖愆祭牲；其血，祭司要灑在壇的周圍。
LEV|7|3|祭司要獻上牠所有的脂肪，把肥尾巴和包著內臟的脂肪，
LEV|7|4|兩個腎和腎上的脂肪，即靠近腎兩旁的脂肪，以及肝上的網油，連同腎一起取下。
LEV|7|5|祭司要把這些燒在壇上，獻給耶和華為火祭，作為贖愆祭。
LEV|7|6|祭司中所有的男丁都可以吃這祭物，要在聖處吃；這是至聖的。
LEV|7|7|贖罪祭怎樣，贖愆祭也是怎樣，都有一樣的條例，用贖愆祭贖罪的祭司要得這祭物。
LEV|7|8|獻燔祭的祭司，無論為誰獻，所獻燔祭牲的皮要歸給那祭司，那是他的。
LEV|7|9|任何素祭，無論是在爐中烤的，用煎鍋或鐵盤做成的，都要歸給獻祭的祭司。
LEV|7|10|任何素祭，無論是用油調和的，是乾的，都要歸 亞倫 的子孫，大家均分。」
LEV|7|11|「獻給耶和華平安祭的條例是這樣：
LEV|7|12|若有人為感謝獻祭，就要把用油調和的無酵餅、抹了油的無酵薄餅，和用油調勻細麵做成的餅，與感謝祭一同獻上。
LEV|7|13|要用有酵的餅，和那為感謝而獻的平安祭，與供物一同獻上。
LEV|7|14|他要從每一種供物中拿一個餅，獻給耶和華為舉祭，是要歸給那灑平安祭牲血的祭司。
LEV|7|15|為感謝而獻的平安祭的肉，要在獻祭當天吃，一點也不可留到早晨。
LEV|7|16|若所獻的是還願祭或甘心祭，要在獻祭當天吃，剩下的，第二天也可以吃。
LEV|7|17|第三天，所剩下的祭肉要用火焚燒。
LEV|7|18|第三天若吃平安祭的肉，必不蒙悅納，所獻的也不算為祭；這祭物是不潔淨的，凡吃這祭物的，必擔當自己的罪孽。
LEV|7|19|「沾了不潔淨之物的肉就不可吃，要用火焚燒。至於其他的肉，凡潔淨的人都可以吃這肉；
LEV|7|20|但不潔淨的人若吃了獻給耶和華平安祭的肉，這人必從民中剪除。
LEV|7|21|若有人摸了不潔之物，無論是人體的不潔淨，或是不潔的牲畜，或是不潔的可憎之物 ，再吃了獻給耶和華平安祭的肉，這人必從民中剪除。」
LEV|7|22|耶和華吩咐 摩西 說：
LEV|7|23|「你要吩咐 以色列 人說：牛、綿羊、山羊的脂肪，你們都不可吃。
LEV|7|24|自然死去的或被野獸撕裂的，那脂肪可以作別的用途，你們卻萬不可吃。
LEV|7|25|任何人吃了獻給耶和華作火祭祭牲的脂肪，這人必從民中剪除。
LEV|7|26|在你們一切的住處，無論是鳥或獸的血，你們都不可吃。
LEV|7|27|無論誰吃了血，這人必從民中剪除。」
LEV|7|28|耶和華吩咐 摩西 說：
LEV|7|29|「你要吩咐 以色列 人說：獻平安祭給耶和華的，要從他的平安祭中取些供物來獻給耶和華。
LEV|7|30|他要親手把獻給耶和華的火祭帶來，要把脂肪和胸帶來，把胸在耶和華面前搖一搖，作為搖祭。
LEV|7|31|祭司要把脂肪燒在壇上，但胸要歸給 亞倫 和他的子孫。
LEV|7|32|你們要從平安祭牲中把右腿作為舉祭，送給祭司。
LEV|7|33|亞倫 子孫中獻平安祭牲的血和脂肪的，要得這右腿，作為他當得的份。
LEV|7|34|因為我從 以色列 人的平安祭中，把這搖祭的胸和這舉祭的腿給 亞倫 祭司和他子孫，作為他們在 以色列 人中永遠當得的份。」
LEV|7|35|這是從耶和華的火祭中取出，作為 亞倫 和他子孫受膏的份，就是 摩西 叫他們前來，給耶和華供祭司職分的那一天開始的。
LEV|7|36|這是在 摩西 膏他們的日子，耶和華吩咐給他們的，作為他們在 以色列 人中世世代代永遠當得的份。
LEV|7|37|這就是燔祭、素祭、贖罪祭、贖愆祭、聖職禮和平安祭的條例，
LEV|7|38|都是耶和華在 西奈山 上吩咐 摩西 的，也是他在 西奈 曠野吩咐 以色列 人獻供物給耶和華的日子所說的。
LEV|8|1|耶和華吩咐 摩西 說：
LEV|8|2|「你領 亞倫 和他兒子前來，並將聖衣、膏油，與贖罪祭的一頭公牛、兩隻公綿羊、一筐無酵餅都一同帶來；
LEV|8|3|又要召集全會眾到會幕的門口。」
LEV|8|4|摩西 就遵照耶和華的吩咐做了，於是會眾聚集在會幕的門口。
LEV|8|5|摩西 對會眾說：「這是耶和華所吩咐當做的事。」
LEV|8|6|摩西 領了 亞倫 和他兒子前來，用水洗他們。
LEV|8|7|他給 亞倫 穿上內袍，束上腰帶，套上外袍，加上以弗得，再束上精緻的帶子，把以弗得繫在他身上。
LEV|8|8|他又給 亞倫 戴上胸袋，把烏陵和土明放在胸袋內。
LEV|8|9|他把禮冠戴在 亞倫 的頭上，禮冠前面安上金牌，成為聖冕，是照耶和華所吩咐 摩西 的。
LEV|8|10|摩西 用膏油抹帳幕和其中所有的，使它們成為聖。
LEV|8|11|他又用膏油在祭壇上彈了七次，抹了壇和壇的一切器皿，以及洗濯盆和盆座，使它們成為聖。
LEV|8|12|他把膏油倒在 亞倫 的頭上膏他，使他成為聖。
LEV|8|13|摩西 帶了 亞倫 的兒子來，給他們穿上內袍，束上腰帶，裹上頭巾，是照耶和華所吩咐 摩西 的。
LEV|8|14|他把贖罪祭的公牛牽來， 亞倫 和他兒子按手在贖罪祭公牛的頭上，
LEV|8|15|就宰了公牛。 摩西 取了血，用指頭抹在祭壇周圍的四個翹角上，使壇潔淨，再把其餘的血倒在壇的底座上，使壇成為聖，為壇贖罪。
LEV|8|16|摩西 把內臟所有的脂肪和肝上的網油，以及兩個腎與腎上的脂肪取出，都燒在壇上。
LEV|8|17|至於公牛，連皮帶肉和糞，他都用火燒在營外，是照耶和華所吩咐 摩西 的。
LEV|8|18|他把燔祭的公綿羊牽來， 亞倫 和他兒子按手在羊的頭上，
LEV|8|19|就宰了公羊。 摩西 把血灑在祭壇的周圍，
LEV|8|20|把羊切成塊，把頭和肉塊，以及脂肪拿去燒，
LEV|8|21|他用水洗了內臟和腿之後，就把全羊燒在壇上，作為馨香的燔祭，是獻給耶和華的火祭，都是照耶和華所吩咐 摩西 的。
LEV|8|22|他又牽來第二隻公綿羊，就是聖職禮的羊， 亞倫 和他兒子按手在羊的頭上，
LEV|8|23|就宰了羊。 摩西 把一些血抹在 亞倫 的右耳垂上，右手的大拇指上和右腳的大腳趾上。
LEV|8|24|他領了 亞倫 的兒子來，把一些血抹在他們的右耳垂上，右手的大拇指上和右腳的大腳趾上。 摩西 把其餘的血灑在壇的周圍。
LEV|8|25|他把脂肪，肥尾巴、內臟所有的脂肪、肝上的網油、兩個腎、腎上的脂肪，和右腿取下，
LEV|8|26|再從耶和華面前那裝無酵餅的籃子中取一個無酵餅、一個油餅和一個薄餅，把這些放在脂肪和右腿上。
LEV|8|27|他把這一切放在 亞倫 和他兒子的手上，在耶和華面前搖一搖，作為搖祭。
LEV|8|28|摩西 從他們的手上把這些祭物拿來，放在壇的燔祭上燒，這就是聖職禮中獻給耶和華馨香的火祭。
LEV|8|29|摩西 拿羊的胸，在耶和華面前搖一搖，作為搖祭，這是聖職禮的羊歸給 摩西 的一份，是照耶和華所吩咐 摩西 的。
LEV|8|30|摩西 取些膏油和壇上的血，彈在 亞倫 和他的衣服上，以及他兒子和他們的衣服上，使 亞倫 和他的衣服，他兒子和他們的衣服都成為聖。
LEV|8|31|摩西 對 亞倫 和他兒子說：「你們要在會幕的門口把肉煮了，在那裏吃這肉和聖職禮中籃子裏的餅，按我所吩咐的說：『這是 亞倫 和他兒子當吃的。』
LEV|8|32|剩下的肉和餅，你們要用火焚燒。
LEV|8|33|這七天，你們不可走出會幕的門口，直等到你們聖職禮的日子滿了，因為授予你們聖職需要七天 。
LEV|8|34|今天所做的，都是耶和華吩咐要做的，好為你們贖罪。
LEV|8|35|這七天，你們要晝夜留在會幕門內，遵守耶和華所吩咐的，免得你們死亡，因為所吩咐我的就是這樣。」
LEV|8|36|於是， 亞倫 和他的兒子就做了耶和華藉著 摩西 所吩咐的一切事。
LEV|9|1|到了第八天， 摩西 召 亞倫 和他兒子，以及 以色列 的眾長老來，
LEV|9|2|對 亞倫 說：「你當取一頭公牛犢作贖罪祭，一隻公綿羊作燔祭，都要沒有殘疾的，獻在耶和華面前。
LEV|9|3|你要對 以色列 人說：『你們當取一隻公山羊作贖罪祭，再取一頭牛犢和一隻小綿羊，都要一歲沒有殘疾的，作燔祭；
LEV|9|4|又當取一頭公牛，一隻公綿羊作平安祭，宰殺獻在耶和華面前，再加上調油的素祭。因為今天耶和華要向你們顯現。』」
LEV|9|5|於是，他們把 摩西 所吩咐的帶到會幕前；全會眾都近前來，站在耶和華面前。
LEV|9|6|摩西 說：「這是耶和華吩咐你們當做的事，耶和華的榮光要向你們顯現。」
LEV|9|7|摩西 對 亞倫 說：「你靠近祭壇前，獻你的贖罪祭和燔祭，為自己與百姓贖罪，再獻上百姓的供物，為他們贖罪，都是照耶和華所吩咐的。」
LEV|9|8|於是， 亞倫 靠近壇前，宰了那頭為自己贖罪的牛犢。
LEV|9|9|亞倫 的兒子把血遞給他，他就把指頭蘸在血中，抹在壇的四個翹角上，再把其餘的血倒在壇的底座上。
LEV|9|10|他把贖罪祭的脂肪和腎，以及肝上的網油，燒在壇上，是照耶和華所吩咐 摩西 的。
LEV|9|11|他用火將肉和皮燒在營外。
LEV|9|12|亞倫 把燔祭牲宰了，他兒子把血遞給他，他就把血灑在壇的周圍。
LEV|9|13|他們又把燔祭一塊一塊地，連頭遞給他，他就燒在壇上。
LEV|9|14|他又洗了內臟和腿，放在壇的燔祭上燒。
LEV|9|15|然後，他奉上百姓的供物。他牽來給百姓作贖罪祭的公山羊，把牠宰了，獻為贖罪祭，和先前的一樣。
LEV|9|16|他也奉上燔祭，按照條例獻上。
LEV|9|17|除了早晨的燔祭以外，他又獻上素祭，用手取了滿滿的一把，燒在壇上。
LEV|9|18|亞倫 宰了那給百姓作平安祭的公牛和公綿羊，他兒子把血遞給他，他就把血灑在壇的周圍；
LEV|9|19|他們把公牛和公綿羊的脂肪、肥尾巴，包著內臟的脂肪，腎和肝上的網油，都遞給他。
LEV|9|20|他們把脂肪放在祭牲的胸上，他就把脂肪燒在壇上。
LEV|9|21|亞倫 把祭牲的胸和右腿在耶和華面前搖一搖，作為搖祭，是照 摩西 所吩咐的。
LEV|9|22|亞倫 向百姓舉手，為他們祝福。他獻了贖罪祭、燔祭、平安祭就下來了。
LEV|9|23|摩西 和 亞倫 進了會幕。他們出來，為百姓祝福；耶和華的榮光向全體百姓顯現。
LEV|9|24|有火從耶和華面前出來，焚燒了壇上的燔祭和脂肪；全體百姓一看見，就都歡呼，臉伏於地。
LEV|10|1|亞倫 的兒子 拿答 和 亞比戶 各拿著自己的香爐，把火放在爐裏，加上香，在耶和華面前獻上凡火，是耶和華沒有吩咐他們的。
LEV|10|2|有火從耶和華面前出來，把他們吞滅，他們就死在耶和華面前。
LEV|10|3|於是， 摩西 對 亞倫 說：「這就是耶和華所吩咐的，說：『我在那親近我的人中要顯為聖；在全體百姓面前，我要得著榮耀。』」 亞倫 就默默不言。
LEV|10|4|摩西 召 亞倫 的叔父 烏薛 的兒子 米沙利 和 以利撒反 前來，對他們說：「過來，把你們的親屬從聖所前抬到營外。」
LEV|10|5|於是，二人過來把屍體連袍子一起抬到營外，是照 摩西 所吩咐的。
LEV|10|6|摩西 對 亞倫 和他兒子 以利亞撒 和 以他瑪 說：「不可蓬頭散髮，也不可撕裂衣服，免得你們死亡，免得耶和華向全會眾發怒。但你們的弟兄 以色列 全家卻要為耶和華發出的火哀哭。
LEV|10|7|你們也不可出會幕的門口，免得你們死亡，因為耶和華的膏油在你們身上。」他們就遵照 摩西 的話去做了。
LEV|10|8|耶和華吩咐 亞倫 說：
LEV|10|9|「你和你兒子進會幕的時候，清酒烈酒都不可喝，免得你們死亡，這要作你們世世代代永遠的定例。
LEV|10|10|你們必須分辨聖的俗的，潔淨的和不潔淨的，
LEV|10|11|也要將耶和華藉 摩西 吩咐 以色列 人的一切律例教導他們。」
LEV|10|12|摩西 對 亞倫 和他剩下的兒子 以利亞撒 和 以他瑪 說：「獻給耶和華的火祭中所剩下的素祭，你們要拿來，在祭壇旁吃這無酵餅，因為它是至聖的。
LEV|10|13|你們要在聖處吃，因為在獻給耶和華的火祭中，這是你和你兒子當得的份；所吩咐我的就是這樣。
LEV|10|14|這搖祭的胸和這舉祭的腿，你要在潔淨的地方和你的兒女一同吃，因為這些是從 以色列 人的平安祭中歸給你，作為你和你兒子當得的份。
LEV|10|15|他們要把舉祭的腿、搖祭的胸和火祭的脂肪一同帶來，在耶和華面前搖一搖，作為搖祭。這些要歸給你和你兒子，作永遠當得的份，都是照耶和華所吩咐的。」
LEV|10|16|那時， 摩西 急切地尋找那隻贖罪祭的公山羊，看哪，牠已經燒掉了。他向 亞倫 剩下的兒子 以利亞撒 和 以他瑪 發怒，說：
LEV|10|17|「你們為何沒有在聖所吃這贖罪祭呢？它是至聖的，是耶和華給你們的，為了除掉會眾的罪孽，在耶和華面前為他們贖罪。
LEV|10|18|看哪，這祭牲的血沒有拿到聖所裏去！你們應當照我所吩咐的，在聖所裏吃這祭肉。」
LEV|10|19|亞倫 對 摩西 說：「看哪，他們今天在耶和華面前獻上贖罪祭和燔祭，但是我卻遭遇這樣的災難。我若今天吃這贖罪祭，耶和華豈能看為美呢？」
LEV|10|20|摩西 聽了，就看為美。
LEV|11|1|耶和華吩咐 摩西 和 亞倫 ，對他們說：
LEV|11|2|「你們要吩咐 以色列 人說，地上一切的走獸中可吃的動物是這些：
LEV|11|3|凡蹄分兩瓣，分趾蹄而又反芻食物的走獸，你們都可以吃。
LEV|11|4|但那反芻或分蹄之中不可吃的是：駱駝，反芻卻不分蹄，對你們是不潔淨的；
LEV|11|5|石獾，反芻卻不分蹄，對你們是不潔淨的；
LEV|11|6|兔子，反芻卻不分蹄，對你們是不潔淨的；
LEV|11|7|豬，蹄分兩瓣，分趾蹄卻不反芻，對你們是不潔淨的。
LEV|11|8|這些獸的肉，你們不可吃；牠們的屍體，你們也不可摸，對你們都是不潔淨的。
LEV|11|9|「水中可吃的是這些：凡在水裏，無論是海或河，有鰭有鱗的，都可以吃。
LEV|11|10|凡在海裏、河裏和水裏滋生的動物，就是在水裏所有的動物，無鰭無鱗的，對你們是可憎的。
LEV|11|11|牠們對你們都是可憎的。你們不可吃牠們的肉；牠們的屍體，也當以為可憎。
LEV|11|12|凡在水裏無鰭無鱗的，對你們是可憎的。
LEV|11|13|「飛鳥中你們當以為可憎，不可吃且可憎的是：鵰、狗頭鵰、紅頭鵰，
LEV|11|14|鷂鷹、小鷹的類群，
LEV|11|15|所有烏鴉的類群，
LEV|11|16|鴕鳥、夜鷹、魚鷹、鷹的類群，
LEV|11|17|鴞鳥、鸕鶿、貓頭鷹，
LEV|11|18|角鴟、鵜鶘、禿鵰，
LEV|11|19|鸛、鷺鷥的類群，戴鵀與蝙蝠。
LEV|11|20|「凡有翅膀卻用四足爬行的群聚動物，對你們是可憎的。
LEV|11|21|只是有翅膀卻用四足爬行的群聚動物中，足上有腿在地上跳的，你們還可以吃；
LEV|11|22|其中你們可以吃的有蝗蟲的類群，螞蚱的類群，蟋蟀的類群和蚱蜢的類群。
LEV|11|23|其餘有翅膀有四足的群聚動物，對你們都是可憎的。
LEV|11|24|「這些都能使你們不潔淨。凡摸牠們屍體的，必不潔淨到晚上。
LEV|11|25|任何人搬動了牠們的屍體，要把衣服洗淨，必不潔淨到晚上。
LEV|11|26|凡蹄分兩瓣卻不分趾或不反芻食物的走獸，對你們是不潔淨的；誰摸了牠們就不潔淨。
LEV|11|27|凡用腳掌行走，四足行走的動物，對你們是不潔淨的；凡摸牠們屍體的，必不潔淨到晚上。
LEV|11|28|誰搬動了牠們的屍體，要把衣服洗淨，必不潔淨到晚上。這些對你們是不潔淨的。
LEV|11|29|「在地上成群的群聚動物中，對你們不潔淨的是這些：鼬鼠、鼫鼠、蜥蜴的類群，
LEV|11|30|壁虎、龍子、守宮、蛇醫、蝘蜓。
LEV|11|31|這些群聚動物對你們都是不潔淨的。在牠們死後，凡摸了牠們屍體的，必不潔淨到晚上。
LEV|11|32|其中死了的，若掉在任何東西上，這東西就不潔淨，無論是木器、衣服、皮革、麻袋，或是任何工作需用的器皿，都要泡在水中，必不潔淨到晚上，然後才是潔淨的。
LEV|11|33|若有一點掉在瓦器裏，裏面的任何東西就不潔淨了； 你們要把這瓦器打破。
LEV|11|34|其中一切可吃的食物，沾到那水的就不潔淨；器皿裏可喝的東西，也必不潔淨。
LEV|11|35|牠們的屍體，只要有一點掉在任何物件上，那物件就不潔淨。無論是烤爐或爐灶，都要打碎；它們不潔淨，而且對你們也不潔淨。
LEV|11|36|但是水泉或池子，就是聚水的地方，仍是潔淨的；凡摸這些屍體的才不潔淨。
LEV|11|37|若牠們的屍體有一點掉在要播的種子上，種子仍是潔淨的；
LEV|11|38|若水已經澆在種子上，牠們的屍體有一點掉在上面，這種子對你們就是不潔淨的了。
LEV|11|39|「你們可吃的走獸中若有死了的，誰摸了牠的屍體，就必不潔淨到晚上。
LEV|11|40|人若吃了那已死的走獸，要把衣服洗淨，必不潔淨到晚上。人若搬動了那已死的牲畜，要把衣服洗淨，必不潔淨到晚上。
LEV|11|41|「凡在地上成群的群聚動物都是可憎的，都不可吃。
LEV|11|42|凡用肚子爬行或用四腳爬行，或是用多足的，地上一切群聚的動物，你們都不可吃，因為是可憎的。
LEV|11|43|你們不可因任何群聚的動物使自己成為可憎的，也不可因牠們成為不潔淨，染了污穢。
LEV|11|44|我是耶和華－你們的上帝。你們要使自己分別為聖，要成為聖，因為我是神聖的。你們不可因地上爬行的群聚動物使自己不潔淨。
LEV|11|45|我是把你們從 埃及 地領出來的耶和華，要作你們的上帝。你們要成為聖，因為我是神聖的。」
LEV|11|46|這是牲畜、飛鳥、水中一切游動的生物和地上一切爬行的動物的條例，
LEV|11|47|為要使你們能分辨潔淨的和不潔淨的，可吃的和不可吃的動物。
LEV|12|1|耶和華吩咐 摩西 說：
LEV|12|2|「你要吩咐 以色列 人說：婦人若懷孕生男孩，就不潔淨七天，像在月經污穢的期間不潔淨一樣。
LEV|12|3|第八天，要給嬰孩行割禮。
LEV|12|4|婦人產後流血的潔淨，要家居三十三天。她潔淨的日子未滿，不可摸聖物，也不可進入聖所。
LEV|12|5|她若生女孩，就不潔淨兩個七天，像經期中一樣。她產後流血的潔淨，要家居六十六天。
LEV|12|6|「潔淨的日子滿了，無論生兒子或女兒，她要把一隻一歲的羔羊作燔祭，一隻雛鴿或一隻斑鳩作贖罪祭，帶到會幕的門口交給祭司。
LEV|12|7|祭司要把這祭物獻在耶和華面前，為她贖罪。這樣，她就從流血中得潔淨了。這是為生男或生女之婦人的條例。
LEV|12|8|婦人的能力若不足，無法獻一隻羔羊，她就要取兩隻斑鳩或兩隻雛鴿，一隻為燔祭，一隻為贖罪祭。祭司要為她贖罪，她就潔淨了。」
LEV|13|1|耶和華吩咐 摩西 和 亞倫 說：
LEV|13|2|「人身上的皮膚若腫脹，或發疹，或有斑點，可能成為痲瘋 的災病，就要把他帶到 亞倫 祭司或 亞倫 的一個作祭司的子孫那裏。
LEV|13|3|祭司要檢查他身上皮膚的患處，若患處的毛已經變白，災病的現象深入身上皮膚內，這就是痲瘋的災病。祭司檢查後，要宣佈他為不潔淨。
LEV|13|4|若這人身上的皮膚有白斑，看起來並沒有深入皮膚內，其上的毛也沒有變白，祭司就要將這病人隔離七天。
LEV|13|5|第七天，祭司要檢查他，看哪，若災病在祭司眼前止住了，沒有在皮膚上擴散，要將他再隔離七天。
LEV|13|6|到了第七天，祭司要再檢查他。看哪，若災病減輕，沒有在皮膚上擴散，祭司就要宣佈他為潔淨，因為他患的不過是疹子。那人要洗自己的衣服，就潔淨了。
LEV|13|7|他給祭司檢查宣佈為潔淨後，疹子若在皮膚上大大擴散，他就要再給祭司檢查。
LEV|13|8|祭司要檢查，看哪，疹子若在皮膚上擴散了，祭司就要宣佈他為不潔淨，是痲瘋病。
LEV|13|9|「人若得了痲瘋的災病，就要把他帶到祭司那裏。
LEV|13|10|祭司要檢查，看哪，若皮膚有白色腫塊，使毛變白，腫塊裏有嫩的新長的肉，
LEV|13|11|這就是他身上皮膚慢性的痲瘋病。祭司要宣佈他為不潔淨，不必將他隔離，因為他已是不潔淨了。
LEV|13|12|若痲瘋在皮膚四處擴散，長滿在患災病之人的皮膚上，據祭司察看，從頭到腳無處不有，
LEV|13|13|祭司就要檢查，看哪，若這病人全身已長滿了痲瘋，就要宣佈他為潔淨；他全身都變白了，他是潔淨的。
LEV|13|14|但他身上一旦出現新長的肉，就不潔淨了。
LEV|13|15|祭司一見新長的肉，就要宣佈他為不潔淨。新長的肉是不潔淨的，這就是痲瘋病。
LEV|13|16|新長的肉若變白了，他就要到祭司那裏。
LEV|13|17|祭司要檢查，看哪，患處若變白了，祭司就要宣佈那患災病的人為潔淨，他就潔淨了。
LEV|13|18|「人身上的皮膚 若長了瘡，卻已經好了，
LEV|13|19|在長瘡之處又發腫變白，或是出現白中帶紅的斑點，就要給祭司檢查。
LEV|13|20|祭司要檢查，看哪，若災病的現象已深入皮膚內，其上的毛也變白了，祭司就要宣佈他為不潔淨，有痲瘋的災病生在瘡中。
LEV|13|21|祭司若檢查，看哪，其上沒有白毛，也沒有深入皮膚內，而且災病減輕，祭司就要將他隔離七天。
LEV|13|22|若在皮膚上大大擴散，祭司就要宣佈他為不潔淨，這是災病。
LEV|13|23|斑點若留在原處，沒有擴散，這就是瘡的疤痕，祭司就要宣佈他為潔淨。
LEV|13|24|「人身上的皮膚若被火燒傷，傷口新長的肉有了斑點，無論是白中帶紅，或是全白，
LEV|13|25|祭司就要檢查，看哪，斑點上的毛若變白了，現象又深入皮膚內，這就是痲瘋長在燒傷處；祭司就要宣佈他為不潔淨，是痲瘋的災病。
LEV|13|26|若祭司檢查，看哪，斑點上沒有白毛，也沒有深入皮膚內，而且災病減輕，祭司就要將他隔離七天。
LEV|13|27|第七天，祭司要檢查他。斑點若在皮膚上大大擴散，祭司就要宣佈他為不潔淨，是患了痲瘋的災病。
LEV|13|28|斑點若留在原處，沒有在皮膚上擴散，並減輕了，它只是燒傷的腫塊，祭司要宣佈他為潔淨，這不過是燒傷後的疤痕。
LEV|13|29|「無論男女，若在頭上或下巴有災病，
LEV|13|30|祭司就要檢查這災病，看哪，若災病的現象深入皮膚內，其上有黃色的細毛，祭司就要宣佈他為不潔淨，這是疥瘡，是頭上或下巴的痲瘋病。
LEV|13|31|祭司要檢查這疥瘡的災病，看哪，現象若未深入皮膚內，其上也沒有黑毛，祭司就要將長疥瘡的人隔離七天。
LEV|13|32|第七天，祭司要檢查這災病，看哪，若疥瘡沒有擴散，其上沒有黃色的毛，疥瘡的現象也沒有深入皮膚內，
LEV|13|33|那人就要剃去鬚髮，但不可剃長疥瘡之處。祭司要將那長疥瘡的人，再隔離七天。
LEV|13|34|第七天，祭司要檢查疥瘡，看哪，疥瘡若沒有在皮膚上擴散，現象也未深入在皮膚內，祭司就要宣佈他為潔淨；那人要洗自己的衣服，就潔淨了。
LEV|13|35|但他被宣佈為潔淨後，疥瘡若在皮膚上大大擴散，
LEV|13|36|祭司就要檢查他。看哪，疥瘡若在皮膚上擴散，祭司就不必找黃色的毛，這人是不潔淨了。
LEV|13|37|若疥瘡在祭司眼前止住了，其上長了黑毛，疥瘡就已痊癒了，那人是潔淨的，祭司要宣佈他為潔淨。
LEV|13|38|「無論男女，身上的皮膚若有斑點，是白色的斑點，
LEV|13|39|祭司就要檢查，看哪，若皮膚的斑點是暗白色的，這是皮膚長了斑；那人是潔淨的。
LEV|13|40|「人的頭髮若掉了，變成禿頭，他是潔淨的。
LEV|13|41|他頭頂的前面若掉了頭髮，以致頂門光禿，他是潔淨的。
LEV|13|42|頭禿處或頂門禿處，若有白中帶紅的災病，這就是痲瘋長在他的頭禿處或頂門禿處。
LEV|13|43|祭司要檢查他，看哪，若頭禿處或頂門禿處的災病腫塊白中帶紅，像身上皮膚痲瘋病的現象一樣，
LEV|13|44|那人就是患了痲瘋病，是不潔淨的。祭司要宣佈他為不潔淨；他的災病是生在頭上。
LEV|13|45|「患有痲瘋災病的人，他的衣服要撕裂，也要蓬頭散髮，遮住上唇，喊著說：『不潔淨！不潔淨！』
LEV|13|46|災病還在他身上的時候，他就是不潔淨的；既然不潔淨，他就要獨居，住在營外。」
LEV|13|47|「衣服若發霉 了，無論是羊毛衣服、麻布衣服，
LEV|13|48|無論是經線、緯線，是麻布的、羊毛的，是皮革，或是任何皮製的物件；
LEV|13|49|若是衣服、皮革、經線、緯線，或是任何皮製的物件呈現綠色或紅色，這就是發霉，必須給祭司檢查。
LEV|13|50|祭司要檢查這霉，把發霉的物件隔離七天。
LEV|13|51|第七天，他要檢查這霉。若霉在衣服上，無論是經線、緯線，或任何用途的皮製物件上擴散，這是侵蝕性的霉，是不潔淨的。
LEV|13|52|發霉的衣服，無論在經線、緯線，羊毛的、麻布的，或是任何皮製物件，都要把它燒掉；因為這是侵蝕性的霉，必須用火焚燒。
LEV|13|53|祭司檢查，看哪，霉若在衣服上，無論是經線、緯線，或在任何的皮製物件上沒有擴散，
LEV|13|54|祭司就要吩咐人把發霉的物件洗了，再隔離七天。
LEV|13|55|洗過之後，祭司要檢查，看哪，若那霉在他眼前沒有變色，霉雖沒有擴散，也是不潔淨的。這是侵蝕性的災病，無論是在正面或反面，都要用火焚燒那物件。
LEV|13|56|祭司若檢查，看哪，那霉在洗過之後已經褪色，他就要從衣服，皮革，或經線、緯線，把發霉的部分撕去。
LEV|13|57|若霉再出現在衣服上，無論是經線、緯線、或在任何皮製物件上，這就是舊霉復發，必須用火將那發霉的物件焚燒。
LEV|13|58|洗過的衣服，或是經線，緯線，或是任何皮製的物件，若霉已經消失了，仍要再洗，這衣服就潔淨了。」
LEV|13|59|這就是衣服發霉的條例。無論是羊毛衣服，麻布衣服，或是經線、緯線，或任何皮製的物件，都按照這條例宣佈為潔淨或不潔淨。
LEV|14|1|耶和華吩咐 摩西 說：
LEV|14|2|「這是患痲瘋病的人得潔淨時的條例：要帶他到祭司那裏，
LEV|14|3|祭司要出到營外，檢查那患痲瘋病的人，看哪，他的痲瘋災病已經痊癒了，
LEV|14|4|祭司就要吩咐人為那求潔淨的人帶兩隻潔淨的活鳥和香柏木、朱紅色紗，以及牛膝草來。
LEV|14|5|祭司要吩咐用瓦器盛清水，把第一隻鳥宰在上面。
LEV|14|6|至於那隻活鳥，祭司要把牠和香柏木、朱紅色紗，以及牛膝草，一同蘸在宰於清水上的鳥血中。
LEV|14|7|他要向那從痲瘋病中得潔淨的人身上彈血七次，宣佈他為潔淨，然後把那活鳥在野地裏放走。
LEV|14|8|求潔淨的人要洗衣服，剃去所有的毛髮，用水洗澡，他就潔淨了。然後，他可以進營，不過仍要在自己的帳棚外居住七天。
LEV|14|9|到了第七天，他要剃所有的毛髮，頭髮、鬍鬚、眼睛的眉毛，他全身的毛都剃了；然後，他要洗衣服，用水洗身，才潔淨了。
LEV|14|10|「第八天，他要取兩隻沒有殘疾的小公羊和一隻沒有殘疾、一歲的小母羊，以及作為素祭的十分之三伊法調了油的細麵和一羅革的油。
LEV|14|11|宣佈潔淨的祭司要將那求潔淨的人，連同這些東西，安置在耶和華面前，會幕的門口。
LEV|14|12|祭司要取一隻小公羊獻為贖愆祭，又取一羅革的油，把它們在耶和華面前搖一搖，作為搖祭；
LEV|14|13|再把小公羊宰於聖處，就是宰贖罪祭牲和燔祭牲的地方。贖愆祭要歸給祭司，與贖罪祭一樣，是至聖的。
LEV|14|14|祭司要取一些贖愆祭牲的血，抹在求潔淨的人的右耳垂上、右手的大拇指上和右腳的大腳趾上。
LEV|14|15|祭司要從那一羅革的油中，取一些倒在自己的左手掌裏，
LEV|14|16|祭司要用右手指蘸在他左手掌的油裏，在耶和華面前用手指彈七次。
LEV|14|17|祭司要把手掌裏剩下的油抹在那求潔淨的人的右耳垂上、右手的大拇指上和右腳的大腳趾上，在贖愆祭牲之血抹過的上面。
LEV|14|18|祭司手掌裏剩下的油要抹在那求潔淨的人的頭上，祭司就在耶和華面前為他贖罪。
LEV|14|19|祭司要獻贖罪祭，為那從不潔淨中得潔淨的人贖罪，然後要宰燔祭牲，
LEV|14|20|祭司要把燔祭和素祭獻在壇上，祭司要為他贖罪，他就潔淨了。
LEV|14|21|「他若貧窮，手頭財力不及，就要取一隻小公羊作贖愆祭，作搖祭為他贖罪。他也要把作為素祭的十分之一伊法調了油的細麵，和一羅革的油，一同取來。
LEV|14|22|他又要照手頭財力所及，取兩隻斑鳩或兩隻雛鴿，一隻作贖罪祭，一隻作燔祭。
LEV|14|23|第八天，為了使自己潔淨，他要把這些祭物帶到耶和華面前，在會幕的門口交給祭司。
LEV|14|24|祭司要把贖愆祭的羔羊和那一羅革的油一同在耶和華面前搖一搖，作為搖祭。
LEV|14|25|祭司要宰贖愆祭的羔羊，取一些贖愆祭牲的血，抹在那求潔淨的人的右耳垂上、右手的大拇指上和右腳的大腳趾上。
LEV|14|26|祭司要把一些油倒在自己的左手掌裏，
LEV|14|27|祭司要用右手指，把他左手掌裏的油在耶和華面前彈七次。
LEV|14|28|祭司要把手掌裏的油抹一些在那求潔淨的人的右耳垂上、右手的大拇指上和右腳的大腳趾上，在贖愆祭牲之血抹過之處的上面。
LEV|14|29|祭司手掌裏剩下的油要抹在那求潔淨的人的頭上，在耶和華面前為他贖罪。
LEV|14|30|那人又要照他手頭財力所及，獻上斑鳩中的一隻或雛鴿中的一隻，
LEV|14|31|照他手頭財力所及，一隻為贖罪祭，一隻為燔祭，與素祭一同獻上。祭司就在耶和華面前為他贖罪。
LEV|14|32|這是為患痲瘋災病，手頭財力不及而求潔淨的人所定的條例。」
LEV|14|33|耶和華吩咐 摩西 和 亞倫 說：
LEV|14|34|「你們到了我所賜給你們為業的 迦南 地，我若使你們所得為業之地的房屋發霉 ，
LEV|14|35|屋主就要去告訴祭司說：『據我看，房屋似乎發霉了。』
LEV|14|36|祭司進去檢查這霉之前，要吩咐把屋內的東西全部搬走，免得屋子裏所有的東西成為不潔淨。然後，祭司要進去檢查房屋。
LEV|14|37|他要檢查這霉，看哪，若屋子牆上的霉有發綠或發紅凹入的斑紋，其現象深入牆內，
LEV|14|38|祭司就要出到屋子的門外，把屋子封鎖七天。
LEV|14|39|第七天，祭司要再去檢查，看哪，霉若在屋子的牆上擴散，
LEV|14|40|祭司要吩咐把發霉的石頭挖出來，扔在城外不潔淨之處。
LEV|14|41|他也要叫人刮屋內的四圍，把刮出來的灰泥倒在城外不潔淨之處。
LEV|14|42|他們要用別的石頭取代挖出來的石頭，用別的灰泥塗抹屋子。
LEV|14|43|「他挖出石頭，刮了屋子，塗抹以後，霉若又在屋子裏出現，
LEV|14|44|祭司就要進去檢查，看哪，霉若在屋子裏擴散，那就是有侵蝕性的霉在屋子裏，是不潔淨的。
LEV|14|45|他要拆毀屋子，把石頭、木料和所有的灰泥都搬到城外不潔淨之處。
LEV|14|46|屋子封鎖的任何時候，進去的人必不潔淨到晚上。
LEV|14|47|在屋子裏躺臥的人必須把衣服洗淨，在屋子裏吃飯的人也必須把衣服洗淨。
LEV|14|48|「屋子塗抹了之後，祭司若進去檢查，看哪，霉沒有在屋內擴散，就要宣佈這房屋為潔淨，因為霉已經消除了。
LEV|14|49|他要為潔淨房屋取兩隻鳥和香柏木、朱紅色紗，以及牛膝草，
LEV|14|50|用瓦器盛清水，把一隻鳥宰在上面。
LEV|14|51|他要把香柏木、牛膝草、朱紅色紗和那一隻活鳥，都蘸在被宰的鳥血和清水中，用來彈屋子七次。
LEV|14|52|他要用鳥血、清水、活鳥、香柏木、牛膝草和朱紅色紗潔淨那房屋。
LEV|14|53|他要把活鳥在城外野地裏放走。他要為房屋贖罪，房屋就潔淨了。」
LEV|14|54|這條例是為痲瘋災病和疥瘡，
LEV|14|55|衣服和房屋發霉，
LEV|14|56|以及皮膚腫脹、發疹、有斑點等，
LEV|14|57|用以分辨何時潔淨，何時不潔淨。這是痲瘋病的條例。
LEV|15|1|耶和華吩咐 摩西 和 亞倫 說：
LEV|15|2|「你們要吩咐 以色列 人，對他們說：人若身體 患了漏症，他因這症就不潔淨了。
LEV|15|3|這就是他因漏症而有的不潔淨：無論是身體流出液體，或身體已經止住不再有液體，他都是不潔淨的。
LEV|15|4|那患漏症的人所躺的床都不潔淨，所坐的任何東西也不潔淨。
LEV|15|5|凡摸他床的人，要洗衣服，用水洗澡，必不潔淨到晚上。
LEV|15|6|人坐了漏症患者坐過的東西，他要洗衣服，用水洗澡，必不潔淨到晚上。
LEV|15|7|人摸了漏症患者，他要洗衣服，用水洗澡，必不潔淨到晚上。
LEV|15|8|若漏症患者吐唾沫在潔淨的人身上，這人要洗衣服，用水洗澡，必不潔淨到晚上。
LEV|15|9|漏症患者所騎的任何鞍子也不潔淨。
LEV|15|10|凡摸了他坐過的任何東西，必不潔淨到晚上；拿了這些東西的，要洗衣服，用水洗澡，必不潔淨到晚上。
LEV|15|11|漏症患者若沒有用水沖洗他的手，無論摸了誰，誰就要洗衣服，用水洗澡，必不潔淨到晚上。
LEV|15|12|漏症患者所摸的瓦器必要打破；他所摸的一切木器必要用水沖洗。
LEV|15|13|「漏症患者的漏症痊癒了，就要為潔淨自己計算七天，也要洗衣服，用清水洗身，就潔淨了。
LEV|15|14|第八天，他要帶兩隻斑鳩或兩隻雛鴿，來到耶和華面前，在會幕門口把鳥交給祭司。
LEV|15|15|祭司要獻上一隻為贖罪祭，一隻為燔祭。祭司要因這人所患的漏症，在耶和華面前為他贖罪。
LEV|15|16|「人若遺精，他要用水洗全身，必不潔淨到晚上。
LEV|15|17|無論是衣服或皮革，若沾染了精液，要用水洗淨，必不潔淨到晚上。
LEV|15|18|女人，若有男人與她同寢，沾染了精液，二人要用水洗澡，必不潔淨到晚上。」
LEV|15|19|「女人月經期間，有血從體內流出，她必不潔淨七天；凡摸她的，必不潔淨到晚上。
LEV|15|20|在不潔淨期間，女人所躺的東西都不潔淨，所坐的任何東西也不潔淨。
LEV|15|21|凡摸她床的，要洗衣服，用水洗澡，必不潔淨到晚上；
LEV|15|22|凡摸她坐過的東西的，要洗衣服，用水洗澡，必不潔淨到晚上；
LEV|15|23|不論是床，或她坐過的東西，人摸了，必不潔淨到晚上。
LEV|15|24|男人若和這女人同寢，沾了她的不潔淨，就不潔淨七天，所躺的床也都不潔淨。
LEV|15|25|「女人若在經期之外仍然流血多日，或是經期過長，她在流血的一切日子都不潔淨，和她在經期的日子不潔淨一樣。
LEV|15|26|在流血的日子，她所躺的床、所坐的任何東西都不潔淨，和在月經期間不潔淨一樣。
LEV|15|27|凡摸這些東西的，就不潔淨；他要洗衣服，用水洗澡，必不潔淨到晚上。
LEV|15|28|這女人的血漏若痊癒了，就要計算七天，然後才潔淨。
LEV|15|29|第八天，她要取兩隻斑鳩或兩隻雛鴿，帶到會幕門口祭司那裏。
LEV|15|30|祭司要獻一隻為贖罪祭，一隻為燔祭。祭司要因這女人血漏的不潔淨，在耶和華面前為她贖罪。
LEV|15|31|「你們要使 以色列 人與他們的不潔淨隔離，免得他們玷污我在他們中間的帳幕，因自己的不潔淨死亡。」
LEV|15|32|這條例是為漏症患者或遺精而不潔淨者，
LEV|15|33|女人經期的不潔，男女患漏症，以及男人與不潔淨女人同寢而立的。
LEV|16|1|亞倫 的兩個兒子靠近耶和華面前，死了。他們死後，耶和華吩咐 摩西 ；
LEV|16|2|耶和華對 摩西 說：「你要吩咐你哥哥 亞倫 ，不可隨時進入聖所的幔子內、到櫃蓋 前，免得他死亡，因為我在櫃蓋上的雲中顯現。
LEV|16|3|亞倫 進聖所要帶這些：一頭公牛犢為贖罪祭，一隻公綿羊為燔祭。
LEV|16|4|他要穿上細麻布聖內袍，把細麻布褲子穿在身上，腰束細麻布帶子，頭戴細麻布禮冠；這些都是聖服。他要用水洗身，然後穿上聖服。
LEV|16|5|他要從 以色列 會眾中取兩隻公山羊為贖罪祭，一隻公綿羊為燔祭。
LEV|16|6|「亞倫要把他自己贖罪祭的公牛獻上，為自己和家人贖罪；
LEV|16|7|也要把兩隻公山羊牽到耶和華面前，安置在會幕的門口。
LEV|16|8|亞倫 要為那兩隻山羊抽籤，一籤歸給耶和華，一籤歸給 阿撒瀉勒 。
LEV|16|9|亞倫 要把那抽中歸給耶和華的山羊牽來獻為贖罪祭，
LEV|16|10|至於抽中歸給 阿撒瀉勒 的山羊，卻要活著安放在耶和華面前，用以贖罪，然後送到曠野去，歸給 阿撒瀉勒 。
LEV|16|11|「 亞倫 要把他自己贖罪祭的公牛獻上，為自己和家人贖罪，他要宰作自己贖罪祭的公牛。
LEV|16|12|他要從耶和華面前的壇上取盛滿火炭的香爐，再拿一捧搗細的香料，把這些都帶入幔子內。
LEV|16|13|在耶和華面前，他要把香放在火上，使香的煙雲遮著法櫃上的蓋子，免得他死亡。
LEV|16|14|他要取一些公牛的血，用手指彈在櫃蓋的前面，就是東面，又在櫃蓋的前面用手指彈血七次。
LEV|16|15|「他要宰那隻為百姓作贖罪祭的公山羊，把羊的血帶入幔子內，把血彈在櫃蓋的上面和前面，好像彈公牛的血一樣。
LEV|16|16|因 以色列 人的不潔淨和過犯，就是他們一切的罪，他要為聖所贖罪；因會幕在他們不潔淨之中，他也要為會幕照樣做。
LEV|16|17|他進聖所贖罪的時候，會幕裏都不准有人，直等到他為自己和家人，以及 以色列 全會眾贖了罪出來。
LEV|16|18|他出來後，要到耶和華面前的祭壇那裏，為壇贖罪。他要取一些公牛的血和公山羊的血，抹在壇周圍的四個翹角上。
LEV|16|19|他也要用手指把血彈在壇上七次，使壇從 以色列 人的不潔淨中得以潔淨，成為聖。」
LEV|16|20|「 亞倫 為聖所和會幕，以及祭壇贖罪後，就要把那隻活的公山羊牽來。
LEV|16|21|他的雙手要按在活的山羊的頭上，承認 以色列 人所有的罪孽過犯，就是他們一切的罪，把這些罪都歸在羊的頭上，再指派一個人把牠送到曠野去。
LEV|16|22|這羊要擔當他們一切的罪孽，帶到無人之地；那人要把羊送到曠野去。
LEV|16|23|「 亞倫 要進入會幕，把他進聖所時所穿的細麻布衣服脫下，放在那裏，
LEV|16|24|又要在聖處用水洗身，穿上衣服出來，把自己的燔祭和百姓的燔祭獻上，為自己和百姓贖罪。
LEV|16|25|贖罪祭牲的脂肪要燒在壇上。
LEV|16|26|那放走山羊歸給 阿撒瀉勒 的人要洗衣服，用水洗身，然後才可以回到營裏。
LEV|16|27|作贖罪祭的公牛和作贖罪祭的公山羊的血被帶入聖所贖罪之後，就要把這牛羊搬到營外，皮、肉、糞都用火焚燒。
LEV|16|28|焚燒的人要洗衣服，用水洗身，然後才可以回到營裏。」
LEV|16|29|「這是你們永遠的定例：每年七月初十，你們要刻苦己心；無論是本地人，是寄居在你們中間的外人，任何工都不可做。
LEV|16|30|因為這日要為你們贖罪，潔淨你們，使你們脫離一切的罪，在耶和華面前得以潔淨。
LEV|16|31|這日你們要守完全安息的安息日，刻苦己心；這是永遠的定例。
LEV|16|32|那受膏接續他父親擔任聖職的祭司要贖罪，穿上細麻布衣服，就是聖衣，
LEV|16|33|為至聖所和會幕贖罪，為祭壇贖罪，並要為祭司和會眾的全體百姓贖罪。
LEV|16|34|這要作你們永遠的定例：因 以色列 人一切的罪，要一年一次為他們贖罪。」於是， 亞倫 照耶和華所吩咐 摩西 的做了 。
LEV|17|1|耶和華吩咐 摩西 說：
LEV|17|2|「你要吩咐 亞倫 和他兒子，以及 以色列 眾人，對他們說，耶和華所吩咐的話是這樣：
LEV|17|3|凡 以色列 家中的人宰公牛，或小綿羊，或山羊，無論是在營內或營外，
LEV|17|4|若不把牲畜牽到會幕門口耶和華的帳幕前，獻給耶和華為供物，所流的血必歸到那人身上。他既使血流出，就要從百姓中剪除。
LEV|17|5|這是為要使 以色列 人把他們在野地裏所宰的祭牲帶來，帶到耶和華前，會幕門口祭司那裏，宰殺這些祭牲，把牠們獻給耶和華為平安祭。
LEV|17|6|祭司要在會幕門口，把血灑在耶和華的祭壇上，把脂肪焚燒，獻給耶和華為馨香的祭。
LEV|17|7|他們不可再宰殺祭牲獻給他們行淫所隨從的山羊鬼魔。這要作他們世世代代永遠的定例。
LEV|17|8|「你要對他們說：凡 以色列 家中的任何人，或寄居在他們中間的外人獻燔祭或祭物，
LEV|17|9|若不帶到會幕門口獻給耶和華，那人必從百姓中剪除。
LEV|17|10|「凡 以色列 家中的任何人，或寄居在他們中間的外人，吃任何的血，我必向那吃血的人變臉，把他從百姓中剪除。
LEV|17|11|因為動物的生命是在血中。我把這血賜給你們，可以在祭壇上為你們的生命贖罪；因為血就是生命，能夠贖罪。
LEV|17|12|因此，我對 以色列 人說：你們都不可吃血；寄居在你們中間的外人也不可吃血。
LEV|17|13|凡 以色列 人，或寄居在他們中間的外人，獵取了可吃的飛禽走獸，必須把牠的血放出來，用土掩蓋。
LEV|17|14|「因一切動物的生命，牠的血就是牠的生命。所以我對 以色列 人說：無論甚麼動物的血，你們都不可吃，因為一切動物的生命就是牠的血。凡吃血的必被剪除。
LEV|17|15|無論是本地人，是寄居的，若吃了自然死去或被野獸撕裂的動物，要洗衣服，用水洗澡，必不潔淨到晚上，晚上就潔淨了。
LEV|17|16|但他若不洗衣服，也不洗身，就要擔當自己的罪孽。」
LEV|18|1|耶和華吩咐 摩西 說：
LEV|18|2|「你要吩咐 以色列 人，對他們說：我是耶和華－你們的上帝。
LEV|18|3|你們不可做你們從前住 埃及 地的人所做的，也不可做我要領你們去的 迦南 地的人所做的。你們不可照他們的習俗行。
LEV|18|4|你們要遵行我的典章，謹守我的律例，按此而行。我是耶和華－你們的上帝。
LEV|18|5|你們要謹守我的律例典章；遵行的人就必因此得生。我是耶和華。
LEV|18|6|「任何人都不可親近骨肉之親，露其下體。我是耶和華。
LEV|18|7|你父親的下體，就是你母親的下體，你不可露；她是你的母親，不可露她的下體。
LEV|18|8|不可露你繼母的下體，就是你父親的下體。
LEV|18|9|你姊妹的下體，或是同父異母的，或是同母異父的，無論生在家或生在外的，都不可露她們的下體。
LEV|18|10|不可露你孫女或外孫女的下體，因為她們的下體就是你自己的下體。
LEV|18|11|你繼母為你父親所生的女兒是你的姊妹，不可露她的下體。
LEV|18|12|不可露你姑母的下體；她是你父親的骨肉之親。
LEV|18|13|不可露你姨母的下體；她是你母親的骨肉之親。
LEV|18|14|不可露你叔伯的下體，不可親近他的妻子；她是你的叔母、伯母。
LEV|18|15|不可露你媳婦的下體，她是你兒子的妻，不可露她的下體。
LEV|18|16|不可露你兄弟妻子的下體，這是你兄弟的下體。
LEV|18|17|不可露婦人的下體，又露她女兒的下體，也不可娶她的孫女或外孫女，露她們的下體；她們是骨肉之親 。這是邪惡的事。
LEV|18|18|你妻子還活著的時候，不可另娶她的姊妹與她作對，露她姊妹的下體。
LEV|18|19|「不可親近經期中不潔淨的女人，露她的下體。
LEV|18|20|不可跟鄰舍的妻交合，因她玷污自己。
LEV|18|21|不可使你兒女經火獻給 摩洛 ，也不可褻瀆你上帝的名。我是耶和華。
LEV|18|22|不可跟男人同寢，像跟女人同寢；這是可憎惡的事。
LEV|18|23|不可跟獸交合，因牠玷污自己。女人也不可站在獸前，與牠交合；這是逆性的事。
LEV|18|24|「在這一切的事上，你們都不可玷污自己，因為我在你們面前所逐出的列國，在這一切的事上玷污了自己。
LEV|18|25|連地也玷污了，我懲罰那地的罪孽，地就吐出它的居民來。
LEV|18|26|但你們要遵守我的律例典章。這一切可憎惡的事，無論是本地人或寄居在你們中間的外人，都不可以做。
LEV|18|27|在你們之前居住那地的人做了這一切可憎惡的事，地就玷污了。
LEV|18|28|不要讓地因你們玷污了它而把你們吐出來，像吐出在你們之前的國一樣。
LEV|18|29|無論是誰，若做了這其中一件可憎惡的事，必從百姓中剪除。
LEV|18|30|你們要遵守我的吩咐，免得你們隨從那些可憎的習俗，就是在你們之前的人所做的，玷污了自己。我是耶和華－你們的上帝。」
LEV|19|1|耶和華吩咐 摩西 說：
LEV|19|2|「你要吩咐 以色列 全會眾，對他們說：你們要成為聖，因為我耶和華－你們的上帝是神聖的。
LEV|19|3|你們各人都當孝敬父母，也要守我的安息日。我是耶和華－你們的上帝。
LEV|19|4|你們不可轉向虛無的神明，也不可為自己鑄造神像。我是耶和華－你們的上帝。
LEV|19|5|「你們宰殺祭牲獻平安祭給耶和華的時候，要獻得使你們可蒙悅納。
LEV|19|6|這祭物要在獻的當天或第二天吃；若有剩到第三天的，就要用火焚燒。
LEV|19|7|第三天若再吃，這祭物是不潔淨的，必不蒙悅納。
LEV|19|8|吃的人必擔當自己的罪孽，因為他褻瀆了耶和華的聖物，這人必從百姓中剪除。
LEV|19|9|「你們在自己的地收割莊稼時，不可割盡田的角落，也不可拾取莊稼所掉落的。
LEV|19|10|不可摘盡葡萄園的葡萄，也不可拾取葡萄園中掉落的葡萄，要把它們留給窮人和寄居的。我是耶和華－你們的上帝。
LEV|19|11|「你們不可偷盜，不可欺騙，也不可彼此說謊。
LEV|19|12|不可指著我的名起假誓，褻瀆你上帝的名。我是耶和華。
LEV|19|13|「不可欺壓你的鄰舍，也不可偷盜。雇工的工錢不可在你那裏過夜，留到早晨。
LEV|19|14|不可咒罵聾子，也不可將絆腳石放在盲人面前。你要敬畏你的上帝。我是耶和華。
LEV|19|15|「你們審判的時候，不可不公正；不可偏護貧窮人，也不可看重有權勢人的臉，總要公平審判你的鄰舍。
LEV|19|16|不可在百姓中到處搬弄是非，不可陷害鄰舍的性命 。我是耶和華。
LEV|19|17|「不可心裏恨你的弟兄；要指摘你的鄰舍，免得因他承擔罪過。
LEV|19|18|不可報仇，也不可埋怨你本國的子民。你要愛鄰如己。我是耶和華。
LEV|19|19|「你們要遵守我的律例。不可使你的牲畜與異類交配；不可在你的田地播下兩樣的種子；也不可穿兩種原料做成的衣服。
LEV|19|20|「若有人與女子同寢交合，而她是婢女，許配了丈夫，尚未被贖或得自由，就要受到懲罰，卻不可把他們處死，因為婢女還沒有得自由。
LEV|19|21|男的要把贖愆祭，就是一隻公綿羊牽到耶和華面前，會幕的門口。
LEV|19|22|祭司要用贖愆祭的羊在耶和華面前為他所犯的罪贖罪，他所犯的罪就必蒙赦免。
LEV|19|23|「你們到了 迦南 地，栽種各樣的果樹，就要把所結的果子當作不潔淨的 ；三年之內，你們要把它視為不潔淨，是不可吃的。
LEV|19|24|但第四年所結的果子全是聖的，用以讚美耶和華 。
LEV|19|25|第五年，你們就可以吃樹上的果子，使樹給你們結出更多的果子。我是耶和華－你們的上帝。
LEV|19|26|「你們不可吃帶血的食物。不可占卜，也不可觀星象。
LEV|19|27|頭的周圍 不可剃，鬍鬚的周圍不可損壞。
LEV|19|28|不可為死人割劃自己的身體，也不可在身上刺花紋。我是耶和華。
LEV|19|29|「不可侮辱你的女兒，使她淪為娼妓，免得這地行淫亂，地就充滿了邪惡。
LEV|19|30|你們要謹守我的安息日，敬畏我的聖所。我是耶和華。
LEV|19|31|「不可轉向招魂的，也不可求問行巫術的，免得被他們玷污。我是耶和華－你們的上帝。
LEV|19|32|「在白髮的人面前，你要站起來，要尊敬老人；要敬畏你的上帝，我是耶和華。
LEV|19|33|「若有外人寄居在你們的地上和你同住，不可欺負他。
LEV|19|34|寄居在你們那裏的外人，你們要看他如本地人，並要愛他如己，因為你們在 埃及 地也作過寄居的。我是耶和華－你們的上帝。
LEV|19|35|「你們審判的時候，不可用不公正的度量衡。
LEV|19|36|你們要用公正的天平、公正的法碼、公正的伊法和公正的欣。我是耶和華－你們的上帝，曾把你們從 埃及 地領出來。
LEV|19|37|你們要謹守我一切的律例典章，遵行它們。我是耶和華。」
LEV|20|1|耶和華吩咐 摩西 說：
LEV|20|2|「你要對 以色列 人說：凡 以色列 人，或是寄居在 以色列 的外人，把自己兒女獻給 摩洛 的，必被處死；本地的百姓要用石頭打死他。
LEV|20|3|我也要向那人變臉，把他從百姓中剪除，因為他把兒女獻給 摩洛 ，玷污了我的聖所，褻瀆了我的聖名。
LEV|20|4|那人把兒女獻給 摩洛 ，本地的百姓若假裝沒看見，不把他處死，
LEV|20|5|我就要向這人和他的家人變臉，把他和所有跟隨他與 摩洛 行淫的人都從百姓中剪除。
LEV|20|6|「人若轉向招魂的和行巫術的，隨從他們行淫，我就要向這人變臉，把他從百姓中剪除。
LEV|20|7|你們要使自己分別為聖，要成為聖，因為我是耶和華－你們的上帝。
LEV|20|8|你們要謹守我的律例，遵行它們；我是使你們分別為聖的耶和華。
LEV|20|9|凡咒罵父母的，必被處死；他咒罵了父母，他的血要歸在他身上。
LEV|20|10|「凡與有夫之婦行姦淫，就是與鄰舍的妻子行姦淫的，姦夫淫婦必被處死。
LEV|20|11|人若與繼母同寢，就是露了父親的下體，二人必被處死，血要歸在他們身上。
LEV|20|12|人若與媳婦同寢，二人必被處死；他們行了亂倫的事，血要歸在他們身上。
LEV|20|13|男人若跟男人同寢，像跟女人同寢，他們二人行了可憎惡的事，必被處死，血要歸在他們身上。
LEV|20|14|人若娶妻，又娶妻子的母親，這是邪惡的事；要把這三人用火焚燒，在你們中間除去這邪惡。
LEV|20|15|人若與獸交合，必被處死；你們也要殺死那獸。
LEV|20|16|女人若與獸親近，與牠交合，你要把那女人和獸殺死；他們必被處死，血要歸在他們身上。
LEV|20|17|「人若娶自己的姊妹，或是同父異母的，或是同母異父的，彼此見了下體，這是可恥的事；他們必在自己百姓眼前被剪除。他露了姊妹的下體，必擔當自己的罪孽。
LEV|20|18|若有人跟經期中的婦人同寢，露了她的下體，暴露婦人的血源，婦人也露了自己的血源，二人必從百姓中剪除。
LEV|20|19|不可露姨母或姑母的下體，因為這是露了骨肉之親的下體，他們必擔當自己的罪孽。
LEV|20|20|人若與叔伯之妻同寢，就露了他叔伯的下體，他們必擔當自己的罪，必沒有子女而死。
LEV|20|21|人若娶了自己兄弟的妻子，就露了他兄弟的下體，這是不潔淨的事，他們必沒有子女。
LEV|20|22|「你們要謹守我一切的律例典章，遵行它們，免得我領你們去住的那地把你們吐出來。
LEV|20|23|我在你們面前所逐出的國民，你們不可隨從他們的風俗。因為他們行了這一切的事，所以我厭惡他們。
LEV|20|24|但我對你們說過，你們要承受他們的土地；我要把這流奶與蜜之地賜給你們，作為你們的產業。我是耶和華－你們的上帝，是把你們從萬民中分別出來的。
LEV|20|25|你們要分辨潔淨和不潔淨的飛禽走獸；不可因我定為不潔淨的飛禽走獸，或爬行在土地上的任何生物，使自己成為可憎惡的。
LEV|20|26|你們要歸我為聖，因為－我耶和華是神聖的；我把你們從萬民中分別出來，作我的子民。
LEV|20|27|「無論男女，是招魂的或行巫術的，他們必被處死。人要用石頭打死他們，血要歸在他們身上。」
LEV|21|1|耶和華對 摩西 說：「你要告訴 亞倫 子孫作祭司的，對他們說：祭司不可為自己百姓中的死人玷污自己，
LEV|21|2|除非是他的骨肉之親，他的父母、兒女、兄弟、
LEV|21|3|或未出嫁還是處女的姊妹，因她是至親，才可以玷污自己。
LEV|21|4|祭司既然在自己百姓中為首，就不可從俗玷污自己 。
LEV|21|5|「不可使頭光禿，不可剃除鬍鬚的邊緣，也不可割劃自己的身體。
LEV|21|6|他們要歸上帝為聖，不可褻瀆他們上帝的名，因為耶和華的火祭，就是上帝的食物，是他們獻的，所以他們要成為聖。
LEV|21|7|「祭司不可娶妓女，或被玷污的女人為妻，也不可娶被休的婦人為妻，因為他是歸上帝為聖的。
LEV|21|8|你要使祭司分別為聖，因為他獻你上帝的食物。你要以他為聖，因為我是使你們分別為聖 的耶和華，是神聖的。
LEV|21|9|「祭司的女兒若行淫玷污自己，就侮辱了父親，要用火將她焚燒。
LEV|21|10|「在弟兄中作大祭司的，頭上倒了膏油，承接聖職，穿了聖衣，不可蓬頭散髮，也不可撕裂衣服；
LEV|21|11|不可挨近任何死屍，即使為了父母也不可玷污自己。
LEV|21|12|他不可出聖所，免得褻瀆了上帝的聖所，因為在他身上有上帝的膏油為聖冕。我是耶和華。
LEV|21|13|他要娶處女為妻。
LEV|21|14|大祭司不可娶寡婦，被休的婦人，或被玷污的妓女為妻；他只可以娶自己百姓中的處女為妻。
LEV|21|15|他不可在自己百姓中侮辱他的兒女，因為我是使他分別為聖的耶和華。」
LEV|21|16|耶和華吩咐 摩西 說：
LEV|21|17|「你吩咐 亞倫 說：你世世代代的後裔，凡有殘疾的都不可近前來獻上帝的食物。
LEV|21|18|因為凡有殘疾的，無論是失明的、瘸腿的、五官不正的、肢體之一過長的、
LEV|21|19|斷腳的、斷手的、
LEV|21|20|駝背的、侏儒的、有眼疾的、長癬的、長疥的，或是睪丸壓傷的，都不可近前來。
LEV|21|21|亞倫 祭司的後裔，凡有殘疾的都不可近前來獻耶和華的火祭。他有殘疾，不可近前來獻上帝的食物。
LEV|21|22|上帝的食物，無論是聖的，或是至聖的，他都可以吃。
LEV|21|23|但他不可進到幔子前，也不可挨近祭壇前，因為他有殘疾，免得他褻瀆我的聖所。我是使他們分別為聖的耶和華。」
LEV|21|24|於是， 摩西 吩咐了 亞倫 和他的兒子，以及 以色列 眾人。
LEV|22|1|耶和華吩咐 摩西 說：
LEV|22|2|「你要吩咐 亞倫 和他子孫說：你們要謹慎處理 以色列 人所分別為聖，歸給我的聖物，免得褻瀆我的聖名。我是耶和華。
LEV|22|3|你要對他們說：你們世世代代的後裔，凡不潔淨，卻挨近 以色列 人所分別為聖，歸給耶和華的聖物，那人必從我面前剪除。我是耶和華。
LEV|22|4|亞倫 的後裔中，凡有痲瘋病的，或患漏症的，都不可吃聖物，直等他潔淨了。無論誰摸了那因屍體而不潔淨的東西，或遺精的人，
LEV|22|5|或摸到任何使他不潔淨的群聚動物或使他不潔淨的人，無論那人有甚麼不潔淨，
LEV|22|6|摸了這些的人必不潔淨到晚上；若不用水洗身，就不可吃聖物。
LEV|22|7|日落的時候，他就潔淨了，然後可以吃聖物，因為這是他的食物。
LEV|22|8|自然死去的或被野獸撕裂的，他不可吃，免得玷污自己。我是耶和華。
LEV|22|9|他們要遵守我的吩咐，免得因褻瀆聖物 ，擔當自己的罪而死。我是使他們分別為聖的耶和華。
LEV|22|10|「任何外人都不可吃聖物；寄居在祭司家的，或雇工，都不可吃聖物。
LEV|22|11|若是祭司用自己的銀錢買來的人，就可以吃聖物；在他家出生的人也可以吃他的食物。
LEV|22|12|祭司的女兒若嫁給外人，就不可吃舉祭的聖物。
LEV|22|13|但祭司的女兒若成為寡婦或被休，又沒有後裔，她回到父家，好像年輕的時候，就可以吃她父親的食物。只是任何外人都不可吃它。
LEV|22|14|若有人誤吃了聖物，要把聖物加上五分之一交給祭司。
LEV|22|15|祭司不可褻瀆 以色列 人獻給耶和華的聖物，
LEV|22|16|免得他們因吃聖物而自取罪孽。我是使他們分別為聖的耶和華。」
LEV|22|17|耶和華吩咐 摩西 說：
LEV|22|18|「你要吩咐 亞倫 和他子孫，以及 以色列 眾人，對他們說： 以色列 家中的人，或在 以色列 中寄居的 ，若要獻供物給耶和華作燔祭，無論是為所許的願或是甘心獻的，
LEV|22|19|就要將一頭公的，沒有殘疾的牛，或綿羊，或山羊獻上，這樣你們才蒙悅納。
LEV|22|20|凡有殘疾的，你們不可獻上，因為這樣你們必不蒙悅納。
LEV|22|21|若有人從牛群或羊群中，將平安祭獻給耶和華，無論是為還所許特別的願，或是甘心獻的，所獻的必須是健康、無任何殘疾的，才蒙悅納。
LEV|22|22|凡瞎眼的、受傷的、斷腿的、潰爛的、長癬的、長疥的，都不可獻給耶和華，不可在壇上作為火祭獻給耶和華。
LEV|22|23|無論是公牛或小綿羊，若一條腿太長或太短，只可作甘心祭獻上；若用來還願，就不蒙悅納。
LEV|22|24|凡睪丸損傷，或壓碎，或破裂，或閹割的，都不可獻給耶和華；不可在你們的地上行這事。
LEV|22|25|從外人的手裏得到任何這類的動物，也不可獻上作你們上帝的食物；因為牠們有缺陷，有殘疾，牠們必不為你們而蒙悅納。」
LEV|22|26|耶和華吩咐 摩西 說：
LEV|22|27|「剛出生的公牛，或綿羊，或山羊，七天當跟著牠的母親；從第八天起，可以當供物作為耶和華的火祭，這是蒙悅納的。
LEV|22|28|無論是牛或羊，不可在同一日宰牠和牠的小牛小羊。
LEV|22|29|你們宰殺祭牲獻感謝祭給耶和華，要獻得使你們可蒙悅納；
LEV|22|30|要在當天吃，一點也不可留到早晨。我是耶和華。
LEV|22|31|「你們要謹守我的誡命，遵行它們。我是耶和華。
LEV|22|32|你們不可褻瀆我的聖名；我在 以色列 人中要被尊為聖。我是使你們分別為聖的耶和華，
LEV|22|33|曾把你們從 埃及 地領出來，作你們的上帝。我是耶和華。」
LEV|23|1|耶和華吩咐 摩西 說：
LEV|23|2|「你要吩咐 以色列 人，對他們說：以下是我的節期，是你們要宣告為聖會的耶和華的節期。」
LEV|23|3|「六日要做工，第七日是完全安息的安息日，要有聖會；你們任何工都不可做。這是在你們一切的住處向耶和華當守的安息日。」
LEV|23|4|「以下是你們要按時宣告為聖會的耶和華的節期。」
LEV|23|5|「正月十四日黃昏的時候 ，是向耶和華守的逾越節。
LEV|23|6|這月的十五日是向耶和華守的除酵節；你們要吃無酵餅七日。
LEV|23|7|第一日要有聖會，任何勞動的工都不可做；
LEV|23|8|要將火祭獻給耶和華七日。第七日要有聖會，任何勞動的工都不可做。」
LEV|23|9|耶和華吩咐 摩西 說：
LEV|23|10|「你要吩咐 以色列 人，對他們說：你們到了我賜給你們的地，收割莊稼的時候，要把初熟莊稼中的一捆拿來給祭司。
LEV|23|11|他要把這捆在耶和華面前搖一搖，使你們蒙悅納。祭司要在安息日的次日把這捆搖一搖。
LEV|23|12|搖這捆的那一日，你們要獻一隻一歲沒有殘疾的小公綿羊，給耶和華作燔祭。
LEV|23|13|同獻的素祭是十分之二伊法調了油的細麵，作為獻給耶和華馨香的火祭；同獻的澆酒祭是四分之一欣酒。
LEV|23|14|無論是餅，是烘熟的穀物，是新穗子，你們都不可吃；直等到你們把這供物帶來獻給你們上帝的那一天，才可以吃。在你們一切的住處，這要成為你們世世代代永遠的定例。」
LEV|23|15|「你們要從安息日的次日，就是獻那捆莊稼為搖祭的那日起，計算足足的七個安息日。
LEV|23|16|到第七個安息日的次日，共計五十天，你們要將新的素祭獻給耶和華。
LEV|23|17|要從你們的住處取十分之二伊法細麵，加酵烤成兩個搖祭的餅，作為初熟之物獻給耶和華。
LEV|23|18|又要將七隻一歲沒有殘疾的羔羊、一頭公牛犢、兩隻公綿羊和餅一同奉上。這些要和素祭和澆酒祭一同作為燔祭獻給耶和華，作馨香的火祭獻給耶和華。
LEV|23|19|你們要獻一隻公山羊為贖罪祭，兩隻一歲的小公綿羊為平安祭。
LEV|23|20|祭司要把這些和初熟莊稼做成的餅，與兩隻小公綿羊一同在耶和華面前搖一搖，作為搖祭。這些獻給耶和華的聖物是歸給祭司的。
LEV|23|21|在這一日，你們要宣告聖會；任何勞動的工都不可做。在你們一切的住處，這要成為你們世世代代永遠的定例。
LEV|23|22|「你們在自己的地收割莊稼時，不可割盡田的角落，也不可拾取莊稼所掉落的，要把它們留給窮人和寄居的。我是耶和華－你們的上帝。」
LEV|23|23|耶和華吩咐 摩西 說：
LEV|23|24|「你要吩咐 以色列 人說：七月初一，你們要守為完全安息的日子，要吹角作紀念，當有聖會。
LEV|23|25|任何勞動的工都不可做；要將火祭獻給耶和華。」
LEV|23|26|耶和華吩咐 摩西 說：
LEV|23|27|「但是，七月初十是贖罪日；你們要守為聖會，刻苦己心，並要將火祭獻給耶和華。
LEV|23|28|在這一日，任何工都不可做；因為這是贖罪日，要在耶和華－你們的上帝面前贖罪。
LEV|23|29|在這一日，凡不刻苦己心的，必從百姓中剪除。
LEV|23|30|凡在這一日做任何工的，我必將他從百姓中除滅。
LEV|23|31|任何工你們都不可做。在你們一切的住處，這要成為你們世世代代永遠的定例。
LEV|23|32|你們要守這日為完全安息的安息日，刻苦己心；從這月初九晚上到次日晚上，你們要守為安息日。」
LEV|23|33|耶和華吩咐 摩西 說：
LEV|23|34|「你要吩咐 以色列 人說：這七月十五日是住棚節，要向耶和華守這節七日。
LEV|23|35|第一日當有聖會，任何勞動的工都不可做。
LEV|23|36|要將火祭獻給耶和華七日。第八日當守聖會，並要獻火祭給耶和華。這是嚴肅會，任何勞動的工都不可做。
LEV|23|37|「這是耶和華的節期，就是你們要宣告為聖會的節期；要將火祭，就是燔祭、素祭、祭物和澆酒祭，按照每日的規定獻給耶和華。
LEV|23|38|除此之外，還有耶和華的安息日，你們獻給耶和華的供物，一切的還願祭，和一切的甘心祭。
LEV|23|39|「但是，從七月十五日起，你們收藏了地的出產之後，要守耶和華的節期七日。第一日為要完全安息，第八日也要完全安息。
LEV|23|40|第一日，你們要拿美好樹上的果子、棕樹枝、樹葉茂密的枝條和河邊的柳枝，在耶和華－你們的上帝面前歡樂七日。
LEV|23|41|每年你們要向耶和華守這節七日。你們在七月裏所守的節，要成為世世代代永遠的定例。
LEV|23|42|你們要住在棚裏七日；凡 以色列 家出生的人都要住在棚裏，
LEV|23|43|好叫你們世世代代知道，我領 以色列 人出 埃及 地的時候，曾使他們住在棚裏。我是耶和華－你們的上帝。」
LEV|23|44|於是， 摩西 向 以色列 人頒佈了耶和華的節期。
LEV|24|1|耶和華吩咐 摩西 說：
LEV|24|2|「你要吩咐 以色列 人，把那搗成的純橄欖油拿來給你，用以點燈，使燈經常點著。
LEV|24|3|在會幕中法櫃前的幔子外， 亞倫 從晚上到早晨要在耶和華面前照管這燈。這要成為你們世世代代永遠的定例。
LEV|24|4|他要在耶和華面前經常照管純金 燈臺上的燈。」
LEV|24|5|「你要取細麵，烤成十二個餅，每個用十分之二伊法。
LEV|24|6|要把餅排成兩行 ，每行六個，供在耶和華面前的純金桌子上。
LEV|24|7|再把純乳香撒在每行餅上，作為紀念，是獻給耶和華為食物的火祭。
LEV|24|8|每個安息日， 亞倫 要把餅不間斷地供在耶和華面前。這是 以色列 人永遠的約。
LEV|24|9|這餅要歸給 亞倫 和他的子孫。他們要在聖處吃這餅，因為在獻給耶和華的火祭中，這餅是至聖的，歸給他作永遠當得的份。」
LEV|24|10|有一個 以色列 婦人的兒子，他父親是 埃及 人。有一日他出去，到 以色列 人中。這 以色列 婦人的兒子和一個 以色列 人在營裏爭吵。
LEV|24|11|以色列 婦人的兒子詛咒，褻瀆了聖名。有人把他送到 摩西 那裏。他的母親名叫 示羅密 ，是 但 支派 底伯利 的女兒。
LEV|24|12|他們把這人收押在監裏，等候耶和華指示的話。
LEV|24|13|耶和華吩咐 摩西 說：
LEV|24|14|「把那詛咒的人帶到營外。凡聽見的人都要把手放在他頭上，全會眾要用石頭打死他。
LEV|24|15|你要吩咐 以色列 人說：凡詛咒上帝的，必要擔當自己的罪。
LEV|24|16|褻瀆耶和華名的，必被處死；全會眾必須用石頭打死他。無論是寄居的，是本地人，他褻瀆聖名的時候必被處死。
LEV|24|17|「打死人的，必被處死；
LEV|24|18|打死牲畜的，必賠上牲畜，以命償命。
LEV|24|19|人若傷害鄰舍以致殘疾，他怎樣做，也要照樣向他做：
LEV|24|20|以傷還傷，以眼還眼，以牙還牙。他怎樣使人有殘疾，也要照樣向他做。
LEV|24|21|打死牲畜的，必賠上牲畜；打死人的，必被處死。
LEV|24|22|無論是寄居的，是本地人，都依照同一條例。我是耶和華－你們的上帝。」
LEV|24|23|於是， 摩西 吩咐 以色列 人，他們就把那詛咒的人帶到營外，用石頭打死。 以色列 人就照耶和華所吩咐 摩西 的做了。
LEV|25|1|耶和華在 西奈山 吩咐 摩西 說：
LEV|25|2|「你要吩咐 以色列 人，對他們說：你們到了我所賜你們那地的時候，地要休耕，向耶和華守安息。
LEV|25|3|你們六年要耕種田地，六年要修整葡萄園，收藏地的出產。
LEV|25|4|第七年，地要守完全安息的安息年，就是向耶和華守安息。你們不可耕種田地，也不可修整葡萄園。
LEV|25|5|不可收割自然生長的莊稼，也不可摘取沒有修剪的葡萄樹上的葡萄。這年，地要完全安息。
LEV|25|6|地在安息年所長出的，要給你和你的奴僕、使女、雇工，以及寄居在你那裏的外人作食物。
LEV|25|7|所有的出產也要給你的牲畜和你地上的走獸作食物。」
LEV|25|8|「你要計算七個安息年，就是七個七年。這就成為你的七個安息年，一共四十九年。
LEV|25|9|七月初十，你要大聲吹角；這是贖罪日，你要在全地吹角。
LEV|25|10|你們要以第五十年為聖年，在全地向所有的居民宣告自由。這是你們的禧年，各人的產業要歸還自己，各人要歸回自己的家。
LEV|25|11|第五十年要作為你們的禧年。你們不可耕種，不可收割自然生長的莊稼，也不可摘取沒有修剪的葡萄樹上的葡萄。
LEV|25|12|因為這是禧年，是你們的聖年；你們要吃地中自然生長的農作物。
LEV|25|13|「這禧年，你們各人的產業要歸還自己。
LEV|25|14|無論你賣甚麼給鄰舍，或從鄰舍的手中買甚麼，彼此不可虧負。
LEV|25|15|你要按照禧年後的年數向鄰舍買；他要按照可收成的年數賣給你；
LEV|25|16|年數越多，價錢就越高；年數越少，價錢就越低，因為他賣給你的是收成的數量。
LEV|25|17|你們彼此不可虧負，只要敬畏你的上帝，因為我是耶和華－你們的上帝。」
LEV|25|18|「你們要遵行我的律例，謹守我的典章，遵行它們，就可以在那地上安然居住。
LEV|25|19|地必出產果實，你們可以吃飽，在那地上安然居住。
LEV|25|20|你們若說：『看哪，第七年我們不耕種，也不收藏農作物，我們吃甚麼呢？』
LEV|25|21|我必在第六年發令賜福給你們，地就長出三年的農作物來。
LEV|25|22|第八年你們要耕種，也要吃陳糧；等到第九年農作物收成的時候，你們還有陳糧吃。」
LEV|25|23|「地不可以賣斷，因為地是我的；你們在我面前是客旅，是寄居的。
LEV|25|24|在你們所得為業的全地，要准許人有權將地贖回。
LEV|25|25|「你的弟兄若漸漸貧窮，賣了他的一些產業，他的至親就要來把弟兄所賣的贖回。
LEV|25|26|若沒有人能為他贖回，他的手頭漸漸寬裕，能夠贖回，
LEV|25|27|就要計算賣後的年數，把剩餘年數的價錢歸還給那買主，他的地業便歸還自己。
LEV|25|28|若他手頭的財力不夠贖回，所賣的地就要留在買主的手裏，直到禧年。到了禧年，地業要歸還賣主。
LEV|25|29|「人若賣城牆內的住宅，賣了以後，一整年內他有權贖回；這是他可以贖回的期限。
LEV|25|30|若他在一整年內不贖回，這有牆之城的房屋就確定永歸買主，直到世世代代；在禧年也不必歸還。
LEV|25|31|但周圍無城牆之村莊的房屋，要看為鄉下的田地，可以贖回；到了禧年就要歸還。
LEV|25|32|至於 利未 人所得為業的城鎮， 利未 人可以隨時贖回他們城鎮中的房屋。
LEV|25|33|在所得為業的城鎮， 利未 人若賣了房屋，又不贖回，到了禧年仍要歸還原主，因為 利未 人城鎮的房屋是他們在 以色列 人中的產業。
LEV|25|34|但是 利未 人各城郊外之地是不可賣的，因為這是他們永遠的產業。」
LEV|25|35|「你的弟兄在你那裏若漸漸貧窮，手頭缺乏，你就要幫補他，使他與你一同生活，像外人和寄居的一樣。
LEV|25|36|不可向他取利息，也不可向他索取高利；要敬畏你的上帝，使你的弟兄與你一同生活。
LEV|25|37|你不可為了利息借錢給他，也不可為了高利而借糧。
LEV|25|38|我是耶和華－你們的上帝，曾領你們從 埃及 地出來，為要把 迦南 地賜給你們，要作你們的上帝。
LEV|25|39|「你的弟兄在你那裏若漸漸貧窮，將自己賣給你，你不可叫他像奴僕服事你。
LEV|25|40|他在你那裏要像雇工和寄居的，服事你直到禧年。
LEV|25|41|他和他兒女要離開你，一同出去，歸回自己的家，回到他祖宗的地業去。
LEV|25|42|因為他們是我的僕人，是我從 埃及 地領出來的。他們不可被賣為奴僕。
LEV|25|43|不可苛刻管轄他，只要敬畏你的上帝。
LEV|25|44|至於你所要的奴僕和使女，可以來自你們四圍的列國，你們可以從他們中買奴僕和使女。
LEV|25|45|那些寄居在你們中間的外人和他們的家屬，就是在你們地上所生的，你們可以從其中買人；他們要作你們的產業。
LEV|25|46|你們可以把他們遺留給你們後代的子孫，作為永遠繼承的產業；你們可以使他們作奴僕。至於你們的弟兄 以色列 人，你們彼此不可苛刻管轄。
LEV|25|47|「住在你那裏的外人或寄居的，若手頭漸漸寬裕，你的弟兄卻漸漸貧窮，將自己賣給那外人或寄居的，或外人家族的一支，
LEV|25|48|賣了以後，有權把自己贖回。他弟兄中的一位可以把他贖回。
LEV|25|49|他的叔伯或叔伯的兒子可以贖他。他家族中的骨肉之親也可以贖他。他自己若手頭漸漸寬裕，也可以贖回自己。
LEV|25|50|他要跟買主計算，從賣自己的那年起，算到禧年；所賣的價錢要按照年數計算，就是雇工跟買主在一起的日子。
LEV|25|51|若剩餘的年數多，就要按著年數從買價中償還他的贖價。
LEV|25|52|若到禧年只剩下幾年，就要按著年數跟買主計算，償還他的贖價。
LEV|25|53|他和買主同住，要像按年雇用的工人，買主不可苛刻管轄他。
LEV|25|54|他若不這樣被贖，到了禧年，仍要和他的兒女一同出去。
LEV|25|55|因為 以色列 人都是我的僕人，他們是我的僕人，是我領他們從 埃及 地出來的。我是耶和華－你們的上帝。」
LEV|26|1|「你們不可為自己造虛無的神明，不可豎立雕刻的偶像或柱像，也不可在你們的地上安放石像，向它跪拜，因為我是耶和華－你們的上帝。
LEV|26|2|你們要謹守我的安息日，敬畏我的聖所。我是耶和華。
LEV|26|3|「你們若遵行我的律例，謹守我的誡命，實行它們，
LEV|26|4|我必按時降雨給你們，使地長出農作物，田野的樹結出果實。
LEV|26|5|你們打穀物要打到摘葡萄的時候，摘葡萄要摘到播種的時候。你們要吃糧食得飽足，在你們的地上安然居住。
LEV|26|6|我要賜平安在地上；你們躺臥，無人驚嚇。我要使你們地上的惡獸消滅，刀劍必不穿越你們的地。
LEV|26|7|你們要追趕仇敵，他們必倒在你們刀下。
LEV|26|8|你們五個人要追趕一百人，一百人要追趕一萬人；仇敵必在你們面前倒在刀下。
LEV|26|9|我要眷顧你們，使你們生養眾多，也要與你們堅立我的約。
LEV|26|10|你們要吃儲存的陳糧，又要為新糧清理陳糧。
LEV|26|11|我要在你們中間立我的帳幕，我的心也不厭惡你們。
LEV|26|12|我要行走在你們中間，作你們的上帝，你們要作我的子民。
LEV|26|13|我是耶和華－你們的上帝，曾將你們從 埃及 地領出來，使你們不再作 埃及 人的奴僕；我曾折斷你們所負的軛，使你們挺身前行。」
LEV|26|14|「你們若不聽從我，不遵行我這一切的誡命，
LEV|26|15|厭棄我的律例，心中厭惡我的典章，不遵行我一切的誡命，背棄了我的約，
LEV|26|16|我就要這樣對待你們：我必使驚惶臨到你們，使你們患癆病，害熱病，以致眼睛失明，身體衰弱。你們要白白撒種，因為仇敵要吃盡你們所種的。
LEV|26|17|我要向你們變臉，使你們敗在仇敵的面前。恨惡你們的必管轄你們；無人追趕，你們卻要逃跑。
LEV|26|18|如果這樣，你們還不聽從我，我就要因你們的罪，加重七倍懲罰你們。
LEV|26|19|我必粉碎你們因勢力而有的驕傲，又要使你們的天堅如鐵，地硬如銅。
LEV|26|20|你們勞力卻白費，因為你們的地沒有出產，地上的樹也不結果實。
LEV|26|21|「你們行事若與我作對，不肯聽從我，我就要因你們的罪，加重七倍災禍擊打你們。
LEV|26|22|我要打發野地的走獸到你們中間，奪去你們的兒女，吞滅你們的牲畜，使你們人數減少，道路荒涼。
LEV|26|23|「如果這樣，你們還不接受管教歸向我，行事與我作對，
LEV|26|24|我就要行事與你們作對，因你們的罪，加重七倍擊打你們。
LEV|26|25|我要使刀劍臨到你們，報復你們的背約。你們若被趕入城中，我要降瘟疫在你們中間，把你們交在仇敵手中。
LEV|26|26|我要斷絕你們糧食的供應 ，使十個女人用一個烤爐給你們烤餅，按配給的定量秤給你們。你們要吃，卻吃不飽。
LEV|26|27|「如果這樣，你們還不聽從我，行事與我作對，
LEV|26|28|我就要向你們發烈怒，行事與你們作對，因你們的罪，加重七倍懲罰你們。
LEV|26|29|你們要吃你們兒子的肉，也要吃你們女兒的肉。
LEV|26|30|我要摧毀你們的丘壇，砍掉你們的香壇，把你們的屍首扔在你們偶像的殘骸上。我的心也必厭惡你們，
LEV|26|31|使你們的城鎮變成廢墟，你們的眾聖所變荒涼，我也不聞你們芬芳的香氣。
LEV|26|32|我要使這地變荒涼，甚至佔領這地的敵人都驚訝。
LEV|26|33|我要把你們驅散到列國中，也要拔刀追趕你們。你們的地要成為荒涼，你們的城鎮要變成廢墟。
LEV|26|34|「當你們在敵人之地的時候，你們的地要在一切荒涼的日子重享安息；在那時候，地要休息，重享安息。
LEV|26|35|地在一切荒涼的日子都要安息，這是你們住在其上的時候所不能得的安息。
LEV|26|36|至於你們倖存的人，我要使他們在敵人之地心中驚慌，甚至風吹落葉的聲音也把他們嚇跑。他們要逃避，像人逃避刀劍，雖無人追趕，卻要跌倒。
LEV|26|37|雖然無人追趕，他們卻要彼此絆倒，像逃避刀劍一樣。你們在仇敵面前必站立不住。
LEV|26|38|你們要在列國中滅亡，敵人之地要吞滅你們，
LEV|26|39|你們倖存的人必因自己的罪孽在敵人之地衰殘，也要因祖先的罪孽衰殘。
LEV|26|40|「他們要承認自己的罪孽和祖先的罪孽，就是背叛我，行事與我作對的過犯。
LEV|26|41|我也行事與他們作對，把他們遣送到敵人之地。那時，他們未受割禮的心若肯謙卑，也服了罪孽的懲罰，
LEV|26|42|我就要記念我與 雅各 的約，記念我與 以撒 的約，與 亞伯拉罕 的約；我也要記念這地。
LEV|26|43|地被他們離棄，因他們不在而荒涼的時候，就要重享安息。他們服了罪孽的懲罰，因為他們厭棄我的典章，心中厭惡我的律例。
LEV|26|44|雖然如此，當他們在敵人之地時，我卻不厭棄他們，不厭惡他們，將他們全然滅絕，也不背棄我與他們的約，因為我是耶和華－他們的上帝。
LEV|26|45|我要為他們的緣故記念我與他們祖先的約；我在列國眼前曾把他們的祖先從 埃及 地領出來，為要作他們的上帝。我是耶和華。」
LEV|26|46|這些律例、典章和法度是耶和華在 西奈山 上藉著 摩西 與 以色列 人立的。
LEV|27|1|耶和華吩咐 摩西 說：
LEV|27|2|「你要吩咐 以色列 人，對他們說：人向耶和華許特別的願，要按照你所估一個人的價錢。
LEV|27|3|你所估的是：二十歲到六十歲男的，按照聖所的舍客勒，估價是五十舍客勒銀子。
LEV|27|4|若是女的，估價是三十舍客勒。
LEV|27|5|五歲到二十歲男的，估價是二十舍客勒，女的十舍客勒。
LEV|27|6|一個月到五歲男的，估價是五舍客勒，女的三舍客勒。
LEV|27|7|六十歲以上男的，估價是十五舍客勒，女的十舍客勒。
LEV|27|8|他若貧窮，不能按照你的估價，就要把他帶到祭司面前，讓祭司為他估價；祭司要按許願者手頭財力所及估價。
LEV|27|9|「許願要獻給耶和華的供物若是牲畜，凡這類獻給耶和華的都要成為聖。
LEV|27|10|不可更換，也不可用另一隻取代，無論是好的換壞的，或是壞的換好的，都不可。若一定要以牲畜取代牲畜，所許的與所取代的都要成為聖。
LEV|27|11|若牲畜不潔淨，不可獻給耶和華為供物，就要把牲畜帶到祭司面前。
LEV|27|12|祭司要估價；牲畜是好是壞，祭司怎樣估定，就是你的估價。
LEV|27|13|許願者若一定要把牠贖回，就要在你的估價上加五分之一。
LEV|27|14|「人將房屋分別為聖，歸給耶和華為聖，祭司就要估價。房屋是好是壞，祭司怎樣估定，就要以他的估價為準。
LEV|27|15|將房屋分別為聖的人，若要贖回房屋，必須付你所估定的價錢，再加上五分之一，房屋才可以歸還給他。
LEV|27|16|「人若將所繼承的一塊田地分別為聖，歸給耶和華，就要按照這地撒種多少來估價；能撒一賀梅珥大麥種子的，是五十舍客勒銀子。
LEV|27|17|他若從禧年起將地分別為聖，就要以你的估價為準。
LEV|27|18|倘若他在禧年以後將地分別為聖，祭司就要按照從那時到下一個禧年所剩的年數推算，從你的估價中減掉。
LEV|27|19|將地分別為聖的人若要把地贖回，必須付你所估定的價錢，再加上五分之一，地才可以歸還給他。
LEV|27|20|他若不贖回那地，或是將地賣給別人，就不能再贖了。
LEV|27|21|到了禧年，那田地要從買主手中退還，歸耶和華為聖，和永獻的地一樣，要歸祭司為業。
LEV|27|22|若分別為聖歸耶和華的田地不是繼承的，而是買來的，
LEV|27|23|祭司就要依照你的估價，推算到禧年。當天，這人要將你所估的歸給耶和華為聖。
LEV|27|24|到了禧年，那田地要退還給賣主，就是繼承那地的原主。
LEV|27|25|凡你所估的價錢都要按照聖所的舍客勒：二十季拉是一舍客勒。
LEV|27|26|「頭生的，就是牲畜中頭生屬耶和華的，人不可再將牠分別為聖，無論是牛是羊都是耶和華的。
LEV|27|27|頭生的牲畜若是不潔淨的，就要按照所估定的價錢，再加上五分之一，把牠贖回。若不贖回，就要按照你的估價把牠賣了。
LEV|27|28|「但一切永獻作當滅的，就是人從他所有永獻給耶和華作當滅的，無論是人，是牲畜，是他繼承的田地，都不可賣，也不可贖。凡永獻作當滅的都歸耶和華為至聖。
LEV|27|29|凡從人中永獻作當滅的都不可贖，必被處死。
LEV|27|30|「地上所有的，無論是地上的種子，是樹上的果子，十分之一是耶和華的，是歸耶和華為聖的。
LEV|27|31|人若要贖回這十分之一，就要另加五分之一。
LEV|27|32|凡牛群羊群中的十分之一，就是一切從牧人杖下經過的，每第十隻要歸耶和華為聖。
LEV|27|33|不可追究是好是壞，也不可取代；若一定要取代，所取代的和本來當獻的牲畜都要成為聖，不可贖回。」
LEV|27|34|這些是耶和華在 西奈山 為 以色列 人所吩咐 摩西 的命令。
NUM|1|1|以色列 人出 埃及 地後第二年二月初一，耶和華在 西奈 曠野，在會幕中吩咐 摩西 說：
NUM|1|2|「你要按宗族、父家、人名的數目計算 以色列 全會眾，數點所有的男丁。
NUM|1|3|以色列 中凡二十歲以上能出去打仗的，你和 亞倫 要按照他們的隊伍數點。
NUM|1|4|每支派要有一個人，就是父家的家長跟你們一起。
NUM|1|5|這是幫助你們的人的名字： 屬 呂便 的， 示丟珥 的兒子 以利蓿 ；
NUM|1|6|屬 西緬 的， 蘇利沙代 的兒子 示路蔑 ；
NUM|1|7|屬 猶大 的， 亞米拿達 的兒子 拿順 ；
NUM|1|8|屬 以薩迦 的， 蘇押 的兒子 拿坦業 ；
NUM|1|9|屬 西布倫 的， 希倫 的兒子 以利押 ；
NUM|1|10|約瑟 子孫、屬 以法蓮 的， 亞米忽 的兒子 以利沙瑪 ；屬 瑪拿西 的， 比大蓿 的兒子 迦瑪列 ；
NUM|1|11|屬 便雅憫 的， 基多尼 的兒子 亞比但 ；
NUM|1|12|屬 但 的， 亞米沙代 的兒子 亞希以謝 ；
NUM|1|13|屬 亞設 的， 俄蘭 的兒子 帕結 ；
NUM|1|14|屬 迦得 的， 丟珥 的兒子 以利雅薩 ；
NUM|1|15|屬 拿弗他利 的， 以南 的兒子 亞希拉 。」
NUM|1|16|這些是從會眾中選出來的父系支派的領袖，是 以色列 部隊的官長。
NUM|1|17|於是， 摩西 和 亞倫 帶著這些按名指定的人，
NUM|1|18|在二月初一召集全會眾。會眾就照他們的宗族、父家、人名的數目，登記二十歲以上的人口。
NUM|1|19|耶和華怎樣吩咐 摩西 ，他就照樣在 西奈 的曠野數點他們。
NUM|1|20|以色列 的長子， 呂便 子孫的後代，照著宗族、父家、人名的數目，他們的人口凡二十歲以上能出去打仗的男丁，
NUM|1|21|呂便 支派被數的共有四萬六千五百名。
NUM|1|22|西緬 子孫的後代，照著宗族、父家、被數 人名的數目，他們的人口凡二十歲以上能出去打仗的男丁，
NUM|1|23|西緬 支派被數的共有五萬九千三百名。
NUM|1|24|迦得 子孫的後代，照著宗族、父家、人名的數目，凡二十歲以上能出去打仗的，
NUM|1|25|迦得 支派被數的共有四萬五千六百五十名。
NUM|1|26|猶大 子孫的後代，照著宗族、父家、人名的數目，凡二十歲以上能出去打仗的，
NUM|1|27|猶大 支派被數的共有七萬四千六百名。
NUM|1|28|以薩迦 子孫的後代，照著宗族、父家、人名的數目，凡二十歲以上能出去打仗的，
NUM|1|29|以薩迦 支派被數的共有五萬四千四百名。
NUM|1|30|西布倫 子孫的後代，照著宗族、父家、人名的數目，凡二十歲以上能出去打仗的，
NUM|1|31|西布倫 支派被數的共有五萬七千四百名。
NUM|1|32|約瑟 子孫屬 以法蓮 子孫的後代，照著宗族、父家、人名的數目，凡二十歲以上能出去打仗的，
NUM|1|33|以法蓮 支派被數的共有四萬零五百名。
NUM|1|34|瑪拿西 子孫的後代，照著宗族、父家、人名的數目，凡二十歲以上能出去打仗的，
NUM|1|35|瑪拿西 支派被數的共有三萬二千二百名。
NUM|1|36|便雅憫 子孫的後代，照著宗族、父家、人名的數目，凡二十歲以上能出去打仗的，
NUM|1|37|便雅憫 支派被數的共有三萬五千四百名。
NUM|1|38|但 子孫的後代，照著宗族、父家、人名的數目，凡二十歲以上能出去打仗的，
NUM|1|39|但 支派被數的共有六萬二千七百名。
NUM|1|40|亞設 子孫的後代，照著宗族、父家、人名的數目，凡二十歲以上能出去打仗的，
NUM|1|41|亞設 支派被數的共有四萬一千五百名。
NUM|1|42|拿弗他利 子孫的後代，照著宗族、父家、人名的數目，凡二十歲以上能出去打仗的，
NUM|1|43|拿弗他利 支派被數的共有五萬三千四百名。
NUM|1|44|這些就是被數點的，是 摩西 、 亞倫 和 以色列 十二個領袖所數點的；每一個領袖代表他們的父家。
NUM|1|45|以色列 人被數點的總數， 以色列 中照著父家，凡二十歲以上能出去打仗的，
NUM|1|46|他們被數點的總數是六十萬三千五百五十名。
NUM|1|47|利未 人卻沒有按照父系支派數在其中。
NUM|1|48|耶和華吩咐 摩西 說：
NUM|1|49|「惟獨 利未 支派你不可數點，也不可在 以色列 人中計算他們的人口。
NUM|1|50|你要派 利未 人管理法櫃的帳幕和其中一切的器具，以及屬帳幕的一切。他們要抬帳幕和其中一切的器具，並要辦理帳幕的事務，在帳幕的四圍安營。
NUM|1|51|帳幕將往前行的時候， 利未 人要拆卸；將駐紮的時候， 利未 人要支搭帳幕。近前來的外人必被處死。
NUM|1|52|以色列 人要按照各自的隊伍安營，各歸本營，各歸本旗。
NUM|1|53|但 利未 人要在法櫃帳幕的四圍安營，免得憤怒臨到 以色列 會眾； 利未 人要負責看守法櫃的帳幕。」
NUM|1|54|以色列 人就這樣做了。凡耶和華所吩咐 摩西 的，他們都照樣做了。
NUM|2|1|耶和華吩咐 摩西 和 亞倫 說：
NUM|2|2|「 以色列 人各人要在自己的旗幟下，按照自己父家的旗號安營，對著會幕的四圍安營。
NUM|2|3|「在東邊，向日出的方向， 猶大 營按照他們的隊伍，在它的旗幟下安營。 猶大 人的領袖是 亞米拿達 的兒子 拿順 ，
NUM|2|4|他的軍隊被數的有七萬四千六百名。
NUM|2|5|在他旁邊安營的是 以薩迦 支派。 以薩迦 人的領袖是 蘇押 的兒子 拿坦業 ，
NUM|2|6|他的軍隊被數的有五萬四千四百名。
NUM|2|7|還有 西布倫 支派， 西布倫 人的領袖是 希倫 的兒子 以利押 ，
NUM|2|8|他的軍隊被數的有五萬七千四百名。
NUM|2|9|凡屬 猶大 營，照他們隊伍被數的共有十八萬六千四百名；他們要作第一隊往前行。
NUM|2|10|「在南邊，按照他們的隊伍是 呂便 營的旗幟。 呂便 人的領袖是 示丟珥 的兒子 以利蓿 ，
NUM|2|11|他的軍隊被數的有四萬六千五百名。
NUM|2|12|在他旁邊安營的是 西緬 支派。 西緬 人的領袖是 蘇利沙代 的兒子 示路蔑 ，
NUM|2|13|他的軍隊被數的有五萬九千三百名。
NUM|2|14|還有 迦得 支派， 迦得 人的領袖是 丟珥 的兒子 以利雅薩 ，
NUM|2|15|他的軍隊被數的有四萬五千六百五十名。
NUM|2|16|凡屬 呂便 營，照他們隊伍被數的共有十五萬一千四百五十名；他們要作第二隊往前行。
NUM|2|17|「會幕與 利未 營在諸營中間往前行。他們怎樣安營就怎樣往前行，各按本位，各歸本旗。
NUM|2|18|「在西邊，按照他們的隊伍是 以法蓮 營的旗幟。 以法蓮 人的領袖是 亞米忽 的兒子 以利沙瑪 ，
NUM|2|19|他的軍隊被數的有四萬零五百名。
NUM|2|20|在他旁邊的是 瑪拿西 支派。 瑪拿西 人的領袖是 比大蓿 的兒子 迦瑪列 ，
NUM|2|21|他的軍隊被數的有三萬二千二百名。
NUM|2|22|還有 便雅憫 支派， 便雅憫 人的領袖是 基多尼 的兒子 亞比但 ，
NUM|2|23|他的軍隊被數的有三萬五千四百名。
NUM|2|24|凡屬 以法蓮 營，照他們隊伍被數的共有十萬八千一百名；他們要作第三隊往前行。
NUM|2|25|「在北邊，按照他們的隊伍是 但 營的旗幟。 但 人的領袖是 亞米沙代 的兒子 亞希以謝 ，
NUM|2|26|他的軍隊被數的有六萬二千七百名。
NUM|2|27|在他旁邊安營的是 亞設 支派。 亞設 人的領袖是 俄蘭 的兒子 帕結 ，
NUM|2|28|他的軍隊被數的有四萬一千五百名。
NUM|2|29|還有 拿弗他利 支派， 拿弗他利 人的領袖是 以南 的兒子 亞希拉 ，
NUM|2|30|他的軍隊被數的有五萬三千四百名。
NUM|2|31|凡屬 但 營被數的共有十五萬七千六百名；他們隨著自己的旗幟行在最後。」
NUM|2|32|以上是 以色列 人按照各自的父家被數的，在諸營中按照各自的隊伍被數的，共有六十萬三千五百五十名。
NUM|2|33|但 利未 人沒有數在 以色列 人中，正如耶和華所吩咐 摩西 的。
NUM|2|34|以色列 人就照著耶和華所吩咐 摩西 的做了，在各自的旗幟下安營，隨著各自的宗族、父家起行。
NUM|3|1|耶和華在 西奈山 與 摩西 說話的日子， 亞倫 和 摩西 的後代如下：
NUM|3|2|這些是 亞倫 兒子的名字，長子 拿答 ，及 亞比戶 、 以利亞撒 、 以他瑪 。
NUM|3|3|這些是 亞倫 兒子的名字，都是受膏的祭司，是 摩西 授聖職使他們擔任祭司職分的。
NUM|3|4|拿答 、 亞比戶 在 西奈 的曠野向耶和華獻上凡火的時候，死在耶和華面前。他們沒有兒子。 以利亞撒 和 以他瑪 在他們的父親 亞倫 面前擔任祭司的職分。
NUM|3|5|耶和華吩咐 摩西 說：
NUM|3|6|「你要帶 利未 支派近前來，站在 亞倫 祭司面前伺候他。
NUM|3|7|他們要替他，又替全會眾，在會幕前執行任務，辦理帳幕的事。
NUM|3|8|他們要看守會幕一切的器具，為 以色列 人執行任務，辦理帳幕的事。
NUM|3|9|你要把 利未 人給 亞倫 和他的兒子；他們是從 以色列 人中選出來完全給他的。
NUM|3|10|你要指派 亞倫 和他的兒子謹守祭司的職分；近前來的外人必被處死。」
NUM|3|11|耶和華吩咐 摩西 說：
NUM|3|12|「看哪，我從 以色列 人中選了 利未 人，代替 以色列 人中所有頭胎的長子； 利未 人要歸我。
NUM|3|13|因為凡頭生的是我的；我在 埃及 地擊殺所有頭生的那日，就把 以色列 中所有頭生的，無論是人或牲畜，都分別為聖歸我；他們定要屬我。我是耶和華。」
NUM|3|14|耶和華在 西奈 的曠野吩咐 摩西 說：
NUM|3|15|「你要照父家、宗族計算 利未 人。凡一個月以上的男子都要數點。」
NUM|3|16|於是 摩西 遵照耶和華的吩咐，按所指示的數點他們。
NUM|3|17|利未 兒子的名字是 革順 、 哥轄 、 米拉利 。
NUM|3|18|按照宗族， 革順 兒子的名字是 立尼 、 示每 。
NUM|3|19|按照宗族， 哥轄 的兒子是 暗蘭 、 以斯哈 、 希伯倫 、 烏薛 。
NUM|3|20|按照宗族， 米拉利 的兒子是 抹利 、 母示 。按照父家，這些都是 利未 人的宗族。
NUM|3|21|屬 革順 的有 立尼 族、 示每 族，他們是 革順 人的宗族。
NUM|3|22|他們被數的，一個月以上所有男子的數目共有七千五百名。
NUM|3|23|這 革順 人的宗族要在西邊，在帳幕後面安營。
NUM|3|24|革順 人父家的領袖是 拉伊勒 的兒子 以利雅薩 。
NUM|3|25|革順 的子孫在會幕中要看守的是帳幕、罩棚、罩棚的蓋、會幕的門簾、
NUM|3|26|帳幕和祭壇周圍院子的帷幔和門簾，以及所有需用的繩子。
NUM|3|27|屬 哥轄 的有 暗蘭 族、 以斯哈 族、 希伯倫 族、 烏薛 族，他們是 哥轄 人的宗族。
NUM|3|28|一個月以上所有男子的數目共有八千六百 名；他們負責看守聖所。
NUM|3|29|哥轄 子孫的宗族要在帳幕的南邊安營。
NUM|3|30|哥轄 人父家宗族的領袖是 烏薛 的兒子 以利撒反 。
NUM|3|31|他們要看守的是約櫃、供桌、燈臺、祭壇、香壇、祭司在聖所內用的器皿、簾子，與一切相關事奉的物件。
NUM|3|32|亞倫 祭司的兒子 以利亞撒 是 利未 人眾領袖的主管，他要監督那些負責看守聖所的人。
NUM|3|33|屬 米拉利 的有 抹利 族、 母示 族，他們是 米拉利 的宗族。
NUM|3|34|他們被數的，一個月以上所有男子的數目共有六千二百名。
NUM|3|35|米拉利 宗族的領袖是 亞比亥 的兒子 蘇列 ，他們要在帳幕的北邊安營。
NUM|3|36|米拉利 子孫的職分是看守帳幕的豎板、橫木、柱子、帶卯眼的座和一切的器具，就是一切相關事奉的物件，
NUM|3|37|以及院子四圍的柱子、其上帶卯眼的座、橛子和繩子。
NUM|3|38|在帳幕前東邊，向日出的方向，安營的是 摩西 、 亞倫 和 亞倫 的兒子。他們負責看守聖所，是為 以色列 人看守的。近前來的外人必被處死。
NUM|3|39|凡被數的 利未 人，就是 摩西 、 亞倫 照耶和華所指示、按宗族所數的，一個月以上所有的男子共有二萬二千名。
NUM|3|40|耶和華對 摩西 說：「你要數點 以色列 人中凡一個月以上頭生的男子，登記他們的名字。
NUM|3|41|我是耶和華。你要揀選 利未 人歸我，代替所有頭生的 以色列 人，也取 利未 人的牲畜代替 以色列 人所有頭生的牲畜。」
NUM|3|42|摩西 就遵照耶和華所吩咐的，把所有 以色列 人頭生的都數點了。
NUM|3|43|按人名的數目，凡一個月以上頭生的男子共有二萬二千二百七十三名。
NUM|3|44|耶和華吩咐 摩西 說：
NUM|3|45|「你要揀選 利未 人代替所有頭生的 以色列 人，也要取 利未 人的牲畜代替 以色列 人的牲畜。 利未 人要歸我，我是耶和華。
NUM|3|46|以色列 人頭生的男子比 利未 人多了二百七十三名，必須把他們贖出來；
NUM|3|47|按照人丁，照聖所的舍客勒，每人當付五舍客勒，一舍客勒是二十季拉。
NUM|3|48|你要把這些多出來的人的贖銀交給 亞倫 和他的兒子。」
NUM|3|49|於是 摩西 從那被 利未 人所贖以外多出來的人取了贖銀。
NUM|3|50|從頭生的 以色列 人所取的銀子，按照聖所的舍客勒，共計一千三百六十五舍客勒。
NUM|3|51|摩西 遵照耶和華指示的話，把贖銀交給 亞倫 和他的兒子，正如耶和華所吩咐的。
NUM|4|1|耶和華吩咐 摩西 和 亞倫 說：
NUM|4|2|「你要照宗族、父家計算 利未 人中 哥轄 子孫的人口，
NUM|4|3|就是從三十歲到五十歲，凡前來任職，在會幕裏事奉的人。
NUM|4|4|這是 哥轄 子孫在會幕裏有關至聖之物的職責。
NUM|4|5|「拔營的時候， 亞倫 和他兒子要進去，把遮掩的幔子取下，用它來遮蓋法櫃，
NUM|4|6|又用精美皮料蓋在上面，鋪上純藍色的布，再把槓穿上。
NUM|4|7|他們要用藍色的布鋪在供餅的桌上，將盤、碟，以及澆酒祭的杯和壺擺在上面；經常供的餅也要留在桌上。
NUM|4|8|他們要在這些東西的上面鋪上朱紅色的布，把精美皮料蓋在上面，再把槓穿上。
NUM|4|9|他們要用藍色的布遮蓋供職用的燈臺、燈臺上的燈盞、燈剪、燈盤，以及所有盛油的器皿；
NUM|4|10|又要用精美皮料把燈臺和燈臺的一切器具包好，放在抬架上。
NUM|4|11|他們要用藍色的布鋪在金壇上，用精美皮料蓋在上面，再把槓穿上。
NUM|4|12|要用藍色的布把聖所供職用的一切器具包好，再用精美皮料蓋在上面，放在抬架上。
NUM|4|13|他們要清理祭壇上的灰，用紫色的布鋪在壇上；
NUM|4|14|又要把供職用的一切器具，就是祭壇一切的器具，火盆、肉叉、鏟子和盤子，都擺在壇上，鋪上精美皮料，再把槓穿上。
NUM|4|15|「拔營的時候， 亞倫 和他兒子把聖所和聖所一切的器具蓋好之後， 哥轄 的子孫才好來抬，免得他們摸聖物而死；這是 哥轄 子孫在會幕裏所當抬的。
NUM|4|16|「祭司 亞倫 的兒子 以利亞撒 所要照管的是點燈的油和香料，以及常獻的素祭和膏油。他要照管整個帳幕和其中所有的，以及聖所和聖所的器具。」
NUM|4|17|耶和華吩咐 摩西 和 亞倫 說：
NUM|4|18|「你們不可使 哥轄 人宗族的這一支從 利未 人中剪除。
NUM|4|19|他們挨近至聖之物的時候，要向他們這樣做，使他們存活，不致死亡； 亞倫 和他的兒子要進去，分派各人當做的，當抬的。
NUM|4|20|但是他們不可進去觀看聖所的拆卸 ，免得死亡。」
NUM|4|21|耶和華吩咐 摩西 說：
NUM|4|22|「你要照父家、宗族計算 革順 子孫的人口；
NUM|4|23|從三十歲到五十歲，凡前來任職，在會幕裏事奉的，都要數點。
NUM|4|24|這是 革順 人宗族的職責，要做的事，要抬的東西如下：
NUM|4|25|他們要抬帳幕的幔子、會幕和會幕的蓋、外層精美皮料的蓋、會幕的門簾、
NUM|4|26|帳幕和祭壇周圍院子的帷幔和門簾、繩子，以及所有需用的器具；一切與這些東西相關的事務，他們要盡職。
NUM|4|27|革順 人的子孫一切的事奉，就是所當抬的，所當做的，都要遵照 亞倫 和他兒子的指示；他們所當抬的，你們要派他們負責。
NUM|4|28|這是 革順 人子孫的宗族在會幕裏的事奉；他們要在 亞倫 祭司的兒子 以他瑪 的手下盡職。」
NUM|4|29|「至於 米拉利 的子孫，你要照宗族、父家數點他們；
NUM|4|30|從三十歲到五十歲，凡前來任職，在會幕裏事奉的，你都要數點。
NUM|4|31|這是他們在會幕裏的事奉，他們負責要抬的是帳幕的豎板、橫木、柱子和帶卯眼的座，
NUM|4|32|院子四圍的柱子和其上帶卯眼的座、橛子、繩子和一切的器具，與一切相關事奉的物件。你們要按名指定他們要抬的器具。
NUM|4|33|這是 米拉利 子孫的宗族在會幕裏的事奉，都在 亞倫 祭司的兒子 以他瑪 的手下。」
NUM|4|34|摩西 、 亞倫 和會眾的領袖按照宗族、父家數點 哥轄 人的子孫；
NUM|4|35|從三十歲到五十歲，凡前來任職，在會幕裏事奉的，
NUM|4|36|按照宗族被數的共有二千七百五十名。
NUM|4|37|這是所有在會幕裏事奉的 哥轄 人宗族中被數的，是 摩西 和 亞倫 遵照耶和華藉 摩西 所指示數點的。
NUM|4|38|革順 子孫被數的，按照宗族、父家，
NUM|4|39|從三十歲到五十歲，凡前來任職，在會幕裏事奉的，
NUM|4|40|按照宗族、父家被數的共有二千六百三十名。
NUM|4|41|這是所有在會幕裏事奉的 革順 子孫宗族中被數的，是 摩西 和 亞倫 遵照耶和華的指示所數點的。
NUM|4|42|米拉利 子孫宗族被數的，按照宗族、父家，
NUM|4|43|從三十歲到五十歲，凡前來任職，在會幕裏事奉的，
NUM|4|44|按照宗族被數的共有三千二百名。
NUM|4|45|這是 米拉利 子孫宗族中被數的，是 摩西 和 亞倫 遵照耶和華藉 摩西 所指示數點的。
NUM|4|46|摩西 、 亞倫 和 以色列 領袖按照宗族、父家數點 利未 人，
NUM|4|47|從三十歲到五十歲，凡前來任職，在會幕裏事奉，做抬物之工的，
NUM|4|48|他們被數的共有八千五百八十名。
NUM|4|49|按照耶和華藉 摩西 所指示的來分派，各人都有自己所做的事、所抬的物；他們就這樣被數點，正如耶和華所吩咐 摩西 的。
NUM|5|1|耶和華吩咐 摩西 說：
NUM|5|2|「你要吩咐 以色列 人，把一切患痲瘋 的、患漏症的和因屍體而不潔淨的，都送到營外去。
NUM|5|3|無論男女你都要送，把他們送到營外，免得他們玷污了他們的營，這是我住在他們中間的地方。」
NUM|5|4|以色列 人就照樣做，把他們送到營外去。耶和華怎樣吩咐 摩西 ， 以色列 人就照樣做了。
NUM|5|5|耶和華吩咐 摩西 說：
NUM|5|6|「你要吩咐 以色列 人：無論男女，若犯了人所常犯的任何罪 ，以致干犯耶和華，那人就有了罪。
NUM|5|7|他要承認所犯的罪，將所虧負人的如數賠償，另外再加五分之一，交給所虧負的人。
NUM|5|8|那人若沒有至親可接受所賠償的，所賠償的就要歸耶和華，交給祭司；另外還要獻一隻贖罪的公羊為他贖罪。
NUM|5|9|以色列 人一切的聖物中，所奉給祭司的一切禮物都要歸給祭司。
NUM|5|10|各人自己的聖物歸自己，給祭司的要歸給祭司。」
NUM|5|11|耶和華吩咐 摩西 說：
NUM|5|12|「你要吩咐 以色列 人，對他們說：若任何人的妻子背離婦道，對丈夫不貞，
NUM|5|13|有人與她同寢交合，這事瞞過她的丈夫，沒有被發現；她玷污自己，沒有證人指控她，也沒有被捉住；
NUM|5|14|丈夫若生了疑忌的心，對妻子起了疑忌，認為她玷污自己；或是丈夫生了疑忌的心，對妻子起了疑忌，雖然她沒有玷污自己，
NUM|5|15|這人要帶妻子到祭司那裏，同時為她帶十分之一伊法大麥麵粉作供物。不可澆上油，也不可加乳香，因為這是疑忌的素祭，是紀念的素祭，使人記得罪孽。
NUM|5|16|「祭司要使那婦人近前來，站在耶和華面前。
NUM|5|17|祭司要把聖水盛在瓦器裏，從帳幕的地上取些塵土，放在水中。
NUM|5|18|祭司要帶那婦人站在耶和華面前，使她蓬頭散髮，再把紀念的素祭，就是疑忌的素祭，放在她的手掌，祭司手裏捧著致詛咒的苦水。
NUM|5|19|祭司要叫婦人起誓，對她說：『若沒有人與你同寢，若你未曾背著丈夫做污穢的事，你就能免去這致詛咒的苦水。
NUM|5|20|但你背著丈夫，玷污自己，跟丈夫以外的人同寢。』
NUM|5|21|祭司叫婦人賭咒起誓，祭司對她說：『當耶和華使你大腿萎縮，肚腹腫脹時，願耶和華使你在你百姓中成為詛咒和咒罵；
NUM|5|22|願這致詛咒的水進入你體內，使你肚腹腫脹，大腿萎縮。』婦人要說：『阿們，阿們。』
NUM|5|23|「祭司要把這詛咒寫在冊上，然後用苦水塗去，
NUM|5|24|又叫婦人喝這致詛咒的苦水，這詛咒的水要進入她裏面，令她痛苦。
NUM|5|25|祭司要從婦人手中取那疑忌的素祭，把素祭在耶和華面前搖一搖，拿到祭壇前；
NUM|5|26|又要從素祭中取出一把，作為紀念，燒在壇上，然後叫婦人喝這水。
NUM|5|27|祭司叫她喝了以後，她若玷污自己，確實對丈夫不貞，這致詛咒的水必進入她裏面，令她痛苦，她的肚腹就要腫脹起來，大腿萎縮；這婦人就在她百姓中成為詛咒。
NUM|5|28|這婦人若沒有玷污自己，是貞潔的，就要免受這災，並且能夠生育。
NUM|5|29|「這是疑忌的條例。妻子背離丈夫玷污自己，
NUM|5|30|或是丈夫生了疑忌的心，對妻子起了疑忌，祭司要使那婦人站在耶和華面前，在她身上照這條例而行。
NUM|5|31|男人可免罪責；女人必須擔當自己的罪孽。」
NUM|6|1|耶和華吩咐 摩西 說：
NUM|6|2|「你要吩咐 以色列 人，對他們說：無論男女，若許了特別的願，就是拿細耳人的願，願意離俗歸耶和華，
NUM|6|3|他就要遠離清酒烈酒，也不可喝任何清酒烈酒做的醋；不可喝任何葡萄汁，也不可吃鮮葡萄和乾葡萄。
NUM|6|4|在一切離俗的日子，任何葡萄樹上所結的，甚至果核和果皮，都不可吃。
NUM|6|5|「在他一切許願離俗的日子，不可用剃刀剃頭。在離俗歸耶和華的日子未滿之前，他要成為聖，要任由頭上的髮綹生長。
NUM|6|6|在他一切離俗歸耶和華的日子，不可挨近死屍。
NUM|6|7|即使他的父母或兄弟姊妹死了，他也不可因他們使自己不潔淨，因為他頭上有離俗歸上帝的記號 。
NUM|6|8|在他一切離俗的日子，他是歸耶和華為聖的。
NUM|6|9|「若在他旁邊忽然有人死了，因而玷污了他離俗的頭，他要在第七日，得潔淨的日子剃頭。
NUM|6|10|第八日，他要把兩隻斑鳩或兩隻雛鴿帶到會幕門口，交給祭司。
NUM|6|11|祭司要獻一隻作贖罪祭，一隻作燔祭，為他贖因屍體而有的罪，並要在當日使他的頭分別為聖。
NUM|6|12|他要另選離俗歸耶和華的日子，牽一隻一歲的小公羊來作贖愆祭。先前的那段日子算為無效，因為他在離俗期間被玷污了。
NUM|6|13|「拿細耳人的條例是這樣的：離俗的日子滿了，祭司要領他到會幕門口，
NUM|6|14|他要將供物獻給耶和華，就是一隻沒有殘疾的一歲小公羊作燔祭，一隻沒有殘疾的一歲小母羊作贖罪祭，和一隻沒有殘疾的公綿羊作平安祭，
NUM|6|15|一籃用油調和的無酵細麵餅和抹了油的無酵薄餅，以及同獻的素祭和澆酒祭。
NUM|6|16|祭司要來到耶和華面前，獻上那人的贖罪祭和燔祭。
NUM|6|17|祭司要把公綿羊和那籃無酵餅獻給耶和華作平安祭，又要獻上同獻的素祭和澆酒祭。
NUM|6|18|拿細耳人要在會幕門口剃離俗的頭，把離俗頭上的髮放在平安祭下的火上。
NUM|6|19|他剃了離俗的頭以後，祭司要取那煮好的公綿羊的一條前腿，連同籃子裏的一塊無酵餅和一塊無酵薄餅，放在他手掌上。
NUM|6|20|祭司要拿這些在耶和華面前搖一搖，作為搖祭；這和所搖的胸、所舉的腿一樣是聖物，是歸給祭司的。然後拿細耳人才可以喝酒。
NUM|6|21|「這是拿細耳人許願的條例，除了他手頭財力所及之外，他要為離俗獻供物給耶和華。他怎樣許願，就當照離俗的條例做。」
NUM|6|22|耶和華吩咐 摩西 說：
NUM|6|23|「你要吩咐 亞倫 和他兒子說：你們要這樣為 以色列 人祝福，對他們說：
NUM|6|24|『願耶和華賜福給你，保護你。
NUM|6|25|願耶和華使他的臉光照你，賜恩給你。
NUM|6|26|願耶和華向你仰臉，賜你平安。』
NUM|6|27|「他們要如此奉我的名為 以色列 人祝福；我也要賜福給他們。」
NUM|7|1|摩西 豎立帳幕後，就用膏抹了帳幕，使它分別為聖，又用膏抹其中的一切器具，以及祭壇和壇上的一切器具，使它們分別為聖。
NUM|7|2|以色列 的領袖，各父家的家長，都前來奉獻。他們是各支派的領袖，管理那些被數的人。
NUM|7|3|他們把自己的供物送到耶和華面前，就是六輛篷車和十二頭公牛。每兩個領袖奉獻一輛車，每個領袖奉獻一頭牛。他們把這些都帶到帳幕前。
NUM|7|4|耶和華對 摩西 說：
NUM|7|5|「你要從他們收下這些，作為會幕事奉的用途，照著 利未 人所事奉的交給他們各人。」
NUM|7|6|於是 摩西 收了車和牛，交給 利未 人。
NUM|7|7|他把兩輛車和四頭牛，照著 革順 子孫所事奉的交給他們，
NUM|7|8|又把四輛車和八頭牛，照著 米拉利 子孫所事奉的交給他們。他們都在 亞倫 祭司的兒子 以他瑪 的手下。
NUM|7|9|但沒有交給 哥轄 子孫任何東西，因為他們所事奉的是聖物，必須抬在肩頭上。
NUM|7|10|用膏抹祭壇的那一天，眾領袖前來為獻壇奉獻；眾領袖都在祭壇前獻供物。
NUM|7|11|耶和華對 摩西 說：「眾領袖為獻壇奉獻供物，每天要有一個領袖前來奉獻。」
NUM|7|12|第一天獻供物的是 猶大 支派的 亞米拿達 的兒子 拿順 。
NUM|7|13|他的供物是：一個重一百三十舍客勒的銀盤，一個重七十舍客勒的銀碗，都是按照聖所的舍客勒，裏面盛滿了調油的細麵作素祭；
NUM|7|14|一個重十舍客勒的金碟子，盛滿了香；
NUM|7|15|一頭公牛犢、一隻公綿羊、一隻一歲的小公羊作燔祭；
NUM|7|16|一隻公山羊作贖罪祭；
NUM|7|17|兩頭公牛、五隻公綿羊、五隻公山羊、五隻一歲的小公羊作平安祭。這是 亞米拿達 的兒子 拿順 的供物。
NUM|7|18|第二天來獻的是 以薩迦 的領袖， 蘇押 的兒子 拿坦業 。
NUM|7|19|他獻為供物的是：一個重一百三十舍客勒的銀盤，一個重七十舍客勒的銀碗，都是按照聖所的舍客勒，裏面盛滿了調油的細麵作素祭；
NUM|7|20|一個重十舍客勒的金碟子，盛滿了香；
NUM|7|21|一頭公牛犢、一隻公綿羊、一隻一歲的小公羊作燔祭；
NUM|7|22|一隻公山羊作贖罪祭；
NUM|7|23|兩頭公牛、五隻公綿羊、五隻公山羊、五隻一歲的小公羊作平安祭。這是 蘇押 的兒子 拿坦業 的供物。
NUM|7|24|第三天是 西布倫 子孫的領袖， 希倫 的兒子 以利押 。
NUM|7|25|他的供物是：一個重一百三十舍客勒的銀盤，一個重七十舍客勒的銀碗，都是按照聖所的舍客勒，裏面盛滿了調油的細麵作素祭；
NUM|7|26|一個重十舍客勒的金碟子，盛滿了香；
NUM|7|27|一頭公牛犢、一隻公綿羊、一隻一歲的小公羊作燔祭；
NUM|7|28|一隻公山羊作贖罪祭；
NUM|7|29|兩頭公牛、五隻公綿羊、五隻公山羊、五隻一歲的小公羊作平安祭。這是 希倫 的兒子 以利押 的供物。
NUM|7|30|第四天是 呂便 子孫的領袖， 示丟珥 的兒子 以利蓿 。
NUM|7|31|他的供物是：一個重一百三十舍客勒的銀盤，一個重七十舍客勒的銀碗，都是按照聖所的舍客勒，裏面盛滿了調油的細麵作素祭；
NUM|7|32|一個重十舍客勒的金碟子，盛滿了香；
NUM|7|33|一頭公牛犢、一隻公綿羊、一隻一歲的小公羊作燔祭；
NUM|7|34|一隻公山羊作贖罪祭；
NUM|7|35|兩頭公牛、五隻公綿羊、五隻公山羊、五隻一歲的小公羊作平安祭。這是 示丟珥 的兒子 以利蓿 的供物。
NUM|7|36|第五天是 西緬 子孫的領袖， 蘇利沙代 的兒子 示路蔑 。
NUM|7|37|他的供物是：一個重一百三十舍客勒的銀盤，一個重七十舍客勒的銀碗，都是按照聖所的舍客勒，裏面盛滿了調油的細麵作素祭；
NUM|7|38|一個重十舍客勒的金碟子，盛滿了香；
NUM|7|39|一頭公牛犢、一隻公綿羊、一隻一歲的小公羊作燔祭；
NUM|7|40|一隻公山羊作贖罪祭；
NUM|7|41|兩頭公牛、五隻公綿羊、五隻公山羊、五隻一歲的小公羊作平安祭。這是 蘇利沙代 的兒子 示路蔑 的供物。
NUM|7|42|第六天是 迦得 子孫的領袖， 丟珥 的兒子 以利雅薩 。
NUM|7|43|他的供物是：一個重一百三十舍客勒的銀盤，一個重七十舍客勒的銀碗，都是按照聖所的舍客勒，裏面盛滿了調油的細麵作素祭；
NUM|7|44|一個重十舍客勒的金碟子，盛滿了香；
NUM|7|45|一頭公牛犢、一隻公綿羊、一隻一歲的小公羊作燔祭；
NUM|7|46|一隻公山羊作贖罪祭；
NUM|7|47|兩頭公牛、五隻公綿羊、五隻公山羊、五隻一歲的小公羊作平安祭。這是 丟珥 的兒子 以利雅薩 的供物。
NUM|7|48|第七天是 以法蓮 子孫的領袖， 亞米忽 的兒子 以利沙瑪 。
NUM|7|49|他的供物是：一個重一百三十舍客勒的銀盤，一個重七十舍客勒的銀碗，都是按照聖所的舍客勒，裏面盛滿了調油的細麵作素祭；
NUM|7|50|一個重十舍客勒的金碟子，盛滿了香；
NUM|7|51|一頭公牛犢、一隻公綿羊、一隻一歲的小公羊作燔祭；
NUM|7|52|一隻公山羊作贖罪祭；
NUM|7|53|兩頭公牛、五隻公綿羊、五隻公山羊、五隻一歲的小公羊作平安祭。這是 亞米忽 的兒子 以利沙瑪 的供物。
NUM|7|54|第八天是 瑪拿西 子孫的領袖， 比大蓿 的兒子 迦瑪列 。
NUM|7|55|他的供物是：一個重一百三十舍客勒的銀盤，一個重七十舍客勒的銀碗，都是按照聖所的舍客勒，裏面盛滿了調油的細麵作素祭；
NUM|7|56|一個重十舍客勒的金碟子，盛滿了香；
NUM|7|57|一頭公牛犢、一隻公綿羊、一隻一歲的小公羊作燔祭；
NUM|7|58|一隻公山羊作贖罪祭；
NUM|7|59|兩頭公牛、五隻公綿羊、五隻公山羊、五隻一歲的小公羊作平安祭。這是 比大蓿 的兒子 迦瑪列 的供物。
NUM|7|60|第九天是 便雅憫 子孫的領袖， 基多尼 的兒子 亞比但 。
NUM|7|61|他的供物是：一個重一百三十舍客勒的銀盤，一個重七十舍客勒的銀碗，都是按照聖所的舍客勒，裏面盛滿了調油的細麵作素祭；
NUM|7|62|一個重十舍客勒的金碟子，盛滿了香；
NUM|7|63|一頭公牛犢、一隻公綿羊、一隻一歲的小公羊作燔祭；
NUM|7|64|一隻公山羊作贖罪祭；
NUM|7|65|兩頭公牛、五隻公綿羊、五隻公山羊、五隻一歲的小公羊作平安祭。這是 基多尼 的兒子 亞比但 的供物。
NUM|7|66|第十天是 但 子孫的領袖， 亞米沙代 的兒子 亞希以謝 。
NUM|7|67|他的供物是：一個重一百三十舍客勒的銀盤，一個重七十舍客勒的銀碗，都是按照聖所的舍客勒，裏面盛滿了調油的細麵作素祭；
NUM|7|68|一個重十舍客勒的金碟子，盛滿了香；
NUM|7|69|一頭公牛犢、一隻公綿羊、一隻一歲的小公羊作燔祭；
NUM|7|70|一隻公山羊作贖罪祭；
NUM|7|71|兩頭公牛、五隻公綿羊、五隻公山羊、五隻一歲的小公羊作平安祭。這是 亞米沙代 的兒子 亞希以謝 的供物。
NUM|7|72|第十一天是 亞設 子孫的領袖， 俄蘭 的兒子 帕結 。
NUM|7|73|他的供物是：一個重一百三十舍客勒的銀盤，一個重七十舍客勒的銀碗，都是按照聖所的舍客勒，裏面盛滿了調油的細麵作素祭；
NUM|7|74|一個重十舍客勒的金碟子，盛滿了香；
NUM|7|75|一頭公牛犢、一隻公綿羊、一隻一歲的小公羊作燔祭；
NUM|7|76|一隻公山羊作贖罪祭；
NUM|7|77|兩頭公牛、五隻公綿羊、五隻公山羊、五隻一歲的小公羊作平安祭。這是 俄蘭 的兒子 帕結 的供物。
NUM|7|78|第十二天是 拿弗他利 子孫的領袖， 以南 兒子 亞希拉 。
NUM|7|79|他的供物是：一個重一百三十舍客勒的銀盤，一個重七十舍客勒的銀碗，都是按照聖所的舍客勒，裏面盛滿了調油的細麵作素祭；
NUM|7|80|一個重十舍客勒的金碟子，盛滿了香；
NUM|7|81|一頭公牛犢、一隻公綿羊、一隻一歲的小公羊作燔祭；
NUM|7|82|一隻公山羊作贖罪祭；
NUM|7|83|兩頭公牛、五隻公綿羊、五隻公山羊、五隻一歲的小公羊作平安祭。這是 以南 的兒子 亞希拉 的供物。
NUM|7|84|用膏抹祭壇的那一天， 以色列 的眾領袖為獻壇所獻的是：銀盤十二個、銀碗十二個、金碟子十二個；
NUM|7|85|一個銀盤重一百三十，一個碗七十。一切器皿的銀子，按照聖所的舍客勒共二千四百舍客勒。
NUM|7|86|十二個金碟子盛滿了香，按照聖所的舍客勒，一個碟子重十舍客勒，所有碟子的金子共一百二十舍客勒。
NUM|7|87|作燔祭的共有公牛十二頭、公羊十二隻、一歲的小公羊十二隻，和同獻的素祭，以及作贖罪祭的公山羊十二隻；
NUM|7|88|作平安祭的共有公牛二十四頭、公綿羊六十隻、公山羊六十隻、一歲的小公羊六十隻。這就是用膏抹壇之後，為獻壇的奉獻。
NUM|7|89|摩西 進會幕要與耶和華說話的時候，聽見法櫃的櫃蓋以上二基路伯中間有對他說話的聲音。耶和華向他說話。
NUM|8|1|耶和華吩咐 摩西 說：
NUM|8|2|「你要吩咐 亞倫 ，對他說：點燈的時候，七盞燈都要照亮燈臺前面。」
NUM|8|3|亞倫 就照樣做了；他點燈，照亮了燈臺前面，正如耶和華所吩咐 摩西 的。
NUM|8|4|燈臺是這樣造的：燈臺是用金子錘出來的，連座帶花都是錘出來的。 摩西 照著耶和華所指示的樣式造了燈臺。
NUM|8|5|耶和華吩咐 摩西 說：
NUM|8|6|「你要從 以色列 人中選出 利未 人來，潔淨他們。
NUM|8|7|你要這樣做來潔淨他們：要用潔淨的水彈在他們身上，又叫他們用剃刀剃刮全身，洗淨衣服，潔淨自己。
NUM|8|8|然後他們要取一頭公牛犢，以及同獻的素祭，就是調油的細麵。你要另取一頭公牛犢作贖罪祭。
NUM|8|9|你要帶 利未 人到會幕前，並且要召集 以色列 全會眾。
NUM|8|10|你要把 利未 人帶到耶和華面前， 以色列 人要為 利未 人按手。
NUM|8|11|亞倫 要從 以色列 人中將 利未 人奉獻 在耶和華面前，作為搖祭，使他們事奉耶和華。
NUM|8|12|利未 人要按手在那兩頭牛的頭上；你要將一頭作贖罪祭，一頭作燔祭，獻給耶和華，為 利未 人贖罪。
NUM|8|13|你也要使 利未 人站在 亞倫 和他兒子面前，將他們奉獻給耶和華，作為搖祭。
NUM|8|14|「你從 以色列 人中將 利未 人分別出來， 利未 人就歸我了。
NUM|8|15|你潔淨了 利未 人，奉獻他們作為搖祭之後，他們就可以進會幕事奉。
NUM|8|16|因為他們是從 以色列 人中全然獻給我的；我選他們歸我，代替 以色列 人中所有頭胎的長子。
NUM|8|17|因為 以色列 人中凡頭生的，無論是人或牲畜，都是我的。我在 埃及 地擊殺所有頭生的那日，已將他們分別為聖歸我。
NUM|8|18|我選 利未 人代替 以色列 人中所有頭生的。
NUM|8|19|我從 以色列 人中將 利未 人給 亞倫 和他的兒子作為賞賜，在會幕中為 以色列 人事奉，又為 以色列 人贖罪，免得 以色列 人因挨近聖所而遭受災禍。」
NUM|8|20|摩西 、 亞倫 和 以色列 全會眾就向 利未 人這樣做。關於 利未 人，凡耶和華怎樣吩咐 摩西 ， 以色列 人就向他們照樣做了。
NUM|8|21|於是 利未 人從罪中潔淨自己，洗淨衣服。 亞倫 將他們奉獻在耶和華面前，作為搖祭，又為他們贖罪，潔淨他們。
NUM|8|22|然後 利未 人進去，在 亞倫 和他兒子面前，在會幕中事奉。關於 利未 人，耶和華怎樣吩咐 摩西 ，他們就向 利未 人照樣做了。
NUM|8|23|耶和華吩咐 摩西 說：
NUM|8|24|「這是有關 利未 人的：二十五歲以上的人都要前來任職，在會幕裏事奉。
NUM|8|25|到了五十歲，他們就要從事奉的工作中退休，不再事奉，
NUM|8|26|只可在會幕裏輔助他們的弟兄盡責，他們自己不再事奉了。關於 利未 人的職責，你要向他們這樣做。」
NUM|9|1|以色列 人出 埃及 地以後，第二年正月，耶和華在 西奈 的曠野吩咐 摩西 說：
NUM|9|2|「 以色列 人應當在所定的日期守逾越節。
NUM|9|3|你們要在本月十四日黃昏的時候 ，在所定的日期守這節，按照一切的律例典章守節。」
NUM|9|4|於是 摩西 吩咐 以色列 人守逾越節。
NUM|9|5|正月十四日黃昏的時候，他們就在 西奈 的曠野守逾越節。凡耶和華所吩咐 摩西 的， 以色列 人都照樣做了。
NUM|9|6|有幾個人因屍體成了不潔淨，不能在那日守逾越節。當天他們到 摩西 、 亞倫 面前。
NUM|9|7|那些人對他說：「我們因屍體而不潔淨，為何禁止我們，不能和 以色列 人在所定的日期獻供物給耶和華呢？」
NUM|9|8|摩西 對他們說：「你們稍等，讓我去聽耶和華對你們有甚麼吩咐。」
NUM|9|9|耶和華吩咐 摩西 說：
NUM|9|10|「你要吩咐 以色列 人說：你們和你們後代中，若有人因屍體成了不潔淨，或出外遠行，仍然要向耶和華守逾越節，
NUM|9|11|他們就要在二月十四日黃昏的時候守節，要吃羔羊，以及無酵餅和苦菜。
NUM|9|12|他們不可留一點食物到早晨；羔羊的骨頭一根也不可折斷。他們要照逾越節的一切律例守這節。
NUM|9|13|但潔淨又不出外遠行的人若不守逾越節，那人要從百姓中剪除，因為他沒有在所定的日期獻供物給耶和華，必須擔當自己的罪。
NUM|9|14|若有寄居在你們那裏的外人要向耶和華守逾越節，他要照逾越節的律例和典章做。無論是寄居的或是本地人，都用同樣的律例。」
NUM|9|15|立起帳幕的那日，有雲彩遮蓋帳幕，就是法櫃的帳幕；從晚上到早晨，雲彩在帳幕上，形狀如火。
NUM|9|16|經常都是這樣：雲彩遮蓋帳幕，夜間雲彩形狀如火。
NUM|9|17|雲彩幾時從帳幕上升， 以色列 人就幾時起行；雲彩在哪裏停住， 以色列 人就在哪裏安營。
NUM|9|18|以色列 人遵照耶和華的指示起行，也遵照耶和華的指示安營。雲彩在帳幕上停留多久，他們就留在營裏多久。
NUM|9|19|雲彩在帳幕上停留許多日子， 以色列 人就遵照耶和華的吩咐不起行。
NUM|9|20|有時雲彩在帳幕上只停了幾天，他們就遵照耶和華的指示留在營裏，也遵照耶和華的指示起行。
NUM|9|21|有時雲彩從晚上留到早晨；早晨雲彩上升，他們就起行。無論是白天是黑夜，當雲彩上升的時候，他們就要起行。
NUM|9|22|雲彩停留在帳幕上，無論是兩天，一個月，或更長的日子， 以色列 人就留在營裏不起行；但雲彩一上升，他們就起行。
NUM|9|23|他們遵照耶和華的指示安營，也遵照耶和華的指示起行。他們遵守耶和華的吩咐，是耶和華藉 摩西 所指示的話。
NUM|10|1|耶和華吩咐 摩西 說：
NUM|10|2|「你要用銀子做兩枝號筒，把它們錘出來，給你用來召集會眾，拔營起行。
NUM|10|3|吹號的時候，全會眾要到你那裏，聚集在會幕的門口。
NUM|10|4|若只吹一枝，眾領袖，就是 以色列 部隊的官長，要到你那裏聚集。
NUM|10|5|你們大聲吹號的時候，東邊安營的要起行。
NUM|10|6|第二次大聲吹號的時候，南邊安營的要起行。起行的時候，要大聲吹號；
NUM|10|7|但召集會眾的時候，你們要吹號，卻不要吹出大聲。
NUM|10|8|亞倫 子孫作祭司的要吹這號筒，作為你們世世代代永遠的定例。
NUM|10|9|當你們在自己的土地上，與欺壓你們的敵人打仗時，要用號筒吹出大聲。你們就在耶和華－你們的上帝面前得蒙記念，也必蒙拯救脫離仇敵。
NUM|10|10|在快樂的日子，節期和初一，獻燔祭與平安祭的時候，你們要吹號筒，在你們的上帝面前作為紀念。我是耶和華－你們的上帝。」
NUM|10|11|第二年二月二十日，雲彩從法櫃的帳幕上升。
NUM|10|12|以色列 人離開 西奈 的曠野，一段一段地往前行，雲彩停在 巴蘭 的曠野。
NUM|10|13|他們遵照耶和華藉 摩西 所指示的，初次往前行。
NUM|10|14|按照隊伍首先起行的是 猶大 營旗幟下的人，帶隊的是 亞米拿達 的兒子 拿順 。
NUM|10|15|以薩迦 支派帶隊的是 蘇押 的兒子 拿坦業 。
NUM|10|16|西布倫 支派帶隊的是 希倫 的兒子 以利押 。
NUM|10|17|帳幕拆卸了， 革順 的子孫和 米拉利 的子孫就抬著帳幕往前行。
NUM|10|18|按照隊伍往前行的是 呂便 營旗幟下的人，帶隊的是 示丟珥 的兒子 以利蓿 。
NUM|10|19|西緬 支派帶隊的是 蘇利沙代 的兒子 示路蔑 。
NUM|10|20|迦得 支派帶隊的是 丟珥 的兒子 以利雅薩 。
NUM|10|21|哥轄 人抬著聖物往前行。他們未到以前，帳幕已經立好了。
NUM|10|22|按照隊伍往前行的是 以法蓮 營旗幟下的人，帶隊的是 亞米忽 的兒子 以利沙瑪 。
NUM|10|23|瑪拿西 支派帶隊的是 比大蓿 的兒子 迦瑪列 。
NUM|10|24|便雅憫 支派帶隊的是 基多尼 的兒子 亞比但 。
NUM|10|25|作全營後衛，按隊伍往前行的是 但 營旗幟下的人，帶隊的是 亞米沙代 的兒子 亞希以謝 。
NUM|10|26|亞設 支派帶隊的是 俄蘭 的兒子 帕結 。
NUM|10|27|拿弗他利 支派帶隊的是 以南 的兒子 亞希拉 。
NUM|10|28|以色列 人就這樣按著隊伍往前行。
NUM|10|29|摩西 對他岳父 ， 米甸 人 流珥 的兒子 何巴 說：「我們要往前行，到耶和華所說的地方；他曾說：『我要將這地賜給你們。』現在請你和我們同去，我們必善待你，因為耶和華已經應許賜福氣給 以色列 人。」
NUM|10|30|何巴 對他說：「我不去，我要回本地本族去。」
NUM|10|31|摩西 說：「請你不要離開我們，因為你知道我們要在曠野安營，你可以當我們的眼目。
NUM|10|32|你若和我們同去，將來耶和華以甚麼福氣恩待我們，我們也必這樣善待你。」
NUM|10|33|以色列 人離開耶和華的山，往前行了三天的路程。耶和華的約櫃在前面行了三天的路程，為他們尋找安歇的地方。
NUM|10|34|他們拔營往前行，日間有耶和華的雲彩在他們上面。
NUM|10|35|約櫃往前行的時候， 摩西 說： 「耶和華啊，求你興起！ 願你的仇敵潰散！ 願恨你的人從你面前逃跑！」
NUM|10|36|約櫃停住的時候，他說： 「 以色列 千萬人的耶和華啊，求你回來 ！」
NUM|11|1|百姓發怨言，惡言傳達到耶和華的耳中。耶和華聽見了就怒氣發作，耶和華的火在他們中間焚燒，燒燬營的外圍。
NUM|11|2|百姓向 摩西 哀求， 摩西 祈求耶和華，火就熄了。
NUM|11|3|那地方就叫做 他備拉 ，因為耶和華的火曾在他們中間焚燒。
NUM|11|4|他們中間的閒雜人動了貪慾的心； 以色列 人又再哭著說：「誰給我們肉吃呢？
NUM|11|5|我們記得在 埃及 的時候，不花錢就可以吃魚，還有黃瓜、西瓜、韭菜、蔥、蒜。
NUM|11|6|現在我們的精力枯乾了。除了這嗎哪以外，在我們眼前甚麼都沒有。」
NUM|11|7|嗎哪好像芫荽子，看上去如同樹脂的樣子。
NUM|11|8|百姓四處走動撿取嗎哪，把它用磨磨碎或用臼搗成粉，在鍋中煮了做成餅，滋味好像油烤餅的滋味。
NUM|11|9|夜間露水降在營中，嗎哪也隨著降下。
NUM|11|10|摩西 聽見百姓家家戶戶在帳棚門口哀哭。因此， 耶和華的怒氣大大發作， 摩西 看了也不高興。
NUM|11|11|摩西 對耶和華說：「你為何苦待僕人？我為何不在你眼前蒙恩，竟把這眾百姓的擔子加在我身上呢？
NUM|11|12|這眾百姓豈是我懷的胎，豈是我生下來的呢？你竟對我說：『把他們抱在懷裏，如養育之父抱著吃奶的嬰孩，一直抱到你起誓應許給他們祖宗的土地去。』
NUM|11|13|我從哪裏拿肉給這眾百姓吃呢？他們都向我哭著說：『給我們肉吃！』
NUM|11|14|我不能獨自帶領這眾百姓，這對我太沉重了。
NUM|11|15|如果你這樣待我，倒不如立刻把我殺了吧！我若在你眼前蒙恩，求你不要讓我再受這樣的苦。」
NUM|11|16|耶和華對 摩西 說：「你要從 以色列 的長老中為我召集七十個人，就是你所認識，作百姓的長老和官長的，領他們到會幕，使他們和你一同站在那裏。
NUM|11|17|我要在那裏降臨，與你說話，把降給你的靈分給他們。他們就和你分擔帶領百姓的擔子，免得你獨自承擔。
NUM|11|18|你要對百姓說：『你們要為了明天使自己分別為聖，你們將有肉吃。因你們哭著說：誰給我們肉吃呢？我們在 埃及 多麼好！這聲音傳到了耶和華的耳中，所以他必給你們肉吃。
NUM|11|19|你們不只吃一天、兩天、五天、十天、二十天，
NUM|11|20|而是整整一個月，直到肉從你們的鼻孔噴出來，使你們厭惡。因為你們厭棄那住在你們中間的耶和華，在他面前哭著說：我們為何出 埃及 呢？』」
NUM|11|21|摩西 說：「跟我在一起的百姓，步行的男人就有六十萬，你還說：『我要把肉賜給他們，使他們可以整整吃一個月。』
NUM|11|22|難道宰了羊群牛群，就夠給他們嗎？或者把海中所有的魚都捕來，就夠給他們嗎？」
NUM|11|23|耶和華對 摩西 說：「耶和華的膀臂 豈是縮短了嗎？現在你要看我的話向你應驗不應驗。」
NUM|11|24|摩西 出去，把耶和華的話告訴百姓，並從百姓的長老中召集七十個人來，叫他們站在會幕的四圍。
NUM|11|25|耶和華在雲中降臨，對 摩西 說話，把降給他的靈分給那七十個長老。靈停在他們身上的時候，他們就說預言，以後卻沒有再說了。
NUM|11|26|但有兩個人仍在營裏，一個名叫 伊利達 ，一個名叫 米達 。他們本是在那些登記的人中，卻沒有到會幕那裏去。靈停在他們身上，他們就在營裏說預言。
NUM|11|27|有一個年輕人跑來告訴 摩西 說：「 伊利達 和 米達 在營裏說預言。」
NUM|11|28|嫩 的兒子 約書亞 ，年輕時就作 摩西 的助手 ，說：「請我主 摩西 禁止他們。」
NUM|11|29|摩西 對他說：「你為我的緣故嫉妒嗎？惟願耶和華的百姓都是先知，願耶和華把他的靈降在他們身上！」
NUM|11|30|於是， 摩西 回到營裏去， 以色列 的長老也回去了。
NUM|11|31|有一陣風從耶和華那裏颳起，把鵪鶉從海上颳來，散落在營地和周圍；一邊約有一天的路程，另一邊也約有一天的路程，離地面約有二肘。
NUM|11|32|百姓起來，整天整夜，甚至次日一整天，都在捕捉鵪鶉。每人至少捉到十賀梅珥，各自擺在營的四圍。
NUM|11|33|但肉在他們牙間還未咀嚼時，耶和華的怒氣向百姓發作，用極重的災禍擊殺百姓。
NUM|11|34|那地方就叫 基博羅‧哈他瓦 ，因為他們在那裏埋葬了貪慾的百姓。
NUM|11|35|百姓從 基博羅‧哈他瓦 起程，到 哈洗錄 ，就住在 哈洗錄 。
NUM|12|1|摩西 娶了 古實 女子為妻。 米利暗 和 亞倫 因他娶了 古實 女子就批評他，
NUM|12|2|他們說：「難道耶和華只與 摩西 說話嗎？他不也與我們說話嗎？」耶和華聽見了。
NUM|12|3|摩西 為人極其謙和，勝過地面上的任何人。
NUM|12|4|忽然，耶和華對 摩西 、 亞倫 和 米利暗 說：「你們三個人都出來，到會幕這裏。」他們三個人就出來了。
NUM|12|5|耶和華在雲柱中降臨，停在會幕門口，叫 亞倫 和 米利暗 。二人就出來，
NUM|12|6|耶和華說：「你們要聽我的話：你們中間若有先知，我－耶和華必在異象中向他顯現，在夢中與他說話；
NUM|12|7|但我的僕人 摩西 不是這樣，他在我全家是盡忠的。
NUM|12|8|我與他面對面說話，清清楚楚，不用謎語，他甚至看見我的形像。你們為何批評我的僕人 摩西 而不懼怕呢？」
NUM|12|9|耶和華向他們怒氣發作，就離開了。
NUM|12|10|當雲彩從帳幕上離開時，看哪， 米利暗 長了痲瘋，像雪那麼白。 亞倫 轉向 米利暗 ，看哪，她長了痲瘋。
NUM|12|11|亞倫 對 摩西 說：「我主啊，求你不要因我們愚昧，因我們犯罪，就將這罪加在我們身上。
NUM|12|12|求你不要使她像那一出母腹、肉已侵蝕了一半的死胎。」
NUM|12|13|於是 摩西 哀求耶和華說：「上帝啊，求你醫治她！」
NUM|12|14|耶和華對 摩西 說：「她父親若吐唾沫在她臉上，她豈不蒙羞七天嗎？現在要把她隔離在營外七天，然後才領她回來。」
NUM|12|15|於是 米利暗 被隔離在營外七天；百姓沒有起程，直等到 米利暗 回來。
NUM|12|16|以後百姓從 哈洗錄 起行，來到 巴蘭 的曠野安營。
NUM|13|1|耶和華吩咐 摩西 說：
NUM|13|2|「你要派人去窺探我所賜給 以色列 人的 迦南 地；每個父系支派要派一個人，是他們中間的族長。」
NUM|13|3|摩西 就遵照耶和華的指示，從 巴蘭 曠野差派他們去；他們都是 以色列 人中的領袖。
NUM|13|4|這是他們的名字： 屬 呂便 支派的， 撒刻 的兒子 沙母亞 。
NUM|13|5|屬 西緬 支派的， 何利 的兒子 沙法 。
NUM|13|6|屬 猶大 支派的， 耶孚尼 的兒子 迦勒 。
NUM|13|7|屬 以薩迦 支派的， 約色 的兒子 以迦 。
NUM|13|8|屬 以法蓮 支派的， 嫩 的兒子 何西阿 。
NUM|13|9|屬 便雅憫 支派的， 拉孚 的兒子 帕提 。
NUM|13|10|屬 西布倫 支派的， 梭底 的兒子 迦疊 。
NUM|13|11|屬 約瑟 支派，就是 瑪拿西 支派的， 穌西 的兒子 迦底 。
NUM|13|12|屬 但 支派的， 基瑪利 的兒子 亞米利 。
NUM|13|13|屬 亞設 支派的， 米迦勒 的兒子 西帖 。
NUM|13|14|屬 拿弗他利 支派的， 縛西 的兒子 拿比 。
NUM|13|15|屬 迦得 支派的， 瑪基 的兒子 臼利 。
NUM|13|16|這些是 摩西 差派去窺探那地之人的名字。 摩西 叫 嫩 的兒子 何西阿 為 約書亞 。
NUM|13|17|摩西 差派他們去窺探 迦南 地，對他們說：「你們上到 尼革夫 那裏，上到山區去，
NUM|13|18|看看那地如何：住那裏的百姓是強是弱，是多是少，
NUM|13|19|他們所住的地是好是壞，所住的城鎮是營地還是堡壘，
NUM|13|20|那地是肥沃還是貧瘠，當中有樹木沒有。你們要放膽，把那地的果子帶些回來。」那時正是葡萄初熟的季節。
NUM|13|21|他們上去窺探那地，從 尋 的曠野到 利合 ，直到 哈馬口 。
NUM|13|22|他們從 尼革夫 上去，到了 希伯崙 。在那裏有 亞衲 族的 亞希幔 人、 示篩 人和 撻買 人。 希伯崙 的建造比 埃及 的 瑣安 早七年。
NUM|13|23|他們到了 以實各谷 ，從那裏砍下葡萄樹枝，上面有一掛葡萄，兩個人用槓抬著，又帶了一些石榴和無花果。
NUM|13|24|以色列 人從那裏砍下一掛葡萄，所以那地方就叫 以實各谷 。
NUM|13|25|他們窺探那地四十天之後，就回來了。
NUM|13|26|他們來到 巴蘭 曠野的 加低斯 ， 摩西 、 亞倫 ，以及 以色列 全會眾那裏，向他們和全會眾報告，又把那地的果子給他們看。
NUM|13|27|他們告訴 摩西 說：「我們到了你派我們去的那地，果然是流奶與蜜之地；這就是那地的果子。
NUM|13|28|但是住那地的百姓很強悍，城鎮又大又堅固，我們也在那裏看見了 亞衲 族人。
NUM|13|29|亞瑪力 人住在 尼革夫 ； 赫 人、 耶布斯 人和 亞摩利 人住在山區； 迦南 人住在沿海一帶和 約旦河 旁。」
NUM|13|30|迦勒 在 摩西 面前安撫百姓，說：「我們立刻上去得那地吧！我們必能征服它。」
NUM|13|31|但那些和他同去的人卻說：「我們不能上去攻打那些百姓，因為他們比我們強大。」
NUM|13|32|於是探子中有人向 以色列 人散佈有關所窺探之地的謠言，說：「我們所走過、所窺探之地是吞沒居民之地，並且我們在那裏所看見的百姓都身材高大。
NUM|13|33|我們在那裏看見巨人，就是巨人中的 亞衲 族人。我們在自己眼中像蚱蜢一樣，而在他們眼中，我們也確是這樣。」
NUM|14|1|全會眾大聲喧嚷，那夜百姓哭號。
NUM|14|2|以色列 眾人向 摩西 和 亞倫 發怨言，全會眾對他們說：「我們寧願死在 埃及 地，寧願死在這曠野！
NUM|14|3|耶和華為甚麼要把我們領到那地，讓我們倒在刀下呢？我們的妻子和孩子必成為擄物。我們回 埃及 去豈不更好嗎？」
NUM|14|4|他們彼此說：「我們不如選一個領袖，回 埃及 去吧！」
NUM|14|5|摩西 和 亞倫 在 以色列 全會眾面前臉伏於地。
NUM|14|6|窺探那地的人中， 嫩 的兒子 約書亞 和 耶孚尼 的兒子 迦勒 撕裂衣服，
NUM|14|7|對 以色列 全會眾說：「我們所走過、所窺探之地是極美之地。
NUM|14|8|耶和華若喜愛我們，就必領我們進入那地，把這流奶與蜜之地賜給我們。
NUM|14|9|但你們不可背叛耶和華，也不要怕那地的百姓，因為他們是我們的食物。保護他們的已經離開他們，耶和華卻與我們同在。不要怕他們！」
NUM|14|10|當全會眾正說著要拿石頭打死他們的時候，耶和華的榮光在會幕中向 以色列 眾人顯現。
NUM|14|11|耶和華對 摩西 說：「這百姓藐視我要到幾時呢？我在他們中間行了這一切神蹟，他們還不信我要到幾時呢？
NUM|14|12|我要用瘟疫擊殺他們，使他們不得承受那地。我要使你成為大國，比他們強大。」
NUM|14|13|摩西 對耶和華說：「 埃及 人必聽見，因你曾施展大能，領這百姓從他們中間出來。
NUM|14|14|埃及 人要告訴這地的居民，他們已經聽見你─耶和華是在這百姓中間，因為你─耶和華面對面 顯示自己，你的雲彩停在他們以上。你日間在雲柱中，夜間在火柱中，在他們的前面行。
NUM|14|15|你若把這百姓殺了，好像殺一個人那樣，那聽見你名聲的列國必說：
NUM|14|16|『耶和華因為不能把這百姓領進他向他們起誓應許之地，所以在曠野把他們殺了。』
NUM|14|17|現在求主顯出大能，照你說過的話說：
NUM|14|18|『耶和華不輕易發怒， 且有豐盛的慈愛。 他赦免罪孽和過犯， 萬不以有罪的為無罪， 必懲罰人的罪， 從父到子，直到三、四代。』
NUM|14|19|求你照你的大慈愛赦免這百姓的罪孽，好像你從 埃及 到如今饒恕這百姓一樣。」
NUM|14|20|耶和華說：「我照著你的話赦免他們。
NUM|14|21|然而，我指著我的永生與遍地充滿了耶和華的榮耀起誓：
NUM|14|22|這些人雖然都看過我的榮耀和我在 埃及 與曠野所行的神蹟，仍然這十次試探我，不聽從我的話，
NUM|14|23|他們絕不能看見我向他們祖宗所起誓應許之地；凡藐視我的，一個也不得看見。
NUM|14|24|惟獨我的僕人 迦勒 ，因他另有一個心志，專心跟從我，我要領他進入他所去過的那地；他的後裔必得那地為業。
NUM|14|25|亞瑪力 人和 迦南 人住在谷中，明天你們要轉回去，沿著 紅海 的路往曠野去。」
NUM|14|26|耶和華對 摩西 和 亞倫 說：
NUM|14|27|「這邪惡的會眾向我發怨言要到幾時呢？ 以色列 人向我發的怨言，我都聽見了。
NUM|14|28|你要告訴他們，耶和華說：『我指著我的永生起誓，我必照你們在我耳中所說的待你們。
NUM|14|29|你們的屍體必倒在這曠野中。你們中間被數點，凡二十歲以上向我發怨言的，
NUM|14|30|必不得進我所起誓應許給你們居住的那地。惟有 耶孚尼 的兒子 迦勒 和 嫩 的兒子 約書亞 才能進去。
NUM|14|31|你們的孩子，就是你們說要成為擄物的，我必領他們進去，他們就得知你們所厭棄的那地。
NUM|14|32|至於你們，你們的屍體必倒在這曠野中；
NUM|14|33|你們的兒女必在曠野遊牧四十年，擔當你們不信的罪 ，直到你們的屍體在曠野消滅為止。
NUM|14|34|按你們窺探那地的四十日，一年抵一日，你們要擔當你們的罪孽四十年，你們就知道我疏遠你們了。』
NUM|14|35|我－耶和華說過，我必這樣對待這一切聚集對抗我的邪惡會眾。他們必在這曠野中消滅，死在這裏。」
NUM|14|36|摩西 所差派去窺探那地的人回來，散佈有關那地的謠言，使全會眾向 摩西 發怨言，
NUM|14|37|這些散佈謠言的人都遭受瘟疫，死在耶和華面前。
NUM|14|38|窺探那地的人中，惟有 嫩 的兒子 約書亞 和 耶孚尼 的兒子 迦勒 得以存活。
NUM|14|39|摩西 把這些話告訴 以色列 眾人，他們都極其悲哀。
NUM|14|40|他們清晨起來，上到山頂，說：「看哪，我們要上到耶和華所說的地方；因為我們犯了罪。」
NUM|14|41|摩西 說：「你們為何要這樣違背耶和華的指示呢？這事必不能順利。
NUM|14|42|不要上去，因為耶和華不在你們中間，恐怕你們在仇敵面前被擊敗。
NUM|14|43|亞瑪力 人和 迦南 人都在你們面前，你們必倒在刀下。因為你們背離不跟從耶和華，耶和華必不與你們同在。」
NUM|14|44|他們卻擅自上到山頂。但耶和華的約櫃和 摩西 都沒有離開營地。
NUM|14|45|於是 亞瑪力 人和住在那山區的 迦南 人下來，擊敗他們，追擊他們直到 何珥瑪 。
NUM|15|1|耶和華吩咐 摩西 說：
NUM|15|2|「你要吩咐 以色列 人，對他們說：你們到了我所賜給你們居住的地，
NUM|15|3|你們要從牛群羊群中取牲畜獻給耶和華為火祭，無論是燔祭或祭物，為要還所許特別的願或甘心祭，或節期的祭，作為獻給耶和華的馨香之祭，
NUM|15|4|那獻供物的要將十分之一伊法細麵和四分之一欣油調和作素祭，獻給耶和華。
NUM|15|5|無論是燔祭或祭物，要為每隻小綿羊預備四分之一欣酒作澆酒祭。
NUM|15|6|要為每隻公綿羊預備十分之二伊法細麵，和三分之一欣油調和作素祭，
NUM|15|7|又用三分之一欣酒作澆酒祭，獻給耶和華為馨香之祭。
NUM|15|8|你預備公牛獻給耶和華作燔祭或祭物，為要還所許特別的願，或平安祭，
NUM|15|9|就要把十分之三伊法細麵和半欣油調和作素祭，和公牛一同獻上，
NUM|15|10|又用半欣酒作澆酒祭，獻給耶和華為馨香的火祭。
NUM|15|11|「獻公牛、或公綿羊、或小綿羊、或小山羊，每隻都要這樣處理；
NUM|15|12|無論你們所獻的數目多少，照著數目每隻都要這樣處理。
NUM|15|13|凡本地人將馨香的火祭獻給耶和華，都要照樣處理。
NUM|15|14|若有外人寄居在你們那裏，或有人世世代代住在你們中間，願意將馨香的火祭獻給耶和華，你們怎樣處理，他也要照樣處理。
NUM|15|15|至於會眾，無論是你們或寄居的外人都要遵守同一條例；這是你們世世代代永遠的定例。在耶和華面前，你們怎樣，寄居的也要怎樣。
NUM|15|16|你們和寄居在你們那裏的外人要遵守同一律法，同一典章。」
NUM|15|17|耶和華吩咐 摩西 說：
NUM|15|18|「你要吩咐 以色列 人，對他們說：你們到了我領你們進去的那地，
NUM|15|19|吃那地的糧食時，要把舉祭獻給耶和華。
NUM|15|20|你們要用初熟的麥子磨麵，做成餅當舉祭獻上。你們要舉上，如同舉禾場的舉祭。
NUM|15|21|你們世世代代要用初熟的麥子磨麵，當舉祭獻給耶和華。
NUM|15|22|「你們若犯了錯，不遵守耶和華所吩咐 摩西 的這一切命令，
NUM|15|23|就是耶和華藉 摩西 一切所命令你們的，從耶和華命令的那日直到你們的世世代代，
NUM|15|24|會眾因沒有察覺而犯了無心之過，全會眾就要將一頭公牛犢作燔祭，遵照典章把素祭和澆酒祭一同獻給耶和華為馨香的祭，又要獻一隻公山羊作贖罪祭。
NUM|15|25|祭司要為 以色列 全會眾贖罪，他們就必蒙赦免，因為這是無心之過。他們要因自己的無心之過，把供物，就是向耶和華當獻的火祭和贖罪祭，帶到耶和華面前。
NUM|15|26|以色列 全會眾和寄居在他們中間的外人就必蒙赦免，因為這是眾百姓的無心之過。
NUM|15|27|「若有一個人無意中犯了罪，他就要獻一隻一歲的母山羊作贖罪祭。
NUM|15|28|這誤犯罪的人因無意中犯了罪，祭司要在耶和華面前為他贖罪，他就必蒙赦免。
NUM|15|29|以色列 中的本地人和寄居在他們中間的外人，若無意中犯了罪，都要遵守同一律法。
NUM|15|30|但那故意犯罪的人，無論是本地人是寄居的，褻瀆了耶和華，這人必從百姓中剪除。
NUM|15|31|因為他藐視耶和華的話，違背耶和華的命令，這人一定要剪除；他的罪孽要歸到自己身上。」
NUM|15|32|以色列 人還在曠野的時候，發現有一個人在安息日撿柴。
NUM|15|33|發現他撿柴的人把他帶到 摩西 、 亞倫 以及全會眾那裏。
NUM|15|34|他們把他收押在監裏，因為還不知道要怎樣懲罰他。
NUM|15|35|耶和華吩咐 摩西 說：「這人應當處死；全會眾要在營外用石頭打死他。」
NUM|15|36|於是全會眾把他帶到營外，用石頭打死他，是照耶和華所吩咐 摩西 的。
NUM|15|37|耶和華對 摩西 說：
NUM|15|38|「你吩咐 以色列 人，對他們說，他們世世代代要在衣服邊上縫繸子，並在邊上的繸子釘一條藍色帶子。
NUM|15|39|你們要佩帶這繸子，好叫你們看見它就記起耶和華一切的命令，並且遵行，不隨從自己內心和眼目的情慾而跟著行淫。
NUM|15|40|這樣，你們就必記得並遵行我一切的命令，成為聖，歸你們的上帝。
NUM|15|41|「我是耶和華－你們的上帝，曾把你們從 埃及 地領出來，要作你們的上帝。我是耶和華－你們的上帝。」
NUM|16|1|利未 的曾孫， 哥轄 的孫子， 以斯哈 的兒子 可拉 ，連同 呂便 子孫中 以利押 的兒子 大坍 和 亞比蘭 ，與 比勒 的兒子 安 ，帶了
NUM|16|2|以色列 人中的二百五十個領袖，就是有名望、從會眾中選出來的人，在 摩西 面前一同起來，
NUM|16|3|聚集攻擊 摩西 、 亞倫 ，說：「你們太過分了！全會眾人人都成為聖，耶和華也在他們中間。你們為甚麼抬高自己，在耶和華的會眾之上呢？」
NUM|16|4|摩西 聽見就臉伏於地，
NUM|16|5|對 可拉 和他所有同夥的人說：「到了早晨，耶和華必指示誰是屬他的，誰是成為聖的，就准許誰親近他。他要叫自己所揀選的人親近他。
NUM|16|6|可拉 和你所有同夥的人哪，你們要這樣做：要拿著香爐，
NUM|16|7|明天在耶和華面前把火盛在爐中，把香放在上面。耶和華揀選誰，誰就成為聖。 利未 的子孫哪，你們太過分了！」
NUM|16|8|摩西 又對 可拉 說：「 利未 的子孫，聽吧！
NUM|16|9|以色列 的上帝將你們從 以色列 會眾中分別出來，使你們親近他，在耶和華的帳幕中事奉，並且站在會眾面前替他們供職。這對你們豈是小事嗎？
NUM|16|10|耶和華已經准許你和你所有的弟兄，就是 利未 的子孫，一同親近他，你們還要求祭司的職分嗎？
NUM|16|11|所以，你和你所有同夥的人聚集是在攻擊耶和華。 亞倫 算甚麼，你們竟向他發怨言？」
NUM|16|12|摩西 派人去叫 以利押 的兒子 大坍 和 亞比蘭 。他們卻說：「我們不上去！
NUM|16|13|你把我們從流奶與蜜之地領出來，讓我們死在曠野，這豈是小事？你還要自立為王管轄我們嗎？
NUM|16|14|你根本沒有領我們到流奶與蜜之地，也沒有給我們田地和葡萄園作為產業。難道你想要挖這些人的眼睛嗎？我們不上去！」
NUM|16|15|摩西 非常生氣，就對耶和華說：「求你不要接受他們的供物。我並沒有奪過他們一匹驢，也沒有害過他們中任何一個人。」
NUM|16|16|摩西 對 可拉 說：「明天，你和你所有同夥的人，以及 亞倫 ，都要站在耶和華面前。
NUM|16|17|你們各人要拿一個香爐，把香放在上面，各人帶香爐到耶和華面前，共二百五十個；你和 亞倫 也各拿自己的香爐。」
NUM|16|18|於是他們各人拿一個香爐，盛著火，加上香，和 摩西 、 亞倫 一同站在會幕的門口。
NUM|16|19|可拉 召集全會眾到會幕門口攻擊 摩西 和 亞倫 。這時，耶和華的榮光向全會眾顯現。
NUM|16|20|耶和華吩咐 摩西 和 亞倫 說：
NUM|16|21|「你們離開這會眾，我好立刻把他們滅絕。」
NUM|16|22|摩西 、 亞倫 臉伏於地，說：「上帝，賜萬人氣息的上帝啊，一人犯罪，你就要向全會眾發怒嗎？」
NUM|16|23|耶和華吩咐 摩西 說：
NUM|16|24|「你吩咐會眾說：『你們遠離 可拉 、 大坍 和 亞比蘭 帳棚的周圍。』」
NUM|16|25|摩西 起來，到 大坍 、 亞比蘭 那裏去； 以色列 的長老也都跟著他去。
NUM|16|26|他吩咐會眾說：「你們離開這些惡人的帳棚吧！不可碰他們的任何東西，免得你們因他們一切的罪而消滅。」
NUM|16|27|於是會眾遠離了 可拉 、 大坍 和 亞比蘭 的帳棚。 大坍 和 亞比蘭 帶著妻子、兒女和小孩子出來，站在自己的帳棚門口。
NUM|16|28|摩西 說：「因這件事，你們就必知道這一切事是耶和華差派我做的，並非出於我的心意。
NUM|16|29|這些人的死若和世人無異，或者他們所遭遇的和其他人相同，那麼耶和華就不曾差派我了。
NUM|16|30|但是，倘若耶和華創作一件新事，使地開了裂口，把他們和一切屬他們的都吞下去，叫他們活活墜落陰間，你們就知道是這些人藐視了耶和華。」
NUM|16|31|摩西 剛說完這些話，他們腳下的地就裂開，
NUM|16|32|地開了裂口，把他們和他們的家眷，以及一切屬 可拉 的人和財物，都吞了下去。
NUM|16|33|他們和一切屬他們的，都活活墜落陰間；地在他們上面又合攏起來，他們就從會眾中滅亡了。
NUM|16|34|在他們四圍的 以色列 眾人聽見他們的叫聲，就都逃跑，說：「恐怕地也要把我們吞下去了！」
NUM|16|35|有火從耶和華那裏出來，吞滅了那上香的二百五十人。
NUM|16|36|耶和華吩咐 摩西 說：
NUM|16|37|「你要對 亞倫 祭司的兒子 以利亞撒 說，把香爐從火中移開，再把炭火撒在別處，因為這些香爐是分別為聖的。
NUM|16|38|要把那些犯罪自喪己命之人的香爐錘成薄片，用以包祭壇；因為這些本是他們在耶和華面前獻過，分別為聖的，可以給 以色列 人作記號。」
NUM|16|39|於是 以利亞撒 祭司把被燒死的人所獻的銅香爐拿來；它們被錘出來，用以包壇，
NUM|16|40|給 以色列 人作紀念，為要叫 亞倫 子孫之外的人不得近前來，在耶和華面前燒香，免得他和 可拉 與同他一夥的人一樣，正如耶和華藉 摩西 所吩咐的。
NUM|16|41|第二天， 以色列 全會眾都向 摩西 、 亞倫 發怨言說：「你們殺了耶和華的百姓了。」
NUM|16|42|會眾聚集攻擊 摩西 、 亞倫 的時候， 摩西 和 亞倫 轉向會幕，看哪，雲彩遮蓋會幕，耶和華的榮光顯現。
NUM|16|43|摩西 、 亞倫 就來到會幕前。
NUM|16|44|耶和華吩咐 摩西 說：
NUM|16|45|「你們離開這會眾，我好立刻把他們滅絕。」他們二人就臉伏於地。
NUM|16|46|摩西 對 亞倫 說：「拿你的香爐，把祭壇的火盛在裏面，加上香，趕快帶到會眾那裏，為他們贖罪。因為有憤怒從耶和華面前發出，瘟疫已經開始了。」
NUM|16|47|亞倫 照 摩西 所說的拿了香爐，跑到會眾中。看哪，瘟疫已經在百姓中開始了。他就加上香，為百姓贖罪。
NUM|16|48|他站在活人和死人之間，瘟疫就止住了。
NUM|16|49|除了因 可拉 事件死的以外，遭瘟疫死的共有一萬四千七百人。
NUM|16|50|亞倫 回到會幕門口 ，到 摩西 那裏，瘟疫已經止住了。
NUM|17|1|耶和華吩咐 摩西 說：
NUM|17|2|「你要吩咐 以色列 人，從他們當中取杖，每父家一根；從他們所有的領袖，按著父家，共取十二根。你要把各人的名字寫在他的杖上，
NUM|17|3|並要把 亞倫 的名字寫在 利未 的杖上，因為各父家的家長都有一根杖。
NUM|17|4|你要把這些杖放在會幕裏法櫃前，我與你們 相會的地方。
NUM|17|5|我所揀選的人，他的杖必發芽。我就平息了 以色列 人向你們所發的怨言，不再達到我這裏。」
NUM|17|6|於是， 摩西 吩咐 以色列 人，他們的眾領袖就把杖給他，一個領袖一根杖，按照父家一個領袖一根杖，共有十二根； 亞倫 的杖也在其中。
NUM|17|7|摩西 把這些杖放在耶和華面前，在法櫃的帳幕裏。
NUM|17|8|第二天， 摩西 進到法櫃的帳幕去，看哪， 利未 族 亞倫 的杖已經發芽，長了花苞，開了花，也結出熟的杏子！
NUM|17|9|摩西 把所有的杖從耶和華面前拿出來，給 以色列 眾人看。他們都看見了，各領袖就把自己的杖拿去。
NUM|17|10|耶和華吩咐 摩西 說：「把 亞倫 的杖放回法櫃前，給這些背叛之子留作記號。你就可以平息他們向我所發的怨言，他們也不會死亡。」
NUM|17|11|摩西 就照樣做了；耶和華怎樣吩咐他，他就照樣做。
NUM|17|12|以色列 人對 摩西 說：「看哪，我們死啦！我們滅亡啦！我們全都滅亡啦！
NUM|17|13|凡挨近耶和華帳幕的，就必死亡。我們都要消滅而死嗎？」
NUM|18|1|耶和華對 亞倫 說：「你和你的兒子，以及你父家的人，要一同擔當干犯聖所的罪孽；你和你的兒子也要擔當干犯祭司職分的罪孽。
NUM|18|2|你也要帶你弟兄 利未 人，就是你父系支派的人前來，與你聯合，服事你。你和你的兒子要一起在法櫃的帳幕前；
NUM|18|3|他們要遵守你的吩咐，負責看守整個帳幕，只是不可挨近聖所的器具和祭壇，免得他們和你們都死亡。
NUM|18|4|他們要與你聯合，負責看守會幕和帳幕一切的事；只是外人不可挨近你們。
NUM|18|5|你們要負責看守聖所和祭壇，免得憤怒再臨到 以色列 人。
NUM|18|6|看哪，我已從 以色列 人中選了你們的弟兄 利未 人，交給你們為賞賜，歸給耶和華，為要在會幕裏事奉。
NUM|18|7|你和你的兒子要謹守祭司的職分，負責一切關於祭壇和幔子內的事。我把祭司的職分賜給你們，作為賞賜好事奉我；凡挨近的外人必被處死。」
NUM|18|8|耶和華吩咐 亞倫 說：「看哪，我已將歸我的舉祭，就是 以色列 人一切分別為聖之物，交給你照管；我把受膏的份賜給你和你的子孫，作為永遠當得的份。
NUM|18|9|這是至聖供物中所給你的，一切獻給我為至聖的素祭、贖罪祭、贖愆祭，其中所有不被火燒的供物，都要歸你和你的子孫。
NUM|18|10|你要把它當作至聖之物吃 ；凡男丁都可以吃。你要以這祭物為聖。
NUM|18|11|這也是你的， 以色列 人所獻的舉祭和搖祭，我已賜給你和你的兒女，作為永遠當得的份；你家中任何潔淨的人都可以吃。
NUM|18|12|凡最好的新油、最好的新酒和五穀，就是 以色列 人獻給耶和華的初熟之物，我都賜給你。
NUM|18|13|凡他們從地上所帶來給耶和華的初熟之物也都要歸給你。你家中任何潔淨的人都可以吃。
NUM|18|14|以色列 中一切永獻的都必歸給你。
NUM|18|15|他們所有奉給耶和華的，無論是人是牲畜，凡頭胎的，都要歸給你；但是人的長子，一定要贖出來。不潔淨牲畜中頭生的，也要贖出來。
NUM|18|16|其中一個月以上所當贖的，要照你的估價，按聖所的舍客勒，付五舍客勒銀子將他贖回，一舍客勒是二十季拉。
NUM|18|17|但是頭生的牛，或頭生的綿羊，或頭生的山羊，卻不可贖，因為牠們都是聖的。要把牠們的血灑在祭壇上，把牠們的脂肪焚燒，當作馨香的火祭獻給耶和華。
NUM|18|18|牠們的肉必歸你，像被搖的胸、被舉的右腿歸你一樣。
NUM|18|19|凡 以色列 人所獻給耶和華聖物中的舉祭，我都賜給你和你的兒女，作為永遠當得的份。這要成為你和你的後裔在耶和華面前永遠的鹽 約。
NUM|18|20|耶和華對 亞倫 說：「你在 以色列 人的境內不可有產業，在他們中間也不可有份。在 以色列 人中，我是你的份，你的產業。
NUM|18|21|「至於 利未 的子孫，看哪，我已賜給他們 以色列 所有出產的十分之一為業，作為他們在會幕中事奉的酬勞。
NUM|18|22|以色列 人不可再挨近會幕，免得他們擔當罪而死。
NUM|18|23|惟獨 利未 人要在會幕中事奉，他們要擔當罪孽，作為你們世世代代永遠的定例。他們在 以色列 人中不可有產業；
NUM|18|24|因為 以色列 人出產的十分之一，就是獻給耶和華為舉祭的，我已賜給 利未 人為業。所以我對他們說，他們不可在 以色列 人中有產業。」
NUM|18|25|耶和華吩咐 摩西 說：
NUM|18|26|「你要吩咐 利未 人，對他們說：你們從 以色列 人中所取的十分之一，就是我給你們為業的，要從這十分之一中取十分之一，作為獻給耶和華的舉祭。
NUM|18|27|這可算為你們的舉祭，如同禾場上的穀，酒池中盛滿的酒。
NUM|18|28|這樣，從 以色列 人中所收取所有的十分之一，你們要從其中取舉祭獻給耶和華；你們要把獻給耶和華的舉祭歸給 亞倫 祭司。
NUM|18|29|你們要將給你們一切禮物中最好的，就是分別為聖的，獻給耶和華為舉祭。
NUM|18|30|你要對 利未 人說：當你們把其中最好的獻上為舉祭之後，這剩下的就算是你們禾場上的農作物，酒池中的酒。
NUM|18|31|你們和你們的家人可以在任何地方吃；這本是你們的賞賜，是你們在會幕裏事奉的酬勞。
NUM|18|32|當你們把其中最好的獻上為舉祭，就不致於因它擔當罪。你們不可玷污 以色列 人的聖物，免得死亡。」
NUM|19|1|耶和華吩咐 摩西 和 亞倫 說：
NUM|19|2|「耶和華所吩咐的律法中，其中一條律例這樣說：要吩咐 以色列 人，把一頭健康、沒有殘疾、未曾負軛的紅母牛牽到你這裏來，
NUM|19|3|交給 以利亞撒 祭司。他要把牛牽到營外，人就在他面前把牛宰了。
NUM|19|4|以利亞撒 祭司要用指頭蘸這牛的血，向會幕前面彈七次。
NUM|19|5|人要在他眼前焚燒這母牛，牛的皮、肉、血和糞都要焚燒。
NUM|19|6|祭司要把香柏木、牛膝草和朱紅色紗都丟在焚燒牛的火中。
NUM|19|7|祭司要洗衣服，用水洗身，然後才可以進營；祭司必不潔淨到晚上。
NUM|19|8|焚燒牛的人也要用水洗衣服，用水洗身，必不潔淨到晚上。
NUM|19|9|一個潔淨的人要收母牛的灰，存放在營外潔淨的地方，為 以色列 會眾留作除污穢的水之用。這是為除罪用的。
NUM|19|10|收取母牛灰的人要洗衣服，必不潔淨到晚上。這要成為 以色列 人和寄居在他們中間的外人永遠的定例。
NUM|19|11|「摸了任何人死屍的，必不潔淨七天。
NUM|19|12|那人要在第三天和第七天潔淨自己，他就潔淨了。若他不在第三天和第七天潔淨自己，他就不潔淨了。
NUM|19|13|凡摸了死屍，就是死了的人的屍體，又不潔淨自己的，就玷污了耶和華的帳幕，這人必從 以色列 中剪除；因為那除污穢的水沒有灑在他身上，他就不潔淨，污穢還在他身上。
NUM|19|14|「若有人死在帳棚裏，條例是這樣：凡進那帳棚的，和所有在帳棚裏的人，都必不潔淨七天。
NUM|19|15|凡敞開的，沒有用繩子紮好蓋子的器皿，也不潔淨。
NUM|19|16|任何人在田野裏摸了被刀殺的，或自然死的，或人的骨頭，或墳墓，就必不潔淨七天。
NUM|19|17|要為這不潔淨的人拿一些燒好的除罪灰放在器皿裏，倒上清水。
NUM|19|18|一個潔淨的人要拿牛膝草蘸在這水中，把水彈在帳棚上，和一切器皿以及帳棚內的人身上，又要彈在那摸了骨頭，或摸了被殺的或自然死的，或摸了墳墓的人身上。
NUM|19|19|那潔淨的人要在第三天和第七天把水彈在不潔淨的人身上，在第七天潔淨那人。那人要洗衣服，用水洗澡，到晚上就潔淨了。
NUM|19|20|但任何不潔淨的人，他若不潔淨自己，那人要從會中剪除，因為他玷污了耶和華的聖所，除污穢的水沒有灑在他身上，他是不潔淨的。
NUM|19|21|這要成為你們永遠的定例。此外，那彈除污穢水的人也要洗衣服。凡碰除污穢水的，必不潔淨到晚上。
NUM|19|22|不潔淨的人所摸的任何東西都不潔淨；摸了這東西的人必不潔淨到晚上。」
NUM|20|1|正月間， 以色列 全會眾到了 尋 的曠野；百姓住在 加低斯 。 米利暗 死在那裏，也葬在那裏。
NUM|20|2|會眾沒有水，就聚集反對 摩西 和 亞倫 。
NUM|20|3|百姓與 摩西 爭鬧，說：「我們恨不得與我們的弟兄一同死在耶和華面前。
NUM|20|4|你們為甚麼領耶和華的會眾到這曠野，使我們和我們的牲畜都死在這裏呢？
NUM|20|5|你們為甚麼領我們從 埃及 上來，把我們帶到這壞的地方呢？這地方不能撒種，沒有無花果樹、葡萄樹、石榴樹，也沒有水喝。」
NUM|20|6|摩西 、 亞倫 離開會眾面前，到會幕的門口，臉伏於地；耶和華的榮光向他們顯現。
NUM|20|7|耶和華吩咐 摩西 說：
NUM|20|8|「你拿著杖去，和你的哥哥 亞倫 召集會眾，在他們眼前吩咐磐石湧出水來，水就會從磐石流出，給會眾和他們的牲畜喝。」
NUM|20|9|於是 摩西 遵照耶和華所吩咐他的，從耶和華面前拿了杖去。
NUM|20|10|摩西 和 亞倫 召集會眾到磐石前。 摩西 對他們說：「聽著，你們這些悖逆的人！我們要叫這磐石流出水來給你們嗎？」
NUM|20|11|摩西 舉起手來，用杖擊打磐石兩下，就有許多水流出來，會眾和他們的牲畜都喝了。
NUM|20|12|但是耶和華對 摩西 、 亞倫 說：「因為你們不信我，沒有在 以色列 人眼前尊我為聖，所以你們必不能領這會眾進入我所要賜給他們的地去。」
NUM|20|13|這就是 米利巴 水，因 以色列 人與耶和華爭鬧，耶和華在他們面前顯為聖。
NUM|20|14|摩西 從 加低斯 差遣使者到 以東 王那裏，說：「你的弟兄 以色列 這樣說：『你知道我們所遭遇的一切困難。
NUM|20|15|我們的祖先曾下到 埃及 ，我們也在 埃及 住了很多年。然而， 埃及 人卻惡待我們和我們的祖先。
NUM|20|16|我們哀求耶和華，他垂聽了我們的聲音，差遣使者把我們從 埃及 領出來。看哪，我們到了你邊界的 加低斯城 。
NUM|20|17|求你讓我們穿越你的地。我們不走田間和葡萄園，也不喝井裏的水。我們只走王的大路，不偏左右，直到過了你的邊界。』」
NUM|20|18|但是， 以東 對他說：「你不可從我這裏穿越！否則，我要帶刀出去攻擊你。」
NUM|20|19|以色列 人對他說：「我們只上大道。如果我和我的牲畜喝了你的水，我必付錢給你。我不求別的事，只求讓我步行過去。」
NUM|20|20|以東 說：「你不可經過！」他就率領一大群軍隊，以強硬的手出來攻擊 以色列 。
NUM|20|21|這樣， 以東 不肯讓 以色列 穿越他的境內， 以色列 就轉去，離開他了。
NUM|20|22|以色列 全會眾從 加低斯 起行，到了 何珥山 。
NUM|20|23|耶和華在 以東 地邊界的 何珥山 對 摩西 、 亞倫 說：
NUM|20|24|「 亞倫 要歸到他祖先 那裏。他必不得進入我所賜給 以色列 人的地，因為你們在 米利巴 水的事上違背了我的指示。
NUM|20|25|你要帶 亞倫 和他的兒子 以利亞撒 上 何珥山 ，
NUM|20|26|把 亞倫 的聖衣脫下，給他的兒子 以利亞撒 穿上。 亞倫 必歸去，死在那裏。」
NUM|20|27|摩西 就遵照耶和華的吩咐去做，他們在全會眾的眼前上了 何珥山 。
NUM|20|28|摩西 把 亞倫 的聖衣脫下，給他的兒子 以利亞撒 穿上， 亞倫 就死在山頂那裏。於是， 摩西 和 以利亞撒 下了山。
NUM|20|29|全會眾見 亞倫 死了， 以色列 全家就為 亞倫 舉哀三十天。
NUM|21|1|住 尼革夫 的 迦南 人的 亞拉得 王，聽說 以色列 從 亞他林 路來，就和 以色列 交戰，擄去他們一些人。
NUM|21|2|以色列 向耶和華許願說：「你若把這百姓真的交在我手中，我就把他們的城鎮徹底毀滅。」
NUM|21|3|耶和華垂聽了 以色列 的聲音，把 迦南 人交出來。 以色列 就把 迦南 人和他們的城鎮徹底毀滅。因此，那地方名叫 何珥瑪 。
NUM|21|4|他們從 何珥山 起行，繞過 以東 地往 紅海 那條路走。在路上，百姓心中煩躁。
NUM|21|5|百姓向上帝和 摩西 發怨言，說：「你們為甚麼把我們從 埃及 領上來 ，使我們死在曠野呢？這裏沒有糧食，沒有水，我們厭惡這淡而無味的食物。」
NUM|21|6|耶和華派火蛇進入百姓當中去咬他們，於是 以色列 中死了許多百姓。
NUM|21|7|百姓到 摩西 那裏，說：「我們有罪了，因為我們向耶和華和你發怨言。求你向耶和華禱告，叫蛇離開我們。」於是 摩西 為百姓禱告。
NUM|21|8|耶和華對 摩西 說：「你要造一條火蛇，掛在杆子上。凡被咬的，一望這蛇就必存活。」
NUM|21|9|摩西 就造了一條銅蛇，掛在杆子上。凡被蛇咬的，一望這銅蛇就活了。
NUM|21|10|以色列 人起行，安營在 阿伯 。
NUM|21|11|又從 阿伯 起行，安營在 以耶‧亞巴琳 ，在 摩押 對面的曠野，向日出的方向。
NUM|21|12|又從那裏起行，安營在 撒烈谷 。
NUM|21|13|從那裏再起行，安營在 亞嫩河 的另一邊。這 亞嫩河 在曠野，從 亞摩利 人的境內流出來； 亞嫩河 是 摩押 的邊界，在 摩押 和 亞摩利 人之間。
NUM|21|14|所以《耶和華的戰記》中提到： 「 蘇法 的 哇哈伯 ， 亞嫩河 谷，
NUM|21|15|以及 亞珥 地區眾河床的斜坡， 都靠近 摩押 的邊境。」
NUM|21|16|以色列 人從那裏起行，到了 比珥 。從前耶和華對 摩西 說：「召集百姓，我要給他們水」，說的就是這井。
NUM|21|17|當時， 以色列 人唱這首歌： 「井啊，湧出水來！ 你們要向它歌唱！
NUM|21|18|這井是領袖用權杖所挖， 是百姓中的貴族用手杖所掘。」 以色列 人從曠野往 瑪他拿 去，
NUM|21|19|從 瑪他拿 到 拿哈列 ，從 拿哈列 到 巴末 ，
NUM|21|20|從 巴末 到 摩押 地的谷，又到那可以瞭望曠野的 毗斯迦山 頂。
NUM|21|21|以色列 差遣使者到 亞摩利 人的王 西宏 那裏，說：
NUM|21|22|「求你讓我們穿越你的地；我們不岔進田間和葡萄園，也不喝井裏的水，只走王的大道，直到過了你的邊界。」
NUM|21|23|但 西宏 不讓 以色列 人穿越他的境內，就召集他的眾百姓出到曠野，要攻擊 以色列 ，到了 雅雜 與 以色列 交戰。
NUM|21|24|以色列 人用刀殺了他，佔領了他的地，從 亞嫩河 到 雅博河 ，直到 亞捫 人的邊界，因為 亞捫 人的邊防堅固。
NUM|21|25|以色列 人奪取這裏所有的城鎮，就住在 亞摩利 人的城鎮中，包括 希實本 和所屬的一切鄉鎮 。
NUM|21|26|希實本 是 亞摩利 王 西宏 的首都； 西宏 曾與先前的 摩押 王交戰，從他手中奪取了他所有的地，直到 亞嫩河 。
NUM|21|27|所以那些作詩歌的說： 你們到 希實本 來吧； 願 西宏 的城被修造建立。
NUM|21|28|因為有火從 希實本 發出， 有火焰從 西宏 的城冒出， 燒燬了 摩押 的 亞珥 ， 亞嫩河 丘壇的主 。
NUM|21|29|摩押 啊，你有禍了！ 基抹 的百姓啊，你們滅亡了！ 基抹 的男子逃亡， 女子被擄， 交給了 亞摩利 王 西宏 。
NUM|21|30|我們射了他們； 希實本 直到 底本 盡都毀滅 。 我們劫掠，直到 挪法 ； 這 挪法 直延到 米底巴 。
NUM|21|31|這樣， 以色列 人就住在 亞摩利 人的地。
NUM|21|32|摩西 差派人去窺探 雅謝 ； 以色列 人佔領了 雅謝 附近的鄉村，趕出那裏的 亞摩利 人。
NUM|21|33|後來， 以色列 人轉回，往上 巴珊 的路去。 巴珊 王 噩 率領他的眾百姓出來，在 以得來 與他們交戰。
NUM|21|34|耶和華對 摩西 說：「不要怕他！因為我已將他和他的眾百姓，以及他的地都交在你手中。你要待他如同待住在 希實本 的 亞摩利 王 西宏 一樣。」
NUM|21|35|於是他們殺了 巴珊 王和他的眾子，以及他的眾百姓，沒有留下一個倖存者，並且佔領了他的地。
NUM|22|1|以色列 人起行，在 摩押 平原， 約旦河 東，對著 耶利哥 安營。
NUM|22|2|西撥 的兒子 巴勒 看見 以色列 向 亞摩利 人所做的一切。
NUM|22|3|摩押 因 以色列 百姓這麼多，非常懼怕。 摩押 因 以色列 人的緣故就憂懼。
NUM|22|4|摩押 對 米甸 的長老說：「現在這群人要舔盡我們四圍的一切，好像牛舔盡田間的草一樣。」 那時， 西撥 的兒子 巴勒 作 摩押 王。
NUM|22|5|他派使者往 大河 附近的 毗奪 去，到 比珥 的兒子 巴蘭 的家鄉 ，召 巴蘭 來，說：「看哪，有一群百姓從 埃及 出來；看哪，他們遮滿地面，住在我的對面。
NUM|22|6|現在請你來，為我詛咒這百姓，因為他們比我強大，或許我能打敗他們，把他們趕出此地。因為我知道，你為誰祝福，誰就得福；你詛咒誰，誰就受詛咒。」
NUM|22|7|摩押 的長老和 米甸 的長老手裏拿著占卜的禮金到 巴蘭 那裏，將 巴勒 的話告訴他。
NUM|22|8|巴蘭 對他們說：「今晚你們在這裏過夜，我必照著耶和華向我說的話給你們答覆。」 摩押 的官員就在 巴蘭 那裏住下。
NUM|22|9|上帝臨到 巴蘭 那裏，說：「你這裏的這些人是誰？」
NUM|22|10|巴蘭 對上帝說：「 摩押 王 西撥 的兒子 巴勒 送信給我：
NUM|22|11|『看哪，從 埃及 出來的百姓遮滿了地面，現在請你來，為我詛咒他們，或許我能打敗他們，把他們趕走。』」
NUM|22|12|上帝對 巴蘭 說：「你不可跟他們去，也不可詛咒這百姓，因為他們是蒙福的。」
NUM|22|13|巴蘭 早晨起來，對 巴勒 的官員說：「你們回本地去吧，因為耶和華不允許我和你們一起去。」
NUM|22|14|摩押 的官員就起來，到 巴勒 那裏，說：「 巴蘭 不肯和我們一起來。」
NUM|22|15|巴勒 又差遣比這些更多，更尊貴的官員。
NUM|22|16|他們來到 巴蘭 那裏，對他說：「 西撥 的兒子 巴勒 這樣說：『請你不要再推辭到我這裏來！
NUM|22|17|我必使你得極大的尊榮，無論你向我要甚麼，我都給你。只求你來為我詛咒這百姓。』」
NUM|22|18|巴蘭 回答 巴勒 的臣僕說：「 巴勒 就是將他滿屋的金銀給我，我也不能做任何大小的事，違背耶和華－我上帝的指示。
NUM|22|19|現在請你們今晚也在這裏住下，我好知道耶和華還要對我說甚麼。」
NUM|22|20|上帝在夜裏臨到 巴蘭 那裏，說：「這些人若來求你，你就起來跟他們去吧，只是你必須照著我對你說的話去做。」
NUM|22|21|巴蘭 早晨起來，備了驢，就和 摩押 的官員一同去了。
NUM|22|22|上帝因他去就怒氣發作；耶和華的使者站在路中間敵對他。他騎著驢，有兩個僕人跟隨他。
NUM|22|23|驢看見耶和華的使者站在路中間，手裏有拔出來的刀，就離開了路，岔入田間。 巴蘭 就打驢，要牠回到路上。
NUM|22|24|耶和華的使者站在葡萄園的窄路上，這邊有牆，那邊也有牆。
NUM|22|25|驢看見耶和華的使者，就往牆擠去，把 巴蘭 的腳擠到牆上； 巴蘭 再打驢。
NUM|22|26|耶和華的使者又往前去，站在狹窄的地方，那裏左右都無路可轉。
NUM|22|27|驢看見耶和華的使者，就伏在 巴蘭 底下。 巴蘭 怒氣發作，用杖打驢。
NUM|22|28|耶和華使驢開口，對 巴蘭 說：「我向你做了甚麼，你竟打我這三次呢？」
NUM|22|29|巴蘭 對驢說：「因為你戲弄我，我恨不得手中有刀，現在就把你殺了。」
NUM|22|30|驢對 巴蘭 說：「我不是你從小直到今天所騎的驢嗎？我平時有這樣待過你嗎？」 巴蘭 說：「沒有。」
NUM|22|31|耶和華使 巴蘭 的眼目明亮，他看見耶和華的使者站在路中間，手裏有拔出來的刀； 巴蘭 就低頭俯伏下拜。
NUM|22|32|耶和華的使者對他說：「你為甚麼這三次打你的驢呢？看哪，我出來敵對你，因為這路在我面前已經偏離了。
NUM|22|33|驢看見我就從我面前迴避了這三次；驢若沒有迴避我，我早把你殺了，留牠存活。」
NUM|22|34|巴蘭 對耶和華的使者說：「我有罪了。我不知道你站在路中間阻擋我；現在你若看為不好，我就回去。」
NUM|22|35|耶和華的使者對 巴蘭 說：「你和這些人去吧！你只要說我對你說的話。」於是 巴蘭 和 巴勒 的官員一同去了。
NUM|22|36|巴勒 聽見 巴蘭 來了，就到 摩押 的城 去迎接他；這城是在邊界的 亞嫩河 旁。
NUM|22|37|巴勒 對 巴蘭 說：「我不是急切地派人到你那裏去召你嗎？你為何不到我這裏來呢？我豈不能使你得尊榮嗎？」
NUM|22|38|巴蘭 對 巴勒 說：「看哪，我已經到你這裏來了！現在我豈能擅自說甚麼呢？上帝將甚麼話放在我口中，我就說甚麼。」
NUM|22|39|巴蘭 和 巴勒 同去，來到 基列‧胡瑣 。
NUM|22|40|巴勒 宰了牛羊為祭物，送給 巴蘭 和陪伴他的官員。
NUM|22|41|到了早晨， 巴勒 領 巴蘭 到 巴末‧巴力 ，從那裏可以看到一部分 以色列 的百姓。
NUM|23|1|巴蘭 對 巴勒 說：「你要在這裏為我築七座壇，又要在這裏為我預備七頭公牛，七隻公羊。」
NUM|23|2|巴勒 照 巴蘭 的話做了。 巴勒 和 巴蘭 在每座壇上獻一頭公牛，一隻公羊。
NUM|23|3|巴蘭 對 巴勒 說：「你站在你的燔祭旁邊，我要往前去，或許耶和華會向我顯現。他指示我甚麼事，我必告訴你。」於是 巴蘭 上到一個光禿的高地。
NUM|23|4|上帝向 巴蘭 顯現。 巴蘭 對他說：「我預備了七座壇，在每座壇上獻了一頭公牛，一隻公羊。」
NUM|23|5|耶和華把話放在 巴蘭 口中，說：「你回到 巴勒 那裏，要這樣說。」
NUM|23|6|他就回到 巴勒 那裏，看哪， 巴勒 和 摩押 的眾官員站在燔祭旁邊。
NUM|23|7|巴蘭 唱起詩歌說： 「 巴勒 領我出 亞蘭 ， 摩押 王領我出東方的山脈： 『來啊，為我詛咒 雅各 ； 來啊，怒罵 以色列 。』
NUM|23|8|上帝沒有詛咒的， 我焉能詛咒？ 耶和華沒有怒罵的， 我豈能怒罵？
NUM|23|9|我從磐石的巔峰看到他， 我從山丘望見他。 看哪，這是獨居的民， 不算在列國中。
NUM|23|10|誰能數點 雅各 的塵土？ 誰能計算 以色列 的塵沙 ？ 我願如正直人之死而死； 我願如正直人之終而終。」
NUM|23|11|巴勒 對 巴蘭 說：「你向我做的是甚麼呢？我帶你來詛咒我的仇敵，看哪，你竟為他們祝福。」
NUM|23|12|他回答說：「耶和華放在我口中的話，我豈能不謹慎地說呢？」
NUM|23|13|巴勒 對他說：「請你跟我到別的地方，在那裏可以看見他們。你只能看見他們的一部分，卻不能看見全部。請你在那裏為我詛咒他們。」
NUM|23|14|於是 巴勒 領 巴蘭 到了 瑣腓 的田野，上了 毗斯迦山 頂 ，築了七座壇，在每座壇上獻一頭公牛，一隻公羊。
NUM|23|15|巴蘭 對 巴勒 說：「你站在你的燔祭旁邊，我要到那邊去看看。」
NUM|23|16|耶和華向 巴蘭 顯現，把話放在他口中，說：「你回到 巴勒 那裏，要這樣說。」
NUM|23|17|他回到 巴勒 那裏，看哪， 巴勒 站在燔祭旁邊， 摩押 的官員也和他在一起。 巴勒 對他說：「耶和華說了甚麼呢？」
NUM|23|18|巴蘭 唱起詩歌說： 「 巴勒 啊，起來，聽； 西撥 的兒子啊，側耳聽我。
NUM|23|19|上帝非人，必不致說謊， 也非人子，必不致後悔。 他說了豈不照著做呢？ 他發了言豈不實現呢？
NUM|23|20|看哪，我奉命祝福； 上帝賜福，我不能扭轉。
NUM|23|21|他未見 雅各 中有災難 ， 也未見 以色列 中有禍患 。 耶和華－他的上帝和他同在； 在他中間有歡呼王的聲音。
NUM|23|22|上帝領他們出 埃及 ， 為 以色列 有如野牛的角。
NUM|23|23|絕沒有法術可以傷 雅各 ， 沒有占卜可以害 以色列 。 現在，人論及 雅各 ，論及 以色列 必說： 『上帝成就了何等的事啊！』
NUM|23|24|看哪，這百姓興起如母獅， 挺身像公獅， 未曾吃獵物， 未曾喝被殺者的血， 絕不躺臥。」
NUM|23|25|巴勒 對 巴蘭 說：「你一點也不要詛咒他們，一點也不要為他們祝福！」
NUM|23|26|巴蘭 回答 巴勒 說：「我不是告訴過你：『凡耶和華所說的，我必須遵行』嗎？」
NUM|23|27|巴勒 對 巴蘭 說：「來，我領你到別的地方，或許上帝喜歡你在那裏為我詛咒他們。」
NUM|23|28|巴勒 就領 巴蘭 到那可瞭望曠野的 毗珥山 頂。
NUM|23|29|巴蘭 對 巴勒 說：「你要在這裏為我築七座壇，又要在這裏為我預備七頭公牛，七隻公羊。」
NUM|23|30|巴勒 就照 巴蘭 的話做，在每座壇上獻一頭公牛，一隻公羊。
NUM|24|1|巴蘭 見耶和華喜歡賜福給 以色列 ，就不像前兩次去求法術，卻面向曠野。
NUM|24|2|巴蘭 舉目，看見 以色列 人照著支派紮營。上帝的靈就臨到他身上，
NUM|24|3|他唱起詩歌說： 「 比珥 的兒子 巴蘭 說， 眼目關閉 的人說，
NUM|24|4|聽見上帝的言語， 得見全能者的異象， 俯伏著，眼睛卻睜開的人說：
NUM|24|5|雅各 啊，你的帳棚何等華美！ 以色列 啊，你的帳幕何其華麗！
NUM|24|6|如連綿的山谷， 如河畔的園子， 如耶和華栽種的沉香樹， 又如水邊的香柏木。
NUM|24|7|水要從他的桶裏流出， 種子要撒在多水之處。 他的王必超越 亞甲 ， 他的國必要振興。
NUM|24|8|上帝領他出 埃及 ， 為他有如野牛的角。 他要吞滅那敵對他的國， 壓碎他們的骨頭， 用箭射透他們。
NUM|24|9|他蹲如公獅， 臥如母獅， 誰敢惹他？ 凡為你祝福的，願他蒙福； 凡詛咒你的，願他受詛咒。」
NUM|24|10|巴勒 向 巴蘭 怒氣發作，就緊握拳頭 。 巴勒 對 巴蘭 說：「我召你來詛咒我的仇敵，看哪，你竟然這三次為他們祝福。
NUM|24|11|如今你趕快回本地去吧！我想使你大得尊榮，看哪，耶和華卻阻止你得尊榮。」
NUM|24|12|巴蘭 對 巴勒 說：「我不是對你所差遣到我那裏的使者說：
NUM|24|13|『 巴勒 就是把他滿屋的金銀給我，我也不能違背耶和華的指示，隨自己的心意做好做歹。耶和華說甚麼，我就說甚麼。』
NUM|24|14|現在，看哪，我要回到我的百姓那裏。來，讓我告訴你這百姓日後要怎樣對待你的百姓。」
NUM|24|15|他就唱起詩歌說： 「 比珥 的兒子 巴蘭 說， 眼目關閉的人說，
NUM|24|16|聽見上帝的言語， 明白至高者的知識， 看見全能者的異象， 俯伏著，眼睛卻睜開的人說：
NUM|24|17|我看見他，卻不在現時； 我望見他，卻不在近處。 有星出於 雅各 ， 有杖從 以色列 興起， 必打破 摩押 的額頭， 必毀壞所有的 塞特 人 。
NUM|24|18|以東 將成為產業， 西珥 將成為它敵人的產業 ； 但 以色列 卻要得勝。
NUM|24|19|有一位出於 雅各 的，必掌大權， 他要除滅城中的倖存者。」
NUM|24|20|巴蘭 看見 亞瑪力 人，就唱起詩歌說： 「 亞瑪力 是諸國之首， 但它終必永遠沉淪 。」
NUM|24|21|巴蘭 看見 基尼 人，就唱起詩歌說： 「你的住處堅固； 你的巢窩造在巖石中。
NUM|24|22|然而 基尼 族 必被吞滅， 直到何時 亞述 把你擄去？ 」
NUM|24|23|巴蘭 又唱起詩歌說： 「哀哉！若上帝做這事， 誰能存活呢？
NUM|24|24|有船隻 從 基提 邊界來到， 要壓制 亞述 ， 要壓制 希伯 ； 他也必永遠沉淪 。」
NUM|24|25|於是 巴蘭 起來，回本地去； 巴勒 也回他的路去了。
NUM|25|1|以色列 人住在 什亭 ，百姓開始與 摩押 女子行淫。
NUM|25|2|這些女子請百姓一同為她們的神明獻祭，百姓吃了祭物，跪拜她們的神明。
NUM|25|3|以色列 與 巴力‧毗珥 聯合，耶和華的怒氣就向 以色列 發作。
NUM|25|4|耶和華對 摩西 說：「拿下百姓中所有的領袖，對著太陽把他們懸掛在我面前，使我向 以色列 所發的怒氣可以平息。」
NUM|25|5|於是 摩西 對 以色列 的審判官說：「你們的人若有與 巴力‧毗珥 聯合的，你們各人就要把他們殺了。」
NUM|25|6|摩西 和 以色列 全會眾在會幕門口哭泣的時候，看哪，有一個 以色列 人，在他們眼前帶著一個 米甸 女子，到他弟兄那裏。
NUM|25|7|亞倫 祭司的孫子， 以利亞撒 的兒子 非尼哈 看見了，就從會眾中起來，手裏拿著槍，
NUM|25|8|跟這 以色列 人進入帳棚，刺穿了二人，就是 以色列 人和那女子的肚腹。這樣， 以色列 人遭受的瘟疫就停止了。
NUM|25|9|遭瘟疫死的，有二萬四千人。
NUM|25|10|耶和華吩咐 摩西 說：
NUM|25|11|「 亞倫 祭司的孫子， 以利亞撒 的兒子 非尼哈 ，使我的憤怒轉離 以色列 人，因為在他們中間，他以我的妒忌為他的妒忌，使我不在妒忌中毀滅 以色列 人。
NUM|25|12|因此，你要說：『看哪，我將我平安的約賜給他。
NUM|25|13|這是他和他的後裔永遠當祭司職任的約，因他為了上帝而妒忌，他為 以色列 人贖罪。』」
NUM|25|14|那與 米甸 女子一起被殺的 以色列 人，名叫 心利 ，是 撒路 的兒子，是 西緬 一個父家的領袖。
NUM|25|15|那被殺的 米甸 女子，名叫 哥斯比 ，是 蘇珥 的女兒； 蘇珥 是 米甸 一個父家的領袖。
NUM|25|16|耶和華吩咐 摩西 說：
NUM|25|17|「你要苦害 米甸 人，擊殺他們；
NUM|25|18|因為他們用詭計苦害你們，在 毗珥 的事上和他們的姊妹， 米甸 領袖的女兒 哥斯比 的事上，欺騙了你們；在瘟疫的日子，這女子因 毗珥 的事件被殺了。」
NUM|26|1|瘟疫過了之後，耶和華對 摩西 和 亞倫 祭司的兒子 以利亞撒 說：
NUM|26|2|「你們要將 以色列 全會眾，按他們的父家，凡二十歲以上能出去為 以色列 打仗的，計算總數。」
NUM|26|3|摩西 和 以利亞撒 祭司在 摩押 平原與 耶利哥 相對的 約旦河 邊吩咐他們說：
NUM|26|4|「計算你們中間從二十歲以上的人數。」正如耶和華所吩咐 摩西 的。 從 埃及 地出來的 以色列 人如下：
NUM|26|5|以色列 的長子是 呂便 。 呂便 的眾子：屬 哈諾 的，有 哈諾 族；屬 法路 的，有 法路 族；
NUM|26|6|屬 希斯倫 的，有 希斯倫 族；屬 迦米 的，有 迦米 族。
NUM|26|7|這就是 呂便 的各族；被數的共有四萬三千七百三十名。
NUM|26|8|法路 的兒子是 以利押 。
NUM|26|9|以利押 的兒子是 尼母利 、 大坍 、 亞比蘭 。這 大坍 、 亞比蘭 ，就是從會中選出來，當 可拉 一夥的人向耶和華爭鬧的時候，一起向 摩西 、 亞倫 爭鬧的；
NUM|26|10|地開了裂口，吞了他們和 可拉 ， 可拉 一夥的人也一同死亡。當時火吞滅了二百五十個人；他們就成為鑑戒。
NUM|26|11|然而 可拉 的眾子沒有死亡。
NUM|26|12|按著宗族， 西緬 的眾子：屬 尼母利 的，有 尼母利 族；屬 雅憫 的，有 雅憫 族；屬 雅斤 的，有 雅斤 族；
NUM|26|13|屬 謝拉 的，有 謝拉 族；屬 掃羅 的，有 掃羅 族。
NUM|26|14|這就是 西緬 的各族，共有二萬二千二百名。
NUM|26|15|按著宗族， 迦得 的眾子：屬 洗分 的，有 洗分 族；屬 哈基 的，有 哈基 族；屬 書尼 的，有 書尼 族；
NUM|26|16|屬 阿斯尼 的，有 阿斯尼 族；屬 以利 的，有 以利 族；
NUM|26|17|屬 亞律 的，有 亞律 族；屬 亞列利 的，有 亞列利 族。
NUM|26|18|這就是 迦得 子孫的各族；他們被數的共有四萬零五百名。
NUM|26|19|猶大 的兒子是 珥 和 俄南 。 珥 和 俄南 死在 迦南 地。
NUM|26|20|按著宗族， 猶大 的眾子：屬 示拉 的，有 示拉 族；屬 法勒斯 的，有 法勒斯 族；屬 謝拉 的，有 謝拉 族。
NUM|26|21|法勒斯 的眾子：屬 希斯崙 的，有 希斯崙 族；屬 哈母勒 的，有 哈母勒 族。
NUM|26|22|這就是 猶大 的各族；他們被數的共有七萬六千五百名。
NUM|26|23|按著宗族， 以薩迦 的眾子：屬 陀拉 的，有 陀拉 族；屬 普瓦 的，有 普瓦 族；
NUM|26|24|屬 雅述 的，有 雅述 族；屬 伸崙 的，有 伸崙 族。
NUM|26|25|這就是 以薩迦 的各族；他們被數的共有六萬四千三百名。
NUM|26|26|按著宗族， 西布倫 的眾子：屬 西烈 的，有 西烈 族；屬 以倫 的，有 以倫 族；屬 雅利 的，有 雅利 族。
NUM|26|27|這就是 西布倫 的各族；他們被數的共有六萬零五百名。
NUM|26|28|按著宗族， 約瑟 的兒子有 瑪拿西 、 以法蓮 。
NUM|26|29|瑪拿西 的眾子：屬 瑪吉 的，有 瑪吉 族； 瑪吉 生 基列 ；屬 基列 的，有 基列 族。
NUM|26|30|這就是 基列 的眾子：屬 伊以謝 的，有 伊以謝 族；屬 希勒 的，有 希勒 族；
NUM|26|31|屬 亞斯烈 的，有 亞斯烈 族；屬 示劍 的，有 示劍 族；
NUM|26|32|屬 示米大 的，有 示米大 族；屬 希弗 的，有 希弗 族。
NUM|26|33|希弗 的兒子 西羅非哈 沒有兒子，只有女兒。 西羅非哈 的女兒的名字是 瑪拉 、 挪阿 、 曷拉 、 密迦 、 得撒 。
NUM|26|34|這就是 瑪拿西 的各族；他們被數的共有五萬二千七百名。
NUM|26|35|這就是按著宗族， 以法蓮 的眾子：屬 書提拉 的，有 書提拉 族；屬 比結 的，有 比結 族；屬 他罕 的，有 他罕 族。
NUM|26|36|這就是 書提拉 的眾子：屬 以蘭 的，有 以蘭 族。
NUM|26|37|這就是 以法蓮 子孫的各族；他們被數的共有三萬二千五百名。按著宗族，以上這些都是 約瑟 的子孫。
NUM|26|38|按著宗族， 便雅憫 的眾子：屬 比拉 的，有 比拉 族；屬 亞實別 的，有 亞實別 族；屬 亞希蘭 的，有 亞希蘭 族；
NUM|26|39|屬 書反 的，有 書反 族；屬 戶反 的，有 戶反 族。
NUM|26|40|比拉 的兒子是 亞勒 、 乃幔 ；屬 亞勒 的 ，有 亞勒 族；屬 乃幔 的，有 乃幔 族。
NUM|26|41|按著宗族，這就是 便雅憫 的子孫；他們被數的共有四萬五千六百名。
NUM|26|42|這就是按著宗族， 但 的眾子：屬 書含 的，有 書含 族。按著宗族，這就是 但 的各族。
NUM|26|43|按照他們被數的， 書含 全宗族共有六萬四千四百名。
NUM|26|44|按著宗族， 亞設 的眾子：屬 音拿 的，有 音拿 族；屬 亦施韋 的，有 亦施韋 族；屬 比利亞 的，有 比利亞 族。
NUM|26|45|比利亞 的眾子：屬 希別 的，有 希別 族；屬 瑪結 的，有 瑪結 族。
NUM|26|46|亞設 的女兒名叫 西拉 。
NUM|26|47|這就是 亞設 子孫的各族；他們被數的共有五萬三千四百名。
NUM|26|48|按著宗族， 拿弗他利 的眾子：屬 雅薛 的，有 雅薛 族；屬 沽尼 的，有 沽尼 族；
NUM|26|49|屬 耶色 的，有 耶色 族；屬 示冷 的，有 示冷 族。
NUM|26|50|按著宗族，這就是 拿弗他利 的各族；他們被數的共有四萬五千四百名。
NUM|26|51|這就是 以色列 人中被數的，共有六十萬零一千七百三十名。
NUM|26|52|耶和華吩咐 摩西 說：
NUM|26|53|「你要按著人名的數目，將地分給這些人為產業。
NUM|26|54|人多的要多給他們產業，人少的要少給他們產業；各照被數的人數分配產業。
NUM|26|55|此外，要以抽籤來分地，按著父系各支派的名字承受產業。
NUM|26|56|要根據抽籤，看人數的多寡，給他們分配產業。」
NUM|26|57|這就是按著宗族，被數的 利未 人：屬 革順 的，有 革順 族；屬 哥轄 的，有 哥轄 族；屬 米拉利 的，有 米拉利 族。
NUM|26|58|這就是 利未 的宗族： 立尼 族、 希伯倫 族、 瑪利 族、 母示 族、 可拉 族。 哥轄 生 暗蘭 。
NUM|26|59|暗蘭 的妻子名叫 約基別 ，是 利未 的女兒，是 利未 在 埃及 所生的。她給 暗蘭 生了 亞倫 、 摩西 ，和他們的姊姊 米利暗 。
NUM|26|60|亞倫 生 拿答 、 亞比戶 、 以利亞撒 、 以他瑪 。
NUM|26|61|拿答 、 亞比戶 在耶和華面前獻凡火的時候死了。
NUM|26|62|利未 人中，凡一個月以上所有被數的男子，共有二萬三千名。他們沒有數在 以色列 人中；因為在 以色列 人中，沒有分給他們產業。
NUM|26|63|這些是 摩西 和 以利亞撒 祭司所數的；他們在 摩押 平原與 耶利哥 相對的 約旦河 邊數點 以色列 人。
NUM|26|64|這些被數的人中，沒有一個是 摩西 和 亞倫 祭司先前在 西奈 曠野所數的 以色列 人，
NUM|26|65|因為耶和華論到他們說：「他們必死在曠野。」所以，除了 耶孚尼 的兒子 迦勒 和 嫩 的兒子 約書亞 以外，他們一個也沒有存留。
NUM|27|1|約瑟 的兒子 瑪拿西 的宗族中，有 瑪拿西 的玄孫， 瑪吉 的曾孫， 基列 的孫子， 希弗 的兒子 西羅非哈 的女兒，名叫 瑪拉 、 挪阿 、 曷拉 、 密迦 、 得撒 。她們前來，
NUM|27|2|站在會幕門口，在 摩西 和 以利亞撒 祭司，以及眾領袖與全會眾面前，說：
NUM|27|3|「我們的父親死在曠野。他沒有與 可拉 同夥聚集攻擊耶和華，是在自己的罪中死的；他沒有兒子。
NUM|27|4|為甚麼因我們的父親沒有兒子就把他的名從他族中除掉呢？求你們在我們父親的兄弟中分給我們產業。」
NUM|27|5|於是， 摩西 將她們的案件呈到耶和華面前。
NUM|27|6|耶和華對 摩西 說：
NUM|27|7|「 西羅非哈 的女兒說得有理。你定要在她們父親的兄弟中，把地分給她們為業，把她們父親的產業傳給她們。
NUM|27|8|你也要吩咐 以色列 人說：『人死了，若沒有兒子，就要把他的產業傳給他的女兒。
NUM|27|9|他若沒有女兒，就要把他的產業給他的兄弟。
NUM|27|10|他若沒有兄弟，就要把他的產業給他父親的兄弟。
NUM|27|11|他父親若沒有兄弟，就要把他的產業給他族中最近的親屬繼承為業。』」這要作 以色列 人的律例典章，是照耶和華所吩咐 摩西 的。
NUM|27|12|耶和華對 摩西 說：「你上這 亞巴琳山脈 ，看我所賜給 以色列 人的地。
NUM|27|13|看了以後，你也必歸到你祖先 那裏，像你哥哥 亞倫 歸去一樣。
NUM|27|14|因為你們在 尋 的曠野，當會眾爭鬧的時候，違背了我的命令，在取水之事上沒有在會眾眼前尊我為聖。」這水就是 尋 的曠野中， 加低斯 的 米利巴 水。
NUM|27|15|摩西 對耶和華說：
NUM|27|16|「願耶和華，賜萬人氣息的上帝，立一個人治理會眾，
NUM|27|17|可以在他們面前出入，引導他們進出，免得耶和華的會眾如同沒有牧人的羊群一般。」
NUM|27|18|耶和華對 摩西 說：「 嫩 的兒子 約書亞 是一個有聖靈的人；你要領他來，為他按手，
NUM|27|19|使他站在 以利亞撒 祭司和全會眾面前，在他們眼前委派他，
NUM|27|20|又將你的尊榮給他一些，好使 以色列 全會眾都聽從他。
NUM|27|21|他要站在 以利亞撒 祭司面前； 以利亞撒 要憑烏陵的判斷，在耶和華面前為他求問。他和 以色列 全會眾都要照 以利亞撒 的指示出入。」
NUM|27|22|於是 摩西 照耶和華所吩咐他的，將 約書亞 領來，使他站在 以利亞撒 祭司和全會眾面前，
NUM|27|23|為他按手，委派他，是照耶和華藉 摩西 所說的。
NUM|28|1|耶和華吩咐 摩西 說：
NUM|28|2|「你要吩咐 以色列 人說：『你們要按時把我的供物，就是獻給我作馨香火祭的食物，獻給我。』
NUM|28|3|要對他們說：『這是當獻給耶和華的火祭：每天兩隻沒有殘疾一歲的小公羊，作為經常獻的燔祭。
NUM|28|4|早晨獻第一隻小公羊，黃昏獻第二隻小公羊；
NUM|28|5|又用十分之一伊法細麵和四分之一欣搗成的油，調和作為素祭。
NUM|28|6|這是在 西奈山 上規定為經常獻的燔祭，是獻給耶和華為馨香的火祭。
NUM|28|7|為每隻小公羊，要有四分之一欣的澆酒祭；在聖所中，你要將醇酒獻給耶和華作澆酒祭。
NUM|28|8|黃昏你獻第二隻小公羊，要照早晨的素祭和同獻的澆酒祭獻上，作為馨香的火祭，獻給耶和華。』」
NUM|28|9|「在安息日，要獻兩隻沒有殘疾，一歲的小公羊、十分之二伊法調了油的細麵為素祭，和同獻的澆酒祭。
NUM|28|10|除了經常獻的燔祭和同獻的澆酒祭之外，這是每一個安息日當獻的燔祭。」
NUM|28|11|「每月初一，要將兩頭公牛犢、一隻公綿羊、七隻沒有殘疾一歲的小公羊，獻給耶和華為燔祭。
NUM|28|12|為每頭公牛，要用十分之三伊法調了油的細麵作為素祭；為那隻公綿羊，要用十分之二伊法調了油的細麵作為素祭；
NUM|28|13|為每隻小公羊，要用十分之一伊法調了油的細麵作為素祭。這是馨香的燔祭，是獻給耶和華的火祭。
NUM|28|14|每頭公牛要有半欣的澆酒祭，每隻公綿羊三分之一欣的澆酒祭，每隻小公羊四分之一欣的澆酒祭。這是一年之中每月初一當獻的燔祭。
NUM|28|15|除了經常獻的燔祭和同獻的澆酒祭之外，又要將一隻公山羊，獻給耶和華為贖罪祭。」
NUM|28|16|「正月十四日是向耶和華守的逾越節。
NUM|28|17|這月十五日是節期，要吃無酵餅七日。
NUM|28|18|第一日要有聖會，任何勞動的工都不可做。
NUM|28|19|要把火祭，就是兩頭公牛犢，一隻公綿羊、七隻一歲的小公羊，都要沒有殘疾的，獻給耶和華為燔祭。
NUM|28|20|要同時獻調了油的細麵為素祭：每頭公牛要獻十分之三伊法；每隻公綿羊要獻十分之二伊法；
NUM|28|21|為那七隻小公羊，每隻要獻十分之一伊法。
NUM|28|22|此外，要獻一隻公山羊作贖罪祭，為你們贖罪。
NUM|28|23|除了早晨經常獻的燔祭之外，你們也要獻這些祭。
NUM|28|24|一連七天，在經常獻的燔祭和同獻的澆酒祭之外，每天要這樣把馨香火祭的食物獻給耶和華。
NUM|28|25|第七日要有聖會，任何勞動的工都不可做。」
NUM|28|26|「七七初熟節，就是你們獻初熟穀物給耶和華為素祭的那一天，要宣告聖會；任何勞動的工都不可做。
NUM|28|27|要將兩頭公牛犢，一隻公綿羊，七隻一歲的小公羊，作為馨香的燔祭獻給耶和華。
NUM|28|28|要同時獻調了油的細麵為素祭：每頭公牛要獻十分之三伊法；每隻公綿羊要獻十分之二伊法；
NUM|28|29|為那七隻小公羊，每隻要獻十分之一伊法。
NUM|28|30|此外，要獻一隻公山羊為你們贖罪。
NUM|28|31|除了經常獻的燔祭和同獻的素祭，你們也要獻上這些沒有殘疾的，和同獻的澆酒祭。」
NUM|29|1|「七月初一，你們當有聖會；任何勞動的工都不可做，是你們當守為吹角的日子。
NUM|29|2|你們要將一頭公牛犢、一隻公綿羊、七隻一歲的小公羊，都是沒有殘疾的，獻給耶和華為馨香的燔祭。
NUM|29|3|要同時獻調了油的細麵為素祭：每頭公牛要獻十分之三伊法；每隻公綿羊要獻十分之二伊法；
NUM|29|4|為那七隻小公羊，每隻要獻十分之一伊法。
NUM|29|5|此外，要獻一隻公山羊作贖罪祭，為你們贖罪。
NUM|29|6|除了初一的燔祭和同獻的素祭、經常獻的燔祭與同獻的素祭，以及同獻的澆酒祭以外，這些都照例作為馨香的火祭獻給耶和華。」
NUM|29|7|「七月初十，你們當有聖會；要刻苦己心，任何工都不可做。
NUM|29|8|要將一頭公牛犢、一隻公綿羊、七隻一歲的小公羊，都是沒有殘疾的，獻給耶和華為馨香的燔祭。
NUM|29|9|要同時獻調了油的細麵為素祭：每頭公牛要獻十分之三伊法；每隻公綿羊要獻十分之二伊法；
NUM|29|10|為那七隻小公羊，每隻要獻十分之一伊法。
NUM|29|11|又要獻一隻公山羊為贖罪祭。這是在贖罪祭和經常獻的燔祭，以及同獻的素祭和澆酒祭以外所獻的。」
NUM|29|12|「七月十五日，你們當有聖會；任何勞動的工都不可做，要向耶和華守節七天。
NUM|29|13|要將十三頭公牛犢、兩隻公綿羊、十四隻一歲的小公羊，都是沒有殘疾的，獻上作火祭，是獻給耶和華馨香的燔祭。
NUM|29|14|要同時獻調了油的細麵為素祭：為那十三頭公牛犢，每頭要獻十分之三伊法；為那兩隻公綿羊，每隻要獻十分之二伊法；
NUM|29|15|為那十四隻小公羊，每隻要獻十分之一伊法。
NUM|29|16|又要獻一隻公山羊為贖罪祭。這是在經常獻的燔祭、同獻的素祭和澆酒祭以外所獻的。
NUM|29|17|「第二日要獻十二頭公牛犢、兩隻公綿羊、十四隻一歲的小公羊，都是沒有殘疾的，
NUM|29|18|並為公牛、公綿羊和小公羊，按數照例奉獻同獻的素祭和澆酒祭。
NUM|29|19|又要獻一隻公山羊為贖罪祭。這是在經常獻的燔祭、同獻的素祭和澆酒祭以外所獻的。
NUM|29|20|「第三日要獻十一頭公牛、兩隻公綿羊、十四隻一歲的小公羊，都是沒有殘疾的，
NUM|29|21|並為公牛、公綿羊和小公羊，按數照例奉獻同獻的素祭和澆酒祭。
NUM|29|22|又要獻一隻公山羊為贖罪祭。這是在經常獻的燔祭、同獻的素祭和澆酒祭以外所獻的。
NUM|29|23|「第四日要獻十頭公牛、兩隻公綿羊、十四隻一歲的小公羊，都是沒有殘疾的，
NUM|29|24|並為公牛、公綿羊和小公羊，按數照例奉獻同獻的素祭和澆酒祭。
NUM|29|25|又要獻一隻公山羊為贖罪祭。這是在經常獻的燔祭、同獻的素祭和澆酒祭以外所獻的。
NUM|29|26|「第五日要獻九頭公牛、兩隻公綿羊、十四隻一歲的小公羊，都是沒有殘疾的，
NUM|29|27|並為公牛、公綿羊和小公羊，按數照例奉獻同獻的素祭和澆酒祭。
NUM|29|28|又要獻一隻公山羊為贖罪祭。這是在經常獻的燔祭、同獻的素祭和澆酒祭以外所獻的。
NUM|29|29|「第六日要獻八頭公牛、兩隻公綿羊、十四隻一歲的小公羊，都是沒有殘疾的，
NUM|29|30|並為公牛、公綿羊和小公羊，按數照例奉獻同獻的素祭和澆酒祭。
NUM|29|31|又要獻一隻公山羊為贖罪祭。這是在經常獻的燔祭、同獻的素祭和澆酒祭以外所獻的。
NUM|29|32|「第七日要獻七頭公牛、兩隻公綿羊、十四隻一歲的小公羊，都是沒有殘疾的，
NUM|29|33|並為公牛、公綿羊和小公羊，按數照例奉獻同獻的素祭和澆酒祭。
NUM|29|34|又要獻一隻公山羊為贖罪祭。這是在經常獻的燔祭、同獻的素祭和澆酒祭以外所獻的。
NUM|29|35|「第八日你們當有嚴肅會；任何勞動的工都不可做；
NUM|29|36|要將一頭公牛、一隻公綿羊、七隻一歲的小公羊，都是沒有殘疾的，獻上作火祭，是獻給耶和華馨香的燔祭。
NUM|29|37|要為公牛、公綿羊和小公羊，按數照例奉獻同獻的素祭和澆酒祭。
NUM|29|38|又要獻一隻公山羊為贖罪祭。這是在經常獻的燔祭、同獻的素祭和澆酒祭以外所獻的。
NUM|29|39|「這些祭要在你們的節期獻給耶和華，都是在所許的願和甘心獻的以外所獻的，作為你們的燔祭、素祭、澆酒祭和平安祭。」
NUM|29|40|於是， 摩西 照耶和華所吩咐他的一切話告訴 以色列 人。
NUM|30|1|摩西 對 以色列 各支派的領袖說：「這是耶和華所吩咐的話：
NUM|30|2|人若向耶和華許願或起誓，要約束自己，就不可食言，必須照口中所出的一切話去做。
NUM|30|3|女子年輕，還在父家的時候，若向耶和華許願，要約束自己，
NUM|30|4|她父親聽見她所許的願和約束自己的話，卻向她默默不言，她所許的願和約束自己的話就都有效。
NUM|30|5|但是，若她父親在聽見的日子不允許她一切所許的願和約束自己的話，這就不算為有效；耶和華也必赦免她，因為她的父親不允許。
NUM|30|6|她若已出嫁，有願在身，或口中出了約束自己的冒失話，
NUM|30|7|她丈夫聽見了，卻在聽見的日子向她默默不言，她所許的願和約束自己的話就都有效。
NUM|30|8|但是，若她丈夫在聽見的日子不允許，丈夫就廢了她所許的願和口中所出約束自己的冒失話；耶和華也必赦免她。
NUM|30|9|寡婦或被休的婦人所許的願，她所有約束自己的話，都是有效的。
NUM|30|10|她若在丈夫家裏許了願或起了誓，要約束自己，
NUM|30|11|丈夫聽見了，卻向她默默不言，沒有不允許，她所許的願和約束自己的話就都有效。
NUM|30|12|她丈夫聽見的日子，若把這些全廢了，她口中一切所許的願或約束自己的話就不算為有效。她丈夫已把這些都廢了，耶和華也必赦免她。
NUM|30|13|凡她所許的願和刻苦約束自己所起的誓，丈夫可以堅立，也可以廢去。
NUM|30|14|倘若她丈夫天天向她默默不言，這就算是堅立她一切所許的願或約束自己的話；因為丈夫在聽見的日子向她默默不言，就算是堅立了這些話。
NUM|30|15|但她丈夫聽見了，以後若再廢了這些話，就要擔當婦人的罪孽。」
NUM|30|16|這是關於丈夫待妻子，父親待女兒，女兒年輕還在父家，耶和華所吩咐 摩西 的條例。
NUM|31|1|耶和華吩咐 摩西 說：
NUM|31|2|「你要為 以色列 人向 米甸 人報仇，然後歸到你祖先 那裏。」
NUM|31|3|摩西 吩咐百姓說：「要在你們中間叫人帶兵器去攻擊 米甸 ，為耶和華向 米甸 報仇。
NUM|31|4|從 以色列 眾支派中，每支派要派一千人去打仗。」
NUM|31|5|於是從 以色列 千萬人中，每支派徵召一千人，一共一萬二千名，帶著兵器預備打仗。
NUM|31|6|摩西 派他們去打仗，每支派一千人；又派 以利亞撒 祭司的兒子 非尼哈 同去； 非尼哈 手裏拿著聖所的器皿和吹號的號筒。
NUM|31|7|他們遵照耶和華所吩咐 摩西 的，與 米甸 打仗，殺了所有的男丁。
NUM|31|8|在所殺的人中，他們殺了 米甸 的王，就是 以未 、 利金 、 蘇珥 、 戶珥 、 利巴 五個 米甸 的王，又用刀殺了 比珥 的兒子 巴蘭 。
NUM|31|9|以色列 人擄了 米甸 的婦女和孩童，搶奪他們一切的牲畜、牛羊和所有的財物，
NUM|31|10|又用火焚燒了他們所住的一切城鎮和所有的營寨。
NUM|31|11|以色列 人把一切擄物和掠物，連人和牲畜都帶走，
NUM|31|12|將俘虜、掠物、擄物帶到 摩押 平原，在 約旦河 邊與 耶利哥 相對的營地，交給 摩西 和 以利亞撒 祭司，以及 以色列 的會眾。
NUM|31|13|摩西 和 以利亞撒 祭司，以及會眾中所有的領袖，都出營迎接他們。
NUM|31|14|摩西 向打仗回來的軍官，就是千夫長和百夫長發怒。
NUM|31|15|摩西 對他們說：「你們要讓這所有的婦女活著嗎？
NUM|31|16|看哪，正是這些婦女，因 巴蘭 的話，在 毗珥 的事上導致 以色列 人背叛耶和華，以致耶和華的會眾遭遇瘟疫。
NUM|31|17|現在，你們要殺所有的男孩，也要把所有曾與男人同房共寢的女子都殺了。
NUM|31|18|但那些未曾與男人同房共寢的女孩，你們可以讓她們存活。
NUM|31|19|你們和你們所擄來的人，要住在營外七天；凡殺了人的，和一切摸了屍體的，要在第三日和第七日潔淨自己。
NUM|31|20|你們也要潔淨一切的衣服，以及用皮革、山羊毛和木頭做的任何東西。」
NUM|31|21|以利亞撒 祭司對打仗回來的士兵說：「耶和華所吩咐 摩西 律法中的條例是這樣：
NUM|31|22|金、銀、銅、鐵、錫、鉛，
NUM|31|23|凡能耐火的，你們要使它經過火，它就潔淨，然而還要用除污穢的水來潔淨它；凡不能耐火的，你們要使它經過水。
NUM|31|24|第七日，你們要洗衣服，才為潔淨，然後可以進營。」
NUM|31|25|耶和華對 摩西 說：
NUM|31|26|「你和 以利亞撒 祭司，以及會眾的各父系家長，要計算所擄掠的人和牲畜的總數。
NUM|31|27|要把所擄掠的分成兩半：一半給那出去打仗的精兵，一半給全會眾。
NUM|31|28|再從那出去打仗的戰士所得的人、牛、驢、羊中，每五百取一，獻給耶和華為貢物。
NUM|31|29|要從他們那一半中取出這些，交給 以利亞撒 祭司，作為耶和華的舉祭。
NUM|31|30|又要從 以色列 人的那一半中，就是從人、牛、驢、羊，各樣牲畜中，每五十取一，交給照管耶和華帳幕的 利未 人。」
NUM|31|31|於是 摩西 和 以利亞撒 祭司遵照耶和華所吩咐 摩西 的做了。
NUM|31|32|除了士兵所奪的財物以外，所擄來的有羊六十七萬五千隻，
NUM|31|33|牛七萬二千頭，
NUM|31|34|驢六萬一千匹；
NUM|31|35|至於人，就是未曾與男人同房共寢的女子，總共三萬二千名。
NUM|31|36|出去打仗之人的那分，就是他們所得的一半，共計羊三十三萬七千五百隻，
NUM|31|37|其中歸耶和華為貢物的羊，六百七十五隻；
NUM|31|38|牛三萬六千頭，其中歸耶和華為貢物的七十二頭；
NUM|31|39|驢三萬零五百匹，其中歸耶和華為貢物的六十一匹；
NUM|31|40|人一萬六千名，其中歸耶和華的三十二名。
NUM|31|41|摩西 把貢物，就是歸給耶和華的舉祭，交給 以利亞撒 祭司，是照耶和華所吩咐 摩西 的。
NUM|31|42|以色列 人所得的另一半，是 摩西 從打仗的人取來分給他們的。
NUM|31|43|會眾的這一半有羊三十三萬七千五百隻，
NUM|31|44|牛三萬六千頭，
NUM|31|45|驢三萬零五百匹，
NUM|31|46|人一萬六千名。
NUM|31|47|無論是人或牲畜， 摩西 都每五十取一，交給照管耶和華帳幕的 利未 人，是照耶和華所吩咐 摩西 的。
NUM|31|48|帶領眾軍隊的軍官，就是千夫長、百夫長，進到 摩西 那裏，
NUM|31|49|對他說：「你的僕人已經計算屬下戰士的總數，一個也沒有少。
NUM|31|50|如今我們把各人所得的金器，就是腳鏈子、手鐲、打印的戒指、耳環、項鏈，都送給耶和華為供物，好在耶和華面前為我們贖罪。」
NUM|31|51|摩西 和 以利亞撒 祭司就收了他們的金子，就是各樣的首飾。
NUM|31|52|千夫長、百夫長所獻給耶和華為舉祭的金子共有一萬六千七百五十舍客勒。
NUM|31|53|打仗的人都把自己所掠奪的各自留下。
NUM|31|54|摩西 和 以利亞撒 祭司收了千夫長、百夫長的金子，就帶進會幕，好使 以色列 人在耶和華面前蒙記念。
NUM|32|1|呂便 子孫和 迦得 子孫的牲畜極其眾多。他們看到 雅謝 地和 基列 地；看哪，這是可牧放牲畜的地方。
NUM|32|2|呂便 子孫和 迦得 子孫就到 摩西 和 以利亞撒 祭司，以及會眾的領袖那裏，說：
NUM|32|3|「 亞他錄 、 底本 、 雅謝 、 寧拉 、 希實本 、 以利亞利 、 示班 、 尼波 、 比穩 ，
NUM|32|4|就是耶和華在 以色列 會眾面前所攻取之地，是可牧放牲畜之地，而你的僕人也有牲畜。」
NUM|32|5|又說：「我們若在你眼前蒙恩，求你把這地給我們為業；不要領我們過 約旦河 。」
NUM|32|6|摩西 對 迦得 子孫和 呂便 子孫說：「難道你們的弟兄去打仗，你們卻留在這裏嗎？
NUM|32|7|你們為甚麼使 以色列 人灰心，不渡過去，進入耶和華所賜給他們的那地呢？
NUM|32|8|我從 加低斯‧巴尼亞 派你們的父執之輩去窺探那地時，他們就曾這樣做過。
NUM|32|9|他們上到 以實各谷 ，窺探了那地之後，竟然使 以色列 人灰心，不願進入耶和華所賜給他們的地。
NUM|32|10|當日，耶和華的怒氣發作，起誓說：
NUM|32|11|『凡從 埃及 上來二十歲以上的人，斷不得看見我對 亞伯拉罕 、 以撒 、 雅各 起誓應許之地，因為他們沒有專心跟從我；
NUM|32|12|惟有 基尼洗 族 耶孚尼 的兒子 迦勒 ，還有 嫩 的兒子 約書亞 可以看見，因為他們專心跟從耶和華。』
NUM|32|13|耶和華的怒氣向 以色列 發作，使他們在曠野飄流四十年，直到在耶和華眼前作惡的那一代都消滅了。
NUM|32|14|看哪，你們這一夥罪人，竟然接續你們父執之輩，再增加耶和華對 以色列 所發的怒氣。
NUM|32|15|你們若轉離不跟從他，他要再把 以色列 人撇在曠野；這樣，你們就使這眾百姓滅亡了。」
NUM|32|16|他們挨近 摩西 ，說：「我們要在這裏為牲畜築圈，為孩童建城。
NUM|32|17|我們自己卻要帶兵器，急速行在 以色列 人的前面，領他們直到他們的地方。我們的孩童可以留在堅固的城內，躲避當地的居民。
NUM|32|18|我們必不回自己的家，直等到 以色列 人各自承受了自己的產業。
NUM|32|19|我們不和他們在 約旦河 那邊分產業，因為我們的產業是在 約旦河 的東邊。」
NUM|32|20|摩西 對他們說：「你們若要這麼做，若要在耶和華面前帶著兵器出去打仗，
NUM|32|21|你們中間所有帶兵器的人都要在耶和華面前過 約旦河 ，直到耶和華把仇敵從他面前趕出去。
NUM|32|22|那地在耶和華面前被征服以後，你們方可回來。這樣，你們向耶和華和 以色列 才算為無罪，這地也必在耶和華面前歸你們為業。
NUM|32|23|倘若你們不這樣做，看哪，你們就得罪了耶和華，當知道你們的罪必找上你們。
NUM|32|24|如今你們可以為孩童建城，為羊群築圈，但你們口所講出來的話，必須實踐。」
NUM|32|25|迦得 子孫和 呂便 子孫對 摩西 說：「你的僕人們必照我主所吩咐的去做。
NUM|32|26|我們的孩子、妻子、牛羊和所有的牲畜都要留在 基列 的各城。
NUM|32|27|但你的僕人，凡能帶兵器上戰場的，都要照我主所說的話，在耶和華面前渡過去打仗。」
NUM|32|28|於是， 摩西 為他們吩咐 以利亞撒 祭司和 嫩 的兒子 約書亞 ，以及 以色列 人各支派父系的領袖。
NUM|32|29|摩西 對他們說：「 迦得 子孫和 呂便 子孫，凡帶兵器在耶和華面前去打仗的，若與你們一同渡過 約旦河 ，那地被你們征服以後，你們就要把 基列 地給他們為業。
NUM|32|30|倘若他們不帶兵器與你們一同渡過去，他們就要在 迦南 地你們中間得產業。」
NUM|32|31|迦得 子孫和 呂便 子孫回答說：「耶和華怎樣吩咐僕人，我們就必照樣做。
NUM|32|32|我們自己必帶著兵器，在耶和華面前渡過去，進入 迦南 地，好使我們在 約旦河 這邊得到我們的產業。」
NUM|32|33|摩西 把 亞摩利 王 西宏 的國和 巴珊 王 噩 的國，就是他們的國土和周圍的城鎮，都給了 迦得 子孫和 呂便 子孫，以及 約瑟 的兒子 瑪拿西 半個支派。
NUM|32|34|迦得 子孫建造了 底本 、 亞他錄 、 亞羅珥 、
NUM|32|35|亞他錄‧朔反 、 雅謝 、 約比哈 、
NUM|32|36|伯‧寧拉 、 伯‧哈蘭 ，都是堅固城，並築有羊圈。
NUM|32|37|呂便 子孫建造了 希實本 、 以利亞利 、 基列亭 、
NUM|32|38|尼波 、 巴力‧免 （名字是改了的）、 西比瑪 ；他們給建造的城另起別名。
NUM|32|39|瑪拿西 的兒子 瑪吉 的子孫往 基列 去，佔了那地，趕出那裏的 亞摩利 人。
NUM|32|40|摩西 把 基列 賜給 瑪拿西 的兒子 瑪吉 ，他就住在那裏。
NUM|32|41|瑪拿西 的子孫 睚珥 佔了 基列 的城鎮，就稱這些城鎮為 哈倭特‧睚珥 。
NUM|32|42|挪巴 佔了 基納 和 基納 的鄉鎮，就照自己的名字稱 基納 為 挪巴 。
NUM|33|1|這是 以色列 人按著隊伍，在 摩西 、 亞倫 的手下，出 埃及 地的行程。
NUM|33|2|摩西 遵照耶和華的指示記錄他們每段行程的起點，這些行程的起點如下：
NUM|33|3|第一個月，就是正月十五日，逾越的第二天，他們從 蘭塞 起行，在所有 埃及 人的眼前抬起頭 來出去了。
NUM|33|4|那時， 埃及 人正埋葬他們的長子，就是耶和華在他們中間所擊殺的；耶和華也懲治了他們的眾神明。
NUM|33|5|以色列 人從 蘭塞 起行，安營在 疏割 。
NUM|33|6|從 疏割 起行，安營在曠野邊上的 以倘 。
NUM|33|7|從 以倘 起行，轉向 巴力‧洗分 對面的 比‧哈希錄 ，安營在 密奪 。
NUM|33|8|從 比‧哈希錄 起行，經過海，進入曠野，在 以倘 的曠野走了三天的路程，就安營在 瑪拉 。
NUM|33|9|從 瑪拉 起行，來到 以琳 ， 以琳 有十二股水泉，七十棵棕樹，就安營在那裏。
NUM|33|10|從 以琳 起行，安營在 紅海 邊。
NUM|33|11|從 紅海 邊起行，安營在 汛 的曠野。
NUM|33|12|從 汛 的曠野起行，安營在 脫加 。
NUM|33|13|從 脫加 起行，安營在 亞錄 。
NUM|33|14|從 亞錄 起行，安營在 利非訂 ；在那裏，百姓沒有水喝。
NUM|33|15|從 利非訂 起行，安營在 西奈 的曠野。
NUM|33|16|從 西奈 的曠野起行，安營在 基博羅‧哈他瓦 。
NUM|33|17|從 基博羅‧哈他瓦 起行，安營在 哈洗錄 。
NUM|33|18|從 哈洗錄 起行，安營在 利提瑪 。
NUM|33|19|從 利提瑪 起行，安營在 臨門‧帕烈 。
NUM|33|20|從 臨門‧帕烈 起行，安營在 立拿 。
NUM|33|21|從 立拿 起行，安營在 勒撒 。
NUM|33|22|從 勒撒 起行，安營在 基希拉他 。
NUM|33|23|從 基希拉他 起行，安營在 沙斐山 。
NUM|33|24|從 沙斐山 起行，安營在 哈拉大 。
NUM|33|25|從 哈拉大 起行，安營在 瑪吉希錄 。
NUM|33|26|從 瑪吉希錄 起行，安營在 他哈 。
NUM|33|27|從 他哈 起行，安營在 他拉 。
NUM|33|28|從 他拉 起行，安營在 密加 。
NUM|33|29|從 密加 起行，安營在 哈摩拿 。
NUM|33|30|從 哈摩拿 起行，安營在 摩西錄 。
NUM|33|31|從 摩西錄 起行，安營在 比尼‧亞干 。
NUM|33|32|從 比尼‧亞干 起行，安營在 曷‧哈及甲 。
NUM|33|33|從 曷‧哈及甲 起行，安營在 約巴他 。
NUM|33|34|從 約巴他 起行，安營在 阿博拿 。
NUM|33|35|從 阿博拿 起行，安營在 以旬‧迦別 。
NUM|33|36|從 以旬‧迦別 起行，安營在 尋 的曠野，就是 加低斯 。
NUM|33|37|從 加低斯 起行，安營在 以東 地邊界的 何珥山 。
NUM|33|38|以色列 人出 埃及 地後四十年，五月初一， 亞倫 祭司遵照耶和華的指示，上 何珥山 ，死在那裏。
NUM|33|39|亞倫 死在 何珥山 的時候一百二十三歲。
NUM|33|40|住在 迦南 地 尼革夫 的 迦南 人 亞拉得 王聽說 以色列 人來了。
NUM|33|41|以色列 人從 何珥山 起行，安營在 撒摩拿 。
NUM|33|42|從 撒摩拿 起行，安營在 普嫩 。
NUM|33|43|從 普嫩 起行，安營在 阿伯 。
NUM|33|44|從 阿伯 起行，安營在 摩押 境內的 以耶‧亞巴琳 。
NUM|33|45|從 以耶‧亞巴琳 起行，安營在 底本‧迦得 。
NUM|33|46|從 底本‧迦得 起行，安營在 亞門‧低比拉太音 。
NUM|33|47|從 亞門‧低比拉太音 起行，安營在 尼波 前面的 亞巴琳山脈 。
NUM|33|48|從 亞巴琳山脈 起行，安營在 約旦河 邊， 耶利哥 對面的 摩押 平原。
NUM|33|49|他們在 摩押 平原，沿著 約旦河 安營，從 伯‧耶施末 直到 亞伯‧什亭 。
NUM|33|50|耶和華在 約旦河 邊， 耶利哥 對面的 摩押 平原吩咐 摩西 說：
NUM|33|51|「你要吩咐 以色列 人說：你們過 約旦河 進 迦南 地的時候，
NUM|33|52|要從你們面前趕出那地所有的居民，摧毀他們一切的石像和鑄成的偶像，也要拆毀他們一切的丘壇。
NUM|33|53|你們要佔領那地，住在那裏，因我已把那地賜給你們為業。
NUM|33|54|你們要按照宗族抽籤，承受土地：人多的要多給他們產業；人少的要少給他們產業。抽到何地給何人，那地就屬於他。你們要按照父系的支派承受產業。
NUM|33|55|倘若你們不把那地的居民從你們面前趕出去，那留下的居民就必成為你們眼中的刺，肋下的荊棘，也必在你們所住的地上擾亂你們；
NUM|33|56|我想要怎樣待他們，也必照樣待你們。」
NUM|34|1|耶和華吩咐 摩西 說：
NUM|34|2|「你要吩咐 以色列 人，對他們說：你們到了 迦南 地，這就是歸你們為業的地， 迦南 地和它四周的邊界：
NUM|34|3|你們的南邊是從 尋 的曠野起，沿著 以東 的邊界；南邊的地界從 鹽海 東邊開始，
NUM|34|4|繞過 亞克拉濱 斜坡的南邊，經過 尋 ，直通到 加低斯‧巴尼亞 的南邊，又通到 哈薩‧亞達 ，經過 押們 ，
NUM|34|5|從 押們 轉向 埃及 溪谷，直通到海。
NUM|34|6|「你們西邊的地界要以 大海 為邊界；這就是你們西邊的地界。
NUM|34|7|「你們北邊的地界要從 大海 開始劃界，直到 何珥山 ，
NUM|34|8|從 何珥山 劃到 哈馬口 ，直通到 西達達 ，
NUM|34|9|又通到 西斐崙 ，直達 哈薩‧以難 。這就是你們北邊的地界。
NUM|34|10|「東邊的地界，你們要從 哈薩‧以難 開始劃界，直到 示番 ，
NUM|34|11|這地界要從 示番 下到 亞延 東邊的 利比拉 ，這地界要下延到 基尼烈海 的東邊，
NUM|34|12|這地界又下到 約旦河 ，直通到 鹽海 。這就是你們的地和它四圍的邊界。」
NUM|34|13|摩西 吩咐 以色列 人說：「這就是耶和華吩咐抽籤給九個半支派承受為業的地。
NUM|34|14|因為 呂便 子孫的支派按著父家、 迦得 子孫的支派按著父家，和 瑪拿西 半個支派已經得到了他們的產業：
NUM|34|15|這兩個半支派已經在 耶利哥 對面， 約旦河 東邊，向日出的方向承受了產業。」
NUM|34|16|耶和華吩咐 摩西 說：
NUM|34|17|「這是為你們分地為業的人的名字： 以利亞撒 祭司和 嫩 的兒子 約書亞 。
NUM|34|18|你要從每個支派中選一個領袖來分配產業。
NUM|34|19|這些人的名字如下： 猶大 支派， 耶孚尼 的兒子 迦勒 。
NUM|34|20|西緬 子孫的支派， 亞米忽 的兒子 示母利 。
NUM|34|21|便雅憫 支派， 基斯倫 的兒子 以利達 。
NUM|34|22|但 子孫支派的領袖， 約利 的兒子 布基 。
NUM|34|23|約瑟 的子孫， 瑪拿西 子孫支派的領袖： 以弗 的兒子 漢尼業 。
NUM|34|24|以法蓮 子孫支派的領袖： 拾弗但 的兒子 基摩利 。
NUM|34|25|西布倫 子孫支派的領袖： 帕納 的兒子 以利撒番 。
NUM|34|26|以薩迦 子孫支派的領袖： 阿散 的兒子 帕鐵 。
NUM|34|27|亞設 子孫支派的領袖： 示羅米 的兒子 亞希忽 。
NUM|34|28|拿弗他利 子孫支派的領袖： 亞米忽 的兒子 比大黑 。」
NUM|34|29|這些就是耶和華所吩咐，在 迦南 地為 以色列 人分產業的人。
NUM|35|1|耶和華在 約旦河 邊， 耶利哥 對面的 摩押 平原吩咐 摩西 說：
NUM|35|2|「你吩咐 以色列 人，要從所得為業的地中把一些城給 利未 人居住，也要把這些城四圍的郊野給 利未 人。
NUM|35|3|這些城鎮要歸他們居住，郊外可以給他們牧放牛羊、牲畜和所有的動物。
NUM|35|4|你們給 利未 人城的郊外，要從城牆量起，四圍往外量一千肘。
NUM|35|5|你們要往東量二千肘，往南量二千肘，往西量二千肘，往北量二千肘為邊界，以城為中心；這城鎮的郊外要歸給他們。」
NUM|35|6|「你們給 利未 人的城鎮中，要設立六座逃城，讓誤殺人的可以逃到那裏。此外還要給他們四十二座城。
NUM|35|7|所以，給 利未 人的城一共有四十八座，連同城的郊外都給他們。
NUM|35|8|從 以色列 人所得的產業中給 利未 人的這些城鎮，多的要多給，少的要少給；各支派要按照所承受為業之地的多少把城鎮給 利未 人。」
NUM|35|9|耶和華吩咐 摩西 說：
NUM|35|10|「你要吩咐 以色列 人，對他們說：你們過了 約旦河 ，進入 迦南 地，
NUM|35|11|要指定幾座城，作為你們的逃城，使誤殺人的可以逃到那裏。
NUM|35|12|這些城要作為逃避報仇者的城，使誤殺人的不至於死，等他站在會眾面前受審判。
NUM|35|13|「你們指定的城，是要作你們的六座逃城。
NUM|35|14|約旦河 東指定三座， 迦南 地也指定三座，作為逃城。
NUM|35|15|這六座城要給 以色列 人和他們中間的外人，以及寄居者，作為逃城，讓誤殺人的可以逃到那裏。
NUM|35|16|「倘若人用鐵器打死人，他是故意殺人的；故意殺人的必被處死。
NUM|35|17|若用手中可以致命的石頭打死人，他是故意殺人的；故意殺人的必被處死。
NUM|35|18|若用手中可以致命的木器打死人，他是故意殺人的；故意殺人的必被處死。
NUM|35|19|報血仇者可以親自殺死那故意殺人的；他一找到兇手，就可以殺死他。
NUM|35|20|人若因怨恨把人推倒，或埋伏等著丟東西砸人，以至於死，
NUM|35|21|或因仇恨用手打死人，打人的必被處死，他是故意殺人的；報血仇者一遇見兇手就可以殺死他。
NUM|35|22|「人若不是出於仇恨，把人推倒，或不是埋伏等著丟東西砸人，
NUM|35|23|或是在不注意的時候，用可以致命的石頭扔在人身上，以至於死，彼此沒有仇恨，也無意害對方，
NUM|35|24|會眾就要照著這些典章，在殺人者和報血仇者中間審判。
NUM|35|25|會眾要救這誤殺人的脫離報血仇者的手，送他回到他曾逃入的逃城那裏。他要住在城中，直到受聖膏的大祭司去世。
NUM|35|26|但誤殺人的，無論甚麼時候，若離開了他所逃入的逃城邊界，
NUM|35|27|報血仇者在逃城邊界外遇見他，把兇手殺了，報血仇者就沒有流人血之罪。
NUM|35|28|因為誤殺人的應該住在逃城裏，直到大祭司去世。大祭司去世以後，誤殺人的才可以回到他所得為業之地。
NUM|35|29|在你們一切的住處，這些都要作為你們世世代代的律例典章。
NUM|35|30|「無論誰殺了人，必須憑幾個證人的口，才可把那故意殺人的處死；只憑一個證人，不足以判人死。
NUM|35|31|那犯死罪的殺人犯，你們不可收贖價來代替他的命；他必須被處死。
NUM|35|32|那逃到逃城的人，你們不可向他收贖價，使他在大祭司未死以先回本地居住。
NUM|35|33|這樣，你們就不會污穢所住之地，因為血能使地污穢；若有血流在地上，除非流那殺人者的血，否則那地就不得潔淨。
NUM|35|34|你們不可玷污所住之地，就是我住在當中的地，因為我－耶和華住在 以色列 人中間。」
NUM|36|1|約瑟 子孫的宗族， 瑪拿西 的孫子， 瑪吉 的兒子 基列 ，他父系宗族的領袖來到 摩西 和作領袖的 以色列 眾父系家長面前，說：
NUM|36|2|「耶和華曾吩咐我主抽籤分地給 以色列 人為業，我主也遵照耶和華的吩咐，把我們兄弟 西羅非哈 的產業給他的女兒。
NUM|36|3|她們若嫁給 以色列 別個支派的人，必拿走我們祖宗所遺留的產業，加在她們丈夫支派的產業上。這樣，我們抽籤所得的產業就要減少了。
NUM|36|4|到了 以色列 人的禧年，她們的產業就必加在她們丈夫支派的產業上。這樣，我們祖宗支派的產業就要減少了。」
NUM|36|5|摩西 照耶和華的指示吩咐 以色列 人說：「 約瑟 子孫支派的人說得有理。
NUM|36|6|關於 西羅非哈 的女兒們，這是耶和華吩咐的話說：『她們可以隨意嫁人，只是必須嫁給同宗，她們父親支派的人。
NUM|36|7|這樣， 以色列 人的產業就不會從這支派轉到另一個支派，因為 以色列 人要各自守住祖宗支派的產業。
NUM|36|8|凡在 以色列 支派中得了產業的女兒，必須嫁給同宗，她們父親支派的人，好使 以色列 人各自承受他們祖宗的產業。
NUM|36|9|產業不可從一個支派轉到另一個支派，因為 以色列 支派的人要各自守住自己的產業。』」
NUM|36|10|耶和華怎樣吩咐 摩西 ， 西羅非哈 的女兒就照樣做。
NUM|36|11|西羅非哈 的女兒 瑪拉 、 得撒 、 曷拉 、 密迦 、 挪阿 都嫁給她們叔伯的兒子。
NUM|36|12|她們嫁給了 約瑟 兒子 瑪拿西 子孫宗族的人；她們的產業保留在同宗，她們父親的支派中。
NUM|36|13|這是耶和華在 約旦河 邊， 耶利哥 對面的 摩押 平原，藉著 摩西 吩咐 以色列 人的命令和典章。
DEUT|1|1|以下是 摩西 在 約旦河 東的曠野， 疏弗 對面的 亞拉巴 ，就是在 巴蘭 、 陀弗 、 拉班 、 哈洗錄 、 底撒哈 之間，向 以色列 眾人所說的話。
DEUT|1|2|從 何烈山 經過 西珥山 到 加低斯‧巴尼亞 要十一天的路程。
DEUT|1|3|第四十年十一月初一， 摩西 照耶和華所吩咐他一切有關 以色列 人的話，都告訴他們。
DEUT|1|4|那時，他已經擊敗了住 希實本 的 亞摩利 王 西宏 和住 亞斯她錄 、 以得來 的 巴珊 王 噩 。
DEUT|1|5|摩西 在 約旦河 東的 摩押 地講解這律法，說：
DEUT|1|6|「耶和華－我們的上帝在 何烈山 吩咐我們說：你們住在這山上已經夠久了。
DEUT|1|7|要起行，轉到 亞摩利 人的山區和附近的地區，就是 亞拉巴 、山區、 謝非拉 、 尼革夫 、沿海一帶， 迦南 人的地和 黎巴嫩 ，直到 大河 ，就是 幼發拉底河 。
DEUT|1|8|看，我將這地擺在你們面前。你們要進去得這地，就是耶和華向你們列祖 亞伯拉罕 、 以撒 、 雅各 起誓要賜給他們和他們後裔為業之地。」
DEUT|1|9|「那時，我對你們說：『我獨自一人無法承擔你們的事。
DEUT|1|10|耶和華－你們的上帝使你們增多。看哪，你們今日好像天上的星那樣多。
DEUT|1|11|惟願耶和華－你們列祖的上帝使你們更增加千倍，照他所應許你們的賜福給你們。
DEUT|1|12|但你們的擔子，你們的重任，以及你們的爭訟，我獨自一人怎能承擔呢？
DEUT|1|13|你們要按著各支派選出有智慧、明辨是非、為人所知的人來，我就立他們為你們的領袖。』
DEUT|1|14|你們回答我說：『你說要做的事很好！』
DEUT|1|15|我就將你們各支派的領袖，就是有智慧、為人所知的人，立他們為領袖，作你們各支派的千夫長、百夫長、五十夫長、十夫長等官長，來管理你們。
DEUT|1|16|「當時，我吩咐你們的審判官說：『你們聽訟，無論是弟兄之間的訴訟，或與寄居者之間的訴訟，都要秉公判斷。
DEUT|1|17|審判的時候不可看人的情面；無論大小，你們都要聽訟。不可因人而懼怕，因為審判是上帝的事。你們當中若有難斷的案件，可以呈到我這裏，讓我來聽訟。』
DEUT|1|18|那時，我已經把你們所當做的事都吩咐你們了。」
DEUT|1|19|「我們照著耶和華－我們上帝所吩咐的，從 何烈山 起行，經過你們所看見那一切大而可怕的曠野，往 亞摩利 人的山區去，到了 加低斯‧巴尼亞 。
DEUT|1|20|我對你們說：『你們已經到了耶和華－我們上帝所賜給我們的 亞摩利 人之山區。
DEUT|1|21|看，耶和華－你的上帝已將那地擺在你面前，你要照耶和華－你列祖的上帝所說的，上去得那地為業。不要懼怕，也不要驚惶。』
DEUT|1|22|你們都來到我這裏，說：『讓我們先派人去，為我們窺探那地，把我們上去該走的路線和該進的城鎮回報我們。』
DEUT|1|23|這話我看為美，就從你們中間選取十二個人，每支派一人。
DEUT|1|24|於是他們起身上山區去，到 以實各谷 ，窺探那地。
DEUT|1|25|他們的手帶著那地的一些果子，下到我們這裏，回報我們說：『耶和華－我們的上帝所賜給我們的是美地。』
DEUT|1|26|「你們卻不肯上去，竟違背了耶和華─你們上帝的指示，
DEUT|1|27|在帳棚內發怨言說：『耶和華因為恨我們，所以將我們從 埃及 地領出來，要把我們交在 亞摩利 人的手中，除滅我們。
DEUT|1|28|我們上哪裏去呢？我們的弟兄使我們膽戰心驚 ，說那裏的百姓比我們又大又高 ，那裏的城鎮又大，城牆又堅固，如天一樣高，並且我們在那裏看見 亞衲 族人。』
DEUT|1|29|我就對你們說：『不要驚惶，也不要怕他們。
DEUT|1|30|在你們前面行的耶和華－你們的上帝必為你們爭戰，正如他在 埃及 ，在你們眼前為你們所做的一樣；
DEUT|1|31|並且你們在曠野所行的一切路上，也看見了耶和華─你們的上帝背著你們，如同人背自己的兒子一樣，直到你們來到這地方。』
DEUT|1|32|你們在這事上卻不信耶和華─你們的上帝。
DEUT|1|33|他一路行在你們前面，為你們尋找安營的地方；他夜間在火中，日間在雲中，指示你們當走的路。」
DEUT|1|34|「耶和華聽見你們的怨言，就發怒，起誓說：
DEUT|1|35|『這邪惡世代的人，一個也不得看見我起誓要賜給你們列祖的美地；
DEUT|1|36|惟有 耶孚尼 的兒子 迦勒 必得看見，並且我要將他所踏過的地賜給他和他的子孫，因為他專心跟從我。』
DEUT|1|37|耶和華也因你們的緣故向我發怒，說：『你也不得進入那地。
DEUT|1|38|那侍候你， 嫩 的兒子 約書亞 必得進入那地。你要勉勵他，因為他要使 以色列 承受那地為業。
DEUT|1|39|你們的孩子，你們說要成為擄物的，就是今日尚不知善惡的兒女，必進入那地。我要將那地賜給他們，他們必得為業。
DEUT|1|40|至於你們，要轉回，從 紅海 的路往曠野去。』
DEUT|1|41|「你們回答我說：『我們得罪了耶和華！現在我們願遵照耶和華─我們上帝一切所吩咐的上去爭戰。』於是你們各人帶著兵器，以為很容易就能上到山區去。
DEUT|1|42|耶和華對我說：『你對他們說：不要上去，也不要爭戰，因我不在你們中間，恐怕你們在仇敵面前被擊敗。』
DEUT|1|43|我就告訴了你們，你們卻不聽從，竟違背耶和華的指示，擅自上到山區去。
DEUT|1|44|住在那山區的 亞摩利 人像蜂群一樣出來迎擊你們，追趕你們，在 西珥 擊敗你們，直到 何珥瑪 。
DEUT|1|45|你們就回來，在耶和華面前哭泣；耶和華卻不聽你們的聲音，也不向你們側耳。
DEUT|1|46|你們照著所停留的日子，在 加低斯 停留了許多日子。」
DEUT|2|1|「我們轉回，從 紅海 的路往曠野去，正如耶和華所吩咐我的。我們在 西珥山 繞行了許多日子。
DEUT|2|2|耶和華對我說：
DEUT|2|3|『你們繞行這山已經夠久了，要轉向北方。
DEUT|2|4|你要吩咐百姓說：你們弟兄 以掃 的子孫住在 西珥 ，你們要經過他們的邊界。他們必懼怕你們，但你們要分外謹慎。
DEUT|2|5|不可向他們挑戰；他們的地，連腳掌可踏之處，我都不給你們，因我已將 西珥山 賜給 以掃 為業。
DEUT|2|6|你們要用錢向他們買糧吃，也要用錢向他們買水喝。
DEUT|2|7|因為耶和華─你的上帝在你手裏所做的一切事上已賜福給你。你走這大曠野，他都知道。這四十年，耶和華─你的上帝與你同在，因此你一無所缺。』
DEUT|2|8|「於是，我們經過我們弟兄 以掃 子孫所住的 西珥 ，從 亞拉巴 的路，經過 以拉他 、 以旬‧迦別 ，轉向 摩押 曠野的路去。
DEUT|2|9|耶和華對我說：『不可侵犯 摩押 ，也不可向他們挑戰。他們的地，我不賜給你為業，因我已將 亞珥 賜給 羅得 的子孫為業。』
DEUT|2|10|先前， 以米 人住在那裏，百姓又大又多，像 亞衲 人一樣高大。
DEUT|2|11|他們跟 亞衲 人一樣，也算是 利乏音 人，但 摩押 人卻稱他們為 以米 人。
DEUT|2|12|從前， 何利 人也住在 西珥 ，但 以掃 的子孫把他們除滅，佔領了他們的地，接續他們在那裏居住，如同 以色列 在耶和華賜給他們為業之地所做的一樣。
DEUT|2|13|『現在，起來，過 撒烈溪 ！』於是我們過了 撒烈溪 。
DEUT|2|14|從離開 加低斯‧巴尼亞 到渡過 撒烈溪 ，這段時期共三十八年，直到這一代的戰士都從營中滅盡，正如耶和華向他們所起的誓。
DEUT|2|15|耶和華的手也攻擊他們，將他們從營中除滅，直到滅盡。
DEUT|2|16|「百姓中所有的戰士滅盡死亡以後，
DEUT|2|17|耶和華吩咐我說：
DEUT|2|18|『你今日要經過 摩押 的邊界 亞珥 ，
DEUT|2|19|走到 亞捫 人之地。不可侵犯他們，也不可向他們挑戰。 亞捫 人的地，我不賜給你們為業，因我已將那地賜給 羅得 的子孫為業。』
DEUT|2|20|那地也算是 利乏音 人之地，因為先前 利乏音 人住在那裏， 亞捫 人稱他們為 散送冥 人。
DEUT|2|21|那裏的百姓又大又多，像 亞衲 人一樣高大，但耶和華從 亞捫 人面前除滅他們， 亞捫 人就佔領他們的地，接續他們在那裏居住。
DEUT|2|22|這正如耶和華從前為住在 西珥 的 以掃 子孫，將 何利 人從他們面前除滅，使他們得了 何利 人的地，接續他們在那裏居住，直到今日一樣。
DEUT|2|23|亞衛 人先前住在鄉村直到 迦薩 ；從 迦斐託 出來的 迦斐託 人將 亞衛 人除滅，接續他們在那裏居住。
DEUT|2|24|你們起來往前去，過 亞嫩谷 。看哪，我已將 亞摩利 人 希實本 王 西宏 和他的地交在你手中，你要開始去得他的地為業，向他挑戰。
DEUT|2|25|從今日起，我要讓天下萬民因你驚慌懼怕，聽見你的名聲，就因你發顫傷慟。」
DEUT|2|26|「我從 基底莫 的曠野派遣使者到 希實本 王 西宏 那裏，用和平的話說：
DEUT|2|27|『求你讓我穿越你的地，我走路的時候，只走大路，不偏左右。
DEUT|2|28|你可以賣糧給我吃，賣水給我喝；只要讓我步行過去，
DEUT|2|29|就如住在 西珥 的 以掃 子孫和住在 亞珥 的 摩押 人待我一樣，等我過了 約旦河 ，進入耶和華－我們上帝所賜給我們的地。』
DEUT|2|30|但 希實本 王 西宏 不肯讓我們從他那裏經過，因為耶和華－你的上帝使他性情頑梗，內心剛硬，為要把他交在你手中，像今日一樣。
DEUT|2|31|耶和華對我說：『看，我已開始把 西宏 和他的地交給你了，你要開始得他的地為業。』
DEUT|2|32|「 西宏 和他的眾百姓出來迎擊我們，在 雅雜 與我們交戰。
DEUT|2|33|耶和華－我們的上帝把他交給我們，我們就殺了他和他的眾兒子，以及他所有的百姓。
DEUT|2|34|那時，我們奪了他一切的城鎮，毀滅各城的男人、女人、孩子，沒有留下一個倖存者。
DEUT|2|35|只有牲畜和所奪各城的財物，我們都取為自己的掠物。
DEUT|2|36|從 亞嫩谷 旁的 亞羅珥 和谷中的城，直到 基列 ，沒有一座城是高得我們不能攻取的；耶和華－我們的上帝把它們全都交給我們了。
DEUT|2|37|只有 亞捫 人之地， 雅博河 沿岸，以及山區的城鎮，你沒有挨近，這全是耶和華－我們上帝所吩咐的。」
DEUT|3|1|「我們又轉回，朝 巴珊 的路上去。 巴珊 王 噩 和他的眾百姓出來迎擊我們，在 以得來 與我們交戰。
DEUT|3|2|耶和華對我說：『不要怕他！因我已把他和他的眾百姓，以及他的地，都交在你手中；你要待他像從前待住在 希實本 的 亞摩利 王 西宏 一樣。』
DEUT|3|3|於是耶和華－我們的上帝也把 巴珊 王 噩 和他的眾百姓都交在我們手中；我們殺了他，沒有給他留下一個倖存者。
DEUT|3|4|那時，我們奪了他一切的城鎮，共六十座，沒有一座城不被我們所奪，這是 亞珥歌伯 的全境， 巴珊 王 噩 的國度。
DEUT|3|5|這些堅固的城都有高的城牆，有門有閂，此外，還有許多無城牆的鄉村。
DEUT|3|6|我們把這些都毀滅了，像從前待 希實本 王 西宏 一樣，毀滅各城的男人、女人、孩子；
DEUT|3|7|只有一切牲畜和城中的財物，我們取為自己的掠物。
DEUT|3|8|那時，我們從兩個 亞摩利 王的手裏把 約旦河 東邊的地奪過來，從 亞嫩谷 直到 黑門山 ，
DEUT|3|9|這 黑門山 ， 西頓 人稱為 西連 ， 亞摩利 人稱為 示尼珥 。
DEUT|3|10|我們奪了平原的各城、 基列 全地、 巴珊 全地，直到 撒迦 和 以得來 ，都是 巴珊 王 噩 國內的城鎮。
DEUT|3|11|利乏音 人所剩下的只有 巴珊 王 噩 。看哪，他的床是鐵床，按照人肘的度量，長九肘，寬四肘，現今不是在 亞捫 人的 拉巴 嗎？」
DEUT|3|12|「那時，我們得了這地。從 亞嫩谷 旁的 亞羅珥 起，連同 基列 山區的一半和境內的城鎮，我都給了 呂便 人和 迦得 人。
DEUT|3|13|基列 其餘的地和 巴珊 全地，就是 噩 的國度，我給了 瑪拿西 半支派。 亞珥歌伯 全境就是 巴珊 全地，也稱為 利乏音 人之地。
DEUT|3|14|瑪拿西 的子孫 睚珥 佔領了 亞珥歌伯 全境，直到 基述 人和 瑪迦 人的邊界，就按自己的名字稱這些地，就是 巴珊 ，為 哈倭特‧睚珥 ，直到今日。
DEUT|3|15|我又將 基列 給了 瑪吉 。
DEUT|3|16|我給了 呂便 人和 迦得 人從 基列 到 亞嫩谷 ，以谷的中央為界，直到 亞捫 人邊界的 雅博河 ；
DEUT|3|17|還有 亞拉巴 和靠近 約旦河 之地，從 基尼烈 直到 亞拉巴海 ，就是 鹽海 ，以及 毗斯迦山 斜坡的山腳東邊之地。
DEUT|3|18|「那時，我吩咐你們說：『耶和華－你們的上帝已將這地賜給你們為業；你們所有的勇士都要帶著兵器，在你們的弟兄 以色列 人前面過去。
DEUT|3|19|但你們的妻子、孩子、牲畜，可以住在我所賜給你們的各城裏，我知道你們有許多牲畜。
DEUT|3|20|等到耶和華讓你們的弟兄像你們一樣，得享太平，他們在 約旦河 另一邊，也得了耶和華－你們的上帝所賜給他們的地，你們各人才可以回到我所賜給你們為業之地。』
DEUT|3|21|那時，我吩咐 約書亞 說：『你親眼看見了耶和華－你們的上帝向這兩個王一切所做的事，耶和華也必向你所要去的各國照樣做。
DEUT|3|22|不要怕他們，因為那為你們爭戰的是耶和華－你們的上帝。』」
DEUT|3|23|「那時，我懇求耶和華說：
DEUT|3|24|『主耶和華啊，你已開始將你的偉大和你大能的手顯給你僕人看。在天上，在地下，有甚麼神明能像你行事，像你有大能的作為呢？
DEUT|3|25|求你讓我過去，看 約旦河 另一邊的美地，就是那佳美的山區和 黎巴嫩 。』
DEUT|3|26|但耶和華因你們的緣故向我發怒，不應允我。耶和華對我說：『你夠了吧！不要再向我提這事。
DEUT|3|27|你上 毗斯迦山 頂去，向東、西、南、北舉目，用你的眼睛觀看，因為你必不能過這 約旦河 。
DEUT|3|28|你卻要吩咐 約書亞 ，勉勵他，使他壯膽，因為他必在這百姓前面過去，使他們承受你所要觀看之地。』
DEUT|3|29|於是我們停留在 伯‧毗珥 對面的谷中。」
DEUT|4|1|「現在， 以色列 啊，聽我所教導你們的律例典章，要遵行，好使你們存活，得以進入耶和華－你們列祖之上帝所賜給你們的地，承受為業。
DEUT|4|2|我吩咐你們的話，你們不可加添，也不可刪減，好叫你們遵守耶和華－你們上帝的命令，就是我所吩咐你們的。
DEUT|4|3|你們已親眼看見耶和華因 巴力‧毗珥 所做的。凡隨從 巴力‧毗珥 的人，耶和華－你的上帝都從你中間除滅了。
DEUT|4|4|只有你們這緊緊跟隨耶和華－你們上帝的人，今日全都存活。
DEUT|4|5|看，我照著耶和華－我的上帝所吩咐我的，將律例和典章教導你們，使你們在所要進去得為業的地上遵行。
DEUT|4|6|你們要謹守遵行；這就是你們在萬民眼前的智慧和聰明。他們聽見這一切律例，必說：『這大國的人真是有智慧，有聰明！』
DEUT|4|7|哪一大國有神明與他們相近，像耶和華－我們的上帝在我們求告他的時候與我們相近呢？
DEUT|4|8|哪一大國有這樣公義的律例典章，像我今日在你們面前所頒佈的這一切律法呢？
DEUT|4|9|「但你要謹慎，殷勤保守你的心靈，免得忘記你親眼所看見的事，又免得在你一生的年日這些事離開你的心，總要把它們傳給你的子子孫孫。
DEUT|4|10|你在 何烈山 站在耶和華－你上帝面前的那日，耶和華對我說：『你為我召集百姓，我要叫他們聽見我的話，使他們活在世上的日子，可以學習敬畏我，又可以教導他們的兒女。』
DEUT|4|11|那時，你們近前來，站在山下；山上有火燃燒，直沖天頂，並有黑暗、密雲、幽暗。
DEUT|4|12|耶和華從火焰中對你們說話，你們聽見說話的聲音，只有聲音，卻沒有看見形像。
DEUT|4|13|他將所吩咐你們當守的約指示你們，就是十條誡命 ，並將誡命寫在兩塊石版上。
DEUT|4|14|那時，耶和華吩咐我將律例典章教導你們，使你們在所要過去得為業的地上遵行。」
DEUT|4|15|「所以，你們為自己的緣故要分外謹慎；因為耶和華在 何烈山 ，從火中對你們說話的那日，你們沒有看見任何形像。
DEUT|4|16|惟恐你們的行為敗壞，為自己雕刻任何形狀的偶像，無論是男像或女像，
DEUT|4|17|或地上任何走獸的像，或任何飛在空中有翅膀的鳥的像，
DEUT|4|18|或地上任何爬行動物的像，或地底下任何水中魚的像。
DEUT|4|19|又恐怕你向天舉目，看見耶和華－你的上帝為天下萬民所擺列的日月星辰，就是天上的萬象，就被誘惑去敬拜它們，事奉它們。
DEUT|4|20|耶和華將你們從 埃及 帶領出來，脫離鐵爐，是要你們成為他產業的子民，像今日一樣。
DEUT|4|21|「耶和華又因你們的緣故向我發怒，起誓不容我過 約旦河 ，不讓我進入耶和華－你上帝所賜你為業的那美地。
DEUT|4|22|我只好死在這地，不能過 約旦河 ；但你們必過去得那美地。
DEUT|4|23|你們要謹慎，免得忘記耶和華－你們的上帝與你們所立的約，為自己雕刻任何形狀的偶像，就是耶和華－你上帝所禁止的，
DEUT|4|24|因為耶和華－你的上帝是吞滅的火，是忌邪 的上帝。
DEUT|4|25|「你們在那地住久了，生子生孫，若行為敗壞，為自己雕刻任何形狀的偶像，行耶和華－你上帝眼中看為惡的事，惹他發怒，
DEUT|4|26|我今日呼天喚地向你們作見證，你們在過 約旦河 得為業的地上必迅速滅亡！你們在那地的日子必不長久，必全然滅絕。
DEUT|4|27|耶和華必將你們分散在萬民中；在耶和華領你們到的列國中，你們剩下的人丁稀少。
DEUT|4|28|在那裏，你們必事奉人手所造的神明，它們是木頭，是石頭，不能看，不能聽，不能吃，不能聞。
DEUT|4|29|你們在那裏必尋求耶和華－你的上帝。你若盡心盡性尋求他，就必尋見。
DEUT|4|30|日後你在患難中，當這一切的事臨到你，你必歸回耶和華－你的上帝，聽從他的話。
DEUT|4|31|耶和華－你的上帝是有憐憫的上帝，他不撇下你，不滅絕你，也不忘記他起誓與你列祖所立的約。
DEUT|4|32|「你去問，在你先前的時代，自從上帝造人在地上以來，從天這邊到天那邊，曾有過或聽過這樣的大事嗎？
DEUT|4|33|有哪些百姓聽見上帝在火中說話的聲音，像你聽見了還能存活呢？
DEUT|4|34|上帝何曾為自己嘗試從別的國中領出一國的子民來，用考驗、神蹟、奇事、戰爭、大能的手、伸出來的膀臂和大可畏的事，像耶和華－你們的上帝在 埃及 ，在你們眼前為你們所做的一切事呢？
DEUT|4|35|這是要顯給你看，使你知道，惟有耶和華他是上帝，除他以外，再沒有別的了。
DEUT|4|36|他從天上使你聽見他的聲音，為要教導你，又在地上使你看見他的烈火，並且聽見他從火中所說的話。
DEUT|4|37|因為他愛你的列祖，揀選他們的後裔 ，親自用大能領你出了 埃及 ，
DEUT|4|38|要將比你強大的列國從你面前趕出，領你進去，把他們的地賜你為業，像今日一樣。
DEUT|4|39|所以，今日你要知道，也要記在心裏，天上地下惟有耶和華他是上帝，再沒有別的了。
DEUT|4|40|我今日吩咐你的律例誡命，你要遵守，使你和你的後裔可以得福，並使你的日子一直在耶和華－你上帝賜你的地上得以長久。」
DEUT|4|41|「那時， 摩西 在 約旦河 東邊，向日出的方向，指定三座城，
DEUT|4|42|使那素無仇恨、無意中殺了鄰舍的兇手，可以逃到這三座城中的一座，就得存活：
DEUT|4|43|屬 呂便 人的是曠野平坦之地的 比悉 ，屬 迦得 人的是 基列 的 拉末 ，屬 瑪拿西 人的是 巴珊 的 哥蘭 。」
DEUT|4|44|這是 摩西 在 以色列 人面前頒佈的律法。
DEUT|4|45|這些法度、律例、典章是 摩西 在 以色列 人出 埃及 後對他們說的，
DEUT|4|46|在 約旦河 東 伯毗珥 對面的谷中，在住 希實本 的 亞摩利 王 西宏 之地；這 西宏 是 摩西 和 以色列 人出 埃及 後所擊殺的。
DEUT|4|47|他們得了他的地，又得了 巴珊 王 噩 的地，就是兩個 亞摩利 王，在 約旦河 東，向日出方向的地：
DEUT|4|48|從 亞嫩谷 旁的 亞羅珥 ，直到 西雲山 ，就是 黑門山 ，
DEUT|4|49|還有 約旦河 東的整個 亞拉巴 ，向日出方向，直到 亞拉巴海 ，靠近 毗斯迦山 斜坡的山腳。
DEUT|5|1|摩西 召集 以色列 眾人，對他們說：「 以色列 啊，要聽我今日在你們耳中所吩咐的律例典章，要學習，謹守遵行。
DEUT|5|2|耶和華－我們的上帝在 何烈山 與我們立約。
DEUT|5|3|這約耶和華不是與我們列祖立的，而是與我們，就是今日在這裏還活著的人立的。
DEUT|5|4|耶和華在山上，從火中，面對面與你們說話。
DEUT|5|5|那時我站在耶和華和你們之間，要將耶和華的話傳給你們，因為你們懼怕那火，沒有上山。他說：
DEUT|5|6|「『我是耶和華－你的上帝，曾將你從 埃及 地為奴之家領出來。
DEUT|5|7|「『除了我以外，你不可有別的神。
DEUT|5|8|「『不可為自己雕刻偶像，也不可做甚麼形像，彷彿上天、下地和地底下水中的百物。
DEUT|5|9|不可跪拜那些像，也不可事奉它們，因為我耶和華－你的上帝是忌邪 的上帝。恨我的，我必懲罰他們的罪，自父及子，直到三、四代；
DEUT|5|10|愛我、守我誡命的，我必向他們施慈愛，直到千代。
DEUT|5|11|「『不可妄稱耶和華－你上帝的名，因為妄稱耶和華名的，耶和華必不以他為無罪。
DEUT|5|12|「『當守安息日為聖日，正如耶和華－你上帝所吩咐的。
DEUT|5|13|六日要勞碌做你一切的工，
DEUT|5|14|但第七日是向耶和華－你的上帝當守的安息日。這一日，你和你的兒女、僕婢、牛、驢、牲畜，以及你城裏寄居的客旅，都不可做任何的工，使你的僕婢可以和你一樣休息。
DEUT|5|15|你要記念你在 埃及 地作過奴僕，耶和華－你的上帝用大能的手和伸出來的膀臂領你從那裏出來。因此，耶和華－你的上帝吩咐你守安息日。
DEUT|5|16|「『當孝敬父母，正如耶和華－你上帝所吩咐的，使你得福，並使你的日子在耶和華－你上帝所賜給你的地上得以長久。
DEUT|5|17|「『不可殺人。
DEUT|5|18|「『不可姦淫。
DEUT|5|19|「『不可偷盜。
DEUT|5|20|「『不可做假見證陷害你的鄰舍。
DEUT|5|21|「『不可貪戀你鄰舍的妻子；也不可貪圖你鄰舍的房屋、田地、僕婢、牛驢，以及他一切所有的。』
DEUT|5|22|「這些話是耶和華在山上，從火焰、密雲、幽暗中，大聲吩咐你們全會眾的，再沒有加添別的話了。他把這些話寫在兩塊石版上，交給我。
DEUT|5|23|山被火焰燒著，你們聽見從黑暗中發出的聲音，那時，你們各支派的領袖和長老都挨近我。
DEUT|5|24|你們說：『看哪，耶和華－我們的上帝將他的榮耀和他的偉大顯給我們看，我們也聽見他從火中發出的聲音。今日我們看到上帝與人說話，人還活著。
DEUT|5|25|現在這大火將要吞滅我們，我們何必死呢？若再聽見耶和華我們上帝的聲音，我們就必死。
DEUT|5|26|凡血肉之軀，有誰像我們一樣，聽見了永生上帝從火中講話的聲音還能活著呢？
DEUT|5|27|求你近前去，聽耶和華－我們上帝所要說的一切話，將耶和華－我們上帝對你說的話都傳給我們，我們就聽從遵行。』
DEUT|5|28|「你們對我說的話，耶和華都聽見了。耶和華對我說：『這百姓對你說的話，我聽見了；他們所說的都對。
DEUT|5|29|惟願他們存這樣的心敬畏我，常遵守我一切的誡命，使他們和他們的子孫永遠得福。
DEUT|5|30|你去對他們說：你們回帳棚去吧！
DEUT|5|31|至於你，可以站在我這裏，我要將一切誡命、律例、典章傳給你。你要教導他們，使他們在我賜他們為業的地上遵行。』
DEUT|5|32|所以，你們要照耶和華－你們上帝所吩咐的謹守遵行，不可偏離左右。
DEUT|5|33|你們要走耶和華－你們的上帝所吩咐的一切道路，使你們可以存活得福，並使你們的日子在所要承受的地上得以長久。」
DEUT|6|1|「這是耶和華－你們的上帝所吩咐要教導你們的誡命、律例、典章，叫你們在所要過去得為業的地上遵行，
DEUT|6|2|好叫你和你的子孫在一生的日子都敬畏耶和華－你的上帝，謹守他的一切律例、誡命，就是我所吩咐你的，使你的日子得以長久。
DEUT|6|3|以色列 啊，你要聽，要謹守遵行，使你可以在那流奶與蜜之地得福，人數極其增多，正如耶和華－你列祖的上帝所應許你的。
DEUT|6|4|「 以色列 啊，你要聽！耶和華－我們的上帝是獨一的主 。
DEUT|6|5|你要盡心、盡性、盡力愛耶和華－你的上帝。
DEUT|6|6|我今日吩咐你的這些話都要記在心上，
DEUT|6|7|也要殷勤教導你的兒女。無論你坐在家裏，走在路上，躺下，起來，都要吟誦。
DEUT|6|8|要繫在手上作記號，戴在額上 作經匣 ；
DEUT|6|9|又要寫在你房屋的門框上和你的城門上。
DEUT|6|10|「耶和華－你的上帝必領你進他向你列祖 亞伯拉罕 、 以撒 、 雅各 起誓要給你的地。那裏有又大又美的城鎮，不是你建造的；
DEUT|6|11|有裝滿各樣美物的房屋，不是你裝滿的；有挖成的水井，不是你挖的；有葡萄園、橄欖園，不是你栽植的；你吃了而且飽足。
DEUT|6|12|你要謹慎，免得你忘記領你從 埃及 地為奴之家出來的耶和華。
DEUT|6|13|你要敬畏耶和華－你的上帝，事奉他，奉他的名起誓。
DEUT|6|14|不可隨從別神，就是你們四圍民族的眾神明，
DEUT|6|15|因為在你中間的耶和華－你的上帝是忌邪 的上帝，恐怕耶和華－你上帝的怒氣向你發作，把你從地上除滅。
DEUT|6|16|「你們不可試探耶和華－你們的上帝，像你們在 瑪撒 那樣試探他。
DEUT|6|17|要謹慎遵守耶和華－你們上帝的誡命，和他所吩咐的法度、律例。
DEUT|6|18|耶和華眼中看為正直和美善的事，你都要遵行，使你得福，可以進去得耶和華向你列祖起誓應許的美地，
DEUT|6|19|可以從你面前趕出你所有的仇敵，正如耶和華所說的。
DEUT|6|20|「日後，你的兒子問你說：『耶和華－我們上帝吩咐你們的法度、律例、典章是甚麼意思呢？』
DEUT|6|21|你要告訴你的兒子說：『我們在 埃及 作過法老的奴僕，耶和華用大能的手將我們從 埃及 領出來。
DEUT|6|22|在我們眼前，他施行重大可怕的神蹟奇事對付 埃及 、法老和他的全家。
DEUT|6|23|他將我們從那裏領出來，為要領我們進入他向我們列祖起誓應許之地，把這地賜給我們。
DEUT|6|24|耶和華又吩咐我們遵行這一切的律例，敬畏耶和華－我們的上帝，使我們一生得福，得以存活，像今日一樣。
DEUT|6|25|我們若照耶和華－我們上帝所吩咐的，在他面前謹守遵行這一切誡命，這就是我們的義了。』」
DEUT|7|1|「耶和華－你的上帝領你進入你要得為業之地，從你面前趕出許多國家，就是比你更強大的七個國家： 赫 人、 革迦撒 人、 亞摩利 人、 迦南 人、 比利洗 人、 希未 人、 耶布斯 人。
DEUT|7|2|當耶和華－你的上帝把他們交給你，你擊殺他們的時候，你要完全消滅他們，不可與他們立約，也不可憐惜他們。
DEUT|7|3|不可與他們結親；不可將你的女兒嫁給他的兒子，也不可叫你的兒子娶他的女兒。
DEUT|7|4|因為他必使你的兒女離棄我，去事奉別神，以致耶和華的怒氣向你們發作，迅速將你除滅。
DEUT|7|5|你們卻要這樣處置他們：拆毀他們的祭壇，打碎他們的柱像，砍斷他們的 亞舍拉 ，用火焚燒他們雕刻的偶像。
DEUT|7|6|「因為你是屬於耶和華－你上帝神聖的子民；耶和華－你的上帝從地面上的萬民中揀選你，作自己寶貴的子民。
DEUT|7|7|耶和華專愛你們，揀選你們，並非因你們人數比任何民族多，其實你們的人數在各民族中是最少的。
DEUT|7|8|因為耶和華愛你們，又因要遵守他向你們列祖所起的誓，耶和華就用大能的手領你們出來，救贖你脫離為奴之家，脫離 埃及 王法老的手。
DEUT|7|9|所以，你知道耶和華－你的上帝，他是上帝，是信實的上帝。他向愛他、守他誡命的人守約施慈愛，直到千代；
DEUT|7|10|向恨他的人，他必當面報應，消滅他們。凡恨他的，他必當面報應，絕不遲延。
DEUT|7|11|所以，你要謹守我今日所吩咐你的誡命、律例、典章，遵行它們。」
DEUT|7|12|「你們若聽從這些典章，謹守遵行，耶和華－你的上帝必照他向你列祖所起的誓，對你守約，施慈愛。
DEUT|7|13|他必愛你，賜福給你，使你人數增多，也必在他向你列祖起誓要給你的地上賜福給你身所生的，你地所產的，你的五穀、新酒和新的油，以及你的牛犢、羔羊。
DEUT|7|14|你必蒙福勝過萬民；你沒有不育的男人和不孕的女人，牲畜也沒有不生育的。
DEUT|7|15|耶和華必使一切的疾病遠離你；你所知道 埃及 各樣的惡疾，他不加在你身上，反要加在所有恨你的人身上。
DEUT|7|16|你要吞滅耶和華－你的上帝交給你的各民族，你的眼目不可顧惜他們。你也不可事奉他們的神明，因為這必成為你的圈套。
DEUT|7|17|「你若心裏說，這些國的人數比我多，我怎能趕出他們呢？
DEUT|7|18|你不必怕他們，要牢牢記住耶和華－你上帝向法老和 埃及 全地所行的事，
DEUT|7|19|你親眼見過的大考驗、神蹟、奇事、大能的手和伸出來的膀臂，都是耶和華－你上帝領你出來所施行的。耶和華－你的上帝也必照樣處置你所懼怕的各民族，
DEUT|7|20|並且耶和華－你的上帝必派瘟疫 攻擊他們，直到那剩下而躲起來的人都從你面前滅亡。
DEUT|7|21|不要因他們驚恐，因為耶和華－你的上帝在你中間是大而可畏的上帝。
DEUT|7|22|耶和華－你的上帝必將這些國從你面前漸漸趕出；你不可迅速把他們消滅，免得野地的走獸多起來危害你。
DEUT|7|23|耶和華－你的上帝必將他們交給你，大大擾亂他們，直到他們被除滅。
DEUT|7|24|他又要將他們的君王交在你手中，你必從天下除去他們的名；必無一人能在你面前站立得住，直到你把他們除滅了。
DEUT|7|25|你們要用火焚燒他們神明的雕刻偶像；不可貪愛偶像上的金銀，也不可私自收起來，免得你因此陷入圈套，因為這是耶和華－你上帝所憎惡的。
DEUT|7|26|你不可把可憎之物帶進你的家，否則，你就像它一樣成為當毀滅的。你要徹底憎恨它，極其厭惡它，因為這是當毀滅的。」
DEUT|8|1|「我今日所吩咐你的一切誡命，你們要謹守遵行，好使你們存活，人數增多，可以進去得耶和華向你們列祖起誓應許的那地。
DEUT|8|2|你要記得，這四十年耶和華─你的上帝在曠野一路引導你，是要磨煉你，考驗你，為要知道你的心如何，是否願意遵守他的誡命。
DEUT|8|3|他磨煉你，任你飢餓，將你和你列祖所不認識的嗎哪賜給你吃，使你知道，人活著，不是單靠食物，乃是靠耶和華口裏所出的一切話。
DEUT|8|4|這四十年，你身上的衣服沒有穿破，你的腳也沒有腫。
DEUT|8|5|你心裏要知道，耶和華─你的上帝管教你，像人管教兒女一樣。
DEUT|8|6|你要謹守耶和華─你上帝的誡命，遵行他的道，敬畏他。
DEUT|8|7|「耶和華─你的上帝必領你進入美地，那地有河流，有泉源和深淵的水從谷中和山上流出。
DEUT|8|8|那地有小麥、大麥、葡萄樹、無花果樹、石榴樹，那地也有橄欖油和蜂蜜。
DEUT|8|9|那地沒有缺乏，你在那裏有食物吃，一無所缺；那地的石頭是鐵，山中可以挖銅。
DEUT|8|10|你吃得飽足，要稱頌耶和華─你的上帝，因為他將那美地賜給你。」
DEUT|8|11|「你要謹慎，免得忘記耶和華─你的上帝，不守他的誡命、典章、律例，就是我今日吩咐你的。
DEUT|8|12|免得你吃得飽足，建造上好的房屋，住在其中，
DEUT|8|13|你的牛羊增多，你的金銀增多，你擁有的一切全都增多，
DEUT|8|14|於是你的心高傲，忘記耶和華─你的上帝。他曾將你從 埃及 地為奴之家領出來，
DEUT|8|15|曾引領你經過那大而可怕的曠野，有火蛇、蠍子、乾旱無水之地。他也曾為你使水從堅硬的磐石中流出來，
DEUT|8|16|又在曠野將你列祖所不認識的嗎哪賜給你吃，為要磨煉你，考驗你，終久使你享福。
DEUT|8|17|你心裏說：『這財富是我的力量、我手的能力得來的。』
DEUT|8|18|你要記得耶和華─你的上帝，因為得財富的能力是他給你的，為要堅守他向你列祖起誓所立的約，像今日一樣。
DEUT|8|19|你若忘記耶和華─你的上帝，隨從別神，事奉它們，敬拜它們，我今日警告你們，你們必定滅亡。
DEUT|8|20|耶和華在你們面前怎樣使列國滅亡，你們也必照樣滅亡，因為你們不聽從耶和華─你們上帝的話。」
DEUT|9|1|「 以色列 啊，你要聽！你今日要過 約旦河 ，進去佔領比你更強大的列國，那裏的城鎮又大，城牆又堅固，如天一樣高。
DEUT|9|2|那裏的百姓是 亞衲 族人，又高又壯，是你所知道的；你也聽說過：『誰能在 亞衲 族人面前站立得住呢？』
DEUT|9|3|你今日應當知道，耶和華─你的上帝在你前面渡過去，如同吞噬的火，要除滅他們，並要在你面前將他們制伏，使你可以趕出他們，速速消滅他們，正如耶和華向你所說的。
DEUT|9|4|「耶和華─你的上帝將他們從你面前趕出以後，你心裏不可說：『耶和華領我得這地是因我的義。』其實，耶和華將這些國家從你面前趕出去是因他們的惡。
DEUT|9|5|你能進去得他們的地，並不是因你的義，也不是因你心裏正直，而是因這些國家的惡，耶和華─你的上帝才把他們從你面前趕出去，為了應驗耶和華向你列祖 亞伯拉罕 、 以撒 、 雅各 起誓應許的話。
DEUT|9|6|「你當知道，耶和華─你的上帝將這美地賜你為業，並不是因你的義；你本是硬著頸項的百姓。
DEUT|9|7|你要記得，不要忘記，你在曠野怎樣惹耶和華－你的上帝發怒。自從你出了 埃及 地的那日，直到你們來到這地方，你們常常悖逆耶和華。
DEUT|9|8|你們在 何烈山 惹耶和華發怒，耶和華對你們動怒，甚至要除滅你們。
DEUT|9|9|我上了山，要領受兩塊石版，就是耶和華與你們立約的版。那時我在山上住了四十晝夜，沒有吃飯，也沒有喝水。
DEUT|9|10|耶和華把那兩塊石版交給我，是上帝用指頭寫成的；版上是耶和華在大會的那一天，在山上從火中對你們所說的一切話。
DEUT|9|11|過了四十晝夜，耶和華把那兩塊石版，就是約版，交給我。
DEUT|9|12|耶和華對我說：『起來，趕快從這裏下去！因為你從 埃及 領出來的百姓已經敗壞了；他們這麼快偏離了我所吩咐的道，為自己鑄造偶像。』
DEUT|9|13|「耶和華對我說：『我看這百姓，看哪，他們是硬著頸項的百姓。
DEUT|9|14|你且由著我，我要除滅他們，從天下塗去他們的名，我要使你成為比他們更大更強的國。』
DEUT|9|15|於是我轉身下山，山上有火燃燒，兩塊約版在我雙手中。
DEUT|9|16|我觀看，看哪，你們得罪了耶和華－你們的上帝，為自己鑄成了一頭牛犢，迅速偏離了耶和華所吩咐你們的道，
DEUT|9|17|我拿著那兩塊石版，從我雙手中扔出去，在你們眼前把它們摔碎了。
DEUT|9|18|因為你們所犯的一切罪，做了耶和華眼中看為惡的事，惹他發怒，我就像從前一樣俯伏在耶和華面前四十晝夜，沒有吃飯，沒有喝水。
DEUT|9|19|我很害怕，因為耶和華向你們大發烈怒，要除滅你們。但那一次耶和華又應允了我。
DEUT|9|20|耶和華也向 亞倫 非常生氣，甚至要除滅他；那時我也為 亞倫 祈禱。
DEUT|9|21|我把那使你們犯罪所鑄的牛犢拿來，用火焚燒，搗碎後再磨成粉末，好像灰塵。我把這灰塵撒在從山上流下來的溪水中。
DEUT|9|22|「你們在 他備拉 、 瑪撒 、 基博羅‧哈他瓦 又惹耶和華發怒。
DEUT|9|23|耶和華叫你們離開 加低斯‧巴尼亞 ，說：『你們上去得我所賜給你們的地。』那時，你們違背了耶和華－你們上帝的指示，不信服他，不聽從他的話。
DEUT|9|24|自從我認識你們的日子以來，你們常常悖逆耶和華。
DEUT|9|25|「我因耶和華說要除滅你們，就在耶和華面前俯伏四十晝夜，像我以前俯伏一樣。
DEUT|9|26|我向耶和華祈禱，說：『主耶和華啊，求你不要滅絕你的百姓，你的產業。他們是你用大能救贖，用你強有力的手從 埃及 領出來的。
DEUT|9|27|求你記念你的僕人 亞伯拉罕 、 以撒 、 雅各 ，不看這百姓的頑梗、邪惡、罪愆，
DEUT|9|28|免得你領我們出來的那地之人說：耶和華因為不能將這百姓領進他所應許之地，又因恨他們，所以領他們出去，要在曠野殺他們。
DEUT|9|29|其實他們是你的百姓，你的產業，是你用大能和伸出的膀臂領出來的。』」
DEUT|10|1|「那時，耶和華對我說：『你要鑿出兩塊石版，和先前的一樣，上山到我這裏來。你也要造一個木櫃。
DEUT|10|2|我要把你先前摔碎的版上所寫的字，寫在這版上；你要把這版放在櫃裏。』
DEUT|10|3|於是我用金合歡木造了一個櫃子，又鑿出兩塊石版，和先前的一樣。我手裏拿著這兩塊版上山。
DEUT|10|4|耶和華將那大會之日、在山上從火中所吩咐你們的十條誡命，照先前所寫的寫在這版上。耶和華把它們交給我。
DEUT|10|5|我轉身下山，將這版放在我所造的櫃裏，現今這版還在那裏，正如耶和華所吩咐我的。
DEUT|10|6|（ 以色列 人從 比羅比尼‧亞干 起行，來到 摩西拉 ， 亞倫 死在那裏，就葬在那裏。他的兒子 以利亞撒 接續他擔任祭司的職分。
DEUT|10|7|他們從那裏起行，來到 谷歌大 ，又從 谷歌大 來到 約巴他 ，有溪水之地。
DEUT|10|8|那時，耶和華將 利未 支派分別出來，抬耶和華的約櫃，又侍立在耶和華面前事奉他，奉他的名祝福，直到今日。
DEUT|10|9|因此， 利未 沒有像他的弟兄有產業，耶和華是他的產業，正如耶和華－你上帝所應許他的。）
DEUT|10|10|「我又像先前一樣在山上停留了四十晝夜。這一次耶和華也應允我，不將你滅絕。
DEUT|10|11|耶和華對我說：『起來，走在百姓前面，領他們進去得我向他們列祖起誓要給他們的地。』」
DEUT|10|12|「 以色列 啊，現在耶和華－你的上帝向你要的是甚麼呢？只要你敬畏耶和華－你的上帝，遵行他一切的道，愛他，盡心盡性事奉耶和華－你的上帝，
DEUT|10|13|遵守耶和華的誡命律例，就是我今日所吩咐你的，為要使你得福。
DEUT|10|14|看哪，天和天上的天，地和地上所有的，都屬耶和華－你的上帝。
DEUT|10|15|然而，耶和華專愛你的列祖，愛他們，從萬民中揀選你們，就是他們的後裔，像今日一樣。
DEUT|10|16|所以你們的心要受割禮，不可再硬著頸項。
DEUT|10|17|因為耶和華－你們的上帝是萬神之神，萬主之主，是偉大、強有力、可畏的上帝，不看人的情面，也不受賄賂。
DEUT|10|18|他為孤兒寡婦伸冤，愛護寄居的，賜給他衣食。
DEUT|10|19|所以你們要愛護寄居的，因為你們在 埃及 地也作過寄居的。
DEUT|10|20|你要敬畏耶和華－你的上帝，事奉他，緊緊跟隨他，奉他的名起誓。
DEUT|10|21|他是你當讚美的，是你的上帝，為你做了大而可畏的事，這些是你親眼見過的。
DEUT|10|22|你的列祖七十人下 埃及 ，現在耶和華－你的上帝卻使你如同天上的星那樣多。」
DEUT|11|1|「你要愛耶和華－你的上帝，天天遵守他的吩咐、律例、典章、誡命。
DEUT|11|2|今日你們應當知道，而不是你們的兒女，因為他們不知道，也沒有見過耶和華─你們上帝的管教、他的偉大、他大能的手和伸出來的膀臂，
DEUT|11|3|以及他在 埃及 向 埃及 王法老和其全地所行的神蹟奇事；
DEUT|11|4|他怎樣對待 埃及 的軍隊、馬和戰車，他們追趕你們的時候，耶和華怎樣用 紅海 的水淹沒他們，消滅了他們，直到今日；
DEUT|11|5|他在曠野怎樣待你們，直到你們來到這地方，
DEUT|11|6|以及他怎樣待 呂便 子孫， 以利押 的兒子 大坍 、 亞比蘭 ，地怎樣在 以色列 人中開了裂口，吞了他們和他們的家眷，帳棚，以及跟他們在一起所有活著的。
DEUT|11|7|惟有你們親眼見過耶和華所做的一切大事。」
DEUT|11|8|「所以，你們要遵守我今日所吩咐的一切誡命，使你們剛強，可以進去得你們所要得的那地，就是你們將過河到那裏要得的，
DEUT|11|9|也使你們的日子，在耶和華向你們列祖起誓要給他們和他們後裔的地上得以長久，那是流奶與蜜之地。
DEUT|11|10|你要進去得為業的那地，不像你出來的 埃及 地。在 埃及 ，你撒種後，要用腳澆灌，像澆灌菜園一樣。
DEUT|11|11|你們要過去得為業的那地乃是有山有谷、天上的雨水滋潤之地，
DEUT|11|12|是耶和華－你上帝所眷顧的地；從歲首到年終，耶和華－你上帝的眼目時常看顧那地。
DEUT|11|13|「你們若留心聽從我今日所吩咐你們的誡命，愛耶和華－你們的上帝，盡心盡性事奉他，
DEUT|11|14|我 必按時降下雨水在你們的地上，就是秋雨和春雨，使你們可以收藏五穀、新酒和新的油，
DEUT|11|15|也必使田野為你的牲畜長出草來；這樣，你必吃得飽足。
DEUT|11|16|你們要謹慎，免得心受誘惑，轉去事奉別神，敬拜它們，
DEUT|11|17|以致耶和華的怒氣向你們發作，使天封閉不下雨，使地不出產，使你們在耶和華所賜給你們的美地上速速滅亡。
DEUT|11|18|「你們要將我這些話存在心裏，留在意念中，繫在手上作記號，戴在額上 作經匣。
DEUT|11|19|你們也要將這些話教導你們的兒女，無論坐在家裏，行在路上，躺下，起來，都要講論，
DEUT|11|20|又要寫在房屋的門框上和你的城門上。
DEUT|11|21|這樣，你們和你們子孫的日子必在耶和華向你們列祖起誓要給他們的地上得以增多，如天地之長久。
DEUT|11|22|你們若留心謹守遵行我所吩咐這一切的誡命，愛耶和華－你們的上帝，遵行他一切的道，緊緊跟隨他，
DEUT|11|23|他必從你們面前趕出這一切國家，你們也要佔領比你們更大更強的國家。
DEUT|11|24|凡你們腳掌所踏之地都必歸於你們；從曠野到 黎巴嫩 ，從 幼發拉底 大河，直到西邊的海，都要成為你們的疆土。
DEUT|11|25|必無一人能在你們面前站立得住；耶和華－你們的上帝必照他所說的，使懼怕驚恐臨到你們所踏的全地。
DEUT|11|26|「看，我今日將祝福與詛咒都陳明在你們面前。
DEUT|11|27|你們若聽從耶和華─你們上帝的誡命，就是我今日所吩咐你們的，就必蒙福。
DEUT|11|28|你們若不聽從耶和華─你們上帝的誡命，偏離我今日所吩咐你們的道，去隨從你們所不認識的別神，就必受詛咒。
DEUT|11|29|當耶和華－你的上帝領你進入要得為業的那地，你就要在 基利心山 上宣佈祝福，在 以巴路山 上宣佈詛咒。
DEUT|11|30|這二座山豈不是在 約旦河 的那邊，日落的方向，在住 亞拉巴 的 迦南 人之地， 吉甲 的前面，靠近 摩利 橡樹嗎？
DEUT|11|31|你們過 約旦河 ，進去得耶和華－你們的上帝所賜你們為業之地；當你們佔領它，在那地居住的時候，
DEUT|11|32|你們要謹守遵行我今日在你們面前頒佈的一切律例典章。」
DEUT|12|1|「你們活在世上的日子，在耶和華─你列祖的上帝所賜你為業的地上，你們要謹守遵行這些律例典章：
DEUT|12|2|你們佔領的國家所事奉他們眾神明的地方，無論是在高山，在小山，在一切的青翠樹下，你們要徹底毀壞；
DEUT|12|3|要拆毀他們的祭壇，打碎他們的柱像，用火焚燒他們的 亞舍拉 ，砍斷他們神明的雕刻偶像，並要從那地方除去他們的名。
DEUT|12|4|你們不可那樣敬拜耶和華－你們的上帝。
DEUT|12|5|但耶和華－你們的上帝在你們各支派中選擇何處作為立他名的居所，你們就要到那裏求問，
DEUT|12|6|將你們的燔祭、祭物、十一奉獻、手中的舉祭、還願祭、甘心祭，以及牛群羊群中頭生的，都帶到那裏。
DEUT|12|7|在那裏，你們和你們的全家都可以在耶和華─你們上帝的面前吃，並且因你們手所做的一切蒙耶和華－你的上帝賜福而歡樂。
DEUT|12|8|你們不可做像我們今日在這裏所做的，各人行自己眼中看為正的一切事；
DEUT|12|9|因為你們現在還沒有進入耶和華－你上帝所賜你的安息，所給你的產業。
DEUT|12|10|你們過了 約旦河 ，住在耶和華─你們上帝給你們承受為業的地；他又使你們得享太平，不受四圍一切仇敵擾亂，使你們安然居住。
DEUT|12|11|那時你們要將我所吩咐你們的燔祭、祭物、十一奉獻、手中的舉祭，和向耶和華許願的一切上好的祭，都帶到耶和華─你們上帝所選擇立他名的居所。
DEUT|12|12|你們和兒女、僕婢，以及住在你們城裏，沒有與你們一起分得產業的 利未 人，都要在耶和華－你們的上帝面前歡樂。
DEUT|12|13|你要謹慎，不可在自己所看中的各處獻燔祭。
DEUT|12|14|惟獨耶和華從你的一個支派中所選擇的地方，你要在那裏獻燔祭，在那裏遵行我一切所吩咐你的。
DEUT|12|15|「然而，你在各城裏都可以照著耶和華－你上帝所賜給你的福分，隨心所欲宰牲吃肉；無論潔淨的人不潔淨的人都可以吃，就如吃羚羊和鹿的肉一樣。
DEUT|12|16|只是血，你不可吃，要把它倒在地上，如同倒水一樣。
DEUT|12|17|你的五穀、新酒和新油的十分之一，或是牛群羊群中頭生的，或是你的許願祭、甘心祭和手中的舉祭，都不可在你的城裏吃，
DEUT|12|18|必須在耶和華－你的上帝面前吃，在耶和華－你上帝所選擇的地方，你和兒女、僕婢，以及住在你城裏的 利未 人都可以吃，並要因你手所做的一切，在耶和華－你上帝面前歡樂。
DEUT|12|19|你要謹慎，在你所住的地上，你永不可離棄 利未 人。
DEUT|12|20|「耶和華－你的上帝照他的應許擴張你疆土的時候，你心裏想要吃肉，說：『我要吃肉』，就可以隨心所欲吃肉。
DEUT|12|21|耶和華－你上帝選擇立他名的地方若離你太遠，你可以照我所吩咐的，將耶和華賜給你的牛羊取些宰了，隨心所欲在你的城裏吃。
DEUT|12|22|其實，就如吃羚羊和鹿的肉一樣，你要這樣吃它，無論潔淨的人不潔淨的人都可以一起吃。
DEUT|12|23|但是你要堅定，不可吃血，因為血是生命；不可將生命與肉一起吃。
DEUT|12|24|你不可吃血，要把它倒在地上，如同倒水一樣。
DEUT|12|25|不可吃血，好讓你和你的子孫可以得福，因為你行了耶和華眼中看為正的事。
DEUT|12|26|只是你分別為聖的物和你所還的願，都要帶到耶和華所選擇的地方去。
DEUT|12|27|你的燔祭，連肉帶血，都要獻在耶和華－你上帝的壇上。祭物的血要倒在耶和華－你上帝的壇上；肉你可以吃。
DEUT|12|28|你要謹守聽從我所吩咐的一切話，好讓你和你的子孫可以永遠得福，因為你行耶和華－你上帝眼中看為善、看為正的事。」
DEUT|12|29|「耶和華－你上帝把你要進去趕出的列國從你面前剪除，並且你得了他們的地為業居住，
DEUT|12|30|那時你要謹慎，在他們從你面前被除滅之後，你不可受引誘隨從他們，也不可求問他們的神明，說：『這些國家怎樣事奉他們的神明，我也要照樣做。』
DEUT|12|31|你不可向耶和華－你的上帝這樣做，因為他們向他們的神明做了耶和華所憎恨、所厭惡的一切事，甚至將自己的兒女用火焚燒，獻給他們的神明。
DEUT|12|32|凡我所吩咐你們的事，你們都要謹守遵行，不可加添，也不可刪減。」
DEUT|13|1|「你中間若有先知或是做夢的人起來，向你顯神蹟奇事，
DEUT|13|2|他對你說的神蹟奇事應驗了，說：『我們去隨從別神，事奉它們吧。』那是你不認識的。
DEUT|13|3|你不可聽那先知或是那做夢之人的話，因為這是耶和華－你們的上帝考驗你們，要知道你們是否盡心盡性愛耶和華－你們的上帝。
DEUT|13|4|你們要順從耶和華－你們的上帝，敬畏他，謹守他的誡命，聽從他的話，事奉他，緊緊跟隨他。
DEUT|13|5|那先知或那做夢的人要被處死，因為他出言悖逆那領你們出 埃及 地、救贖你脫離為奴之家的耶和華－你們的上帝，要引誘你離開耶和華－你上帝吩咐你要行的道。這樣，你就把惡從你中間除掉。
DEUT|13|6|「你的同胞兄弟，或是你的兒女，或是你懷中的妻，或是如同自己性命的朋友，若暗中引誘你，說：『我們去事奉別神吧。』那是你和你列祖所不認識的，
DEUT|13|7|你四圍列國的神明，無論是離你近或離你遠，從地這邊到地那邊，
DEUT|13|8|你都不可附和他，也不要聽從他。你的眼不可顧惜他，不可憐憫他，也不可袒護他。
DEUT|13|9|你務必殺他；你先下手，然後眾百姓才下手，把他處死。
DEUT|13|10|要用石頭打死他，因為他想引誘你離開那領你出 埃及 地為奴之家的耶和華－你的上帝。
DEUT|13|11|全 以色列 都要聽見而害怕，不敢在你中間再行這樣的惡事了。
DEUT|13|12|「若你聽見人說，在耶和華－你上帝所賜給你居住的城鎮中的一座，
DEUT|13|13|有些無賴之徒從你中間出來，引誘本城的居民，說：『我們去事奉別神吧。』那是你們不認識的，
DEUT|13|14|你就要調查，探聽，細心詢問。看哪，是真的，確實有這可憎的事在你中間發生，
DEUT|13|15|你務必用刀殺那城裏的居民，把城裏所有的，連牲畜都用刀滅盡。
DEUT|13|16|你要把從城裏所奪取的一切財物堆在廣場中，用火將那城和其中奪取的一切財物全燒給耶和華－你的上帝。那城要永遠成為廢墟，不得重建。
DEUT|13|17|那當毀滅的物一點都不可黏你的手，好讓耶和華轉回，不向你發烈怒，卻恩待你，憐憫你，照他向你列祖所起的誓使你人數增多；
DEUT|13|18|因為你聽從耶和華－你上帝的話，遵守我今日所吩咐你的一切誡命，行耶和華－你上帝眼中看為正的事。」
DEUT|14|1|「你們是耶和華─你們上帝的兒女。不可為了死人割劃自己，也不可使額上 光禿；
DEUT|14|2|因為你是屬於耶和華－你上帝神聖的子民，耶和華從地面上的萬民中揀選了你，作自己寶貴的子民。」
DEUT|14|3|「凡可憎的物， 你都不可吃。
DEUT|14|4|可吃的牲畜是：牛、綿羊、山羊、
DEUT|14|5|鹿、羚、麃子、野山羊、瞪羚、羚羊、山綿羊。
DEUT|14|6|凡蹄分兩瓣，分趾蹄而又反芻食物的牲畜，你們都可以吃。
DEUT|14|7|但那反芻或分蹄之中不可吃的是：駱駝、兔子、石獾，雖然反芻卻不分蹄，對你們是不潔淨的；
DEUT|14|8|豬，雖然分蹄卻不反芻，對你們也是不潔淨的。牠們的肉，你們一點都不可吃；牠們的屍體，你們也不可摸。
DEUT|14|9|「水中可吃的是這些：凡有鰭有鱗的都可以吃；
DEUT|14|10|凡無鰭無鱗的都不可吃，對你們是不潔淨的。
DEUT|14|11|「凡潔淨的鳥，你們都可以吃。
DEUT|14|12|不可吃的是：鵰、狗頭鵰、紅頭鵰、
DEUT|14|13|鸇、小鷹、鷂鷹的類群，
DEUT|14|14|各種烏鴉的類群、
DEUT|14|15|鴕鳥、夜鷹、魚鷹、鷹的類群、
DEUT|14|16|鴞鳥、貓頭鷹、角鴟、
DEUT|14|17|鵜鶘、禿鵰、鸕鶿、
DEUT|14|18|鸛、鷺鷥的類群、戴鵀與蝙蝠。
DEUT|14|19|凡有翅膀卻爬行的群聚動物對你們是不潔淨的，都不可吃。
DEUT|14|20|凡潔淨的鳥，你們都可以吃。
DEUT|14|21|「凡自然死去的動物，你們都不可吃，可以給城裏寄居的人吃，或賣給外人，因為你是屬於耶和華－你上帝神聖的子民。 「不可用母山羊的奶來煮牠的小山羊。」
DEUT|14|22|「每年，你務必從你播種的一切收成，田地所出產的，取十分之一獻上。
DEUT|14|23|要在耶和華－你上帝面前，就是他選擇那裏作為他名居所的地方，吃你所獻十分之一的五穀、新酒和新的油，以及牛群羊群中頭生的，好讓你天天學習敬畏耶和華－你的上帝。
DEUT|14|24|當耶和華－你的上帝賜福給你的時候，耶和華－你上帝選擇立他名的地方若離你太遠，路途太長，使你不能把這東西帶到那裏去，
DEUT|14|25|你可以把它換成銀子，把銀子包起來，拿在手中，往耶和華－你上帝所選擇的地方去。
DEUT|14|26|在那裏，你可以隨心所欲用銀子或買牛羊，或買清酒烈酒，或買任何你心所想的。你和你的全家要在耶和華－你上帝面前吃喝歡樂。
DEUT|14|27|「住在你城裏的 利未 人，你不可離棄他，因為他在你那裏沒有分得產業。
DEUT|14|28|每三年的最後一年，你要把那一年收成的十分之一取出來，積存在你的城中；
DEUT|14|29|那沒有與你一起分得產業的 利未 人，和城裏的寄居者，以及孤兒寡婦，都可以前來，吃得飽足，好讓耶和華－你的上帝在你手裏所做的一切事上賜福給你。」
DEUT|15|1|「每七年的最後一年，你要施行豁免。
DEUT|15|2|豁免的方式是這樣：凡債主要把手裏所借給鄰舍的全豁免，不可向鄰舍和弟兄追討，因為耶和華的豁免已經宣告了。
DEUT|15|3|你可以向外邦人追討；但你弟兄欠你的，無論是甚麼，你都要放手豁免。
DEUT|15|4|其實，在你中間不會有貧窮人；因為在耶和華－你上帝所賜你為業的地上，耶和華必大大賜福給你。
DEUT|15|5|只要你留心聽從耶和華－你上帝的話，謹守遵行我今日所吩咐你這一切的命令，
DEUT|15|6|因為耶和華－你的上帝會照他所應許你的賜福給你，你必借給許多國家，卻不需要去借貸；你要管轄許多國家，它們卻不能管轄你。
DEUT|15|7|「在耶和華－你上帝所賜給你的地上，任何一座城裏，你弟兄中若有一個貧窮人，你不可硬著心，袖手不幫助你貧窮的弟兄。
DEUT|15|8|你總要伸手幫助他，照他所缺乏的借給他，補他的不足。
DEUT|15|9|你要謹慎，不可心起惡念，說：『第七年的豁免年快到了』，你就冷眼看你貧窮的弟兄，甚麼都不給他。他若為你的緣故求告耶和華，你就有罪了。
DEUT|15|10|你要慷慨解囊，給他的時候不要心疼，因為耶和華－你的上帝必為這事，在你一切的工作上和你手所做的一切賜福給你。
DEUT|15|11|因為地上的貧窮人永遠不會斷絕，所以我吩咐你說：『總要伸手幫助你地上困苦貧窮的弟兄。』」
DEUT|15|12|「你弟兄中，若有一個 希伯來 男人或 希伯來 女人賣給你，已服事你六年，到了第七年就要讓他自由離開你。
DEUT|15|13|你讓他自由離開的時候，不可讓他空手而去，
DEUT|15|14|要從你的羊群、禾場、壓酒池中取一些，慷慨地送給他；耶和華－你的上帝怎樣賜福給你，你也要照樣給他。
DEUT|15|15|要記得你在 埃及 地作過奴僕，耶和華－你的上帝救贖了你。為此，我今日將這事吩咐你。
DEUT|15|16|他若對你說：『我不願意離開你』，因為他愛你和你的家，並且他在你那裏很好，
DEUT|15|17|你要拿錐子在門上穿透他的耳朵，他就永遠成為你的奴僕了。你待婢女也要這樣。
DEUT|15|18|你讓他從你那裏自由離開的時候，不要看作困難，因為他已服事你六年，相當於雇工雙倍的工錢。這樣，耶和華－你的上帝必在你所做的一切事上賜福給你。」
DEUT|15|19|「你牛群羊群中頭生的，凡是公的，都要分別為聖，歸給耶和華－你的上帝。頭生的牛，不可用牠來耕作；頭生的羊，不可剪牠的毛。
DEUT|15|20|這頭生的，你和你全家每年要到耶和華所選擇的地方，在耶和華－你上帝面前吃。
DEUT|15|21|這頭生的若有殘疾，瘸腿的或瞎眼的，若有任何嚴重缺陷，都不可獻給耶和華－你的上帝。
DEUT|15|22|你們可以在城裏吃，潔淨的人和不潔淨的人都可以吃，就如吃羚羊和鹿一樣。
DEUT|15|23|只是牠的血，你不可吃，要倒在地上，如同倒水一樣。」
DEUT|16|1|「你要守亞筆月，向耶和華－你的上帝守逾越節，因為在亞筆月，耶和華－你的上帝在夜間領你出 埃及 。
DEUT|16|2|你當在那裏，耶和華選擇作為他名居所的地方，從羊群牛群中，將逾越節的祭牲獻給耶和華－你的上帝。
DEUT|16|3|這祭牲不可和有酵的東西一起吃。因為你曾匆忙離開 埃及 地，你要吃無酵餅，就是困苦餅七日，好讓你一生的年日記得你從 埃及 地出來的那一日。
DEUT|16|4|在你全境內，七日不可見到酵母。第一日晚上所獻的肉，一點也不可留到早晨。
DEUT|16|5|你不可在耶和華－你上帝所賜的各城中，任何一座城裏，獻逾越節的祭，
DEUT|16|6|只可在那裏，耶和華－你上帝選擇作為他名居所的地方，在晚上日落的時候，就是你出 埃及 的時候，獻逾越節的祭。
DEUT|16|7|你要在耶和華－你上帝所選擇的地方把肉烤來吃，次日早晨就回到你的帳棚去。
DEUT|16|8|你要吃無酵餅六日，第七日要向耶和華－你的上帝守嚴肅會，不可做工。」
DEUT|16|9|「你要計算七個七日：從你用鐮刀開始收割莊稼時算起，一共七個七日。
DEUT|16|10|你要向耶和華－你的上帝守七七節，按照耶和華－你上帝所賜你的福，獻上你手裏的甘心祭。
DEUT|16|11|你和你的兒女、僕婢，以及住在你城裏的 利未 人、在你中間寄居的和孤兒寡婦，都要在那裏，耶和華－你上帝選擇作為他名居所的地方，在耶和華－你上帝面前歡樂。
DEUT|16|12|你要記得你在 埃及 作過奴僕，也要謹守遵行這些律例。」
DEUT|16|13|「你收藏了禾場和壓酒池的出產以後，就要守住棚節七日。
DEUT|16|14|在節期中，你和你的兒女、僕婢，以及住在你城裏的 利未 人、寄居的和孤兒寡婦，都要歡樂。
DEUT|16|15|在耶和華所選擇的地方，你要向耶和華－你的上帝守節七日，因為耶和華－你的上帝要在你一切的收成上和你手裏所做的一切賜福給你，你就非常歡樂。
DEUT|16|16|「你所有的男丁要在除酵節、七七節、住棚節，一年三次，在耶和華－你上帝所選擇的地方朝見他，不可空手朝見耶和華。
DEUT|16|17|各人要按自己手中的能力，照耶和華－你上帝所賜你的福，奉獻禮物。」
DEUT|16|18|「你要在耶和華－你上帝所賜的各城中，為各支派設立審判官和官長。他們要按公義的判斷審判百姓，
DEUT|16|19|不可屈枉正直，不可看人的情面，也不可接受賄賂，因為賄賂能使智慧人的眼睛變瞎，又能曲解義人的證詞。
DEUT|16|20|公正！你要追求公正，好使你存活，承受耶和華－你上帝所賜你的地。」
DEUT|16|21|「你為耶和華－你的上帝築壇，不可在壇旁栽種任何樹木作 亞舍拉 ，
DEUT|16|22|也不可為自己設立柱像，這是耶和華－你的上帝所憎恨的。」
DEUT|17|1|「凡有殘疾，有任何惡疾的牛羊，你都不可獻給耶和華－你的上帝，因為這是耶和華－你上帝所憎惡的。
DEUT|17|2|「在你中間，在耶和華－你上帝所賜你的各城中，任何一座城裏，若有男人或女人做了耶和華－你上帝眼中看為惡的事，違背了他的約，
DEUT|17|3|去事奉別神，敬拜它們，或拜太陽，或拜月亮，或拜天上的萬象，是我 不曾吩咐的。
DEUT|17|4|有人告訴你，你也聽見了，就要細心探聽。看哪，是真的，確實有這可憎的事在 以色列 中發生，
DEUT|17|5|你就要將行這惡事的男人或女人拉到城門外，用石頭把這男人或女人處死。
DEUT|17|6|要憑兩個證人或三個證人的口，才可以把他處死，不可只憑一個證人的口處死他。
DEUT|17|7|證人要先動手，然後眾百姓也動手把他處死。這樣，你就把惡從你中間除掉。
DEUT|17|8|「你城中若有難以判斷的案件，涉及流血，訴訟，或毆打等爭訟的事，你就要起來，上到那裏，耶和華－你上帝所選擇的地方，
DEUT|17|9|去見 利未 家的祭司和當時的審判官，求問他們，他們必將判決指示你。
DEUT|17|10|他們在耶和華所選擇的地方指示你的判決，你要執行，謹守遵行他們一切所教導你的。
DEUT|17|11|要按照所教導你的律法、所告訴你的典章去執行；他們指示你的判決，你不可偏離左右。
DEUT|17|12|若有人擅自行事，不聽從那侍立在耶和華－你上帝那裏事奉的祭司，或不聽從審判官，那人就要處死。這樣，你就把惡從 以色列 中除掉。
DEUT|17|13|眾百姓聽見了都要害怕，不再擅自行事了。」
DEUT|17|14|「你到了耶和華－你上帝所賜你的地，得了那地居住在其中的時候，若說：『我要立王治理我，像我四圍所有的國家一樣』，
DEUT|17|15|你一定要立耶和華－你上帝所揀選的人為你的王。要從你弟兄中立一人為你的王，不可立你弟兄之外的外邦人治理你。
DEUT|17|16|只是王不可為自己加添馬匹，也不可為加添馬匹使百姓回 埃及 去，因耶和華曾對你們說：『不可再回那條路去。』
DEUT|17|17|王不可為自己多立妃嬪，免得他的心偏離；也不可為自己多積金銀。
DEUT|17|18|他登了國度的王位之後，要在 利未 家的祭司面前，將這律法書為自己抄寫一份在書卷上。
DEUT|17|19|這書要存在他那裏，他一生的年日要誦讀，好使他學習敬畏耶和華－他的上帝，謹守遵行這律法書上的一切話和這些律例，
DEUT|17|20|免得他的心向弟兄高傲，偏離了這誡命，或向右或向左。這樣，他和他的子孫就可以長久作王治理 以色列 。」
DEUT|18|1|「 利未 家的祭司和 利未 全支派在 以色列 中沒有分得產業；他們可以吃耶和華的火祭，那是他的產業。
DEUT|18|2|他在弟兄中沒有產業；耶和華是他的產業，正如耶和華所應許他的。
DEUT|18|3|祭司從百姓當得的權益是這樣：凡獻牛或羊為祭物的，要把前腿、兩腮和胃給祭司。
DEUT|18|4|初收的五穀、新酒和新的油，以及初剪的羊毛，也要給他。
DEUT|18|5|因為耶和華－你的上帝從你眾支派中揀選他，使他和他子孫永遠奉耶和華的名侍立，事奉。
DEUT|18|6|「 利未 人若離開他在 以色列 中所居住的任何一座城，一心願意到耶和華所選擇的地方，
DEUT|18|7|就要在那裏奉耶和華－他上帝的名事奉，正如他的眾弟兄 利未 人在耶和華面前侍立一樣。
DEUT|18|8|除了賣祖產所得的以外，他們 要吃同等分量的祭物。」
DEUT|18|9|「你到了耶和華－你上帝所賜你之地，不可學那些國家行可憎惡的事。
DEUT|18|10|你中間不可有人使兒女經火，也不可有占卜的、觀星象的、行法術的 、行邪術的、
DEUT|18|11|施符咒的、招魂的、行巫術的和求問死人的。
DEUT|18|12|凡做這些事的都是耶和華所憎惡的；因這可憎惡的事，耶和華－你的上帝把他們從你面前趕出去。
DEUT|18|13|你要向耶和華－你的上帝作完全人。
DEUT|18|14|你所要趕出的那些國家都聽從觀星象的和占卜的，但是耶和華－你的上帝從來不准你這樣做。」
DEUT|18|15|「耶和華－你的上帝要從你弟兄中給你興起一位先知像我，你們要聽他。
DEUT|18|16|這正如你在 何烈山 大會的那日向耶和華－你的上帝所求的一切，說：『求你不要再叫我聽見耶和華－我上帝的聲音，也不要再叫我看見這大火，免得我死亡。』
DEUT|18|17|耶和華對我說：『他們說得對。
DEUT|18|18|我必在他們弟兄中給他們興起一位先知像你。我要將當說的話放在他口裏；他要將我一切所吩咐的都告訴他們。
DEUT|18|19|誰不聽從他奉我名所說的話，我必親自向他追究。
DEUT|18|20|若有先知擅自奉我的名說了我未曾吩咐他說的話，或是奉別神的名說話，那先知就必處死。』
DEUT|18|21|你心裏若說：『我們怎能知道那話是耶和華未曾吩咐的呢？』
DEUT|18|22|先知奉耶和華的名說話，所說的若沒有實現，或不應驗，這話就是耶和華未曾吩咐的，而是那先知擅自說的，你不必怕他。」
DEUT|19|1|「耶和華－你的上帝將列國剪除，他們的地耶和華－你上帝已賜給你，你又趕出他們，並且住在他們的城鎮和房屋，
DEUT|19|2|那時，你要在耶和華－你上帝所賜你為業的地上，為自己指定三座城。
DEUT|19|3|你要預備道路，將耶和華－你上帝使你承受為業的地分為三區，使任何一個殺人的可以逃到那裏去。
DEUT|19|4|「殺人的逃到那裏得以存活的案例是這樣：凡素無仇恨，無意中殺了鄰舍的，
DEUT|19|5|就如人與鄰舍同入林中伐木，手拿斧子一砍，本想砍下樹木，斧頭卻脫了把，飛落在鄰舍身上，以致那人死去，這人就可以逃到那些城中的一座，得以存活，
DEUT|19|6|免得報血仇的心中發火，去追趕那殺了人的，因為路途遙遠就能追上他，把他殺死。其實他是不該死的，因為他與被殺者素無仇恨。
DEUT|19|7|所以我吩咐你說，要為自己指定三座城。
DEUT|19|8|耶和華－你的上帝若照他向你列祖所起的誓擴張你的疆土，將所應許賜你列祖的全地給你，
DEUT|19|9|你若謹守遵行我今日所吩咐的這一切誡命，愛耶和華－你的上帝，天天遵行他的道，就要在這三座城之外，再添三座城，
DEUT|19|10|免得無辜人的血流在耶和華－你上帝所賜你為業的地中間，血就歸到你身上了。
DEUT|19|11|「若有人恨他的鄰舍，埋伏等著，起來擊殺他，把他殺死，然後逃到這些城中的一座，
DEUT|19|12|他本城的長老就要派人去，從那裏把他帶出來，交在報血仇者的手中，把他處死。
DEUT|19|13|你的眼不可顧惜他，要從 以色列 中除掉流無辜血的罪，使你得福。」
DEUT|19|14|「在耶和華－你上帝所賜你承受為業，所分得的地上，不可挪移你鄰舍的地界，因為這是前人所定的。」
DEUT|19|15|「人無論犯甚麼罪，作甚麼惡，不可單憑一個人的見證，總要憑兩個證人的口或三個證人的口才可定案。
DEUT|19|16|若有人懷惡意，起來作證，控告他人犯法，
DEUT|19|17|這兩個爭訟的人就要站在耶和華面前，和當時的祭司與審判官面前，
DEUT|19|18|審判官要細心調查。看哪，證人作的是偽證，要用偽證陷害弟兄，
DEUT|19|19|你們就要對付他如同他想要對付的弟兄一樣。這樣，你就把惡從你中間除掉。
DEUT|19|20|其他的人聽見就害怕，不敢在你中間再行這樣的惡事了。
DEUT|19|21|你的眼不可顧惜，要以命償命，以眼還眼，以牙還牙，以手還手，以腳還腳。」
DEUT|20|1|「你出去與仇敵作戰，若看見馬匹、戰車，以及比你更多的士兵，不要怕他們，因為領你出 埃及 地的耶和華－你的上帝與你同在。
DEUT|20|2|你們將要上陣的時候，祭司要來，向士兵宣告，
DEUT|20|3|對他們說：『 以色列 啊，要聽！你們今日將要與仇敵作戰，不要心驚膽戰，不要懼怕戰兢，也不要因他們驚慌，
DEUT|20|4|因為與你們同去的是耶和華－你們的上帝，他要為你們與仇敵作戰，拯救你們。』
DEUT|20|5|官長也要向士兵宣告說：『誰建了新的房屋尚未奉獻，他可以回家去，免得他陣亡，別人去奉獻。
DEUT|20|6|誰栽植了葡萄園尚未享用所結的果子，他可以回家去，免得他陣亡，別人去享用。
DEUT|20|7|誰與女子訂了婚尚未迎娶，他可以回家去，免得他陣亡，別人去娶。』
DEUT|20|8|官長要繼續對士兵說：『誰懼怕，心驚膽戰，可以回家去，免得他弟兄的心像他的心一樣消沉。』
DEUT|20|9|官長向士兵宣告完畢，軍官就率領士兵去了。
DEUT|20|10|「你來到一座城，要攻城之前，先向它宣告和平。
DEUT|20|11|那城若願意以和平回應，給你開城，城裏所有的人就要為你做苦工，服事你。
DEUT|20|12|若那城拒絕和平，卻要與你打仗，你就要圍困那城。
DEUT|20|13|耶和華－你的上帝把那城交在你手裏時，你就要用刀殺盡城裏的男丁。
DEUT|20|14|至於婦女、孩童、牲畜和城裏所有的，你都可以取為自己的掠物。從仇敵所掠奪的，就是耶和華－你上帝所賜給你的，你都可以享用。
DEUT|20|15|離你很遠的各城，就是不屬於這些國家的城鎮，你都要這樣對待他們。
DEUT|20|16|但是這些民族的城鎮，就是耶和華－你上帝所賜給你的產業，其中凡有氣息的，一個都不可存留。
DEUT|20|17|你要照耶和華－你上帝所吩咐的，將這些 赫 人、 亞摩利 人、 迦南 人、 比利洗 人、 希未 人、 耶布斯 人全都滅絕，
DEUT|20|18|免得他們教導你們去行一切可憎惡的事，就是他們向自己神明所行的，使你們得罪耶和華－你們的上帝。
DEUT|20|19|「你若圍困一座城，需要攻打許多日子才能奪取，就不可用斧頭砍壞樹木。你可以吃樹上的果子，卻不可把樹砍下來。田間的樹木豈是人，讓你去圍攻的嗎？
DEUT|20|20|只有那些你知道不能生產食物的樹才可以毀壞；你可以把它們砍下來造攻城的工具，攻打那與你打仗的城，直到把城攻下。」
DEUT|21|1|「在耶和華－你上帝所賜你為業的地上，若發現有人被殺，暴屍野地，不知道是誰殺的，
DEUT|21|2|長老和審判官 就要出去，從屍體那裏量起，量到四圍的城鎮，
DEUT|21|3|看哪一座城最靠近這屍體，那城的幾位長老就要取一頭未曾耕地、未曾負軛的母牛犢；
DEUT|21|4|那城的長老要把這母牛犢牽到流著溪水、未曾耕耘、未曾撒種的山谷去，在谷中打斷牠的頸項。
DEUT|21|5|利未 人祭司要近前來，因為耶和華－你的上帝揀選他們來事奉他，奉耶和華的名祝福，並且有任何的爭訟和毆打，都由他們的口判決。
DEUT|21|6|離屍體最近的那座城的每位長老要在山谷中，在頸項被打斷的母牛犢上面洗手，
DEUT|21|7|聲明說：『我們的手未曾流這人的血；我們的眼也未曾看見這事。
DEUT|21|8|耶和華啊，求你赦免你所救贖的百姓 以色列 ，不要讓無辜的血歸在你的百姓 以色列 中間。』這樣，他們流血的罪就必得赦免。
DEUT|21|9|你行了耶和華眼中看為正的事，就可以從你中間除掉無辜的血。」
DEUT|21|10|「你出去與仇敵作戰的時候，耶和華－你的上帝將他交在你手中，你就擄了他為俘虜。
DEUT|21|11|若你在被擄的人中看見美麗的女子，喜歡她，要娶她為妻，
DEUT|21|12|就可以帶她到你家去。她要剪頭髮，修指甲，
DEUT|21|13|脫去被擄時所穿的衣服，住在你家裏為自己父母哀哭一個月。然後，你就可以與她同房；你作她的丈夫，她作你的妻子。
DEUT|21|14|以後你若不喜歡她，就要讓她自由離開，絕不可為錢把她賣了，也不可把她當奴隸看待，因為你已經佔有過她。」
DEUT|21|15|「人若有兩個妻子，一個是他寵愛的，另一個是失寵的 ，她們都給他生了兒子，但長子是他失寵妻子生的；
DEUT|21|16|到了分產業給兒子的時候，不可將自己寵愛的妻子所生的兒子立為長子，在他失寵妻子所生的長子之上。
DEUT|21|17|他必須認失寵妻子所生的兒子為長子，在所有的產業中給他雙分，因為這兒子是他壯年時生的，長子的名分應當是他的。」
DEUT|21|18|「人若有頑梗忤逆的兒子，不聽從父母的話，他們雖然懲戒他，他還是不聽從他們，
DEUT|21|19|父母就要抓住他，帶他出去到當地的城門，本城的長老那裏，
DEUT|21|20|對本城的長老說：『我們這個兒子頑梗忤逆，不聽從我們的話，是貪食好酒的人。』
DEUT|21|21|然後，城裏的眾人就要用石頭將他打死。這樣，你就把惡從你中間除掉，全 以色列 聽見了都要害怕。」
DEUT|21|22|「人若犯了死罪被處死，你把他掛在木頭上，
DEUT|21|23|不可讓屍體留在木頭上過夜，一定要當日把他埋葬，因為被掛的人是上帝所詛咒的。你不可玷污耶和華－你上帝所賜你為業的地。」
DEUT|22|1|「你若看見弟兄的牛或羊迷了路，不可避開牠們，總要把牠們牽回來交給你的弟兄。
DEUT|22|2|你弟兄若離你遠，或是你不認識他，你就要牽到你家，留在你那裏，等你的弟兄來尋找就還給他。
DEUT|22|3|你弟兄所失落的，無論是驢，衣服，或任何東西，你若發現，都要這樣做，不能避開。
DEUT|22|4|你若看見你弟兄的牛或驢在路上跌倒了，不可避開牠們，總要幫助他把牛或驢拉起來。
DEUT|22|5|「婦女不可穿戴男子所穿戴的，男人也不可穿婦女的衣服，因為這樣做是耶和華－你上帝所憎惡的。
DEUT|22|6|「你若路上看見鳥窩，無論在樹上或地上，裏頭有小鳥或有蛋，母鳥伏在小鳥或蛋上，你不可連母鳥帶小鳥一起拿去。
DEUT|22|7|總要放母鳥走，只可以取小鳥。這樣你就可以享福，日子得以長久。
DEUT|22|8|「你若建造新房屋，要在屋頂安欄杆，免得有人從屋頂掉下來，血就歸於你家。
DEUT|22|9|「不可在你的葡萄園裏栽種別的種子，免得你栽種所結的和葡萄園的果子都成了聖物。
DEUT|22|10|不可並用牛和驢來耕地。
DEUT|22|11|不可穿羊毛和細麻混合做成的衣服。
DEUT|22|12|「你要在所披外衣的四個邊上縫繸子。」
DEUT|22|13|「人若娶妻，與她同房後恨惡她，
DEUT|22|14|捏造她行可恥的事，把醜名加在她身上，說：『我娶了這女人，親近她，卻發現她沒有貞潔的憑據』。
DEUT|22|15|女方的父母就要把這女子貞潔的憑據拿出去，到城門的本城長老那裏。
DEUT|22|16|女方的父親要對長老說：『我把女兒嫁給這人，他卻恨惡她，
DEUT|22|17|看哪，他捏造可恥的事，說：我發現你女兒沒有貞潔的憑據。但是，這就是我女兒貞潔的憑據。』父母要把那布鋪在本城長老的面前。
DEUT|22|18|那城的長老要拿住那人，懲罰他，
DEUT|22|19|罰他一百銀子，給女方的父親，因為他把醜名加在 以色列 一個少女身上。這女子仍是他的妻子，那人終身不可休她。
DEUT|22|20|但若這事是真的，找不到女子貞潔的憑據，
DEUT|22|21|他們就要把這女子帶到她父家的門口，城裏的人要用石頭打死她，因為她在父家犯了淫亂，在 以色列 中做了可恥的事。這樣，你就把惡從你中間除掉。
DEUT|22|22|「若發現有人與有夫之婦同寢，就要將姦夫淫婦一起處死。這樣，你就把惡從 以色列 中除掉。
DEUT|22|23|「若一女子是處女，已經許配了人，有男子在城裏遇見她，與她同寢，
DEUT|22|24|你們就要把這二人帶到那城的城門口，用石頭打死他們。處死女子是因為她雖然在城裏， 卻沒有喊叫；處死男子是因為他玷污了鄰舍的妻子。這樣，你就把惡從你中間除掉。
DEUT|22|25|「若有男子在野地遇見已經許配人的女子，抓住她與她同寢，只要處死那與女子同寢的男子。
DEUT|22|26|不可對女子處刑，這女子沒有該死的罪。這案件就好比人起來攻擊鄰舍，把他殺了一樣。
DEUT|22|27|因為男子是在野地遇見她，這已經許配了人的女子雖然喊叫，卻沒有人救她。
DEUT|22|28|「若有男子遇見沒有許配人的少女，抓住她與她同寢，被人發現，
DEUT|22|29|這男子就要拿五十銀子給女子的父親，並要娶她為妻，終身不可休她，因為他玷污了這女子。
DEUT|22|30|「人不可娶繼母為妻，不可掀開父親衣服的下邊 。」
DEUT|23|1|「凡外腎損傷的，或被閹割的，不可入耶和華的會。
DEUT|23|2|「私生子不可入耶和華的會；甚至到第十代，也不可入耶和華的會。
DEUT|23|3|「 亞捫 人或 摩押 人不可入耶和華的會；甚至到第十代，也永不可入耶和華的會。
DEUT|23|4|因為你們出 埃及 的時候，他們沒有拿食物和水在路上迎接你們，並且雇了 美索不達米亞 的 毗奪 人， 比珥 的兒子 巴蘭 來詛咒你。
DEUT|23|5|然而耶和華－你的上帝不願聽 巴蘭 ，耶和華－你的上帝為你使詛咒變為祝福，因為耶和華－你的上帝愛你。
DEUT|23|6|你一生一世永不可為他們求平安和福氣。
DEUT|23|7|「不可憎惡 以東 人，因為他是你的弟兄。不可憎惡 埃及 人，因為你曾在他的地上作過寄居的。
DEUT|23|8|他們所生的第三代子孫可以入耶和華的會。」
DEUT|23|9|「你出兵攻打敵人，要遠離一切惡事。
DEUT|23|10|「你中間若有人因夜間夢遺而不潔淨，就要出到營外，不可入營。
DEUT|23|11|到了傍晚，他要用水洗澡，等到日落才可以入營。
DEUT|23|12|「你要在營外劃定一個地方，你可以出去在那裏方便。
DEUT|23|13|在你器械中當有一把鍬；你出營外便溺以後，要用它挖洞，轉身掩蓋排泄物。
DEUT|23|14|因為耶和華－你的上帝在你營中走動，要拯救你，將仇敵交給你，所以你的營應當聖潔，免得他見你那裏有污穢之物就轉身離開你。」
DEUT|23|15|「你不可把從主人身邊逃到你那裏的奴僕，交回給他的主人，
DEUT|23|16|要讓他在你那裏與你同住，由他在你的城鎮中選擇一個自己喜歡的地方居住，不可欺負他。
DEUT|23|17|「 以色列 的女子中不可作神廟娼妓； 以色列 的男子中也不可作神廟娼妓。
DEUT|23|18|妓女和男娼 的賞金，都不可帶進耶和華－你上帝的殿中還願，因為兩者都是耶和華－你上帝所憎惡的。
DEUT|23|19|「你借給你弟兄的，無論是錢財是糧食，或任何可生利息的財物，都不可取利。
DEUT|23|20|借給外邦人可以取利，但借給你的弟兄就不可取利；好讓耶和華－你的上帝在你去得為業的地上和你手裏所做的一切，賜福給你。
DEUT|23|21|「你向耶和華－你的上帝許願，不可遲延還願，因為耶和華－你的上帝必定向你追討，你就有罪了。
DEUT|23|22|你若不許願，倒沒有罪。
DEUT|23|23|你嘴唇所說的，你親口承諾的，要照你甘心向耶和華－你上帝許的願謹守遵行。
DEUT|23|24|「你進入鄰舍的葡萄園，可以隨意吃葡萄，直到飽足，卻不可裝在器皿中。
DEUT|23|25|你進入鄰舍的莊稼中，可以用手摘麥穗，卻不可用鐮刀割取莊稼。」
DEUT|24|1|「人若娶妻，作了她的丈夫，發現她有不合宜的事不喜歡她，而寫休書交在她手中，打發她離開夫家，
DEUT|24|2|婦人若離開夫家以後，去嫁別人，
DEUT|24|3|後夫若恨惡她，寫休書交在她手中，打發她離開夫家，又或者娶她為妻的後夫死了，
DEUT|24|4|那休她的前夫就不可在婦人玷污之後再娶她為妻，因為這是耶和華所憎惡的。不可使耶和華－你上帝所賜為業之地蒙受玷污。
DEUT|24|5|「人若娶了新娘，不可從軍出征，也不可派他辦理任何事情。他可以在家清閒一年，使他所娶的妻快活。
DEUT|24|6|「不可拿人的石磨或上面的磨石作抵押，因為這是拿人的命作抵押。
DEUT|24|7|「若發現有人綁架 以色列 人中的一個弟兄，把他當奴隸對待，或把他賣了，那綁架人的就必處死。這樣，你就把惡從你中間除掉。
DEUT|24|8|「關於痲瘋 的災病，你們要謹慎，照 利未 家的祭司一切所指教你們的留心遵行。我怎樣吩咐他們，你們要照樣遵行。
DEUT|24|9|要記得，在你們出 埃及 後的路途中，耶和華－你的上帝向 米利暗 所做的事。
DEUT|24|10|「你借給鄰舍，無論是甚麼，不可進他家拿抵押品。
DEUT|24|11|要站在外面，等那借貸的人把抵押品拿出來交給你。
DEUT|24|12|他若是困苦的人，你不可用他的抵押品蓋著睡覺。
DEUT|24|13|日落的時候，總要把抵押品還給他，讓他用那件外衣蓋著睡覺，他就為你祝福。這在耶和華－你的上帝面前就是你的義行了。
DEUT|24|14|「困苦貧窮的雇工，無論是你的弟兄，或是住在你境內，在你城裏寄居的，你都不可欺負他 。
DEUT|24|15|要當日給他工錢，不可等到日落，因為他困苦，需要靠工錢過活，免得他因你的緣故求告耶和華，罪就歸於你了。
DEUT|24|16|「不可因兒子處死父親，也不可因父親處死兒子；各人要因自己的罪被處死。
DEUT|24|17|「不可對寄居的和孤兒屈枉正直，也不可拿寡婦的衣服作抵押。
DEUT|24|18|要記得你曾在 埃及 作過奴僕，耶和華－你的上帝從那裏救贖了你，所以我吩咐你遵行這事。
DEUT|24|19|「你在田間收割莊稼，若忘了一捆在田間，就不要再回去拿，要留給寄居的、孤兒和寡婦；好讓耶和華－你的上帝在你手裏所做的一切，賜福給你。
DEUT|24|20|你打了橄欖樹，枝上剩下的不可再打，要留給寄居的、孤兒和寡婦。
DEUT|24|21|你摘葡萄園的葡萄，掉落的不可拾取，要留給寄居的、孤兒和寡婦。
DEUT|24|22|你要記得你曾在 埃及 地作過奴僕，所以我吩咐你遵行這事。
DEUT|25|1|「人與人若有爭訟，要求審判，當宣判義人為義，惡人有罪的時候，
DEUT|25|2|惡人若該受責打，審判官就要叫他當著面，伏在地上，按他的罪照數責打。
DEUT|25|3|只能打四十下，不可加多；多過這數目就是在你眼中作賤你的弟兄了。
DEUT|25|4|「牛在踹穀的時候，不可籠住牠的嘴。」
DEUT|25|5|「兄弟住在一起，若其中一個死了，沒有兒子，死者的妻子就不可出去嫁給陌生人。她丈夫的兄弟應當盡兄弟的本分，娶她為妻，與她同房。
DEUT|25|6|婦人生的長子要歸在已故兄弟的名下，免得他的名在 以色列 中塗去了。
DEUT|25|7|那人若不情願娶他兄弟的妻子，他兄弟的妻子就要上到城門長老那裏，說：『我丈夫的兄弟拒絕在 以色列 中為他的兄弟留名，不願意為我盡兄弟的本分。』
DEUT|25|8|本城的長老就要召那人來，跟他談話。若他堅持說：『我不情願娶她。』
DEUT|25|9|他兄弟的妻子就要在長老眼前來到那人跟前，脫下他腳上的鞋，吐唾沫在他臉上，回應說：『凡不為兄弟建立家室的都要這樣待他。』
DEUT|25|10|在 以色列 中，他要以『脫鞋之家』聞名。」
DEUT|25|11|「若有人和弟兄爭鬥，其中一人的妻子近前去，為了救丈夫脫離那打丈夫之人的手，伸手抓住那人的下體，
DEUT|25|12|你就要砍斷婦人的手，你的眼不可顧惜。
DEUT|25|13|「你袋中不可有一大一小兩樣的法碼。
DEUT|25|14|你家裏不可有一大一小兩樣的伊法 。
DEUT|25|15|當用準確公正的法碼和伊法，好使你的日子在耶和華－你上帝所賜你的地上得以長久。
DEUT|25|16|因為行這一切不義之事的人都是耶和華－你上帝所憎惡的。」
DEUT|25|17|「你要記得你們出 埃及 的時候， 亞瑪力 在路上怎樣對待你，
DEUT|25|18|在路上迎擊你，趁你疲乏困倦時擊殺所有在你後面軟弱的人；並不敬畏上帝。
DEUT|25|19|所以，當耶和華－你的上帝使你不被四圍一切仇敵擾亂，在耶和華－你上帝賜你為業的地上得享平靜的時候，你要把 亞瑪力 的名從天下塗去；你不可忘記這事。」
DEUT|26|1|「你進去得了耶和華－你上帝所賜你為業的地，並且居住在那裏的時候，
DEUT|26|2|就要從耶和華－你上帝所賜你的地上，將收成的各種初熟土產取一些來，盛在筐子裏，帶到那裏，耶和華－你上帝選擇作為他名居所的地方，
DEUT|26|3|到當時的祭司那裏，對他說：『我今日向耶和華－你的上帝宣認，我已來到耶和華向我們列祖起誓要賜給我們的地。』
DEUT|26|4|祭司就從你手裏把筐子接過來，供在耶和華－你上帝的祭壇前。
DEUT|26|5|你要在耶和華－你上帝面前告白說：『我的祖先原是一個流亡的 亞蘭 人，帶著稀少的人丁下到 埃及 寄居。在那裏，他卻成了又大又強、人數眾多的國。
DEUT|26|6|埃及 人惡待我們，迫害我們，將苦工加在我們身上。
DEUT|26|7|於是我們哀求耶和華我們列祖的上帝。耶和華聽見我們的聲音，看見我們所受的困苦、勞役和欺壓，
DEUT|26|8|耶和華就用大能的手和伸出來的膀臂，以及大而可畏的事和神蹟奇事，領我們出了 埃及 ，
DEUT|26|9|將我們領進這地方，把這流奶與蜜之地賜給我們。
DEUT|26|10|耶和華啊，看哪，現在我把你所賜我地上初熟的土產供上。』隨後你要把筐子供在耶和華－你上帝面前，向耶和華－你的上帝下拜。
DEUT|26|11|你和 利未 人，以及在你中間寄居的，要因耶和華－你上帝所賜你和你家的一切福分歡樂。
DEUT|26|12|「每逢第三年，就是捐十分之一的那年，你從你一切土產中取了十分之一，要分給 利未 人、寄居的、孤兒和寡婦，使他們在你的城鎮中可以吃得飽足。
DEUT|26|13|你又要在耶和華－你上帝面前說：『我已將聖物從家裏拿出來，給了 利未 人、寄居的、孤兒和寡婦，是遵照你吩咐我的一切命令。你的命令，我沒有違背，也沒有忘記。
DEUT|26|14|我守喪的時候，沒有吃這聖物，不潔淨的時候，也沒有拿出來，又沒有把它獻給死人。我聽從了耶和華－我上帝的話，都照你一切所吩咐的做了。
DEUT|26|15|求你從天上，從你的聖所垂看，賜福給你的百姓 以色列 和你向我們列祖起誓所賜給我們的這片土地，就是流奶與蜜之地。』」
DEUT|26|16|「耶和華－你的上帝今日吩咐你遵行這些律例典章，所以你要盡心盡性謹守遵行。
DEUT|26|17|你今日宣認耶和華為你的上帝，承諾遵行他的道，謹守他的律例、誡命、典章，聽從他的話。
DEUT|26|18|耶和華今日照他所應許你的，也認你為他寶貴的子民，叫你謹守他的一切誡命，
DEUT|26|19|要使你得稱讚、美名、尊榮，超乎他所造的萬國之上，並且照他所應許的，使你歸耶和華－你的上帝為神聖的子民。」
DEUT|27|1|摩西 和 以色列 的眾長老吩咐百姓說：「你們要遵守我今日所吩咐的一切誡命。
DEUT|27|2|你們過了 約旦河 ，到耶和華－你上帝所賜給你的地，當日要豎立幾塊大石頭，塗上石灰。
DEUT|27|3|當你過了河，進入耶和華－你上帝所賜給你流奶與蜜之地，正如耶和華－你列祖的上帝所應許你的，你要把這律法的一切話寫在石頭上。
DEUT|27|4|你們過了 約旦河 ，就要在 基利心山 上照我今日所吩咐的，把這些石頭豎立起來，塗上石灰。
DEUT|27|5|你在那裏要為耶和華－你的上帝築一座石壇，卻不可動用鐵器在石頭上。
DEUT|27|6|要用沒有鑿過的石頭築耶和華－你上帝的壇，在壇上將燔祭獻給耶和華－你的上帝，
DEUT|27|7|又要獻平安祭，在那裏吃，在耶和華－你的上帝面前歡樂。
DEUT|27|8|你要將這律法的一切話清楚地寫在石頭上。」
DEUT|27|9|摩西 和 利未 家的祭司吩咐 以色列 眾人說：「 以色列 啊，你要靜默傾聽！你今日已成為耶和華－你上帝的子民了。
DEUT|27|10|你要聽從耶和華－你上帝的話，遵行他的誡命律例，就是我今日所吩咐你的。」
DEUT|27|11|當日， 摩西 吩咐百姓說：
DEUT|27|12|「你們過了 約旦河 ， 西緬 、 利未 、 猶大 、 以薩迦 、 約瑟 和 便雅憫 等支派的人要站在 基利心山 上為百姓祝福。
DEUT|27|13|呂便 、 迦得 、 亞設 、 西布倫 、 但 和 拿弗他利 等支派的人要站在 以巴路山 上宣佈詛咒。
DEUT|27|14|利未 人要大聲對 以色列 眾人說：
DEUT|27|15|「『凡製造耶和華所憎惡的偶像，無論是雕刻的，是鑄造的，就是工匠用手造的，或暗中設置的，這人必受詛咒！』眾百姓要回應說：『阿們！』
DEUT|27|16|「『輕慢父母的，必受詛咒！』眾百姓要說：『阿們！』
DEUT|27|17|「『挪移鄰舍地界的，必受詛咒！』眾百姓要說：『阿們！』
DEUT|27|18|「『引領瞎子走錯路的，必受詛咒！』眾百姓要說：『阿們！』
DEUT|27|19|「『對寄居的、孤兒和寡婦屈枉正直的，必受詛咒！』眾百姓要說：『阿們！』
DEUT|27|20|「『與繼母同寢的，必受詛咒！因為他掀開父親衣服的下邊。』眾百姓要說：『阿們！』
DEUT|27|21|「『與獸交合的，必受詛咒！』眾百姓要說：『阿們！』
DEUT|27|22|「『與同父異母，或同母異父的姊妹同寢的，必受詛咒！』眾百姓要說：『阿們！』
DEUT|27|23|「『與岳母同寢的，必受詛咒！』眾百姓要說：『阿們！』
DEUT|27|24|「『暗中擊殺鄰舍的，必受詛咒！』眾百姓要說：『阿們！』
DEUT|27|25|「『受賄賂擊殺人而流無辜之血的，必受詛咒！』眾百姓要說：『阿們！』
DEUT|27|26|「『不堅守遵行這律法之話的，必受詛咒！』眾百姓要說：『阿們！』」
DEUT|28|1|「你若留心聽從耶和華－你上帝的話，謹守遵行他的一切誡命，就是我今日所吩咐你的，他必使你超乎地上的萬國之上。
DEUT|28|2|你若聽從耶和華－你上帝的話，這一切的福氣必臨到你身上，追隨你：
DEUT|28|3|你在城裏必蒙福，在田間也必蒙福。
DEUT|28|4|你身所生的，你地所產的，你牲畜所生的，牛犢、羔羊，都必蒙福。
DEUT|28|5|你的筐子和你的揉麵盆都必蒙福。
DEUT|28|6|你出也蒙福，入也蒙福。
DEUT|28|7|「耶和華必使那起來攻擊你的仇敵在你面前潰敗。他們從一條路來攻擊你，必在你面前從七條路逃跑。
DEUT|28|8|在你倉房裏，以及你手所做的一切，耶和華必發令賜福給你。耶和華－你上帝也必在所賜你的地上賜福給你。
DEUT|28|9|你若謹守耶和華－你上帝的誡命，遵行他的道，他必照他向你所起的誓立你為自己神聖的子民。
DEUT|28|10|地上的萬民見你歸在耶和華的名下，就必懼怕你。
DEUT|28|11|在耶和華向你列祖起誓應許賜你的土地上，他必使你身所生的，牲畜所生的，地所產的，都豐富有餘。
DEUT|28|12|耶和華必為你敞開天上的寶庫，按時降雨在你的地上。他必賜福你手裏所做的一切。你必借給許多國家，卻不必去借貸。
DEUT|28|13|你若聽從耶和華－你上帝的誡命，就是我今日所吩咐你的，謹守遵行，耶和華就必使你作首不作尾，居上不居下，
DEUT|28|14|只要你不偏左右，不背離我今日所吩咐你的一切話，也不隨從別神，事奉它們。」
DEUT|28|15|「你若不聽從耶和華－你上帝的話，不謹守遵行他的一切誡命律例，就是我今日所吩咐你的，這一切的詛咒必臨到你身上，追隨你：
DEUT|28|16|你在城裏必受詛咒，在田間也必受詛咒。
DEUT|28|17|你的筐子和你的揉麵盆都必受詛咒。
DEUT|28|18|你身所生的，你地所產的，以及牛犢、羔羊，都必受詛咒。
DEUT|28|19|你出也受詛咒，入也受詛咒。
DEUT|28|20|耶和華因你作惡離棄他，必在你手裏所做的一切，使詛咒、困擾、責罰臨到你，直到你被除滅，直到你迅速滅亡。
DEUT|28|21|耶和華必使瘟疫緊貼著你，直到他把你從所進去得為業的地上滅絕。
DEUT|28|22|耶和華要用癆病、熱病、發炎、高燒、刀劍 、焚風 和霉爛攻擊你；這些要追趕你，直到你滅亡。
DEUT|28|23|你頭上的天要變成銅，下面的地要化為鐵。
DEUT|28|24|耶和華要使那降在你地上的雨變為灰塵，塵土從天落在你身上，直到你被除滅。
DEUT|28|25|「耶和華必使你在仇敵面前潰敗。你從一條路去攻擊他們，必從七條路逃跑。地上萬國必因你而驚駭。
DEUT|28|26|你的屍首必給空中的飛鳥和地上的走獸作食物，卻無人鬨趕。
DEUT|28|27|耶和華必用 埃及 人的瘡、潰瘍、癬和疥攻擊你，使你不得醫治。
DEUT|28|28|耶和華必用癲狂、眼瞎、心驚攻擊你。
DEUT|28|29|你必在午間摸索，好像盲人在黑暗中摸索。你的道路必不亨通，天天受人欺壓、搶奪，無人搭救。
DEUT|28|30|你聘了妻子，別人必與她同寢；你建了房屋，卻不得住在其內；你栽植了葡萄園，卻不得享用所結的果子。
DEUT|28|31|你的牛在你眼前宰了，你吃不到牠的肉；你的驢在你眼前被人搶奪，卻討不回來；你的羊被敵人拿走，無人幫助你。
DEUT|28|32|你的兒女被交給別國的民；你的眼目終日切望，甚至失明，你的手卻無能為力。
DEUT|28|33|你地所產的和你勞力所得的，必被你所不認識的百姓吃盡。你天天只被欺負，受壓制，
DEUT|28|34|甚至你因眼中所見的景象而瘋狂。
DEUT|28|35|耶和華必攻擊你，使你膝上腿上，從腳掌到頭頂，都長滿了毒瘡，無法醫治。
DEUT|28|36|「耶和華必將你和你所立統治你的王，領到你和你列祖不認識的國去；在那裏你必事奉別神，就是木頭和石頭。
DEUT|28|37|你在耶和華趕你到的萬民中，要令人驚駭，成為笑柄，被人譏誚。
DEUT|28|38|你撒在田裏的種子雖多，收的卻少，因為蝗蟲把它吃光了。
DEUT|28|39|你栽植修整葡萄園，卻沒有酒喝，也不得儲存，因為蟲子把它吃了。
DEUT|28|40|你全境有橄欖樹，卻得不到油抹身，因為你的橄欖都掉光了。
DEUT|28|41|你生兒育女，卻不屬於你，因為他們必被擄去。
DEUT|28|42|你所有的樹木和你地裏的出產必被蝗蟲吃盡了。
DEUT|28|43|在你中間寄居的必上升高過你，高而又高；你必下降，低而又低。
DEUT|28|44|他必借給你，你卻不能借給他；他必作首，你必作尾。
DEUT|28|45|這一切的詛咒必臨到你，追趕你，趕上你，直到把你除滅，因為你不聽從耶和華－你上帝的話，不遵守他吩咐的誡命律例。
DEUT|28|46|這些詛咒必在你和你後裔身上成為神蹟奇事，直到永遠！
DEUT|28|47|因為你富裕的時候，不以歡喜快樂的心事奉耶和華－你的上帝，
DEUT|28|48|所以你必在飢餓、乾渴、赤身、缺乏中事奉仇敵，那是耶和華派來攻擊你的。他必把鐵軛加在你的頸項上，直到把你除滅。
DEUT|28|49|耶和華要從遠方、地極之處帶一國來，如鷹飛來攻擊你；這國的語言，你聽不懂。
DEUT|28|50|這國的人面貌兇惡，不給長者面子，也不恩待年輕人。
DEUT|28|51|他們必吃你牲畜所生的和你土地所產的，直到你被除滅。你的五穀、新酒和新的油，以及牛犢、羔羊，他都不給你留下，直到使你滅亡。
DEUT|28|52|他們必在你的各城圍困你，直到你在全地所倚靠、高大堅固的城牆都倒塌。他們必在耶和華－你上帝所賜給你全地的各城圍困你。
DEUT|28|53|你在仇敵圍困的窘迫中，必吃你本身所生的，就是耶和華－你上帝所賜給你的兒女之肉。
DEUT|28|54|你中間，連那溫和文雅的人都必冷眼惡待自己的兄弟和懷中的妻子，以及他所剩下其餘的兒女，
DEUT|28|55|不把所吃兒女的肉分一點給他們任何一個人，因為在被仇敵圍困、陷入窘迫的各城中，他已經一無所剩了。
DEUT|28|56|你中間柔順嬌嫩的婦人，甚至因柔順嬌嫩腳不肯踏地的婦人，也必冷眼惡待她懷中的丈夫和自己的兒女。
DEUT|28|57|在被仇敵圍困、陷入窘迫的城鎮中，她因缺乏一切，就要暗中把從她兩腿中間出來的胞衣和所生下的兒女吃了。
DEUT|28|58|「這書上所寫律法的一切話，是叫你敬畏耶和華－你上帝尊榮可畏的名，你若不謹守遵行，
DEUT|28|59|耶和華就必將奇異的災害，就是嚴重持久的災害和長期難治的疾病，加在你和你後裔的身上。
DEUT|28|60|他必使你所畏懼、 埃及 一切的疾病臨到你，緊貼著你，
DEUT|28|61|沒有寫在這律法書上的各樣疾病、災害，耶和華也必降在你身上，直到你被除滅。
DEUT|28|62|你們雖然曾像天上的星那樣多，卻因不聽從耶和華－你上帝的話，所剩的人丁就稀少了。
DEUT|28|63|耶和華先前怎樣喜愛善待你們，使你們增多，耶和華也要照樣喜愛消滅你們，使你們滅絕。你們必從所要進去得為業的地上被拔除。
DEUT|28|64|耶和華必把你們分散在萬民中，從地的這邊到地的另一邊，在那裏你必事奉你和你列祖不認識的神明，就是木頭和石頭。
DEUT|28|65|在那些國中，你必得不到安寧，腳掌也沒有安歇之處；耶和華卻要使你在那裏心中發顫，眼目失明，精神沮喪。
DEUT|28|66|你的一生懸空不安；你晝夜恐懼，生命沒有保障。
DEUT|28|67|你因心中的恐懼，眼睛所見的景象，早晨必說：『但願現在是晚上！』晚上必說：『但願現在是早晨！』
DEUT|28|68|耶和華要用船把你送回 埃及 去，走那我曾告訴你不再看見的路；在那裏你們必賣身給你的仇敵作奴婢，卻沒有人要買。」
DEUT|29|1|耶和華在 何烈山 與 以色列 人立約以外，這是耶和華在 摩押 地吩咐 摩西 與 以色列 人立約的話。
DEUT|29|2|摩西 召全 以色列 來，對他們說：「耶和華在 埃及 地，在你們眼前向法老和他眾臣僕，以及他的全地所做的一切事，你們都看見了，
DEUT|29|3|就是你親眼看見的大考驗，那些神蹟和大奇事。
DEUT|29|4|但耶和華到今日還沒有使你們心能明白，眼能看見，耳能聽見。
DEUT|29|5|我領你們在曠野四十年，你們身上的衣服沒有穿破，腳上的鞋也沒有穿壞；
DEUT|29|6|你們沒有吃餅，也沒有喝清酒烈酒，好讓你們知道『我─耶和華是你們的上帝』。
DEUT|29|7|你們來到這地方， 希實本 王 西宏 和 巴珊 王 噩 出來迎擊我們，與我們交戰，我們擊敗了他們，
DEUT|29|8|取了他們的地，給 呂便 支派、 迦得 支派和 瑪拿西 半支派為業。
DEUT|29|9|所以你們要謹守這約的話，遵行它們，好使你們在一切所做的事上亨通。
DEUT|29|10|「今日你們全都要站在耶和華－你們的上帝面前，就是各領袖、族長 、長老、官長、 以色列 所有的男子、
DEUT|29|11|你們的妻子兒女、你營中寄居的，從為你砍柴到為你挑水的人，
DEUT|29|12|為要使你進入耶和華－你上帝的約，就是耶和華－你上帝今日向你起誓所立的；
DEUT|29|13|這樣，他今日要立你作他的子民，他作你的上帝，是照他向你所應許的，又照他向你列祖 亞伯拉罕 、 以撒 、 雅各 所起的誓。
DEUT|29|14|我不單單與你們立這約，起這誓，
DEUT|29|15|就是今日與我們一同站在耶和華－我們上帝面前的，而且也包括今日不在我們這裏的人。
DEUT|29|16|「你們知道，我們曾住過 埃及 地，也經過列國，從他們中間穿越。
DEUT|29|17|你們也見過他們的可憎之物，他們木、石、金、銀的偶像。
DEUT|29|18|惟恐你們中間有人，或男或女，或宗族或支派，今日心裏偏離耶和華－我們的上帝，去事奉那些國的神明，又怕你們中間有根長出苦菜和茵蔯來。
DEUT|29|19|這樣的人聽見這詛咒的話，心裏還慶幸，說：『我雖然隨著頑固的心行事，卻還是平安無事。』以致有水的和無水的都消滅了。
DEUT|29|20|耶和華必不願饒恕他；耶和華的怒氣與妒忌必向他如煙冒出，將這書上所寫的一切詛咒都加在他身上，耶和華也要從天下塗去他的名。
DEUT|29|21|耶和華又必照著寫在律法書上，約中的一切詛咒，將他從 以色列 眾支派中分別出來，使他遭受禍害。
DEUT|29|22|你們的後代，就是接續你們興起的子孫，和遠方來的外邦人，看見這地的災禍，以及耶和華所降於這地的疾病，
DEUT|29|23|遍地都被硫磺和鹽所侵蝕，不能耕種，沒有出產，連草都長不出來，好像耶和華在怒氣和憤怒中所傾覆的 所多瑪 、 蛾摩拉 、 押瑪 、 洗扁 一樣，
DEUT|29|24|萬國必說：『耶和華為甚麼向此地這樣做呢？為甚麼要大發烈怒呢？』
DEUT|29|25|人必說：『這是因為這地的人離棄了耶和華─他們列祖的上帝領他們出 埃及 地的時候與他們所立的約，
DEUT|29|26|去事奉別神，敬拜他們所不認識的神明，這是耶和華未曾允許的。
DEUT|29|27|所以耶和華的怒氣向這地發作，將這書上所寫的一切詛咒都降在這地上。
DEUT|29|28|耶和華在怒氣、憤怒、大惱恨中將他們從本地拔出來，扔到別的地上，像今日一樣。』
DEUT|29|29|「隱祕的事是屬耶和華─我們上帝的，但明顯的事是永遠屬我們和我們子孫的，為要叫我們遵行這律法上的一切話。」
DEUT|30|1|「當這一切的事，就是我擺在你面前的祝福和詛咒臨到你的時候，你在耶和華－你上帝趕逐你去的萬國中，心裏回想這些事，
DEUT|30|2|你和你的子孫若盡心盡性歸向耶和華－你的上帝，照我今日一切所吩咐你的，聽從他的話，
DEUT|30|3|耶和華－你的上帝就必憐憫你，使你這被擄的子民歸回。耶和華－你的上帝必轉回，從分散你到的萬民中把你召集回來。
DEUT|30|4|你就是被趕逐到天涯，耶和華－你的上帝也必從那裏召集你，從那裏領你回來。
DEUT|30|5|耶和華－你的上帝必領你進入你列祖所得的地，你必得著這地為業。他必善待你，使你增多，勝過你的列祖。
DEUT|30|6|耶和華－你的上帝要使你的心和你後裔的心受割禮，好叫你盡心盡性愛耶和華－你的上帝，使你可以存活。
DEUT|30|7|耶和華－你的上帝必將這一切詛咒加在你仇敵和恨惡你、迫害你的人身上。
DEUT|30|8|你必回轉，聽從耶和華的話，遵行他的一切誡命，就是我今日所吩咐你的。
DEUT|30|9|耶和華－你的上帝必使你手裏所做的一切，以及你身所生的，牲畜所生的，土地所產的都豐富有餘，而且順利；耶和華必再喜愛善待你，正如他喜愛你的列祖一樣，
DEUT|30|10|只要你聽從耶和華－你上帝的話，謹守這律法書上所寫的誡命律例，盡心盡性歸向耶和華－你的上帝。」
DEUT|30|11|「我今日所吩咐你的誡命，對你並不困難，也不太遠；
DEUT|30|12|不是在天上，使你說：『誰為我們上天去取來給我們，使我們聽了可以遵行呢？』
DEUT|30|13|也不是在海的那邊，使你說：『誰為我們渡海到另一邊，去取來給我們，使我們聽了可以遵行呢？』
DEUT|30|14|因這話離你很近，就在你口中，在你心裏，使你可以遵行。
DEUT|30|15|「看，我今日將生死禍福擺在你面前。
DEUT|30|16|我今日所吩咐你的 ，就是要愛耶和華－你的上帝，遵行他的道，謹守他的誡命、律例、典章，使你可以存活，增多，而且耶和華－你的上帝必在你所要進去得為業的地上賜福給你。
DEUT|30|17|倘若你的心偏離，不肯聽從，卻被引誘去敬拜別神，事奉它們，
DEUT|30|18|我今日向你們申明，你們必定滅亡；在你過 約旦河 進去得為業的地上，你的日子必不長久。
DEUT|30|19|我今日呼天喚地向你作見證：我已經將生與死，祝福與詛咒，擺在你面前。所以你要揀選生命，好使你和你的後裔都得存活。
DEUT|30|20|要愛耶和華－你的上帝，聽從他的話，緊緊跟隨他，因為他是你的生命，必使你的日子得以長久，可以在耶和華向你列祖 亞伯拉罕 、 以撒 、 雅各 起誓要給他們的地上居住。」
DEUT|31|1|摩西 去把這些話吩咐 以色列 眾人 ，
DEUT|31|2|對他們說：「我已經一百二十歲了，現在不能照常出入。耶和華曾對我說：『你不得過這 約旦河 。』
DEUT|31|3|耶和華－你的上帝必在你面前過河，把這些國從你面前除滅，你就必得他們的地。 約書亞 要在你面前過河，是照耶和華所吩咐的。
DEUT|31|4|耶和華必對待他們，如同從前待他所除滅的 亞摩利 人的王 西宏 與 噩 ，以及他們的國一樣。
DEUT|31|5|耶和華必將他們交在你們面前，你們要照我所吩咐的一切命令待他們。
DEUT|31|6|你們當剛強壯膽，不要害怕，也不要畏懼他們，因為耶和華－你的上帝必與你同去；他必不撇下你，也不丟棄你。」
DEUT|31|7|摩西 召了 約書亞 來，在 以色列 眾人眼前對他說：「你當剛強壯膽！因為你要和這百姓一同進入 耶和華向他們列祖起誓要給他們的地，你也要使他們承受那地為業。
DEUT|31|8|耶和華必在你前面行，他必親自與你同在，必不撇下你，也不丟棄你。你不要懼怕，也不要驚惶。」
DEUT|31|9|摩西 寫下這律法，交給抬耶和華約櫃的 利未 人祭司和 以色列 的眾長老。
DEUT|31|10|摩西 吩咐他們說：「每逢七年的最後一年，就是定期的豁免年，在住棚節的時候，
DEUT|31|11|當 以色列 眾人來到耶和華－你上帝所選擇的地方朝見他的時候，你要在 以色列 眾人面前念這律法給他們聽。
DEUT|31|12|要召集百姓，男人、女人、孩子，和在你城裏寄居的，叫他們都得以聽見，好學習敬畏耶和華－你們的上帝，謹守遵行這律法的一切話。
DEUT|31|13|他們的兒女，就是那未曾認識的，也可以聽，學習敬畏耶和華－你們的上帝；你們一生的日子，在你們過 約旦河 得為業的地上，都要這樣做。」
DEUT|31|14|耶和華對 摩西 說：「看哪，你的死期已近了。要召 約書亞 來，和你一起站在會幕裏，我好吩咐他。」於是 摩西 和 約書亞 去站在會幕裏。
DEUT|31|15|耶和華在會幕裏，在雲柱中顯現，雲柱停在會幕門口的上面。
DEUT|31|16|耶和華對 摩西 說：「看哪，你必和你的祖先同睡。這百姓要起來，在他們所要去的地上，在那地的人中，隨從外邦的神明行淫，離棄我，違背我與他們所立的約。
DEUT|31|17|那時，我的怒氣必向他們發作，我必離棄他們，轉臉不顧他們，以致他們被吞滅，並有許多的禍患災難臨到他們。在那日，人必說：『這些禍患臨到我，豈不是因為我的上帝不在我中間嗎？』
DEUT|31|18|在那日，因人偏向別神所行的一切惡事，我必定轉臉不顧。
DEUT|31|19|現在你們要寫下這首歌，教導 以色列 人，放在他們口中，使這首歌成為我指責 以色列 人的見證。
DEUT|31|20|因為我將他們領進我向他們列祖起誓應許那流奶與蜜之地，他們在那裏吃得飽足，長得肥胖，就偏向別神，事奉它們，藐視我，背棄我的約。
DEUT|31|21|當許多禍患災難臨到他們的時候，這首歌必在他們面前作見證，因為他們後裔的口必吟誦不忘。我未領他們到我所起誓應許之地以先，他們所懷的意念我都知道了。」
DEUT|31|22|當日 摩西 就寫了一首歌，教導 以色列 人。
DEUT|31|23|耶和華吩咐 嫩 的兒子 約書亞 說：「你當剛強壯膽，因為你必領 以色列 人進入我所起誓應許他們的地，我必與你同在。」
DEUT|31|24|當 摩西 把這律法的話寫完在書上，到完成的時候，
DEUT|31|25|摩西 吩咐抬耶和華約櫃的 利未 人說：
DEUT|31|26|「把這律法書拿來，放在耶和華－你們上帝的約櫃旁，可以在那裏作指責你們的見證。
DEUT|31|27|因為我知道你們是悖逆的，是硬著頸項的。看哪，我今日還活著與你們同在，你們尚且悖逆耶和華，何況我死後呢？
DEUT|31|28|你們要召集你們支派的眾長老和官長到我這裏來，我好把這些話說給他們聽，並且呼喚天地見證他們的不是。
DEUT|31|29|我知道我死後你們必全然敗壞，偏離我所吩咐你們的道。日後必有禍患臨到你們，因為你們做了耶和華眼中看為惡的事，以你們手中所做的惹他發怒。」
DEUT|31|30|摩西 把這首歌的話，從頭到尾吟誦給 以色列 全會眾聽。
DEUT|32|1|「諸天哪，要側耳聽我說話； 願地聆聽我口中的言語。
DEUT|32|2|我的教導要淋漓如雨， 我的言語要滴落如露， 如細雨降在嫩草上， 如甘霖降在蔬菜中。
DEUT|32|3|因為我要宣揚耶和華的名， 你們要把偉大歸給我們的上帝。
DEUT|32|4|「他是磐石，他的作為完全， 他一切所行的都公平； 他是信實無偽的上帝， 又公義，又正直。
DEUT|32|5|這乖僻彎曲的世代 向他行了敗壞的事； 因著他們的弊病， 不再是他的兒女。
DEUT|32|6|愚昧無知的百姓啊， 你們這樣報答耶和華嗎？ 他豈不是你的父，創造了你嗎？ 他造了你，堅立你。
DEUT|32|7|你當回想上古之日， 思念歷代之年； 問你的父親，他必告訴你； 問你的長者，他必向你述說。
DEUT|32|8|至高者將地業賜給列國， 將世人分開， 他按照神明 的數目， 為萬民劃定疆界。
DEUT|32|9|因為耶和華的份是他的百姓， 他的產業就是 雅各 。
DEUT|32|10|「耶和華在曠野之地， 在空曠，野獸吼叫之荒地遇見他， 就環繞他，看顧他， 保護他，如同保護眼中的瞳人。
DEUT|32|11|鷹怎樣攪動巢窩， 在雛鷹上面飛翔， 展開雙翅接住雛鷹， 背在兩翼之上，
DEUT|32|12|耶和華也照樣獨自引導他， 並無外邦神明與他同在。
DEUT|32|13|耶和華使他馳騁在地的高處， 他吃田間的出產； 耶和華使他從巖石中吃蜜， 從堅石中吸油，
DEUT|32|14|也吃牛的乳酪、羊的奶、 羔羊的脂肪， 巴珊 所出的公綿羊和山羊， 和上好的麥子。 你要喝葡萄汁釀的美酒。
DEUT|32|15|「 耶書崙 漸漸肥胖，能踼跳。 你長得肥胖，粗壯，豐潤。 他離棄造他的上帝， 輕看救他的磐石。
DEUT|32|16|他們用外邦神明惹上帝妒忌， 以可憎之物惹他發怒。
DEUT|32|17|他們祭祀鬼魔，而非上帝， 是他們不認識的神明， 是近來新興的， 是你們列祖所不畏懼的。
DEUT|32|18|你輕忽生你的磐石， 忘記生產你的上帝。
DEUT|32|19|「耶和華看見了， 因他兒女惹動他就拋棄他們，
DEUT|32|20|說：『我要轉臉離開他們， 看他們的結局如何。 他們是極乖謬的世代， 是不忠實的兒女。
DEUT|32|21|他們以那不是上帝的激起我妒忌， 以虛無的神明 惹我發怒。 我也要以不成國的激起你們嫉妒， 我要以愚頑的國惹起你們發怒。
DEUT|32|22|因為我的怒火焚燒， 直燒到極深的陰間， 吞噬地和地的出產， 連山的根基也燒著了。
DEUT|32|23|「『我要把禍患堆在他們身上， 我用盡我的箭射向他們：
DEUT|32|24|餓死人的饑荒、 灼人的熱症、 痛苦的災害。 我要叫野獸用牙齒咬他們， 叫土中爬行的用毒液害他們。
DEUT|32|25|外有刀劍使人喪亡， 內有驚恐， 少男少女是如此， 吃奶的、白髮的也是如此。
DEUT|32|26|我曾說，我要粉碎他們， 使他們的名 從人間消失。
DEUT|32|27|惟恐仇敵挑釁， 他們的敵人誤解， 說，我們的手得勝了， 這一切並非耶和華做的。』
DEUT|32|28|「因為他們是缺乏智謀的國家， 他們裏面毫無聰明。
DEUT|32|29|惟願他們有智慧，能明白這事， 他們就會想到自己的結局。
DEUT|32|30|若非他們的磐石賣了他們， 若非耶和華交出他們， 一人豈能追趕千人， 二人焉能使萬人逃跑呢？
DEUT|32|31|甚至我們的仇敵都承認， 他們的磐石不如我們的磐石。
DEUT|32|32|他們的葡萄樹是 所多瑪 的葡萄樹， 是 蛾摩拉 田園所長的； 他們的葡萄是毒葡萄， 整串都是苦的。
DEUT|32|33|他們的酒是大蛇的毒液， 是毒蛇劇烈的毒汁。
DEUT|32|34|「這豈不都存放在我這裏， 封存在我庫房中嗎？
DEUT|32|35|伸冤報應在我 ， 到了時候他們會失腳。 因為他們遭難的日子近了， 他們的厄運快要臨到。
DEUT|32|36|耶和華見他的百姓毫無能力， 無論是為奴的、自由的，都沒有存留， 就必為他們伸冤， 為自己的僕人發憐憫。
DEUT|32|37|他必說：『他們的神明， 他們所投靠的磐石，在哪裏呢？
DEUT|32|38|吃了他們祭牲脂肪的， 喝了他們澆酒祭之酒的， 叫那些神明站出來幫助你們， 作為你們的保障吧！
DEUT|32|39|「『如今，看！我，惟有我是上帝 ； 我以外並無別神。 我使人死，我使人活； 我擊傷人，也醫治人， 沒有人能從我手中救出來。
DEUT|32|40|我向天舉手， 我憑我的永生起誓說：
DEUT|32|41|我若磨我閃亮的刀， 我的手掌握審判權， 就必報復我的敵人， 報應那些恨我的人。
DEUT|32|42|我要使我的箭飲血而醉， 就是被殺被擄之人的血； 我的刀也要吃肉， 就是仇敵披髮頭顱 的肉。』
DEUT|32|43|「列國啊，當與耶和華的子民一同歡呼 ； 因為他要為他僕人 所流的血伸冤， 報應他的敵人 ， 救贖他的土地和他的子民 。」
DEUT|32|44|摩西 和 嫩 的兒子 約書亞 前來把這首歌的一切話吟誦給百姓聽。
DEUT|32|45|摩西 向 以色列 眾人吟誦完了這一切話，
DEUT|32|46|對他們說：「我今日以這一切話警戒你們，你們都要記在心中，要吩咐你們的子孫謹守遵行這律法上一切的話。
DEUT|32|47|因為這不是與你們無關的空話，而是你們的生命；因遵行這話，你們的日子必在你們過 約旦河 得為業的地上得以長久。」
DEUT|32|48|就在那日，耶和華吩咐 摩西 說：
DEUT|32|49|「你上 摩押 地的 亞巴琳山脈 ，到面對 耶利哥 的 尼波山 去，看我所要賜給 以色列 人為業的 迦南 地。
DEUT|32|50|你必死在你所登的山上，歸到你祖先 那裏，像你哥哥 亞倫 死在 何珥山 上，歸到他祖先 那裏一樣。
DEUT|32|51|因為你們在 以色列 人中得罪了我，在 尋 的曠野， 加低斯 的 米利巴 水那裏，在 以色列 人中沒有尊我為聖。
DEUT|32|52|我所賜給 以色列 人的地，你只可從對面觀看，卻不得進到那裏去。」
DEUT|33|1|這是神人 摩西 未死以前為 以色列 人的祝福。
DEUT|33|2|他說： 「耶和華從 西奈 來， 從 西珥 向他們顯現， 從 巴蘭山 發出光輝； 從萬萬聖者中來臨 ， 從他右手向他們發出烈火的律法 。
DEUT|33|3|他實在疼愛萬民。 他的眾聖徒都在你手中， 他們坐在你的腳下， 領受你的言語。」
DEUT|33|4|摩西 將律法傳給我們， 作為 雅各 會眾的產業。
DEUT|33|5|「耶和華 在 耶書崙 作王； 百姓的眾領袖和 以色列 各支派一同歡聚。
DEUT|33|6|願 呂便 存活，不致死亡， 雖然他的人丁稀少。
DEUT|33|7|關於 猶大 ，他這麼說： 『耶和華啊，求你垂聽 猶大 的聲音， 引導他歸回他的百姓中。 他曾用手為自己爭戰， 你必幫助他攻擊敵人。』
DEUT|33|8|關於 利未 ，他說： 『願你的土明和烏陵都在你的虔誠人那裏 。 你在 瑪撒 曾考驗他， 在 米利巴 水與他爭論。
DEUT|33|9|關於自己的父母，他說：我未曾關注。 他的弟兄，他不承認， 他的兒女，他也不認識， 因為 利未 人遵行你的話， 謹守你的約。
DEUT|33|10|他們將你的典章教導 雅各 ， 將你的律法教導 以色列 。 他們奉上香讓你聞， 把全牲的燔祭獻在你壇上。
DEUT|33|11|求耶和華賜福給他的財物 ， 悅納他手裏的工作。 求你刺透起來攻擊他的人的腰， 使那些恨惡他的人不再起來。』
DEUT|33|12|關於 便雅憫 ，他說： 『耶和華所親愛的必同耶和華安然居住， 耶和華終日庇護他， 他也住在耶和華兩肩之中 。』
DEUT|33|13|關於 約瑟 ，他說： 『願他的地蒙耶和華賜福， 得天上的甘露， 地下的泉源；
DEUT|33|14|得太陽下的美果， 月光中的佳穀；
DEUT|33|15|得古老山嶽的至寶， 永恆山嶺的寶物；
DEUT|33|16|得地的寶物和其中所充滿的， 得住在荊棘中者的喜悅。 願這些福都臨到 約瑟 的頭上， 臨到那與兄弟有分別之人的頭頂上。
DEUT|33|17|他是牛群中頭生的， 大有威嚴； 他的雙角是野牛的角， 用以牴觸萬民，直到地極。 這對角是 以法蓮 的萬萬， 這對角是 瑪拿西 的千千。』
DEUT|33|18|關於 西布倫 ，他說： 『 西布倫 哪，你出外可以歡喜。 以薩迦 啊，你在帳棚裏可以快樂。
DEUT|33|19|他們要召集萬民到山上， 在那裏獻公義的祭。 因為他們要吸取海裏的財富， 沙中隱藏的珍寶。』
DEUT|33|20|關於 迦得 ，他說： 『那使 迦得 擴張的，當受稱頌！ 迦得 臥如母獅， 撕裂膀臂和頭皮。
DEUT|33|21|他為自己看中了最好的， 因為那是為掌權者所存留的一份。 他與百姓的領袖同來 ， 執行耶和華的公義 和耶和華為 以色列 所立的典章。』
DEUT|33|22|關於 但 ，他說： 『 但 是小獅子， 從 巴珊 跳出來。』
DEUT|33|23|關於 拿弗他利 ，他說： 『 拿弗他利 啊，你享足恩寵， 滿得耶和華的福， 可以得西方和南方為業。』
DEUT|33|24|關於 亞設 ，他說： 『願 亞設 在眾子中蒙福 ， 願他得他弟兄的喜悅， 可以把腳蘸在油中。
DEUT|33|25|你的門閂是鐵的，是銅的。 只要你有多少日子，你就有多少力量 。』
DEUT|33|26|「 耶書崙 哪，沒有誰能比上帝！ 他騰雲，大顯威榮， 從天空來幫助你。
DEUT|33|27|亙古的上帝是避難所， 下面有永久的膀臂。 他從你面前趕走仇敵， 說：『毀滅吧！』
DEUT|33|28|因此， 以色列 獨自安然居住， 雅各 的泉源在五穀新酒之地， 他的天也滴下露水。
DEUT|33|29|以色列 啊，你有福了！ 蒙耶和華拯救的百姓啊，誰能像你？ 他是幫助你的盾牌， 是你威榮的刀劍。 你的仇敵要屈身就你； 你卻要踐踏他們的背脊 。」
DEUT|34|1|摩西 從 摩押 平原登上 尼波山 ，到了 耶利哥 對面的 毗斯迦山 頂。耶和華把全地指給他看：從 基列 到 但 ，
DEUT|34|2|拿弗他利 全地， 以法蓮 、 瑪拿西 的地， 猶大 全地直到西邊的海，
DEUT|34|3|尼革夫 ，從棕樹城 耶利哥 的平原到 瑣珥 。
DEUT|34|4|耶和華對他說：「這就是我向 亞伯拉罕 、 以撒 、 雅各 起誓應許之地，說：『我必將這地賜給你的後裔。』現在我使你親眼看見了，你卻不得過到那裏去。」
DEUT|34|5|於是耶和華的僕人 摩西 死在 摩押 地那裏，正如耶和華所說的。
DEUT|34|6|耶和華將他葬在 摩押 地， 伯‧毗珥 對面的谷中，只是到今日，沒有人知道他的墳墓。
DEUT|34|7|摩西 死的時候一百二十歲，眼目沒有昏花，力量沒有衰退。
DEUT|34|8|以色列 人在 摩押 平原為 摩西 哀哭了三十天，為 摩西 哀哭居喪的日期才結束。
DEUT|34|9|嫩 的兒子 約書亞 ，因為 摩西 曾為他按手，他就被智慧的靈充滿。 以色列 人聽從他，照著耶和華所吩咐 摩西 的去做。
DEUT|34|10|以後， 以色列 中再沒有興起一位先知像 摩西 的，他是耶和華面對面所認識的。
DEUT|34|11|耶和華差派他在 埃及 地，向法老和他的一切臣僕，以及他的全地，行了各樣神蹟奇事，
DEUT|34|12|又在 以色列 眾人眼前顯出大能的手，行了一切大而可畏的事。
JOSH|1|1|耶和華的僕人 摩西 死了以後，耶和華對 摩西 的助手 嫩 的兒子 約書亞 說：
JOSH|1|2|「我的僕人 摩西 死了。現在你要起來，和眾百姓過這 約旦河 ，往我所要賜給 以色列 人的地去。
JOSH|1|3|凡你們腳掌所踏之地，我都照我所應許 摩西 的話賜給你們了。
JOSH|1|4|從曠野和這 黎巴嫩 ，直到 大河 ，就是 幼發拉底河 ， 赫 人的全地，又到 大海 日落的方向，都要作你們的疆土。
JOSH|1|5|你一生的日子，必無人能在你面前站立得住。我怎樣與 摩西 同在，也必照樣與你同在；我必不撇下你，也不丟棄你。
JOSH|1|6|你當剛強壯膽，因為你必使這百姓承受那地為業，就是我向他們列祖起誓要給他們的地。
JOSH|1|7|只要剛強，大大壯膽，謹守遵行我僕人 摩西 所吩咐你的一切律法，不可偏離左右，使你無論往哪裏去， 都可以順利。
JOSH|1|8|這律法書不可離開你的口，總要晝夜思想 ，好使你謹守遵行這書上所寫的一切話。如此，你的道路就可以亨通，凡事順利。
JOSH|1|9|我豈沒有吩咐你嗎？你當剛強壯膽，不要懼怕，也不要驚惶，因為你無論往哪裏去，耶和華你的上帝必與你同在。」
JOSH|1|10|於是， 約書亞 吩咐百姓的官長說：
JOSH|1|11|「你們要走遍營中，吩咐百姓說：『當預備食物， 因為三日之內你們要過這 約旦河 ，進去得耶和華－你們上帝賜給你們為業之地。』」
JOSH|1|12|約書亞 對 呂便 人、 迦得 人和 瑪拿西 半支派的人說：
JOSH|1|13|「你們要記得耶和華的僕人 摩西 所吩咐你們的話說：『耶和華－你們的上帝使你們得享安寧，必將這地賜給你們。』
JOSH|1|14|你們的妻子、孩子和牲畜可以留在 約旦河 東、 摩西 所給你們的地。但你們中間所有大能的勇士都要帶著兵器，在你們的弟兄前面過去，你們要幫助他們。
JOSH|1|15|等到耶和華使你們的弟兄和你們一樣得享平靜，並且得著耶和華－你們上帝所賜他們為業之地的時候，你們才可以回到你們所得之地，承受為業，就是耶和華的僕人 摩西 在 約旦河 東、向日出的方向所給你們的地。」
JOSH|1|16|他們回答 約書亞 說：「凡你吩咐我們的，我們都必做；凡你差我們去的地方，我們都必去。
JOSH|1|17|我們在一切事上怎樣聽從 摩西 ，也必照樣聽從你。惟願耶和華－你的上帝與你同在，像與 摩西 同在一樣。
JOSH|1|18|無論甚麼人違背你的命令，不聽從你所吩咐他的一切話，就必處死。你只要剛強壯膽！」
JOSH|2|1|嫩 的兒子 約書亞 從 什亭 暗中派兩個人作探子，說：「你們去窺探那地和 耶利哥 。」於是二人去了，來到一個名叫 喇合 的妓女家裏，在那裏睡覺。
JOSH|2|2|有人告訴 耶利哥 王說：「看哪，今夜有 以色列 人到這裏來窺探此地。」
JOSH|2|3|耶利哥 王派人到 喇合 那裏， 說：「你要交出那來到你這裏、進了你家的人，因為他們來是要窺探全地。」
JOSH|2|4|但女人已把二人藏起來，卻說：「那兩個人確實到我這裏來過，他們從哪裏來，我卻不知道。
JOSH|2|5|天黑、要關城門的時候，他們就出去了。他們往哪裏去我也不知道。你們趕快去追他們，就必追上。」
JOSH|2|6|其實，這女人已經領二人上了屋頂，把他們藏在她擺列在屋頂的的亞麻梗中。
JOSH|2|7|那些人就往 約旦河 的路上追趕他們，直到渡口。追趕他們的人一出去，城門就關了。
JOSH|2|8|二人還沒有睡之前，女人就上屋頂，到他們那裏，
JOSH|2|9|對他們說：「我知道耶和華已經把這地賜給你們了，並且我們也都懼怕你們。這地所有的居民在你們面前都融化了。
JOSH|2|10|因為我們聽見你們出 埃及 的時候，耶和華怎樣在你們前面使 紅海 的水乾了，並且你們怎樣處置 約旦河 東的兩個 亞摩利 王， 西宏 和 噩 ，把他們完全消滅。
JOSH|2|11|我們一聽見就膽戰心驚 ，人人因你們的緣故勇氣全失。耶和華－你們的上帝是天上地下的上帝。
JOSH|2|12|現在我既然恩待你們，求你們指著耶和華向我起誓，你們也要恩待我的父家。請你們給我一個確實的憑據，
JOSH|2|13|要救活我的父母、兄弟、姊妹，和所有屬他們的，拯救我們的性命脫離死亡。」
JOSH|2|14|那二人對她說：「我們願意以性命來替你們死。你們若不洩漏我們這件事，當耶和華將這地賜給我們的時候，我們必以慈愛和誠信待你。」
JOSH|2|15|於是女人用繩子把二人從窗戶縋下去，因為她的屋子是在城牆邊上，她也住在城牆上。
JOSH|2|16|她對他們說：「你們暫且往山上去，免得追趕的人遇見你們。要在那裏躲藏三天，等追趕的人回來，你們才可以走自己的路。」
JOSH|2|17|二人對她說：「你叫我們所起的誓與我們無關，
JOSH|2|18|除非，看哪，當我們來到這地的時候，你把這條朱紅線繩子繫在縋我們下去的窗戶上，並要叫你的父母、兄弟和你父的全家都聚集在你家中。
JOSH|2|19|凡離開你家門往街上去的，他的血必歸到自己頭上，與我們無關；凡在你家裏的，若有人下手害他，他的血就歸到我們頭上。
JOSH|2|20|你若洩漏我們這件事，你叫我們所起的誓 就與我們無關了。」
JOSH|2|21|女人說：「就照你們的話吧！」於是她送他們走了，就把朱紅繩子繫在窗戶上。
JOSH|2|22|二人離開，到山上去，在那裏停留三天，直等到追趕的人回去。追趕的人一路尋找，卻找不著。
JOSH|2|23|二人回來，下了山，過了河，來到 嫩 的兒子 約書亞 那裏，向他報告他們所遭遇的一切事。
JOSH|2|24|他們對 約書亞 說：「耶和華果然將那全地交在我們手中了，並且那地所有的居民在我們面前都融化了。」
JOSH|3|1|約書亞 清早起來，和 以色列 眾人起行，離開 什亭 ，來到 約旦河 ，過河以前住在那裏。
JOSH|3|2|過了三天，官長走遍營中，
JOSH|3|3|吩咐百姓說：「當你們看見 利未 家的祭司抬著耶和華－你們上帝的約櫃的時候，你們就要起行離開所住的地方，跟著約櫃走，
JOSH|3|4|使你們知道所當走的路，因為這條路是你們從來沒有走過的。只是你們要與約櫃相隔約二千肘，不可太靠近約櫃。」
JOSH|3|5|約書亞 吩咐百姓說：「你們要使自己分別為聖，因為明天耶和華必在你們中間行奇事。」
JOSH|3|6|約書亞 對祭司說：「你們抬起約櫃，在百姓的前面過去。」於是他們抬起約櫃，走在百姓前面。
JOSH|3|7|耶和華對 約書亞 說：「從今日起，我必使你在 以色列 眾人眼前被尊為大，使他們知道我怎樣與 摩西 同在，也必照樣與你同在。
JOSH|3|8|你要吩咐抬約櫃的祭司說：『你們到了 約旦河 的水邊，要在 約旦河 中站著。』」
JOSH|3|9|約書亞 對 以色列 人說：「你們近前，到這裏來，聽耶和華－你們上帝的話。」
JOSH|3|10|約書亞 說：「你們因這事會知道永生的上帝在你們中間，他必從你們面前趕出 迦南 人、 赫 人、 希未 人、 比利洗 人、 革迦撒 人、 亞摩利 人、 耶布斯 人。
JOSH|3|11|看哪！全地之主的約櫃必在你們的前面過去，到 約旦河 裏。
JOSH|3|12|現在， 你們要從 以色列 支派中選出十二個人，每支派一人。
JOSH|3|13|當抬耶和華全地之主約櫃的祭司，腳掌踏入 約旦河 水裏的時候， 約旦河 的水，就是從上往下流的水，必然中斷，豎立成壘。」
JOSH|3|14|百姓起行離開帳棚過 約旦河 的時候，抬約櫃的祭司在百姓的前面。
JOSH|3|15|那時正是收割的日子， 約旦河 的水漲滿兩岸。抬約櫃的人到了 約旦河 ，抬約櫃的祭司腳一入水邊，
JOSH|3|16|那從上往下流的水就在很遠的地方，在 撒拉但 旁邊的 亞當城 那裏停住，豎立成壘；那往 亞拉巴海 ，就是 鹽海 下流的水全然中斷。於是，百姓在 耶利哥 的對面過了河。
JOSH|3|17|抬耶和華約櫃的祭司在 約旦河 中的乾地上穩穩站著， 以色列 眾人都從乾地上過去，直到全國都過了 約旦河 。
JOSH|4|1|當全國都過了 約旦河 ，耶和華對 約書亞 說：
JOSH|4|2|「你要從百姓中選出十二個人，每支派一人，
JOSH|4|3|吩咐他們說：『你們從這裏，從 約旦河 中祭司的腳穩穩站立的地方，取十二塊石頭 ，一起帶過去，放在你們今夜住宿的地方。』」
JOSH|4|4|於是 約書亞 召集了他從 以色列 人中所選的十二個人，每支派一人。
JOSH|4|5|約書亞 對他們說：「你們要過去，到 約旦河 中，耶和華－你們上帝的約櫃前面，按 以色列 人支派的數目，每人各取一塊石頭扛在肩上。
JOSH|4|6|這些石頭在你們中間將成為記號。日後，你們的子孫問你們說：『這些石頭對你們有甚麼意思呢？』
JOSH|4|7|你們就對他們說：『這是因為 約旦河 的水在耶和華的約櫃前中斷；約櫃過 約旦河 的時候， 約旦河 的水就中斷了。這些石頭要作 以色列 人永遠的紀念。』」
JOSH|4|8|以色列 人就照 約書亞 所吩咐的做了。他們按 以色列 人支派的數目，從 約旦河 中取了十二塊石頭，正如耶和華所吩咐 約書亞 的。他們把石頭帶過去，到他們所住宿的地方，就放在那裏。
JOSH|4|9|約書亞 另外把十二塊石頭立在 約旦河 的中間，在抬約櫃祭司的腳站立的地方；直到今日，石頭還在那裏。
JOSH|4|10|抬約櫃的祭司站在 約旦河 的中間，直到耶和華命令 約書亞 告訴百姓的一切事辦完為止，正如 摩西 所吩咐 約書亞 的一切話。 於是，百姓急速過了河。
JOSH|4|11|全體百姓都過了河之後，耶和華的約櫃和祭司才過去，到百姓的前面。
JOSH|4|12|呂便 人、 迦得 人、 瑪拿西 半支派的人都照 摩西 所吩咐他們的，帶著兵器在 以色列 人的前面過去。
JOSH|4|13|約有四萬帶兵器的軍隊在耶和華面前過去，到 耶利哥 的平原，準備上陣。
JOSH|4|14|在那日，耶和華使 約書亞 在 以色列 眾人眼前被尊為大。在他一生的年日中，百姓敬服他，像從前敬服 摩西 一樣。
JOSH|4|15|耶和華對 約書亞 說：
JOSH|4|16|「你吩咐抬法櫃的祭司從 約旦河 上來。」
JOSH|4|17|約書亞 就吩咐祭司說：「你們從 約旦河 上來。」
JOSH|4|18|抬耶和華約櫃的祭司從 約旦河 中上來，腳掌一落乾地， 約旦河 的水就流回原處，仍舊漲滿兩岸。
JOSH|4|19|正月初十，百姓從 約旦河 上來，就在 耶利哥 東邊的 吉甲 安營。
JOSH|4|20|約書亞 把他們從 約旦河 取來的那十二塊石頭立在 吉甲 ，
JOSH|4|21|對 以色列 人說：「日後，你們的子孫問他們的父親說：『這些石頭是甚麼意思呢？』
JOSH|4|22|你們就讓你們的子孫知道，說：『 以色列 人曾走乾地過這 約旦河 。』
JOSH|4|23|因為耶和華－你們的上帝在你們前面使 約旦河 的水乾了，直到你們過來，就如耶和華－你們的上帝從前在我們前面使 紅海 乾了，直到我們過來一樣，
JOSH|4|24|要使地上萬民都知道，耶和華的手大有能力，也要使你們天天敬畏耶和華－你們的上帝。」
JOSH|5|1|約旦河 西 亞摩利 人的眾王和靠海 迦南 人的眾王，聽見耶和華在 以色列 人前面使 約旦河 的水乾了，直到他們過了河 ，眾王因 以色列 人的緣故都膽戰心驚，勇氣全失。
JOSH|5|2|那時，耶和華對 約書亞 說：「你要造火石刀，第二次為 以色列 人行割禮。」
JOSH|5|3|約書亞 就造了火石刀，在 哈爾拉勒山 為 以色列 人行割禮。
JOSH|5|4|約書亞 行割禮的原因是這樣：從 埃及 出來的眾百姓，所有能打仗的男丁，出了 埃及 以後，都死在曠野的路上。
JOSH|5|5|這些從 埃及 出來的眾百姓都受過割禮；但是那些出 埃及 以後，在曠野的路上所生的眾百姓卻沒有受過割禮。
JOSH|5|6|以色列 人在曠野走了四十年，直到那從 埃及 出來，全國能打仗的人都消滅了，因為他們沒有聽從耶和華的話。耶和華曾向他們起誓，必不容許他們看見耶和華向他們列祖起誓要給我們的地，就是流奶與蜜之地。
JOSH|5|7|他們的子孫，就是耶和華興起接續他們的，都沒有受過割禮；因為在路上他們沒有受割禮， 約書亞 就為他們行割禮。
JOSH|5|8|全國的人都受了割禮，留在營中自己的地方，直到痊癒。
JOSH|5|9|耶和華對 約書亞 說：「我今日將 埃及 的羞辱從你們身上除掉了。」因此，那地方名叫 吉甲 ，直到今日。
JOSH|5|10|以色列 人在 吉甲 安營。正月十四日晚上，他們在 耶利哥 的平原守逾越節。
JOSH|5|11|逾越節的第二日，他們吃了當地的出產，就在那一天，吃了無酵餅和烘過的穀物。
JOSH|5|12|他們吃了當地出產的第二日，嗎哪就停止了。 以色列 人不再有嗎哪了。那一年，他們就吃 迦南 地的出產。
JOSH|5|13|約書亞 靠近 耶利哥 的時候，舉目觀看，看哪，有一個人站在他對面，手裏拿著拔出來的刀。 約書亞 到他那裏，對他說：「你是屬我們的，還是屬我們敵人的呢？」
JOSH|5|14|他說：「不，我現在來是要作耶和華軍隊的元帥。」 約書亞 就臉伏於地下拜，說：「我主有甚麼話，請吩咐僕人吧！」
JOSH|5|15|耶和華軍隊的元帥對 約書亞 說：「把你腳上的鞋脫下來，因為你所站的地方是聖的。」 約書亞 就照著做了。
JOSH|6|1|耶利哥 的城門因 以色列 人的緣故，關得嚴緊，無人出入。
JOSH|6|2|耶和華對 約書亞 說：「看，我已經把 耶利哥城 和 耶利哥 王，以及大能的勇士，都交在你手中。
JOSH|6|3|你們要圍繞這城，所有的士兵繞城一次，六日你都要這樣做。
JOSH|6|4|七個祭司要拿七個羊角走在約櫃前。到了第七日，你們要圍繞這城七次，祭司也要吹角。
JOSH|6|5|羊角聲拖長的時候，你們一聽見角聲，眾百姓要大聲呼喊，城牆就必倒塌，各人要往前直上。」
JOSH|6|6|嫩 的兒子 約書亞 召了祭司來，對他們說：「你們抬起約櫃來，要有七個祭司拿七個羊角在耶和華的約櫃前。」
JOSH|6|7|他又對百姓說：「你們向前去圍繞那城，帶兵器的要在耶和華的約櫃前過去。」
JOSH|6|8|按照 約書亞 對百姓所說的，七個祭司拿了七個羊角在耶和華面前過去，他們吹著角，耶和華的約櫃在他們後面跟著。
JOSH|6|9|帶兵器的走在吹角的祭司前面，後隊跟著約櫃走，號角繼續在吹。
JOSH|6|10|約書亞 吩咐百姓說：「你們不可呼喊，不可讓人聽見你們的聲音，連一句話也不可出你們的口，直到我對你們說『呼喊』的那日，你們才呼喊。」
JOSH|6|11|這樣， 約書亞 使耶和華的約櫃圍繞那城，把城繞了一次。然後，眾人回到營裏，就在營裏住宿。
JOSH|6|12|約書亞 清早起來，祭司又抬起耶和華的約櫃。
JOSH|6|13|七個祭司拿七個羊角，走在耶和華的約櫃前，他們吹著角；帶兵器的走在他們前面，後隊跟著耶和華的約櫃走，號角繼續在吹。
JOSH|6|14|第二日，他們再把城圍繞一次，就回營裏去。六日都是這樣做。
JOSH|6|15|第七日清早黎明時，他們起來，以同樣的方式圍繞城七次；惟獨這一日他們圍繞城七次。
JOSH|6|16|到了第七次，祭司吹角的時候， 約書亞 對百姓說：「呼喊吧，因為耶和華已經把城交給你們了！
JOSH|6|17|這城和其中所有的都要永獻給耶和華作當毀滅的，只有妓女 喇合 與她家中所有的可以存活，因為她隱藏了我們所派的使者。
JOSH|6|18|但你們務必謹慎，不可取那當滅的物，免得你們受詛咒，取了那當滅的物，使 以色列 全營成為詛咒而遭受災禍。
JOSH|6|19|只有金子、銀子和銅鐵的器皿都要歸耶和華為聖，放入耶和華的庫房中。」
JOSH|6|20|於是百姓呼喊，祭司吹角。百姓一聽見角聲就大聲呼喊，城牆隨著倒塌。百姓上去進城，各人往前直上，把城奪取。
JOSH|6|21|他們把城中所有的，無論男女老少，牛羊和驢，都用刀殺盡。
JOSH|6|22|約書亞 對窺探這地的兩個人說：「你們進那妓女的家，照你們向她所起的誓，將那女人和她所有的都從那裏帶出來。」
JOSH|6|23|兩個作過探子的青年進去，把 喇合 與她的父母、兄弟，和她所有的帶出來，他們把她所有的親屬都帶出來，安置在 以色列 的營外。
JOSH|6|24|他們用火焚燒了那城和其中所有的，只有金子、銀子和銅鐵的器皿都放在耶和華殿的庫房中。
JOSH|6|25|至於妓女 喇合 和她父家，以及她所有的， 約書亞 保存了他們的性命。她就住在 以色列 中，直到今日，因為她隱藏了 約書亞 派來窺探 耶利哥 的使者。
JOSH|6|26|當時， 約書亞 叫眾人起誓說：「凡興起重修這 耶利哥城 的，當在耶和華面前受詛咒。 他立根基的時候，必喪長子， 安城門的時候，必喪幼子。」
JOSH|6|27|耶和華與 約書亞 同在， 約書亞 的名聲傳遍全地。
JOSH|7|1|以色列 人在當滅之物上犯了罪。 猶大 支派中， 謝拉 的曾孫， 撒底 的孫子， 迦米 的兒子 亞干 取了當滅之物，耶和華的怒氣就向 以色列 人發作。
JOSH|7|2|約書亞 從 耶利哥 派人往 伯特利 東邊，靠近 伯‧亞文 的 艾城 去，對他們說：「你們上去窺探那地。」那些人就上去窺探 艾城 。
JOSH|7|3|他們回到 約書亞 那裏，對他說：「眾百姓不必都上去，只要二、三千人上去就能攻取 艾城 ；不必勞動眾百姓都上去，因為他們人少。」
JOSH|7|4|於是百姓中約有三千人上那裏去，但他們竟在 艾城 的人面前逃跑。
JOSH|7|5|艾城 的人擊殺他們約三十六人，從城門前追趕他們，直到 示巴琳 ，在下坡的地方擊敗他們。他們都膽戰心驚，融化如水。
JOSH|7|6|約書亞 和 以色列 的長老就撕裂衣服，在耶和華的約櫃前臉伏於地，直到晚上。他們把灰撒在頭上。
JOSH|7|7|約書亞 說：「唉！主耶和華啊，你為甚麼領這百姓過 約旦河 ，把我們交在 亞摩利 人手中，使我們滅亡呢？我們不如住在 約旦河 的那邊！
JOSH|7|8|主啊，求求你， 以色列 人既在仇敵面前轉身逃跑，我還有甚麼可說的呢？
JOSH|7|9|迦南 人和這地所有的居民聽見了就必圍困我們，把我們的名從地上除去。那時，你為你至大的名要怎樣做呢？」
JOSH|7|10|耶和華對 約書亞 說：「起來！你的臉為何這樣俯伏呢？
JOSH|7|11|以色列 犯了罪，又違背了我所吩咐他們的約，又取了當滅之物。他們又偷竊，又行詭詐，又把那當滅的物與自己的器皿放在一起。
JOSH|7|12|因此， 以色列 人在仇敵面前站立不住。他們在仇敵面前轉身逃跑，因為他們成了當滅的物。你們若不把當滅的物從你們中間除掉，我就不再與你們同在了。
JOSH|7|13|你起來，去叫百姓分別為聖，說：『你們要為了明天使自己分別為聖，因為耶和華－ 以色列 的上帝這樣說： 以色列 啊，在你中間有當滅的物；你們若不把你們中間當滅之物除掉，你在仇敵面前必站立不住！』
JOSH|7|14|到了早晨，你們要按著支派近前來。耶和華所選的支派，要按著宗族近前來；耶和華所選的宗族，要按著家族近前來；耶和華所選的家族，要按著男丁，一個一個近前來。
JOSH|7|15|被選的人有當滅之物在他那裏，他和他所有的必被火焚燒，因為他違背了耶和華的約，又因他在 以色列 中做了愚妄的事。」
JOSH|7|16|於是， 約書亞 清早起來，召 以色列 按著支派近前來。選出來的是 猶大 支派。
JOSH|7|17|他召 猶大 的宗族近前來，選出來的是 謝拉 宗族。他召 謝拉 宗族，按著男丁 ，一個一個近前來，選出來的是 撒底 。
JOSH|7|18|他召 撒底 的家族，按著男丁，一個一個近前來，就選出 猶大 支派， 謝拉 的曾孫， 撒底 的孫子， 迦米 的兒子 亞干 。
JOSH|7|19|約書亞 對 亞干 說：「我兒，我勸你將榮耀歸給耶和華－ 以色列 的上帝，在他面前認罪，把你所做的事告訴我，不可向我隱瞞。」
JOSH|7|20|亞干 回答 約書亞 說：「我實在得罪了耶和華－ 以色列 的上帝。這是我所做的：
JOSH|7|21|我在所奪取的財物中看見一件美好的 示拿 外袍，二百舍客勒銀子，一條重五十舍客勒的金子。我貪愛這些物件，就拿去了。看哪，這些東西都埋在我帳棚內的地裏，銀子在外袍底下。」
JOSH|7|22|約書亞 就派使者跑到 亞干 的帳棚裏。看哪，那件外袍藏在他的帳棚裏，銀子在外袍底下。
JOSH|7|23|他們從帳棚裏把這些東西取出來，拿到 約書亞 和 以色列 眾人 那裏，倒在耶和華面前。
JOSH|7|24|約書亞 和 以色列 眾人把 謝拉 的曾孫 亞干 和那銀子、那件外袍、那條金子，以及 亞干 的兒女、牛、驢、羊、帳棚，和他所有的，都帶著上到 亞割谷 去。
JOSH|7|25|約書亞 說：「你為甚麼給我們招惹災禍呢？今日耶和華必使你遭受災禍。」於是 以色列 眾人用石頭打死他，用火焚燒他們，把石頭扔在其上。
JOSH|7|26|眾人在 亞干 身上堆了一大堆石頭，直存到今日。於是耶和華轉意，不發他的烈怒。因此，那地方名叫 亞割谷 ，直到今日。
JOSH|8|1|耶和華對 約書亞 說：「不要懼怕，也不要驚惶。你起來，率領所有作戰的士兵上 艾城 去。看，我已經把 艾城 的王和他的百姓、他的城，以及他的地，都交在你手裏。
JOSH|8|2|你怎樣處置 耶利哥 和 耶利哥 的王，也當照樣處置 艾城 和 艾城 的王。只是城內所奪的財物和牲畜，你們可以取為自己的掠物。你要在城的後面設下伏兵。
JOSH|8|3|於是， 約書亞 和所有作戰的士兵都起來，上 艾城 去。 約書亞 選了三萬大能的勇士，夜間派遣他們前去，
JOSH|8|4|吩咐他們說：「看，你們要在城的後面埋伏，不可離城太遠，各人都要準備。
JOSH|8|5|我與我所帶領的眾士兵要向城前進。城裏的人像上一次那樣出來迎擊我們的時候，我們就在他們面前逃跑。
JOSH|8|6|他們會出來追趕我們，直到我們引誘他們遠離那城。因為他們必說：『這些人像上次那樣在我們面前逃跑。』所以我們要在他們面前逃跑 。
JOSH|8|7|那時，你們就從埋伏的地方起來，奪取那城，因為耶和華－你們的上帝必把城交在你們的手裏。
JOSH|8|8|你們奪了城以後，要放火燒城，照耶和華的話去做。看，這是我吩咐你們的。」
JOSH|8|9|於是， 約書亞 派遣他們前去。他們行軍到埋伏的地方，伏在 伯特利 和 艾城 的中間，就是 艾城 的西邊。這夜， 約書亞 在士兵中間過夜。
JOSH|8|10|約書亞 清早起來，點齊士兵。他和 以色列 的長老在百姓前面上 艾城 去。
JOSH|8|11|所有跟他一起作戰的士兵都上去，向前逼近，來到城前，就在 艾城 北邊安營。 約書亞 與 艾城 之間隔著一個山谷。
JOSH|8|12|他選了約五千人，安排他們埋伏在 伯特利 和 艾城 的中間，就是 艾城 的西邊。
JOSH|8|13|於是，他們佈署軍隊，就是城北的全軍和城西的伏兵。當夜 約書亞 進入山谷之中。
JOSH|8|14|艾城 的王看見了，就和城裏的人清早起來，急忙出去，他和所有的士兵到了所定的地點，在 亞拉巴 前，迎擊 以色列 ，與之交戰；王並不知道城的後面有伏兵。
JOSH|8|15|約書亞 和 以色列 眾人在他們面前裝敗，往曠野的路逃跑。
JOSH|8|16|城內所有的百姓都被召來追趕他們。 艾城 的人追趕 約書亞 的時候，就被引誘遠離了城。
JOSH|8|17|艾城 和 伯特利 沒有一人不出來追趕 以色列 人的。他們撇下敞開的城門，去追趕 以色列 人。
JOSH|8|18|耶和華對 約書亞 說：「你向 艾城 伸出手裏的標槍，因為我要把那城交在你手裏。」 約書亞 就向那城伸出手裏的標槍。
JOSH|8|19|他一伸手，伏兵立刻從埋伏的地方衝出來，直攻入城，奪了它，立刻放火燒城。
JOSH|8|20|艾城 的人回頭，往後一看，看哪，城中煙氣沖天，他們向這邊或那邊都無處可逃。往曠野逃跑的百姓就轉身攻擊那些追趕他們的人。
JOSH|8|21|約書亞 和 以色列 眾人見伏兵已經奪了城，城中煙氣上騰，就轉身擊殺 艾城 的人。
JOSH|8|22|伏兵也出城追擊他們，他們就被 以色列 人前後夾攻，四面受敵。於是 以色列 人擊殺他們，沒有留下一個倖存者，也沒有一個逃脫。
JOSH|8|23|以色列 人生擒了 艾城 的王，把他解到 約書亞 那裏。
JOSH|8|24|以色列 人在田間和曠野殺盡了追趕他們的 艾城 所有的居民。他們全倒在刀下，直到滅盡。 以色列 眾人就回到 艾城 ，用刀殺了城中的人。
JOSH|8|25|當日殺死的人，連男帶女共有一萬二千，這也是 艾城 所有的人。
JOSH|8|26|約書亞 沒有收回手裏所伸出來的標槍，直到他滅絕 艾城 所有的居民。
JOSH|8|27|只是牲畜和城內所奪的財物， 以色列 人都照耶和華所吩咐 約書亞 的話，取為自己的掠物。
JOSH|8|28|約書亞 焚燒 艾城 ，使城成為永遠的廢墟，直到今日還是荒涼。
JOSH|8|29|他把 艾城 的王掛在樹上，直到晚上。日落的時候， 約書亞 吩咐人把屍首從樹上取下來，丟在城門口，並在屍首上堆了一大堆石頭，直存到今日。
JOSH|8|30|那時， 約書亞 在 以巴路山 上為耶和華－ 以色列 的上帝築一座壇。
JOSH|8|31|這壇是照耶和華的僕人 摩西 吩咐 以色列 人，用沒有動過鐵器的整塊石頭所築的，正如 摩西 律法書上所寫的。他們在這壇上給耶和華奉獻燔祭，又宰牲作為平安祭。
JOSH|8|32|約書亞 在那裏，當著 以色列 人面前，將 摩西 所寫的律法抄寫在石頭上。
JOSH|8|33|以色列 眾人，無論是本地人或寄居的，都和他們的長老、官長和審判官，站在約櫃兩旁，在抬耶和華約櫃的 利未 家的祭司面前，一半對著 基利心山 ，一半對著 以巴路山 ，照耶和華的僕人 摩西 先前所吩咐的，為 以色列 百姓祝福。
JOSH|8|34|隨後， 約書亞 將律法上祝福和詛咒的話，照著律法書上一切所寫的，宣讀一遍。
JOSH|8|35|摩西 所吩咐的一切話， 約書亞 在 以色列 全會眾和婦女、孩童，以及住在他們中間的外人面前，沒有一句不宣讀的。
JOSH|9|1|約旦河 西，住山區、低地和沿 大海 一帶直到 黎巴嫩 的諸王，就是 赫 人、 亞摩利 人、 迦南 人、 比利洗 人、 希未 人、 耶布斯 人的諸王，聽見這事，
JOSH|9|2|就都聚集，同心合意要與 約書亞 和 以色列 人作戰。
JOSH|9|3|基遍 的居民聽見 約書亞 向 耶利哥 和 艾城 所做的事，
JOSH|9|4|就設詭計，假扮使者 出去。他們拿舊布袋和破裂補過的舊皮酒袋馱在驢上，
JOSH|9|5|將補過的舊鞋穿在腳上，把舊衣服穿在身上，作食物的餅都又乾又長了霉 。
JOSH|9|6|他們到 吉甲 營中 約書亞 那裏，對他和 以色列 人說：「我們是從遠地來的，現在求你與我們立約。」
JOSH|9|7|以色列 人對 希未 人說：「或許你是住在我附近的。若是這樣，我怎能和你立約呢？」
JOSH|9|8|他們對 約書亞 說：「我們是你的僕人。」 約書亞 對他們說：「你們是甚麼人？是從哪裏來的？」
JOSH|9|9|他們對他說：「你的僕人是因耶和華－你上帝的名從極遠之地來的。我們聽見他的名聲，他在 埃及 所做的一切，
JOSH|9|10|以及他向 約旦河 東的兩個 亞摩利 王， 希實本 王 西宏 和在 亞斯她錄 的 巴珊 王 噩 所做的一切。
JOSH|9|11|我們的長老和我們當地所有的居民對我們說：『你們手裏要帶著路上用的乾糧去迎接 以色列 人，對他們說：我們是你們的僕人。現在求你們與我們立約。』
JOSH|9|12|我們出來要往你們這裏來的那日，這從我們家裏帶出來的餅是熱的；看哪，現在這餅又乾又長了霉。
JOSH|9|13|這些皮酒袋，我們盛酒的時候還是新的；看哪，現在已經破裂了。我們這些衣服和鞋，因為路途非常遙遠，也都穿舊了。」
JOSH|9|14|以色列 人收下他們的一些食物，但是沒有求問耶和華的指示。
JOSH|9|15|於是 約書亞 與他們建立和好關係，與他們立約，讓他們存活；會眾的領袖也向他們起誓。
JOSH|9|16|以色列 人與他們立約之後，過了三天才聽說他們是近鄰，住在附近。
JOSH|9|17|以色列 人起行，第三天就到了他們的城鎮，他們的城鎮是 基遍 、 基非拉 、 比錄 和 基列‧耶琳 。
JOSH|9|18|因為會眾的領袖已經指著耶和華－ 以色列 的上帝向他們起誓，所以 以色列 人不擊殺他們。全會眾就向領袖發怨言。
JOSH|9|19|眾領袖對全會眾說：「我們已經指著耶和華－ 以色列 的上帝向他們起誓，現在我們不能碰他們。
JOSH|9|20|我們要這樣對待他們，讓他們存活，免得因我們向他們所起的誓而憤怒臨到我們。」
JOSH|9|21|領袖對會眾說：「讓他們活著吧。」於是他們照領袖所說的，為全會眾作劈柴挑水的人。
JOSH|9|22|約書亞 召了他們來，對他們說：「你們為甚麼欺騙我們說：『我們離你們很遠』呢？其實你們就住在我們附近。
JOSH|9|23|現在你們當受詛咒！你們中間必不斷有人作奴僕，為我上帝的殿作劈柴挑水的人。」
JOSH|9|24|他們回答 約書亞 說：「因為確實有人告訴你的僕人，耶和華－你的上帝曾吩咐他的僕人 摩西 ，把這全地賜給你們，並要在你們面前除滅這地所有的居民。我們因你們的緣故很怕自己喪命，就做了這事。
JOSH|9|25|現在，看哪，我們在你手中，你看怎樣待我們是好的，是對的，就這樣做吧！」
JOSH|9|26|於是 約書亞 就這樣對待他們，他救了他們脫離 以色列 人的手， 以色列 人沒有殺他們。
JOSH|9|27|那日， 約書亞 分派他們到耶和華選擇的地方，為會眾和耶和華的壇劈柴挑水，直到今日。
JOSH|10|1|耶路撒冷 王 亞多尼‧洗德 聽見 約書亞 奪了 艾城 ，徹底毀滅，處置 艾城 和 艾城 的王像處置 耶利哥 和 耶利哥 的王一樣，又聽見 基遍 的居民與 以色列 人立了和約，住在他們中間，
JOSH|10|2|耶路撒冷 人就很懼怕，因為 基遍 是一座大城，如京城一樣，比 艾城 更大，並且城內的人都是勇士。
JOSH|10|3|耶路撒冷 王 亞多尼‧洗德 派人去見 希伯崙 王 何咸 、 耶末 王 毗蘭 、 拉吉 王 雅非亞 和 伊磯倫 王 底璧 ，說：
JOSH|10|4|「求你們上來幫助我，我們好攻打 基遍 ，因為它與 約書亞 和 以色列 人立了和約。」
JOSH|10|5|於是五個 亞摩利 王，就是 耶路撒冷 王、 希伯崙 王、 耶末 王、 拉吉 王和 伊磯倫 王，聯合上去，率領他們所有的軍隊，對著 基遍 安營，要攻打 基遍 。
JOSH|10|6|基遍 人就派人到 吉甲 的營中 約書亞 那裏，說：「不要袖手不顧你的僕人，求你趕快上來拯救我們，幫助我們，因為住山區 亞摩利 人的諸王已經聯合來攻擊我們。」
JOSH|10|7|於是 約書亞 和所有跟他一起作戰的士兵，以及大能的勇士，從 吉甲 上去。
JOSH|10|8|耶和華對 約書亞 說：「不要怕他們， 因為我已將他們交在你手裏，他們沒有一人能在你面前站立得住。」
JOSH|10|9|約書亞 就連夜從 吉甲 上去，猛然襲擊他們。
JOSH|10|10|耶和華使他們在 以色列 人面前潰亂。 約書亞 在 基遍 大大擊殺他們，在 伯‧和崙 的上坡路上追趕他們，擊殺他們，直到 亞西加 和 瑪基大 。
JOSH|10|11|他們在 以色列 人面前逃跑。正在 伯‧和崙 下坡的時候，耶和華從天上降下大冰雹 在他們身上，直降到 亞西加 ，打死他們。被冰雹打死的，比 以色列 人用刀殺死的還多。
JOSH|10|12|當耶和華將 亞摩利 人交給 以色列 人的那一日， 約書亞 向耶和華說話，在 以色列 人眼前說： 「太陽啊，停在 基遍 ； 月亮啊，停在 亞雅崙谷 。」
JOSH|10|13|太陽就停住，月亮就止住， 直到國民向敵人報仇。 這事豈不是寫在《雅煞珥書》上嗎？太陽停在天空當中，沒有急速下落，約有一整天。
JOSH|10|14|在這日以前，這日以後，耶和華聽人的聲音，沒有像這日的，這是因為耶和華為 以色列 作戰。
JOSH|10|15|約書亞 和跟他一起的 以色列 眾人回到 吉甲 的營中。
JOSH|10|16|那五個王逃跑，躲在 瑪基大 洞裏。
JOSH|10|17|有人告訴 約書亞 說：「那五個王已經找到了，都躲在 瑪基大 洞裏。」
JOSH|10|18|約書亞 說：「你們把幾塊大石頭滾到洞口，派人在那裏看守他們。
JOSH|10|19|你們卻不可停留，要追趕你們的仇敵，從後面攻擊他們，不讓他們進到自己的城鎮，因為耶和華－你們的上帝已經把他們交在你們手裏。」
JOSH|10|20|約書亞 和 以色列 人徹底擊敗他們，直到把他們滅盡，只剩下少許的人逃進堅固的城。
JOSH|10|21|眾百姓就安然回到 瑪基大 營中 ，到 約書亞 那裏。沒有人敢向 以色列 人饒舌。
JOSH|10|22|約書亞 說：「打開洞口，把那五個王從洞裏帶出來，到我這裏。」
JOSH|10|23|眾人就這樣做，把那五個王，就是 耶路撒冷 王、 希伯崙 王、 耶末 王、 拉吉 王和 伊磯倫 王，從洞裏帶出來，到 約書亞 那裏。
JOSH|10|24|他們帶出那五個王到 約書亞 那裏的時候， 約書亞 就召了 以色列 眾人來，對和他同去的軍官說：「你們近前來，把腳踏在這些王的頸項上。」他們就近前來，把腳踏在這些王的頸項上。
JOSH|10|25|約書亞 對他們說：「你們不要懼怕，也不要驚惶。當剛強壯膽，因為耶和華必這樣處置你們要攻打的所有仇敵。」
JOSH|10|26|隨後， 約書亞 把這五個王殺死，掛在五棵樹上。他們就被掛在樹上，直到晚上。
JOSH|10|27|日落的時候， 約書亞 吩咐人把屍首從樹上取下來，丟在他們躲過的洞裏，把幾塊大石頭放在洞口，直存到今日。
JOSH|10|28|當日， 約書亞 奪了 瑪基大 ，用刀擊殺城中的人和王，把城中所有人完全滅盡，沒有留下一個倖存者。他處置 瑪基大 王，像從前處置 耶利哥 王一樣。
JOSH|10|29|約書亞 和跟他一起的 以色列 眾人從 瑪基大 往 立拿 去，攻打 立拿 。
JOSH|10|30|耶和華將 立拿 和 立拿 的王也交在 以色列 人手裏。 約書亞 攻打這城，用刀擊殺了城中所有的人，沒有留下一個倖存者。他處置 立拿 王，像從前處置 耶利哥 王一樣。
JOSH|10|31|約書亞 和跟他一起的 以色列 眾人從 立拿 往 拉吉 去，對著 拉吉 安營，攻打這城。
JOSH|10|32|耶和華將 拉吉 交在 以色列 人的手裏。第二日 約書亞 就奪了 拉吉 ，用刀擊殺了城中所有的人，正如他向 立拿 一切所做的。
JOSH|10|33|那時 基色 王 何蘭 上來幫助 拉吉 ， 約書亞 就把他和他的百姓都擊殺了，沒有留下一個倖存者。
JOSH|10|34|約書亞 和跟他一起的 以色列 眾人從 拉吉 往 伊磯倫 去，對著 伊磯倫 安營，攻打這城。
JOSH|10|35|當日 約書亞 就奪了城，用刀擊殺了城中的人。那日， 約書亞 把城中所有的人完全滅盡，正如他向 拉吉 一切所做的。
JOSH|10|36|約書亞 和跟他一起的 以色列 眾人從 伊磯倫 上 希伯崙 去，攻打這城，
JOSH|10|37|奪了 希伯崙 ，用刀擊敗 希伯崙 、它的王和屬它的一切城鎮，以及城中所有的人；他沒有留下一個倖存者，正如他向 伊磯倫 所做的，把城中所有的人完全滅盡。
JOSH|10|38|約書亞 和跟他一起的 以色列 眾人回到 底璧 ，攻打這城，
JOSH|10|39|奪了 底璧 和屬它的一切城鎮，又擒獲它的王，用刀把城中所有的人完全滅盡，沒有留下一個倖存者。他處置 底璧 和它的王，像從前處置 希伯崙 ，處置 立拿 和它的王一樣。
JOSH|10|40|這樣， 約書亞 擊敗全地的人，就是山區、 尼革夫 、低地、山坡的人，和那裏的眾王，沒有留下一個倖存者。他把凡有氣息的完全滅盡，正如耶和華－ 以色列 的上帝所吩咐的。
JOSH|10|41|約書亞 從 加低斯‧巴尼亞 攻到 迦薩 ，又攻打 歌珊 全地，直到 基遍 。
JOSH|10|42|約書亞 一舉擊敗了這些王，奪了他們的地，因為耶和華－ 以色列 的上帝為 以色列 作戰。
JOSH|10|43|於是 約書亞 和跟他一起的 以色列 眾人回到 吉甲 的營中。
JOSH|11|1|夏瑣 王 耶賓 聽見了，就派人到 瑪頓 王 約巴 、 伸崙 王、 押煞 王，
JOSH|11|2|和北方山區、 基尼烈 南邊的 亞拉巴 、低地、西邊 多珥 山岡 的諸王，
JOSH|11|3|以及東方和西方的 迦南 人、山區的 亞摩利 人、 赫 人、 比利洗 人、 耶布斯 人，和 黑門山 下 米斯巴 地的 希未 人那裏。
JOSH|11|4|他們和他們的眾軍都出來，一大隊人馬，多如海邊的沙，並有極多的戰車戰馬。
JOSH|11|5|眾王組成聯軍，來到 米倫 水邊一同安營，要與 以色列 作戰。
JOSH|11|6|耶和華對 約書亞 說：「你不要怕他們。明日這時，我必把他們全部交給 以色列 人殺滅。你要砍斷他們馬的蹄筋，用火焚燒他們的戰車。」
JOSH|11|7|於是 約書亞 和所有跟他一起作戰的士兵，來到 米倫 水邊，突然攻擊他們。
JOSH|11|8|耶和華將他們交在 以色列 人手裏， 以色列 人就擊殺他們，追趕他們到 西頓 大城，到 米斯利弗‧瑪音 ，直到東邊 米斯巴 的山谷。 以色列 人擊殺他們，沒有留下一個倖存者。
JOSH|11|9|約書亞 照耶和華所吩咐他的去做，砍斷他們馬的蹄筋，用火焚燒他們的戰車。
JOSH|11|10|那時， 約書亞 轉回，奪了 夏瑣 ，用刀殺了 夏瑣 王。先前 夏瑣 在這些王國中是為首的。
JOSH|11|11|以色列 人用刀擊殺城中所有的人，把他們完全滅盡；凡有氣息的，沒有留下一個。 約書亞 又用火焚燒 夏瑣 。
JOSH|11|12|約書亞 奪了這些王的一切城鎮，擒獲了這些王，用刀殺了他們，把他們完全滅盡，正如耶和華的僕人 摩西 所吩咐的。
JOSH|11|13|至於造在山岡上的城鎮，除了 夏瑣 以外， 以色列 人都沒有焚燒。 約書亞 只焚燒了 夏瑣 。
JOSH|11|14|從那些城鎮所奪的財物和牲畜， 以色列 人都取為自己的掠物。至於所有的人，他們都用刀殺了，直到滅盡；凡有氣息的，沒有留下一個。
JOSH|11|15|耶和華怎樣吩咐他的僕人 摩西 ， 摩西 就這樣吩咐 約書亞 ， 約書亞 也照樣做了。凡耶和華所吩咐 摩西 的， 約書亞 沒有一件偏離不做的。
JOSH|11|16|約書亞 奪了那全地，就是山區、整個 尼革夫 、 歌珊 全地、低地、 亞拉巴 、 以色列 的山區和山下的低地，
JOSH|11|17|從上 西珥 的 哈拉山 ，直到 黑門山 下面 黎巴嫩 平原的 巴力‧迦得 。他擒獲了那裏的眾王，把他們殺死。
JOSH|11|18|約書亞 和這些王作戰了很長的一段日子。
JOSH|11|19|除了 希未 人 基遍 的居民之外，沒有一城與 以色列 人講和，都是 以色列 人作戰奪來的。
JOSH|11|20|因為耶和華的意思是要使他們的心剛硬，來與 以色列 人作戰，好使他們全被殺滅，不蒙憐憫，反被除滅，正如耶和華所吩咐 摩西 的。
JOSH|11|21|那時 約書亞 來到，剪除了住山區、 希伯崙 、 底璧 、 亞拿伯 、整個 猶大 山區和 以色列 山區的 亞衲 族人。 約書亞 把他們和他們的城鎮盡都毀滅。
JOSH|11|22|以色列 人的地中沒有留下一個 亞衲 族人，只有一些還留在 迦薩 、 迦特 和 亞實突 。
JOSH|11|23|這樣， 約書亞 照著耶和華所吩咐 摩西 的一切話奪了那全地，就按著 以色列 支派所得的份把地分給他們為業。於是國中太平，沒有戰爭了。
JOSH|12|1|這些是 以色列 人在 約旦河 東，向日出的方向，從 亞嫩谷 直到 黑門山 ，以及東邊 亞拉巴 的整個地區所擊殺的王和所得的地：
JOSH|12|2|有住 希實本 的 亞摩利 王 西宏 ，他統治的地從 亞嫩谷 邊的 亞羅珥 起，包括谷中之城和 基列 的一半，直到 亞捫 人邊界的 雅博河 ，
JOSH|12|3|以及從東邊的 亞拉巴 ，直到 基尼烈海 ，又向東通過 伯‧耶施末 的路，直到 亞拉巴 的海，就是 鹽海 ，再往南直到 毗斯迦山 斜坡的山腳。
JOSH|12|4|又有 巴珊 王 噩 ，他是 利乏音 人所剩下的，住在 亞斯她錄 和 以得來 。
JOSH|12|5|他統治的地是 黑門山 、 撒迦 、 巴珊 全地，直到 基述 人和 瑪迦 人的邊界，以及 基列 的一半，直到 希實本 王 西宏 的邊界。
JOSH|12|6|這兩個王是耶和華的僕人 摩西 和 以色列 人所擊殺的。耶和華的僕人 摩西 把他們的地賜給 呂便 人、 迦得 人和 瑪拿西 半支派的人為業。
JOSH|12|7|這些是 約書亞 和 以色列 人在 約旦河 西所擊殺的諸王，他們的地從 黎巴嫩 平原的 巴力‧迦得 ，直上到 西珥 的 哈拉山 。 約書亞 按著 以色列 支派所得的份把這地分給他們為業，
JOSH|12|8|就是 赫 人、 亞摩利 人、 迦南 人、 比利洗 人、 希未 人、 耶布斯 人的地，包括山區、低地、 亞拉巴 、山坡、曠野和 尼革夫 。
JOSH|12|9|這些王是： 耶利哥 王一人， 靠近 伯特利 的 艾城 王一人，
JOSH|12|10|耶路撒冷 王一人， 希伯崙 王一人，
JOSH|12|11|耶末 王一人， 拉吉 王一人，
JOSH|12|12|伊磯倫 王一人， 基色 王一人，
JOSH|12|13|底璧 王一人， 基德 王一人，
JOSH|12|14|何珥瑪 王一人， 亞拉得 王一人，
JOSH|12|15|立拿 王一人， 亞杜蘭 王一人，
JOSH|12|16|瑪基大 王一人， 伯特利 王一人，
JOSH|12|17|他普亞 王一人， 希弗 王一人，
JOSH|12|18|亞弗 王一人， 拉沙崙 王一人，
JOSH|12|19|瑪頓 王一人， 夏瑣 王一人，
JOSH|12|20|伸崙‧米崙 王一人 ， 押煞 王一人，
JOSH|12|21|他納 王一人， 米吉多 王一人，
JOSH|12|22|基低斯 王一人， 靠近 迦密 的 約念 王一人，
JOSH|12|23|多珥 山岡 的 多珥 王一人， 吉甲 的 戈印 王一人，
JOSH|12|24|得撒 王一人， 共三十一個王。
JOSH|13|1|約書亞 年紀老邁，耶和華對他說：「你年紀老邁了，還有極多剩下的未得之地。
JOSH|13|2|這是剩下的地： 非利士 人的全境和一切屬於 基述 人的，
JOSH|13|3|是從 埃及 東邊的 西曷河 往北，直到 以革倫 的邊界，算是屬 迦南 人的地，那裏有 非利士 人五個領袖統治 迦薩 人、 亞實突 人、 亞實基倫 人、 迦特 人、 以革倫 人；還有屬於 亞衛 人的，
JOSH|13|4|在南邊；還有 迦南 人的全地，以及 西頓 人的 米亞拉 到 亞弗 ，直到 亞摩利 人的邊界；
JOSH|13|5|還有 迦巴勒 人的地，以及向日出方向的 黎巴嫩 全地，從 黑門山 下的 巴力‧迦得 ，直到 哈馬口 ；
JOSH|13|6|從 黎巴嫩 直到 米斯利弗‧瑪音 ，一切山區的居民，就是所有的 西頓 人，我必在 以色列 人面前趕走他們。你只管照我所吩咐的，抽籤將這地分給 以色列 人為業。
JOSH|13|7|現在你要把這地分給九個支派和 瑪拿西 半個支派為業。
JOSH|13|8|呂便 、 迦得 二支派已經和 瑪拿西 另外半個支派得了產業，就是耶和華的僕人 摩西 在 約旦河 東所賜給他們的：
JOSH|13|9|從 亞嫩谷 邊的 亞羅珥 和谷中之城， 米底巴 的整個平原，直到 底本 ；
JOSH|13|10|還有在 希實本 作王的 亞摩利 王 西宏 的諸城，直到 亞捫 人的邊界；
JOSH|13|11|還有 基列 ， 基述 人和 瑪迦 人的邊界，整個 黑門山 、整個 巴珊 ，直到 撒迦 ；
JOSH|13|12|還有在 亞斯她錄 和 以得來 作王的 巴珊 王 噩 的整個國土， 噩 是 利乏音 人惟一存留的。 摩西 擊敗了這些人，把他們趕走。
JOSH|13|13|以色列 人卻沒有趕走 基述 人和 瑪迦 人； 基述 人和 瑪迦 人仍住在 以色列 中，直到今日。
JOSH|13|14|只是 利未 支派， 摩西 沒有分產業給他們。他們的產業是獻給耶和華－ 以色列 上帝的火祭，正如耶和華對他們說的。
JOSH|13|15|摩西 按著 呂便 支派的宗族分產業給他們。
JOSH|13|16|他們的地界是 亞嫩谷 邊的 亞羅珥 和谷中之城，靠近 米底巴 的整個平原；
JOSH|13|17|還有 希實本 和屬 希實本 平原的各城， 底本 、 巴末‧巴力 、 伯‧巴力‧勉 、
JOSH|13|18|雅雜 、 基底莫 、 米法押 、
JOSH|13|19|基列亭 、 西比瑪 、谷中山岡上的 細列‧沙轄 、
JOSH|13|20|伯‧毗珥 、 毗斯迦山 斜坡、 伯‧耶施末 ；
JOSH|13|21|還有平原的各城，和 亞摩利 王 西宏 的整個國土。這 西宏 曾在 希實本 作王， 摩西 把他和 米甸 的族長 以未 、 利金 、 蘇珥 、 戶珥 、 利巴 擊殺了；他們都是屬 西宏 的領袖，曾住在這地。
JOSH|13|22|以色列 人殺了這些人時，也用刀殺了 比珥 的兒子占卜的 巴蘭 。
JOSH|13|23|呂便 人的地界就是 約旦河 和靠近 約旦河 的地。以上是 呂便 人按著宗族所得為業的城鎮和所屬的村莊。
JOSH|13|24|摩西 按著 迦得 支派的宗族分產業給他們。
JOSH|13|25|他們的地界是 雅謝 和 基列 的各城，以及 亞捫 人之地的一半，直到 拉巴 前面的 亞羅珥 ；
JOSH|13|26|還有從 希實本 到 拉抹‧米斯巴 和 比多寧 ，又從 瑪哈念 到 底璧 的邊界，
JOSH|13|27|和谷中的 伯‧亞蘭 、 伯‧寧拉 、 疏割 、 撒分 ，就是 希實本 王 西宏 國土中其餘的地，以及 約旦河 與靠近 約旦河 的地，直到 基尼烈海 的邊緣，都在 約旦河 東。
JOSH|13|28|以上是 迦得 人按著宗族所得為業的城鎮和所屬的村莊。
JOSH|13|29|摩西 分產業給 瑪拿西 半支派，這是按著 瑪拿西 半支派的宗族分的。
JOSH|13|30|他們的地界是從 瑪哈念 起，包括整個 巴珊 全地，就是 巴珊 王 噩 的整個國土，以及在 巴珊 、 睚珥 的一切城鎮，共六十個；
JOSH|13|31|還有 基列 的一半，以及 巴珊 國的王 噩 的 亞斯她錄 和 以得來 兩座城。這些地是按著宗族分給 瑪拿西 兒子 瑪吉 子孫的，就是給 瑪吉 一半子孫的。
JOSH|13|32|以上是 摩西 在 約旦河 東， 耶利哥 對面的 摩押 平原所分配的產業。
JOSH|13|33|只是 利未 支派， 摩西 沒有把產業分給他們。耶和華－ 以色列 的上帝是他們的產業，正如耶和華對他們說的。
JOSH|14|1|這是 以色列 人在 迦南 地所得的產業，就是祭司 以利亞撒 和 嫩 的兒子 約書亞 ，以及 以色列 人各支派父系的領袖所分給他們的。
JOSH|14|2|他們照耶和華藉 摩西 所吩咐的，抽籤分產業給九個半支派。
JOSH|14|3|摩西 在 約旦河 東已經分了產業給另外兩個半支派。但是，他在他們中間沒有分產業給 利未 人。
JOSH|14|4|因 約瑟 的子孫成了兩個支派，就是 瑪拿西 和 以法蓮 。雖然他們沒有分地給 利未 人，卻給 利未 人城鎮居住，以及城鎮的郊外供他們牧養牲畜，安置財物。
JOSH|14|5|耶和華怎樣吩咐 摩西 ， 以色列 人就照樣做，把地分了。
JOSH|14|6|猶大 人來到 吉甲 ， 約書亞 那裏， 基尼洗 族 耶孚尼 的兒子 迦勒 對 約書亞 說：「耶和華在 加低斯‧巴尼亞 指著我和你對神人 摩西 所說的話，你都知道。
JOSH|14|7|耶和華的僕人 摩西 從 加低斯‧巴尼亞 差派我窺探這地的時候，我剛四十歲。我把心裏的話向他報告。
JOSH|14|8|雖然同我上去的眾弟兄使百姓膽戰心驚，我仍然專心跟從耶和華－我的上帝。
JOSH|14|9|那日， 摩西 起誓說：『你腳所踏之地必要歸你和你的子孫永遠為業，因為你專心跟從耶和華－我的上帝。』
JOSH|14|10|現在，看哪，耶和華照他所說的使我活了這四十五年。當 以色列 人在曠野飄流的時候，耶和華曾對 摩西 說了這話。現在，看哪，我已經八十五歲了。
JOSH|14|11|現今我還很健壯，像 摩西 差派我去的那天一樣；無論是戰爭，是出入，我現在的力量和那時的力量一樣。
JOSH|14|12|請你將耶和華那日所說的這山區給我。那日你也曾聽說，這裏有 亞衲 族人，以及寬大堅固的城，或許耶和華會照他所說的與我同在，我就把他們趕出去。」
JOSH|14|13|於是 約書亞 為 耶孚尼 的兒子 迦勒 祝福，把 希伯崙 給他為業。
JOSH|14|14|所以 希伯崙 成了 基尼洗 族 耶孚尼 的兒子 迦勒 的產業，直到今日，因為他專心跟從耶和華－ 以色列 的上帝。
JOSH|14|15|希伯崙 從前名叫 基列‧亞巴 ； 亞巴 是 亞衲 族最尊貴的人。於是國中太平，沒有戰爭了。
JOSH|15|1|猶大 支派按著宗族抽籤所得之地是在最南端，到 以東 的邊界，往南直到 尋 的曠野。
JOSH|15|2|他們南邊的地界是從 鹽海 的頂端，就是朝南的海灣開始，
JOSH|15|3|通到 亞克拉濱 斜坡的南邊，經過 尋 ，上到 加低斯‧巴尼亞 的南邊，又經過 希斯崙 ，上到 亞達珥 ，轉到 甲加 ，
JOSH|15|4|再經過 押們 ，順著 埃及 溪谷，這地界直通到海為止。這就是你們 南邊的地界。
JOSH|15|5|東邊的地界是從 鹽海 到 約旦河 口。北邊的地界是從 約旦河 口的海灣開始，
JOSH|15|6|這地界上到 伯‧曷拉 ，經過 伯‧亞拉巴 的北邊，這地界上到 呂便 之子 波罕 的磐石。
JOSH|15|7|這地界是從 亞割谷 往北上到 底璧 ，直向 亞都冥 斜坡對面的 吉甲 ，就是河的南邊，這地界再經過 隱‧示麥 泉，直通到 隱‧羅結 。
JOSH|15|8|這地界又上到 欣嫩子谷 ， 耶布斯 斜坡的南方， 耶布斯 就是 耶路撒冷 ，這地界又上到 欣嫩谷 西邊對面的山頂，就是在 利乏音谷 的最北端。
JOSH|15|9|這地界又從山頂延伸到 尼弗多亞 水泉，通到 以弗崙山 的城鎮，這地界又延伸到 巴拉 ， 巴拉 就是 基列‧耶琳 。
JOSH|15|10|這地界又從 巴拉 往西繞到 西珥山 ，經過 耶琳山 斜坡的北邊， 耶琳 就是 基撒崙 ，從那裏又下到 伯‧示麥 ，經過 亭拿 ，
JOSH|15|11|這地界通到 以革倫 斜坡的北邊。這地界又延伸到 施基崙 ，經過 巴拉山 到 雅比聶 ，這地界直通到海為止。
JOSH|15|12|西邊的地界就是 大海 和沿海一帶之地。這是 猶大 人按著宗族所得之地四圍的邊界。
JOSH|15|13|約書亞 照耶和華所指示的，把 猶大 人中的一份土地，就是 基列‧亞巴 ，分給 耶孚尼 的兒子 迦勒 。 亞巴 是 亞衲 族的祖先， 基列‧亞巴 就是 希伯崙 。
JOSH|15|14|迦勒 從那裏趕出 亞衲 的三族，就是 亞衲 族的 示篩 人、 亞希幔 人和 撻買 人。
JOSH|15|15|他又從那裏上去，攻擊 底璧 的居民，這 底璧 從前名叫 基列‧西弗 。
JOSH|15|16|迦勒 說：「誰能攻打 基列‧西弗 ，奪取那城，我就把我女兒 押撒 嫁給他。」
JOSH|15|17|迦勒 兄弟 基納斯 的兒子 俄陀聶 奪取了那城， 迦勒 就把女兒 押撒 嫁給他。
JOSH|15|18|押撒 來的時候，催促丈夫向她父親要一塊田。 押撒 一下驢， 迦勒 就對她說：「你要甚麼？」
JOSH|15|19|她說：「求你給我福分；你既然把我安置在 尼革夫 地，求你也給我水泉。」她父親就把上泉和下泉都賜給她。
JOSH|15|20|這是 猶大 支派按著宗族所得的產業。
JOSH|15|21|猶大 支派最南端，靠近 以東 邊界的城鎮，是 甲薛 、 以得 、 雅姑珥 、
JOSH|15|22|基拿 、 底摩拿 、 亞大達 、
JOSH|15|23|基低斯 、 夏瑣 、 以提楠 、
JOSH|15|24|西弗 、 提鍊 、 比亞綠 、
JOSH|15|25|夏瑣‧哈大他 、 加略‧希斯崙 ， 加略‧希斯崙 就是 夏瑣 ，
JOSH|15|26|亞曼 、 示瑪 、 摩拉大 、
JOSH|15|27|哈薩‧迦大 、 黑實門 、 伯‧帕列 、
JOSH|15|28|哈薩‧書亞 、 別是巴 、 比斯約他 、
JOSH|15|29|巴拉 、 以因 、 以森 、
JOSH|15|30|伊勒多臘 、 基失 、 何珥瑪 、
JOSH|15|31|洗革拉 、 麥瑪拿 、 三撒拿 、
JOSH|15|32|利巴勿 、 實忻 、 亞因 、 臨門 ，共二十九座城，還有所屬的村莊。
JOSH|15|33|在低地有 以實陶 、 瑣拉 、 亞實拿 、
JOSH|15|34|撒挪亞 、 隱‧干寧 、 他普亞 、 以楠 、
JOSH|15|35|耶末 、 亞杜蘭 、 梭哥 、 亞西加 、
JOSH|15|36|沙拉音 、 亞底他音 、 基底拉 、 基底羅他音 ，共十四座城，還有所屬的村莊。
JOSH|15|37|又有 洗楠 、 哈大沙 、 麥大‧迦得 、
JOSH|15|38|底連 、 米斯巴 、 約帖 、
JOSH|15|39|拉吉 、 波斯加 、 伊磯倫 、
JOSH|15|40|迦本 、 拉幔 、 基提利 、
JOSH|15|41|基低羅 、 伯‧大袞 、 拿瑪 、 瑪基大 ，共十六座城，還有所屬的村莊。
JOSH|15|42|又有 立拿 、 以帖 、 亞珊 、
JOSH|15|43|益弗他 、 亞實拿 、 尼悉 、
JOSH|15|44|基伊拉 、 亞革悉 、 瑪利沙 ，共九座城，還有所屬的村莊。
JOSH|15|45|又有 以革倫 和所屬的鄉鎮 與村莊，
JOSH|15|46|從 以革倫 直到海，一切靠近 亞實突 之地，以及所屬的村莊、
JOSH|15|47|亞實突 和所屬的鄉鎮與村莊， 迦薩 和所屬的鄉鎮與村莊，到 埃及 溪谷，直到 大海 以及沿海一帶之地。
JOSH|15|48|在山區有 沙密 、 雅提珥 、 梭哥 、
JOSH|15|49|大拿 、 基列‧薩拿 ， 基列‧薩拿 就是 底璧 ，
JOSH|15|50|亞拿伯 、 以實提莫 、 亞念 、
JOSH|15|51|歌珊 、 何崙 、 基羅 ，共十一座城，還有所屬的村莊。
JOSH|15|52|又有 亞拉 、 度瑪 、 以珊 、
JOSH|15|53|雅農 、 伯‧他普亞 、 亞非加 、
JOSH|15|54|宏他 、 基列‧亞巴 ， 基列‧亞巴 就是 希伯崙 ， 洗珥 ，共九座城，還有所屬的村莊。
JOSH|15|55|又有 瑪雲 、 迦密 、 西弗 、 淤他 、
JOSH|15|56|耶斯列 、 約甸 、 撒挪亞 、
JOSH|15|57|該隱 、 基比亞 、 亭拿 ，共十座城，還有所屬的村莊。
JOSH|15|58|又有 哈忽 、 伯‧夙 、 基突 、
JOSH|15|59|瑪臘 、 伯‧亞諾 、 伊勒提君 ，共六座城，還有所屬的村莊。
JOSH|15|60|又有 基列‧巴力 ， 基列‧巴力 就是 基列‧耶琳 ， 拉巴 ，共兩座城，還有所屬的村莊。
JOSH|15|61|在曠野有 伯‧亞拉巴 、 密丁 、 西迦迦 、
JOSH|15|62|匿珊 、 鹽城 、 隱‧基底 ，共六座城，還有所屬的村莊。
JOSH|15|63|至於住 耶路撒冷 的 耶布斯 人， 猶大 人不能把他們趕出去。於是， 耶布斯 人與 猶大 人同住在 耶路撒冷 ，直到今日。
JOSH|16|1|約瑟 的子孫抽籤所得之地是從靠近 耶利哥 的 約旦河 起，以 耶利哥 東邊的河水為邊界，經過曠野，從 耶利哥 上去，直到 伯特利 的山區；
JOSH|16|2|從 伯特利 又到 路斯 ，經過 亞基 人的邊界，直到 亞大錄 ；
JOSH|16|3|又往西，下到 押利提 人的邊界，到 下伯‧和崙 的邊界，到 基色 ，直通到海為止。
JOSH|16|4|約瑟 的兒子 瑪拿西 、 以法蓮 得了地業。
JOSH|16|5|以法蓮 子孫的地界，按著宗族所得的如下：他們地業的東界，是從 亞大錄‧亞達 到 上伯‧和崙 ，
JOSH|16|6|這地界直通到海。在北邊，這地界是從 密米他 ，向東繞到 他納‧示羅 ，又經過 雅挪哈 的東邊，
JOSH|16|7|從 雅挪哈 下到 亞大錄 和 拿拉 ，再到 耶利哥 ，直到 約旦河 為止。
JOSH|16|8|這地界又從 他普亞 ，順著 加拿河 往西延伸，直通到海為止。這就是 以法蓮 支派按著宗族所得的地業。
JOSH|16|9|在 瑪拿西 人地業的一切城鎮和所屬的村莊中，也保留一些城鎮給 以法蓮 的子孫。
JOSH|16|10|他們卻沒有趕出住在 基色 的 迦南 人。 迦南 人就住在 以法蓮 人中，成為服勞役的僕人，直到今日。
JOSH|17|1|瑪拿西 是 約瑟 的長子，這是他的支派抽籤所得之地。 瑪拿西 的長子， 基列 的父親 瑪吉 ，因為是勇士，就得了 基列 和 巴珊 。
JOSH|17|2|瑪拿西 其餘的子孫，就是 亞比以謝 的子孫， 希勒 的子孫， 亞斯烈 的子孫， 示劍 的子孫， 希弗 的子孫， 示米大 的子孫，都按著宗族抽籤得了地。這都是 約瑟 的兒子 瑪拿西 子孫中各宗族的男丁。
JOSH|17|3|瑪拿西 的玄孫， 瑪吉 的曾孫， 基列 的孫子， 希弗 的兒子 西羅非哈 沒有兒子，只有女兒。他的女兒名叫 瑪拉 、 挪阿 、 曷拉 、 密迦 、 得撒 。
JOSH|17|4|她們來到 以利亞撒 祭司和 嫩 的兒子 約書亞 以及眾領袖面前，說：「耶和華曾吩咐 摩西 在我們兄弟中分產業給我們。」於是 約書亞 照耶和華的指示，在她們叔伯中，把產業分給她們。
JOSH|17|5|除了 約旦河 東的 基列 和 巴珊 地之外，還有十份的地業是屬於 瑪拿西 的，
JOSH|17|6|因為 瑪拿西 支派的女子也在男子中分得產業。 基列 地屬於 瑪拿西 其餘的子孫。
JOSH|17|7|瑪拿西 的地界是從 亞設 起，到 示劍 前面的 密米他 ，往右 到 隱‧他普亞 居民之地。
JOSH|17|8|他普亞 地歸於 瑪拿西 ，只是 瑪拿西 邊界的 他普亞城 卻歸於 以法蓮 子孫。
JOSH|17|9|這地界從那裏下到 加拿河 。河南邊的城鎮雖然在 瑪拿西 境內，卻是屬於 以法蓮 的。 瑪拿西 的地界是在河的北邊直通到海為止。
JOSH|17|10|南邊屬於 以法蓮 ，北邊屬於 瑪拿西 ，以海為界；北邊達到 亞設 ，東邊達到 以薩迦 。
JOSH|17|11|瑪拿西 在 以薩迦 和 亞設 境內，有 伯‧善 和所屬的鄉鎮， 以伯蓮 和所屬的鄉鎮， 多珥 和所屬鄉鎮的居民；還有 隱‧多珥 和所屬鄉鎮的居民， 他納 和所屬鄉鎮的居民， 米吉多 和所屬鄉鎮的居民，共三個山岡 。
JOSH|17|12|只是 瑪拿西 的子孫不能趕出這些城鎮的居民， 迦南 人仍堅持住在那地。
JOSH|17|13|以色列 人強盛的時候，就叫 迦南 人做苦工，沒有把他們全然趕走。
JOSH|17|14|約瑟 的子孫對 約書亞 說：「耶和華到如今這樣賜福給我，我百姓眾多，你為甚麼只給我抽一籤，分一份的土地為業呢？」
JOSH|17|15|約書亞 對他們說：「如果你百姓眾多，而 以法蓮 山區太窄小，那麼你可以上 比利洗 人和 利乏音 人之地的樹林中，在那裏開墾。」
JOSH|17|16|約瑟 的子孫說：「那山區容不下我們，而且住平原的 迦南 人，就是住 伯‧善 和所屬的鄉鎮，以及住在 耶斯列 平原的人，都有鐵的戰車。」
JOSH|17|17|約書亞 對 約瑟 家，就是 以法蓮 和 瑪拿西 人，說：「你百姓眾多，並且強大，不可只有一籤而已。
JOSH|17|18|那山區也要歸你，雖然是樹林，你可以去開墾，邊緣之地也必歸你。 迦南 人縱然強盛，有鐵的戰車，你也能把他們趕出去。」
JOSH|18|1|以色列 全會眾都聚集在 示羅 ，把會幕設立在那裏。那地已經被他們征服了。
JOSH|18|2|以色列 人中剩下七個支派還沒有分得他們的地業。
JOSH|18|3|約書亞 對 以色列 人說：「耶和華－你們列祖的上帝所賜給你們的地，你們耽延不去得，要到幾時呢？
JOSH|18|4|你們每支派要選三個人，我好派他們去，他們要起身走遍那地，按照各支派應得的地業寫明，然後回到我這裏來。
JOSH|18|5|他們要把地分成七份。 猶大 在南方，住在他的境內。 約瑟 家在北方，住在他們的境內。
JOSH|18|6|你們把地劃成七份之後，就要把所寫的帶到我這裏來。我要在耶和華－我們的上帝面前，為你們抽籤。
JOSH|18|7|利未 人在你們中間沒有分得地業，因為耶和華祭司的職分就是他們的產業。 迦得 支派、 呂便 支派和 瑪拿西 半支派已經在 約旦河 東得了地業，是耶和華的僕人 摩西 給他們的。」
JOSH|18|8|那些去劃地的人起來正要去的時候， 約書亞 吩咐他們說：「你們去走遍那地，把地劃分以後，就回到我這裏來。我要在 示羅 這裏，在耶和華面前為你們抽籤。」
JOSH|18|9|那些人就去了，走遍那地，按照城鎮把地劃成七份，寫在冊上，回到 示羅 營中 約書亞 那裏。
JOSH|18|10|約書亞 就在 示羅 ，在耶和華面前為他們抽籤。 約書亞 按照 以色列 人的支派，在那裏把地分給他們。
JOSH|18|11|便雅憫 支派，按著宗族抽籤所得之地，是在 猶大 子孫和 約瑟 子孫之間。
JOSH|18|12|他們北邊的地界是從 約旦河 起，上到 耶利哥 斜坡的北邊，再往西上到山區，直到 伯‧亞文 的曠野。
JOSH|18|13|這地界從那裏往南經過 路斯 ，直到 路斯 的斜坡， 路斯 就是 伯特利 ，又下到 亞他錄‧亞達 ，直到 下伯‧和崙 南邊的山。
JOSH|18|14|這地界往西延伸，又轉向南，從 伯‧和崙 南邊對面的山，直通到 猶大 人的城 基列‧巴力 ， 基列‧巴力 就是 基列‧耶琳 。這就是西邊的地界。
JOSH|18|15|南邊是從 基列‧耶琳 的頂端為起點，這地界往西 通到 尼弗多亞 水泉，
JOSH|18|16|這地界又下到 欣嫩子谷 對面山的邊緣，就是 利乏音谷 的北邊；又下到 欣嫩谷 ，沿著 耶布斯 斜坡的南邊，下到 隱‧羅結 ；
JOSH|18|17|又往北轉彎，通到 隱‧示麥 ，直到 亞都冥 斜坡對面的 基利綠 ，又下到 呂便 之子 波罕 的磐石，
JOSH|18|18|又往北經過 亞拉巴 對面的斜坡 ，下到 亞拉巴 。
JOSH|18|19|這地界又經過 伯‧曷拉 斜坡的北邊，直通到 鹽海 的北灣，就是 約旦河 的南端為止。這就是南邊的地界。
JOSH|18|20|東邊的地界是 約旦河 。這是 便雅憫 人按著宗族，照著他們四圍的邊界所得的地業。
JOSH|18|21|便雅憫 支派按著宗族所得的城鎮就是： 耶利哥 、 伯‧曷拉 、 伊麥‧基悉 、
JOSH|18|22|伯‧亞拉巴 、 洗瑪臉 、 伯特利 、
JOSH|18|23|亞文 、 巴拉 、 俄弗拉 、
JOSH|18|24|基法‧阿摩尼 、 俄弗尼 和 迦巴 ，共十二座城，以及所屬的村莊；
JOSH|18|25|又有 基遍 、 拉瑪 、 比錄 、
JOSH|18|26|米斯巴 、 基非拉 、 摩撒 、
JOSH|18|27|利堅 、 伊利毗勒 、 他拉拉 、
JOSH|18|28|洗拉 、 以利弗 、 耶布斯 ， 耶布斯 就是 耶路撒冷 ， 基比亞 、 基列 ，共十四座城，以及所屬的村莊。這是 便雅憫 人按著宗族所得的地業。
JOSH|19|1|第二籤是 西緬 ，是 西緬 支派的人按著宗族抽出的，他們所得的地業是在 猶大 人地業的中間。
JOSH|19|2|他們所得為業之地是： 別是巴 ，或名 示巴 ， 摩拉大 、
JOSH|19|3|哈薩‧書亞 、 巴拉 、 以森 、
JOSH|19|4|伊勒多臘 、 比土力 、 何珥瑪 、
JOSH|19|5|洗革拉 、 伯‧瑪加博 、 哈薩‧蘇撒 、
JOSH|19|6|伯‧利巴勿 、 沙魯險 ，共十三座城，還有所屬的村莊；
JOSH|19|7|又有 亞因 、 利門 、 以帖 、 亞珊 ，共四座城，還有所屬的村莊；
JOSH|19|8|以及這些城鎮周圍一切的村莊，直到 巴拉‧比珥 ，就是 尼革夫 的 拉瑪 。這是 西緬 支派的人按著宗族所得的地業。
JOSH|19|9|西緬 人的地業取自 猶大 人的土地，因為 猶大 人所得的份過多，所以 西緬 人從 猶大 人的地業中取了地業。
JOSH|19|10|第三籤是 西布倫 人按著宗族抽到的。他們地業的邊界延伸到 撒立 。
JOSH|19|11|他們的地界往西，上到 瑪拉拉 ，達到 大巴設 ，又達到 約念 前面的河。
JOSH|19|12|又從 撒立 往東轉到向日出的方向，經過 吉斯綠‧他泊 的邊界，到 大比拉 ，又上到 雅非亞 。
JOSH|19|13|又從那裏往東，經過 迦特‧希弗 ，到 以特‧加汛 ，通到 臨門 ，延伸到 尼亞 。
JOSH|19|14|這地界在北邊繞過 尼亞 ，到 哈拿頓 ，直通到 伊弗他‧伊勒谷 ，
JOSH|19|15|包括 加他 、 拿哈拉 、 伸崙 、 以大拉 、 伯利恆 ，共十二座城，還有所屬的村莊。
JOSH|19|16|這些城鎮和所屬的村莊是 西布倫 人按著宗族所得的地業。
JOSH|19|17|第四籤是 以薩迦 ，是 以薩迦 人按著宗族抽出的。
JOSH|19|18|他們的地界是到 耶斯列 、 基蘇律 、 書念 、
JOSH|19|19|哈弗連 、 示按 、 亞拿哈拉 、
JOSH|19|20|拉璧 、 基善 、 亞別 、
JOSH|19|21|利篾 、 隱‧干寧 、 隱‧哈大 、 伯‧帕薛 。
JOSH|19|22|這地界達到 他泊 、 沙哈洗瑪 、 伯‧示麥 ，他們的地界直通到 約旦河 為止，共十六座城，還有所屬的村莊。
JOSH|19|23|這些城鎮和所屬的村莊是 以薩迦 支派的人按著宗族所得的地業。
JOSH|19|24|第五籤是 亞設 支派的人按著宗族抽出的。
JOSH|19|25|他們的地界是 黑甲 、 哈利 、 比田 、 押煞 、
JOSH|19|26|亞拉米勒 、 亞末 、 米沙勒 ，往西達到 迦密 ，又到 希曷‧立納 ，
JOSH|19|27|又轉到向日出方向的 伯‧大袞 ，達到 細步綸 ；又往北到 伊弗他‧伊勒谷 ，到 伯‧以墨 和 尼業 ，也通到 迦步勒 的左邊 ，
JOSH|19|28|又到 義伯崙 、 利合 、 哈們 、 加拿 ，直到 西頓 大城。
JOSH|19|29|這地界轉到 拉瑪 ，直到堅固的 推羅城 。這地界又轉到 何薩 ，靠近 亞革悉 一帶的地方 ，直通到海為止。
JOSH|19|30|又有 烏瑪 、 亞弗 、 利合 ，共二十二座城，還有所屬的村莊。
JOSH|19|31|這些城鎮和所屬的村莊是 亞設 支派的人按著宗族所得的地業。
JOSH|19|32|第六籤是 拿弗他利 人，是 拿弗他利 人按著宗族抽出的。
JOSH|19|33|他們的地界是從 希利弗 ，從 撒拿音 的橡樹、 亞大米‧尼吉 和 雅比聶 ，直到 拉共 ，直通到 約旦河 為止。
JOSH|19|34|這地界往西轉到 亞斯納‧他泊 ，從那裏通到 戶割 ，南邊達到 西布倫 ，西邊達到 亞設 ，向日出的方向達到 約旦河 的 猶大 。
JOSH|19|35|堅固的城有 西丁 、 側耳 、 哈末 、 拉甲 、 基尼烈 、
JOSH|19|36|亞大瑪 、 拉瑪 、 夏瑣 、
JOSH|19|37|基低斯 、 以得來 、 隱‧夏瑣 、
JOSH|19|38|以利穩 、 密大‧伊勒 、 和璉 、 伯‧亞納 、 伯‧示麥 ，共十九座城，還有所屬的村莊。
JOSH|19|39|這些城鎮和所屬的村莊是 拿弗他利 支派的人按著宗族所得的地業。
JOSH|19|40|但 支派，按著宗族，抽到第七籤。
JOSH|19|41|他們地業的邊界是 瑣拉 、 以實陶 、 伊珥‧示麥 、
JOSH|19|42|沙拉賓 、 亞雅崙 、 伊提拉 、
JOSH|19|43|以倫 、 亭拿 、 以革倫 、
JOSH|19|44|伊利提基 、 基比頓 、 巴拉 、
JOSH|19|45|伊胡得 、 比尼‧比拉 、 迦特‧臨門 、
JOSH|19|46|美‧耶昆 、 拉昆 ，以及 約帕 對面的地界。
JOSH|19|47|當 但 的子孫失去他們疆土的時候，就上去攻取 利善 ，用刀擊殺城中的人，得了那城，住在城中，以他們祖先 但 的名字將 利善 改名為 但 。
JOSH|19|48|這些城鎮和所屬的村莊是 但 支派的人按著宗族所得的地業。
JOSH|19|49|以色列 人按著疆土完成了地業的分配，就在他們中間把地給 嫩 的兒子 約書亞 為業。
JOSH|19|50|他們照著耶和華的指示，把 約書亞 所要的城，就是 以法蓮 山區的 亭拿‧西拉 給了他。 約書亞 修建那城，住在城中。
JOSH|19|51|這就是 以利亞撒 祭司和 嫩 的兒子 約書亞 ，以及 以色列 人各支派父系的領袖，在 示羅 會幕的門口，耶和華面前抽籤所分的地業。這樣， 他們就完成了分地的事。
JOSH|20|1|耶和華吩咐 約書亞 說：
JOSH|20|2|「你吩咐 以色列 人說：『你們要照我藉 摩西 所吩咐你們的，為自己設立逃城，
JOSH|20|3|使那無意中誤殺人的，可以逃到那裏。這些要作為你們逃避報血仇者的城。
JOSH|20|4|殺人者要逃到這些城中的一座，站在城門口，把他的事情陳訴給那城的長老聽。他們就要接他入城，給他地方，讓他住在他們中間。
JOSH|20|5|若是報血仇者追上了他，長老不可把他交在報血仇者的手裏，因為他是無意中殺了鄰舍的，並非過去彼此之間有仇恨。
JOSH|20|6|他要住在那城裏，直到他站在會眾面前受審判；等到當時的大祭司死後，殺人者才可以回到本城本家，就是他所逃出來的那城。』」
JOSH|20|7|於是， 以色列 人劃分 拿弗他利 山區 加利利 的 基低斯 、 以法蓮 山區的 示劍 和 猶大 山區的 基列‧亞巴 ， 基列‧亞巴 就是 希伯崙 。
JOSH|20|8|他們在 約旦河 的另一邊，就是 耶利哥 的東邊，從 呂便 支派中，在曠野的平原設立 比悉 ，從 迦得 支派中設立 基列 的 拉末 ，從 瑪拿西 支派中設立 巴珊 的 哥蘭 。
JOSH|20|9|這都是為 以色列 眾人和在他們中間寄居的外人所指定的城鎮，使凡誤殺人者可以逃到那裏，不至於死在報血仇者的手中，直到他站在會眾面前受審判 。
JOSH|21|1|利未 人的眾族長近前來到 以利亞撒 祭司和 嫩 的兒子 約書亞 ，以及 以色列 人各支派父系的領袖那裏，
JOSH|21|2|在 迦南 地的 示羅 對他們說：「從前耶和華曾藉著 摩西 吩咐給我們城鎮居住，以及城鎮的郊外供我們牧養牲畜。」
JOSH|21|3|於是 以色列 人照耶和華的指示，從自己的地業中，把這些城鎮和城鎮的郊外給了 利未 人。
JOSH|21|4|哥轄 族抽了籤。 利未 人中 亞倫 祭司的子孫，從 猶大 支派、 西緬 支派、 便雅憫 支派的地業中，抽籤得了十三座城。
JOSH|21|5|哥轄 其餘的子孫，從 以法蓮 支派、 但 支派、 瑪拿西 半支派宗族的地業中，抽籤得了十座城。
JOSH|21|6|革順 的子孫，從 以薩迦 支派、 亞設 支派、 拿弗他利 支派、住 巴珊 的 瑪拿西 半支派宗族的地業中，抽籤得了十三座城。
JOSH|21|7|米拉利 的子孫，按著宗族，從 呂便 支派、 迦得 支派、 西布倫 支派的地業中，得了十二座城。
JOSH|21|8|以色列 人照耶和華藉 摩西 所吩咐的，把這些城鎮和城鎮的郊外，抽籤給 利未 人。
JOSH|21|9|他們從 猶大 支派和 西緬 支派的地業中，給了以下所記名字的各城，
JOSH|21|10|就是給 利未 人 哥轄 宗族的 亞倫 子孫，因為他們抽到第一籤：
JOSH|21|11|把 猶大 山區的 基列‧亞巴 ，就是 希伯崙 ，和四圍的郊野給了他們。 亞巴 是 亞衲 族的祖先。
JOSH|21|12|但是，這城的田地和所屬的村莊卻給了 耶孚尼 的兒子 迦勒 為業。
JOSH|21|13|他們把 希伯崙 ，就是誤殺人的逃城和城的郊外，給了 亞倫 祭司的子孫；又給了 立拿 和城的郊外、
JOSH|21|14|雅提珥 和城的郊外、 以實提莫 和城的郊外、
JOSH|21|15|何崙 和城的郊外、 底璧 和城的郊外、
JOSH|21|16|亞因 和城的郊外、 淤他 和城的郊外，以及 伯‧示麥 和城的郊外，共九座城，都是從這二支派中分出來的。
JOSH|21|17|又從 便雅憫 支派的地業中給了 基遍 和城的郊外、 迦巴 和城的郊外、
JOSH|21|18|亞拿突 和城的郊外，以及 亞勒們 和城的郊外，共四座城。
JOSH|21|19|亞倫 子孫作祭司的共有十三座城，以及城的郊外。
JOSH|21|20|利未 人 哥轄 的宗族，就是 哥轄 其餘的子孫，抽籤所得的城是從 以法蓮 支派來的。
JOSH|21|21|他們把 以法蓮 山區的 示劍 ，就是誤殺人的逃城和城的郊外給了 哥轄 其餘的子孫；又給了 基色 和城的郊外、
JOSH|21|22|基伯先 和城的郊外，以及 伯‧和崙 和城的郊外，共四座城。
JOSH|21|23|又從 但 支派的地業中給了 伊利提基 和城的郊外、 基比頓 和城的郊外、
JOSH|21|24|亞雅崙 和城的郊外，以及 迦特‧臨門 和城的郊外，共四座城。
JOSH|21|25|又從 瑪拿西 半支派的地業中給了 他納 和城的郊外，以及 迦特‧臨門 和城的郊外，共兩座城。
JOSH|21|26|哥轄 其餘的子孫共有十座城，以及城的郊外。
JOSH|21|27|利未 人宗族中 革順 的子孫，從 瑪拿西 半支派的地業中所得的是 巴珊 的 哥蘭 ，就是誤殺人的逃城和城的郊外，以及 比‧施提拉 和城的郊外，共兩座城。
JOSH|21|28|從 以薩迦 支派的地業中所得的是 基善 和城的郊外、 大比拉 和城的郊外、
JOSH|21|29|耶末 和城的郊外，以及 隱‧干寧 和城的郊外，共四座城。
JOSH|21|30|從 亞設 支派的地業中所得的是 米沙勒 和城的郊外、 押頓 和城的郊外、
JOSH|21|31|黑甲 和城的郊外，以及 利合 和城的郊外，共四座城。
JOSH|21|32|從 拿弗他利 支派的地業中所得的是 加利利 的 基低斯 ，就是誤殺人的逃城和城的郊外、 哈末‧多珥 和城的郊外，以及 加珥坦 和城的郊外，共三座城。
JOSH|21|33|革順 人按著宗族共有十三個城，以及城的郊外。
JOSH|21|34|其餘的 利未 人，就是 米拉利 的子孫，按著宗族從 西布倫 支派的地業中所得的是 約念 和城的郊外、 加珥他 和城的郊外、
JOSH|21|35|丁拿 和城的郊外，以及 拿哈拉 和城的郊外，共四座城。
JOSH|21|36|從 呂便 支派的地業中所得的是 比悉 和城的郊外、 雅雜 和城的郊外、
JOSH|21|37|基底莫 和城的郊外，以及 米法押 和城的郊外，共四座城。
JOSH|21|38|從 迦得 支派的地業中所得的是 基列 的 拉末 ，就是誤殺人的逃城和城的郊外、 瑪哈念 和城的郊外、
JOSH|21|39|希實本 和城的郊外，以及 雅謝 和城的郊外，共四座城。
JOSH|21|40|利未 宗族其餘的人，就是 米拉利 的子孫，按著宗族抽籤所得的，共十二座城。
JOSH|21|41|利未 人在 以色列 人的地業中所得的城，共四十八個，還有城的郊外。
JOSH|21|42|這些城的四圍都有郊野，每個城都是如此。
JOSH|21|43|這樣，耶和華將從前向他們列祖起誓要給他們的全地賜給 以色列 人，他們就得了為業，住在其中。
JOSH|21|44|耶和華照著向他們列祖起誓所應許的一切，賜給他們全境安寧。他們所有的仇敵，沒有一個能在他們面前站立得住。耶和華把所有仇敵都交在他們手中。
JOSH|21|45|耶和華應許賜福給 以色列 家的話，一句都沒有落空，全都應驗了。
JOSH|22|1|此後， 約書亞 召了 呂便 人、 迦得 人和 瑪拿西 半支派的人來，
JOSH|22|2|對他們說：「耶和華的僕人 摩西 所吩咐你們的，你們都遵守了；我吩咐你們的話，你們也都聽從了。
JOSH|22|3|你們這許多日子，都沒有撇棄你們的弟兄，直到今日，並且遵守了耶和華你們上帝所吩咐的命令。
JOSH|22|4|如今耶和華－你們的上帝已經照著他所應許的，使你們的弟兄得享安寧。你們現在可以返回自己的帳棚，回到耶和華的僕人 摩西 在 約旦河 東所賜給你們為業之地。
JOSH|22|5|只是務要謹守遵行耶和華的僕人 摩西 所吩咐你們的誡命和律法，愛耶和華－你們的上帝，行他一切的道，守他的誡命，緊緊跟隨他，盡心盡性事奉他。」
JOSH|22|6|於是 約書亞 為他們祝福，送他們回去，他們就回到自己的帳棚去了。
JOSH|22|7|摩西 在 巴珊 曾把地業分給 瑪拿西 的半支派；然後 約書亞 在 約旦河 的西岸，在他們弟兄中，又把地業分給 瑪拿西 的另外半支派。 約書亞 送他們回帳棚的時候，為他們祝福，
JOSH|22|8|對他們說：「你們要把許多財物，許多牲畜，和金、銀、銅、鐵，以及許多衣服，帶回你們的帳棚去，要把你們從仇敵奪來的東西分給你們的眾弟兄。」
JOSH|22|9|於是 呂便 人、 迦得 人、 瑪拿西 半支派的人從 迦南 地的 示羅 起行，離開 以色列 人，回到他們已得為業的 基列 地，就是他們照耶和華藉 摩西 所吩咐而得的。
JOSH|22|10|呂便 人、 迦得 人和 瑪拿西 半支派的人到了 迦南 地的 約旦河 一帶地方，就在 約旦河 那裏築了一座壇，一座高大壯觀的壇。
JOSH|22|11|以色列 人聽見了，說：「看哪， 呂便 人、 迦得 人、 瑪拿西 半支派的人在 迦南 地對面， 約旦河 一帶地方， 以色列 人的境內，築了一座壇。」
JOSH|22|12|以色列 人一聽見，全會眾的 以色列 人就聚集在 示羅 ，要上去攻打他們。
JOSH|22|13|以色列 人派 以利亞撒 祭司的兒子 非尼哈 ，往 基列 地，到 呂便 人、 迦得 人和 瑪拿西 半支派的人那裏。
JOSH|22|14|和他同去的還有十個領袖， 以色列 每個支派在父家中各派一個領袖，這些人每一個在 以色列 族系中都是父家的領袖。
JOSH|22|15|他們來到 基列 地，到 呂便 人、 迦得 人和 瑪拿西 半支派的人那裏，對他們說：
JOSH|22|16|「耶和華全會眾這樣說：『你們今日離棄耶和華不跟從他，干犯 以色列 的上帝，悖逆耶和華，為自己築了一座壇，你們所犯的是何等的罪！
JOSH|22|17|從前我們在 毗珥 犯的罪孽，導致瘟疫臨到耶和華的會眾，甚至到今日都還沒有洗淨，這還算小事嗎？
JOSH|22|18|你們今日竟然離棄耶和華不跟從他！你們今日既然悖逆耶和華，明日他必向 以色列 全會眾發怒。
JOSH|22|19|若你們認為所得為業之地不潔淨，可以過來，到耶和華之地，就是耶和華的帳幕所居住之地，在我們中間得地業。你們卻不可悖逆耶和華，也不可背叛我們，在耶和華－我們上帝的壇以外為自己築壇。
JOSH|22|20|從前 謝拉 的曾孫 亞干 豈不是在那當滅的物上犯了罪，導致憤怒臨到 以色列 全會眾嗎？死在他所犯的罪中的，不只是他一個人而已！』」
JOSH|22|21|於是 呂便 人、 迦得 人、 瑪拿西 半支派的人回答 以色列 族系的領袖，說：
JOSH|22|22|「大能者上帝耶和華！大能者上帝耶和華！他已知道，願 以色列 人也知道，我們若有悖逆的行為，或是干犯耶和華，你今日就不要讓我們活著！
JOSH|22|23|若我們為自己築壇，離棄耶和華不跟從他，或將燔祭、素祭、平安祭獻在壇上，願耶和華親自追究。
JOSH|22|24|不是這樣！我們做這事的原因是懼怕將來你們的子孫對我們的子孫說：『你們與耶和華－ 以色列 的上帝有甚麼關係呢？
JOSH|22|25|因為耶和華以 約旦河 作我們和你們 呂便 人、 迦得 人的交界，所以你們在耶和華裏無份。』這樣，你們的子孫就使我們的子孫不再敬畏耶和華了。
JOSH|22|26|因此我們說：『不如為自己築一座壇，不是為獻燔祭，也不是為獻別樣的祭，
JOSH|22|27|而是為你我之間和後代子孫之間作證據，好使我們也在耶和華面前獻我們的燔祭、平安祭和別樣的祭來事奉他，免得你們的子孫將來對我們的子孫說，你們在耶和華裏無份。』
JOSH|22|28|所以我們說：『將來他們若對我們，或對我們的子孫這樣說，我們就可以回答說：你們看，我們列祖所築的壇是耶和華壇的樣式，這並不是為獻燔祭，也不是為獻別樣的祭，而是作為你們和我們之間的證據。』
JOSH|22|29|除了耶和華－我們上帝帳幕前的壇以外，我們絕沒有意思要為著獻燔祭、素祭和別樣的祭而另外築一座壇，悖逆耶和華，今日離棄不跟從他。」
JOSH|22|30|非尼哈 祭司與會眾中的領袖，就是與他同來那些 以色列 族系的領袖，聽見 呂便 人、 迦得 人、 瑪拿西 人所說的話，就都看為美。
JOSH|22|31|以利亞撒 祭司的兒子 非尼哈 對 呂便 人、 迦得 人、 瑪拿西 人說：「今日我們知道耶和華在我們中間，因為你們沒有向他犯悖逆的罪。現在你們把 以色列 人從耶和華的手中救出來了。」
JOSH|22|32|以利亞撒 祭司的兒子 非尼哈 與眾領袖離開了 呂便 人和 迦得 人，從 基列 地回 迦南 地，到了 以色列 人那裏，就把這事向他們回報。
JOSH|22|33|以色列 人看這事為美； 以色列 人就稱頌上帝，不再說要上去攻打 呂便 人和 迦得 人，毀壞他們所住的地了。
JOSH|22|34|呂便 人和 迦得 人給這壇起了名，因為這壇在我們之間見證耶和華是上帝。
JOSH|23|1|耶和華使 以色列 人從四圍所有的仇敵中得享安寧，已經有很多日子了。 約書亞 年紀老邁，
JOSH|23|2|就召了全 以色列 的眾長老、領袖、審判官和官長來，對他們說：「我年紀已經老邁。
JOSH|23|3|耶和華－你們的上帝因你們的緣故向這些國家所做的一切，你們都親眼看見了，那為你們作戰的是耶和華－你們的上帝。
JOSH|23|4|看，我已經把所剩下的列國，連同從 約旦河 起到 大海 日落的方向，我所剪除的列國，都抽籤分給你們各支派為業了。
JOSH|23|5|耶和華－你們的上帝必將他們從你們面前趕出去，使他們離開你們，你們就必得他們的地為業，正如耶和華－你們的上帝向你們所應許的。
JOSH|23|6|你們要大大壯膽，謹守遵行寫在 摩西 律法書上的一切話，不可偏離左右。
JOSH|23|7|不可與你們中間所剩下的這些國家往來。你們不可提他們神明的名，不可指著它們起誓，不可事奉它們，也不可敬拜它們。
JOSH|23|8|只要緊緊跟隨耶和華－你們的上帝，就像你們直到今日所做的。
JOSH|23|9|因為耶和華已經把又大又強的列國從你們面前趕出；直到今日，沒有一人能在你們面前站立得住。
JOSH|23|10|你們一人必追趕千人，因為耶和華－你們的上帝照他向你們所應許的，為你們作戰。
JOSH|23|11|你們要分外謹慎，愛耶和華－你們的上帝。
JOSH|23|12|你們若斷然轉離，緊緊跟隨你們中間所剩下的這些國家，彼此結親，互相往來，
JOSH|23|13|就要確實知道，耶和華－你們的上帝必不再將他們從你們面前趕出；他們卻要成為你們的羅網、圈套、肋上的鞭、眼中的刺，直到你們在耶和華－你們上帝所賜的這美地上滅亡。
JOSH|23|14|「看哪，我今日要走世人必走的路了。你們要一心一意知道，耶和華－你們上帝所應許要賜給你們的一切福氣，沒有一件落空，都應驗在你們身上了。
JOSH|23|15|耶和華－你們的上帝所應許的一切福氣怎樣臨到你們身上，耶和華也必照樣使各樣災禍臨到你們身上，直到他把你們從耶和華－你們上帝所賜給你們的這美地上除滅。
JOSH|23|16|你們若違背耶和華－你們上帝吩咐你們所守的約，去事奉別神，敬拜它們，耶和華的怒氣必向你們發作，使你們在他所賜給你們的美地上迅速滅亡。」
JOSH|24|1|約書亞 召集 以色列 的眾支派到 示劍 ，他召了 以色列 的長老、領袖、審判官和官長來；他們都站在上帝面前。
JOSH|24|2|約書亞 對眾百姓說：「耶和華－ 以色列 的上帝如此說：『古時你們的列祖，就是 亞伯拉罕 和 拿鶴 的父親 他拉 ，住在 大河 那邊事奉別神。
JOSH|24|3|我將你們的祖宗 亞伯拉罕 從 大河 那邊帶出來，領他走遍 迦南 全地，又使他的子孫眾多。我把 以撒 賜給他，
JOSH|24|4|我又把 雅各 和 以掃 賜給 以撒 ，將 西珥山 賜給 以掃 為業。但 雅各 和他的子孫下到 埃及 去了。
JOSH|24|5|我差遣 摩西 和 亞倫 ，照我在 埃及 中間所做的，降災與 埃及 ，然後把你們領出來。
JOSH|24|6|我領你們的祖宗出 埃及 ，你們就到了 紅海 。 埃及 人帶領戰車騎兵，追趕你們的祖宗到 紅海 。
JOSH|24|7|你們的祖宗哀求耶和華，他就用黑暗把你們和 埃及 人隔開了，又使海水衝向 埃及 人，淹沒他們。我在 埃及 所做的，你們都親眼見過。你們在曠野住了很多日子。
JOSH|24|8|我領你們到 約旦河 東 亞摩利 人所住之地。他們與你們爭戰，我把他們交在你們手中，你們就得了他們的地為業。我也在你們面前滅絕他們。
JOSH|24|9|那時， 摩押 王 西撥 的兒子 巴勒 起來攻擊 以色列 人，派人去召 比珥 的兒子 巴蘭 來詛咒你們。
JOSH|24|10|但我不願聽 巴蘭 ，所以他反而為你們連連祝福。這樣，我救了你們脫離他的手。
JOSH|24|11|你們過了 約旦河 ，來到 耶利哥 。 耶利哥 人、 亞摩利 人、 比利洗 人、 迦南 人、 赫 人、 革迦撒 人、 希未 人、 耶布斯 人都與你們爭戰，我卻把他們交在你們手裏。
JOSH|24|12|我派遣瘟疫 在你們前面，將 亞摩利 人的兩個王從你們面前趕出，並不是用你的刀，也不是用你的弓。
JOSH|24|13|我賜給你們的地，不是你們開墾的；我賜給你們的城鎮，不是你們建造的。你們卻住在其中，又得吃那不是你們栽植的葡萄園和橄欖園的果子。』
JOSH|24|14|「現在你們要敬畏耶和華，誠心誠意事奉他，除掉你們列祖在 大河 那邊和在 埃及 事奉的神明，事奉耶和華。
JOSH|24|15|若你們認為事奉耶和華不好，今日就可以選擇所要事奉的：是你們列祖在 大河 那邊所事奉的神明，或是你們所住這地 亞摩利 人的神明呢？至於我和我家，我們必定事奉耶和華。」
JOSH|24|16|百姓回答說：「我們絕不離棄耶和華去事奉別神。
JOSH|24|17|因為耶和華－我們的上帝曾領我們和我們的祖宗從 埃及 地為奴之家出來，在我們眼前行了那些大神蹟，並在我們所行的一切路上，和所經過的各民族中保護了我們。
JOSH|24|18|耶和華又把各民族和住此地的 亞摩利 人都從我們面前趕出去。所以，我們也必事奉耶和華，因為他是我們的上帝。」
JOSH|24|19|約書亞 對百姓說：「你們不能事奉耶和華，因為他是神聖的上帝，是忌邪 的上帝，必不赦免你們的過犯罪惡。
JOSH|24|20|你們若離棄耶和華去事奉外邦的神明，耶和華在降福之後，必轉而降禍給你們，把你們滅絕。」
JOSH|24|21|百姓對 約書亞 說：「不，我們要事奉耶和華。」
JOSH|24|22|約書亞 對百姓說：「你們選擇耶和華，要事奉他，你們自己作證吧！」他們說：「我們願意作證。」
JOSH|24|23|「現在，你們要除掉你們中間外邦的神明，專心歸向耶和華－ 以色列 的上帝。」
JOSH|24|24|百姓對 約書亞 說：「我們必事奉耶和華－我們的上帝，聽從他的話。」
JOSH|24|25|那日， 約書亞 就與百姓立約，在 示劍 為他們制定律例典章。
JOSH|24|26|約書亞 把這些話寫在上帝的律法書上，又拿一塊大石頭立在橡樹下耶和華聖所的旁邊。
JOSH|24|27|約書亞 對眾百姓說：「看哪，這石頭可以向我們作見證，因為它聽見了耶和華所吩咐我們的一切話；這石頭將向你們作見證，免得你們背叛你們的上帝。」
JOSH|24|28|於是 約書亞 解散百姓，各自回到自己的地業去了。
JOSH|24|29|這些事以後，耶和華的僕人， 嫩 的兒子 約書亞 死了，那時他一百一十歲。
JOSH|24|30|以色列 人把他葬在他自己地業的境內， 以法蓮 山區的 亭拿‧西拉 ，在 迦實山 的北邊。
JOSH|24|31|約書亞 在世的日子和他死了以後，那些知道耶和華為 以色列 所做一切事的長老還在世的時候， 以色列 人事奉耶和華。
JOSH|24|32|以色列 人把從 埃及 所帶來 約瑟 的骸骨安葬在 示劍 ，就是 雅各 從前用一百可錫塔 向 示劍 的父親 哈抹 的眾子所買的那塊地；這塊地就成了 約瑟 子孫的產業。
JOSH|24|33|亞倫 的兒子 以利亞撒 也死了，他們把他葬在他兒子 非尼哈 所得 以法蓮 山區的小山上 。
JUDG|1|1|約書亞 死後， 以色列 人求問耶和華說：「我們中間誰當首先上去攻打 迦南 人，與他們爭戰呢？」
JUDG|1|2|耶和華說：「 猶大 要先上去。看哪，我已將那地交在他手中。」
JUDG|1|3|猶大 對他哥哥 西緬 說：「請你同我上到我抽籤所得之地，與 迦南 人爭戰；我也同你去你抽籤所得之地。」於是 西緬 與他同去。
JUDG|1|4|猶大 就上去，耶和華把 迦南 人和 比利洗 人交在他們手中。他們在 比色 擊殺了一萬人。
JUDG|1|5|他們在 比色 遇見 亞多尼‧比色 ，與他爭戰，擊敗了 迦南 人和 比利洗 人。
JUDG|1|6|亞多尼‧比色 逃跑，他們追趕他，捉住他，砍斷他大拇指和大腳趾。
JUDG|1|7|亞多尼‧比色 說：「從前有七十個王，大拇指和大腳趾都被我砍斷，在我桌子底下拾取零碎食物。現在上帝照著我所做的報應我了。」他們把 亞多尼‧比色 帶到 耶路撒冷 ，他就死在那裏。
JUDG|1|8|猶大 人攻打 耶路撒冷 ，奪取了它，用刀殺城內的人，並且放火燒城。
JUDG|1|9|後來 猶大 人下去，與住山區、 尼革夫 和低地的 迦南 人爭戰。
JUDG|1|10|猶大 去攻打住 希伯崙 的 迦南 人，殺了 示篩 、 亞希幔 、 撻買 。 希伯崙 從前名叫 基列‧亞巴 。
JUDG|1|11|猶大 從那裏去攻擊 底壁 的居民。 底壁 從前名叫 基列‧西弗 。
JUDG|1|12|迦勒 說：「誰能攻打 基列‧西弗 ，奪取那城，我就把我女兒 押撒 嫁給他。」
JUDG|1|13|迦勒 的弟弟 基納斯 的兒子 俄陀聶 奪取了那城， 迦勒 就把女兒 押撒 嫁給他。
JUDG|1|14|押撒 來的時候，催促丈夫 向她父親要一塊田。 押撒 一下驢， 迦勒 就對她說：「你要甚麼？」
JUDG|1|15|她對 迦勒 說：「求你賜我福分；你既然把 尼革夫 給了我，求你也給我水泉。」 迦勒 就把上泉和下泉都賜給她。
JUDG|1|16|摩西 的岳父是 基尼 人，他的子孫與 猶大 人一起上到棕樹城，往 亞拉得 以南的 猶大 曠野 去，住在百姓當中 。
JUDG|1|17|猶大 和他哥哥 西緬 同去，擊殺了住 洗法 的 迦南 人，將城徹底毀滅。因此，那城名叫 何珥瑪 。
JUDG|1|18|猶大 攻取了 迦薩 和所屬的領土， 亞實基倫 和所屬的領土， 以革倫 和所屬的領土。
JUDG|1|19|耶和華與 猶大 同在， 猶大 取得了山區，卻不能趕出平原的居民，因為他們有鐵的戰車。
JUDG|1|20|以色列 人照 摩西 所說的，把 希伯崙 給了 迦勒 。 迦勒 從那裏趕出 亞衲 的三支後裔。
JUDG|1|21|至於住 耶路撒冷 的 耶布斯 人， 便雅憫 人沒有把他們趕出。於是， 耶布斯 人與 便雅憫 人同住在 耶路撒冷 ，直到今日。
JUDG|1|22|約瑟 家也上到 伯特利 去，耶和華與他們同在。
JUDG|1|23|約瑟 家去窺探 伯特利 ，那城起先名叫 路斯 。
JUDG|1|24|探子看見一個人從城裏出來，就對他說：「請你把進城的路指示我們，我們會厚待你。」
JUDG|1|25|那人把進城的路指示他們。他們就用刀擊殺了城中的居民，卻放走那人和他的全家。
JUDG|1|26|那人往 赫 人之地去，建造了一座城，起名叫 路斯 。那城到如今還叫這名。
JUDG|1|27|瑪拿西 沒有趕出 伯˙善 和所屬鄉鎮 的居民， 他納 和所屬鄉鎮的居民， 多珥 和所屬鄉鎮的居民， 以伯蓮 和所屬鄉鎮的居民， 米吉多 和所屬鄉鎮的居民； 迦南 人仍堅持住在這地。
JUDG|1|28|以色列 強盛的時候，就叫 迦南 人做苦工，沒有把他們全然趕走。
JUDG|1|29|以法蓮 沒有趕出住 基色 的 迦南 人。於是 迦南 人仍住在 基色 ，在 以法蓮 中間。
JUDG|1|30|西布倫 沒有趕出 基倫 的居民和 拿哈拉 的居民。於是 迦南 人仍住在 西布倫 中間，成了服勞役的人。
JUDG|1|31|亞設 沒有趕出 亞柯 的居民和 西頓 的居民，以及 亞黑拉 、 亞革悉 、 黑巴 、 亞弗革 和 利合 的居民。
JUDG|1|32|亞設 人因為沒有趕出那地的居民 迦南 人，就住在他們中間。
JUDG|1|33|拿弗他利 沒有趕出 伯˙示麥 和 伯˙亞納 的居民。於是 拿弗他利 就住在那地的居民 迦南 人中，而 伯˙示麥 和 伯˙亞納 的居民卻成了為他們服勞役的人。
JUDG|1|34|亞摩利 人強逼 但 人住在山區，不准他們下到平原。
JUDG|1|35|亞摩利 人仍堅持住在 希烈山 、 亞雅崙 和 沙賓 ；然而 約瑟 家權勢強盛的時候，他們成為服勞役的人。
JUDG|1|36|亞摩利 人 的地界是從 亞克拉濱 斜坡，從 西拉 延伸而上。
JUDG|2|1|耶和華的使者從 吉甲 上到 波金 ，說：「我領你們從 埃及 上來，帶你們到我向你們列祖起誓應許之地。我曾說：『我永不廢棄我與你們的約。
JUDG|2|2|你們不可與這地的居民立約，要拆毀他們的祭壇。』你們竟沒有聽從我的話。你們為何這樣做呢！
JUDG|2|3|因此我說：『我必不將他們從你們面前趕出。他們必作你們肋下的荊棘 ，他們的神明必成為你們的圈套。』」
JUDG|2|4|耶和華的使者向 以色列 眾人說這些話的時候，百姓放聲大哭。
JUDG|2|5|於是他們給那地方起名叫 波金 ，並在那裏向耶和華獻祭。
JUDG|2|6|約書亞 解散百姓， 以色列 人回到自己的地業，佔各自的地。
JUDG|2|7|約書亞 在世的日子和他死了以後，那些見過耶和華為 以色列 所做一切大事的長老還在世的時候，百姓都事奉耶和華。
JUDG|2|8|耶和華的僕人， 嫩 的兒子 約書亞 死了，那時他一百一十歲。
JUDG|2|9|以色列 人把他葬在他自己地業的境內， 以法蓮 山區的 亭拿‧希烈 ，在 迦實山 的北邊。
JUDG|2|10|那世代的人也都歸到自己的列祖。後來興起的另一世代不認識耶和華，也不知道他為 以色列 所做的事。
JUDG|2|11|以色列 人行耶和華眼中看為惡的事，去事奉諸 巴力 。
JUDG|2|12|他們離棄領他們出 埃及 地的耶和華－他們列祖的上帝，去隨從別神，就是四圍列國的神明，向它們叩拜，惹耶和華發怒。
JUDG|2|13|他們離棄了耶和華，去事奉 巴力 和 亞斯她錄 。
JUDG|2|14|耶和華的怒氣向 以色列 發作，把他們交在搶奪他們的人手中，又把他們交給四圍仇敵的手中 ，以致他們在仇敵面前再也不能站立得住。
JUDG|2|15|他們無論往何處去，耶和華的手都以災禍攻擊他們，正如耶和華所說的，又如耶和華向他們所起的誓；他們就極其困苦。
JUDG|2|16|耶和華興起士師，士師就拯救他們脫離搶奪他們之人的手。
JUDG|2|17|然而，他們卻不聽從士師，竟隨從別神而行淫，向它們叩拜。他們列祖所行的道，所聽從耶和華的命令，他們都速速偏離了，並不照樣遵行。
JUDG|2|18|耶和華為他們興起士師，耶和華與士師同在。士師在世的一切日子，耶和華拯救他們脫離仇敵的手。耶和華因他們受欺壓迫害所發出的哀聲，就憐憫他們。
JUDG|2|19|但士師一死，他們又轉去行惡，比他們祖宗更壞，去隨從別神，事奉叩拜它們，總不放棄他們的惡習和頑梗的行為。
JUDG|2|20|於是耶和華的怒氣向 以色列 發作，說：「因為這國違背我吩咐他們列祖當守的約，不聽從我的話，
JUDG|2|21|約書亞 死的時候所剩下的各國，我必不再從他們面前趕出任何一個，
JUDG|2|22|為要藉此考驗 以色列 是否肯謹守遵行耶和華的道，像他們列祖一樣地謹守。」
JUDG|2|23|耶和華留下那些國家，不將他們速速趕出，也不把他們交在 約書亞 的手中。
JUDG|3|1|耶和華留下這些國家，為要考驗所有未曾經歷 迦南 任何戰役的 以色列 人，
JUDG|3|2|只是為了要 以色列 人的後代認識戰爭，教導他們，尤其那些未曾認識這些事的人。
JUDG|3|3|留下的有 非利士 的五個領袖，所有的 迦南 人， 西頓 人，以及從 巴力‧黑門山 到 哈馬口 ，住 黎巴嫩山 的 希未 人。
JUDG|3|4|他們是為了要考驗 以色列 ，好知道他們是否肯聽從耶和華藉 摩西 吩咐他們列祖的命令。
JUDG|3|5|以色列 人住在 迦南 人、 赫 人、 亞摩利 人、 比利洗 人、 希未 人、 耶布斯 人中間，
JUDG|3|6|娶他們的女兒，將自己的女兒嫁給他們的兒子，並事奉他們的神明。
JUDG|3|7|以色列 人行耶和華眼中看為惡的事，忘記耶和華－他們的上帝，去事奉諸 巴力 和 亞舍拉 ，
JUDG|3|8|所以耶和華的怒氣向 以色列 發作，把他們交給 美索不達米亞 王 古珊‧利薩田 的手中。 以色列 人服事 古珊‧利薩田 八年。
JUDG|3|9|以色列 人呼求耶和華，耶和華就為 以色列 人興起一位拯救者來救他們，就是 迦勒 的弟弟 基納斯 的兒子 俄陀聶 。
JUDG|3|10|耶和華的靈降在他身上，他就作了 以色列 的士師。他出去爭戰，耶和華將 亞蘭 王 古珊‧利薩田 交在他手中，他的手戰勝了 古珊‧利薩田 。
JUDG|3|11|於是這地太平四十年。 基納斯 的兒子 俄陀聶 死了。
JUDG|3|12|以色列 人又行耶和華眼中看為惡的事。耶和華使 摩押 王 伊磯倫 強大，攻擊 以色列 ，因為他們行耶和華眼中看為惡的事。
JUDG|3|13|伊磯倫 召集 亞捫 人和 亞瑪力 人到他那裏，他就去攻打 以色列 ，佔據了棕樹城。
JUDG|3|14|於是 以色列 人服事 摩押 王 伊磯倫 十八年。
JUDG|3|15|以色列 人呼求耶和華，耶和華就為他們興起一位拯救者， 便雅憫 人 基拉 的兒子 以笏 ，他是個慣用左手的人 。 以色列 人託他送禮物給 摩押 王 伊磯倫 。
JUDG|3|16|以笏 打造了一把兩刃的劍，長一短肘 ，綁在右腿上衣服裏面。
JUDG|3|17|他把禮物獻給 摩押 王 伊磯倫 。 伊磯倫 是個很肥胖的人。
JUDG|3|18|以笏 獻完禮物的時候，就把抬禮物的人送走。
JUDG|3|19|但他自己卻從靠近 吉甲 的雕像那裏轉回來，說：「王啊，我有一件機密的事要奏告你。」王說：「迴避吧！」於是所有侍立在他左右的人都退去了。
JUDG|3|20|以笏 來到王那裏，那時他獨自一人坐在陰涼的頂樓。 以笏 說：「我有上帝的話向你報告。」王就從座位上站起來。
JUDG|3|21|以笏 伸出左手，從右腿上拔出劍來，刺入王的肚腹。
JUDG|3|22|劍柄連同劍刃都刺進去了，肥肉夾住了劍刃。他沒有把劍從王的肚腹拔出來，糞便就流出來了 。
JUDG|3|23|以笏 出到門廊，把王關在樓門裏面，就上了鎖。
JUDG|3|24|以笏 出來之後，王的僕人就來了。他們觀看，看哪，樓門鎖住，就說：「他必是在陰涼的房間裏大解。」
JUDG|3|25|他們等得不耐煩，看哪，樓門仍然不開，就拿鑰匙打開樓門，看哪，他們的主人已經倒在地上死了。
JUDG|3|26|他們耽延的時候， 以笏 就逃跑了。他經過雕像那裏，逃到 西伊拉 。
JUDG|3|27|他到了那裏，就在 以法蓮 山區吹角。 以色列 人跟隨他從山區下來，他在他們前面引路，
JUDG|3|28|對他們說：「緊跟著我！因為耶和華已經把你們的仇敵 摩押 交在你們手中。」於是他們跟著他下去，佔據了 摩押 對面 約旦河 的渡口，不准一人過去。
JUDG|3|29|那時，他們擊殺了約一萬 摩押 人，都是強壯的勇士，連一個也沒有逃脫。
JUDG|3|30|那日， 摩押 在 以色列 手下制伏了。於是這地太平八十年。
JUDG|3|31|以笏 之後，有 亞拿 的兒子 珊迦 ，他用趕牛的棍子打死六百 非利士 人。他也拯救了 以色列 。
JUDG|4|1|以笏 死後， 以色列 人又行耶和華眼中看為惡的事。
JUDG|4|2|耶和華把他們交給在 夏瑣 作王的 迦南 王 耶賓 手中；他的將軍是 西西拉 ，住在 夏羅設‧哈歌印 。
JUDG|4|3|以色列 人呼求耶和華，因為 耶賓 王有鐵的戰車九百輛，並且殘酷欺壓 以色列 人二十年。
JUDG|4|4|有一位女先知 底波拉 ，是 拉比多 的妻子，當時作 以色列 的士師。
JUDG|4|5|她住在 以法蓮 山區 拉瑪 和 伯特利 的中間，在 底波拉 的棕樹下。 以色列 人都上到她那裏去聽審判。
JUDG|4|6|她派人從 拿弗他利 的 基低斯 把 亞比挪菴 的兒子 巴拉 召來，對他說：「耶和華－ 以色列 的上帝吩咐你：『你要率領一萬 拿弗他利 人和 西布倫 人上 他泊山 去。
JUDG|4|7|我必使 耶賓 的將軍 西西拉 率領他的戰車和全軍往 基順河 ，到你那裏去，我必把他交在你手中。』」
JUDG|4|8|巴拉 對她說：「你若同我去，我就去；你若不同我去，我就不去。」
JUDG|4|9|底波拉 說：「我一定會與你同去，然而你在所行的路上必得不著榮耀，因為耶和華要把 西西拉 交給一個婦人的手裏。」於是 底波拉 起來，與 巴拉 一同往 基低斯 去了。
JUDG|4|10|巴拉 召集 西布倫 人和 拿弗他利 人到 基低斯 ，跟他上去的有一萬人。 底波拉 也同他上去。
JUDG|4|11|摩西 岳父 何巴 的後裔， 基尼 人 希百 離開了 基尼 族，到靠近 基低斯 的 撒拿音 橡樹旁支搭帳棚。
JUDG|4|12|有人告訴 西西拉 ：「 亞比挪菴 的兒子 巴拉 已經上了 他泊山 。」
JUDG|4|13|西西拉 就召集所有的鐵戰車九百輛和隨從的全軍，從 夏羅設‧哈歌印 出來，到了 基順河 。
JUDG|4|14|底波拉 對 巴拉 說：「起來，今日就是耶和華把 西西拉 交在你手中的日子。耶和華豈不在你前面行嗎?」於是 巴拉 下了 他泊山 ，跟隨他的有一萬人。
JUDG|4|15|耶和華使 西西拉 和他一切的戰車，以及全軍潰亂，在 巴拉 面前倒在刀下。 西西拉 下了車，徒步逃跑。
JUDG|4|16|巴拉 追趕戰車、軍隊，直到 夏羅設‧哈歌印 。 西西拉 的全軍都倒在刀下，一個也沒有留下。
JUDG|4|17|只有 西西拉 徒步逃跑到 基尼 人 希百 之妻 雅億 的帳棚，因為 夏瑣 王 耶賓 與 基尼 人的 希百 家和平共處。
JUDG|4|18|雅億 出來迎接 西西拉 ，對他說：「請我主進來，進到我這裏來，不要怕。」 西西拉 就進了她的帳棚， 雅億 用被子將他蓋住。
JUDG|4|19|西西拉 對 雅億 說：「我渴了，求你給我一點水喝。」 雅億 就打開裝奶的皮袋，給他喝，再把他蓋住。
JUDG|4|20|西西拉 對 雅億 說：「請你站在帳棚門口，若有人來問你說：『有人在這裏嗎？』你就說：『沒有。』」
JUDG|4|21|西西拉 疲乏沉睡了。 希百 的妻 雅億 取了帳棚的橛子，手拿著錘子，靜悄悄地到他那裏，將橛子從他的太陽穴釘進去，直釘到地裏。 西西拉 就死了。
JUDG|4|22|看哪， 巴拉 追趕 西西拉 ， 雅億 出來迎接他，對他說：「來，我給你看你要找的人。」他就進入帳棚，看哪， 西西拉 已經倒在地上死了，橛子還在他的太陽穴中。
JUDG|4|23|那日，上帝在 以色列 人面前制伏了 迦南 王 耶賓 。
JUDG|4|24|從此， 以色列 人的手對 迦南 王 耶賓 越來越強硬，直到將 迦南 王 耶賓 剪除。
JUDG|5|1|那日， 底波拉 和 亞比挪菴 的兒子 巴拉 唱歌，說：
JUDG|5|2|「 以色列 有領袖率領 ， 百姓甘心犧牲自己， 你們當稱頌耶和華！
JUDG|5|3|「君王啊，要聽！王子啊，要側耳！ 我要，我要向耶和華歌唱； 我要歌頌耶和華－ 以色列 的上帝。
JUDG|5|4|「耶和華啊，你從 西珥 出來， 從 以東 田野向前行， 地震動 天滴下， 雲也滴下雨水。
JUDG|5|5|眾山在耶和華面前搖動， 西奈山 在耶和華－ 以色列 上帝面前也搖動。
JUDG|5|6|「在 亞拿 之子 珊迦 的時候， 在 雅億 的日子， 大道無人行走， 過路人繞道而行。
JUDG|5|7|以色列 農村荒蕪， 空無一人， 直到我 底波拉 興起， 興起作 以色列 之母！
JUDG|5|8|以色列 人選擇新的諸神， 戰爭就臨到城門。 以色列 四萬人中， 看得見盾牌槍矛嗎？
JUDG|5|9|我心嚮往 以色列 的領袖， 他們在民中甘心犧牲自己。 你們應當稱頌耶和華！
JUDG|5|10|「騎淺色母驢的、 坐繡花毯子的、 行走在路上的， 你們都當思想！
JUDG|5|11|打水的聲音勝過弓箭的響聲， 那裏，人要述說耶和華公義的作為， 他對 以色列 鄉民公義的作為。 「那時，耶和華的子民下到城門。
JUDG|5|12|「 底波拉 啊，興起！興起！ 當興起，興起，唱歌！ 巴拉 啊，你當興起！ 亞比挪菴 的兒子啊，當俘擄你的俘虜！
JUDG|5|13|那時，貴族中的倖存者前進， 耶和華的百姓為我前進攻擊勇士。
JUDG|5|14|源自 亞瑪力 的人從 以法蓮 下來 ， 跟著你，你的族人 便雅憫 ； 有領袖從 瑪吉 下來， 手握官員權杖的從 西布倫 下來。
JUDG|5|15|以薩迦 的領袖與 底波拉 一起； 巴拉 怎樣， 以薩迦 也怎樣； 他跟隨 巴拉 衝下平原。 呂便 支派 有胸懷大志的人。
JUDG|5|16|你為何坐在羊圈內， 聽羊群中吹笛的聲音呢？ 呂便 支派具心有大謀的人。
JUDG|5|17|基列 安居在 約旦河 東。 但 為何住在船上呢？ 亞設 在海邊居住， 它在港口安居。
JUDG|5|18|西布倫 是拚命敢死的百姓， 拿弗他利 在田野的高處也是如此。 　
JUDG|5|19|「君王都來爭戰； 那時 迦南 諸王在 米吉多 水旁的 他納 爭戰， 卻得不到擄掠的銀錢。
JUDG|5|20|星宿從天上爭戰， 從它們的軌道攻擊 西西拉 。
JUDG|5|21|基順 的急流沖走他們， 古老的急流， 基順 的急流。 我的靈啊，努力前進！
JUDG|5|22|「那時馬蹄踢踏， 壯馬奔馳飛騰。
JUDG|5|23|「耶和華的使者說：『要詛咒 米羅斯 ， 重重詛咒其中的居民， 因為他們不來幫助耶和華， 不來幫助耶和華攻擊壯士。』
JUDG|5|24|「願 基尼 人 希百 的妻子 雅億 比眾婦人多得福氣， 比帳棚中的婦人更蒙福祉。
JUDG|5|25|西西拉 求水， 雅億 給他奶， 用貴重的碗裝乳酪給他。
JUDG|5|26|雅億 左手拿著帳棚的橛子， 右手拿著工匠的錘子， 擊打 西西拉 ，打碎他的頭， 打破穿透他的太陽穴。
JUDG|5|27|西西拉 在她腳下曲身，仆倒，躺臥， 在她腳下曲身，仆倒； 他在哪裏曲身，就在哪裏仆倒，死亡。
JUDG|5|28|「 西西拉 的母親從窗戶裏往外觀看， 她在窗格子中哀號： 『他的戰車為何遲遲未歸？ 他的車輪為何走得那麼慢呢？』
JUDG|5|29|她聰明的宮女回答她， 她也自言自語說：
JUDG|5|30|『或許他們得了戰利品而分， 每個壯士得了一兩個女子？ 西西拉 得了彩衣為擄物， 得了繡花的彩衣為掠物， 這兩面繡花的彩衣， 披在頸項上作為戰利品。』
JUDG|5|31|「耶和華啊，願你的仇敵都這樣滅亡！ 願愛你的人如太陽上升，大發光輝！」 於是這地太平四十年。
JUDG|6|1|以色列 人又行耶和華眼中看為惡的事，耶和華就把他們交在 米甸 手裏七年。
JUDG|6|2|米甸 的手戰勝 以色列 ； 以色列 人躲避 米甸 人，就在山中挖洞穴，挖洞建營寨。
JUDG|6|3|每當 以色列 人撒種之後， 米甸 、 亞瑪力 和東邊的人都上來攻打他們，
JUDG|6|4|對著他們安營，毀壞那地的農作物，直到 迦薩 ，沒有給 以色列 留下食物，牛、羊、驢也沒有留下。
JUDG|6|5|因為那些人帶著他們的牲畜和帳棚上來，像蝗蟲那樣多；人和駱駝無數，都進入境內，毀壞全地。
JUDG|6|6|以色列 因 米甸 的緣故極其窮乏， 以色列 人就呼求耶和華。
JUDG|6|7|以色列 人因 米甸 的緣故呼求耶和華的時候，
JUDG|6|8|耶和華就差遣先知到 以色列 人那裏，對他們說：「耶和華－ 以色列 的上帝如此說：『我曾領你們從 埃及 上來，從為奴之家出來，
JUDG|6|9|救你們脫離 埃及 人的手，脫離一切欺壓你們之人的手。我從你們面前趕出他們，把他們的地賜給你們。
JUDG|6|10|我對你們說，我是耶和華－你們的上帝。你們住在 亞摩利 人的地，不可敬畏他們的神明，但你們卻不聽從我的話。』」
JUDG|6|11|耶和華的使者到了 俄弗拉 ，坐在 亞比以謝 族 約阿施 的橡樹下。 約阿施 的兒子 基甸 正在醡酒池那裏打麥子，為了躲避 米甸 人。
JUDG|6|12|耶和華的使者向 基甸 顯現，對他說：「大能的勇士啊，耶和華與你同在！」
JUDG|6|13|基甸 對他說：「主啊，請容許我說，耶和華若與我們同在，我們怎麼會遭遇這一切事呢？我們的列祖告訴我們：『耶和華領我們從 埃及 上來』，他那奇妙的作為在哪裏呢？現在耶和華卻丟棄了我們，把我們交在 米甸 人的手掌中。」
JUDG|6|14|耶和華轉向 基甸 ，說：「去，靠著你這能力拯救 以色列 脫離 米甸 人的手掌。我豈不是已經差遣了你嗎？」
JUDG|6|15|基甸 對他說：「主啊，請容許我說，我怎能拯救 以色列 呢？看哪，我這一支在 瑪拿西 支派中是最貧寒的，我在我父家又是最微小的。」
JUDG|6|16|耶和華對他說：「我與你同在，你就必擊敗 米甸 ，如擊打一個人。」
JUDG|6|17|基甸 對他說：「我若在你眼前蒙恩，求你給我一個證據，證明是你在跟我說話。
JUDG|6|18|求你不要離開這裏，等我回來，將供物帶來，供在你面前。」他說：「我必等你回來。」
JUDG|6|19|基甸 去預備一隻小山羊，用一伊法細麵做了無酵餅，將肉放在籃子裏，將湯盛在壺中，帶到他那裏，在橡樹下獻上。
JUDG|6|20|上帝的使者對 基甸 說：「將肉和無酵餅放在這磐石上，把湯倒出來。」他就照樣做了。
JUDG|6|21|耶和華的使者伸出手裏的杖，杖頭一碰到肉和無酵餅，就有火從磐石中出來，吞滅了肉和無酵餅。耶和華的使者就從他眼前消失了。
JUDG|6|22|基甸 見他是耶和華的使者，就說：「哎呀！主耶和華啊！因為我真的面對面看見了耶和華的使者。」
JUDG|6|23|耶和華對他說：「安心吧，不要怕，你不會死。」
JUDG|6|24|於是 基甸 在那裏為耶和華築了一座壇，起名叫「耶和華沙龍」 。這壇至今還在 亞比以謝 族的 俄弗拉 。
JUDG|6|25|那夜，耶和華對 基甸 說：「你要把你父親的公牛，就是 那七歲的第二頭公牛取來，並拆毀你父親為 巴力 築的壇，砍下壇旁的 亞舍拉 ，
JUDG|6|26|在這堡壘頂上整整齊齊地為耶和華－你的上帝築一座壇，將第二頭公牛獻為燔祭，用你所砍下的 亞舍拉 當柴。」
JUDG|6|27|基甸 就從他僕人中選了十個人，照耶和華吩咐他的做了。他因怕父家和本城的人，不敢在白天做這事，就在夜間做。
JUDG|6|28|城裏的人清早起來，看哪， 巴力 的壇被拆毀，壇旁的 亞舍拉 被砍下，第二頭公牛獻在築好的壇上，
JUDG|6|29|就彼此問：「這是誰做的事呢？」他們尋找查訪之後，就說：「這是 約阿施 的兒子 基甸 做的事。」
JUDG|6|30|城裏的人對 約阿施 說：「把你的兒子交出來，我們要處死他，因為他拆毀了 巴力 的壇，砍下了壇旁的 亞舍拉 。」
JUDG|6|31|約阿施 對站著敵對他的眾人說：「你們是為 巴力 辯護嗎？你們要救它嗎？誰為它辯護，就在早晨把誰處死吧！ 巴力 如果是上帝，有人拆毀了它的壇，就讓它為自己辯護吧！」
JUDG|6|32|所以那日人稱 基甸 為 耶路巴力 ，意思是：「他拆毀了 巴力 的壇，讓 巴力 與他爭辯吧。」
JUDG|6|33|那時，所有的 米甸 人、 亞瑪力 人和東邊的人都聚集在一起，過了河，在 耶斯列 平原安營。
JUDG|6|34|耶和華的靈降在 基甸 身上；他吹角， 亞比以謝 族都聚集跟隨他。
JUDG|6|35|他派使者走遍 瑪拿西 ， 瑪拿西 人也聚集跟隨他。他又派使者到 亞設 、 西布倫 、 拿弗他利 ，他們也都上來會合。
JUDG|6|36|基甸 對上帝說：「你如果真的照你所說的，藉我的手拯救 以色列 ，
JUDG|6|37|看哪，我把一團羊毛放在禾場上，若單是羊毛上有露水，遍地都是乾的，我就知道你必照你所說的，藉我的手拯救 以色列 。」
JUDG|6|38|一切果然發生了。次日早晨 基甸 起來，把羊毛擰一擰，從羊毛中擠出露水來，裝滿一碗的水。
JUDG|6|39|基甸 又對上帝說：「求你不要向我發怒，我再說一次，讓我用羊毛再試一次，但願羊毛是乾的，遍地都有露水。」
JUDG|6|40|這夜，上帝也照樣做，遍地都有露水，只有羊毛是乾的。
JUDG|7|1|耶路巴力 ，就是 基甸 ，和所有跟隨他的人早晨起來，在 哈律泉 旁安營。 米甸 營在他北邊，靠近 摩利岡 的平原。
JUDG|7|2|耶和華對 基甸 說：「跟隨你的人太多，我不能把 米甸 交在他們手中，免得 以色列 向我自誇，說：『是我自己的手救了我。』
JUDG|7|3|現在你要向這百姓宣告說：『凡懼怕戰兢的，可以離開 基列山 回去。』」於是有二萬二千人回去，只剩下一萬人。
JUDG|7|4|耶和華對 基甸 說：「人還是太多。你要帶他們下到水旁，我好在那裏為你試試他們。我指著誰對你說：『這人可以跟你去』，他就可以跟你去；我指著誰對你說：『這人不可跟你去』，他就不可跟你去。」
JUDG|7|5|基甸 就帶百姓下到水旁。耶和華對 基甸 說：「凡用舌頭舔水像狗一樣舔的，要使他單獨站在一處；那些用雙膝跪下喝水的，也要使他單獨站在一處。」
JUDG|7|6|用手捧到嘴邊舔水的數目有三百人，其餘的百姓都用雙膝跪下喝水。
JUDG|7|7|耶和華對 基甸 說：「我要用這舔水的三百人拯救你們，把 米甸 交在你手中；其餘的百姓都可以各回自己的地方去。」
JUDG|7|8|百姓手裏拿著食物和角；其餘的 以色列 人， 基甸 都打發他們各自回到自己的帳棚，只留下這三百人。 米甸 營在他下邊的平原上。
JUDG|7|9|那夜，耶和華對 基甸 說：「起來，下去攻營，因我已把它交在你手中。
JUDG|7|10|倘若你害怕下去，可以帶你的僕人 普拉 下到那營裏去，
JUDG|7|11|你必聽見他們所說的，這樣你的手就有力量下去攻營。」於是 基甸 帶著僕人 普拉 下到軍營裏帶著兵器的人邊上。
JUDG|7|12|米甸 人、 亞瑪力 人和所有東邊的人都散佈在平原，如同蝗蟲那樣多。他們的駱駝無數，多如海邊的沙。
JUDG|7|13|基甸 到了那裏，看哪，有一人把夢告訴同伴說：「看哪，我做了一個夢。看哪，一個大麥餅滾入 米甸 營中，來到帳幕，把帳幕撞倒，帳幕就翻轉倒塌了。」
JUDG|7|14|同伴回答說：「這不是別的，而是 以色列 人 約阿施 的兒子 基甸 的刀。上帝已把 米甸 和全軍都交在他手中了。」
JUDG|7|15|基甸 聽見這夢的敘述和夢的解釋，就敬拜上帝。他回到 以色列 營中，說：「起來吧！耶和華已把 米甸 軍隊交在你們手中了。」
JUDG|7|16|於是 基甸 將三百人分成三隊，把角和空瓶交在每個人手中，瓶內有火把。
JUDG|7|17|他對他們說：「看著我，你們要照樣做。看哪，我來到營邊，我怎樣做，你們也要照樣做。
JUDG|7|18|我和所有跟隨我的人吹角的時候，你們也要在營的四圍吹角，喊叫：『為耶和華！為 基甸 ！』」
JUDG|7|19|基甸 和跟隨他的一百人，在半夜之初換崗哨的時候來到營旁。他們就吹角，打破手中的瓶；
JUDG|7|20|三隊的人都吹角，打破瓶子。他們左手拿著火把，右手拿著吹的角，喊叫：「耶和華和 基甸 的刀！」
JUDG|7|21|他們圍著軍營，各人站在自己的地方；全營的人都逃竄，一面喊，一面逃跑。
JUDG|7|22|三百人就吹角，耶和華使全營的人用刀自相擊殺。全營的人逃往 西利拉 的 伯‧哈示他 ，一直逃到靠近 他巴 的 亞伯‧米何拉 。
JUDG|7|23|從 拿弗他利 、 亞設 和 瑪拿西 全地來的 以色列 人被召來，追趕 米甸 人。
JUDG|7|24|基甸 也派人走遍 以法蓮 山區，說：「你們下來迎擊 米甸 人，在他們的前面沿著 約旦河 把守渡口，直到 伯‧巴拉 。」於是 以法蓮 眾人聚集，沿著 約旦河 把守渡口，直到 伯‧巴拉 。
JUDG|7|25|他們捉住了 米甸 的兩個領袖， 俄立 和 西伊伯 。他們在 俄立 磐石上殺了 俄立 ，在 西伊伯 酒池那裏殺了 西伊伯 。他們追趕 米甸 人，把 俄立 和 西伊伯 的首級帶到 約旦河 對岸，到 基甸 那裏。
JUDG|8|1|以法蓮 人對 基甸 說：「你去與 米甸 爭戰，沒有召我們同去，你為甚麼這樣待我們呢？」他們就和 基甸 激烈地爭吵。
JUDG|8|2|基甸 對他們說：「我現在所做的怎麼與你們所做的相比呢？ 以法蓮 拾取剩下的葡萄不強過 亞比以謝 族所摘的葡萄嗎？
JUDG|8|3|上帝已把 米甸 的兩個領袖 俄立 和 西伊伯 交在你們手中；我所做的怎能與你們所做的相比呢？」 基甸 說了這話，他們對他的怒氣就消了。
JUDG|8|4|基甸 和跟隨他的三百人來到 約旦河 ，渡了過去；他們雖然疲乏，還是追趕。
JUDG|8|5|基甸 對 疏割 人說：「請你們拿幾塊餅來給跟隨我的百姓，因為他們疲乏了。我正在追擊 米甸 王 西巴 和 撒慕拿 。」
JUDG|8|6|疏割 人的領袖回答說：「 西巴 和 撒慕拿 的手掌現在已經在你手裏，因此我們該將餅送給你的軍隊嗎？」
JUDG|8|7|基甸 說：「好吧！耶和華將 西巴 和 撒慕拿 交在我手之後，我必用曠野的荊棘和枳條鞭打你們。」
JUDG|8|8|基甸 從那裏上到 毗努伊勒 ，對那裏的人也提出同樣的請求； 毗努伊勒 人給他的答覆跟 疏割 人的答覆一樣。
JUDG|8|9|他也對 毗努伊勒 人說：「我平平安安回來的時候，必拆毀這城樓。」
JUDG|8|10|那時 西巴 和 撒慕拿 ，以及跟隨他們的軍隊都在 加各 ，約有一萬五千人，是東邊的人全軍所剩下的，因為拿刀戰死的約有十二萬人。
JUDG|8|11|基甸 從 挪巴 和 約比哈 的東邊，從住帳棚人 的路上去，趁 米甸 的軍兵以為安全的時候攻擊他們。
JUDG|8|12|西巴 和 撒慕拿 逃跑； 基甸 追趕他們，捉住 米甸 的兩個王 西巴 和 撒慕拿 ，使他們全軍潰散。
JUDG|8|13|約阿施 的兒子 基甸 從戰場，沿著 希列斯 斜坡回來，
JUDG|8|14|捉住 疏割 人的一個少年，查問他。他就為 基甸 寫下 疏割 的領袖和長老的名字，共七十七人。
JUDG|8|15|基甸 到了 疏割 人那裏，說：「你們從前譏笑我說：『 西巴 和 撒慕拿 的手掌現在已經在你手裏，因此我們該將餅送給跟隨你的疲乏的人嗎？』看哪， 西巴 和 撒慕拿 在這裏。」
JUDG|8|16|於是他拿住城內的長老，用曠野的荊棘和枳條責打 疏割 人。
JUDG|8|17|他又拆了 毗努伊勒 的城樓，殺了城裏的人。
JUDG|8|18|基甸 對 西巴 和 撒慕拿 說：「你們在 他泊山 所殺的人是甚麼樣子的？」他們說：「他們很像你，個個都有王子的樣子。」
JUDG|8|19|基甸 說：「他們都是我的兄弟，我母親的兒子。我指著永生的耶和華起誓，你們若存留他們的性命，我就不殺你們了。」
JUDG|8|20|他對他的長子 益帖 說：「你起來殺他們！」但是這少年害怕，不敢拔刀，因為他還是個少年。
JUDG|8|21|西巴 和 撒慕拿 說：「你自己起來殺我們吧！因為人如何，力量也如何。」 基甸 就起來，殺了 西巴 和 撒慕拿 ，取了他們駱駝頸項上的月牙圈。
JUDG|8|22|以色列 人對 基甸 說：「你既然救我們脫離 米甸 的手，願你治理我們，你的兒子孫子也治理我們。」
JUDG|8|23|基甸 對他們說：「我不治理你們，我的兒子也不治理你們，耶和華會治理你們。」
JUDG|8|24|基甸 又對他們說：「我有一件事求你們，請你們各人把所奪的耳環給我。」因敵人都戴金耳環，他們是 以實瑪利 人。
JUDG|8|25|以色列 人說：「我們情願送給你！」他們就鋪開一件外衣，各人將所奪的耳環丟在上面。
JUDG|8|26|基甸 所要求的金耳環，重一千七百舍客勒金子。此外還有 米甸 王所戴的月牙圈、耳環，和所穿的紫色衣服，以及駱駝頸項上的鏈子。
JUDG|8|27|基甸 以此造了一個以弗得，設立在他的本城 俄弗拉 。全 以色列 就在那裏拜這以弗得行淫，這就成了 基甸 和他全家的圈套。
JUDG|8|28|這樣， 米甸 就被 以色列 人制伏了，再也不能抬頭。 基甸 還在的日子，這地太平四十年。
JUDG|8|29|約阿施 的兒子 耶路巴力 回去，住在自己家裏。
JUDG|8|30|基甸 有七十個親生的兒子，因為他有許多妻子。
JUDG|8|31|他在 示劍 的妾也為他生了一個兒子， 基甸 給他起名叫 亞比米勒 。
JUDG|8|32|約阿施 的兒子 基甸 年紀老邁而死，葬在 亞比以謝 族的 俄弗拉 ，他父親 約阿施 的墳墓裏。
JUDG|8|33|基甸 死後， 以色列 人又去隨從諸 巴力 而行淫，以 巴力‧比利土 為他們的神明。
JUDG|8|34|以色列 人不記得耶和華－他們的上帝，就是那位拯救他們脫離四圍仇敵之手的，
JUDG|8|35|也不照著 耶路巴力 ，就是 基甸 向 以色列 所施的恩惠善待他的家。
JUDG|9|1|耶路巴力 的兒子 亞比米勒 到 示劍 他的母舅那裏，對他們和他外祖父全家的人說：
JUDG|9|2|「請你們問 示劍 所有的居民：『是 耶路巴力 的眾兒子七十人都治理你們好，還是一人治理你們好呢？』你們要記得，我是你們的骨肉。」
JUDG|9|3|他的母舅們為他把這一切話說給 示劍 所有的居民聽，他們的心就傾向 亞比米勒 ，因為他們說：「他是我們的弟兄。」
JUDG|9|4|他們從 巴力‧比利土 的廟中取了七十銀子給 亞比米勒 ， 亞比米勒 用這些錢雇了一些無賴匪徒跟隨他。
JUDG|9|5|他來到 俄弗拉 他父親的家，在一塊磐石上把他的兄弟，就是 耶路巴力 的七十個兒子都殺了，只剩下 耶路巴力 的小兒子 約坦 ，因為他躲了起來。
JUDG|9|6|示劍 所有的居民和全 伯‧米羅 都聚集在一起，到 示劍 橡樹旁的柱子那裏，立 亞比米勒 為王。
JUDG|9|7|有人將這事告訴 約坦 ，他就去站在 基利心山 頂上，高聲喊叫，對他們說：「 示劍 的居民哪，你們要聽我，上帝也就會聽你們。
JUDG|9|8|有一次，樹木要膏一王治理他們，就去對橄欖樹說：『請你來作王治理我們！』
JUDG|9|9|橄欖樹對它們說：『我豈可停止生產使神明和人得尊榮的油，而行走飄搖在眾樹之上呢？』
JUDG|9|10|樹木對無花果樹說：『請你來作王治理我們！』
JUDG|9|11|無花果樹對它們說：『我豈可停止結甜美的果子，而行走飄搖在眾樹之上呢？』
JUDG|9|12|樹木對葡萄樹說：『請你來作王治理我們！』
JUDG|9|13|葡萄樹對它們說：『我豈可停止出產使神明和人歡樂的新酒，而行走飄搖在眾樹之上呢。』
JUDG|9|14|眾樹對荊棘說：『請你來作王治理我們！』
JUDG|9|15|荊棘對眾樹說：『你們若真的要膏我作王治理你們，就要來到我的蔭下尋求庇護；不然，願火從荊棘裏出來，吞滅 黎巴嫩 的香柏樹。』
JUDG|9|16|「現在你們若以誠實正直立 亞比米勒 為王，若善待 耶路巴力 和他的家，若照他手所做的回報他─
JUDG|9|17|從前我父為你們爭戰，冒生命的危險救你們脫離 米甸 的手，
JUDG|9|18|但是你們如今起來攻擊我的父家，在一塊磐石上把他的七十個兒子全殺了，又立他使女所生的兒子 亞比米勒 為 示劍 居民的王，因為他是你們的弟兄─
JUDG|9|19|你們如今若以誠實正直對待 耶路巴力 和他的家，就可以因 亞比米勒 歡樂，他也可以因你們歡樂；
JUDG|9|20|不然，願火從 亞比米勒 發出，吞滅 示劍 居民和 伯‧米羅 ，又願火從 示劍 居民和 伯‧米羅 發出，吞滅 亞比米勒 。」
JUDG|9|21|約坦 因躲避他的兄弟 亞比米勒 就逃跑，去到 比珥 ，住在那裏。
JUDG|9|22|亞比米勒 治理 以色列 三年。
JUDG|9|23|上帝派邪靈到 亞比米勒 和 示劍 居民中間， 示劍 居民就以詭詐待 亞比米勒 。
JUDG|9|24|這是要使 耶路巴力 七十個兒子受害所流的血，歸於他們的兄弟 亞比米勒 ，因他殺害他們，也歸於那些出手幫助他殺害兄弟的 示劍 居民。
JUDG|9|25|示劍 居民在山頂上設下埋伏，等候 亞比米勒 。凡沿著那條路，從他們那裏經過的人，他們就搶劫。有人把這事告訴 亞比米勒 。
JUDG|9|26|以別 的兒子 迦勒 和他的弟兄經過，來到 示劍 ， 示劍 居民都信任他。
JUDG|9|27|他們出到田間，摘下葡萄，踹酒，作樂。他們進入他們神明的廟中吃喝，詛咒 亞比米勒 。
JUDG|9|28|以別 的兒子 迦勒 說：「 亞比米勒 是誰，我們 示劍 人是誰，叫我們服事他呢？他不是 耶路巴力 的兒子嗎？他的助手不是 西布勒 嗎？你們應當服事 示劍 的父親 哈抹 的後裔！我們為何要服事 亞比米勒 呢？
JUDG|9|29|惟願這民歸到我的手下，我就除掉 亞比米勒 。」他就對 亞比米勒 說：「增加你的軍兵，出來吧！」
JUDG|9|30|西布勒 市長聽見 以別 的兒子 迦勒 的話，就怒氣大發。
JUDG|9|31|他悄悄地派一些使者到 亞比米勒 那裏，說：「看哪， 以別 的兒子 迦勒 和他的弟兄到了 示劍 。看哪，他們煽動那城攻擊你。
JUDG|9|32|現在，你和跟隨你的百姓要夜間起來，在田間埋伏。
JUDG|9|33|早晨太陽一出，你就趁早攻城。看哪， 迦勒 和跟隨他的百姓出來攻擊你的時候，你就全力對付他們。」
JUDG|9|34|於是， 亞比米勒 和跟隨他的眾百姓夜間起來，兵分四隊，埋伏攻擊 示劍 。
JUDG|9|35|以別 的兒子 迦勒 出去，站在城門口。 亞比米勒 和跟隨他的百姓從埋伏之處起來。
JUDG|9|36|迦勒 看見百姓，就對 西布勒 說：「看哪，有百姓從山頂上下來。」 西布勒 對他說：「你把山的影子看作是人了。」
JUDG|9|37|迦勒 又繼續講，他說：「看哪，有百姓從地的高處下來，又有一隊從 米惡尼尼 橡樹 的路前來。」
JUDG|9|38|西布勒 對他說：「你所誇口的在哪裏呢？你曾說：『 亞比米勒 是誰，叫我們服事他呢？』這不是你所藐視的百姓嗎？你現在出去，與他們交戰吧！」
JUDG|9|39|於是 迦勒 率領 示劍 居民出去，與 亞比米勒 交戰。
JUDG|9|40|亞比米勒 追趕 迦勒 ， 迦勒 在他面前逃跑。有許多人被刺傷仆倒，直到城門口。
JUDG|9|41|亞比米勒 住在 亞魯瑪 。 西布勒 趕出 迦勒 和他的弟兄，不准他們住在 示劍 。
JUDG|9|42|次日，百姓出到田間，有人告訴 亞比米勒 ，
JUDG|9|43|他就帶領百姓，把他們分成三隊，埋伏在田間窺探。看哪， 示劍 居民從城裏出來，他就起來擊殺他們。
JUDG|9|44|亞比米勒 和跟隨他的一隊向前衝，站在城門口；另外兩隊直衝向田間，擊殺了眾人。
JUDG|9|45|亞比米勒 攻城一整天，將城奪取，殺了其中的百姓，把城拆毀，撒上了鹽。
JUDG|9|46|示劍 城樓裏所有的居民聽見了，就進入 伊勒‧比利土 廟的地窖裏。
JUDG|9|47|有人告訴 亞比米勒 ， 示劍 城樓裏所有的居民都聚在一起。
JUDG|9|48|亞比米勒 和所有跟隨他的百姓都上 撒們山 去。 亞比米勒 手拿斧子，砍下一根樹枝，舉起來，扛在肩上，對跟隨他的百姓說：「你們看我做甚麼，就趕快照樣做。」
JUDG|9|49|眾百姓也都各砍一根樹枝，跟 亞比米勒 走，把樹枝堆在地窖上，放火燒地窖。這樣， 示劍 城樓裏所有的人都死了，男女約有一千。
JUDG|9|50|亞比米勒 到 提備斯 ，對著 提備斯 安營，攻取了那城。
JUDG|9|51|城中有一座堅固的樓；城裏所有的居民，無論男女，都逃到那裏，關上門，上了樓頂。
JUDG|9|52|亞比米勒 到了樓前，攻打它。他挨近樓門，要放火焚燒。
JUDG|9|53|有一個婦人把一塊上磨石拋在 亞比米勒 的頭上，打破了他的頭蓋骨。
JUDG|9|54|他就急忙叫拿他兵器的青年來，對他說：「拔出你的刀來，殺了我吧！免得有人提到我說：『他被一個婦人殺了。』」於是那青年把他刺透，他就死了。
JUDG|9|55|以色列 人見 亞比米勒 死了，就各回自己的地方去了。
JUDG|9|56|這樣，上帝報應了 亞比米勒 向他父親所做的惡事，就是殺了自己七十個兄弟。
JUDG|9|57|示劍 人的一切惡事，上帝也都報應在他們頭上； 耶路巴力 的兒子 約坦 的詛咒都臨到他們身上了。
JUDG|10|1|亞比米勒 以後， 陀拉 興起，拯救 以色列 ，他是 朵多 的孫子， 普瓦 的兒子， 以薩迦 人，住在 以法蓮 山區的 沙密 。
JUDG|10|2|陀拉 作 以色列 的士師二十三年。他死了，葬在 沙密 。
JUDG|10|3|陀拉 以後有 基列 人 睚珥 興起，作 以色列 的士師二十二年。
JUDG|10|4|他有三十個兒子，騎著三十匹驢駒。他們有三十座城，叫作 哈倭特‧睚珥 ，直到如今，都在 基列 地。
JUDG|10|5|睚珥 死了，葬在 加們 。
JUDG|10|6|以色列 人又行耶和華眼中看為惡的事，去事奉諸 巴力 和 亞斯她錄 ，以及 亞蘭 的神明、 西頓 的神明、 摩押 的神明、 亞捫 人的神明、 非利士 人的神明。他們離棄耶和華，不事奉他。
JUDG|10|7|耶和華的怒氣向 以色列 發作，把他們交給 非利士 人和 亞捫 人的手中。
JUDG|10|8|從那年起，他們欺壓迫害 以色列 人，在 約旦河 東， 亞摩利 人境內， 基列 一帶所有的 以色列 人，長達十八年。
JUDG|10|9|亞捫 人渡過 約旦河 去攻打 猶大 和 便雅憫 ，以及 以法蓮 家族。 以色列 的處境非常困苦。
JUDG|10|10|以色列 人哀求耶和華說：「我們得罪了你，因為我們離棄了我們的上帝，去事奉諸 巴力 。」
JUDG|10|11|耶和華對 以色列 人說：「我豈沒有救你們脫離 埃及 人、 亞摩利 人、 亞捫 人和 非利士 人嗎？
JUDG|10|12|西頓 人、 亞瑪力 人和 馬雲 人 欺壓你們，你們哀求我，我也拯救你們脫離他們的手。
JUDG|10|13|你們竟離棄我去事奉別神！所以我不再救你們了。
JUDG|10|14|你們去哀求你們所選擇的神明；你們遭遇急難的時候，讓它們救你們吧！」
JUDG|10|15|以色列 人對耶和華說：「我們犯罪了，照你看為好的待我們，只求你今日拯救我們吧！」
JUDG|10|16|以色列 人就除掉他們中間的外邦神明，事奉耶和華。耶和華因 以色列 所受的苦難而心裏焦急。
JUDG|10|17|亞捫 人被召來，在 基列 安營； 以色列 人也聚集，在 米斯巴 安營。
JUDG|10|18|基列 百姓中的領袖彼此說：「誰領先出去攻打 亞捫 人，誰就作 基列 所有居民的領袖。」
JUDG|11|1|基列 人 耶弗他 是個大能的勇士，是妓女的兒子。 基列 生了 耶弗他 。
JUDG|11|2|基列 的妻子也給他生了幾個兒子。他妻子生的兒子長大後，就把 耶弗他 趕出去，說：「你不可在我們父家繼承產業，因為你是別的女人生的兒子。」
JUDG|11|3|耶弗他 就逃離他的兄弟，住在 陀伯 地。有些無賴的人聚集在他那裏，與他一同出入。
JUDG|11|4|過了些日子， 亞捫 人攻打 以色列 。
JUDG|11|5|亞捫 人攻打 以色列 的時候， 基列 的長老去請 耶弗他 從 陀伯 地回來。
JUDG|11|6|他們對 耶弗他 說：「請你來作我們的指揮官，好讓我們跟 亞捫 人打仗。」
JUDG|11|7|耶弗他 對 基列 的長老說：「你們不是恨我，把我趕出父家嗎？現在你們遭遇急難，為何到我這裏來呢？」
JUDG|11|8|基列 的長老對 耶弗他 說：「現在我們回到你這裏，是要請你同我們去跟 亞捫 人打仗，作 基列 所有居民的領袖。」
JUDG|11|9|耶弗他 對 基列 的長老說：「若你們請我回去跟 亞捫 人打仗，耶和華把他們交給我，我就作你們的領袖。」
JUDG|11|10|基列 的長老對 耶弗他 說：「有耶和華在你我之間作證，我們必定照你的話做。」
JUDG|11|11|於是 耶弗他 與 基列 的長老同去，百姓就立 耶弗他 作他們的領袖和指揮官。 耶弗他 在 米斯巴 將他一切的事陳述在耶和華面前。
JUDG|11|12|耶弗他 派使者到 亞捫 人的王那裏，說：「你與我有甚麼相干，竟來到我這裏攻打我的地呢？」
JUDG|11|13|亞捫 人的王對 耶弗他 的使者說：「因為 以色列 從 埃及 上來的時候佔據我的地，從 亞嫩河 到 雅博河 ，直到 約旦河 。現在你要和平歸還這些地方！」
JUDG|11|14|耶弗他 又派使者到 亞捫 人的王那裏，
JUDG|11|15|對他說：「 耶弗他 如此說： 以色列 並沒有佔據 摩押 地和 亞捫 人的地。
JUDG|11|16|以色列 人從 埃及 上來，是經過曠野到 紅海 ，來到 加低斯 。
JUDG|11|17|那時， 以色列 派使者去 以東 王那裏，說：『求你讓我穿越你的地。』 以東 王卻不聽。 以色列 又照樣派使者去 摩押 王那裏，他也不肯。於是 以色列 人就住在 加低斯 。
JUDG|11|18|他們又經過曠野，繞過 以東 地和 摩押 地，到 摩押 地的東邊 ，在 亞嫩河 邊安營，並沒有進入 摩押 的境內，因為 亞嫩河 是 摩押 的邊界。
JUDG|11|19|以色列 派使者去 亞摩利 王，就是 希實本 王 西宏 那裏； 以色列 對他說：『求你讓我們穿越你的地，到我自己的地方去。』
JUDG|11|20|西宏 卻不信任 以色列 ，不讓他們穿越他的疆界。他召集了他的眾百姓在 雅雜 安營，與 以色列 爭戰。
JUDG|11|21|耶和華－ 以色列 的上帝將 西宏 和他的眾百姓都交在 以色列 手中， 以色列 人就擊殺他們，佔領了那地居民 亞摩利 人的全地。
JUDG|11|22|他們佔領了 亞摩利 人所有的疆土，從 亞嫩河 到 雅博河 ，從曠野直到 約旦河 。
JUDG|11|23|耶和華－ 以色列 的上帝如今從他百姓 以色列 面前趕出 亞摩利 人，你竟要佔領它嗎？
JUDG|11|24|你不是已經得了你的神明 基抹 賜給你的地為業嗎？耶和華－我們的上帝在我們面前所趕出的，我們也要得它為業。
JUDG|11|25|現在你比 西撥 的兒子 摩押 王 巴勒 還強嗎？他真的曾與 以色列 爭執，或是真的與他們爭戰了嗎？
JUDG|11|26|以色列 人住 希實本 和所屬的鄉鎮， 亞羅珥 和所屬的鄉鎮，以及沿著 亞嫩河 的一切城鎮，已經有三百年了。在這期間，你們為甚麼不取回呢？
JUDG|11|27|我並沒有得罪你，你卻要攻打我，加害於我。願審判人的耶和華今日在 以色列 人和 亞捫 人之間判斷是非。」
JUDG|11|28|但 亞捫 人的王不聽 耶弗他 傳達給他的話。
JUDG|11|29|耶和華的靈降在 耶弗他 身上，他就經過 基列 和 瑪拿西 ，經過 基列 的 米斯巴 ，又從 基列 的 米斯巴 過到 亞捫 人那裏。
JUDG|11|30|耶弗他 向耶和華許願，說：「你若真的將 亞捫 人交在我手中，
JUDG|11|31|我從 亞捫 人那裏平平安安回來的時候，無論誰先從我家門出來迎接我，就要歸給耶和華，我必將他獻上作為燔祭。」
JUDG|11|32|於是 耶弗他 往 亞捫 人那裏去，與他們爭戰。耶和華將他們交在他手中，
JUDG|11|33|他就徹底擊敗他們，從 亞羅珥 到 米匿 ，直到 亞備勒‧基拉明 ，攻取了二十座城。這樣， 亞捫 人就在 以色列 人面前被制伏了。
JUDG|11|34|耶弗他 回 米斯巴 去，到了自己的家，看哪，他女兒拿著手鼓跳舞出來迎接他。她是 耶弗他 的獨生女，除她以外，沒有別的兒女。
JUDG|11|35|耶弗他一看見她，就撕裂衣服，說：「哀哉！我的女兒啊，你使我非常悲痛，叫我十分為難了。因為我已經向耶和華開了口，不能收回。」
JUDG|11|36|他女兒對他說：「我的父親啊，你既向耶和華開了口，就當照你口中所說的向我行，因為耶和華已經在你的仇敵 亞捫 人身上為你報了仇。」
JUDG|11|37|她又對父親說：「我只求你這一件事，給我兩個月，讓我和同伴下到山裏，好為我的童貞哀哭。」
JUDG|11|38|耶弗他 說：「你去吧！」他就讓她離開兩個月。她和同伴去了，在山裏為她的童貞哀哭。
JUDG|11|39|過了兩個月，她回到父親那裏，父親就照所許的願向她行了。她從來沒有親近男人。於是 以色列 中有個風俗，
JUDG|11|40|每年按著日期 以色列 的女子要去為 基列 人 耶弗他 的女兒哀哭四天。
JUDG|12|1|以法蓮 人被召來，渡河來到 撒分 。他們對 耶弗他 說：「你去與 亞捫 人爭戰，為甚麼沒有召我們同去呢？我們必用火將你和你的家燒了。」
JUDG|12|2|耶弗他 對他們說：「我和我的百姓與 亞捫 人有極大的衝突；我曾召你們來，你們卻沒有來救我脫離他們的手。
JUDG|12|3|我見你們不來救我，就拚了命前去攻打 亞捫 人，耶和華就將他們交在我手中。你們今日為甚麼上我這裏來攻打我呢？」
JUDG|12|4|於是 耶弗他 召集 基列 所有的人，要與 以法蓮 人爭戰。 基列 人擊殺 以法蓮 人，因 以法蓮 人曾說：「你們 基列 人在 以法蓮 和 瑪拿西 中，不過是 以法蓮 逃亡的人而已。」
JUDG|12|5|基列 人把守 約旦河 的渡口，不許 以法蓮 人過去。逃跑的 以法蓮 人若說：「讓我過河。」 基列 人就問他說：「你是不是 以法蓮 人？」他若說：「不是」，
JUDG|12|6|基列 人就對他說：「你說『示播列』。」 以法蓮 人因為發音不準，就會說成「西播列」。 基列 人就捉住他，在 約旦河 的渡口把他殺了。那時， 以法蓮 人被殺的有四萬二千人。
JUDG|12|7|耶弗他 作 以色列 的士師六年。 基列 人 耶弗他 死了，葬在 基列 的城裏 。
JUDG|12|8|耶弗他 以後，有 伯利恆 人 以比讚 作 以色列 的士師。
JUDG|12|9|他有三十個兒子。他把三十個女兒都嫁出去了，也為他的兒子從外面娶了三十個媳婦。他作 以色列 的士師七年。
JUDG|12|10|以比讚 死了，葬在 伯利恆 。
JUDG|12|11|以比讚 以後，有 西布倫 人 以倫 作 以色列 的士師，他作 以色列 的士師十年。
JUDG|12|12|西布倫 人 以倫 死了，葬在 西布倫 地的 亞雅崙 。
JUDG|12|13|以倫 以後，有 比拉頓 人 希列 的兒子 押頓 作 以色列 的士師。
JUDG|12|14|他有四十個兒子，三十個孫子，騎著七十匹驢駒。 押頓 作 以色列 的士師八年。
JUDG|12|15|比拉頓 人 希列 的兒子 押頓 死了，葬在 以法蓮 地的 比拉頓 ，就在 亞瑪力 人的山區。
JUDG|13|1|以色列 人又行耶和華眼中看為惡的事，耶和華將他們交在 非利士 人手中四十年。
JUDG|13|2|那時，有一個 但 支派的 瑣拉 人，名叫 瑪挪亞 。他的妻子不懷孕，不生育。
JUDG|13|3|耶和華的使者向那婦人顯現，對她說：「看哪，以前你不懷孕，不生育，如今你必懷孕生一個兒子。
JUDG|13|4|現在你要謹慎，清酒烈酒都不可喝，任何不潔之物都不可吃，
JUDG|13|5|看哪，你必懷孕，生一個兒子。不可用剃刀剃他的頭，因為這孩子一出母胎就歸給上帝作拿細耳人。他必開始拯救 以色列 脫離 非利士 人的手。」
JUDG|13|6|那婦人來對丈夫說：「有一個神人到我這裏來，他的容貌如上帝使者的容貌，非常可畏。我沒有問他從哪裏來，他也沒有把他的名字告訴我。
JUDG|13|7|他對我說：『看哪，你要懷孕，生一個兒子 。現在，清酒烈酒都不可喝，任何不潔之物都不可吃，因為這孩子從出母胎一直到死的那一天，要歸給上帝作拿細耳人。』」
JUDG|13|8|瑪挪亞 祈求耶和華說：「主啊，求你再差遣那神人到我們這裏來，指示我們對這將要生的孩子該怎樣作。」
JUDG|13|9|上帝垂聽了 瑪挪亞 的聲音。那婦人坐在田間的時候，上帝的使者又到她那裏，但是她的丈夫 瑪挪亞 沒有同她在一起。
JUDG|13|10|婦人急忙跑去告訴丈夫，對他說：「看哪，那日到我這裏來的人又向我顯現了。」
JUDG|13|11|瑪挪亞 起來，跟隨他的妻子來到那人那裏，對他說：「你就是跟這婦人說話的那個人嗎？」他說：「是我。」
JUDG|13|12|瑪挪亞 說：「現在，願你的話應驗！這孩子該如何管教呢？他當做甚麼呢？」
JUDG|13|13|耶和華的使者對 瑪挪亞 說：「我告訴這婦人的一切事，她都要遵守。
JUDG|13|14|葡萄樹所結的不可吃，清酒烈酒都不可喝，任何不潔之物也不可吃。凡我所吩咐的，她都當遵守。」
JUDG|13|15|瑪挪亞 對耶和華的使者說：「請容許我們留你下來，好為你預備一隻小山羊。」
JUDG|13|16|耶和華的使者對 瑪挪亞 說：「你雖然留我，我卻不吃你的食物。你若預備燔祭，就當獻給耶和華。」因 瑪挪亞 不知道他是耶和華的使者。
JUDG|13|17|瑪挪亞 對耶和華的使者說：「請問大名？好讓我們在你的話應驗的時候尊敬你。」
JUDG|13|18|耶和華的使者對他說：「你何必問我的名字呢？我的名字是奇妙的。」
JUDG|13|19|瑪挪亞 取一隻小山羊和素祭，在磐石上獻給耶和華。他行奇妙的事， 瑪挪亞 和他的妻子觀看，
JUDG|13|20|火焰從壇上往上升，耶和華的使者也在壇上的火焰中升上去了。 瑪挪亞 和他的妻子看見，就臉伏於地。
JUDG|13|21|耶和華的使者不再向 瑪挪亞 和他的妻子顯現了。那時， 瑪挪亞 才知道他是耶和華的使者。
JUDG|13|22|瑪挪亞 對他的妻子說：「我們一定會死，因為我們看見了上帝。」
JUDG|13|23|他的妻子卻對他說：「耶和華若有意要我們死，就不會從我們手中接受燔祭和素祭，不會將這一切事指示我們，這時也不會讓我們聽到這話。」
JUDG|13|24|後來婦人生了一個兒子，給他起名叫 參孫 。孩子漸漸長大，耶和華賜福給他。
JUDG|13|25|在 瑣拉 和 以實陶 之間的 瑪哈尼‧但 ，耶和華的靈開始感動 參孫 。
JUDG|14|1|參孫 下到 亭拿 ，在 亭拿 看見一個女子，是 非利士 人的女兒。
JUDG|14|2|他上來告訴他父母說：「我在 亭拿 看見一個女子，是 非利士 人的女兒，現在請你們給我娶她為妻。」
JUDG|14|3|他父母對他說：「在你弟兄的女兒中，或在本族所有的人中，難道沒有女子嗎？你何必在未受割禮的 非利士 人中去娶妻呢？」 參孫 對他父親說：「請你給我娶那女子，因為我喜歡她。」
JUDG|14|4|他的父母並不知道這事是出於耶和華，因為他在找機會攻擊 非利士 人。那時， 非利士 人轄制 以色列 人。
JUDG|14|5|參孫 跟他父母下 亭拿 去，他們到了 亭拿 的葡萄園。看哪，有一隻少壯獅子對著他吼叫。
JUDG|14|6|耶和華的靈大大感動 參孫 ，他就手無寸鐵撕裂獅子，如撕裂小山羊一樣。他做這事，並沒有告訴他的父母親。
JUDG|14|7|參孫 下去跟那女子說話，看著就喜歡她。
JUDG|14|8|過了些日子，他回來要娶那女子，繞道去看獅子的殘骸，看哪，有一群蜜蜂在獅子的屍體內，也有蜜在裏面。
JUDG|14|9|他就取了蜜，放在手掌上，邊走邊吃。他到了父母那裏，給他們蜜，他們也吃了。但他沒有告訴他們，這蜜是從獅子的屍體內取來的。
JUDG|14|10|他父親下到女子那裏去。 參孫 在那裏擺設宴席， 因為這是當時年輕人的習俗。
JUDG|14|11|他們看見 參孫 ，就請了三十個人陪伴他。
JUDG|14|12|參孫 對他們說：「我給你們出個謎語，你們若能在七日宴席之內，猜出謎底告訴我，我就給你們三十件細麻內衣和三十套更換的衣服。
JUDG|14|13|但你們若不能告訴我，你們就給我三十件細麻內衣和三十套更換的衣服。」他們對他說：「請把謎語說給我們聽。」
JUDG|14|14|參孫 對他們說： 「吃的從吃者出來； 甜的從強者出來」。 三日之久，他們都猜不出謎語來。
JUDG|14|15|第七日 ，他們對 參孫 的妻子說：「你哄騙你的丈夫，為我們探出謎底來，否則我們就用火燒你和你的父家。你們請我們來，是不是要奪走我們所有的呢？」
JUDG|14|16|參孫 的妻子在丈夫面前哭哭啼啼說：「你只是恨我，並不愛我。你給我本族的人出謎語，卻不把謎底告訴我。」 參孫 對她說：「看哪，連我的父母我都沒有說，我怎麼可以告訴你呢？」
JUDG|14|17|在七日宴席中，她一直在丈夫面前哭哭啼啼。第七日， 參孫 因妻子的催逼就把謎底告訴了她。她把謎底告訴了她本族的人。
JUDG|14|18|第七日日落以前，那城裏的人對 參孫 說： 「有甚麼比蜜還甜呢？ 有甚麼比獅子更強呢？」 參孫 對他們說： 「你們若不用我的母牛犢耕地， 就無法猜出我的謎底來。」
JUDG|14|19|耶和華的靈大大感動 參孫 ，他就下到 亞實基倫 ，擊殺了三十個人，奪了他們身上的衣服，把衣服給了猜出謎語的人。 參孫 怒氣大發，就上他父親的家去了。
JUDG|14|20|參孫 的妻子就歸了 參孫 的一個同伴，就是作過他伴郎的。
JUDG|15|1|過了些日子，在割麥子的時候， 參孫 帶著一隻小山羊去探望他的妻子，說：「我要進內室到我妻子那裏。」他岳父不許他進去。
JUDG|15|2|他岳父說：「我以為你極其恨她，因此我把她給了你的同伴。她妹妹不是比她更美麗嗎？你可以娶來代替她！」
JUDG|15|3|參孫 對他們說：「這一次我若加害 非利士 人，就不算是我的錯了。」
JUDG|15|4|於是 參孫 去捉了三百隻狐狸，把牠們的尾巴一對一對地綁住，再將火把綁在兩條尾巴中間。
JUDG|15|5|他點著火把，把狐狸放進 非利士 人直立的莊稼，把堆積的禾捆和直立的莊稼，葡萄園、橄欖園全都燒了。
JUDG|15|6|非利士 人說：「這事是誰做的呢？」有人說：「是 亭拿 人的女婿 參孫 做的，因為他岳父把他的妻子給了他的同伴。」於是 非利士 人上去，用火燒了女子和她的父親。
JUDG|15|7|參孫 對他們說：「你們既然這麼做，我必向你們報仇才肯罷休。」
JUDG|15|8|參孫 狠狠擊殺他們，把他們連腿帶腰都砍了。過後，他就下去，住在 以坦巖 的石洞裏。
JUDG|15|9|非利士 人上去，安營在 猶大 ，侵犯 利希 。
JUDG|15|10|猶大 人說：「你們為何上來攻擊我們呢？」他們說：「我們上來是要捆綁 參孫 ，照他向我們所做的對待他。」
JUDG|15|11|於是，三千 猶大 人下到 以坦巖 的石洞裏，對 參孫 說：「 非利士 人轄制我們，你不知道嗎？你向我們做的是甚麼事呢？」他說：「他們向我怎樣做，我也要向他們怎樣做。」
JUDG|15|12|猶大 人對他說：「我們下來是要捆綁你，把你交在 非利士 人手中。」 參孫 說：「你們要向我起誓，你們自己不殺害我。」
JUDG|15|13|他們說：「我們絕不殺你，只把你捆綁，交在 非利士 人手中。」於是他們用兩條新繩綁住 參孫 ，把他從 以坦巖 帶上去。
JUDG|15|14|參孫 到了 利希 ， 非利士 人對著他喊叫。耶和華的靈大大感動 參孫 ，他手臂上的繩子就像著火的麻一樣，綁他的繩子從他手上脫落下來。
JUDG|15|15|他找到一塊未乾的驢腮骨，就伸手拾起來，用它殺了一千人。
JUDG|15|16|參孫 說： 「用驢腮骨， 一堆又一堆 ； 用驢腮骨， 我殺了一千人。」
JUDG|15|17|說完這話，就把那腮骨從手裏拋出去。因此，那地叫作 拉末‧利希 。
JUDG|15|18|參孫 非常口渴，就求告耶和華說：「你既藉僕人的手施行這麼大的拯救，現在我要渴死，落在未受割禮的人手中嗎？」
JUDG|15|19|上帝就使 利希 的窪地裂開，從中湧出水來。 參孫 喝了，精神恢復。因此那泉名叫 隱‧哈歌利 ，直到今日它仍在 利希 。
JUDG|15|20|在 非利士 人轄制的時候， 參孫 作 以色列 的士師二十年。
JUDG|16|1|參孫 到了 迦薩 ，在那裏看見一個妓女，就與她親近。
JUDG|16|2|有人告訴 迦薩 人說：「 參孫 到這裏來了！」他們就包圍起來，整夜在城門埋伏等著他。他們整夜靜悄悄地，說：「等到天一亮我們就殺他。」
JUDG|16|3|參孫 睡到半夜，在半夜起來，抓住城門的門扇和兩個門框，把它們和門閂一起拆下來，扛在肩上，抬到 希伯崙 前面的山頂上。
JUDG|16|4|這事以後， 參孫 在 梭烈谷 愛上了一個女子，名叫 大利拉 。
JUDG|16|5|非利士 人的領袖上去，到那女子那裏，對她說：「請你哄騙 參孫 ，探出他為何有這麼大的力氣，以及我們要用甚麼方法才能勝他，將他捆綁制伏。我們就每人給你一千一百塊銀子。」
JUDG|16|6|大利拉 對 參孫 說：「請你告訴我，你為何有這麼大的力氣，要用甚麼方法才能捆綁制伏你。」
JUDG|16|7|參孫 對她說：「若用七條未乾的新繩子捆綁我，我就像平常人一樣軟弱。」
JUDG|16|8|於是 非利士 人的領袖拿了七條未乾的新繩子來，交給她，她就用繩子捆綁 參孫 。
JUDG|16|9|當時，埋伏的人正在她的內室等著。她對 參孫 說：「 參孫 ， 非利士 人來捉你了！」 參孫 就掙斷繩子，繩子如遇到火的麻線斷裂一樣。這樣，人還是不知道他的力量從哪裏來。
JUDG|16|10|大利拉 對 參孫 說：「看哪，你欺騙我，對我說謊。現在請你告訴我，要用甚麼方法才能捆綁你。」
JUDG|16|11|參孫 對她說：「若用未曾用過的新繩子捆綁我，我就像平常人一樣軟弱。」
JUDG|16|12|大利拉 就用新繩子捆綁他，對他說：「 參孫 ， 非利士 人來捉你了！」當時，埋伏的人在內室等著。 參孫 掙斷手臂上的繩子，如掙斷一條線一樣。
JUDG|16|13|大利拉 對 參孫 說：「你到現在還是欺騙我，對我說謊。請你告訴我，要用甚麼方法才能捆綁你。」 參孫 對她說：「只要用織布的線將我頭上的七條髮綹編織起來就可以了」。
JUDG|16|14|於是 大利拉 用梭子將他的髮綹釘住，對他說：「 參孫 ， 非利士 人來捉你了！」 參孫 從睡中醒來，將織布機上的梭子和織布的線一齊都拔出來了。
JUDG|16|15|大利拉 對 參孫 說：「你既不與我同心，怎麼能說『我愛你』呢？你這三次欺騙我，不告訴我，你為甚麼有這麼大的力氣。」
JUDG|16|16|大利拉 天天用話催逼他，糾纏他，他就心裏煩得要死，
JUDG|16|17|終於把心中的一切都告訴她。 參孫 對她說：「從來沒有人用剃刀剃我的頭，因為我一出母胎就歸給上帝作拿細耳人。若有人剃了我的頭髮，我的力氣就會離開我，我就像平常人一樣軟弱。」
JUDG|16|18|大利拉 見他說出了心中的一切，就派人去召 非利士 人的領袖，說：「請再上來一次，因為他已經說出了心中的一切。」於是 非利士 人的領袖手裏拿著銀子，上到她那裏。
JUDG|16|19|大利拉 哄 參孫 睡在她的膝上，叫一個人來剃掉 參孫 頭上的七條髮綹。於是 大利拉 開始制伏 參孫 ，他的力氣就離開他了。
JUDG|16|20|大利拉 說：「 參孫 ， 非利士 人來捉你了！」 參孫 從睡中醒來，說：「我要像前幾次一樣脫身而去。」他卻不知道耶和華已經離開他了。
JUDG|16|21|非利士 人逮住他，挖了他的眼睛，帶他下到 迦薩 ，用銅鏈鎖住他，叫他在監獄裏推磨。
JUDG|16|22|然而他的頭髮被剃以後，又開始長起來了。
JUDG|16|23|非利士 人的領袖聚集，要向他們的神明 大袞 獻大祭，並且慶祝，說：「我們的神明把我們的仇敵 參孫 交在我們手中了。」
JUDG|16|24|眾人看見 參孫 ，就讚美他們的神明說：「我們的神明把那毀壞我們的地、殺害我們許多人的仇敵交在我們手中了。」
JUDG|16|25|他們心裏高興的時候，就說：「叫 參孫 來，逗我們歡樂。」於是他們把 參孫 從監獄裏提出來，在他們面前戲耍。他們叫他站在兩根柱子中間。
JUDG|16|26|參孫 對牽他手的童僕說：「讓我摸摸支撐這廟宇的柱子，我要靠一靠。」
JUDG|16|27|那時廟宇內充滿男女， 非利士 人的眾領袖也都在那裏，屋頂上約有三千男女觀看 參孫 逗他們歡樂。
JUDG|16|28|參孫 求告耶和華說：「主耶和華啊，求你眷念我。上帝啊，就這一次，求你賜給我力量，使我向 非利士 人報那挖我雙眼的仇。」
JUDG|16|29|參孫 抱住中間支撐廟宇的兩根柱子，左手抱一根，右手抱一根。
JUDG|16|30|然後他說：「讓我與 非利士 人一起死吧！」他盡力彎腰，廟宇就倒塌了，壓住領袖和廟宇內的眾人。這樣， 參孫 死的時候所殺的人比活著所殺的還多。
JUDG|16|31|他的兄弟和他父親的全家都下去收他的屍首，抬上去，葬在 瑣拉 和 以實陶 中間、他父親 瑪挪亞 的墳墓裏。 參孫 作 以色列 的士師二十年。
JUDG|17|1|以法蓮 山區有一個人，名叫 米迦 。
JUDG|17|2|他對母親說：「你的一千一百塊銀子被人拿走了，為此你發咒起誓，也說給我聽。看哪，銀子在我這裏，是我拿的。」他母親說：「願我兒蒙耶和華賜福！」
JUDG|17|3|米迦 把這一千一百塊銀子還他母親。他母親說：「我把這銀子分別為聖，親手獻給耶和華，為我兒子造一尊雕刻的像，以及一尊鑄成的像。現在我把銀子交給你。」
JUDG|17|4|米迦 把銀子還他母親，他母親把二百塊銀子交給銀匠，去造一尊雕刻的像，以及一尊鑄成的像，安置在 米迦 的房子裏。
JUDG|17|5|米迦 這個人有了神堂，又造了以弗得和家中的神像，派他的一個兒子作祭司。
JUDG|17|6|那時， 以色列 中沒有王，各人照自己眼中看為對的去做。
JUDG|17|7|猶大 的 伯利恆 有一個年輕人，是 猶大 族的人。他是 利未 人，寄居在那裏。
JUDG|17|8|這人離開 猶大 的 伯利恆城 ，要找一個可住的地方。他來到 以法蓮 山區 米迦 的家，還要往前走。
JUDG|17|9|米迦 對他說：「你從哪裏來？」他說：「我從 猶大 的 伯利恆 來。我是 利未 人，要找一個可住的地方。」
JUDG|17|10|米迦 說：「你就住在我這裏吧！我以你為父為祭司，每年給你十塊銀子和一套衣服，以及生活所需的食物。」 利未 人就來了。
JUDG|17|11|利未 人願意和這人同住；他待這年輕人如自己的兒子一樣。
JUDG|17|12|米迦 授這年輕的 利未 人祭司的職任，他就住在 米迦 的家裏。
JUDG|17|13|米迦 說：「現在我知道耶和華必恩待我，因為我有 利未 人作我的祭司。」
JUDG|18|1|那時， 以色列 中沒有王。 但 支派的人還在覓地居住，因為直到那日，他們還沒有在 以色列 支派中抽籤得地為業。
JUDG|18|2|但 人從 瑣拉 和 以實陶 派本族中的五個勇士，去窺探偵察那地，對他們說：「你們去偵察那地。」他們來到 以法蓮 山區 米迦 的家中，就在那裏住宿。
JUDG|18|3|他們臨近 米迦 的家，聽出那年輕的 利未 人的口音，就繞到那裏，對他說：「誰領你到這裏來？你在這裏做甚麼？你在這裏得了甚麼？」
JUDG|18|4|他對他們說：「 米迦 如此如此待我，他雇用我，我就作了他的祭司。」
JUDG|18|5|他們對他說：「請你求問上帝，使我們知道所走的道路是否通達。」
JUDG|18|6|祭司對他們說：「你們平平安安去吧，你們所行的道路是在耶和華面前的。」
JUDG|18|7|五人就走了，來到 拉億 ，見那裏的人安居，像 西頓 人的生活一樣安寧無慮，那地無人羞辱他們，無人奪取侵略。他們離 西頓 人很遠，與世無爭 。
JUDG|18|8|五人回到 瑣拉 和 以實陶 他們的弟兄那裏。他們的弟兄對他們說：「你們怎麼了？」
JUDG|18|9|他們說：「起來，我們上去攻打他們吧！我們已經窺探了那地，看哪，那地非常好。你們還要待在這裏嗎？不要再遲延了，立刻出發去得那地為業吧！
JUDG|18|10|你們去，必來到安居的百姓和兩邊遼闊的地。上帝已將那地方交在你們手中了；那裏不缺地上的任何東西。」
JUDG|18|11|於是 但 族的六百人，各帶兵器，從 瑣拉 和 以實陶 出發，
JUDG|18|12|上到 猶大 的 基列‧耶琳 ，在那裏安營。因此那地方名叫 瑪哈尼‧但 ，直到今日。看哪，它在 基列‧耶琳 的西邊。
JUDG|18|13|他們從那裏往 以法蓮 山區去，來到 米迦 的家。
JUDG|18|14|先前窺探 拉億 地的五個人對他們的弟兄說：「你們知道嗎？這些屋子裏有以弗得和家中的神像，以及一尊雕刻的像與一尊鑄成的像。現在你們要知道該怎麼做。」
JUDG|18|15|五人轉身，進入 米迦 的家，來到那年輕 利未 人的房間，向他問安。
JUDG|18|16|六百 但 人各帶兵器，站在門口。
JUDG|18|17|那窺探這地的五個人上前去，進入裏面，拿走雕刻的像、以弗得、家中的神像，以及鑄成的像。祭司和帶兵器的六百人一同站在門口。
JUDG|18|18|當五個人進入 米迦 的家，拿走雕刻的像、以弗得、家中的神像，以及鑄成的像，祭司對他們說：「你們做甚麼呢？」
JUDG|18|19|他們對他說：「不要作聲，用手摀口，跟我們去吧！我們必以你為父為祭司。你作一家的祭司好呢？還是作 以色列 一支派一族的祭司好呢？」
JUDG|18|20|祭司心裏歡喜，拿著以弗得和家中的神像，以及雕刻的像，跟這些百姓走了。
JUDG|18|21|他們轉身離開那裏，把孩子、牲畜、財物安排在前頭。
JUDG|18|22|他們離了 米迦 的家已遠， 米迦 家附近的鄰居被召來，追趕 但 人。
JUDG|18|23|他們呼叫 但 人， 但 人回頭對 米迦 說：「你召集這許多人來做甚麼呢？」
JUDG|18|24|米迦 說：「你們把我所造的神像，還有祭司，都帶走了，我還有甚麼呢？你怎麼還對我說『你在做甚麼』呢？」
JUDG|18|25|但 人對 米迦 說：「你不要讓我們再聽見你的聲音，恐怕這群惱怒成性的人會攻擊你們，你和你的全家就會喪命。」
JUDG|18|26|但 人仍走他們的路。 米迦 見他們的勢力比自己強，就轉身回家去了。
JUDG|18|27|但 人把 米迦 造的神像和他的祭司帶走，來到 拉億 安寧無慮的百姓那裏，用刀殺了他們，放火燒了那城。
JUDG|18|28|沒有人來搭救，因為這城離 西頓 很遠，他們又與世無爭；這城在靠近 伯‧利合 的平原。 但 人建造這城，在那裏居住，
JUDG|18|29|並照著他們祖先 以色列 之子 但 的名字，給這城起名叫 但 。原先這城名叫 拉億 。
JUDG|18|30|但 人為自己設立了那雕刻的像。 摩西 的孫子， 革舜 的兒子 約拿單 和他的子孫作 但 支派的祭司，直到那地遭擄掠的日子。
JUDG|18|31|上帝的家在 示羅 多少日子， 但 人為自己設立 米迦 所雕刻的像也在 但 多少日子。
JUDG|19|1|當 以色列 中沒有王的時候，有一個 利未 人寄居 以法蓮 山區的邊界，他娶了一個 猶大伯利恆 的女子為妾。
JUDG|19|2|這妾對丈夫生氣 ，離開丈夫，回到 猶大伯利恆 的父家，在那裏住了四個月。
JUDG|19|3|她的丈夫起來，帶著一個僕人、兩匹驢跟著她去，要用好話勸她回來。女子就帶丈夫進到父親家裏。女子的父親看見了他，就歡歡喜喜地迎接他。
JUDG|19|4|這岳父，就是女子的父親，留他住了三天。他們在那裏吃喝，住宿。
JUDG|19|5|第四日，他們清早起來， 利未 人起身要走，女子的父親對女婿說：「先吃點東西，加添心力，然後你們才走。」
JUDG|19|6|於是二人坐下，一同吃喝。女子的父親對那人說：「請你答應再住一夜，使你的心舒暢。」
JUDG|19|7|那人起身要走，他岳父挽留他，他就留下，在那裏又住了一夜。
JUDG|19|8|第五日，他清早起來要走，女子的父親說：「來，請加添心力，留到太陽偏西吧。」於是二人一同再吃。
JUDG|19|9|那人同他的妾和僕人起身要走，但他岳父，就是女子的父親，對他說：「看哪，太陽下山，天快晚了，你們再住一夜吧。看哪，太陽偏西了，就在這裏住宿，使你的心舒暢，明天你們一早起來上路，回你的帳棚去。」
JUDG|19|10|那人不願再住一夜，就備上兩匹驢，帶著他的妾起身走了，來到 耶布斯 的對面， 耶布斯 就是 耶路撒冷 。
JUDG|19|11|將近 耶布斯 的時候，太陽快下山了，僕人對主人說：「來吧，我們進這 耶布斯 人的城，在這裏住宿。」
JUDG|19|12|主人對他說：「我們不可進入外邦人的城，那不是 以色列 人的地方，我們越過這裏到 基比亞 去吧。」
JUDG|19|13|他又對僕人說：「來，讓我們到 基比亞 或 拉瑪 的一個地方住宿。」
JUDG|19|14|於是他們越過那裏往前走，將到 便雅憫 的 基比亞 的時候，太陽已經下山了。
JUDG|19|15|他們進入 基比亞 要在那裏住宿。他來坐在城裏的廣場上，但沒有人接待他們到家裏住宿。
JUDG|19|16|看哪，晚上有一個老人從田間做工回來。他是 以法蓮 山區的人，寄居在 基比亞 ；那地方的人是 便雅憫 人。
JUDG|19|17|老人舉目看見那過路的人在城裏的廣場上，就說：「你從哪裏來？要到哪裏去？」
JUDG|19|18|他對他說：「我們從 猶大 的 伯利恆 過來，要到 以法蓮 山區的邊界去。我是那裏的人，去了 猶大 的 伯利恆 ，現在要到耶和華的家去，卻沒有人接待我到他的家。
JUDG|19|19|其實我有飼料草料可以餵驢，我和你的使女，以及與我們在一起的僕人都有餅有酒，甚麼都不缺。」
JUDG|19|20|老人說：「願你平安！你所需用的我都會給你們，只是不可在廣場上過夜。」
JUDG|19|21|於是老人領他到家裏，餵上驢。他們洗了腳，就吃喝起來。
JUDG|19|22|他們心裏歡樂的時候，看哪，城中的無賴圍住房子，連連叩門，對老人，這家的主人說：「把那進你家的人帶出來，我們要與他交合。」
JUDG|19|23|這家的主人出來對他們說：「弟兄們，不要做這樣的惡事。這人既然進了我的家，你們就不要做這樣可恥的事。
JUDG|19|24|看哪，我有個女兒還是處女，還有這人的妾，我把她們領出來任由你們污辱她們，就照你們看為好的對待她們吧！但對這人你們不要做這樣可恥的事。」
JUDG|19|25|那些人卻不肯聽從他。那人抓住他的妾，把她拉出去給他們。他們強姦了她，整夜凌辱她，直到早晨，天色快亮才放她走。
JUDG|19|26|到了早晨，婦人回來，仆倒在留她主人住宿的那人的家門前，直到天亮。
JUDG|19|27|早晨，她的主人起來開了門，出去要上路。看哪，那婦人，他的妾倒在屋子門前，雙手搭在門檻上。
JUDG|19|28|他對婦人說：「起來，我們走吧！」婦人卻沒有回應。那人就將她馱在驢上，起身回自己的地方去了。
JUDG|19|29|到了家裏，他拿刀，抓住他的妾，把她的屍身切成十二塊，分送到 以色列 全境。
JUDG|19|30|凡看見的人都說：「自從 以色列 人離開 埃及 地上來，直到今日，像這樣的事還沒有發生過，也沒有見過。大家應當想一想，商討一下再說。」
JUDG|20|1|於是 以色列 眾人從 但 到 別是巴 ，以及從 基列 地出來，如同一人，聚集在 米斯巴 耶和華那裏。
JUDG|20|2|以色列 各支派中眾百姓的領袖，都站在上帝百姓的會中。拿刀的步兵共有四十萬。
JUDG|20|3|便雅憫 人聽見 以色列 人上了 米斯巴 。 以色列 人說：「請說，這惡事是怎麼發生的呢？」
JUDG|20|4|那 利未 人，就是被害婦人的丈夫，回答說：「我和我的妾來到 便雅憫 的 基比亞 住宿。
JUDG|20|5|基比亞 人夜間起來攻擊我，包圍我住的屋子。他們想要殺我，並把我的妾污辱致死。
JUDG|20|6|我把我的妾切成塊，分送到 以色列 得為業的全地，因為 基比亞 人在 以色列 中做了邪惡可恥的事。
JUDG|20|7|看哪，你們大家， 以色列 人哪，在此提出你們的建議和對策吧！」
JUDG|20|8|眾百姓都起來如同一人，說：「我們誰也不回自己的帳棚，誰也不回自己的家去！
JUDG|20|9|現在，我們要這樣對付 基比亞 ，照所抽的籤去攻打他們。
JUDG|20|10|我們要在 以色列 各支派中，一百人選十人，一千人選一百人，一萬人選一千人，為那到 便雅憫 的 迦巴 去的士兵運糧；因為 基比亞 在 以色列 中行了可恥的事。」
JUDG|20|11|於是 以色列 眾人彼此聯合如同一人，聚集攻擊那城。
JUDG|20|12|以色列 眾支派派人去，問 便雅憫 支派的各家說：「你們中間怎麼做了這樣的惡事呢？
JUDG|20|13|現在你們要把 基比亞 的那些無賴交出來，我們好處死他們，從 以色列 中除掉這惡。」 便雅憫 人卻不肯聽從他們弟兄 以色列 人的話。
JUDG|20|14|便雅憫 人從各城聚集到 基比亞 ，出來要與 以色列 人打仗。
JUDG|20|15|那日， 便雅憫 人從各城裏徵召了拿刀的士兵，共有二萬六千，另外還從 基比亞 居民中徵召七百個精兵。
JUDG|20|16|全軍中有特選的七百個精兵，都是慣用左手的，個個能用機弦甩石，毫髮不差。
JUDG|20|17|以色列 人，除了 便雅憫 之外，共徵召了四十萬拿刀的，個個都是戰士。
JUDG|20|18|以色列 人起來，上到 伯特利 去求問上帝說：「我們中間誰當首先上去與 便雅憫 人爭戰呢？」耶和華說：「 猶大 先上去。」
JUDG|20|19|以色列 人早晨起來，對著 基比亞 安營。
JUDG|20|20|以色列 人出來與 便雅憫 人打仗， 以色列 人在 基比亞 對著他們擺陣。
JUDG|20|21|便雅憫 人從 基比亞 出來，當日把 以色列 中二萬二千人殺倒在地。
JUDG|20|22|以色列 人的士兵鼓起勇氣，在第一日擺陣的地方又擺陣。
JUDG|20|23|因 以色列 人上去，在耶和華面前哀哭，直到晚上。他們求問耶和華說：「我可以再出兵與我弟兄 便雅憫 人打仗嗎？」耶和華說：「可以上去攻打他們。」
JUDG|20|24|第二日， 以色列 人就上前攻擊 便雅憫 人。
JUDG|20|25|便雅憫 人也在第二日從 基比亞 出來與他們交戰，又把 以色列 人一萬八千個拿刀的士兵殺倒在地。
JUDG|20|26|以色列 眾人和全體士兵上到 伯特利 ，坐在耶和華面前哭泣。那日，他們禁食直到晚上，又在耶和華面前獻燔祭和平安祭。
JUDG|20|27|以色列 人去求問耶和華；那時，上帝的約櫃在那裏。
JUDG|20|28|那時， 亞倫 的孫子， 以利亞撒 的兒子 非尼哈 侍立在約櫃前。他們說：「我可以再出去與我弟兄 便雅憫 人打仗嗎？還是停戰呢？」耶和華說：「你們可以上去，因為明日我必把他交在你手中。」
JUDG|20|29|以色列 在 基比亞 的四圍設下埋伏。
JUDG|20|30|第三日， 以色列 人又上去攻擊 便雅憫 人，在 基比亞 前擺陣，與前兩次一樣。
JUDG|20|31|便雅憫 人也出來迎敵，就被引誘出城外。在田間的兩條路上，一條通往 伯特利 ，一條通往 基比亞 ，他們像前兩次一樣，動手殺了約三十個 以色列 人。
JUDG|20|32|便雅憫 人說：「他們仍像以前一樣敗在我們面前。」但 以色列 人說：「讓我們逃跑，引誘他們離開城到路上來。」
JUDG|20|33|以色列 眾人都起來，在 巴力‧他瑪 擺陣， 以色列 的伏兵從 馬利‧迦巴 埋伏的地方衝上前去。
JUDG|20|34|全 以色列 中的一萬精兵來到 基比亞 前，戰爭十分激烈。 便雅憫 人卻不知道災禍臨近了。
JUDG|20|35|耶和華在 以色列 面前擊打 便雅憫 。那日， 以色列 人殲滅二萬五千一百個 便雅憫 人，都是拿刀的士兵。
JUDG|20|36|便雅憫 人看到自己戰敗了。 以色列 人因為信任在 基比亞 前所設的伏兵，就在 便雅憫 人面前假裝撤退。
JUDG|20|37|伏兵迅速闖進 基比亞 ；他們繼續前進，用刀殺死全城的人。
JUDG|20|38|以色列 人預先與伏兵約定在城內放火，以上騰的煙為信號。
JUDG|20|39|以色列 人從陣上撤退， 便雅憫 人動手殺死 以色列 人，約有三十個，就說：「他們仍像以前一樣敗在我們面前。」
JUDG|20|40|當煙如柱一般從城中上騰的時候， 便雅憫 人回頭，看哪，全城已經濃煙沖天了。
JUDG|20|41|以色列 人又轉身回來， 便雅憫 人就很驚惶，因為看見災禍臨到自己了。
JUDG|20|42|他們在 以色列 人面前轉身往曠野逃跑，戰況對他們不利，那從城裏出來的也去夾攻，殺滅他們。
JUDG|20|43|以色列 人圍攻 便雅憫 人，追趕他們，在他們歇腳之處，直到向日出方向的 基比亞 的對面，踐踏他們。
JUDG|20|44|便雅憫 人倒下的有一萬八千名，這些全都是勇士。
JUDG|20|45|其餘的人轉身往曠野逃跑，到 臨門巖 去。 以色列 人在路上殺了五千人，如拾穗一樣，緊追他們直到 基頓 ，又殺了二千人。
JUDG|20|46|那日 便雅憫 人倒下的有二萬五千名，這些全都是拿刀的勇士。
JUDG|20|47|有六百人轉身往曠野逃跑，到了 臨門巖 ，在 臨門巖 住了四個月。
JUDG|20|48|以色列 人又轉回去攻擊 便雅憫 人，凡經過的各城，其中的人和牲畜都用刀殺了，又放火燒了所經過的一切城鎮。
JUDG|21|1|以色列 人在 米斯巴 曾起誓說：「我們中誰都不把女兒嫁給 便雅憫 人。」
JUDG|21|2|以色列 人來到 伯特利 ，坐在那裏直到晚上，在上帝面前放聲大哭，
JUDG|21|3|說：「耶和華－ 以色列 的上帝啊，為何 以色列 中會發生這樣的事，使 以色列 今日缺了一個支派呢？」
JUDG|21|4|次日，百姓清早起來，在那裏築了一座壇，獻燔祭和平安祭。
JUDG|21|5|以色列 人說：「 以色列 各支派中，誰沒有同會眾一起上到耶和華那裏呢？」因為 以色列 人曾起重誓說：「凡不上 米斯巴 到耶和華那裏的，必被處死。」
JUDG|21|6|以色列 人憐憫他們的弟兄 便雅憫 ，說：「如今 以色列 中斷絕一個支派了。
JUDG|21|7|我們既然向耶和華起誓說，必不把我們的女兒嫁給 便雅憫 人，現在我們該怎麼辦，使他們剩下的人可以娶妻呢？」
JUDG|21|8|他們又說：「 以色列 支派中誰沒有上 米斯巴 到耶和華那裏呢？」看哪， 基列 的 雅比 沒有一人進營到會眾那裏，
JUDG|21|9|百姓被數點的時候，看哪， 基列 的 雅比 居民沒有一人在那裏。
JUDG|21|10|會眾就派一萬二千名大勇士，吩咐他們說：「你們去用刀把 基列 的 雅比 居民連婦女帶孩子都殺了。
JUDG|21|11|這是你們當做的事：要把所有男人和曾與男人同房共寢的女人全都殺了。」
JUDG|21|12|他們在 基列 的 雅比 居民中，找到四百個未曾與男人同房共寢的處女，就帶她們到 迦南 地的 示羅 營裏。
JUDG|21|13|全會眾派人到 臨門巖 的 便雅憫 人那裏，與他們講和。
JUDG|21|14|當時 便雅憫 人回來了， 以色列 人就把所留下， 基列 的 雅比 活著的女子嫁給他們，可是還是不夠。
JUDG|21|15|百姓憐憫 便雅憫 人，因為耶和華使 以色列 支派中有一個缺口。
JUDG|21|16|會眾中的長老說：「 便雅憫 中的女子既然都除滅了，我們該怎麼辦，使剩下的人可以娶妻呢？」
JUDG|21|17|他們又說：「 便雅憫 逃脫的人應當有地業，免得 以色列 中的一個支派被塗去。
JUDG|21|18|只是我們不能把自己的女兒嫁給他們。」因為 以色列 人曾起誓說：「把女兒嫁給 便雅憫 人的必受詛咒。」
JUDG|21|19|他們又說：「看哪，一年一度耶和華的節期正在 示羅 舉行。」 示羅 位於 利波拿 的南邊， 伯特利 的北邊，從 伯特利 往 示劍 大路的東邊。
JUDG|21|20|他們吩咐 便雅憫 人說：「你們去，躲在葡萄園中，
JUDG|21|21|觀看；看哪，若 示羅 的女子出來跳舞，你們就從葡萄園出來，各人從 示羅 的女子中搶一個為妻，然後到 便雅憫 地去。
JUDG|21|22|他們的父親或兄弟若來與我們爭論，我們就對他們說：『請看我們的情面恩待這些人吧！因為我們在戰爭的時候沒有給他們任何人留下女子為妻。這次也不是你們給他們的，若是你們給的，就算有罪了。』」
JUDG|21|23|於是 便雅憫 人就照樣做了，按照他們的人數，把從跳舞女子中搶來的娶為妻子，帶回自己的地業，重建城鎮，居住在其中。
JUDG|21|24|那時 以色列 人離開那裏，各自回到自己的支派、宗族；他們從那裏起行，各自回到自己的地業去了。
JUDG|21|25|那時， 以色列 中沒有王，各人照自己眼中看為對的去做。
RUTH|1|1|士師統治的時候，國中有饑荒。在 猶大 的 伯利恆 ，有一個人帶著妻子和兩個兒子往 摩押 地去寄居。
RUTH|1|2|這人名叫 以利米勒 ，他的妻子名叫 拿娥米 ；他兩個兒子，一個名叫 瑪倫 ，一個名叫 基連 ，都是 猶大伯利恆 的 以法他 人。他們到了 摩押 地，就住在那裏。
RUTH|1|3|後來 拿娥米 的丈夫 以利米勒 死了，剩下她和兩個兒子。
RUTH|1|4|兩個兒子娶了 摩押 女子，一個名叫 俄珥巴 ，第二個名叫 路得 ，在那裏住了約有十年。
RUTH|1|5|瑪倫 和 基連 二人也死了，剩下 拿娥米 ，沒有丈夫，也沒有兒子。
RUTH|1|6|拿娥米 與兩個媳婦起身，要從 摩押 地回去，因為她在 摩押 地聽見耶和華眷顧自己的百姓，賜糧食給他們。
RUTH|1|7|她和兩個媳婦就起行，離開所住的地方，上路回 猶大 地去。
RUTH|1|8|拿娥米 對兩個媳婦說：「你們各自回娘家去吧！願耶和華恩待你們，像你們待已故的人和我一樣。
RUTH|1|9|願耶和華使你們各自在新的丈夫家中得歸宿！」於是 拿娥米 與她們親吻，她們就放聲大哭，
RUTH|1|10|對她說：「不，我們要與你一同回你的百姓那裏去。」
RUTH|1|11|拿娥米 說：「我的女兒啊，回去吧！為何要跟我去呢？我還能生兒子作你們的丈夫嗎？
RUTH|1|12|我的女兒啊，回去吧！我年紀老了，不能再有丈夫。就算我還有希望，今夜有丈夫，而且也生了兒子，
RUTH|1|13|你們豈能等著他們長大呢？你們能守住自己不嫁人嗎？我的女兒啊，不要這樣。我比你們更苦，因為耶和華伸手擊打我。」
RUTH|1|14|兩個媳婦又放聲大哭， 俄珥巴 與婆婆吻別，但是 路得 卻緊跟著 拿娥米 。
RUTH|1|15|拿娥米 說：「看哪，你嫂嫂已經回她的百姓和她的神明那裏去了，你也跟你嫂嫂回去吧！」
RUTH|1|16|路得 說： 「不要勸我離開你， 轉去不跟隨你。 你往哪裏去， 我也往哪裏去； 你在哪裏住， 我也在哪裏住； 你的百姓就是我的百姓； 你的上帝就是我的上帝。
RUTH|1|17|你死在哪裏， 我也死在哪裏，葬在哪裏。 只有死能使你我分離； 不然，願耶和華重重懲罰我！」
RUTH|1|18|拿娥米 見 路得 決意要跟自己去，就不再對她說甚麼了。
RUTH|1|19|於是二人同行，來到 伯利恆 。她們到了 伯利恆 ，全城因她們騷動起來。婦女們說：「這是 拿娥米 嗎？」
RUTH|1|20|拿娥米 對她們說： 「不要叫我 拿娥米 ， 要叫我 瑪拉 ， 因為全能者使我受盡了苦。
RUTH|1|21|我滿滿地出去， 耶和華使我空空地回來。 耶和華使我受苦， 全能者降禍於我。 你們為何還叫我 拿娥米 呢？」
RUTH|1|22|拿娥米 從 摩押 地回來了，她的媳婦 摩押 女子 路得 跟她在一起。她們到了 伯利恆 ，正是開始收割大麥的時候。
RUTH|2|1|拿娥米 有一個親戚，是她丈夫 以利米勒 本族的人，名叫 波阿斯 ，是個大財主。
RUTH|2|2|摩押 女子 路得 對 拿娥米 說：「讓我到田裏去拾取麥穗，我在誰的眼中蒙恩，就跟在誰的身後。」 拿娥米 說：「女兒啊，你去吧。」
RUTH|2|3|路得 就去了。她來到田間，在收割的人身後拾取麥穗。她恰巧來到 以利米勒 本族的人 波阿斯 那塊田裏。
RUTH|2|4|看哪， 波阿斯 正從 伯利恆 來，對收割的人說：「願耶和華與你們同在！」他們對他說：「願耶和華賜福給你！」
RUTH|2|5|波阿斯 對監督收割的僕人說：「那是誰家的女子？」
RUTH|2|6|監督收割的僕人回答說：「她是 摩押 女子，跟隨 拿娥米 從 摩押 地回來的。
RUTH|2|7|她說：『請你容許我拾取麥穗，在收割的人身後撿禾捆中掉落的麥穗。』她就來了，從早晨直到如今，除了在屋子裏坐一會兒，她都留在這裏。」
RUTH|2|8|波阿斯 對 路得 說：「女兒啊，聽我說，不要到別人田裏去拾取麥穗，也不要離開這裏，要緊跟著我的女僕們。
RUTH|2|9|你要看好我的僕人正在哪塊田收割，就跟著女僕們去。我已經吩咐僕人不可侵犯你。你渴了，可以到水缸那裏喝僕人打來的水。」　
RUTH|2|10|路得 就臉伏於地叩拜，對他說：「我既是外邦女子，怎麼會在你眼中蒙恩，使你這樣照顧我呢？」
RUTH|2|11|波阿斯 回答她說：「自從你丈夫死後，凡你向婆婆所行的，以及你離開父母和你的出生地，到素不相識的百姓中，這些事人都告訴我了。
RUTH|2|12|願耶和華照你所行的報償你。你來投靠在耶和華－ 以色列 上帝的翅膀下，願你滿得他的報償。」
RUTH|2|13|路得 說：「我主啊，願我在你眼前蒙恩。我雖然不及你的一個婢女，你還安慰我，對你的婢女說關心的話。」
RUTH|2|14|吃飯的時候， 波阿斯 對 路得 說：「你到這裏來吃些餅，把你的一塊蘸在醋裏。」 路得 就在收割的人旁邊坐下。 波阿斯 把烘了的穗子遞給她。她吃飽了，還有剩餘的。
RUTH|2|15|她又起來拾取麥穗， 波阿斯 吩咐僕人說：「她即使在禾捆中拾取麥穗，也不可羞辱她。
RUTH|2|16|你們還要從捆裏抽一些出來，留給她拾取，不可責備她。」
RUTH|2|17|這樣， 路得 在田間拾取麥穗，直到晚上。她把所拾取的麥穗打了約有一伊法的大麥。
RUTH|2|18|路得 把所拾取的帶進城去給婆婆看，又把她吃飽所剩的拿出來，給了婆婆。
RUTH|2|19|婆婆問她說：「你今日在哪裏拾取麥穗？在哪裏做工呢？願那照顧你的得福。」 路得 告訴婆婆，她在誰那裏做工，說：「我今日在一個名叫 波阿斯 的人那裏做工。」
RUTH|2|20|拿娥米 對媳婦說：「願那人蒙耶和華賜福，因為他不斷地恩待活人死人。」 拿娥米 又對她說：「那人是我們本族的人，是一個可以贖我們產業的至親。」
RUTH|2|21|摩押 女子 路得 說：「他還對我說：『你要緊跟著我的僕人拾取麥穗，直到他們把我所有的莊稼收割完畢。』」
RUTH|2|22|拿娥米 對媳婦 路得 說：「女兒啊，你要跟著他的女僕出去，免得你在別人的田間受人騷擾。」
RUTH|2|23|於是 路得 緊跟著 波阿斯 的女僕拾取麥穗，直到大麥和小麥收割完畢。 路得 仍與婆婆同住。
RUTH|3|1|路得 的婆婆 拿娥米 對她說：「女兒啊，我不該為你找個歸宿，使你享福嗎？
RUTH|3|2|你與 波阿斯 的女僕常在一處，現在， 波阿斯 不是我們的親人嗎？看哪，他今夜將在禾場簸大麥。
RUTH|3|3|你要沐浴抹膏，穿上外衣，下到禾場，一直到那人吃喝完了，都不要讓他認出你來。
RUTH|3|4|他躺下的時候，你看準他躺臥的地方，就進去掀露他的腳，躺臥在那裏，他必告訴你所當做的事。」
RUTH|3|5|路得 說：「凡你所吩咐我的，我必遵行。」
RUTH|3|6|路得 就下到禾場，照她婆婆吩咐她的一切去做。
RUTH|3|7|波阿斯 吃喝完了，心情暢快，就去躺臥在麥堆旁邊。 路得 悄悄走來，掀露他的腳，躺臥在那裏。
RUTH|3|8|到了半夜，那人驚醒，翻過身來，看哪，有個女子躺在他的腳旁。
RUTH|3|9|他就說：「你是誰？」 路得 說：「我是你的使女 路得 。請你用你衣服的邊來遮蓋你的使女，因為你是可以贖我產業的至親。」
RUTH|3|10|波阿斯 說：「女兒啊，願你蒙耶和華賜福。你後來的忠誠比先前的更美，因為無論貧富的年輕人，你都沒有跟從。
RUTH|3|11|女兒啊，現在不要懼怕，凡你所說的，我必為你做，因為我城裏的百姓都知道你是個賢德的女子。
RUTH|3|12|現在，我的確是一個可以贖你產業的至親，可是還有一個人比我更親。
RUTH|3|13|你今夜在這裏住宿，明早他若肯為你盡至親的本分，很好，就由他吧！倘若他不肯，我指著永生的耶和華起誓，我必為你盡上至親的本分。你只管躺到早晨。」
RUTH|3|14|路得 就在他腳旁躺到早晨，在人還無法彼此辨認的時候就起來了。 波阿斯 說：「不可讓人知道有女子到禾場來。」　
RUTH|3|15|他又對 路得 說：「把你所披的外衣拿來，握緊它。」她就握緊外衣， 波阿斯 量了六簸箕的大麥，幫 路得 扛上，他就進城去了 。」
RUTH|3|16|路得 回到婆婆那裏，婆婆說：「女兒啊，怎麼樣了 ？」 路得 就把那人向她所做的一切都告訴了婆婆，
RUTH|3|17|又說：「那人給了我這六簸箕的大麥，對我說：『你不可空手回去見婆婆。』」
RUTH|3|18|婆婆說：「女兒啊，等著吧，看這事結果如何，因為那人今日不辦妥這事，必不罷休。」
RUTH|4|1|波阿斯 上到城門，坐在那裏，看哪， 波阿斯 所說那個可以贖產業的至親經過。 波阿斯 說：「某某先生，請你轉回來，坐在這裏。」他就轉回來坐下。
RUTH|4|2|波阿斯 又請了本城的十個長老來，對他們說：「請你們坐在這裏。」他們就都坐下。
RUTH|4|3|波阿斯 對那至親說：「從 摩押 地回來的 拿娥米 ，現在要賣我們弟兄 以利米勒 的那塊地。
RUTH|4|4|我想我應該向你說清楚：你可以買那塊地，當著在座的眾人和我百姓的長老面前，你若要贖就贖吧！倘若你不贖 就告訴我，讓我知道，因為除了你以外，沒有人可以先贖，在你之後才輪到我。」那人說：「我要贖。」
RUTH|4|5|波阿斯 說：「你從 拿娥米 和 摩押 女子 路得 手中買這地的時候，也當買死人的妻子，使死人在產業上留名。」
RUTH|4|6|那至親說：「這樣我就不能贖了，免得對我的產業有損。你儘管去贖我所當贖的吧，我不能贖了！」
RUTH|4|7|從前，在 以色列 中要確認任何交易，無論是贖業或買賣，一方必須脫鞋給另一方。 以色列 中都以此為證。
RUTH|4|8|那至親對 波阿斯 說：「你自己買吧！」於是把鞋脫了下來。
RUTH|4|9|波阿斯 對長老和所有在場的百姓說：「你們今日都是證人；凡屬 以利米勒 ，以及 基連 和 瑪倫 的，我都從 拿娥米 手中買下來了。
RUTH|4|10|我也娶 瑪倫 的妻子 摩押 女子 路得 ，好讓死人可以在產業上留名，免得他的名在本族本鄉的城門中消失了。你們今日都是證人。」
RUTH|4|11|在城門坐著的所有百姓和長老說：「我們都是證人。願耶和華使進你家的這女子，像建立 以色列 家的 拉結 和 利亞 二人一樣。又願你在 以法他 得亨通，在 伯利恆 有名聲。
RUTH|4|12|願耶和華從這年輕女子賜你後裔，使你的家像 她瑪 從 猶大 所生 法勒斯 的家一樣。」
RUTH|4|13|於是， 波阿斯 娶了 路得 為妻，與她同房。耶和華使她懷孕生了一個兒子。
RUTH|4|14|婦女們對 拿娥米 說：「耶和華是應當稱頌的！因為他今日沒有使你斷絕可以贖產業的至親。願這孩子在 以色列 中得名聲。
RUTH|4|15|他必振奮你的精神，奉養你的晚年，因為他是愛慕你的媳婦所生的。有這樣的媳婦，比有七個兒子更好！」
RUTH|4|16|拿娥米 接過孩子來，抱在懷中撫養他。
RUTH|4|17|鄰居的婦人給孩子起名，說：「 拿娥米 得了一個孩子了！」她們就給他起名叫 俄備得 。 俄備得 是 耶西 的父親，是 大衛 的祖父。
RUTH|4|18|這是 法勒斯 的後代： 法勒斯 生 希斯崙 ；
RUTH|4|19|希斯崙 生 蘭 ； 蘭 生 亞米拿達 ；
RUTH|4|20|亞米拿達 生 拿順 ； 拿順 生 撒門 ；
RUTH|4|21|撒門 生 波阿斯 ； 波阿斯 生 俄備得 ；
RUTH|4|22|俄備得 生 耶西 ； 耶西 生 大衛 。
1SAM|1|1|以法蓮 山區有一個 拉瑪 的 瑣非 人 ，名叫 以利加拿 ，他是 蘇弗 的玄孫， 託戶 的曾孫， 以利戶 的孫子， 耶羅罕 的兒子，是 以法蓮 人。
1SAM|1|2|他有兩個妻子：一個名叫 哈拿 ，另一個名叫 毗尼拿 。 毗尼拿 有孩子， 哈拿 卻沒有孩子。
1SAM|1|3|這人每年從本城上到 示羅 ，敬拜萬軍之耶和華，向他獻祭。在那裏有 以利 的兩個兒子 何弗尼 和 非尼哈 當耶和華的祭司。
1SAM|1|4|每逢獻祭的日子， 以利加拿 把祭肉分給他的妻子 毗尼拿 和 毗尼拿 所生的兒女。
1SAM|1|5|他給 哈拿 的卻是雙分，因為他愛 哈拿 。耶和華卻不使 哈拿 生育。
1SAM|1|6|她的對頭 毗尼拿 因耶和華不使 哈拿 生育，就常常惹她發怒，要使她生氣。
1SAM|1|7|年年都是如此。每當她上到耶和華殿的時候， 毗尼拿 就這樣惹她發怒，以致她哭泣不吃飯。
1SAM|1|8|她丈夫 以利加拿 對她說：「 哈拿 ，你為何哭泣？為何不吃飯？為何傷心難過呢？有我不比有十個兒子更好嗎？」
1SAM|1|9|他們在 示羅 吃喝完了， 哈拿 就站起來。祭司 以利 坐在耶和華殿門框旁邊的位子上。
1SAM|1|10|哈拿 心裏愁苦，就痛痛哭泣，向耶和華祈禱。
1SAM|1|11|她許願說：「萬軍之耶和華啊，你若垂顧你使女的苦情，眷念不忘你的使女，賜你的使女一個子嗣，我必使他終生歸給耶和華，不用剃刀剃他的頭。」
1SAM|1|12|哈拿 在耶和華面前不住地祈禱， 以利 注意她的嘴。
1SAM|1|13|哈拿 心中默禱，只動嘴唇，聽不到她的聲音，因此 以利 以為她喝醉了。
1SAM|1|14|以利 對她說：「你要醉到幾時呢？不要再喝酒了！」
1SAM|1|15|哈拿 回答說：「我主啊，不是這樣。我是心裏愁苦的婦人，清酒烈酒都沒有喝，只在耶和華面前傾心吐意。
1SAM|1|16|不要將你的使女看作不正經的女子。我因極其難過和生氣，所以一直禱告到如今。」
1SAM|1|17|以利 回答說：「平平安安地回去吧。願 以色列 的上帝允准你向他所求的！」
1SAM|1|18|哈拿 說：「願你的婢女在你眼前蒙恩。」於是婦人上路，去吃飯，臉上不再帶愁容了。
1SAM|1|19|他們清早起來，在耶和華面前敬拜，就回去，往 拉瑪 自己的家裏。 以利加拿 和妻子 哈拿 同房，耶和華顧念 哈拿 。
1SAM|1|20|時候到了， 哈拿 懷孕生了一個兒子， 哈拿 給他起名叫 撒母耳 ，說：「這是我從耶和華那裏求來的。」
1SAM|1|21|以利加拿 和他全家都上去，要向耶和華獻年祭和還願祭。
1SAM|1|22|哈拿 卻沒有上去，因為她對丈夫說：「等孩子斷了奶，我就帶他上去朝見耶和華，讓他永遠住在那裏。」
1SAM|1|23|她丈夫 以利加拿 對她說：「就照你看為好的去做吧！可以留到兒子斷了奶，願耶和華應驗他的話。」於是婦人留在家裏乳養兒子，直到斷了奶。
1SAM|1|24|斷奶之後，她就帶著孩子，連同一頭三歲的公牛 ，一伊法細麵 ，一皮袋酒，上 示羅 耶和華的殿去。那時，孩子還小。
1SAM|1|25|他們宰了公牛，就領孩子到 以利 面前。
1SAM|1|26|婦人說：「我主啊，請容許我說，我向你，我的主起誓，從前在你這裏站著祈求耶和華的那婦人就是我。
1SAM|1|27|我祈求為要得這孩子，耶和華已將我向他所求的賜給我了。
1SAM|1|28|所以，我將這孩子獻給耶和華，使他終生歸給耶和華。」 他就在那裏敬拜耶和華。
1SAM|2|1|哈拿 禱告說： 「我的心因耶和華快樂， 我的角因耶和華高舉。 我的口向仇敵張開； 我因你的救恩歡欣。
1SAM|2|2|「沒有一位聖者像耶和華， 除你以外沒有別的了， 也沒有磐石像我們的上帝。
1SAM|2|3|不要誇口說驕傲的話， 也不要口出狂妄的言語， 因耶和華是有知識的上帝， 人的行為被他衡量。
1SAM|2|4|勇士的弓折斷， 跌倒的人以力量束腰。
1SAM|2|5|飽足的人作雇工求食； 飢餓的人也不再飢餓。 不生育的生了七個； 兒女多的反倒孤獨。
1SAM|2|6|耶和華使人死，也使人活， 使人下陰間，也使人往上升。
1SAM|2|7|耶和華使人貧窮，也使人富足； 使人降卑，也使人升高。
1SAM|2|8|他從灰塵裏抬舉貧寒人， 從糞堆中提拔貧窮人， 使他們與貴族同坐， 繼承榮耀的座位。 地的柱子屬耶和華， 他將世界立在其上。
1SAM|2|9|「他必保護他聖民的腳步， 但惡人卻在黑暗中毀滅， 因為人不是靠力量得勝。
1SAM|2|10|與耶和華相爭的，必被打碎； 他必從天上打雷攻擊他們。 耶和華審判地極的人， 將力量賜給所立的王， 高舉受膏者的角。」
1SAM|2|11|以利加拿 往 拉瑪 回自己的家去了。那孩子在 以利 祭司面前事奉耶和華。
1SAM|2|12|以利 的兩個兒子是無賴，不認識耶和華。
1SAM|2|13|這二祭司對待百姓的規矩是這樣：凡有人獻祭，正煮肉的時候，祭司的僕人就手拿三齒的叉子來，
1SAM|2|14|將叉子往盆裏，或鍋裏，或釜裏，或壺裏一插，插上來的肉，祭司都拿了去。他們對所有上到 示羅 的 以色列 人都這樣做。
1SAM|2|15|甚至在未燒脂肪之前，祭司的僕人就來對獻祭的人說：「把肉給祭司，讓他烤吧。他不要拿你煮過的肉，要生的。」
1SAM|2|16|獻祭的人若說：「他們必須先燒脂肪，然後你才可以隨意拿。」僕人就說：「不，你立刻給我，不然我就要搶了。」
1SAM|2|17|這些年輕人的罪在耶和華面前非常嚴重，因為這些人藐視耶和華的祭物。
1SAM|2|18|那時， 撒母耳 還是孩子，穿著細麻布的以弗得，侍立在耶和華面前。
1SAM|2|19|他母親每年為他做一件小外袍，同丈夫上來獻年祭的時候帶來給他。
1SAM|2|20|以利 為 以利加拿 和他妻子祝福，說：「願耶和華由這婦人再賜你後裔，代替從耶和華求來的孩子。」他們就回自己的地方去了。
1SAM|2|21|耶和華眷顧 哈拿 ，她就懷孕生了三個兒子，兩個女兒。那孩子 撒母耳 在耶和華面前漸漸長大。
1SAM|2|22|以利 年紀老邁，聽見他兩個兒子對 以色列 眾人所做一切的事，又聽見他們與會幕門前伺候的婦人同寢，
1SAM|2|23|就對他們說：「你們為何做這樣的事呢？我從這眾百姓聽見了你們的惡行。
1SAM|2|24|我兒啊，不可這樣！我聽到耶和華的百姓傳出你們不好的名聲 。
1SAM|2|25|人若得罪人，有上帝 可以裁決；人若得罪耶和華，誰能為他代求呢？」然而他們還是不聽父親的話，因為耶和華想要他們死。
1SAM|2|26|撒母耳 這孩子漸漸長大，耶和華與人越發喜愛他。
1SAM|2|27|有神人來見 以利 ，對他說：「耶和華如此說：『你祖宗的家在 埃及 法老家 的時候，我不是向他們顯現嗎？
1SAM|2|28|在 以色列 眾支派中，我不是揀選他作我的祭司，上我的祭壇，燒香，在我面前穿以弗得嗎？我不是將 以色列 人所獻的火祭都賜給你祖宗的家嗎？
1SAM|2|29|你們為何踐踏我所吩咐獻在我居所的祭物和供物呢 ？你為何尊重你的兒子過於尊重我，將我百姓 以色列 所獻美好的祭物都拿去養肥你們自己呢？』
1SAM|2|30|因此，耶和華－ 以色列 的上帝說：『我確實說過，你和你祖宗的家必永遠行在我面前，但現在耶和華卻說，我絕不會這樣做。因為尊重我的，我必尊重他；藐視我的，他必被輕視。
1SAM|2|31|看哪，日子將到，我要折斷你的膀臂和你祖宗家的膀臂，使你家中沒有一個老年人。
1SAM|2|32|你在 以色列 人享福的時候必看見我居所的衰敗 ，你家中必永遠沒有一個老年人。
1SAM|2|33|你家中的人，我沒有從我壇前剪除的，必使你眼睛失明，心中憂傷。你家中所添的人口都必夭折。
1SAM|2|34|你的兩個兒子 何弗尼 、 非尼哈 所遭遇的事是給你的預兆：他們二人必在同一日死亡。
1SAM|2|35|我要為自己立一個忠心的祭司，他行事必照我的心、如我的意。我要為他建立堅固的家，他必天天行走在我受膏者的面前。
1SAM|2|36|你家所剩下的人都必來叩拜他，求一塊銀子，一個餅，說：求你給我一個祭司的職分，好使我得點餅吃。』」
1SAM|3|1|那孩子 撒母耳 在 以利 面前事奉耶和華。在那些日子，耶和華的言語稀少，不常有異象。
1SAM|3|2|那時， 以利 在自己的地方睡覺；他眼目開始昏花，不能看見。
1SAM|3|3|上帝的燈還沒有熄滅， 撒母耳 睡在耶和華的殿內，上帝的約櫃就在那裏。
1SAM|3|4|耶和華呼喚 撒母耳 ， 撒母耳 說：「我在這裏！」
1SAM|3|5|他跑到 以利 那裏，說：「你叫我嗎？我在這裏。」 以利 說：「我沒有叫你，回去睡吧。」他就回去睡了。
1SAM|3|6|耶和華又呼喚 撒母耳 。 撒母耳 起來，到 以利 那裏，說：「你叫我嗎？我在這裏。」 以利 說：「我兒，我沒有叫你，回去睡吧。」
1SAM|3|7|那時 撒母耳 還未認識耶和華，耶和華的話也未曾向他啟示。
1SAM|3|8|耶和華第三次再呼喚 撒母耳 。 撒母耳 起來，到 以利 那裏，說：「你叫我嗎？我在這裏。」 以利 才明白是耶和華呼喚這小孩。
1SAM|3|9|以利 對 撒母耳 說：「你回去睡吧。他若再叫你，你就說：『耶和華啊，請說，僕人敬聽！』」 撒母耳 就回去，仍睡在原處。
1SAM|3|10|耶和華來站著，像前幾次呼喚：「 撒母耳 ！ 撒母耳 ！」 撒母耳 說：「請說，僕人敬聽！」
1SAM|3|11|耶和華對 撒母耳 說：「看哪，我在 以色列 中必行一件事，凡聽見的人都必雙耳齊鳴。
1SAM|3|12|我指著 以利 家所說的話，到了時候，必從頭到尾應驗在 以利 身上。
1SAM|3|13|我曾告訴他，我必永遠懲罰他的家，因為他知道自己的兒子作惡，褻瀆上帝 ，卻不禁止他們。
1SAM|3|14|所以我向 以利 家起誓：『 以利 家的罪孽，就是獻祭物和供物，也永不得贖。』」
1SAM|3|15|撒母耳 睡到天亮，就開了耶和華殿的門。 撒母耳 害怕，不敢將異象告訴 以利 。
1SAM|3|16|以利 呼喚 撒母耳 說：「我兒 撒母耳 ！」 撒母耳 說：「我在這裏！」
1SAM|3|17|以利 說：「他對你說了甚麼話，你不要向我隱瞞。你若將他對你所說的話向我隱瞞一句，願上帝重重懲罰你。」
1SAM|3|18|撒母耳 就把一切話都告訴 以利 ，並沒有隱瞞。 以利 說：「他是耶和華，願他照他看為好的去做。」
1SAM|3|19|撒母耳 長大了，耶和華與他同在，使他所說的話一句都不落空。
1SAM|3|20|從 但 到 別是巴 ，所有的 以色列 人都知道耶和華立 撒母耳 為先知。
1SAM|3|21|耶和華又在 示羅 顯現，因為耶和華在 示羅 藉他的話向 撒母耳 啟示他自己。
1SAM|4|1|撒母耳 的話傳遍了全 以色列 。 以色列 人出去與 非利士 人打仗，安營在 以便‧以謝 ， 非利士 人安營在 亞弗 。
1SAM|4|2|非利士 人向 以色列 人擺陣。兩軍交戰的時候， 以色列 人敗在 非利士 人面前； 非利士 人在戰場上殺了他們約四千人。
1SAM|4|3|百姓回到營裏， 以色列 的長老說：「耶和華今日為何使我們敗在 非利士 人面前呢？我們要將耶和華的約櫃從 示羅 抬到我們這裏來，好讓他來到我們中間，救我們脫離敵人的手掌。」
1SAM|4|4|於是百姓派人到 示羅 ，從那裏將坐在二基路伯上萬軍之耶和華的約櫃抬來。 以利 的兩個兒子 何弗尼 、 非尼哈 也與上帝的約櫃同來。
1SAM|4|5|耶和華的約櫃到了營中，全 以色列 就大聲歡呼，連地都震動。
1SAM|4|6|非利士 人聽見歡呼的聲音，就說：「為何 希伯來 人在營裏這麼大聲歡呼呢？」他們知道耶和華的約櫃到了營中。
1SAM|4|7|非利士 人就懼怕，說：「有神明到了他們營中。」又說：「我們有禍了！從來不曾有這樣的事。
1SAM|4|8|我們有禍了！誰能救我們脫離這些大能之神明的手呢？從前在曠野用各樣災禍擊打 埃及 人的，就是這些神明。
1SAM|4|9|非利士 人哪，要剛強，要作大丈夫，免得作 希伯來 人的奴僕，如同他們作你們的奴僕一樣。你們要作大丈夫，與他們爭戰。」
1SAM|4|10|非利士 人進攻， 以色列 人敗了，各往自己的家逃跑。被殺的人很多， 以色列 倒下的步兵有三萬。
1SAM|4|11|上帝的約櫃被擄去， 以利 的兩個兒子 何弗尼 、 非尼哈 也都被殺了。
1SAM|4|12|有一個 便雅憫 人從戰場上逃跑，衣服撕裂，頭蒙灰塵，當日來到 示羅 。
1SAM|4|13|他到了的時候，看哪， 以利 正坐在路旁的位子上觀望，為上帝的約櫃心裏擔憂。那人進城報信，全城的人就都呼喊起來。
1SAM|4|14|以利 聽見呼喊的聲音就說：「這喧嚷的聲音是甚麼呢？」那人急忙來報信給 以利 。
1SAM|4|15|那時 以利 九十八歲了，兩眼發直，不能看見。
1SAM|4|16|那人對 以利 說：「我是從戰場上來的，今日剛從戰場上逃回來。」 以利 說：「我兒，事情怎樣了？」
1SAM|4|17|報信的回答說：「 以色列 人在 非利士 人面前逃跑，百姓中被殺的很多！你的兩個兒子 何弗尼 和 非尼哈 也都死了，並且上帝的約櫃已經被擄去了。」
1SAM|4|18|他一提到上帝的約櫃， 以利 就從城門旁自己的位子上往後跌倒，折斷頸項而死，因為他年紀老邁，身體沉重。 以利 作 以色列 的士師四十年。
1SAM|4|19|以利 的媳婦， 非尼哈 的妻子懷孕將到產期，她聽見上帝的約櫃被擄，公公和丈夫都死了，就曲身生產，極其疼痛。
1SAM|4|20|她將要死的時候，旁邊站著的婦人們對她說：「不要怕！你生了男孩了。」她不回答，也不放在心上。
1SAM|4|21|她給孩子起名叫 以迦博 ，說：「榮耀離開 以色列 了！」這是因為上帝的約櫃被擄去，又因為她公公和丈夫都死了。
1SAM|4|22|她又說：「榮耀離開 以色列 ，因為上帝的約櫃被擄去了。」
1SAM|5|1|非利士 人擄去上帝的約櫃，從 以便‧以謝 帶到 亞實突 。
1SAM|5|2|非利士 人擄了上帝的約櫃，帶進 大袞 廟，放在 大袞 的旁邊。
1SAM|5|3|次日， 亞實突 人清早起來，看哪， 大袞 仆倒在耶和華的約櫃前，臉伏於地，他們就扶起 大袞 ，把它放回原處。
1SAM|5|4|又次日，他們清早起來，看哪， 大袞 仆倒在耶和華的約櫃前，臉伏於地，並且 大袞 的頭和兩手都在門檻上折斷，只剩下 大袞 的軀幹。
1SAM|5|5|因此， 大袞 的祭司和所有進 大袞 廟的人，都不踏 亞實突 的 大袞 廟的門檻，直到今日。
1SAM|5|6|耶和華的手重重擊打 亞實突 人，使他們恐懼，使 亞實突 和 亞實突 周圍的人都生痔瘡。
1SAM|5|7|亞實突 人見這情況，就說：「 以色列 上帝的約櫃不可留在我們這裏，因為他的手重重擊打我們和我們的神明 大袞 」。
1SAM|5|8|他們就派人去請 非利士 的眾領袖來聚集，對他們說：「我們向 以色列 上帝的約櫃應當怎樣做呢？」他們說：「可以把 以色列 上帝的約櫃運到 迦特 去。」於是他們把 以色列 上帝的約櫃運到那裏。
1SAM|5|9|運到之後，耶和華的手擊打那城，使那城的人非常驚慌，無論大小都生痔瘡。
1SAM|5|10|他們就把上帝的約櫃送到 以革倫 。上帝的約櫃到了 以革倫 ， 以革倫 人就呼喊說：「他們把 以色列 上帝的約櫃運到我這裏，要害我和我的百姓！」
1SAM|5|11|於是他們派人去請 非利士 的眾領袖來，說：「請你們把 以色列 上帝的約櫃送回原處，免得害死我和我的百姓！」原來上帝的手重重攻擊那城，死亡的恐懼瀰漫全城，
1SAM|5|12|沒有死的人都受痔瘡的折磨。城裏的哀聲上達於天。
1SAM|6|1|耶和華的約櫃在 非利士 人之地七個月。
1SAM|6|2|非利士 人召了祭司和占卜的來，說：「我們向耶和華的約櫃應當怎樣做呢？請指示我們要用甚麼方法把約櫃送回原處。」
1SAM|6|3|他們說：「若要將 以色列 上帝的約櫃送回去，不可空手送回，一定要給他獻賠罪的禮物，然後你們才可以得痊癒，並且知道他的手為何不離開你們。」
1SAM|6|4|非利士 人說：「應當用甚麼獻為賠罪的禮物呢？」他們說：「當按照 非利士 領袖的數目，獻五個金痔瘡和五個金老鼠，因為你們眾人和領袖所遭遇的都是一樣的災禍。
1SAM|6|5|當製造你們痔瘡的像和毀壞田地老鼠的像，並要將榮耀歸給 以色列 的上帝，或者他向你們和你們的神明，以及你們的田地，把手放輕些。
1SAM|6|6|你們為何硬著心，像 埃及 人和法老硬著心一樣呢？上帝豈不是嚴厲對付 埃及 ，使 埃及 人釋放 以色列 人，他們就走了嗎？
1SAM|6|7|現在你們應當造一輛新車，把兩頭未曾負軛，還在哺乳的母牛套在車上，趕牛犢離開母牛，回家去。
1SAM|6|8|你們要把耶和華的約櫃放在車上，把所獻賠罪的金器裝在匣子裏，放在櫃旁，送走櫃子，讓它去。
1SAM|6|9|你們要觀察：車若直行過 以色列 的邊界，上到 伯‧示麥 去，這大災禍就是耶和華降在我們身上的；若不然，我們就知道，這不是他的手擊打我們，而是我們偶然遭遇的。」
1SAM|6|10|非利士 人就照樣做了。他們取了兩頭哺乳的母牛套在車上，把牛犢關在家裏，
1SAM|6|11|把耶和華的約櫃和裝金老鼠以及金痔瘡像的匣子都放在車上。
1SAM|6|12|牛直行大路，在往 伯‧示麥 的一條大道上，一面走一面叫，不偏左右。 非利士 的領袖跟在後面，直到 伯‧示麥 的地界。
1SAM|6|13|那時， 伯‧示麥 人正在平原收割麥子，舉目看見約櫃，就歡歡喜喜地迎見它。
1SAM|6|14|車到了 伯‧示麥 人 約書亞 的田間，就在那裏停了。在那裏有一塊大磐石，他們把車的木頭劈了，把兩頭母牛獻給耶和華為燔祭。
1SAM|6|15|利未 人將耶和華的約櫃和櫃子旁邊裝金器的匣子拿下來，放在大磐石上。當日 伯‧示麥 人獻上燔祭，又獻其他祭物給耶和華。
1SAM|6|16|非利士 人的五個領袖看見了，當日就回 以革倫 去。
1SAM|6|17|非利士 人獻給耶和華作賠罪的金痔瘡像如下：一個為 亞實突 ，一個為 迦薩 ，一個為 亞實基倫 ，一個為 迦特 ，一個為 以革倫 。
1SAM|6|18|金老鼠的數目是按照 非利士 五個領袖的城鎮，就是堅固的城鎮和鄉村，以及大磐石。這磐石是安放耶和華約櫃的，到今日還在 伯‧示麥 人 約書亞 的田間。
1SAM|6|19|耶和華擊殺 伯‧示麥 人，因為他們觀看他的約櫃。他擊殺了百姓七十人 。百姓因耶和華大大擊殺他們，就哀哭了。
1SAM|6|20|伯‧示麥 人說：「誰能在耶和華這位聖潔的上帝面前侍立呢？這約櫃可以從我們這裏上到誰那裏去呢？」
1SAM|6|21|於是他們派使者到 基列‧耶琳 的居民那裏，說：「 非利士 人將耶和華的約櫃送回來了，你們下來將約櫃接了，上到你們那裏去吧！」
1SAM|7|1|基列‧耶琳 人就來了，將耶和華的約櫃接上去，抬到山上 亞比拿達 的家中，將他兒子 以利亞撒 分別為聖，看守耶和華的約櫃。
1SAM|7|2|從約櫃留在 基列‧耶琳 的那天起，經過了許多日子，有二十年； 以色列 全家都哀哭歸向耶和華。
1SAM|7|3|撒母耳 對 以色列 全家說：「你們若全心回轉歸向耶和華，就要從你們中間除掉外邦的神明和 亞斯她錄 ，預備你們的心歸向耶和華，單單事奉他，他必救你們脫離 非利士 人的手。」
1SAM|7|4|以色列 人就除掉諸 巴力 和 亞斯她錄 ，單單事奉耶和華。
1SAM|7|5|撒母耳 說：「要召集 以色列 眾人到 米斯巴 去，我好為你們向耶和華禱告。」
1SAM|7|6|他們就聚集在 米斯巴 ，打水澆在耶和華面前。當日他們禁食，說：「我們得罪了耶和華。」 撒母耳 在 米斯巴 作 以色列 人的士師。
1SAM|7|7|非利士 人聽見 以色列 人聚集在 米斯巴 ， 非利士 的領袖就上來要攻擊 以色列 。 以色列 人聽見，就懼怕 非利士 人。
1SAM|7|8|以色列 人對 撒母耳 說：「願你不住為我們呼求耶和華－我們的上帝，救我們脫離 非利士 人的手。」
1SAM|7|9|撒母耳 就把一隻吃奶的羔羊獻給耶和華作全牲的燔祭，為 以色列 人呼求耶和華，耶和華就應允他。
1SAM|7|10|撒母耳 正獻燔祭的時候， 非利士 人前來要與 以色列 爭戰。當日，耶和華打雷，發出極大的聲音，使 非利士 人潰亂，他們就敗在 以色列 面前。
1SAM|7|11|以色列 人從 米斯巴 出來，追趕 非利士 人，擊殺他們，直到 伯‧甲 的下邊。
1SAM|7|12|撒母耳 拿一塊石頭立在 米斯巴 和 善 的中間，給石頭起名叫 以便‧以謝 ，說：「到如今耶和華都幫助我們。」
1SAM|7|13|因此， 非利士 人被制伏了，不再入侵 以色列 境內。 撒母耳 有生之年，耶和華的手攻擊 非利士 人。
1SAM|7|14|非利士 人所奪取 以色列 的城鎮，從 以革倫 直到 迦特 ，都歸回 以色列 了。 以色列 也從 非利士 人手中收回這些城所屬的地界。那時 以色列 與 亞摩利 人和平相處。
1SAM|7|15|撒母耳 一生作 以色列 的士師。
1SAM|7|16|他每年巡行到 伯特利 、 吉甲 、 米斯巴 ，在這些地方審判 以色列 人。
1SAM|7|17|隨後他回到 拉瑪 ，因為他的家在那裏；他在那裏審判 以色列 人，並且在那裏為耶和華築了一座壇。
1SAM|8|1|撒母耳 年紀老邁，就立他的兒子作 以色列 的士師。
1SAM|8|2|他的長子名叫 約珥 ，次子名叫 亞比亞 ；他們在 別是巴 作士師。
1SAM|8|3|他的兒子不行他的道，貪圖財利，收取賄賂，屈枉正直。
1SAM|8|4|以色列 的長老都聚集在 拉瑪 ，來到 撒母耳 那裏，
1SAM|8|5|對他說：「看哪，你年紀老了，你的兒子又不行你的道。現在請你為我們立一個王治理我們，像列國一樣。」
1SAM|8|6|撒母耳 不喜悅他們說「立一個王治理我們」，他就向耶和華禱告。
1SAM|8|7|耶和華對 撒母耳 說：「你只管聽從百姓向你說的一切話，因為他們不是厭棄你，而是厭棄我，不要我作他們的王。
1SAM|8|8|自從我領他們出 埃及 的日子到如今，他們離棄我，事奉別神；正像他們從前所做的一切事，現在他們也照樣向你做了。
1SAM|8|9|現在你只管聽從他們的話，不過要嚴厲警告他們，告訴他們將來王會用甚麼方式管轄他們。」
1SAM|8|10|撒母耳 將耶和華一切的話轉告求他立王的百姓。
1SAM|8|11|他說：「管轄你們的王必用這樣的方式：他必派你們的兒子為他駕車，趕馬，在他的戰車前奔跑。
1SAM|8|12|他要為自己立千夫長、五十夫長；耕種他的田地，收割他的莊稼；打造他的兵器和車上的器械。
1SAM|8|13|他必叫你們的女兒為他製造香膏，作廚師與烤餅的，
1SAM|8|14|也必取你們最好的田地、葡萄園、橄欖園，賜給他的臣僕。
1SAM|8|15|你們的糧食和葡萄園所出產的，他必徵收十分之一給他的官員和臣僕，
1SAM|8|16|又必叫你們的僕人婢女，健壯的青年和你們的驢為他做工。
1SAM|8|17|你們的羊群，他必徵收十分之一，你們自己也必作他的僕人。
1SAM|8|18|那日，你們必因自己所選的王哀求耶和華，但那日耶和華卻不應允你們。」
1SAM|8|19|百姓卻不肯聽 撒母耳 的話，說：「不！我們一定要一個王治理我們，
1SAM|8|20|使我們像列國一樣，有王治理我們，率領我們，為我們爭戰。」
1SAM|8|21|撒母耳 聽見百姓這一切話，就稟告給耶和華聽。
1SAM|8|22|耶和華對 撒母耳 說：「你只管聽從他們的話，為他們立一個王。」 撒母耳 對 以色列 人說：「去，你們各歸各城吧！」
1SAM|9|1|有一個 便雅憫 人名叫 基士 ，是 便雅憫 人 亞斐亞 的玄孫， 比歌拉 的曾孫， 洗羅 的孫子， 亞別 的兒子，是個大能的勇士 。
1SAM|9|2|他有一個兒子名叫 掃羅 ，又健壯、又英俊，在 以色列 人中沒有一個可以與他相比；他比眾百姓高出一個頭 。
1SAM|9|3|掃羅 的父親 基士 丟失了幾匹母驢，他就吩咐兒子 掃羅 說：「起來，帶一個僕人去尋找驢子。」
1SAM|9|4|掃羅 走過 以法蓮 山區，又過 沙利沙 地，都沒有找著。他們走過 沙琳 地，驢不在那裏，又走過 便雅憫 地，也沒有找到。
1SAM|9|5|到了 蘇弗 地， 掃羅 對跟隨他的僕人說：「我們不如回去，免得我父親不為驢掛慮，反為我們擔憂。」
1SAM|9|6|僕人對他說：「看哪，這城裏有一位神人，受人敬重，凡他所說的全都應驗。現在讓我們到他那裏去，或者他能指示我們當走的路。」
1SAM|9|7|掃羅 對僕人說：「看哪，我們若去，送甚麼給那人呢？我們袋子裏的食物都吃完了，也沒有禮物可以送給神人，我們還有些甚麼呢？」
1SAM|9|8|僕人又回答 掃羅 說：「看哪，我手裏還有四分之一舍客勒的銀子，可以送給神人，請他指示我們當走的路。」
1SAM|9|9|從前 以色列 中，若有人去求問上帝，就這麼說：「來，我們到先見那裏去吧！」因現在的先知，從前稱為先見。
1SAM|9|10|掃羅 對僕人說：「好主意！來，我們去吧。」於是他們往神人所住的城裏去了。
1SAM|9|11|他們上坡要進城，遇見幾個少女出來打水，就問她們說：「先見有沒有在這裏呢？」
1SAM|9|12|她們回答說：「有的，看哪，他就在你們前面。快！他今日正來到城裏，因為今日百姓要在丘壇獻祭。
1SAM|9|13|你們一進城，他還沒有上丘壇吃祭物之前，就會遇見他。因為他沒有到，百姓不能吃，必須等他先為祭物祝謝，然後受邀的人才可以吃。現在就上去吧，因為這時候你們會遇見他。」
1SAM|9|14|他們就上到那城，進入城中的時候，看哪， 撒母耳 正迎著他們來，要上丘壇去。
1SAM|9|15|掃羅 還沒有到的前一日，耶和華已經對 撒母耳 啟示說：
1SAM|9|16|「明日這時候，我必使一個人從 便雅憫 地到你這裏來，你要膏他作我百姓 以色列 的君王。他必救我的百姓脫離 非利士 人的手，因為我眷顧我的百姓 ，他們的哀聲已上達於我。」
1SAM|9|17|撒母耳 看見 掃羅 的時候，耶和華對他說：「看哪，這就是我對你所說的人，他必治理我的百姓。」
1SAM|9|18|掃羅 在城門中走到 撒母耳 跟前，說：「請告訴我，先見的家在哪裏？」
1SAM|9|19|撒母耳 回答掃羅說：「我就是先見。你在我前面先上丘壇去，因為你們今日必跟我同席。明日早晨我送你走，會把你心裏一切的事都告訴你。
1SAM|9|20|至於你前三日所丟失的幾匹母驢，你心裏不必掛慮，都已經找到了。 以色列 眾人所仰慕的是誰呢？不是仰慕你和你父的全家嗎？」
1SAM|9|21|掃羅 回答說：「我不是 以色列 支派中最小的 便雅憫 人嗎？我的家族不是 便雅憫 支派中最小的家族嗎？你為何對我說這樣的話呢？」
1SAM|9|22|撒母耳 領 掃羅 和他的僕人進了大廳，使他們在受邀的人中坐首位；受邀者約有三十個。
1SAM|9|23|撒母耳 對廚師說：「我交給你的那一份祭肉，吩咐你收存的，現在可以拿來。」
1SAM|9|24|廚師就舉起祭肉的腿和腿上的部分 ，擺在 掃羅 面前。 撒母耳 說：「看哪，所存留的擺在你面前了。吃吧！因為這是為你保留到這特定的時候的，好讓你說，是我請了這百姓來，」 當日， 掃羅 就與 撒母耳 同席。
1SAM|9|25|他們從丘壇下來進城， 撒母耳 和 掃羅 在房頂上說話。
1SAM|9|26|次日他們清早起來。黎明的時候， 撒母耳 呼叫在房頂上的 掃羅 ，說：「起來，我好送你回去。」 掃羅 就起來，和 撒母耳 二人一同到外面去。
1SAM|9|27|二人下到城邊， 撒母耳 對 掃羅 說：「你要吩咐僕人先走，僕人走了以後， 你要留在這裏，這時候我要將上帝的話傳給你聽。」
1SAM|10|1|撒母耳 拿一瓶膏油倒在 掃羅 的頭上，親吻他，說：「耶和華豈不是膏你作他產業的君王嗎？
1SAM|10|2|你今日離開我之後，會在 便雅憫 境內的 謝撒 ，靠近 拉結 的墳墓，遇見兩個人。他們會對你說：『你要找的幾匹母驢已經找到了。看哪，你父親不為驢子的事掛慮，反為你擔憂，說：我為兒子該做些甚麼呢？』
1SAM|10|3|你從那裏往前走，到了 他泊 的橡樹那裏，會遇見三個往 伯特利 去敬拜上帝的人：一個帶著三隻小山羊，一個帶著三個餅，一個帶著一皮袋酒。
1SAM|10|4|他們會向你問安，給你兩個餅，你就從他們手中接過來。
1SAM|10|5|然後你要到上帝的山去，在那裏有 非利士 的駐軍。你到了城裏的時候，會遇見一隊先知從丘壇下來，前面有鼓瑟的、擊鼓的、吹笛的、彈琴的，他們都受感說話。
1SAM|10|6|耶和華的靈必大大感動你，你就與他們一同受感說話，轉變成另一個人。
1SAM|10|7|這徵兆臨到你，你就要趁機做該做的事，因為上帝與你同在。
1SAM|10|8|你要在我以先下到 吉甲 。看哪，我必下到你那裏獻燔祭和平安祭。你要等候七日，等我到你那裏指示你當做的事。」
1SAM|10|9|掃羅 轉身離開 撒母耳 ，上帝就改變他，賜給他另一顆心。當日這一切徵兆都應驗了。
1SAM|10|10|他們來到那座山，看哪，有一隊先知遇見 掃羅 。上帝的靈大大感動他，他就在先知中受感說話。
1SAM|10|11|所有先前認識 掃羅 的人看見了，看哪，他和先知一同受感說話，百姓就彼此說：「 基士 的兒子遇見了甚麼呢？ 掃羅 也在先知中嗎？」
1SAM|10|12|那地方有一個人說：「這些人的父親是誰呢？」因此就有一句俗語說：「 掃羅 也在先知中嗎？」
1SAM|10|13|掃羅 受感說完了話，就上丘壇去了。
1SAM|10|14|掃羅 的叔叔問 掃羅 和他的僕人說：「你們到哪裏去了？」他說：「我們找驢子去了。但我們找不到，就去了 撒母耳 那裏。」
1SAM|10|15|掃羅 的叔叔說：「告訴我 撒母耳 對你們說了些甚麼。」
1SAM|10|16|掃羅 對他的叔叔說：「他明明告訴我們，驢子已經找到了。」至於 撒母耳 所說君王的事， 掃羅 沒有告訴叔叔。
1SAM|10|17|撒母耳 召集百姓到 米斯巴 耶和華那裏。
1SAM|10|18|他對 以色列 眾人說：「耶和華－ 以色列 的上帝如此說：『我領 以色列 出 埃及 ，救你們脫離 埃及 人的手，以及脫離欺壓你們各國之人的手。』
1SAM|10|19|你們今日卻厭棄救你們脫離一切災禍和患難的上帝，對他說：『求你立一個王治理我們。』現在你們應當按支派和宗族站在耶和華面前。」
1SAM|10|20|於是， 撒母耳 叫 以色列 眾支派近前來抽籤，抽到了 便雅憫 支派。
1SAM|10|21|然後，他叫 便雅憫 支派按宗族近前來，抽到了 瑪特利 族，接著又抽到了 基士 的兒子 掃羅 。眾人尋找他卻找不到，
1SAM|10|22|就再問耶和華說：「那人來到這裏了沒有？」耶和華說：「看哪，他藏在物品堆中。」
1SAM|10|23|眾人就跑去從那裏領他出來。他站在百姓中間，比眾百姓高出一個頭。
1SAM|10|24|撒母耳 對眾百姓說：「你們看到了耶和華所揀選的人嗎？眾百姓中沒有人可以與他相比。」眾百姓就歡呼說：「願王萬歲！」
1SAM|10|25|撒母耳 將君王的典章對百姓說明，又記在書上，放在耶和華面前，然後 撒母耳 遣散眾百姓，各回自己的家去了。
1SAM|10|26|掃羅 也往 基比亞 自己的家去，有一群心中被上帝感動的勇士跟隨他。
1SAM|10|27|但有些無賴之輩說：「這人怎麼能救我們呢？」他們就藐視他，不送禮物給他。 掃羅 卻保持沉默。
1SAM|11|1|亞捫 人 拿轄 上來，對著 基列 的 雅比 安營。 雅比 眾人對 拿轄 說：「你與我們立約，我們就服事你。」
1SAM|11|2|亞捫 人 拿轄 對他們說：「你們若由我挖出你們各人的右眼，以此凌辱 以色列 眾人，我就與你們立約。」
1SAM|11|3|雅比 的長老對他說：「求你寬容我們七日，等我們派人到 以色列 的全境去。若沒有人來救我們，我們就出來歸順你。」
1SAM|11|4|使者到了 掃羅 住的 基比亞 ，把這事說給百姓聽，眾百姓就都放聲大哭。
1SAM|11|5|看哪， 掃羅 正從田間趕牛回來，說：「百姓為甚麼哭呢？」眾人把 雅比 人的話告訴他。
1SAM|11|6|掃羅 聽見這些話，就被上帝的靈催逼，大發怒氣。
1SAM|11|7|他把一對牛切成小塊，吩咐使者傳送到 以色列 全境，說：「凡不出來跟隨 掃羅 和 撒母耳 的，就必這樣待他的牛。」耶和華使百姓懼怕，他們就都出來如同一人。
1SAM|11|8|掃羅 在 比色 數點他們： 以色列 人有三十萬， 猶大 人有三萬。
1SAM|11|9|他們對那些來的使者說：「你們要對 基列 的 雅比 人這樣說，明天太陽快到中午的時候，你們必得解救。」使者回去告訴 雅比 人，他們就歡喜了。
1SAM|11|10|於是 雅比 人對 亞捫 人說：「明日我們出來歸順你們，可以照你們看為好的待我們。」
1SAM|11|11|第二日， 掃羅 把百姓分為三隊，在清晨換崗哨的時候入侵 亞捫 人的軍營，擊殺他們直到中午的時候。逃脫的人都分散了，甚至沒有兩個人同在一起。
1SAM|11|12|百姓對 撒母耳 說：「那說『 掃羅 豈能作我們的王』的是誰呢？把他們交出來，我們好處死他們。」
1SAM|11|13|掃羅 說：「今日耶和華在 以色列 中施行拯救，所以今日不可處死人。」
1SAM|11|14|撒母耳 對百姓說：「來，我們到 吉甲 去，在那裏開始新的王國。」
1SAM|11|15|眾百姓到了 吉甲 那裏，在耶和華面前擁立 掃羅 為王，又在耶和華面前獻平安祭。 掃羅 和 以色列 眾人在那裏都非常歡喜。
1SAM|12|1|撒母耳 對 以色列 眾人說：「看哪，我已聽了你們對我所說一切的話，為你們立了一個王。
1SAM|12|2|現在，看哪，有這王行走在你們前面。我已年老髮白，看哪，我的兒子都在你們這裏。我從幼年直到今日都行走在你們前面。
1SAM|12|3|我在這裏，你們要在耶和華和他的受膏者面前為我作證，我奪過誰的牛，搶過誰的驢，欺負過誰，虐待過誰，從誰手裏收過賄賂而蒙蔽自己的眼目呢？若有，我必償還。」
1SAM|12|4|眾人說：「你未曾欺負我們，虐待我們，也未曾從任何人手裏收過任何東西。」
1SAM|12|5|撒母耳 對他們說：「你們在我手裏沒有找著甚麼，有耶和華在你們中間作證，也有他的受膏者今日作證。」他們說 ：「願耶和華作證。」
1SAM|12|6|撒母耳 對百姓說：「從前立 摩西 和 亞倫 ，又領你們祖先出 埃及 地的是耶和華。
1SAM|12|7|現在你們要站住，讓我在耶和華面前，以耶和華向你們和你們祖先所行一切公義的事來和你們爭辯。
1SAM|12|8|從前 雅各 到了 埃及 ，後來你們的祖先呼求耶和華，耶和華就差遣 摩西 和 亞倫 領你們的祖先出 埃及 ，來到這地方居住。
1SAM|12|9|他們卻忘記耶和華－他們的上帝，他就把他們交給 夏瑣 將軍 西西拉 的手中，以及 非利士 人和 摩押 王的手中 。於是這些人常來攻擊他們。
1SAM|12|10|他們呼求耶和華說：『我們離棄了耶和華去事奉諸 巴力 和 亞斯她錄 ，我們有罪了。現在求你救我們脫離仇敵的手，我們必事奉你。』
1SAM|12|11|耶和華就差遣 耶路巴力 、 比但 、 耶弗他 、 撒母耳 救你們脫離四圍仇敵的手，你們才安然居住。
1SAM|12|12|你們見 亞捫 人的王 拿轄 來攻擊你們，就對我說：『不，要有一個王治理我們。』其實耶和華－你們的上帝是你們的王。
1SAM|12|13|現在，看哪，這就是你們所選的、你們所求的王。看哪，耶和華已經為你們立王了。
1SAM|12|14|你們若敬畏耶和華，事奉他，聽從他的話，不違背耶和華的命令，你們和治理你們的王也都跟從耶和華－你們的上帝就好了。
1SAM|12|15|倘若不聽從耶和華的話，違背他的命令，耶和華的手必攻擊你們，像從前攻擊你們祖先一樣。
1SAM|12|16|現在你們要站住，看耶和華在你們眼前要行的一件大事。
1SAM|12|17|這不是割麥子的時候嗎？我求告耶和華，他必打雷降雨，讓你們知道並且看出，你們為自己求立王的事在耶和華眼前是犯大罪了。」
1SAM|12|18|於是 撒母耳 求告耶和華，耶和華就在這日打雷降雨，眾百姓就非常懼怕耶和華和 撒母耳 。
1SAM|12|19|眾百姓對 撒母耳 說：「請你為僕人向耶和華－你的上帝禱告，免得我們死亡，因為我們求立王的事，正是罪上加罪了。」
1SAM|12|20|撒母耳 對百姓說：「不要懼怕！你們雖然行了這惡，卻不要偏離耶和華，只要盡心事奉他。
1SAM|12|21|不可偏離去隨從那沒有益處、不能救人的虛無的神明 ，因為它們是虛無的。
1SAM|12|22|耶和華必因他大名的緣故不撇棄他的子民，因為耶和華喜悅你們作他的子民。
1SAM|12|23|至於我，我如果停止為你們禱告，就得罪耶和華了，我絕不會這樣做。我必以善道正路指教你們。
1SAM|12|24|但你們要敬畏耶和華，誠誠實實地盡心事奉他，因你們要留意，他向你們所行的事何等大。
1SAM|12|25|你們若不斷作惡，你們和你們的王必一同滅亡。」
1SAM|13|1|掃羅 登基的時候年三十 歲，作 以色列 王二年 。
1SAM|13|2|掃羅 從 以色列 中選出三千人：二千跟隨 掃羅 在 密抹 和 伯特利 山區，一千跟隨 約拿單 在 便雅憫 的 基比亞 。其餘的百姓， 掃羅 打發他們各自回自己的帳棚去了。
1SAM|13|3|約拿單 攻擊 非利士 人在 迦巴 的駐軍， 非利士 人聽見了這事。 掃羅 就在遍地吹角，說：「讓 希伯來 人都聽見。」
1SAM|13|4|以色列 眾人聽見 掃羅 攻擊 非利士 的駐軍，又聽見 以色列 為 非利士 人所憎惡，百姓就跟隨 掃羅 ，在 吉甲 集合。
1SAM|13|5|非利士 人集合，要與 以色列 人作戰。他們有戰車三萬輛，騎兵六千，士兵像海邊的沙那樣多。他們上來，在 伯‧亞文 東邊的 密抹 安營。
1SAM|13|6|以色列 人見自己危急，軍隊被圍攻，百姓就藏在山洞、叢林、巖隙、地窖和深坑中。
1SAM|13|7|有些 希伯來 人過了 約旦河 ，逃到 迦得 和 基列 地。 掃羅 還在 吉甲 ，所有的人都戰戰兢兢地跟隨他。
1SAM|13|8|掃羅 照著 撒母耳 所定的日期等了七日。但是， 撒母耳 還沒有來到 吉甲 ，百姓就離開 掃羅 散去了。
1SAM|13|9|於是 掃羅 說：「把燔祭和平安祭帶到我這裏來。」 掃羅 就獻上燔祭。
1SAM|13|10|他剛獻完燔祭，看哪， 撒母耳 就到了。 掃羅 出去迎接他，向他問安。
1SAM|13|11|撒母耳 說：「你做了甚麼事啊？」 掃羅 說：「因為我見百姓離開我散去，你又不照所定的日期來到，而且 非利士 人已在 密抹 集合；
1SAM|13|12|我說：『現在 非利士 人已經下到 吉甲 來攻擊我，可是我還沒有向耶和華禱告。』所以我就勉強獻上燔祭。」
1SAM|13|13|撒母耳 對 掃羅 說：「你做了糊塗事了，沒有遵守耶和華－你上帝吩咐你的命令。不然，耶和華會在 以色列 中堅立你的國度，直到永遠。
1SAM|13|14|現在你的國度必不長久。耶和華已經尋著一個合他心意的人，立他作百姓的君王，因為你沒有遵守耶和華所吩咐你的。」
1SAM|13|15|撒母耳 就起來，從 吉甲 上到 便雅憫 的 基比亞 。 掃羅 數點跟隨他的百姓，約有六百人。
1SAM|13|16|掃羅 和他兒子 約拿單 ，以及跟隨他們的百姓，都住在 便雅憫 的 迦巴 ， 非利士 人卻在 密抹 安營。
1SAM|13|17|有突擊隊從 非利士 營中出來，分成三隊：一隊往 俄弗拉 到 書亞 地去，
1SAM|13|18|一隊往 伯‧和崙 去，一隊往邊界，下望朝著曠野的 洗波音谷 。
1SAM|13|19|那時， 以色列 全地找不到一個鐵匠，因為 非利士 人說：「恐怕 希伯來 人製造刀槍。」
1SAM|13|20|以色列 眾人要磨鋤、犁、斧、鏟，就各自下到 非利士 人那裏去磨。
1SAM|13|21|磨鋤或犁的價錢是三分之二舍客勒，磨斧或修整刺棒的價錢是三分之一舍客勒。
1SAM|13|22|所以到了戰爭的日子，所有跟隨 掃羅 和 約拿單 的百姓找不到一個手裏有刀有槍的，惟 掃羅 和他兒子 約拿單 有。
1SAM|13|23|非利士 人的一隊駐軍出來，到 密抹 的隘口。
1SAM|14|1|有一日， 掃羅 的兒子 約拿單 對拿他兵器的青年說：「來，我們過去到 非利士 的駐軍那裏。」但他沒有告訴父親。
1SAM|14|2|掃羅 在 基比亞 的郊外，坐在 米磯崙 的石榴樹下，跟隨他的百姓約有六百人。
1SAM|14|3|在那裏有 亞希突 的兒子 亞希亞 ，穿著以弗得。 亞希突 是 以迦博 的哥哥， 非尼哈 的兒子， 以利 的孫子。 以利 從前在 示羅 作耶和華的祭司。 約拿單 去了，百姓卻不知道。
1SAM|14|4|約拿單 要從隘口過到 非利士 駐軍那裏去。這隘口兩邊各有一座齒狀峭壁：一座名叫 播薛 ，另一座名叫 西尼 ；
1SAM|14|5|一座向北，對著 密抹 ，一座向南，對著 迦巴 。
1SAM|14|6|約拿單 對拿兵器的青年說：「來，我們過去到那些未受割禮之人的駐軍那裏，或者耶和華為我們施展能力，因為耶和華使人得勝，不在乎人多人少 。」
1SAM|14|7|拿兵器的對他說：「隨你的心意做吧。你上去，看哪，我一定跟隨你，與你同心。」
1SAM|14|8|約拿單 說：「看哪，我們要過去到那些人那裏，在他們那裏展現我們自己。
1SAM|14|9|他們若對我們這麼說：『站住，等我們到你們那裏去』，我們就站在原地，不上他們那裏去；
1SAM|14|10|但他們若這麼說：『上到我們這裏來吧』，我們就上去，因為耶和華把他們交在我們手裏了。這就是我們的憑據。」
1SAM|14|11|二人就讓 非利士 的駐軍看見。 非利士 人說：「看哪， 希伯來 人從躲藏的洞穴裏出來了！」
1SAM|14|12|站崗的士兵對 約拿單 和拿兵器的人說：「上到這裏來，我們有一件事要告訴你們。」 約拿單 就對拿兵器的人說：「跟我上去，因為耶和華把他們交在 以色列 人手裏了。」
1SAM|14|13|約拿單 手腳並用爬上去，拿兵器的人跟隨他。 非利士 人仆倒在 約拿單 面前，拿兵器的人跟著他，殺死他們。
1SAM|14|14|約拿單 和拿兵器的人第一次擊殺的約有二十人，都在一畝 地的半犁溝之內。
1SAM|14|15|於是在軍營、在田野、在眾百姓中，人心惶惶，駐軍和突擊隊都戰兢；地也震動，這是從上帝那裏來的驚恐 。
1SAM|14|16|在 便雅憫 的 基比亞 ， 掃羅 的哨兵觀看，看哪， 非利士 全軍潰亂，四處亂竄。
1SAM|14|17|掃羅 就對跟隨他的百姓說：「你們去數點人數，看是誰從我們這裏出去。」他們一數點，看哪， 約拿單 和拿兵器的人不在其中。
1SAM|14|18|那時上帝的約櫃 在 以色列 人那裏。 掃羅 對 亞希亞 說：「你把上帝的約櫃請到這裏來。」
1SAM|14|19|掃羅 正與祭司說話的時候， 非利士 營中的騷亂越來越劇烈； 掃羅 就對祭司說：「停手吧！」
1SAM|14|20|掃羅 和所有跟隨他的百姓都集合，來到戰場，看哪， 非利士 人用刀互相擊殺，大大混亂。
1SAM|14|21|那先前由四方來跟隨 非利士 人、在他們營中的 希伯來 人，現在也轉過來幫助跟隨 掃羅 和 約拿單 的 以色列 人了。
1SAM|14|22|那藏在 以法蓮 山區的 以色列 眾人聽說 非利士 人逃跑，就出來緊緊地追擊他們。
1SAM|14|23|那日，耶和華使 以色列 人得勝，戰爭一直打到 伯‧亞文 。
1SAM|14|24|那日， 以色列 人非常困憊，因為 掃羅 叫百姓起誓說：「凡不等到晚上我向敵人報完了仇就吃東西的，必受詛咒。」因此所有的百姓都沒有嘗食物。
1SAM|14|25|所有的百姓 進入樹林，見地面上有蜜。
1SAM|14|26|百姓進了樹林，看哪，有蜜流出來，卻沒有人敢用手取蜜入口，因為百姓怕那誓言。
1SAM|14|27|約拿單 沒有聽見他父親叫百姓起誓，所以他伸出手中的杖，以杖頭蘸在蜂房裏，用手取回送入口內，他的眼睛就明亮了。
1SAM|14|28|百姓中有一人對他說：「你父親曾叫百姓嚴嚴地起誓說，今日吃東西的人必受詛咒；因此百姓就疲乏了。」
1SAM|14|29|約拿單 說：「我父親給這地添麻煩了。你們看，我嘗了這一點蜜，眼睛就明亮了。
1SAM|14|30|今日百姓若隨意吃了從仇敵奪來的東西，現在擊殺的 非利士 人豈不更多嗎？」
1SAM|14|31|這日， 以色列 人擊殺 非利士 人，從 密抹 直到 亞雅崙 。但百姓非常疲乏，
1SAM|14|32|就急著撲向掠物，奪取牛羊和牛犢，宰於地上，連肉帶血吃了。
1SAM|14|33|有人告訴 掃羅 說：「看哪，百姓吃帶血的肉，得罪耶和華了。」 掃羅 說：「你們行了詭詐，今日把一塊大石頭滾到我這裏來吧。」
1SAM|14|34|掃羅 又說：「你們分散到百姓中，對他們說，你們各人把牛羊牽到我這裏來宰了吃，不可吃帶血的肉得罪耶和華。」那夜，所有的百姓把自己手中的牛 牽到那裏宰了。
1SAM|14|35|掃羅 為耶和華築了一座壇，這是他開始為耶和華築的壇。
1SAM|14|36|掃羅 說：「我們要在夜裏下去追趕 非利士 人，搶掠他們，直到天亮，不給他們留下一人。」眾百姓說：「你看怎樣好就做吧！」祭司說：「我們要先在這裏親近上帝。」
1SAM|14|37|掃羅 求問上帝說：「我可以下去追趕 非利士 人嗎？你把他們交在 以色列 人手裏嗎？」這日上帝沒有回答他。
1SAM|14|38|掃羅 說：「百姓中的眾領袖，你們都要近前來到這裏，查明今日這罪是怎樣發生的。
1SAM|14|39|我指著拯救 以色列 的永生的耶和華起誓，就是我兒子 約拿單 犯了罪，他也必被處死。」但眾百姓中無人回答他。
1SAM|14|40|掃羅 對 以色列 眾人說：「你們站在一邊，我與我兒子 約拿單 也站在一邊。」百姓對 掃羅 說：「你看怎樣好就做吧！」
1SAM|14|41|掃羅 向耶和華－ 以色列 的上帝禱告說：「求你指示正確的答案。」抽中的是 掃羅 和 約拿單 ，百姓盡都無事。
1SAM|14|42|掃羅 說：「你們再抽籤，看是我，還是我兒子 約拿單 。」抽中的是 約拿單 。
1SAM|14|43|掃羅 對 約拿單 說：「你告訴我，你做了甚麼事？」 約拿單 說：「我只是用手中的杖，以杖頭蘸了一點蜜嘗嘗，看哪，我就要死嗎？」
1SAM|14|44|掃羅 說：「 約拿單 哪，你一定要死！若不然，願上帝重重懲罰我。」
1SAM|14|45|百姓對 掃羅 說：「 約拿單 在 以色列 中大行拯救，豈可死呢？絕對不可！我們指著永生的耶和華起誓，連他的一根頭髮也不可落地，因為他今日與上帝一同做事。」於是百姓救 約拿單 免了死亡。
1SAM|14|46|掃羅 上去，不追趕 非利士 人， 非利士 人也回本地去了。
1SAM|14|47|掃羅 執掌 以色列 的國權，攻打他四圍所有的仇敵，就是 摩押 人、 亞捫 人、 以東 人和 瑣巴 諸王，以及 非利士 人。他無論往何處去，都打敗他們。
1SAM|14|48|掃羅 奮勇作戰，擊敗 亞瑪力 人，救了 以色列 脫離搶掠他們之人的手。
1SAM|14|49|掃羅 的兒子是 約拿單 、 亦施韋 、 麥基‧舒亞 。他的兩個女兒：長女名叫 米拉 ，次女名叫 米甲 。
1SAM|14|50|掃羅 的妻子名叫 亞希暖 ，是 亞希瑪斯 的女兒。 掃羅 軍隊的元帥名叫 押尼珥 ，是 掃羅 的叔叔 尼珥 的兒子。
1SAM|14|51|掃羅 的父親 基士 ， 押尼珥 的父親 尼珥 ，都是 亞別 的兒子。
1SAM|14|52|掃羅 有生之年常與 非利士 人激烈爭戰，他看到任何有能力的人或勇士，都招募來跟隨他。
1SAM|15|1|撒母耳 對 掃羅 說：「耶和華差遣我膏你為王，治理他的百姓 以色列 ，現在你要聽從耶和華的話。
1SAM|15|2|萬軍之耶和華如此說：『 以色列 人從 埃及 上來的時候，在路上 亞瑪力 人怎樣待他們，怎樣抵擋他們，我都要懲罰。
1SAM|15|3|現在你要去攻打 亞瑪力 人，滅盡他們所有的，不可憐惜他們，將男女、孩童、吃奶的，以及牛、羊、駱駝和驢全都殺死。』」
1SAM|15|4|於是 掃羅 在 提拉因 召集百姓，數點他們，共有二十萬步兵和一萬 猶大 人。
1SAM|15|5|掃羅 到了 亞瑪力 的京城，在谷中設下埋伏。
1SAM|15|6|掃羅 對 基尼 人說：「你們離開 亞瑪力 人下去吧，免得我把你們和 亞瑪力 人一同殺滅，因為 以色列 眾人從 埃及 上來的時候，你們曾恩待他們。」於是 基尼 人離開了 亞瑪力 人。
1SAM|15|7|掃羅 攻打 亞瑪力 人，從 哈腓拉 直到 埃及 東邊的 書珥 ，
1SAM|15|8|生擒了 亞瑪力 王 亞甲 ，用刀殺盡 亞瑪力 的眾百姓。
1SAM|15|9|掃羅 和百姓卻憐惜 亞甲 ，愛惜上好的牛、羊、牛犢、羔羊，以及一切美物，不肯滅絕。但是凡看不上眼和沒有價值的，他們盡都殺了。
1SAM|15|10|耶和華的話臨到 撒母耳 說：
1SAM|15|11|「我立 掃羅 為王，我感到遺憾，因為他轉去不跟從我，不遵守我的命令。」 撒母耳 就很生氣，終夜哀求耶和華。
1SAM|15|12|撒母耳 清早起來，去見 掃羅 。有人告訴 撒母耳 說：「 掃羅 到了 迦密 ，看哪，他在那裏為自己立了紀念碑，又轉身下到 吉甲 。」
1SAM|15|13|撒母耳 到了 掃羅 那裏， 掃羅 對他說：「願耶和華賜福給你，耶和華的命令我已遵守了。」
1SAM|15|14|撒母耳 說：「我耳中聽見有羊叫、牛鳴的聲音，又是甚麼呢？」
1SAM|15|15|掃羅 說：「這是百姓從 亞瑪力 人那裏帶來的，因為他們愛惜上好的牛羊，要獻給耶和華－你的上帝。其餘的，我們都滅盡了。」
1SAM|15|16|撒母耳 對 掃羅 說：「住口吧！等我把耶和華昨夜向我所說的話告訴你。」 掃羅 說：「請說。」
1SAM|15|17|撒母耳 說：「你雖然看自己為小，你豈不是作了 以色列 諸支派的元首嗎？耶和華膏你作了 以色列 的王。
1SAM|15|18|耶和華差遣你，吩咐你說：『你去除滅那些犯罪的 亞瑪力 人，攻打他們，直到把他們完全滅盡。』
1SAM|15|19|你為何沒有聽從耶和華的話呢？你為何急著撲向掠物，行耶和華眼中看為惡的事呢？」
1SAM|15|20|掃羅 對 撒母耳 說：「我聽從了耶和華的話，行了耶和華派我行的路，擒了 亞瑪力 王 亞甲 來，滅盡了 亞瑪力 人。
1SAM|15|21|百姓卻從掠物中取了牛羊，是當滅之物中最好的，要在 吉甲 獻給耶和華－你的上帝。」
1SAM|15|22|撒母耳 說： 「耶和華喜愛燔祭和祭物， 豈如喜愛人聽從他的話呢？ 看哪，聽命勝於獻祭， 順從勝於公羊的脂肪。
1SAM|15|23|悖逆與占卜的罪相等， 頑梗與拜偶像的罪孽相同。 因為你厭棄耶和華的命令， 耶和華也厭棄你作王。」
1SAM|15|24|掃羅 對 撒母耳 說：「我有罪了！我違背了耶和華的指示和你的命令；因為我懼怕百姓，聽從了他們的話。
1SAM|15|25|現在求你赦免我的罪，同我回去，我好敬拜耶和華。」
1SAM|15|26|撒母耳 對 掃羅 說：「我不同你回去，因為你厭棄耶和華的命令，耶和華也厭棄你作 以色列 的王。」
1SAM|15|27|撒母耳 轉身要走， 掃羅 抓住他外袍的衣角，外袍就斷裂了。
1SAM|15|28|撒母耳 對他說：「今日耶和華使 以色列 國與你斷絕，把這國賜給另一個比你更好的人。
1SAM|15|29|以色列 的大能者必不說謊，也不後悔，因為他不是世人，絕不後悔。」
1SAM|15|30|掃羅 說：「我有罪了。現在求你在我百姓的長老和 以色列 人面前尊重我，同我回去，我好敬拜耶和華－你的上帝。」
1SAM|15|31|於是 撒母耳 轉身跟隨 掃羅 回去， 掃羅 就敬拜耶和華。
1SAM|15|32|撒母耳 說：「把 亞瑪力 王 亞甲 帶到我這裏來。」 亞甲 就歡歡喜喜地來到他面前，說：「死亡的苦難必定過去了。」
1SAM|15|33|撒母耳 說：「你既用刀使婦人喪子，你母親在婦人中也必照樣喪子。」於是， 撒母耳 在 吉甲 耶和華面前把 亞甲 砍碎了。
1SAM|15|34|撒母耳 回了 拉瑪 。 掃羅 上他所住的 基比亞 ，回自己的家去了。
1SAM|15|35|撒母耳 直到死的日子，再沒有見 掃羅 。但 撒母耳 為 掃羅 悲傷，因為耶和華遺憾立 掃羅 為 以色列 的王。
1SAM|16|1|耶和華對 撒母耳 說：「我既厭棄 掃羅 作 以色列 的王，你為他悲傷要到幾時呢？你將膏油盛滿了角；來，我差遣你到 伯利恆 人 耶西 那裏去，因為我在他兒子中已看中了一個為我作王的。」
1SAM|16|2|撒母耳 說：「我怎麼能去呢？ 掃羅 一聽見，就會殺我。」耶和華說：「你可以手裏牽一頭小母牛去，說：『我來是要向耶和華獻祭。』
1SAM|16|3|你要請 耶西 來一同獻祭，我會指示你當做的事。我對你說的那個人，你要為我膏他。」
1SAM|16|4|撒母耳 遵照耶和華的話去做，來到 伯利恆 ，城裏的長老都戰戰兢兢出來迎接他，有人問他說：「你是為平安來的嗎？」
1SAM|16|5|他說：「為平安來的，我來是要向耶和華獻祭。你們要使自己分別為聖，來跟我一同獻祭。」 撒母耳 把 耶西 和他眾兒子分別為聖，請他們來一同獻祭。
1SAM|16|6|他們來的時候， 撒母耳 看見 以利押 ，就心裏說，耶和華的受膏者一定在耶和華面前了。
1SAM|16|7|耶和華卻對 撒母耳 說：「不要只看他的外貌和他身材高大，我不揀選他。因為耶和華不像人看人，人是看外貌 ，耶和華是看內心。」
1SAM|16|8|耶西 叫 亞比拿達 從 撒母耳 面前經過， 撒母耳 說：「耶和華也不揀選他。」
1SAM|16|9|耶西 又叫 沙瑪 經過， 撒母耳 說：「耶和華也不揀選他。」
1SAM|16|10|耶西 叫他七個兒子都從 撒母耳 面前經過， 撒母耳 對 耶西 說：「這些都不是耶和華所揀選的。」
1SAM|16|11|撒母耳 對 耶西 說：「你的兒子都在這裏了嗎？」他說：「還有一個最小的，看哪，他正在放羊。」 撒母耳 對 耶西 說：「你派人去叫他來；他若不來這裏，我們必不坐席。」
1SAM|16|12|耶西 就派人去叫他來。他面色紅潤，雙目清秀，容貌俊美。耶和華說：「起來，膏他，因為這就是他了。」
1SAM|16|13|撒母耳 就用角裏的膏油，在他的兄長中膏了他。從這日起，耶和華的靈就大大感動 大衛 。 撒母耳 起身回 拉瑪 去了。
1SAM|16|14|耶和華的靈離開 掃羅 ，有邪靈從耶和華那裏來擾亂他。
1SAM|16|15|掃羅 的臣僕對他說：「看哪，有邪靈從上帝那裏來擾亂你。
1SAM|16|16|我們的主可以吩咐你面前的臣僕，去找一個善於彈琴的來。上帝那裏來的邪靈臨到你身上的時候，他用手彈琴，你就會感覺爽快。」
1SAM|16|17|掃羅 對臣僕說：「你們給我找一個善於彈琴的，帶到我這裏來。」
1SAM|16|18|僕人中有一個回答說：「看哪，我曾見 伯利恆 人 耶西 的一個兒子善於彈琴，是大能的勇士，說話合宜，容貌俊美，耶和華也與他同在。」
1SAM|16|19|於是 掃羅 差遣使者到 耶西 那裏，說：「叫你放羊的兒子 大衛 到我這裏來。」
1SAM|16|20|耶西 把幾個餅和一皮袋酒，以及一隻小山羊，馱在驢上，由兒子 大衛 的手送給 掃羅 。
1SAM|16|21|大衛 到了 掃羅 那裏，就侍立在 掃羅 面前。 掃羅 很喜歡他，他就作了 掃羅 拿兵器的人。
1SAM|16|22|掃羅 派人到 耶西 那裏，說：「讓 大衛 侍立在我面前，因為他在我眼前蒙了恩寵。」
1SAM|16|23|從上帝那裏來的邪靈臨到 掃羅 身上的時候， 大衛 就拿琴，用手彈奏，使 掃羅 舒暢，感覺爽快，那邪靈就離開他了。
1SAM|17|1|非利士 人召集他們的軍隊來爭戰。他們聚集在 猶大 的 梭哥 ，在 梭哥 和 亞西加 中間的 以弗‧大憫 安營。
1SAM|17|2|掃羅 和 以色列 人也聚集，在 以拉谷 安營，擺陣迎戰，要與 非利士 人打仗。
1SAM|17|3|非利士 人站在這邊的山上， 以色列 人站在那邊的山上，當中有谷。
1SAM|17|4|從 非利士 營中出來一個挑戰的人，名叫 歌利亞 ，是 迦特 人，身高六肘一虎口。
1SAM|17|5|他頭戴銅盔，身穿鎧甲，甲重五千舍客勒銅。
1SAM|17|6|他腿上有銅護膝，兩肩之中背負銅矛。
1SAM|17|7|他的槍桿粗如織布機的軸，槍頭的鐵重六百舍客勒。有一個拿盾牌的人走在他前面。
1SAM|17|8|歌利亞 站著，對 以色列 的軍隊喊叫，對他們說：「你們出來擺陣作戰是為了甚麼呢？我不是 非利士 人嗎？你們不是 掃羅 的僕人嗎？你們選一個人出來，叫他下來到我這裏吧。
1SAM|17|9|他若能與我決鬥，把我殺死，我們就作你們的奴隸；我若勝了他，把他殺死，你們就作我們的奴隸，服事我們。」
1SAM|17|10|那 非利士 人又說：「我今日向 以色列 的軍隊罵陣。你們叫一個人出來，跟我決鬥吧。」
1SAM|17|11|掃羅 和 以色列 眾人聽見 非利士 人這些話就驚惶，非常害怕。
1SAM|17|12|大衛 是 猶大 伯利恆 的 以法他 人 耶西 的兒子， 耶西 有八個兒子。在 掃羅 的時候，這人年老，在眾人中受敬重 。
1SAM|17|13|耶西 最大的三個兒子跟隨 掃羅 出征。出征的三個兒子名字是：長子 以利押 ，次子 亞比拿達 ，三子 沙瑪 。
1SAM|17|14|大衛 是最小的，最大的三個兒子跟隨 掃羅 。
1SAM|17|15|大衛 有時離開 掃羅 ，回 伯利恆 為他父親放羊。
1SAM|17|16|那 非利士 人早晚都出來站著，共四十日。
1SAM|17|17|耶西 對他兒子 大衛 說：「你拿一伊法烘了的穗子和十個餅，跑到營裏去，交給你的哥哥，
1SAM|17|18|再拿這十塊奶餅，送給他們的千夫長，並要問你哥哥好，向他們要個憑據回來。」
1SAM|17|19|掃羅 和 大衛 的三個哥哥，以及 以色列 眾人，都在 以拉谷 與 非利士 人打仗。
1SAM|17|20|大衛 早晨起來，把羊交託一個看守的人，照 耶西 所吩咐的帶著食物去了。到了軍營，軍隊剛出到戰場，吶喊叫陣。
1SAM|17|21|以色列 人和 非利士 人都擺列陣勢，彼此相對。
1SAM|17|22|大衛 把東西留在看守物件的人手中，跑到戰場，問他哥哥好。
1SAM|17|23|他與他們說話的時候，看哪，那挑戰的人，就是 迦特 的 非利士 人 歌利亞 ，從 非利士 隊伍中上來，說了同樣的話， 大衛 聽見了。
1SAM|17|24|以色列 眾人看見那人就非常害怕，從他面前逃跑。
1SAM|17|25|以色列 人說：「這上來的人你看見了嗎？他上來是要向 以色列 人罵陣。若有人能殺他，王必賞賜他大財，將自己的女兒嫁給他，並在 以色列 人中免除他父家納糧服役。」
1SAM|17|26|大衛 對站在旁邊的人說：「若有人殺這 非利士 人，除掉 以色列 人的羞辱，他會怎樣呢？這未受割禮的 非利士 人是誰，竟敢向永生上帝的軍隊罵陣！」
1SAM|17|27|百姓照同樣的話對他說：「若有人殺了那人，必這樣待他。」
1SAM|17|28|大衛 的長兄 以利押 聽見 大衛 與他們所說的話，就向他發怒，說：「你下來做甚麼呢？在曠野的那幾隻羊，你交託誰了呢？我知道你的驕傲和你心裏的惡意，你下來只是為了看戰爭！」
1SAM|17|29|大衛 說：「我現在做了甚麼呢？只是問一句話也不可以嗎？」
1SAM|17|30|大衛 離開他轉向別人，問了同樣的事，百姓也照先前的話回答他。
1SAM|17|31|有人聽見 大衛 所說的話，就在 掃羅 面前報告； 掃羅 就派人叫他來。
1SAM|17|32|大衛 對 掃羅 說：「人不必因那 非利士 人灰心。你的僕人要去與他決鬥。」
1SAM|17|33|掃羅 對 大衛 說：「你不能去與那 非利士 人決鬥，因為你年紀太輕，他從小就是戰士。」
1SAM|17|34|大衛 對 掃羅 說：「你僕人為父親放羊，有時獅子來了，有時熊來了，從群中抓走一隻羔羊。
1SAM|17|35|我就追趕牠，擊打牠，把羔羊從牠口中救出來。牠起來攻擊我，我就揪牠的鬍子，打死牠。
1SAM|17|36|你僕人曾打死獅子和熊，這未受割禮的 非利士 人必像獅子和熊一樣，因為他向永生上帝的軍隊罵陣。」
1SAM|17|37|大衛 又說：「耶和華救我脫離獅子和熊的爪，他必救我脫離這 非利士 人的手。」 掃羅 對 大衛 說：「你去吧！耶和華必與你同在。」
1SAM|17|38|掃羅 把自己的戰衣給 大衛 穿上，將銅盔戴在他頭上，又給他穿上鎧甲。
1SAM|17|39|大衛 佩刀在戰衣上，試著走走看。因 大衛 沒有試過，就對 掃羅 說：「我穿戴這些不能走路，因為我沒有試過。」於是他脫下身上的這些軍裝。
1SAM|17|40|他手中拿杖，又在溪中挑選了五塊光滑的石子，放在袋裏，就是牧人帶的囊裏，手裏拿著甩石的機弦，迎向那 非利士 人。
1SAM|17|41|那 非利士 人漸漸走近 大衛 ，拿盾牌的人在他前面。
1SAM|17|42|非利士 人觀看，見了 大衛 ，就藐視他，因為他年輕，面色紅潤，容貌俊美。
1SAM|17|43|非利士 人對 大衛 說：「你拿著杖到我這裏來，我豈是狗嗎？」 非利士 人就指著自己的神明詛咒 大衛 。
1SAM|17|44|非利士 人又對 大衛 說：「來吧！我要把你的肉給空中的飛鳥和田野的走獸。」
1SAM|17|45|大衛 對 非利士 人說：「你來攻擊我，是靠著刀槍和銅矛，但我來攻擊你，是靠著萬軍之耶和華的名，就是你所辱罵、帶領 以色列 軍隊的上帝。
1SAM|17|46|今日耶和華必將你交在我手裏。我必殺你，砍下你的頭，今日我要把 非利士 軍兵的屍體給空中的飛鳥和地上的野獸，使全地的人都知道以色列中有上帝，
1SAM|17|47|又使這裏的全會眾知道，耶和華使人得勝，不是用刀用槍，因為戰爭全在乎耶和華。他必將你們交在我們手裏。」
1SAM|17|48|那 非利士 人起來，迎向 大衛 ，走近前來。 大衛 急忙往戰場，迎向 非利士 人跑去。
1SAM|17|49|大衛 伸手入囊中，從裏面掏出一塊石子來，用機弦甩去，擊中 非利士 人的前額，石子進入額內，他就仆倒，面伏於地。
1SAM|17|50|這樣， 大衛 用機弦和石子勝了那 非利士 人，擊中了他，把他殺死； 大衛 手中沒有刀。
1SAM|17|51|大衛 跑去，站在那 非利士 人身旁，把他的刀從鞘中拔出來，殺死他，用刀割下他的頭。 非利士 眾人看見他們的勇士死了，就都逃跑。
1SAM|17|52|以色列 人和 猶大 人就起來吶喊，追趕 非利士 人，直到 該 和 以革倫 的城門。被殺的 非利士 人倒在路上，從 沙拉音 直到 迦特 和 以革倫 。
1SAM|17|53|以色列 人追趕 非利士 人回來，搶奪了他們的軍營。
1SAM|17|54|大衛 拿著那 非利士 人的頭帶到 耶路撒冷 ，卻把那 非利士 人的軍裝放在自己的帳棚裏。
1SAM|17|55|掃羅 看見 大衛 去迎戰 非利士 人，就問 押尼珥 元帥說：「 押尼珥 ，那年輕人是誰的兒子？」 押尼珥 說：「王啊，我在你面前起誓，我不知道。」
1SAM|17|56|王說：「你可以問問那孩子是誰的兒子。」
1SAM|17|57|大衛 打死那 非利士 人回來， 押尼珥 領他到 掃羅 面前， 大衛 手中拿著 非利士 人的頭。
1SAM|17|58|掃羅 問他說：「年輕人，你是誰的兒子？」 大衛 說：「我是你僕人 伯利恆 人 耶西 的兒子。」
1SAM|18|1|大衛 對 掃羅 說完了話， 約拿單 的心與 大衛 的心深相契合。 約拿單 愛 大衛 ，如同愛自己的性命。
1SAM|18|2|那日 掃羅 留住 大衛 ，不讓他回父家。
1SAM|18|3|約拿單 愛 大衛 如同愛自己的性命，就與他立約。
1SAM|18|4|約拿單 從身上脫下外袍，給了 大衛 ，又把戰衣、刀、弓、腰帶都給了他。
1SAM|18|5|掃羅 無論差遣 大衛 往何處去，他都做事精明。 掃羅 立他作軍隊的指揮官，眾百姓和 掃羅 的臣僕都看為美。
1SAM|18|6|大衛 打死了那 非利士 人，同眾人回來的時候，婦女們從 以色列 各城裏出來，歡歡喜喜，打鼓奏樂，唱歌跳舞，迎接 掃羅 王。
1SAM|18|7|眾婦女歡樂唱和，說： 「 掃羅 殺死千千， 大衛 殺死萬萬。」
1SAM|18|8|掃羅 非常憤怒，不喜歡這話。他說：「將萬萬歸給 大衛 ，千千歸給我，只剩下王國沒有給他！」
1SAM|18|9|從這日起， 掃羅 就敵視 大衛 。
1SAM|18|10|次日，從上帝來的邪靈緊抓住 掃羅 ，他就在家中胡言亂語。 大衛 照常彈琴， 掃羅 手裏拿著槍。
1SAM|18|11|掃羅 把槍一擲，心裏說：「我要將 大衛 刺透，釘在牆上。」 大衛 閃避了他兩次。
1SAM|18|12|掃羅 懼怕 大衛 ，因為耶和華離開自己，與 大衛 同在。
1SAM|18|13|所以 掃羅 叫 大衛 離開自己，立他為千夫長，他就領兵出入。
1SAM|18|14|大衛 所做的每一件事都精明，耶和華也與他同在。
1SAM|18|15|掃羅 見 大衛 做事精明，就更怕他。
1SAM|18|16|但 以色列 和 猶大 眾人都愛 大衛 ，因為他領他們出入。
1SAM|18|17|掃羅 對 大衛 說：「看哪，我將大女兒 米拉 嫁給你，只要你作我的勇士，為耶和華爭戰。」 掃羅 心裏說：「我不好親手害他，要藉 非利士 人的手害他。」
1SAM|18|18|大衛 對 掃羅 說：「我是誰，我是甚麼出身，我父家在 以色列 中算甚麼，豈敢作王的女婿呢？」
1SAM|18|19|掃羅 的女兒 米拉 到了當嫁給 大衛 的時候， 掃羅 卻將她嫁給了 米何拉 人 亞得列 。
1SAM|18|20|掃羅 的女兒 米甲 愛 大衛 。有人告訴 掃羅 ，這件事在 掃羅 眼中看為合宜。
1SAM|18|21|掃羅 心裏說：「我把這女兒嫁給 大衛 ，作他的圈套，好藉 非利士 人的手害他。」所以 掃羅 第二次對 大衛 說：「你今日可以作我的女婿。」
1SAM|18|22|掃羅 吩咐臣僕：「你們暗中對 大衛 說：『看哪，王喜歡你，王的臣僕也都愛戴你，現在你就作王的女婿吧。』」
1SAM|18|23|掃羅 的臣僕照這話說給 大衛 聽。 大衛 說：「你們把作王的女婿看為小事嗎？我是貧窮卑微的人。」
1SAM|18|24|掃羅 的臣僕回奏說， 大衛 說了這樣的話。
1SAM|18|25|掃羅 說：「你們要對 大衛 這樣說：『王不要甚麼聘禮，只要一百 非利士 人的包皮，好在王的仇敵身上報仇。』」 掃羅 的意圖是要 大衛 落在 非利士 人的手中。
1SAM|18|26|掃羅 的臣僕把這話告訴 大衛 ， 大衛 就歡喜作王的女婿。日期還沒有到，
1SAM|18|27|大衛 和跟隨他的人起來前往，殺了二百 非利士 人，將包皮足數交給王，為要作王的女婿。於是 掃羅 將女兒 米甲 嫁給 大衛 。
1SAM|18|28|掃羅 見耶和華與 大衛 同在，女兒 米甲 又愛 大衛 ，
1SAM|18|29|就更怕 大衛 ，常常與 大衛 為敵。
1SAM|18|30|每逢 非利士 的軍官出來打仗， 大衛 做事比 掃羅 任何臣僕更精明，因此他的名極受尊重。
1SAM|19|1|掃羅 吩咐他兒子 約拿單 和眾臣僕要殺 大衛 ，但 掃羅 的兒子 約拿單 卻很喜愛 大衛 。
1SAM|19|2|約拿單 告訴 大衛 說：「我父 掃羅 想要殺你，現在你要小心，明日早晨留在一個僻靜的地方藏起來。
1SAM|19|3|我會出去，到你所藏的田裏，站在我父親旁邊，與父親談論到你。我看情形怎樣，會告訴你。」
1SAM|19|4|約拿單 向他父親 掃羅 說 大衛 的好話，對他說：「王不可得罪王的僕人 大衛 ，因為他未曾得罪你，他所行的對你都很有益處。
1SAM|19|5|他拚了命殺那 非利士 人，並且耶和華為全 以色列 大施拯救。那時你看見，也很歡喜，現在為何要犯罪，流無辜人的血，無緣無故殺 大衛 呢？」
1SAM|19|6|掃羅 聽了 約拿單 的話，就指著永生的耶和華起誓：「我絕不殺他。」
1SAM|19|7|約拿單 叫 大衛 來，把這一切事告訴他。 約拿單 帶他去見 掃羅 ，他就像以前一樣侍立在 掃羅 面前。
1SAM|19|8|此後又有戰爭， 大衛 出去與 非利士 人打仗。他大大擊敗他們，他們就在他面前逃跑。
1SAM|19|9|從耶和華來的邪靈又降在 掃羅 身上， 掃羅 手裏拿槍坐在屋裏， 大衛 正用手彈琴。
1SAM|19|10|掃羅 想要用槍刺透 大衛 ，把他釘在牆上，他卻躲開 掃羅 ， 掃羅 的槍刺入牆內。當夜 大衛 逃走，躲起來了。
1SAM|19|11|掃羅 派一些使者到 大衛 的房屋那裏守著他，等到天亮要殺他。 大衛 的妻子 米甲 對 大衛 說：「你今夜若不逃命，明日就要被殺。」
1SAM|19|12|於是 米甲 將 大衛 從窗戶縋下去，讓他走； 大衛 就逃走，躲起來了。
1SAM|19|13|米甲 把家中的神像放在床上，頭枕在山羊毛的枕頭上，用衣服蓋起來。
1SAM|19|14|掃羅 派一些使者去捉拿 大衛 ， 米甲 說：「他病了。」
1SAM|19|15|掃羅 又派一些使者去看 大衛 ，說：「把他連床一起抬到我這裏，我好殺他。」
1SAM|19|16|使者進去，看哪，神像在床上，頭枕在山羊毛的枕頭上。
1SAM|19|17|掃羅 對 米甲 說：「你為甚麼這樣欺騙我，放我仇敵逃走呢？」 米甲 對 掃羅 說：「他對我說：『你放我走吧，我何必要殺你呢？』」
1SAM|19|18|大衛 逃跑躲避，來到 拉瑪 的 撒母耳 那裏，把 掃羅 向他所行的事全告訴他。他和 撒母耳 就去，住在 拿約 。
1SAM|19|19|有人告訴 掃羅 說：「看哪， 大衛 在 拉瑪 的 拿約 」。
1SAM|19|20|掃羅 派一些使者去捉拿 大衛 。去的人見一隊先知受感說話， 撒母耳 站在當中領導他們， 掃羅 派去的使者也受上帝的靈感動說話。
1SAM|19|21|有人把這事告訴 掃羅 ，他又派另一些使者去，他們也受感說話。 掃羅 第三次派使者去，他們也受感說話。
1SAM|19|22|然後 掃羅 親自往 拉瑪 去，到了 西沽 的大井，問人說：「 撒母耳 和 大衛 在哪裏？」有人說：「看哪，在 拉瑪 的 拿約 。」
1SAM|19|23|他就往那裏去，到了 拉瑪 的 拿約 。上帝的靈也臨到他，他一面走一面受感說話，直到 拉瑪 的 拿約 。
1SAM|19|24|他也脫了衣服，也在 撒母耳 面前受感說話，一日一夜赤身躺臥。因此有人說：「 掃羅 也在先知中嗎？」
1SAM|20|1|大衛 從 拉瑪 的 拿約 逃跑，來到 約拿單 面前，對他說：「我做了甚麼，有甚麼罪孽，在你父親面前犯了甚麼罪，他竟要尋索我的性命呢？」
1SAM|20|2|約拿單 對他說：「絕無此事！你必不至於死。看哪，我父做事，無論大小，沒有不告訴我的。我父親為甚麼要隱瞞我這件事呢？不會這樣的！」
1SAM|20|3|大衛 又起誓說：「你父親確實知道我在你眼前蒙恩。所以他說，『這事不要讓 約拿單 知道，免得他愁煩。』我指著永生的耶和華起誓，又指著你的性命起誓，我離死只差一步而已。」
1SAM|20|4|約拿單 對 大衛 說：「你心裏所求的，我必為你成就。」
1SAM|20|5|大衛 對 約拿單 說：「看哪，明日是初一，我必須與王同席用餐，求你讓我去藏在田野，直到第三日傍晚。
1SAM|20|6|你父親若見我不在席上，你就說：『 大衛 懇求我允許他趕回本城 伯利恆 去，因為他全家在那裏獻年祭。』
1SAM|20|7|你父親若說好，你的僕人就平安了；他若大怒，你就知道他決意行惡。
1SAM|20|8|求你施恩於僕人，因你在耶和華面前曾與僕人立約。我若有罪孽，你就親自殺死我，何必把我交給你父親呢？」
1SAM|20|9|約拿單 說：「絕無此事！我若確實知道我父親決意害你，怎麼會不告訴你呢？」
1SAM|20|10|大衛 對 約拿單 說：「你父親若嚴厲回答你，誰來告訴我呢？」
1SAM|20|11|約拿單 對 大衛 說：「來，讓我們到田野去。」二人就往田野去了。
1SAM|20|12|約拿單 對 大衛 說：「願耶和華－ 以色列 的上帝作證。明日約在這時候，或第三日，我一探出我父親的心意，看哪，若對 大衛 是好意，我怎麼會不派人來告訴你呢？
1SAM|20|13|我父親若有意害你，而我不告訴你，送你平安地離開，願耶和華重重懲罰 約拿單 。願耶和華與你同在，如同從前與我父親同在一樣。
1SAM|20|14|你要照耶和華的慈愛恩待我，不但我活著的時候免我死亡，
1SAM|20|15|就是耶和華從地面逐一剪除 大衛 仇敵的時候，你也永不可向我家斷絕恩惠。」
1SAM|20|16|於是 約拿單 與 大衛 家立約：「願耶和華從 大衛 仇敵 的手來追討。」
1SAM|20|17|約拿單 因愛 大衛 如同愛自己的性命，就叫他再起誓。
1SAM|20|18|約拿單 對他說：「明日是初一，你的座位空著，人必察覺你不在。
1SAM|20|19|到第三日，就要走一段長路下去 ，去到你遇事那天所藏的地方，在 以色 磐石 的旁邊等候。
1SAM|20|20|我會向磐石旁邊射三箭，如同射箭靶一樣。
1SAM|20|21|看哪，我會派僮僕，說：『去把箭找來。』我若對僮僕喊說：『看哪，箭在你的這邊，把箭拿來』，你就可以平安回來；我指著永生的耶和華起誓，你一定沒有事。
1SAM|20|22|我若對孩子說：『看哪，箭在你的前方』，你就要離開，因為是耶和華差你去的。
1SAM|20|23|至於你和我，我們所說的話，看哪，耶和華在你我中間作證，直到永遠。」
1SAM|20|24|大衛 就去藏在田野。到了初一，王要坐席用餐。
1SAM|20|25|王照常坐在靠牆的位子上， 約拿單 在對面 ， 押尼珥 坐在 掃羅 旁邊， 大衛 的座位卻是空的。
1SAM|20|26|這日 掃羅 沒有說甚麼，因為他說：「 大衛 或許有事，偶染不潔，還未得潔淨。」
1SAM|20|27|初二， 大衛 的座位還空著。 掃羅 對他兒子 約拿單 說：「 耶西 的兒子為何昨日、今日都沒有來用餐呢？」
1SAM|20|28|約拿單 回答 掃羅 說：「 大衛 懇求我允許他回 伯利恆 去，
1SAM|20|29|說：『求你讓我去，因為我家在城裏有獻祭的事，我哥哥吩咐我去。如今我若在你眼前蒙恩，求你讓我去見我的兄弟。』所以 大衛 沒有來赴王的筵席。」
1SAM|20|30|掃羅 向 約拿單 怒氣大發，對他說：「你這頑梗悖逆之婦人所生的，我怎麼會不知道你選擇 耶西 的兒子 ，自取羞辱，也使你母親露體蒙羞呢？
1SAM|20|31|只要 耶西 的兒子還活在世上一天，你和你的國必保不住。現在你要派人去，把他帶到我這裏來，因為他是該死的。」
1SAM|20|32|約拿單 回答父親 掃羅 說：「他為甚麼該死呢？他做了甚麼呢？」
1SAM|20|33|掃羅 向 約拿單 擲槍要刺他， 約拿單 就知道他父親決意要殺死 大衛 。
1SAM|20|34|於是 約拿單 氣憤憤地從席上起來。他在初二這天沒有吃飯，因為他為 大衛 愁煩，又因為他父親羞辱了他。
1SAM|20|35|次日早晨， 約拿單 按著與 大衛 約定的時候到田野去，有一個小僮僕跟隨他。
1SAM|20|36|約拿單 對僮僕說：「你跑去把我所射的箭找來。」僮僕跑去， 約拿單 就把箭射在僮僕的前方。
1SAM|20|37|僮僕到了 約拿單 落箭之地， 約拿單 呼叫僮僕說：「箭不是在你的前方嗎？」
1SAM|20|38|約拿單 又呼叫僮僕說：「快去，不要站在那裏！」僮僕就撿起箭來，回到主人那裏。
1SAM|20|39|僮僕不知道這是甚麼意思，只有 約拿單 和 大衛 知道這事。
1SAM|20|40|約拿單 把他的弓箭交給僮僕，吩咐他說：「你拿到城裏去。」
1SAM|20|41|僮僕一去， 大衛 就從南邊 出來，俯伏在地，拜了三拜。他們彼此親吻，一起哭泣， 大衛 哭得更悲哀。
1SAM|20|42|約拿單 對 大衛 說：「你平平安安地去吧！因為我們二人曾指著耶和華的名起誓說：『願耶和華在你我中間，以及你我後裔中間作證，直到永遠。』」 大衛 就起身走了， 約拿單 也回城裏去了。
1SAM|21|1|大衛 到了 挪伯 的 亞希米勒 祭司那裏， 亞希米勒 戰戰兢兢地出來迎接他，對他說：「你為甚麼獨自一人，沒有人跟隨你呢？」
1SAM|21|2|大衛 對 亞希米勒 祭司說：「王吩咐我一件事，對我說：『我差遣你，吩咐你的這件事，不可讓任何人知道。』因此我已告訴一些僕人到某處去 。
1SAM|21|3|現在你手中有甚麼？請你給我五個餅或是可以找到的食物。」
1SAM|21|4|祭司對 大衛 說：「我手中沒有普通的餅，只有聖餅，只能給沒有親近婦人的年輕人。」
1SAM|21|5|大衛 回答祭司說：「我們確實沒有親近婦人，如同往常我出征的時候一樣。平常行路，僕人的身體 都還分別為聖，何況今日豈不更使自己分別為聖嗎？」
1SAM|21|6|祭司拿聖餅給他，因為在那裏沒有別的餅，只有那從耶和華面前撤下的供餅，就是換上熱餅的日子取下來的。
1SAM|21|7|當日，有 掃羅 的一個臣僕在那裏，他留在耶和華的面前，名叫 多益 ，是 以東 人，作 掃羅 的畜牧長。
1SAM|21|8|大衛 對 亞希米勒 說：「你手中有沒有槍或刀？因為王的事緊急，連刀劍兵器我都沒有帶。」
1SAM|21|9|祭司說：「你在 以拉谷 所殺的 非利士 人 歌利亞 的那刀，看哪，裹在布中，放在以弗得後邊。你若要可以拿去，除此以外，再沒有別的了。」 大衛 說：「沒有甚麼可以跟它比的了！請你給我。」
1SAM|21|10|那日 大衛 起來，躲避 掃羅 ，逃到 迦特 王 亞吉 那裏。
1SAM|21|11|亞吉 的臣僕對他說：「這不是那地的國王 大衛 嗎？那裏的人跳舞唱和： 『 掃羅 殺死千千， 大衛 殺死萬萬』， 不是指著他說的嗎？」
1SAM|21|12|大衛 把這些話放在心裏，就很懼怕 迦特 王 亞吉 。
1SAM|21|13|於是他在眾人眼前一反常態，在他們中間 裝瘋作癲，在城門的門扇上胡寫亂畫，任由唾沫流在鬍子上。
1SAM|21|14|亞吉 對臣僕說：「看哪，你們看這人瘋了，為甚麼帶他到我這裏來呢？
1SAM|21|15|我豈缺少瘋子，你們竟然帶這人到我面前瘋癲嗎？這個人可以進我的家嗎？」
1SAM|22|1|大衛 離開那裏，逃到 亞杜蘭 洞。他的兄弟和他父親全家聽見了，都下到他那裏去。
1SAM|22|2|凡生活窘迫的、欠債的、心裏苦惱的都聚集到 大衛 那裏，他就作他們的領袖，跟隨他的約有四百人。
1SAM|22|3|大衛 從那裏往 摩押 的 米斯巴 去，對 摩押 王說：「請你讓我父母搬來，跟你們在一起，等我知道上帝要為我怎樣做。」
1SAM|22|4|大衛 領他父母到 摩押 王面前。 大衛 住山寨一切的日子，他父母也都住在 摩押 王那裏。
1SAM|22|5|先知 迦得 對 大衛 說：「你不要住在山寨，要到 猶大 地去。」 大衛 就去，來到 哈列 的樹林。
1SAM|22|6|掃羅 聽見 大衛 和跟隨他之人的下落， 掃羅 正在 基比亞 ，坐在山頂 的柳樹下，手裏拿著槍，眾臣僕侍立在左右。
1SAM|22|7|掃羅 對左右侍立的臣僕說：「 便雅憫 人哪，聽著！ 耶西 的兒子也能把田地和葡萄園賜給你們各人嗎？他能立你們各人作千夫長和百夫長嗎？
1SAM|22|8|你們竟都結黨害我！我兒子與 耶西 的兒子立約的時候，無人告訴我；我兒子挑唆我的臣僕謀害我，像今日這樣，也無人告訴我，為我憂慮。」
1SAM|22|9|那時 以東 人 多益 站在 掃羅 的臣僕中，回答說：「我曾看見 耶西 的兒子往 挪伯 去，到了 亞希突 的兒子 亞希米勒 那裏。
1SAM|22|10|亞希米勒 為他求問耶和華，給他食物，又把 非利士 人 歌利亞 的刀給了他。」
1SAM|22|11|王就派人把 亞希突 的兒子 亞希米勒 祭司和他父親的全家，就是在 挪伯 的祭司都召了來，他們都來到王那裏。
1SAM|22|12|掃羅 說：「 亞希突 的兒子，聽著！」他說：「我主，我在這裏。」
1SAM|22|13|掃羅 對他說：「你為甚麼與 耶西 的兒子結黨害我，把食物和刀給他，又為他求問上帝，使他起來謀害我，像今日這樣？」
1SAM|22|14|亞希米勒 回答王說：「王的眾臣僕中有誰比 大衛 忠心呢？他是王的女婿，又是你的侍衛長 ，並且是你宮中受敬重的人。
1SAM|22|15|我今日才開始為他求問上帝嗎？絕非如此！王不要歸罪於我和我父全家，因為這事，無論大小，僕人都不知情。」
1SAM|22|16|王說：「 亞希米勒 ，你和你父全家都是該死的！」
1SAM|22|17|王吩咐左右的侍衛說：「你們轉身去殺耶和華的祭司吧！因為他們幫助 大衛 ，知道 大衛 逃跑卻不告訴我。」但王的臣僕都不願動手殺耶和華的祭司。
1SAM|22|18|王吩咐 多益 說：「你轉身去殺祭司吧！」 以東 人 多益 就轉身去殺祭司，那日殺了穿細麻布以弗得的，共八十五人，
1SAM|22|19|又用刀把祭司城 挪伯 中的男女、孩童和吃奶的都殺了，又用刀殺了牛、羊和驢子。
1SAM|22|20|亞希突 的兒子 亞希米勒 有一個兒子逃脫了；他名叫 亞比亞他 ，逃到 大衛 那裏。
1SAM|22|21|亞比亞他 把 掃羅 殺耶和華祭司的事告訴 大衛 。
1SAM|22|22|大衛 對 亞比亞他 說：「那日我見 以東 人 多益 在那裏，就知道他一定會告訴 掃羅 。你父的全家喪命，都是因我的緣故。
1SAM|22|23|你可以住在我這裏，不要懼怕。因為尋索你命的也要尋索我的命，你在我這裏可得保護。」
1SAM|23|1|有人告訴 大衛 說：「看哪， 非利士 人攻擊 基伊拉 ，搶奪禾場。」
1SAM|23|2|大衛 求問耶和華說：「我可以去嗎？我可以去攻打那些 非利士 人嗎？」耶和華對 大衛 說：「你可以去攻打 非利士 人，拯救 基伊拉 。」
1SAM|23|3|大衛 的人對他說：「看哪，我們在 猶大 這裏尚且懼怕，何況到 基伊拉 去攻打 非利士 人的軍隊呢？」
1SAM|23|4|大衛 又再求問耶和華，耶和華回答說：「你起身下 基伊拉 去，我必將 非利士 人交在你手裏。」
1SAM|23|5|於是 大衛 和他的人往 基伊拉 去，與 非利士 人打仗，大大擊敗他們，奪取他們的牲畜。這樣， 大衛 救了 基伊拉 的居民。
1SAM|23|6|亞希米勒 的兒子 亞比亞他 逃往 基伊拉 到 大衛 那裏的時候，手裏拿著以弗得。
1SAM|23|7|有人告訴 掃羅 ， 大衛 到了 基伊拉 。 掃羅 說：「上帝將他交在我手裏了，因為他進了有門有閂的城，把自己關起來了。」
1SAM|23|8|於是 掃羅 召集眾百姓，要下去攻打 基伊拉 ，圍困 大衛 和他的人。
1SAM|23|9|大衛 知道 掃羅 設計陷害他，就對 亞比亞他 祭司說：「把以弗得拿過來。」
1SAM|23|10|大衛 說：「耶和華－ 以色列 的上帝啊，你僕人確實聽見 掃羅 設法要到 基伊拉 來，為我的緣故毀滅這城。
1SAM|23|11|基伊拉 人會把我交在 掃羅 手裏嗎？ 掃羅 會下來，正如你僕人所聽見的嗎？耶和華－ 以色列 的上帝啊，求你指示僕人！」耶和華說：「他會下來。」
1SAM|23|12|大衛 又說：「 基伊拉 人會把我和我的人交在 掃羅 手裏嗎？」耶和華說：「他們會交出來。」
1SAM|23|13|於是 大衛 和他的人約有六百名起身離開 基伊拉 ，往他們所能去的地方去。有人告訴 掃羅 ， 大衛 離開 基伊拉 逃走了， 掃羅 就停止出發了。
1SAM|23|14|大衛 住在曠野的山寨裏，在 西弗 曠野的山區。 掃羅 天天尋索 大衛 ，上帝卻不將 大衛 交在他手裏。
1SAM|23|15|大衛 看到 掃羅 出來尋索他的命。那時，他住在 西弗 曠野的樹林裏 ；
1SAM|23|16|掃羅 的兒子 約拿單 起身，到樹林裏去見 大衛 ，使他的手倚靠上帝得以堅固，
1SAM|23|17|對他說：「不要懼怕！我父 掃羅 的手無法害你 ，你必作 以色列 的王，我必作你的宰相。我父 掃羅 也知道這事。」
1SAM|23|18|於是二人在耶和華面前立約。 大衛 仍住在樹林裏， 約拿單 就回家去了。
1SAM|23|19|西弗 人上 基比亞 到 掃羅 那裏，說：「 大衛 不是在我們那裏，在樹林裏的山寨中，在荒野 南邊的 哈基拉山 藏著嗎？
1SAM|23|20|現在，王啊，請隨你的心願要下來，就請下來；至於我們，一定會把他交在王的手裏。」
1SAM|23|21|掃羅 說：「願耶和華賜福給你們，因為你們體恤我。
1SAM|23|22|請你們回去，再確定一下，調查並看清楚他落腳的地方，是誰看見他在那裏 ，因為有人告訴我他很狡猾。
1SAM|23|23|你們要看清楚，調查他藏匿的每一個地方，回來給我確實的報告，我就與你們同去。他若在境內，我必從 猶大 的千門萬戶中搜出他來。」
1SAM|23|24|西弗 人動身，在 掃羅 以先往 西弗 去。 大衛 和他的人卻在 瑪雲 曠野，在荒野南邊的 亞拉巴 。
1SAM|23|25|掃羅 和他的人去尋索 大衛 。有人告訴 大衛 ，他就下到巖石那裏，留在 瑪雲 的曠野。 掃羅 聽見了，就在 瑪雲 的曠野追趕 大衛 。
1SAM|23|26|掃羅 在山的這一邊走， 大衛 和他的人在山的那一邊。 大衛 急忙躲避 掃羅 ， 掃羅 和他的人正四面圍住 大衛 和他的人，要捉拿他們。
1SAM|23|27|有使者來對 掃羅 說：「 非利士 人入境搶掠，請快快回去！」
1SAM|23|28|於是 掃羅 不再追趕 大衛 ，回去迎擊 非利士 人。因此那地方名叫 西拉‧哈瑪希羅結 。
1SAM|23|29|大衛 從那裏上去，住在 隱‧基底 的山寨裏。
1SAM|24|1|掃羅 追趕 非利士 人回來，有人告訴他說：「看哪， 大衛 在 隱‧基底 的曠野。」
1SAM|24|2|掃羅 就從全 以色列 中挑選三千精兵，往 野山羊磐石 的東邊 去，尋索 大衛 和他的人。
1SAM|24|3|到了路旁的羊圈，在那裏有個洞， 掃羅 進去大解。 大衛 和他的人正藏在洞裏的深處。
1SAM|24|4|大衛 的人對 大衛 說：「看哪，這日子到了！耶和華曾對你說：『看哪，我要將你的仇敵交在你手裏，你可以照你看為好的對待他。』」 大衛 就起來，悄悄地割下 掃羅 外袍的衣角。
1SAM|24|5|隨後 大衛 心中自責，因為他割下了 掃羅 的衣角。
1SAM|24|6|他對他的人說：「耶和華絕不允許我對我的主，耶和華的受膏者做這事，伸手害他，因為他是耶和華的受膏者。」
1SAM|24|7|大衛 用這話勸阻他的人，不許他們起來害 掃羅 。 掃羅 起來，從洞裏出去，預備上路。
1SAM|24|8|然後 大衛 也起來，從洞裏出去，呼喚 掃羅 說：「我主，我王！」 掃羅 回頭觀看， 大衛 就屈身，臉伏於地下拜。
1SAM|24|9|大衛 對 掃羅 說：「你為何聽信人的讒言，說『看哪， 大衛 想要害你』呢？
1SAM|24|10|看哪，今日你親眼看見，在洞中耶和華將你交在我手裏。有人要我殺你，我卻愛惜你，說：『我不敢伸手害我的主，因為他是耶和華的受膏者。』
1SAM|24|11|我父啊，請看，看你外袍的衣角在我手中。我割下你外袍的衣角，卻沒有殺你。你知道，並且看見我沒有惡意要悖逆你。你雖然要獵取我的命，我卻沒有得罪你。
1SAM|24|12|願耶和華在你我中間判斷，願耶和華在你身上為我伸冤，我卻不親手加害於你。
1SAM|24|13|古人有句俗語說：『惡事出於惡人。』我卻不親手加害於你。
1SAM|24|14|以色列 王出來要尋找誰呢？你要追趕誰呢？不過是一條死狗，一隻跳蚤而已。
1SAM|24|15|願耶和華作仲裁者，在你我中間判斷。願他鑒察，為我伸冤，救我脫離你的手。」
1SAM|24|16|大衛 向 掃羅 說完了這些話， 掃羅 說：「我兒 大衛 ，這是你的聲音嗎？」於是 掃羅 放聲大哭，
1SAM|24|17|對 大衛 說：「你比我公義，因為你以善待我，我卻以惡待你。
1SAM|24|18|今日你已顯明是以善待我，因為耶和華將我交在你手裏，你卻沒有殺我。
1SAM|24|19|人若遇見仇敵，豈肯放他平安上路呢？願耶和華因你今日向我所做的，以善回報你。
1SAM|24|20|現在，看哪，我知道你一定會作王， 以色列 的國必要堅立在你手裏。
1SAM|24|21|現在你要指著耶和華向我起誓，你必不剪除我的後裔，必不從我父家除去我的名。」
1SAM|24|22|於是 大衛 向 掃羅 起誓， 掃羅 就回家去， 大衛 和他的人也上山寨去了。
1SAM|25|1|撒母耳 死了， 以色列 眾人聚集，為他哀哭，把他葬在 拉瑪 他的家裏。 大衛 動身，下到 巴蘭 的曠野。
1SAM|25|2|在 瑪雲 有一個人，他的產業在 迦密 。這人是一個大富翁，有三千隻綿羊，一千隻山羊；他正在 迦密 剪羊毛。
1SAM|25|3|這人名叫 拿八 ，他的妻子名叫 亞比該 。 拿八 的妻子有美好的見識，又有美麗的容貌，但 拿八 為人剛愎兇惡，是 迦勒 族的人。
1SAM|25|4|大衛 在曠野聽見 拿八 正在剪羊毛，
1SAM|25|5|就派十個僕人，對他們說：「你們上 迦密 到 拿八 那裏，提我的名向他問安。
1SAM|25|6|你們要如此說：『願你來年平安 ，願你家平安，願你一切所有的都平安。
1SAM|25|7|現在我聽說你有剪羊毛的人，你的牧人和我們在一起，他們在 迦密 一切的日子，我們沒有欺負過他們，他們也未曾失去甚麼。
1SAM|25|8|你問你的僕人，他們會告訴你。願我的僕人在你眼前得歡心，因為我們是在好日子來的。請你隨手分點食物給僕人和你兒子 大衛 。』」
1SAM|25|9|大衛 的僕人到了，就提 大衛 的名，把這一切話告訴 拿八 ，他們就停頓下來。
1SAM|25|10|拿八 回答 大衛 的僕人說：「 大衛 是誰？ 耶西 的兒子是誰？今日悖逆主人奔逃的僕人很多。
1SAM|25|11|我豈可把飲食，以及我為剪羊毛的人所宰的肉給那些我不知道從哪裏來的人呢？」
1SAM|25|12|大衛 的僕人轉身從原路回去，照這一切的話告訴 大衛 。
1SAM|25|13|大衛 對他的人說：「你們各人都要佩上刀！」各人就都佩上刀， 大衛 也佩上刀。跟隨 大衛 上去的約有四百人，留下二百人看守物件。
1SAM|25|14|拿八 的一個僕人告訴 拿八 的妻子 亞比該 說：「看哪， 大衛 從曠野派使者來向我主人問安，主人卻辱罵他們。
1SAM|25|15|但是那些人待我們真好；我們在田野與他們一切來往的日子，沒有受他們欺負，也未曾失去甚麼。
1SAM|25|16|我們在他們那裏牧羊，一切的日子他們晝夜保護我們 。
1SAM|25|17|現在，你當知道，看怎樣做才好。不然，禍患必定臨到我主人和他全家。他性情兇暴，無人敢與他說話。」
1SAM|25|18|亞比該 急忙將二百個餅，兩皮袋酒，五隻宰好的羊，五細亞烘熟的穗子，一百個葡萄乾餅，二百個無花果餅，都馱在驢上，
1SAM|25|19|對僕人說：「你們在我前面走，看哪，我跟著你們去。」她卻沒有告訴丈夫 拿八 。
1SAM|25|20|亞比該 騎著驢，正下山坡，看哪， 大衛 和他的人正迎著 亞比該 下來，她就去迎接他們。
1SAM|25|21|大衛 曾說：「我在曠野為那人看守他一切所有的，以致他未失去任何一樣東西，實在是徒然了！他竟然向我以惡報善。
1SAM|25|22|凡屬 拿八 的男丁，我若留一個到明日早晨，願上帝重重懲罰 大衛 ！」
1SAM|25|23|亞比該 看見 大衛 ，就急忙下驢，在 大衛 面前臉伏於地叩拜。
1SAM|25|24|她俯伏在 大衛 的腳前，說：「我主啊，願這罪歸於我！求你容許使女向你進言，更求你聽使女的話。
1SAM|25|25|我主不必理會 拿八 這性情兇暴的人，他就像他的名字一樣；他名叫 拿八 ，為人也真是愚頑。至於我，你的使女並沒有看見我主所派來的僕人。
1SAM|25|26|現在，我主啊，耶和華既然阻止你親手報仇，避免流人的血，我指著永生的耶和華起誓，又指著你的性命起誓：『現在，願你的仇敵和謀害我主的人都像 拿八 一樣。』
1SAM|25|27|現在求我主把婢女送來的禮物給跟隨我主的僕人。
1SAM|25|28|求你原諒使女的冒犯。耶和華必為我主建立堅固的家，因為我主為耶和華爭戰，並且你一生的日子查不出有甚麼惡來。
1SAM|25|29|雖有人起來追逼你，要尋索你的性命，我主的性命在耶和華－你的上帝那裏，如同藏在生命的寶藏中。至於你仇敵的性命，耶和華必甩去，如用機弦甩石一樣。
1SAM|25|30|耶和華照所應許你的福氣賜給我主，立你作 以色列 王的時候，
1SAM|25|31|我主就不至於因為親手報仇，流了無辜人的血，而心裏不安，良心有虧了。耶和華賜福給我主的時候，求你記得你的使女。」
1SAM|25|32|大衛 對 亞比該 說：「耶和華－ 以色列 的上帝是應當稱頌的，因為他今日派你來迎接我。
1SAM|25|33|你和你的見識也配得稱讚，因為你今日攔阻我親手報仇、流人的血。
1SAM|25|34|我指著阻止我加害於你的耶和華－ 以色列 永生的上帝起誓，若不是你很快地來迎接我，到早晨天亮的時候，凡屬 拿八 的男丁，必定一個也不留。」
1SAM|25|35|大衛 從 亞比該 手中收了她帶來的禮物，對她說：「平平安安上你的家去吧！你看，我看了你的情面，聽了你的話。」
1SAM|25|36|亞比該 到 拿八 那裏，看哪，他在家裏擺設宴席，如同王的宴席。 拿八 心情舒暢，酩酊大醉。所以 亞比該 大小事都沒有告訴他，直等到早晨天亮的時候。
1SAM|25|37|到了早晨， 拿八 酒醒了，他的妻子把這些事都告訴他，他就發心臟病快死了，僵如石頭。
1SAM|25|38|過了十天，耶和華擊打 拿八 ，他就死了。
1SAM|25|39|大衛 聽見 拿八 死了，就說：「耶和華是應當稱頌的，因為我從 拿八 手中受了羞辱，他為我伸冤，又阻止他的僕人行惡；耶和華使 拿八 的惡歸到他自己頭上。」於是 大衛 派人去向 亞比該 說，要娶她為妻。
1SAM|25|40|大衛 的僕人來到 迦密 ，到 亞比該 那裏，對她說：「 大衛 派我們到你這裏，要娶你作他的妻子。」
1SAM|25|41|亞比該 起來叩拜，俯伏在地，說：「看哪，你的使女情願作婢女，為我主的僕人洗腳。」
1SAM|25|42|亞比該 立刻起身，騎上驢，五個女僕跟著她走。她跟從 大衛 的使者去，就作了 大衛 的妻子。
1SAM|25|43|大衛 先前娶了 耶斯列 人 亞希暖 ，她們二人都作了他的妻子。
1SAM|25|44|掃羅 已把他的女兒 米甲 ，就是 大衛 的妻子，給了 迦琳 人 拉億 的兒子 帕提 為妻。
1SAM|26|1|西弗 人來到 基比亞 ，到 掃羅 那裏，說：「 大衛 不是在荒野 東邊 的 哈基拉山 藏著嗎？」
1SAM|26|2|掃羅 動身，帶領 以色列 人中挑選的三千精兵下到 西弗 的曠野，要在那裏尋索 大衛 。
1SAM|26|3|掃羅 在荒野東邊的 哈基拉山 ，在路旁安營。那時 大衛 住在曠野，看見 掃羅 到曠野來追趕他，
1SAM|26|4|大衛 就派人去探聽，知道 掃羅 果然來了。
1SAM|26|5|大衛 起來，到 掃羅 安營的地方，看見 掃羅 和 尼珥 的兒子 押尼珥 元帥躺臥之處； 掃羅 睡在軍營裏，士兵安營在他周圍。
1SAM|26|6|大衛 對 赫 人 亞希米勒 和 洗魯雅 的兒子 約押 的兄弟 亞比篩 說：「誰同我下到 掃羅 營裏去？」 亞比篩 說：「我同你下去。」
1SAM|26|7|於是 大衛 和 亞比篩 夜間到了士兵那裏；看哪， 掃羅 睡在軍營裏，他的槍在頭旁，插在地上。 押尼珥 和士兵睡在他周圍。
1SAM|26|8|亞比篩 對 大衛 說：「上帝將你的仇敵交在你手裏，現在讓我拿槍把他刺透在地上，一刺就成，不用再刺他了。」
1SAM|26|9|大衛 對 亞比篩 說：「不可殺害他！有誰伸手害耶和華的受膏者而無罪呢？」
1SAM|26|10|大衛 又說：「我指著永生的耶和華起誓，他或被耶和華擊殺，或死期到了，或出戰陣亡，
1SAM|26|11|耶和華絕不允許我伸手害耶和華的受膏者。現在你可以把他頭旁的槍和水壺拿來，我們就走。」
1SAM|26|12|大衛 從 掃羅 的頭旁拿了槍和水壺，他們就走了。沒有人看見，沒有人知道，也沒有人醒過來。他們都睡著了，因為耶和華使他們沉睡了。
1SAM|26|13|大衛 過到另一邊去，遠遠地站在山頂上，與他們相離很遠。
1SAM|26|14|大衛 呼叫百姓和 尼珥 的兒子 押尼珥 說：「 押尼珥 ，你為何不回答呢？」 押尼珥 回答說：「你是誰？竟敢呼喚王呢？」
1SAM|26|15|大衛 對 押尼珥 說：「你不是個大丈夫嗎？ 以色列 中誰能比你呢？百姓中有一個人進來要害死你主你王，你為何沒有保護你主你王呢？
1SAM|26|16|你做的這件事不好！我指著永生的耶和華起誓，你們都是該死的，因為你們沒有保護你們的主，就是耶和華的受膏者。現在你看，王頭旁的槍和水壺在哪裏？」
1SAM|26|17|掃羅 認出 大衛 的聲音，就說：「我兒 大衛 ，這是你的聲音嗎？」 大衛 說：「我主我王啊，是我的聲音。」
1SAM|26|18|又說：「我主為何要追趕僕人呢？我做了甚麼？我手做了甚麼惡事呢？
1SAM|26|19|現在求我主我王聽僕人的話：若是耶和華激發你來攻擊我，願耶和華悅納供物；若是出於人，願他們在耶和華面前受詛咒，因為他們今日趕逐我，不讓我在耶和華的產業中有分，說：『你去事奉別神吧！』
1SAM|26|20|現在不要使我的血流在遠離耶和華面的地上。因為 以色列 王出來，只不過是尋找一隻跳蚤，如同人在山上獵取一隻鷓鴣。」
1SAM|26|21|掃羅 說：「我有罪了！我兒 大衛 ，回來吧！我必不再加害於你，因為你今日看我的性命為寶貴。看哪，我是個糊塗人，大大錯了。」
1SAM|26|22|大衛 回答說：「看哪，這是王的槍，可以吩咐一個僕人過來拿去。
1SAM|26|23|今日耶和華將王交在我手裏，我卻不肯伸手害耶和華的受膏者。耶和華必照各人的公義誠實報應他。
1SAM|26|24|看哪，我今日看重你的性命，願耶和華也照樣看重我的性命，並且拯救我脫離一切患難。」
1SAM|26|25|掃羅 對 大衛 說：「我兒 大衛 ，願你得福！你必做大事，也必得勝。」於是 大衛 上路， 掃羅 也回自己的地方去了。
1SAM|27|1|大衛 心裏說：「總有一天我會死在 掃羅 手裏，現在我最好逃到 非利士 人的地去， 掃羅 就會絕望，不會繼續在 以色列 全境內尋索我了。這樣，我才可以脫離他的手。」
1SAM|27|2|於是 大衛 動身，和跟隨他的六百人投奔 瑪俄 的兒子 迦特 王 亞吉 去了。
1SAM|27|3|大衛 和他的兩個妻子，就是 耶斯列 人 亞希暖 和作過 拿八 妻子的 迦密 人 亞比該 ，以及他的人，連同各人的眷屬，都住在 迦特 的 亞吉 那裏。
1SAM|27|4|有人告訴 掃羅 ：「 大衛 逃到 迦特 。」 掃羅 就不再尋索他了。
1SAM|27|5|大衛 對 亞吉 說：「我若蒙你看得起，求你在郊外的城鎮中賜我一個地方，讓我住在那裏。僕人何必與王同住京城呢？」
1SAM|27|6|當日 亞吉 把 洗革拉 賜給他，因此 洗革拉 屬於 猶大 王，直到今日。
1SAM|27|7|大衛 在 非利士 人的地，住的期間有一年四個月。
1SAM|27|8|大衛 和他的人上去，侵奪 基述 人、 基色 人、 亞瑪力 人，這些是從 帖蘭 經過 書珥 直到 埃及 地的居民 。
1SAM|27|9|大衛 攻擊那地，無論男女沒有留下一個活口，又奪獲牛、羊、驢、駱駝和衣服，回來到 亞吉 那裏。
1SAM|27|10|亞吉 說：「今日你們沒有去搶奪甚麼地方吧 ？」 大衛 說：「侵奪了 猶大 、 耶拉篾 、 基尼 等地的南方。」
1SAM|27|11|無論男女， 大衛 沒有留下一個活口帶到 迦特 來。他說：「恐怕他們把我們的事告訴人，說：『 大衛 如此做了。』」這是他住在 非利士 人之地一切日子的慣例。
1SAM|27|12|亞吉 信了 大衛 ，說：「 大衛 已經使本族 以色列 人憎惡他，所以他必永遠作我的僕人了。」
1SAM|28|1|那時， 非利士 人召集軍隊，要與 以色列 打仗。 亞吉 對 大衛 說：「你當知道，你和你的人都要隨我出征。」
1SAM|28|2|大衛 對 亞吉 說：「好，僕人所能做的事，王都知道。」 亞吉 對 大衛 說：「好，我立你終生作我 的侍衛。」
1SAM|28|3|那時 撒母耳 已經死了， 以色列 眾人為他哀哭，把他葬在他的本城 拉瑪 。 掃羅 曾在國內驅除招魂的和行巫術的人。
1SAM|28|4|非利士 人集合，來到 書念 安營； 掃羅 集合 以色列 眾人在 基利波 安營。
1SAM|28|5|掃羅 看見 非利士 的軍隊，就懼怕，心中大大戰兢。
1SAM|28|6|掃羅 求問耶和華，耶和華卻不藉夢，或烏陵，或先知回答他。
1SAM|28|7|掃羅 吩咐臣僕說：「為我找一個招魂的婦人，我好去問她。」臣僕對他說：「看哪，在 隱‧多珥 有一個招魂的婦人。」
1SAM|28|8|於是 掃羅 改了裝，穿上別的衣服，帶著兩個人，夜裏去見那婦人。 掃羅 說：「請你用招魂的法術，把我所告訴你的死人，為我招上來。」
1SAM|28|9|婦人對他說：「看哪，你知道 掃羅 所做的，他從國中剪除招魂的和行巫術的。你為何為我的性命設下羅網，要害死我呢？」
1SAM|28|10|掃羅 向婦人指著耶和華起誓說：「我指著永生的耶和華起誓，你必不因這事受罰。」
1SAM|28|11|婦人說：「我為你招誰上來呢？」他說：「為我招 撒母耳 上來。」
1SAM|28|12|婦人看見 撒母耳 ，就大聲喊叫。婦人對 掃羅 說：「你是 掃羅 ，為甚麼欺騙我呢？」
1SAM|28|13|王對婦人說：「不要懼怕，你看見甚麼呢？」婦人對 掃羅 說：「我看見有神明從地裏上來。」
1SAM|28|14|掃羅 說：「他是怎樣的形狀？」婦人說：「有一個老人上來，身穿長袍。」 掃羅 知道是 撒母耳 ，就屈身，臉伏於地下拜。
1SAM|28|15|撒母耳 對 掃羅 說：「你為甚麼攪擾我，招我上來呢？」 掃羅 說：「我十分為難，因為 非利士 人攻擊我，上帝離開我，不再藉先知或夢回答我。因此請你上來，好指示我應當怎樣做。」
1SAM|28|16|撒母耳 說：「耶和華已經離開你，與你為敵，你何必問我呢？
1SAM|28|17|耶和華照他藉我所說的話為他自己 實現了。耶和華已經從你手裏奪去國權，賜給別人，就是 大衛 。
1SAM|28|18|因為你沒有聽從耶和華的話，沒有執行他對 亞瑪力 人的惱怒，所以今日耶和華向你做這事。
1SAM|28|19|耶和華也必將你和 以色列 交在 非利士 人手裏。明日你和你兒子們必與我在一處了；耶和華也必將 以色列 的軍兵交在 非利士 人手裏。」
1SAM|28|20|掃羅 突然全身仆倒在地，因為 撒母耳 的話令他十分懼怕。他毫無氣力，因為他一日一夜都沒有吃甚麼。
1SAM|28|21|婦人到 掃羅 面前，見他極其驚恐，對他說：「看哪，婢女聽從了你，不顧惜自己的性命，遵從你吩咐我的話。
1SAM|28|22|現在求你也聽婢女的話，讓我在你面前擺上一點食物，你吃了才有氣力上路。」
1SAM|28|23|掃羅 不肯，說：「我不吃。」但他的僕人和那婦人再三勸他，他才聽他們的話，從地上起來，坐在床上。
1SAM|28|24|婦人急忙把家裏的一隻肥牛犢宰了，又拿麵來揉，烤成無酵餅，
1SAM|28|25|擺在 掃羅 和他僕人面前。他們吃了，當夜就起身走了。
1SAM|29|1|非利士 人聚集他們所有的軍隊到 亞弗 ； 以色列 人在 耶斯列 的泉旁安營。
1SAM|29|2|非利士 人的領袖各率隊伍，或百或千的前進； 大衛 和他的人同 亞吉 跟在後邊前進。
1SAM|29|3|非利士 人的領袖說：「這些 希伯來 人在這裏做甚麼呢？」 亞吉 對 非利士 人的領袖說：「這不是 以色列 王 掃羅 的臣僕 大衛 嗎？他在我這裏有些年日了。自從他投降直到今日，我未曾見他有甚麼過錯。」
1SAM|29|4|非利士 人的領袖向 亞吉 發怒，對他說：「叫這人回去！叫他回到你指派他的地方去，不可讓他同我們出征，免得他在陣上反成為我們的敵人。他用甚麼與他主人復和呢？豈不是用我們這些人的首級嗎？
1SAM|29|5|有人跳舞唱和說： 『 掃羅 殺死千千， 大衛 殺死萬萬』， 不就是這個 大衛 嗎？」
1SAM|29|6|亞吉 叫 大衛 來，對他說：「我指著永生的耶和華起誓，你是個正直人。你隨我在軍中出入，我也很滿意。自從你投奔我到如今，我未曾看見你有甚麼過失，但是眾領袖看你不順眼。
1SAM|29|7|現在你平平安安地回去，不要做 非利士 人領袖眼中看為惡的事。」
1SAM|29|8|大衛 對 亞吉 說：「但我做了甚麼呢？自從僕人到你面前，直到今日，你查出我有甚麼過錯，使我不去攻擊我主我王的仇敵呢？」
1SAM|29|9|亞吉 回答 大衛 說：「我知道你在我眼中是好人，如同上帝的使者一樣，只是 非利士 人的領袖說：『這人不可同我們上戰場。』
1SAM|29|10|現在，你和跟隨你來的，就是你主人的僕人，清晨要早早起來，回到我所指派你的地方去，不要把中傷的話放在心上，因為你在我面前很好 。你們清晨早早起來，天一亮就回去吧！」
1SAM|29|11|於是 大衛 和他的人清晨早早起來，回到 非利士 人的地去。 非利士 人也上 耶斯列 去了。
1SAM|30|1|第三日， 大衛 和他的人到了 洗革拉 。 亞瑪力 人已經侵奪 尼革夫 和 洗革拉 。他們攻破 洗革拉 ，用火焚燒。
1SAM|30|2|他們擄去城內的婦女和城中的大小人口，一個都沒有殺，全都帶走，他們就上路去了。
1SAM|30|3|大衛 和他的人到了那城，看哪，城已被火燒燬，他們的妻子兒女都被擄去了。
1SAM|30|4|大衛 和跟隨他的百姓就放聲大哭，直到沒有氣力再哭。
1SAM|30|5|大衛 的兩個妻子， 耶斯列 人 亞希暖 和作過 拿八 妻子的 迦密 人 亞比該 ，也被擄去了。
1SAM|30|6|大衛 非常焦急，因為眾百姓為自己的兒女痛心，說要用石頭打死他。 大衛 卻倚靠耶和華－他的上帝，堅定自己。
1SAM|30|7|大衛 對 亞希米勒 的兒子 亞比亞他 祭司說：「請你把以弗得拿來給我。」 亞比亞他 就把以弗得拿給 大衛 。
1SAM|30|8|大衛 求問耶和華說：「我追趕這群人，是否追得上呢？」耶和華對他說：「你可以追，一定追得上，也一定救得回來。」
1SAM|30|9|於是， 大衛 出發，他和跟隨他的六百人來到 比梭溪 ，那些不能前去的就留在那裏。
1SAM|30|10|大衛 帶著四百人往前追趕；有二百人疲乏，不能過 比梭溪 ，留在那裏。
1SAM|30|11|這四百人在田野遇見一個 埃及 人，就帶他到 大衛 面前，給他餅吃，給他水喝，
1SAM|30|12|又給他一塊無花果餅，兩個葡萄乾餅。他吃了，精神就恢復了，因為他三日三夜沒有吃餅，沒有喝水。
1SAM|30|13|大衛 對他說：「你是誰的人？你從哪裏來？」他說：「我是 埃及 的青年，是 亞瑪力 人的奴僕。因為我三天前生病，我主人就把我撇棄了。
1SAM|30|14|我們侵奪了 基利提 的南方和屬 猶大 的地，以及 迦勒 地的南方，又用火燒了 洗革拉 。」
1SAM|30|15|大衛 對他說：「你肯領我們下到那群人那裏嗎？」他說：「你要向我指著上帝起誓，你不殺我，也不把我交在我主人手裏，我就領你下到那群人那裏。」
1SAM|30|16|那人領 大衛 下去，看哪，他們分散在全地面，吃喝跳舞，因為他們從 非利士 人的地和 猶大 地擄來的財物非常多。
1SAM|30|17|大衛 擊殺他們，從黎明直到次日晚上，除了四百個騎駱駝逃走的青年之外，一個也沒有逃脫。
1SAM|30|18|亞瑪力 人所擄去的財物， 大衛 全都奪回，並救回他的兩個妻子。
1SAM|30|19|凡 亞瑪力 人所擄去的，無論大小、兒女、掠物和一切被擄去的， 大衛 全都奪回來。
1SAM|30|20|大衛 所奪來的牛群羊群，有人趕在群畜前面，說：「這是 大衛 的掠物。」
1SAM|30|21|大衛 到了那疲乏不能跟隨、留在 比梭溪 的二百人那裏。他們出來迎接 大衛 和跟隨他的百姓。 大衛 上前向他們問安。
1SAM|30|22|跟隨 大衛 去的人中，每一個惡人和無賴都說：「這些人既然沒有和我同去，我們所奪的財物就不分給他們，只把他們各人的妻子兒女給他們，讓他們帶回去就好了。」
1SAM|30|23|大衛 說：「我的弟兄，耶和華所賜給我們的，你們不可這麼做，因為他保佑了我們，把那群來攻擊我們的人交在我們手裏。
1SAM|30|24|誰肯在這事上聽你們呢？上陣的分得多少，留下看守物件的也分得多少，大家應當平分。」
1SAM|30|25|從那日起， 大衛 定此為 以色列 的律例典章，直到今日。
1SAM|30|26|大衛 到了 洗革拉 ，從掠物中取些送給他的朋友，就是 猶大 的長老，說：「看哪，這是從耶和華仇敵那裏奪來的，送給你們作禮物。」
1SAM|30|27|有在 伯特利 的， 尼革夫 之 拉末 的， 雅提珥 的，
1SAM|30|28|有在 亞羅珥 的， 息末 的， 以實提莫 的，
1SAM|30|29|有在 拉哈勒 的， 耶拉篾 各城的， 基尼 各城的，
1SAM|30|30|有在 何珥瑪 的， 坡拉珊 的， 亞撻 的，
1SAM|30|31|有在 希伯崙 的，以及 大衛 和跟隨他的人經常進出之處的。
1SAM|31|1|非利士 人攻打 以色列 。 以色列 人在 非利士 人面前逃跑，很多人 在 基利波山 被殺仆倒。
1SAM|31|2|非利士 人緊追 掃羅 和他的兒子，殺了 掃羅 的兒子 約拿單 、 亞比拿達 、 麥基‧舒亞 。
1SAM|31|3|攻擊 掃羅 的戰事激烈，弓箭手追上他，他被弓箭手射中，傷勢很重 。
1SAM|31|4|掃羅 吩咐拿他兵器的人說：「你拔出刀來，把我刺死，免得那些未受割禮的人來刺我，凌辱我。」但拿兵器的人不肯，因為他非常懼怕。於是 掃羅 拿起刀來，伏在刀上。
1SAM|31|5|拿兵器的人見 掃羅 已死，也伏在刀上跟他一起死。
1SAM|31|6|這樣， 掃羅 和他三個兒子，與拿他兵器的人，以及他所有的人 ，都在那日一起死了。
1SAM|31|7|住平原那邊和 約旦河 那邊的 以色列 人，見 以色列 軍兵逃跑， 掃羅 和他兒子都死了，就棄城逃跑。 非利士 人前來住在其中。
1SAM|31|8|次日， 非利士 人來剝那些被殺之人的衣服，看見 掃羅 和他三個兒子仆倒在 基利波山 。
1SAM|31|9|他們割下他的首級，剝了他的盔甲，派人到 非利士 人之地的四境，報信給他們廟裏的偶像和百姓。
1SAM|31|10|他們將 掃羅 的盔甲放在 亞斯她錄 廟裏，把他的屍身釘在 伯‧珊 的城牆上。
1SAM|31|11|基列 的 雅比 居民聽見 非利士 人向 掃羅 所行的事，
1SAM|31|12|他們所有的勇士就起身，走了一夜，把 掃羅 和他兒子的屍身從 伯‧珊 城牆上取下來，送到 雅比 ，在那裏用火燒了，
1SAM|31|13|把骸骨葬在 雅比 的柳樹下，並且禁食七日。
2SAM|1|1|掃羅 死後， 大衛 擊殺 亞瑪力 人回來，在 洗革拉 住了兩天。
2SAM|1|2|第三天，看哪，有一人從 掃羅 的營裏出來，衣服撕裂，頭蒙灰塵，到 大衛 面前伏地叩拜。
2SAM|1|3|大衛 對他說：「你從哪裏來？」他說：「我從 以色列 的營裏逃來。」
2SAM|1|4|大衛 又對他說：「事情怎麼樣？請你告訴我。」他說：「士兵從陣上逃跑，也有許多士兵仆倒死亡， 掃羅 和他兒子 約拿單 也死了。」
2SAM|1|5|大衛 問報信的青年說：「你怎麼知道 掃羅 和他兒子 約拿單 死了呢？」
2SAM|1|6|報信的青年說：「我恰巧到 基利波山 ，看哪， 掃羅 靠在自己的槍上，看哪，有戰車、騎兵緊緊地追他。
2SAM|1|7|他回頭看見我，就呼叫我。我說：『我在這裏。』
2SAM|1|8|他問我說：『你是甚麼人？』我說：『我是 亞瑪力 人。』
2SAM|1|9|他對我說：『請你站到我這裏來，把我殺死，因為我非常痛苦，只剩下一口氣。』
2SAM|1|10|我就站到他那裏，殺了他，因為我知道他一倒下就活不了。然後，我把他頭上的冠冕和臂上的鐲子拿到我主這裏來。」
2SAM|1|11|大衛 就抓著自己的衣服，把衣服撕裂，所有跟隨他的人也都如此。
2SAM|1|12|他們為 掃羅 和他兒子 約拿單 ，以及耶和華的百姓和 以色列 家的人悲哀哭泣，禁食到晚上，因為他們都倒在刀下。
2SAM|1|13|大衛 問報信的青年說：「你是哪裏人？」他說：「我是一個寄居者的兒子，是 亞瑪力 人。」
2SAM|1|14|大衛 對他說：「你動手殺害耶和華的受膏者，怎麼不畏懼呢？」
2SAM|1|15|大衛 叫了一個僕人來，說：「來，殺了他！」僕人擊殺他，他就死了。
2SAM|1|16|大衛 對他說：「你的血歸到你自己頭上，因為你親口作證控訴自己，說：『我殺了耶和華的受膏者。』」
2SAM|1|17|大衛 作了這首哀歌，哀悼 掃羅 和他兒子 約拿單 ，
2SAM|1|18|並吩咐人把這首「弓歌」教導 猶大 人，看哪，它寫在《雅煞珥書》上：
2SAM|1|19|以色列 啊，尊榮者在你的高處被殺！ 大英雄竟然仆倒！
2SAM|1|20|不要在 迦特 報告， 不要在 亞實基倫 街上傳揚， 免得 非利士 的女子歡喜， 免得未受割禮之人的女子歡樂。
2SAM|1|21|基利波山 哪，願你那裏沒有雨，沒有露！ 願你的田地無土產可作供物！ 因為英雄的盾牌在那裏受辱， 掃羅 的盾牌沒有抹油。
2SAM|1|22|在被殺者的血前， 在勇士的脂肪前， 約拿單 的弓絕不退縮， 掃羅 的刀斷不虛回。
2SAM|1|23|掃羅 和 約拿單 生時相悅相愛， 死時也不分離。 他們比鷹更快， 比獅子還強。
2SAM|1|24|以色列 的女子啊，當為 掃羅 哭泣！ 他曾使你們穿朱紅色的美衣， 使你們衣服有黃金的妝飾。
2SAM|1|25|英雄竟然在陣上仆倒！ 約拿單 竟然在你的高處被殺！
2SAM|1|26|我兄 約拿單 哪，我為你悲傷！ 我甚喜愛你！ 你對我的愛何等奇妙， 過於婦女的愛情。
2SAM|1|27|英雄竟然仆倒！ 兵器竟然廢棄！
2SAM|2|1|此後， 大衛 求問耶和華說：「我可以上 猶大 的一個城去嗎？」耶和華對他說：「可以上去。」 大衛 說：「我上哪一個城去呢？」耶和華說：「 希伯崙 。」
2SAM|2|2|於是 大衛 和他的兩個妻子，一個是 耶斯列 人 亞希暖 ，一個是作過 迦密 人 拿八 妻子的 亞比該 ，都上那裏去了。
2SAM|2|3|大衛 也把跟隨他的人和他們各人的眷屬一同帶上去，住在 希伯崙 的城鎮中。
2SAM|2|4|猶大 人來，在那裏膏 大衛 作 猶大 家的王。 有人告訴 大衛 說：「埋葬 掃羅 的是 基列 的 雅比 人。」
2SAM|2|5|大衛 就派使者到 基列 的 雅比 人那裏，對他們說：「願耶和華賜福給你們！因為你們忠心對待你們的主 掃羅 ，埋葬了他。
2SAM|2|6|你們既做了這事，願耶和華以慈愛和信實待你們，我也要為此厚待你們。
2SAM|2|7|現在，你們的主 掃羅 死了， 猶大 家也已經膏我作他們的王，你們的手要堅強，要作英勇的人。」
2SAM|2|8|掃羅 軍隊的元帥， 尼珥 的兒子 押尼珥 ，曾將 掃羅 的兒子 伊施．波設 帶過河，到 瑪哈念 ，
2SAM|2|9|立他作王，治理 基列 、 亞書利 、 耶斯列 、 以法蓮 、 便雅憫 和 以色列 眾人。
2SAM|2|10|掃羅 的兒子 伊施．波設 登基的時候年四十歲，作 以色列 王二年，但是 猶大 家卻隨從 大衛 。
2SAM|2|11|大衛 在 希伯崙 作 猶大 家的王，共七年六個月。
2SAM|2|12|尼珥 的兒子 押尼珥 和 掃羅 的兒子 伊施．波設 的僕人從 瑪哈念 出來，往 基遍 去。
2SAM|2|13|洗魯雅 的兒子 約押 和 大衛 的僕人也出來，在 基遍 池旁與他們相遇；一隊坐在池的這邊，一隊坐在池的那邊。
2SAM|2|14|押尼珥 對 約押 說：「讓年輕人起來，在我們面前較量一下吧！」 約押 說：「讓他們起來吧。」
2SAM|2|15|他們就起來，點了人數過來：屬 掃羅 兒子 伊施．波設 的有 便雅憫 人十二名， 大衛 的僕人也有十二名。
2SAM|2|16|每人抓住對方的頭，用刀刺對方的肋旁，一同仆倒。所以，那地叫做 希利甲‧哈素林 ，就在 基遍 。
2SAM|2|17|那日戰況激烈， 押尼珥 和 以色列 人敗在 大衛 的僕人面前。
2SAM|2|18|在那裏有 洗魯雅 的三個兒子： 約押 、 亞比篩 、 亞撒黑 。 亞撒黑 的腳快如野地裏的羚羊；
2SAM|2|19|亞撒黑 追趕 押尼珥 ，直追趕他不偏左右。
2SAM|2|20|押尼珥 回頭說：「 亞撒黑 ，是你嗎？」他說：「是我。」
2SAM|2|21|押尼珥 對他說：「你轉左或轉右，去抓一個年輕人，剝去他的戰衣吧。」 亞撒黑 卻不肯轉開而不追趕他。
2SAM|2|22|押尼珥 又對 亞撒黑 說：「轉開，不要再追我了！我何必把你擊殺在地上呢？我若殺了你，怎麼有臉見你哥哥 約押 呢？」
2SAM|2|23|亞撒黑 仍不肯轉開， 押尼珥 就用回馬槍 刺入他的肚腹，甚至槍從背後穿出， 亞撒黑 就仆倒在那裏，當場死了。眾人趕到 亞撒黑 仆倒而死的地方，就都站住。
2SAM|2|24|約押 和 亞比篩 追趕 押尼珥 。日落的時候，他們到了通往 基遍 曠野的路旁， 基亞 對面的 亞瑪山 。
2SAM|2|25|便雅憫 人聚集在 押尼珥 後面，成為一隊，站在一座山頂上。
2SAM|2|26|押尼珥 呼叫 約押 說：「刀劍豈可永遠吞噬呢？你豈不知，結局必是痛苦的嗎？你要等到何時才叫百姓回去，不追趕他們的弟兄呢？」
2SAM|2|27|約押 說：「我指著永生的上帝起誓：你若沒有這麼說，百姓就必繼續追趕弟兄，直到早晨 。」
2SAM|2|28|於是 約押 吹角，眾百姓就站住，不再追趕 以色列 人，也不再打仗了。
2SAM|2|29|押尼珥 和他的人整夜行過 亞拉巴 。他們過了 約旦河 ，走過 畢倫 ，到了 瑪哈念 。
2SAM|2|30|約押 追趕 押尼珥 回來，聚集眾百姓， 大衛 的僕人中缺少了十九個人和 亞撒黑 。
2SAM|2|31|但 大衛 的僕人殺了 押尼珥 的人， 便雅憫 人三百六十名。
2SAM|2|32|他們把 亞撒黑 送到 伯利恆 ，葬在他父親的墳墓裏。 約押 和他的人走了一整夜，天亮的時候他們才到 希伯崙 。
2SAM|3|1|掃羅 家和 大衛 家爭戰許久。 大衛 家日見強盛， 掃羅 家卻日見衰弱。
2SAM|3|2|大衛 在 希伯崙 生了幾個兒子：長子 暗嫩 是 耶斯列 人 亞希暖 所生的；
2SAM|3|3|次子 基利押 是作過 迦密 人 拿八 的妻子 亞比該 所生的；三子 押沙龍 是 基述 王 達買 的女兒 瑪迦 所生的；
2SAM|3|4|四子 亞多尼雅 是 哈及 所生的；五子 示法提雅 是 亞比她 所生的；
2SAM|3|5|六子 以特念 是 大衛 的妻子 以格拉 所生的。 大衛 這六個兒子都是在 希伯崙 生的。
2SAM|3|6|掃羅 家和 大衛 家爭戰的時候， 押尼珥 在 掃羅 家大有權勢。
2SAM|3|7|掃羅 有一妃子，名叫 利斯巴 ，是 愛亞 的女兒。一日， 伊施．波設 對 押尼珥 說：「你為甚麼與我父的妃子同寢呢？」
2SAM|3|8|押尼珥 因 伊施．波設 的話非常生氣，說：「我豈是狗的頭，向著 猶大 呢？我今日忠心對待你父 掃羅 的家和他的弟兄、朋友，不將你交在 大衛 手裏，今日你竟為這婦人責備我嗎？
2SAM|3|9|願上帝重重懲罰 押尼珥 ！我要照著耶和華起誓應許 大衛 的話為他成就，
2SAM|3|10|廢去 掃羅 家的國度，建立 大衛 的王位，使他治理 以色列 和 猶大 ，從 但 直到 別是巴 。」
2SAM|3|11|伊施．波設 懼怕 押尼珥 ，一句話也不能回答。
2SAM|3|12|押尼珥 派使者到 大衛 所在的地方 ，說：「這地歸誰呢？」又說：「你與我立約，看哪，我必幫助你，使全 以色列 都擁護你。」
2SAM|3|13|大衛 說：「好！我與你立約。但有一件事我要求你，你來見我面的時候，除非把 掃羅 的女兒 米甲 帶來，就不必來見我的面了。」
2SAM|3|14|大衛 派使者到 掃羅 的兒子 伊施．波設 那裏，說：「你要把我的妻子 米甲 歸還我；她是我從前用一百 非利士 人的包皮所聘定的。」
2SAM|3|15|伊施．波設 就派人去，把 米甲 從 拉億 的兒子，她丈夫 帕鐵 那裏帶來。
2SAM|3|16|米甲 的丈夫跟著她，一面走一面哭，直跟到 巴戶琳 。 押尼珥 對他說：「你回去吧！」 帕鐵 就回去了。
2SAM|3|17|押尼珥 與 以色列 長老商議，說：「從前你們企盼 大衛 作王治理你們，
2SAM|3|18|現在你們可以這樣做了。因為耶和華曾論到 大衛 說：『我必藉我僕人 大衛 的手，救我民 以色列 脫離 非利士 人和眾仇敵的手。』」
2SAM|3|19|押尼珥 也說給 便雅憫 人聽。 押尼珥 又到 希伯崙 ，把 以色列 人和 便雅憫 全家所看為好的，說給 大衛 聽。
2SAM|3|20|押尼珥 帶著二十個人來到 希伯崙大衛 那裏， 大衛 就為 押尼珥 和他帶來的人擺設宴席。
2SAM|3|21|押尼珥 對 大衛 說：「我要起身去召集全 以色列 ，來到我主我王這裏，與你立約，你就可以照你的心願作王，統治一切。」於是 大衛 送走 押尼珥 ，他就平安地去了。
2SAM|3|22|看哪， 大衛 的僕人和 約押 突擊回來，帶回許多掠物。那時 押尼珥 不在 希伯崙大衛 那裏，因 大衛 已經送他走，他也平安地去了。
2SAM|3|23|約押 和跟隨他的全軍到了，有人告訴 約押 說：「 尼珥 的兒子 押尼珥 來到王這裏，王送走他，他也平安地去了。」
2SAM|3|24|約押 到王那裏，說：「你這是做甚麼呢？看哪， 押尼珥 來到你這裏，你為何送他走，讓他去了呢？
2SAM|3|25|你知道， 尼珥 的兒子 押尼珥 來，是要騙你，要打聽你的出入，知道你一切所行的事。」
2SAM|3|26|約押 從 大衛 那裏出來，派些使者去追 押尼珥 ，從 西拉井 那裏帶他回來， 大衛 卻不知道。
2SAM|3|27|押尼珥 回到 希伯崙 ， 約押 領他到城門中間，要與他私下交談，就在那裏刺穿了他的肚腹。他就死了，因為他流了 約押 兄弟 亞撒黑 的血。
2SAM|3|28|這事以後， 大衛 聽見了，說：「流 尼珥 兒子 押尼珥 的血，我和我的國在耶和華面前永遠是無辜的。
2SAM|3|29|願這血歸到 約押 頭上和他父的全家；又願 約押 家不斷有患漏症的，長痲瘋 的，架柺杖而行的 ，仆倒在刀下的，缺乏食物的。」
2SAM|3|30|約押 和他弟弟 亞比篩 殺了 押尼珥 ，是因為在 基遍 戰爭的時候， 押尼珥 殺了他們的弟弟 亞撒黑 。
2SAM|3|31|大衛 對 約押 和跟隨他的眾百姓說：「你們當撕裂衣服，腰束麻布，在 押尼珥 前面哀哭。」 大衛 王也跟在棺木後面。
2SAM|3|32|他們把 押尼珥 葬在 希伯崙 。王在 押尼珥 的墓旁放聲大哭，眾百姓也都哭了。
2SAM|3|33|王為 押尼珥 舉哀，說： 押尼珥 怎麼會像愚頑人一樣地死呢？
2SAM|3|34|你手未曾被捆綁，腳未曾被腳鐐鎖住。 你仆倒，如仆倒在兇惡之子手下一樣。 於是眾百姓又為 押尼珥 哀哭。
2SAM|3|35|白天的時候，眾百姓來勸 大衛 吃飯，但 大衛 起誓說：「我若在太陽未下山以前吃飯，或吃任何東西，願上帝重重懲罰我！」
2SAM|3|36|眾百姓知道了就看為好。凡王所做的，眾百姓都看為好。
2SAM|3|37|那日， 以色列 眾百姓才知道殺 尼珥 的兒子 押尼珥 並非出於王意。
2SAM|3|38|王對臣僕說：「你們豈不知今日在 以色列 中倒了一個作元帥的大人物嗎？
2SAM|3|39|我雖然受膏為王，今日還是軟弱。 洗魯雅 的兩個兒子，這些人比我強硬。願耶和華照著惡人所行的惡報應他。」
2SAM|4|1|掃羅 的兒子 伊施．波設 聽見 押尼珥 死在 希伯崙 ，手就發軟，全 以色列 也都驚惶。
2SAM|4|2|掃羅 的兒子 伊施．波設 有兩個軍官，一個叫 巴拿 ，第二個叫 利甲 ，都是 便雅憫 支派 比錄 人 臨門 的兒子；因為 比錄 也算是屬於 便雅憫 的。
2SAM|4|3|比錄 人先前逃到 基他音 ，在那裏寄居，直到今日。
2SAM|4|4|掃羅 的兒子 約拿單 有一個兒子，名叫 米非波設 ，是瘸腿的。 掃羅 和 約拿單 的消息從 耶斯列 傳來的時候，他才五歲。他的奶媽抱著他逃跑；因為跑得太急，孩子掉在地上，腿就瘸了。
2SAM|4|5|比錄 人 臨門 的兩個兒子 利甲 和 巴拿 出去，天正熱的時候到了 伊施．波設 的家。那時， 伊施．波設 在睡午覺。
2SAM|4|6|婦人進到房子中間，要取麥子。 利甲 和他的哥哥 巴拿 刺穿了 伊施．波設 的肚腹，然後逃跑了。
2SAM|4|7|他們進到房子的時候， 伊施．波設 正躺在臥房的床上，他們就把他殺死，割了他的首級，拿著首級在 亞拉巴 的路上走了一整夜。
2SAM|4|8|他們把 伊施．波設 的首級拿到 希伯崙 大衛 那裏，對王說：「王的仇敵 掃羅 曾尋索你的性命。看哪，這是他兒子 伊施．波設 的首級；耶和華今日為我主我王在 掃羅 和他後裔身上報了仇。」
2SAM|4|9|大衛 回答 比錄 人 臨門 的兒子 利甲 和他哥哥 巴拿 說：「我指著救我性命脫離一切苦難、永生的耶和華起誓：
2SAM|4|10|從前有人告訴我說：『看哪， 掃羅 死了。』他自以為報好消息，我就拿住他，把他殺在 洗革拉 ，作為他報消息的賞賜。
2SAM|4|11|更何況惡人把義人殺在他家的床上，我豈不從你們手中追討他的血，從地上除滅你們嗎？」
2SAM|4|12|於是 大衛 吩咐僕人把他們殺了，砍斷他們的手腳，掛在 希伯崙 的池旁。然後，他們把 伊施．波設 的首級葬在 希伯崙押尼珥 的墳墓裏。
2SAM|5|1|以色列 眾支派來到 希伯崙 見 大衛 ，說：「看哪，我們是你的骨肉。
2SAM|5|2|從前 掃羅 作我們王的時候，率領 以色列 人出入的是你。耶和華也曾對你說：『你必牧養我的百姓 以色列 ，你必作 以色列 的君王。』」
2SAM|5|3|於是 以色列 的眾長老都來到 希伯崙 見王 。 大衛 在 希伯崙 ，在耶和華面前與他們立約，他們就膏 大衛 作 以色列 的王。
2SAM|5|4|大衛 登基的時候年三十歲，作王四十年。
2SAM|5|5|他在 希伯崙 作 猶大 王七年六個月，在 耶路撒冷 作 以色列 和 猶大 王三十三年。
2SAM|5|6|王和他的人到了 耶路撒冷 ，要攻打住那地方的 耶布斯 人。 耶布斯 人對 大衛 說：「你必不能進到這裏，就是盲人、瘸子都可以把你擊退。」就是說：「 大衛 絕不能進到這裏。」
2SAM|5|7|然而 大衛 攻取了 錫安 的堡壘，就是 大衛 的城。
2SAM|5|8|當日， 大衛 說：「誰攻打 耶布斯 人，就要從水道上去，攻打我心裏所恨惡的 瘸子、盲人。」因此有人說：「盲人和瘸子不得進殿裏去。」
2SAM|5|9|大衛 住在堡壘裏，給它起名叫 大衛城 。 大衛 又從 米羅 往內，周圍建築。
2SAM|5|10|大衛 日見強大，耶和華－萬軍之上帝與他同在。
2SAM|5|11|推羅 王 希蘭 派使者把香柏木運到 大衛 那裏，又派木匠和石匠給 大衛 建造宮殿。
2SAM|5|12|大衛 知道耶和華堅立他作 以色列 王，又為自己百姓 以色列 的緣故，使他的國興盛。
2SAM|5|13|大衛 離開 希伯崙 之後，在 耶路撒冷 又立后妃，又生兒女。
2SAM|5|14|在 耶路撒冷 所生的孩子的名字是 沙母亞 、 朔罷 、 拿單 、 所羅門 、
2SAM|5|15|益轄 、 以利書亞 、 尼斐 、 雅非亞 、
2SAM|5|16|以利沙瑪 、 以利雅大 、 以利法列 。
2SAM|5|17|非利士 人聽見 大衛 受膏作 以色列 王， 非利士 眾人就上來尋索 大衛 。 大衛 聽見了，就下到堡壘去。
2SAM|5|18|非利士 人來了，散佈在 利乏音谷 。
2SAM|5|19|大衛 求問耶和華說：「我可以上去攻打 非利士 人嗎？你將他們交在我手裏嗎？」耶和華對 大衛 說：「你可以上去，我必將 非利士 人交在你手裏。」
2SAM|5|20|大衛 來到 巴力‧毗拉心 ，在那裏擊敗了 非利士 人。他說：「耶和華在我面前沖破敵人，如水沖破一樣。」因此他稱那地方為 巴力‧毗拉心 。
2SAM|5|21|非利士 人把偶像拋棄在那裏， 大衛 和他的人拿去了。
2SAM|5|22|非利士 人又上來，散佈在 利乏音谷 。
2SAM|5|23|大衛 求問耶和華；耶和華說：「不要直上，要繞到他們後頭，從桑樹林對面攻打他們。
2SAM|5|24|你聽見桑樹梢上有腳步的聲音，就要急速前去，因為那時耶和華已經出去，在你前頭攻打 非利士 人的軍隊了。」
2SAM|5|25|大衛 就遵照耶和華所吩咐的去做，攻打 非利士 人，從 迦巴 直到 基色 。
2SAM|6|1|大衛 又聚集 以色列 中所有挑選的人，共三萬名。
2SAM|6|2|大衛 起身，和跟隨他的眾百姓前往，要從 巴拉‧猶大 那裏將上帝的約櫃接上來；這約櫃是以坐在二基路伯上萬軍之耶和華的名所命名的。
2SAM|6|3|他們將上帝的約櫃從山岡上 亞比拿達 的家裏抬出來，放在新車上； 亞比拿達 的兒子 烏撒 和 亞希約 趕這新車。
2SAM|6|4|他們將上帝的約櫃從山岡上 亞比拿達 家裏抬出來 ， 亞希約 在約櫃前行走。
2SAM|6|5|大衛 和 以色列 全家在耶和華面前，隨著松木製造的各樣樂器 和琴、瑟、鼓、鈸、鑼跳舞。
2SAM|6|6|到了 拿艮 的禾場，因為牛失前蹄 ， 烏撒 就伸手扶住上帝的約櫃。
2SAM|6|7|耶和華的怒氣向 烏撒 發作；上帝因這冒犯在那裏擊打他，他就死在那裏，在上帝的約櫃旁。
2SAM|6|8|大衛 因耶和華突然衝出撞死 烏撒 就生氣，稱那地方為 毗列斯‧烏撒 ，直到今日。
2SAM|6|9|那日， 大衛 懼怕耶和華，說：「耶和華的約櫃怎可到我這裏來呢？」
2SAM|6|10|於是 大衛 不願將耶和華的約櫃接進 大衛城 他自己的地方，卻轉送到 迦特 人 俄別‧以東 的家中。
2SAM|6|11|耶和華的約櫃停在 迦特 人 俄別‧以東 家中三個月，耶和華賜福給 俄別‧以東 和他的全家。
2SAM|6|12|有人告訴 大衛 王說：「耶和華因約櫃的緣故賜福給 俄別‧以東 的家和一切屬他的。」 大衛 就去，歡歡喜喜地將上帝的約櫃從 俄別‧以東 家中接上來，到 大衛城 裏。
2SAM|6|13|抬耶和華約櫃的人走了六步， 大衛 就獻牛與肥畜為祭。
2SAM|6|14|大衛 穿著細麻布以弗得，在耶和華面前極力跳舞。
2SAM|6|15|這樣， 大衛 和 以色列 全家歡呼吹角，將耶和華的約櫃接了上來。
2SAM|6|16|耶和華的約櫃進 大衛城 的時候， 掃羅 的女兒 米甲 從窗戶裏往外觀看，見 大衛 王在耶和華面前踴躍跳舞，心裏就輕視他。
2SAM|6|17|眾人將耶和華的約櫃請進去，安放在所預備的地方，就是 大衛 為它搭的帳幕中。 大衛 在耶和華面前獻燔祭和平安祭。
2SAM|6|18|大衛 獻完了燔祭和平安祭，就奉萬軍之耶和華的名祝福百姓，
2SAM|6|19|並且分給 以色列 眾人，所有的百姓，無論男女，每人一個餅，一個棗子餅 ，一個葡萄餅。眾人就各自回家去了。
2SAM|6|20|大衛 回去要為家裏的人祝福， 掃羅 的女兒 米甲 出來迎接他，說：「 以色列 王今日有好大的榮耀啊！他今日在臣僕的使女眼前露體，如同一個無賴赤身露體一樣，」
2SAM|6|21|大衛 對 米甲 說：「這是在耶和華面前的。耶和華已揀選我，在你父和你父的全家之上，立我作耶和華百姓 以色列 的君王，所以我在耶和華面前跳舞，
2SAM|6|22|我也必更加卑微，自己看為低賤 。至於你所說的那些使女，她們反而尊重我。」
2SAM|6|23|掃羅 的女兒 米甲 ，直到死的那日沒有孩子。
2SAM|7|1|王住在自己宮中，耶和華使他平靜，不被四圍的仇敵擾亂。
2SAM|7|2|王對 拿單 先知說：「你看，我住在香柏木的宮中，上帝的約櫃卻停在幔子裏。」
2SAM|7|3|拿單 對王說：「你可以完全照你的心意去做，因為耶和華與你同在。」
2SAM|7|4|當夜耶和華的話臨到 拿單 ，說：
2SAM|7|5|「你去對我僕人 大衛 說：『耶和華如此說：你要建造殿宇給我居住嗎？
2SAM|7|6|自從我領 以色列 人從 埃及 上來，直到今日，我未曾住過殿宇，卻在會幕和帳幕中行走。
2SAM|7|7|凡我同 以色列 人所走的地方，我何曾向 以色列 任何一個領袖 ，就是我吩咐牧養我百姓 以色列 的，說過這話：你們為何不給我建造香柏木的殿宇呢？』
2SAM|7|8|現在，你要對我僕人 大衛這樣 說：『萬軍之耶和華如此說：我從羊圈中將你召來，叫你不再牧放羊群，立你作我百姓 以色列 的君王。
2SAM|7|9|你無論往哪裏去，我都與你同在，剪除你所有的仇敵。我必使你得大名，好像世上偉人的名一樣。
2SAM|7|10|我必為我百姓 以色列 選定一個地方，栽植他們，使他們住自己的地方，不再受攪擾；兇惡之子也不像從前那樣苦待他們，
2SAM|7|11|並不像我命令士師治理我百姓 以色列 的日子。我必使你平靜，不受任何仇敵攪擾，並且耶和華應許你，耶和華必為你建立家室。
2SAM|7|12|當你壽數滿足、與你祖先同睡的時候，我必使你身所生的後裔接續你；我也必堅定他的國。
2SAM|7|13|他必為我的名建造殿宇，我必堅定他國度的王位，直到永遠。
2SAM|7|14|我要作他的父，他要作我的子；他若犯了罪，我必用人的杖，用世人的鞭責罰他。
2SAM|7|15|但我的慈愛仍不離開他，像離開在你面前所廢的 掃羅 一樣。
2SAM|7|16|你的家和你的國必在你 面前永遠堅立，你的王位也必堅定，直到永遠。』」
2SAM|7|17|拿單 就按這一切話，照這一切異象告訴 大衛 。
2SAM|7|18|於是 大衛 王進去，坐在耶和華面前，說：「主耶和華啊，我是誰，我的家算甚麼，你竟帶領我到這地步呢？
2SAM|7|19|主耶和華啊，這在你眼中還看為小，你又說到你僕人的家將來的情況。主耶和華啊，這豈是人的常理嗎？
2SAM|7|20|大衛 還有甚麼可以對你說呢？主耶和華啊，你是知道你僕人的。
2SAM|7|21|你行這一切大事，使你的僕人明白，是因你應許的緣故，也照著你的心意。
2SAM|7|22|因此，主耶和華啊，你本為大；照我們耳中一切所聽見的，沒有可比你的，除你以外再沒有上帝。
2SAM|7|23|誰像你的百姓 以色列 呢？上帝親自去救贖世上的一國 ，作自己的子民，顯出他的大名；為了你的地，從列國和他們的神明中，在你親自從埃及贖出來的子民面前，為自己行了大而可畏的事 。
2SAM|7|24|你曾堅立你的百姓 以色列 作你的子民，直到永遠；你－耶和華也作他們的上帝。
2SAM|7|25|現在，耶和華上帝啊，你所應許僕人和僕人家的話，求你堅定，直到永遠；求你照你所說的而行。
2SAM|7|26|願人永遠尊你的名為大，說：『萬軍之耶和華是治理 以色列 的上帝。』這樣，你僕人 大衛 的家必在你面前堅立。
2SAM|7|27|萬軍之耶和華－ 以色列 的上帝啊，因你啟示你的僕人說：『我必為你建立家室』，所以僕人大膽向你如此祈禱。
2SAM|7|28|現在，主耶和華啊，惟有你是上帝！你的話是真實的，你也應許將這福氣賜給僕人。
2SAM|7|29|現在，求你賜福給你僕人的家，可以永存在你面前。主耶和華啊，因為這是你所應許的。願你的福分永遠賜給你僕人的家，使之蒙福！」
2SAM|8|1|此後， 大衛 攻打 非利士 人，制伏了他們。 大衛 從 非利士 人手中奪取了京城的治理權 。
2SAM|8|2|他又攻打 摩押 人，使他們躺臥在地上，用繩來量，量二繩的殺了，量一繩的活著。 摩押 人就臣服 大衛 ，向他進貢。
2SAM|8|3|利合 的兒子 瑣巴 王 哈大底謝 往 幼發拉底河 去，要奪回他的國權， 大衛 就攻打他，
2SAM|8|4|俘擄了他的騎兵一千七百人，步兵二萬人。 大衛 把所有戰馬的蹄筋砍斷，只留下一百輛戰車。
2SAM|8|5|大馬士革 的 亞蘭 人來幫助 瑣巴 王 哈大底謝 ， 大衛 殺了 亞蘭 人二萬二千。
2SAM|8|6|於是 大衛 在 大馬士革 的 亞蘭 設立軍營， 亞蘭 人就臣服 大衛 ，向他進貢。 大衛 無論往哪裏去，耶和華都使他得勝。
2SAM|8|7|大衛奪了 哈大底謝 臣僕擁有的金盾牌，帶到 耶路撒冷 。
2SAM|8|8|大衛 王又從 哈大底謝 的 比他 和 比羅他 二城奪取了許多的銅。
2SAM|8|9|哈馬 王 陀以 聽見 大衛 擊敗 哈大底謝 的全軍，
2SAM|8|10|就派他兒子 約蘭 到 大衛 王那裏，向他請安，為他祝福，因他與 哈大底謝 爭戰，並且擊敗了他；原來 哈大底謝 與 陀以 常常爭戰。 約蘭 手裏帶了金銀銅的器皿來。
2SAM|8|11|大衛 王把這些器皿分別為聖，連同他制伏各國所分別為聖的金銀，獻給耶和華，
2SAM|8|12|就是從 亞蘭 、 摩押 、 亞捫 人、 非利士 人、 亞瑪力 人，以及從 利合 的兒子 瑣巴 王 哈大底謝 所掠之物。
2SAM|8|13|大衛 得了名聲。當他回來的時候，在 鹽谷 擊殺了一萬八千 以東 人。
2SAM|8|14|大衛 在 以東 設立軍營；他在全 以東 設立軍營， 以東 人就都臣服他。 大衛 無論往哪裏去，耶和華都使他得勝。
2SAM|8|15|大衛 作全 以色列 的王，又向眾百姓秉公行義。
2SAM|8|16|洗魯雅 的兒子 約押 作元帥； 亞希律 的兒子 約沙法 作史官；
2SAM|8|17|亞希突 的兒子 撒督 和 亞比亞他 的兒子 亞希米勒 作祭司； 西萊雅 作書記；
2SAM|8|18|耶何耶大 的兒子 比拿雅 管轄 基利提 人和 比利提 人。 大衛 的眾子都作祭司。
2SAM|9|1|大衛 說：「 掃羅 家還有剩下的人沒有？我要因 約拿單 的緣故向他施恩。」
2SAM|9|2|掃羅 家有一個僕人名叫 洗巴 ，有人叫他來到 大衛 那裏。王對他說：「你是 洗巴 嗎？」他說：「僕人是。」
2SAM|9|3|王說：「 掃羅 家還有沒有剩下的人？我要照上帝的慈愛恩待他。」 洗巴 對王說：「還有 約拿單 的一個兒子，雙腿是瘸的。」
2SAM|9|4|王對他說：「他在哪裏？」 洗巴 對王說：「看哪，他在 羅‧底巴 ， 亞米利 的兒子 瑪吉 家裏。」
2SAM|9|5|於是 大衛 王派人去，從 羅‧底巴 ， 亞米利 的兒子 瑪吉 家裏召了他來。
2SAM|9|6|掃羅 的孫子， 約拿單 的兒子 米非波設 來到 大衛 那裏，臉伏於地叩拜。 大衛 說：「 米非波設 ！」 米非波設 說：「看哪，僕人在此。」
2SAM|9|7|大衛 對他說：「你不要懼怕，我必因你父親 約拿單 的緣故向你施恩，把你祖父 掃羅 的一切田地都歸還你，你也可以常與我同席吃飯。」
2SAM|9|8|米非波設 叩拜，說：「你的僕人算甚麼，不過如死狗一般，竟蒙你這樣眷顧！」
2SAM|9|9|王召了 掃羅 的僕人 洗巴 來，對他說：「我已把屬 掃羅 和他的一切家產都賜給你主人的兒子了。
2SAM|9|10|你，你的眾子和僕人要為你主人的兒子耕種田地，把所收穫的拿來供他食用；你主人的兒子 米非波設 卻要常與我同席吃飯。」 洗巴 有十五個兒子和二十個僕人。
2SAM|9|11|洗巴 對王說：「凡我主我王吩咐僕人的，僕人都必遵行。」於是 米非波設 與王 同席吃飯，如王的兒子一樣。
2SAM|9|12|米非波設 有一個小兒子，名叫 米迦 。凡住在 洗巴 家裏的人都作了 米非波設 的僕人。
2SAM|9|13|米非波設 住在 耶路撒冷 ，常與王同席吃飯。他兩腿都是瘸的。
2SAM|10|1|此後， 亞捫 人的王死了，他兒子 哈嫩 接續他作王。
2SAM|10|2|大衛 說：「 哈嫩 的父親 拿轄 怎樣向我施恩，我也要怎樣向 哈嫩 施恩。」於是 大衛 派臣僕為他的父親安慰他。當 大衛 的臣僕到了 亞捫 人的境內，
2SAM|10|3|亞捫 人的領袖對他們的主 哈嫩 說：「 大衛 派人來安慰你，你看他是要尊敬你父親嗎？ 大衛 派臣僕到你這裏，不是為了要窺探偵察，而傾覆這城嗎？」
2SAM|10|4|哈嫩 就抓住 大衛 的臣僕，把他們的鬍鬚剃去一半，又割斷他們下半截的袍子，露出下體，然後放了他們。
2SAM|10|5|有人告訴 大衛 ，他就派人去迎接他們，因為這些人覺得很羞恥。王說：「可以住在 耶利哥 ，等到鬍鬚長出來再回來。」
2SAM|10|6|亞捫 人看到 大衛 憎惡他們，就派人去雇用 伯‧利合 的 亞蘭 人和 瑣巴 的 亞蘭 人，步兵二萬，以及 瑪迦 王的人一千、 陀伯 人一萬二千。
2SAM|10|7|大衛 聽見了，就派 約押 和所有勇猛的軍隊出去。
2SAM|10|8|亞捫 人出來，在城門前擺陣； 瑣巴 與 利合 的 亞蘭 人、 陀伯 人，以及 瑪迦 人另外在郊野擺陣。
2SAM|10|9|約押 看見戰陣對著他前後擺列，就把從 以色列 所有精兵中挑選出來的，擺陣迎戰 亞蘭 人。
2SAM|10|10|他把其餘的兵交在他兄弟 亞比篩 手裏， 亞比篩 就擺陣迎戰 亞捫 人。
2SAM|10|11|約押 對 亞比篩說：「 亞蘭 人若強過我，你就來幫助我； 亞捫 人若強過你，我就去幫助你。
2SAM|10|12|你要剛強，我們要為自己的百姓，為我們上帝的城鎮奮勇。願耶和華照他所看為好的去做！」
2SAM|10|13|於是， 約押 和跟隨他的士兵前進攻打 亞蘭 人； 亞蘭 人在他面前逃跑。
2SAM|10|14|亞捫 人見 亞蘭 人逃跑，他們也在 亞比篩 面前逃跑進城。 約押 就離開 亞捫 人，回 耶路撒冷 去了。
2SAM|10|15|亞蘭 人見自己被 以色列 打敗，就集合起來。
2SAM|10|16|哈大底謝 派人去，把 大河 那邊的 亞蘭 人調來；他們到了 希蘭 ，由 哈大底謝 的將軍 朔法 在他們前面率領。
2SAM|10|17|有人告訴 大衛 ，他就聚集 以色列 眾人過 約旦河 ，來到 希蘭 。 亞蘭 人迎著 大衛 擺陣，與他打仗。
2SAM|10|18|亞蘭 人在 以色列 人面前逃跑。 大衛 殺了 亞蘭 七百輛戰車的士兵，四萬騎兵 ，又擊殺 亞蘭 的將軍 朔法 ，他就死在那裏。
2SAM|10|19|哈大底謝 屬下的諸王見自己被 以色列 打敗，就與 以色列 講和，臣服他們。於是 亞蘭 人害怕，不再幫助 亞捫 人了。
2SAM|11|1|過了一年，正是諸王出戰的時候， 大衛 派 約押 率領臣僕和 以色列 眾人出去。他們打敗 亞捫 人，圍攻 拉巴 。 大衛 仍然留在 耶路撒冷 。
2SAM|11|2|黃昏的時候， 大衛 從床上起來，在王宮的平頂上散步。他從平頂上看見一個婦人沐浴，這婦人容貌非常美麗。
2SAM|11|3|大衛 派人打聽那婦人是誰。有人說：「她不是 以連 的女兒， 赫 人 烏利亞 的妻子 拔示巴 嗎？」
2SAM|11|4|大衛 派使者去把婦人接來；她來到大衛那裏，那時她的月經剛潔淨， 大衛 與她同寢。她就回家去了。
2SAM|11|5|那婦人懷了孕，派人去告訴 大衛 說：「我懷孕了。」
2SAM|11|6|大衛 派人告訴 約押 ：「你派 赫 人 烏利亞 到我這裏來。」 約押 就派 烏利亞 到 大衛 那裏。
2SAM|11|7|烏利亞 來到 大衛那裏， 大衛 問 約押 好，也問士兵好，又問戰爭的情況。
2SAM|11|8|大衛 對 烏利亞 說：「下到你家去，洗洗腳吧！」 烏利亞 出了王宮，隨後王送他一份禮物。
2SAM|11|9|烏利亞 卻和他主人所有的僕人一同睡在王宮門口，沒有下到他家去。
2SAM|11|10|有人告訴 大衛 說：「 烏利亞 沒有下到他的家。」 大衛 就對 烏利亞 說：「你不是從遠路上來嗎？為甚麼不下到你家去呢？」
2SAM|11|11|烏利亞 對 大衛 說：「約櫃， 以色列 和 猶大 都留在棚裏，我主 約押 和我主的僕人都在田野安營，我豈可回家吃喝，與妻子同房呢？我指著王和王的性命起誓：『我絕不做這事！』」
2SAM|11|12|大衛 對 烏利亞 說：「你今日仍留在這裏，明日我打發你去。」於是 烏利亞 那日留在 耶路撒冷 。次日，
2SAM|11|13|大衛 召了 烏利亞 來，叫他在自己面前吃喝，使他喝醉。黃昏的時候， 烏利亞 出去，躺臥在自己的床上；與他主的僕人在一起，並沒有下到他的家去。
2SAM|11|14|早晨， 大衛 寫信給 約押 ，交 烏利亞 親手帶去。
2SAM|11|15|他在信內寫著說：「要派 烏利亞 到戰爭激烈的前線去，然後你們撤退離開他，使他被擊殺而死。」
2SAM|11|16|約押 偵察城的時候，知道敵人哪裏有勇士，就派 烏利亞 到那地方。
2SAM|11|17|城裏的人出來和 約押 打仗， 大衛 的僕人中有幾個士兵被殺， 赫 人 烏利亞 也死了。
2SAM|11|18|於是， 約押 派人去將戰爭的一切事奏告 大衛 ，
2SAM|11|19|又吩咐使者說：「你把戰爭的一切事對王說完了，
2SAM|11|20|王若發怒，對你說：『你們打仗為甚麼挨近城呢？豈不知敵人會從城牆上射箭嗎？
2SAM|11|21|從前擊殺 耶路比設 的兒子 亞比米勒 的是誰呢？豈不是一個婦人從城牆上拋下一塊上磨石來，打在他身上，他就死在 提備斯 嗎？你們為甚麼挨近城牆呢？』你就說：『你的僕人 赫 人 烏利亞 也死了。』」
2SAM|11|22|使者就去，照著 約押 所吩咐的一切話來奏告 大衛 。
2SAM|11|23|使者對 大衛 說：「敵人強過我們，出到郊外攻打我們，我們把他們趕回到城門口。
2SAM|11|24|弓箭手從城牆上射你的僕人，射死幾個王的僕人，你的僕人 赫 人 烏利亞 也死了。」
2SAM|11|25|大衛 向使者說：「你對 約押 這樣說：『不要為這事難過，因為刀劍可能吞滅這人或那人。你只管竭力攻城，將城傾覆。』你要勉勵 約押 。」
2SAM|11|26|烏利亞 的妻聽見丈夫 烏利亞 死了，就為丈夫哀哭。
2SAM|11|27|居喪的日子過了， 大衛 派人把她接到宮裏，她就作了 大衛 的妻子，給 大衛 生了一個兒子。但 大衛 做的這事，耶和華的眼中看為惡。
2SAM|12|1|耶和華差遣 拿單 到 大衛 那裏。 拿單 到了他那裏，對他說：「在一座城裏有兩個人，一個是富翁，一個是窮人。
2SAM|12|2|富翁有極多的牛群羊群；
2SAM|12|3|窮人除了所買來養活的一隻小母羊之外，一無所有。小羊在他家裏和他兒女一同長大，吃他所吃的，喝他所喝的，睡在他懷中，在他看來如同女兒一樣。
2SAM|12|4|有一客人來到這富翁那裏，富翁捨不得從自己的牛群羊群中取一隻招待來到他那裏的旅客，卻取了窮人的小母羊，招待來到他那裏的人。」
2SAM|12|5|大衛 就非常惱怒那人，對 拿單 說：「我指著永生的耶和華起誓，做這事的人該死！
2SAM|12|6|他必須償還小母羊四倍，因為他做這事，沒有憐憫的心。」
2SAM|12|7|拿單 對 大衛 說：「你就是那人！耶和華－ 以色列 的上帝如此說：『我膏你作 以色列 的王，我救你脫離 掃羅 的手；
2SAM|12|8|我將你主人的家業賜給你，將你主人的妃嬪交在你懷裏，又將 以色列 和 猶大 家賜給你；若還嫌少，我也會如此這般加倍賜給你。
2SAM|12|9|你為甚麼藐視耶和華的命令，做他眼中看為惡的事呢？你用刀擊殺 赫 人 烏利亞 ，又娶了他的妻子為妻，借 亞捫 人的刀殺死他。
2SAM|12|10|現在刀劍必永不離開你的家，因你藐視我，娶了 赫 人 烏利亞 的妻子為妻。』
2SAM|12|11|耶和華如此說：『看哪，我必從你家中興起災禍攻擊你；我必在你眼前把你的妃嬪賜給你身邊的人，他要在光天化日下與你的妃嬪同寢。
2SAM|12|12|你在暗中做那事，我卻要在 以色列 眾人面前，在日光之下做這事。』」
2SAM|12|13|大衛 對 拿單 說：「我得罪耶和華了！」 拿單 說：「耶和華已經除去你的罪，你必不至於死。
2SAM|12|14|只是在這事上，你大大藐視耶和華 ，因此，你生的孩子必定要死。」
2SAM|12|15|拿單 就回家去了。 耶和華擊打 烏利亞 的妻子為 大衛 生的孩子，他就得了重病。
2SAM|12|16|大衛 為這孩子懇求上帝。 大衛 刻苦禁食，到裏面去，躺在地上過夜。
2SAM|12|17|他家中的老臣來到他旁邊，要把他從地上扶起來，他卻不肯，也不同他們吃飯。
2SAM|12|18|到第七日，孩子死了。 大衛 的臣僕不敢告訴他孩子死了，因他們說：「看哪，孩子還活著的時候，我們勸他，他尚且不聽我們的話，我們怎麼能告訴他孩子死了，讓他做出不好的事呢？」
2SAM|12|19|大衛 見臣僕彼此低聲說話，就知道孩子死了。他問臣僕說：「孩子死了嗎？」他們說：「死了。」
2SAM|12|20|大衛 就從地上起來，沐浴，抹膏，換了衣服，進耶和華的殿敬拜。然後他回宮，吩咐人為他擺飯，他就吃了。
2SAM|12|21|臣僕對他說：「你所做的是甚麼事呢？孩子活著的時候，你為他禁食哭泣；孩子死了，你卻起來吃飯。」
2SAM|12|22|大衛 說：「孩子還活著，我禁食哭泣，因為我想，或許耶和華憐憫我，會讓孩子活下來。
2SAM|12|23|現在孩子死了，我何必禁食呢？我能使他回來嗎？我必往他那裏去，他卻不能回到我這裏來。」
2SAM|12|24|大衛 安慰他的妻子 拔示巴 ，與她同房，她就生了兒子，給他起名叫 所羅門 。耶和華喜愛他，
2SAM|12|25|就藉 拿單 先知賜他一個名字，叫 耶底底亞 ；這是為了耶和華的緣故。
2SAM|12|26|約押 攻打 亞捫 人的 拉巴 ，攻佔了京城。
2SAM|12|27|約押 派使者到 大衛 那裏，說：「我攻打 拉巴 ， 也攻佔了水城。
2SAM|12|28|現在你要召集其餘的軍兵，安營圍攻這城，攻佔它，免得我攻佔這城，人就以我的名叫這城。」
2SAM|12|29|於是 大衛 召集全軍，往 拉巴 去攻城，就攻佔了它。
2SAM|12|30|他也奪了 米勒公 頭上所戴的冠冕，其上的金子重一他連得，又嵌著寶石。這冠冕就戴在 大衛 頭上。 大衛 又從城裏奪了許多財物，
2SAM|12|31|把城裏的百姓拉出來，叫他們用鋸，用鐵耙，用鐵斧做工，派他們在磚窯中服役； 大衛 待 亞捫 各城的居民都是如此。於是， 大衛 和全軍都回 耶路撒冷 去了。
2SAM|13|1|後來發生了一件事。 大衛 的兒子 押沙龍 有一個美貌的妹妹，名叫 她瑪 。 大衛 的兒子 暗嫩 愛上了她。
2SAM|13|2|暗嫩 為他妹妹 她瑪 苦戀成疾，因為 她瑪 還是處女， 暗嫩 眼看難以向她行事。
2SAM|13|3|暗嫩 有一個密友，名叫 約拿達 ，是 大衛 長兄 示米亞 的兒子。這 約拿達 為人極其狡猾。
2SAM|13|4|他對 暗嫩 說：「王的兒子啊，你何不告訴我，為何你一天比一天憔悴呢？」 暗嫩 對他說：「我愛上了我兄弟 押沙龍 的妹妹 她瑪 。」
2SAM|13|5|約拿達 對他說：「你躺在床上裝病，等你父親來看你，就對他說：『請讓我妹妹 她瑪 來，給我東西吃，在我眼前預備食物，使我可以看見，好從她手裏接過來吃。』」
2SAM|13|6|於是 暗嫩 躺著裝病，王來看他。 暗嫩 對王說：「請讓我妹妹 她瑪 來，在我眼前為我做兩個餅，我好從她手裏接過來吃。」
2SAM|13|7|大衛 就派人去宮裏，到 她瑪 那裏，說：「你到你哥哥 暗嫩 的屋裏去，為他預備食物。」
2SAM|13|8|她瑪 就到她哥哥 暗嫩 的屋裏，那時 暗嫩 正躺著。 她瑪 拿了麵團揉麵，在他眼前做餅，把餅烤熟了。
2SAM|13|9|她瑪 拿了鍋子，在他面前把餅倒出來，他卻不肯吃。 暗嫩 說：「每一個人都離開我，出去吧！」眾人就都離開他，出去了。
2SAM|13|10|暗嫩 對 她瑪 說：「你把食物拿進臥房，我好從你手裏接過來吃。」 她瑪 就把所做的餅拿進臥房，到她哥哥 暗嫩 那裏。
2SAM|13|11|她瑪 上前去給他吃，他就拉住 她瑪 ，對她說：「我妹妹，你來與我同寢。」
2SAM|13|12|她瑪 對他說：「哥哥，不可以！不要玷辱我！ 以色列 中不可以這樣做，你不要做這醜事！
2SAM|13|13|我蒙受恥辱，該往那裏去呢？至於你，你在 以色列 中也成了一個愚頑人。現在你可以求王，他必不禁止我歸你。」
2SAM|13|14|但 暗嫩 不肯聽她的話，因他比她更有力，就玷辱她，與她同寢。
2SAM|13|15|隨後， 暗嫩 極其恨她，恨她的心比先前愛她的心更甚，就對她說：「你起來，去吧！」
2SAM|13|16|她瑪 對 暗嫩 說：「不要這樣！你趕我出去的這惡比你剛才向我所做的更嚴重！」但 暗嫩 不肯聽她，
2SAM|13|17|就叫伺候自己的僕人來，說：「把這女子從我這裏趕出去！她一出去，你就閂上門。」
2SAM|13|18|那時 她瑪 穿著彩衣，因為沒有出嫁的公主都穿這樣的外袍。 暗嫩 的僕人把她趕出去，她一出去，僕人就閂上門。
2SAM|13|19|她瑪 把灰塵撒在頭上，撕裂所穿的彩衣，以手抱頭，一面走一面哭喊。
2SAM|13|20|她胞兄 押沙龍 對她說：「你哥哥 暗嫩 與你親近了嗎？妹妹，現在暫且不要作聲，他是你的哥哥，不要把這事放在心上。」 她瑪 就孤孤單單地住在她胞兄 押沙龍 的家裏。
2SAM|13|21|大衛 王聽見這一切的事，就非常憤怒。
2SAM|13|22|押沙龍 卻不和 暗嫩 說好說歹；因為 暗嫩 玷辱他妹妹 她瑪 ，所以 押沙龍 恨惡他。
2SAM|13|23|過了二年，有人在靠近 以法蓮 的 巴力‧夏瑣 為 押沙龍 剪羊毛。 押沙龍 請了王所有的兒子來。
2SAM|13|24|押沙龍 來到王那裏，說：「看哪，有人正為你的僕人剪羊毛，請王和王的臣僕與你的僕人同去。」
2SAM|13|25|王對 押沙龍 說：「不，我兒，我們不必都去，免得成了你的負擔。」 押沙龍 再三請王，王仍是不肯去，只為他祝福。
2SAM|13|26|押沙龍 說：「王若不去，請讓我哥哥 暗嫩 與我們同去。」王對他說：「為何要他與你同去呢？」
2SAM|13|27|押沙龍 再三求王，王就派 暗嫩 和王所有的兒子與他同去。
2SAM|13|28|押沙龍 吩咐僕人說：「你們注意， 暗嫩 開懷暢飲的時候，我對你們說擊殺 暗嫩 ，你們就殺他。不要懼怕，這不是我吩咐你們的嗎？你們要剛強，作勇士！」
2SAM|13|29|押沙龍 的僕人就照 押沙龍 所吩咐的，向 暗嫩 行了。王所有的兒子都起來，各人騎上騾子逃跑了。
2SAM|13|30|他們還在路上，就有風聲傳到 大衛 那裏，說：「 押沙龍 擊殺了王所有的兒子，沒有留下一個。」
2SAM|13|31|王就起來，撕裂衣服，躺在地上。王的臣僕全都撕裂衣服，站在旁邊。
2SAM|13|32|大衛 的長兄 示米亞 的兒子 約拿達 說：「我主，不要以為他們把所有的年輕人，就是王的兒子都殺了，只有 暗嫩 一個人死了。自從 暗嫩 玷辱了 押沙龍 的妹妹 她瑪 那日， 押沙龍 已經決定這事了。
2SAM|13|33|現在，我主我王，不要把這事放在心上，以為王所有的兒子都死了。其實，只有 暗嫩 一人死了。」
2SAM|13|34|押沙龍 逃跑了。守望的年輕人舉目觀看，看哪，有許多人從 何羅念 山坡的路上來。
2SAM|13|35|約拿達 對王說：「看哪，王的兒子都來了，正如你僕人所說的，事情就這樣發生了。」
2SAM|13|36|話剛說完，看哪，王的兒子都到了，放聲大哭。王和他的眾臣僕也都號咷痛哭。
2SAM|13|37|押沙龍 逃到 亞米忽 的兒子 基述 王 達買 那裏去了。 大衛 天天為他兒子悲哀。
2SAM|13|38|押沙龍 逃到 基述 去了，在那裏住了三年。
2SAM|13|39|王想要出去對付 押沙龍 的心化解了 ，因為王對 暗嫩 之死這事已經得了安慰。
2SAM|14|1|洗魯雅 的兒子 約押 知道王心裏想念 押沙龍 。
2SAM|14|2|他派人往 提哥亞 去，從那裏叫了一個有智慧的婦人來，對她說：「請你裝作居喪的人，穿上喪服，不用膏抹身，裝作為死者悲哀多日的婦人。
2SAM|14|3|你到王那裏，對王如此如此說。」於是 約押 把當說的話放在她口中。
2SAM|14|4|提哥亞 婦人到王面前 ，臉伏於地叩拜，說：「王啊，求你拯救！」
2SAM|14|5|王對她說：「你有甚麼事呢？」她說：「我實在是個寡婦，我丈夫死了。
2SAM|14|6|婢女有兩個兒子，二人在田間打架，沒有人從中勸解，一個擊殺另一個，把他打死了。
2SAM|14|7|看哪，全家族都起來攻擊婢女，說：『把那打死兄弟的交出來，我們好處死他，為他所打死的兄弟償命，滅絕那承受家業的。』這樣，他們要把我剩下的炭火滅盡，不給我丈夫留名或留後在地面上。」
2SAM|14|8|王對婦人說：「你回家去吧！我必為你下個命令。」
2SAM|14|9|提哥亞 婦人又對王說：「我主我王，願這罪孽歸我和我的父家，與王和王的位無關。」
2SAM|14|10|王說：「有人說話難為你，你就帶他到我這裏來，他必不再攪擾你。」
2SAM|14|11|婦人說：「願王對耶和華－你的上帝發誓，不許報血仇的人施行毀滅，免得他們滅絕我的兒子。」王說：「我指著永生的耶和華起誓：你的兒子連一根頭髮也不致落在地上。」
2SAM|14|12|婦人說：「求我主我王容許婢女再說一句話。」王說：「你說吧！」
2SAM|14|13|婦人說：「王為何起意做這事，要害上帝的百姓呢？王不使那逃亡的人回來，王說這話就證實自己錯了！
2SAM|14|14|我們都必死，如同水潑在地上，不能收回。上帝不會讓人不死，但仍設法 使逃亡的人不致成為趕出、回不來的人。
2SAM|14|15|現在我來將這話告訴我主我王，是因百姓使我懼怕。婢女想：『不如告訴王，或者王會成就使女所求的。
2SAM|14|16|人要把我和我兒子從上帝的地業上一同除滅，王必應允救使女脫離他的手。』
2SAM|14|17|婢女想：『我主我王的話必安慰我』；因為我主我王能辨別是非，如同上帝的使者一樣。惟願耶和華－你的上帝與你同在！」
2SAM|14|18|王回答婦人說：「我問你一句話，你一點也不可瞞我。」婦人說：「我主我王，請說。」
2SAM|14|19|王說：「這一切莫非是 約押 的手指使你的嗎？」婦人回答說：「我敢在我主我王面前起誓：我主我王所說的一切不偏左右，這是王的僕人 約押 吩咐我的，這一切話是他放在婢女口中的。
2SAM|14|20|王的僕人 約押 做這事，為要扭轉局面。我主的智慧卻如上帝使者的智慧，能知地上一切的事。」
2SAM|14|21|王對 約押 說：「看哪，我應允這事。你去，把那年輕人 押沙龍 帶回來。」
2SAM|14|22|約押 臉伏於地叩拜，為王祝福，說：「王既應允僕人這件事，僕人今日知道在我主我王眼前蒙恩寵了。」
2SAM|14|23|於是 約押 起身往 基述 去，把 押沙龍 帶回 耶路撒冷 。
2SAM|14|24|王說：「讓他回自己的家去，不要來見我的面。」 押沙龍 就回自己的家去，沒有見王的面。
2SAM|14|25|全 以色列 中，無人像 押沙龍 那樣俊美，得人稱讚，從腳底到頭頂毫無瑕疵。
2SAM|14|26|他的頭髮很重，每到年底剪髮一次，所剪下來的，按王的秤稱一稱，重二百舍客勒。
2SAM|14|27|押沙龍 生了三個兒子，一個女兒。女兒名叫 她瑪 ，是個容貌美麗的女子。
2SAM|14|28|押沙龍 住在 耶路撒冷 ，足足有二年沒有見王的面。
2SAM|14|29|押沙龍 派人去叫 約押 來，要託他到王那裏去， 約押 卻不肯來。 押沙龍 第二次派人去叫他，他仍不肯來。
2SAM|14|30|於是 押沙龍 對僕人說：「你們看， 約押 有一塊田靠近我的田，其中有大麥，你們去放火把它燒了。」 押沙龍 的僕人就去放火燒了那田。
2SAM|14|31|於是 約押 起來，到了 押沙龍 家裏，對他說：「你的僕人為何放火燒我的田呢？」
2SAM|14|32|押沙龍 對 約押 說：「看哪，我派人去請你來，好託你到王那裏去，說：『我為何從 基述 回來呢？我仍在那裏比較好。』現在讓我去見王的面；我若有罪孽，就任憑王殺了我吧。」
2SAM|14|33|於是 約押 到王那裏，奏告王，王就叫 押沙龍 來。 押沙龍 到王那裏，在王面前臉伏於地，王就親吻 押沙龍 。
2SAM|15|1|此後， 押沙龍 為自己預備車馬，又派五十人在他前頭奔跑。
2SAM|15|2|押沙龍 常常早晨起來，站在城門的路旁，任何人有爭訟要去求王判決， 押沙龍 就叫他過來，說：「你是哪一城的人？」他說：「僕人是 以色列 某支派的人。」
2SAM|15|3|押沙龍 就對他說：「看，你的案件合情合理，無奈王沒有委派人聽你申訴。」
2SAM|15|4|押沙龍 又說：「恨不得我作這地的審判官！ 凡有爭訟的人可以到我這裏來，我必秉公判斷。」
2SAM|15|5|若有人近前來要拜 押沙龍 ， 押沙龍 就伸手拉住他，親吻他。
2SAM|15|6|以色列 中，凡到王那裏求判決的， 押沙龍 都這麼做。這樣， 押沙龍 暗中贏得了 以色列 人的心。
2SAM|15|7|過了四年 ， 押沙龍 對王說：「求你准我往 希伯崙 去，還我向耶和華所許的願。
2SAM|15|8|因為僕人住在 亞蘭 的 基述 時，曾許願說：『耶和華若使我再回 耶路撒冷 ，我必事奉他 。』」
2SAM|15|9|王對他說：「你平安地去吧！」 押沙龍 就動身，往 希伯崙 去了。
2SAM|15|10|押沙龍 派密使走遍 以色列 各支派，說：「你們一聽見角聲就說：『 押沙龍 在 希伯崙 作王了！』」
2SAM|15|11|押沙龍 在 耶路撒冷 請了二百人與他同去，都是誠心誠意去的，一點也不知道實情。
2SAM|15|12|押沙龍 獻祭的時候，派人去把 大衛 的謀士， 基羅 人 亞希多弗 從他本城 基羅 請來 。於是叛亂越發強大，因為隨從 押沙龍 的百姓日漸增多。
2SAM|15|13|報信的人來到 大衛 那裏，說：「 以色列 人的心都歸向 押沙龍 了！」
2SAM|15|14|大衛 就對 耶路撒冷 所有跟隨他的臣僕說：「起來，我們逃吧！否則，我們來不及逃避 押沙龍 。要快點離開，免得他很快追上我們，加害於我們，用刀擊殺城裏的人。」
2SAM|15|15|王的臣僕對王說：「我主我王所決定的一切，看哪，僕人都願遵行。」
2SAM|15|16|於是王出去了，他的全家都跟隨他，但留下十個妃嬪看守宮殿。
2SAM|15|17|王出去，眾百姓都跟隨他；到了最後一座屋子 ，他們就停下來。
2SAM|15|18|王的眾臣僕都在他旁邊過去。 基利提 人、 比利提 人，和從 迦特 跟隨王來的六百個 迦特 人，也都在王面前過去。
2SAM|15|19|王對 迦特 人 以太 說：「你是外邦人，從你本地逃來的，為甚麼與我們同去呢？你回去留在新王那裏吧！
2SAM|15|20|你昨天才到，我今日怎好叫你與我們一同流亡，而我卻要到處飄流呢？回去吧，你帶你的弟兄回去吧！願主用慈愛信實待你 。」
2SAM|15|21|以太 回答王說：「我指著永生的耶和華起誓，又敢在王面前起誓：無論生死，王在哪裏，你的僕人也必在哪裏。」
2SAM|15|22|大衛 對 以太 說：「去，過去吧！」於是 迦特 人 以太 帶著所有跟隨他的人和孩子過去了。
2SAM|15|23|眾百姓過去時，當地的人全都放聲大哭。王過了 汲淪溪 ，眾百姓就往曠野的路上去了。
2SAM|15|24|看哪， 撒督 和所有抬上帝約櫃的 利未 人也一同來了。他們將上帝的約櫃放下， 亞比亞他 上來 ，直到眾百姓從城裏出來走過去為止。
2SAM|15|25|王對 撒督 說：「你將上帝的約櫃請回城去。我若在耶和華眼前蒙恩，他必使我回來，再見到約櫃和他的居所。
2SAM|15|26|倘若他說：『我不喜愛你』；我在這裏，就照他眼中看為好的待我！」
2SAM|15|27|王對 撒督 祭司說：「你不是先見嗎？你可以平安地回城，你兒子 亞希瑪斯 和 亞比亞他 的兒子 約拿單 ，你們二人的兒子可以與你們同去。
2SAM|15|28|看，我在曠野的渡口那裏等，直到你們來報信給我。」
2SAM|15|29|於是 撒督 和 亞比亞他 將上帝的約櫃請回 耶路撒冷 ，他們就留在那裏。
2SAM|15|30|大衛 蒙頭赤腳走上 橄欖山 的斜坡，一面上一面哭。所有跟隨他的百姓也都各自蒙頭哭著上去；
2SAM|15|31|有人告訴 大衛 說 ：「 亞希多弗 也在叛黨之中，隨從 押沙龍 。」 大衛 說：「耶和華啊，求你使 亞希多弗 的計謀變為愚拙！」
2SAM|15|32|大衛 到了山頂，敬拜上帝的地方，看哪， 亞基 人 戶篩 衣服撕裂，頭蒙灰塵來迎見他。
2SAM|15|33|大衛 對他說：「你若與我一同過去，必拖累我；
2SAM|15|34|你若回城去，對 押沙龍 說：『王啊，我願作你的僕人。我向來作你父親的僕人，現在我也願意作你的僕人。』你就可以為我破壞 亞希多弗 的計謀。
2SAM|15|35|撒督 和 亞比亞他 二位祭司豈不都在你那裏嗎？你在王宮裏聽見甚麼，就要告訴 撒督 和 亞比亞他 二位祭司。
2SAM|15|36|看哪， 撒督 的兒子 亞希瑪斯 ， 亞比亞他 的兒子 約拿單 ，也跟二位祭司在那裏。凡你們所聽見的事，可以託這二人來向我報告。」
2SAM|15|37|於是， 大衛 的朋友 戶篩 進了城， 押沙龍 也進了 耶路撒冷 。
2SAM|16|1|大衛 剛過山頂，看哪， 米非波設 的僕人 洗巴 拉著裝好鞍子的兩匹驢，驢上馱著二百個麵餅，一百個葡萄餅，一百個夏天的果餅，一皮袋酒來迎接他。
2SAM|16|2|王對 洗巴 說：「你的這些東西是甚麼意思呢？」 洗巴 說：「驢是給王的家眷騎的，麵餅和夏天的果餅是給年輕人吃的，酒是給在曠野疲乏的人喝的。」
2SAM|16|3|王說：「你主人的兒子在哪裏呢？」 洗巴 對王說：「看哪，他留在 耶路撒冷 ，因他說：『 以色列 家今日必將我父的國歸還我。』」
2SAM|16|4|王對 洗巴 說：「看哪，凡屬 米非波設 的都是你的了。」 洗巴 說：「我叩拜我主我王，願我在你眼前蒙恩寵。」
2SAM|16|5|大衛 王到了 巴戶琳 ，看哪，有一個人從那裏出來，是 掃羅 家族中 基拉 的兒子，名叫 示每 。他一面走一面咒罵，
2SAM|16|6|又向 大衛 王和王的眾臣僕扔石頭；眾百姓和勇士都在王的左右。
2SAM|16|7|示每 這樣咒罵說：「你這好流人血的，你這無賴，滾吧！滾吧！
2SAM|16|8|你流了 掃羅 全家的血，接續他作王，耶和華把這罪歸在你身上。耶和華將這國交在你兒子 押沙龍 的手中。看哪，你咎由自取，因為你是好流人血的人。」
2SAM|16|9|洗魯雅 的兒子 亞比篩 對王說：「這死狗為何咒罵我主我王呢？讓我過去，割下他的頭來。」
2SAM|16|10|王說：「 洗魯雅 的兒子，我與你們有何相干呢？他這樣咒罵是因耶和華吩咐他：『你要咒罵 大衛 。』如此，誰敢說：『你為甚麼這樣做呢？』」
2SAM|16|11|大衛 又對 亞比篩 和眾臣僕說：「看哪，我親生的兒子尚且尋索我的性命，何況現在這 便雅憫 人呢？由他咒罵吧！因為這是耶和華吩咐他的。
2SAM|16|12|或者耶和華見我遭難 ，因我今日被這人咒罵而向我施恩。」
2SAM|16|13|於是 大衛 和他的人在路上走。 示每 走在 大衛 對面的山坡，一面走一面咒罵，又向他扔石頭，揚起塵土。
2SAM|16|14|王和跟隨他的眾百姓來了，非常疲乏，就在那裏歇息。
2SAM|16|15|押沙龍 和 以色列 眾百姓來到 耶路撒冷 ， 亞希多弗 也與他同來。
2SAM|16|16|大衛 的朋友 亞基 人 戶篩 來到 押沙龍 那裏，對他說：「願王萬歲！願王萬歲！」
2SAM|16|17|押沙龍 對 戶篩 說：「你這樣做是忠誠對待你的朋友嗎？為甚麼不與你的朋友同去呢？」
2SAM|16|18|戶篩 對 押沙龍 說：「不，誰是耶和華和這百姓，以及 以色列 眾人所揀選的，我必歸順他，留在他那裏。
2SAM|16|19|再者，我當服事誰呢？豈不是前王的兒子嗎？我怎樣服事你父親，也必照樣服事你。」
2SAM|16|20|押沙龍 對 亞希多弗 說：「你們出個主意，我們該怎麼做？」
2SAM|16|21|亞希多弗 對 押沙龍 說：「你父親所留下看守宮殿的妃嬪，你可以與她們親近。 以色列 眾人聽見你敢惹你父親憎惡你，凡歸順你人的手就更堅強了。」
2SAM|16|22|於是他們為 押沙龍 在屋頂上支搭帳棚， 押沙龍 就在 以色列 眾人眼前，與他父親的妃嬪親近。
2SAM|16|23|那時 亞希多弗 所出的主意好像人從上帝求問得來的話一樣；他給 大衛 ，給 押沙龍 所出的一切主意，都是這樣。
2SAM|17|1|亞希多弗 對 押沙龍 說：「請讓我挑選一萬二千人，今夜起身追趕 大衛 。
2SAM|17|2|我必趁他疲乏手軟的時候追上他，使他驚惶。跟隨他的眾百姓必都逃跑，我就只殺王一個人。
2SAM|17|3|我必使眾百姓都歸順你，正如眾人歸順你所追殺的人一樣 ，眾百姓就都平安無事了。」
2SAM|17|4|這話在 押沙龍 和 以色列 眾長老的眼中都看為好。
2SAM|17|5|押沙龍 說：「把 亞基 人 戶篩 也召來，我們也要聽他怎麼說。」
2SAM|17|6|戶篩 到了 押沙龍 那裏， 押沙龍 向他說：「 亞希多弗 說了這樣的話，我們要照他的話做嗎？若不可，你就說吧！」
2SAM|17|7|戶篩 對 押沙龍 說：「 亞希多弗 這次所出的主意不好。」
2SAM|17|8|戶篩 又說：「你知道，你父親和他的人都是勇士，他們心裏惱怒，如同田野中失去小熊的母熊一樣；而且你父親是個戰士，必不和百姓一同住宿。
2SAM|17|9|看哪，他現今或藏在一個坑中或在別處，若我們 有人首先被殺，聽見的必說：『跟隨 押沙龍 的百姓被殺了。』
2SAM|17|10|雖有勇士膽大如獅子，他的心也必定融化，因為全 以色列 都知道你父親是英雄，跟隨他的人都是勇士。
2SAM|17|11|依我之計，要把如同海邊的沙那樣多的 以色列 眾人，從 但 直到 別是巴 ，聚集到你這裏來，由你親自率領他們出戰。
2SAM|17|12|我們到他那裏，在任何地方遇見他，就突然臨到他，如同露水滴在泥土上。這樣，他和所有跟隨他的人，一個也不留。
2SAM|17|13|他若撤退到一座城， 以色列 眾人必帶繩子去那城，把城拉到河裏，甚至連一塊小石子也找不到。」
2SAM|17|14|押沙龍 和 以色列 眾人都說：「 亞基 人 戶篩 的計謀比 亞希多弗 的更好！」這是因為耶和華定意破壞 亞希多弗 的良謀，為的是耶和華要降禍給 押沙龍 。
2SAM|17|15|戶篩 對 撒督 和 亞比亞他 二位祭司說：「 亞希多弗 為 押沙龍 和 以色列 的長老出的主意是如此如此，我出的主意是如此如此。
2SAM|17|16|現在你們要急速派人去告訴 大衛 說：『今夜不可在曠野的渡口住宿，務要過河，免得王和所有跟隨他的百姓都被吞滅。』」
2SAM|17|17|約拿單 和 亞希瑪斯 在 隱‧羅結 等候，不敢進城，恐怕被人看見。有一個婢女出來，把這話告訴他們，他們就去報信給 大衛 王。
2SAM|17|18|然而有一個僮僕看見他們，就去告訴 押沙龍 。他們二人急忙離開，跑到 巴戶琳 一個人的家裏。那人院中有一口井，他們就下到那裏。
2SAM|17|19|那家的婦人用蓋蓋上井口，又在上頭鋪上碎麥，事情就沒有洩漏。
2SAM|17|20|押沙龍 的僕人來到婦人的家，說：「 亞希瑪斯 和 約拿單 在哪裏？」婦人對他們說：「他們過了河了。」僕人搜尋，卻找不著，就回 耶路撒冷 去了。
2SAM|17|21|他們走後，二人從井裏上來，去告訴 大衛 王。他們對 大衛 說：「 亞希多弗 出這樣的主意要害你，你們起來，快快過河。」
2SAM|17|22|於是 大衛 和所有跟隨他的百姓都起來，過 約旦河 。到了天亮，無一人不過 約旦河 的。
2SAM|17|23|亞希多弗 見他的計謀不被接納，就備上驢，動身歸回本城，到了自己的家。他留下遺囑給他的家，就上吊死了，葬在他父親的墳墓裏。
2SAM|17|24|大衛 到了 瑪哈念 ， 押沙龍 和跟隨他的 以色列 眾人也都過了 約旦河 。
2SAM|17|25|押沙龍 立 亞瑪撒 作元帥，取代 約押 。 亞瑪撒 是 以實瑪利 人 以特拉 的兒子。 以特拉 曾與 拿轄 的女兒 亞比該 親近；這 亞比該 與 約押 的母親 洗魯雅 是姊妹。
2SAM|17|26|押沙龍 和 以色列 人安營在 基列 地。
2SAM|17|27|大衛 到了 瑪哈念 ， 亞捫 族的 拉巴 人 拿轄 的兒子 朔比 ， 羅‧底巴 人 亞米利 的兒子 瑪吉 ，來自 羅基琳 的 基列 人 巴西萊 ，
2SAM|17|28|帶著被褥、盆、瓦器，還有小麥、大麥、麥麵、烤熟的穀穗、豆子、紅豆、炒豆、
2SAM|17|29|蜂蜜、奶油、綿羊、奶餅，供給 大衛 和跟隨他的人吃，因為他們想：「百姓在曠野中，必定又飢渴又疲乏。」
2SAM|18|1|大衛 數點跟隨他的百姓，立千夫長、百夫長率領他們。
2SAM|18|2|大衛 把軍兵分為三隊 ：三分之一在 約押 手下，三分之一在 洗魯雅 的兒子 約押 弟弟 亞比篩 手下，三分之一在 迦特 人 以太 手下。王對軍兵說：「我必與你們一同出戰。」
2SAM|18|3|軍兵卻說：「你不可出戰。若是我們逃跑，敵人不會把心放在我們身上；我們陣亡一半，敵人也不會把心放在我們身上。但現在你一人抵過我們萬人，所以你最好留在城裏支援我們。」
2SAM|18|4|王對他們說：「你們看怎樣好，我就怎樣做。」於是王站在城門旁，所有的軍兵成百成千地挨次出戰去了。
2SAM|18|5|王囑咐 約押 、 亞比篩 、 以太 說：「你們要為我的緣故寬待那年輕人 押沙龍 。」王為 押沙龍 的事囑咐眾將領的話，所有的軍兵都聽見了。
2SAM|18|6|軍兵出到田野迎戰 以色列 ，在 以法蓮 的樹林裏交戰。
2SAM|18|7|在那裏， 以色列 百姓敗在 大衛 的臣僕面前。那日在那裏陣亡的很多，共有二萬人。
2SAM|18|8|戰爭蔓延到整個地面，那日被樹林吞噬的軍兵比被刀劍吞噬的更多。
2SAM|18|9|押沙龍 剛好遇見了 大衛 的臣僕。 押沙龍 騎著騾子，從大橡樹密枝底下經過，他的頭被橡樹夾住，懸掛在空中 ，所騎的騾子就離他去了。
2SAM|18|10|有個人看見，就告訴 約押 說：「看哪，我看見 押沙龍 掛在橡樹上了。」
2SAM|18|11|約押 對報信的人說：「看哪，你既看見了，為甚麼不當場把他擊殺在地呢？我必賞你十個銀子和一條帶子。」
2SAM|18|12|那人對 約押 說：「即使我手裏得了一千銀子，也不敢伸手害王的兒子，因為我們聽見王囑咐你、 亞比篩 、 以太 說：『你們要謹慎，不可害那年輕人 押沙龍 。』
2SAM|18|13|我若冒著生命危險做這傻事 ，無論何事都瞞不過王，你自己也必遠遠站在一旁。」
2SAM|18|14|約押 說：「我不能在你面前這樣耗下去！」 約押 手拿三枝短槍，趁 押沙龍 在橡樹上 還活著，就刺透他的心。
2SAM|18|15|給 約押 拿兵器的十個青年圍著 押沙龍 ，擊殺他，將他殺死。
2SAM|18|16|約押 吹角，軍兵就回來，不去追趕 以色列 人，因為 約押 制止了軍兵。
2SAM|18|17|他們拿下 押沙龍 ，把他丟在樹林中一個大坑裏，上頭堆起一大堆石頭。 以色列 眾人都逃跑，各回自己的帳棚去了。
2SAM|18|18|押沙龍 活著的時候，曾在 王谷 立了一根柱子，因他說：「我沒有兒子為我留名。」他就以自己的名字稱那柱子為 押沙龍碑 ，直到今日。
2SAM|18|19|撒督 的兒子 亞希瑪斯 說：「讓我跑去報信給王，耶和華已經為王伸冤，使他脫離仇敵的手了。」
2SAM|18|20|約押 對他說：「你今日不可作報信的人，改日再去報信；因為今日王的兒子死了，所以你不可去報信。」
2SAM|18|21|約押 對 古實 人說：「你去把你所看見的告訴王。」 古實 人向 約押 叩拜後，就跑去了。
2SAM|18|22|撒督 的兒子 亞希瑪斯 又對 約押 說：「無論怎樣，讓我隨著 古實 人跑去吧！」 約押 說：「我兒，你報這信息，既不得賞賜，何必要跑去呢？」
2SAM|18|23|他說：「無論怎樣，我要跑去。」 約押 對他說：「你跑去吧！」 亞希瑪斯 就從平原的路往前跑，越過了 古實 人。
2SAM|18|24|大衛 正坐在內外城門之間。守望的人上到城牆，在城門的頂上舉目觀看，看哪，有一個人獨自跑來。
2SAM|18|25|守望的人就大聲告訴王。王說：「他若獨自來，必是報口信的。」那人跑得越來越近了。
2SAM|18|26|守望的人又見一人跑來，就對守城門的人喊說：「看哪，又有一人獨自跑來。」王說：「這也是報信的。」
2SAM|18|27|守望的人說：「我看前面那人的跑法，好像 撒督 的兒子 亞希瑪斯 的跑法。」王說：「他是個好人，是來報好消息的。」
2SAM|18|28|亞希瑪斯 向王呼叫說：「平安了！」他就臉伏於地向王叩拜，說：「耶和華－你的上帝是應當稱頌的，他已把些那舉手攻擊我主我王的人交出來了。」
2SAM|18|29|王說：「年輕人 押沙龍 平安嗎？」 亞希瑪斯 說：「 約押 派王的僕人，就是你的僕人時，我看見一陣大騷動，卻不知道是甚麼事。」
2SAM|18|30|王說：「你退去，站在這裏。」他就退去，站著。
2SAM|18|31|看哪， 古實 人也來到，說：「有信息報給我主我王！耶和華今日為你伸冤，使你脫離一切起來攻擊你之人的手。」
2SAM|18|32|王對 古實 人說：「年輕人 押沙龍 平安嗎？」 古實 人說：「願我主我王的仇敵，和一切起來惡意要害你的人，都像那年輕人一樣。」
2SAM|18|33|王戰抖，就上城門的樓房去痛哭，一面走一面說：「我兒 押沙龍 啊！我兒，我兒 押沙龍 啊！我恨不得替你死， 押沙龍 啊，我兒！我兒！」
2SAM|19|1|有人告訴 約押 ：「看哪，王為 押沙龍 悲哀哭泣。」
2SAM|19|2|那日眾軍兵聽說王為他兒子悲傷，他們得勝的日子變成悲哀了。
2SAM|19|3|那日軍兵暗暗地進城，如同戰場上逃跑、羞愧的士兵一般。
2SAM|19|4|王蒙著臉，大聲哭號說：「我兒 押沙龍 啊！ 押沙龍 ，我兒，我兒啊！」
2SAM|19|5|約押 進了宮到王那裏，說：「你今日使你眾臣僕的臉面羞愧了！他們今日救了你的性命和你兒女妻妾的性命，
2SAM|19|6|你卻愛那些恨你的人，恨那些愛你的人。今日你擺明了不以將帥、臣僕為念。我今日看得出，若 押沙龍 活著，我們今日全都死了，你就高興了。
2SAM|19|7|現在你要起來，出去安慰你臣僕的心。我指著耶和華起誓：你若不出去，今夜必沒有一人跟你在一起了。這禍患比你從幼年到如今所遭受的更嚴重！」
2SAM|19|8|於是王起來，坐在城門口。有人告訴眾軍兵說：「看哪，王坐在城門口。」眾軍兵就都到王的面前。 那時， 以色列 人已經逃跑，各回自己的帳棚去了。
2SAM|19|9|以色列 眾支派的百姓都議論紛紛，說：「王曾救我們脫離仇敵的手，又救我們脫離 非利士 人的手，現在他為了 押沙龍 逃離這地了。
2SAM|19|10|我們所膏治理我們的 押沙龍 已經陣亡。現在你們為甚麼沉默，不請王回來呢？」
2SAM|19|11|大衛 王派人到 撒督 和 亞比亞他 二位祭司那裏，說：「你們當向 猶大 長老說：『 以色列 眾人已經有話到了王那裏 ，你們為甚麼最後才請王回宮呢？
2SAM|19|12|你們是我的弟兄，是我的骨肉，為甚麼最後才請王回來呢？』
2SAM|19|13|你們要對 亞瑪撒 說：『你不是我的骨肉嗎？我若不立你在我面前取代 約押 永久作元帥，願上帝重重懲罰我！』」
2SAM|19|14|這樣，他挽回了 猶大 眾人的心，如同一人。他們就派人到王那裏，說：「請王和王的眾臣僕回來。」
2SAM|19|15|王回來了，到 約旦河 。 猶大 人來到 吉甲 ，去迎接王，請王過 約旦河 。
2SAM|19|16|來自 巴戶琳 的 便雅憫 人 基拉 的兒子 示每 急忙與 猶大 人一同下去迎接 大衛 王。
2SAM|19|17|跟從 示每 的有一千個 便雅憫 人，還有 掃羅 家的僕人 洗巴 和他十五個兒子、二十個隨從僕人，他們都趕緊過 約旦河 到王的面前。
2SAM|19|18|渡船就渡王的家眷過河 ，照王看為好的去做。 王過 約旦河 的時候， 基拉 的兒子 示每 俯伏在王面前，
2SAM|19|19|對王說：「我主我王離開 耶路撒冷 的那日，僕人行了悖逆的事，現在求我主不要因此加罪於僕人，不要記得，也不要放在心上。
2SAM|19|20|僕人明知自己有罪，看哪， 約瑟 全家之中，今日我首先下來迎接我主我王。」
2SAM|19|21|洗魯雅 的兒子 亞比篩 回答說：「 示每 既然咒罵耶和華的受膏者，不應當為這緣故處死他嗎？」
2SAM|19|22|大衛 說：「 洗魯雅 的兒子，我與你們有何相干，你們今日要跟我作對嗎？今日在 以色列 中豈可把任何人處死呢？我豈不知今日我是 以色列 的王嗎？」
2SAM|19|23|於是王對 示每 說：「你必不死。」王就向他起誓。
2SAM|19|24|掃羅 的孫子 米非波設 也下去迎接王。他自從王離開的那一日，直到王平安回 耶路撒冷 的日子，沒有修腳，沒有剃鬍鬚，也沒有洗衣服。
2SAM|19|25|他來迎接王的時候 ，王對他說：「 米非波設 ，你為甚麼沒有與我同去呢？」
2SAM|19|26|他說：「我主我王啊，我的僕人欺騙了我。那日僕人想要備驢騎上，與王同去，因為僕人是瘸腿的。
2SAM|19|27|他卻在我主我王面前毀謗僕人。然而我主我王如同上帝的使者一樣，你看怎樣好，就怎樣做吧！
2SAM|19|28|因為我祖全家的人，在我主我王面前不過是該死的人，王卻使僕人列在王的席上吃飯的人當中，我現在還有甚麼權利能向王請求呢？」
2SAM|19|29|王對他說：「你何必再提你的事呢？我說，你與 洗巴 要平分土地。」
2SAM|19|30|米非波設 對王說：「我主我王既然平安地回宮，甚至讓 洗巴 全都拿去也沒關係。」
2SAM|19|31|基列 人 巴西萊 從 羅基琳 下來，要護送王過 約旦河 ，就跟王一同過 約旦河 。
2SAM|19|32|巴西萊 年紀老邁，已經八十歲了。王住在 瑪哈念 的時候，他拿食物來供給王，因他是個大富翁。
2SAM|19|33|王對 巴西萊 說：「你與我一同渡過去，我要在 耶路撒冷 我的身邊奉養你。」
2SAM|19|34|巴西萊 對王說：「我還能活多少年日，可以與王一同上 耶路撒冷 呢？
2SAM|19|35|今日我已八十歲了，還能辨別美醜嗎？僕人還能嘗出飲食的滋味嗎？還能聽男女歌唱的聲音嗎？僕人何必拖累我主我王呢？
2SAM|19|36|僕人護送王過 約旦河 只是一件小事，王何必用這樣的賞賜來報答我呢？
2SAM|19|37|請讓我回去，死在我本城，葬在我父母的墓旁。看哪，這裏有 金罕 作王的僕人，讓他同我主我王過去，你看怎樣好，就怎樣對待他吧。」
2SAM|19|38|王說：「 金罕 可以與我一同過去，我必照你看為好的待他。你要我做的，我都會為你做。」
2SAM|19|39|於是眾百姓過了 約旦河 ，王也過去了。王親吻 巴西萊 ，為他祝福， 巴西萊 就回自己的地方去了。
2SAM|19|40|王渡過去 ，到了 吉甲 ， 金罕 也跟他過去。 猶大 眾百姓和 以色列 百姓的一半也都送王過去。
2SAM|19|41|看哪， 以色列 眾人來到王那裏，對王說：「我們的弟兄 猶大 人為甚麼暗暗地送王和王的家眷，以及所有跟隨王的人，過 約旦河 呢？」
2SAM|19|42|猶大 眾人回答 以色列 人說：「因為王與我們是親屬，你們為何因這事發怒呢？我們靠王吃了甚麼呢？王真正給了我們甚麼賞賜呢？」
2SAM|19|43|以色列 人回答 猶大 人說：「我們與王有十倍的關係，就是在 大衛 身上，我們也比你們更有權利 。你們為何藐視我們呢？我們不是最先提議請王回來的嗎？」但 猶大 人的話比 以色列 人的話更強硬。
2SAM|20|1|在那裏恰巧有一個無賴，名叫 示巴 ，是 便雅憫 人 比基利 的兒子。他吹角，說： 「我們與 大衛 無份， 與 耶西 的兒子無關。 以色列 啊，各回自己的帳棚去吧！」
2SAM|20|2|於是 以色列 眾人都離棄 大衛 去跟隨 比基利 的兒子 示巴 ，但 猶大 人從 約旦河 直到 耶路撒冷 ，都緊緊跟隨他們的王。
2SAM|20|3|大衛 王來到 耶路撒冷 ，進了宮，就把從前留下看守宮殿的十個妃嬪軟禁在冷宮，養活她們，卻不與她們親近。她們被關起來，活著如同寡婦，直到死的日子。
2SAM|20|4|王對 亞瑪撒 說：「你要在三日之內召集 猶大 人到我這裏來，你自己也要留在這裏。」
2SAM|20|5|亞瑪撒 就去召集 猶大 人，不過他卻耽延，過了王所定的期限。
2SAM|20|6|大衛 對 亞比篩 說：「現在 比基利 的兒子 示巴 對我們的危害恐怕比 押沙龍 更大。你要帶領你主的一些僕人追趕他，免得他得了堅固的城鎮，在我們眼前逃脫 。」
2SAM|20|7|約押 的人和 基利提 人、 比利提 人，以及所有的勇士都跟著 亞比篩 ，從 耶路撒冷 出去追趕 比基利 的兒子 示巴 。
2SAM|20|8|他們到了 基遍 的大石頭那裏， 亞瑪撒 來迎接他們。那時 約押 穿著戰衣，腰束佩刀的帶子，刀在鞘內。 約押 前行時，刀從鞘內掉出來。
2SAM|20|9|約押 對 亞瑪撒 說：「我的弟兄，你平安嗎？」他就用右手抓住 亞瑪撒 的鬍子，要親吻他。
2SAM|20|10|亞瑪撒 沒有防備 約押 手裏拿著的刀； 約押 用刀刺入他的肚腹，他的腸子流在地上， 約押 沒有再刺，他就死了。 約押 和他弟弟 亞比篩 往前追趕 比基利 的兒子 示巴 。
2SAM|20|11|有 約押 的一個僕人站在 亞瑪撒 屍體的旁邊，說：「誰喜愛 約押 ，誰歸順 大衛 ，就當跟隨 約押 。」
2SAM|20|12|亞瑪撒 渾身是血，躺在路中間。那人見眾百姓都站住，就把 亞瑪撒 的屍體從路上移到田間，把衣服蓋在他身上，因為他看見眾人經過時都站住。
2SAM|20|13|屍體從路上移走之後，眾人就都跟隨 約押 去追趕 比基利 的兒子 示巴 。
2SAM|20|14|示巴 走遍 以色列 各支派，直到 伯‧瑪迦 的 亞比拉 ；所有精選的人 都聚集跟隨他。
2SAM|20|15|跟隨 約押 的眾百姓到了 伯‧瑪迦 的 亞比拉 ，圍困 示巴 ，對著城建土堆，與城郭相對。他們猛撞城牆，要使城倒塌。
2SAM|20|16|一個有智慧的婦人從城上呼叫：「聽啊，聽啊，請你們告訴 約押 ：『近前來到這裏，我好與你說話。』」
2SAM|20|17|約押 就近前到她那裏，婦人對他說：「你是 約押 嗎？」他說：「我是。」婦人對他說：「請你聽使女的話。」 約押 說：「我正在聽。」
2SAM|20|18|婦人說：「古時有話說，當在 亞比拉 求問，事情就可以解決。
2SAM|20|19|我在 以色列 中是和平、忠誠的。你現在想要毀壞這城， 以色列 的根源 ，為何你要吞滅耶和華的產業呢？」
2SAM|20|20|約押 回答說：「不，我絕不吞滅和毀壞！
2SAM|20|21|話不是這麼說的，只是因為有一個 以法蓮 山區的人，就是 比基利 的兒子名叫 示巴 ，他舉手攻擊 大衛 王；你們只要把他一人交出來，我就離城而去。」婦人對 約押 說：「看哪，他的首級必從城牆上丟給你。」
2SAM|20|22|婦人憑她的智慧去勸眾百姓，他們就割下 比基利 的兒子 示巴 的首級，丟給 約押 。 約押 吹角，眾人就離城散開，各回自己的帳棚去了。 約押 回 耶路撒冷 ，到王那裏。
2SAM|20|23|約押 統管 以色列 全軍； 耶何耶大 的兒子 比拿雅 統管 基利提 人和 比利提 人；
2SAM|20|24|亞多蘭 管理勞役的人； 亞希律 的兒子 約沙法 作史官；
2SAM|20|25|示法 作書記； 撒督 和 亞比亞他 作祭司；
2SAM|20|26|睚珥 人 以拉 也作 大衛 的祭司。
2SAM|21|1|大衛 在位年間有饑荒，一連三年， 大衛 求問耶和華，耶和華說：「 掃羅 和他家犯了流人血之罪，因為他殺死了 基遍 人。」
2SAM|21|2|大衛 王召了 基遍 人來，跟他們說話。 基遍 人不是 以色列 人，而是 亞摩利 人中所剩下的人。 以色列 人曾向他們起誓， 掃羅 卻為 以色列 人和 猶大 人大發熱心，追殺他們，為了要消滅他們。
2SAM|21|3|大衛 對 基遍 人說：「我當為你們做甚麼呢？要用甚麼贖這罪，使你們為耶和華的產業祝福呢？」
2SAM|21|4|基遍 人對他說：「我們和 掃羅 以及他家的事與金銀無關，也不要因我們的緣故殺任何 以色列 人。」 大衛 說：「你們怎樣說，我就為你們怎樣做。」
2SAM|21|5|他們對王說：「那謀害我們、要消滅我們、使我們不得住 以色列 境內的人，
2SAM|21|6|請把他的子孫七人交給我們，我們好在耶和華面前，把他們懸掛在 基比亞 ，就是耶和華揀選 掃羅 的地方。」王說：「我必交給你們。」
2SAM|21|7|王顧惜 掃羅 的孫子， 約拿單 的兒子 米非波設 ，因為在 大衛 和 掃羅 的兒子 約拿單 之間，有指著耶和華的誓言。
2SAM|21|8|王卻把 愛亞 的女兒 利斯巴 為 掃羅 所生的兩個兒子 亞摩尼 和 米非波設 ，以及 掃羅 的女兒 米拉 為 米何拉 人 巴西萊 兒子 亞得列 所生的五個兒子
2SAM|21|9|交在 基遍 人的手裏。 基遍 人在耶和華面前把他們懸掛在山上，這七人就一起死了。他們被殺的時候正是收割的頭幾天，就是開始收割大麥的時候。
2SAM|21|10|愛亞 的女兒 利斯巴 用麻布舖在磐石上搭棚，從收割的開始直到天降雨在屍體上，她白日不許空中的飛鳥落在屍體上，夜間不讓田野的走獸前來。
2SAM|21|11|有人把 掃羅 的妃子 愛亞 女兒 利斯巴 所做的事告訴 大衛 。
2SAM|21|12|大衛 就去，從 基列 的 雅比 人那裏把 掃羅 和他兒子 約拿單 的骸骨搬來。先前 非利士 人在 基利波 殺了 掃羅 ，把屍體懸掛在 伯‧珊 的廣場上，後來 基列 的 雅比 人把屍體偷走。
2SAM|21|13|大衛 把 掃羅 和他兒子 約拿單 的骸骨從那裏搬上來，又收殮了被懸掛的那些人的骸骨。
2SAM|21|14|他們將 掃羅 和他兒子 約拿單 的骸骨葬在 便雅憫 的 洗拉 ，在 掃羅 父親 基士 的墳墓裏。他們遵照王所吩咐的一切做了。此後上帝垂聽了為那地的祈求。
2SAM|21|15|非利士 人與 以色列 人打仗。 大衛 帶領僕人下去，與 非利士 人交戰， 大衛 就疲乏了。
2SAM|21|16|巨人族的後裔 以實‧比諾 說要殺 大衛 ；他的銅槍重三百舍客勒，腰間又佩著新刀 。
2SAM|21|17|但 洗魯雅 的兒子 亞比篩 幫助 大衛 攻擊 非利士 人，殺死了他。當日， 大衛 的人向 大衛 起誓說：「你不可再與我們一同出戰，免得 以色列 的燈熄滅了。」
2SAM|21|18|後來，在 歌伯 又與 非利士 人打仗，那時 戶沙 人 西比該 殺了巨人族的後裔 撒弗 。
2SAM|21|19|他們又在 歌伯 與 非利士 人打仗， 伯利恆 人 雅雷 的兒子 伊勒哈難 殺了 迦特 人 歌利亞 ；這人的槍桿粗如織布機的軸。
2SAM|21|20|又有一次，他們在 迦特 打仗。那裏有一個身材高大的人，雙手各有六根手指，雙腳各有六根腳趾，共有二十四根；他也是巨人族的後裔。
2SAM|21|21|他向 以色列 罵陣， 大衛 的哥哥 示米亞 的兒子 約拿單 就殺了他。
2SAM|21|22|這四個人是 迦特 巨人族的後裔，都仆倒在 大衛 和他僕人的手下。
2SAM|22|1|當耶和華救 大衛 脫離所有仇敵和 掃羅 之手的日子，他用這詩的歌詞向耶和華說話。
2SAM|22|2|他說： 耶和華是我的巖石、我的山寨、我的救主、
2SAM|22|3|我的上帝、我的磐石、我所投靠的。 他是我的盾牌，是拯救我的角， 是我的碉堡，是我的避難所， 是我的救主，救我脫離兇暴的。
2SAM|22|4|我要求告當讚美的耶和華， 我必從仇敵手中被救出來。
2SAM|22|5|死亡的波浪環繞我， 毀滅的急流驚嚇我，
2SAM|22|6|陰間的繩索纏繞我， 死亡的圈套臨到我。
2SAM|22|7|我在急難中求告耶和華， 向我的上帝呼求。 他從殿中聽了我的聲音； 我的呼求進入他的耳中。
2SAM|22|8|那時，因他發怒地就搖撼震動； 天的根基也戰抖搖撼。
2SAM|22|9|他的鼻孔冒煙上騰； 他的口發火焚燒，連煤炭也燒著了。
2SAM|22|10|他使天下垂，親自降臨； 黑雲在他腳下。
2SAM|22|11|他乘坐基路伯飛行， 在風的翅膀上顯現。
2SAM|22|12|他以黑暗和聚集的水、 天空的密雲為四圍的行宮。
2SAM|22|13|因他發出光輝， 火炭都燒著了。
2SAM|22|14|耶和華在天上打雷； 至高者發出聲音。
2SAM|22|15|他射出箭來，使仇敵四散； 發出閃電，擊潰他們。
2SAM|22|16|耶和華的斥責一發，鼻孔的氣一出， 海底就顯現，大地的根基也暴露。
2SAM|22|17|他從高天伸手抓住我， 把我從大水中拉上來。
2SAM|22|18|他救我脫離我的強敵， 脫離那些恨我的人， 因為他們比我強盛。
2SAM|22|19|我遭遇災難的日子，他們來攻擊我； 但耶和華是我的倚靠。
2SAM|22|20|他領我到寬闊之處， 他救拔我，因他喜愛我。
2SAM|22|21|耶和華必按我的公義報答我， 按我手中的清潔賞賜我。
2SAM|22|22|因為我遵守耶和華的道， 未曾作惡離開我的上帝。
2SAM|22|23|他的一切典章在我面前， 他的律例我也未曾丟棄。
2SAM|22|24|我在他面前作了完全人， 我也持守自己遠離罪孽。
2SAM|22|25|所以耶和華按我的公義， 在他眼前按我的清潔賞賜我。
2SAM|22|26|慈愛的人，你以慈愛待他； 完全的人，你以完善待他；
2SAM|22|27|清潔的人，你以清潔待他； 歪曲的人，你以彎曲待他。
2SAM|22|28|困苦的百姓，你必拯救； 但你的眼目察看高傲的人，使他們降卑。
2SAM|22|29|耶和華啊，你是我的燈； 耶和華必照明我的黑暗。
2SAM|22|30|我藉著你衝入敵軍， 藉著我的上帝跳過城牆。
2SAM|22|31|至於上帝，他的道是完全的； 耶和華的話是純淨的。 凡投靠他的，他就作他們的盾牌。
2SAM|22|32|除了耶和華，誰是上帝呢？ 除了我們的上帝，誰是磐石呢？
2SAM|22|33|上帝是我堅固的保障， 他為我開完全的路。
2SAM|22|34|他使我的腳快如母鹿， 使我站穩在高處。
2SAM|22|35|他教導我的手能爭戰， 我的膀臂能開銅造的弓。
2SAM|22|36|你賜救恩給我作盾牌， 你的庇護 使我為大。
2SAM|22|37|你使我腳步寬闊， 我的腳踝未曾滑跌。
2SAM|22|38|我追趕我的仇敵，消滅他們； 若不將他們滅絕，我總不歸回。
2SAM|22|39|我滅絕了他們， 打傷了他們，使他們站不起來； 他們都倒在我的腳下。
2SAM|22|40|你曾以力量束我的腰，使我能爭戰； 也曾使那起來攻擊我的，都服在我以下。
2SAM|22|41|你又使我的仇敵在我面前轉身逃跑， 使我能殲滅那恨我的人。
2SAM|22|42|他們仰望，卻無人拯救； 就是呼求耶和華，他也不應允。
2SAM|22|43|我搗碎他們，如同地上的灰塵； 踐踏壓碎他們，如同街上的泥土。
2SAM|22|44|你救我脫離我百姓 的紛爭， 保護我作列國的元首； 我素不認識的百姓必事奉我。
2SAM|22|45|外邦人要向我投降， 一聽見我的名聲就必順從我。
2SAM|22|46|外邦人要喪膽， 戰戰兢兢地出營寨。
2SAM|22|47|耶和華永遠活著。 願我的磐石被稱頌， 願上帝－救我的磐石受尊崇。
2SAM|22|48|這位上帝為我伸冤， 使萬民服在我以下。
2SAM|22|49|他救我脫離仇敵， 又把我舉起，高過那些起來攻擊我的人， 救我脫離殘暴的人。
2SAM|22|50|耶和華啊，因此我要在列國中稱謝你， 歌頌你的名。
2SAM|22|51|耶和華賜極大的救恩給他所立的王， 施慈愛給他的受膏者， 就是給 大衛 和他的後裔，直到永遠！
2SAM|23|1|以下是 大衛 末了的話： 「 耶西 的兒子 大衛 的話， 得居高位的， 雅各 的上帝所膏的， 以色列 所喜愛的詩人的話。
2SAM|23|2|耶和華的靈藉著我說話， 他的言語在我的舌頭上。
2SAM|23|3|以色列 的上帝說， 以色列 的磐石向我說： 『那以公義治理人， 以敬畏上帝來治理的，
2SAM|23|4|他必像晨光， 如無雲清晨的日出， 如雨後的光輝， 在嫩草地上。』
2SAM|23|5|我的家在上帝面前不是如此嗎？ 上帝與我立永遠的約， 這約既全備又穩妥。 我的一切救恩和我一切所想望的， 他豈不成全嗎？
2SAM|23|6|但無賴全都像被丟棄的荊棘； 它們不能用手去拿；
2SAM|23|7|碰它們的人必須用鐵器和槍桿， 它們必在那裏被火燒盡。」
2SAM|23|8|大衛 勇士的名字如下： 哈革摩尼 人 約設‧巴設 ，他是三勇士之首；他又名叫 伊斯尼 人 亞底挪 ，曾一次就殺了八百人 。
2SAM|23|9|跟隨 大衛 的三勇士中，其次是 亞何亞 人 朵多 的兒子 以利亞撒 。從前 非利士 人聚集要打仗，他們向 非利士 人罵陣。 以色列 人上去的時候，
2SAM|23|10|他起來擊殺 非利士 人，直到手臂疲乏，手黏住刀把。那日耶和華大獲全勝，百姓跟在 以利亞撒 後面只顧奪取掠物。
2SAM|23|11|再其次是 哈拉 人 亞基 的兒子 沙瑪 。一次， 非利士 人聚集在 利希 ，在一塊長滿紅豆的田裏，百姓在 非利士 人面前逃跑。
2SAM|23|12|沙瑪 卻站在那田的中間，防守那田，擊敗了 非利士 人。耶和華大獲全勝。
2SAM|23|13|開始收割的時候，三個 侍衛 下到 亞杜蘭洞 ，到 大衛 那裏。 非利士 的軍兵在 利乏音谷 安營。
2SAM|23|14|那時 大衛 在山寨， 非利士 人的駐軍在 伯利恆 。
2SAM|23|15|大衛 渴想著說：「但願有人從 伯利恆 城門旁的井裏打水來給我喝！」
2SAM|23|16|這三個勇士就闖過 非利士 人的軍營，從 伯利恆 城門旁的井裏打水，拿來給 大衛 喝。他卻不肯喝，將水澆在耶和華面前，
2SAM|23|17|說：「耶和華啊，我絕不做這事！這三個人冒生命的危險，這不是他們的血嗎？」 大衛 不肯喝這水。這是三個勇士所做的事。
2SAM|23|18|洗魯雅 的兒子， 約押 的兄弟 亞比篩 是這三個勇士的領袖；他曾舉槍殺了三百人，就在三個勇士中得了名。
2SAM|23|19|他在這三個 勇士中是最有名望的，所以作他們的領袖，只是不及前三個勇士。
2SAM|23|20|耶何耶大 的兒子 比拿雅 是來自 甲薛 的勇士，曾行了大事。他殺了 摩押 人 亞利伊勒 的兩個兒子，又在下雪的時候下到坑裏去，殺了一隻獅子。
2SAM|23|21|他又殺了一個魁梧的 埃及 人； 埃及 人手裏拿著槍。 比拿雅 只拿著棍子下到他那裏去，從 埃及 人手裏奪過槍來，用那槍殺死了他。
2SAM|23|22|這些是 耶何耶大 的兒子 比拿雅 所做的事，就在三個勇士裏得了名。
2SAM|23|23|他比那三十個勇士 更有名望，只是不及前三個勇士。 大衛 立他作護衛長。
2SAM|23|24|三十個勇士中有 約押 的兄弟 亞撒黑 ， 伯利恆 人 朵多 的兒子 伊勒哈難 ，
2SAM|23|25|哈律 人 沙瑪 ， 哈律 人 以利加 ，
2SAM|23|26|帕勒提 人 希利斯 ， 提哥亞 人 益吉 的兒子 以拉 ，
2SAM|23|27|亞拿突 人 亞比以謝 ， 戶沙 人 米本乃 ，
2SAM|23|28|亞何亞 人 撒們 ， 尼陀法 人 瑪哈萊 ，
2SAM|23|29|尼陀法 人 巴拿 的兒子 希立 ， 便雅憫 族 基比亞 人 利拜 的兒子 以太 ，
2SAM|23|30|比拉頓 人 比拿雅 ， 迦實溪 人 希太 ，
2SAM|23|31|亞拉巴 人 亞比‧亞本 ， 巴魯米 人 押斯瑪弗 ，
2SAM|23|32|沙本 人 以利雅哈巴 ， 雅善 兒子中的 約拿單 ，
2SAM|23|33|哈拉 人 沙瑪 ， 哈拉 人 沙拉 的兒子 亞希暗 ，
2SAM|23|34|瑪迦 人 亞哈拜 的兒子 以利法列 ， 基羅 人 亞希多弗 的兒子 以連 ，
2SAM|23|35|迦密 人 希斯萊 ， 亞巴 人 帕萊 ，
2SAM|23|36|瑣巴 人 拿單 的兒子 以甲 ， 迦得 人 巴尼 ，
2SAM|23|37|亞捫 人 洗勒 ， 比錄 人 拿哈萊 ，是給 洗魯雅 的兒子 約押 拿兵器的，
2SAM|23|38|以帖 人 以拉 ， 以帖 人 迦立 ，
2SAM|23|39|赫 人 烏利亞 ，共三十七人。
2SAM|24|1|耶和華的怒氣又向 以色列 發作，激起 大衛 來對付他們，說：「去，數點 以色列 人和 猶大 人。」
2SAM|24|2|大衛 對跟隨他的 約押 元帥說：「你來回走遍 以色列 眾支派，從 但 直到 別是巴 ，數點百姓，我好知道百姓的數目。」
2SAM|24|3|約押 對王說：「願耶和華－你的上帝使百姓的數目增加百倍，使我主我王親眼得見。我主我王何必要做這事呢？」
2SAM|24|4|但王堅持他對 約押 和眾軍官的命令。 約押 和眾軍官就從王面前出去，數點 以色列 的百姓。
2SAM|24|5|他們過 約旦河 ，在 迦得谷 中、城的右邊 亞羅珥 安營，與 雅謝 相對。
2SAM|24|6|他們來到 基列 ，到了 他停‧合示 地 ，又來到 但‧雅安 ，繞到 西頓 。
2SAM|24|7|他們來到 推羅 的堡壘，以及 希未 人和 迦南 人的各城，又出來，到 猶大尼革夫 的 別是巴 。
2SAM|24|8|他們來回走遍全地，過了九個月又二十天，就回到 耶路撒冷 。
2SAM|24|9|約押 向王報告百姓的總數： 以色列 拿刀的勇士有八十萬； 猶大 有五十萬人。
2SAM|24|10|大衛 數點百姓以後，心中自責。大衛向耶和華說：「我做這事大大有罪了。耶和華啊，現在求你除掉僕人的罪孽，因我所做的非常愚昧。」
2SAM|24|11|大衛 早晨起來，耶和華的話臨到 迦得 先知，就是 大衛 的先見，說：
2SAM|24|12|「你去告訴 大衛 ：『耶和華如此說：我向你提出三樣，隨你選擇一樣，我好降給你。』」
2SAM|24|13|於是 迦得 來到 大衛 那裏告訴他，問他：「你要國中有七 年的饑荒呢？或是你在敵人面前逃跑，被追趕三個月呢？或是在你國中有三日的瘟疫呢？現在你要考慮思量，我怎樣去回覆那差我來的。」
2SAM|24|14|大衛 對 迦得 說：「我很為難。我們寧願落在耶和華的手裏，因為他有豐盛的憐憫；我不願落在人的手裏。」
2SAM|24|15|於是，耶和華降瘟疫給 以色列 。自早晨到所定的時候，從 但 直到 別是巴 ，百姓中死了七萬人。
2SAM|24|16|天使向 耶路撒冷 伸手要毀滅這城的時候，耶和華改變心意，不降那災難，就對那在百姓中施行毀滅的天使說：「夠了！住手吧！」耶和華的使者正在 耶布斯 人 亞勞拿 的禾場那裏。
2SAM|24|17|大衛 看見那在百姓中施行毀滅的天使，就向耶和華說：「看哪，我犯了罪，行了惡，但這群羊做了甚麼呢？願你的手攻擊我和我的父家。」
2SAM|24|18|當日， 迦得 來到 大衛 那裏，對他說：「你上去，在 耶布斯 人 亞勞拿 的禾場上為耶和華立一座壇。」
2SAM|24|19|大衛 就照著 迦得 的話，照著耶和華所吩咐的上去了。
2SAM|24|20|亞勞拿 觀看，看見王和臣僕向他走過來。 亞勞拿 就出去，臉伏於地，向王下拜。
2SAM|24|21|亞勞拿 說：「我主我王為何來到僕人這裏呢？」 大衛 說：「我要買你這禾場，為耶和華築一座壇，使瘟疫在百姓中停止。」
2SAM|24|22|亞勞拿 對 大衛 說：「我主我王，你眼中看為好，就拿去獻祭。看，這裏有牛可以作燔祭，有打糧的器具和套牛的軛可以當作柴。
2SAM|24|23|王啊，這一切， 亞勞拿 都獻給王。」 亞勞拿 又對王說：「願耶和華－你的上帝悅納你。」
2SAM|24|24|王對 亞勞拿 說：「不，我一定要按價錢向你買；我不能用白白得來的東西作燔祭獻給耶和華－我的上帝。」 大衛 就用五十舍客勒銀子買了那禾場與牛。
2SAM|24|25|大衛 在那裏為耶和華築了一座壇，獻燔祭和平安祭。耶和華垂聽了為那地的祈求，瘟疫就在 以色列 中停止了。
1KGS|1|1|大衛 王年紀老邁，雖然蓋著外袍，仍不夠暖和。
1KGS|1|2|臣僕對他說：「不如為我主我王找一個年輕的少女，侍立在王面前，照顧王，睡在王的懷中，好使我主我王得暖。」
1KGS|1|3|於是他們在 以色列 全境尋找美貌的少女，找到了一個 書念 女子 亞比煞 ，帶到王那裏。
1KGS|1|4|這少女極其美貌，她照顧王，伺候王，王卻沒有與她親近。
1KGS|1|5|那時， 哈及 的兒子 亞多尼雅 妄自尊大，說：「我要作王」，就為自己預備座車、騎兵，又派五十人在他前頭奔跑。
1KGS|1|6|他父親從來沒有責怪他，說：「你為何這麼做？」他非常俊美，生在 押沙龍 之後。
1KGS|1|7|亞多尼雅 與 洗魯雅 的兒子 約押 和 亞比亞他 祭司商議；他們就順從 亞多尼雅 ，幫助他。
1KGS|1|8|但 撒督 祭司、 耶何耶大 的兒子 比拿雅 、 拿單 先知、 示每 、 利以 ，以及 大衛 自己的勇士 都不順從 亞多尼雅 。
1KGS|1|9|亞多尼雅 在 隱‧羅結 旁 瑣希列 磐石那裏獻牛羊、肥犢為祭，請了他的眾兄弟，就是王的眾兒子，以及所有作王臣僕的 猶大 人。
1KGS|1|10|但他沒有邀請 拿單 先知、 比拿雅 和勇士們，以及他的弟弟 所羅門 。
1KGS|1|11|拿單 對 所羅門 的母親 拔示巴 說：「 哈及 的兒子 亞多尼雅 作王了，你沒有聽見嗎？我們的主 大衛 卻不知道。
1KGS|1|12|現在，來，我給你出個主意，好保全你和你兒子 所羅門 的性命。
1KGS|1|13|你去，進到 大衛 王那裏，對他說：『我主我王啊，你不是曾向使女起誓說：你兒子 所羅門 必接續我作王，他必坐在我的王位上嗎？ 亞多尼雅 怎麼作了王呢？』
1KGS|1|14|看哪，你還在那裏與王說話的時候，我會隨後進去，證實你的話。」
1KGS|1|15|拔示巴 進入內室，到王那裏。那時，王很老了， 書念 女子 亞比煞 正伺候著王。
1KGS|1|16|拔示巴 向王屈身下拜，王說：「你要甚麼？」
1KGS|1|17|她對王說：「我主啊，你曾向使女指著耶和華－你的上帝起誓：『你兒子 所羅門 必接續我作王，他必坐在我的王位上。』
1KGS|1|18|現在，看哪， 亞多尼雅 作王了，你 ，我主我王卻不知道。
1KGS|1|19|他獻許多牛羊、肥犢為祭，請了王的眾兒子和 亞比亞他 祭司，以及 約押 元帥，他卻沒有請王的僕人 所羅門 。
1KGS|1|20|但你 ，我主我王啊， 以色列 眾人的眼目都仰望你，等你告訴他們，在我主我王之後誰坐你的王位。
1KGS|1|21|若不然，我主我王與祖先同睡的時候，我和我兒子 所羅門 必列為罪犯了。」
1KGS|1|22|看哪， 拔示巴 還與王說話的時候， 拿單 先知也進來了。
1KGS|1|23|有人奏告王說：「看哪， 拿單 先知來了。」 拿單 進到王面前，臉伏於地，向王叩拜。
1KGS|1|24|拿單 說：「我主我王，你果真說過『 亞多尼雅 必接續我作王，他要坐在我的王位上』嗎？
1KGS|1|25|他今日下去，獻了許多牛羊、肥犢為祭，請了王的眾兒子和軍官們，以及 亞比亞他 祭司；看哪，他們正在 亞多尼雅 面前吃喝，說：『 亞多尼雅 王萬歲！』
1KGS|1|26|至於我，就是你的僕人，和 撒督 祭司、 耶何耶大 的兒子 比拿雅 、王的僕人 所羅門 ，他都沒有請。
1KGS|1|27|這事果真出於我主我王嗎？王卻沒有告訴僕人們，在我主我王之後誰坐你的王位。」
1KGS|1|28|大衛 王回答說：「召 拔示巴 到我這裏來。」 拔示巴 就來，站在王面前。
1KGS|1|29|王起誓說：「我指著救我性命脫離一切苦難的永生的耶和華起誓。
1KGS|1|30|我既然指著耶和華－ 以色列 的上帝向你起誓說：你兒子 所羅門 必接續我作王，他必繼承我坐在我的王位上，我今日必這樣做。」
1KGS|1|31|於是， 拔示巴 屈身，臉伏於地，向王叩拜，說：「我主 大衛 王萬歲！」
1KGS|1|32|大衛 王又說：「召 撒督 祭司、 拿單 先知、 耶何耶大 的兒子 比拿雅 到我這裏來！」他們就都來到王面前。
1KGS|1|33|王對他們說：「要帶領你們主的僕人，讓我兒子 所羅門 騎我自己的騾子，送他下到 基訓 。
1KGS|1|34|在那裏， 撒督 祭司和 拿單 先知要膏他作 以色列 的王；你們也要吹角，說：『 所羅門 王萬歲！』
1KGS|1|35|你們要跟隨他上來，使他坐在我的王位上，他要接續我作王。我已立他作 以色列 和 猶大 的君王。」
1KGS|1|36|耶何耶大 的兒子 比拿雅 回應王說：「阿們！願耶和華－我主我王的上帝這樣說。
1KGS|1|37|耶和華怎樣與我主我王同在，願他照樣與 所羅門 同在，使他的王位比我主 大衛 王的王位更大。」
1KGS|1|38|於是， 撒督 祭司、 拿單 先知、 耶何耶大 的兒子 比拿雅 ，以及 基利提 人和 比利提 人都下去，讓 所羅門 騎上 大衛 王的騾子，送他到 基訓 。
1KGS|1|39|撒督 祭司從帳幕中取了盛膏油的角來，膏 所羅門 。他們就吹角，眾百姓都說：「 所羅門 王萬歲！」
1KGS|1|40|眾百姓跟隨他上來，吹著笛，大大歡呼，地被他們的聲音震裂。
1KGS|1|41|亞多尼雅 和所有的賓客剛吃完，聽見這聲音； 約押 聽見角聲就說：「城中為何有這響聲呢？」
1KGS|1|42|他正說話的時候，看哪， 亞比亞他 祭司的兒子 約拿單 來了。 亞多尼雅 說：「進來吧！你是個賢明的人，必是來報好消息的。」
1KGS|1|43|約拿單 回答 亞多尼雅 說：「我們的主 大衛 王已經立 所羅門 為王了！
1KGS|1|44|王派 撒督 祭司、 拿單 先知、 耶何耶大 的兒子 比拿雅 ，以及 基利提 人和 比利提 人和 所羅門 一起去，叫他騎上王的騾子。
1KGS|1|45|撒督 祭司和 拿單 先知已經在 基訓 膏他作王了。他們從那裏歡呼著上來，城都震動，這就是你們所聽見的聲音。
1KGS|1|46|所羅門 也已經登上國度的王位了。
1KGS|1|47|王的臣僕也來為我們的主 大衛 王祝福，說：『願上帝使 所羅門 的名比你的名更尊榮，使他的王位比你的王位更大。』王在床上屈身敬拜，
1KGS|1|48|王也這樣說：『耶和華－ 以色列 的上帝是應當稱頌的，因他今日賞賜一個人坐在我的王位上，我也親眼看見了。』」
1KGS|1|49|亞多尼雅 所有的賓客都戰兢，起來，各走各路去了。
1KGS|1|50|亞多尼雅 懼怕 所羅門 ，就起來，去抓住祭壇的翹角。
1KGS|1|51|有人告訴 所羅門 說：「看哪， 亞多尼雅 懼怕 所羅門 王。看哪，他抓住祭壇的翹角，說：『願 所羅門 王先向我起誓，必不用刀殺死僕人。』」
1KGS|1|52|所羅門 說：「他若作賢明的人，連一根頭髮也不致落在地上；他若作惡，必要死亡。」
1KGS|1|53|於是 所羅門 王派人叫 亞多尼雅 從壇上下來，他就來向 所羅門 王下拜。 所羅門 對他說：「你回家去吧！」
1KGS|2|1|大衛 的死期臨近了，就吩咐他兒子 所羅門 說：
1KGS|2|2|「我要走世人必走的路了。你當剛強，作大丈夫，
1KGS|2|3|遵守耶和華－你上帝所吩咐的，照著 摩西 律法上所寫的行耶和華的道，謹守他的律例、誡命、典章、法度，好讓你無論做甚麼，不拘往何處去，盡都亨通。
1KGS|2|4|耶和華必成就他所說關於我的話，說：『你的子孫若謹慎自己的行為，盡心盡意憑信實行在我面前，就不斷有人坐 以色列 的王位。』
1KGS|2|5|你也知道 洗魯雅 的兒子 約押 向我所做的事，他對付 以色列 的兩個元帥， 尼珥 的兒子 押尼珥 和 益帖 的兒子 亞瑪撒 ，殺了他們。他在太平之時，如同戰爭一般，流這二人的血，把這戰爭的血染了他腰間束的帶和腳上穿的鞋。
1KGS|2|6|所以你要照你的智慧去做，不讓他白髮安然下陰間。
1KGS|2|7|你當恩待 基列 人 巴西萊 的眾兒子，請他們常與你同席吃飯，因為我躲避你哥哥 押沙龍 的時候，他們親近我。
1KGS|2|8|看哪，在你這裏有來自 巴戶琳 的 便雅憫 人， 基拉 的兒子 示每 。我到 瑪哈念 去的那日，他用狠毒的言語咒罵我。後來他卻下 約旦河 迎接我，我就指著耶和華向他起誓說：『我必不用刀殺死你。』
1KGS|2|9|但現在你不要以他為無罪。你是有智慧的人，必知道怎樣待他，使他白髮流血下陰間。」
1KGS|2|10|大衛 與他祖先同睡，葬在 大衛城 。
1KGS|2|11|大衛 作 以色列 王四十年：在 希伯崙 作王七年，在 耶路撒冷 作王三十三年。
1KGS|2|12|所羅門 坐他父親 大衛 的王位，他的國度非常穩固。
1KGS|2|13|哈及 的兒子 亞多尼雅 到 所羅門 的母親 拔示巴 那裏， 拔示巴 問他說：「你是為平安來的嗎？」他說：「為平安來的。」
1KGS|2|14|他又說：「我有話對你說。」 拔示巴 說：「你說吧。」
1KGS|2|15|亞多尼雅 說：「你知道這國原是歸我的，全 以色列 也都期望我作王。然而，這國反歸了我兄弟，因這國歸了他是出乎耶和華。
1KGS|2|16|現在我有一件事求你，請你不要推辭。」 拔示巴 對他說：「你說吧。」
1KGS|2|17|他說：「求你請 所羅門 王把 書念 女子 亞比煞 賜我為妻，因他必不拒絕你。」
1KGS|2|18|拔示巴 說：「好，我必為你對王提說。」
1KGS|2|19|於是， 拔示巴 來到 所羅門 王那裏，要為 亞多尼雅 說話。王起來迎接，向她下拜，然後坐在自己的位上，又為王的母親設一座位，她就坐在王的右邊。
1KGS|2|20|拔示巴 說：「我要向你提出一個小小的請求，請你不要回絕我。」王對她說：「母親，請提出來，我必不回絕你。」
1KGS|2|21|拔示巴 說：「請你把 書念 女子 亞比煞 賜給你哥哥 亞多尼雅 為妻。」
1KGS|2|22|所羅門 王回答母親說：「為何替 亞多尼雅 求 書念 女子 亞比煞 呢？可以為他求王國吧！他是我的兄長，不但為他，也為 亞比亞他 祭司和 洗魯雅 的兒子 約押 求吧！ 」
1KGS|2|23|所羅門 王指著耶和華起誓說：「 亞多尼雅 講這話是自己送命，不然，願上帝重重懲罰我。
1KGS|2|24|耶和華堅立我，使我坐在父親 大衛 的王位上，照著他所應許的為我建立家室；現在我指著永生的耶和華起誓， 亞多尼雅 今日必被處死。」
1KGS|2|25|於是 所羅門 王派 耶何耶大 的兒子 比拿雅 去擊殺 亞多尼雅 ，他就死了。
1KGS|2|26|王對 亞比亞他 祭司說：「你回 亞拿突 歸自己的田地去吧！你本是該死的，但因你在我父親 大衛 面前抬過主耶和華的約櫃，又與我父親同受一切苦難，所以我今日不殺死你。」
1KGS|2|27|所羅門 就革除 亞比亞他 ，不讓他作耶和華的祭司。這就應驗了耶和華在 示羅 論 以利 家所說的話。
1KGS|2|28|雖然 約押 沒有擁護 押沙龍 ，卻擁護了 亞多尼雅 ；這消息傳到 約押 那裏，他就逃到耶和華的帳幕，抓住祭壇的翹角。
1KGS|2|29|有人告訴 所羅門 王：「 約押 逃到耶和華的帳幕，看哪，他在祭壇的旁邊。」 所羅門 就派 耶何耶大 的兒子 比拿雅 ，說：「去，殺了他。」
1KGS|2|30|比拿雅 來到耶和華的帳幕，對 約押 說：「王這樣吩咐：『你出來吧！』」他說：「不，我要死在這裏。」 比拿雅 就去回覆王，說：「 約押 這樣說，他這樣回答我。」
1KGS|2|31|王對他說：「你可以照著他的話去做，殺了他，把他葬了，好叫 約押 流無辜人血的罪不歸在我和我的父家。
1KGS|2|32|耶和華必使 約押 的血歸到他自己頭上，因為他擊殺兩個比他又公義又良善的人，就是 尼珥 的兒子 以色列 的元帥 押尼珥 和 益帖 的兒子 猶大 的元帥 亞瑪撒 ，用刀殺了他們，我父親 大衛 卻不知道。
1KGS|2|33|這二人的血必歸到 約押 和他後裔頭上，直到永遠；惟有 大衛 和他的後裔，以及他的家與王位，必從耶和華那裏得平安，直到永遠。」
1KGS|2|34|於是 耶何耶大 的兒子 比拿雅 上去，擊殺 約押 ，殺死他，把他葬在曠野 約押 自己的家裏。
1KGS|2|35|王就立 耶何耶大 的兒子 比拿雅 作元帥，代替 約押 ，又使 撒督 祭司代替 亞比亞他 。
1KGS|2|36|王派人召 示每 來，對他說：「你要在 耶路撒冷 為自己建造房屋，住在那裏，不可從那裏出來到任何地方去。
1KGS|2|37|你當確實知道，你何日出來過 汲淪溪 ，就必定死！你的血必歸到自己頭上。」
1KGS|2|38|示每 對王說：「這話很好！我主我王怎樣說，僕人必照樣做。」於是 示每 住在 耶路撒冷 許多日子。
1KGS|2|39|過了三年， 示每 的兩個奴僕逃到 瑪迦 的兒子 迦特 王 亞吉 那裏去。有人告訴 示每 說：「看哪，你的奴僕在 迦特 。」
1KGS|2|40|示每 起來，備上驢，往 迦特 到 亞吉 那裏去找他的奴僕，從 迦特 帶他的奴僕回來。
1KGS|2|41|有人告訴 所羅門 ：「 示每 出 耶路撒冷 到 迦特 去，又回來了。」
1KGS|2|42|王就派人召 示每 來，對他說：「我豈不是叫你指著耶和華起誓，並且警告你說『你當確實知道，你何日出來到任何地方去，就必定死』嗎？你也對我說：『這話很好，我必聽從。』
1KGS|2|43|你為何不遵守你對耶和華的誓言和我吩咐你的命令呢？」
1KGS|2|44|王又對 示每 說：「你向我父親 大衛 所做的一切惡事，你自己心裏都知道，耶和華必使你的罪惡歸到你自己的頭上。
1KGS|2|45|但 所羅門 王必蒙福， 大衛 的王位必在耶和華面前堅立，直到永遠。」
1KGS|2|46|於是王吩咐 耶何耶大 的兒子 比拿雅 ，他就出去，擊殺 示每 ， 示每 就死了。這樣，國度在 所羅門 的手中鞏固了。
1KGS|3|1|所羅門 與 埃及 王法老結親，娶了法老的女兒，接她進入 大衛城 ，直等到建完了自己的宮和耶和華的殿，以及 耶路撒冷 周圍的城牆。
1KGS|3|2|當那些日子，百姓仍在丘壇獻祭，因為還沒有為耶和華的名建殿。
1KGS|3|3|所羅門 愛耶和華，遵行他父親 大衛 的律例，只是還在丘壇獻祭燒香。
1KGS|3|4|所羅門 王到 基遍 ，在那裏獻祭，因為 基遍 有極大的丘壇。 所羅門 在那壇上獻了一千祭牲為燔祭。
1KGS|3|5|在 基遍 ，耶和華夜間在夢中向 所羅門 顯現；上帝說：「你願我賜你甚麼，你可以求。」
1KGS|3|6|所羅門 說：「你曾向你僕人我父親 大衛 大施慈愛，因為他用忠信、公義、正直的心行在你面前。你又為他存留大慈愛，賜他一個兒子坐在他的王位上，正如今日一樣。
1KGS|3|7|現在，耶和華－我的上帝啊，你使僕人接續我父親 大衛 作王；但我是幼小的孩子，不知道應當怎樣出入。
1KGS|3|8|僕人住在你揀選的百姓中，這百姓之多，多得不可點，不可算。
1KGS|3|9|所以求你賜僕人善於了解的心，可以判斷你的百姓，辨別是非。不然，誰能判斷你這麼多的百姓呢？」
1KGS|3|10|所羅門 因為求這事，就蒙主喜悅。
1KGS|3|11|上帝對他說：「你既然求這事，不為自己求壽、求富，也不求滅絕你仇敵的性命，只求能明辨，可以聽訟，
1KGS|3|12|看哪，我會照你的話去做，看哪，我會賜你智慧和明辨的心，在你以前沒有像你的，在你以後也沒有興起像你的。
1KGS|3|13|你沒有求的，我也賜給你，就是富足、尊榮，使你在世一切的日子，列王中沒有一個能比你的。
1KGS|3|14|你若遵行我的道，謹守我的律例、誡命，正如你父親 大衛 所行的，我必使你長壽。」
1KGS|3|15|所羅門 醒了，看哪，是個夢。他就來到 耶路撒冷 ，站在耶和華的約櫃前，獻燔祭和平安祭，又為眾臣僕擺設宴席。
1KGS|3|16|那時，有兩個妓女來，站在王面前。
1KGS|3|17|一個婦人說：「我主啊，我和這婦人同住一屋。她在屋子裏的時候，我生了一個孩子。
1KGS|3|18|我生了以後第三天，這婦人也生了。我們是一起的，屋子裏除了我們二人之外，再沒有別人在屋子裏。
1KGS|3|19|夜間，這婦人的兒子死了，因為她壓在她的兒子身上。
1KGS|3|20|她半夜起來，趁你使女睡著的時候，從我旁邊把我兒子抱走，放在她懷裏，又把她死的兒子放在我懷裏。
1KGS|3|21|清早，我起來要給我的兒子吃奶，看哪，他死了；早晨我仔細察看他，看哪，他不是我所生的兒子。」
1KGS|3|22|另一個婦人說：「不！我的兒子是活的，你的兒子是死的。」但這一個說：「不！你的兒子是死的，我的兒子是活的。」她們就在王面前爭吵。
1KGS|3|23|王說：「這婦人說：『這是我的兒子，他是活的，你的兒子是死的。』那婦人說：『不！你的兒子是死的，我的兒子是活的。』」
1KGS|3|24|王就說：「給我拿刀來！」人就把刀拿到王面前來。
1KGS|3|25|王說：「把活孩子劈成兩半，一半給這婦人，一半給那婦人。」
1KGS|3|26|活孩子的母親為自己的兒子心急如焚，對王說：「求我主把活孩子給那婦人吧，萬不可殺死他！」那婦人說：「這孩子也不歸我，也不歸你，你們就劈了吧！」
1KGS|3|27|王回應說：「把活孩子給這婦人，萬不可殺死他，因為這婦人是他的母親。」
1KGS|3|28|全 以色列 聽見王這樣判斷，就都敬畏王，因為他們看見他心中有上帝的智慧，能夠斷案。
1KGS|4|1|所羅門 作全 以色列 的王。
1KGS|4|2|這些是他的官員： 撒督 的兒子 亞撒利雅 作祭司，
1KGS|4|3|示沙 的兩個兒子 以利何烈 、 亞希亞 作書記， 亞希律 的兒子 約沙法 作史官，
1KGS|4|4|耶何耶大 的兒子 比拿雅 作元帥， 撒督 和 亞比亞他 作祭司，
1KGS|4|5|拿單 的兒子 亞撒利雅 作宰相， 拿單 的兒子 撒布得 作祭司和王的顧問，
1KGS|4|6|亞希煞 作管家， 亞比大 的兒子 亞多尼蘭 掌管服勞役的工人。
1KGS|4|7|所羅門 在全 以色列 有十二個官員，供給王和王室的食物，每年各人供給一個月。
1KGS|4|8|這些是他們的名字：在 以法蓮 山區有 便‧戶珥 ；
1KGS|4|9|在 瑪迦斯 、 沙賓 、 伯‧示麥 、 以倫‧伯‧哈南 有 便‧底甲 ；
1KGS|4|10|在 亞魯泊 有 便‧希悉 ，他管理 梭哥 和 希弗 全地；
1KGS|4|11|在 多珥 山岡 有 便‧亞比拿達 ，他娶了 所羅門 的女兒 她法 為妻；
1KGS|4|12|在 他納 和 米吉多 ，以及靠近 撒拉他拿 、 耶斯列 下邊的 伯‧善 全地，從 伯‧善 到 亞伯‧米何拉 直到 約緬 的另一邊有 亞希律 的兒子 巴拿 ；
1KGS|4|13|在 基列 的 拉末 有 便‧基別 ，他管理在 基列 的 瑪拿西 子孫 睚珥 的城鎮， 巴珊 的 亞珥歌伯 地的六十座大城，各有城牆和銅閂；
1KGS|4|14|在 瑪哈念 有 易多 的兒子 亞希拿達 ；
1KGS|4|15|在 拿弗他利 有 亞希瑪斯 ，他也娶了 所羅門 的一個女兒 巴實抹 為妻；
1KGS|4|16|在 亞設 和 亞祿 有 戶篩 的兒子 巴拿 ；
1KGS|4|17|在 以薩迦 有 帕路亞 的兒子 約沙法 ；
1KGS|4|18|在 便雅憫 有 以拉 的兒子 示每 ；
1KGS|4|19|在 基列 地，就是 亞摩利 王 西宏 和 巴珊 王 噩 之地，有 烏利 的兒子 基別 ，他一個官員管理這地 。
1KGS|4|20|猶大 人和 以色列 人如同海邊的沙那樣多，都吃喝快樂。
1KGS|4|21|所羅門 統治諸國，從 大河 到 非利士 地，直到 埃及 的邊界。 所羅門 在世的日子，這些國都向他進貢，服事他。
1KGS|4|22|所羅門 每日所用的食物：三十歌珥細麵，六十歌珥粗麵，
1KGS|4|23|十頭肥牛，二十頭草場的牛，一百隻羊，還有鹿、羚羊、麃子，以及肥禽。
1KGS|4|24|所羅門 管理整個 大河 西邊，從 提弗薩 直到 迦薩 ，以及 大河 西邊的諸王，屬他的四境盡都平安。
1KGS|4|25|所羅門 在世的日子，從 但 到 別是巴 ， 猶大 和 以色列 各人都在自己的葡萄樹下和無花果樹下安然居住。
1KGS|4|26|所羅門 擁有給戰車用的四萬個 馬棚，還有一萬二千名騎兵。
1KGS|4|27|這些官員各按自己的月份供給 所羅門 王，以及一切與他同席之人的食物，一無所缺。
1KGS|4|28|他們各按其分，把給馬與快馬吃的大麥和乾草送到指定的地方去。
1KGS|4|29|上帝賜給 所羅門 極大的智慧和聰明，以及寬闊的心，如同海邊的沙。
1KGS|4|30|所羅門 的智慧超過所有東方人的智慧，和 埃及 人一切的智慧。
1KGS|4|31|他的智慧勝過萬人，勝過 以斯拉 人 以探 ，以及 瑪曷 的兒子 希幔 、 甲各 、 達大 。他的名聲傳遍四圍的列國。
1KGS|4|32|他作箴言三千句，詩歌一千零五首。
1KGS|4|33|他講論草木，從 黎巴嫩 的香柏樹直到牆上長的牛膝草，又講論飛禽、走獸、爬行動物和魚類。
1KGS|4|34|地上凡曾聽過他智慧的君王，都派人來；萬民都有人來聽 所羅門 的智慧。
1KGS|5|1|推羅 王 希蘭 是 大衛 平生的好友。 希蘭 聽見 以色列 人膏 所羅門 接續他父親作王，就派臣僕到他那裏。
1KGS|5|2|所羅門 也派人到 希蘭 那裏，說：
1KGS|5|3|「你知道我父親 大衛 因四圍的戰爭，不能為耶和華－他上帝的名建殿，直等到耶和華使仇敵都服在他腳下。
1KGS|5|4|現在耶和華－我的上帝使我四圍太平，沒有仇敵，沒有災禍。
1KGS|5|5|看哪，我吩咐要為耶和華－我上帝的名建殿，是照耶和華向我父親 大衛 說的：『我必使你兒子接續你，坐你的王位，他必為我的名建殿。』
1KGS|5|6|現在，請吩咐人在 黎巴嫩 為我砍伐香柏木，我的僕人必幫助你的僕人。至於你僕人的工錢，我必照你所定的給你。你知道，在我們中間沒有人像 西頓 人那樣擅長砍伐樹木。」
1KGS|5|7|希蘭 聽見 所羅門 的話，就很高興，說：「今日耶和華是應當稱頌的，因為他賜給 大衛 一個有智慧的兒子，治理這眾多的百姓。」
1KGS|5|8|希蘭 送信給 所羅門 ，說：「你派人向我所提的那事，我已聽見了；論到香柏木和松木，我必照你一切的心願去做。
1KGS|5|9|我的僕人必把這木料從 黎巴嫩 運到海裏，我會把它們紮成筏子浮在海上，運到你告訴我的地方，在那裏拆開，你就可以收取；你也要照我的心願做，把食物給我的家。」
1KGS|5|10|於是 希蘭 照 所羅門 的心願，給他香柏木和松木；
1KGS|5|11|所羅門 給 希蘭 二萬歌珥麥子，二十歌珥 搗成的油，作他家的食物。 所羅門 每年都是這樣給 希蘭 。
1KGS|5|12|耶和華照著所應許的賜智慧給 所羅門 。 希蘭 與 所羅門 和平相處，二人彼此立約。
1KGS|5|13|所羅門 王從全 以色列 挑取服勞役的人，徵來的人有三萬，
1KGS|5|14|派他們輪流每月一萬人上 黎巴嫩 去；一個月在 黎巴嫩 ，兩個月在家裏。 亞多尼蘭 管理他們。
1KGS|5|15|所羅門 有七萬扛抬的，八萬在山上鑿石頭的。
1KGS|5|16|此外， 所羅門 有三千三百個監督工作的官長，監管百姓做工。
1KGS|5|17|王下令，他們就鑿出又大又貴重的石頭來，用以立殿的根基。
1KGS|5|18|所羅門 的工匠和 希蘭 的工匠，以及 迦巴勒 人，把石頭鑿好，預備了木料和石頭來建殿。
1KGS|6|1|以色列 人出 埃及 地後四百八十年， 所羅門 作 以色列 王第四年西弗月，就是二月，他開工建造耶和華的殿。
1KGS|6|2|所羅門 王為耶和華所建的殿，長六十肘，寬二十肘，高三十肘。
1KGS|6|3|殿的正堂前走廊長二十肘，與殿的寬度一樣，殿前寬十肘；
1KGS|6|4|他為殿做了有框嵌壁式的窗戶。
1KGS|6|5|靠著殿牆，圍著外殿和內殿的牆，周圍建造了廂房；
1KGS|6|6|下層寬五肘，中層寬六肘，第三層寬七肘。他在殿牆的周圍造坎，免得梁木插入殿牆裏。
1KGS|6|7|殿是用山中鑿成的石頭建的，所以建殿的時候，鎚子、斧子和別樣鐵器的響聲都沒有聽見。
1KGS|6|8|在殿右邊當中的廂房有門，可以從螺旋梯上到中層，再從中層上到第三層。
1KGS|6|9|所羅門 完成殿的建造。他用香柏木作梁木和橫板，遮蓋殿頂。
1KGS|6|10|靠著整個殿所造的廂房，每層高五肘，香柏木的梁板擱在殿的牆坎上。
1KGS|6|11|耶和華的話臨到 所羅門 ，說：
1KGS|6|12|「論到你所建的這殿，你若遵行我的律例，謹守我的典章，遵從我的一切誡命，行在其中，我必向你應驗我所應許你父親 大衛 的話。
1KGS|6|13|我必住在 以色列 人中間，並不丟棄我的百姓 以色列 。」
1KGS|6|14|所羅門 完成殿的建造。
1KGS|6|15|他用香柏木板建造殿的內牆，從殿的地到牆頂 都貼上木板，又用松木板鋪地。
1KGS|6|16|他在殿的後部建了一間內殿，長二十肘，從地到牆 用香柏木板，作為至聖所。
1KGS|6|17|殿，就在內殿的前面 ，長四十肘。
1KGS|6|18|殿裏一點石頭都不顯露，一概用香柏木遮蔽；香柏木上刻著野瓜和綻開的花。
1KGS|6|19|他在殿的中間預備內殿，在那裏安放耶和華的約櫃。
1KGS|6|20|內殿 長二十肘，寬二十肘，高二十肘，都貼上純金。他又用香柏木做壇。
1KGS|6|21|所羅門 用純金貼殿內，又用金鏈子掛在內殿前，內殿也貼上金子。
1KGS|6|22|整個殿都貼上金子，直到貼滿；內殿前的整個壇，也都包上金子。
1KGS|6|23|他在內殿裏用橄欖木做兩個基路伯，各高十肘。
1KGS|6|24|這基路伯的一個翅膀長五肘，另一個翅膀長五肘，從一個翅膀尖到另一個翅膀尖共有十肘；
1KGS|6|25|第二個基路伯也是十肘；兩個基路伯的尺寸、形狀都一樣。
1KGS|6|26|這一個基路伯高十肘，第二個基路伯也是如此。
1KGS|6|27|他把兩個基路伯安在內殿中間。基路伯的翅膀是張開的，這基路伯的一個翅膀挨著這邊的牆，第二個基路伯的一個翅膀挨著那邊的牆，向內的兩個翅膀在殿中間彼此相接。
1KGS|6|28|二基路伯都包上金子。
1KGS|6|29|殿周圍的牆上全都刻著基路伯、棕樹和綻開的花，內外都是如此。
1KGS|6|30|殿的地板都貼上金子，內外都是如此。
1KGS|6|31|他用橄欖木製造內殿的入口、門楣和五邊形的門柱。
1KGS|6|32|在橄欖木做的兩門扇上刻著基路伯、棕樹和綻開的花，都貼上金子。基路伯和棕樹上也灑上金子。
1KGS|6|33|他又為外殿的入口，用橄欖木製造門柱，是四邊形的。
1KGS|6|34|他用松木做兩扇門。這一扇有兩葉摺疊，第二扇也有兩葉 摺疊。
1KGS|6|35|上面刻著基路伯、棕樹和綻開的花，雕刻物都均勻地貼上金子。
1KGS|6|36|他又用三層鑿成的石頭、香柏木一層建造內院。
1KGS|6|37|所羅門 在位第四年西弗月，立了耶和華殿的根基。
1KGS|6|38|到十一年布勒月，就是八月，殿和一切屬殿的都按著樣式造成。他建殿共用了七年。
1KGS|7|1|所羅門 為自己建造宮殿，十三年方才建成整座宮殿。
1KGS|7|2|他建造 黎巴嫩林宮 ，長一百肘，寬五十肘，高三十肘，有四行香柏木柱，柱上有香柏木橫梁；
1KGS|7|3|廂房以上覆蓋著香柏木，在四十五根柱子之上，每行十五根。
1KGS|7|4|窗戶有三排，三排的窗與窗相對。
1KGS|7|5|所有的門和門柱都有四方形的框，共有三行，彼此相對。
1KGS|7|6|他建造有柱子的廳，長五十肘，寬三十肘。在這前面有走廊，前面有柱子和頂蓋 。
1KGS|7|7|他又建造一個有座位的廳，就是審判廳，他在那裏審判；這廳的地板從這邊到那邊都鋪上香柏木。
1KGS|7|8|廳後面的院內有 所羅門 自己住的宮殿，都用同樣的建造方式。 所羅門 又為所娶法老的女兒建造一座宮，建造方式與這廳一樣。
1KGS|7|9|建造這一切所用的石頭都是貴重的，按著尺寸鑿成，用鋸子裏外鋸齊；從根基直到房檐，從外頭直到大院，都是如此。
1KGS|7|10|根基是貴重的大石頭，有長十肘的，有長八肘的；
1KGS|7|11|上面有香柏木和按著尺寸鑿成的貴重石頭。
1KGS|7|12|大院周圍有鑿成的石頭三層、香柏木板一層，都照耶和華殿的內院和殿的走廊的樣式。
1KGS|7|13|所羅門 王派人從 推羅 把 戶蘭 接來。
1KGS|7|14|他是 拿弗他利 支派中一個寡婦的兒子，父親是 推羅 人，是作銅匠的。 戶蘭 滿有智慧、聰明、技能，善作各樣的銅器。他來到 所羅門 王那裏，為王做一切的工。
1KGS|7|15|戶蘭 製造兩根銅柱，一根高十八肘，第二根柱子用繩子量，周圍是十二肘 ；
1KGS|7|16|他做了兩個柱頂安在柱上，是用銅鑄造的，一個柱頂高五肘，第二個柱頂也高五肘。
1KGS|7|17|柱子頂上有裝飾的網子和編成的鏈子，一個柱頂有七個，第二個柱頂也有七個。
1KGS|7|18|他做了柱子 ，第一根柱子的柱頂上，周圍有兩行網子在柱子 上面遮蓋柱頂，第二根柱頂也是這樣做。
1KGS|7|19|走廊柱子頂上的柱頂高四肘，刻著百合花。
1KGS|7|20|兩根柱子上面有柱頂，柱頂靠近網子的圓凸面上，有石榴的行列環繞著，共二百個，第二個柱頂也是如此。
1KGS|7|21|他把兩根柱子立在殿的走廊前：右邊立一根，起名叫 雅斤 ；左邊立一根，起名叫 波阿斯 。
1KGS|7|22|柱頂上刻著百合花。這樣，柱子的工程就完畢了。
1KGS|7|23|他又鑄一個銅海，周圍是圓的，直徑十肘，高五肘，用繩子量周圍是三十肘。
1KGS|7|24|銅海邊緣下面的周圍有野瓜的形狀，每肘十個，共兩行，繞著銅海，是造銅海的時候鑄上去的。
1KGS|7|25|銅海安在十二頭銅牛上：三頭向北，三頭向西，三頭向南，三頭向東。銅海安在牛上，牛尾都向內。
1KGS|7|26|銅海厚一掌，邊如杯邊，像百合花，容量是二千罷特。
1KGS|7|27|他用銅製造十個盆座，每座長四肘，寬四肘，高三肘。
1KGS|7|28|銅座的造法是這樣：周圍各有嵌邊，嵌邊裝在框架中。
1KGS|7|29|裝在框架中的嵌邊上有獅子和牛，以及基路伯。框架上有小座，獅子和牛的上面和下面有錘成的花紋浮雕。
1KGS|7|30|每座有四個銅輪和銅軸，它有四個支架在盆以下，這些支架是鑄成的，各邊都有花紋。
1KGS|7|31|它的口在柱頂裏，向上高一肘，口是圓的，做法如座一樣，直徑是一肘半，口上也有雕工。嵌邊是方形的，不是圓的。
1KGS|7|32|四個輪子在嵌邊以下，輪軸與座相連，每輪高一肘半。
1KGS|7|33|輪的樣式如同車的輪子；軸、輞、輻、轂都是鑄成的。
1KGS|7|34|每個座四邊有四個盆形的支架，這些支架是與座從一整塊鑄成的。
1KGS|7|35|座頂有圓架，高半肘；座頂有支柱和嵌邊，是與座從一整塊鑄成的。
1KGS|7|36|他在支柱和嵌邊上，每個空處刻上基路伯、獅子和棕樹，周圍有花紋。
1KGS|7|37|他按照這樣的做法造了十個盆座，它們的鑄法、尺寸、樣式全都相同。
1KGS|7|38|他又造十個銅盆，每盆的容量四十罷特，直徑四肘。在十個座上，每座安設一盆。
1KGS|7|39|他把五個安置在殿的右邊，五個安置在殿的左邊，又把銅海安置在殿的右旁，在東南邊。
1KGS|7|40|戶蘭 又造了盆、鏟子和盤子。這樣， 戶蘭 為 所羅門 王做完了耶和華殿一切的工：
1KGS|7|41|兩根柱子和柱子頂上兩個如碗的柱頂，以及蓋著如碗柱頂的兩個網子；
1KGS|7|42|四百個石榴，安在兩個網子上，每網兩行石榴，蓋著柱子上面兩個如碗的柱頂；
1KGS|7|43|十個盆座和其上的十個盆；
1KGS|7|44|銅海和其下的十二頭牛；
1KGS|7|45|盆、鏟子、盤子。 戶蘭 給 所羅門 王為耶和華殿造的這一切器皿都是用光亮的銅，
1KGS|7|46|是王在 約旦 平原、 疏割 和 撒拉但 中間的泥巴地鑄成的。
1KGS|7|47|所羅門 允許這一切器皿不過秤，因為所用的銅太多，重量無法計算。
1KGS|7|48|所羅門 又為耶和華的殿造了各樣的器皿：金壇和獻供餅的金供桌；
1KGS|7|49|內殿前的純金燈臺，右邊五個，左邊五個，以及其上的花、燈盞、燈剪，都是金的；
1KGS|7|50|純金的杯、鉗子、盤子、勺子 、火盆，以及聖殿的最裏面，就是至聖所的門樞和外殿的門樞，都是金的。
1KGS|7|51|所羅門 王做完了耶和華殿一切的工，就把他父親 大衛 分別為聖的金銀和器皿都帶來，放在耶和華殿的庫房裏。
1KGS|8|1|那時， 所羅門 召集 以色列 的長老、各支派的領袖和 以色列 人的族長到 耶路撒冷 ， 所羅門 王那裏，要把耶和華的約櫃從 大衛城 ，就是 錫安 ，接上來。
1KGS|8|2|以他念月，就是七月，在節期時，所有的 以色列 人都聚集到 所羅門 王那裏。
1KGS|8|3|以色列 眾長老一來到，祭司就抬起約櫃。
1KGS|8|4|祭司和 利未 人將耶和華的約櫃請上來，又把會幕和會幕一切的聖器皿都帶上來。
1KGS|8|5|所羅門 王和聚集到他那裏的 以色列 全會眾一同在約櫃前獻牛羊為祭，多得不可勝數，無法計算。
1KGS|8|6|祭司將耶和華的約櫃請進內殿，就是至聖所，安置在兩個基路伯的翅膀底下約櫃的地方。
1KGS|8|7|基路伯張開翅膀在約櫃上面的地方，從上面遮住約櫃和抬櫃的槓。
1KGS|8|8|這槓很長，從內殿前的聖所可以看見槓頭，從外面卻看不見。這槓直到今日還在那裏。
1KGS|8|9|約櫃裏沒有別的，只有兩塊石版，就是 以色列 人出 埃及 地，耶和華與他們立約的時候， 摩西 在 何烈山 放在那裏的。
1KGS|8|10|祭司從聖所出來的時候，有雲充滿耶和華的殿，
1KGS|8|11|祭司因雲彩的緣故不能站立供職，因為耶和華的榮光充滿了耶和華的殿。
1KGS|8|12|那時， 所羅門 說： 「耶和華曾說要住在幽暗之處 。
1KGS|8|13|我的確為你建了一座雄偉的殿宇， 作為你永遠居住的地方。」
1KGS|8|14|王轉過臉來為 以色列 全會眾祝福， 以色列 全會眾都站立。
1KGS|8|15|所羅門 說：「耶和華－ 以色列 的上帝是應當稱頌的！因他親口向我父 大衛 應許的，也親手成就了；他曾說：
1KGS|8|16|『自從那日我領我百姓 以色列 出 埃及 以來，我未曾在 以色列 各支派中選擇一城，在那裏為我的名建造殿宇，但我揀選 大衛 治理我的百姓 以色列 。』
1KGS|8|17|我父 大衛 的心意是要為耶和華－ 以色列 上帝的名建殿。
1KGS|8|18|耶和華卻對我父 大衛 說：『你有心為我的名建殿，這心意是好的；
1KGS|8|19|但你不可建殿，惟有你親生的兒子才可為我的名建殿。』
1KGS|8|20|現在耶和華實現了他所應許的話，使我接續我父 大衛 坐 以色列 的王位，正如耶和華所說的，我也為耶和華－ 以色列 上帝的名建造了這殿。
1KGS|8|21|我也在那裏為約櫃預備一處。約櫃那裏有耶和華的約，就是他領我們列祖出 埃及 地的時候，與他們所立的約。」
1KGS|8|22|所羅門 當著 以色列 全會眾，站在耶和華的壇前，向天舉手，
1KGS|8|23|說：「耶和華－ 以色列 的上帝啊，天上地下沒有神明可與你相比！你向那些盡心行在你面前的僕人守約施慈愛，
1KGS|8|24|這約是你向你僕人 大衛 守的，是你應許他的。你親口應許，親手成就，正如今日一樣。
1KGS|8|25|耶和華－ 以色列 的上帝啊，你向你僕人我父 大衛 應許說：『你的子孫若謹慎自己的行為，在我面前行事像你所行的一樣，就不斷有人在我面前坐 以色列 的王位。』現在求你信守這話。
1KGS|8|26|以色列 的上帝啊，現在求你成就向你僕人我父 大衛 所應許的話。
1KGS|8|27|「上帝果真住在地上嗎？看哪，天和天上的天尚且不足容納你，何況我所建的這殿呢？
1KGS|8|28|惟求耶和華－我的上帝垂顧僕人的禱告祈求，俯聽僕人今日在你面前的祈禱呼求。
1KGS|8|29|願你的眼目晝夜看顧這殿，就是你說要作為你名的居所；求你垂聽禱告，你僕人向此處的禱告。
1KGS|8|30|你僕人和你百姓 以色列 向此處祈禱的時候，求你在你天上的居所垂聽，垂聽而赦免。
1KGS|8|31|「人若得罪鄰舍，有人強迫他，要他起誓，他來到這殿，在你的壇前起誓，
1KGS|8|32|求你在天上垂聽、處理，向你的僕人施行審判，定惡人有罪，照他所行的報應在他頭上；定義人為義，照他的義賞賜他。
1KGS|8|33|「你的百姓 以色列 若得罪你，敗在仇敵面前，卻又歸向你，宣認你的名，在這殿裏向你祈求禱告，
1KGS|8|34|求你在天上垂聽，赦免你百姓 以色列 的罪，使他們歸回你賜給他們列祖的地。
1KGS|8|35|「你的百姓若得罪了你，你使天閉塞不下雨；他們若向此處禱告，宣認你的名，因你的懲罰而離開他們的罪，
1KGS|8|36|求你在天上垂聽，赦免你僕人你百姓 以色列 的罪，將當行的善道教導他們，並降雨在你的地，就是你賜給你百姓為業之地。
1KGS|8|37|「這地若有饑荒、瘟疫、焚風 、霉爛、蝗蟲、螞蚱，或有仇敵圍困這地的 城門，無論遭遇甚麼災禍疾病，
1KGS|8|38|你的百姓 以色列 ，或眾人或一人，內心知道有禍，向這殿舉手，無論祈求甚麼，禱告甚麼，
1KGS|8|39|求你在天上你的居所垂聽、赦免、處理。因為你知道人心，惟有你知道世人的心，求你照各人所行的一切待他們，
1KGS|8|40|使他們在你賜給我們列祖的土地上一生一世敬畏你。
1KGS|8|41|「論到不屬你百姓 以色列 的外邦人，若為你的名從遠方而來，
1KGS|8|42|他們因聽見你的大名和大能的手，以及伸出來的膀臂，來向這殿禱告，
1KGS|8|43|求你在天上你的居所垂聽，照著外邦人向你所求的一切而行，使地上萬民都認識你的名，敬畏你，像你的百姓 以色列 一樣，又使他們知道我所建造的是稱為你名下的殿。
1KGS|8|44|「你的百姓若奉你的派遣出去，無論往何處與仇敵爭戰，他們若向耶和華所選擇的城，以及我為你名所建造的這殿禱告，
1KGS|8|45|求你在天上垂聽他們的禱告祈求，為他們伸張正義。
1KGS|8|46|「你的百姓若得罪你，因為沒有人不犯罪，你向他們發怒，把他們交在仇敵面前，擄他們的人把他們帶到仇敵之地，或遠或近，
1KGS|8|47|他們若在被擄之地那裏回心轉意，在擄掠者之地悔改，向你懇求說：『我們有罪了，我們悖逆了，我們作惡了』；
1KGS|8|48|他們若在擄他們的仇敵之地盡心盡性歸向你，又向自己的地，就是你賜給他們列祖的地和你所選擇的城，以及我為你名所建造的這殿禱告，
1KGS|8|49|求你在天上你的居所垂聽他們的禱告祈求，為他們伸張正義，
1KGS|8|50|饒恕得罪你的子民，赦免他們向你所犯一切的過犯，使他們在擄他們的人面前蒙憐憫。
1KGS|8|51|因為他們是你的子民，你的產業，是你從 埃及 ，從鐵爐中領出來的。
1KGS|8|52|願你的眼目看顧僕人和你百姓 以色列 的祈求；他們無論何時向你呼求，願你垂聽。
1KGS|8|53|主耶和華啊，你將他們從地上萬民中分別出來作你的產業，是照著你領我們列祖出 埃及 的時候，藉你僕人 摩西 所應許的。」
1KGS|8|54|所羅門 在耶和華的壇前屈膝跪著，向天舉手；他在耶和華面前禱告祈求完畢的時候，就起來，
1KGS|8|55|站著，大聲為 以色列 全會眾祝福，說：
1KGS|8|56|「耶和華是應當稱頌的！因為他照著一切所應許的賜平安給他的百姓 以色列 ，凡藉他僕人 摩西 應許賜福的話，一句都沒有落空。
1KGS|8|57|願耶和華－我們的上帝與我們同在，像與我們列祖同在一樣，不撇下我們，不丟棄我們，
1KGS|8|58|使我們的心歸向他，遵行他一切的道，謹守他吩咐我們列祖的誡命、律例、典章。
1KGS|8|59|願我在耶和華面前祈求的這些話，晝夜靠近耶和華－我們的上帝，好讓他每日為他僕人和他百姓 以色列 伸張正義，
1KGS|8|60|使地上的萬民都知道惟獨耶和華是上帝，沒有別的了。
1KGS|8|61|所以你們當向耶和華－我們的上帝存純正的心，遵行他的律例，謹守他的誡命，如同今日一樣。」
1KGS|8|62|王和全 以色列 一同在耶和華面前獻祭。
1KGS|8|63|所羅門 向耶和華獻平安祭，二萬二千頭牛，十二萬隻羊。這樣，王和全 以色列 為耶和華的殿行了奉獻之禮。
1KGS|8|64|當日，王因耶和華殿前的銅壇太小，容不下燔祭、素祭和平安祭牲的脂肪，就將耶和華殿前院子的中間分別為聖，在那裏獻燔祭、素祭和平安祭牲的脂肪。
1KGS|8|65|那時 所羅門 守節，從 哈馬口 直到 埃及 溪谷的 以色列 眾人都與他同在一起，成了一個盛大的會，在耶和華－我們的上帝面前七日又七日，共十四日。
1KGS|8|66|第八日，王遣散百姓；他們都為王祝福。他們為耶和華向他僕人 大衛 和他百姓 以色列 所施的一切恩惠都心中喜樂，愉快地各回自己的帳棚去了。
1KGS|9|1|所羅門 建造耶和華的殿和王宮，以及一切所想要建造的都完畢了，
1KGS|9|2|耶和華第二次向 所羅門 顯現，如先前在 基遍 向他顯現一樣。
1KGS|9|3|耶和華對他說：「我已聽了你在我面前的禱告和祈求，將你所建的這殿分別為聖，使我的名永遠立在那裏；我的眼、我的心也必時常在那裏。
1KGS|9|4|你若以純正的心和正直行在我面前，效法你父 大衛 所行的，遵行我一切所吩咐你的，謹守我的律例典章，
1KGS|9|5|我就必堅固你在 以色列 國度的王位，直到永遠，正如我應許你父 大衛 說：『你的子孫必不斷有人坐 以色列 的王位。』
1KGS|9|6|倘若你們和你們的子孫轉去不跟從我，不守我擺在你們面前的誡命律例，去事奉別神，敬拜它們，
1KGS|9|7|我就必把 以色列 從我賜給他們的地上剪除，也必從我面前捨棄那為我名所分別為聖的殿，使 以色列 在萬民中成為笑柄，被人譏誚。
1KGS|9|8|這殿雖然崇高 ，將來凡經過的人必驚訝，嗤笑，說：『耶和華為何向這地和這殿如此行呢？』
1KGS|9|9|人必說：『因為此地的人離棄領他們祖先出 埃及 地的耶和華－他們的上帝，去親近別神，敬拜事奉它們，所以耶和華使這一切災禍臨到他們。』」
1KGS|9|10|所羅門 建造耶和華殿和王宮這兩座殿宇，用了二十年才完成。
1KGS|9|11|推羅 王 希蘭 曾照 所羅門 所要的資助他香柏木、松木和金子， 所羅門 王就把 加利利 地的二十座城給了 希蘭 。
1KGS|9|12|希蘭 從 推羅 出來，察看 所羅門 給他的城鎮，看不順眼，
1KGS|9|13|就說：「我兄啊，你給我的是甚麼城鎮呢？」他就給這些城鎮起名叫 迦步勒 地，直到今日。
1KGS|9|14|希蘭 曾給 所羅門 一百二十他連得金子。
1KGS|9|15|所羅門 王挑取服勞役的工人，為要建造耶和華的殿、自己的宮、 米羅 、 耶路撒冷 的城牆、 夏瑣 、 米吉多 和 基色 。
1KGS|9|16|先前 埃及 王法老上來攻取 基色 ，用火焚燒，殺了城內居住的 迦南 人，把城賜給他的女兒，就是 所羅門 的妻子，作為嫁妝。
1KGS|9|17|所羅門 建造 基色 、 下伯‧和崙 、
1KGS|9|18|巴拉 ，和位於境內曠野的 達莫 。
1KGS|9|19|所羅門 建造一切的儲貨城、戰車城、戰馬城，以及他所想要建造的，在 耶路撒冷 、 黎巴嫩 和自己治理全國中的一切建設。
1KGS|9|20|至於所有剩下的百姓，不屬 以色列 人的 亞摩利 人、 赫 人、 比利洗 人、 希未 人、 耶布斯 人，
1KGS|9|21|那些 以色列 人在當地不能滅盡的人， 所羅門 徵召他們剩下的後代作服勞役的奴僕，直到今日。
1KGS|9|22|惟有 以色列 人， 所羅門 不使他們作奴僕，而是作他的戰士、臣僕、官長、軍官、戰車長、騎兵長。
1KGS|9|23|這些是 所羅門 工程的五百五十個監工，他們在百姓中監管作工的人。
1KGS|9|24|法老的女兒從 大衛城 上到 所羅門 為她建造的宮裏。那時， 所羅門 才建造 米羅 。
1KGS|9|25|所羅門 每年三次在他為耶和華所築的壇上獻燔祭和平安祭，又在耶和華面前的壇上燒香。這樣，他完成了建殿。
1KGS|9|26|所羅門 王在 以東 地 紅海 邊，靠近 以祿 的 以旬‧迦別 製造船隻。
1KGS|9|27|希蘭 派他的僕人，就是熟悉航海的船員，與 所羅門 的僕人一同坐船航海。
1KGS|9|28|他們到了 俄斐 ，從那裏得了四百二十他連得金子，運到 所羅門 王那裏。
1KGS|10|1|示巴 女王聽見 所羅門 因耶和華的名所得的名聲，就來要用難題考問 所羅門 。
1KGS|10|2|她帶著很多的隨從來到 耶路撒冷 ，有駱駝馱著香料、極多金子和寶石。她來到 所羅門 那裏，向他提出心中所有的問題。
1KGS|10|3|所羅門 回答了她所有的問題，沒有一個問題太難，王不能向她解答的。
1KGS|10|4|示巴 女王看見 所羅門 一切的智慧，和他所建造的宮殿，
1KGS|10|5|席上的食物，坐著的群臣，侍立的僕人，他們的服裝，和他的司酒長，以及他在耶和華殿裏所獻的燔祭 ，就詫異得神不守舍。
1KGS|10|6|她對王說：「我在本國所聽到的話，論到你的事和你的智慧是真的！
1KGS|10|7|我本來不信那些話，及至我來親眼看見了，看哪，人所告訴我的還不到一半，你的智慧和你的福分超過我所聽見的傳聞。
1KGS|10|8|你的人 是有福的！你這些僕人常侍立在你面前、聽你智慧的話是有福的！
1KGS|10|9|耶和華－你的上帝是應當稱頌的！他喜愛你，使你坐 以色列 的王位，因為他永遠愛 以色列 ，所以立你作王，使你秉公行義。」
1KGS|10|10|於是， 示巴 女王把一百二十他連得金子、極多的香料和寶石送給 所羅門 王；送來的香料，從來沒有像 示巴 女王送給他的那麼多。
1KGS|10|11|希蘭 的船隻也從 俄斐 運了金子來，又從 俄斐 運了許多檀香木和寶石來。
1KGS|10|12|王用檀香木為耶和華的殿和王宮做欄杆，又為歌唱的人做琴瑟。以後再沒有這樣的檀香木運進來，也再沒有人見過，直到如今。
1KGS|10|13|所羅門 王除了照自己的厚意餽贈 示巴 女王之外，凡她所提出的一切要求， 所羅門 王都送給她。於是女王和她臣僕轉回，到本國去了。
1KGS|10|14|所羅門 每年所得的金子，重六百六十六他連得；
1KGS|10|15|另外還有來自商人 和做生意的商品，以及 阿拉伯 諸王和各地省長的。
1KGS|10|16|所羅門 王用錘出來的金子打成二百面盾牌，每面盾牌用六百舍客勒金子；
1KGS|10|17|又用錘出來的金子打成三百面小盾牌，每面小盾牌用三彌那金子。王把它們放在 黎巴嫩林宮 裏。
1KGS|10|18|王又製造一個大的象牙寶座，包上純金。
1KGS|10|19|寶座有六層臺階，座的後背是圓的，座位之處兩旁有扶手，靠近扶手有兩隻獅子站立。
1KGS|10|20|六層臺階上有十二隻獅子站立，分站左邊和右邊；任何國度都沒有這樣做的。
1KGS|10|21|所羅門 王一切的飲器都是金的， 黎巴嫩林宮 裏所有的器皿都是純金的。在 所羅門 的日子，銀子算不了甚麼。
1KGS|10|22|王有 他施 船隻與 希蘭 的船隻一同航海， 他施 船隻每三年一次把金、銀、象牙、猿猴、孔雀 運回來。
1KGS|10|23|所羅門 王的財寶與智慧勝過地上的眾王。
1KGS|10|24|全地都求見 所羅門 的面，要聽上帝放在他心裏的智慧。
1KGS|10|25|他們各帶貢物，就是銀器、金器、衣服、兵器、香料、馬、騾子，每年都有一定的數量。
1KGS|10|26|所羅門 聚集戰車騎兵；他有一千四百輛戰車，一萬二千名騎兵，安置在屯車城，在 耶路撒冷 的王那裏。
1KGS|10|27|王在 耶路撒冷 使銀子多如石頭，香柏木多如 謝非拉 的桑樹。
1KGS|10|28|所羅門 的馬是從 埃及 和 科威 運來的，是王的商人按著定價從 科威 買來的。
1KGS|10|29|從 埃及 進口的戰車，每輛六百舍客勒銀子，馬每匹一百五十舍客勒； 赫 人眾王和 亞蘭 諸王的戰車和馬，也是經由他們的手出口的。
1KGS|11|1|所羅門 王在法老的女兒之外，又寵愛許多外邦女子，就是 摩押 女子、 亞捫 女子、 以東 女子、 西頓 女子、 赫 人女子。
1KGS|11|2|論到這些國的人，耶和華曾吩咐 以色列 人說：「你們不可跟他們通婚，他們也不可跟你們在一起，因為他們一定會誘惑你們的心去隨從他們的神明。」 所羅門 卻為了愛，緊緊跟從他們。
1KGS|11|3|所羅門 娶七百個公主，三百個妃嬪。這些妻妾誘惑他的心。
1KGS|11|4|所羅門 年老的時候，他的妻妾誘惑他的心去隨從別神，不像他父親 大衛 以純正的心順服耶和華－他的上帝。
1KGS|11|5|所羅門 隨從 西頓 人的女神 亞斯她錄 和 亞捫 人可憎的 米勒公 。
1KGS|11|6|所羅門 行耶和華眼中看為惡的事，不像他父親 大衛 專心順從耶和華。
1KGS|11|7|那時， 所羅門 為 摩押 可憎的 基抹 和 亞捫 人可憎的 摩洛 ，在 耶路撒冷 對面的山上建造丘壇。
1KGS|11|8|他為所有的妻妾，就是那些向自己神明燒香獻祭的外邦女子，也是這樣做。
1KGS|11|9|耶和華向 所羅門 發怒，因為他的心偏離了向他顯現兩次的耶和華－ 以色列 的上帝。
1KGS|11|10|耶和華曾吩咐他這件事，不可隨從別神，他卻沒有遵守耶和華所吩咐的。
1KGS|11|11|所以耶和華對他說：「你既然是這樣，不遵守我所吩咐你守的約和律例，我必定把國度撕裂離開你，將它賜給你的大臣。
1KGS|11|12|然而，因你父親 大衛 的緣故，我不在你的日子行這事，而要從你兒子的手中撕裂這國。
1KGS|11|13|只是我不撕裂全國，卻要因我僕人 大衛 和我所選擇的 耶路撒冷 ，保留一個支派給你的兒子。」
1KGS|11|14|耶和華使 以東 人 哈達 興起，作 所羅門 的敵人；他是 以東 王的後裔。
1KGS|11|15|大衛 在 以東 的時候， 約押 元帥上去埋葬陣亡的人，殺了 以東 所有的男丁。
1KGS|11|16|約押 和 以色列 眾人在 以東 住了六個月，直到把 以東 的男丁盡都剪除。
1KGS|11|17|那時 哈達 還是幼童；他和他父親的臣僕，以及幾個 以東 人逃往 埃及 。
1KGS|11|18|他們從 米甸 起行，到了 巴蘭 ，再從 巴蘭 帶著幾個人來到 埃及 ，到 埃及 王法老那裏。法老給他房屋，吩咐給他糧食，又把地賜給他。
1KGS|11|19|哈達 在法老眼前大蒙恩寵，法老就把王后 答比匿 的妹妹嫁給他。
1KGS|11|20|答比匿 的妹妹給 哈達 生了一個兒子，叫 基努拔 。 答比匿 使 基努拔 在法老的宮裏斷奶， 基努拔 就與法老的眾子一同住在法老的宮裏。
1KGS|11|21|哈達 在 埃及 聽見 大衛 與他祖先同睡， 約押 元帥也死了，就對法老說：「請你讓我走，我要回本國去。」
1KGS|11|22|法老對他說：「你在我這裏有甚麼缺乏？看哪，你竟想要回你本國去！」他說：「我沒有缺乏甚麼，只是懇求王准我回去。」
1KGS|11|23|上帝又使 以利亞大 的兒子 利遜 興起，作 所羅門 的敵人。他曾逃避主人 瑣巴 王 哈大底謝 。
1KGS|11|24|大衛 擊殺 瑣巴 人的時候， 利遜 召集了一群人，自己作他們的領袖。他們往 大馬士革 ，住在那裏，在 大馬士革 建立王國。
1KGS|11|25|所羅門 活著的時候，除了 哈達 為患之外， 利遜 也作 以色列 的敵人。他憎恨 以色列 ，作了 亞蘭 人的王。
1KGS|11|26|尼八 的兒子 耶羅波安 也舉起手來攻擊王。他是 所羅門 的臣僕， 以法蓮 支派的 洗利達 人；他母親是個寡婦，名叫 洗魯阿 。
1KGS|11|27|他舉手攻擊王是因先前 所羅門 建造 米羅 ，修補他父親 大衛城 缺口的這件事。
1KGS|11|28|耶羅波安 是個大有才能的人。 所羅門 見這青年殷勤，就派他監管 約瑟 家所有服勞役的工人。
1KGS|11|29|那時， 耶羅波安 出了 耶路撒冷 ， 示羅 人 亞希雅 先知在路上遇見他； 亞希雅 身上穿著一件新衣。田野中只有他們二人，沒有其他的人。
1KGS|11|30|亞希雅 拿起穿在自己身上的新衣，把它撕成十二片，
1KGS|11|31|對 耶羅波安 說：「你可以拿十片。耶和華－ 以色列 的上帝如此說：『看哪，我必從 所羅門 手裏撕裂這國，把十個支派賜給你。
1KGS|11|32|我因我僕人 大衛 和我在 以色列 眾支派中所選擇的 耶路撒冷城 的緣故，仍為 所羅門 留一個支派。
1KGS|11|33|因為他們 離棄我，敬拜 西頓 人的女神 亞斯她錄 、 摩押 的神明 基抹 和 亞捫 人的神明 米勒公 ，沒有像他父親 大衛 一樣遵從我的道，行我眼中看為正的事，守我的律例典章。
1KGS|11|34|但我不從他手裏奪走整個國家，卻使他在活著的日子作君王，是因我所揀選的僕人 大衛 遵守我的誡命律例。
1KGS|11|35|我必從他兒子手裏將王國奪走，賜給你十個支派，
1KGS|11|36|只留一個支派給他的兒子，使我僕人 大衛 在我所選擇立我名的 耶路撒冷城 那裏，在我面前常有燈光。
1KGS|11|37|我選你，使你照你心裏一切所願的作王，成為 以色列 的王。
1KGS|11|38|你若聽從我一切所吩咐你的，遵行我的道，行我眼中看為正的事，謹守我的律例誡命，像我僕人 大衛 所行的，我就與你同在，為你立堅固的家，像我為 大衛 所立的一樣，將 以色列 賜給你。
1KGS|11|39|我必因這事使 大衛 的後裔遭受患難，但不是永遠的。』」
1KGS|11|40|所羅門 想要殺 耶羅波安 ， 耶羅波安 起身逃往 埃及 。他到了 埃及 王 示撒 那裏，就住在 埃及 ，直到 所羅門 死了。
1KGS|11|41|所羅門 其餘的事，凡他所做的和他的智慧，不都寫在《所羅門記》上嗎？
1KGS|11|42|所羅門 在 耶路撒冷 作全 以色列 的王四十年。
1KGS|11|43|所羅門 與他祖先同睡，葬在他父親 大衛 的城裏，他兒子 羅波安 接續他作王。
1KGS|12|1|羅波安 往 示劍 去，因 以色列 眾人都到了 示劍 ，要立他作王。
1KGS|12|2|尼八 的兒子 耶羅波安 先前躲避 所羅門 王，逃往 埃及 ，住在那裏。他還在 埃及 ，聽見了這事 ，
1KGS|12|3|以色列 人派人去請他來。 耶羅波安 就和 以色列 全會眾來，與 羅波安 談話，說：
1KGS|12|4|「你父親使我們負重軛，現在求你減輕你父親所加給我們的苦工和重軛，我們就服事你。」
1KGS|12|5|羅波安 對他們說：「你們走吧，過三天再來見我。」百姓就走了。
1KGS|12|6|羅波安 的父親 所羅門 在世的日子，有侍立在他面前的長者， 羅波安 王和他們商議，說：「你們出個主意，好把話帶回給這百姓。」
1KGS|12|7|他們對他說：「現在王若像僕人一樣服事這百姓，用好話回覆他們，他們就永遠作王的僕人了。」
1KGS|12|8|王不採納長者給他出的主意，卻和那些與他一同長大、在他面前侍立的年輕人商議。
1KGS|12|9|他對他們說：「這百姓對我說：『你父親使我們負重軛，求你減輕一些。』你們出個甚麼主意，我們好把話帶回給他們。」
1KGS|12|10|那些與他一同長大的年輕人對他說：「這百姓對王說：『你父親使我們負重軛，求你給我們減輕一些。』王要對他們如此說：『我的小指頭比我父親的腰還粗呢！
1KGS|12|11|我父親使你們負重軛，現在我必使你們負更重的軛！我父親用鞭子懲罰你們，我要用蠍子懲罰你們！』」
1KGS|12|12|耶羅波安 和眾百姓遵照王所說「你們第三天再來見我」的話，第三天來到 羅波安 那裏。
1KGS|12|13|王嚴厲地回答百姓，不採納長者給他出的主意。
1KGS|12|14|他照著年輕人所出的主意對他們說：「我父親使你們負重軛，我必使你們負更重的軛！我父親用鞭子懲罰你們，我卻要用蠍子懲罰你們！」
1KGS|12|15|王不依從百姓，因這事件是出於耶和華，為要應驗耶和華藉 示羅 人 亞希雅 對 尼八 的兒子 耶羅波安 所說的話。
1KGS|12|16|以色列 眾人見王不依從他們，百姓就回話給王，說： 「我們在 大衛 中有甚麼份呢？ 我們在 耶西 的兒子中沒有產業！ 以色列 啊，回你的帳棚去吧！ 大衛 啊，現在你顧自己的家吧！」 於是， 以色列 人都回自己的帳棚去了；
1KGS|12|17|至於住 猶大 城鎮的 以色列 人， 羅波安 仍作他們的王。
1KGS|12|18|羅波安 王派監管勞役的 亞多蘭 去， 以色列 眾人用石頭打他，他就死了。 羅波安 王急忙上車，逃回 耶路撒冷 去了。
1KGS|12|19|這樣， 以色列 背叛 大衛 家，直到今日。
1KGS|12|20|以色列 眾人聽見 耶羅波安 回來了，就派人去請他到會眾那裏，立他作全 以色列 的王。除了 猶大 支派，沒有跟從 大衛 家的。
1KGS|12|21|羅波安 來到 耶路撒冷 ，召集了 猶大 全家和 便雅憫 支派的人共十八萬，都是精選的戰士，要與 以色列 家打仗，好將王國奪回，歸 所羅門 的兒子 羅波安 。
1KGS|12|22|但上帝的話臨到神人 示瑪雅 ，說：
1KGS|12|23|「你去告訴 所羅門 的兒子 猶大 王 羅波安 ， 猶大 和 便雅憫 全家，以及其餘的百姓，說：
1KGS|12|24|『耶和華如此說：你們不可上去與你們的弟兄 以色列 人打仗。你們各自回家去吧！因為這事是出於我。』」眾人就聽從耶和華的話，遵照耶和華的話回去了。
1KGS|12|25|耶羅波安 在 以法蓮 山區建了 示劍 ，住在其中，又從 示劍 出去，建了 毗努伊勒 。
1KGS|12|26|耶羅波安 心裏說：「現在，這國恐怕仍會歸 大衛 家；
1KGS|12|27|這百姓若上 耶路撒冷 去，在耶和華的殿裏獻祭，他們的心必歸向他們的主 猶大 王 羅波安 。他們會殺了我，仍歸 猶大 王 羅波安 。」
1KGS|12|28|耶羅波安 王就籌劃，鑄造了兩個金牛犢，對眾百姓說：「你們上 耶路撒冷 去實在夠久了。 以色列 啊，看哪，這是領你出 埃及 地的神明。」
1KGS|12|29|他把一個安置在 伯特利 ，另一個安置在 但 。
1KGS|12|30|這事使百姓陷入罪裏，因為他們甚至到 但 去拜那牛犢。
1KGS|12|31|耶羅波安 在一些丘壇建神殿，立不屬 利未 人的平民百姓為祭司。
1KGS|12|32|耶羅波安 定八月十五日為節期，像在 猶大 的節期一樣，自己上壇獻祭。他在 伯特利 這樣做，向他所鑄的牛犢獻祭，又把他所立丘壇的祭司安置在 伯特利 。
1KGS|12|33|他在八月十五日，就是他自己心中所定的月份，在 伯特利 上到自己所造的祭壇；他為 以色列 人定了一個節期，親自上壇燒香。
1KGS|13|1|看哪，有一個神人遵照耶和華的話從 猶大 來到 伯特利 。 耶羅波安 正站在壇旁燒香；
1KGS|13|2|神人遵照耶和華的話向壇呼叫，說：「壇哪，壇哪！耶和華如此說：『看哪， 大衛 家必生一個兒子，名叫 約西亞 ，他必將在你上面燒香的丘壇祭司，宰殺在你上面，人的骨頭也必燒在你上面。』」
1KGS|13|3|當日，神人設個預兆，說：「這是耶和華說的預兆：『看哪，這壇必破裂，壇上的灰必傾倒出來。』」
1KGS|13|4|耶羅波安 王聽見神人向 伯特利 的壇呼叫的話，就從壇上伸手，說：「拿住他！」王向神人所伸的手卻萎縮了，不能彎回。
1KGS|13|5|壇也破裂了，壇上的灰傾倒出來，正如神人遵照耶和華的話所設的預兆。
1KGS|13|6|王對神人說：「請你為我禱告，向耶和華－你的上帝懇求恩惠，使我的手復原。」於是神人向耶和華懇求，王的手就復原了，如平常一樣。
1KGS|13|7|王對神人說：「請你跟我回宮，讓你恢復心力，我必給你賞賜。」
1KGS|13|8|神人對王說：「你就是把你一半的王宮給我，我也不跟你進去，也不在這地方吃飯喝水，
1KGS|13|9|因為耶和華的話這樣吩咐我說：『不可吃飯喝水，也不可從你去的原路回來。』」
1KGS|13|10|於是神人從別的路回去，不從他到 伯特利 來的原路回去。
1KGS|13|11|有一個老先知住在 伯特利 ，他的兒子來，把神人當日在 伯特利 所做的一切事和他向王所說的話，都告訴了父親。
1KGS|13|12|父親對他們說：「神人從哪條路去了呢？」他的兒子都看到 從 猶大 來的神人所去的路。
1KGS|13|13|老先知吩咐兒子說：「你們為我備驢。」他們備好了驢，他就騎上，
1KGS|13|14|去追神人，遇見神人坐在橡樹底下，就對他說：「你是不是從 猶大 來的神人？」他說：「是我。」
1KGS|13|15|老先知對他說：「請你跟我一起回家吃飯。」
1KGS|13|16|神人說：「我不能跟你回去，與你同行，也不能在這地方跟你一起吃飯喝水，
1KGS|13|17|因為有耶和華的話吩咐我說：『你在那裏不可吃飯喝水，也不可從你去的原路回來。』」
1KGS|13|18|老先知對他說：「我也是先知，和你一樣。有天使遵照耶和華的話對我說：『你去帶他一同回你的家，給他吃飯喝水。』」老先知在欺騙他。
1KGS|13|19|於是神人跟老先知回去，在他家裏吃飯喝水。
1KGS|13|20|他們坐席的時候，耶和華的話臨到那帶神人回來的先知，
1KGS|13|21|他就對從 猶大 來的神人宣告說：「耶和華如此說：『你既違背耶和華的指示，不遵守耶和華－你上帝的命令，
1KGS|13|22|反倒回來，在耶和華禁止你吃飯喝水的地方吃了飯喝了水，因此你的屍體必不得葬在你祖先的墳墓裏。』」
1KGS|13|23|神人吃喝完了，老先知為他帶回來的先知備驢。
1KGS|13|24|神人就去了，在路上有隻獅子遇見他，把他咬死。他的屍體倒在路上，驢站在屍體旁邊，獅子也站在屍體旁邊。
1KGS|13|25|看哪，有人經過，看見屍體倒在路上，獅子站在屍體旁邊，就來到老先知所住的城裏述說這事。
1KGS|13|26|那帶神人回來的先知聽見了，就說：「這是那違背了耶和華指示的神人，所以耶和華把他交給獅子；獅子撕裂他，咬死他，正如耶和華對他說的話。」
1KGS|13|27|老先知吩咐他兒子說：「你們為我備驢。」他們就備了驢。
1KGS|13|28|他去了，發現神人的屍體倒在路上，驢和獅子站在屍體旁邊，獅子卻沒有吃屍體，也沒有撕裂驢。
1KGS|13|29|老先知把神人的屍體抬起，馱在驢上，帶回自己的城裏，要為他哀哭，為他安葬。
1KGS|13|30|老先知把屍體葬在自己的墳裏，為他哀哭，說：「哀哉！我的弟兄啊！」
1KGS|13|31|安葬之後，老先知對他兒子說：「我死了，你們要把我葬在神人所葬的墳裏，使我的屍骨在他的屍骨旁邊，
1KGS|13|32|因為他遵照耶和華的話，指著 伯特利 的壇和 撒瑪利亞 各城丘壇神殿所宣告的話必定應驗。」
1KGS|13|33|這事以後， 耶羅波安 仍不離開他的惡道，立平民百姓為丘壇的祭司；凡願意的，他都分別為聖，立為丘壇的祭司。
1KGS|13|34|這事使 耶羅波安 的家陷入罪裏，甚至他的家被剪除，從地面上消滅了。
1KGS|14|1|那時， 耶羅波安 的兒子 亞比雅 病了。
1KGS|14|2|耶羅波安 對他的妻子說：「你起來改裝，使人認不出你是 耶羅波安 的妻子。你往 示羅 去，看哪，那裏有先知 亞希雅 ，他曾告訴我說，你必作這百姓的王。
1KGS|14|3|現在你手裏要帶十個餅、幾個薄餅和一瓶蜜到他那裏去，他必告訴你，孩子會怎樣。」
1KGS|14|4|耶羅波安 的妻子就照樣做，起身往 示羅 去，到了 亞希雅 的家。 亞希雅 因年紀老邁，兩眼發直，不能看見。
1KGS|14|5|耶和華對 亞希雅 說：「看哪， 耶羅波安 的妻子來問你她兒子的事，因她兒子病了，你當如此如此告訴她。她進來的時候會扮成別的婦人。」
1KGS|14|6|她剛進門， 亞希雅 聽見她的腳步聲，就說：「 耶羅波安 的妻子，進來吧！你為何扮成別的婦人呢？我奉差遣將凶信告訴你。
1KGS|14|7|你回去告訴 耶羅波安 說：『耶和華－ 以色列 的上帝如此說：我從百姓中提拔了你，立你作我百姓 以色列 的君王，
1KGS|14|8|將 大衛 家的國撕裂，賜給你，你卻不效法我僕人 大衛 ，遵守我的誡命，全心順從我，行我眼中看為正的事。
1KGS|14|9|你反倒行惡，比在你之前所有的人更嚴重；你離開了我，為自己立了別神，鑄了偶像，惹我發怒，將我丟在背後。
1KGS|14|10|因此，看哪，我必使災禍臨到 耶羅波安 的家，把屬 耶羅波安 的男丁，無論是奴役的、自由的，都從 以色列 中剪除。我必除滅 耶羅波安 的家，如同人掃除糞土，直到消滅。
1KGS|14|11|凡屬 耶羅波安 的人，死在城中的必被狗吃，死在田野的必被空中的鳥吃。這是耶和華說的。』
1KGS|14|12|你起身回家去吧！你的腳一進城，孩子就死了。
1KGS|14|13|以色列 眾人必為他哀哭，為他安葬。凡屬 耶羅波安 的人，只有他可以葬入墳墓，因為在 耶羅波安 的家中，只有他向耶和華－ 以色列 的上帝表現出好的行為。
1KGS|14|14|耶和華必另立一王治理 以色列 ，這一天，他必剪除 耶羅波安 的家；甚麼時候呢？現在就是了。
1KGS|14|15|耶和華必擊打 以色列 ，使他們搖動，像水中的蘆葦一樣，又將他們從耶和華賜給他們列祖的美地上拔出來，分散在 大河 那邊，因為他們造了 亞舍拉 ，惹耶和華發怒。
1KGS|14|16|因 耶羅波安 所犯的罪，又因他使 以色列 陷入罪裏，耶和華必將 以色列 交出來。」
1KGS|14|17|耶羅波安 的妻子起身回去，到了 得撒 ，剛到門檻，孩子就死了。
1KGS|14|18|以色列 眾人為他安葬，為他哀哭，正如耶和華藉他僕人 亞希雅 先知所說的話。
1KGS|14|19|耶羅波安 其餘的事，他怎樣打仗，怎樣作王，看哪，都寫在《以色列諸王記》上。
1KGS|14|20|耶羅波安 作王二十二年，就與他祖先同睡，他兒子 拿答 接續他作王。
1KGS|14|21|所羅門 的兒子 羅波安 作 猶大 王。他登基的時候年四十一歲，在 耶路撒冷 ，就是耶和華從 以色列 眾支派中所選擇立他名的城，作王十七年。 羅波安 的母親名叫 拿瑪 ，是 亞捫 人。
1KGS|14|22|猶大 人行耶和華眼中看為惡的事，以所犯的罪惹動他的妒忌，比他們的祖先所犯的一切更嚴重。
1KGS|14|23|因為他們在各高岡上，各青翠樹下築丘壇，立柱像和 亞舍拉 。
1KGS|14|24|國中也有男的廟妓。他們效法耶和華在 以色列 人面前所趕出的外邦人，行一切可憎惡的事。
1KGS|14|25|羅波安 王第五年， 埃及 王 示撒 上來攻打 耶路撒冷 ，
1KGS|14|26|奪了耶和華殿和王宮裏的寶物，盡都帶走，又奪走 所羅門 製造的一切金盾牌。
1KGS|14|27|羅波安 王製造銅盾牌代替那些金盾牌，交給看守王宮宮門的護衛長看管。
1KGS|14|28|每逢王進耶和華的殿，護衛兵就舉起這些盾牌；隨後仍將盾牌送回護衛室。
1KGS|14|29|羅波安 其餘的事，凡他所做的，不都寫在《猶大列王記》上嗎？
1KGS|14|30|羅波安 與 耶羅波安 時常交戰。
1KGS|14|31|羅波安 與他祖先同睡，與他祖先同葬在 大衛城 。他母親名叫 拿瑪 ，是 亞捫 人，他兒子 亞比央 接續他作王。
1KGS|15|1|尼八 的兒子 耶羅波安 王十八年， 亞比央 登基作 猶大 王，
1KGS|15|2|在 耶路撒冷 作王三年。他母親名叫 瑪迦 ，是 押沙龍 的女兒。
1KGS|15|3|亞比央 行他父親從前所犯一切的罪，他的心不像他曾祖父 大衛 以純正的心順服耶和華－他的上帝。
1KGS|15|4|然而耶和華－他的上帝因 大衛 的緣故，仍使大衛在 耶路撒冷 有燈光，立他兒子接續他作王，又堅立 耶路撒冷 。
1KGS|15|5|因為 大衛 除了 赫 人 烏利亞 那件事，都行耶和華眼中看為正的事，一生沒有違背耶和華一切所吩咐的。
1KGS|15|6|羅波安 在世的日子常與 耶羅波安 交戰。
1KGS|15|7|亞比央 其餘的事，凡他所做的，不都寫在《猶大列王記》上嗎？ 亞比央 常與 耶羅波安 交戰。
1KGS|15|8|亞比央 與他祖先同睡，葬在 大衛城 ，他兒子 亞撒 接續他作王。
1KGS|15|9|以色列 王 耶羅波安 第二十年， 亞撒 登基作 猶大 王，
1KGS|15|10|在 耶路撒冷 作王四十一年。他祖母名叫 瑪迦 ，是 押沙龍 的女兒。
1KGS|15|11|亞撒 效法他的高祖父 大衛 行耶和華眼中看為正的事，
1KGS|15|12|從國中除去男的廟妓，又除掉他祖先所造的一切偶像。
1KGS|15|13|他甚至廢了他祖母 瑪迦 太后的位，因 瑪迦 造了可憎的 亞舍拉 。 亞撒 砍下她的偶像，在 汲淪溪 邊燒了，
1KGS|15|14|只是丘壇還沒有廢去。 亞撒 一生向耶和華存純正的心。
1KGS|15|15|亞撒 將他父親所分別為聖與自己所分別為聖的金銀和器皿都奉到耶和華的殿裏。
1KGS|15|16|亞撒 和 以色列 王 巴沙 在世的日子常常交戰。
1KGS|15|17|以色列 王 巴沙 上來攻擊 猶大 ，修築 拉瑪 ，不許人從 猶大 王 亞撒 那裏出入。
1KGS|15|18|於是 亞撒 把耶和華殿和王宮府庫裏所剩下的金銀都交在他臣僕手中，派他們到住在 大馬士革 的 亞蘭 王，就是 希旬 的孫子， 他伯利門 的兒子 便‧哈達 那裏去，說：
1KGS|15|19|「你父曾與我父立約，我與你也要這樣立約。看哪，我把金銀送給你作禮物，請你廢掉你與 以色列 王 巴沙 所立的約，使他從我這裏撤退。」
1KGS|15|20|便‧哈達 聽從了 亞撒 王，就派遣他的軍官去攻打 以色列 的城鎮，攻下了 以雲 、 但 、 亞伯‧伯‧瑪迦 、全 基尼烈 、 拿弗他利 全地。
1KGS|15|21|巴沙 聽見了，就停工不修築 拉瑪 ，仍住在 得撒 。
1KGS|15|22|於是 亞撒 王向 猶大 眾人宣佈，不准任何人推辭，吩咐他們運走 巴沙 修築 拉瑪 所用的石頭和木料。 亞撒 王用它們來修築 便雅憫 的 迦巴 和 米斯巴 。
1KGS|15|23|亞撒 其餘的事，他英勇的事蹟，凡他所做的，以及他所建築的城鎮，不都寫在《猶大列王記》上嗎？只是 亞撒 年老的時候患有腳疾。
1KGS|15|24|亞撒 與他祖先同睡，與他祖先同葬在 大衛城 ，他兒子 約沙法 接續他作王。
1KGS|15|25|猶大 王 亞撒 第二年， 耶羅波安 的兒子 拿答 登基作 以色列 王二年，
1KGS|15|26|拿答 行耶和華眼中看為惡的事，行他父親所行的道，犯他父親使 以色列 陷入罪裏的那罪。
1KGS|15|27|以薩迦 人 亞希雅 的兒子 巴沙 背叛 拿答 ，在 非利士 人的 基比頓 殺了他，那時 拿答 和 以色列 眾人正圍困 基比頓 。
1KGS|15|28|猶大 王 亞撒 第三年， 巴沙 殺了 拿答 ，篡了他的位。
1KGS|15|29|巴沙 一作王就殺了 耶羅波安 全家， 耶羅波安 家凡有氣息的，一個也沒有留下，都殺滅了，正如耶和華藉他僕人 示羅 人 亞希雅 所說的話。
1KGS|15|30|這是因為 耶羅波安 所犯的罪，他使 以色列 陷入罪裏，激怒了耶和華－ 以色列 的上帝。
1KGS|15|31|拿答 其餘的事，凡他所做的，不都寫在《以色列諸王記》上嗎？
1KGS|15|32|亞撒 和 以色列 王 巴沙 在世的日子常常交戰。
1KGS|15|33|猶大 王 亞撒 第三年， 亞希雅 的兒子 巴沙 在 得撒 登基，作全 以色列 的王二十四年。
1KGS|15|34|他行耶和華眼中看為惡的事，行 耶羅波安 所行的道，犯他使 以色列 陷入罪裏的那罪。
1KGS|16|1|耶和華的話臨到 哈拿尼 的兒子 耶戶 ，責備 巴沙 說：
1KGS|16|2|「我既從塵埃中提拔你，立你作我百姓 以色列 的君王，你竟行 耶羅波安 所行的道，使我的百姓 以色列 陷入罪裏，以他們的罪惹我發怒，
1KGS|16|3|看哪，我必除盡 巴沙 和他的家，使你的家像 尼八 的兒子 耶羅波安 的家一樣。
1KGS|16|4|凡屬 巴沙 的人，死在城中的必被狗吃，死在田野的必被空中的鳥吃。」
1KGS|16|5|巴沙 其餘的事，凡他所做的和他英勇的事蹟，不都寫在《以色列諸王記》上嗎？
1KGS|16|6|巴沙 與他祖先同睡，葬在 得撒 ，他兒子 以拉 接續他作王。
1KGS|16|7|耶和華的話臨到 哈拿尼 的兒子 耶戶 先知，責備 巴沙 和他的家，因他行耶和華眼中看為惡的一切事，以他手所做的惹耶和華發怒，像 耶羅波安 的家一樣，又因他殺了 耶羅波安 全家。
1KGS|16|8|猶大 王 亞撒 第二十六年， 巴沙 的兒子 以拉 在 得撒 登基，作 以色列 王二年。
1KGS|16|9|他的大臣 心利 ，就是管理他一半戰車的軍官背叛他。當他在 得撒 ，在王宮的管家 亞雜 家裏喝醉的時候，
1KGS|16|10|心利 進去擊殺他，把他殺死，篡了他的位。這是 猶大 王 亞撒 第二十七年的事。
1KGS|16|11|心利 一坐上王位就殺了 巴沙 全家，連他的親屬和朋友，一個男丁也沒有留下。
1KGS|16|12|心利 滅絕 巴沙 全家，正如耶和華藉 耶戶 先知責備 巴沙 的話。
1KGS|16|13|這是因為 巴沙 和他兒子 以拉 的一切罪，就是他們使 以色列 陷入罪裏的那罪，以虛無的神明 惹耶和華－ 以色列 的上帝發怒。
1KGS|16|14|以拉 其餘的事，凡他所做的，不都寫在《以色列諸王記》上嗎？
1KGS|16|15|猶大 王 亞撒 第二十七年， 心利 在 得撒 作王七日。那時軍兵正安營圍攻 非利士 人的 基比頓 。
1KGS|16|16|軍兵在營中聽說 心利 已經背叛，殺了王， 以色列 眾人當日就在營中立 暗利 元帥作 以色列 王。
1KGS|16|17|暗利 率領 以色列 眾人，從 基比頓 上去，圍困 得撒 。
1KGS|16|18|心利 見城被攻陷，就進了王宮的堡壘，放火焚燒宮殿，自焚而死。
1KGS|16|19|這是因為他犯罪，行耶和華眼中看為惡的事，行 耶羅波安 所行的道，犯他使 以色列 陷入罪裏的那罪。
1KGS|16|20|心利 其餘的事和他背叛的事，不都寫在《以色列諸王記》上嗎？
1KGS|16|21|那時， 以色列 百姓分為兩半：一半隨從 基納 的兒子 提比尼 ，要擁立他作王；另一半隨從 暗利 。
1KGS|16|22|但隨從 暗利 的百姓勝過隨從 基納 兒子 提比尼 的百姓。 提比尼 死了， 暗利 就作了王。
1KGS|16|23|猶大 王 亞撒 第三十一年， 暗利 登基作 以色列 王十二年；他在 得撒 作王六年。
1KGS|16|24|暗利 用二他連得銀子向 撒瑪 買了 撒瑪利亞山 ，在山上建城，按著山的原主 撒瑪 的名，給所建的城起名叫 撒瑪利亞 。
1KGS|16|25|暗利 行耶和華眼中看為惡的事，比他以前所有的王作惡更嚴重。
1KGS|16|26|因為他行了 尼八 的兒子 耶羅波安 所行的道，犯他使 以色列 陷入罪裏的那罪，以虛無的神明惹耶和華－ 以色列 的上帝發怒。
1KGS|16|27|暗利 其餘的事，他所做的和所顯出的英勇事蹟，不都寫在《以色列諸王記》上嗎？
1KGS|16|28|暗利 與他祖先同睡，葬在 撒瑪利亞 ，他兒子 亞哈 接續他作王。
1KGS|16|29|猶大 王 亞撒 第三十八年， 暗利 的兒子 亞哈 登基作 以色列 王。 暗利 的兒子 亞哈 在 撒瑪利亞 作 以色列 王二十二年。
1KGS|16|30|暗利 的兒子 亞哈 行耶和華眼中看為惡的事，比他以前所有的王更嚴重。
1KGS|16|31|他犯了 尼八 的兒子 耶羅波安 所犯的罪，還當作是小事，又娶了 西頓 王 謁巴力 的女兒 耶洗別 為妻，去事奉 巴力 ，敬拜它，
1KGS|16|32|又在 撒瑪利亞 建 巴力廟 ，在廟裏為 巴力 築壇。
1KGS|16|33|亞哈 又造 亞舍拉 ，他所做的惹耶和華－ 以色列 的上帝發怒，比他以前所有的 以色列 王更嚴重。
1KGS|16|34|亞哈 的日子， 伯特利 人 希伊勒 重修 耶利哥 。立根基的時候，他喪了長子 亞比蘭 ；安門的時候，他喪了幼子 西割 ，正如耶和華藉 嫩 的兒子 約書亞 所說的話。
1KGS|17|1|住在 基列 的 提斯比 人 以利亞 對 亞哈 說：「我指著所事奉永生的耶和華－ 以色列 的上帝起誓，這幾年我若不禱告，必不降露水，也不下雨。」
1KGS|17|2|耶和華的話臨到 以利亞 ，說：
1KGS|17|3|「你離開這裏往東去，躲在 約旦河 東邊的 基立溪 旁。
1KGS|17|4|你要喝那溪裏的水，我已吩咐烏鴉在那裏供養你。」
1KGS|17|5|於是 以利亞 去了，他遵照耶和華的話做，去住在 約旦河 東的 基立溪 旁。
1KGS|17|6|烏鴉早上給他叼餅和肉來，晚上也有餅和肉，他又喝溪裏的水。
1KGS|17|7|過了些日子溪水乾了，因為雨沒有下在地上。
1KGS|17|8|耶和華的話臨到他，說：
1KGS|17|9|「你起身到 西頓 的 撒勒法 去，住在那裏，看哪，我已吩咐那裏的一個寡婦供養你。」
1KGS|17|10|以利亞 就起身往 撒勒法 去。他到了城門，看哪，有一個寡婦在那裏撿柴。 以利亞 呼喚她說：「請你用器皿取點水來給我喝。」
1KGS|17|11|她去取水的時候， 以利亞 又呼喚她說：「請你手裏也拿點餅來給我。」
1KGS|17|12|她說：「我指著永生的耶和華－你的上帝起誓，我沒有餅，罈內只有一把麵，瓶裏只有一點油。看哪，我去找兩根柴，帶回家為我和我兒子做餅。我們吃了，就等死吧！」
1KGS|17|13|以利亞 對她說：「不要怕！你去照你所說的做吧！只要先為我做一個小餅，拿來給我，然後為你和你的兒子做餅；
1KGS|17|14|因為耶和華－ 以色列 的上帝如此說：『罈內的麵必不用盡，瓶裏的油必不短缺，直到耶和華使雨降在地上的日子。』」
1KGS|17|15|婦人就照 以利亞 的話去做。她和 以利亞 ，以及她家中的人，吃了許多日子。
1KGS|17|16|罈內的麵果然沒有用盡，瓶裏的油也不短缺，正如耶和華藉 以利亞 所說的話。
1KGS|17|17|這事以後，那婦人，就是那家的女主人，她的兒子病了，病得很重，甚至沒有氣息。
1KGS|17|18|婦人對 以利亞 說：「神人哪，我跟你有甚麼關係，你竟到我這裏來，使上帝記起我的罪，以致我的兒子死了呢？」
1KGS|17|19|以利亞 對她說：「把你兒子交給我。」 以利亞 就從婦人懷中接過孩子來，抱到他所住的頂樓，放在自己的床上。
1KGS|17|20|他求告耶和華說：「耶和華－我的上帝啊，我寄居在這寡婦的家裏，你卻降禍於她，使她的兒子死了嗎？」
1KGS|17|21|以利亞 三次伏在孩子的身上，求告耶和華說：「耶和華－我的上帝啊，求你使這孩子的生命歸回給他吧！」
1KGS|17|22|耶和華聽了 以利亞 的呼求，孩子的生命歸回給他，他就活了。
1KGS|17|23|以利亞 把孩子從樓上抱下來，進了房間交給他母親，說：「看，你的兒子活了！」
1KGS|17|24|婦人對 以利亞 說：「現在我知道你是神人，耶和華藉你口所說的話是真的。」
1KGS|18|1|過了許多日子，到了第三年，耶和華的話臨到 以利亞 ，說：「你去，讓 亞哈 看見你，我要降雨在地面上。」
1KGS|18|2|以利亞 就去，要讓 亞哈 見到他。那時， 撒瑪利亞 的饑荒非常嚴重。
1KGS|18|3|亞哈 召來他的管家 俄巴底 。 俄巴底 非常敬畏耶和華。
1KGS|18|4|耶洗別 殺耶和華先知的時候， 俄巴底 把一百個先知藏了，每五十人藏在一個洞裏，拿餅和水供養他們。
1KGS|18|5|亞哈 對 俄巴底 說：「我們要走遍這地，到一切水泉旁和一切溪邊，或者能找到青草，可以救活馬和騾子，免得喪失一些牲畜。」
1KGS|18|6|於是二人分地巡查， 亞哈 獨自走一路， 俄巴底 獨自走另一路。
1KGS|18|7|俄巴底 在路上時，看哪， 以利亞 遇見他。 俄巴底 認出他來，就臉伏於地，說：「你是我主 以利亞 嗎？」
1KGS|18|8|以利亞 對他說：「我是。你去，告訴你主人說：『看哪， 以利亞 在這裏。』」
1KGS|18|9|俄巴底 說：「僕人犯了甚麼罪，你竟要把我交在 亞哈 手裏，使他殺我呢？
1KGS|18|10|我指著永生的耶和華－你的上帝起誓，無論哪一邦哪一國，我主都派人去找你。若他們說：『不在這裏』，他就叫那邦那國的人起誓說，他們實在找不到你。
1KGS|18|11|現在你說：『你去告訴你主人說，看哪， 以利亞 在這裏』；
1KGS|18|12|恐怕我一離開你，耶和華的靈就把你提到我所不知道的地方去。這樣，我去告訴 亞哈 ，他若找不到你，就必殺我。僕人是自幼敬畏耶和華的。
1KGS|18|13|耶洗別 殺耶和華先知的時候，我把耶和華的一百個先知藏了，每五十人藏在一個洞裏，拿餅和水供養他們，難道沒有人把我做的這事告訴我主嗎？
1KGS|18|14|現在你說：『你去告訴你主人說，看哪， 以利亞 在這裏』，他一定會殺我。」
1KGS|18|15|以利亞 說：「我指著所事奉永生的萬軍之耶和華起誓，我今日要讓 亞哈 見到我。」
1KGS|18|16|於是 俄巴底 去迎見 亞哈 ，告訴他這事。 亞哈 就去見 以利亞 。
1KGS|18|17|亞哈 見了 以利亞 ，就說：「真的是你嗎？你這使 以色列 遭殃的人！」
1KGS|18|18|以利亞 說：「使 以色列 遭殃的不是我，而是你和你的父家，因為你們離棄耶和華的誡命 ，去隨從 巴力 。
1KGS|18|19|現在你要派人去召集 以色列 眾人，以及 耶洗別 所供養的四百五十個 巴力 的先知和四百個 亞舍拉 的先知，叫他們都上 迦密山 到我這裏來。」
1KGS|18|20|亞哈 就派人到 以色列 眾人那裏，召集先知上 迦密山 。
1KGS|18|21|以利亞 近前來對眾百姓說：「你們心持二意要到幾時呢？如果耶和華是上帝，就當順從耶和華；如果是 巴力 ，就當順從 巴力 。」百姓一言不答。
1KGS|18|22|以利亞 對百姓說：「作耶和華先知的只剩下我一個； 巴力 的先知卻有四百五十人。
1KGS|18|23|請給我們兩頭牛犢， 巴力 的先知可以為自己挑選一頭牛犢，切成小塊，放在柴上，不要點火；我也預備一頭牛犢放在柴上，也不點火。
1KGS|18|24|你們求告你們神明的名，我也求告耶和華的名。那應允禱告降火的就是上帝。」眾百姓回答說：「好主意。」
1KGS|18|25|以利亞 對 巴力 的先知說：「因為你們人多，先挑選一頭牛犢，預備好了，求告你們神明的名，卻不要點火。」
1KGS|18|26|他們把所給他們的牛犢預備好了，從早晨到中午，求告 巴力 的名說：「 巴力 啊，求你應允我們！」卻沒有聲音，也沒有回應。他們就在所築的壇四圍蹦跳。
1KGS|18|27|到了正午， 以利亞 嘲笑他們，說：「大聲求告吧！因為它是神明，它或許在默想，或許正忙著 ，或許在路上，或許在睡覺，它該醒過來了。」
1KGS|18|28|他們大聲求告，按著他們的儀式，用刀槍刺割自己，直到渾身流血。
1KGS|18|29|中午過去了，他們狂呼亂叫，直到獻晚祭的時候，卻沒有聲音，沒有回應的，也沒有理睬的。
1KGS|18|30|以利亞 對眾百姓說：「你們到我這裏來。」眾百姓就到他那裏，他把那已經毀壞了的耶和華的壇修好。
1KGS|18|31|以利亞 按照 雅各 子孫支派的數目，取了十二塊石頭；耶和華的話曾臨到 雅各 ，說：「你的名要叫 以色列 。」
1KGS|18|32|以利亞 用這些石頭為耶和華的名築一座壇，在壇的四圍挖溝，可容納二細亞穀種。
1KGS|18|33|他又在壇上擺好了柴，把牛犢切成小塊放在柴上，說：「你們用四個桶盛滿水，倒在燔祭和柴上。」
1KGS|18|34|他又說：「倒第二次。」他們就倒第二次。他又說：「倒第三次。」他們就倒第三次。
1KGS|18|35|水流到壇的四圍，溝裏也滿了水。
1KGS|18|36|到了獻晚祭的時候，先知 以利亞 近前來，說：「耶和華－ 亞伯拉罕 、 以撒 、 以色列 的上帝啊，求你今日使人知道你是 以色列 的上帝，我是你的僕人，我遵照你的話做這一切事。
1KGS|18|37|求你應允我，耶和華啊，應允我，使這百姓知道你－耶和華是上帝，是你叫他們回心轉意的。」
1KGS|18|38|於是，耶和華降下火來，燒盡燔祭、木柴、石頭、塵土，又燒乾了溝裏的水。
1KGS|18|39|眾百姓看見了，就臉伏於地，說：「耶和華是上帝！耶和華是上帝！」
1KGS|18|40|以利亞 對他們說：「拿住 巴力 的先知，不讓任何人逃走！」眾人就拿住他們。 以利亞 帶他們到 基順河 邊，在那裏殺了他們。
1KGS|18|41|以利亞 對 亞哈 說：「你現在可以上去吃喝，因為有暴雨的響聲了。」
1KGS|18|42|亞哈 就上去吃喝。 以利亞 上了 迦密山 頂，屈身在地，把臉伏在兩膝之中。
1KGS|18|43|他對僕人說：「你上去，向海觀看。」僕人就上去觀看，說：「沒有甚麼。」 以利亞 說：「你再去。」如此七次。
1KGS|18|44|第七次，僕人說：「看哪，有一小片雲從海裏上來，好像人的手掌那麼大。」 以利亞 說：「你上去告訴 亞哈 ，當套車下去，免得被雨阻擋。」
1KGS|18|45|霎時間，天因風雲黑暗，降下大雨。 亞哈 就坐上車，往 耶斯列 去了。
1KGS|18|46|耶和華的手按在 以利亞 身上，他就束上腰，奔在 亞哈 前頭，一路到 耶斯列 。
1KGS|19|1|亞哈 把 以利亞 一切所做的和他用刀殺眾先知的事都告訴 耶洗別 。
1KGS|19|2|耶洗別 就派使者到 以利亞 那裏，說：「明日約這時候，我若不使你的性命像那些人的性命一樣，願神明重重懲罰我。」
1KGS|19|3|以利亞 害怕 ，就起來逃命，到了 猶大 的 別是巴 ，把僕人留在那裏。
1KGS|19|4|他自己在曠野走了一日的路程，來到一棵羅騰 樹下，就坐在那裏求死，說：「耶和華啊，現在夠了！求你取我的性命吧，因為我不比我的祖先好。」
1KGS|19|5|他躺在羅騰樹下睡著了。看哪，有一個天使拍他，對他說：「起來吃吧！」
1KGS|19|6|他觀看，看哪，頭旁有燒熱的石頭烤的餅和一壺水，他就吃了喝了，又再躺下。
1KGS|19|7|耶和華的使者回來，第二次拍他，說：「起來吃吧！因為你要走的路很遠。」
1KGS|19|8|他就起來吃了喝了，仗著這飲食的力走了四十晝夜，到了上帝的山，就是 何烈山 。
1KGS|19|9|他在那裏進了一個洞，在洞中過夜。看哪，耶和華的話臨到他，說：「 以利亞 ，你在這裏做甚麼？」
1KGS|19|10|他說：「我為耶和華－萬軍之上帝大發熱心，因為 以色列 人背棄了你的約，毀壞了你的壇，用刀殺了你的先知，只剩下我一人，他們還要追殺我。」
1KGS|19|11|耶和華說：「你出來站在山上，在耶和華面前。」看哪，耶和華從那裏經過。在耶和華面前有烈風大作，山崩石裂，耶和華卻不在風中；風後有地震，耶和華也不在其中；
1KGS|19|12|地震後有火，耶和華也不在火中；火以後，有輕微細小的聲音。
1KGS|19|13|以利亞 聽見，就用外衣蒙臉，出來站在洞口。聽啊，有聲音向他說：「 以利亞 ，你在這裏做甚麼？」
1KGS|19|14|他說：「我為耶和華－萬軍之上帝大發熱心，因為 以色列 人背棄了你的約，毀壞了你的壇，用刀殺了你的先知，只剩下我一人，他們還要追殺我。」
1KGS|19|15|耶和華對他說：「去吧，從原路回去，往 大馬士革 的曠野去。到了那裏，你要膏 哈薛 作 亞蘭 王，
1KGS|19|16|又膏 寧示 的孫子 耶戶 作 以色列 王，並膏 亞伯‧米何拉 人 沙法 的兒子 以利沙 作先知接續你。
1KGS|19|17|將來逃過 哈薛 之刀的，必被 耶戶 所殺；逃過 耶戶 之刀的，必被 以利沙 所殺。
1KGS|19|18|但我在 以色列 中留下七千人，是未曾向 巴力 屈膝，未曾親吻 巴力 的。」
1KGS|19|19|於是， 以利亞 離開那裏走了，遇見 沙法 的兒子 以利沙 ；他正在耕田，在他前頭有十二對牛，自己趕著第十二對。 以利亞 經過他，把自己的外衣搭在他身上。
1KGS|19|20|以利沙 就離開牛，跑到 以利亞 那裏，說：「請你讓我先與父母吻別，然後我就跟隨你。」 以利亞 對他說：「因我對你所做的事，你去吧，然後回來。 」
1KGS|19|21|以利沙 離開他回去，宰了一對牛，用套牛的器具煮肉給百姓吃，隨後就起身跟隨 以利亞 ，服事他。
1KGS|20|1|亞蘭 王 便‧哈達 召集他的全軍，率領三十二個王，帶著馬和戰車，上來圍困 撒瑪利亞 ，要攻打它。
1KGS|20|2|他派使者進城到 以色列 王 亞哈 那裏，對他說：「 便‧哈達 如此說：
1KGS|20|3|『你的金銀都要歸我，你妻妾兒女中最美的也要歸我。』」
1KGS|20|4|以色列 王回答說：「我主我王啊，就照著你的話，我和我所有的都歸你。」
1KGS|20|5|使者又來說：「 便‧哈達 如此說：『我已派人到你那裏，要你把你的金銀、妻妾、兒女都歸我。』
1KGS|20|6|但明日約在這時候，我還要派臣僕到你那裏，搜查你的家和你僕人的家，你眼中一切所喜愛的都由他們的手拿走。」
1KGS|20|7|以色列 王召了國內所有的長老來，說：「你們要知道，看哪，這人是來找麻煩的！他派人到我這裏來，要我的妻妾、兒女和金銀，我並沒有拒絕他。」
1KGS|20|8|所有的長老和眾百姓對王說：「不要聽從他，也不要答應他。」
1KGS|20|9|以色列 王對 便‧哈達 的使者說：「你們告訴我主我王說：『王頭一次派人向僕人所要的一切，僕人都依從，但這事我不能依從。』」使者就去回覆 便‧哈達 。
1KGS|20|10|便‧哈達 又派人到 亞哈 那裏，說：「 撒瑪利亞 的塵土若足夠跟從我的軍兵每人手拿一把，願神明重重懲罰我！」
1KGS|20|11|以色列 王回答說：「你們告訴他說，『剛束上腰帶的，不要像已卸下的那樣誇口。』」
1KGS|20|12|便‧哈達 和諸王正在帳幕裏喝酒，聽見這話，就對他臣僕說：「擺陣吧！」他們就擺陣攻城。
1KGS|20|13|看哪，一個先知靠近 以色列 王 亞哈 ，說：「耶和華如此說：『這一大群人你看見了嗎？看哪，今日我必把他們交在你手裏，你就知道我是耶和華。』」
1KGS|20|14|亞哈 說：「藉著誰呢？」他說：「耶和華如此說：『藉著跟從省長的年輕人。』」 亞哈 說：「誰要開戰呢？」他說：「你！」
1KGS|20|15|於是 亞哈 數點跟從省長的年輕人，共二百三十二名，然後又數點 以色列 的眾軍兵，共七千名。
1KGS|20|16|中午，他們出了城； 便‧哈達 和幫助他的三十二個王正在帳幕裏暢飲。
1KGS|20|17|跟從省長的年輕人先出城。 便‧哈達 派人去，他們回報說：「有人從 撒瑪利亞 出來了。」
1KGS|20|18|他說：「他們若為求和出來，要活捉他們，若為打仗出來，也要活捉他們。」
1KGS|20|19|跟從省長的年輕人，和跟隨他們的軍兵，都出了城，
1KGS|20|20|各人遇見敵人就擊殺。 亞蘭 人逃跑， 以色列 人追趕他們； 亞蘭 王 便‧哈達 騎著馬和騎兵一同逃跑。
1KGS|20|21|以色列 王出城攻擊 馬和戰車，大大擊殺 亞蘭 人。
1KGS|20|22|那先知靠近 以色列 王，對他說：「去吧，你當自強，看清楚，也要知道你所要做的事，因為再過一年， 亞蘭 王會上來攻擊你。」
1KGS|20|23|亞蘭 王的臣僕對他說：「他們的神是山神，所以他們勝過我們。但在平原與他們打仗，我們一定勝過他們。
1KGS|20|24|王當做這樣的事，把諸王革去，派軍官代替他們，
1KGS|20|25|又照著王喪失軍兵的數目，再招募一支軍隊，馬補馬，車補車。然後在平原與他們打仗，我們一定勝過他們。」王就聽臣僕的話，照樣去做。
1KGS|20|26|過了一年， 便‧哈達 果然召集 亞蘭 人上 亞弗 去，要與 以色列 人打仗。
1KGS|20|27|以色列 人也召集軍兵，預備食物，去迎戰 亞蘭 人。 以色列 人對著他們安營，好像兩小群的山羊； 亞蘭 人卻佈滿了地面。
1KGS|20|28|有神人靠近，對 以色列 王說：「耶和華如此說：『 亞蘭 人既說我－耶和華是山神，不是平原之神，我必將這一大群人全都交在你手中，你們就知道我是耶和華。』」
1KGS|20|29|以色列 人與 亞蘭 人相對安營七日，到第七日兩軍開戰。那一日 以色列 人殺了 亞蘭 的十萬步兵，
1KGS|20|30|其餘的都逃向 亞弗 ，到了城裏，城牆倒塌，壓死了剩下的二萬七千人。 便‧哈達 也逃入城內，藏在嚴密的內室裏。
1KGS|20|31|他的臣僕對他說：「看哪，我們聽說 以色列 家的王都是仁慈的王；讓我們腰束麻布，頭套繩索，出去到 以色列 王那裏，也許他會存留王的性命。」
1KGS|20|32|於是他們腰束麻布，頭套繩索，來到 以色列 王那裏，說：「王的僕人 便‧哈達 說：『求王饒我一命。』」 亞哈 說：「他還活著嗎？他是我的兄弟。」
1KGS|20|33|這些人正在探測吉凶，就立即抓住他的話說：「 便‧哈達 是王的兄弟！」王說：「你們去請他來。」 便‧哈達 出來到王那裏，王就請他上車。
1KGS|20|34|便‧哈達 對王說：「我父從你父那裏所奪的城鎮，我必歸還給你。你可以在 大馬士革 為你自己設立街市，像我父在 撒瑪利亞 所設立的一樣。」 亞哈 說：「我照此立約，放你回去。」王就與他立約，放了他。
1KGS|20|35|有一個人是先知的門徒，遵照耶和華的話對他同伴說：「你打我吧！」那人不肯打他。
1KGS|20|36|他就對那人說：「你既不聽從耶和華的話，看哪，你一離開我，必有獅子咬死你。」那人一離開他，果然遇見獅子，把他咬死了。
1KGS|20|37|先知的門徒又遇見一個人，對他說：「你打我吧！」那人就打他，把他打傷。
1KGS|20|38|那先知就去了，用頭巾蒙眼，改了裝，在路旁等候王。
1KGS|20|39|王從那裏經過，他向王呼叫說：「僕人出戰的時候，看哪，有人轉過來，帶了一個人到我這裏來，說：『你要看守這人，若他真的失蹤了，你的性命必代替他的性命，否則，你就要交出一他連得銀子來。』
1KGS|20|40|僕人正在到處忙碌的時候，那人就不見了。」 以色列 王對他說：「你自己決定了，就必照樣判你。」
1KGS|20|41|他急忙除掉蒙眼的頭巾， 以色列 王就認出他是一個先知。
1KGS|20|42|他對王說：「耶和華如此說：『因你把我決定要消滅的人從你手中放走，所以你的命必代替他的命，你的百姓必代替他的百姓。』」
1KGS|20|43|於是 以色列 王生氣，憂悶地回 撒瑪利亞 ，到自己的宮去了。
1KGS|21|1|這些事以後，又有一事。 耶斯列 人 拿伯 在 耶斯列 有一個葡萄園，靠近 撒瑪利亞 ， 亞哈 王的宮。
1KGS|21|2|亞哈 對 拿伯 說：「把你的葡萄園給我作菜園，因為它靠近我的宮，我就把更好的葡萄園換給你。你若要銀子，我就按著價錢給你。」
1KGS|21|3|拿伯 對 亞哈 說：「耶和華不准我把我祖先留下的產業給你。」
1KGS|21|4|亞哈 因 耶斯列 人 拿伯 說「我不把我祖先留下的產業給你」，就生氣，憂悶地回宮，躺在床上，臉轉向內，也不吃飯。
1KGS|21|5|耶洗別 王后來對他說：「你為甚麼心裏這樣生氣，不吃飯呢？」
1KGS|21|6|他對王后說：「我向 耶斯列 人 拿伯 說：『把你的葡萄園按價錢賣給我，或是你願意，我可以把別的葡萄園換給你。』他卻說：『我不把我的葡萄園給你。』」
1KGS|21|7|耶洗別 王后對王說：「你現在是不是治理 以色列 國呢？只管起來，心裏暢暢快快地吃飯，我會把 耶斯列 人 拿伯 的葡萄園給你。」
1KGS|21|8|於是王后以 亞哈 的名義寫信，蓋上王的印，把信送給那些與 拿伯 同城居住的長老和貴族。
1KGS|21|9|她在信上寫著說：「你們當宣告禁食，叫 拿伯 坐在百姓的高位上，
1KGS|21|10|又叫兩個無賴坐在 拿伯 對面，作證告他說：『你詛咒了上帝和王。』然後把他拉出去用石頭打死。」
1KGS|21|11|那些與 拿伯 同城居住的長老和貴族，照 耶洗別 送給他們的信去做。正如她送的信上所寫，
1KGS|21|12|他們宣告禁食，叫 拿伯 坐在百姓的高位上。
1KGS|21|13|有兩個無賴來，坐在 拿伯 對面。無賴當著百姓作證告他說：「 拿伯 詛咒上帝和王了！」眾人就把他拉到城外，用石頭打他，他就死了。
1KGS|21|14|於是他們派人到 耶洗別 那裏，說：「 拿伯 被石頭打死了。」
1KGS|21|15|耶洗別 聽見 拿伯 被石頭打死，就對 亞哈 說：「你起來，去取得 耶斯列 人 拿伯 不肯出價賣給你的葡萄園吧！因為 拿伯 不在了，他已經死了。」
1KGS|21|16|亞哈 聽見 拿伯 死了，就起來，下去要取得 耶斯列 人 拿伯 的葡萄園。
1KGS|21|17|耶和華的話臨到 提斯比 人 以利亞 ，說：
1KGS|21|18|「你起來，去見在 撒瑪利亞 的 以色列 王 亞哈 。看哪，他下去要取得 拿伯 的葡萄園，他正在那園裏。
1KGS|21|19|你要對他說：『耶和華如此說：你殺了人，還要取得他的產業嗎？』又要對他說：『耶和華如此說：狗在何處舔 拿伯 的血，狗也必在何處舔你的血。』」
1KGS|21|20|亞哈 對 以利亞 說：「我的仇敵啊，你找到我了嗎？」他說：「我找到你了。因為你出賣自己，行了耶和華眼中看為惡的事。
1KGS|21|21|耶和華說：『看哪，我必使災禍臨到你，把你除滅。 以色列 中凡屬 亞哈 的男丁，無論是奴役的、自由的，我都要剪除。
1KGS|21|22|我必使你的家像 尼八 的兒子 耶羅波安 的家，又像 亞希雅 的兒子 巴沙 的家，因為你惹我發怒，又使 以色列 陷入罪裏。』
1KGS|21|23|論到 耶洗別 ，耶和華說：『狗必在 耶斯列 的城郭 吃 耶洗別 。
1KGS|21|24|凡屬 亞哈 的人，死在城中的必被狗吃，死在田野的必被空中的鳥吃。』」
1KGS|21|25|（只是從來沒有像 亞哈 的，因他受 耶洗別 王后的唆使，出賣自己，行了耶和華眼中看為惡的事。
1KGS|21|26|他行了最可憎的事，隨從偶像，正如耶和華在 以色列 人面前趕出的 亞摩利 人所行的一切。）
1KGS|21|27|亞哈 聽見這些話，就撕裂衣服，禁食，貼身穿著麻布，也睡在麻布上，沮喪地走來走去。
1KGS|21|28|耶和華的話臨到 提斯比 人 以利亞 ，說：
1KGS|21|29|「 亞哈 在我面前這樣謙卑，你看見了嗎？因為他在我面前謙卑，所以在他的日子，我不降這禍；到他兒子的時候，我必降這禍於他的家。」
1KGS|22|1|亞蘭 和 以色列 之間連續三年沒有戰爭。
1KGS|22|2|到了第三年， 猶大 王 約沙法 下去見 以色列 王。
1KGS|22|3|以色列 王對臣僕說：「你們不知道 基列 的 拉末 是屬我們的嗎？我們豈可不採取行動，把它從 亞蘭 王手裏奪回來呢？」
1KGS|22|4|亞哈 問 約沙法 說：「你肯同我去攻打 基列 的 拉末 嗎？」 約沙法 對 以色列 王說：「你我不分彼此，我的軍隊就是你的軍隊，我的馬就是你的馬。」
1KGS|22|5|約沙法 對 以色列 王說：「請你先求問耶和華的話。」
1KGS|22|6|於是 以色列 王召集先知，約有四百人，問他們說：「我可以上去攻打 基列 的 拉末 嗎？還是不要上去呢？」他們說：「可以上去，因為主必將那城交在王的手裏。」
1KGS|22|7|約沙法 說：「這裏還有沒有耶和華的先知，我們好求問他呢？」
1KGS|22|8|以色列 王對 約沙法 說：「還有一個人，是 音拉 的兒子 米該雅 ，我們可以託他求問耶和華。只是我真的很恨他，因為他對我說預言，從不說吉言，總是說凶信。」 約沙法 說：「請王不要這麼說。」
1KGS|22|9|以色列 王召了一個官員來，說：「你快去，把 音拉 的兒子 米該雅 召來。」
1KGS|22|10|以色列 王和 猶大 王 約沙法 在 撒瑪利亞 城門前的禾場，各穿朝服，坐在寶座上，所有的先知都在他們面前說預言。
1KGS|22|11|基拿拿 的兒子 西底家 造了鐵角，說：「耶和華如此說：『你要用這些角牴觸 亞蘭 人，直到將他們滅盡。』」
1KGS|22|12|所有的先知也都這樣預言說：「可以上 基列 的 拉末 去，必然得勝，因為耶和華必將那城交在王的手中。」
1KGS|22|13|那去召 米該雅 的使者對他說：「看哪，眾先知都異口同聲向王說吉言，你也跟他們說一樣的話，說吉言吧！」
1KGS|22|14|米該雅 說：「我指著永生的耶和華起誓，耶和華向我說甚麼，我就說甚麼。」
1KGS|22|15|米該雅 來到王那裏，王問他：「 米該雅 ，我們可以上去攻打 基列 的 拉末 嗎？還是不要上去呢？」他對王說：「你可以上去，必然得勝，耶和華必將那城交在王的手中。」
1KGS|22|16|王對他說：「我要你發誓多少次，你才會奉耶和華的名向我說實話呢？」
1KGS|22|17|米該雅 說：「我看見 以色列 眾人散佈在山上，如同沒有牧人的羊群一般。耶和華說：『這些人沒有主人，他們可以平安地各自回家去。』」
1KGS|22|18|以色列 王對 約沙法 說：「我豈沒有告訴你，這人對我說預言，從不說吉言，只說凶信嗎？」
1KGS|22|19|米該雅 說：「因此你要聽耶和華的話！我看見耶和華坐在寶座上，天上的萬軍侍立在他左右。
1KGS|22|20|耶和華說：『誰去引誘 亞哈 上 基列 的 拉末 去陣亡呢？』這個這樣說，那個那樣說。
1KGS|22|21|隨後有一個靈出來，站在耶和華面前，說：『我去引誘他。』
1KGS|22|22|耶和華問他：『用甚麼方法呢？』他說：『我要出去，在他眾先知的口中成為謊言的靈。』耶和華說：『這樣，你去引誘他，必能成功。你出去，照樣做吧！』
1KGS|22|23|現在，看哪，耶和華使謊言的靈入了你所有的這些先知的口，並且耶和華已經宣告要降禍於你。」
1KGS|22|24|基拿拿 的兒子 西底家 前來，打 米該雅 一巴掌，說：「耶和華的靈從哪裏離開我向你說話呢？」
1KGS|22|25|米該雅 說：「看哪，你進入嚴密的內室躲藏的那日，就必看見。」
1KGS|22|26|以色列 王說：「把 米該雅 帶走，交回給 亞們 市長和 約阿施 王子。
1KGS|22|27|你們要說：『王如此說，把這個人關在監獄裏，使他受苦，吃不飽喝不足，直等到我平安回來。』」
1KGS|22|28|米該雅 說：「你若真的能平安回來，那就是耶和華沒有藉我說這話了。」他又說：「眾百姓啊，你們都要聽！」
1KGS|22|29|以色列 王和 猶大 王 約沙法 上 基列 的 拉末 去。
1KGS|22|30|以色列 王對 約沙法 說：「我要改裝上陣，你可以仍穿王袍。」 以色列 王就改裝上陣去了。
1KGS|22|31|亞蘭 王吩咐他的三十二個戰車長說：「你們不要與他們的大將或小兵交戰，只要單單攻擊 以色列 王。」
1KGS|22|32|那些戰車長看見 約沙法 就說：「這一定是 以色列 王！」他們轉過去與他交戰， 約沙法 就呼喊起來。
1KGS|22|33|戰車長見他不是 以色列 王，就轉身不追他了。
1KGS|22|34|有一人開弓，並不知情，箭恰巧射入 以色列 王鎧甲的縫裏。王對駕車的說：「我受重傷了，你掉過車來，載我離開戰場！」
1KGS|22|35|那日，戰況越來越猛，有人扶著王站在戰車上，面對 亞蘭 人。到了傍晚，王就死了，血從傷處流入車底。
1KGS|22|36|約在日落的時候，有喊聲傳遍軍中，說：「大家各歸本城，各歸本地吧！」
1KGS|22|37|王死了，人把他送到 撒瑪利亞 ，葬在 撒瑪利亞 。
1KGS|22|38|他們在 撒瑪利亞 的水池旁洗他的車，有狗來舔他的血，有妓女在那裏洗澡，正如耶和華所說的話。
1KGS|22|39|亞哈 其餘的事，凡他所做的、他所修造的象牙宮和所建築的一切城鎮，不都寫在《以色列諸王記》上嗎？
1KGS|22|40|亞哈 與他祖先同睡，他兒子 亞哈謝 接續他作王。
1KGS|22|41|以色列 王 亞哈 第四年， 亞撒 的兒子 約沙法 登基作 猶大 王。
1KGS|22|42|約沙法 登基的時候年三十五歲，在 耶路撒冷 作王二十五年。他母親名叫 阿蘇巴 ，是 示利希 的女兒。
1KGS|22|43|約沙法 效法他父親 亞撒 所行的道，不偏離左右，行耶和華眼中看為正的事。只是丘壇還沒有廢去，百姓仍在那裏獻祭燒香。
1KGS|22|44|約沙法 與 以色列 王和平相處。
1KGS|22|45|約沙法 其餘的事和他所行的英勇事蹟，以及他的戰役，不都寫在《猶大列王記》上嗎？
1KGS|22|46|約沙法 把他父親 亞撒 的日子所剩下男的廟妓都從國中除去了。
1KGS|22|47|那時 以東 沒有立王，由總督治理。
1KGS|22|48|約沙法 造了 他施 船隻，要往 俄斐 去，把金子運來，卻沒有啟航，因為船在 以旬‧迦別 毀壞了。
1KGS|22|49|亞哈 的兒子 亞哈謝 對 約沙法 說：「讓我的僕人和你的僕人坐船同去吧！」 約沙法 卻不肯。
1KGS|22|50|約沙法 與他祖先同睡，與他祖先同葬在 大衛城 ，他兒子 約蘭 接續他作王。
1KGS|22|51|猶大 王 約沙法 第十七年， 亞哈 的兒子 亞哈謝 在 撒瑪利亞 登基作 以色列 王；他作 以色列 王二年。
1KGS|22|52|他行耶和華眼中看為惡的事，行他父母的道，又行 尼八 的兒子 耶羅波安 的道，使 以色列 陷入罪裏。
1KGS|22|53|他事奉 巴力 ，敬拜它，惹耶和華－ 以色列 的上帝發怒，正如他父親一切所行的。
2KGS|1|1|亞哈 死後， 摩押 背叛 以色列 。
2KGS|1|2|亞哈謝 在 撒瑪利亞 ，一日從樓上的欄杆跌下來，就病了。於是他派使者，對他們說：「你們去問 以革倫 的神明 巴力‧西卜 ，我這病是否能痊癒。」
2KGS|1|3|但耶和華的使者對 提斯比 人 以利亞 說：「你起來，上去迎見 撒瑪利亞 王的使者，對他們說：『你們去問 以革倫 的神明 巴力‧西卜 ，是因為 以色列 中沒有上帝嗎？』
2KGS|1|4|所以耶和華如此說：『你必不能下你所上的床，因為你一定會死！』」 以利亞 就去了。
2KGS|1|5|使者回到王那裏，王對他們說：「你們為甚麼回來了呢？」
2KGS|1|6|他們對王說：「有一個人上來迎見我們，對我們說：『去，回到差你們來的王那裏，對他說：耶和華如此說，你派人去問 以革倫 的神明 巴力‧西卜 ，是因為 以色列 中沒有上帝嗎？所以你必不能下所上的床，你一定會死。』」
2KGS|1|7|王對他們說：「上來迎見你們，告訴你們這些話的人是甚麼樣子呢？」
2KGS|1|8|他們對王說：「這人身穿毛衣 ，腰束皮帶。」王說：「他一定是 提斯比 人 以利亞 。」
2KGS|1|9|於是，王派了一個五十夫長，帶領五十人到 以利亞 那裏。他上來，看哪， 以利亞 正坐在山頂上。五十夫長對他說：「神人哪，王吩咐你下來！」
2KGS|1|10|以利亞 回答五十夫長說：「我若是神人，願火從天上降下來，吞滅你和你的五十個人！」於是有火從天上降下來，吞滅五十夫長和他的五十個人。
2KGS|1|11|王又派另一個五十夫長，帶領五十人到 以利亞 那裏。五十夫長對他說：「神人哪，王這樣吩咐，快快下來！」
2KGS|1|12|以利亞 回答他們說：「我若是神人，願火從天上降下來，吞滅你和你的五十個人！」於是上帝的火 從天上降下來，吞滅五十夫長和他的五十個人。
2KGS|1|13|王第三次又派一個五十夫長，帶領五十人去。第三個五十夫長上去，雙膝跪在 以利亞 面前，哀求他說：「神人哪，願我的性命和你這五十個僕人的性命在你眼中看為寶貴！
2KGS|1|14|看哪，已經有火從天上降下來，吞滅前兩次來的五十夫長和他們的五十個人，現在願我的性命在你眼中看為寶貴！」
2KGS|1|15|耶和華的使者對 以利亞 說：「你跟他下去，不要怕他！」 以利亞 就起來，跟他下到王那裏去。
2KGS|1|16|他對王說：「耶和華如此說：『你派人去問 以革倫 的神明 巴力‧西卜 ，是因為 以色列 中沒有上帝可以讓你求問他的話嗎？所以你必不能下所上的床，你一定會死！』」
2KGS|1|17|亞哈謝 死了，正如耶和華藉 以利亞 所說的話。 猶大 王 約沙法 的兒子 約蘭 第二年， 亞哈謝 的兄弟 約蘭 接續他作王，因 亞哈謝 沒有兒子。
2KGS|1|18|亞哈謝 其餘所做的事，不都寫在《以色列諸王記》上嗎？
2KGS|2|1|耶和華要用旋風接 以利亞 升天的時候， 以利亞 與 以利沙 從 吉甲 往前行。
2KGS|2|2|以利亞 對 以利沙 說：「耶和華差遣我往 伯特利 去，你可以留在這裏。」 以利沙 說：「我指著永生的耶和華，又指著你的性命起誓，我必不離開你。」於是二人下到 伯特利 。
2KGS|2|3|在 伯特利 的先知的門徒出來，到 以利沙 那裏，對他說：「耶和華今日要接你的師父離開你 ，你知不知道？」他說：「我知道，你們不要作聲。」
2KGS|2|4|以利亞 對 以利沙 說：「耶和華差遣我往 耶利哥 去，你可以留在這裏。」 以利沙 說：「我指著永生的耶和華，又指著你的性命起誓，我必不離開你。」於是二人到了 耶利哥 。
2KGS|2|5|在 耶利哥 的先知的門徒來靠近 以利沙 ，對他說：「耶和華今日要接你的師父離開你，你知不知道？」他說：「我知道，你們不要作聲。」
2KGS|2|6|以利亞 對 以利沙 說：「耶和華差遣我往 約旦河 去，你可以留在這裏。」 以利沙 說：「我指著永生的耶和華，又指著你的性命起誓，我必不離開你。」於是二人一同往前行。
2KGS|2|7|有五十個先知的門徒同去，遠遠地站在他們對面；他們二人在 約旦河 邊站住。
2KGS|2|8|以利亞 捲起自己的外衣，用來打水，水就左右分開，二人走乾地過去。
2KGS|2|9|過去之後， 以利亞 對 以利沙 說：「我未被接去離開你以前，你要我為你做甚麼，只管求。」 以利沙 說：「願感動你的靈雙倍感動我。」
2KGS|2|10|以利亞 說：「你求的是一件難事。我被接去離開你的時候，你若看見我，就必得著；若不然，就得不著了。」
2KGS|2|11|他們邊走邊說話的時候，看哪，有火馬和火焰車出現，把二人隔開， 以利亞 就乘旋風升天去了。
2KGS|2|12|以利沙 看見，就呼叫說：「我父啊！我父啊！ 以色列 的戰車騎兵啊！」 以利沙 不再看見他的時候，就把自己的衣服撕為兩片。
2KGS|2|13|他拾起 以利亞 身上掉下來的外衣，回去站在 約旦河 邊。
2KGS|2|14|他用 以利亞 身上掉下來的外衣打水，說：「耶和華－ 以利亞 的上帝在哪裏呢？」打水之後，水也左右分開， 以利沙 就過去了。
2KGS|2|15|在 耶利哥 的先知的門徒從對面看見他，說：「感動 以利亞 的靈臨到 以利沙 身上了。」他們就來迎接他，俯伏於地，向他下拜，
2KGS|2|16|對他說：「看哪，僕人這裏有五十個壯士，請你讓他們去尋找你師父，或者耶和華的靈將他提起來，投在某山某谷。」 以利沙 說：「你們不必派人去。」
2KGS|2|17|他們再三催促，直到他不好意思，就說：「你們派人去吧！」他們就派了五十個人去，尋找了三天，也沒有找著他。
2KGS|2|18|以利沙 仍然留在 耶利哥 ，他們回到他那裏，他對他們說：「我不是告訴你們不必去嗎？」
2KGS|2|19|耶利哥城 的人對 以利沙 說：「看哪，這城的地勢美好，正如我主所看見的，只是水質惡劣，地也沒有生產。」
2KGS|2|20|以利沙 說：「你們拿一個新的瓶子來，裏面裝鹽。」他們就拿給他。
2KGS|2|21|他出去到了水源，把鹽倒在那裏，說：「耶和華如此說：『我治好了這水，從那裏不會再有死亡和不生產的事了。』」
2KGS|2|22|於是那水治好了，直到今日，正如 以利沙 所說的話。
2KGS|2|23|以利沙 從那裏上 伯特利 去。正上路的時候，有些孩童從城裏出來，譏笑他，對他說：「禿頭的，上去吧！禿頭的，上去吧！」
2KGS|2|24|他轉過身來瞪著他們，奉耶和華的名詛咒他們。於是有兩隻母熊從林中出來，撕裂他們當中的四十二個孩童。
2KGS|2|25|以利沙 從 伯特利 上 迦密山 ，又從那裏回到 撒瑪利亞 。
2KGS|3|1|猶大 王 約沙法 第十八年， 亞哈 的兒子 約蘭 在 撒瑪利亞 登基，作 以色列 王十二年。
2KGS|3|2|他行耶和華眼中看為惡的事，但不致像他父母所行的，因為他除掉他父所造 巴力 的柱像。
2KGS|3|3|然而，他依戀 尼八 的兒子 耶羅波安 使 以色列 陷入罪裏的那罪，總不離開。
2KGS|3|4|摩押 王 米沙 牧養許多羊，曾向 以色列 王進貢十萬羔羊和十萬公綿羊的毛。
2KGS|3|5|亞哈 死後， 摩押 王背叛 以色列 王。
2KGS|3|6|那時 約蘭 王出 撒瑪利亞 ，數點 以色列 眾人。
2KGS|3|7|他向前行，派人到 猶大 王 約沙法 那裏，說：「 摩押 王背叛我，你肯同我去攻打 摩押 嗎？」 約沙法 說：「我肯上去，你我不分彼此，我的軍隊就是你的軍隊，我的馬就是你的馬。」
2KGS|3|8|然後 約沙法 說：「我們從哪條路上去呢？」 約蘭 說：「從 以東 曠野的路上去。」
2KGS|3|9|於是， 以色列 王和 猶大 王，以及 以東 王，都一同去。他們繞行了七日的路程，軍隊和所帶的牲畜都沒有水喝。
2KGS|3|10|以色列 王說：「哀哉！耶和華召集我們這三王，是要交在 摩押 人的手裏。」
2KGS|3|11|約沙法 說：「這裏不是有耶和華的先知嗎？我們可以託他求問耶和華。」 以色列 王的一個大臣回答說：「這裏有 沙法 的兒子 以利沙 ，就是從前服事 以利亞 的 。」
2KGS|3|12|約沙法 說：「他必有耶和華的話。」於是 以色列 王、 約沙法 和 以東 王都下去見他。
2KGS|3|13|以利沙 對 以色列 王說：「我跟你有甚麼關係呢？去問你父親的先知和你母親的先知吧！」 以色列 王對他說：「不，因為耶和華召集我們這三王，是要交在 摩押 人的手裏。」
2KGS|3|14|以利沙 說：「我指著所事奉永生的萬軍之耶和華起誓，我若不看 猶大 王 約沙法 的情面，必不理你，不睬你。
2KGS|3|15|現在你們給我找一個彈琴的人來。」彈琴的人彈奏的時候，耶和華的手就按在 以利沙 身上。
2KGS|3|16|他就說：「耶和華如此說：『你們要在這谷中到處挖溝。』
2KGS|3|17|因為耶和華如此說：『你們雖不見風，也不見雨，這谷卻必滿了水，使你們和你們的牛羊牲畜都有水喝。』
2KGS|3|18|在耶和華眼中這還算是小事，他也必將 摩押 人交在你們手中。
2KGS|3|19|你們必攻破一切堡壘和美好的城鎮，砍伐各種好樹，塞住一切水泉，用石頭毀壞一切良田。」
2KGS|3|20|到了早晨，約在獻祭的時候，看哪，有水從 以東 而來，遍地就滿了水。
2KGS|3|21|摩押 眾人聽見這三王上來要與他們打仗，凡能束上腰帶的，無論老少，都被召集站在邊界上。
2KGS|3|22|摩押 人清早起來，日光照在水上，他們看見對面水紅如血，
2KGS|3|23|就說：「這是血啊！必是三王互相擊殺，全都滅亡了。 摩押 人哪，我們現在去搶奪財物吧！」
2KGS|3|24|摩押 人到了 以色列 營， 以色列 人起來攻打他們，他們就在 以色列 人面前逃跑。 以色列 人追殺 摩押 人，直殺入 摩押 境內 。
2KGS|3|25|他們拆毀 摩押 的城鎮，各人拋石頭填滿一切良田，塞住一切水泉，砍伐各種好樹，只剩下 吉珥‧哈列設 的石牆，但甩石的兵仍然包圍攻打那城。
2KGS|3|26|摩押 王見戰事激烈，對他不利，就率領七百個拿刀的兵，想突圍逃到 以東 王那裏，卻沒有成功。
2KGS|3|27|於是他在城牆上，把那應當接續他作王的長子獻為燔祭。 有極大的憤怒臨到 以色列 ，於是三王離開 摩押 王，各自回本地去了。
2KGS|4|1|有個先知門徒的妻子哀求 以利沙 說：「你的僕人，我丈夫死了，他敬畏耶和華是你所知道的。現在有債主來，要帶走我的兩個孩子給他作奴隸。」
2KGS|4|2|以利沙 對她說：「我可以為你做甚麼呢？告訴我，你家裏有甚麼？」她說：「婢女家中除了一瓶油之外，甚麼也沒有。」
2KGS|4|3|以利沙 說：「你到外面去向所有的鄰舍借器皿，要空的器皿，不要少借。
2KGS|4|4|然後你回家，關上門，你和你兒子在裏面把油倒在所有的器皿裏，倒滿了就放在一邊。」
2KGS|4|5|於是婦人離開 以利沙 去了。她關上門，把自己和兒子關在家裏。他們把器皿拿給她，她就倒油。
2KGS|4|6|器皿都滿了，她對兒子說：「再給我拿器皿來。」兒子對她說：「沒有器皿了。」油就止住了。
2KGS|4|7|婦人去告訴神人，神人說：「你去賣了油還債，你和你兩個兒子可以靠著所剩的過活。」
2KGS|4|8|一日， 以利沙 經過 書念 ，在那裏有一個富有的婦人強留他吃飯。此後， 以利沙 每次經過就轉到那裏去吃飯。
2KGS|4|9|婦人對丈夫說：「看哪，我知道那常從我們這裏經過的是神聖的神人。
2KGS|4|10|我們可以為他蓋一間有牆的小閣樓，裏面安放床榻、桌子、椅子、燈臺。每當他來到我們這裏，就可以住在那裏。」
2KGS|4|11|一日， 以利沙 來到那裏，轉進那閣樓，躺臥在那裏。
2KGS|4|12|以利沙 吩咐僕人 基哈西 說：「你叫這 書念 婦人來。」他把婦人叫了來，婦人就站在 以利沙 面前。
2KGS|4|13|以利沙 吩咐僕人說：「你對她說：『看哪，你為我們費了許多心思，我可以為你做甚麼呢？我可以為你向王或元帥求甚麼呢？』」她說：「我已住在自己百姓之中。」
2KGS|4|14|以利沙 說：「究竟可以為她做甚麼呢？」 基哈西 說：「她真的沒有兒子，她丈夫也老了。」
2KGS|4|15|以利沙 說：「叫她回來。」於是他叫了她來，她就站在門口。
2KGS|4|16|以利沙 說：「明年這時候 ，你必抱一個兒子。」她說：「神人，我主啊，不要這樣欺哄婢女。」
2KGS|4|17|婦人果然懷孕，到了明年那時候，生了一個兒子，正如 以利沙 向她所說的。
2KGS|4|18|孩子長大，一日出去到他父親和收割的人那裏。
2KGS|4|19|他對父親說：「我的頭啊，我的頭啊！」他父親對僕人說：「把他抱到他母親那裏。」
2KGS|4|20|僕人抱去，交給他母親。孩子坐在母親的膝上，到中午就死了。
2KGS|4|21|他母親上去，把他放在神人的床上，關了門出來，
2KGS|4|22|呼叫她丈夫說：「你叫一個僕人給我牽一匹驢來，我要趕去見神人，然後回來。」
2KGS|4|23|丈夫說：「今日不是初一，也不是安息日，你為何要到他那裏去呢？」婦人說：「平安無事。」
2KGS|4|24|於是她備上驢，對僕人說：「走，趕緊走，除非我吩咐你，不要為了我而慢下來。」
2KGS|4|25|婦人往 迦密山 去，到了神人那裏。 神人遠遠看見她，對僕人 基哈西 說：「看哪， 書念 的婦人來了！
2KGS|4|26|現在你跑去迎接她，對她說，你平安嗎？你丈夫平安嗎？孩子平安嗎？」她說：「平安。」
2KGS|4|27|婦人上了山，到神人那裏，就抱住神人的腳。 基哈西 前來要推開她，神人說：「由她吧！因為她心裏愁苦。但耶和華向我隱瞞這事，沒有告訴我。」
2KGS|4|28|婦人說：「我何嘗向我主求過兒子呢？我豈不是說過，不要欺哄我嗎？」
2KGS|4|29|以利沙 吩咐 基哈西 說：「你束上腰，手拿我的杖前去。若遇見人，不要向他問安，人若向你問安，也不要回答。要把我的杖放在孩子臉上。」
2KGS|4|30|孩子的母親說：「我指著永生的耶和華，又指著你的性命起誓，我必不離開你。」於是 以利沙 起身，隨著她去了。
2KGS|4|31|基哈西 在他們以先去了，把杖放在孩子臉上，卻沒有聲音，也沒有動靜。 基哈西 回去，迎見 以利沙 ，告訴他說：「孩子還沒有醒過來。」
2KGS|4|32|以利沙 進了屋子，看哪，孩子死了，放在自己的床上。
2KGS|4|33|他進去，關上門，只有他們兩個人，他就向耶和華祈禱。
2KGS|4|34|他上去伏在孩子身上，口對口，眼對眼，手對手。他伏在孩子身上，孩子的身體就漸漸暖和了。
2KGS|4|35|然後他下來，在屋裏來回走了一趟，又上去伏在孩子身上。孩子打了七個噴嚏，眼睛就睜開了。
2KGS|4|36|以利沙 叫 基哈西 說：「你叫這 書念 婦人來。」於是他叫了她來。婦人來到 以利沙 那裏， 以利沙 說：「把你兒子抱起來。」
2KGS|4|37|婦人就進來，在 以利沙 腳前俯伏於地，向他下拜，然後抱起她兒子出去了。
2KGS|4|38|以利沙 回到 吉甲 ，那地正有饑荒。先知的門徒坐在他面前，他吩咐僕人說：「你把大鍋放在火上，給先知的門徒熬湯。」
2KGS|4|39|有一個人去到田野摘菜，發現一棵野瓜藤，就摘了滿滿一兜的野瓜回來，切了放進熬湯的鍋中，並不知道那是甚麼。
2KGS|4|40|他們把湯倒出來給大家吃。他們吃湯裏東西的時候，喊叫說：「神人哪，鍋子裏的東西會死人！」所以他們不能吃了。
2KGS|4|41|以利沙 說：「拿點麵來。」他把麵撒在鍋中，說：「倒出來，給大家吃吧！」鍋中就沒有毒了。
2KGS|4|42|有一個人從 巴力‧沙利沙 來，帶著初熟果子的食物、二十個大麥做的餅和新麥穗，裝在袋子裏送給神人。神人說：「把這些給大家吃。」
2KGS|4|43|僕人說：「這些豈可擺在一百人面前呢？」 以利沙 說：「你只管給大家吃吧！因為耶和華如此說，他們必吃了，還有剩下的。」
2KGS|4|44|僕人就擺在他們面前，他們吃了，還有剩下，正如耶和華所說的。
2KGS|5|1|亞蘭 王的元帥 乃縵 在他主人面前是一個偉大的人，得王的喜悅，因為耶和華曾藉他使 亞蘭 人得勝。他雖然是大能的勇士，卻染上了痲瘋 。
2KGS|5|2|亞蘭 人成群出征的時候，從 以色列 地擄了一個小女孩，她就服事 乃縵 的妻子。
2KGS|5|3|她對女主人說：「我希望主人去見 撒瑪利亞 的先知，他必能治好主人的痲瘋。」
2KGS|5|4|乃縵 去告訴他主人說，從 以色列 地來的女孩如此如此說。
2KGS|5|5|亞蘭 王說：「你可以去，我也會送信給 以色列 王。」於是 乃縵 手裏帶十他連得銀子、六千舍客勒金子和十套衣裳去了。
2KGS|5|6|他帶著這信給 以色列 王，說：「現在你接到這信，看哪，我派臣僕 乃縵 到你這裏來，你要治好他的痲瘋。」
2KGS|5|7|以色列 王讀了信就撕裂衣服，說：「我豈是上帝，能使人死使人活呢？這人竟派人來，叫我治好一個人的痲瘋。你們要知道，看，這人是找機會來跟我吵架的。」
2KGS|5|8|神人 以利沙 聽見 以色列 王撕裂衣服，就派人到王那裏，說：「你為甚麼撕裂衣服呢？讓那人到我這裏來，他會知道 以色列 中有先知。」
2KGS|5|9|於是 乃縵 帶著車馬到了 以利沙 的家，站在門前。
2KGS|5|10|以利沙 派一個使者，對 乃縵 說：「去，在 約旦河 中沐浴七次，你的肉就必復原，你會得潔淨。」
2KGS|5|11|乃縵 卻發怒走了。他說：「看哪，我以為他必定會出來，到我這裏，站著求告耶和華－他上帝的名，在患處上搖手，治好這痲瘋。
2KGS|5|12|大馬士革 的 亞瑪拿河 和 法珥法河 豈不比 以色列 的一切水更好嗎？我難道不可以在那裏沐浴而得潔淨嗎？」於是他生氣，轉身走了。
2KGS|5|13|他的僕人近前來，對他說：「我父啊，先知若吩咐你做一件大事，你豈不做嗎？何況是吩咐你去沐浴，得潔淨呢？」
2KGS|5|14|於是 乃縵 下去，照著神人的話，在 約旦河 裏浸了七次。他的肉復原，好像小孩的肉，他就潔淨了。
2KGS|5|15|乃縵 帶著所有跟隨他的人，回到神人那裏，站在他面前，說：「看哪，我知道，除了 以色列 ，全地沒有上帝。現在請你收下僕人的禮物。」
2KGS|5|16|以利沙 說：「我指著所事奉永生的耶和華起誓，我必不接受。」 乃縵 再三請他收下，他卻不肯。
2KGS|5|17|乃縵 說：「你若不肯，請把兩匹騾子能馱的土賜給僕人，僕人必不再把燔祭或祭物獻給別神，只獻給耶和華。
2KGS|5|18|惟有一件事，願耶和華饒恕你僕人：我主人進 臨門 廟在那裏叩拜的時候，他總是扶著我的手，所以我也在 臨門 廟叩拜。我在 臨門 廟叩拜的這事，願耶和華饒恕你僕人。」
2KGS|5|19|以利沙 對他說：「你平安地回去吧！」 乃縵 離開他去了。走了一小段路，
2KGS|5|20|神人 以利沙 的僕人 基哈西 說：「看哪，我主人不願從這 亞蘭 人 乃縵 手裏接受他帶來的禮物，我指著永生的耶和華起誓，我必跑去追上他，向他拿些東西。」
2KGS|5|21|於是 基哈西 去追 乃縵 。 乃縵 看見有人追來，就下車迎著他，說：「都平安嗎？」
2KGS|5|22|他說：「都平安！我主人派我來說：『看哪，現在有兩個年輕人，是先知的門徒，從 以法蓮 山區來到我這裏，請你給他們一他連得銀子，兩套衣裳。』」
2KGS|5|23|乃縵 說：「好啊，請收下二他連得。」他再三請求，就把二他連得銀子裝在兩個袋子裏，連同兩套衣裳交給兩個僕人；他們就在 基哈西 前頭抬著走。
2KGS|5|24|到了山岡， 基哈西 從他們手中接過來，放在屋裏，打發這些人走了。
2KGS|5|25|基哈西 進去，站在主人面前。 以利沙 對他說：「 基哈西 ，你從哪裏來？」他說：「僕人哪裏也沒去。」
2KGS|5|26|以利沙 對他說：「那人下車轉過來迎著你的時候，我的心豈沒有去呢？這豈是接受銀子，接受衣裳、橄欖園、葡萄園、牛羊、僕婢的時候呢？
2KGS|5|27|因此， 乃縵 的痲瘋必緊隨你和你的後裔，直到永遠。」 基哈西 從 以利沙 面前出去，就長了痲瘋，像雪一樣。
2KGS|6|1|先知的門徒對 以利沙 說：「看哪，我們在你面前居住的地方，那裏對我們太窄小了。
2KGS|6|2|讓我們往 約旦河 去，各人從那裏取一根木料，在那裏為自己建造居住的地方。」他說：「你們去吧！」
2KGS|6|3|有一人說：「請你與僕人同去。」他說：「我可以去。」
2KGS|6|4|於是 以利沙 與他們同去。到了 約旦河 ，他們砍伐樹木。
2KGS|6|5|有一人砍樹的時候，斧子的頭掉在水裏，他就喊著說：「不好了！我主啊，斧子是借來的。」
2KGS|6|6|神人說：「掉在哪裏了？」他把那地方指給 以利沙 看。 以利沙 砍了一塊木頭，拋在水裏，就使斧子的頭浮上來了。
2KGS|6|7|以利沙 說：「拿起來吧！」那人就伸手拿起來了。
2KGS|6|8|亞蘭 王與 以色列 作戰，他和臣僕商議說：「我要在某處某處安營 。」
2KGS|6|9|神人派人到 以色列 王那裏，說：「你要小心，不要從某處經過，因為 亞蘭 人下到那裏去了。」
2KGS|6|10|以色列 王派人到神人告訴他的地方去。神人警告他，他就在那裏有所防備，不止一兩次。
2KGS|6|11|亞蘭 王因這事心裏氣憤，召了臣僕來，對他們說：「我們當中有誰幫助 以色列 王，你們不告訴我嗎？」
2KGS|6|12|有一個臣僕說：「不，我主，我王！只有 以色列 中的先知 以利沙 ，把王在臥房所說的話告訴 以色列 王。」
2KGS|6|13|王說：「你們去查看他在哪裏，我好派人去捉拿他。」有人告訴王說：「看哪，他在 多坍 。」
2KGS|6|14|王就派遣車馬和大軍往那裏去，夜間他們到了，圍困那城。
2KGS|6|15|神人的僕人清早起來出去，看哪，車馬軍兵圍困了城。僕人對神人說：「不好了！我主啊，我們該怎麼辦呢？」
2KGS|6|16|神人說：「不要懼怕！因與我們同在的比與他們同在的更多。」
2KGS|6|17|以利沙 禱告說：「耶和華啊，求你開他的眼目，使他能看見。」耶和華開了這年輕人的眼目，他就看見了，看哪，滿山有火馬和火焰車圍繞 以利沙 。
2KGS|6|18|亞蘭 人下到 以利沙 那裏， 以利沙 向耶和華禱告說：「求你擊打這國，使他們眼目失明。」耶和華就照 以利沙 的話，擊打他們，使他們眼目失明。
2KGS|6|19|以利沙 對他們說：「這不是那條路，也不是那座城。你們跟我走，我必領你們到你們要尋找的人那裏。」於是他領他們到了 撒瑪利亞 。
2KGS|6|20|他們進了 撒瑪利亞 ， 以利沙 說：「耶和華啊，求你開這些人的眼目，使他們能看見。」耶和華開了他們的眼目，他們就看見了，看哪，是在 撒瑪利亞城 中。
2KGS|6|21|以色列 王看見他們，就對 以利沙 說：「我父啊，我真的可以擊殺他們嗎？」
2KGS|6|22|他說：「不可擊殺！這些人豈是你用刀用弓擄來給你擊殺的呢？當在他們面前擺設飲食給他們吃喝，讓他們回到他們主人那裏。」
2KGS|6|23|王為他們預備了盛大的宴席。他們吃喝完了，王就送他們回到他們主人那裏。此後， 亞蘭 的軍隊不再侵犯 以色列 地了。
2KGS|6|24|此後， 亞蘭 王 便‧哈達 召集他的全軍，上來圍困 撒瑪利亞 。
2KGS|6|25|看哪，被圍困的時候， 撒瑪利亞 有大饑荒，甚至一個驢頭值八十舍客勒，四分之一卡布 的鴿子糞值五舍客勒。
2KGS|6|26|一日， 以色列 王在城牆上經過，有一個婦人向他呼叫說：「我主，我王啊！求你幫助。」
2KGS|6|27|王說：「耶和華不幫助你，我從哪裏幫助你呢？是從禾場，或從壓酒池嗎？」
2KGS|6|28|王對婦人說：「你有甚麼事？」她說：「這婦人對我說：『把你的兒子交出來，我們今日可以吃他，明日可以吃我的兒子。』
2KGS|6|29|我們就煮了我的兒子吃了。次日我對她說：『要把你的兒子交出來，我們可以吃。』她卻把她的兒子藏起來。」
2KGS|6|30|王聽見婦人的話，就撕裂衣服；那時，王在城牆上經過，百姓看見了，看哪，王貼身穿著麻布。
2KGS|6|31|王說：「我今日若容許 沙法 的兒子 以利沙 的頭還留在他身上，願上帝重重懲罰我！」
2KGS|6|32|那時， 以利沙 正坐在家中，有長老與他同坐。王派一個人先去，使者還沒有到， 以利沙 對長老說：「你們看，這兇手之子派人來斬我的頭。你們注意，當使者來到，你們就關上門，把他關在門外。在他後頭不就是他主人的腳步聲嗎？」
2KGS|6|33|正與他們說話的時候，看哪，使者 下到他那裏，說：「看哪，這災禍是從耶和華來的，我何必再仰望耶和華呢？」
2KGS|7|1|以利沙 說：「你們要聽耶和華的話，耶和華如此說：明日約這時候，在 撒瑪利亞 城門口，一細亞細麵只賣一舍客勒，二細亞大麥也賣一舍客勒。」
2KGS|7|2|有一個攙扶王的軍官回答神人說：「看哪，即使耶和華打開天上的窗戶，也不可能有這事。」 以利沙 說：「看哪，你必親眼看見，在那裏卻吃不到甚麼。」
2KGS|7|3|在城門口有四個長痲瘋的人，他們彼此說：「我們為何坐在這裏等死呢？
2KGS|7|4|我們若說要進城去，城裏有饑荒，我們必死在那裏。若我們在這裏坐著不動，也必死。現在，來吧，我們去向 亞蘭 人的軍隊投降。若他們饒我們的命，我們就活著；若殺我們，我們就死吧！」
2KGS|7|5|黃昏的時候，他們起來往 亞蘭 人的軍營去；到了營邊，看哪，沒有一人在那裏。
2KGS|7|6|因為主使 亞蘭 人的軍隊聽見戰車戰馬的聲音，大軍的聲音，他們就彼此說：「看哪，這必是 以色列 王雇用 赫 人諸王和 埃及 諸王來攻擊我們。」
2KGS|7|7|所以，在黃昏的時候他們起來逃跑，撇下帳棚、馬、驢，把軍營留在原處，只顧逃命。
2KGS|7|8|那些長痲瘋的人到了營邊，進了一座帳棚，吃了喝了，從當中拿走金銀和衣服，收藏起來。他們又回來，進了另一座帳棚，從當中拿走財物去收藏。
2KGS|7|9|那時，他們彼此說：「我們所做的不對了！這一天是有好消息的日子，我們竟不作聲！若等到天亮，我們就有罪了。現在，來，我們去向王室報信吧！」
2KGS|7|10|他們就去叫守城門的人，告訴他們說：「我們到了 亞蘭 人的軍營，看哪，沒有一人在那裏，也無人聲，只有拴著的馬和驢，帳棚都留在原處。」
2KGS|7|11|守城門的人就呼叫，他們向城內的王室報信。
2KGS|7|12|王夜間起來，對臣僕說：「我告訴你們 亞蘭 人向我們做的事。他們知道我們飢餓，所以離營，埋伏在田野，說：『 以色列 人出城的時候，我們活捉他們，我們就可以進到城裏去。』」
2KGS|7|13|王的一個臣僕回答說：「不如叫人從城裏剩下的馬中取五匹，看哪，這些馬像 以色列 大眾一樣 ，快要滅亡了；我們派人去窺探吧！」
2KGS|7|14|於是他們取了兩輛車和馬，王派人去跟蹤 亞蘭 人的軍隊，說：「你們去窺探吧。」
2KGS|7|15|他們去跟蹤 亞蘭 人，直到 約旦河 。看哪，整條路上都是 亞蘭 人匆忙逃跑時所丟棄的衣服和器具，使者就回來向王報告。
2KGS|7|16|百姓就出去，擄掠 亞蘭 人的軍營。於是一細亞細麵只賣一舍客勒，二細亞大麥也賣一舍客勒，正如耶和華所說的。
2KGS|7|17|王派攙扶他的那軍官在城門指揮，百姓在城門把他踩死了，正如神人在王下到他那裏的時候所說的。
2KGS|7|18|神人曾對王說：「明日約這時候，在 撒瑪利亞 城門口，二細亞大麥只賣一舍客勒，一細亞細麵也賣一舍客勒。」
2KGS|7|19|那軍官回答神人說：「看哪，即使耶和華打開天上的窗戶，也不可能有這事。」神人說：「看哪，你必親眼看見，在那裏卻吃不到甚麼。」
2KGS|7|20|這話果然應驗在他身上，因為百姓在城門把他踩死了。
2KGS|8|1|以利沙 曾對他救活的孩子的母親說：「你和你的全家要起身，往你可住的地方去住，因為耶和華已令饑荒降在這地七年。」
2KGS|8|2|婦人就起身，照神人的話去做，帶著全家往 非利士 人的地去，寄居了七年。
2KGS|8|3|過了七年，那婦人從 非利士 人的地回來，就出去為自己的房屋田地哀求王。
2KGS|8|4|那時王正與神人的僕人 基哈西 談話，說：「你把 以利沙 所做的一切大事告訴我。」
2KGS|8|5|基哈西 告訴王 以利沙 如何使死人復活，看哪， 以利沙 所救活的孩子的母親正為自己的房屋田地來哀求王。 基哈西 說：「我主我王，這就是那婦人，這是她的兒子，就是 以利沙 所救活的。」
2KGS|8|6|王問那婦人，她就把事情告訴王。於是王為她派一個官員，說：「凡屬這婦人的都還給她，自從她離開本地直到今日，她田地的出產也都還給她。」
2KGS|8|7|以利沙 來到 大馬士革 ， 亞蘭 王 便‧哈達 正患病。有人告訴王說：「神人來到這裏了。」
2KGS|8|8|王就吩咐 哈薛 說：「你帶著禮物去見神人，託他求問耶和華，我這病能不能好？」
2KGS|8|9|於是 哈薛 用四十匹駱駝，馱著 大馬士革 的各樣美物為禮物，去迎見 以利沙 。 哈薛 到了那裏，站在他面前，說：「你兒子 亞蘭 王 便‧哈達 派我到你這裏，問說：『我這病會不會好？』」
2KGS|8|10|以利沙 對 哈薛 說：「你回去告訴他說：『你一定會好。』但耶和華指示我，他必定會死。」
2KGS|8|11|神人定睛看著 哈薛 ，直到他感到羞愧。神人就哭了。
2KGS|8|12|哈薛 說：「我主為甚麼哭？」他說：「因為我知道你必虐待 以色列 人，用火焚燒他們的堡壘，用刀殺死他們的壯丁，摔死他們的嬰孩，剖開他們的孕婦。」
2KGS|8|13|哈薛 說：「僕人算甚麼，不過是一條狗，怎麼能行這大事呢？」 以利沙 說：「耶和華指示我，你必作 亞蘭 王。」
2KGS|8|14|哈薛 離開 以利沙 ，回到他主人那裏。主人對他說：「 以利沙 對你說了甚麼？」他說：「他告訴我你必能好。」
2KGS|8|15|次日， 哈薛 拿被子浸在水中，蒙住王的臉，王就死了。於是 哈薛 篡了他的位。
2KGS|8|16|亞哈 的兒子 以色列 王 約蘭 第五年－ 約沙法 曾作 猶大 王 － 猶大 王 約沙法 的兒子 約蘭 登基作了 猶大 王。
2KGS|8|17|約蘭 登基的時候年三十二歲，在 耶路撒冷 作王八年。
2KGS|8|18|他行 以色列 諸王的道，正如 亞哈 家所行的，因他娶了 亞哈 的女兒為妻，行耶和華眼中看為惡的事。
2KGS|8|19|耶和華卻因他僕人 大衛 的緣故，不肯滅絕 猶大 ，要照他所應許的，永遠賜燈光給 大衛 和他的子孫。
2KGS|8|20|約蘭 在位期間， 以東 背叛，自己立王治理他們，脫離 猶大 的權勢。
2KGS|8|21|約蘭 率領他所有的戰車過到 撒益 去。他夜間起來，攻打圍困他的 以東 人和戰車長； 猶大 軍兵逃跑，各回自己的帳棚去了；
2KGS|8|22|這樣， 以東 背叛，脫離 猶大 的管轄，直到今日。那時 立拿 也背叛了。
2KGS|8|23|約蘭 其餘的事，凡他所做的，不都寫在《猶大列王記》上嗎？
2KGS|8|24|約蘭 與他祖先同睡，與他祖先同葬在 大衛城 ，他兒子 亞哈謝 接續他作王。
2KGS|8|25|亞哈 的兒子 以色列 王 約蘭 第十二年， 猶大 王 約蘭 的兒子 亞哈謝 登基。
2KGS|8|26|他登基的時候年二十二歲，在 耶路撒冷 作王一年。他母親名叫 亞她利雅 ，是 以色列 王 暗利 的孫女。
2KGS|8|27|亞哈謝 行 亞哈 家的道，行耶和華眼中看為惡的事，與 亞哈 家一樣，因為他是 亞哈 家的女婿。
2KGS|8|28|他與 亞哈 的兒子 約蘭 同往 基列 的 拉末 去，與 亞蘭 王 哈薛 交戰。 亞蘭 人打傷了 約蘭 ，
2KGS|8|29|約蘭 王回到 耶斯列 ，醫治在 拉末 與 亞蘭 王 哈薛 打仗時，被 亞蘭 人擊打所受的傷。 約蘭 的兒子 猶大 王 亞哈謝 因為 亞哈 的兒子 約蘭 病了，就下到 耶斯列 看望他。
2KGS|9|1|以利沙 先知叫了一個先知的門徒來，吩咐他：「你束上腰，手拿這瓶膏油往 基列 的 拉末 去。
2KGS|9|2|你到了那裏，要在那裏尋找 寧示 的孫子， 約沙法 的兒子 耶戶 。你去，使他從弟兄中起來，帶他進最裏面的內室，
2KGS|9|3|把瓶裏的膏油倒在他頭上，說：『耶和華如此說：我膏你作 以色列 王。』然後你就開門逃跑，不要等候。」
2KGS|9|4|於是那青年，那年輕的先知往 基列 的 拉末 去了。
2KGS|9|5|他到了那裏，看哪，眾軍官都坐著，就說：「長官，我有話對你說。」 耶戶 說：「你要對我們哪一個說呢？」他說：「長官，我要對你說。」
2KGS|9|6|耶戶 就起來，進了內室，那青年把膏油倒在他頭上，對他說：「耶和華－ 以色列 的上帝如此說：『我膏你作耶和華百姓 以色列 的王。
2KGS|9|7|你要擊殺你主人 亞哈 的全家，我好在 耶洗別 身上，為我僕人眾先知和耶和華所有僕人的血伸冤。
2KGS|9|8|亞哈 全家都必滅亡，凡屬 亞哈 的男丁，無論是奴役的、自由的，我必從 以色列 中剪除。
2KGS|9|9|我必使 亞哈 的家像 尼八 兒子 耶羅波安 的家，又像 亞希雅 兒子 巴沙 的家。
2KGS|9|10|至於 耶洗別 ，狗必在 耶斯列 田裏吃她，無人埋葬。』」於是那青年就開門逃跑了。
2KGS|9|11|耶戶 出來，回到他主人的臣僕那裏，有一人問他說：「平安嗎？這瘋狂的人為甚麼到你這裏來呢？」他對他們說：「你們認得那人，也知道他在胡說。」
2KGS|9|12|他們說：「說謊！告訴我們吧。」他說：「他如此如此對我說：『耶和華如此說：我膏你作 以色列 的王。』」
2KGS|9|13|他們各人就急忙把自己的衣服鋪在臺階的上層，在 耶戶 的下面；他們吹角，說：「 耶戶 作王了！」
2KGS|9|14|這樣， 寧示 的孫子， 約沙法 的兒子 耶戶 背叛了 約蘭 。先前 約蘭 和 以色列 眾人因為 亞蘭 王 哈薛 的緣故，把守 基列 的 拉末 。
2KGS|9|15|後來 約蘭 王回到 耶斯列 ，醫治他與 亞蘭 王 哈薛 打仗時，被 亞蘭 人擊打所受的傷。 耶戶 說：「若你們有這樣的意思，就不要讓人溜出城，到 耶斯列 去報信。」
2KGS|9|16|於是 耶戶 駕戰車往 耶斯列 去，因為 約蘭 臥病在那裏。 猶大 王 亞哈謝 已經下去看望他。
2KGS|9|17|有一個守望的人站在 耶斯列 的城樓上，看見 耶戶 帶著一隊人來，就說：「我看見一隊人。」 約蘭 說：「派一個騎兵去迎接他們，問說：『平安嗎？』」
2KGS|9|18|騎兵就去迎接 耶戶 ，說：「王如此說：『平安嗎？』」耶戶說：「平安不平安跟你有甚麼關係呢？轉身跟在我後面吧！」守望的人說：「使者到了他們那裏，卻不回來。」
2KGS|9|19|王又派第二個騎兵去。這人到了他們那裏，說：「王如此說：『平安嗎？』」 耶戶 說：「平安不平安跟你有甚麼關係呢？轉身跟在我後面吧！」
2KGS|9|20|守望的人又說：「他到了他們那裏，也不回來。車駕得很兇猛，好像 寧示 的孫子 耶戶 在駕車。」
2KGS|9|21|約蘭 吩咐說：「套車！」人就給他套車。 以色列 王 約蘭 和 猶大 王 亞哈謝 各坐自己的車出去迎接 耶戶 ，在 耶斯列 人 拿伯 的田那裏遇見他。
2KGS|9|22|約蘭 見 耶戶 就說：「 耶戶 ，平安嗎？」 耶戶 說：「你母親 耶洗別 的淫行邪術這樣多，怎麼能平安呢？」
2KGS|9|23|約蘭 用手轉過車來逃跑，對 亞哈謝 說：「 亞哈謝 啊，反了！」
2KGS|9|24|耶戶 全力拉弓，射中 約蘭 兩臂中間，箭從心窩穿出， 約蘭 就仆倒在車上。
2KGS|9|25|耶戶 對他的軍官 畢甲 說：「把他拋在 耶斯列 人 拿伯 的田裏。你當記得，你我一同駕車跟隨他父親 亞哈 的時候，耶和華對 亞哈 說了預言，
2KGS|9|26|耶和華說：『我昨日看見 拿伯 的血和他眾子的血，我發誓我必在這塊田上報應你。』這是耶和華說的。現在你要照著耶和華的話，把他拋在這田裏。」
2KGS|9|27|猶大 王 亞哈謝 看見了，就沿著 伯．哈干 的路逃跑。 耶戶 追趕他，說：「把這人也擊殺在車上，在靠近 以伯蓮 的 姑珥 坡上 。」他逃到 米吉多 ，就死在那裏。
2KGS|9|28|他的臣僕用車把他的屍體運回 耶路撒冷 ，與他祖先同葬在 大衛城 ，他自己的墳墓裏。
2KGS|9|29|亞哈 的兒子 約蘭 第十一年， 亞哈謝 登基作了 猶大 王。
2KGS|9|30|耶戶 到了 耶斯列 。 耶洗別 聽見了，就畫眼影、梳頭，從窗戶往外觀看。
2KGS|9|31|耶戶 進了城門， 耶洗別 說：「殺主人的 心利 啊，平安嗎？」
2KGS|9|32|耶戶 向窗戶抬頭，說：「有誰順從我？誰？」有兩三個太監向外看他。
2KGS|9|33|耶戶 說：「把她拋下來！」他們就把她拋下來。她的血濺在牆上和馬上， 耶戶 踐踏在她身上。
2KGS|9|34|耶戶 進去，吃了喝了，說：「你們去處理這被詛咒的婦人，埋了她，因為她是王的女兒。」
2KGS|9|35|他們去了，要埋葬她，卻只找到她的頭骨和腳，以及手掌。
2KGS|9|36|他們回來報告 耶戶 ， 耶戶 說：「這正應驗耶和華藉他僕人 提斯比 人 以利亞 所說的話，說：『在 耶斯列 田裏，狗必吃 耶洗別 的肉，
2KGS|9|37|耶洗別 的屍體必在 耶斯列 田裏的地面上如同糞土，甚至沒有人可說：這是 耶洗別 。』」
2KGS|10|1|亞哈 有七十個兒子在 撒瑪利亞 。 耶戶 寫信送到 撒瑪利亞 ，給 耶斯列 的領袖和長老 ，以及教養 亞哈 眾兒子的人，說：
2KGS|10|2|「你們主人的眾兒子既然在你們那裏，你們又有戰車、馬匹、兵器、堅固城，現在你們接了這信，
2KGS|10|3|可以在你們主人的眾兒子中選一個賢能正直的，使他坐他父親的王位，你們也可以為你們主人的家作戰。」
2KGS|10|4|他們卻非常懼怕，說：「看哪，兩個王在他面前尚且站立不住，我們怎能站立得住呢？」
2KGS|10|5|王宮總管、市長和長老，並教養眾兒子的人，派人到 耶戶 那裏，說：「我們是你的僕人，凡你所吩咐的，我們都必遵行。我們不立誰作王，你看怎樣好就怎樣做吧。」
2KGS|10|6|耶戶 寫第二封信給他們，說：「你們若歸順我，聽從我的話，明日這時候，要帶著你們主人眾兒子的首級，來到 耶斯列 我這裏。」那時王的兒子七十人都住在城中教養他們的那些尊貴人家裏。
2KGS|10|7|信一到他們那裏，他們就把王的七十個兒子殺了，將首級裝在筐裏，送到 耶斯列 ， 耶戶 那裏。
2KGS|10|8|有使者來告訴 耶戶 說：「他們把王眾兒子的首級送來了。」 耶戶 說：「把首級分成兩堆，放在城門口，直到早晨。」
2KGS|10|9|次日早晨， 耶戶 出來，站著對眾百姓說：「你們都是公義的！看哪，我背叛了我的主人，把他殺了，但這所有的人又是誰殺的呢？
2KGS|10|10|由此可知，耶和華指著 亞哈 家所說的話一句也沒有落空，因為耶和華實現了他藉他僕人 以利亞 所說的話。」
2KGS|10|11|凡 亞哈 家在 耶斯列 所剩下的，他的大臣、密友、祭司， 耶戶 全都殺了，沒有留下一個倖存者。
2KGS|10|12|耶戶 起身往 撒瑪利亞 去。路途中，在牧人聚集的 伯．艾克特 ，
2KGS|10|13|耶戶 遇見 猶大 王 亞哈謝 的兄弟，說：「你們是誰？」他們說：「我們是 亞哈謝 的兄弟，現在下去要向王和太后的眾兒子問安。」
2KGS|10|14|耶戶 說：「活捉他們！」人就活捉了他們，把他們殺在 伯．艾克特 的坑邊，共四十二人，一個也沒有留下。
2KGS|10|15|耶戶 從那裏往前行，遇見 利甲 的兒子 約拿達 來迎接他， 耶戶 向他問安，對他說：「你的心 ，像我的心待你的心那樣正直嗎？」 約拿達 說：「是。」 耶戶 說：「若是這樣，請你伸出手來。」他伸出手， 耶戶 就拉他上車。
2KGS|10|16|耶戶 說：「你和我同去，看我為耶和華怎樣熱心。」於是他們請他坐在車上。
2KGS|10|17|到了 撒瑪利亞 ， 耶戶 把 亞哈 家在 撒瑪利亞 剩下的人全都殺了，直到滅盡，正如耶和華對 以利亞 所說的話。
2KGS|10|18|耶戶 召集眾百姓，對他們說：「 亞哈 事奉 巴力 還不夠熱心， 耶戶 更要熱心。
2KGS|10|19|現在你們召集 巴力 的眾先知和所有拜 巴力 的人，以及 巴力 的眾祭司，都到我這裏來，一個也不可缺少，因為我要給 巴力 獻大祭；凡不來的必不得活。」 耶戶 行詭詐，為要消滅拜 巴力 的人。
2KGS|10|20|耶戶 說：「要為 巴力 召集嚴肅會！」於是他們宣告了。
2KGS|10|21|耶戶 派人走遍 以色列 ；凡拜 巴力 的人都來齊了，沒有留下一個不來的。他們進了 巴力 廟， 巴力 廟中前後都擠滿了人。
2KGS|10|22|耶戶 對掌管服裝的人說：「拿出袍子來，給所有拜 巴力 的人穿。」他就拿出禮服來給了他們。
2KGS|10|23|耶戶 和 利甲 的兒子 約拿達 進了 巴力 廟，對拜 巴力 的人說：「你們要搜查察看，不可以有耶和華的僕人在你們這裏，只可以有拜 巴力 的人。」
2KGS|10|24|他們進去，獻上祭物和燔祭． 耶戶 先安排八十人在廟外，說：「我把這些人交在你們手中，誰放走其中一人，誰就要以命償命！」
2KGS|10|25|耶戶 獻完了燔祭，就對護衛兵和眾軍官說：「進去殺他們，不要讓一人逃脫！」護衛兵和軍官用刀殺了他們，將屍體拋出去，然後進入 巴力 廟的堡壘，
2KGS|10|26|將 巴力 廟中的柱像都 拿出來焚燒。
2KGS|10|27|他們毀壞 巴力 的柱像，拆毀了 巴力 廟當廁所，直到今日。
2KGS|10|28|這樣， 耶戶 在 以色列 中消滅了 巴力 。
2KGS|10|29|只是 耶戶 不離開 尼八 的兒子 耶羅波安 使 以色列 人陷入罪裏的那罪，就是拜 伯特利 和 但 的金牛犢。
2KGS|10|30|耶和華對 耶戶 說：「因你辦好我眼中看為正的事，照我的心意待 亞哈 家，你的子孫必接續你坐 以色列 的王位，直到第四代。」
2KGS|10|31|只是 耶戶 不盡心遵守耶和華－ 以色列 上帝的律法，不離開 耶羅波安 使 以色列 人陷入罪裏的那罪。
2KGS|10|32|在那些日子，耶和華開始削弱 以色列 。 哈薛 在 以色列 各邊界攻擊他們，
2KGS|10|33|就是 約旦河 東 基列 全地，從靠近 亞嫩谷 邊的 亞羅珥 起，包括 基列 和 巴珊 ，就是 迦得 人、 呂便 人、 瑪拿西 人的地。
2KGS|10|34|耶戶 其餘的事，凡他所做的和他英勇的事蹟，不都寫在《以色列諸王記》上嗎？
2KGS|10|35|耶戶 與他祖先同睡，葬在 撒瑪利亞 ，他兒子 約哈斯 接續他作王。
2KGS|10|36|耶戶 在 撒瑪利亞 作 以色列 王二十八年。
2KGS|11|1|亞哈謝 的母親 亞她利雅 見她兒子死了，就起來剿滅王室所有的後裔。
2KGS|11|2|但 約蘭 王的女兒， 亞哈謝 的妹妹 約示巴 ，將 亞哈謝 的兒子 約阿施 從被殺的王子中偷出來，把他和他的奶媽藏在臥房裏，躲避了 亞她利雅 ，沒有被殺。
2KGS|11|3|亞她利雅 治理這地的時候， 約阿施 和他的奶媽在耶和華的殿裏藏了六年。
2KGS|11|4|第七年， 耶何耶大 派人叫 迦利 人和護衛兵的眾百夫長來，領他們進耶和華的殿，與他們立約，使他們在耶和華殿裏起誓，又把王的兒子指給他們看，
2KGS|11|5|吩咐他們說：「你們要這樣做：你們當中在安息日值班的，三分之一要把守王宮，
2KGS|11|6|三分之一要在 蘇珥門 ，三分之一要在護衛兵院的後門；你們要這樣輪流把守王宮。
2KGS|11|7|你們安息日所有不值班的兩隊人員要在耶和華的殿裏護衛王；
2KGS|11|8|各人手拿兵器，四圍保護王。凡擅自闖入你們行列的，要被處死。王出入的時候，你們當跟隨他。」
2KGS|11|9|眾百夫長就照著 耶何耶大 祭司一切所吩咐的去做，各帶自己的人，無論安息日值班或不值班的，都到 耶何耶大 祭司那裏。
2KGS|11|10|祭司就把耶和華殿裏所藏 大衛 王的槍和盾牌交給百夫長。
2KGS|11|11|護衛兵手中各拿兵器，在祭壇和殿那裏，從殿南到殿北，站在王的四圍。
2KGS|11|12|耶何耶大 領 約阿施 出來，給他戴上冠冕，把律法書交給他，膏他作王；眾人都鼓掌說：「願王萬歲！」
2KGS|11|13|亞她利雅 聽見護衛兵和百姓的聲音，就進耶和華的殿，到百姓那裏。
2KGS|11|14|她觀看，看哪，王照儀式站在柱旁，百夫長和號手在王旁邊，國中的眾百姓歡樂吹號。 亞她利雅 就撕裂衣服，喊著說：「反了！反了！」
2KGS|11|15|耶何耶大 祭司吩咐管軍兵的百夫長，對他們說：「把她從行列之間趕出去，凡跟隨她的必用刀殺死！」因為祭司說：「不可在耶和華殿裏殺她。」
2KGS|11|16|他們就下手拿住她；她進入通往王宮的 馬門 ，就在那裏被殺。
2KGS|11|17|耶何耶大 使王和百姓與耶和華立約，作耶和華的子民，又使王與百姓立約。
2KGS|11|18|於是國中的眾百姓都到 巴力 廟去，拆毀了廟，徹底打碎祭壇和偶像，又在壇前把 巴力 的祭司 瑪坦 殺了。 耶何耶大 祭司派官員看守耶和華的殿，
2KGS|11|19|又率領百夫長， 迦利 人和護衛兵，以及國中的眾百姓，請王從耶和華的殿下來，由護衛兵的門進入王宮，他就坐上王位。
2KGS|11|20|國中的眾百姓都歡樂，合城也都平靜。他們已將 亞她利雅 在王宮那裏用刀殺了。
2KGS|11|21|約阿施 登基的時候年方七歲。
2KGS|12|1|耶戶 第七年， 約阿施 登基，在 耶路撒冷 作王四十年。他母親名叫 西比亞 ，是 別是巴 人。
2KGS|12|2|約阿施 在 耶何耶大 祭司教導他的一切日子，行耶和華眼中看為正的事。
2KGS|12|3|只是丘壇還沒有廢去，百姓仍在丘壇獻祭燒香。
2KGS|12|4|約阿施 對眾祭司說：「凡獻到耶和華殿分別為聖的銀子，無論是人的贖價，各人生命的贖價， 或自願獻給耶和華殿的銀子，
2KGS|12|5|祭司可以各自從認識的人收取，用來修理殿的破壞之處，就是在那裏發現的一切破壞之處。」
2KGS|12|6|然而，到了 約阿施 王第二十三年，祭司仍未修理殿的破壞之處。
2KGS|12|7|所以 約阿施 王召了 耶何耶大 祭司和眾祭司來，對他們說：「你們怎麼不修理殿的破壞之處呢？現在，不要再從認識的人收銀子了，但要為了殿的破壞之處，把銀子交出來。」
2KGS|12|8|眾祭司答應不再收百姓的銀子，也不再修理殿的破壞之處。
2KGS|12|9|耶何耶大 祭司取了一個櫃子，在櫃蓋上鑽了一個洞，放在祭壇旁，在進耶和華殿的右邊；守門的祭司將獻到耶和華殿的一切銀子投在櫃裏。
2KGS|12|10|他們見櫃裏的銀子多了，就叫王的書記和大祭司上來，將耶和華殿裏所得的銀子數點了，包起來。
2KGS|12|11|他們把秤好了的銀子交在管理耶和華殿督工的手裏，督工就支付給木匠和建造耶和華殿的工人，
2KGS|12|12|瓦匠和石匠，又買木料和鑿成的石頭，用來修理耶和華殿的破壞之處，以及其他修理殿的各項費用。
2KGS|12|13|但這些獻到耶和華殿的銀子，並沒有用來造耶和華殿裏的銀杯、鉗子、盤子、號筒和其他的金銀器皿。
2KGS|12|14|他們把這銀子交給工人，用來整修耶和華的殿。
2KGS|12|15|他們不用跟這些經手接受銀子去支付工人的人算賬，因為這些人辦事誠實。
2KGS|12|16|贖愆祭和贖罪祭的銀子沒有獻到耶和華的殿裏，都歸給祭司。
2KGS|12|17|那時， 亞蘭 王 哈薛 上來攻打 迦特 ，攻取了它。 哈薛 就定意上來攻打 耶路撒冷 。
2KGS|12|18|猶大 王 約阿施 將他祖先 猶大 王 約沙法 、 約蘭 、 亞哈謝 所分別為聖的物和自己所分別為聖的物，以及耶和華殿與王宮府庫裏所有的金子都送給 亞蘭 王 哈薛 ； 哈薛 就不上 耶路撒冷 來了。
2KGS|12|19|約阿施 其餘的事，凡他所做的，不都寫在《猶大列王記》上嗎？
2KGS|12|20|約阿施 的臣僕起來背叛，在下到 悉拉 路上的 米羅 宮那裏把他殺了。
2KGS|12|21|殺他的臣僕就是 示米押 的兒子 約撒拔 和 朔默 的兒子 約薩拔 。他與祖先同葬在 大衛城 ，他兒子 亞瑪謝 接續他作王。
2KGS|13|1|亞哈謝 的兒子 猶大 王 約阿施 第二十三年， 耶戶 的兒子 約哈斯 在 撒瑪利亞 登基作 以色列 王十七年。
2KGS|13|2|約哈斯 行耶和華眼中看為惡的事，效法 尼八 的兒子 耶羅波安 使 以色列 陷入罪裏的那罪，總不離開。
2KGS|13|3|於是，耶和華的怒氣向 以色列 發作，將他們屢次交在 亞蘭 王 哈薛 和他兒子 便‧哈達 的手裏。
2KGS|13|4|約哈斯 懇求耶和華，耶和華就應允他，因為耶和華看見 以色列 所受的欺壓，因 亞蘭 王欺壓他們。
2KGS|13|5|耶和華賜給 以色列 一位拯救者，使他們脫離 亞蘭 人的手，於是 以色列 人仍舊安居在自己的帳棚裏。
2KGS|13|6|然而他們不離開 耶羅波安 家使 以色列 陷入罪裏的那罪，仍行在罪中，並且在 撒瑪利亞 留下 亞舍拉 。
2KGS|13|7|亞蘭 王滅絕 約哈斯 的軍隊，踐踏他們如禾場上的塵沙，只給 約哈斯 留下五十騎兵，十輛戰車，一萬步兵。
2KGS|13|8|約哈斯 其餘的事，凡他所做的和他英勇的事蹟，不都寫在《以色列諸王記》上嗎？
2KGS|13|9|約哈斯 與他祖先同睡，葬在 撒瑪利亞 ，他兒子 約阿施 接續他作王。
2KGS|13|10|猶大 王 約阿施 第三十七年， 約哈斯 的兒子 約阿施 在 撒瑪利亞 登基作 以色列 王十六年。
2KGS|13|11|他行耶和華眼中看為惡的事，不離開 尼八 的兒子 耶羅波安 使 以色列 陷入罪裏的一切罪，仍行在罪中。
2KGS|13|12|約阿施 其餘的事，凡他所做的和他與 猶大 王 亞瑪謝 交戰的英勇事蹟，不都寫在《以色列諸王記》上嗎？
2KGS|13|13|約阿施 與他祖先同睡， 耶羅波安 坐上他的王位。 約阿施 與 以色列 諸王一同葬在 撒瑪利亞 。
2KGS|13|14|以利沙 得了致命的病， 以色列 王 約阿施 下來看他，伏在他臉上哭泣，說：「我父啊！我父啊！ 以色列 的戰車和騎兵啊！」
2KGS|13|15|以利沙 對他說：「把弓箭拿來。」王就拿了弓箭來。
2KGS|13|16|以利沙 對 以色列 王說：「你用手開弓。」王就用手開弓。 以利沙 按手在王的手上，
2KGS|13|17|說：「打開朝東的窗戶。」他就打開。 以利沙 說：「射箭！」他就射箭。 以利沙 說：「這是耶和華得勝的箭，是戰勝 亞蘭 人的箭，因為你必在 亞弗 攻打 亞蘭 人，直到滅盡他們。」
2KGS|13|18|以利沙 又說：「拿幾枝箭來。」他就拿了來。 以利沙 對 以色列 王說：「打地吧！」他打了三次，就停止了。
2KGS|13|19|神人向他發怒，說：「你應當擊打五六次，就能攻打 亞蘭 人直到滅盡；現在你只能打敗 亞蘭 人三次。」
2KGS|13|20|以利沙 死了，人把他埋葬了。新的一年， 摩押 人成群結隊入侵境內。
2KGS|13|21|有人正在埋葬死人，看哪，他們看見一群人來，就把死人拋在 以利沙 的墳墓裏，逃跑了。死人一碰到 以利沙 的骸骨，就活過來，用腳站了起來。
2KGS|13|22|約哈斯 在位年間， 亞蘭 王 哈薛 屢次欺壓 以色列 。
2KGS|13|23|耶和華卻因與 亞伯拉罕 、 以撒 、 雅各 所立的約，仍施恩給 以色列 人，憐憫他們，眷顧他們，不肯滅盡他們，直到現在 仍不趕逐他們離開自己面前。
2KGS|13|24|亞蘭 王 哈薛 死了，他兒子 便‧哈達 接續他作王。
2KGS|13|25|從前 哈薛 和 約阿施 的父親 約哈斯 交戰，攻取了些城鎮，現在 約哈斯 的兒子 約阿施 三次打敗 哈薛 的兒子 便‧哈達 ，從他手中收回了 以色列 的城鎮。
2KGS|14|1|約哈斯 的兒子 以色列 王 約阿施 第二年， 猶大 王 約阿施 的兒子 亞瑪謝 登基。
2KGS|14|2|他登基的時候年二十五歲，在 耶路撒冷 作王二十九年。他母親名叫 約耶但 ，是 耶路撒冷 人。
2KGS|14|3|亞瑪謝 行耶和華眼中看為正的事，但不如他祖先 大衛 。他效法他父親 約阿施 一切所行的。
2KGS|14|4|只是丘壇還沒有廢去，百姓仍在丘壇獻祭燒香。
2KGS|14|5|王國在他手裏鞏固的時候，他就把殺他父王的臣僕殺了，
2KGS|14|6|卻沒有處死殺王兇手的兒子，正如 摩西 律法書上耶和華所吩咐的說：「不可因子殺父，也不可因父殺子，各人要為自己的罪而死。」
2KGS|14|7|亞瑪謝 在 鹽谷 殺了一萬 以東 人，又在戰役中攻取了 西拉 ，稱它為 約帖 ，直到今日。
2KGS|14|8|那時， 亞瑪謝 派使者到 耶戶 的孫子， 約哈斯 的兒子 以色列 王 約阿施 那裏，說：「來，讓我們面對面較量吧！」
2KGS|14|9|以色列 王 約阿施 派人去見 猶大 王 亞瑪謝 ，說：「 黎巴嫩 的蒺藜派人去見 黎巴嫩 的香柏樹，說：『將你的女兒嫁給我的兒子。』但有一隻野獸經過 黎巴嫩 ，把蒺藜踐踏了。
2KGS|14|10|你果然打敗了 以東 ，就心高氣傲。你以此為榮，就待在自己家裏算了吧，為何要惹禍，使自己和 猶大 一同敗亡呢？」
2KGS|14|11|亞瑪謝 卻不肯聽從。於是 以色列 王 約阿施 上來，在 猶大 的 伯‧示麥 與 猶大 王 亞瑪謝 面對面較量。
2KGS|14|12|猶大 敗在 以色列 面前，他們逃跑，各人逃回自己的帳棚去了。
2KGS|14|13|以色列 王 約阿施 在 伯‧示麥 擒住 亞哈謝 的孫子， 約阿施 的兒子 猶大 王 亞瑪謝 ，就來到 耶路撒冷 ，拆毀 耶路撒冷 的城牆，從 以法蓮門 直到 角門 共四百肘。
2KGS|14|14|他又拿了耶和華殿裏與王宮府庫裏所有的金銀和器皿，並帶著人質，回 撒瑪利亞 去了。
2KGS|14|15|約阿施 其餘所做的事和他英勇的事蹟，以及他與 猶大 王 亞瑪謝 交戰的事，不都寫在《以色列諸王記》上嗎？
2KGS|14|16|約阿施 與他祖先同睡，與 以色列 諸王一同葬在 撒瑪利亞 ，他兒子 耶羅波安 接續他作王。
2KGS|14|17|約哈斯 的兒子 以色列 王 約阿施 死後， 猶大 王 約阿施 的兒子 亞瑪謝 又活了十五年。
2KGS|14|18|亞瑪謝 其餘的事，不都寫在《猶大列王記》上嗎？
2KGS|14|19|耶路撒冷 有人背叛 亞瑪謝 ， 亞瑪謝 逃往 拉吉 ；他們卻派人追到 拉吉 ，在那裏殺了他。
2KGS|14|20|有人用馬將他馱回，葬在 耶路撒冷 ，與他祖先一同葬在 大衛城 。
2KGS|14|21|猶大 眾百姓立 亞撒利雅 接續他父親 亞瑪謝 作王，那時他年十六歲。
2KGS|14|22|亞瑪謝 王與他祖先同睡之後， 亞撒利雅 收復 以拉他 回歸 猶大 ，又重新整修。
2KGS|14|23|約阿施 的兒子 猶大 王 亞瑪謝 第十五年， 以色列 王 約阿施 的兒子 耶羅波安 在 撒瑪利亞 登基，作王四十一年。
2KGS|14|24|他行耶和華眼中看為惡的事，不離開 尼八 的兒子 耶羅波安 使 以色列 陷入罪裏的一切罪。
2KGS|14|25|他收回 以色列 邊界之地，從 哈馬口 直到 亞拉巴海 ，正如耶和華－ 以色列 的上帝藉他僕人 迦特．希弗 人 亞米太 的兒子 約拿 先知所說的。
2KGS|14|26|因耶和華看見 以色列 非常艱苦的困境；沒有奴役的，沒有自由的，也沒有人來幫助 以色列 。
2KGS|14|27|耶和華並沒有說要將 以色列 的名從天下塗抹，卻要藉 約阿施 的兒子 耶羅波安 拯救他們。
2KGS|14|28|耶羅波安 其餘的事，凡他所做的和他英勇的事蹟，他怎樣作戰，怎樣收復 大馬士革 和先前屬 猶大 的 哈馬 回歸 以色列 ，不都寫在《以色列諸王記》上嗎？
2KGS|14|29|耶羅波安 與他祖先 以色列 諸王同睡，他兒子 撒迦利雅 接續他作王。
2KGS|15|1|以色列 王 耶羅波安 第二十七年， 猶大 王 亞瑪謝 的兒子 亞撒利雅 登基。
2KGS|15|2|他登基的時候年十六歲，在 耶路撒冷 作王五十二年。他母親名叫 耶可利雅 ，是 耶路撒冷 人。
2KGS|15|3|亞撒利雅 行耶和華眼中看為正的事，效法他父親 亞瑪謝 一切所行的。
2KGS|15|4|只是丘壇還沒有廢去，百姓仍在丘壇獻祭燒香。
2KGS|15|5|耶和華降災於王，使他長了痲瘋，直到死的那日。他住在隔離的行宮裏，他兒子 約坦 管理王的家，治理這地的百姓。
2KGS|15|6|亞撒利雅 其餘的事，凡他所做的，不都寫在《猶大列王記》上嗎？
2KGS|15|7|亞撒利雅 與他祖先同睡，與他祖先同葬在 大衛城 ，他兒子 約坦 接續他作王。
2KGS|15|8|猶大 王 亞撒利雅 第三十八年， 耶羅波安 的兒子 撒迦利雅 登基，在 撒瑪利亞 作 以色列 王六個月。
2KGS|15|9|他行耶和華眼中看為惡的事，效法他祖先所行的，不離開 尼八 的兒子 耶羅波安 使 以色列 陷入罪裏的那罪。
2KGS|15|10|雅比 的兒子 沙龍 背叛他，在百姓面前 擊殺他，篡了他的位。
2KGS|15|11|撒迦利雅 其餘的事，看哪，都寫在《以色列諸王記》上。
2KGS|15|12|這就是耶和華應許 耶戶 的話：「你的子孫必坐 以色列 的王位，直到第四代。」這事果然發生了。
2KGS|15|13|猶大 王 烏西雅 第三十九年， 雅比 的兒子 沙龍 登基，在 撒瑪利亞 作王一個月。
2KGS|15|14|迦底 的兒子 米拿現 從 得撒 上 撒瑪利亞 ，殺了 雅比 的兒子 沙龍 ，篡了他的位。
2KGS|15|15|沙龍 其餘的事和他陰謀背叛的事，看哪，都寫在《以色列諸王記》上。
2KGS|15|16|那時， 米拿現 從 得撒 起擊殺 提斐薩 和城中所有的人，以及它周圍的地區，因為他們沒有給他開城門。他擊殺他們，剖開其中所有的孕婦。
2KGS|15|17|猶大 王 亞撒利雅 第三十九年， 迦底 的兒子 米拿現 登基，在 撒瑪利亞 作 以色列 王十年。
2KGS|15|18|他行耶和華眼中看為惡的事，終生不離開 尼八 的兒子 耶羅波安 使 以色列 陷入罪裏的那罪。
2KGS|15|19|亞述 王 普勒 來攻擊這地， 米拿現 給他一千他連得銀子，為了請 普勒 幫助他鞏固他所掌握的國度。
2KGS|15|20|米拿現 向 以色列 所有的富豪索取銀子，要他們各出五十舍客勒，交給 亞述 王。於是 亞述 王回去了，不在境內停留。
2KGS|15|21|米拿現 其餘的事，凡他所做的，不都寫在《以色列諸王記》上嗎？
2KGS|15|22|米拿現 與他祖先同睡，他兒子 比加轄 接續他作王。
2KGS|15|23|猶大 王 亞撒利雅 第五十年， 米拿現 的兒子 比加轄 登基，在 撒瑪利亞 作 以色列 王二年。
2KGS|15|24|他行耶和華眼中看為惡的事，不離開 尼八 的兒子 耶羅波安 使 以色列 陷入罪裏的那罪。
2KGS|15|25|比加轄 的將軍， 利瑪利 的兒子 比加 背叛他，在 撒瑪利亞 王宮的堡壘殺了他。 亞珥歌伯 和 亞利耶 並 基列 的五十人幫助 比加 ； 比加 擊殺他，篡了他的位。
2KGS|15|26|比加轄 其餘的事，凡他所做的，看哪，都寫在《以色列諸王記》上。
2KGS|15|27|猶大 王 亞撒利雅 第五十二年， 利瑪利 的兒子 比加 登基，在 撒瑪利亞 作 以色列 王二十年。
2KGS|15|28|他行耶和華眼中看為惡的事，不離開 尼八 的兒子 耶羅波安 使 以色列 陷入罪裏的那罪。
2KGS|15|29|在 以色列 王 比加 的日子， 亞述 王 提革拉‧毗列色 來奪取 以雲 、 亞伯‧伯‧瑪迦 、 亞挪 、 基低斯 、 夏瑣 、 基列 、 加利利 和 拿弗他利 全地，把這些地方的居民都擄到 亞述 去了。
2KGS|15|30|烏西雅 的兒子 約坦 第二十年， 以拉 的兒子 何細亞 背叛 利瑪利 的兒子 比加 ，擊殺他，篡了他的位。
2KGS|15|31|比加 其餘的事，凡他所做的，看哪，都寫在《以色列諸王記》上。
2KGS|15|32|利瑪利 的兒子 以色列 王 比加 第二年， 猶大 王 烏西雅 的兒子 約坦 登基。
2KGS|15|33|他登基的時候年二十五歲，在 耶路撒冷 作王十六年。他母親名叫 耶路沙 ，是 撒督 的女兒。
2KGS|15|34|約坦 行耶和華眼中看為正的事，效法他父親 烏西雅 一切所行的。
2KGS|15|35|只是丘壇還沒有廢去，百姓仍在丘壇獻祭燒香。 約坦 建了耶和華殿的 上門 。
2KGS|15|36|約坦 其餘的事，凡他所做的，不都寫在《猶大列王記》上嗎？
2KGS|15|37|在那些日子，耶和華開始差 亞蘭 王 利汛 和 利瑪利 的兒子 比加 去攻擊 猶大 。
2KGS|15|38|約坦 與他祖先同睡，與他祖先同葬在 大衛城 ，他兒子 亞哈斯 接續他作王。
2KGS|16|1|利瑪利 的兒子 比加 第十七年， 猶大 王 約坦 的兒子 亞哈斯 登基。
2KGS|16|2|他登基的時候年二十歲，在 耶路撒冷 作王十六年。他不像他祖先 大衛 行耶和華－他上帝眼中看為正的事，
2KGS|16|3|卻行 以色列 諸王的道，又照著耶和華從 以色列 人面前趕出的外邦人所行可憎的事，使他的兒子經火，
2KGS|16|4|並在丘壇上、山岡上、各青翠樹下獻祭燒香。
2KGS|16|5|那時， 亞蘭 王 利汛 和 利瑪利 的兒子 以色列 王 比加 上來攻打 耶路撒冷 ，圍困 亞哈斯 ，卻不能打勝。
2KGS|16|6|當時 亞蘭 王 利汛 收復 以拉他 回歸 亞蘭 ，把 猶大 人從 以拉他 趕出去。 以東 人來到 以拉他 ，住在那裏，直到今日。
2KGS|16|7|亞哈斯 派使者到 亞述 王 提革拉‧毗列色 那裏，說：「我是你的僕人，你的兒子。現在 亞蘭 王和 以色列 王攻擊我，求你上來，救我脫離他們的手。」
2KGS|16|8|亞哈斯 將耶和華殿裏和王宮府庫裏所有的金銀都送給 亞述 王為禮物。
2KGS|16|9|亞述 王答應了他，上去攻打 大馬士革 ，攻下了城，殺了 利汛 ，把居民擄到 吉珥 。
2KGS|16|10|亞哈斯 王到 大馬士革 迎接 亞述 王 提革拉‧毗列色 ，在 大馬士革 看見一座壇。 亞哈斯 王把壇的規模和樣式，以及作法的細節，送到 烏利亞 祭司那裏。
2KGS|16|11|烏利亞 祭司照著 亞哈斯 王從 大馬士革 所送來的一切，在 亞哈斯 王還未從 大馬士革 回來之前，築了一座壇。
2KGS|16|12|王從 大馬士革 回來，看見壇，走近壇前，在壇上獻祭。
2KGS|16|13|他燒燔祭和素祭，獻澆酒祭，將平安祭牲的血灑在壇上。
2KGS|16|14|他移動耶和華面前的銅壇，從殿的前面，新壇和耶和華殿的中間，搬到新壇的北邊。
2KGS|16|15|亞哈斯 王吩咐 烏利亞 祭司說：「早晨的燔祭、晚上的素祭，王的燔祭、素祭，國內眾百姓的燔祭、素祭、澆酒祭都要燒在大壇上。燔祭牲和其他祭牲的血全都要灑在這壇上。至於銅壇，我要作求問之用。」
2KGS|16|16|烏利亞 祭司就照著 亞哈斯 王所吩咐的一切做了。
2KGS|16|17|亞哈斯 王把盆座四面的嵌邊拆下來，把盆從座上挪下來，又將銅海從馱銅海的銅牛上搬下來，放在石板鋪的地上。
2KGS|16|18|他為了 亞述 王的緣故，在耶和華的殿裏移動 殿裏為安息日所蓋的遮棚 和王從外面進來的入口。
2KGS|16|19|亞哈斯 其餘所做的事，不都寫在《猶大列王記》上嗎？
2KGS|16|20|亞哈斯 與他祖先同睡， 與他祖先同葬在 大衛城 ，他兒子 希西家 接續他作王。
2KGS|17|1|猶大 王 亞哈斯 第十二年， 以拉 的兒子 何細亞 在 撒瑪利亞 登基作 以色列 王九年。
2KGS|17|2|他行耶和華眼中看為惡的事，只是不像在他以前的 以色列 諸王。
2KGS|17|3|亞述 王 撒縵以色 上來攻擊 何細亞 ， 何細亞 就服事他，向他進貢。
2KGS|17|4|何細亞 背叛，派使者到 埃及 王 梭 那裏 ，不照往年所行的向 亞述 王進貢。 亞述 王知道了，就逮捕他，把他囚在監裏。
2KGS|17|5|亞述 王上來攻擊 以色列 全地，上到 撒瑪利亞 ，圍困這城三年。
2KGS|17|6|何細亞 第九年， 亞述 王攻取了 撒瑪利亞 ，把 以色列 人擄到 亞述 ，安置在 哈臘 與 歌散 的 哈博河 邊，以及 瑪代 人的城鎮。
2KGS|17|7|這是因為 以色列 人得罪了那領他們出 埃及 地、脫離 埃及 王法老之手的耶和華－他們的上帝，去敬畏別神，
2KGS|17|8|隨從耶和華在 以色列 人面前所趕出外邦人的風俗和 以色列 諸王所立的規條。
2KGS|17|9|以色列 人暗中行不正的事，違背耶和華－他們的上帝，在他們所有的城鎮，從瞭望樓直到堅固城，建築丘壇；
2KGS|17|10|在各高岡上、各青翠樹下立柱像和 亞舍拉 ；
2KGS|17|11|在各丘壇上燒香，效法耶和華在他們面前趕出的外邦人所行的，又行惡事，惹耶和華發怒。
2KGS|17|12|他們事奉偶像，耶和華對他們說：「你們不可做這事。」
2KGS|17|13|耶和華藉眾先知、先見勸戒 以色列 和 猶大 說：「當離開你們的惡行，謹守我的誡命律例，遵行我吩咐你們祖先、藉我僕人眾先知所傳給你們的一切律法。」
2KGS|17|14|他們卻不聽從，竟硬著頸項，像他們祖先一樣，不信服耶和華－他們的上帝。
2KGS|17|15|他們厭棄他的律例，和他與他們列祖所立的約，以及他勸戒他們的話，去隨從虛無的神明 ，自己成為虛妄，效法周圍的列國，就是耶和華囑咐他們不可效法的。
2KGS|17|16|他們離棄耶和華－他們上帝的一切誡命，為自己鑄造了兩個牛犢的像，立了 亞舍拉 ，敬拜天上的萬象，事奉 巴力 ，
2KGS|17|17|使他們的兒女經火，占卜，行法術，出賣自己，行耶和華眼中看為惡的事，惹他發怒。
2KGS|17|18|所以耶和華向 以色列 大大發怒，從自己面前趕出他們，只剩下 猶大 一個支派。
2KGS|17|19|但是， 猶大 也不遵守耶和華－他們上帝的誡命，效法 以色列 所立的規條。
2KGS|17|20|耶和華就厭棄 以色列 所有的後裔，使他們受苦，把他們交在搶奪他們的人手中，直到他把他們從自己面前趕出去。
2KGS|17|21|當他使 以色列 從 大衛 家分離出來的時候，他們立 尼八 的兒子 耶羅波安 作王。 耶羅波安 引誘 以色列 不隨從耶和華，陷入大罪中。
2KGS|17|22|以色列 人行 耶羅波安 所犯的一切罪，總不離開，
2KGS|17|23|以致耶和華把他們從自己面前趕出去，正如他藉他僕人眾先知所說的。這樣， 以色列 人從自己的土地被擄到 亞述 ，直到今日。
2KGS|17|24|亞述 王從 巴比倫 、 古他 、 亞瓦 、 哈馬 和 西法瓦音 遷移人來，安置在 撒瑪利亞 的城鎮，代替 以色列 人；他們就佔據了 撒瑪利亞 ，住在城中。
2KGS|17|25|他們開始住在那裏的時候，不敬畏耶和華，所以耶和華叫獅子進入他們中間，咬死了一些人。
2KGS|17|26|有人對 亞述 王說：「你所遷移安置在 撒瑪利亞 城鎮的各國的人，他們不知道那地之上帝的規矩，所以他叫獅子進入他們中間。看哪，獅子咬死了他們，因為他們不知道那地之上帝的規矩。」
2KGS|17|27|亞述 王吩咐說：「當派一個從那裏擄來的祭司回去，叫他住在那裏，將那地之上帝的規矩指導他們。」
2KGS|17|28|於是有一個從 撒瑪利亞 擄去的祭司回來，住在 伯特利 ，教導他們怎樣敬畏耶和華。
2KGS|17|29|然而，各國的人在所住的城裏為自己製造神像，安置在 撒瑪利亞 人所建有丘壇的廟中。
2KGS|17|30|巴比倫 人造 疏割‧比訥 像； 古他 人造 匿甲 像； 哈馬 人造 亞示瑪 像；
2KGS|17|31|亞瓦 人造 匿哈 和 他珥他 像； 西法瓦音 人用火焚燒兒女，獻給 西法瓦音 的神明 亞得米勒 和 亞拿米勒 。
2KGS|17|32|他們懼怕耶和華，卻從他們中間立丘壇的祭司，在丘壇的廟中為他們獻祭。
2KGS|17|33|他們懼怕耶和華，但又事奉自己的神明，從何邦遷來，就隨從那裏的風俗，
2KGS|17|34|直到如今仍照先前的風俗去行。 他們不敬畏耶和華，不遵守耶和華吩咐 雅各 後裔的律例、典章、律法、誡命； 雅各 就是從前耶和華起名叫 以色列 的。
2KGS|17|35|耶和華曾與他們立約，吩咐他們說：「不可敬畏別神，不可跪拜事奉它們，也不可向它們獻祭。
2KGS|17|36|惟有那用大能和伸出來的膀臂領你們出 埃及 地的耶和華，你們當敬畏他，向他跪拜，向他獻祭。
2KGS|17|37|他給你們寫的律例、典章、律法、誡命，你們應當永遠謹守遵行。你們不可敬畏別神。
2KGS|17|38|你們不可忘記我與你們所立的約，也不可敬畏別神。
2KGS|17|39|只要敬畏耶和華－你們的上帝，他必救你們脫離一切仇敵的手。」
2KGS|17|40|他們卻不聽從，仍照先前的風俗去行。
2KGS|17|41|這樣，這些國家又懼怕耶和華，又事奉他們的偶像。他們子子孫孫也都照樣行，效法他們的祖宗，直到今日。
2KGS|18|1|以拉 的兒子 以色列 王 何細亞 第三年， 猶大 王 亞哈斯 的兒子 希西家 登基。
2KGS|18|2|他登基的時候年二十五歲，在 耶路撒冷 作王二十九年。他母親名叫 亞比 ，是 撒迦利雅 的女兒。
2KGS|18|3|希西家 行耶和華眼中看為正的事，效法他祖先 大衛 一切所行的。
2KGS|18|4|他廢去丘壇，毀壞柱像，砍下 亞舍拉 ，打碎 摩西 所造的銅蛇，因為到那時 以色列 人仍向銅蛇燒香。人叫銅蛇為 尼忽士但 。
2KGS|18|5|希西家 倚靠耶和華－ 以色列 的上帝，在他之前和在他之後的 猶大 列王中沒有一個像他一樣的。
2KGS|18|6|因為他緊緊跟隨耶和華，謹守耶和華所吩咐 摩西 的誡命，總不離開。
2KGS|18|7|耶和華與他同在，他無論往何處去盡都亨通。他背叛 亞述 王，不服事他。
2KGS|18|8|希西家 攻擊 非利士 人，直到 迦薩 ，以及所屬的領土，從瞭望樓到堅固城。
2KGS|18|9|希西家 王第四年，也就是 以拉 的兒子 以色列 王 何細亞 第七年， 亞述 王 撒縵以色 上來圍困 撒瑪利亞 。
2KGS|18|10|過了三年，他們攻取了城。 希西家 第六年， 以色列 王 何細亞 第九年， 撒瑪利亞 被攻取了。
2KGS|18|11|亞述 王把 以色列 人擄到 亞述 ，安置在 哈臘 與 歌散 的 哈博河 邊，以及 瑪代 人的城鎮。
2KGS|18|12|這是因為他們不聽從耶和華－他們的上帝的話，違背了他的約；他們既不聽從，也不遵行耶和華僕人 摩西 一切所吩咐的。
2KGS|18|13|希西家 王十四年， 亞述 王 西拿基立 上來攻擊 猶大 的一切堅固的城，將城攻取。
2KGS|18|14|猶大 王 希西家 派人到 拉吉 ， 亞述 王那裏，說：「我錯了，求你撤退離開我；凡你罰我的，我必承當。」於是 亞述 王罰 猶大 王 希西家 三百他連得銀子，三十他連得金子。
2KGS|18|15|希西家 把耶和華殿裏和王宮府庫裏所有的銀子都給了他。
2KGS|18|16|那時， 猶大 王 希西家 將耶和華殿門上的金子和他自己包在柱子上的金子都刮下來，給了 亞述 王。
2KGS|18|17|亞述 王從 拉吉 差遣元帥 、太監長 和將軍 率領大軍前往 耶路撒冷 ，到 希西家 王那裏去。他們上來，到 耶路撒冷 。他們上來之後，站在 上池 的水溝旁，在往漂布地的大路上。
2KGS|18|18|他們呼叫王， 希勒家 的兒子 以利亞敬 宮廷總管， 舍伯那 書記和 亞薩 的兒子 約亞 史官就出來見他們。
2KGS|18|19|將軍對他們說：「你們去告訴 希西家 ，大王 亞述 王如此說：『你倚靠甚麼，讓你如此自信滿滿？
2KGS|18|20|你說，你有打仗的計謀和能力，我看不過是空話。你到底倚靠誰，竟敢背叛我呢？
2KGS|18|21|現在，看哪，你自己所倚靠的 埃及 是那斷裂的葦杖，人若倚靠這杖，它就刺進他的手，穿透它。 埃及 王法老向所有倚靠他的人都是這樣。
2KGS|18|22|你們若對我說：我們倚靠耶和華－我們的上帝， 希西家 豈不是將上帝的丘壇和祭壇廢去，並且吩咐 猶大 和 耶路撒冷 的人說：你們當在 耶路撒冷 這壇前敬拜嗎？
2KGS|18|23|現在你與我主 亞述 王打賭，我給你兩千匹馬，看你能否派得出騎士來騎牠們。
2KGS|18|24|若不然，怎能使我主臣僕中最小的一個軍官轉臉而逃呢？你難道要倚靠 埃及 的戰車和騎兵嗎？
2KGS|18|25|現在我上來攻擊毀滅這地方，豈不是出於耶和華嗎？耶和華吩咐我說，你上去攻擊這地，毀滅它吧！』」
2KGS|18|26|希勒家 的兒子 以利亞敬 ， 舍伯那 和 約亞 對將軍說：「求你用 亞蘭 話對僕人說，因為我們聽得懂；不要用 猶大 話對我們說，免得傳到城牆上百姓的耳中。」
2KGS|18|27|將軍對他們說：「我主差遣我來，豈是單對你和你的主人說這些話嗎？不也是對這些坐在城牆上、要與你們一同吃自己糞、喝自己尿的人說的嗎？」
2KGS|18|28|於是 亞述 將軍站著，用 猶大 話大聲喊著說：「你們當聽大王 亞述 王的話，
2KGS|18|29|王如此說：『你們不要被 希西家 欺哄了，因他不能救你們脫離我的手。
2KGS|18|30|不要聽憑 希西家 說服你們倚靠耶和華，他說，耶和華必要拯救我們，這城必不交在 亞述 王的手中。』
2KGS|18|31|你們不要聽 希西家 的話！因 亞述 王如此說：『你們要與我講和，出來投降我，各人就可以吃自己葡萄樹和無花果樹的果子，喝自己井裏的水，
2KGS|18|32|等我來領你們到一個地方，與你們本地一樣，就是有五穀和新酒之地，有糧食和葡萄園之地，有橄欖樹和蜂蜜之地，好使你們存活，不至於死。不要聽 希西家 的話，因為他誤導你們說：耶和華必拯救我們。
2KGS|18|33|列國的神明有哪一個曾救它本國脫離 亞述 王的手呢？
2KGS|18|34|哈馬 、 亞珥拔 的神明在哪裏呢？ 西法瓦音 、 希拿 、 以瓦 的神明在哪裏呢？ 它們曾救 撒瑪利亞 脫離我的手嗎？
2KGS|18|35|這些國的神明有誰曾救自己的國脫離我的手呢？難道耶和華能救 耶路撒冷 脫離我的手嗎？』」
2KGS|18|36|百姓靜默不言，一句不答，因為 希西家 王曾吩咐說：「不要回答他。」
2KGS|18|37|當下， 希勒家 的兒子 以利亞敬 宮廷總管、 舍伯那 書記和 亞薩 的兒子 約亞 史官，都撕裂衣服，來到 希西家 那裏，將 亞述 將軍的話告訴他。
2KGS|19|1|希西家 王聽見了，就撕裂衣服，披上麻布，進了耶和華的殿。
2KGS|19|2|他差遣 以利亞敬 宮廷總管和 舍伯那 書記，並祭司中年長的，都披上麻布，到 亞摩斯 的兒子 以賽亞 先知那裏去。
2KGS|19|3|他們對他說：「 希西家 如此說：『今日是急難、懲罰、凌辱的日子，就如嬰孩快要出生，卻沒有力氣生產。
2KGS|19|4|或許耶和華－你的上帝聽見 亞述 將軍一切的話，就是他主人 亞述 王差他來辱罵永生上帝的話，耶和華－你的上帝就斥責所聽見的這些話。求你為倖存的餘民揚聲禱告。』」
2KGS|19|5|希西家 王的臣僕來到 以賽亞 那裏的時候，
2KGS|19|6|以賽亞 對他們說：「要對你們的主人這樣說，耶和華如此說：『你聽見 亞述 王的僕人褻瀆我的話，不要懼怕。
2KGS|19|7|看哪，我必驚動他的心 ，他要聽見風聲就歸回本地，在那裏我必使他倒在刀下。』」
2KGS|19|8|亞述 將軍聽見 亞述 王已拔營離開 拉吉 ，就啟程返回，正遇見 亞述 王去攻打 立拿 。
2KGS|19|9|亞述 王聽見有人談論 古實 王 特哈加 說：「看哪，他出來要與你爭戰。」於是 亞述 王又差使者去見 希西家 ，說：
2KGS|19|10|「你們要對 猶大 王 希西家 如此說：『不要聽你所倚靠的上帝欺哄你說： 耶路撒冷 必不交在 亞述 王的手中。
2KGS|19|11|看哪，你總聽說 亞述 諸王向列國所行的是盡行滅絕，難道你能倖免嗎？
2KGS|19|12|我祖先所毀滅的，就是 歌散 、 哈蘭 、 利色 和 提‧拉撒 的 伊甸 人；這些國的神明何曾拯救他們呢？
2KGS|19|13|哈馬 的王， 亞珥拔 的王， 西法瓦音城 的王， 希拿 和 以瓦 的王，都在哪裏呢？』」
2KGS|19|14|希西家 從使者手裏接過書信，讀完了，就上耶和華的殿，在耶和華面前展開書信。
2KGS|19|15|希西家 向耶和華禱告說：「坐在基路伯之上耶和華－ 以色列 的上帝啊，你，惟有你是地上萬國的上帝，你創造了天和地。
2KGS|19|16|耶和華啊，求你側耳而聽；耶和華啊，求你睜眼而看，聽 西拿基立 差遣使者辱罵永生上帝的話。
2KGS|19|17|耶和華啊， 亞述 諸王果然使列國和列國之地變為荒蕪，
2KGS|19|18|將列國的神像扔在火裏，因為它們不是上帝，是人手所造的，是木頭、石頭，所以被滅絕了。
2KGS|19|19|耶和華－我們的上帝啊，現在求你救我們脫離 亞述 王的手，使地上萬國都知道惟獨你－耶和華是上帝！」
2KGS|19|20|亞摩斯 的兒子 以賽亞 差人去見 希西家 ，說：「耶和華－ 以色列 的上帝如此說：你因 亞述 王 西拿基立 的事向我祈求，我已聽見了。
2KGS|19|21|耶和華論他這樣說： 『少女 錫安 藐視你，嘲笑你； 耶路撒冷 向你搖頭。
2KGS|19|22|『你辱罵誰，褻瀆誰， 揚起聲來，高舉眼目攻擊誰呢？ 你攻擊的是 以色列 的聖者。
2KGS|19|23|你藉你的使者辱罵主說： 我率領許多戰車登上高山， 到 黎巴嫩 的頂端； 我要砍伐其中高大的香柏樹 和上好的松樹； 我必進到極遙遠的住所， 進入最茂盛的森林裏。
2KGS|19|24|我已經在外邦挖井喝水； 我必用腳掌踏乾 埃及 一切的河流。
2KGS|19|25|『你豈沒有聽見 我早先所定、古時所立、現今實現的事嗎？ 就是讓你去毀壞堅固的城鎮，使它們變為廢墟；
2KGS|19|26|城裏的居民力量微小， 他們驚惶羞愧； 像野草，像青菜， 如房頂上的草， 又如未長成而枯乾的禾稼。
2KGS|19|27|『你坐下，你出去，你進來， 你向我發烈怒，我都知道。
2KGS|19|28|因你向我發烈怒， 你的狂傲上達我耳中， 我要用鉤子鉤住你的鼻子， 將嚼環放在你口裏， 使你從原路轉回去。』
2KGS|19|29|「這是給你的預兆：你們今年要吃野生的，明年也要吃自長的；後年，你們就要耕種收割，栽葡萄園，吃其中的果子。
2KGS|19|30|猶大 家所逃脫剩餘的，仍要往下扎根，向上結果。
2KGS|19|31|必有剩餘的民從 耶路撒冷 而出，有逃脫的人從 錫安山 而來。萬軍之耶和華的熱心必成就這事。
2KGS|19|32|「所以耶和華論 亞述 王如此說：他必不得來到這城，也不在這裏射箭，不得拿盾牌到城前，也不建土堆攻城。
2KGS|19|33|他從哪條路來，必從那條路回去，必不得來到這城。這是耶和華說的。
2KGS|19|34|因我為自己的緣故，又為我僕人 大衛 的緣故，必保護拯救這城。」
2KGS|19|35|當夜，耶和華的使者出去，在 亞述 營中殺了十八萬五千人。清早有人起來，看哪，都是死屍。
2KGS|19|36|亞述 王 西拿基立 就拔營回去，住在 尼尼微 。
2KGS|19|37|一日，他在他的神明 尼斯洛 廟裏叩拜，他兒子 亞得米勒 和 沙利色 用刀殺了他，然後逃到 亞拉臘 地；他兒子 以撒．哈頓 接續他作王。
2KGS|20|1|那些日子， 希西家 病得要死， 亞摩斯 的兒子 以賽亞 先知來見他，對他說：「耶和華如此說：『你當留遺囑給你的家，因為你必死，不能活了。』」
2KGS|20|2|希西家 轉臉朝牆，向耶和華禱告說：
2KGS|20|3|「耶和華啊，求你記念我在你面前怎樣存完全的心，按誠實行事，又做你眼中看為善的事。」 希西家 就痛哭。
2KGS|20|4|以賽亞 出來，還沒有離開中院，耶和華的話就臨到他，說：
2KGS|20|5|「你回去告訴我百姓的君王 希西家 說：耶和華－你祖先 大衛 的上帝如此說：『我聽見了你的禱告，看見了你的眼淚。看哪，我必醫治你；到第三日，你必上到耶和華的殿。
2KGS|20|6|我必加添你十五年的壽數，並且我要救你和這城脫離 亞述 王的手。我為自己和我僕人 大衛 的緣故，必保護這城。』」
2KGS|20|7|以賽亞 說：「取一塊無花果餅來。」人就取了來，貼在瘡上，王就痊癒了。
2KGS|20|8|希西家 對 以賽亞 說：「耶和華必醫治我，到第三日我能上耶和華的殿，有甚麼預兆呢？」
2KGS|20|9|以賽亞 說：「耶和華必成就他所說的這話。這是耶和華給你的預兆：你要日影向前進十度呢？或是要往後退十度呢？」
2KGS|20|10|希西家 說：「日影向前進十度容易；不，讓日影往後退十度吧。」
2KGS|20|11|以賽亞 先知求告耶和華，耶和華就使 亞哈斯 日晷上照下來的日影，往後退了十度。
2KGS|20|12|那時， 巴拉但 的兒子， 巴比倫 王 米羅達‧巴拉但 聽見 希西家 生病了，就送書信和禮物給他。
2KGS|20|13|希西家 聽使者的話 ，就將自己一切寶庫裏的金子、銀子、香料、貴重的膏油和他軍械庫裏的兵器，以及他所有的財寶，都給他們看；在他家中和全國之內， 希西家 沒有一樣東西不給他們看的。
2KGS|20|14|於是 以賽亞 先知到 希西家 王那裏去，對他說：「這些人說了些甚麼？他們從哪裏來見你？」 希西家 說：「他們從遠方的 巴比倫 來。」
2KGS|20|15|以賽亞 說：「他們在你家裏看見了甚麼？」 希西家 說：「凡我家中所有的，他們都看見了；我財寶中沒有一樣東西不給他們看的。」
2KGS|20|16|以賽亞 對 希西家 說：「你要聽耶和華的話：
2KGS|20|17|耶和華說：『看哪，日子將到，凡你家裏所有的，並你祖先積蓄到如今的一切，都要被擄到 巴比倫 去，不留下一樣；
2KGS|20|18|從你本身所生的孩子，其中必有被擄到 巴比倫 王宮當太監的。』」
2KGS|20|19|希西家 對 以賽亞 說：「你所說耶和華的話甚好。」因為他想：「在我有生之年豈不是有太平和安穩嗎？」
2KGS|20|20|希西家 其餘的事和他一切英勇的事蹟，他怎樣造池、挖溝、引水入城，不都寫在《猶大列王記》上嗎？
2KGS|20|21|希西家 與他祖先同睡，他兒子 瑪拿西 接續他作王。
2KGS|21|1|瑪拿西 登基的時候年十二歲，在 耶路撒冷 作王五十五年。他母親名叫 協西巴 。
2KGS|21|2|瑪拿西 行耶和華眼中看為惡的事，效法耶和華在 以色列 人面前趕出的列國那些可憎的事。
2KGS|21|3|他重新建築他父親 希西家 所毀壞的丘壇，又為 巴力 築壇，造 亞舍拉 ，效法 以色列 王 亞哈 所行的，敬拜天上的萬象，事奉它們。
2KGS|21|4|他在耶和華殿中築壇，耶和華曾指著這殿說：「我必立我的名在 耶路撒冷 。」
2KGS|21|5|他在耶和華殿的兩個院子為天上的萬象築壇，
2KGS|21|6|並使他的兒子經火，又觀星象，行法術，求問招魂的和行巫術的，多行耶和華眼中看為惡的事，惹他發怒。
2KGS|21|7|他又把自己所造的 亞舍拉 雕像立在殿內，耶和華曾對 大衛 和他兒子 所羅門 說：「我在 以色列 眾支派中所選擇的 耶路撒冷 和這殿，必立我的名，直到永遠。
2KGS|21|8|只要 以色列 人謹守遵行我一切所吩咐的和我僕人 摩西 所吩咐的一切律法，我就不再使他們的腳挪移，離開我所賜給他們列祖之土地。」
2KGS|21|9|他們卻不聽從，並且 瑪拿西 引誘他們行惡，比耶和華在 以色列 人面前所滅的列國更嚴重。
2KGS|21|10|耶和華藉他僕人眾先知說：
2KGS|21|11|「因 猶大 王 瑪拿西 行這些可憎的惡事，比先前 亞摩利 人所行的一切更壞，使 猶大 人拜偶像，陷入罪裏，
2KGS|21|12|所以耶和華－ 以色列 的上帝如此說：看哪，我必降禍於 耶路撒冷 和 猶大 ，凡聽見的人都必雙耳齊鳴。
2KGS|21|13|我必用量 撒瑪利亞 的準繩和 亞哈 家的鉛垂線拉在 耶路撒冷 之上；我必擦拭 耶路撒冷 ，如人擦盤子，把盤子翻過來。
2KGS|21|14|我必撇棄我產業中的餘民，把他們交在仇敵手中，使他們成為所有仇敵的擄物和掠物，
2KGS|21|15|因為自從他們的祖先出 埃及 的那日直到今日，他們常行我眼中看為惡的事，惹我發怒。」
2KGS|21|16|瑪拿西 行耶和華眼中看為惡的事，使 猶大 陷入罪裏，又流許多無辜人的血，直到這血充滿了 耶路撒冷 ，從這邊到那邊。
2KGS|21|17|瑪拿西 其餘的事，凡他所做的和他所犯的罪，不都寫在《猶大列王記》上嗎？
2KGS|21|18|瑪拿西 與他祖先同睡，葬在自己王宮的園子， 烏撒 園裏，他兒子 亞們 接續他作王。
2KGS|21|19|亞們 登基的時候年二十二歲，在 耶路撒冷 作王二年。他母親名叫 米舒利密 ，是 約提巴 人 哈魯斯 的女兒。
2KGS|21|20|亞們 行耶和華眼中看為惡的事，效法他父親 瑪拿西 所行的。
2KGS|21|21|他行他父親一切所行的道，事奉他父親所事奉的偶像，敬拜它們，
2KGS|21|22|離棄耶和華－他列祖的上帝，不遵行耶和華的道。
2KGS|21|23|亞們 的臣僕背叛他，在宮裏殺了王。
2KGS|21|24|但這地的百姓殺了所有背叛 亞們 王的人；這地的百姓立他兒子 約西亞 接續他作王。
2KGS|21|25|亞們 其餘所做的事，不都寫在《猶大列王記》上嗎？
2KGS|21|26|亞們 葬在 烏撒 園內自己的墳墓裏，他兒子 約西亞 接續他作王。
2KGS|22|1|約西亞 登基的時候年八歲，在 耶路撒冷 作王三十一年。他母親名叫 耶底大 ，是 波斯加 人 亞大雅 的女兒。
2KGS|22|2|約西亞 行耶和華眼中看為正的事，行他祖先 大衛 一切所行的道，不偏左右。
2KGS|22|3|約西亞 王十八年，王派 米書蘭 的孫子， 亞薩利雅 的兒子 沙番 書記上耶和華殿去，說：
2KGS|22|4|「你上到 希勒家 大祭司那裏，請他把奉獻到耶和華殿的銀子，就是門口的守衛從百姓中收來的銀子，結算清楚，
2KGS|22|5|交在管理耶和華殿督工的手裏，由他們支付給在耶和華殿裏做工的人，好修理殿的破壞之處，
2KGS|22|6|就是木匠、工人和瓦匠，又買木料和鑿成的石頭，來整修殿宇。
2KGS|22|7|但他們不用跟這些經手接受銀子的人算帳，因為這些人辦事誠實。」
2KGS|22|8|希勒家 大祭司對 沙番 書記說：「我在耶和華殿裏發現了律法書。」 希勒家 把書遞給 沙番 ， 沙番 就讀了。
2KGS|22|9|沙番 書記到王那裏，把這事回覆王說：「你的僕人已把殿裏所發現的銀子倒出來，交在管理耶和華殿督工的手裏了。」
2KGS|22|10|沙番 書記又向王報告說：「 希勒家 祭司遞給我一卷書。」 沙番 就在王面前朗讀那書。
2KGS|22|11|王聽見律法書上的話，就撕裂衣服。
2KGS|22|12|王吩咐 希勒家 祭司與 沙番 的兒子 亞希甘 、 米該亞 的兒子 亞革波 、 沙番 書記和王的臣僕 亞撒雅 ，說：
2KGS|22|13|「你們去，以所發現這書上的話，為我、為百姓、為全 猶大 求問耶和華；因為我們祖先沒有聽從這書上的話，沒有遵照一切所寫有關我們的 去行，耶和華就向我們大發烈怒。」
2KGS|22|14|於是， 希勒家 祭司和 亞希甘 、 亞革波 、 沙番 、 亞撒雅 都去見 戶勒大 女先知，她是掌管禮服的 沙龍 的妻子； 沙龍 是 哈珥哈斯 的孫子， 特瓦 的兒子。 戶勒大 住在 耶路撒冷 第二區。他們向她請教。
2KGS|22|15|她對他們說：「耶和華－ 以色列 的上帝如此說：『你們可以回覆那派你們來見我的人說，
2KGS|22|16|耶和華如此說：看哪，我必照著 猶大 王所讀那書上的一切話，降禍於這地方和其上的居民。
2KGS|22|17|因為他們離棄我，向別神燒香，用他們手所做的一切惹我發怒，所以我的憤怒必向這地方發作，總不止息。』
2KGS|22|18|然而，派你們來求問耶和華的 猶大 王，你們要這樣回覆他：『耶和華－ 以色列 的上帝如此說：至於你所聽見的話，
2KGS|22|19|就是聽見我指著這地方和其上的居民說，要使這地方變為荒蕪、百姓受詛咒的話，你的心就軟化，在耶和華面前謙卑下來，撕裂衣服，向我哭泣，因此我應允你。這是耶和華說的。
2KGS|22|20|因此，看哪，我必使你歸到你祖先那裏，平安地進入墳墓；我要降於這地方的一切災禍，你不會親眼看見。』」他們就去把這話回覆王。
2KGS|23|1|王派人召集 猶大 和 耶路撒冷 的眾長老來。
2KGS|23|2|王和 猶大 眾人、 耶路撒冷 的居民、祭司、先知，以及所有的百姓，無論大小，都一同上到耶和華的殿去；王把耶和華殿裏所發現的約書上一切的話讀給他們聽。
2KGS|23|3|王站在柱子旁邊，在耶和華面前立約，要盡心盡性跟從耶和華，遵守他的誡命、法度、律例，實行這書上所寫這約的話。全體百姓都願遵守所立的約。
2KGS|23|4|王吩咐 希勒家 大祭司和副祭司，以及把守殿門的，把那些為 巴力 和 亞舍拉 ，以及天上萬象所造的器皿，都從耶和華殿裏搬出來，在 耶路撒冷 外 汲淪 的田間燒了，把灰拿到 伯特利 去。
2KGS|23|5|從前 猶大 列王所立拜偶像的祭司，在 猶大 城鎮的丘壇和 耶路撒冷 周圍燒香，現在王都廢去，他們是向 巴力 和日、月、行星，以及天上萬象燒香的人。
2KGS|23|6|他把 亞舍拉 從耶和華殿裏搬到 耶路撒冷 外的 汲淪溪 ，在 汲淪溪 邊焚燒，打碎成灰，把灰撒在平民的墳上。
2KGS|23|7|他又拆毀耶和華殿裏男的廟妓的屋子，就是婦女在那裏為 亞舍拉 編織衣服的屋子。
2KGS|23|8|他從 猶大 的城鎮將眾祭司帶來，從 迦巴 直到 別是巴 ，玷污祭司燒香的丘壇。他又拆毀城門旁的丘壇，這丘壇是在 約書亞 市長的城門前，在人進城門的左邊。
2KGS|23|9|只是丘壇的祭司不登 耶路撒冷 耶和華的壇，僅在他們弟兄中間吃無酵餅。
2KGS|23|10|他又玷污 欣嫩子谷 的 陀斐特 ，不許人在那裏使兒女經火獻給 摩洛 。
2KGS|23|11|他把在耶和華殿門旁、靠近 拿單‧米勒 官員走廊的屋子， 猶大 列王獻給太陽的馬廢去，且用火焚燒獻給太陽的戰車。
2KGS|23|12|猶大 列王在 亞哈斯 樓房頂上所築的壇和 瑪拿西 在耶和華殿兩院中所築的壇，王都拆毀，從那裏移走 ，把灰倒在 汲淪溪 中。
2KGS|23|13|從前 以色列 王 所羅門 在 耶路撒冷 東邊、 邪僻山 南邊為 西頓 人可憎的 亞斯她錄 、 摩押 人可憎的 基抹 、 亞捫 人可憎的 米勒公 所築的丘壇，王都玷污了，
2KGS|23|14|又打碎柱像，砍下 亞舍拉 ，用人的骨頭填滿那地方。
2KGS|23|15|此外，在 伯特利 丘壇的壇，就是 尼八 的兒子 耶羅波安 所築、使 以色列 人陷入罪裏的，他也把這壇和丘壇都拆毀了，又焚燒丘壇 ，打碎成灰，並焚燒了 亞舍拉 。
2KGS|23|16|約西亞 轉頭，看見山上的墳墓，就派人取出墳墓裏的骸骨，燒在壇上，玷污了壇，正如從前 耶羅波安 在節期中站在壇旁時，耶和華藉神人所宣告的話。 約西亞 轉頭看見了宣告這些話的神人的墳墓。
2KGS|23|17|他說：「我看見的這碑是甚麼呢？」那城裏的人對他說：「這是神人的墳墓，他從 猶大 來，宣告了王向 伯特利 的壇所做的這些事。」
2KGS|23|18|約西亞 說：「讓他安息吧！不要挪移他的骸骨。」他們就保存了他的骸骨和從 撒瑪利亞 來的那先知的骸骨。
2KGS|23|19|從前 以色列 諸王在 撒瑪利亞 的城鎮所建一切惹動怒氣的丘壇的廟， 約西亞 也都廢去了，正如他在 伯特利 所做的。
2KGS|23|20|他又把在那裏所有丘壇的祭司都殺在壇上，並在壇上燒人的骨頭。於是他回 耶路撒冷 去了。
2KGS|23|21|王吩咐眾百姓說：「你們當照這約書上所寫的，向耶和華－你們的上帝守逾越節。」
2KGS|23|22|自從士師治理 以色列 ，到 以色列 諸王、 猶大 列王在位的一切日子，從來沒有守過這樣的逾越節，
2KGS|23|23|只有在 約西亞 王十八年，才在 耶路撒冷 向耶和華守這逾越節。
2KGS|23|24|此外，在 猶大 地和 耶路撒冷 所見那些招魂的、行巫術的，家中的神像和偶像，以及一切可憎之物， 約西亞 盡都除掉，實行了 希勒家 祭司在耶和華殿裏所發現的律法書上所寫的話。
2KGS|23|25|在 約西亞 以前，沒有王像他盡心、盡性、盡力地歸向耶和華，遵行 摩西 的一切律法；在他以後，也沒有興起一個王像他。
2KGS|23|26|然而，耶和華向 猶大 所發猛烈的怒氣仍不止息，因為 瑪拿西 種種的惡事激怒了他。
2KGS|23|27|耶和華說：「我也必將 猶大 從我面前趕出，如同趕出 以色列 一樣。我必撇棄我從前所選擇的這城 耶路撒冷 和我所說我的名必留在那裏的殿。」
2KGS|23|28|約西亞 其餘的事，凡他所做的，不都寫在《猶大列王記》上嗎？
2KGS|23|29|約西亞 的日子， 埃及 王法老 尼哥 上到 幼發拉底河 ，到 亞述 王那裏； 約西亞 王去迎擊他。 埃及 王在 米吉多 看見 約西亞 ，就殺了他。
2KGS|23|30|他的臣僕用車把他的屍體從 米吉多 送到 耶路撒冷 ，葬在他自己的墳墓裏。這地的百姓選 約西亞 的兒子 約哈斯 ，膏立他，接續他父親作王。
2KGS|23|31|約哈斯 登基的時候年二十三歲，在 耶路撒冷 作王三個月。他母親名叫 哈慕她 ，是 立拿 人 耶利米 的女兒。
2KGS|23|32|約哈斯 行耶和華眼中看為惡的事，效法他祖先一切所行的。
2KGS|23|33|法老 尼哥 把 約哈斯 監禁在 哈馬 地的 利比拉 ，不許他在 耶路撒冷 作王 ，又罰這地一百他連得銀子，一他連得金子。
2KGS|23|34|法老 尼哥 立 約西亞 的兒子 以利亞敬 接續他父親 約西亞 作王，給他改名叫 約雅敬 ，卻把 約哈斯 帶到 埃及 ，他就死在那裏。
2KGS|23|35|約雅敬 進貢金銀給法老，照著法老的指示在這地徵收銀子，向這地的百姓按各人的能力索取金銀，要送給法老 尼哥 。
2KGS|23|36|約雅敬 登基的時候年二十五歲，在 耶路撒冷 作王十一年。他母親名叫 西布大 ，是 魯瑪 人 毗大雅 的女兒。
2KGS|23|37|約雅敬 行耶和華眼中看為惡的事，效法他祖先一切所行的。
2KGS|24|1|約雅敬 的日子， 巴比倫 王 尼布甲尼撒 上來； 約雅敬 服事他三年，以後又背叛他。
2KGS|24|2|耶和華派 迦勒底 、 亞蘭 、 摩押 和 亞捫 人的軍隊來攻擊 約雅敬 ；耶和華派他們來攻擊 猶大 ，要毀滅它，正如耶和華藉他僕人眾先知所說的話。
2KGS|24|3|這事臨到 猶大 ，誠然是出於耶和華的命令 ，要把 猶大 從自己面前趕出去，是因 瑪拿西 所犯的一切罪，
2KGS|24|4|又因他流無辜人的血，使無辜人的血充滿 耶路撒冷 ；耶和華不願赦免。
2KGS|24|5|約雅敬 其餘的事，凡他所做的，不都寫在《猶大列王記》上嗎？
2KGS|24|6|約雅敬 與他祖先同睡，他兒子 約雅斤 接續他作王。
2KGS|24|7|埃及 王不再從他的國出征，因為 巴比倫 王把 埃及 王所管之地，從 埃及 溪谷直到 幼發拉底河 都奪去了。
2KGS|24|8|約雅斤 登基的時候年十八歲，在 耶路撒冷 作王三個月。他母親名叫 尼護施她 ，是 耶路撒冷 人 以利拿單 的女兒。
2KGS|24|9|約雅斤 行耶和華眼中看為惡的事，效法他父親一切所行的。
2KGS|24|10|那時， 巴比倫 王 尼布甲尼撒 的軍兵上到 耶路撒冷 ，城被圍困。
2KGS|24|11|當他的軍兵圍困城的時候， 巴比倫 王 尼布甲尼撒 親自來到 耶路撒冷 。
2KGS|24|12|猶大 王 約雅斤 和他母親、臣僕、王子、官員一同出來，向 巴比倫 王投降。 巴比倫 王俘擄了他，那時是 巴比倫 王第八年。
2KGS|24|13|巴比倫 王把耶和華殿裏和王宮裏一切的寶物從那裏拿走，又把 以色列 王 所羅門 所造耶和華殿裏一切的金器都毀壞了，正如耶和華所說的。
2KGS|24|14|他把全 耶路撒冷 眾領袖和所有大能的勇士，共一萬人，連同所有的木匠和鐵匠都擄了去，只留下這地最貧窮的百姓。
2KGS|24|15|他把 約雅斤 和他的母親、后妃、官員，以及這地的貴族，都從 耶路撒冷 擄到 巴比倫 去了，
2KGS|24|16|又把所有的勇士七千人，木匠和鐵匠一千人，全是能上陣的勇士，都擄到 巴比倫 去了。
2KGS|24|17|巴比倫 王立 約雅斤 的叔父 瑪探雅 取代他作王，給 瑪探雅 改名叫 西底家 。
2KGS|24|18|西底家 登基的時候年二十一歲，在 耶路撒冷 作王十一年。他母親名叫 哈慕她 ，是 立拿 人 耶利米 的女兒。
2KGS|24|19|西底家 行耶和華眼中看為惡的事，正如 約雅敬 一切所行的。
2KGS|24|20|因此，耶和華向 耶路撒冷 和 猶大 發怒，以致把他們從自己面前趕出去。 西底家 背叛 巴比倫 王。
2KGS|25|1|西底家 作王第九年十月初十， 巴比倫 王 尼布甲尼撒 率領全軍前來攻擊 耶路撒冷 ，對城安營，四圍築堡壘攻城。
2KGS|25|2|城被圍困，直到 西底家 王十一年。
2KGS|25|3|四月初九，城裏的饑荒非常嚴重，當地的百姓都沒有糧食。
2KGS|25|4|城被攻破，士兵全都在夜間從靠近王的花園、兩城牆中間的門逃跑。 迦勒底 人正在四圍攻城，王就往 亞拉巴 逃去。
2KGS|25|5|迦勒底 的軍隊追趕王，在 耶利哥 的平原追上他；他的全軍都離開他潰散了。
2KGS|25|6|迦勒底 人就拿住王，帶他到 利比拉 的 巴比倫 王那裏；他們就判他的罪。
2KGS|25|7|他們在 西底家 眼前殺了他的兒女，挖了 西底家 的眼睛，用銅鏈鎖著他，帶到 巴比倫 去。
2KGS|25|8|巴比倫 王 尼布甲尼撒 十九年五月初七， 巴比倫 王的臣僕 尼布撒拉旦 護衛長進入 耶路撒冷 ，
2KGS|25|9|他焚燒了耶和華的殿、王宮和 耶路撒冷 一切的房屋；用火焚燒所有大戶人家的房屋。
2KGS|25|10|跟從護衛長的 迦勒底 全軍拆毀了 耶路撒冷 四圍的城牆。
2KGS|25|11|那時 尼布撒拉旦 護衛長將城裏剩下的百姓和那些投降 巴比倫 王的人，以及其餘的眾人，都擄去了。
2KGS|25|12|但護衛長留下一些當地最窮的人，叫他們修整葡萄園，耕種田地。
2KGS|25|13|耶和華殿的銅柱並殿內的盆座和銅海， 迦勒底 人都打碎了，把那些銅運到 巴比倫 去。
2KGS|25|14|他們又帶走鍋、鏟子、鉗子、勺子和供奉用的一切銅器；
2KGS|25|15|火盆和碗，無論金的銀的，護衛長都帶走了；
2KGS|25|16|還有 所羅門 為耶和華殿所造的兩根柱子、一個銅海和盆座，這一切器皿的銅多得無法可秤。
2KGS|25|17|這一根柱子高十八肘，柱上有銅頂，銅頂高三肘；銅頂的周圍有網子和石榴，也都是銅的。第二根柱子與此相同，也有網子。
2KGS|25|18|護衛長拿住 西萊雅 大祭司、 西番亞 副祭司和門口的三個守衛，
2KGS|25|19|又從城中拿住一個管理士兵的官 ，並在城裏所找到王面前的五個親信，和召募當地百姓之將軍的書記官，以及在城中找到的六十個當地百姓。
2KGS|25|20|尼布撒拉旦 護衛長把這些人帶到 利比拉 的 巴比倫 王那裏。
2KGS|25|21|巴比倫 王擊殺他們，在 哈馬 地的 利比拉 把他們處死。這樣， 猶大 人就被擄去離開本地。
2KGS|25|22|至於 猶大 地剩下的百姓，就是 巴比倫 王 尼布甲尼撒 所留下的， 巴比倫 王立了 沙番 的孫子， 亞希甘 的兒子 基大利 作他們的省長。
2KGS|25|23|所有的軍官和屬他們的人聽見 巴比倫 王立了 基大利 作省長， 尼探雅 的兒子 以實瑪利 、 加利亞 的兒子 約哈難 、 尼陀法 人 單戶蔑 的兒子 西萊雅 、 瑪迦 人的兒子 雅撒尼亞 ，和屬他們的人，都來到 米斯巴 的 基大利 那裏。
2KGS|25|24|基大利 向他們和屬他們的人起誓說：「你們不必懼怕 迦勒底 臣僕，只管住在這地，服事 巴比倫 王，就可以得福。」
2KGS|25|25|七月中，王室後裔 以利沙瑪 的孫子， 尼探雅 的兒子 以實瑪利 帶著十個人來，擊殺了 基大利 和同他在 米斯巴 的 猶大 人與 迦勒底 人，把他們殺死。
2KGS|25|26|於是眾人，無論大小，連同軍官，因為懼怕 迦勒底 人，都起身逃到 埃及 去了。
2KGS|25|27|巴比倫 王 以未‧米羅達 作王的元年，就是 猶大 王 約雅斤 被擄後三十七年，十二月二十七日，他使 猶大 王 約雅斤 抬起頭來，提他出監，
2KGS|25|28|對他說好話，使他的位高過與他一同被擄在 巴比倫 眾王的位；
2KGS|25|29|又給他脫了囚服，使他終身常在 巴比倫 王面前吃飯。
2KGS|25|30|王賜給他日常需用的食物，每日一份，終身都是這樣。
1CHR|1|1|亞當 ， 塞特 ， 以挪士 ，
1CHR|1|2|該南 ， 瑪勒列 ， 雅列 ，
1CHR|1|3|以諾 ， 瑪土撒拉 ， 拉麥 ，
1CHR|1|4|挪亞 ， 閃 ， 含 ， 雅弗 。
1CHR|1|5|雅弗 的兒子是 歌篾 、 瑪各 、 瑪代 、 雅完 、 土巴 、 米設 和 提拉 。
1CHR|1|6|歌篾 的兒子是 亞實基拿 、 低法 和 陀迦瑪 。
1CHR|1|7|雅完 的兒子是 以利沙 、 他施 、 基提 和 羅單 人 。
1CHR|1|8|含 的兒子是 古實 、 麥西 、 弗 和 迦南 。
1CHR|1|9|古實 的兒子是 西巴 、 哈腓拉 、 撒弗他 、 拉瑪 和 撒弗提迦 。 拉瑪 的兒子是 示巴 和 底但 。
1CHR|1|10|古實 又生 寧錄 ，他是地上第一個勇士。
1CHR|1|11|麥西 生 路低 人、 亞拿米 人、 利哈比 人、 拿弗土希 人、
1CHR|1|12|帕斯魯細 人、 迦斯路希 人和 迦斐託 人； 非利士 人是從 迦斐託 人 出來的。
1CHR|1|13|迦南 生了長子 西頓 ，又生 赫
1CHR|1|14|和 耶布斯 人、 亞摩利 人、 革迦撒 人、
1CHR|1|15|希未 人、 亞基 人、 西尼 人、
1CHR|1|16|亞瓦底 人、 洗瑪利 人和 哈馬 人。
1CHR|1|17|閃 的兒子是 以攔 、 亞述 、 亞法撒 、 路德 、 亞蘭 、 烏斯 、 戶勒 、 基帖 和 米設 。
1CHR|1|18|亞法撒 生 沙拉 ； 沙拉 生 希伯 。
1CHR|1|19|希伯 生了兩個兒子：一個名叫 法勒 ，因為那時人分地居住； 法勒 的兄弟名叫 約坍 。
1CHR|1|20|約坍 生 亞摩答 、 沙列 、 哈薩瑪非 、 耶拉 、
1CHR|1|21|哈多蘭 、 烏薩 、 德拉 、
1CHR|1|22|以巴錄 、 亞比瑪利 、 示巴 、
1CHR|1|23|阿斐 、 哈腓拉 和 約巴 。這些都是 約坍 的兒子。
1CHR|1|24|閃 ， 亞法撒 ， 沙拉 ，
1CHR|1|25|希伯 ， 法勒 ， 拉吳 ，
1CHR|1|26|西鹿 ， 拿鶴 ， 他拉 ，
1CHR|1|27|亞伯蘭 ， 亞伯蘭 就是 亞伯拉罕 。
1CHR|1|28|亞伯拉罕 的兒子是 以撒 和 以實瑪利 。
1CHR|1|29|以實瑪利 的後代如下： 以實瑪利 的長子是 尼拜約 ，又有 基達 、 亞德別 、 米比衫 、
1CHR|1|30|米施瑪 、 度瑪 、 瑪撒 、 哈大 、 提瑪 、
1CHR|1|31|伊突 、 拿非施 和 基底瑪 。這些都是 以實瑪利 的兒子。
1CHR|1|32|亞伯拉罕 的妾 基土拉 所生的兒子，就是 心蘭 、 約珊 、 米但 、 米甸 、 伊施巴 和 書亞 。 約珊 的兒子是 示巴 和 底但 。
1CHR|1|33|米甸 的兒子是 以法 、 以弗 、 哈諾 、 亞比大 和 以勒大 。這些都是 基土拉 的子孫。
1CHR|1|34|亞伯拉罕 生 以撒 ； 以撒 的兒子是 以掃 和 以色列 。
1CHR|1|35|以掃 的兒子是 以利法 、 流珥 、 耶烏施 、 雅蘭 和 可拉 。
1CHR|1|36|以利法 的兒子是 提幔 、 阿抹 、 洗玻 、 迦坦 、 基納斯 、 亭納 和 亞瑪力 。
1CHR|1|37|流珥 的兒子是 拿哈 、 謝拉 、 沙瑪 和 米撒 。
1CHR|1|38|西珥 的兒子是 羅坍 、 朔巴 、 祭便 、 亞拿 、 底順 、 以察 和 底珊 。
1CHR|1|39|羅坍 的兒子是 何利 和 荷幔 ； 羅坍 的妹妹是 亭納 。
1CHR|1|40|朔巴 的兒子是 亞勒文 、 瑪拿轄 、 以巴錄 、 示非 和 阿南 。 祭便 的兒子是 愛亞 和 亞拿 。
1CHR|1|41|亞拿 的兒子是 底順 。 底順 的兒子是 哈默蘭 、 伊是班 、 益蘭 和 基蘭 。
1CHR|1|42|以察 的兒子是 辟罕 、 撒番 ，和 亞干 。 底珊 的兒子是 烏斯 和 亞蘭 。
1CHR|1|43|以色列 人未有君王治理之前，這些是在 以東 地作王的。有 比珥 的兒子 比拉 ，他的城名叫 亭哈巴 。
1CHR|1|44|比拉 死了， 波斯拉 人 謝拉 的兒子 約巴 接續他作王。
1CHR|1|45|約巴 死了， 提幔 人之地的 戶珊 接續他作王。
1CHR|1|46|戶珊 死了， 比達 的兒子 哈達 接續他作王， 哈達 曾在 摩押 地擊敗 米甸 人，他的城名叫 亞未得 。
1CHR|1|47|哈達 死了， 瑪士利加 人 桑拉 接續他作王。
1CHR|1|48|桑拉 死了， 大河 邊的 利河伯 人 掃羅 接續他作王。
1CHR|1|49|掃羅 死了， 亞革波 的兒子 巴勒‧哈南 接續他作王。
1CHR|1|50|巴勒‧哈南 死了， 哈達 接續他作王，他的城名叫 巴伊 。他的妻子名叫 米希她別 ，是 米‧薩合 的孫女， 瑪特列 的女兒。
1CHR|1|51|哈達 死了。 以東 的族長有： 亭納 族長、 亞勒瓦 族長、 耶帖 族長、
1CHR|1|52|阿何利巴瑪 族長、 以拉 族長、 比嫩 族長、
1CHR|1|53|基納斯 族長、 提幔 族長、 米比薩 族長、
1CHR|1|54|瑪基疊 族長、 以蘭 族長。這些都是 以東 的族長。
1CHR|2|1|以色列 的兒子是 呂便 、 西緬 、 利未 、 猶大 、 以薩迦 、 西布倫 、
1CHR|2|2|但 、 約瑟 、 便雅憫 、 拿弗他利 、 迦得 和 亞設 。
1CHR|2|3|猶大 的兒子是 珥 、 俄南 和 示拉 ，這三人是 迦南 女子 拔．書亞 所生的。 猶大 的長子 珥 在耶和華眼中看為惡，耶和華就殺死了他。
1CHR|2|4|猶大 的媳婦 她瑪 為 猶大 生了 法勒斯 和 謝拉 。 猶大 共有五個兒子。
1CHR|2|5|法勒斯 的兒子是 希斯崙 和 哈母勒 。
1CHR|2|6|謝拉 的兒子是 心利 、 以探 、 希幔 、 甲各 和 大拉 ，共五人。
1CHR|2|7|迦米 的兒子是 亞迦 ，他在當滅的物上犯了罪，連累了 以色列 人。
1CHR|2|8|以探 的兒子是 亞撒利雅 。
1CHR|2|9|希斯崙 所生的兒子是 耶拉篾 、 蘭 和 基路拜 。
1CHR|2|10|蘭 生 亞米拿達 ； 亞米拿達 生 拿順 ， 拿順 是 猶大 人的領袖。
1CHR|2|11|拿順 生 撒門 ； 撒門 生 波阿斯 ；
1CHR|2|12|波阿斯 生 俄備得 ； 俄備得 生 耶西 ；
1CHR|2|13|耶西 生長子 以利押 ，次子 亞比拿達 ，三子 示米亞 ，
1CHR|2|14|四子 拿坦業 ，五子 拉代 ，
1CHR|2|15|六子 阿鮮 ，七子 大衛 。
1CHR|2|16|他們的姊妹是 洗魯雅 和 亞比該 。 洗魯雅 的兒子是 亞比篩 、 約押 和 亞撒黑 ，共三人。
1CHR|2|17|亞比該 生 亞瑪撒 ； 亞瑪撒 的父親是 以實瑪利 人 益帖 。
1CHR|2|18|希斯崙 的兒子 迦勒 娶 阿蘇巴 和 耶略 為妻， 阿蘇巴 的兒子是 耶設 、 朔罷 和 押墩 。
1CHR|2|19|阿蘇巴 死了， 迦勒 又娶 以法她 ，生了 戶珥 。
1CHR|2|20|戶珥 生 烏利 ； 烏利 生 比撒列 。
1CHR|2|21|後來， 希斯崙 六十歲時娶了 基列 的父親 瑪吉 的女兒，與她同房； 瑪吉 的女兒為他生了 西割 ；
1CHR|2|22|西割 生 睚珥 。 睚珥 在 基列 地有二十三座城。
1CHR|2|23|後來 基述 和 亞蘭 奪了 哈倭特．睚珥 ，以及 基納 和所屬的鄉鎮 ，共六十個。這些城鎮的人全都是 基列 的父親 瑪吉 的子孫。
1CHR|2|24|希斯崙 在 迦勒‧以法他 死後，他的妻子 亞比雅 為他生了 提哥亞 的父親 亞施戶 。
1CHR|2|25|希斯崙 的長子 耶拉篾 的兒子有長子 蘭 、 布拿 、 阿連 、 阿鮮 和 亞希雅 。
1CHR|2|26|耶拉篾 又娶一妻名叫 亞她拉 ，是 阿南 的母親。
1CHR|2|27|耶拉篾 的長子 蘭 的兒子有 瑪斯 、 雅憫 和 以結 。
1CHR|2|28|阿南 的兒子是 沙買 和 雅大 。 沙買 的兒子是 拿答 和 亞比述 。
1CHR|2|29|亞比述 的妻子名叫 亞比孩 ，為他生了 亞辦 和 摩利 。
1CHR|2|30|拿答 的兒子是 西列 和 亞遍 ； 西列 死了，沒有兒子。
1CHR|2|31|亞遍 的兒子是 以示 ； 以示 的兒子是 示珊 ； 示珊 的兒子是 亞來 。
1CHR|2|32|沙買 的兄弟 雅大 的兒子是 益帖 和 約拿單 ； 益帖 死了，沒有兒子。
1CHR|2|33|約拿單 的兒子是 比勒 和 撒薩 。這些都是 耶拉篾 的子孫。
1CHR|2|34|示珊 沒有兒子，只有女兒。 示珊 有一個僕人名叫 耶哈 ，是 埃及 人。
1CHR|2|35|示珊 把女兒嫁給僕人 耶哈 ，她為他生了 亞太 。
1CHR|2|36|亞太 生 拿單 ； 拿單 生 撒拔 ；
1CHR|2|37|撒拔 生 以弗拉 ； 以弗拉 生 俄備得 ；
1CHR|2|38|俄備得 生 耶戶 ； 耶戶 生 亞撒利雅 ；
1CHR|2|39|亞撒利雅 生 希利斯 ； 希利斯 生 以利亞薩 ；
1CHR|2|40|以利亞薩 生 西斯買 ； 西斯買 生 沙龍 ；
1CHR|2|41|沙龍 生 耶加米雅 ； 耶加米雅 生 以利沙瑪 。
1CHR|2|42|耶拉篾 的兄弟 迦勒 的眾兒子：長子是 米沙 ， 米沙 是 西弗 的父親，還有 希伯倫 的父親 瑪利沙 的眾兒子。
1CHR|2|43|希伯倫 的兒子是 可拉 、 他普亞 、 利肯 和 示瑪 。
1CHR|2|44|示瑪 生 拉含 ，是 約干 之祖。 利肯 生 沙買 。
1CHR|2|45|沙買 的兒子是 瑪雲 ； 瑪雲 是 伯‧夙 的父親。
1CHR|2|46|迦勒 的妾 以法 生 哈蘭 、 摩撒 和 迦謝 ； 哈蘭 生 迦卸 。
1CHR|2|47|雅代 的兒子是 利健 、 約坦 、 基珊 、 毗力 、 以法 和 沙亞弗 。
1CHR|2|48|迦勒 的妾 瑪迦 生 示別 和 特哈拿 ，
1CHR|2|49|又生 麥瑪拿 的父親 沙亞弗 ，又生 抹比拿 和 基比亞 的父親 示法 。 迦勒 的女兒是 押撒 。
1CHR|2|50|這些都是 迦勒 的子孫。 以法她 的長子 戶珥 的子孫： 基列‧耶琳 之祖 朔巴 ，
1CHR|2|51|伯利恆 之祖 薩瑪 ， 伯‧迦得 之祖 哈勒 。
1CHR|2|52|基列‧耶琳 之祖 朔巴 的子孫是 哈羅以 和一半的 米努哈 人 。
1CHR|2|53|基列‧耶琳 的宗族有 以帖 人、 布特 人、 舒瑪 人、 密來 人，又從這些宗族生出 瑣拉 人和 以實陶 人。
1CHR|2|54|薩瑪 的子孫有 伯利恆 人、 尼陀法 人、 亞他綠‧伯‧約押 人、一半的 瑪拿哈 人、 瑣利 人。
1CHR|2|55|住 雅比斯 的文士的宗族有 特拉 人、 示米押 人和 蘇甲 人。這些都是 利甲 家之祖 哈末 所生的 基尼 人。
1CHR|3|1|大衛 在 希伯崙 所生的兒子如下：長子 暗嫩 是 耶斯列 人 亞希暖 生的。次子 但以利 是 迦密 人 亞比該 生的。
1CHR|3|2|三子 押沙龍 是 基述 王 達買 的女兒 瑪迦 生的。四子 亞多尼雅 是 哈及 生的。
1CHR|3|3|五子 示法提雅 是 亞比她 生的。六子 以特念 是 大衛 的妻子 以格拉 生的。
1CHR|3|4|這六人都是 大衛 在 希伯崙 生的。 大衛 在 希伯崙 作王七年六個月，在 耶路撒冷 作王三十三年。
1CHR|3|5|大衛 在 耶路撒冷 所生的兒子是 示米亞 、 朔罷 、 拿單 和 所羅門 。這四人是 亞米利 的女兒 拔‧書亞 生的。
1CHR|3|6|還有 益轄 、 以利沙瑪 、 以利法列 、
1CHR|3|7|挪迦 、 尼斐 、 雅非亞 、
1CHR|3|8|以利沙瑪 、 以利雅大 、 以利法列 ，共九人。
1CHR|3|9|這些全都是 大衛 的兒子，妃嬪的兒子不在其內； 她瑪 是他們的妹妹。
1CHR|3|10|所羅門 的後裔如下： 羅波安 ，他的兒子 亞比雅 ，他的兒子 亞撒 ，他的兒子 約沙法 ，
1CHR|3|11|他的兒子 約蘭 ，他的兒子 亞哈謝 ，他的兒子 約阿施 ，
1CHR|3|12|他的兒子 亞瑪謝 ，他的兒子 亞撒利雅 ，他的兒子 約坦 ；
1CHR|3|13|他的兒子 亞哈斯 ，他的兒子 希西家 ，他的兒子 瑪拿西 ，
1CHR|3|14|他的兒子 亞們 ，他的兒子 約西亞 ，
1CHR|3|15|他的長子 約哈難 ，次子 約雅敬 ，三子 西底家 ，四子 沙龍 。
1CHR|3|16|約雅敬 的後裔：他的兒子 耶哥尼雅 ，他的兒子 西底家 。
1CHR|3|17|被擄的 耶哥尼雅 的後裔如下：他的兒子 撒拉鐵 、
1CHR|3|18|瑪基蘭 、 毗大雅 、 示拿薩 、 耶加米 、 何沙瑪 和 尼大比雅 。
1CHR|3|19|毗大雅 的兒子是 所羅巴伯 和 示每 。 所羅巴伯 的兒子是 米書蘭 和 哈拿尼雅 ， 示羅密 是他們的妹妹；
1CHR|3|20|還有 哈舒巴 、 阿黑 、 比利家 、 哈撒底 、 于沙‧希悉 ，共五人。
1CHR|3|21|哈拿尼雅 的兒子是 毗拉提 和 耶篩亞 。還有 利法雅 的眾兒子， 亞珥難 的眾兒子， 俄巴底亞 的眾兒子， 示迦尼 的眾兒子。
1CHR|3|22|示迦尼 的後裔： 示瑪雅 ， 示瑪雅 的兒子 哈突 、 以甲 、 巴利亞 、 尼利雅 、 沙法 ，共六人。
1CHR|3|23|尼利雅 的兒子是 以利約乃 、 希西家 、 亞斯利干 ，共三人。
1CHR|3|24|以利約乃 的兒子是 何大雅 、 以利亞實 、 毗萊雅 、 阿谷 、 約哈難 、 第萊雅 、 阿拿尼 ，共七人。
1CHR|4|1|猶大 的兒子是 法勒斯 、 希斯崙 、 迦米 、 戶珥 和 朔巴 。
1CHR|4|2|朔巴 的兒子 利亞雅 生 雅哈 ； 雅哈 生 亞戶買 和 拉哈 。這些是 瑣拉 人的宗族。
1CHR|4|3|以坦 之祖 是 耶斯列 、 伊施瑪 和 伊得巴 ；他們的妹妹名叫 哈悉勒玻尼 。
1CHR|4|4|基多 之祖是 毗努伊勒 。 戶沙 之祖是 以謝珥 。這些都是 伯利恆 之祖， 以法她 的長子 戶珥 的後裔。
1CHR|4|5|提哥亞 的父親 亞施戶 有兩個妻子， 希拉 和 拿拉 。
1CHR|4|6|拿拉 為 亞施戶 生 亞戶撒 、 希弗 、 提米尼 和 哈轄斯他利 。這些都是 拿拉 的兒子。
1CHR|4|7|希拉 生的是 洗列 、 瑣轄 和 伊提南 。
1CHR|4|8|哥斯 生 亞諾 、 瑣比巴 和 哈崙 的兒子 亞哈黑 的宗族。
1CHR|4|9|雅比斯 比他眾兄弟更尊貴，他母親給他起名叫 雅比斯 ，意思說：「我生他甚是痛苦。」
1CHR|4|10|雅比斯 求告 以色列 的上帝說：「甚願你賜福與我，擴張我的疆界，你的手常與我同在，保佑我不遭患難，不受艱苦。」上帝就應允他所求的。
1CHR|4|11|書哈 的兄弟 基綠 生 米黑 ， 米黑 是 伊施屯 的父親。
1CHR|4|12|伊施屯 生 伯拉巴 、 巴西亞 和 珥．拿轄 之祖 提欣拿 。這些都是 利迦 人。
1CHR|4|13|基納斯 的兒子是 俄陀聶 和 西萊雅 。 俄陀聶 的兒子是 哈塔 。
1CHR|4|14|憫挪太 生 俄弗拉 ； 西萊雅 生 革‧夏納欣 之祖 約押 。他們都是工匠。
1CHR|4|15|耶孚尼 的兒子 迦勒 的後裔： 以路 、 以拉 和 拿安 。 以拉 的兒子是 基納斯 。
1CHR|4|16|耶哈利勒 的兒子是 西弗 、 西法 、 提利 和 亞撒列 。
1CHR|4|17|以斯拉 的兒子是 益帖 、 米列 、 以弗 和 雅倫 。 米列 所娶法老的女兒 比提雅 的後裔如下：她懷了 米利暗 、 沙買 ，和 以實提摩 之祖 益巴 。 米列 的 猶大 妻子生 基多 之祖 雅列 ， 梭哥 之祖 希伯 ，和 撒挪亞 之祖 耶古鐵 。
1CHR|4|18|
1CHR|4|19|拿含 的妹妹， 荷第雅 的妻子所生的是 達利亞 ， 迦米 人 基伊拉 和 瑪迦 人 以實提摩 的祖先。
1CHR|4|20|示門 的兒子是 暗嫩 、 林拿 、 便‧哈南 和 提倫 。 以示 的兒子是 梭黑 和 便‧梭黑 。
1CHR|4|21|猶大 的兒子 示拉 的後裔： 利迦 之祖 珥 ， 瑪利沙 之祖 拉大 ，和住在 伯‧亞實比 織細麻布的各宗族。
1CHR|4|22|還有 約敬 、 哥西巴 人、 約阿施 ，和那在 摩押 娶妻，回到 利恆 的 薩拉 。這都是古時的記載。
1CHR|4|23|這些人都是陶匠，是 尼他應 和 基底拉 的居民。他們住在王那裏，為王做工。
1CHR|4|24|西緬 的後裔如下： 尼母利 、 雅憫 、 雅立 、 謝拉 和 掃羅 ；
1CHR|4|25|他的兒子 沙龍 ，他的兒子 米比衫 ，他的兒子 米施瑪 ；
1CHR|4|26|米施瑪 的後裔：他的兒子 哈母利 ，他的兒子 撒刻 ，他的兒子 示每 。
1CHR|4|27|示每 有十六個兒子和六個女兒，但他兄弟的兒女不多，他們各家族也不如 猶大 族那樣人丁興旺。
1CHR|4|28|西緬 人住在 別是巴 、 摩拉大 、 哈薩‧書亞 、
1CHR|4|29|辟拉 、 以森 、 陀臘 、
1CHR|4|30|彼土利 、 何珥瑪 、 洗革拉 、
1CHR|4|31|伯‧瑪加博 、 哈薩‧蘇撒 、 伯‧比利 和 沙拉音 ，這些城鎮直到 大衛 作王的時候都是屬 西緬 人的；
1CHR|4|32|還有所屬的村莊 以坦 、 亞因 、 臨門 、 陀健 、 亞珊 ，共五個城鎮；
1CHR|4|33|連同環繞這些城鎮的一切鄉村，直到 巴力 。這是他們的住處，他們都有家譜。
1CHR|4|34|還有 米所巴 、 雅米勒 、 亞瑪謝 的兒子 約沙 、
1CHR|4|35|約珥 ，和 亞薛 的曾孫， 西萊雅 的孫子， 約示比 的兒子 耶戶 。
1CHR|4|36|還有 以利約乃 、 雅哥巴 、 約朔海 、 亞帥雅 、 亞底業 、 耶西篾 、 比拿雅 、
1CHR|4|37|細撒 ； 細撒 是 示非 的兒子， 示非 是 亞龍 的兒子， 亞龍 是 耶大雅 的兒子， 耶大雅 是 申利 的兒子， 申利 是 示瑪雅 的兒子。
1CHR|4|38|以上所記的人名都是作族長的，他們父系的家屬大量增加。
1CHR|4|39|他們往平原東邊 基多口 去，尋找牧放羊群的草場，
1CHR|4|40|找到了肥沃優美的草場，又寬闊又平靜安寧之地；從前住那裏的是 含 族的人。
1CHR|4|41|以上紀錄上有名的人，在 猶大 王 希西家 的日子，來攻擊 含 族人的帳棚和那裏所有的 米烏尼 人，把他們滅盡，就住在他們的地方，直到今日，因為那裏有草場可以牧放羊群。
1CHR|4|42|這些 西緬 人中有五百人上 西珥山 ，率領他們的是 以示 的兒子 毗拉提 、 尼利雅 、 利法雅 和 烏薛 。
1CHR|4|43|他們殺了 亞瑪力 剩下的殘存之民，就住在那裏，直到今日。
1CHR|5|1|以色列 的長子 呂便 的後裔。 呂便 玷污了父親的床，他長子的名分就歸了 以色列 的兒子 約瑟 的後裔；因此，家譜就不按出生順序登錄。
1CHR|5|2|雖然 猶大 比他兄弟強盛，君王也從他而出，然而長子的名分卻歸 約瑟 。
1CHR|5|3|以色列 長子 呂便 的後裔如下： 哈諾 、 法路 、 希斯倫 和 迦米 。
1CHR|5|4|約珥 的後裔：他的兒子 示瑪雅 ，他的兒子 歌革 ，他的兒子 示每 ，
1CHR|5|5|他的兒子 米迦 ，他的兒子 利亞雅 ，他的兒子 巴力 ，
1CHR|5|6|他的兒子 備拉 ；這 備拉 作 呂便 支派的領袖，被 亞述 王 提革拉‧毗列色 擄去。
1CHR|5|7|他的弟兄照著宗族，按著家譜作族長的是 耶利 、 撒迦利雅 、
1CHR|5|8|比拉 ； 比拉 是 亞撒 的兒子， 亞撒 是 示瑪 的兒子， 示瑪 是 約珥 的兒子； 約珥 住在 亞羅珥 ，直到 尼波 和 巴力‧免 。
1CHR|5|9|他也住在東邊，直到 幼發拉底河 這邊的曠野邊界，因為他們在 基列 地牲畜增多。
1CHR|5|10|掃羅 年間，他們與 夏甲 人爭戰， 夏甲 人倒在他們手下，他們就在 基列 東邊的全地，住在 夏甲 人的帳棚裏。
1CHR|5|11|迦得 的後裔在 呂便 對面，住在 巴珊 地，延伸到 撒迦 ：
1CHR|5|12|有作族長的 約珥 ，有作副族長的 沙番 ，還有 雅乃 和住在 巴珊 的 沙法 。
1CHR|5|13|按著家族，他們的弟兄是 米迦勒 、 米書蘭 、 示巴 、 約賴 、 雅干 、 細亞 和 希伯 ，共七人。
1CHR|5|14|這些都是 亞比孩 的兒子； 亞比孩 是 戶利 的兒子， 戶利 是 耶羅亞 的兒子， 耶羅亞 是 基列 的兒子， 基列 是 米迦勒 的兒子， 米迦勒 是 耶示篩 的兒子， 耶示篩 是 耶哈多 的兒子， 耶哈多 是 布斯 的兒子；
1CHR|5|15|古尼 的孫子， 押比疊 的兒子 亞希 是他們的族長。
1CHR|5|16|他們住在 基列 、 巴珊 和所屬的鄉鎮，以及 沙崙 一切的郊野，直到四圍的交界。
1CHR|5|17|這些人在 猶大 王 約坦 和 以色列 王 耶羅波安 年間，都載入家譜。
1CHR|5|18|呂便 人、 迦得 人和 瑪拿西 半支派的人，能拿盾牌和刀劍、拉弓、出征善戰的勇士共有四萬四千七百六十名。
1CHR|5|19|他們與 夏甲 人、 伊突 人、 拿非施 人、 挪答 人打仗。
1CHR|5|20|他們在打仗的時候得了上帝的幫助， 夏甲 人和所有跟隨 夏甲 人的人都交在他們手中；因為他們在陣上呼求上帝，倚賴他，他就應允他們。
1CHR|5|21|他們擄掠了 夏甲 人的牲畜，有五萬匹駱駝，二十五萬隻羊，二千匹驢，又有十萬人；
1CHR|5|22|被殺仆倒的很多，因為這戰爭是出乎上帝。他們就住在 夏甲 人的地上，直到被擄的時候。
1CHR|5|23|瑪拿西 半支派的人住在那地，從 巴珊 延到 巴力‧黑門 、 示尼珥 和 黑門山 ，他們人數增多 。
1CHR|5|24|他們的族長如下： 以弗 、 以示 、 以利業 、 亞斯列 、 耶利米 、 何達威雅 和 雅疊 ；他們都是大能的勇士，有名的人，是作族長的。
1CHR|5|25|但他們得罪了他們列祖的上帝，隨從當地百姓的神明而行淫，這百姓就是上帝在他們面前所除滅的。
1CHR|5|26|因此， 以色列 的上帝激發 亞述 王 普勒 ，就是 亞述 王 提革拉‧毗列色 的心，他擄掠了 呂便 人、 迦得 人、 瑪拿西 半支派的人，把他們帶到 哈臘 、 哈博 、 哈拉 與 歌散河 邊，直到今日。
1CHR|6|1|利未 的後裔： 革順 、 哥轄 和 米拉利 。
1CHR|6|2|哥轄 的兒子是 暗蘭 、 以斯哈 、 希伯倫 和 烏薛 。
1CHR|6|3|暗蘭 的兒女是 亞倫 、 摩西 和 米利暗 。 亞倫 的兒子是 拿答 、 亞比戶 、 以利亞撒 和 以他瑪 。
1CHR|6|4|以利亞撒 生 非尼哈 ； 非尼哈 生 亞比書 ；
1CHR|6|5|亞比書 生 布基 ； 布基 生 烏西 ；
1CHR|6|6|烏西 生 西拉希雅 ； 西拉希雅 生 米拉約 ；
1CHR|6|7|米拉約 生 亞瑪利雅 ； 亞瑪利雅 生 亞希突 ；
1CHR|6|8|亞希突 生 撒督 ； 撒督 生 亞希瑪斯 ；
1CHR|6|9|亞希瑪斯 生 亞撒利雅 ； 亞撒利雅 生 約哈難 ；
1CHR|6|10|約哈難 生 亞撒利雅 ， 亞撒利雅 在 所羅門 建造的 耶路撒冷 殿中擔任祭司的職分；
1CHR|6|11|亞撒利雅 生 亞瑪利雅 ； 亞瑪利雅 生 亞希突 ；
1CHR|6|12|亞希突 生 撒督 ； 撒督 生 沙龍 ；
1CHR|6|13|沙龍 生 希勒家 ； 希勒家 生 亞撒利雅 ；
1CHR|6|14|亞撒利雅 生 西萊雅 ； 西萊雅 生 約薩答 。
1CHR|6|15|當耶和華藉 尼布甲尼撒 的手擄掠 猶大 和 耶路撒冷 的時候， 約薩答 也被擄去。
1CHR|6|16|利未 的後裔： 革順 、 哥轄 和 米拉利 。
1CHR|6|17|革順 的兒子名叫 立尼 和 示每 。
1CHR|6|18|哥轄 的兒子是 暗蘭 、 以斯哈 、 希伯倫 和 烏薛 。
1CHR|6|19|米拉利 的兒子是 抹利 和 母示 。這是按著父系所分 利未 人的宗族。
1CHR|6|20|屬 革順 的：他的兒子 立尼 ，他的兒子 雅哈 ，他的兒子 薪瑪 ，
1CHR|6|21|他的兒子 約亞 ，他的兒子 易多 ，他的兒子 謝拉 ，他的兒子 耶特賴 。
1CHR|6|22|哥轄 的後裔：他的兒子 亞米拿達 ，他的兒子 可拉 ，他的兒子 亞惜 ，
1CHR|6|23|他的兒子 以利加拿 ，他的兒子 以比雅撒 ，他的兒子 亞惜 ，
1CHR|6|24|他的兒子 他哈 ，他的兒子 烏列 ，他的兒子 烏西雅 ，他的兒子 少羅 。
1CHR|6|25|以利加拿 的兒子是 亞瑪賽 、 亞希摩 、
1CHR|6|26|以利加拿 。 以利加拿 的後裔：他的兒子 瑣菲 ，他的兒子 拿哈 ，
1CHR|6|27|他的兒子 以利押 ，他的兒子 耶羅罕 ，他的兒子 以利加拿 ，他的兒子 撒母耳 。
1CHR|6|28|撒母耳 的兒子是長子 約珥 和次子 亞比亞 。
1CHR|6|29|米拉利 的後裔： 抹利 ，他的兒子 立尼 ，他的兒子 示每 ，他的兒子 烏撒 ，
1CHR|6|30|他的兒子 示米亞 ，他的兒子 哈基雅 ，他的兒子 亞帥雅 。
1CHR|6|31|這些是約櫃安設之後， 大衛 派在耶和華殿中管理歌唱事奉的人。
1CHR|6|32|他們在會幕前負責歌唱的事奉，及至 所羅門 在 耶路撒冷 建造了耶和華的殿，他們就按著班次供職。
1CHR|6|33|供職的人和他們的子孫如下： 哥轄 的子孫中有歌唱的 希幔 ； 希幔 是 約珥 的兒子， 約珥 是 撒母耳 的兒子，
1CHR|6|34|撒母耳 是 以利加拿 的兒子， 以利加拿 是 耶羅罕 的兒子， 耶羅罕 是 以利業 的兒子， 以利業 是 陀亞 的兒子，
1CHR|6|35|陀亞 是 蘇弗 的兒子， 蘇弗 是 以利加拿 的兒子， 以利加拿 是 瑪哈 的兒子， 瑪哈 是 亞瑪賽 的兒子，
1CHR|6|36|亞瑪賽 是 以利加拿 的兒子， 以利加拿 是 約珥 的兒子， 約珥 是 亞撒利雅 的兒子， 亞撒利雅 是 西番雅 的兒子，
1CHR|6|37|西番雅 是 他哈 的兒子， 他哈 是 亞惜 的兒子， 亞惜 是 以比雅撒 的兒子， 以比雅撒 是 可拉 的兒子，
1CHR|6|38|可拉 是 以斯哈 的兒子， 以斯哈 是 哥轄 的兒子， 哥轄 是 利未 的兒子， 利未 是 以色列 的兒子。
1CHR|6|39|希幔 的弟兄 亞薩 在 希幔 的右邊供職； 亞薩 是 比利家 的兒子， 比利家 是 示米亞 的兒子，
1CHR|6|40|示米亞 是 米迦勒 的兒子， 米迦勒 是 巴西雅 的兒子， 巴西雅 是 瑪基雅 的兒子，
1CHR|6|41|瑪基雅 是 伊特尼 的兒子， 伊特尼 是 謝拉 的兒子， 謝拉 是 亞大雅 的兒子，
1CHR|6|42|亞大雅 是 以探 的兒子， 以探 是 薪瑪 的兒子， 薪瑪 是 示每 的兒子，
1CHR|6|43|示每 是 雅哈 的兒子， 雅哈 是 革順 的兒子， 革順 是 利未 的兒子。
1CHR|6|44|他們的弟兄 米拉利 的子孫，在他們左邊供職的有 以探 ； 以探 是 基示 的兒子， 基示 是 亞伯底 的兒子， 亞伯底 是 瑪鹿 的兒子，
1CHR|6|45|瑪鹿 是 哈沙比雅 的兒子， 哈沙比雅 是 亞瑪謝 的兒子， 亞瑪謝 是 希勒家 的兒子，
1CHR|6|46|希勒家 是 暗西 的兒子， 暗西 是 巴尼 的兒子， 巴尼 是 沙麥 的兒子，
1CHR|6|47|沙麥 是 末力 的兒子， 末力 是 母示 的兒子， 母示 是 米拉利 的兒子， 米拉利 是 利未 的兒子。
1CHR|6|48|他們的弟兄 利未 人也被派辦理上帝殿中帳幕的一切事務。
1CHR|6|49|亞倫 和他的子孫在燔祭壇和香壇上獻祭燒香，辦理至聖所一切的事，為 以色列 贖罪，正如上帝僕人 摩西 所吩咐的一切。
1CHR|6|50|亞倫 的後裔如下：他的兒子 以利亞撒 ，他的兒子 非尼哈 ，他的兒子 亞比書 ，
1CHR|6|51|他的兒子 布基 ，他的兒子 烏西 ，他的兒子 西拉希雅 ，
1CHR|6|52|他的兒子 米拉約 ，他的兒子 亞瑪利雅 ，他的兒子 亞希突 ，
1CHR|6|53|他的兒子 撒督 ，他的兒子 亞希瑪斯 。
1CHR|6|54|他們的住處按著境內的營寨如下： 亞倫 的子孫 哥轄 族先抽籤得地，
1CHR|6|55|得了 猶大 地的 希伯崙 和四圍的郊野；
1CHR|6|56|只是這城的田地和所屬的村莊都為 耶孚尼 的兒子 迦勒 所得。
1CHR|6|57|亞倫 的子孫所得逃城如下： 希伯崙 、 立拿 與其郊野、 雅提珥 、 以實提莫 與其郊野、
1CHR|6|58|希崙 與其郊野、 底璧 與其郊野、
1CHR|6|59|亞珊 與其郊野、 伯‧示麥 與其郊野。
1CHR|6|60|他們也從 便雅憫 支派中得了 迦巴 與其郊野、 阿勒篾 與其郊野、 亞拿突 與其郊野。他們宗族所得的城共十三座。
1CHR|6|61|哥轄 族其餘的人抽籤，按支派的宗族，從半個支派，就是 瑪拿西 半支派中得了十座城。
1CHR|6|62|革順 族按著宗族，從 以薩迦 支派、 亞設 支派、 拿弗他利 支派、 巴珊 內的 瑪拿西 支派中，得了十三座城。
1CHR|6|63|米拉利 族按著宗族抽籤，從 呂便 支派、 迦得 支派、 西布倫 支派中，得了十二座城。
1CHR|6|64|以色列 人把這些城與其郊野給了 利未 人。
1CHR|6|65|以色列 人用抽籤的方式，從 猶大 人、 西緬 人、 便雅憫 人三支派中，把以上提到名字的城給了他們。
1CHR|6|66|哥轄 子孫中有幾個宗族從 以法蓮 支派中也得了城鎮作為他們的區域。
1CHR|6|67|他們在 以法蓮 山區所得的逃城： 示劍 與其郊野、 基色 與其郊野、
1CHR|6|68|約緬 與其郊野、 伯‧和崙 與其郊野、
1CHR|6|69|亞雅崙 與其郊野、 迦特‧臨門 與其郊野。
1CHR|6|70|哥轄 其餘的子孫從 瑪拿西 半支派中得了 亞乃 與其郊野、 比連 與其郊野。
1CHR|6|71|革順 子孫從 瑪拿西 半支派中得了 巴珊 的 哥蘭 與其郊野、 亞斯她錄 與其郊野；
1CHR|6|72|從 以薩迦 支派中得了 基低斯 與其郊野、 大比拉 與其郊野、
1CHR|6|73|拉末 與其郊野、 亞年 與其郊野；
1CHR|6|74|從 亞設 支派中得了 瑪沙 與其郊野、 押頓 與其郊野、
1CHR|6|75|戶割 與其郊野、 利合 與其郊野；
1CHR|6|76|從 拿弗他利 支派中得了 加利利 的 基低斯 與其郊野、 哈們 與其郊野、 基列亭 與其郊野。
1CHR|6|77|米拉利 其餘的子孫從 西布倫 支派中得了 臨摩挪 與其郊野、 他泊 與其郊野；
1CHR|6|78|又在 耶利哥 的 約旦河 東，從 呂便 支派中得了曠野的 比悉 與其郊野、 雅雜 與其郊野，
1CHR|6|79|基底莫 與其郊野、 米法押 與其郊野；
1CHR|6|80|又從 迦得 支派中得了 基列 的 拉末 與其郊野、 瑪哈念 與其郊野、
1CHR|6|81|希實本 與其郊野、 雅謝 與其郊野。
1CHR|7|1|以薩迦 的後裔： 陀拉 、 普瓦 、 雅述 和 伸崙 ，共四人。
1CHR|7|2|陀拉 的後裔： 烏西 、 利法雅 、 耶勒 、 雅買 、 易伯散 和 示母利 ，都是 陀拉 的族長，在他們世代中是大能的勇士。到 大衛 年間，他們的人數共有二萬二千六百名。
1CHR|7|3|烏西 的後裔： 伊斯拉希 ， 伊斯拉希 的兒子 米迦勒 、 俄巴底亞 、 約珥 和 伊示雅 ，共五人，全都是族長。
1CHR|7|4|他們所率領的，按著家譜，照著父家，可作戰的軍隊共有三萬六千人，因為他們的妻子和兒子眾多。
1CHR|7|5|他們的弟兄在 以薩迦 各族中的大能勇士，登記在家譜中的全部共有八萬七千人。
1CHR|7|6|便雅憫 ： 比拉 、 比結 和 耶疊 ，共三人。
1CHR|7|7|比拉 的兒子： 以斯本 、 烏西 、 烏薛 、 耶利末 和 以利 ，共五人，都是族長，是大能的勇士。登記在家譜中的人共有二萬二千零三十四人。
1CHR|7|8|比結 的兒子： 細米拉 、 約阿施 、 以利以謝 、 以利約乃 、 暗利 、 耶列末 、 亞比雅 、 亞拿突 和 亞拉篾 ；這些全都是 比結 的兒子。
1CHR|7|9|登記在家譜中，按家譜的族長，大能的勇士，共有二萬零二百人。
1CHR|7|10|耶疊 的後裔： 比勒罕 ， 比勒罕 的兒子 耶烏施 、 便雅憫 、 以笏 、 基拿拿 、 細坦 、 他施 和 亞希沙哈 。
1CHR|7|11|這些全都是 耶疊 的後裔，都是族長，是大能的勇士，能上陣打仗的共有一萬七千二百人。
1CHR|7|12|還有 以珥 的兒子 書品 和 戶品 ，以及 亞黑 的兒子 戶伸 。
1CHR|7|13|拿弗他利 的後裔： 雅薛 、 沽尼 、 耶色 和 沙龍 ，都是 辟拉 的子孫。
1CHR|7|14|瑪拿西 的兒子 亞斯烈 是他的妾 亞蘭 女子所生的；她又生了 瑪吉 ，是 基列 的父親。
1CHR|7|15|瑪吉 為 戶品 和 書品 各娶了一妻，他的姊妹名叫 瑪迦 。第二個名叫 西羅非哈 ； 西羅非哈 只有女兒。
1CHR|7|16|瑪吉 的妻子 瑪迦 生了一個兒子， 瑪迦 給他起名叫 毗利施 。 毗利施 的弟弟名叫 示利施 ； 示利施 的兒子是 烏蘭 和 利金 。
1CHR|7|17|烏蘭 的兒子是 比但 。這些都是 基列 的子孫； 基列 是 瑪吉 的兒子， 瑪吉 是 瑪拿西 的兒子。
1CHR|7|18|基列 的妹妹 哈摩利吉 生了 伊施荷 、 亞比以謝 和 瑪拉 。
1CHR|7|19|示米大 的兒子是 亞現 、 示劍 、 利克希 和 阿尼安 。
1CHR|7|20|以法蓮 的後裔： 書提拉 ，他的兒子 比列 ，他的兒子 他哈 ，他的兒子 以拉大 ，他的兒子 他哈 ，
1CHR|7|21|他的兒子 撒拔 ，他的兒子 書提拉 。 以法蓮 又生 以謝 和 以列 ；這二人因為下去奪取 迦特 人的牲畜，被本地的 迦特 人殺了。
1CHR|7|22|他們的父親 以法蓮 為他們悲哀了多日，他的兄弟都來安慰他。
1CHR|7|23|以法蓮 與妻子同房，妻子懷孕生了一子， 以法蓮 因為家裏遭禍，就給這兒子起名叫 比利亞 。
1CHR|7|24|他的女兒名叫 舍伊拉 ， 舍伊拉 建築了 上伯‧和崙 、 下伯‧和崙 和 烏羨‧舍伊拉 。
1CHR|7|25|他的兒子 利法 和 利悉 ，他的兒子 他拉 ，他的兒子 他罕 ，
1CHR|7|26|他的兒子 拉但 ，他的兒子 亞米忽 ，他的兒子 以利沙瑪 ，
1CHR|7|27|他的兒子 嫩 ，他的兒子 約書亞 。
1CHR|7|28|以法蓮 人的地業和住處是 伯特利 和所屬的鄉鎮，東邊 拿蘭 ，西邊 基色 和所屬的鄉鎮， 示劍 和所屬的鄉鎮，直到 艾雅 和所屬的鄉鎮；
1CHR|7|29|還有靠近 瑪拿西 人的邊界， 伯‧善 和所屬的鄉鎮， 他納 和所屬的鄉鎮， 米吉多 和所屬的鄉鎮， 多珥 和所屬的鄉鎮。 以色列 兒子 約瑟 的子孫住在這些地方。
1CHR|7|30|亞設 的後裔： 音拿 、 亦施瓦 、 亦施韋 和 比利亞 ，還有他們的妹妹 西拉 。
1CHR|7|31|比利亞 的兒子是 希別 和 瑪結 ； 瑪結 是 比撒威 的父親。
1CHR|7|32|希別 生 雅弗勒 、 朔默 、 何坦 和他們的妹妹 書雅 。
1CHR|7|33|雅弗勒 的兒子是 巴薩 、 賓哈 和 亞施法 ；這些都是 雅弗勒 的兒子。
1CHR|7|34|朔默 的兒子是 亞希 、 羅迦 、 耶戶巴 和 亞蘭 。
1CHR|7|35|朔默 的兄弟 希連 的兒子是 瑣法 、 音那 、 示利斯 和 亞抹 。
1CHR|7|36|瑣法 的兒子是 書亞 、 哈尼弗 、 書阿勒 、 比利 、 音拉 、
1CHR|7|37|比悉 、 河得 、 珊瑪 、 施沙 、 益蘭 和 比拉 。
1CHR|7|38|益帖 的兒子是 耶孚尼 、 毗斯巴 和 亞拉 。
1CHR|7|39|烏拉 的兒子是 亞拉 、 漢尼業 和 利寫 。
1CHR|7|40|這些全都是 亞設 的子孫，都是族長，是精壯大能的勇士，也是領袖中的領袖。登記在家譜中，能上陣打仗的共有二萬六千人。
1CHR|8|1|便雅憫 生長子 比拉 ，次子 亞實別 ，三子 亞哈拉 ，
1CHR|8|2|四子 挪哈 ，五子 拉法 。
1CHR|8|3|比拉 的兒子是 亞大 、 基拉 、 亞比忽 、
1CHR|8|4|亞比書 、 乃幔 、 亞何亞 、
1CHR|8|5|基拉 、 示孚汛 和 戶蘭 。
1CHR|8|6|以忽 的後裔如下，他們是 迦巴 居民的族長，曾被擄到 瑪拿轄 ：
1CHR|8|7|乃幔 、 亞希亞 、 基拉 ；他擄了他們，又生了 烏撒 和 亞希忽 。
1CHR|8|8|沙哈連 休了兩個妻子 戶伸 和 巴拉 之後，在 摩押 地生了兒子。
1CHR|8|9|他與妻子 賀得 生了 約巴 、 洗比雅 、 米沙 、 瑪拉干 、
1CHR|8|10|耶烏斯 、 沙迦 和 米瑪 ；這些是他的兒子，都是族長。
1CHR|8|11|戶伸 為他生了 亞比突 和 以利巴力 。
1CHR|8|12|以利巴力 的兒子是 希伯 、 米珊 和 沙麥 ； 沙麥 建立 阿挪 、 羅德 和所屬的鄉鎮。
1CHR|8|13|比利亞 和 示瑪 是 亞雅崙 居民的族長，他們驅逐了 迦特 的居民。
1CHR|8|14|亞希約 、 沙煞 、 耶列末 、
1CHR|8|15|西巴第雅 、 亞拉得 、 亞得 、
1CHR|8|16|米迦勒 、 伊施巴 和 約哈 都是 比利亞 的兒子。
1CHR|8|17|西巴第雅 、 米書蘭 、 希西基 、 希伯 、
1CHR|8|18|伊施米萊 、 伊斯利亞 和 約巴 都是 以利巴力 的兒子。
1CHR|8|19|雅金 、 細基利 、 撒底 、
1CHR|8|20|以利乃 、 洗勒太 、 以利業 、
1CHR|8|21|亞大雅 、 比拉雅 和 申拉 都是 示每 的兒子。
1CHR|8|22|伊施班 、 希伯 、 以利業 、
1CHR|8|23|亞伯頓 、 細基利 、 哈難 、
1CHR|8|24|哈拿尼雅 、 以攔 、 安陀提雅 、
1CHR|8|25|伊弗底雅 、 毗努伊勒 都是 沙煞 的兒子。
1CHR|8|26|珊示萊 、 示哈利 、 亞他利雅 、
1CHR|8|27|雅利西 、 以利亞 和 細基利 都是 耶羅罕 的兒子。
1CHR|8|28|這些人按照他們的家譜都是族長，是領袖，都住在 耶路撒冷 。
1CHR|8|29|在 基遍 住的有 基遍 的父親 耶利 ，他的妻子名叫 瑪迦 ；
1CHR|8|30|他的長子是 亞伯頓 ，還有 蘇珥 、 基士 、 巴力 、 拿答 、
1CHR|8|31|基多 、 亞希約 和 撒迦 。
1CHR|8|32|米基羅 生 示米暗 。這些人在他們弟兄的對面，和他們的弟兄同住在 耶路撒冷 。
1CHR|8|33|尼珥 生 基士 ； 基士 生 掃羅 ； 掃羅 生 約拿單 、 麥基‧舒亞 、 亞比拿達 和 伊施巴力 。
1CHR|8|34|約拿單 的兒子是 米力‧巴力 ； 米力‧巴力 生 米迦 。
1CHR|8|35|米迦 的兒子是 毗敦 、 米勒 、 他利亞 和 亞哈斯 ；
1CHR|8|36|亞哈斯 生 耶何阿達 ； 耶何阿達 生 亞拉篾 、 亞斯瑪威 和 心利 ； 心利 生 摩撒 ；
1CHR|8|37|摩撒 生 比尼亞 ； 比尼亞 的兒子是 拉法 ， 拉法 的兒子是 以利亞薩 ， 以利亞薩 的兒子是 亞悉 。
1CHR|8|38|亞悉 有六個兒子，他們的名字是 亞斯利干 、 波基路 、 以實瑪利 、 示亞利雅 、 俄巴底雅 和 哈難 ；這些全都是 亞悉 的兒子。
1CHR|8|39|亞悉 兄弟 以設 的兒子：長子是 烏蘭 ，次子是 耶烏施 ，三子是 以利法列 。
1CHR|8|40|烏蘭 的兒子都是大能的勇士，是弓箭手，他們有許多的子孫，共一百五十名，都是 便雅憫 人。
1CHR|9|1|以色列 眾人按家譜登記，看哪，都寫在《以色列諸王記》上。 猶大 人因背叛被擄到 巴比倫 。
1CHR|9|2|從 巴比倫 先回來，住在自己地業城鎮中的有 以色列 人、祭司、 利未 人和殿役。
1CHR|9|3|住在 耶路撒冷 的有 猶大 人、 便雅憫 人、 以法蓮 人和 瑪拿西 人：
1CHR|9|4|猶大 兒子 法勒斯 的子孫中有 烏太 ， 烏太 是 亞米忽 的兒子， 亞米忽 是 暗利 的兒子， 暗利 是 音利 的兒子， 音利 是 巴尼 的兒子；
1CHR|9|5|示羅 人中有長子 亞帥雅 和他的眾兒子；
1CHR|9|6|謝拉 的子孫中有 耶烏利 和他的弟兄，共六百九十人；
1CHR|9|7|便雅憫 人中有 哈西努亞 的曾孫， 何達威雅 的孫子， 米書蘭 的兒子 撒路 ；
1CHR|9|8|又有 耶羅罕 的兒子 伊比內雅 ； 米基立 的孫子， 烏西 的兒子 以拉 ； 伊比尼雅 的曾孫， 流珥 的孫子， 示法提雅 的兒子 米書蘭 ；
1CHR|9|9|和他們的弟兄，按著家譜登記，共有九百五十六名；這些人都是族長。
1CHR|9|10|祭司中有 耶大雅 、 耶何雅立 、 雅斤 ，
1CHR|9|11|還有管理上帝殿的 亞撒利雅 ， 亞撒利雅 是 希勒家 的兒子， 希勒家 是 米書蘭 的兒子， 米書蘭 是 撒督 的兒子， 撒督 是 米拉約 的兒子， 米拉約 是 亞希突 的兒子。
1CHR|9|12|還有 瑪基雅 的曾孫， 巴施戶珥 的孫子， 耶羅罕 的兒子 亞大雅 ；又有 瑪賽 ， 瑪賽 是 亞第業 的兒子， 亞第業 是 雅希細拉 的兒子， 雅希細拉 是 米書蘭 的兒子， 米書蘭 是 米實利密 的兒子， 米實利密 是 音麥 的兒子。
1CHR|9|13|他們和他們的弟兄都是族長，共有一千七百六十人，都善於做上帝殿的事工。
1CHR|9|14|利未 人 米拉利 的子孫中有 哈沙比雅 的曾孫， 押利甘 的孫子， 哈述 的兒子 示瑪雅 ；
1CHR|9|15|有 拔巴甲 、 黑勒施 、 加拉 和 亞薩 的曾孫， 細基利 的孫子， 米迦 的兒子 瑪探雅 ；
1CHR|9|16|又有 耶杜頓 的曾孫， 加拉 的孫子， 示瑪雅 的兒子 俄巴底 ，還有 以利加拿 的孫子， 亞撒 的兒子 比利家 。他們都住在 尼陀法 人的村莊。
1CHR|9|17|守衛是 沙龍 、 亞谷 、 達們 、 亞希幔 和他們的弟兄； 沙龍 是領袖。
1CHR|9|18|從前這些人看守朝東的王門，如今是 利未 人營中的守衛。
1CHR|9|19|可拉 的曾孫， 以比雅撒 的孫子， 可利 的兒子 沙龍 ，和他父家的弟兄 可拉 人管理事務，看守會幕的門。他們的祖宗曾管理耶和華的軍營，把守營的入口。
1CHR|9|20|從前 以利亞撒 的兒子 非尼哈 管理他們，耶和華也與他同在。
1CHR|9|21|米施利米雅 的兒子 撒迦利雅 是看守會幕門口的。
1CHR|9|22|被選作門口守衛的總共有二百一十二名。他們在自己的村莊，按著家譜登記，是 大衛 和 撒母耳 先見所派擔當這受託之職任的。
1CHR|9|23|他們和他們的子孫看守耶和華殿的門，就是會幕的門口。
1CHR|9|24|在東西南北，四方 都有守衛。
1CHR|9|25|他們的弟兄住在村莊，每七日來與他們換班。
1CHR|9|26|這些守衛的四個領袖都是 利未 人，各有受託的職任，看守上帝殿的房間和寶庫。
1CHR|9|27|他們住在上帝殿的四圍，受託看守聖殿，負責每日早晨開門。
1CHR|9|28|利未 人中有人管理所使用的器皿，拿出拿入都按數目點算。
1CHR|9|29|又有人管理器具和聖所一切的器皿，以及細麵、酒、油、乳香和香料。
1CHR|9|30|祭司的子孫中有人用香料做膏油。
1CHR|9|31|利未 人 瑪他提雅 是 可拉 族 沙龍 的長子，他受託做烤餅。
1CHR|9|32|他們弟兄 哥轄 子孫中，有人負責每安息日排列供餅。
1CHR|9|33|歌唱的有 利未 人的族長，住在殿的房間，晝夜供職，不做別樣的工。
1CHR|9|34|以上都是 利未 人的族長，按各世系作領袖，他們都住在 耶路撒冷 。
1CHR|9|35|在 基遍 住的有 基遍 的父親 耶利 ，他的妻子名叫 瑪迦 ；
1CHR|9|36|他的長子是 亞伯頓 ，還有 蘇珥 、 基士 、 巴力 、 尼珥 、 拿答 、
1CHR|9|37|基多 、 亞希約 、 撒迦利雅 和 米基羅 。
1CHR|9|38|米基羅 生 示米暗 。這些人在他們弟兄的對面，和他們的弟兄同住在 耶路撒冷 。
1CHR|9|39|尼珥 生 基士 ； 基士 生 掃羅 ； 掃羅 生 約拿單 、 麥基‧舒亞 、 亞比拿達 和 伊施巴力 。
1CHR|9|40|約拿單 的兒子是 米力‧巴力 ； 米力‧巴力 生 米迦 。
1CHR|9|41|米迦 的兒子是 毗敦 、 米勒 、 他利亞 和 亞哈斯 。
1CHR|9|42|亞哈斯 生 雅拉 ； 雅拉 生 亞拉篾 、 亞斯瑪威 和 心利 ； 心利 生 摩撒 ；
1CHR|9|43|摩撒 生 比尼亞 ； 比尼亞 的兒子是 利法雅 ， 利法雅 的兒子是 以利亞薩 ， 以利亞薩 的兒子是 亞悉 。
1CHR|9|44|亞悉 有六個兒子，他們的名字是 亞斯利干 、 波基路 、 以實瑪利 、 示亞利雅 、 俄巴底雅 和 哈難 ；這些都是 亞悉 的兒子。
1CHR|10|1|非利士 人攻打 以色列 。 以色列 人在 非利士 人面前逃跑，很多人 在 基利波山 被殺仆倒。
1CHR|10|2|非利士 人緊追 掃羅 和他的兒子，殺了 掃羅 的兒子 約拿單 、 亞比拿達 、 麥基‧舒亞 。
1CHR|10|3|攻擊 掃羅 的戰事激烈， 掃羅 被弓箭手射中，被他們射傷。
1CHR|10|4|掃羅 吩咐拿他兵器的人說：「你拔出刀來，把我刺死，免得那些未受割禮的人來凌辱我。」但拿兵器的人非常懼怕，不肯刺他。於是 掃羅 拿起刀來，伏在刀上。
1CHR|10|5|拿兵器的人見 掃羅 已死，也伏在刀上死了。
1CHR|10|6|這樣， 掃羅 和他三個兒子，以及他的全家都一起陣亡了。
1CHR|10|7|住平原的 以色列 眾人見 以色列 軍兵 逃跑， 掃羅 和他兒子都死了，就棄城逃跑。 非利士 人前來，佔據了他們的城。
1CHR|10|8|次日， 非利士 人來剝那些被殺之人的衣服，看見 掃羅 和他兒子仆倒在 基利波山 。
1CHR|10|9|他們剝了他的軍裝，拿著他的首級和盔甲，派人到 非利士 人之地的四境，報信給他們的偶像和百姓。
1CHR|10|10|他們將 掃羅 的盔甲放在他們神明的廟裏，把他的首級釘在 大袞 廟中。
1CHR|10|11|基列 的 雅比 居民聽見 非利士 人向 掃羅 所行的一切事，
1CHR|10|12|他們中間所有的勇士就起身，把 掃羅 和他兒子的屍身送到 雅比 ，把他們的屍骨葬在 雅比 的橡樹下，禁食七日。
1CHR|10|13|這樣， 掃羅 為了他的不忠死了；因為他干犯耶和華，沒有遵守耶和華的話，又因他求問招魂的婦人，
1CHR|10|14|不求問耶和華，所以耶和華使他被殺，把王國給了 耶西 的兒子 大衛 。
1CHR|11|1|以色列 眾人聚集到 希伯崙 見 大衛 ，說：「看哪，我們是你的骨肉。
1CHR|11|2|從前 掃羅 作王的時候，率領 以色列 人出入的是你；耶和華－你的上帝也曾對你說：『你必牧養我的百姓 以色列 ，你必作我百姓 以色列 的君王。』」
1CHR|11|3|於是 以色列 的眾長老都來到 希伯崙 見王。 大衛 在 希伯崙 ，在耶和華面前與他們立約，他們就膏 大衛 作 以色列 的王，正如耶和華藉 撒母耳 所說的話。
1CHR|11|4|大衛 和 以色列 眾人到了 耶路撒冷 ，就是 耶布斯 ；那時 耶布斯 人住在那裏。
1CHR|11|5|耶布斯 人對 大衛 說：「你必不能進到這裏。」然而 大衛 攻取了 錫安 的堡壘，就是 大衛 的城。
1CHR|11|6|大衛 說：「誰先攻打 耶布斯 人，必作領袖，作元帥。」 洗魯雅 的兒子 約押 先上去，就作了領袖。
1CHR|11|7|大衛 住在堡壘裏，所以那堡壘叫作 大衛城 。
1CHR|11|8|大衛 又從 米羅 起，四圍建築城牆，其餘的由 約押 修建。
1CHR|11|9|大衛 日見強大，萬軍之耶和華與他同在。
1CHR|11|10|以下是跟隨 大衛 勇士的領袖；他們奮勇幫助他得到國度，並照著耶和華吩咐 以色列 的話，與 以色列 眾人一同立他作王。
1CHR|11|11|大衛 勇士的名單如下： 哈革摩尼 的兒子 雅朔班 ，他是軍官的統領 ，曾一次舉槍殺了三百人。
1CHR|11|12|其次是 亞何亞 人 朵多 的兒子 以利亞撒 ，他是三個勇士裏的一個。
1CHR|11|13|他從前與 大衛 在 巴斯‧大憫 ， 非利士 人聚集要打仗。那裏有一塊長滿大麥的田。百姓在 非利士 人面前逃跑，
1CHR|11|14|他們 卻站在那塊田的中間，防守那田，擊敗了 非利士 人。耶和華大獲全勝。
1CHR|11|15|三十個領袖中的三個人下到磐石那裏，進了 亞杜蘭洞 見 大衛 ； 非利士 的軍隊在 利乏音谷 安營。
1CHR|11|16|那時 大衛 在山寨， 非利士 人的駐軍在 伯利恆 。
1CHR|11|17|大衛 渴想著說：「但願有人從 伯利恆 城門旁的井裏打水來給我喝！」
1CHR|11|18|這三個勇士就闖過 非利士 人的軍營，從 伯利恆 城門旁的井裏打水，拿來給 大衛 喝。 大衛 卻不肯喝，將水澆在耶和華面前，
1CHR|11|19|說：「我的上帝啊，我絕不做這事！這些人冒死去打水，這水是他們用生命換來的，我怎能喝他們的血呢？」 大衛 不肯喝這水。這是三個勇士所做的事。
1CHR|11|20|約押 的兄弟 亞比篩 是這三個 勇士的領袖；他曾舉槍殺了三百人，就在三個勇士中得了名。
1CHR|11|21|他在這三個勇士裏比其他兩個更有名望，所以作他們的領袖，只是不及前三個勇士。
1CHR|11|22|耶何耶大 的兒子 比拿雅 是來自 甲薛 的勇士，曾行了大事。他殺了 摩押 人 亞利伊勒 的兩個兒子，又在下雪的時候下到坑裏去，殺了一隻獅子。
1CHR|11|23|他又殺了一個身高五肘的 埃及 人； 埃及 人手裏拿著槍，槍桿粗如織布機的軸。 比拿雅 只拿著棍子下到他那裏去，從 埃及 人手裏奪過槍來，用那槍殺死了他。
1CHR|11|24|這些是 耶何耶大 的兒子 比拿雅 所做的事，就在三個勇士裏得了名。
1CHR|11|25|看哪，他比那三十個勇士更有名望，只是不及前三個勇士。 大衛 立他作護衛長。
1CHR|11|26|軍中的勇士有 約押 的兄弟 亞撒黑 ， 伯利恆 人 朵多 的兒子 伊勒哈難 ，
1CHR|11|27|哈律 人 沙瑪 ， 比倫 人 希利斯 ，
1CHR|11|28|提哥亞 人 益吉 的兒子 以拉 ， 亞拿突 人 亞比以謝 ，
1CHR|11|29|戶沙 人 西比該 ， 亞何亞 人 以來 ，
1CHR|11|30|尼陀法 人 瑪哈萊 ， 尼陀法 人 巴拿 的兒子 希立 ，
1CHR|11|31|便雅憫 族 基比亞 人 利拜 的兒子 以太 ， 比拉頓 人 比拿雅 ，
1CHR|11|32|迦實溪 人 戶萊 ， 亞拉巴 人 亞比 ，
1CHR|11|33|巴路米 人 押斯瑪弗 ， 沙本 人 以利雅哈巴 ，
1CHR|11|34|基孫 人 哈深 的眾兒子， 哈拉 人 沙基 的兒子 約拿單 ，
1CHR|11|35|哈拉 人 沙甲 的兒子 亞希暗 ， 吾珥 的兒子 以利法勒 ，
1CHR|11|36|米基拉 人 希弗 ， 比倫 人 亞希雅 ，
1CHR|11|37|迦密 人 希斯羅 ， 伊斯拜 的兒子 拿萊 ，
1CHR|11|38|拿單 的兄弟 約珥 ， 哈基利 的兒子 彌伯哈 ，
1CHR|11|39|亞捫 人 洗勒 ， 比錄 人 拿哈萊 ，他是給 洗魯雅 的兒子 約押 拿兵器的，
1CHR|11|40|以帖 人 以拉 ， 以帖 人 迦立 ，
1CHR|11|41|赫 人 烏利亞 ， 亞萊 的兒子 撒拔 ，
1CHR|11|42|呂便 人 示撒 的兒子 亞第拿 ，是 呂便 支派中的一個領袖，率領三十人，
1CHR|11|43|瑪迦 的兒子 哈難 ， 彌特尼 人 約沙法 ，
1CHR|11|44|亞施他拉 人 烏西亞 ， 亞羅珥 人 何坦 的兒子 沙瑪 和 耶利 ，
1CHR|11|45|提洗 人 申利 的兒子 耶疊 和他的兄弟 約哈 ，
1CHR|11|46|瑪哈未 人 以利業 ， 伊利拿安 的兒子 耶利拜 和 約沙未雅 ， 摩押 人 伊特瑪 、
1CHR|11|47|以利業 、 俄備得 ，以及 米瑣八 人 雅西業 。
1CHR|12|1|以下是 大衛 因 基士 的兒子 掃羅 的緣故被放逐到 洗革拉 的時候，到他那裏幫助他打仗的勇士；
1CHR|12|2|他們是弓箭手，能左右甩石，開弓射箭，都是 便雅憫 人 掃羅 同族的弟兄：
1CHR|12|3|為首的是 亞希以謝 ，其次是 約阿施 ，都是 基比亞 人 示瑪 的兒子。還有 亞斯瑪威 的兒子 耶薛 和 毗力 ， 比拉迦 ， 亞拿突 人 耶戶 ，
1CHR|12|4|基遍 人 以實買雅 ，他在三十人中是勇士，管理這三十人，又有 耶利米 ， 雅哈悉 ， 約哈難 ， 基底拉 人 約撒拔 ，
1CHR|12|5|伊利烏賽 ， 耶利末 ， 比亞利雅 ， 示瑪利雅 ， 哈律弗 人 示法提雅 ，
1CHR|12|6|可拉 人 以利加拿 、 耶西亞 、 亞薩列 、 約以謝 、 雅朔班 ，
1CHR|12|7|基多 人 耶羅罕 的兒子 猶拉 和 西巴第雅 。
1CHR|12|8|迦得 人中有人到曠野的山寨投奔 大衛 ，都是大能的勇士，能拿盾牌和槍的戰士。他們的面貌好像獅子，敏捷如山上的鹿。
1CHR|12|9|第一 以薛 ，第二 俄巴底雅 ，第三 以利押 ，
1CHR|12|10|第四 彌施瑪拿 ，第五 耶利米 ，
1CHR|12|11|第六 亞太 ，第七 以利業 ，
1CHR|12|12|第八 約哈難 ，第九 以利薩巴 ，
1CHR|12|13|第十 耶利米 ，第十一 末巴奈 。
1CHR|12|14|這些都是 迦得 人中的軍官，小的能抵一百人，大的能抵一千人 。
1CHR|12|15|正月， 約旦河 水漲過兩岸的時候，他們過河，使所有住河谷的人東奔西逃。
1CHR|12|16|便雅憫 人和 猶大 人中有人來到山寨 大衛 那裏。
1CHR|12|17|大衛 出去迎接他們，回答他們說：「你們若和平地來幫助我，我的心就與你們契合；但你們若把我這雙手無辜的人賣給敵人，願我們列祖的上帝察看責罰。」
1CHR|12|18|那時軍官 的領袖 亞瑪撒 受靈的感動說： 「 大衛 啊，我們歸向你！ 耶西 的兒子啊，我們幫助你！ 願你平平安安， 願幫助你的也都平安！ 因為你的上帝幫助你。」 大衛 就收留他們，派他們作軍官。
1CHR|12|19|大衛 從前與 非利士 人同去，要與 掃羅 爭戰，有些 瑪拿西 人來投奔 大衛 。其實他們並沒有幫助 非利士 人，因為 非利士 人的領袖商議，打發他回去，說：「恐怕 大衛 拿我們的首級去向他的主人 掃羅 投誠。」
1CHR|12|20|大衛 往 洗革拉 去的時候，有 瑪拿西 人的千夫長 押拿 、 約撒拔 、 耶疊 、 米迦勒 、 約撒拔 、 以利戶 、 洗勒太 都來投奔他。
1CHR|12|21|他們幫助 大衛 攻擊敵軍；因為他們都是大能的勇士，又作軍官。
1CHR|12|22|那時天天有人來幫助 大衛 ，以致成了強大的軍隊，如上帝的軍隊一樣。
1CHR|12|23|以下是來到 希伯崙 見 大衛 ，要照耶和華的話把 掃羅 的國位歸給 大衛 的武裝士兵的數目：
1CHR|12|24|猶大 人，拿盾牌和槍的武裝戰士有六千八百人。
1CHR|12|25|西緬 人中，能上陣的大能勇士有七千一百人。
1CHR|12|26|利未 人中，有四千六百人。
1CHR|12|27|耶何耶大 是 亞倫 家的領袖，跟從他的有三千七百人。
1CHR|12|28|還有大能的青年勇士 撒督 ，同他本族的二十二個軍官。
1CHR|12|29|便雅憫 人中， 掃羅 同族的弟兄也有三千人；直到現在他們大部分仍然效忠 掃羅 家。
1CHR|12|30|以法蓮 人中，在本族中著名的大能勇士有二萬零八百人。
1CHR|12|31|瑪拿西 半支派，冊上有名來擁立 大衛 作王的，有一萬八千人。
1CHR|12|32|以薩迦 人中，通達時務，知道 以色列 所當行，同族弟兄也都聽從他們命令的族長有二百人。
1CHR|12|33|西布倫 中，能上陣用各樣作戰的兵器、不生二心幫助打仗的有五萬人。
1CHR|12|34|拿弗他利 中，有一千個軍官；跟從他們、拿盾牌和槍的有三萬七千人。
1CHR|12|35|但 人中，能擺陣的有二萬八千六百人。
1CHR|12|36|亞設 中，能上陣打仗的有四萬人。
1CHR|12|37|約旦河 東的 呂便 人、 迦得 人、 瑪拿西 半支派，拿各樣兵器打仗的有十二萬人。
1CHR|12|38|以上都是能列隊上陣的戰士，他們都全心來到 希伯崙 ，要擁立 大衛 作全 以色列 的王。 以色列 其餘的人也都一心要擁立 大衛 作王。
1CHR|12|39|他們在那裏三日，與 大衛 一同吃喝，因為他們同族的弟兄已經為他們預備好了。
1CHR|12|40|他們附近的人，以及 以薩迦 、 西布倫 、 拿弗他利 人，都將食物，許多麵餅、無花果餅、乾葡萄、酒、油，用驢、駱駝、騾子、牛馱來，又帶了許多的牛和羊來，因為在 以色列 中充滿了歡樂。
1CHR|13|1|大衛 與千夫長、百夫長，以及所有的領袖商議。
1CHR|13|2|大衛 對 以色列 全會眾說：「你們若以為好，見這事是出於耶和華－我們的上帝，我們就派人到遠近各處去見仍留在 以色列 各地我們的弟兄，以及住在有郊野之城的祭司和 利未 人，使他們都到我們這裏來聚集。
1CHR|13|3|我們要把上帝的約櫃接到這裏來；因為在 掃羅 年間，我們沒有去尋求約櫃 。」
1CHR|13|4|全會眾都說可以這麼做，因這事在眾百姓眼中都看為好。
1CHR|13|5|於是， 大衛 把 以色列 眾人從 埃及 的 西曷河 直到 哈馬口 都召集了來，要從 基列‧耶琳 將上帝的約櫃接來。
1CHR|13|6|大衛 率領 以色列 眾人上到 巴拉 ，就是屬 猶大 的 基列‧耶琳 ，要將耶和華上帝的約櫃從那裏接上來，他坐在二基路伯之上，這約櫃是以他的名來命名的。
1CHR|13|7|他們將上帝的約櫃從 亞比拿達 的家裏抬出來，放在新車上，由 烏撒 和 亞希約 趕車。
1CHR|13|8|大衛 和 以色列 眾人在上帝面前隨著詩歌、琴、瑟、鼓、鈸、號，極力跳舞。
1CHR|13|9|到了 基頓 的禾場，因為牛失前蹄 ， 烏撒 就伸手扶住約櫃。
1CHR|13|10|耶和華的怒氣向 烏撒 發作，因他伸手扶住約櫃而擊殺他，他就死在那裏，在上帝面前。
1CHR|13|11|大衛 因耶和華突然衝出撞死 烏撒 就生氣，稱那地方為 毗列斯‧烏撒 ，直到今日。
1CHR|13|12|那日， 大衛 懼怕上帝，說：「我怎能將上帝的約櫃接到我這裏來呢？」
1CHR|13|13|於是 大衛 不將約櫃接進 大衛城 他自己的地方，卻轉送到 迦特 人 俄別‧以東 的家中。
1CHR|13|14|上帝的約櫃停在 俄別‧以東 家中三個月，耶和華賜福給 俄別‧以東 的家和他一切所有的。
1CHR|14|1|推羅 王 希蘭 派使者把香柏木運到 大衛 那裏，又派石匠和木匠給 大衛 建造宮殿。
1CHR|14|2|大衛 知道耶和華堅立他作 以色列 王，又為自己百姓 以色列 的緣故，使他的國興盛。
1CHR|14|3|大衛 在 耶路撒冷 又立后妃，又生兒女。
1CHR|14|4|在 耶路撒冷 所生的孩子名字是 沙母亞 、 朔罷 、 拿單 、 所羅門 、
1CHR|14|5|益轄 、 以利書亞 、 以法列 、
1CHR|14|6|挪迦 、 尼斐 、 雅非亞 、
1CHR|14|7|以利沙瑪 、 比利雅大 、 以利法列 。
1CHR|14|8|非利士 人聽見 大衛 受膏作全 以色列 的王， 非利士 眾人就上來尋索 大衛 。 大衛 聽見了，就出去迎敵。
1CHR|14|9|非利士 人來了，侵犯 利乏音谷 。
1CHR|14|10|大衛 求問上帝說：「我可以上去攻打 非利士 人嗎？你將他們交在我手裏嗎？」耶和華對他說：「你可以上去，我必將他們交在你手裏。」
1CHR|14|11|非利士 人上到 巴力‧毗拉心 ， 大衛 在那裏擊敗他們。 大衛 說：「上帝藉我的手沖破敵人，如水沖破一樣。」因此那地方稱為 巴力‧毗拉心 。
1CHR|14|12|非利士 人把神像拋棄在那裏， 大衛 吩咐人用火焚燒了。
1CHR|14|13|非利士 人又侵犯 利乏音谷 。
1CHR|14|14|大衛 再求問上帝。上帝對他說：「不要從他們後頭追上去，要繞道離開他們，從桑樹林對面攻打他們。
1CHR|14|15|你聽見桑樹梢上有腳步的聲音，那時你就要出戰，因為上帝已經出去，在你前頭攻打 非利士 人的軍隊了。」
1CHR|14|16|大衛 就遵照上帝所吩咐的去做，攻打 非利士 人的軍隊，從 基遍 直到 基色 。
1CHR|14|17|於是 大衛 的名傳揚到萬邦，耶和華使萬國都懼怕他。
1CHR|15|1|大衛 在 大衛城 為自己建造宮殿，又為上帝的約櫃預備地方，支搭帳幕。
1CHR|15|2|那時 大衛 說：「除了 利未 人之外，無人可抬上帝的約櫃，因為耶和華揀選他們抬上帝的約櫃，永遠事奉他。」
1CHR|15|3|大衛 召集 以色列 眾人到 耶路撒冷 ，要將耶和華的約櫃接到他所預備的地方。
1CHR|15|4|大衛 又召集 亞倫 的子孫和 利未 人：
1CHR|15|5|哥轄 子孫中有領袖 烏列 和他的弟兄一百二十人，
1CHR|15|6|米拉利 子孫中有領袖 亞帥雅 和他的弟兄二百二十人，
1CHR|15|7|革順 子孫中有領袖 約珥 和他的弟兄一百三十人，
1CHR|15|8|以利撒反 子孫中有領袖 示瑪雅 和他的弟兄二百人，
1CHR|15|9|希伯倫 子孫中有領袖 以利業 和他的弟兄八十人，
1CHR|15|10|烏薛 子孫中有領袖 亞米拿達 和他的弟兄一百一十二人。
1CHR|15|11|大衛 召來 撒督 和 亞比亞他 二位祭司，以及 利未 人 烏列 、 亞帥雅 、 約珥 、 示瑪雅 、 以利業 、 亞米拿達 ，
1CHR|15|12|對他們說：「你們是 利未 人的族長，你們和你們的弟兄應當使自己分別為聖，好將耶和華－ 以色列 上帝的約櫃接到我所預備的地方。
1CHR|15|13|因為你們上一次沒有抬這約櫃，並且我們沒有按規矩求問耶和華－我們的上帝，所以他衝出來攻擊我們。」
1CHR|15|14|於是祭司和 利未 人使自己分別為聖，將耶和華－ 以色列 上帝的約櫃接上來。
1CHR|15|15|利未 子孫用槓，把上帝的約櫃抬在肩上，正如 摩西 按照耶和華的話所吩咐的。
1CHR|15|16|大衛 吩咐 利未 人的領袖派他們歌唱的弟兄用琴瑟和鈸的樂器奏樂，歡歡喜喜地大聲歌頌。
1CHR|15|17|於是 利未 人派 約珥 的兒子 希幔 和他弟兄中 比利家 的兒子 亞薩 ，以及他們同族弟兄 米拉利 子孫裏 古沙雅 的兒子 以探 。
1CHR|15|18|其次還有跟隨他們的弟兄 撒迦利雅 、 便‧雅薛 、 示米拉末 、 耶歇 、 烏尼 、 以利押 、 比拿雅 、 瑪西雅 、 瑪他提雅 、 以利斐利戶 、 彌克尼雅 ，以及門口的守衛 俄別‧以東 和 耶利 。
1CHR|15|19|歌唱的 希幔 、 亞薩 和 以探 ，敲銅鈸，聲音響亮；
1CHR|15|20|撒迦利雅 、 雅薛 、 示米拉末 、 耶歇 、 烏尼 、 以利押 、 瑪西雅 、 比拿雅 鼓瑟，調用女音；
1CHR|15|21|瑪他提雅 、 以利斐利戶 、 彌克尼雅 、 俄別‧以東 、 耶利 、 亞撒西雅 用琴指揮，調用第八。
1CHR|15|22|基拿尼雅 是 利未 人聖詠團的領袖，又教導人唱歌，因為他精通此事。
1CHR|15|23|比利家 和 以利加拿 是約櫃的守衛。
1CHR|15|24|示巴尼 、 約沙法 、 拿坦業 、 亞瑪賽 、 撒迦利雅 、 比拿亞 、 以利以謝 眾祭司在上帝的約櫃前吹號。 俄別‧以東 和 耶希亞 也是約櫃的守衛。
1CHR|15|25|於是， 大衛 和 以色列 的長老，以及千夫長都去，歡歡喜喜地將耶和華的約櫃從 俄別‧以東 家中接上來。
1CHR|15|26|上帝賜恩給抬耶和華約櫃的 利未 人，他們就獻上七頭公牛，七隻公羊。
1CHR|15|27|大衛 和所有抬約櫃的 利未 人，以及聖詠團的領袖 基拿尼雅 和歌唱的人，都穿著細麻布外袍； 大衛 另外穿著細麻布以弗得。
1CHR|15|28|這樣， 以色列 眾人歡呼、吹角、吹號、敲鈸、鼓瑟、彈琴，聲音響亮，將耶和華的約櫃接上來。
1CHR|15|29|耶和華的約櫃進 大衛城 的時候， 掃羅 的女兒 米甲 從窗戶裏往外觀看，見 大衛 王踴躍跳舞，心裏就輕視他。
1CHR|16|1|眾人將上帝的約櫃請進去，安放在 大衛 為它搭的帳幕中，就在上帝面前獻燔祭和平安祭。
1CHR|16|2|大衛 獻完了燔祭和平安祭，就奉耶和華的名祝福百姓，
1CHR|16|3|並且分給每一個 以色列 人，無論男女，每人一個餅，一個棗子餅 ，一個葡萄餅。
1CHR|16|4|大衛 派幾個 利未 人在耶和華的約櫃前事奉，頌揚，稱謝，讚美耶和華－ 以色列 的上帝：
1CHR|16|5|為首的是 亞薩 ，其次是 撒迦利雅 、 耶利 、 示米拉末 、 耶歇 、 瑪他提雅 、 以利押 、 比拿雅 、 俄別‧以東 、 耶利 ；他們鼓瑟彈琴， 亞薩 敲鈸，聲音響亮；
1CHR|16|6|比拿雅 和 雅哈悉 二位祭司常在上帝的約櫃前吹號。
1CHR|16|7|那日， 大衛 初次指派 亞薩 和他的弟兄稱謝耶和華。
1CHR|16|8|你們要稱謝耶和華，求告他的名， 在萬民中傳揚他的作為！
1CHR|16|9|要向他唱詩，向他歌頌， 述說他一切奇妙的作為！
1CHR|16|10|要誇耀他的聖名！ 願尋求耶和華的人心中歡喜！
1CHR|16|11|要尋求耶和華與他的能力， 時常尋求他的面。
1CHR|16|12|他僕人 以色列 的後裔， 他所揀選 雅各 的子孫哪， 要記念他奇妙的作為和他的奇事， 並他口中的判語。
1CHR|16|13|
1CHR|16|14|他是耶和華－我們的上帝， 全地都有他的判斷。
1CHR|16|15|要記念他的約，直到永遠； 記念他吩咐的話，直到千代，
1CHR|16|16|就是他與 亞伯拉罕 所立的約， 向 以撒 所起的誓。
1CHR|16|17|他將這約向 雅各 定為律例， 向 以色列 定為永遠的約，
1CHR|16|18|說：「我必將 迦南 地賜給你， 作你們應得的產業。」
1CHR|16|19|當時，你們人丁有限， 數目稀少，在那地寄居。
1CHR|16|20|他們從這邦遊到那邦， 從這國去到另一民族。
1CHR|16|21|他不容人欺負他們， 為他們的緣故責備君王：
1CHR|16|22|「不可傷害我的受膏者， 也不可惡待我的先知。」
1CHR|16|23|全地都要向耶和華歌唱！ 天天傳揚他的救恩！
1CHR|16|24|在列國中述說他的榮耀！ 在萬民中述說他的奇事！
1CHR|16|25|因耶和華本為大，當受極大的讚美； 他在萬神之上，當受敬畏。
1CHR|16|26|因萬民的神明都屬虛無； 惟獨耶和華創造諸天。
1CHR|16|27|有尊榮和威嚴在他面前， 有能力和喜樂在他自己的地方。
1CHR|16|28|民中的萬族啊，要將榮耀、能力歸給耶和華， 都歸給耶和華！
1CHR|16|29|要將耶和華的名所當得的榮耀歸給他， 拿供物來獻在他面前； 當敬拜神聖榮耀的耶和華 。
1CHR|16|30|全地都要在他面前戰抖！ 世界堅定，不得動搖。
1CHR|16|31|願天歡喜，願地快樂！ 願人在列國中說： 「耶和華作王了！」
1CHR|16|32|願海和其中所充滿的澎湃！ 願田和其中所有的都歡樂！
1CHR|16|33|那時，林中的樹木都要在耶和華面前歡呼， 因為他來要審判全地。
1CHR|16|34|你們要稱謝耶和華，因他本為善， 他的慈愛永遠長存！
1CHR|16|35|你們要說： 「拯救我們的上帝啊，求你拯救我們， 聚集我們，救我們脫離列國， 我們好頌揚你的聖名， 以讚美你為誇勝。
1CHR|16|36|耶和華－ 以色列 的上帝是應當稱頌的， 從亙古直到永遠。」 全體百姓都說：「阿們！」並且讚美耶和華。
1CHR|16|37|大衛 把 亞薩 和他的弟兄留在耶和華的約櫃那裏，經常在約櫃前事奉，天天盡本分供職，
1CHR|16|38|又有 俄別‧以東 和他的弟兄六十八人； 耶杜頓 的兒子 俄別‧以東 ，以及 何薩 作門口的守衛。
1CHR|16|39|還有 撒督 祭司和他弟兄眾祭司在 基遍 的丘壇、耶和華的帳幕前，
1CHR|16|40|在燔祭壇上，每日早晚，照著寫在耶和華律法書上所吩咐 以色列 的，經常獻燔祭給耶和華。
1CHR|16|41|與他們一同的還有 希幔 、 耶杜頓 ，和其餘被選、名字錄在冊上的，為要稱謝耶和華，因他的慈愛永遠長存。
1CHR|16|42|希幔 、 耶杜頓 同他們吹號、敲鈸，聲音響亮，並用其他樂器配合，歌頌上帝。 耶杜頓 的子孫作門口的守衛。
1CHR|16|43|於是眾百姓各自回家， 大衛 也回去為家人祝福。
1CHR|17|1|大衛 住在自己宮中，對 拿單 先知說：「看哪，我住在香柏木的宮中，耶和華的約櫃卻在幔子裏。」
1CHR|17|2|拿單 對 大衛 說：「你可以完全照你的心意去做，因為上帝與你同在。」
1CHR|17|3|當夜上帝的話臨到 拿單 ，說：
1CHR|17|4|「你去對我僕人 大衛 說：『耶和華如此說：你不可建造殿宇給我居住。
1CHR|17|5|自從我領 以色列 人上來，直到今日，我未曾住過殿宇；我從這會幕到那會幕，從這帳幕到那帳幕 。
1CHR|17|6|凡我同 以色列 人所走的地方，我何曾向 以色列 的一個士師，就是我吩咐牧養我百姓的，說過這話：你們為何不給我建造香柏木的殿宇呢？』
1CHR|17|7|現在，你要對我僕人 大衛 這樣說：『萬軍之耶和華如此說：我從羊圈中將你召來，叫你不再牧放羊群，立你作我百姓 以色列 的君王。
1CHR|17|8|你無論往哪裏去，我都與你同在，剪除你所有的仇敵。我必使你得大名，好像世上偉人的名一樣。
1CHR|17|9|我必為我百姓 以色列 選定一個地方，栽植他們，使他們住自己的地方，不再受攪擾；兇惡之子也不再像從前那樣擾亂他們，
1CHR|17|10|並不像我命令士師治理我百姓 以色列 的日子。我必制伏你所有的仇敵，並且我應許你 ，耶和華必為你建立家室。
1CHR|17|11|當你壽數滿足歸你祖先的時候，我必使你的後裔，你自己的兒子接續你；我也必堅定他的國。
1CHR|17|12|他必為我建造殿宇，我必堅定他的王位，直到永遠。
1CHR|17|13|我要作他的父，他要作我的子；我必不使我的慈愛離開他，像離開在你以前的那位一樣。
1CHR|17|14|我要永遠堅立他在我的家和我的國裏；他的王位也必堅定，直到永遠。』」
1CHR|17|15|拿單 就按這一切話，照這一切異象告訴 大衛 。
1CHR|17|16|於是 大衛 王進去，坐在耶和華面前，說：「耶和華上帝啊，我是誰，我的家算甚麼，你竟帶領我到這地步呢？
1CHR|17|17|上帝啊，這在你眼中還看為小，你又說到你僕人的家將來的情況。耶和華上帝啊，你看顧我好像看顧尊貴的人。
1CHR|17|18|你加於僕人的尊榮， 大衛 還有甚麼可以對你說呢？你是知道你僕人的。
1CHR|17|19|耶和華啊，因你僕人的緣故，也照著你的心意，你行這一切大事，為了顯明這一切偉大的事。
1CHR|17|20|耶和華啊，照我們耳中一切所聽見的，沒有可比你的，除你以外再沒有上帝。
1CHR|17|21|世上有何國能比你的百姓 以色列 呢？上帝親自去救贖世上的一國 ，作自己的子民，又行大而可畏的事，顯出你的大名，在你從 埃及 贖出來的子民面前驅逐了列國。
1CHR|17|22|你使你的百姓 以色列 作你的子民，直到永遠；你－耶和華也作他們的上帝。
1CHR|17|23|現在，耶和華啊，你所應許僕人和僕人家的話，求你堅定，直到永遠；求你照你所說的而行。
1CHR|17|24|願你的名永遠堅立，被尊為大，人要說：『萬軍之耶和華－ 以色列 的上帝，是 以色列 的上帝。』這樣，你僕人 大衛 的家必在你面前堅立。
1CHR|17|25|我的上帝啊，因你啟示你的僕人，要為他建立家室，所以僕人大膽在你面前祈禱。
1CHR|17|26|現在，耶和華啊，惟有你是上帝！你應許將這福氣賜給僕人。
1CHR|17|27|現在，你喜悅賜福給僕人的家，可以永存在你面前。耶和華啊，因你已經賜福，還要賜福到永遠。」
1CHR|18|1|此後， 大衛 攻打 非利士 人，制伏了他們，從 非利士 人手中奪取了 迦特 和所屬的鄉鎮。
1CHR|18|2|他又攻打 摩押 ， 摩押 人就臣服 大衛 ，向他進貢。
1CHR|18|3|瑣巴 王 哈大底謝 往 幼發拉底河 去，要鞏固自己的國權。 大衛 攻打他，直到 哈馬 ，
1CHR|18|4|奪了他的戰車一千，俘擄了騎兵七千人，步兵二萬人。 大衛 把所有戰馬的蹄筋砍斷，只留下一百輛戰車。
1CHR|18|5|大馬士革 的 亞蘭 人來幫助 瑣巴 王 哈大底謝 ， 大衛 殺了 亞蘭 人二萬二千。
1CHR|18|6|於是 大衛 在 大馬士革 的 亞蘭 地設立軍營 ， 亞蘭 人就臣服 大衛 ，向他進貢。 大衛 無論往哪裏去，耶和華都使他得勝。
1CHR|18|7|大衛 奪了 哈大底謝 臣僕擁有的金盾牌，帶到 耶路撒冷 。
1CHR|18|8|大衛 又從 哈大底謝 的 提巴 和 均 二城奪取了許多的銅；後來 所羅門 用這些銅製造銅海、銅柱和銅器。
1CHR|18|9|哈馬 王 陀烏 聽見 大衛 擊敗 瑣巴 王 哈大底謝 的全軍，
1CHR|18|10|就派他兒子 哈多蘭 到 大衛 王那裏，向他請安，為他祝福，因他與 哈大底謝 爭戰，並且擊敗了他；原來 哈大底謝 與 陀烏 常常爭戰。 哈多蘭 帶了金銀銅的各樣器皿來。
1CHR|18|11|大衛 王把這些器皿，以及從各國奪來的金銀，就是從 以東 、 摩押 、 亞捫 人、 非利士 人、 亞瑪力 所奪來的，都分別為聖獻給耶和華。
1CHR|18|12|洗魯雅 的兒子 亞比篩 在 鹽谷 擊殺了一萬八千 以東 人。
1CHR|18|13|大衛 在 以東 設立軍營， 以東 人就都臣服他。 大衛 無論往哪裏去，耶和華都使他得勝。
1CHR|18|14|大衛 作全 以色列 的王，又向眾百姓秉公行義。
1CHR|18|15|洗魯雅 的兒子 約押 作元帥； 亞希律 的兒子 約沙法 作史官；
1CHR|18|16|亞希突 的兒子 撒督 和 亞比亞他 的兒子 亞希米勒 作祭司； 沙威沙 作書記；
1CHR|18|17|耶何耶大 的兒子 比拿雅 管轄 基利提 人和 比利提 人。 大衛 的眾兒子都在王的左右作領袖。
1CHR|19|1|此後， 亞捫 人的王 拿轄 死了，他兒子接續他作王。
1CHR|19|2|大衛 說：「 哈嫩 的父親 拿轄 怎樣向我施恩，我也要怎樣向 哈嫩 施恩。」於是 大衛 派使者為他的父親安慰他。 大衛 的臣僕到了 亞捫 人的境內來見 哈嫩 ，要安慰他。
1CHR|19|3|但 亞捫 人的領袖對 哈嫩 說：「 大衛 派人來安慰你，你看他是要尊敬你父親嗎？他的臣僕來見你，不是為了要窺探偵察，而傾覆這地嗎？」
1CHR|19|4|哈嫩 就抓住 大衛 的臣僕，剃去他們的鬍鬚，又割斷他們下半截的衣服，露出臀部，然後放了他們。
1CHR|19|5|他們走了，有人把臣僕所遭遇的事告訴 大衛 ，他就派人去迎接他們，因為這些人覺得很羞恥。王說：「可以住在 耶利哥 ，等到鬍鬚長出來再回來。」
1CHR|19|6|亞捫 人看到 大衛 憎惡他們， 哈嫩 和 亞捫 人就派人拿一千他連得銀子，從 美索不達米亞 、 亞蘭‧瑪迦 、 瑣巴 雇用戰車和騎兵。
1CHR|19|7|他們雇了三萬二千輛戰車，以及 瑪迦 王和他的軍兵；這些部隊來安營在 米底巴 前。 亞捫 人也從他們的城裏出來，聚集預備作戰。
1CHR|19|8|大衛 聽見了，就派 約押 和所有勇猛的軍隊出去。
1CHR|19|9|亞捫 人出來，在城門前擺陣，前來的諸王另在郊野擺陣。
1CHR|19|10|約押 看見戰陣對著他前後擺列，就把從 以色列 所有精兵中挑選出來的，擺陣迎戰 亞蘭 人。
1CHR|19|11|他把其餘的兵交在他兄弟 亞比篩 手裏，他們就擺陣迎戰 亞捫 人。
1CHR|19|12|約押 說：「 亞蘭 人若強過我，你就來幫助我； 亞捫 人若強過你，我就去幫助你。
1CHR|19|13|你要剛強，我們要為自己的百姓，為我們上帝的城鎮奮勇。願耶和華照他所看為好的去做！」
1CHR|19|14|於是， 約押 和跟隨他的士兵前進攻打 亞蘭 人； 亞蘭 人在他面前逃跑。
1CHR|19|15|亞捫 人見 亞蘭 人逃跑，他們也在 約押 的兄弟 亞比篩 面前逃跑進城。 約押 就回 耶路撒冷 去了。
1CHR|19|16|亞蘭 人見自己被 以色列 打敗，就派使者把 大河 那邊的 亞蘭 人調來，由 哈大底謝 的將軍 朔法 在他們前面率領。
1CHR|19|17|有人告訴 大衛 ，他就聚集 以色列 眾人過 約旦河 ，來到 亞蘭 人那裏，迎著他們擺陣。 大衛 擺陣攻擊 亞蘭 人， 亞蘭 人就與他打仗。
1CHR|19|18|亞蘭 人在 以色列 人面前逃跑。 大衛 殺了 亞蘭 七千輛戰車的士兵，四萬步兵，又殺死 亞蘭 的將軍 朔法 。
1CHR|19|19|哈大底謝 的臣僕見自己被 以色列 打敗，就與 大衛 講和，臣服他。於是 亞蘭 人不願再幫助 亞捫 人了。
1CHR|20|1|到了年初，諸王出征的時候， 約押 率領軍兵蹂躪 亞捫 人的地，前來圍攻 拉巴 ； 大衛 仍住在 耶路撒冷 。 約押 攻打 拉巴 ，把它毀壞。
1CHR|20|2|大衛 奪了 米勒公 所戴的冠冕，其上的金子重一他連得，又嵌著寶石。這冠冕就戴在 大衛 頭上。 大衛 又從城裏奪了許多財物，
1CHR|20|3|把城裏的百姓拉出來，放在鋸下，或鐵耙下，或斧 的下面； 大衛 待 亞捫 各城的居民都是如此。於是， 大衛 和全軍都回 耶路撒冷 去了。
1CHR|20|4|後來， 以色列 人在 基色 與 非利士 人打仗。 戶沙 人 西比該 殺了巨人族的後裔 細派 ， 非利士 人就被制伏了。
1CHR|20|5|他們又與 非利士 人打仗。 睚珥 的兒子 伊勒哈難 殺了 迦特 人 歌利亞 的兄弟 拉哈米 ；這人的槍桿粗如織布機的軸。
1CHR|20|6|又有一次，他們在 迦特 打仗。那裏有一個身材高大的人，手指腳趾都是六根，共有二十四根；他也是巨人族的後裔。
1CHR|20|7|他向 以色列 罵陣， 大衛 的哥哥 示米亞 的兒子 約拿單 就殺了他。
1CHR|20|8|這些人是 迦特 巨人族的後裔，都仆倒在 大衛 和他僕人的手下。
1CHR|21|1|撒但起來攻擊 以色列 ，激起 大衛 數點以色列人。
1CHR|21|2|大衛 對 約押 和百姓的領袖說：「去，數點 以色列 人，從 別是巴 直到 但 ，回來告訴我，我好知道他們的數目。」
1CHR|21|3|約押 說：「願耶和華使他的百姓比現在加增百倍。我主我王啊，他們不都是我主的僕人嗎？我主為何吩咐行這事，為何使 以色列 陷入罪裏呢？」
1CHR|21|4|但王堅持他對 約押 的命令。 約押 就出去，來回走遍 以色列 ，然後回到 耶路撒冷 。
1CHR|21|5|約押 向 大衛 報告百姓的總數：全 以色列 拿刀的有一百一十萬人； 猶大 拿刀的有四十七萬人。
1CHR|21|6|惟有 利未 人和 便雅憫 人沒有算在其中，因為 約押 厭惡王的這命令。
1CHR|21|7|這件事在上帝眼中看為惡，上帝就降災給 以色列 。
1CHR|21|8|大衛 對上帝說：「我做這事大大有罪了。現在求你除掉僕人的罪孽，因為我所做的非常愚昧。」
1CHR|21|9|耶和華吩咐 迦得 ， 大衛 的先見，說：
1CHR|21|10|「你去告訴 大衛 說：『耶和華如此說：我列出三樣災禍給你，隨你選擇一樣，我好降與你。』」
1CHR|21|11|於是， 迦得 來到 大衛 那裏，對他說：「耶和華如此說：『你可以隨意選擇：
1CHR|21|12|三年的饑荒，或敗在敵人面前，被敵人的刀追殺三個月，或在國中三日有耶和華的刀，就是瘟疫，讓耶和華的使者在 以色列 全境施行毀滅呢？』現在你要想一想，我怎樣去回覆那差我來的。」
1CHR|21|13|大衛 對 迦得 說：「我很為難。我寧願落在耶和華的手裏，因為他有豐盛的憐憫；我不願落在人的手裏。」
1CHR|21|14|於是，耶和華降瘟疫給 以色列 ， 以色列 中死了七萬人。
1CHR|21|15|上帝派遣使者去毀滅 耶路撒冷 ，剛要毀滅的時候，耶和華看見就改變心意，不降這災了。他吩咐那滅城的天使說：「夠了，住手吧！」耶和華的使者正站在 耶布斯 人 阿珥楠 的禾場那裏。
1CHR|21|16|大衛 舉目，看見耶和華的使者站在天和地之間，手裏有拔出來的刀，伸在 耶路撒冷 以上。 大衛 和長老都披上麻布，臉伏於地。
1CHR|21|17|大衛 向上帝說：「吩咐數點百姓的不是我嗎？是我犯了罪，行了大惡，但這群羊做了甚麼呢？耶和華－我的上帝啊，願你的手攻擊我和我的父家，不要降瘟疫給你的百姓。」
1CHR|21|18|耶和華的使者吩咐 迦得 去告訴 大衛 ，叫他上去，在 耶布斯 人 阿珥楠 的禾場上為耶和華立一座壇。
1CHR|21|19|大衛 就照著 迦得 奉耶和華名所說的話上去。
1CHR|21|20|阿珥楠 回頭看見天使，跟他在一起的四個兒子都藏起來了， 阿珥楠 繼續打麥子。
1CHR|21|21|大衛 到了 阿珥楠 那裏， 阿珥楠 觀看，看見 大衛 ，就從禾場上出去，臉伏於地，向他下拜。
1CHR|21|22|大衛 對 阿珥楠 說：「你把這禾場的地方給我，照著十足的價錢賣給我，我好在其上為耶和華築一座壇，使瘟疫在百姓中停止。」
1CHR|21|23|阿珥楠 對 大衛 說：「請用這禾場吧，願我主我王照你眼中看為好的去做。看，我提供牛作燔祭，打糧的器具作柴，麥子作素祭，這一切我全都提供。」
1CHR|21|24|大衛 王對 阿珥楠 說：「不，我一定要按十足的價錢買；因我不能用你的東西獻給耶和華，也不能用白得之物獻為燔祭。」
1CHR|21|25|於是 大衛 為那個地方付了六百舍客勒重的金子給 阿珥楠 。
1CHR|21|26|大衛 在那裏為耶和華築了一座壇，獻燔祭和平安祭，求告耶和華。耶和華就應允他，使火從天降在燔祭壇上。
1CHR|21|27|耶和華吩咐使者，他就收刀入鞘。
1CHR|21|28|那時， 大衛 見耶和華在 耶布斯 人 阿珥楠 的禾場上應允了他，就在那裏獻祭。
1CHR|21|29|摩西 在曠野所造之耶和華的帳幕和燔祭壇，當時都在 基遍 的丘壇，
1CHR|21|30|只是 大衛 不能前去求問上帝，因為他懼怕耶和華使者的刀。
1CHR|22|1|大衛 說：「這是耶和華上帝的殿，這是 以色列 獻燔祭的壇。」
1CHR|22|2|大衛 吩咐人召集住 以色列 地的寄居者，又派石匠鑿石頭，要建造上帝的殿。
1CHR|22|3|大衛 預備許多鐵，要做門上的釘子和鉤子，又預備許多銅，多得無法可秤；
1CHR|22|4|還有無數的香柏木，因為 西頓 人和 推羅 人給 大衛 運了許多香柏木來。
1CHR|22|5|大衛 說：「我兒子 所羅門 還年幼脆弱，要為耶和華建造的殿宇必須高大輝煌，使名聲榮耀傳遍萬國，所以我要為殿預備。」於是， 大衛 在未死之前預備了許多材料。
1CHR|22|6|大衛 召了他兒子 所羅門 來，吩咐他為耶和華－ 以色列 的上帝建造殿宇。
1CHR|22|7|大衛 對 所羅門 說：「我兒啊，我心裏本想為耶和華－我上帝的名建造殿宇，
1CHR|22|8|可是耶和華的話臨到我說：『你流了許多的血，打了多次大仗；你不可為我的名建造殿宇，因為你在我面前使許多血流在地上。
1CHR|22|9|看哪，你要生一個兒子，他必成為安寧的人；我必使他得享安寧，不被四圍仇敵擾亂。他的名字要叫 所羅門 ，在他的日子，我必使 以色列 平安康泰。
1CHR|22|10|他必為我的名建造殿宇。他要作我的子，我要作他的父。我必堅定他國度的王位，使他治理 以色列 ，直到永遠。』
1CHR|22|11|我兒啊，現今願耶和華與你同在，使你亨通，建造耶和華－你上帝的殿，正如他指著你所說的。
1CHR|22|12|但願耶和華賜你聰明智慧，好按著他吩咐你的去治理 以色列 ，遵行耶和華－你上帝的律法。
1CHR|22|13|那時候，你若謹守遵行耶和華藉 摩西 吩咐 以色列 的律例典章，就得亨通。你當剛強壯膽，不要懼怕，也不要驚惶。
1CHR|22|14|看哪，我辛苦地為耶和華的殿預備了十萬他連得金子，一百萬他連得銀子，銅和鐵多得無法可秤；我也預備了木頭、石頭，你還可以增添。
1CHR|22|15|你有許多工匠，就是石匠、木匠，和一切能做各樣工的巧匠，
1CHR|22|16|以及無數的金銀銅鐵。你當起來做工，願耶和華與你同在。」
1CHR|22|17|大衛 又吩咐 以色列 的眾官長幫助他兒子 所羅門 ：
1CHR|22|18|「耶和華－你們的上帝不是與你們同在嗎？他不是使你們四圍都平安嗎？因他已將這地的居民交在我手中，這地已在耶和華與他百姓面前制伏了。
1CHR|22|19|現在你們應當立定心意，尋求耶和華－你們的上帝。你們當起來建造耶和華上帝的聖所，好將耶和華的約櫃和上帝神聖的器皿都搬進為耶和華的名建造的殿裏。」
1CHR|23|1|大衛 年紀老邁，日子滿足，就立他兒子 所羅門 作 以色列 的王。
1CHR|23|2|大衛 召集 以色列 的眾領袖、祭司和 利未 人。
1CHR|23|3|利未 人三十歲以上的都被數點，他們男丁的數目共有三萬八千；
1CHR|23|4|其中有二萬四千人管理耶和華殿的事務，有六千人作官長和審判官，
1CHR|23|5|有四千人作門口的守衛，又有四千人頌讚耶和華，用 大衛 造的樂器來頌讚。
1CHR|23|6|大衛 把 利未 人 革順 、 哥轄 、 米拉利 的子孫分了班次。
1CHR|23|7|屬 革順 的有 拉但 和 示每 。
1CHR|23|8|拉但 的長子是 耶歇 ，還有 西坦 和 約珥 ，共三人。
1CHR|23|9|示每 的兒子是 示羅密 、 哈薛 、 哈蘭 三人。這是 拉但 族的族長。
1CHR|23|10|示每 的兒子是 雅哈 、 細拿 、 耶烏施 、 比利亞 ，這四人是 示每 的兒子。
1CHR|23|11|雅哈 是長子， 細撒 是次子。但 耶烏施 和 比利亞 的子孫不多，所以算為一族。
1CHR|23|12|哥轄 的兒子是 暗蘭 、 以斯哈 、 希伯倫 、 烏薛 ，共四人。
1CHR|23|13|暗蘭 的兒子是 亞倫 和 摩西 。 亞倫 被分別出來，把至聖之物分別為聖，使他和他的子孫在耶和華面前燒香、事奉他，奉他的名祝福，直到永遠。
1CHR|23|14|至於神人 摩西 ，他的子孫記名在 利未 支派下。
1CHR|23|15|摩西 的兒子是 革舜 和 以利以謝 。
1CHR|23|16|革舜 的兒子，長子是 細布業 ；
1CHR|23|17|以利以謝 的兒子，長子是 利哈比雅 。 以利以謝 沒有別的兒子，但 利哈比雅 的子孫很多。
1CHR|23|18|以斯哈 的兒子，長子是 示羅密 。
1CHR|23|19|希伯倫 的兒子，長子是 耶利雅 ，次子是 亞瑪利亞 ，三子是 雅哈悉 ，四子是 耶加面 。
1CHR|23|20|烏薛 的兒子，長子是 米迦 ，次子是 耶西雅 。
1CHR|23|21|米拉利 的兒子是 抹利 和 母示 。 抹利 的兒子是 以利亞撒 和 基士 。
1CHR|23|22|以利亞撒 死了，沒有兒子，只有女兒，他們本族 基士 的幾個兒子娶了她們為妻。
1CHR|23|23|母示 的兒子是 末力 、 以得 、 耶列末 ，共三人。
1CHR|23|24|以上是 利未 子孫作族長的，按著父系、照著男丁的數目，二十歲以上登記的，都辦理耶和華殿的事務。
1CHR|23|25|大衛 說：「耶和華－ 以色列 的上帝已經使他的百姓得享安寧，他永遠住在 耶路撒冷 。
1CHR|23|26|因此， 利未 人不必再抬帳幕和其中所使用的一切器皿了。」
1CHR|23|27|照著 大衛 臨終的話， 利未 人二十歲以上的都被數點。
1CHR|23|28|他們的職務是作 亞倫 子孫的幫手，在耶和華的殿事奉，照管院子和屋子，潔淨一切聖物，辦理上帝殿的事務。
1CHR|23|29|他們負責預備供餅、素祭的細麵和無酵薄餅，或用盤烤，或用油調和的祭物，確認其數量和大小。
1CHR|23|30|每日早晚、安息日、初一，以及節期，按數照例，經常獻燔祭給耶和華的時候，他們站立稱謝讚美耶和華。
1CHR|23|31|
1CHR|23|32|他們照管會幕和聖所，服事他們的弟兄 亞倫 的子孫，辦理耶和華殿的事務。
1CHR|24|1|亞倫 子孫的班次如下： 亞倫 的兒子是 拿答 、 亞比戶 、 以利亞撒 、 以他瑪 。
1CHR|24|2|拿答 和 亞比戶 死在他們父親之先，沒有留下兒子；因此， 以利亞撒 和 以他瑪 擔任祭司的職分。
1CHR|24|3|大衛 和 以利亞撒 的子孫 撒督 ，以及 以他瑪 的子孫 亞希米勒 ，把他們按照任務分成班次，
1CHR|24|4|發現 以利亞撒 子孫中作領袖的，比 以他瑪 子孫中作領袖的更多，就分班如下： 以利亞撒 的子孫中有十六個族長， 以他瑪 的子孫中有八個族長。
1CHR|24|5|他們抽籤分配，彼此一樣。在聖所和上帝面前作領袖的有 以利亞撒 的子孫，也有 以他瑪 的子孫。
1CHR|24|6|作書記的 利未 人 拿坦業 的兒子 示瑪雅 在王和領袖，與 撒督 祭司、 亞比亞他 的兒子 亞希米勒 ，以及祭司和 利未 人的族長面前記錄他們的名字；在 以利亞撒 的子孫中取一族，在 以他瑪 的子孫中也取一族。
1CHR|24|7|抽籤的時候，第一籤抽到的是 耶何雅立 ，第二是 耶大雅 ，
1CHR|24|8|第三是 哈琳 ，第四是 梭琳 ，
1CHR|24|9|第五是 瑪基雅 ，第六是 米雅民 ，
1CHR|24|10|第七是 哈歌斯 ，第八是 亞比雅 ，
1CHR|24|11|第九是 耶書亞 ，第十是 示迦尼 ，
1CHR|24|12|第十一是 以利亞實 ，第十二是 雅金 ，
1CHR|24|13|第十三是 胡巴 ，第十四是 耶是比押 ，
1CHR|24|14|第十五是 璧迦 ，第十六是 音麥 ，
1CHR|24|15|第十七是 希悉 ，第十八是 哈闢悉 ，
1CHR|24|16|第十九是 毗他希雅 ，第二十是 以西結 ，
1CHR|24|17|第二十一是 雅斤 ，第二十二是 迦末 ，
1CHR|24|18|第二十三是 第來雅 ，第二十四是 瑪西亞 。
1CHR|24|19|這就是他們事奉的班次，要照耶和華－ 以色列 的上帝藉他們祖宗 亞倫 所吩咐的條例，進入耶和華的殿辦理事務。
1CHR|24|20|利未 其餘的子孫如下： 暗蘭 的子孫中有 書巴業 ； 書巴業 的子孫中有 耶希底亞 。
1CHR|24|21|屬 利哈比雅 ， 利哈比雅 的兒子中有長子 伊示雅 。
1CHR|24|22|屬 以斯哈 人的有 示羅摩 ； 示羅摩 的子孫中有 雅哈 。
1CHR|24|23|希伯倫 的兒子中有長子 耶利雅 ，次子 亞瑪利亞 ，三子 雅哈悉 ，四子 耶加面 。
1CHR|24|24|烏薛 的子孫中有 米迦 ； 米迦 的子孫中有 沙密 。
1CHR|24|25|米迦 的兄弟是 伊示雅 ； 伊示雅 的子孫中有 撒迦利雅 。
1CHR|24|26|米拉利 的兒子是 抹利 和 母示 ； 雅西雅 的子孫中有 比挪 ；
1CHR|24|27|米拉利 的子孫中有屬 雅西雅 的 比挪 、 朔含 、 撒刻 、 伊比利 。
1CHR|24|28|屬 抹利 的有 以利亞撒 ； 以利亞撒 沒有兒子。
1CHR|24|29|屬 基士 ， 基士 的子孫中有 耶拉篾 。
1CHR|24|30|母示 的兒子是 末力 、 以得 、 耶利末 。按著宗族，這些都是 利未 的子孫。
1CHR|24|31|他們在 大衛 王和 撒督 ，以及 亞希米勒 與祭司和 利未 人的族長面前也抽籤，正如他們弟兄 亞倫 的子孫一樣。各族的族長與最年輕的兄弟都一樣。
1CHR|25|1|大衛 和事奉團隊的眾領袖分派 亞薩 、 希幔 ，以及 耶杜頓 的子孫唱歌 ，以彈琴、鼓瑟、敲鈸伴奏。他們供職的人數如下：
1CHR|25|2|亞薩 的兒子 撒刻 、 約瑟 、 尼探雅 、 亞薩利拉 ， 亞薩 的兒子都在 亞薩 的指導下，遵王的指示唱歌。
1CHR|25|3|屬 耶杜頓 ， 耶杜頓 的兒子 基大利 、 西利 、 耶篩亞 、 示每 、 哈沙比雅 、 瑪他提雅 共六人，都在他們父親 耶杜頓 的指導下唱歌，以彈琴伴奏，稱謝，頌讚耶和華。
1CHR|25|4|屬 希幔 ， 希幔 的兒子是 布基雅 、 瑪探雅 、 烏薛 、 細布業 、 耶利末 、 哈拿尼雅 、 哈拿尼 、 以利亞他 、 基大利提 、 羅幔提‧以謝 、 約施比加沙 、 瑪羅提 、 何提 、 瑪哈秀 。
1CHR|25|5|這些都是 希幔 的兒子； 希幔 奉上帝之命作王的先見，吹角頌讚。上帝賜給 希幔 十四個兒子，三個女兒，
1CHR|25|6|他們都在父親的指導下，在耶和華的殿唱歌，以敲鈸、彈琴、鼓瑟伴奏，遵從王的指示，在上帝的殿裏事奉。 亞薩 、 耶杜頓 、 希幔 ，
1CHR|25|7|他們和他們的弟兄學習頌讚耶和華，精通者的數目共有二百八十八人。
1CHR|25|8|這些人無論大小，為師的、為徒的，都一同抽籤分了班次。
1CHR|25|9|抽籤的時候，第一籤抽到的是 亞薩 的兒子 約瑟 。第二是 基大利 ；他和他兄弟，以及兒子共十二人。
1CHR|25|10|第三是 撒刻 ，他兒子和他兄弟共十二人。
1CHR|25|11|第四是 伊洗利 ，他兒子和他兄弟共十二人。
1CHR|25|12|第五是 尼探雅 ，他兒子和他兄弟共十二人。
1CHR|25|13|第六是 布基雅 ，他兒子和他兄弟共十二人。
1CHR|25|14|第七是 耶薩利拉 ，他兒子和他兄弟共十二人。
1CHR|25|15|第八是 耶篩亞 ，他兒子和他兄弟共十二人。
1CHR|25|16|第九是 瑪探雅 ，他兒子和他兄弟共十二人。
1CHR|25|17|第十是 示每 ，他兒子和他兄弟共十二人。
1CHR|25|18|第十一是 亞薩烈 ，他兒子和他兄弟共十二人。
1CHR|25|19|第十二是 哈沙比雅 ，他兒子和他兄弟共十二人。
1CHR|25|20|第十三是 書巴業 ，他兒子和他兄弟共十二人。
1CHR|25|21|第十四是 瑪他提雅 ，他兒子和他兄弟共十二人。
1CHR|25|22|第十五是 耶列末 ，他兒子和他兄弟共十二人。
1CHR|25|23|第十六是 哈拿尼雅 ，他兒子和他兄弟共十二人。
1CHR|25|24|第十七是 約施比加沙 ，他兒子和他兄弟共十二人。
1CHR|25|25|第十八是 哈拿尼 ，他兒子和他兄弟共十二人。
1CHR|25|26|第十九是 瑪羅提 ，他兒子和他兄弟共十二人。
1CHR|25|27|第二十是 以利亞他 ，他兒子和他兄弟共十二人。
1CHR|25|28|第二十一是 何提 ，他兒子和他兄弟共十二人。
1CHR|25|29|第二十二是 基大利提 ，他兒子和他兄弟共十二人。
1CHR|25|30|第二十三是 瑪哈秀 ，他兒子和他兄弟共十二人。
1CHR|25|31|第二十四是 羅幔提‧以謝 ，他兒子和他兄弟共十二人。
1CHR|26|1|門口守衛的班次如下： 可拉 族 以比雅撒 的子孫中，有 可利 的兒子 米施利米雅 。
1CHR|26|2|米施利米雅 的長子是 撒迦利亞 ，次子是 耶疊 ，三子是 西巴第雅 ，四子是 耶提聶 ，
1CHR|26|3|五子是 以攔 ，六子是 約哈難 ，七子是 以利約乃 。
1CHR|26|4|俄別‧以東 的長子是 示瑪雅 ，次子是 約薩拔 ，三子是 約亞 ，四子是 沙甲 ，五子是 拿坦業 ，
1CHR|26|5|六子是 亞米利 ，七子是 以薩迦 ，八子是 毗烏利太 ，因為上帝賜福給 俄別‧以東 。
1CHR|26|6|他的兒子 示瑪雅 生了幾個兒子，都是大能的勇士，管理父親的家。
1CHR|26|7|示瑪雅 的兒子是 俄得尼 、 利法益 、 俄備得 、 以利薩巴 。 以利薩巴 的兄弟 以利戶 和 西瑪迦 是能人。
1CHR|26|8|這些都是 俄別‧以東 的子孫，他們和他們的兒子，以及兄弟，都是善於辦事的能人。屬 俄別‧以東 的共六十二人。
1CHR|26|9|米施利米雅 的兒子和兄弟都是能人，共十八人。
1CHR|26|10|米拉利 子孫中的 何薩 有幾個兒子：為首的是 申利 ；他原不是長子，是他父親立他為首的，
1CHR|26|11|次子是 希勒家 ，三子是 底巴利雅 ，四子是 撒迦利亞 。 何薩 的兒子和兄弟共十三人。
1CHR|26|12|這些是門口守衛的班次，各隨他們的班長，與他們的兄弟一同在耶和華殿裏按班供職。
1CHR|26|13|他們無論大小，都按著父系抽籤，分守各門。
1CHR|26|14|抽到東門的是 示利米雅 ；他的兒子 撒迦利亞 是精明的謀士，抽到北門。
1CHR|26|15|俄別‧以東 守南門，他的兒子守倉庫。
1CHR|26|16|書聘 與 何薩 守西門，在靠近 沙利基 門、通往上去的街道上，守衛與守衛相對。
1CHR|26|17|東門有六個 利未 人 ，北門每日有四人，南門每日有四人，庫房有兩人輪流替換。
1CHR|26|18|至於走廊，在西面街道上有四人，在走廊上有兩人。
1CHR|26|19|以上是 可拉 子孫和 米拉利 子孫門口守衛的班次。
1CHR|26|20|利未 人中有 亞希雅 管理上帝殿的庫房和聖物的庫房。
1CHR|26|21|拉但 子孫中， 革順 族屬 拉但 、作族長的是 革順 族屬 拉但 的 耶希伊利 。
1CHR|26|22|耶希伊利 的兒子 西坦 和他兄弟 約珥 管理耶和華殿的庫房。
1CHR|26|23|暗蘭 人、 以斯哈 人、 希伯倫 人、 烏薛 人也有職務。
1CHR|26|24|摩西 的孫子， 革舜 的兒子 細布業 管理庫房。
1CHR|26|25|還有他的弟兄： 以利以謝 ， 以利以謝 的兒子 利哈比雅 ， 利哈比雅 的兒子 耶篩亞 ， 耶篩亞 的兒子 約蘭 ， 約蘭 的兒子 細基利 ， 細基利 的兒子 示羅密 。
1CHR|26|26|這 示羅密 和他的兄弟管理一切庫房的聖物，就是 大衛 王和眾族長、千夫長、百夫長，以及軍官所分別為聖之物。
1CHR|26|27|他們把打仗時奪取的一些財物分別為聖，用來修造耶和華的殿。
1CHR|26|28|凡 撒母耳 先見、 基士 的兒子 掃羅 、 尼珥 的兒子 押尼珥 、 洗魯雅 的兒子 約押 分別為聖的，一切分別為聖之物都歸 示羅密 和他的兄弟掌管。
1CHR|26|29|以斯哈 人有 基拿尼雅 和他眾兒子作官長和審判官，管理 以色列 對外的事務。
1CHR|26|30|希伯倫 人有 哈沙比雅 和他弟兄一千七百人，都是能人，在 約旦河 西監督 以色列 人，辦理耶和華的一切工作和王的事務。
1CHR|26|31|希伯倫 人中有 耶利雅 作族長。 大衛 作王第四十年在各族各家從事尋訪，在 基列 的 雅謝 ，從這族中發現大能的勇士。
1CHR|26|32|耶利雅 的弟兄有二千七百人，都是能人，又是族長； 大衛 王派他們在 呂便 人、 迦得 人、 瑪拿西 半支派中管理上帝和王的一切事務。
1CHR|27|1|以色列 人的族長、千夫長、百夫長和官長都分配班次，每班二萬四千人，整年按月輪流出入，按班次服事王。
1CHR|27|2|正月第一班的班長是 撒巴第業 的兒子 雅朔班 ；他班內有二萬四千人。
1CHR|27|3|他是 法勒斯 的後裔，統管正月軍隊所有的官長。
1CHR|27|4|二月的班長是 亞何亞 人 朵代 ，他的班有總長 密基羅 ；他班內有二萬四千人。
1CHR|27|5|三月第三班的班長是 耶何耶大 祭司長的兒子 比拿雅 ；他班內有二萬四千人。
1CHR|27|6|這 比拿雅 是那三十人中的勇士，管理那三十人；他班內又有他兒子 暗米薩拔 。
1CHR|27|7|四月第四班的班長是 約押 的兄弟 亞撒黑 。接續他的是他兒子 西巴第雅 ；他班內有二萬四千人。
1CHR|27|8|五月第五班的班長是 伊斯拉 人 珊合 ；他班內有二萬四千人。
1CHR|27|9|六月第六班的班長是 提哥亞 人 益吉 的兒子 以拉 ；他班內有二萬四千人。
1CHR|27|10|七月第七班的班長是 以法蓮 族 比倫 人 希利斯 ；他班內有二萬四千人。
1CHR|27|11|八月第八班的班長是 謝拉 族 戶沙 人 西比該 ；他班內有二萬四千人。
1CHR|27|12|九月第九班的班長是 便雅憫 族 亞拿突 人 亞比以謝 ；他班內有二萬四千人。
1CHR|27|13|十月第十班的班長是 謝拉 族 尼陀法 人 瑪哈萊 ；他班內有二萬四千人。
1CHR|27|14|十一月第十一班的班長是 以法蓮 族 比拉頓 人 比拿雅 ；他班內有二萬四千人。
1CHR|27|15|十二月第十二班的班長是 俄陀聶 族 尼陀法 人 黑玳 ；他班內有二萬四千人。
1CHR|27|16|管理 以色列 眾支派的如下：管 呂便 人的是 細基利 的兒子 以利以謝 ；管 西緬 人的是 瑪迦 的兒子 示法提雅 ；
1CHR|27|17|管 利未 的是 基摩利 的兒子 哈沙比雅 ；管 亞倫 子孫的是 撒督 ；
1CHR|27|18|管 猶大 的是 大衛 的一個哥哥 以利戶 ；管 以薩迦 的是 米迦勒 的兒子 暗利 ；
1CHR|27|19|管 西布倫 的是 俄巴第雅 的兒子 伊施瑪雅 ；管 拿弗他利 的是 亞斯列 的兒子 耶利摩 ；
1CHR|27|20|管 以法蓮 的是 阿撒細雅 的兒子 何細亞 ；管 瑪拿西 半支派的是 毗大雅 的兒子 約珥 ；
1CHR|27|21|管 基列 地 瑪拿西 半支派的是 撒迦利亞 的兒子 易多 ；管 便雅憫 的是 押尼珥 的兒子 雅西業 ；
1CHR|27|22|管 但 的是 耶羅罕 的兒子 亞薩列 。以上是 以色列 眾支派的領袖。
1CHR|27|23|以色列 人二十歲以下的， 大衛 沒有記其數目；因耶和華曾應許，必加增 以色列 人如天上的星那樣多。
1CHR|27|24|洗魯雅 的兒子 約押 開始數點，卻還沒有數完。為了這事，烈怒臨到 以色列 ，數點的數目也沒有寫在《大衛王記》上。
1CHR|27|25|管理王的庫房的是 亞疊 的兒子 押斯馬威 。管理田野、城鎮、村莊、堡壘之倉庫的是 烏西雅 的兒子 約拿單 。
1CHR|27|26|管理耕田種地的是 基綠 的兒子 以斯利 。
1CHR|27|27|管理葡萄園的是 拉瑪 人 示每 。管理葡萄園酒窖的是 實弗米 人 撒巴底 。
1CHR|27|28|管理 謝非拉 橄欖樹和桑樹的是 基第利 人 巴勒‧哈南 。管理油庫的是 約阿施 。
1CHR|27|29|管理 沙崙 牧放牛群的是 沙崙 人 施提萊 。管理山谷牧養牛群的是 亞第萊 的兒子 沙法 。
1CHR|27|30|管理駱駝群的是 以實瑪利 人 阿比勒 。管理驢群的是 米崙 人 耶希底亞 。管理羊群的是 夏甲 人 雅悉 。
1CHR|27|31|這些都是為 大衛 王管理產業的領袖。
1CHR|27|32|大衛 的叔父 約拿單 作謀士；這人有智慧，又作書記。 哈摩尼 的兒子 耶歇 陪伴王的眾兒子。
1CHR|27|33|亞希多弗 作王的謀士。 亞基 人 戶篩 作王的顧問。
1CHR|27|34|亞希多弗 之後，有 比拿雅 的兒子 耶何耶大 ，以及 亞比亞他 接續他。 約押 作王的元帥。
1CHR|28|1|大衛 召集 以色列 所有的領袖，各支派的領袖、輪班服事王的官長、千夫長、百夫長、掌管王和王子一切產業牲畜的、宮廷官員、勇士，和所有大能的勇士，都到 耶路撒冷 來。
1CHR|28|2|大衛 王站起來，說：「我的弟兄，我的百姓啊，請聽我說！我心裏本想建造殿宇，安放耶和華的約櫃，作為我們上帝的腳凳，並且我已經預備了建造的材料。
1CHR|28|3|只是上帝對我說：『你不可為我的名建造殿宇，因你是戰士，流了人的血。』
1CHR|28|4|然而，耶和華－ 以色列 的上帝在我父的全家揀選我作 以色列 的王，直到永遠。因他揀選 猶大 為領袖，在 猶大 家中揀選我父家，在我父的眾兒子裏喜悅我，立我作全 以色列 的王。
1CHR|28|5|耶和華賜我許多兒子，在我兒子中揀選我兒子 所羅門 坐耶和華國度的王位，治理 以色列 。
1CHR|28|6|耶和華對我說：『你兒子 所羅門 必建造我的殿和院宇，因為我揀選他作我的子，我也必作他的父。
1CHR|28|7|他若恆久遵行我的誡命典章如今日一樣，我就必堅定他的國，直到永遠。』
1CHR|28|8|現今在 以色列 眾人眼前，在耶和華的會中，在我們上帝的垂聽下，你們務要遵行並尋求耶和華－你們上帝的一切誡命，如此你們就可以承受這美地，並留給你們的子孫，永遠為業。
1CHR|28|9|「我兒 所羅門 哪，你當認識耶和華－你父的上帝，全心樂意地事奉他，因為耶和華鑒察眾人的心，知道一切心思意念。你若尋求他，他必使你尋見；你若離棄他，他必永遠丟棄你。
1CHR|28|10|現在你當謹慎，因耶和華揀選你建造殿宇作為聖所。你當剛強去做。」
1CHR|28|11|大衛 指示他兒子 所羅門 有關殿的走廊、屋子、庫房、樓房、內殿和櫃蓋 之處的樣式，
1CHR|28|12|被靈感動所得的一切樣式：耶和華殿的院子、周圍一切的房屋、上帝殿的庫房和聖物庫房；
1CHR|28|13|祭司和 利未 人的班次，耶和華殿裏各樣事奉的工作，耶和華殿裏一切事奉用的器皿，
1CHR|28|14|以及各樣事奉所用金器的重量，和各樣事奉所用銀器的重量，
1CHR|28|15|金燈臺和金燈的重量，按每一個燈臺和燈的重量；銀燈臺和銀燈的重量，按每一個燈臺和燈的重量，都按照每一個燈臺的用途；
1CHR|28|16|每張供餅桌子的金子重量，和銀桌子的銀子重量，
1CHR|28|17|純金的肉叉子、盤子，和壺的重量，金碗，按每個金碗的重量，和銀碗，按每個銀碗的重量，
1CHR|28|18|純金香壇的重量，金基路伯座車的樣式，基路伯張開翅膀，遮蓋耶和華的約櫃。
1CHR|28|19|大衛 說：「這一切，所有工作的樣式，是耶和華用手寫的文件使我明白的。」
1CHR|28|20|大衛 又對他兒子 所羅門 說：「你當剛強壯膽去做！不要懼怕，也不要驚惶，因為耶和華上帝，我的上帝與你同在。他必不撇下你，也不丟棄你，直到耶和華殿的工作都完畢。
1CHR|28|21|看哪，有祭司和 利未 人的班次，為要辦理上帝殿各樣的事務，又有擅長做各樣事務的人，樂意在各樣工作上幫助你，並且領袖和眾百姓也都聽從你的一切命令。」
1CHR|29|1|大衛 王對全會眾說：「我兒子 所羅門 是上帝特選的，還年幼脆弱，但這工程浩大，因這殿不是為人，而是為耶和華上帝建造的。
1CHR|29|2|我為我上帝的殿已經盡力，預備金子做金器，銀子做銀器，銅做銅器，鐵做鐵器，木做木器，還有紅瑪瑙、可鑲嵌的寶石、彩石、各樣的寶石和許多大理石。
1CHR|29|3|此外，因我愛慕我上帝的殿，在預備建造聖殿的一切材料之外，又將我自己積蓄的金銀獻給我上帝的殿，
1CHR|29|4|就是三千他連得 俄斐 金子、七千他連得純銀，用來貼殿的牆；
1CHR|29|5|金子做金器，銀子做銀器，並藉工匠的手做一切的工。今日有誰願意將自己獻給耶和華呢？」
1CHR|29|6|於是，眾族長和 以色列 各支派的領袖、千夫長、百夫長，以及監管王工作的官長，都樂意奉獻。
1CHR|29|7|他們為上帝殿的工程獻上五千他連得又一萬達利克 金子，一萬他連得銀子，一萬八千他連得銅，十萬他連得鐵。
1CHR|29|8|凡有寶石的都送入耶和華殿的庫房，由 革順 人 耶歇 的手管理。
1CHR|29|9|因這些人全心樂意獻給耶和華，百姓就歡喜， 大衛 王也大大歡喜。
1CHR|29|10|大衛 在全會眾眼前稱頌耶和華； 大衛 說：「耶和華－ 以色列 的上帝，我們的父，你是應當稱頌的，直到永永遠遠！
1CHR|29|11|耶和華啊，尊大、能力、榮耀、勝利、威嚴都是你的；天上地下的一切都是你的；耶和華啊，國度是你的，並且你為至高，為萬有之首。
1CHR|29|12|豐富尊榮都從你而來，你也治理萬物。在你手裏有大能大力，你的手使人尊大強盛。
1CHR|29|13|我們的上帝啊，現在我們稱謝你，讚美你榮耀之名！
1CHR|29|14|「我算甚麼，我的百姓算甚麼，竟然能夠如此樂意奉獻？因為萬物都從你而來，我們把從你的手得來的獻給你。
1CHR|29|15|我們在你面前是客旅，是寄居的，與我們的列祖一樣。我們在世的日子如影子，沒有盼望。
1CHR|29|16|耶和華－我們的上帝啊，我們預備這許多材料，要為你的聖名建造殿宇，都是從你的手而來，都是屬你的。
1CHR|29|17|我的上帝啊，我知道你察驗人心，喜悅正直；我以正直的心樂意獻上這一切。現在我歡喜見你的百姓在此樂意奉獻給你。
1CHR|29|18|耶和華－我們列祖 亞伯拉罕 、 以撒 、 以色列 的上帝啊，求你使你的百姓心中常存這樣的心思意念，堅定他們的心歸向你，
1CHR|29|19|又求你賜我兒子 所羅門 全心遵守你的命令、法度、律例，成就這一切的事，用我所預備的建造殿宇。」
1CHR|29|20|大衛 對全會眾說：「你們應當稱頌耶和華－你們的上帝。」於是全會眾稱頌耶和華－他們列祖的上帝，低頭向耶和華和王下拜。
1CHR|29|21|次日，他們向耶和華獻平安祭和燔祭，獻一千頭公牛，一千隻公綿羊，一千隻羔羊，以及同獻的澆酒祭，並為 以色列 眾人獻許多的祭。
1CHR|29|22|那日，他們在耶和華面前吃喝，大大歡樂。 他們再次立 大衛 的兒子 所羅門 作王，膏他歸耶和華作君王，又膏 撒督 作祭司。
1CHR|29|23|於是 所羅門 坐在耶和華所賜的王位上，接續他父親 大衛 作王；他萬事亨通，全 以色列 都聽從他。
1CHR|29|24|眾領袖和勇士，以及 大衛 王的眾兒子，都順服 所羅門 王。
1CHR|29|25|耶和華使 所羅門 在 以色列 眾人眼前非常尊大，賜他君王的威嚴，勝過他以前任何一位 以色列 王。
1CHR|29|26|耶西 的兒子 大衛 作全 以色列 的王。
1CHR|29|27|他作 以色列 王的時期共四十年：在 希伯崙 作王七年，在 耶路撒冷 作王三十三年。
1CHR|29|28|他死的時候年紀老邁，日子滿足，享盡榮華富貴。他的兒子 所羅門 接續他作王。
1CHR|29|29|大衛 王自始至終的事蹟，看哪，都寫在 撒母耳 先見的書上、 拿單 先知的書上和 迦得 先見的書上，
1CHR|29|30|包括他治國的一切和他英勇的事蹟，以及他和 以色列 與世上列國所經歷的事。
2CHR|1|1|大衛 的兒子 所羅門 鞏固他的國度；耶和華－他的上帝與他同在，使他極其尊大。
2CHR|1|2|所羅門 吩咐全 以色列 ，就是千夫長、百夫長、審判官、全 以色列 的眾領袖和族長前來。
2CHR|1|3|所羅門 率領全會眾往 基遍 的丘壇去，因那裏有上帝的會幕，就是耶和華的僕人 摩西 在曠野所造的。
2CHR|1|4|只是上帝的約櫃， 大衛 已經從 基列‧耶琳 接到他所預備的地方，因他曾在 耶路撒冷 為約櫃支搭了帳幕，
2CHR|1|5|把 戶珥 的孫子， 烏利 的兒子 比撒列 所造的銅壇擺在 基遍 耶和華的會幕前。 所羅門 和會眾求告耶和華。
2CHR|1|6|所羅門 上到耶和華面前會幕的銅壇那裏，在壇上獻一千祭牲為燔祭。
2CHR|1|7|當夜，上帝向 所羅門 顯現，對他說：「你願我賜你甚麼，你可以求。」
2CHR|1|8|所羅門 對上帝說：「你曾向我父親 大衛 大施慈愛，使我接續他作王。
2CHR|1|9|耶和華上帝啊，現在求你實現向我父親 大衛 所應許的話；因你立我作這百姓的王，他們如同地上的塵沙那樣多。
2CHR|1|10|現在，求你賜我智慧聰明，好在這百姓面前出入；不然，誰能判斷你這麼多的百姓呢？」
2CHR|1|11|上帝對 所羅門 說：「你有這心意，不求資財、豐富、尊榮，也不求滅絕恨你之人的性命，又不求長壽；我既立你作我百姓的王，你只求智慧聰明，好審判我的百姓，
2CHR|1|12|我必賜你智慧聰明，也必賜你資財、豐富、尊榮，在你以前的列王未曾有過，在你以後也不會再有。」
2CHR|1|13|於是， 所羅門 從 基遍 丘壇會幕前回到 耶路撒冷 ，治理 以色列 。
2CHR|1|14|所羅門 聚集戰車騎兵；他有一千四百輛戰車，一萬二千名騎兵，安置在屯車城，在 耶路撒冷 的王那裏。
2CHR|1|15|王在 耶路撒冷 使金銀多如石頭，香柏木多如 謝非拉 的桑樹。
2CHR|1|16|所羅門 的馬是從 埃及 和 科威 運來的，是王的商人按著定價從 科威 買來的。
2CHR|1|17|他們從 埃及 進口戰車，每輛六百舍客勒銀子，馬每匹一百五十舍客勒； 赫 人眾王和 亞蘭 諸王的戰車和馬，也是經由他們的手出口的。
2CHR|2|1|所羅門 吩咐要為耶和華的名建造殿宇，又為自己的王國建造宮殿。
2CHR|2|2|所羅門 徵召七萬名扛抬的，八萬個在山上鑿石頭的人，三千六百個監工。
2CHR|2|3|所羅門 派人去見 推羅 王 希蘭 ，說：「你曾運香柏木給我父親 大衛 建造宮殿居住，請你也這樣待我。
2CHR|2|4|看哪，我要為耶和華－我上帝的名建造殿宇，分別為聖獻給他，在他面前燒芬芳的香，經常獻供餅，每早晚、安息日、初一，以及耶和華－我們上帝所定的節期獻燔祭。這是 以色列 人永遠的定例。
2CHR|2|5|我所要建造的殿宇宏大，因為我們的上帝至大，超乎眾神。
2CHR|2|6|天和天上的天，尚且不足他居住，誰能為他建造殿宇呢？我是誰，能為他建造殿宇嗎？不過在他面前燒香而已！
2CHR|2|7|現在請你派一個巧匠來，就是善用金、銀、銅、鐵，和紫色、朱紅色、藍色線做工，並精於雕刻之工的巧匠，與跟我一起在 猶大 和 耶路撒冷 、我父親 大衛 所預備的巧匠一同做工；
2CHR|2|8|又請你從 黎巴嫩 運香柏木、松木、檀香木到我這裏來，因我知道你的僕人擅長砍伐 黎巴嫩 的樹木。看哪，我的僕人必幫助你的僕人，
2CHR|2|9|好為我預備許多的木料，因我要建造的殿宇高大出奇。
2CHR|2|10|看哪，我必給你僕人，就是砍伐樹木的伐木工，二萬歌珥壓碎的小麥 ，二萬歌珥大麥，二萬罷特酒，二萬罷特油。」
2CHR|2|11|推羅 王 希蘭 寫信回答 所羅門 說：「耶和華因為愛他的百姓，所以立你作他們的王。」
2CHR|2|12|又說：「創造天和地的耶和華－ 以色列 的上帝是應當稱頌的！他賜給 大衛 王一個有智慧的兒子，使他有見識，有聰明，可以為耶和華建造殿宇，又為自己的王國建造宮殿。
2CHR|2|13|「現在我派一個精巧聰明的人去，他是我的師父 戶蘭 ，
2CHR|2|14|是 但 支派一個婦人的兒子，父親是 推羅 人。他善用金、銀、銅、鐵、石、木，和紫色、藍色、細麻和朱紅色線製造各物，並精於雕刻，又能設計各樣交給他做的圖案。我派這人與你的巧匠和你父親－我主 大衛 的巧匠一同做工。
2CHR|2|15|我主所說的小麥、大麥、酒、油，請運來給眾僕人。
2CHR|2|16|我們必照你所需用的，從 黎巴嫩 砍伐樹木，紮成筏子，浮海運到 約帕 ；你可以從那裏運到 耶路撒冷 。」
2CHR|2|17|所羅門 仿照他父親 大衛 數點所有在 以色列 地寄居的外邦人，共有十五萬三千六百名。
2CHR|2|18|他叫其中的七萬人作扛抬，八萬人在山上鑿石頭，三千六百人監督百姓工作。
2CHR|3|1|所羅門 在 耶路撒冷 開工建造耶和華的殿，就在耶和華向他父親 大衛 顯現的 摩利亞山 上， 耶布斯 人 阿珥楠 的禾場， 大衛 指定的地方。
2CHR|3|2|所羅門 作王第四年二月初二 開工建造。
2CHR|3|3|所羅門 所建築的上帝殿的根基是這樣：長六十肘，寬二十肘，都按著古時的尺寸。
2CHR|3|4|前面的 走廊長二十肘，與殿的寬度一樣，高一百二十肘；裏面貼上純金。
2CHR|3|5|大殿的牆都用松木板遮蔽，又貼上純金，上面刻著棕樹和鏈子。
2CHR|3|6|他用寶石裝飾這殿，使殿華美；金子都是 巴瓦音 的金子。
2CHR|3|7|他用金子貼殿和殿的棟梁、門檻、牆壁、門扇；牆上刻著基路伯。
2CHR|3|8|他建造至聖所，長二十肘，與殿的寬度一樣，寬二十肘，都貼上純金，共用了六百他連得金子。
2CHR|3|9|金的釘子重五十舍客勒。樓房都貼上金子。
2CHR|3|10|他又在至聖所用雕刻的手藝造兩個基路伯，包上金子。
2CHR|3|11|兩個基路伯的翅膀共長二十肘。這基路伯的一個翅膀長五肘，挨著殿這邊的牆；另一個翅膀也長五肘，與那基路伯翅膀相接。
2CHR|3|12|那基路伯的一個翅膀長五肘，挨著殿那邊的牆；另一個翅膀也長五肘，與這基路伯的翅膀相接。
2CHR|3|13|這兩個基路伯張開翅膀，共長二十肘，用腳站立，臉面向殿。
2CHR|3|14|他又用藍色、紫色、朱紅色線和細麻織幔子，在其上繡基路伯。
2CHR|3|15|他在殿前造了兩根柱子，高三十五肘；柱子上面的柱頂高五肘。
2CHR|3|16|他造鏈子在內殿裏，安在柱頂上，又做一百個石榴，安在鏈子上。
2CHR|3|17|他把兩根柱子立在殿前，一根在右邊，一根在左邊；右邊的起名叫 雅斤 ，左邊的起名叫 波阿斯 。
2CHR|4|1|他造一座銅壇，長二十肘，寬二十肘，高十肘。
2CHR|4|2|他又鑄一個銅海，周圍是圓的，直徑十肘，高五肘，用繩子量周圍是三十肘。
2CHR|4|3|銅海下面的周圍有牛的樣式，有十肘，繞著銅海；牛有兩行，是造銅海的時候鑄上去的。
2CHR|4|4|銅海安在十二頭銅牛上：三頭向北，三頭向西，三頭向南，三頭向東。銅海安在牛上，牛尾都向內。
2CHR|4|5|銅海厚一掌，邊如杯邊，像百合花，容量是三千罷特。
2CHR|4|6|他又造十個盆：五個放在右邊，五個放在左邊，作洗滌之用。獻燔祭所用之物都洗在盆內；但銅海是為祭司洗滌用的。
2CHR|4|7|他照所定的樣式造十個金燈臺，放在殿裏：五個在右邊，五個在左邊。
2CHR|4|8|他造十張桌子，放在殿裏：五張在右邊，五張在左邊。他又造一百個金碗。
2CHR|4|9|他建造祭司院和大院，以及院門，門扇包上銅。
2CHR|4|10|他把銅海安在殿的右邊，就是東南邊。
2CHR|4|11|戶蘭 又造了盆、鏟子和盤子。這樣， 戶蘭 為 所羅門 王做完了上帝殿的工：
2CHR|4|12|兩根柱子和柱子頂上兩個如碗的柱頂，以及蓋著如碗柱頂的兩個網子；
2CHR|4|13|四百個石榴，安在兩個網子上，每網兩行石榴，蓋著柱子上面兩個如碗的柱頂。
2CHR|4|14|他造盆座，又造其上的盆；
2CHR|4|15|銅海和其下的十二頭牛；
2CHR|4|16|盆、鏟子、肉叉。巧匠 戶蘭 給 所羅門 王為耶和華殿造的這一切器皿都是用磨亮的銅，
2CHR|4|17|是王在 約旦 平原、 疏割 和 撒利但 中間的泥巴地鑄成的。
2CHR|4|18|所羅門 造這一切器皿，數量很多，銅的重量無法計算。
2CHR|4|19|所羅門 又為上帝的殿造了各樣的器皿：金壇和獻供餅的供桌；
2CHR|4|20|純金的燈臺和燈盞，可以照定例點在內殿前；
2CHR|4|21|燈臺上的花和燈盞，以及燈剪，都是金的，而且是純金的；
2CHR|4|22|純金的鉗子、盤子、勺子、火盆。至於殿門和至聖所的門扇，以及殿的門扇，都是金的。
2CHR|5|1|所羅門 王做完了耶和華殿一切的工，就把他父親 大衛 分別為聖的金銀和一切器皿都帶來，放在上帝殿的庫房裏。
2CHR|5|2|於是， 所羅門 召集 以色列 的長老、各支派的領袖和 以色列 人的族長到 耶路撒冷 ，要把耶和華的約櫃從 大衛城 ，就是 錫安 ，接上來。
2CHR|5|3|在七月節期的時候，所有的 以色列 人都聚集到王那裏。
2CHR|5|4|以色列 眾長老一來到， 利未 人就抬起約櫃。
2CHR|5|5|祭司和 利未 人將約櫃請上來，又把會幕和會幕一切的聖器皿都帶上來。
2CHR|5|6|所羅門 王和聚集到他那裏的 以色列 全會眾都在約櫃前獻牛羊為祭，多得不可勝數，無法計算。
2CHR|5|7|祭司將耶和華的約櫃請進內殿，就是至聖所，安置在兩個基路伯的翅膀底下約櫃自己的地方。
2CHR|5|8|基路伯張開翅膀在約櫃上面的地方，從上面遮住約櫃和抬櫃的槓。
2CHR|5|9|這槓很長，從內殿前的約櫃可以看見槓頭，從外面卻看不見。這槓直到今日還在那裏。
2CHR|5|10|約櫃裏沒有別的，只有兩塊石版，就是 以色列 人出 埃及 ，耶和華與他們立約的時候， 摩西 在 何烈山 所放的。
2CHR|5|11|當時，所有在那裏的祭司，不論哪個班次供職的，都使自己分別為聖。祭司從聖所出來的時候，
2CHR|5|12|所有歌唱的 利未 人， 亞薩 、 希幔 、 耶杜頓 ，和他們的眾兒子、眾弟兄都穿細麻布衣服，站在祭壇的東邊敲鈸，鼓瑟，彈琴，和他們一起的還有一百二十個吹號的祭司。
2CHR|5|13|吹號的、歌唱的都合一齊聲，讚美稱謝耶和華。他們配合號筒、鐃鈸和其他樂器，揚聲讚美耶和華： 「耶和華本為善， 他的慈愛永遠長存！」 那時，耶和華的殿充滿了雲彩。
2CHR|5|14|祭司因雲彩的緣故不能站立供職，因為耶和華的榮光充滿了上帝的殿。
2CHR|6|1|那時， 所羅門 說： 「耶和華曾說要住在幽暗之處。
2CHR|6|2|我為你建了一座雄偉的殿宇， 作為你永遠居住的地方。」
2CHR|6|3|王轉過臉來為 以色列 全會眾祝福， 以色列 全會眾都站立。
2CHR|6|4|所羅門 說：「耶和華－ 以色列 的上帝是應當稱頌的！因他親口向我父 大衛 應許的，也親手成就了；他曾說：
2CHR|6|5|『自從那日我領我百姓出 埃及 地以來，我未曾在 以色列 各支派中選擇一城，在那裏為我的名建造殿宇，也未曾揀選一人作我百姓 以色列 的君王。
2CHR|6|6|但我選擇 耶路撒冷 ，使我的名留在那裏，又揀選 大衛 治理我的百姓 以色列 。』
2CHR|6|7|我父 大衛 的心意是要為耶和華－ 以色列 上帝的名建殿。
2CHR|6|8|耶和華卻對我父 大衛 說：『你有心為我的名建殿，這心意是好的；
2CHR|6|9|但你不可建殿，惟有你親生的兒子才可為我的名建殿。』
2CHR|6|10|現在耶和華實現了他所應許的話，使我接續我父 大衛 坐 以色列 的王位，正如耶和華所說的，我也為耶和華－ 以色列 上帝的名建造了這殿。
2CHR|6|11|我將約櫃安置在那裏，櫃內有耶和華的約，就是他與 以色列 人所立的約。」
2CHR|6|12|所羅門 當著 以色列 全會眾，站在耶和華的壇前，舉起手來。
2CHR|6|13|所羅門 曾造一個銅臺，長五肘，寬五肘，高三肘，放在院中。他站在臺上，當著 以色列 全會眾雙膝跪下，向天舉手，
2CHR|6|14|說：「耶和華－ 以色列 的上帝啊，天上地下沒有神明可與你相比！你向那些盡心行在你面前的僕人守約施慈愛，
2CHR|6|15|這約是你向你僕人 大衛 守的，是你應許他的。你親口應許，親手成就，正如今日一樣。
2CHR|6|16|耶和華－ 以色列 的上帝啊，你向你僕人我父 大衛 應許說：『你的子孫若謹慎自己的行為，遵行我的律法，像你在我面前所行的，就不斷有人在我面前坐 以色列 的王位。』現在求你信守這話。
2CHR|6|17|耶和華－ 以色列 的上帝啊，現在求你成就向你僕人 大衛 所應許的話。
2CHR|6|18|「上帝果真與世人同住在地上嗎？看哪，天和天上的天尚且不足容納你，何況我所建的這殿呢？
2CHR|6|19|惟求耶和華－我的上帝垂顧僕人的禱告祈求，俯聽僕人在你面前的祈禱呼求。
2CHR|6|20|願你的眼目晝夜看顧這殿，就是你應許立為你名的居所；求你垂聽禱告，你僕人向此處的禱告。
2CHR|6|21|你僕人和你百姓 以色列 向此處祈禱的時候，求你從天上你的居所垂聽，垂聽而赦免。
2CHR|6|22|「人若得罪鄰舍，有人強迫他，要他起誓，他來到這殿，在你的壇前起誓，
2CHR|6|23|求你從天上垂聽、處理，向你的僕人施行審判，定惡人有罪，照他所行的報應在他頭上；定義人為義，照他的義賞賜他。
2CHR|6|24|「你的百姓 以色列 若得罪你，敗在仇敵面前，卻又歸向你，宣認你的名，在這殿裏向你祈求禱告，
2CHR|6|25|求你從天上垂聽，赦免你百姓 以色列 的罪，使他們歸回你賜給他們和他們列祖之地。
2CHR|6|26|「你的百姓若得罪了你，你使天閉塞不下雨；他們若向此處禱告，宣認你的名，因你的懲罰而離開他們的罪，
2CHR|6|27|求你在天上垂聽，赦免你僕人你百姓 以色列 的罪，將當行的善道教導他們，並降雨在你的地，就是你賜給你百姓為業之地。
2CHR|6|28|「這地若有饑荒、瘟疫、焚風 、霉爛、蝗蟲、螞蚱，或有仇敵圍困這地的城門，無論遭遇甚麼災禍疾病，
2CHR|6|29|你的百姓 以色列 ，或眾人或一人，自覺災禍困苦，向這殿舉手，無論祈求甚麼，禱告甚麼，
2CHR|6|30|求你從天上你的居所垂聽赦免。因為你知道人心，惟有你知道世人的心，求你照各人所行的一切待他們，
2CHR|6|31|使他們在你賜給我們列祖的土地上一生一世敬畏你，遵行你的道。
2CHR|6|32|「論到不屬你百姓 以色列 的外邦人，若為你的大名和大能的手，以及伸出來的膀臂，從遠方而來，來向這殿禱告，
2CHR|6|33|求你從天上你的居所垂聽，照著外邦人向你所求的一切而行，使地上萬民都認識你的名，敬畏你，像你的百姓 以色列 一樣，又使他們知道我所建造的是稱為你名下的殿。
2CHR|6|34|「你的百姓若奉你的派遣出去，無論往何處與仇敵爭戰，他們若向你所選擇的這城和我為你名所建造的殿禱告，
2CHR|6|35|求你從天上垂聽他們的禱告祈求，為他們伸張正義。
2CHR|6|36|「你的百姓若得罪你，因為沒有人不犯罪，你向他們發怒，把他們交在仇敵面前，擄他們的人把他們帶到或遠或近之地；
2CHR|6|37|他們若在被擄之地那裏回心轉意，在被擄之地悔改，向你懇求說：『我們有罪了，我們悖逆了，我們作惡了』；
2CHR|6|38|他們若在被擄之地盡心盡性歸向你，又向自己的地，就是你賜給他們列祖的地和你所選擇的城，以及我為你名所建造的這殿禱告，
2CHR|6|39|求你從天上你的居所垂聽他們的禱告祈求，為他們伸張正義，赦免你的百姓向你犯的罪。
2CHR|6|40|我的上帝啊，現在求你睜眼看，側耳聽在此處所獻的禱告。
2CHR|6|41|「耶和華上帝啊，現在求你興起， 與你有能力的約櫃同入安歇之所。 耶和華上帝啊，願你的祭司披上救恩， 願你的聖民蒙福歡樂。
2CHR|6|42|耶和華上帝啊，求你不要厭棄你的受膏者， 要記得向你僕人 大衛 所施的慈愛。」
2CHR|7|1|所羅門 祈禱完畢，就有火從天降下來，燒盡燔祭和祭物。耶和華的榮光充滿了殿；
2CHR|7|2|因耶和華的榮光充滿了耶和華的殿，所以祭司不能進耶和華的殿。
2CHR|7|3|那火降下、耶和華的榮光在殿上的時候， 以色列 眾人看見，就在石板地俯伏敬拜，稱謝耶和華： 「耶和華本為善， 他的慈愛永遠長存！」
2CHR|7|4|王和眾百姓在耶和華面前獻祭。
2CHR|7|5|所羅門 王獻二萬二千頭牛，十二萬隻羊為祭。這樣，王和眾百姓為上帝的殿行了奉獻之禮。
2CHR|7|6|祭司各供其職侍立， 利未 人拿著耶和華的樂器，就是 大衛 王所造、為要頌讚耶和華的樂器，因他的慈愛永遠長存；他們為 大衛 的讚美詩奏樂；祭司在眾人面前吹號， 以色列 眾人都站立。
2CHR|7|7|所羅門 因他所造的銅壇容不下燔祭、素祭和脂肪，就將耶和華殿前院子的中間分別為聖，在那裏獻燔祭和平安祭牲的脂肪。
2CHR|7|8|那時 所羅門 守節七日，從 哈馬口 直到 埃及 溪谷的 以色列 眾人都與他同在一起，成了一個極其盛大的會。
2CHR|7|9|第八日他們舉行嚴肅會，行奉獻壇的禮七日，守節七日。
2CHR|7|10|七月二十三日，王差遣百姓回自己的帳棚去；他們為耶和華向 大衛 和 所羅門 ，以及他百姓 以色列 所施的恩惠，心裏都歡喜快樂。
2CHR|7|11|所羅門 建完了耶和華的殿和王宮；在耶和華的殿和王宮的工程上，凡他心中所要做的，都順利做成了。
2CHR|7|12|夜間耶和華向 所羅門 顯現，對他說：「我已聽了你的禱告，也選擇這地方歸我作獻祭的殿宇。
2CHR|7|13|我若使天閉塞不下雨，或使蝗蟲吃這地的出產，或降瘟疫在我子民中，
2CHR|7|14|這稱為我名下的子民，若是謙卑自己，禱告，尋求我的面，轉離他們的惡行，我必從天上垂聽，赦免他們的罪，醫治他們的地。
2CHR|7|15|我必睜眼看，側耳聽在此處所獻的禱告。
2CHR|7|16|現在我已選擇這殿，分別為聖，使我的名永在其中；我的眼、我的心也必時常在那裏。
2CHR|7|17|你若行在我面前，效法你父 大衛 所行的，遵行我一切所吩咐你的，謹守我的律例典章，
2CHR|7|18|我就必堅固你國度的王位，正如我與你父 大衛 所立的約，說：『你的子孫必不斷有人治理 以色列 。』
2CHR|7|19|「倘若你們轉去，離棄我擺在你們面前的律例誡命，去事奉別神，敬拜它們，
2CHR|7|20|我就必把 以色列 人從我賜給他們的地上連根拔起，也必從我面前捨棄那為我名所分別為聖的殿，使它在萬民中成為笑柄，被人譏誚。
2CHR|7|21|這殿雖然崇高，將來凡經過的人必驚訝說：『耶和華為何向這地和這殿如此行呢？』
2CHR|7|22|人必說：『因為此地的人離棄領他們祖先出 埃及 地的耶和華－他們的上帝，去親近別神，敬拜事奉它們，所以耶和華使這一切災禍臨到他們。』」
2CHR|8|1|所羅門 建造耶和華的殿和王宮，用了二十年才完成。
2CHR|8|2|所羅門 修築 希蘭 送給他的城鎮，使 以色列 人住在那裏。
2CHR|8|3|所羅門 往 哈馬‧瑣巴 去，攻取了那地方。
2CHR|8|4|所羅門 建造曠野的 達莫 ，建造 哈馬 一切的儲貨城，
2CHR|8|5|又建造 上伯‧和崙 、 下伯‧和崙 ，成為有牆、門、閂的堡壘城。
2CHR|8|6|所羅門 建造 巴拉 和一切的儲貨城、戰車城、戰馬城，以及他所想要建造的，在 耶路撒冷 、 黎巴嫩 ，和自己所治理全國中的一切建設。
2CHR|8|7|至於所有剩下的百姓，不屬 以色列 的 赫 人、 亞摩利 人、 比利洗 人、 希未 人、 耶布斯 人，
2CHR|8|8|那些 以色列 人在當地不能滅盡的人， 所羅門 徵召他們剩下的後代服勞役，直到今日。
2CHR|8|9|惟有 以色列 人， 所羅門 不使他們當奴僕做工，而是作他的戰士、軍官、戰車長、騎兵長。
2CHR|8|10|這些是 所羅門 王的監工，共有二百五十名百姓的監工。
2CHR|8|11|所羅門 把法老的女兒遷出 大衛城 ，上到他為她建造的宮裏，因 所羅門 說：「耶和華約櫃所到之處都是聖地，所以我的妻子不可住在 以色列 王 大衛 的宮裏。」
2CHR|8|12|那時， 所羅門 在走廊前他所築的耶和華的壇上，向耶和華獻燔祭，
2CHR|8|13|又遵照 摩西 的吩咐，在安息日、初一，以及每年在除酵節、七七節、住棚節三個節期，獻每日所當獻上的祭。
2CHR|8|14|所羅門 照著他父親 大衛 所定的條例，分派祭司的班次，擔任他們的職務，又分派 利未 人的任務，負責頌讚，並在祭司面前做每日當做的事，又派門口的守衛按著班次看守各門，因為神人 大衛 是這樣吩咐的。
2CHR|8|15|王對眾祭司和 利未 人的吩咐，無論是管理庫房或任何事務，他們都不違背。
2CHR|8|16|所羅門 所有的工作都準備就緒，從立耶和華殿的根基直到完工的日子。耶和華的殿就完成了。
2CHR|8|17|那時， 所羅門 往 以東 地海岸的 以旬‧迦別 和 以祿 去。
2CHR|8|18|希蘭 派他的臣僕，把船隻和熟悉航海的僕人送到 所羅門 那裏。他們同 所羅門 的僕人到了 俄斐 ，從那裏得了四百五十他連得金子，運到 所羅門 王那裏。
2CHR|9|1|示巴 女王聽見 所羅門 的名聲，就來到 耶路撒冷 ，要用難題考問 所羅門 。她帶著很多的隨從，有駱駝馱著香料、許多金子和寶石。她來到 所羅門 那裏，向他提出心中所有的問題。
2CHR|9|2|所羅門 回答了她所有的問題，沒有一個問題太難，是 所羅門 不能向她解答的。
2CHR|9|3|示巴 女王看見 所羅門 的智慧和他所建造的宮殿，
2CHR|9|4|席上的食物，坐著的群臣，侍立的僕人和他們的服裝，司酒長和他們的服裝，以及他上耶和華殿的臺階 ，就詫異得神不守舍。
2CHR|9|5|她對王說：「我在本國所聽到的話，論到你的事和你的智慧是真的！
2CHR|9|6|我本來不信那些話，及至我來親眼看見了，看哪，人所告訴我的，還不及你豐富智慧的一半，超過我所聽見的傳聞。
2CHR|9|7|你的人是有福的！你這些常侍立在你面前、聽你智慧話的僕人是有福的！
2CHR|9|8|耶和華－你的上帝是應當稱頌的！他喜愛你，使你坐他的王位，為耶和華－你的上帝作王；因為你的上帝愛 以色列 ，要永遠堅立它，所以立你作他們的王，使你秉公行義。」
2CHR|9|9|於是 示巴 女王把一百二十他連得金子、極多的香料和寶石送給 所羅門 王；從來沒有像 示巴 女王送給 所羅門 王那麼多的香料。
2CHR|9|10|希蘭 的僕人和 所羅門 的僕人也從 俄斐 運了金子來，又運了檀香木和寶石來。
2CHR|9|11|王用檀香木為耶和華的殿和王宮做階梯，又為歌唱的人做琴瑟； 猶大 地從來沒有見過這樣的。
2CHR|9|12|所羅門 王除了回贈 示巴 女王所帶來的，凡她所提出的一切要求， 所羅門 王都送給她。於是女王和她臣僕轉回，到本國去了。
2CHR|9|13|所羅門 每年所得的金子，重六百六十六他連得，
2CHR|9|14|另外還有從商人和貿易所收到的，以及 阿拉伯 諸王和各地的省長進貢給 所羅門 的金銀。
2CHR|9|15|所羅門 王用錘出來的金子打成二百面盾牌，每面盾牌用六百舍客勒錘出來的金子；
2CHR|9|16|又用錘出來的金子打成三百面小盾牌，每面小盾牌用三百舍客勒金子。王把它們放在 黎巴嫩林宮 裏。
2CHR|9|17|王又製造一個大的象牙寶座，包上純金。
2CHR|9|18|寶座有六層臺階，又有金腳凳，與寶座相連。座位之處兩旁有扶手，靠近扶手有兩隻獅子站立。
2CHR|9|19|六層臺階上有十二隻獅子站立，分站左邊和右邊；任何國度都沒有這樣做的。
2CHR|9|20|所羅門 王一切的飲器都是金的， 黎巴嫩林宮 裏所有的器皿都是純金的。在 所羅門 的日子，銀子算不了甚麼。
2CHR|9|21|因王的船隻與 希蘭 的僕人一同往 他施 去， 他施 船隻每三年一次把金、銀、象牙、猿猴、孔雀 運回來。
2CHR|9|22|所羅門 王的財寶與智慧勝過地上的眾王。
2CHR|9|23|地上的眾王都求見 所羅門 的面，要聽上帝放在他心裏的智慧。
2CHR|9|24|他們各帶貢物，就是銀器、金器、衣服、兵器、香料、馬、騾子，每年都有一定的數量。
2CHR|9|25|所羅門 擁有給戰車和馬用的四千個棚子，還有一萬二千名騎兵，安置在屯車城，在 耶路撒冷 的王那裏。
2CHR|9|26|所羅門 統管諸王，從 大河 到 非利士 人的地，直到 埃及 的邊界。
2CHR|9|27|王在 耶路撒冷 使銀子多如石頭，香柏木多如 謝非拉 的桑樹。
2CHR|9|28|有人從 埃及 和各國為 所羅門 把馬匹運來。
2CHR|9|29|所羅門 其餘的事，自始至終，不都寫在 拿單 先知的書上和 示羅 人 亞希雅 的《預言書》上，以及 易多 先見論 尼八 兒子 耶羅波安 的《默示書》上嗎？
2CHR|9|30|所羅門 在 耶路撒冷 作全 以色列 的王四十年。
2CHR|9|31|所羅門 與他祖先同睡，葬在他父親 大衛 的城裏，他兒子 羅波安 接續他作王。
2CHR|10|1|羅波安 往 示劍 去，因 以色列 眾人都到了 示劍 ，要立他作王。
2CHR|10|2|尼八 的兒子 耶羅波安 先前躲避 所羅門 王，逃往 埃及 ，住在那裏；他聽見這事，就從 埃及 回來。
2CHR|10|3|以色列 人派人去請他來。 耶羅波安 就和 以色列 眾人來，與 羅波安 談話，說：
2CHR|10|4|「你父親使我們負重軛，現在求你減輕你父親所加給我們的苦工和重軛，我們就服事你。」
2CHR|10|5|羅波安 對他們說：「過三天再來見我吧！」百姓就走了。
2CHR|10|6|羅波安 的父親 所羅門 在世的時候，有侍立在他面前的長者， 羅波安 王和他們商議，說：「你們出個主意，好把話帶回給這百姓。」
2CHR|10|7|他們對他說：「王若恩待這百姓，使他們喜悅，跟他們說好話，他們就永遠作王的僕人了。」
2CHR|10|8|王不採納長者給他出的主意，卻和那些與他一同長大、在他面前侍立的年輕人商議。
2CHR|10|9|他對他們說：「這百姓對我說：『你父親使我們負重軛，求你減輕一些。』你們出個甚麼主意，我們好把話帶回給他們。」
2CHR|10|10|那些與他一同長大的年輕人對他說：「這些百姓對王說：『你父親使我們負重軛，求你給我們減輕一些。』王要對他們如此說：『我的小指頭比我父親的腰還粗呢！
2CHR|10|11|我父親使你們負重軛，現在我必使你們負更重的軛！我父親用鞭子懲罰你們，我卻要用蠍子！』」
2CHR|10|12|耶羅波安 和眾百姓遵照王所說「你們第三天再來見我」的話，第三天來到 羅波安 那裏。
2CHR|10|13|王嚴厲地回答他們。 羅波安 王不採納長者所出的主意，
2CHR|10|14|卻照著年輕人所出的主意對他們說：「我 使你們負重軛，我必使你們負更重的軛！我父親用鞭子懲罰你們，我卻要用蠍子！」
2CHR|10|15|王不依從百姓，因這事件是出於上帝，為要應驗耶和華藉 示羅 人 亞希雅 對 尼八 的兒子 耶羅波安 所說的話。
2CHR|10|16|以色列 眾人見王不依從他們，百姓就回覆王說： 「我們在 大衛 中有甚麼分呢？ 我們在 耶西 的兒子中沒有產業！ 以色列 啊，各回自己的帳棚去吧！ 大衛 啊，現在你顧自己的家吧！」 於是， 以色列 眾人都回自己的帳棚去了；
2CHR|10|17|至於住 猶大 城鎮的 以色列 人， 羅波安 仍作他們的王。
2CHR|10|18|羅波安 王派監管勞役的 哈多蘭 去， 以色列 人用石頭打他，他就死了。 羅波安 王急忙上車，逃回 耶路撒冷 去了。
2CHR|10|19|這樣， 以色列 背叛 大衛 家，直到今日。
2CHR|11|1|羅波安 來到 耶路撒冷 ，召集 猶大 家和 便雅憫 家，共十八萬人，都是精選的戰士，要與 以色列 爭戰，好將國奪回再歸自己。
2CHR|11|2|但耶和華的話臨到神人 示瑪雅 ，說：
2CHR|11|3|「你去告訴 所羅門 的兒子 猶大 王 羅波安 和住 猶大 、 便雅憫 的 以色列 眾人，說：
2CHR|11|4|『耶和華如此說：你們不可上去與你們的弟兄爭戰。各自回家去吧！因為這事是出於我。』」眾人就聽從耶和華的話回去，不去與 耶羅波安 爭戰。
2CHR|11|5|羅波安 住在 耶路撒冷 ，在 猶大 為防禦修築城鎮，
2CHR|11|6|他修築 伯利恆 、 以坦 、 提哥亞 、
2CHR|11|7|伯‧夙 、 梭哥 、 亞杜蘭 、
2CHR|11|8|迦特 、 瑪利沙 、 西弗 、
2CHR|11|9|亞多萊音 、 拉吉 、 亞西加 、
2CHR|11|10|瑣拉 、 亞雅崙 、 希伯崙 。這都是 猶大 和 便雅憫 的堅固城。
2CHR|11|11|羅波安 又鞏固這些堡壘，在其中安置軍官，儲備糧食、油和酒。
2CHR|11|12|他在各城裏預備盾牌和槍，使城極其堅固。 猶大 和 便雅憫 都歸了他。
2CHR|11|13|全 以色列 的祭司和 利未 人都從四方來歸 羅波安 。
2CHR|11|14|利未 人放棄他們的郊野和產業，來到 猶大 與 耶路撒冷 ，因為 耶羅波安 和他的兒子拒絕他們，不許他們擔任祭司事奉耶和華。
2CHR|11|15|耶羅波安 為丘壇，為山羊鬼魔，為自己所造的牛犢設立祭司。
2CHR|11|16|以色列 各支派中，凡立定心意尋求耶和華－ 以色列 上帝的，都隨從 利未 人來到 耶路撒冷 獻祭給耶和華－他們列祖的上帝。
2CHR|11|17|這就鞏固了 猶大 王國，使 所羅門 的兒子 羅波安 強盛三年，因為這三年他們遵行 大衛 和 所羅門 的道。
2CHR|11|18|羅波安 娶 大衛 兒子 耶利末 的女兒 瑪哈拉 為妻，又娶 耶西 兒子 以利押 的女兒 亞比孩 為妻，
2CHR|11|19|從她生了幾個兒子，就是 耶烏施 、 示瑪利雅 和 撒罕 。
2CHR|11|20|後來他又娶 押沙龍 的女兒 瑪迦 ，從她生了 亞比雅 、 亞太 、 細撒 和 示羅密 。
2CHR|11|21|羅波安 有十八個妻和六十個妾，生了二十八個兒子，六十個女兒；他卻愛 押沙龍 的女兒 瑪迦 ，過於愛其他的妻妾。
2CHR|11|22|羅波安 立 瑪迦 的兒子 亞比雅 作太子，在他兄弟中為首，因為要立他作王。
2CHR|11|23|羅波安 辦事精明，把他眾兒子分散在 猶大 和 便雅憫 全地各堅固城裏，賜他們大量的糧食，又給他們娶許多妻子。
2CHR|12|1|羅波安 的王國穩固，他強盛的時候就離棄耶和華的律法，全 以色列 都跟從他。
2CHR|12|2|羅波安 王第五年， 埃及 王 示撒 上來攻打 耶路撒冷 ，因為他們背叛了耶和華。
2CHR|12|3|示撒 帶著一千二百輛戰車，六萬名騎兵，以及跟隨他從 埃及 出來的 路比 人、 蘇基 人和 古實 人的軍隊，多得不可勝數。
2CHR|12|4|他攻取了 猶大 的堅固城，來到 耶路撒冷 。
2CHR|12|5|那時， 猶大 的領袖因為 示撒 的緣故聚集在 耶路撒冷 ，有先知 示瑪雅 去見 羅波安 和眾領袖，對他們說：「耶和華如此說：『你們離棄了我，所以我也離棄你們，把你們交在 示撒 手裏。』」
2CHR|12|6|於是 以色列 的領袖和王都謙卑說：「耶和華是公義的。」
2CHR|12|7|耶和華見他們謙卑，耶和華的話就臨到 示瑪雅 ，說：「他們既謙卑，我必不滅絕他們；我要使他們暫時得拯救，不藉著 示撒 的手將我的怒氣倒在 耶路撒冷 。
2CHR|12|8|然而他們必作 示撒 的僕人，好叫他們知道，服事我與服事地上邦國有何分別。」
2CHR|12|9|於是， 埃及 王 示撒 上來攻取 耶路撒冷 ，奪了耶和華殿和王宮裏的寶物，盡都帶走，又奪走 所羅門 製造的金盾牌。
2CHR|12|10|羅波安 王製造銅盾牌代替那些金盾牌，交給看守王宮宮門的護衛長看管。
2CHR|12|11|每逢王進耶和華的殿，護衛兵就來，舉起這些盾牌；隨後仍將盾牌送回護衛室。
2CHR|12|12|王謙卑的時候，耶和華的怒氣就轉消了，不全然滅盡，並且在 猶大 中，情況也有好轉。
2CHR|12|13|羅波安 王自強，在 耶路撒冷 作王。他登基的時候年四十一歲，在 耶路撒冷 ，就是耶和華從 以色列 眾支派中所選擇立他名的城，作王十七年。 羅波安 的母親名叫 拿瑪 ，是 亞捫 人。
2CHR|12|14|羅波安 行惡，因他沒有立定心意尋求耶和華。
2CHR|12|15|羅波安 的事蹟，自始至終不都寫在 示瑪雅 先知和 易多 先見的《史記》上嗎？ 羅波安 與 耶羅波安 時常交戰。
2CHR|12|16|羅波安 與他祖先同睡，葬在 大衛城 ，他的兒子 亞比雅 接續他作王。
2CHR|13|1|耶羅波安 王十八年， 亞比雅 登基作 猶大 王，
2CHR|13|2|在 耶路撒冷 作王三年。他母親名叫 米該亞 ，是 基比亞 人 烏列 的女兒 。 亞比雅 常與 耶羅波安 交戰。
2CHR|13|3|有一次 亞比雅 率領四十萬精選的士兵出戰，他們都是勇敢的戰士； 耶羅波安 也率領八十萬精選的大能勇士，迎著 亞比雅 擺陣。
2CHR|13|4|亞比雅 站在 以法蓮 山區中的 洗瑪臉山 上，說：「 耶羅波安 和 以色列 眾人哪，要聽我說！
2CHR|13|5|耶和華－ 以色列 的上帝曾立鹽約，將 以色列 國永遠賜給 大衛 和他的子孫，你們不知道嗎？
2CHR|13|6|但 大衛 兒子 所羅門 的臣僕、 尼八 的兒子 耶羅波安 起來背叛他的主人。
2CHR|13|7|有些無賴的歹徒聚集跟從他，逞強攻擊 所羅門 的兒子 羅波安 ；那時 羅波安 還年輕，心志軟弱，不能抵擋他們。
2CHR|13|8|「現在你們說要抗拒 大衛 子孫手下所治理的耶和華的國，你們的人數眾多，你們那裏又有 耶羅波安 為你們所造當作神明的金牛犢。
2CHR|13|9|你們不是驅逐耶和華的祭司 亞倫 的後裔和 利未 人嗎？不是照著外邦人的惡俗為自己立祭司嗎？無論何人牽一頭公牛犢、七隻公綿羊將自己分別出來，就可作虛無神明的祭司。
2CHR|13|10|至於我們，耶和華是我們的上帝，我們並沒有離棄他。我們有事奉耶和華的祭司，都是 亞倫 的後裔，並有 利未 人各盡其職。
2CHR|13|11|他們每日早晚向耶和華獻燔祭，燒芬芳的香，又在純金的 供桌上擺供餅，每晚點燃金燈臺上的燈盞，因為我們遵守耶和華－我們上帝的命令，但你們卻離棄了他。
2CHR|13|12|看哪，率領我們的是上帝，又有他的祭司拿號向你們吹出響聲。 以色列 人哪，不要與耶和華－你們列祖的上帝爭戰，因你們必不能得勝。」
2CHR|13|13|耶羅波安 卻在 猶大 人的後頭設伏兵。這樣， 以色列 人在 猶大 人的前頭，伏兵在 猶大 人的後頭。
2CHR|13|14|猶大 人轉過來，看哪，前後都有戰事，就呼求耶和華，祭司也吹號。
2CHR|13|15|於是 猶大 人吶喊。 猶大 人吶喊的時候，上帝就擊打 耶羅波安 和 以色列 眾人，使他們敗在 亞比雅 與 猶大 人面前。
2CHR|13|16|以色列 人在 猶大 人面前逃跑，上帝將他們交在 猶大 人手裏。
2CHR|13|17|亞比雅 和他的軍兵大大擊殺 以色列 人， 以色列 人被殺仆倒的精兵有五十萬。
2CHR|13|18|那時， 以色列 人被制伏了。 猶大 人得勝，因為他們倚靠耶和華－他們列祖的上帝。
2CHR|13|19|亞比雅 追趕 耶羅波安 ，攻取了他的幾座城，就是 伯特利 和所屬的鄉鎮 ， 耶沙拿 和所屬的鄉鎮， 以法拉音 和所屬的鄉鎮。
2CHR|13|20|亞比雅 在世的時候， 耶羅波安 不再強盛；耶和華擊打他，他就死了。
2CHR|13|21|亞比雅 卻漸漸強盛。他娶了十四個妻妾，生了二十二個兒子，十六個女兒。
2CHR|13|22|亞比雅 其餘的事和他的言行都寫在 易多 先知的評傳上。
2CHR|14|1|亞比雅 與他祖先同睡，葬在 大衛城 ，他的兒子 亞撒 接續他作王。 亞撒 在位期間，國中太平十年。
2CHR|14|2|亞撒 行耶和華－他上帝眼中看為善為正的事，
2CHR|14|3|除掉外邦的祭壇和丘壇，打碎柱像，砍下 亞舍拉 ，
2CHR|14|4|吩咐 猶大 人尋求耶和華－他們列祖的上帝，遵行他的律法和誡命，
2CHR|14|5|又在 猶大 各城鎮除掉丘壇和香壇。在他治理下，國中太平。
2CHR|14|6|他在 猶大 建造了幾座堅固城。那些年間，國中太平，沒有戰爭，因為耶和華賜他平安。
2CHR|14|7|他對 猶大 人說：「我們要建造這些城鎮，四圍築牆，蓋城樓，安門，做閂；地仍屬於我們，因為我們尋求耶和華－我們的上帝；我們尋求他，他就賜我們四境平安。」於是他們建造城鎮，諸事亨通。
2CHR|14|8|亞撒 的軍兵，出自 猶大 拿盾牌拿槍的三十萬人，出自 便雅憫 拿小盾牌拉弓的二十八萬人；這些全都是大能的勇士。
2CHR|14|9|古實 人 謝拉 率領一百萬軍兵，三百輛戰車，出來攻擊 猶大 人，到了 瑪利沙 。
2CHR|14|10|亞撒 出去迎戰，在 瑪利沙 的 洗法谷 彼此擺陣。
2CHR|14|11|亞撒 呼求耶和華－他的上帝說：「耶和華啊，在強弱之間，惟有你能幫助。耶和華－我們的上帝啊，求你幫助我們，因為我們仰賴你，奉你的名來抵擋這大軍。耶和華啊，你是我們的上帝，不要讓人勝過你。」
2CHR|14|12|於是耶和華擊打 古實 人，使他們敗在 亞撒 和 猶大 人面前， 古實 人就逃跑了。
2CHR|14|13|亞撒 和跟隨他的軍兵追趕他們，直到 基拉耳 。 古實 人被殺的很多，無法復原，因為他們在耶和華與他軍兵面前被擊潰。 猶大 人奪了許多財物，
2CHR|14|14|又攻打 基拉耳 四圍一切的城鎮；城中的人都懼怕耶和華。 猶大 人擄掠了一切的城鎮，因其中的財物很多，
2CHR|14|15|又毀壞了群畜的圈，奪取許多的羊和駱駝，就回 耶路撒冷 去了。
2CHR|15|1|上帝的靈臨到 俄德 的兒子 亞撒利雅 。
2CHR|15|2|他出來迎接 亞撒 ，對他說：「 亞撒 ， 猶大 和 便雅憫 眾人哪，要聽我說：你們若順從耶和華，耶和華必與你們同在；你們若尋求他，就必尋見；你們若離棄他，他必離棄你們。
2CHR|15|3|以色列 人不信真神，沒有訓誨的祭司，也沒有律法，已經許多日子了。
2CHR|15|4|但他們在急難的時候歸向耶和華－ 以色列 的上帝，尋求他，他就被他們尋見。
2CHR|15|5|那時，出入的人不得平安，各地的居民都遭大亂；
2CHR|15|6|他們被破壞殆盡，這國攻擊那國，這城攻擊那城，因為上帝用各樣災難擾亂他們。
2CHR|15|7|現在你們要剛強，不要手軟，因你們所行的必得賞賜。」
2CHR|15|8|亞撒 聽見這些話和 俄德 先知的預言，就壯起膽來，在 猶大 和 便雅憫 全地，以及 以法蓮 山區所奪的各城，把其中的可憎之物盡都除掉，又在耶和華殿的走廊前重新修築耶和華的壇。
2CHR|15|9|他又召集 猶大 和 便雅憫 眾人，以及他們中間寄居的 以法蓮 人、 瑪拿西 人、 西緬 人。有許多 以色列 人歸順 亞撒 ，因為他們看見耶和華－他的上帝與他同在。
2CHR|15|10|亞撒 作王第十五年三月，他們都聚集在 耶路撒冷 。
2CHR|15|11|那日他們從所取的擄物中，將七百頭牛和七千隻羊獻給耶和華。
2CHR|15|12|他們立約，要盡心盡性尋求耶和華－他們列祖的上帝。
2CHR|15|13|凡不尋求耶和華－ 以色列 上帝的，無論大小、男女，必被處死。
2CHR|15|14|他們就大聲歡呼，吹號吹角，向耶和華起誓。
2CHR|15|15|猶大 眾人為所起的誓歡喜，因他們盡心起誓，盡意尋求耶和華，耶和華就被他們尋見，且賜他們四境平安。
2CHR|15|16|亞撒 王甚至廢了他祖母 瑪迦 太后的位，因 瑪迦 造了可憎的 亞舍拉 。 亞撒 砍下她的偶像，搗得粉碎，在 汲淪溪 邊燒了，
2CHR|15|17|只是丘壇還沒有從 以色列 中廢去，然而 亞撒 一生有純正的心。
2CHR|15|18|亞撒 將他父親所分別為聖與自己所分別為聖的金銀和器皿都奉到上帝的殿裏。
2CHR|15|19|亞撒 作王直到第三十五年，都沒有戰事。
2CHR|16|1|亞撒 作王第三十六年， 以色列 王 巴沙 上來攻擊 猶大 ，修築 拉瑪 ，不許人從 猶大 王 亞撒 那裏出入。
2CHR|16|2|於是 亞撒 從耶和華殿和王宮的府庫裏拿出金銀來，送給住在 大馬士革 的 亞蘭 王 便‧哈達 ，說：
2CHR|16|3|「你父曾與我父立約，我與你也要這樣立約。看哪，我把金銀送給你，請你廢掉你與 以色列 王 巴沙 所立的約，使他從我這裏撤退。」
2CHR|16|4|便‧哈達 聽從了 亞撒 王，就派遣他的軍官去攻打 以色列 的城鎮。他們攻下了 以雲 、 但 、 亞伯‧瑪音 和 拿弗他利 一切的儲貨城。
2CHR|16|5|巴沙 聽見了，就停工不修築 拉瑪 ，任由他的工程停止。
2CHR|16|6|於是 亞撒 王率領 猶大 眾人，運走 巴沙 修築 拉瑪 所用的石頭和木料，用以修築 迦巴 和 米斯巴 。
2CHR|16|7|那時， 哈拿尼 先見來見 猶大 王 亞撒 ，對他說：「因你仰賴 亞蘭 王，沒有仰賴耶和華－你的上帝，所以 亞蘭 王的軍兵逃脫了你的手。
2CHR|16|8|古實 人和 路比 人的軍隊不是非常強大嗎？他們的戰車騎兵不是極多嗎？只因你仰賴耶和華，他就將他們交在你手裏。
2CHR|16|9|因為耶和華的眼目遍察全地，要堅固向他存純正之心的人。你在這事上行得愚昧；因此，以後你必有戰爭。」
2CHR|16|10|亞撒 惱恨先見，為了這事向他發怒，將他囚在監裏。那時 亞撒 也虐待一些百姓。
2CHR|16|11|亞撒 自始至終的事蹟，看哪，都寫在《猶大和以色列諸王記》上。
2CHR|16|12|亞撒 作王三十九年的時候患了腳疾，非常嚴重。他生病的時候沒有求耶和華，只求醫生。
2CHR|16|13|他作王四十一年死了，與他祖先同睡，
2CHR|16|14|葬在 大衛城 自己所鑿的墳墓裏。人把他放在床上，床上堆滿各樣馨香的香料，就是按做香的作法調和的香料，又為他生一堆大火誌哀。
2CHR|17|1|亞撒 的兒子 約沙法 接續他作王，奮勇自強，防備 以色列 。
2CHR|17|2|他安置軍兵在 猶大 一切堅固城裏，又安置駐軍在 猶大 地和他父親 亞撒 所得 以法蓮 的城鎮中。
2CHR|17|3|耶和華與 約沙法 同在，因為他行他祖先 大衛 從前所行的道，不去尋求諸 巴力 ，
2CHR|17|4|只尋求他父親的上帝，遵行他的誡命，不效法 以色列 人的行為。
2CHR|17|5|所以耶和華堅定 約沙法 手中的國， 猶大 眾人給他進貢； 約沙法 大有財富和尊榮。
2CHR|17|6|他樂意遵行耶和華的道，並且從 猶大 再次除掉一切丘壇和 亞舍拉 。
2CHR|17|7|他作王第三年，差遣官員 便‧亥伊勒 、 俄巴底 、 撒迦利雅 、 拿坦業 、 米該亞 往 猶大 各城去教導百姓。
2CHR|17|8|跟他們一同去的有 利未 人 示瑪雅 、 尼探雅 、 西巴第雅 、 亞撒黑 、 示米拉末 、 約拿單 、 亞多尼雅 、 多比雅 、 駝‧巴多尼雅 ；跟他們一同的又有 以利沙瑪 和 約蘭 二位祭司。
2CHR|17|9|他們在 猶大 教導，帶著耶和華的律法書，走遍 猶大 各城教導百姓。
2CHR|17|10|猶大 四圍地上的邦國都懼怕耶和華，不敢與 約沙法 爭戰。
2CHR|17|11|有些 非利士 人送禮物，進貢銀子給 約沙法 。 阿拉伯 人也送他七千七百隻公綿羊，七千七百隻公山羊。
2CHR|17|12|約沙法 日漸強大，他在 猶大 建造堡壘和儲貨城。
2CHR|17|13|他在 猶大 城鎮中有許多工程，在 耶路撒冷 又有戰士，就是大能的勇士。
2CHR|17|14|他們按著父家的數目如下： 猶大 族的千夫長以 押拿 為首，率領三十萬大能的勇士；
2CHR|17|15|其次是 約哈難 千夫長，率領二十八萬；
2CHR|17|16|其次是 細基利 的兒子 亞瑪斯雅 ，他是一個自願奉獻給耶和華的人，率領二十萬大能的勇士。
2CHR|17|17|便雅憫 族有大能的勇士 以利雅大 ，率領二十萬拿弓箭和盾牌的人；
2CHR|17|18|其次是 約薩拔 ，率領十八萬預備打仗的人。
2CHR|17|19|這些都是伺候王的，還有王在全 猶大 的堅固城所安置的不在其內。
2CHR|18|1|約沙法 大有財富和尊榮，他與 亞哈 結親。
2CHR|18|2|過了幾年，他下到 撒瑪利亞 去見 亞哈 ； 亞哈 為他和跟從他的人宰了許多牛羊，勸他一同上去攻打 基列 的 拉末 。
2CHR|18|3|以色列 王 亞哈 問 猶大 王 約沙法 說：「你肯同我去攻打 基列 的 拉末 嗎？」他回答說：「你我不分彼此，我的軍隊就是你的軍隊，我們必與你一同去爭戰。」
2CHR|18|4|約沙法 對 以色列 王說：「請你先求問耶和華的話。」
2CHR|18|5|於是 以色列 王召集先知四百人，問他們說：「我可以上去攻打 基列 的 拉末 嗎？還是不要上去呢？」他們說：「可以上去，因為上帝必將那城交在王的手裏。」
2CHR|18|6|約沙法 說：「這裏還有沒有耶和華的先知，我們好求問他呢？」
2CHR|18|7|以色列 王對 約沙法 說：「還有一個人，是 音拉 的兒子 米該雅 ，我們可以託他求問耶和華。只是我真的很恨他，因為他對我說預言，從不說吉言，總是說凶信。」 約沙法 說：「請王不要這麼說。」
2CHR|18|8|以色列 王就召了一個官員來，說：「你快去，把 音拉 的兒子 米該雅 召來。」
2CHR|18|9|以色列 王和 猶大 王 約沙法 在 撒瑪利亞 城門前的禾場，各穿朝服，坐在寶座上，所有的先知都在他們面前說預言。
2CHR|18|10|基拿拿 的兒子 西底家 為自己造了鐵角，說：「耶和華如此說：『你要用這些角牴觸 亞蘭 人，直到將他們滅盡。』」
2CHR|18|11|所有的先知也都這樣預言說：「可以上 基列 的 拉末 去，必然得勝，因為耶和華必將那城交在王的手中。」
2CHR|18|12|那去召 米該雅 的使者對他說：「看哪，眾先知都異口同聲向王說吉言，你也跟他們說一樣的話，說吉言吧！」
2CHR|18|13|米該雅 說：「我指著永生的耶和華起誓，我的上帝說甚麼，我就說甚麼。」
2CHR|18|14|米該雅 來到王那裏，王問他：「 米該雅 啊，我們可以上去攻打 基列 的 拉末 嗎？還是不要上去呢？」他說：「可以上去，必然得勝，敵人必交在你們手裏。」
2CHR|18|15|王對他說：「我要你發誓多少次，你才會奉耶和華的名向我說實話呢？」
2CHR|18|16|米該雅 說：「我看見 以色列 眾人散佈在山上，如同沒有牧人的羊群一般。耶和華說：『這些人沒有主人，他們可以平安地各自回家去。』」
2CHR|18|17|以色列 王對 約沙法 說：「我豈沒有告訴你，這人對我說預言，從不說吉言，只說凶信嗎？」
2CHR|18|18|米該雅 說：「因此你們要聽耶和華的話！我看見耶和華坐在寶座上，天上的萬軍侍立在他左右。
2CHR|18|19|耶和華 說：『誰去引誘 以色列 王 亞哈 上 基列 的 拉末 去陣亡呢？』這個這樣說，那個那樣說。
2CHR|18|20|隨後有一個靈出來，站在耶和華面前，說：『我去引誘他。』耶和華問他：『用甚麼方法呢？』
2CHR|18|21|他說：『我要出去，在他眾先知的口中成為謊言的靈。』耶和華說：『這樣，你去引誘他，必能成功。你出去，照樣做吧！』
2CHR|18|22|現在，看哪，耶和華使謊言的靈入了你的這些先知的口，並且耶和華已經宣告要降禍於你。」
2CHR|18|23|基拿拿 的兒子 西底家 前來打 米該雅 一巴掌，說：「耶和華的靈從哪裏離開我向你說話呢？」
2CHR|18|24|米該雅 說：「看哪，你進入嚴密的內室躲藏的那日，就必看見。」
2CHR|18|25|以色列 王說：「把 米該雅 帶走，交回給 亞們 市長和 約阿施 王子。
2CHR|18|26|你們要說：『王如此說：把這個人關在監獄裏，使他受苦，吃不飽喝不足，直等到我平安回來。』」
2CHR|18|27|米該雅 說：「你若真的能平安回來，那就是耶和華沒有藉我說話了。」他又說：「眾百姓啊，你們都要聽！」
2CHR|18|28|以色列 王和 猶大 王 約沙法 上 基列 的 拉末 去。
2CHR|18|29|以色列 王對 約沙法 說：「我要改裝上陣，你可以仍穿王服。」於是 以色列 王改裝，他們上陣去了。
2CHR|18|30|亞蘭 王吩咐他的戰車長說：「你們不要與他們的大將或小兵交戰，只要單單攻擊 以色列 王。」
2CHR|18|31|那些戰車長看見 約沙法 就說：「這一定是 以色列 王！」他們轉過去與他交戰。 約沙法 一呼喊，耶和華就幫助他，上帝使他們轉離他。
2CHR|18|32|戰車長見他不是 以色列 王，就轉身不追他了。
2CHR|18|33|有一人開弓，並不知情，箭恰巧射入 以色列 王鎧甲的縫裏。王對駕車的說：「我受重傷了，你掉過車來，載我離開戰場！」
2CHR|18|34|那日，戰況越來越猛， 以色列 王勉強站在戰車上，面對 亞蘭 人，直到傍晚。日落的時候，王就死了。
2CHR|19|1|猶大 王 約沙法 平安回 耶路撒冷 ，到自己的宮裏。
2CHR|19|2|哈拿尼 的兒子 耶戶 先見出來迎接 約沙法 王，對他說：「你怎麼可以幫助惡人，愛那恨耶和華的人呢？因此耶和華的憤怒臨到你了。
2CHR|19|3|然而你還有善行，因你從國中除掉 亞舍拉 ，立定心意尋求上帝。」
2CHR|19|4|約沙法 住在 耶路撒冷 ，以後又出巡民間，從 別是巴 直到 以法蓮 山區，引導百姓歸向耶和華－他們列祖的上帝。
2CHR|19|5|他在國中，在 猶大 一切堅固城設立審判官，各城都是如此。
2CHR|19|6|他對審判官說：「你們應當謹慎所做的事，因為你們審判不是為人，而是為耶和華。在審判的事上，他必與你們同在。
2CHR|19|7|現在，你們應當敬畏耶和華，謹慎辦事，因為耶和華－我們的上帝沒有不義，不看人的情面，也不受賄賂。」
2CHR|19|8|約沙法 從 利未 人和祭司，以及 以色列 族長中，也委派人在 耶路撒冷 為耶和華施行審判，為 耶路撒冷 的居民聽訟斷案 。
2CHR|19|9|約沙法 吩咐他們說：「你們當這樣，以敬畏耶和華、誠實和純正的心辦事。
2CHR|19|10|你們住在各城的弟兄，若有爭訟的案件呈到你們這裏，或為流血，或犯律法、誡命、律例、典章，你們要警戒他們，免得他們得罪耶和華，以致憤怒臨到你們和你們的弟兄；你們當這樣行，就沒有罪了。
2CHR|19|11|看哪，凡屬耶和華的事，有 亞瑪利雅 祭司長管理你們；凡屬王的事，有 猶大 家的領袖 以實瑪利 的兒子 西巴第雅 管理你們；在你們面前有 利未 人作官長。你們應當壯膽辦事，願耶和華與善人同在。」
2CHR|20|1|此後， 摩押 人和 亞捫 人，連同一些 米烏尼 人 來攻擊 約沙法 。
2CHR|20|2|有人來報告 約沙法 說：「從海的那邊， 以東 有大軍來攻擊你，看哪，他們在 哈洗遜‧他瑪 ，就是 隱‧基底 。」
2CHR|20|3|約沙法 懼怕，就定意尋求耶和華，在全 猶大 宣告禁食。
2CHR|20|4|於是 猶大 人聚集，求耶和華幫助，甚至他們從 猶大 各城前來尋求耶和華。
2CHR|20|5|約沙法 站在 猶大 和 耶路撒冷 的會眾中，在耶和華殿新的院子前，
2CHR|20|6|說：「耶和華－我們列祖的上帝啊，你不是天上的上帝嗎？你不是萬邦萬國的主宰嗎？在你手中有大能大力，無人能抵擋你。
2CHR|20|7|我們的上帝啊，你不是曾在你百姓 以色列 面前驅逐這地的居民，將這地賜給你朋友 亞伯拉罕 的後裔永遠為業嗎？
2CHR|20|8|他們住在這地，又為你的名建造聖所，說：
2CHR|20|9|『若有禍患臨到我們，或刀兵的懲罰，或瘟疫饑荒，我們在急難的時候，站在這殿前向你呼求，你必垂聽並且拯救，因為你的名在這殿裏。』
2CHR|20|10|現在，看哪， 以色列 人出 埃及 地的時候，你不容許 以色列 人侵犯 亞捫 人、 摩押 人和 西珥山 人， 以色列 人就離開他們，不滅絕他們。
2CHR|20|11|看哪，他們這樣回報我們，要來驅逐我們離開你賜給我們為業之地。
2CHR|20|12|我們的上帝啊，你不懲罰他們嗎？因為我們無力抵擋這來攻擊我們的大軍。我們不知道該怎麼做，我們的眼目單仰望你。」
2CHR|20|13|猶大 眾人和他們的孩童、妻子、兒女都站在耶和華面前。
2CHR|20|14|那時，耶和華的靈在會眾中臨到 利未 人 亞薩 的後裔 雅哈悉 ，他是 瑪探雅 的玄孫， 耶利 的曾孫， 比拿雅 的孫子， 撒迦利雅 的兒子。
2CHR|20|15|他說：「 猶大 眾人、 耶路撒冷 的居民和 約沙法 王啊，你們要留心聽，耶和華對你們如此說：『不要因這大軍恐懼驚惶，因為勝敗不在乎你們，而是在乎上帝。
2CHR|20|16|明日你們要下去迎敵；看哪，他們從 洗斯坡 上來，你們必在 耶魯伊勒 曠野前的谷口遇見他們。
2CHR|20|17|猶大 和 耶路撒冷 人哪，這次你們不要爭戰，要擺陣站著，看耶和華為你們施行拯救。不要恐懼，也不要驚惶。明日當出去迎敵，因為耶和華與你們同在。』」
2CHR|20|18|約沙法 屈身，臉伏於地， 猶大 眾人和 耶路撒冷 的居民也俯伏在耶和華面前，敬拜耶和華。
2CHR|20|19|哥轄 子孫和 可拉 子孫的 利未 人都起來，用極大的聲音讚美耶和華－ 以色列 的上帝。
2CHR|20|20|清晨，眾人早起往 提哥亞 的曠野去。出去的時候， 約沙法 站著說：「 猶大 人和 耶路撒冷 的居民哪，要聽我說：信靠耶和華－你們的上帝就必站立得穩；信賴他的先知就必亨通。」
2CHR|20|21|約沙法 與百姓商議，就設立歌唱的人，頌讚耶和華，使他們穿上聖潔的禮服，走在軍隊前讚美耶和華： 「當稱謝耶和華， 因他的慈愛永遠長存！」
2CHR|20|22|他們開始唱歌讚美的時候，耶和華派伏兵擊殺那來攻擊 猶大 的 亞捫 人、 摩押 人和 西珥山 人，他們就被打敗了。
2CHR|20|23|亞捫 人和 摩押 人起來，擊殺住 西珥山 的人，把他們滅盡；滅盡住 西珥山 的人之後，他們又彼此自相擊殺。
2CHR|20|24|猶大 人來到曠野的瞭望樓，向那大軍觀看，看哪，遍地都是屍體，沒有一個逃脫的。
2CHR|20|25|約沙法 和他的百姓就來收取掠物，找到許多牲畜 、財物、衣服 和珍寶。他們取掠物歸為己有，直到無法攜帶；因為掠物太多，他們足足收取了三日。
2CHR|20|26|第四日，眾人聚集在 比拉迦谷 ，在那裏稱頌耶和華；因此那地方名叫 比拉迦谷 ，直到今日。
2CHR|20|27|在 約沙法 率領下， 猶大 人和 耶路撒冷 人都歡歡喜喜地回 耶路撒冷 ，耶和華使他們因戰勝仇敵而喜樂。
2CHR|20|28|他們彈琴、鼓瑟、吹號來到 耶路撒冷 ，進了耶和華的殿。
2CHR|20|29|地上所有的邦國聽見耶和華打敗 以色列 的仇敵，就都懼怕上帝。
2CHR|20|30|這樣， 約沙法 的國得享太平，因為上帝賜他四境平安。
2CHR|20|31|約沙法 作 猶大 王，登基的時候年三十五歲，在 耶路撒冷 作王二十五年。他母親名叫 阿蘇巴 ，是 示利希 的女兒。
2CHR|20|32|約沙法 效法他父親 亞撒 所行的道，不偏離左右，行耶和華眼中看為正的事。
2CHR|20|33|只是丘壇還沒有廢去，百姓也沒有立定心意歸向他們列祖的上帝。
2CHR|20|34|約沙法 其餘的事，看哪，自始至終都寫在 哈拿尼 的兒子 耶戶 的書上，這些事也記載在《以色列諸王記》上。
2CHR|20|35|此後， 猶大 王 約沙法 與 以色列 王 亞哈謝 結盟； 亞哈謝 多行惡事。
2CHR|20|36|他們合夥造船要往 他施 去，就在 以旬‧迦別 造船。
2CHR|20|37|瑪利沙 人 多大瓦 的兒子 以利以謝 向 約沙法 預言說：「因你與 亞哈謝 結盟，耶和華必破壞你所造的。」後來那些船果然毀壞，不能往 他施 去了。
2CHR|21|1|約沙法 與他祖先同睡，與他祖先同葬在 大衛城 ，他的兒子 約蘭 接續他作王。
2CHR|21|2|約蘭 有幾個兄弟，就是 約沙法 的兒子 亞撒利雅 、 耶歇 、 撒迦利雅 、 亞撒列夫 、 米迦勒 、 示法提雅 ；這些都是 以色列 王 約沙法 的兒子。
2CHR|21|3|他們的父親把許多禮物，金銀財寶和 猶大 的堅固城賜給他們，卻把國賜給 約蘭 ，因為他是長子。
2CHR|21|4|約蘭 起來治理他父親的國，奮勇自強，用刀殺了他所有的兄弟和 以色列 的幾個領袖。
2CHR|21|5|約蘭 登基的時候年三十二歲，在 耶路撒冷 作王八年。
2CHR|21|6|他行 以色列 諸王的道，正如 亞哈 家所行的，因他娶了 亞哈 的女兒為妻，行耶和華眼中看為惡的事。
2CHR|21|7|耶和華卻因自己與 大衛 所立的約，不肯滅絕 大衛 的家，要照他所應許的，永遠賜燈光給 大衛 和他的子孫。
2CHR|21|8|約蘭 在位期間， 以東 背叛，自己立王治理他們，脫離 猶大 的權勢。
2CHR|21|9|約蘭 就率領他的軍官和所有的戰車過去。他夜間起來，攻打圍困他的 以東 人和戰車長。
2CHR|21|10|這樣， 以東 背叛，脫離 猶大 的權勢，直到今日。那時， 立拿 也背叛了，脫離它的權勢，因為 約蘭 離棄耶和華－他列祖的上帝。
2CHR|21|11|他又在 猶大 山嶺 建造丘壇，使 耶路撒冷 的居民行淫，誘惑 猶大 。
2CHR|21|12|以利亞 先知寫信給 約蘭 說：「耶和華－你祖先 大衛 的上帝如此說：『因為你不行你父 約沙法 和 猶大 王 亞撒 的道，
2CHR|21|13|反而行 以色列 諸王的道，使 猶大 和 耶路撒冷 居民行淫，像 亞哈 家行淫一樣，又殺了你父家比你好的那些兄弟。
2CHR|21|14|看哪，耶和華必降大災於你的百姓和你的妻妾、兒女，以及你一切所有的。
2CHR|21|15|至於你，你必患許多的病 ，你的腸子也必生許多的病，日漸沉重，直到腸子墜落下來。』」
2CHR|21|16|耶和華激發 非利士 人和靠近 古實 人的 阿拉伯 人的心來攻擊 約蘭 。
2CHR|21|17|他們上來攻擊 猶大 ，侵入境內，擄掠了王宮裏所有的財物和他的妻妾、兒女，除了他的小兒子 約哈斯 之外，沒有留下一個兒子。
2CHR|21|18|這一切事以後，耶和華擊打 約蘭 ，使他的腸子患不能醫治的病。
2CHR|21|19|這病纏綿日久，過了二年，腸子墜落下來，他就病重而死。他的百姓沒有為他生火誌哀，像從前為他祖先生火一樣。
2CHR|21|20|約蘭 登基的時候年三十二歲，在 耶路撒冷 作王八年。他逝世無人思慕，眾人把他葬在 大衛城 ，只是不在列王的墳墓裏。
2CHR|22|1|耶路撒冷 的居民立 約蘭 的小兒子 亞哈謝 接續他作王，因為跟隨 阿拉伯 人來攻營的軍兵把 亞哈謝 所有的兄長都殺了； 猶大 王 約蘭 的兒子 亞哈謝 就作了王。
2CHR|22|2|亞哈謝 登基的時候年四十二歲 ，在 耶路撒冷 作王一年。他母親名叫 亞她利雅 ，是 暗利 的孫女。
2CHR|22|3|亞哈謝 也行 亞哈 家的道，因為他母親給他主謀，使他行惡。
2CHR|22|4|他行耶和華眼中看為惡的事，像 亞哈 家一樣；因他父親死後，他們給他主謀，使他敗壞。
2CHR|22|5|他也聽從他們的計謀，與 以色列 王 亞哈 的兒子 約蘭 同往 基列 的 拉末 去，與 亞蘭 王 哈薛 交戰。 亞蘭 人打傷了 約蘭 ，
2CHR|22|6|他回到 耶斯列 ，醫治在 拉末 與 亞蘭 王 哈薛 打仗時被擊打所受的傷。 約蘭 的兒子 猶大 王 亞哈謝 因為 亞哈 的兒子 約蘭 病了，就下到 耶斯列 看望他。
2CHR|22|7|亞哈謝 去見 約蘭 而遇害，這是出乎上帝；因為他一到就同 約蘭 出去攻擊 寧示 的孫子 耶戶 ；這 耶戶 是耶和華所膏，使他剪除 亞哈 家的。
2CHR|22|8|耶戶 向 亞哈 家施行懲罰的時候，遇見 猶大 的眾領袖和 亞哈謝 的姪子們正服事 亞哈謝 ，就把他們都殺了。
2CHR|22|9|亞哈謝 躲在 撒瑪利亞 ， 耶戶 尋找他，眾人把他拿住，送到 耶戶 那裏，就殺了他。他們把他埋葬，因他們說，他是那盡心尋求耶和華之 約沙法 的兒子。這樣， 亞哈謝 的家無力保住國權。
2CHR|22|10|亞哈謝 的母親 亞她利雅 見她兒子死了，就起來剿滅 猶大 王室所有的後裔。
2CHR|22|11|但王的女兒 約示巴 將 亞哈謝 的兒子 約阿施 從那被殺的王子中偷出來，把他和他的奶媽藏在臥房裏。 約示巴 是 約蘭 王的女兒， 亞哈謝 的妹妹，祭司 耶何耶大 的妻子。她藏了 約阿施 ，躲避 亞她利雅 ，免受殺害。
2CHR|22|12|亞她利雅 治理這地的時候， 約阿施 和他們一同在上帝殿裏藏了六年。
2CHR|23|1|第七年， 耶何耶大 奮勇自強，叫了 耶羅罕 的兒子 亞撒利雅 、 約哈難 的兒子 以實瑪利 、 俄備得 的兒子 亞撒利雅 、 亞大雅 的兒子 瑪西雅 ，和 細基利 的兒子 以利沙法 等眾百夫長，與他們立約。
2CHR|23|2|他們走遍 猶大 ，從 猶大 各城召集 利未 人和 以色列 的眾族長到 耶路撒冷 來。
2CHR|23|3|全會眾在上帝殿裏與王立約。 耶何耶大 對他們說：「看哪，王的兒子必作王，正如耶和華指著 大衛 子孫所應許的。
2CHR|23|4|你們要這樣做：在安息日值班的祭司和 利未 人，三分之一要把守各門，
2CHR|23|5|三分之一要在王宮，三分之一要在 根基門 ；眾百姓都要在耶和華殿的院內。
2CHR|23|6|除了祭司和供職的 利未 人之外，不准別人進耶和華的殿；只有他們可以進去，因為他們是神聖的。眾百姓都要遵守耶和華所吩咐的。
2CHR|23|7|利未 人要手中各拿兵器，四圍保護王；凡擅自進殿的，要被處死。王出入的時候，你們當跟隨他。」
2CHR|23|8|利未 人和 猶大 眾人都照著 耶何耶大 祭司一切所吩咐的去做，各帶自己的人，無論安息日值班或不值班的都來，因為 耶何耶大 祭司不許他們下班。
2CHR|23|9|耶何耶大 祭司就把上帝殿裏所藏 大衛 王的槍和大小盾牌交給百夫長，
2CHR|23|10|又分派眾百姓手中各拿兵器，在祭壇和殿那裏，從殿南到殿北，站在王的四圍；
2CHR|23|11|他們領 約阿施 出來，給他戴上冠冕，把律法書交給他，立他作王。 耶何耶大 和他的兒子們膏他，他們說：「願王萬歲！」
2CHR|23|12|亞她利雅 聽見百姓奔走讚美王的聲音，就進耶和華的殿，到百姓那裏。
2CHR|23|13|她觀看，看哪，王站在殿門的柱旁，百夫長和號手在王旁邊，國中的眾百姓都歡樂吹號，又有歌唱的人用樂器領人歌唱讚美。 亞她利雅 就撕裂衣服，喊著說：「反了！反了！」
2CHR|23|14|耶何耶大 祭司帶領管軍兵的百夫長出來，對他們說：「把她從行列之間趕出去，凡跟隨她的必用刀殺死！」因為祭司說：「不可在耶和華殿裏殺她。」
2CHR|23|15|他們就下手拿住她；她進入通往王宮的 馬門 ，他們就在那裏把她殺了。
2CHR|23|16|耶何耶大 與眾百姓，又與王立約，要作耶和華的子民。
2CHR|23|17|於是眾百姓到 巴力 廟去，拆毀了廟，打碎祭壇和偶像，又在壇前把 巴力 的祭司 瑪坦 殺了。
2CHR|23|18|耶何耶大 派官員在 利未 家的祭司手下看守耶和華的殿，他們是 大衛 所分派的，在耶和華殿中照 摩西 律法上所寫，獻燔祭給耶和華，又按 大衛 所定的，歡樂歌唱。
2CHR|23|19|耶何耶大 又設立守衛把守耶和華殿的各門，無論因何事而不潔淨的人，都不准進去。
2CHR|23|20|他又率領百夫長和貴族，與民間的官長，以及國中的眾百姓，請王從耶和華的殿下來，由 上門 正中進入王宮，使王坐在國度的王位上。
2CHR|23|21|國中的眾百姓都歡樂，合城也都平靜。他們已將 亞她利雅 用刀殺了。
2CHR|24|1|約阿施 登基的時候年方七歲，在 耶路撒冷 作王四十年。他母親名叫 西比亞 ，是 別是巴 人。
2CHR|24|2|耶何耶大 祭司在世的日子， 約阿施 行耶和華眼中看為正的事。
2CHR|24|3|耶何耶大 為他娶了兩個妻子，他生兒育女。
2CHR|24|4|此後， 約阿施 有心重修耶和華的殿，
2CHR|24|5|就召集祭司和 利未 人，吩咐他們說：「你們要往 猶大 各城去，向 以色列 眾人徵收銀子，按每年的需要整修你們上帝的殿；你們要急速辦理這事。」但 利未 人沒有急速辦理。
2CHR|24|6|王召了 耶何耶大 祭司長來，對他說：「從前耶和華的僕人 摩西 ，為法櫃的帳幕與 以色列 會眾所定的捐獻，你為何不叫 利未 人照這例向 猶大 和 耶路撒冷 徵收呢？」
2CHR|24|7|因為那惡婦 亞她利雅 的兒子們曾拆毀上帝的殿，又用耶和華殿中分別為聖的物供奉諸 巴力 。
2CHR|24|8|於是王下令造一個櫃子，放在耶和華殿的門外，
2CHR|24|9|又通告 猶大 和 耶路撒冷 ，要將上帝僕人 摩西 在曠野所吩咐 以色列 的捐獻送來給耶和華。
2CHR|24|10|眾領袖和百姓都歡歡喜喜帶捐獻來，投入櫃中，直到投滿。
2CHR|24|11|利未 人見銀子多了，把櫃子抬到王所派的官長面前；這時王的書記和祭司長的助手就會來把櫃子倒空，然後放回原處。日日都是這樣做，積蓄的銀子很多。
2CHR|24|12|王與 耶何耶大 把銀子交給耶和華殿裏辦事的人，他們就雇了石匠、木匠重修耶和華的殿，又雇了鐵匠、銅匠整修耶和華的殿。
2CHR|24|13|工人做工，修理工程在他們手中漸漸完成，他們將上帝的殿修理得如同從前一樣，非常堅固。
2CHR|24|14|他們做完了，就把多餘的銀子拿到王與 耶何耶大 面前，用以製造耶和華殿供奉所用的器皿和調羹，以及金銀的器皿。 耶何耶大 在世的日子，眾人經常在耶和華殿裏獻燔祭。
2CHR|24|15|耶何耶大 年紀老邁，日子滿足而死，死的時候年一百三十歲。
2CHR|24|16|眾人把他與列王同葬在 大衛城 ，因為他在 以色列 中為上帝和他的殿做了美善的事。
2CHR|24|17|耶何耶大 死後， 猶大 的眾領袖來叩拜王，那時王就聽了他們。
2CHR|24|18|他們離棄耶和華－他們列祖上帝的殿，去事奉 亞舍拉 和偶像；因他們這罪，就有憤怒臨到 猶大 和 耶路撒冷 。
2CHR|24|19|但上帝仍差遣先知到他們那裏，引導他們歸向耶和華。先知警戒他們，他們卻不肯聽。
2CHR|24|20|那時，上帝的靈感動 耶何耶大 的兒子 撒迦利亞 祭司，他就站在上面，對百姓說：「上帝如此說：『你們為何干犯耶和華的誡命，以致不得亨通呢？因為你們離棄耶和華，所以他也離棄你們。』」
2CHR|24|21|眾人謀害 撒迦利亞 ，照著王的吩咐，在耶和華殿的院內用石頭打死他。
2CHR|24|22|這樣， 約阿施 王不記念 撒迦利亞 的父親 耶何耶大 向自己所施的恩，殺了他的兒子。 撒迦利亞 臨死的時候說：「願耶和華鑒察伸冤！」
2CHR|24|23|年底的時候， 亞蘭 的軍兵上來攻擊 約阿施 ，來到 猶大 和 耶路撒冷 ，殺了百姓中的眾領袖，把所掠取的財物全送到 大馬士革 王那裏。
2CHR|24|24|亞蘭 的軍兵雖只來了一小隊人，耶和華卻將極大的軍隊交在他們手裏；因為 猶大 人離棄耶和華－他們列祖的上帝，所以 亞蘭 人懲罰 約阿施 。
2CHR|24|25|亞蘭 人離開 約阿施 的時候，他患重病 ；他的臣僕背叛他，要報 耶何耶大 祭司兒子 的流血之仇，在床上殺了他。他就死了，葬在 大衛城 ，只是不葬在列王的墳墓裏。
2CHR|24|26|背叛他的是 亞捫 婦人 示米押 的兒子 撒拔 和 摩押 婦人 示米利 的兒子 約薩拔 。
2CHR|24|27|至於他的兒子們和他所受的眾多警戒，以及他重修上帝殿的事，看哪，都寫在《列王評傳》上。他的兒子 亞瑪謝 接續他作王。
2CHR|25|1|亞瑪謝 登基的時候年二十五歲，在 耶路撒冷 作王二十九年。他母親名叫 約耶但 ，是 耶路撒冷 人。
2CHR|25|2|亞瑪謝 行耶和華眼中看為正的事，只是沒有純正的心。
2CHR|25|3|他的王國一鞏固，就把殺他父王的臣僕殺了，
2CHR|25|4|卻沒有處死他們的兒子，這是照 摩西 律法書上耶和華所吩咐的說：「不可因子殺父，也不可因父殺子，各人要為自己的罪而死。」
2CHR|25|5|亞瑪謝 召集 猶大 人，按著父家為全 猶大 和 便雅憫 設立千夫長、百夫長，又數點人數，從二十歲以上，能拿槍拿盾牌出去打仗的精兵共有三十萬；
2CHR|25|6|又用一百他連得銀子，從 以色列 招募了十萬大能的勇士。
2CHR|25|7|有一個神人來見 亞瑪謝 ，對他說：「王啊，不要帶領 以色列 的軍兵與你同去，因為耶和華不和 以色列 ，和任何 以法蓮 的子孫同在。
2CHR|25|8|你若一定要去，就奮勇作戰吧！但上帝必使你敗在敵人面前，因為上帝能助人得勝，也能使人落敗。」
2CHR|25|9|亞瑪謝 問神人：「我給了 以色列 軍隊的那一百他連得銀子怎麼樣呢？」神人回答：「耶和華會把比這些更多的賜給你。」
2CHR|25|10|於是 亞瑪謝 把那從 以法蓮 來的軍兵分別出來，叫他們到自己的地方去。他們非常惱怒 猶大 ，氣憤地回自己的地方去了。
2CHR|25|11|亞瑪謝 壯起膽來，率領他的軍隊到 鹽谷 ，殺了一萬 西珥 人。
2CHR|25|12|猶大 人又生擒了一萬人，把他們帶到 西拉 山頂上，從 西拉 山頂扔下去，把他們全都摔碎了。
2CHR|25|13|但 亞瑪謝 所打發回去、不許一同出征的那些軍兵劫掠 猶大 各城，從 撒瑪利亞 直到 伯‧和崙 ，殺了三千人，搶了許多財物。
2CHR|25|14|亞瑪謝 擊殺 以東 人回來以後，他把 西珥 人的神像帶回，立為自己的神明，在它們面前叩拜燒香。
2CHR|25|15|耶和華的怒氣向 亞瑪謝 發作，差派一個先知去見他，對他說：「這些神明不能救自己的百姓脫離你的手，你為何尋求它們呢？」
2CHR|25|16|先知與王說話的時候，王對他說：「難道我們立你作王的謀士嗎？你住口吧！為何要挨打呢？」先知就止住了，卻說：「我知道上帝已定意要消滅你，因為你行這事，不聽從我的勸戒。」
2CHR|25|17|猶大 王 亞瑪謝 經商議後，就派人去見 耶戶 的孫子， 約哈斯 的兒子 以色列 王 約阿施 ，說：「來，讓我們面對面較量吧！」
2CHR|25|18|以色列 王 約阿施 派人去見 猶大 王 亞瑪謝 ，說：「 黎巴嫩 的蒺藜派人去見 黎巴嫩 的香柏樹，說：『將你的女兒嫁給我的兒子。』但有一隻野獸經過 黎巴嫩 ，把蒺藜踐踏了。
2CHR|25|19|你說，看哪，你打敗了 以東 ，就心高氣傲，以此為榮。現在，你待在家裏算了吧，為何要惹禍使自己和 猶大 一同敗亡呢？」
2CHR|25|20|亞瑪謝 卻不肯聽從。這是出乎上帝，好將他們交在敵人手裏，因為他們尋求 以東 的神明。
2CHR|25|21|於是 以色列 王 約阿施 上來，在 猶大 的 伯‧示麥 與 猶大 王 亞瑪謝 面對面較量。
2CHR|25|22|猶大 敗在 以色列 面前，他們逃跑，各人逃回自己的帳棚去了。
2CHR|25|23|以色列 王 約阿施 在 伯‧示麥 擒住 約哈斯 的孫子， 約阿施 的兒子 猶大 王 亞瑪謝 ，把他帶到 耶路撒冷 ，又拆毀 耶路撒冷 的城牆，從 以法蓮門 直到 角門 共四百肘。
2CHR|25|24|他帶著 俄別‧以東 所看守上帝殿裏的一切金銀和器皿，與王宮裏的財寶，又帶著人質，回 撒瑪利亞 去了。
2CHR|25|25|約哈斯 的兒子 以色列 王 約阿施 死後， 猶大 王 約阿施 的兒子 亞瑪謝 又活了十五年。
2CHR|25|26|亞瑪謝 其餘的事，自始至終，看哪，不都寫在《猶大和以色列諸王記》上嗎？
2CHR|25|27|自從 亞瑪謝 離棄耶和華之後，在 耶路撒冷 有人背叛他，他就逃往 拉吉 ；他們卻派人追到 拉吉 ，在那裏殺了他。
2CHR|25|28|有人用馬將他馱回，把他與祖先一同葬在 猶大 的城 。
2CHR|26|1|猶大 眾百姓立 烏西雅 接續他父親 亞瑪謝 作王，那時他年十六歲。
2CHR|26|2|亞瑪謝 王與他祖先同睡之後， 烏西雅 收復 以祿 回歸 猶大 ，又重新修建。
2CHR|26|3|烏西雅 登基的時候年十六歲，在 耶路撒冷 作王五十二年。他母親名叫 耶可利雅 ，是 耶路撒冷 人。
2CHR|26|4|烏西雅 行耶和華眼中看為正的事，效法他父親 亞瑪謝 一切所行的。
2CHR|26|5|撒迦利亞 是一個通曉上帝默示的人 ，他在世的日子， 烏西雅 定意尋求上帝； 烏西雅 尋求耶和華的日子，上帝使他亨通。
2CHR|26|6|他出去攻擊 非利士 人，拆毀了 迦特 、 雅比尼 和 亞實突 的城牆，又在 非利士 人中，在 亞實突 境內建築城鎮。
2CHR|26|7|上帝幫助他攻擊 非利士 人和住在 姑珥‧巴力 的 阿拉伯 人，以及 米烏尼 人。
2CHR|26|8|米烏尼 人 向 烏西雅 進貢。他的名聲傳到 埃及 ，因他非常強盛。
2CHR|26|9|烏西雅 在 耶路撒冷 的 角門 和 谷門 ，以及城牆轉角之處建築城樓，非常堅固。
2CHR|26|10|他在曠野建築瞭望樓，又挖了許多井，因為他在 謝非拉 和平原有很多牲畜。他在山區和肥沃的土地雇用耕種田地和修整葡萄園的人，因為他喜愛土地。
2CHR|26|11|烏西雅 又有軍兵，照書記 耶利 和官長 瑪西雅 所數點的，在王的一個將軍 哈拿尼雅 手下，分隊出戰。
2CHR|26|12|族長和大能勇士的總數共二千六百人，
2CHR|26|13|他們手下的軍兵共三十萬七千五百人，都大有能力，善於作戰，幫助王攻擊仇敵。
2CHR|26|14|烏西雅 為全軍預備盾牌、頭盔、鎧甲、槍、弓和甩石的機弦，
2CHR|26|15|又在 耶路撒冷 叫巧匠設計機器，安在城樓和角樓上，用以射箭，投擲大石。 烏西雅 的名聲傳到遠方，因為他得了非凡的幫助，極其強盛。
2CHR|26|16|烏西雅 既強盛，就心高氣傲，以致敗壞。他干犯耶和華－他的上帝，進耶和華的殿，要在香壇上燒香。
2CHR|26|17|亞撒利雅 祭司率領八十名勇敢的耶和華的祭司，跟隨他進去。
2CHR|26|18|他們阻止 烏西雅 王，對他說：「 烏西雅 啊，給耶和華燒香不是你的事，而是 亞倫 子孫的事，他們是分別為聖來燒香的祭司。你出聖殿吧！因為你犯了罪，耶和華上帝必不使你得尊榮。」
2CHR|26|19|烏西雅 發怒，手拿香爐要燒香。他在耶和華殿中香壇旁向眾祭司發怒的時候，他的額頭在眾祭司面前忽然長出痲瘋 。
2CHR|26|20|亞撒利雅 祭司長和眾祭司轉向他，看哪，他的額頭長出痲瘋，就催他離開那裏；他自己也急速出去，因為耶和華降災於他。
2CHR|26|21|烏西雅 王患痲瘋直到死的那日；他因為染上痲瘋，就住在隔離的行宮裏，與耶和華的殿隔絕。他兒子 約坦 管理王的家，治理這地的百姓。
2CHR|26|22|烏西雅 其餘的事，自始至終， 亞摩斯 的兒子 以賽亞 先知都記錄下來。
2CHR|26|23|烏西雅 與他祖先同睡，與他祖先同葬在田間的王陵；因為人說，他是長痲瘋的。他的兒子 約坦 接續他作王。
2CHR|27|1|約坦 登基的時候年二十五歲，在 耶路撒冷 作王十六年。他母親名叫 耶路沙 ，是 撒督 的女兒。
2CHR|27|2|約坦 行耶和華眼中看為正的事，效法他父親 烏西雅 一切所行的，只是他不入耶和華的殿。百姓仍舊行敗壞的事。
2CHR|27|3|約坦 建造耶和華殿的 上門 ，在 俄斐勒 城牆上有很多建設，
2CHR|27|4|又在 猶大 山區建造城鎮，在樹林中建築營寨和瞭望樓。
2CHR|27|5|約坦 與 亞捫 人的王打仗，勝了他們。那年 亞捫 人向他進貢一百他連得銀子，一萬歌珥小麥，一萬歌珥大麥；第二年、第三年 亞捫 人也這樣做。
2CHR|27|6|約坦 日漸強盛，因為他在耶和華－他上帝面前行正道。
2CHR|27|7|約坦 其餘的事和一切戰役，以及他的行為，看哪，都寫在《以色列和猶大列王記》上。
2CHR|27|8|他登基的時候年二十五歲，在 耶路撒冷 作王十六年。
2CHR|27|9|約坦 與他祖先同睡，葬在 大衛城 ，他兒子 亞哈斯 接續他作王。
2CHR|28|1|亞哈斯 登基的時候年二十歲，在 耶路撒冷 作王十六年。他不像他祖先 大衛 行耶和華眼中看為正的事，
2CHR|28|2|卻行 以色列 諸王的道，又鑄造諸 巴力 的像，
2CHR|28|3|照著耶和華從 以色列 人面前趕出的外邦人所行可憎的事，在 欣嫩子谷 燒香，用火焚燒他的兒女，
2CHR|28|4|又在丘壇上、山岡上、各青翠樹下獻祭燒香。
2CHR|28|5|耶和華－他的上帝將他交在 亞蘭 王手裏。 亞蘭 王打敗他，從他擄走了許多人，帶到 大馬士革 去。上帝又將他交在 以色列 王手裏， 以色列 王向他大行殺戮。
2CHR|28|6|利瑪利 的兒子 比加 一日之內在 猶大 殺了十二萬人，都是勇士，因為他們離棄了耶和華－他們列祖的上帝。
2CHR|28|7|有一個叫 細基利 的 以法蓮 勇士，殺了 瑪西雅 王子、 押斯利甘 宮廷總管和 以利加拿 宰相。
2CHR|28|8|以色列 人擄了他們的弟兄，連婦人帶兒女共二十萬，又掠取了許多財物，把這些掠物帶到 撒瑪利亞 去。
2CHR|28|9|但那裏有耶和華的一個先知，名叫 俄德 ，出來迎接往 撒瑪利亞 去的軍兵，對他們說：「看哪，耶和華－你們列祖的上帝惱怒 猶大 人，將他們交在你們手裏，你們竟怒氣沖天，向他們大行殺戮。
2CHR|28|10|如今你們又有意強逼 猶大 人和 耶路撒冷 人作你們的奴婢，你們豈不是也得罪了耶和華－你們的上帝嗎？
2CHR|28|11|現在你們當聽我說，要將從你們弟兄中擄來的釋放回去，因耶和華的烈怒已臨到你們了。」
2CHR|28|12|於是， 以法蓮 人的幾個領袖，就是 約哈難 的兒子 亞撒利雅 、 米實利末 的兒子 比利家 、 沙龍 的兒子 耶希西家 、 哈得萊 的兒子 亞瑪撒 ，起來攔阻從戰場上回來的人，
2CHR|28|13|對他們說：「你們不可把這些被擄的人帶到這裏，因我們已經得罪耶和華了。你們還想加增我們的罪惡過犯嗎？因為我們的罪過深重，已經有烈怒臨到 以色列 了。」
2CHR|28|14|於是帶兵器的人將擄來的人口和掠取的財物都留在眾領袖和全會眾面前。
2CHR|28|15|以上提名的那些人就起來，照顧被擄的人；其中凡赤身的，就從所掠取的財物中拿出衣服和鞋來，給他們穿，又給他們吃喝，用膏抹他們；其中凡軟弱的，就使他們騎驢，送到棕樹城 耶利哥 他們弟兄那裏。然後，他們就回 撒瑪利亞 去了。
2CHR|28|16|那時， 亞哈斯 王派人去求 亞述 諸王 來幫助他，
2CHR|28|17|因為 以東 人又來攻擊 猶大 ，擄掠俘虜。
2CHR|28|18|非利士 人也來侵佔 謝非拉 和 猶大 的 尼革夫 的城鎮，攻取了 伯‧示麥 、 亞雅崙 、 基低羅 、 梭哥 和所屬的鄉鎮、 亭拿 和所屬的鄉鎮、 瑾鎖 和所屬的鄉鎮，就住在那裏。
2CHR|28|19|因為 以色列 王 亞哈斯 在 猶大 放肆，大大干犯耶和華，所以耶和華使 猶大 卑微。
2CHR|28|20|亞述 王 提革拉‧毗列色 來攻擊他，不幫助他，反倒欺負他。
2CHR|28|21|亞哈斯 從耶和華殿裏和王宮中，以及眾領袖家中取財寶送給 亞述 王，也無濟於事。
2CHR|28|22|這 亞哈斯 王在急難的時候，越發得罪耶和華。
2CHR|28|23|他向那攻擊他的 大馬士革 的神明獻祭，說：「因為 亞蘭 王的神明幫助他們，我也要向這些神明獻祭，好讓它們幫助我。」但那些神明卻使他和全 以色列 敗亡。
2CHR|28|24|亞哈斯 聚集上帝殿裏的器皿，把上帝殿裏的器皿都打碎了，並且封鎖耶和華殿的門，又在 耶路撒冷 各處的轉角為自己建築祭壇。
2CHR|28|25|他在 猶大 各城建立丘壇，向別神燒香，惹耶和華－他列祖的上帝發怒。
2CHR|28|26|亞哈斯 其餘的事和他一切的行為，自始至終，看哪，都寫在《猶大和以色列諸王記》上。
2CHR|28|27|亞哈斯 與他祖先同睡，葬在 耶路撒冷 城裏，卻沒有送入 以色列 諸王的墳墓。他的兒子 希西家 接續他作王。
2CHR|29|1|希西家 登基的時候年二十五歲，在 耶路撒冷 作王二十九年。他母親名叫 亞比雅 ，是 撒迦利雅 的女兒。
2CHR|29|2|希西家 行耶和華眼中看為正的事，效法他祖先 大衛 一切所行的。
2CHR|29|3|元年正月，他開了耶和華殿的門，重新整修。
2CHR|29|4|他召祭司和 利未 人來，聚集在東邊的廣場，
2CHR|29|5|對他們說：「 利未 人哪，當聽我說：現在你們要將自己分別為聖，又將耶和華－你們列祖上帝的殿分別為聖，從聖所中除去污穢之物。
2CHR|29|6|因我們的祖先犯了罪，行耶和華－我們上帝眼中看為惡的事，離棄他，轉臉背向耶和華的居所。
2CHR|29|7|他們又封鎖走廊的門，吹滅燈火，不在聖所中向 以色列 的上帝燒香，或獻燔祭。
2CHR|29|8|耶和華的憤怒臨到 猶大 和 耶路撒冷 ，使他們恐懼，令人驚駭，使人嗤笑，正如你們親眼所見的。
2CHR|29|9|看哪，我們的祖宗倒在刀下，我們的妻子兒女也為此被擄掠。
2CHR|29|10|現在我心中有意與耶和華－ 以色列 的上帝立約，好使他的烈怒轉離我們。
2CHR|29|11|我的眾子啊，現在不要懈怠；因為耶和華揀選你們站在他面前事奉他，作他的僕人，向他燒香。」
2CHR|29|12|於是， 利未 人起來，當中有 哥轄 的子孫， 亞瑪賽 的兒子 瑪哈 、 亞撒利雅 的兒子 約珥 ； 米拉利 的子孫， 亞伯底 的兒子 基士 、 耶哈利勒 的兒子 亞撒利雅 ； 革順 人， 薪瑪 的兒子 約亞 、 約亞 的兒子 伊甸 ；
2CHR|29|13|以利撒反 的子孫 申利 和 耶利 ； 亞薩 的子孫， 撒迦利雅 和 瑪探雅 ；
2CHR|29|14|希幔 的子孫 耶歇 和 示每 ； 耶杜頓 的子孫 示瑪雅 和 烏薛 。
2CHR|29|15|他們聚集他們的弟兄，將自己分別為聖，照著耶和華的話和王的吩咐，進去潔淨耶和華的殿。
2CHR|29|16|祭司進入耶和華的內殿要潔淨殿，把耶和華殿中所發現一切污穢之物都搬出去，搬到耶和華殿的院子，由 利未 人接走，搬出去到外頭的 汲淪溪 。
2CHR|29|17|從正月初一開始分別為聖，初八就來到耶和華殿的走廊。他們又用了八日使耶和華的殿分別為聖，到正月十六日才完成。
2CHR|29|18|於是，他們到裏面去見 希西家 王，說：「我們已將耶和華的全殿和燔祭壇，以及壇的一切器皿、供餅的供桌，與供桌的一切器皿都潔淨了；
2CHR|29|19|並且連 亞哈斯 王在位犯罪的時候所廢棄的器皿，我們也都預備齊全，分別為聖，看哪，它們都在耶和華的祭壇前。」
2CHR|29|20|希西家 王清早起來，召集城裏的領袖都上耶和華的殿。
2CHR|29|21|他們牽了七頭公牛，七隻公羊，七隻羔羊，七隻公山羊，要為國、為殿、為 猶大 作贖罪祭。王吩咐 亞倫 的子孫眾祭司在耶和華的壇上獻祭。
2CHR|29|22|他們宰了公牛，祭司將血接來，灑在壇上；他們宰了公羊，把血灑在壇上，又宰了羔羊，也把血灑在壇上。
2CHR|29|23|他們把那些作贖罪祭的公山羊牽到王和會眾面前，按手在公山羊上。
2CHR|29|24|祭司宰了羊，將血獻在壇上作贖罪祭，為全 以色列 贖罪，因為王吩咐要為全 以色列 獻上燔祭和贖罪祭。
2CHR|29|25|王又派 利未 人在耶和華殿中敲鈸，鼓瑟，彈琴，正如 大衛 和王的先見 迦得 ，以及 拿單 先知所吩咐的，就是耶和華藉先知所吩咐的。
2CHR|29|26|利未 人拿 大衛 的樂器，祭司拿號，一同站立。
2CHR|29|27|希西家 吩咐在壇上獻燔祭，開始獻燔祭的時候，他們就唱讚美耶和華的歌，吹號，並用 以色列 王 大衛 的樂器伴奏。
2CHR|29|28|全會眾都敬拜，歌唱的歌唱，吹號的吹號，如此直到燔祭獻完了。
2CHR|29|29|獻完了祭，王和所有在場跟隨他的人都俯伏敬拜。
2CHR|29|30|希西家 王與眾領袖吩咐 利未 人用 大衛 和 亞薩 先見的詩詞頌讚耶和華，他們歡歡喜喜地頌讚，低頭敬拜。
2CHR|29|31|希西家 回應說：「如今你們既承接聖職歸耶和華，就要前來把祭物和感謝祭奉到耶和華的殿裏。」會眾就奉上祭物和感謝祭，凡甘心樂意的也奉上燔祭。
2CHR|29|32|會眾所奉的燔祭數目如下：七十頭公牛，一百隻公羊，二百隻羔羊，這些全都是要作燔祭獻給耶和華的；
2CHR|29|33|又有分別為聖之物，就是六百頭公牛，三千隻綿羊。
2CHR|29|34|但祭司太少，不能剝盡所有燔祭牲的皮，所以他們的弟兄 利未 人幫助他們，直等獻祭的事完畢，直到其他的祭司也分別為聖了；因 利未 人以正直的心分別為聖，勝過祭司。
2CHR|29|35|燔祭和平安祭牲的脂肪，以及與燔祭同獻的澆酒祭很多。這樣，耶和華殿中的事務俱都齊備了。
2CHR|29|36|希西家 和眾百姓都因上帝為百姓所預備的而喜樂，因為這事辦得很迅速。
2CHR|30|1|希西家 派人去見 以色列 和 猶大 眾人，又寫信給 以法蓮 和 瑪拿西 人，要他們到 耶路撒冷 耶和華的殿，向耶和華－ 以色列 的上帝守逾越節，
2CHR|30|2|因為王和眾領袖，以及 耶路撒冷 全會眾已經商議，要在二月份守逾越節。
2CHR|30|3|那時他們不能守，因為分別為聖的祭司不夠，百姓也還沒有聚集在 耶路撒冷 。
2CHR|30|4|這事在王與全會眾眼中都看為合宜。
2CHR|30|5|於是他們下令，通告全 以色列 ，從 別是巴 直到 但 ，吩咐百姓都來，在 耶路撒冷 向耶和華－ 以色列 的上帝守逾越節，因為他們已經許久沒有照所寫的守這節了 。
2CHR|30|6|信差遵著王命，拿著王和眾領袖所發的信，送達全 以色列 和 猶大 ，說：「 以色列 人哪，當轉向耶和華－ 亞伯拉罕 、 以撒 、 以色列 的上帝，好叫他轉向你們這些脫離 亞述 諸王之手的餘民。
2CHR|30|7|不要效法你們的祖先和你們的弟兄；他們干犯耶和華－他們列祖的上帝，以致耶和華使他們令人驚駭，正如你們所見的。
2CHR|30|8|現在，不要像你們祖先硬著頸項，只要歸順耶和華，進入他的聖所，就是永遠成聖的居所，又要事奉耶和華－你們的上帝，好使他的烈怒轉離你們。
2CHR|30|9|你們若轉向耶和華，你們的弟兄和兒女必在擄掠他們的人面前蒙憐憫，得以歸回這地，因為耶和華－你們的上帝有恩惠，有憐憫。你們若轉向他，他必不會轉臉不顧你們。」
2CHR|30|10|信差從這城跑到那城，傳遍了 以法蓮 和 瑪拿西 之地，直到 西布倫 ；那裏的人卻戲笑他們，譏誚他們。
2CHR|30|11|然而 亞設 、 瑪拿西 、 西布倫 中也有人謙卑自己，來到 耶路撒冷 。
2CHR|30|12|上帝也按手在 猶大 人身上，使他們一心遵行王與眾領袖照著耶和華的話所發的命令。
2CHR|30|13|二月時，許多百姓聚集在 耶路撒冷 ，成為一個盛大的會，要守除酵節。
2CHR|30|14|他們起來，把 耶路撒冷 的祭壇和燒香的壇盡都除去，扔在 汲淪溪 中。
2CHR|30|15|二月十四日，他們宰了逾越節的羔羊。祭司與 利未 人覺得慚愧，就使自己分別為聖，把燔祭奉到耶和華的殿中。
2CHR|30|16|他們遵照神人 摩西 的律法，按定例站在自己的地方；祭司從 利未 人手裏接過血來，灑出去。
2CHR|30|17|會眾中有許多人尚未分別為聖，所以 利未 人為所有不潔的人宰逾越節的羔羊，使他們歸耶和華為聖。
2CHR|30|18|從 以法蓮 、 瑪拿西 、 以薩迦 、 西布倫 來的許多百姓尚未自潔，他們卻吃逾越節的羔羊，不合所寫的條例。 希西家 為他們禱告說：「求至善的耶和華饒恕
2CHR|30|19|那凡專心尋求上帝耶和華－他列祖的上帝，卻未照聖所潔淨禮自潔的人。」
2CHR|30|20|耶和華應允 希西家 ，醫治了百姓。
2CHR|30|21|在 耶路撒冷 的 以色列 人守除酵節七日，大大喜樂。 利未 人和祭司為耶和華演奏響亮的樂器，天天頌讚耶和華。
2CHR|30|22|希西家 慰勞所有精通禮儀，事奉耶和華的 利未 人。於是眾人吃節期的筵席七日，又獻平安祭，並且稱謝耶和華－他們列祖的上帝。
2CHR|30|23|全會眾商議，要再守節七日；於是他們歡歡喜喜地又守節七日。
2CHR|30|24|猶大 王 希西家 賜給會眾一千頭公牛，七千隻羊；眾領袖也賜給會眾一千頭公牛，一萬隻羊，並有許多祭司將自己分別為聖。
2CHR|30|25|猶大 全會眾、祭司、 利未 人和從 以色列 來的全會眾，以及那些從 以色列 地來的和住在 猶大 的寄居的人，盡都喜樂。
2CHR|30|26|這樣，在 耶路撒冷 大有喜樂，因自從 以色列 王 大衛 的兒子 所羅門 以來，在 耶路撒冷 從未有過這樣的喜樂。
2CHR|30|27|那時，祭司和 利未 人起來，為百姓祝福。他們的聲音蒙上帝垂聽，他們的禱告達到他天上的聖所。
2CHR|31|1|這一切事都完畢以後，在那裏的 以色列 眾人就到 猶大 的城鎮，打碎柱像，砍斷 亞舍拉 ，又在 猶大 、 便雅憫 、 以法蓮 、 瑪拿西 遍地把丘壇和祭壇完全拆毀。於是 以色列 眾人各回各城，各歸自己產業的地去了。
2CHR|31|2|希西家 分派祭司和 利未 人的班次，使祭司和 利未 人照各自的班次，按各自的職分獻燔祭和平安祭，又在耶和華殿 的門內事奉，稱謝頌讚耶和華。
2CHR|31|3|王又從自己的產業中分出一份來作燔祭，就是早晚的燔祭，和安息日、初一，以及節期的燔祭，都是按耶和華律法上所記載的。
2CHR|31|4|他又吩咐住 耶路撒冷 的百姓將祭司和 利未 人所應得的份給他們，使他們堅守耶和華的律法。
2CHR|31|5|命令一出， 以色列 人就把初熟的五穀、新酒、新油、蜜和田地的出產多多送來；他們把各樣出產的十分之一大量送來。
2CHR|31|6|住 猶大 各城的 以色列 人和 猶大 人也將牛羊的十分之一，以及分別為聖歸耶和華－他們上帝之物，就是十分取一之物，盡都送來，積成一堆一堆；
2CHR|31|7|他們從三月開始堆積，到七月才完成。
2CHR|31|8|希西家 和眾領袖來，看見這些堆積物，就稱頌耶和華，又為耶和華的百姓 以色列 祝福。
2CHR|31|9|希西家 向祭司和 利未 人查問這些堆積物。
2CHR|31|10|撒督 家的 亞撒利雅 祭司長告訴他說：「自從禮物開始送到耶和華的殿以來，我們不但吃飽，而且剩下的很多；因為耶和華賜福給他的百姓，所剩下的才這樣豐盛。」
2CHR|31|11|希西家 吩咐要在耶和華殿裏預備倉房，他們就預備了。
2CHR|31|12|他們誠心將禮物，十分取一之物，就是分別為聖之物，都搬入倉內。 利未 人 歌楠雅 主管這事，他的兄弟 示每 是副主管。
2CHR|31|13|耶歇 、 亞撒細雅 、 拿哈 、 亞撒黑 、 耶利摩 、 約撒拔 、 以列 、 伊斯瑪基雅 、 瑪哈 、 比拿雅 都是督辦，在 歌楠雅 和他兄弟 示每 的手下，是 希西家 王和管理上帝殿的 亞撒利雅 所委派的。
2CHR|31|14|守東門的 利未 人 音拿 的兒子 可利 ，掌管獻給上帝的甘心祭，發放獻給耶和華的禮物和至聖的物。
2CHR|31|15|在祭司的各城裏，在他手下忠心協助他的有 伊甸 、 (王民)雅(王民) 、 耶書亞 、 示瑪雅 、 亞瑪利雅 、 示迦尼雅 ，都按著班次分給他們的弟兄，無論大小，
2CHR|31|16|不論是否登錄在家譜，凡三歲以上的男丁，每日進耶和華殿、按班次供職事奉的，都分給他，
2CHR|31|17|也發放給按父家登錄在家譜的祭司；又按班次職任分給二十歲以上的 利未 人，
2CHR|31|18|又按家譜的登記，分給他們的小孩、妻子、兒女，給全體會眾；因為他們忠誠，將自己分別為聖。
2CHR|31|19|住在各城郊野 亞倫 的子孫、按名受委任的人，要把應得的份給祭司中所有的男丁和載入家譜的 利未 人。
2CHR|31|20|希西家 在全 猶大 都這樣辦理，在耶和華－他上帝面前行良善、正直、忠誠的事。
2CHR|31|21|凡他所行的，無論是開始辦上帝殿的事，是遵律法守誡命，是尋求他的上帝，他都盡心去做，無不亨通。
2CHR|32|1|在這些虔誠的事以後， 亞述 王 西拿基立 來侵犯 猶大 ，圍困堅固城，想要攻破它們。
2CHR|32|2|希西家 見 西拿基立 來，定意要攻打 耶路撒冷 ，
2CHR|32|3|就與領袖和勇士商議，塞住城外的泉源；他們都幫助他。
2CHR|32|4|於是許多百姓聚集，塞住一切泉源，以及國中流通的小河，說：「 亞述 諸王來，為何讓他們得著許多水呢？」
2CHR|32|5|希西家 奮勇自強，修築所有毀壞的城牆，升高城樓，又在城外築另一片城牆，堅固 大衛城 的 米羅 ，製造許多兵器和盾牌。
2CHR|32|6|他設立軍事將領管理百姓，召集他們在城門的廣場，勉勵他們，說：
2CHR|32|7|「你們當剛強壯膽，不要因 亞述 王和跟隨他的大軍恐懼驚慌，因為與我們同在的，比與他們同在的更大。
2CHR|32|8|與他們同在的是血肉之臂，但與我們同在的是耶和華－我們的上帝，他必幫助我們，為我們爭戰。」百姓因 猶大 王 希西家 的話就得到鼓勵。
2CHR|32|9|此後， 亞述 王 西拿基立 和跟隨他的全軍攻打 拉吉 ，派臣僕到 耶路撒冷 見 猶大 王 希西家 和所有在 耶路撒冷 的 猶大 人，說：
2CHR|32|10|「 亞述 王 西拿基立 如此說：『你們倚靠甚麼，還留在 耶路撒冷 受困嗎？
2CHR|32|11|希西家 說：耶和華－我們的上帝必救我們脫離 亞述 王的手，這不是誘惑你們，使你們受飢渴而死嗎？
2CHR|32|12|希西家 豈不是將耶和華的丘壇和祭壇廢去，並且吩咐 猶大 與 耶路撒冷 的人說：你們當在一個壇前敬拜，在其上燒香嗎？
2CHR|32|13|我與我祖先向列邦民族所行的，你們豈不知道嗎？列邦的神明何嘗能救自己的國脫離我的手呢？
2CHR|32|14|我祖先所滅的那些國的神明，有誰能救自己的百姓脫離我的手呢？難道你們的上帝能救你們脫離我的手嗎？
2CHR|32|15|現在，不要讓 希西家 這樣欺騙你們，誘惑你們，也不要相信他，因為沒有一國一邦的神明能救自己的百姓脫離我的手和我祖先的手，你們的上帝也絕不能救你們脫離我的手。』」
2CHR|32|16|西拿基立 的臣僕還說了一些話來毀謗耶和華上帝和他的僕人 希西家 。
2CHR|32|17|西拿基立 也寫信毀謗耶和華－ 以色列 的上帝，說：「列邦的神明既不能救自己的百姓脫離我的手， 希西家 的上帝也不能救他的百姓脫離我的手。」
2CHR|32|18|亞述 王的臣僕用 猶大 話向 耶路撒冷 城牆上的百姓大聲呼喊，要恐嚇他們，擾亂他們，以便取城。
2CHR|32|19|他們談論 耶路撒冷 的上帝，如同談論世上人手所造的神明一樣。
2CHR|32|20|希西家 王和 亞摩斯 的兒子 以賽亞 先知為此禱告，向天呼求。
2CHR|32|21|耶和華就差遣一個使者進入 亞述 王的營中，把所有大能的勇士、官長和將領盡都滅了。 亞述 王滿面羞愧地回到本國，進了他神明的廟中，他幾個親生的兒子在那裏用刀殺了他。
2CHR|32|22|這樣，耶和華救 希西家 和 耶路撒冷 的居民脫離 亞述 王 西拿基立 的手，也脫離一切仇敵的手，又賜他們四境平安 。
2CHR|32|23|有許多人到 耶路撒冷 將供物獻與耶和華，又將寶物送給 猶大 王 希西家 。自此之後， 希西家 在列國人的眼中受人尊崇。
2CHR|32|24|那些日子， 希西家 病得要死，就向耶和華禱告，耶和華應允他，賜他一個預兆。
2CHR|32|25|希西家 卻沒有照他所蒙的恩回報，因他心裏驕傲，所以憤怒要臨到他，臨到 猶大 和 耶路撒冷 。
2CHR|32|26|但 希西家 和 耶路撒冷 的居民為了心裏驕傲，就一同謙卑，以致耶和華的憤怒在 希西家 的日子沒有臨到他們。
2CHR|32|27|希西家 大有財富和尊榮，他為自己建造府庫，收藏金銀、寶石、香料、盾牌和各樣的寶器，
2CHR|32|28|又建造倉房，收藏五穀、新酒和新的油，又為各類牲畜蓋棚立圈，
2CHR|32|29|並且為自己建立城鎮，也擁有許多的羊群牛群，因為上帝賜他極多的財產。
2CHR|32|30|這 希西家 也塞住 基訓 的上源，引水直下，流在 大衛城 的西邊。 希西家 所行的事盡都亨通。
2CHR|32|31|但當 巴比倫 諸侯差遣使者來見 希西家 ，詢問國中所發生的奇事時，上帝離開他，要考驗他，好知道他心裏的一切。
2CHR|32|32|希西家 其餘的事和他的善行，看哪，都寫在 亞摩斯 的兒子 以賽亞 先知的《默示書》上和《猶大和以色列諸王記》上。
2CHR|32|33|希西家 與他祖先同睡，葬在 大衛 子孫陵墓的斜坡上。他死的時候， 猶大 眾人和 耶路撒冷 的居民都向他致敬。他的兒子 瑪拿西 接續他作王。
2CHR|33|1|瑪拿西 登基的時候年十二歲，在 耶路撒冷 作王五十五年。
2CHR|33|2|他行耶和華眼中看為惡的事，效法耶和華在 以色列 人面前趕出的列國那些可憎的事。
2CHR|33|3|他重新建築他父親 希西家 所拆毀的丘壇，為諸 巴力 築壇，造 亞舍拉 ，又敬拜天上的萬象，事奉它們。
2CHR|33|4|他在耶和華殿中築壇，耶和華曾指著這殿說：「我的名必永遠在 耶路撒冷 。」
2CHR|33|5|他在耶和華殿的兩個院子為天上的萬象築壇，
2CHR|33|6|並在 欣嫩子谷 使他的兒子經火，又觀星象，行法術，行邪術，求問招魂的和行巫術的，多行耶和華眼中看為惡的事，惹他發怒。
2CHR|33|7|他在上帝殿內立雕刻的偶像；上帝曾對 大衛 和他兒子 所羅門 說：「我在 以色列 眾支派中所選擇的 耶路撒冷 和這殿，必立我的名，直到永遠。
2CHR|33|8|只要 以色列 人謹守遵行我藉 摩西 吩咐他們的一切律法、律例、典章，我就不再使他們的腳挪移，離開我所賜給他們列祖之土地。」
2CHR|33|9|瑪拿西 引誘 猶大 和 耶路撒冷 的居民行惡，比耶和華在 以色列 人面前所滅的列國更嚴重。
2CHR|33|10|耶和華警戒 瑪拿西 和他的百姓，他們卻不聽。
2CHR|33|11|所以耶和華使 亞述 王的將領來攻擊他們，用手銬銬住 瑪拿西 ，用銅鏈鎖住他，把他帶到 巴比倫 去。
2CHR|33|12|他在急難的時候懇求耶和華－他的上帝，並在他列祖的上帝面前極其謙卑。
2CHR|33|13|他祈禱耶和華，耶和華就應允他，垂聽他的禱告，使他歸回 耶路撒冷 ，仍坐王位。 瑪拿西 這才知道惟獨耶和華是上帝。
2CHR|33|14|此後， 瑪拿西 在 大衛城 外，從谷內 基訓 西邊直到 魚門 口，建築城牆，環繞 俄斐勒 ；這牆建得很高。他又在 猶大 各堅固城內設立將領。
2CHR|33|15|他除掉外邦人的神像與耶和華殿中的偶像，又將他在耶和華殿的山上和 耶路撒冷 所築的各壇都拆毀，拋在城外。
2CHR|33|16|他重修耶和華的祭壇，在壇上獻平安祭和感謝祭，並吩咐 猶大 人事奉耶和華－ 以色列 的上帝。
2CHR|33|17|百姓卻仍在丘壇上獻祭，不過，他們只獻給耶和華－他們的上帝。
2CHR|33|18|瑪拿西 其餘的事和他向上帝的禱告，以及先見奉耶和華－ 以色列 上帝的名警戒他的話，看哪，都在《以色列諸王記》上。
2CHR|33|19|他的禱告，上帝怎樣應允他，他未謙卑以前的一切罪愆過犯，以及在何處建築丘壇，設立 亞舍拉 和雕刻的偶像，看哪，都寫在 何賽 的書上。
2CHR|33|20|瑪拿西 與他祖先同睡，葬在自己的宮中，他兒子 亞們 接續他作王。
2CHR|33|21|亞們 登基的時候年二十二歲，在 耶路撒冷 作王二年。
2CHR|33|22|他行耶和華眼中看為惡的事，效法他父親 瑪拿西 所行的，祭祀他父親 瑪拿西 所雕刻的一切偶像，事奉它們，
2CHR|33|23|但他不像他父親 瑪拿西 在耶和華面前那樣謙卑下來。這 亞們 的罪越犯越大。
2CHR|33|24|他的臣僕背叛他，在宮裏殺了他。
2CHR|33|25|但這地的百姓殺了所有背叛 亞們 王的人；這地的百姓立他兒子 約西亞 接續他作王。
2CHR|34|1|約西亞 登基的時候年八歲，在 耶路撒冷 作王三十一年。
2CHR|34|2|他行耶和華眼中看為正的事，行他祖先 大衛 所行的道，不偏左右。
2CHR|34|3|他作王第八年，尚且年輕，就尋求他祖先 大衛 的上帝。到了十二年，他開始潔淨 猶大 和 耶路撒冷 ，除掉丘壇、 亞舍拉 、雕刻的像和鑄造的像。
2CHR|34|4|眾人在他面前拆毀諸 巴力 的壇，砍斷壇上高高的香壇，又把 亞舍拉 和雕刻的像，以及鑄造的像打碎成灰，撒在向偶像獻祭之人的墳上，
2CHR|34|5|把祭司的骸骨燒在他們的壇上，潔淨了 猶大 和 耶路撒冷 。
2CHR|34|6|他又在 瑪拿西 、 以法蓮 、 西緬 、 拿弗他利 各城和四圍的廢墟 ，
2CHR|34|7|拆毀祭壇，把 亞舍拉 和雕刻的像打碎成灰，砍斷 以色列 全地所有的香壇。於是他回 耶路撒冷 去了。
2CHR|34|8|約西亞 王十八年，這地和殿潔淨了之後，他派 亞薩利雅 的兒子 沙番 、 瑪西雅 市長、 約哈斯 的兒子 約亞 史官去整修耶和華－他上帝的殿。
2CHR|34|9|他們去見 希勒家 大祭司，把奉到上帝殿的銀子交給他；這銀子是看守殿門的 利未 人從 瑪拿西 、 以法蓮 ，和 以色列 所有倖存的人，以及 猶大 、 便雅憫 眾人和 耶路撒冷 的居民收來的。
2CHR|34|10|他們把這銀子交給耶和華殿裏督工的，由他們轉交整修耶和華殿的工匠，
2CHR|34|11|就是交給木匠和石匠，好為 猶大 王所毀壞的殿，買鑿成的石頭和作鉤子與棟梁的木料。
2CHR|34|12|這些人辦事誠實，管理他們的是 利未 人 米拉利 的子孫 雅哈 和 俄巴底 ，又有 哥轄 人 撒迦利亞 和 米書蘭 ；還有所有善於奏樂的 利未 人。
2CHR|34|13|他們監督扛抬的人，督導一切做各樣工的人。 利未 人中也有作書記、官員、守衛的。
2CHR|34|14|他們把奉到耶和華殿的銀子運出來的時候， 希勒家 祭司發現了耶和華藉 摩西 所傳的律法書。
2CHR|34|15|希勒家 對 沙番 書記說：「我在耶和華殿裏發現了律法書。」 希勒家 把書遞給 沙番 。
2CHR|34|16|沙番 把書拿到王那裏，又把這事回覆王說：「凡交給僕人的手所辦的事，他們都辦好了。
2CHR|34|17|耶和華殿裏所發現的銀子已經倒出來，交在督工和工匠的手裏了。」
2CHR|34|18|沙番 書記又向王報告說：「 希勒家 祭司遞給我一卷書。」 沙番 就在王面前朗讀那書。
2CHR|34|19|王聽見律法的話，就撕裂衣服。
2CHR|34|20|王吩咐 希勒家 與 沙番 的兒子 亞希甘 、 米迦 的兒子 亞比頓 、 沙番 書記和王的臣僕 亞撒雅 ，說：
2CHR|34|21|「你們去，以所發現這書上的話，為我、為 以色列 和 猶大 倖存的人求問耶和華；因為我們的祖先沒有遵守耶和華的話，沒有照這書上所記的一切去做，耶和華的烈怒就倒在我們身上。」
2CHR|34|22|於是， 希勒家 和王的人 都去見 戶勒大 女先知，她是掌管禮服的 沙龍 的妻子， 沙龍 是 哈斯拉 的孫子， 特瓦 的兒子。 戶勒大 住在 耶路撒冷 第二區。他們向她說明來意。
2CHR|34|23|她對他們說：「耶和華－ 以色列 的上帝如此說：『你們可以回覆那派你們來見我的人說，
2CHR|34|24|耶和華如此說：看哪，我必照著在 猶大 王面前所讀那書上記載的一切詛咒，降禍於這地方和其上的居民。
2CHR|34|25|因為他們離棄我，向別神燒香，用他們手所做的一切惹我發怒，所以我的憤怒必倒在這地方，總不止息。』
2CHR|34|26|然而，派你們來求問耶和華的 猶大 王，你們要這樣回覆他：『耶和華－ 以色列 的上帝如此說：至於你所聽見的話，
2CHR|34|27|就是聽見我指著這地方和其上居民所說的話，你的心就軟化，在我面前謙卑下來，撕裂衣服，向我哭泣，因此我應允你。這是耶和華說的。
2CHR|34|28|看哪，我必使你歸到你祖先那裏，平安地進入墳墓，我要降於這地方和其上居民的一切災禍，你不會親眼看見。』」他們就去把這話回覆王。
2CHR|34|29|王派人召集 猶大 和 耶路撒冷 的眾長老來。
2CHR|34|30|王和 猶大 眾人、 耶路撒冷 的居民、祭司、 利未 人，以及所有的百姓，無論大小，都一同上到耶和華的殿去；王把殿裏所發現的約書上面一切的話讀給他們聽。
2CHR|34|31|王站在自己的位上，在耶和華面前立約，要盡心盡性跟從耶和華，遵守他的誡命、法度、律例，實行這書上所記這約的話；
2CHR|34|32|又使所有住 耶路撒冷 和 便雅憫 的人都服從這約。於是 耶路撒冷 的居民都遵行上帝，就是他們列祖之上帝的約。
2CHR|34|33|約西亞 從 以色列 各處把一切可憎之物盡都除掉，使 以色列 境內的人都事奉耶和華－他們的上帝。 約西亞 在世的日子，眾人都跟從耶和華－他們列祖的上帝，總不離開。
2CHR|35|1|約西亞 在 耶路撒冷 向耶和華守逾越節。正月十四日，他們宰了逾越節的羔羊。
2CHR|35|2|王分派祭司各盡其職，又勉勵他們辦耶和華殿中的事。
2CHR|35|3|他對那歸耶和華為聖、教導 以色列 眾人的 利未 人說：「你們將聖約櫃安放在 以色列 王 大衛 兒子 所羅門 建造的殿裏，不必再用肩扛抬。現在你們要服事耶和華－你們的上帝和他的百姓 以色列 。
2CHR|35|4|你們應當按著父家，照著班次，遵照 以色列 王 大衛 和他兒子 所羅門 所寫的，預備自己。
2CHR|35|5|要按著你們百姓的弟兄、父家的班次，侍立在聖所；每父家的班次中要有幾個 利未 人。
2CHR|35|6|要宰逾越節的羔羊，將自己分別為聖，為你們的弟兄預備，好遵守耶和華藉 摩西 所吩咐的話。」
2CHR|35|7|約西亞 從群畜中賜給所有在場的百姓，三萬隻小綿羊和小山羊，三千頭牛，作逾越節的祭物；這些都是出自王的產業。
2CHR|35|8|約西亞 的眾領袖也樂意把祭牲給百姓、祭司和 利未 人；管理上帝殿的 希勒家 、 撒迦利亞 、 耶歇 ，把二千六百隻羔羊和三百頭牛給祭司作逾越節的祭物。
2CHR|35|9|利未 人的族長 歌楠雅 和他兩個兄弟 示瑪雅 、 拿坦業 ，與 哈沙比雅 、 耶利 、 約撒拔 ，把五千隻羔羊和五百頭牛給 利未 人作逾越節的祭物。
2CHR|35|10|這樣，事奉的工作都安排好了，照王所吩咐的，祭司站在自己的位上， 利未 人按著班次侍立。
2CHR|35|11|他們宰了逾越節的羔羊，祭司從他們手裏接過血來 灑出去； 利未 人剝皮，
2CHR|35|12|把燔祭拿走，再按著父家的班次分給眾百姓，照 摩西 書上所寫的獻給耶和華；獻牛也是這樣。
2CHR|35|13|他們按著常例，用火烤逾越節的羔羊。至於其他的聖物，他們用盆，用鍋，用釜煮了，速速地送給眾百姓。
2CHR|35|14|然後他們為自己和祭司預備祭物，因為作祭司的 亞倫 子孫獻燔祭和脂肪，直到晚上。所以 利未 人為自己和作祭司的 亞倫 子孫預備。
2CHR|35|15|歌唱的 亞薩 子孫，照著 大衛 、 亞薩 、 希幔 和王的先見 耶杜頓 所吩咐的，站在自己的位上。守門的看守各門，不用離開他們的職守，因為他們的弟兄 利未 人給他們預備。
2CHR|35|16|當日，一切供奉耶和華、守逾越節，以及在耶和華壇上獻燔祭的事，都照 約西亞 王的吩咐預備好了。
2CHR|35|17|那時，在場的 以色列 人都守逾越節，又守除酵節七日。
2CHR|35|18|自從 撒母耳 先知的日子以來，在 以色列 中沒有守過這樣的逾越節， 以色列 諸王也沒有守過像 約西亞 、祭司、 利未 人、所有住 猶大 和 以色列 的人，以及 耶路撒冷 居民所守的逾越節。
2CHR|35|19|這逾越節是 約西亞 作王十八年時守的。
2CHR|35|20|約西亞 為殿做完這一切事以後， 埃及 王 尼哥 上來，要攻打靠近 幼發拉底河 的 迦基米施 ； 約西亞 出去迎擊他。
2CHR|35|21|他派使者來見 約西亞 ，說：「 猶大 王啊，我跟你有甚麼相干呢？我今日來不是要攻打你，而是要攻打與我爭戰之家，並且上帝吩咐我從速行事。你不要干預與我同在的上帝，免得他毀滅你。」
2CHR|35|22|約西亞 卻不轉臉離開他，反而改裝要與他打仗。他不聽從上帝藉 尼哥 的口所說的話，就來到 米吉多 平原爭戰。
2CHR|35|23|弓箭手射中 約西亞 王。王對他的臣僕說：「我受了重傷，你們載我離開戰場吧！」
2CHR|35|24|他的臣僕扶他下了戰車，上了他的副座車，送他到 耶路撒冷 。他就死了，葬在他祖先的墳墓裏。全 猶大 和 耶路撒冷 都哀悼 約西亞 。
2CHR|35|25|耶利米 為 約西亞 作哀歌，所有歌唱的男女也唱哀歌，追悼 約西亞 ，直到今日。他們在 以色列 中以此為定例；看哪，這些哀歌寫在《哀歌書》上。
2CHR|35|26|約西亞 其餘的事和他遵照耶和華律法上所記而行的善事，
2CHR|35|27|以及他自始至終所行的，看哪，都寫在《以色列和猶大列王記》上。
2CHR|36|1|這地的百姓立 約西亞 的兒子 約哈斯 在 耶路撒冷 接續他父親作王。
2CHR|36|2|約哈斯 登基的時候年二十三歲，在 耶路撒冷 作王三個月。
2CHR|36|3|埃及 王在 耶路撒冷 廢了他，又罰這地一百他連得銀子，一他連得金子。
2CHR|36|4|埃及 王 尼哥 立 約哈斯 的哥哥 以利雅敬 作 猶大 和 耶路撒冷 的王，給他改名叫 約雅敬 。 尼哥 卻將他的弟弟 約哈斯 帶到 埃及 去。
2CHR|36|5|約雅敬 登基的時候年二十五歲，在 耶路撒冷 作王十一年。他行耶和華－他上帝眼中看為惡的事。
2CHR|36|6|巴比倫 王 尼布甲尼撒 上來攻擊他，用銅鏈鎖著他，要把他帶到 巴比倫 去。
2CHR|36|7|尼布甲尼撒 又將耶和華殿裏的一些器皿帶到 巴比倫 ，放在 巴比倫 自己的宮裏 。
2CHR|36|8|約雅敬 其餘的事和他所行可憎的事，以及發生在他身上的事，看哪，都寫在《以色列和猶大列王記》上，他兒子 約雅斤 接續他作王。
2CHR|36|9|約雅斤 登基的時候年八歲 ，在 耶路撒冷 作王三個月十天，他行耶和華眼中看為惡的事。
2CHR|36|10|過了一年， 尼布甲尼撒 王差遣人將 約雅斤 和耶和華殿裏寶貴的器皿帶到 巴比倫 ，然後立 約雅斤 的叔父 西底家 作 猶大 和 耶路撒冷 的王。
2CHR|36|11|西底家 登基的時候年二十一歲，在 耶路撒冷 作王十一年。
2CHR|36|12|他行耶和華－他上帝眼中看為惡的事，沒有謙卑聽從 耶利米 先知所傳達耶和華的話。
2CHR|36|13|尼布甲尼撒 王曾叫他指著上帝起誓，他卻背叛，硬著頸項，內心頑固，不歸向耶和華－ 以色列 的上帝。
2CHR|36|14|眾祭司長和百姓也多多犯罪，效法列國一切可憎的事，玷污耶和華在 耶路撒冷 分別為聖的殿。
2CHR|36|15|耶和華－他們列祖的上帝因為愛惜自己的百姓和居所，一再差遣使者去警戒他們。
2CHR|36|16|他們卻嘲笑上帝的使者，藐視他的話，譏誚他的先知，以致耶和華向他的百姓大發烈怒，甚至無法可救。
2CHR|36|17|所以，耶和華使 迦勒底 人的王來攻擊他們，在他們聖殿裏用刀殺了他們的壯丁，不憐憫他們的少男少女、老人長者。耶和華把所有的人都交在他手裏。
2CHR|36|18|他把上帝殿裏一切的大小器皿與耶和華殿裏的財寶，以及王和眾領袖的財寶，全都帶到 巴比倫 去。
2CHR|36|19|迦勒底 人焚燒了上帝的殿，拆毀 耶路撒冷 的城牆，用火燒了城裏所有的宮殿，毀壞了城裏一切寶貴的器皿。
2CHR|36|20|凡脫離刀劍的倖存者， 迦勒底 王都擄到 巴比倫 去，作他和他子孫的僕婢，直到 波斯 國興起。
2CHR|36|21|這就應驗耶和華藉 耶利米 的口所說的話：地得享安息；在荒涼的日子，地就守安息，直到滿了七十年。
2CHR|36|22|波斯 王 居魯士 元年，耶和華為要應驗藉 耶利米 的口所說的話，就激發 波斯 王 居魯士 的心，使他下詔書通告全國，說：
2CHR|36|23|「 波斯 王 居魯士 如此說：耶和華－天上的上帝已將地上萬國賜給我，又委派我在 猶大 的 耶路撒冷 為他建造殿宇。你們中間凡作他子民的可以上去，願耶和華－他的上帝與他同在。」
EZRA|1|1|波斯 王 居魯士 元年，耶和華為要應驗藉 耶利米 的口所說的話，就激發 波斯 王 居魯士 的心，使他下詔書通告全國，說：
EZRA|1|2|「 波斯 王 居魯士 如此說：耶和華天上的上帝已將地上萬國賜給我，又委派我在 猶大 的 耶路撒冷 為他建造殿宇。
EZRA|1|3|你們中間凡作他子民的，可以上 猶大 的 耶路撒冷 去，重建耶和華－ 以色列 上帝的殿，他是在 耶路撒冷 的上帝；願上帝與這人同在。
EZRA|1|4|凡存留的人，無論寄居何處，那地的人要用金銀、財物、牲畜幫助他，還要為 耶路撒冷 上帝的殿甘心獻上禮物。」
EZRA|1|5|於是， 猶大 和 便雅憫 的族長、祭司、 利未 人，凡是心被上帝感動的人都起來，要上 耶路撒冷 去建造耶和華的殿。
EZRA|1|6|四圍所有的人都拿銀器 、金子、財物、牲畜、珍寶支持他們 ，此外還有甘心獻的一切禮物 。
EZRA|1|7|居魯士 王也把耶和華殿的器皿拿出來，這些器皿是 尼布甲尼撒 從 耶路撒冷 掠取，放在自己神明廟中的。
EZRA|1|8|波斯 王 居魯士 派 米提利達 司庫把這些器皿拿出來，點交給 猶大 的領袖 設巴薩 。
EZRA|1|9|它們的數目如下：金盤三十個，銀盤一千個，刀二十九把，
EZRA|1|10|金碗三十個，備用銀碗四百一十個，其他器皿一千件。
EZRA|1|11|金銀器皿共有五千四百件。被擄的人從 巴比倫 上 耶路撒冷 的時候， 設巴薩 把這一切都帶了上來。
EZRA|2|1|這些是從被擄之地上來的省民， 巴比倫 王 尼布甲尼撒 把他們擄到 巴比倫 ，他們重返 耶路撒冷 和 猶大 ，各歸本城。
EZRA|2|2|他們是同 所羅巴伯 、 耶書亞 、 尼希米 、 西萊雅 、 利來雅 、 末底改 、 必珊 、 米斯拔 、 比革瓦伊 、 利宏 、 巴拿 一起回來的。 以色列 百姓的人數如下：
EZRA|2|3|巴錄 的子孫二千一百七十二名；
EZRA|2|4|示法提雅 的子孫三百七十二名；
EZRA|2|5|亞拉 的子孫七百七十五名；
EZRA|2|6|巴哈‧摩押 的後裔，就是 耶書亞 和 約押 的子孫二千八百一十二名；
EZRA|2|7|以攔 的子孫一千二百五十四名；
EZRA|2|8|薩土 的子孫九百四十五名；
EZRA|2|9|薩改 的子孫七百六十名；
EZRA|2|10|巴尼 的子孫六百四十二名；
EZRA|2|11|比拜 的子孫六百二十三名；
EZRA|2|12|押甲 的子孫一千二百二十二名；
EZRA|2|13|亞多尼干 的子孫六百六十六名；
EZRA|2|14|比革瓦伊 的子孫二千零五十六名；
EZRA|2|15|亞丁 的子孫四百五十四名；
EZRA|2|16|亞特 的後裔，就是 希西家 的子孫九十八名；
EZRA|2|17|比賽 的子孫三百二十三名；
EZRA|2|18|約拉 的子孫一百一十二名；
EZRA|2|19|哈順 的子孫二百二十三名；
EZRA|2|20|吉罷珥 人九十五名；
EZRA|2|21|伯利恆 人一百二十三名；
EZRA|2|22|尼陀法 人五十六名；
EZRA|2|23|亞拿突 人一百二十八名；
EZRA|2|24|亞斯瑪弗 人四十二名；
EZRA|2|25|基列‧耶琳 人、 基非拉 人、 比錄 人共七百四十三名；
EZRA|2|26|拉瑪 人和 迦巴 人共六百二十一名；
EZRA|2|27|默瑪 人一百二十二名；
EZRA|2|28|伯特利 人和 艾 人共二百二十三名；
EZRA|2|29|尼波 人五十二名；
EZRA|2|30|末必 人一百五十六名；
EZRA|2|31|另一個 以攔 的子孫一千二百五十四名；
EZRA|2|32|哈琳 的子孫三百二十名；
EZRA|2|33|羅德 人、 哈第 人、 阿挪 人共七百二十五名；
EZRA|2|34|耶利哥 人三百四十五名；
EZRA|2|35|西拿 人三千六百三十名。
EZRA|2|36|祭司： 耶書亞 家 耶大雅 的子孫九百七十三名；
EZRA|2|37|音麥 的子孫一千零五十二名；
EZRA|2|38|巴施戶珥 的子孫一千二百四十七名；
EZRA|2|39|哈琳 的子孫一千零一十七名。
EZRA|2|40|利未 人： 何達威雅 的後裔，就是 耶書亞 和 甲篾 的子孫七十四名。
EZRA|2|41|歌唱的： 亞薩 的子孫一百二十八名。
EZRA|2|42|門口的守衛： 沙龍 的子孫、 亞特 的子孫、 達們 的子孫、 亞谷 的子孫、 哈底大 的子孫、 朔拜 的子孫，共一百三十九名。
EZRA|2|43|殿役： 西哈 的子孫、 哈蘇巴 的子孫、 答巴俄 的子孫、
EZRA|2|44|基綠 的子孫、 西亞 的子孫、 巴頓 的子孫、
EZRA|2|45|利巴拿 的子孫、 哈迦巴 的子孫、 亞谷 的子孫、
EZRA|2|46|哈甲 的子孫、 薩買 的子孫、 哈難 的子孫、
EZRA|2|47|吉德 的子孫、 迦哈 的子孫、 利亞雅 的子孫、
EZRA|2|48|利汛 的子孫、 尼哥大 的子孫、 迦散 的子孫、
EZRA|2|49|烏撒 的子孫、 巴西亞 的子孫、 比賽 的子孫、
EZRA|2|50|押拿 的子孫、 米烏寧 的子孫、 尼普心 的子孫、
EZRA|2|51|巴卜 的子孫、 哈古巴 的子孫、 哈忽 的子孫、
EZRA|2|52|巴洗律 的子孫、 米希大 的子孫、 哈沙 的子孫、
EZRA|2|53|巴柯 的子孫、 西西拉 的子孫、 答瑪 的子孫、
EZRA|2|54|尼細亞 的子孫、 哈提法 的子孫。
EZRA|2|55|所羅門 僕人的後裔： 瑣太 的子孫、 瑣斐列 的子孫、 比路大 的子孫、
EZRA|2|56|雅拉 的子孫、 達昆 的子孫、 吉德 的子孫、
EZRA|2|57|示法提雅 的子孫、 哈替 的子孫、 玻黑列‧哈斯巴音 的子孫、 亞米 的子孫。
EZRA|2|58|殿役和 所羅門 僕人的後裔共三百九十二名。
EZRA|2|59|從 特‧米拉 、 特‧哈薩 、 基綠 、 亞頓 、 音麥 上來，不能證明他們的父系家族和後裔是否屬 以色列 的如下：
EZRA|2|60|第萊雅 的子孫、 多比雅 的子孫、 尼哥大 的子孫，共六百五十二名。
EZRA|2|61|祭司中， 哈巴雅 的子孫、 哈哥斯 的子孫、 巴西萊 的子孫， 巴西萊 因為娶了 基列 人 巴西萊 的女兒為妻，所以就以此為名。
EZRA|2|62|這些人在族譜之中尋查自己的譜系，卻尋不著，因此算為不潔，不得作祭司。
EZRA|2|63|省長對他們說，不可吃至聖的物，直到有會用烏陵和土明的祭司興起來。
EZRA|2|64|全會眾共有四萬二千三百六十名。
EZRA|2|65|此外，還有他們的僕婢七千三百三十七名，又有歌唱的男女二百名。
EZRA|2|66|他們有七百三十六匹馬，二百四十五匹騾子，
EZRA|2|67|四百三十五匹駱駝，六千七百二十匹驢。
EZRA|2|68|有些族長到了 耶路撒冷 耶和華的殿，為上帝的殿甘心獻上禮物，要在原有的根基上重新建造。
EZRA|2|69|他們量力捐入工程的庫房，有六萬一千達利克 金子，五千彌那銀子，以及一百件祭司的禮服。
EZRA|2|70|於是祭司、 利未 人、百姓中的一些人、歌唱的、門口的守衛、殿役，各住在自己的城裏； 以色列 眾人都住在自己的城裏。
EZRA|3|1|到了七月， 以色列 人住在自己的城裏；那時他們如同一人，聚集在 耶路撒冷 。
EZRA|3|2|約薩達 的兒子 耶書亞 和他的弟兄眾祭司，以及 撒拉鐵 的兒子 所羅巴伯 和他的弟兄，都起來建築 以色列 上帝的壇，要照神人 摩西 律法書上所寫的，在壇上獻燔祭。
EZRA|3|3|他們在原有的根基上築壇，因為他們懼怕鄰邦民族，又在其上向耶和華早晚獻燔祭，
EZRA|3|4|並照律法書上所寫的守住棚節，按數照例每日獻所當獻的燔祭。
EZRA|3|5|此後，他們獻常獻的燔祭，並在初一和耶和華一切分別為聖的節期獻祭，又向耶和華獻各人的甘心祭。
EZRA|3|6|從七月初一起，雖然耶和華殿的根基尚未立定，他們開始向耶和華獻燔祭。
EZRA|3|7|他們把銀子給石匠、木匠，把糧食、酒、油給 西頓 人、 推羅 人，好將香柏樹從 黎巴嫩 浮海運到 約帕 ，是照 波斯 王 居魯士 所允准他們的。
EZRA|3|8|他們到了 耶路撒冷 上帝殿的第二年，二月的時候， 撒拉鐵 的兒子 所羅巴伯 ， 約薩達 的兒子 耶書亞 和其餘的弟兄，就是祭司和 利未 人，以及所有被擄歸回 耶路撒冷 的人，就開工建造；他們派二十歲以上的 利未 人，監督建造耶和華殿的工作。
EZRA|3|9|於是 何達威雅 的後裔，就是 耶書亞 和他的子孫與弟兄、 甲篾 和他的子孫，他們和 利未 人 希拿達 的子孫與弟兄，都起來如同一人，監督那些在上帝殿裏做工的人。
EZRA|3|10|工匠立耶和華殿根基的時候，祭司穿禮服吹號， 利未 人 亞薩 的子孫敲鈸，都照 以色列 王 大衛 親手所定的，站著讚美耶和華。
EZRA|3|11|他們彼此唱和，讚美稱謝耶和華： 「他本為善， 他向 以色列 永施慈愛。」 他們讚美耶和華的時候，眾百姓大聲呼喊，因為耶和華殿的根基已經立定。
EZRA|3|12|然而有許多祭司、 利未 人和族長，就是見過先前那殿的老年人，現在親眼看見這殿立了根基，就大聲哭號，也有許多人大聲歡呼，
EZRA|3|13|百姓不能分辨歡呼的聲音或哭號的聲音，因為百姓大聲呼喊，聲音連遠處都可聽到。
EZRA|4|1|猶大 和 便雅憫 的敵人聽說被擄歸回的人為耶和華－ 以色列 的上帝建造殿宇，
EZRA|4|2|就去見 所羅巴伯 和族長，對他們說：「請讓我們與你們一同建造，因為我們也與你們一樣尋求你們的上帝。自從 亞述 王 以撒‧哈頓 帶我們上這地的日子以來，我們常向上帝獻祭。」
EZRA|4|3|但 所羅巴伯 、 耶書亞 和其餘 以色列 的族長對他們說：「我們建造上帝的殿與你們無關，因為我們要照 波斯 王 居魯士 所吩咐的，自己為耶和華－ 以色列 的上帝協力建造。」
EZRA|4|4|那地的人就在 猶大 百姓建造的時候，使他們的手發軟，擾亂他們。
EZRA|4|5|從 波斯 王 居魯士 年間，直到 波斯 王 大流士 在位的時候，那些人賄賂謀士，要破壞他們的計劃。
EZRA|4|6|亞哈隨魯 在位，他的國度剛開始的時候，他們上書控告 猶大 和 耶路撒冷 的居民。
EZRA|4|7|亞達薛西 年間， 比施蘭 、 米特利達 、 他別 和他們 的同僚上書奏告 波斯 王 亞達薛西 。奏文是用 亞蘭 文寫的，以 亞蘭 文呈上。
EZRA|4|8|利宏 省長、 伸帥 書記也上奏 亞達薛西 王，控告 耶路撒冷 如下
EZRA|4|9|（那時， 利宏 省長、 伸帥 書記和他們其餘的同僚，法官、官員、軍官、 波斯 官員 、 亞基衛 人、 巴比倫 人，和 書珊迦 人，就是 以攔 人 ，
EZRA|4|10|以及被 亞斯那巴 大人遷移、安置在 撒瑪利亞城 和 大河 西邊一帶地方其餘的人。現在 ，
EZRA|4|11|這是他們上奏 亞達薛西 王奏文的抄本）：「 河西 的臣僕上奏 亞達薛西 王，現在
EZRA|4|12|請王知道，從王那裏上到我們這裏的 猶太 人，已經抵達 耶路撒冷 。他們正在重建這反叛惡劣的城，已經完成了城牆，正要修復根基。
EZRA|4|13|如今請王知道，這城若再建造，城牆完工，他們就不再進貢、納糧、繳稅，王的國庫必受虧損。
EZRA|4|14|如今，我們吃的鹽既然全是宮廷的鹽，就不忍見王吃虧，因此奏告於王，
EZRA|4|15|請王考察先王史籍，必會在史籍上查知這城是反叛的城，對列王和各省有害；自古以來，城中常有悖逆的事，因此這城曾被拆毀。
EZRA|4|16|我們謹奏王知，這城若再建造，城牆完工， 河西 之地王就無份了。」
EZRA|4|17|那時王諭覆 利宏 省長、 伸帥 書記和他們其餘的同僚，就是住 撒瑪利亞 和 河西 一帶地方的人，說：「願你們平安。現在
EZRA|4|18|你們所呈給我們的奏本，已經清楚地在我面前讀了。
EZRA|4|19|我已下令考查，得知這城自古以來果然背叛列王，其中常有反叛悖逆的事。
EZRA|4|20|也曾有強大的君王治理 耶路撒冷 ，統管 河西 全地，人就給他們進貢、納糧、繳稅。
EZRA|4|21|現在你們要下令叫這些人停工，使這城不得建造，等到我再降旨。
EZRA|4|22|你們當謹慎辦這事，不可遲延，何必讓損害加重，使王受虧損呢？」
EZRA|4|23|亞達薛西 王上諭的抄本在 利宏 和 伸帥 書記，以及他們的同僚面前宣讀，他們就急忙往 耶路撒冷 去見 猶太 人，用勢力和強權叫他們停工。
EZRA|4|24|於是，在 耶路撒冷 上帝殿的工程就停止了，直停到 波斯 王 大流士 第二年。
EZRA|5|1|那時， 哈該 先知和 易多 的孫子 撒迦利亞 ，兩個先知奉 以色列 上帝的名向 猶大 和 耶路撒冷 的 猶太 人說預言。
EZRA|5|2|於是 撒拉鐵 的兒子 所羅巴伯 和 約薩達 的兒子 耶書亞 起來，開始建造 耶路撒冷 上帝的殿，有上帝的先知在那裏幫助他們。
EZRA|5|3|當時 河西 的 達乃 總督和 示他‧波斯乃 ，以及他們的同僚來對 猶太 人這樣說：「誰降旨讓你們建造這殿，完成這建築呢？」
EZRA|5|4|於是我們告訴他們建造這建築物的人叫甚麼名字。
EZRA|5|5|但上帝的眼目看顧 猶太 人的長老，以致沒有人叫他們停工，直到奏文上告 大流士 ，得著他對這事的回諭。
EZRA|5|6|這是 河西 的 達乃 總督和 示他‧波斯乃 ，以及他們的同僚，就是住 河西 的官員 ，上書奏告 大流士 王的抄本，
EZRA|5|7|他們上書給王的奏文，其中寫著：「願 大流士 王諸事平安。
EZRA|5|8|請王知道，我們往 猶大 省去，到了至大上帝的殿。這殿是用鑿成的石頭建造的，梁木插入牆內。這項工程進行迅速，在他們手中順利。
EZRA|5|9|於是我們問那些長老，對他們這樣說：『誰降旨讓你們建造這殿，完成這建築呢？』
EZRA|5|10|我們又問他們的名字，要記下他們領袖的名字，奏告於王。
EZRA|5|11|他們這樣回答我們說：『我們是天和地之上帝的僕人，重建多年前所建造的殿，就是 以色列 一位偉大的君王建造完成的。
EZRA|5|12|但因我們祖先惹天上的上帝發怒，上帝把他們交在 迦勒底 人 巴比倫 王 尼布甲尼撒 的手中，他就拆毀這殿，又把百姓擄到 巴比倫 。
EZRA|5|13|然而 巴比倫 王 居魯士 元年，他降旨允准建造上帝的這殿。
EZRA|5|14|上帝殿中的金銀器皿，就是 尼布甲尼撒 從 耶路撒冷 殿中掠取帶到 巴比倫 廟裏的， 居魯士 王從 巴比倫 廟裏取出來，交給派為省長，名叫 設巴薩 的，
EZRA|5|15|對他說：可以將這些器皿帶去，放在 耶路撒冷 的殿中，在原處建造上帝的殿。
EZRA|5|16|於是那位 設巴薩 來建立 耶路撒冷 上帝殿的根基。但從那時直到如今，這殿尚未修建完畢。』
EZRA|5|17|現在，王若以為好，請查閱 巴比倫 王的檔案庫，看 居魯士 王有沒有降旨允准在 耶路撒冷 建造上帝的殿。請降旨指示我們王對這件事的心意。」
EZRA|6|1|於是 大流士 王降旨，要尋察典籍庫，就是在 巴比倫 藏檔案之處；
EZRA|6|2|在 瑪代 省 亞馬他城 的宮內尋得一卷，其中這樣寫著，「紀錄如下：
EZRA|6|3|居魯士 王元年，王降旨論到在 耶路撒冷 上帝的殿，要建造這殿作為獻祭之處，堅固它的根基。殿高六十肘，寬六十肘，
EZRA|6|4|要用三層鑿成的石頭，一層木頭 ，經費可出於王的庫房。
EZRA|6|5|至於上帝殿的金銀器皿，就是 尼布甲尼撒 從 耶路撒冷 的殿中掠取帶到 巴比倫 的，必須歸還，帶回 耶路撒冷 的殿中，各按原處放在上帝的殿裏。」
EZRA|6|6|「現在， 河西 的 達乃 總督和 示他‧波斯乃 ，以及他們的同僚，就是住 河西 的官員，你們當遠離那裏。
EZRA|6|7|不要攔阻這上帝殿的工作，任由 猶太 人的省長和長老在原處建造上帝的這殿。
EZRA|6|8|我又降旨，吩咐你們為建造上帝的殿當向 猶太 人的長老這樣行：從王的財產中，由 河西 所繳納的貢銀，迅速支付這些人，免得工程停頓。
EZRA|6|9|他們向天上的上帝獻燔祭所需用的公牛犢、公綿羊、小綿羊，以及麥子、鹽、酒、油，都要照 耶路撒冷 祭司的話，每日供給他們，不得有誤；
EZRA|6|10|好叫他們獻馨香的祭給天上的上帝，又為王和王眾子的壽命祈禱。
EZRA|6|11|我再降旨，無論誰更改這命令，必從他房屋中拆出一根梁木，把他舉起，懸在其上，又使他的房屋為此成為糞堆。
EZRA|6|12|任何王或百姓若伸手更改這命令，拆毀在 耶路撒冷 上帝的這殿，願那立他名在那裏的上帝將他們滅絕。我 大流士 降這諭旨，你們要速速遵行。」
EZRA|6|13|於是， 河西 的 達乃 總督和 示他‧波斯乃 ，以及他們的同僚，急速遵行 大流士 王所頒的命令。
EZRA|6|14|猶太 人的長老因 哈該 先知和 易多 的孫子 撒迦利亞 的預言，就建造這殿，凡事順利。他們遵照 以色列 上帝的命令和 波斯 王 居魯士 、 大流士 、 亞達薛西 的諭旨，建造完畢。
EZRA|6|15|大流士 王第六年，亞達月初三，這殿完工了。
EZRA|6|16|以色列 人、祭司和 利未 人，以及其餘被擄歸回的人都歡歡喜喜地為上帝的這殿行奉獻禮。
EZRA|6|17|他們為這上帝殿的奉獻禮獻了一百頭公牛，二百隻公綿羊，四百隻小綿羊，又照 以色列 支派的數目獻十二隻公山羊，作 以色列 眾人的贖罪祭。
EZRA|6|18|他們派祭司按著班次， 利未 人也按著班次在 耶路撒冷 事奉上帝，正如 摩西 律法書上所寫的。
EZRA|6|19|正月十四日，被擄歸回的人守逾越節。
EZRA|6|20|祭司和 利未 人一同自潔，他們全都潔淨了。 利未 人為被擄歸回的眾人和他們的弟兄眾祭司，並為自己宰逾越節的羔羊。
EZRA|6|21|從被擄之地歸回的 以色列 人，並所有歸附他們、除掉這地外邦人的污穢、尋求耶和華－ 以色列 上帝的人，都吃這羔羊。
EZRA|6|22|他們歡歡喜喜地守除酵節七日，因為耶和華使他們歡喜。耶和華又使 亞述 王的心轉向他們，堅固他們的手，去做上帝－ 以色列 上帝殿的工。
EZRA|7|1|這些事以後， 波斯 王 亞達薛西 在位的時候，有個人叫 以斯拉 ，他是 西萊雅 的兒子， 西萊雅 是 亞撒利雅 的兒子， 亞撒利雅 是 希勒家 的兒子，
EZRA|7|2|希勒家 是 沙龍 的兒子， 沙龍 是 撒督 的兒子， 撒督 是 亞希突 的兒子，
EZRA|7|3|亞希突 是 亞瑪利雅 的兒子， 亞瑪利雅 是 亞撒利雅 的兒子， 亞撒利雅 是 米拉約 的兒子，
EZRA|7|4|米拉約 是 西拉希雅 的兒子， 西拉希雅 是 烏西 的兒子， 烏西 是 布基 的兒子，
EZRA|7|5|布基 是 亞比書 的兒子， 亞比書 是 非尼哈 的兒子， 非尼哈 是 以利亞撒 的兒子， 以利亞撒 是 亞倫 大祭司的兒子。
EZRA|7|6|這 以斯拉 從 巴比倫 上來，他是一個文士，精通耶和華－ 以色列 上帝所賜 摩西 的律法。王允准他一切所求的，因為耶和華－他上帝的手幫助他。
EZRA|7|7|亞達薛西 王第七年，有些 以色列 人、一些祭司、 利未 人、歌唱的、門口的守衛、殿役，上 耶路撒冷 去。
EZRA|7|8|王第七年五月， 以斯拉 到了 耶路撒冷 。
EZRA|7|9|正月初一，他從 巴比倫 起程，五月初一就到了 耶路撒冷 ，因為他上帝施恩的手幫助他。
EZRA|7|10|以斯拉 立志考究遵行耶和華的律法，又將律例典章教導 以色列 人。
EZRA|7|11|亞達薛西 王賜給精通耶和華誡命和 以色列 律例的文士 以斯拉 祭司的諭旨，抄本如下：
EZRA|7|12|「諸王之王 亞達薛西 ，達於精通天上之上帝律法的 以斯拉 祭司文士等等：現在
EZRA|7|13|住在我國中的 以色列 百姓、祭司、 利未 人，凡願意上 耶路撒冷 去的，我降旨准他們與你同去。
EZRA|7|14|既然王與七個謀士派你去，照你手中上帝的律法視察 猶大 和 耶路撒冷 的景況；
EZRA|7|15|你又帶著王和謀士樂意獻給住 耶路撒冷 、 以色列 上帝的金銀，
EZRA|7|16|和你在 巴比倫 全省所得的一切金銀，以及百姓、祭司甘心獻給 耶路撒冷 他們上帝殿的禮物，
EZRA|7|17|那麼，你就當用這銀子急速買公牛、公綿羊、小綿羊，和同獻的素祭、澆酒祭，獻在 耶路撒冷 你們上帝殿的壇上。
EZRA|7|18|剩下的金銀，你和你的弟兄看怎樣好，就怎樣用，但總要遵照你們上帝的旨意。
EZRA|7|19|你要帶著交託給你、在上帝殿中事奉用的器皿，到 耶路撒冷 上帝面前。
EZRA|7|20|你上帝殿裏若再有需用的經費，是你負責供應的，可以從王的寶庫裏支取。
EZRA|7|21|「我 亞達薛西 王又降旨達於 河西 所有的司庫：『精通天上之上帝律法的 以斯拉 祭司文士無論向你們要甚麼，你們要速速辦理，
EZRA|7|22|直至一百他連得銀子，一百柯珥 麥子，一百罷特酒，一百罷特油，鹽不限其數。
EZRA|7|23|凡天上之上帝所吩咐的，當為天上之上帝的殿切實辦理。何必使憤怒臨到王和王眾子的國呢？
EZRA|7|24|我再吩咐你們：至於任何祭司、 利未 人、歌唱的、門口的守衛和殿役，以及在上帝的這殿事奉的人，不可要求他們進貢，納糧，繳稅。』
EZRA|7|25|「你， 以斯拉 啊，要照著你上帝賜你的智慧，指派所有明白你上帝律法的人作官長、審判官，治理 河西 所有的百姓，教導不明白上帝律法的人。
EZRA|7|26|凡不遵行你上帝律法和王命令的人，當速速定他的罪，或處死，或充軍，或抄家，或囚禁。」
EZRA|7|27|以斯拉 說：「耶和華－我們列祖的上帝是應當稱頌的！因他使王起這心願，使 耶路撒冷 耶和華的殿得榮耀，
EZRA|7|28|他又在王和謀士，以及王所有大能的軍官面前施恩於我。我因耶和華－我上帝的手的幫助，得以堅強，從 以色列 中召集領袖，與我一同上來。」
EZRA|8|1|這些是 亞達薛西 王在位的時候，同我從 巴比倫 上來的族長和他們的家譜：
EZRA|8|2|屬 非尼哈 的子孫有 革順 ；屬 以他瑪 的子孫有 但以理 ；屬 大衛 的子孫有 哈突 ；
EZRA|8|3|屬 示迦尼 的子孫；屬 巴錄 的子孫有 撒迦利亞 ，同著他按家譜計算，男丁一百五十人；
EZRA|8|4|屬 巴哈‧摩押 的子孫有 西拉希雅 的兒子 以利約乃 ，同著他有男丁二百人；
EZRA|8|5|屬 薩土 的子孫有 雅哈悉 的兒子 示迦尼 ，同著他有男丁三百人；
EZRA|8|6|屬 亞丁 的子孫有 約拿單 的兒子 以別 ，同著他有男丁五十人；
EZRA|8|7|屬 以攔 的子孫有 亞他利雅 的兒子 耶篩亞 ，同著他有男丁七十人；
EZRA|8|8|屬 示法提雅 的子孫有 米迦勒 的兒子 西巴第雅 ，同著他有男丁八十人；
EZRA|8|9|屬 約押 的子孫有 耶歇 的兒子 俄巴底亞 ，同著他有男丁二百一十八人；
EZRA|8|10|屬 巴尼 的子孫有 約細斐 的兒子 示羅密 ，同著他有男丁一百六十人；
EZRA|8|11|屬 比拜 的子孫有 比拜 的兒子 撒迦利亞 ，同著他有男丁二十八人；
EZRA|8|12|屬 押甲 的子孫有 哈加坦 的兒子 約哈難 ，同著他有男丁一百一十人；
EZRA|8|13|屬 亞多尼干 的子孫，就是晚到的，他們的名字是 以利法列 、 耶利 、 示瑪雅 ，同著他們有男丁六十人；
EZRA|8|14|屬 比革瓦伊 的子孫有 烏太 和 撒刻 ，同著他們有男丁七十人。
EZRA|8|15|我召集這些人在流入 亞哈瓦 的河旁邊，我們在那裏紮營三日。我查看百姓和祭司，發現並沒有 利未 人在那裏，
EZRA|8|16|就派人到 以利以謝 、 亞列 、 示瑪雅 、 以利拿單 、 雅立 、 以利拿單 、 拿單 、 撒迦利亞 、 米書蘭 等領袖，以及 約雅立 和 以利拿單 教師那裏。
EZRA|8|17|我吩咐他們往 迦西斐雅 地方去見那裏的領袖 易多 ，又告訴他們當向 易多 和他的弟兄，就是 迦西斐雅 那地方的殿役說甚麼話，好為我們上帝的殿帶事奉的人來。
EZRA|8|18|蒙我們上帝施恩的手幫助我們，他們在 以色列 的曾孫， 利未 的孫子， 抹利 的後裔中帶了一個精明的人來，就是 示利比 ，還有他的眾子與兄弟共十八人。
EZRA|8|19|另外，還有 哈沙比雅 ，同著他有 米拉利 的子孫 耶篩亞 ，以及他的眾子和兄弟共二十人。
EZRA|8|20|從前 大衛 和眾領袖派殿役服事 利未 人，現在從這殿役中也帶了二百二十人來，全都是按名指定的。
EZRA|8|21|那時，我在 亞哈瓦河 邊宣告禁食，為要在我們上帝面前刻苦己心，求他使我們和我們的孩子，以及一切所有的，都得平坦的道路。
EZRA|8|22|我以求王撥步兵騎兵幫助我們抵擋路上的仇敵為羞愧，因我們曾對王說：「我們上帝施恩的手必幫助凡尋求他的，但他的能力和憤怒必攻擊凡離棄他的。」
EZRA|8|23|我們為此禁食祈求我們的上帝，他就應允我們。
EZRA|8|24|我分派十二位祭司長，就是 示利比 、 哈沙比雅 和與他們一起的兄弟十人，
EZRA|8|25|把王和謀士、軍官，並在那裏的 以色列 眾人為我們上帝殿所獻的金銀和器皿，都秤了交給他們。
EZRA|8|26|我秤了交在他們手中的有六百五十他連得銀子，一百他連得銀器，一百他連得金子，
EZRA|8|27|二十個金碗，值一千達利克，上等光亮的銅器皿兩個，珍貴如金。
EZRA|8|28|我對他們說：「你們歸耶和華為聖，器皿也歸為聖；金銀是甘心獻給耶和華－你們列祖之上帝的。
EZRA|8|29|你們要警醒看守，直到你們在祭司長和 利未 族長，以及 以色列 的各族長面前，在 耶路撒冷 耶和華殿的庫房內，把這些過了秤。」
EZRA|8|30|於是，祭司和 利未 人把秤過的金銀和器皿接過來，要帶到 耶路撒冷 我們上帝的殿裏。
EZRA|8|31|正月十二日，我們從 亞哈瓦河 邊起行，要往 耶路撒冷 去。我們上帝的手保佑我們，救我們脫離仇敵和路上埋伏之人的手。
EZRA|8|32|我們到了 耶路撒冷 ，在那裏住了三日。
EZRA|8|33|第四日，金銀和器皿都在我們上帝的殿裏過了秤，交在 烏利亞 的兒子 米利末 祭司的手中。同著他的有 非尼哈 的兒子 以利亞撒 ，還有 利未 人 耶書亞 的兒子 約撒拔 和 賓內 的兒子 挪亞底 。
EZRA|8|34|那時，這一切都點過秤過了，重量全寫在冊上。
EZRA|8|35|從被擄之地歸回的人向 以色列 的上帝獻燔祭，為 以色列 眾人獻十二頭公牛，九十六隻公綿羊，七十七隻小綿羊，又獻十二隻公山羊作贖罪祭，這些全都是獻給耶和華的燔祭。
EZRA|8|36|被擄歸回的人把王的諭旨交給王的總督與 河西 的省長，他們就支助百姓和上帝的殿。
EZRA|9|1|這些事完成以後，眾領袖來接近我，說：「 以色列 百姓、祭司和 利未 人沒有棄絕 迦南 人、 赫 人、 比利洗 人、 耶布斯 人、 亞捫 人、 摩押 人、 埃及 人和 亞摩利 人等列邦民族所行可憎的事。
EZRA|9|2|因他們為自己和兒子娶了這些外邦女子，以致聖潔的種籽和列邦民族混雜，而且領袖和官長在這事上是罪魁。」
EZRA|9|3|我一聽見這事，就撕裂衣服和外袍，拔了頭髮和鬍鬚，驚惶地坐著。
EZRA|9|4|凡為 以色列 上帝言語戰兢的人，都因被擄歸回之人所犯的罪，聚集到我這裏來。我驚惶地坐著，直到獻晚祭的時候。
EZRA|9|5|獻晚祭的時候我從愁煩中起來，穿著撕裂的衣服和外袍，雙膝跪下，向耶和華－我的上帝舉手，
EZRA|9|6|說： 「我的上帝啊，我抱愧蒙羞，不敢向你－我的上帝仰面，因為我們的罪孽多到滅頂，我們的罪惡滔天。
EZRA|9|7|從我們祖先的日子直到今日，我們的罪惡深重；因我們的罪孽，我們和君王、祭司都交在鄰國諸王的手中，被殺害，擄掠，搶奪，臉上蒙羞，正如今日的景況。
EZRA|9|8|現在耶和華－我們的上帝暫且向我們施恩，為我們留下一些殘存之民，使我們如釘子釘在他的聖所，讓我們的上帝光照我們的眼目，使我們在受轄制之中稍微復興。
EZRA|9|9|我們是奴僕，然而在受轄制之中，我們的上帝沒有丟棄我們，在 波斯 諸王面前向我們施恩，叫我們復興，能重建我們上帝的殿，修補毀壞之處，使我們在 猶大 和 耶路撒冷 有城牆。
EZRA|9|10|「我們的上帝啊，既然如此，現在我們還有甚麼話可說呢？因為我們離棄了你的誡命，
EZRA|9|11|就是你藉你僕人眾先知所吩咐的，說：『你們要去得為業之地是污穢之地，因列邦民族的污穢和可憎的事，叫這地從這邊到那邊都充滿了污穢。
EZRA|9|12|現在，不可把你們的女兒嫁給他們的兒子，也不可為你們的兒子娶他們的女兒，永不可求他們的平安和他們的利益，這樣你們就可以強盛，吃這地的美物，並把這地留給你們的子孫永遠為業。』
EZRA|9|13|我們因自己的惡行和大罪，遭遇這一切的事，但你－我們的上帝懲罰我們輕於我們罪所當得的，又為我們留下這些殘存之民。
EZRA|9|14|我們豈可再違背你的誡命，與行這些可憎之事的民族結親呢？若我們這樣行，你豈不向我們發怒，將我們滅絕，以致沒有一個餘民或殘存之民嗎？
EZRA|9|15|耶和華－ 以色列 的上帝啊，你是公義的，我們才能剩下這些殘存之民，正如今日的景況。看哪，我們在你面前有罪惡，因此無人能在你面前站立得住。」
EZRA|10|1|以斯拉 禱告，認罪，哭泣，俯伏在上帝殿前的時候，有 以色列 中的男女和孩童聚集到 以斯拉 那裏，成了一個盛大的會，百姓無不痛哭。
EZRA|10|2|以攔 的子孫， 耶歇 的兒子 示迦尼 對 以斯拉 說：「我們娶了這地的外邦女子，干犯了我們的上帝，然而現在 以色列 人在這事上還有指望。
EZRA|10|3|現在，我們要與我們的上帝立約，送走所有的妻子和她們所生的，照著主和那些因我們上帝誡命戰兢之人所議定的，按律法去行。
EZRA|10|4|起來，這是你當辦的事，我們必支持你，你當奮勇而行。」
EZRA|10|5|以斯拉 就起來，叫祭司長和 利未 人，以及 以色列 眾人起誓，要照這話去做；他們就起了誓。
EZRA|10|6|以斯拉 從上帝殿前起來，進入 以利亞實 的兒子 約哈難 的屋裏，到了那裏不吃飯，也不喝水，為被擄歸回之人所犯的罪悲傷。
EZRA|10|7|他們通告 猶大 和 耶路撒冷 ，叫所有被擄歸回的人聚集在 耶路撒冷 。
EZRA|10|8|凡不遵照領袖和長老所議定，三日之內不來的，就必毀壞他所有的財產，把他從被擄歸回之人的會中開除。
EZRA|10|9|於是， 猶大 和 便雅憫 眾人三日之內都聚集在 耶路撒冷 。那時是九月，那月的二十日，眾百姓坐在上帝殿前的廣場，因這事，又因下大雨，就都戰抖。
EZRA|10|10|以斯拉 祭司站起來，對他們說：「你們有罪了，因為你們娶了外邦女子，增添 以色列 的罪惡。
EZRA|10|11|現在當向耶和華－你們列祖的上帝認罪，遵行他的旨意，離開這地的百姓和外邦女子。」
EZRA|10|12|全會眾大聲回答說：「好！我們必照著你的話去做。
EZRA|10|13|只是百姓眾多，又逢大雨的季節，我們沒有氣力站在外面；這也不是一兩天可以辦完的事，因我們在這事上犯了大罪。
EZRA|10|14|讓我們的領袖代表全會眾留在那裏。我們城鎮中凡娶外邦女子的，當按所定的日期，會同本城的長老和審判官前來，直到辦完這事，上帝的烈怒轉離我們 。」
EZRA|10|15|惟有 亞撒黑 的兒子 約拿單 ， 特瓦 的兒子 雅哈謝 反對這事，並有 米書蘭 和 利未 人 沙比太 支持他們。
EZRA|10|16|被擄歸回的人就如此做了。 以斯拉 祭司按著父家指名選派一些族長 。十月初一，他們一同坐下來查辦這事，
EZRA|10|17|到正月初一，才查清所有娶外邦女子的人數。
EZRA|10|18|在祭司中查出娶外邦女子的： 耶書亞 的子孫中，有 約薩達 的兒子，和他兄弟 瑪西雅 、 以利以謝 、 雅立 、 基大利 ，
EZRA|10|19|他們承諾要送走他們的妻子。他們因有罪，就獻羊群中的一隻公綿羊贖罪；
EZRA|10|20|音麥 的子孫中，有 哈拿尼 、 西巴第雅 ；
EZRA|10|21|哈琳 的子孫中，有 瑪西雅 、 以利雅 、 示瑪雅 、 耶歇 、 烏西雅 ；
EZRA|10|22|巴施戶珥 的子孫中，有 以利約乃 、 瑪西雅 、 以實瑪利 、 拿坦業 、 約撒拔 、 以利亞薩 。
EZRA|10|23|利未 人中，有 約撒拔 、 示每 、 基拉雅 ， 基拉雅 就是 基利他 ，還有 毗他希雅 、 猶大 、 以利以謝 。
EZRA|10|24|歌唱的人中有 以利亞實 。門口的守衛中，有 沙龍 、 提聯 、 烏利 。
EZRA|10|25|以色列 人 巴錄 的子孫中，有 拉米 、 耶西雅 、 瑪基雅 、 米雅民 、 以利亞撒 、 瑪基雅 、 比拿雅 。
EZRA|10|26|以攔 的子孫中，有 瑪他尼 、 撒迦利亞 、 耶歇 、 押底 、 耶列末 、 以利雅 。
EZRA|10|27|薩土 的子孫中，有 以利約乃 、 以利亞實 、 瑪他尼 、 耶列末 、 撒拔 、 亞西撒 。
EZRA|10|28|比拜 的子孫中，有 約哈難 、 哈拿尼雅 、 薩拜 、 亞勒 。
EZRA|10|29|巴尼 的子孫中，有 米書蘭 、 瑪鹿 、 亞大雅 、 雅述 、 示押 、 拉末 。
EZRA|10|30|巴哈‧摩押 的子孫中，有 阿底拿 、 基拉 、 比拿雅 、 瑪西雅 、 瑪他尼 、 比撒列 、 賓內 、 瑪拿西 。
EZRA|10|31|哈琳 的子孫中，有 以利以謝 、 伊示雅 、 瑪基雅 、 示瑪雅 、 西緬 、
EZRA|10|32|便雅憫 、 瑪鹿 、 示瑪利雅 。
EZRA|10|33|哈順 的子孫中，有 瑪特乃 、 瑪達他 、 撒拔 、 以利法列 、 耶利買 、 瑪拿西 、 示每 。
EZRA|10|34|巴尼 的子孫中，有 瑪玳 、 暗蘭 、 烏益 、
EZRA|10|35|比拿雅 、 比底雅 、 基祿 、
EZRA|10|36|瓦尼雅 、 米利末 、 以利亞實 、
EZRA|10|37|瑪他尼 、 瑪特乃 、 雅掃 、
EZRA|10|38|巴尼 、 賓內 、 示每 、
EZRA|10|39|示利米雅 、 拿單 、 亞大雅 、
EZRA|10|40|瑪拿底拜 、 沙賽 、 沙賴 、
EZRA|10|41|亞薩利 、 示利米雅 、 示瑪利雅 、
EZRA|10|42|沙龍 、 亞瑪利雅 、 約瑟 。
EZRA|10|43|尼波 的子孫中，有 耶利 、 瑪他提雅 、 撒拔 、 西比拿 、 雅玳 、 約珥 、 比拿雅 。
EZRA|10|44|這些人全都娶了外邦女子，其中也有生了兒女的 。
NEH|1|1|哈迦利亞 的兒子 尼希米 的言語如下： 亞達薛西 王二十年基斯流月，我在 書珊 城堡中。
NEH|1|2|那時，我有一個兄弟 哈拿尼 ，同幾個人從 猶大 來。我問他們那些被擄歸回、剩下殘存的 猶太 人和 耶路撒冷 的情況。
NEH|1|3|他們對我說：「那些被擄歸回剩下的餘民在 猶大 省那裏遭大難，受凌辱； 耶路撒冷 的城牆被拆毀，城門被火焚燒。」
NEH|1|4|我聽見這話，就坐下哭泣，悲哀幾日，在天上的上帝面前禁食祈禱，
NEH|1|5|說：「唉，耶和華－天上大而可畏的上帝，向愛你、守你誡命的人守約施慈愛的上帝啊，
NEH|1|6|願你睜眼看，側耳聽你僕人今日晝夜在你面前，為你眾僕人 以色列 人的祈禱，承認我們 以色列 人向你所犯的罪；我與我父家都犯了罪。
NEH|1|7|我們向你所行的非常敗壞，沒有遵守你吩咐你僕人 摩西 的誡命、律例、典章。
NEH|1|8|求你記念所吩咐你僕人 摩西 的話，說：『你們若犯罪，我就把你們分散在萬民中；
NEH|1|9|但你們若歸向我，謹守遵行我的誡命，你們被趕散的人雖在天涯，我也必從那裏將他們召集回來，帶到我所選擇立為我名居所的地方。』
NEH|1|10|他們是你的僕人和你的百姓，是你用大力和大能的手所救贖的。
NEH|1|11|唉，主啊，求你側耳聽你僕人的祈禱，聽喜愛敬畏你名眾僕人的祈禱，使你僕人今日亨通，在這人面前蒙恩。」 我是王的酒政。
NEH|2|1|亞達薛西 王二十年尼散月，酒擺在王面前 ，我拿起酒來奉給王。我在王面前從來沒有愁容。
NEH|2|2|王對我說：「你既沒有病，為甚麼面帶愁容呢？這不是別的，必是你心中愁煩。」於是我非常懼怕。
NEH|2|3|我對王說：「願王萬歲！我祖先墳墓所在的那城荒涼，城門被火焚燒，我豈能面無愁容呢？」
NEH|2|4|王對我說：「你想求甚麼？」於是我向天上的上帝祈禱。
NEH|2|5|我對王說：「王若以為好，僕人若在王面前蒙恩，求王差遣我往 猶大 ，到我祖先墳墓所在的那城去，我好重新建造。」
NEH|2|6|那時王后坐在王的旁邊，王對我說：「你要去多久？幾時回來？」王看這事為好，就派我去。我給王定了日期。
NEH|2|7|我又對王說：「王若以為好，求王賜我詔書，通知 河西 的省長准我經過，直到 猶大 ；
NEH|2|8|又賜詔書，通知管理王園林的 亞薩 ，叫他給我木材，作為殿的營樓之門、城牆，和我自己要住的房屋的橫梁。」王就允准我，因為我上帝施恩的手幫助我。
NEH|2|9|王派了軍官和騎兵護送我。我到了 河西 的省長那裏，將王的詔書交給他們。
NEH|2|10|和倫 人 參巴拉 和作臣僕的 亞捫 人 多比雅 ，聽見有人來為 以色列 人爭取利益，就很惱怒。
NEH|2|11|我到了 耶路撒冷 ，在那裏停留了三天。
NEH|2|12|夜間我和跟隨我的幾個人起來；但上帝感動我心要為 耶路撒冷 做的事，我並沒有告訴人。只有我自己騎的牲口，沒有別的牲口在我那裏。
NEH|2|13|當夜，我出了 谷門 ，往 野狗泉 去，到了 糞廠門 ，察看 耶路撒冷 的城牆，城牆被拆毀，城門被火焚燒。
NEH|2|14|我又往前，到了 泉門 ，又到 王池 ，但所騎的牲口沒有地方可以過去。
NEH|2|15|於是我夜間沿溪而上，察看城牆，又轉身進入 谷門 ，就回來了。
NEH|2|16|我往哪裏去，我做甚麼事，官長都不知道。我也沒有告訴 猶大 人、祭司、貴族、官長和其餘做工的人。
NEH|2|17|以後，我對他們說：「我們所遭的難， 耶路撒冷 怎樣荒涼，城門被火焚燒，你們都看見了。來吧，讓我們重建 耶路撒冷 的城牆，免得再受凌辱！」
NEH|2|18|我告訴他們我上帝施恩的手怎樣幫助我，以及王向我所說的話。他們就說：「我們起來建造吧！」於是他們使自己的手堅強，做這美好的工作。
NEH|2|19|但 和倫 人 參巴拉 、作臣僕的 亞捫 人 多比雅 和 阿拉伯 人 基善 聽見就嗤笑我們，藐視我們，說：「你們所做的這事是甚麼呢？要背叛王嗎？」
NEH|2|20|我回答他們的話，對他們說：「天上的上帝必使我們亨通。我們作他僕人的，要起來建造；你們卻在 耶路撒冷 無份、無權、無名號 。」
NEH|3|1|那時， 以利亞實 大祭司和他的弟兄眾祭司起來建立 羊門 ，將門分別為聖，安立門扇，直到 哈米亞樓 。他們又將它分別為聖，直到 哈楠業樓 。
NEH|3|2|在他旁邊建造的是 耶利哥 人。在他旁邊建造的是 音利 的兒子 撒刻 。
NEH|3|3|哈西拿 的子孫建立 魚門 ，架橫梁、安門扇，裝閂和鎖。
NEH|3|4|在他們旁邊修造的是 哈哥斯 的孫子， 烏利亞 的兒子 米利末 。在他們旁邊修造的是 米示薩別 的孫子， 比利迦 的兒子 米書蘭 。在他們旁邊修造的是 巴拿 的兒子 撒督 。
NEH|3|5|在他們旁邊修造的是 提哥亞 人；但是他們的貴族不用肩 扛他們主人的工作。
NEH|3|6|巴西亞 的兒子 耶何耶大 與 比所玳 的兒子 米書蘭 修造 古門 ，架橫梁，安門扇，裝閂和鎖。
NEH|3|7|在他們旁邊修造的是 基遍 人 米拉提 、 米倫 人 雅頓 、 基遍 人，和 河西 總督所管的 米斯巴 人。
NEH|3|8|在他旁邊修造的是 哈海雅 的兒子 烏薛 銀匠。在他旁邊修造的是做香料的 哈拿尼雅 。他們修復 耶路撒冷 ，直到 寬牆 。
NEH|3|9|在他們旁邊修造的是管理 耶路撒冷 城區的一半、 戶珥 的兒子 利法雅 。
NEH|3|10|在他們旁邊的是 哈路抹 的兒子 耶大雅 在自己房屋的對面修造。在他旁邊修造的是 哈沙尼 的兒子 哈突 。
NEH|3|11|哈琳 的兒子 瑪基雅 和 巴哈‧摩押 的兒子 哈述 修造下一段和 爐樓 。
NEH|3|12|在他旁邊修造的是管理 耶路撒冷 城區的另一半、 哈羅黑 的兒子 沙龍 和他的女兒們。
NEH|3|13|哈嫩 和 撒挪亞 的居民修造 谷門 ；他們立門，安門扇，裝閂和鎖，又修造城牆一千肘，直到 糞廠門 。
NEH|3|14|管理 伯‧哈基琳 區、 利甲 的兒子 瑪基雅 修造 糞廠門 ；他立門，安門扇，裝閂和鎖。
NEH|3|15|管理 米斯巴 區、 各‧荷西 的兒子 沙崙 修造 泉門 ；他立門，蓋門頂，安門扇，裝閂和鎖，又修造靠近王的花園 西羅亞池 的城牆，直到那從 大衛城 下來的臺階。
NEH|3|16|接續他修造的是管理 伯‧夙 區的一半、 押卜 的兒子 尼希米 ，直到 大衛 墳地的對面，又到人造池，到達勇士的房屋。
NEH|3|17|接續他修造的是 利未 人 巴尼 的兒子 利宏 。在他旁邊的是管理 基伊拉 區一半的 哈沙比雅 為本區修造。
NEH|3|18|接續他修造的是他們弟兄中管理 基伊拉 區的另一半、 希拿達 的兒子 賓內 。
NEH|3|19|在他旁邊的是管理 米斯巴 、 耶書亞 的兒子 以謝珥 修造武庫的上坡對面、城牆轉彎處的那一段。
NEH|3|20|接續他的是 薩拜 的兒子 巴錄 竭力修造下一段，從轉彎處，直到 以利亞實 大祭司的府門。
NEH|3|21|接續他的是 哈哥斯 的孫子， 烏利亞 的兒子 米利末 修造下一段，從 以利亞實 的府門，直到 以利亞實 府的盡頭。
NEH|3|22|接續他修造的是住平原的祭司。
NEH|3|23|接續他的是 便雅憫 與 哈述 在自己房屋的對面修造。接續他的是 亞難尼 的孫子， 瑪西雅 的兒子 亞撒利雅 在自己房屋的旁邊修造。
NEH|3|24|接續他的是 希拿達 的兒子 賓內 修造下一段，從 亞撒利雅 的房屋直到轉彎處，又到城角。
NEH|3|25|烏賽 的兒子 巴拉 修造轉彎處的對面和靠近護衛院、王宮上層凸出來的城樓。接續他的是 巴錄 的兒子 毗大雅 ，
NEH|3|26|（殿役住在 俄斐勒 ，直到朝東 水門 的對面和凸出來的城樓。）
NEH|3|27|接續他的是 提哥亞 人又修造一段，對著那凸出來的大城樓，直到 俄斐勒 的城牆。
NEH|3|28|從 馬門 往上，祭司各在自己房屋的對面修造。
NEH|3|29|接續他的是 音麥 的兒子 撒督 在自己房屋的對面修造。接續他修造的是 東門 的守衛、 示迦尼 的兒子 示瑪雅 。
NEH|3|30|接續他的是 示利米雅 的兒子 哈拿尼雅 和 薩拉 的第六個兒子 哈嫩 修造下一段。接續他的是 比利迦 的兒子 米書蘭 在自己房屋的對面修造。
NEH|3|31|接續他的是 瑪基雅 銀匠修造，直到殿役和商人的房屋，對著 集合門 ，直到角樓。
NEH|3|32|銀匠與商人在角樓和 羊門 之間修造。
NEH|4|1|參巴拉 聽見我們建造城牆就發怒，非常惱恨，並嗤笑 猶太 人。
NEH|4|2|他對他的弟兄和 撒瑪利亞 的軍兵說：「這些軟弱的 猶太 人做甚麼呢？要為自己重建嗎 ？要獻祭嗎？要一日完工嗎？要使土堆裏火燒過的石頭再有用嗎？」
NEH|4|3|亞捫 人 多比雅 在一旁說：「他們所修造的石牆，就是狐狸上去也必崩裂。」
NEH|4|4|我們的上帝啊，求你垂聽，因為我們被藐視。求你使他們的毀謗歸於他們自己頭上，使他們在被擄之地成為掠物。
NEH|4|5|不要遮掩他們的罪孽，不要使他們的罪惡從你面前塗去，因為他們在修造的人前面惹你發怒。
NEH|4|6|這樣，我們修造城牆，整個城牆就連接起來，到一半高，因為百姓一心做工。
NEH|4|7|參巴拉 、 多比雅 、 阿拉伯 人、 亞捫 人和 亞實突 人聽見 耶路撒冷 城牆正在修造，破裂的地方開始進行修補，就非常憤怒。
NEH|4|8|大家同謀要來攻打 耶路撒冷 ，使城混亂。
NEH|4|9|然而，我們向我們的上帝禱告，又因他們的緣故，就派人站崗，晝夜防備他們。
NEH|4|10|但 猶大 有話說： 「扛抬的人力氣衰弱， 瓦礫太多， 我們自己不可能 建造城牆。」
NEH|4|11|我們的敵人說：「趁他們不知道，看不見的時候，我們進入他們中間，殺了他們，使工作停止。」
NEH|4|12|那靠近敵人居住的 猶太 人十次從各處來見我們，說：「你們必須回到我們那裏。」
NEH|4|13|我叫百姓站在城牆後邊低窪的空處，使百姓各按宗族站著，拿刀、拿槍、拿弓。
NEH|4|14|我察看了，就起來對貴族、官長和其餘的百姓說：「不要怕他們！當記得主是大而可畏的。你們要為你們的弟兄、兒女、妻子、家園爭戰。」
NEH|4|15|仇敵聽見我們知道了他們的計謀，上帝也破壞他們的計謀，我們就都回到城牆那裏，各做各的工。
NEH|4|16|從那日起，我的僕人一半做工，一半拿槍、拿盾牌、拿弓、穿鎧甲，官長都站在 猶大 全家的後邊。
NEH|4|17|他們建造城牆；扛抬材料的人扛抬的時候，一手做工，一手拿兵器。
NEH|4|18|建造的人都腰間佩刀建造，吹角的人在我旁邊。
NEH|4|19|我對貴族、官長和其餘的百姓說：「這工程浩大，範圍遼闊，我們在城牆上彼此相離很遠。
NEH|4|20|你們一聽見角聲在哪裏，就聚集到我們那裏去。我們的上帝必為我們爭戰。」
NEH|4|21|於是，我們做這工程，一半的人拿槍，從天亮直到星宿出現的時候。
NEH|4|22|那時，我又對百姓說：「各人和他的僕人當在 耶路撒冷 過夜，好為我們夜間守衛，白晝做工。」
NEH|4|23|這樣，我和弟兄僕人，以及跟從我的衛兵都不脫衣服，各人打水時 也拿著自己的兵器。
NEH|5|1|百姓和他們的妻子大大呼號，埋怨他們的弟兄 猶太 人。
NEH|5|2|有的說：「我們和兒女人口眾多，必須得糧食吃，才能活下去。」
NEH|5|3|有的說：「我們典押了田地、葡萄園、房屋，才得糧食充飢。」
NEH|5|4|有的說：「我們借了錢付田地和葡萄園的稅給王。
NEH|5|5|現在，我們的身體與我們弟兄的身體是一樣的，我們的兒女與他們的兒女沒有差別。看哪，我們卻要迫使兒女作人的奴婢。我們有些女兒已被搶走了，我們卻無能為力，因為我們的田地和葡萄園已經歸了別人。」
NEH|5|6|我聽見他們的呼號和這些話，就非常憤怒。
NEH|5|7|我心裏作了決定，就斥責貴族和官長，對他們說：「你們各人借錢給弟兄，竟然索取利息！」於是我召開大會攻擊他們。
NEH|5|8|我對他們說：「我們已盡力贖回我們的弟兄，就是賣到列國的 猶太 人；你們還要賣弟兄，讓我們去買回來嗎？」他們就靜默不語，無話可答。
NEH|5|9|我又說：「你們做的這事不對！你們行事不是應該敬畏我們的上帝，免得列國我們的仇敵毀謗我們嗎？
NEH|5|10|我和我的弟兄僕人也要把銀錢糧食借給百姓，大家都當免除利息。
NEH|5|11|就在今日，你們要把他們的田地、葡萄園、橄欖園、房屋，以及向他們所取銀錢的利息 、糧食、新酒和新油都歸還他們。」
NEH|5|12|貴族和官長說：「我們必歸還，不再向他們索取，必照你所說的去做。」我就召了祭司來，叫貴族和官長起誓，必照這話去做。
NEH|5|13|我也抖著胸前的衣袋，說：「凡不實行這話的，願上帝照樣抖他離開他的家和他勞碌得來的，直到抖空了。」全會眾都說：「阿們！」又讚美耶和華。百姓就照著這話去做。
NEH|5|14|自從我奉派作 猶大 地省長的那日，就是從 亞達薛西 王二十年直到三十二年，共十二年之久，我與我弟兄都沒有吃省長的俸祿。
NEH|5|15|在我以前的省長加重百姓的負擔，向百姓索取糧食和酒，以及四十舍客勒銀子 ，甚至他們的僕人也轄制百姓，但我因敬畏上帝不這樣做。
NEH|5|16|我也努力修造城牆。我們並沒有購置田地，我所有的僕人也都聚集在那裏做工。
NEH|5|17|除了從四圍列國來的人以外，有 猶太 人和官長一百五十人與我同席。
NEH|5|18|每日預備一頭公牛，六隻肥羊，又為我預備飛禽；每十日一次多多預備各樣的酒。雖然如此，我並不索取省長的俸祿，因為這百姓負的勞役很重。
NEH|5|19|我的上帝啊，求你記念我為這百姓所做的一切，施恩於我。
NEH|6|1|參巴拉 、 多比雅 、 阿拉伯 人 基善 和我們其餘的仇敵聽見我已經建造了城牆，沒有破裂之處在其中，那時我還沒有在城門安門扇；
NEH|6|2|參巴拉 和 基善 就派人來見我，說：「請你來，我們在 阿挪 平原的村莊見面。」其實，他們想要害我。
NEH|6|3|於是我派使者到他們那裏，說：「我正在進行大的工程，不能下去。我怎麼能離開，下去見你們，而讓工程停頓呢？」
NEH|6|4|他們這樣派人來見我四次，我都用這話回答他們。
NEH|6|5|參巴拉 第五次同樣派僕人來見我，手裏拿著未封的信，
NEH|6|6|信上寫著：「列國中有風聲， 基善 也說，你和 猶太 人謀反，所以你建造城牆。據說，你要作他們的王，
NEH|6|7|並且你派先知在 耶路撒冷 指著你宣講說，『在 猶大 有王。』如今這些話必傳給王知，現在請你來，我們一起商議。」
NEH|6|8|我就派人到他那裏，說：「你所說的這些事，一概沒有，是你心裏捏造的。」
NEH|6|9|他們全都要使我們懼怕，說：「他們的手必軟弱，不能工作，以致不能完工。」現在，求你堅固我的手。
NEH|6|10|我到了 米希大別 的孫子， 第來雅 的兒子 示瑪雅 家裏；那時，他閉門不出。他說：「我們可以在上帝的殿裏，就在殿的中間會面，鎖住殿門，因為他們要來殺你，要在夜裏來殺你。」
NEH|6|11|我說：「像我這樣的人豈會逃跑呢？像我這樣的人豈能進入殿裏保全生命呢？我不進去！」
NEH|6|12|我看清楚了，看哪，上帝並沒有派他，是他自己說預言攻擊我，是 多比雅 和 參巴拉 收買了他；
NEH|6|13|收買他的目的是要叫我懼怕，依從他犯罪，留下一個壞名聲，好讓他們毀謗我。
NEH|6|14|我的上帝啊，求你記得 多比雅 、 參巴拉 、 挪亞底 女先知和其餘的先知，因他們行這些事，要叫我懼怕。
NEH|6|15|以祿月二十五日，城牆修完了，共修了五十二天。
NEH|6|16|我們所有的仇敵聽見了，四圍的列國就懼怕，愁眉不展，因為他們知道這工作得以完成，是出於我們的上帝。
NEH|6|17|而且，在那些日子， 猶大 的貴族屢次寄信給 多比雅 ， 多比雅 也回信給他們。
NEH|6|18|在 猶大 有許多人與 多比雅 結盟，因為他是 亞拉 的兒子 示迦尼 的女婿，並且他的兒子 約哈難 娶了 比利迦 的兒子 米書蘭 的女兒。
NEH|6|19|他們也在我面前說 多比雅 的好話，又把我的話傳給他。 多比雅 常寄信來，要叫我懼怕。
NEH|7|1|城牆修完，我安了門扇，門口的守衛、歌唱的和 利未 人都已派定。
NEH|7|2|我吩咐我的兄弟 哈拿尼 和城堡的官長 哈拿尼雅 管理 耶路撒冷 ，因為 哈拿尼雅 是一個忠信的人，敬畏上帝過於眾人。
NEH|7|3|我對他們說：「等到太陽熱的時候才可開 耶路撒冷 的城門；要派 耶路撒冷 的居民，各按班次在自己房屋的前面站崗。他們還在站崗的時候，就要關門上閂。」
NEH|7|4|城又寬又大，城中的百姓卻稀少，房屋也還沒有建造。
NEH|7|5|我的上帝感動我的心，我就召集貴族、官長和百姓，要登記家譜。我找到第一次上來之人的家譜，發現上面寫著：
NEH|7|6|這些是從被擄之地上來的省民， 巴比倫 王 尼布甲尼撒 把他們擄去，他們重返 耶路撒冷 和 猶大 ，各歸本城。
NEH|7|7|他們是同 所羅巴伯 、 耶書亞 、 尼希米 、 亞撒利雅 、 拉米 、 拿哈瑪尼 、 末底改 、 必珊 、 米斯毗列 、 比革瓦伊 、 尼宏 、 巴拿 一起回來的。 以色列 百姓的人數如下：
NEH|7|8|巴錄 的子孫二千一百七十二名；
NEH|7|9|示法提雅 的子孫三百七十二名；
NEH|7|10|亞拉 的子孫六百五十二名；
NEH|7|11|巴哈‧摩押 的後裔，就是 耶書亞 和 約押 的子孫二千八百一十八名；
NEH|7|12|以攔 的子孫一千二百五十四名；
NEH|7|13|薩土 的子孫八百四十五名；
NEH|7|14|薩改 的子孫七百六十名；
NEH|7|15|賓內 的子孫六百四十八名；
NEH|7|16|比拜 的子孫六百二十八名；
NEH|7|17|押甲 的子孫二千三百二十二名；
NEH|7|18|亞多尼干 的子孫六百六十七名；
NEH|7|19|比革瓦伊 的子孫二千零六十七名；
NEH|7|20|亞丁 的子孫六百五十五名；
NEH|7|21|亞特 的後裔，就是 希西家 的子孫九十八名；
NEH|7|22|哈順 的子孫三百二十八名；
NEH|7|23|比賽 的子孫三百二十四名；
NEH|7|24|哈拉 的子孫一百一十二名；
NEH|7|25|基遍 人九十五名；
NEH|7|26|伯利恆 人和 尼陀法 人共一百八十八名；
NEH|7|27|亞拿突 人一百二十八名；
NEH|7|28|伯‧亞斯瑪弗 人四十二名；
NEH|7|29|基列‧耶琳 人、 基非拉 人、 比錄 人共七百四十三名；
NEH|7|30|拉瑪 人和 迦巴 人共六百二十一名；
NEH|7|31|默瑪 人一百二十二名；
NEH|7|32|伯特利 人和 艾 人共一百二十三名；
NEH|7|33|別的 尼波 人五十二名；
NEH|7|34|另一個 以攔 子孫一千二百五十四名；
NEH|7|35|哈琳 的子孫三百二十名；
NEH|7|36|耶利哥 人三百四十五名；
NEH|7|37|羅德 人、 哈第 人、 阿挪 人共七百二十一名；
NEH|7|38|西拿 人三千九百三十名。
NEH|7|39|祭司： 耶書亞 家， 耶大雅 的子孫九百七十三名；
NEH|7|40|音麥 的子孫一千零五十二名；
NEH|7|41|巴施戶珥 的子孫一千二百四十七名；
NEH|7|42|哈琳 的子孫一千零一十七名。
NEH|7|43|利未 人： 何達威 的後裔，就是 耶書亞 和 甲篾 的子孫七十四名。
NEH|7|44|歌唱的： 亞薩 的子孫一百四十八名。
NEH|7|45|門口的守衛： 沙龍 的子孫、 亞特 的子孫、 達們 的子孫、 亞谷 的子孫、 哈底大 的子孫、 朔拜 的子孫，共一百三十八名。
NEH|7|46|殿役： 西哈 的子孫、 哈蘇巴 的子孫、 答巴俄 的子孫、
NEH|7|47|基綠 的子孫、 西亞 的子孫、 巴頓 的子孫、
NEH|7|48|利巴拿 的子孫、 哈迦巴 的子孫、 薩買 的子孫、
NEH|7|49|哈難 的子孫、 吉德 的子孫、 迦哈 的子孫、
NEH|7|50|利亞雅 的子孫、 利汛 的子孫、 尼哥大 的子孫、
NEH|7|51|迦散 的子孫、 烏撒 的子孫、 巴西亞 的子孫、
NEH|7|52|比賽 的子孫、 米烏寧 的子孫、 尼普心 的子孫、
NEH|7|53|巴卜 的子孫、 哈古巴 的子孫、 哈忽 的子孫、
NEH|7|54|巴洗律 的子孫、 米希大 的子孫、 哈沙 的子孫、
NEH|7|55|巴柯 的子孫、 西西拉 的子孫、 答瑪 的子孫、
NEH|7|56|尼細亞 的子孫、 哈提法 的子孫。
NEH|7|57|所羅門 僕人的後裔： 瑣太 的子孫、 瑣斐列 的子孫、 比路大 的子孫、
NEH|7|58|雅拉 的子孫、 達昆 的子孫、 吉德 的子孫、
NEH|7|59|示法提雅 的子孫、 哈替 的子孫、 玻黑列‧哈斯巴音 的子孫、 亞們 的子孫。
NEH|7|60|殿役和 所羅門 僕人的後裔共三百九十二名。
NEH|7|61|從 特‧米拉 、 特‧哈薩 、 基綠 、 亞頓 、 音麥 上來，不能證明他們的父系家族和後裔是否屬 以色列 的如下：
NEH|7|62|第萊雅 的子孫、 多比雅 的子孫、 尼哥大 的子孫，共六百四十二名。
NEH|7|63|祭司中， 哈巴雅 的子孫、 哈哥斯 的子孫、 巴西萊 的子孫， 巴西萊 因為娶了 基列 人 巴西萊 的女兒為妻，所以就以此為名。
NEH|7|64|這些人在族譜之中尋查自己的譜系，卻尋不著，因此算為不潔，不得作祭司。
NEH|7|65|省長對他們說，不可吃至聖的物，直到有會用烏陵和土明的祭司興起來。
NEH|7|66|全會眾共有四萬二千三百六十名。
NEH|7|67|此外，還有他們的僕婢七千三百三十七名，又有歌唱的男女二百四十五名。
NEH|7|68|他們有七百三十六匹馬，二百四十五匹騾子，
NEH|7|69|四百三十五匹駱駝，六千七百二十匹驢。
NEH|7|70|有些族長為工程捐助。省長捐入庫房中的有一千達利克 金子，五十個碗，五百三十件祭司的禮服。
NEH|7|71|有些族長捐入工程的庫房，有二萬達利克金子，二千二百彌那銀子。
NEH|7|72|其餘百姓所捐的有二萬達利克金子，二千彌那銀子，六十七件祭司的禮服。
NEH|7|73|於是祭司、 利未 人、門口的守衛、歌唱的、百姓中的一些人、殿役，並 以色列 眾人，都住在自己的城裏。 到了七月， 以色列 人住在自己的城裏。
NEH|8|1|那時，眾百姓如同一人聚集在 水門 前的廣場，請 以斯拉 文士將耶和華吩咐 以色列 的 摩西 的律法書帶來。
NEH|8|2|七月初一， 以斯拉 祭司將律法書帶到聽了能明白的男女會眾面前。
NEH|8|3|他在 水門 前的廣場，從清早到中午，在男女和能明白的人面前讀這律法書，眾百姓都側耳而聽。
NEH|8|4|以斯拉 文士站在為這事特製的木臺上。站在他旁邊的有 瑪他提雅 、 示瑪 、 亞奈雅 、 烏利亞 和 希勒家 ；站在他右邊的有 瑪西雅 ；站在他左邊的有 毗大雅 、 米沙利 、 瑪基雅 、 哈順 、 哈拔大拿 、 撒迦利亞 和 米書蘭 。
NEH|8|5|以斯拉 站在上面，在眾百姓眼前展開這書。他一展開，眾百姓都站起來。
NEH|8|6|以斯拉 稱頌耶和華至大的上帝，眾百姓都舉手應聲說：「阿們！阿們！」他們低頭，俯伏在地，敬拜耶和華。
NEH|8|7|耶書亞 、 巴尼 、 示利比 、 雅憫 、 亞谷 、 沙比太 、 荷第雅 、 瑪西雅 、 基利他 、 亞撒利雅 、 約撒拔 、 哈難 、 毗萊雅 和 利未 人使百姓明白律法；百姓都站在自己的地方。
NEH|8|8|他們清清楚楚地念上帝的律法書，講明意思，使百姓明白所念的。
NEH|8|9|尼希米 省長、 以斯拉 祭司文士，和教導百姓的 利未 人對眾百姓說：「今日是耶和華－你們上帝的聖日，不要悲哀，也不要哭泣。」這是因為眾百姓聽見律法書上的話都哭了。
NEH|8|10|尼希米 對他們說：「你們去吃肥美的，喝甘甜的，有不能預備的就分給他，因為今日是我們主的聖日。你們不要憂愁，因靠耶和華而得的喜樂是你們的力量。」
NEH|8|11|於是 利未 人叫眾百姓安靜，說：「安靜，因今日是聖日，不要憂愁。」
NEH|8|12|眾百姓去吃喝，也分給別人，都大大喜樂，因為他們明白所教導他們的話。
NEH|8|13|次日，眾百姓的族長、祭司和 利未 人都聚集到 以斯拉 文士那裏，要明白律法書上的話。
NEH|8|14|他們發現律法書上寫著，耶和華藉 摩西 吩咐 以色列 人要在七月的節期中住在棚裏，
NEH|8|15|並要在各城和 耶路撒冷 傳揚宣告說：「你們當出去，上山，把橄欖樹、野橄欖樹、番石榴樹、棕樹和各樣茂密樹的枝子取來，照著所寫的搭棚。」
NEH|8|16|於是百姓出去，取了樹枝來，各人在自己的房頂上、院子裏、上帝殿的院內、 水門 的廣場和 以法蓮門 的廣場搭棚。
NEH|8|17|從被擄之地歸回的全會眾就搭棚，住在棚裏。從 嫩 的兒子 約書亞 的時候直到這日， 以色列 人沒有這樣行。他們都大大喜樂。
NEH|8|18|從第一天直到末一天， 以斯拉 天天朗讀上帝的律法書。他們守節七日，第八日照例有嚴肅會。
NEH|9|1|這月二十四日， 以色列 人聚集禁食，他們披麻蒙灰。
NEH|9|2|以色列 的後裔與所有的外邦人分別出來，站著承認自己的罪和祖先的罪孽。
NEH|9|3|那日的四分之一，他們站在自己的地方念耶和華－他們上帝的律法書，又在那日的四分之一認罪，敬拜耶和華－他們的上帝。
NEH|9|4|耶書亞 、 巴尼 、 甲篾 、 示巴尼 、 布尼 、 示利比 、 巴尼 、 基拿尼 站在 利未 人的臺階上，大聲哀求耶和華－他們的上帝。
NEH|9|5|利未 人 耶書亞 、 甲篾 、 巴尼 、 哈沙尼 、 示利比 、 荷第雅 、 示巴尼 、 毗他希雅 說：「起來，稱頌耶和華－你們的上帝，永世無盡：『你榮耀之名是應當稱頌的，超乎一切稱頌和讚美。
NEH|9|6|「『你，惟獨你是耶和華！你造了天和天上的天，以及天上的萬象，地和地上的萬物，海和海中所有的；一切的生命全都是你賞賜的。天軍都敬拜你。
NEH|9|7|你是耶和華上帝，曾揀選 亞伯蘭 ，領他出 迦勒底 的 吾珥 ，給他改名叫 亞伯拉罕 。
NEH|9|8|你發現他在你面前心裏忠誠，就與他立約，要把 迦南 人、 赫 人、 亞摩利 人、 比利洗 人、 耶布斯 人、 革迦撒 人之地賜給他的後裔，並且你也實現了你的話，因為你是公義的。
NEH|9|9|「『你曾看見我們祖先在 埃及 所受的困苦，垂聽他們在 紅海 邊的哀求，
NEH|9|10|施行神蹟奇事在法老和他所有臣僕，以及他國中眾百姓身上，因為你知道他們向我們祖先行事狂傲。你也得了名聲，正如今日一樣。
NEH|9|11|你在我們祖先面前把海分開，使他們走過海中乾地，將追趕他們的人拋在深海，如石頭拋在大水中。
NEH|9|12|白晝你用雲柱引導他們，黑夜你用火柱照亮他們當行的路。
NEH|9|13|你降臨在 西奈山 ，從天上與他們說話，賜給他們正直的典章、真實的律法、美好的律例與誡命，
NEH|9|14|又使他們知道你的聖安息日，並藉你僕人 摩西 傳給他們誡命、律例、律法。
NEH|9|15|你從天上賜下糧食給他們充飢，使水從磐石流出給他們解渴。你吩咐他們進去，得你起誓應許要賜給他們的地。
NEH|9|16|「『但我們的祖先行事狂傲，硬著頸項不聽從你的誡命。
NEH|9|17|他們不肯順從，也不記念你在他們中間所行的奇事，竟硬著頸項，居心悖逆，自立領袖，要回 埃及 他們為奴之地 。但你是樂意饒恕人，有恩惠，有憐憫，不輕易發怒，有豐盛慈愛的上帝，並沒有丟棄他們。
NEH|9|18|他們雖然為自己鑄了一頭牛犢，說，這就是領你出 埃及 的神明，因而犯了褻瀆的大罪，
NEH|9|19|你還是有豐富的憐憫，不把他們丟棄在曠野。白晝，雲柱不離開他們，仍引導他們行路；黑夜，火柱仍照亮他們當行的路。
NEH|9|20|你賜下你良善的靈教導他們，沒有收回嗎哪不給他們吃，仍賜水給他們解渴。
NEH|9|21|在曠野四十年，你養育他們，他們一無所缺，衣服沒有穿破，腳也沒有腫。
NEH|9|22|你將列國和諸民族交給他們，把那些角落分給他們，他們就得了 西宏 之地，就是 希實本 王之地，和 巴珊 王 噩 之地。
NEH|9|23|你使他們的子孫多如天上的星，帶他們到你對他們祖先說要進去得為業之地。
NEH|9|24|這樣，這些子孫進去得了那地。你在他們面前制伏那地的居民 迦南 人，把 迦南 人和他們的君王，以及那地的民族，都交在他們手裏，讓他們任意處置。
NEH|9|25|他們得了堅固的城鎮、肥沃的土地，取了裝滿各樣美物的房屋、挖成的水井、葡萄園、橄欖園，以及許多果樹。他們就吃了，而且飽足，身體肥胖，因你的大恩活得快樂。
NEH|9|26|「『然而，他們不順從，竟背叛你，將你的律法丟在背後，又殺害那些勸他們回轉歸向你的眾先知，犯了褻瀆的大罪。
NEH|9|27|所以你將他們交在敵人的手中，敵人就折磨他們。他們遭難的時候哀求你，你就從天上垂聽，照你豐富的憐憫賜給他們拯救者，救他們脫離敵人的手。
NEH|9|28|但他們得享太平之後，又在你面前行惡，所以你丟棄他們，交在仇敵的手中，仇敵就轄制他們；然而他們轉回哀求你，你就從天上垂聽，屢次照你的憐憫拯救他們，
NEH|9|29|你警戒他們，要使他們歸順你的律法。他們卻行事狂傲，不聽從你的誡命，干犯你的典章，人若遵行就必因此存活。他們頑梗地扭轉肩頭，硬著頸項，不肯聽從。
NEH|9|30|但你多年寬容他們，又以你的靈藉眾先知勸戒他們，他們仍不側耳而聽，所以你將他們交在列邦民族的手中。
NEH|9|31|然而因你豐富的憐憫，你不全然滅絕他們，也不丟棄他們，因為你是有恩惠、有憐憫的上帝。
NEH|9|32|「『現在，我們的上帝啊，你是至大、至能、至可畏、守約施慈愛的上帝；我們的君王、官長、祭司、先知、祖先和你的眾百姓，從 亞述 諸王的時候直到今日所遭遇的一切苦難，求你不要看為小事。
NEH|9|33|在一切臨到我們的事上，你是公義的，因為你所行的是信實，我們所做的是邪惡。
NEH|9|34|我們的君王、官長、祭司、祖先都不遵守你的律法，不聽從你的誡命和你警戒他們的話。
NEH|9|35|他們在本國領受你大恩的時候，在你所賜給他們這廣大肥沃之地不事奉你，也不轉離他們的惡行。
NEH|9|36|看哪，我們今日成了奴僕！你賜給我們祖先享受土產和美物的地，看哪，我們在這地上竟作了奴僕！
NEH|9|37|這地許多的出產都歸了諸王，就是你因我們的罪派來轄制我們的。他們任意轄制我們的身體和牲畜，我們遭了大難。』」
NEH|9|38|因這一切，我們立確實的約，寫在冊上。我們的領袖、 利未 人和祭司都用了印。
NEH|10|1|用印的是 哈迦利亞 的兒子 尼希米 省長、 西底家 ；
NEH|10|2|還有 西萊雅 、 亞撒利雅 、 耶利米 、
NEH|10|3|巴施戶珥 、 亞瑪利雅 、 瑪基雅 、
NEH|10|4|哈突 、 示巴尼 、 瑪鹿 、
NEH|10|5|哈琳 、 米利末 、 俄巴底亞 、
NEH|10|6|但以理 、 近頓 、 巴錄 、
NEH|10|7|米書蘭 、 亞比雅 、 米雅民 、
NEH|10|8|瑪西亞 、 璧該 、 示瑪雅 等祭司；
NEH|10|9|又有 利未 人 亞散尼 的兒子 耶書亞 、 希拿達 的子孫 賓內 、 甲篾 ，
NEH|10|10|他們的弟兄 示巴尼 、 荷第雅 、 基利他 、 毗萊雅 、 哈難 、
NEH|10|11|米迦 、 利合 、 哈沙比雅 、
NEH|10|12|撒刻 、 示利比 、 示巴尼 、
NEH|10|13|荷第雅 、 巴尼 、 比尼努 ；
NEH|10|14|還有百姓中的領袖 巴錄 、 巴哈‧摩押 、 以攔 、 薩土 、 巴尼 、
NEH|10|15|布尼 、 押甲 、 比拜 、
NEH|10|16|亞多尼雅 、 比革瓦伊 、 亞丁 、
NEH|10|17|亞特 、 希西家 、 押朔 、
NEH|10|18|荷第雅 、 哈順 、 比賽 、
NEH|10|19|哈拉 、 亞拿突 、 尼拜 、
NEH|10|20|抹比押 、 米書蘭 、 希悉 、
NEH|10|21|米示薩別 、 撒督 、 押杜亞 、
NEH|10|22|毗拉提 、 哈難 、 亞奈雅 、
NEH|10|23|何細亞 、 哈拿尼雅 、 哈述 、
NEH|10|24|哈羅黑 、 毗利哈 、 朔百 、
NEH|10|25|利宏 、 哈沙拿 、 瑪西雅 、
NEH|10|26|亞希雅 、 哈難 、 亞難 、
NEH|10|27|瑪鹿 、 哈琳 、 巴拿 。
NEH|10|28|其餘的百姓、祭司、 利未 人、門口的守衛、歌唱的、殿役，所有與鄰邦民族分別出來、歸服上帝律法的，以及他們的妻子、兒女，凡有知識、能明白的，
NEH|10|29|都隨從他們貴族的弟兄發咒起誓，要遵行上帝藉他僕人 摩西 所賜的律法，謹守遵行耶和華－我們主的一切誡命、典章、律例。
NEH|10|30|我們不把我們的女兒嫁給這地的居民，也不為我們的兒子娶他們的女兒。
NEH|10|31|這地的民族若在安息日，或甚麼聖日，帶了貨物或糧食來賣，我們必不買。每逢第七年必不耕種，凡欠我們債的必不追討。
NEH|10|32|我們又為自己定例，每年各人捐獻三分之一舍客勒，作為我們上帝殿之用：
NEH|10|33|為供餅、常獻的素祭和燔祭，安息日、初一、節期所獻的祭和聖物， 以色列 的贖罪祭，以及我們上帝殿裏一切工作之用。
NEH|10|34|我們的祭司、 利未 人和百姓都抽籤，每年按父家定期將奉獻的木柴帶到我們上帝的殿裏，照著律法上所寫的，燒在耶和華－我們上帝的壇上。
NEH|10|35|每年我們又將地上初熟的土產和各樣樹上初熟的果子，都奉到耶和華的殿裏。
NEH|10|36|我們又照律法上所寫的，將我們頭胎的兒子和首生的牛羊都奉到我們上帝的殿，交給在上帝殿裏供職的祭司；
NEH|10|37|並將初熟麥子所磨的麵和舉祭、各樣樹上的果子、新酒與新油奉給祭司，收在我們上帝殿的庫房裏，又把我們土地所產的十分之一奉給 利未 人，因 利未 人在我們一切城鎮的土產中當取十分之一。
NEH|10|38|利未 人取十分之一的時候， 亞倫 的子孫中當有一個祭司與 利未 人同在。 利未 人也當從十分之一中取十分之一，奉到我們上帝的殿，收在庫房的倉裏。
NEH|10|39|因 以色列 人和 利未 人要把禮物，就是五穀、新酒和新油，帶到收存聖所器皿的倉裏，供職的祭司、門口的守衛、歌唱的都在那裏。我們絕不會不顧我們上帝的殿。
NEH|11|1|百姓的領袖住在 耶路撒冷 。其餘的百姓抽籤，每十人中選一人來住在聖城 耶路撒冷 ，另外九人住在別的城鎮。
NEH|11|2|凡甘心樂意住在 耶路撒冷 的，百姓都為他們祝福。
NEH|11|3|以色列 人、祭司、 利未 人、殿役和 所羅門 僕人的後裔都住在 猶大 的城鎮，各在自己城內的地業中。本省的領袖住在 耶路撒冷 的如下：
NEH|11|4|住在 耶路撒冷 的有一些 猶大 人和 便雅憫 人。 猶大 人中有 法勒斯 的子孫 亞他雅 ； 亞他雅 是 烏西雅 的兒子， 烏西雅 是 撒迦利雅 的兒子， 撒迦利雅 是 亞瑪利雅 的兒子， 亞瑪利雅 是 示法提雅 的兒子， 示法提雅 是 瑪勒列 的兒子；
NEH|11|5|又有 瑪西雅 ； 瑪西雅 是 巴錄 的兒子， 巴錄 是 谷‧何西 的兒子， 谷‧何西 是 哈賽雅 的兒子， 哈賽雅 是 亞大雅 的兒子， 亞大雅 是 約雅立 的兒子， 約雅立 是 撒迦利雅 的兒子， 撒迦利雅 是 示羅尼 的兒子；
NEH|11|6|住在 耶路撒冷 所有 法勒斯 的子孫共四百六十八名，都是勇士。
NEH|11|7|便雅憫 人中有 撒路 ； 撒路 是 米書蘭 的兒子， 米書蘭 是 約葉 的兒子， 約葉 是 毗大雅 的兒子， 毗大雅 是 哥賴雅 的兒子， 哥賴雅 是 瑪西雅 的兒子， 瑪西雅 是 以鐵 的兒子， 以鐵 是 耶篩亞 的兒子；
NEH|11|8|其次有 迦拜 、 撒來 ，共九百二十八名。
NEH|11|9|細基利 的兒子 約珥 是他們的長官； 哈西努亞 的兒子 猶大 是 耶路撒冷 的副長官。
NEH|11|10|祭司中有 約雅立 的兒子 耶大雅 ，又有 雅斤 ，
NEH|11|11|還有管理上帝殿的 西萊雅 ； 西萊雅 是 希勒家 的兒子， 希勒家 是 米書蘭 的兒子， 米書蘭 是 撒督 的兒子， 撒督 是 米拉約 的兒子， 米拉約 是 亞希突 的兒子；
NEH|11|12|還有他們的弟兄在殿裏供職的，共八百二十二名；又有 亞大雅 ； 亞大雅 是 耶羅罕 的兒子， 耶羅罕 是 毗拉利 的兒子， 毗拉利 是 暗洗 的兒子， 暗洗 是 撒迦利亞 的兒子， 撒迦利亞 是 巴施戶珥 的兒子， 巴施戶珥 是 瑪基雅 的兒子；
NEH|11|13|還有他的弟兄作族長的，共二百四十二名；又有 亞瑪帥 ； 亞瑪帥 是 亞薩列 的兒子， 亞薩列 是 亞哈賽 的兒子， 亞哈賽 是 米實利末 的兒子， 米實利末 是 音麥 的兒子；
NEH|11|14|還有他們的弟兄，大能的勇士共一百二十八名； 哈基多琳 的兒子 撒巴第業 是他們的長官。
NEH|11|15|利未 人中有 示瑪雅 ； 示瑪雅 是 哈述 的兒子， 哈述 是 押利甘 的兒子， 押利甘 是 哈沙比雅 的兒子， 哈沙比雅 是 布尼 的兒子；
NEH|11|16|又有 利未 人的族長 沙比太 和 約撒拔 管理上帝殿外面的事務；
NEH|11|17|祈禱的時候， 瑪他尼 是主禮，開始稱謝； 瑪他尼 是 米迦 的兒子， 米迦 是 撒底 的兒子， 撒底 是 亞薩 的兒子；又有 瑪他尼 弟兄中的 八布迦 為副；還有 押大 ； 押大 是 沙母亞 的兒子， 沙母亞 是 加拉 的兒子， 加拉 是 耶杜頓 的兒子；
NEH|11|18|在聖城所有的 利未 人共二百八十四名。
NEH|11|19|門口的守衛是 亞谷 和 達們 ，以及他們的弟兄，看守各門，共一百七十二名。
NEH|11|20|其餘的 以色列 人、祭司、 利未 人都住在 猶大 一切的城鎮，各在自己的地業中。
NEH|11|21|殿役卻住在 俄斐勒 ； 西哈 和 基斯帕 管理他們。
NEH|11|22|在 耶路撒冷 ， 利未 人的長官，管理上帝殿事務的是歌唱者 亞薩 的子孫 烏西 ； 烏西 是 巴尼 的兒子， 巴尼 是 哈沙比雅 的兒子， 哈沙比雅 是 瑪他尼 的兒子， 瑪他尼 是 米迦 的兒子。
NEH|11|23|王為歌唱者下命令，確定他們每日當辦的事 。
NEH|11|24|猶大 的兒子 謝拉 的子孫， 米示薩別 的兒子 毗他希雅 輔助王辦理百姓一切的事。
NEH|11|25|至於村莊和所屬的田地，有 猶大 人住在 基列‧亞巴 和所屬的鄉鎮 、 底本 和所屬的鄉鎮、 葉甲薛 和所屬的村莊、
NEH|11|26|耶書亞 、 摩拉大 、 伯‧帕列 、
NEH|11|27|哈薩‧書亞 、 別是巴 和所屬的鄉鎮、
NEH|11|28|洗革拉 、 米哥拿 和所屬的鄉鎮、
NEH|11|29|隱‧臨門 、 瑣拉 、 耶末 、
NEH|11|30|撒挪亞 、 亞杜蘭 和屬它們的村莊、 拉吉 和所屬的田地、 亞西加 和所屬的鄉鎮；他們所住的地方是從 別是巴 直到 欣嫩谷 。
NEH|11|31|便雅憫 人從 迦巴 起，住在 密抹 、 亞雅 、 伯特利 和所屬的鄉鎮、
NEH|11|32|亞拿突 、 挪伯 、 亞難雅 、
NEH|11|33|夏瑣 、 拉瑪 、 基他音 、
NEH|11|34|哈第 、 洗編 、 尼八拉 、
NEH|11|35|羅德 、 阿挪 、 革‧夏納欣 。
NEH|11|36|在 猶大 地區的 利未 人中，有些已歸屬 便雅憫 。
NEH|12|1|這些是同 撒拉鐵 的兒子 所羅巴伯 以及 耶書亞 一起上來的祭司和 利未 人： 西萊雅 、 耶利米 、 以斯拉 、
NEH|12|2|亞瑪利雅 、 瑪鹿 、 哈突 、
NEH|12|3|示迦尼 、 利宏 、 米利末 、
NEH|12|4|易多 、 近頓 、 亞比雅 、
NEH|12|5|米雅民 、 瑪底雅 、 璧迦 、
NEH|12|6|示瑪雅 、 約雅立 、 耶大雅 、
NEH|12|7|撒路 、 亞木 、 希勒家 、 耶大雅 ；這些人在 耶書亞 的時代作祭司和他們弟兄的領袖。
NEH|12|8|利未 人有 耶書亞 、 賓內 、 甲篾 、 示利比 、 猶大 、 瑪他尼 ； 瑪他尼 和他的弟兄負責讚美詩歌。
NEH|12|9|他們的弟兄 八布迦 和 烏尼 按照班次站在他們的對面。
NEH|12|10|耶書亞 生 約雅金 ， 約雅金 生 以利亞實 ， 以利亞實 生 耶何耶大 ，
NEH|12|11|耶何耶大 生 約拿單 ， 約拿單 生 押杜亞 。
NEH|12|12|在 約雅金 的時代，祭司作族長的， 西萊雅 族有 米拉雅 ， 耶利米 族有 哈拿尼雅 ，
NEH|12|13|以斯拉 族有 米書蘭 ， 亞瑪利雅 族有 約哈難 ，
NEH|12|14|米利古 族有 約拿單 ， 示巴尼 族有 約瑟 ，
NEH|12|15|哈琳 族有 押拿 ， 米拉約 族有 希勒愷 ，
NEH|12|16|易多 族有 撒迦利亞 ， 近頓 族有 米書蘭 ，
NEH|12|17|亞比雅 族有 細基利 ， 米拿民 族， 摩亞底 族有 毗勒太 ，
NEH|12|18|璧迦 族有 沙母亞 ， 示瑪雅 族有 約拿單 ，
NEH|12|19|約雅立 族有 瑪特乃 ， 耶大雅 族有 烏西 ，
NEH|12|20|撒來 族有 加萊 ， 亞木 族有 希伯 ，
NEH|12|21|希勒家 族有 哈沙比雅 ， 耶大雅 族有 拿坦業 。
NEH|12|22|在 以利亞實 、 耶何耶大 、 約哈難 、 押杜亞 的時代， 利未 人的族長都記在冊上，祭司也一樣，直到 波斯 王 大流士 在位的時候。
NEH|12|23|利未 人作族長的記在史籍上，一直記到 以利亞實 的兒子 約哈難 的時代。
NEH|12|24|利未 人的族長是 哈沙比雅 、 示利比 、 甲篾 的兒子 耶書亞 ，他們的弟兄站在他們的對面，照神人 大衛 的命令按著班次讚美稱謝。
NEH|12|25|瑪他尼 、 八布迦 、 俄巴底亞 、 米書蘭 、 達們 、 亞谷 是門口的守衛，在庫房的門口站崗。
NEH|12|26|這些人都在 約撒達 的孫子， 耶書亞 的兒子 約雅金 和 尼希米 省長，以及 以斯拉 祭司文士的時代供職。
NEH|12|27|為 耶路撒冷 城牆行奉獻禮的時候，眾人把各處的 利未 人召到 耶路撒冷 ，要以稱謝、歌唱、敲鈸、鼓瑟、彈琴，喜樂地行奉獻禮。
NEH|12|28|歌唱的人從 耶路撒冷 的周圍聚集，從 尼陀法 人的村莊、
NEH|12|29|伯‧吉甲 ，以及 迦巴 和 亞斯瑪弗 的田地而來；因為歌唱的人在 耶路撒冷 四圍為自己建立了村莊。
NEH|12|30|祭司和 利未 人就潔淨自己，也潔淨百姓，以及城門和城牆。
NEH|12|31|我帶 猶大 的領袖上城牆，把稱謝的人分為兩大隊，在城牆上往右邊的 糞廠門 行進，
NEH|12|32|在他們後面行進的有 何沙雅 與 猶大 一半的領袖，
NEH|12|33|又有 亞撒利雅 、 以斯拉 、 米書蘭 、
NEH|12|34|猶大 、 便雅憫 、 示瑪雅 、 耶利米 。
NEH|12|35|還有祭司的子孫，吹號的有 撒迦利亞 ； 撒迦利亞 是 約拿單 的兒子， 約拿單 是 示瑪雅 的兒子， 示瑪雅 是 瑪他尼 的兒子， 瑪他尼 是 米該亞 的兒子， 米該亞 是 撒刻 的兒子， 撒刻 是 亞薩 的兒子；
NEH|12|36|又有 撒迦利亞 的弟兄 示瑪雅 、 亞撒利 、 米拉萊 、 基拉萊 、 瑪艾 、 拿坦業 、 猶大 、 哈拿尼 ，各拿著神人 大衛 的樂器，由 以斯拉 文士在前面引領。
NEH|12|37|他們經過 泉門 往前，登 大衛城 的臺階，上城牆的斜坡，從 大衛 宮殿之上，直到朝東的 水門 。
NEH|12|38|第二隊稱謝的人要往反方向而行。我和一半的百姓在城牆上跟隨他們，從 爐樓 之上，直到 寬牆 ；
NEH|12|39|又過了 以法蓮門 、 古門 、 魚門 、 哈楠業樓 、 哈米亞樓 ，直到 羊門 ，就在 護衛門 站住。
NEH|12|40|於是，這兩隊稱謝的人連同我和一半跟隨我的官長，站在上帝的殿裏。
NEH|12|41|還有 以利亞金 、 瑪西雅 、 米拿民 、 米該亞 、 以利約乃 、 撒迦利亞 、 哈楠尼亞 等吹號的祭司；
NEH|12|42|又有 瑪西雅 、 示瑪雅 、 以利亞撒 、 烏西 、 約哈難 、 瑪基雅 、 以攔 和 以謝 。歌唱的大聲唱歌，有 伊斯拉希雅 作指揮。
NEH|12|43|那日，眾人獻上豐盛的祭物，並且歡樂，因為上帝使他們大大歡樂，連婦女帶孩童也都歡樂，甚至從遠處都可聽到 耶路撒冷 的歡聲。
NEH|12|44|當日，有些人受派管理庫房，把舉祭、初熟之物，和所取的十一奉獻，按各城的田地，照律法所定，歸給祭司和 利未 人的份，都收在庫房裏。 猶大 人因祭司和 利未 人供職就歡樂。
NEH|12|45|祭司和 利未 人遵守上帝所吩咐的，守潔淨禮。歌唱的和門口的守衛照著 大衛 和他兒子 所羅門 的命令也如此行。
NEH|12|46|古時，在 大衛 和 亞薩 的日子，有歌唱者的指揮，也有讚美稱謝上帝的詩歌。
NEH|12|47|在 所羅巴伯 和 尼希米 的時代， 以色列 眾人把歌唱者和門口的守衛每日當得的份供給他們，又把給 利未 人的分別出來； 利未 人又把給 亞倫 子孫的分別出來。
NEH|13|1|在那日，百姓聽到人朗讀 摩西 的律法書，發現書上寫著， 亞捫 人和 摩押 人永不可入上帝的會；
NEH|13|2|因為他們沒有拿食物和水來迎接 以色列 人，卻雇了 巴蘭 詛咒他們，但我們的上帝使那詛咒變為祝福。
NEH|13|3|以色列 人聽見這律法，就與所有不同族群的人分別出來。
NEH|13|4|在這之前，與 多比雅 結親的 以利亞實 祭司，受派管理我們上帝殿中的庫房，
NEH|13|5|為 多比雅 預備了一間大屋子，就是從前收存素祭、乳香、器皿，和照例供給 利未 人、歌唱者、門口守衛的五穀、新酒和新油的十分之一，以及歸祭司之舉祭的屋子。
NEH|13|6|當這一切事發生的時候，我不在 耶路撒冷 ，因為 巴比倫 王 亞達薛西 三十二年，我回到王那裏。過了多日，我又向王告假。
NEH|13|7|我來到 耶路撒冷 ，才知道 以利亞實 為 多比雅 所做、在上帝殿的院內為他預備屋子的那件惡事。
NEH|13|8|我非常憤怒，就把 多比雅 的一切家具都從屋子裏拋出去。
NEH|13|9|我又吩咐人潔淨這屋子，然後將上帝殿的器皿、素祭和乳香搬回那裏。
NEH|13|10|我發現 利未 人當得的份無人供給他們，甚至供職的 利未 人與歌唱的都各奔回自己的田地去了。
NEH|13|11|我就斥責官長說：「你們為何不顧上帝的殿呢？」於是我召集 利未 人，使他們在自己的崗位上供職。
NEH|13|12|猶大 眾人就把五穀、新酒和新油的十分之一送入庫房。
NEH|13|13|我派 示利米雅 祭司、 撒督 文士和 利未 人 毗大雅 作司庫管理庫房，副手是 哈難 ； 哈難 是 撒刻 的兒子， 撒刻 是 瑪他尼 的兒子；這些人都是忠實的，他們的職務是分派他們弟兄所當得的份。
NEH|13|14|我的上帝啊，求你因這事記念我，不要塗去我為上帝的殿與其中的禮儀所獻的忠心。
NEH|13|15|那些日子，我在 猶大 見有人在安息日踹醡酒池，搬運禾捆馱在驢上，又把酒、葡萄、無花果和各樣的擔子在安息日扛入 耶路撒冷 ，我就在他們賣食物的那日警戒他們。
NEH|13|16|有一些住在城裏的 推羅 人也把魚和各樣貨物運進來，甚至在 耶路撒冷 ，在安息日賣給 猶大 人。
NEH|13|17|我就斥責 猶大 的貴族，對他們說：「你們怎麼會做這惡事干犯安息日呢！
NEH|13|18|你們祖先豈不是這樣做，以致我們的上帝使一切災禍臨到我們和這城嗎？你們竟干犯安息日，使憤怒越發臨到 以色列 ！」
NEH|13|19|安息日前一日黃昏的時候，我吩咐人把 耶路撒冷 城門鎖上；我又吩咐，不過安息日不准開門。我也派幾個僕人在城門口站崗，免得有人在安息日挑擔子進城。
NEH|13|20|於是商人和販賣各樣貨物的人，有一兩次在 耶路撒冷 城外過夜。
NEH|13|21|我警告他們說：「你們為何在城牆前過夜呢？若再這樣，我必下手辦你們。」從此以後，他們在安息日就不再來了。
NEH|13|22|我吩咐 利未 人潔淨自己來守城門，使安息日分別為聖。我的上帝啊，求你因這事記念我，照你豐盛的慈愛憐憫我。
NEH|13|23|那些日子，我又看見 猶太 人娶了 亞實突 、 亞捫 和 摩押 的女子為妻。
NEH|13|24|他們的兒女，一半說 亞實突 話，或其他種族的方言，不會說 猶大 話。
NEH|13|25|我就斥責他們，詛咒他們，打了他們幾個人，拔下他們的鬍鬚，叫他們指著上帝起誓：「你們不可把自己的女兒嫁給外邦人的兒子，也不可為自己和兒子娶他們的女兒。
NEH|13|26|以色列 王 所羅門 不也在這樣的事上犯罪嗎？在許多國家中並沒有一位王像他，蒙他上帝喜愛，上帝立他作王治理全 以色列 。然而，連他也被外邦女子引誘犯罪。
NEH|13|27|我們豈能聽憑你們行這一切大惡，娶外邦女子干犯我們的上帝呢？」
NEH|13|28|以利亞實 大祭司的孫子， 耶何耶大 的一個兒子是 和倫 人 參巴拉 的女婿，我就把他從我這裏趕出去。
NEH|13|29|我的上帝啊，求你記得他們的罪，因為他們玷污了祭司的職分，違背祭司和 利未 人的約。
NEH|13|30|這樣，我潔淨他們，使他們脫離屬外邦人的一切；我又分派祭司和 利未 人的班次，使他們各盡其職，
NEH|13|31|按定期奉獻木柴和初熟的土產。我的上帝啊，求你記念我，施恩於我。
ESTH|1|1|這事發生在 亞哈隨魯 的時代， 亞哈隨魯 從 印度 直到 古實 統治一百二十七個省，
ESTH|1|2|就是 亞哈隨魯 王在 書珊 城堡中坐國度王位的那些日子。
ESTH|1|3|他在位第三年，為所有官員和臣僕擺設宴席，有 波斯 和 瑪代 的權貴，各省的貴族與領袖在他面前。
ESTH|1|4|他把他榮耀國度的豐富和他偉大威嚴的尊貴給他們看了許多日子，共一百八十天。
ESTH|1|5|這些日子滿了，王又為所有住 書珊 城堡的百姓，無論大小，在御花園的院子裏擺設宴席七日。
ESTH|1|6|院子裏有白色棉和藍色線，用細麻繩、紫色繩繫在白玉石柱的銀環上，又有金銀的床榻擺在紅、白、黃、黑大理石鑲嵌的地上。
ESTH|1|7|用金器皿盛酒，有很多不同的器皿，照王的厚意提供豐富的御酒。
ESTH|1|8|飲酒有規定，不准勉強人 ，因為王吩咐宮裏所有的臣宰，讓人各隨己意。
ESTH|1|9|瓦實提 王后在 亞哈隨魯 王的宮內也為婦女擺設宴席。
ESTH|1|10|第七日， 亞哈隨魯 王飲酒，心中快樂，就吩咐在他面前侍立的七個太監 米戶幔 、 比斯他 、 哈波拿 、 比革他 、 亞拔他 、 西達 、 甲迦 ，
ESTH|1|11|請 瓦實提 王后頭戴王后的冠冕到王面前，讓各民族和官員觀看她的美貌，因為她容貌美麗。
ESTH|1|12|瓦實提 王后卻不肯遵照太監所傳的王命前來，所以王非常憤怒，怒火中燒。
ESTH|1|13|按王的常規，辦事必先詢問知例明法的人。那時，王詢問通達時務的智慧人，
ESTH|1|14|就是在王左右常見王面、在國中坐高位的 波斯 和 瑪代 的七個大臣， 甲示拿 、 示達 、 押瑪他 、 他施斯 、 米力 、 瑪西拿 、 米慕干 ：
ESTH|1|15|「 瓦實提 王后不遵照太監所傳的王命，照例應當怎樣辦理呢？」
ESTH|1|16|米慕干 在王和眾官長面前回答說：「 瓦實提 王后這事，不但得罪王，並且有害於 亞哈隨魯 王各省的臣民。
ESTH|1|17|因為王后這事必傳到眾婦人那裏，她們就會藐視自己的丈夫，說：『 亞哈隨魯 王吩咐 瓦實提 王后到王面前，她卻不來。』
ESTH|1|18|今日 波斯 和 瑪代 的眾夫人聽見王后這事，必向王所有的官長照樣說，如此必造成無數的藐視和憤怒。
ESTH|1|19|王若以為好，請降諭旨，寫在 波斯 和 瑪代 人的條例中，永不更改，不准 瓦實提 再到 亞哈隨魯 王面前，把她王后的位分賜給比她更好的妃子。
ESTH|1|20|王的諭旨一傳遍全國，國土縱然遼闊，凡作妻子的，無論丈夫是尊貴或卑賤，都必尊敬他。」
ESTH|1|21|王和眾官長都以這話為美，王就照 米慕干 的建議去做。
ESTH|1|22|王下詔書，用各省的文字、各族的語言通知各省，使凡作丈夫的在家中作主，各說本地的語言 。
ESTH|2|1|這些事以後， 亞哈隨魯 王的憤怒平息，就想起 瓦實提 和她所做的，以及自己怎樣降旨辦她。
ESTH|2|2|於是王的侍臣對王說：「請派人為王尋找美貌的少女；
ESTH|2|3|請王派官員在國中各省招聚所有美貌的少女到 書珊 城堡的女院，交給王所派掌管女子的太監 希該 ，給她們香膏塗抹。
ESTH|2|4|王眼中看為好的女子可以立為王后，代替 瓦實提 。」王以這話為美，就照樣做。
ESTH|2|5|書珊 城堡中有一個 猶太 人名叫 末底改 ，是 便雅憫 人 基士 的曾孫， 示每 的孫子， 睚珥 的兒子。
ESTH|2|6|從前 巴比倫 王 尼布甲尼撒 把 猶大 王 耶哥尼雅 和百姓從 耶路撒冷 擄來， 末底改 也在被擄的人當中。
ESTH|2|7|末底改 撫養他叔叔的女兒 哈大沙 ，就是 以斯帖 ，因為她沒有父母。這女子容貌美麗；她父母死了， 末底改 收她為自己的女兒。
ESTH|2|8|王的諭旨和敕令傳出之後，許多女子被招聚到 書珊 城堡，交給掌管女子的 希該 ； 以斯帖 也被送入王宮，交給 希該 。
ESTH|2|9|希該 眼中寵愛 以斯帖 ，就恩待她，急忙給她塗抹的香膏和當得的份，又從王宮裏挑選七個宮女來服事她，使她和她的宮女搬入女院上好的房屋。
ESTH|2|10|以斯帖 未曾將自己的籍貫宗族告訴人，因為 末底改 囑咐她不可叫人知道。
ESTH|2|11|末底改 天天在女院前徘徊，要知道 以斯帖 是否平安，過得如何。
ESTH|2|12|眾女子照例先塗抹身體十二個月：六個月用沒藥油，六個月用香料和塗抹的香膏。滿了日期，每個女子挨次進去朝見 亞哈隨魯 王。
ESTH|2|13|女子進去朝見王是這樣：從女院到王宮的時候，凡她所要的都必給她帶進去。
ESTH|2|14|晚上她進去，次日回到另一個女院，交給掌管妃嬪的太監 沙甲 。除非王喜愛她，再提名召她，她就不再進去見王。
ESTH|2|15|末底改 的叔叔 亞比孩 的女兒，就是 末底改 收為自己女兒的 以斯帖 ，按次序要進去朝見王的時候，除了掌管女子的太監 希該 所分派給她的，她別無所求。凡看見 以斯帖 的都喜歡她。
ESTH|2|16|亞哈隨魯 王第七年十月，就是提別月， 以斯帖 被引入宮中朝見王。
ESTH|2|17|王愛 以斯帖 過於眾女子，她在王面前蒙寵愛勝過眾少女。王把王后的冠冕戴在她頭上，立她為王后，代替 瓦實提 。
ESTH|2|18|王為所有的官長和臣僕擺設大宴席，稱為 以斯帖 的宴席，又豁免各省的租稅，並照王的厚意大頒賞賜。
ESTH|2|19|第二次招聚少女的時候， 末底改 坐在朝門。
ESTH|2|20|以斯帖 遵照 末底改 所囑咐的，沒有將籍貫宗族告訴人； 以斯帖 照 末底改 的吩咐去做，正如受他撫養的時候一樣。
ESTH|2|21|那時候， 末底改 坐在朝門，王有兩個守門的太監， 辟探 和 提列 ，惱恨 亞哈隨魯 王，想要下手害他。
ESTH|2|22|末底改 知道了這件事，就告訴 以斯帖 王后。 以斯帖 以 末底改 的名向王報告。
ESTH|2|23|這事經過查究後發現是真的，二人就被掛在木頭上。這事在王面前記錄在史籍上。
ESTH|3|1|這些事以後， 亞哈隨魯 王使 亞甲 人 哈米大他 的兒子 哈曼 尊大，提升了他，叫他的爵位超過所有與他同朝的官長。
ESTH|3|2|在朝門，王所有的臣僕都跪拜 哈曼 ，因為王如此吩咐，但 末底改 不跪不拜。
ESTH|3|3|在朝門，王的臣僕對 末底改 說：「你為何違背王的命令呢？」
ESTH|3|4|他們天天勸他，他還是不聽，他們就告訴 哈曼 ，要看 末底改 的事是否站得住，因他已經告訴他們自己是 猶太 人。
ESTH|3|5|哈曼 見 末底改 不跪不拜，就非常憤怒。
ESTH|3|6|有人把 末底改 的宗族告訴 哈曼 。 哈曼 看下手只害 末底改 一人是小事，還圖謀要滅絕 亞哈隨魯 王全國所有的 猶太 人，就是 末底改 的宗族。
ESTH|3|7|亞哈隨魯 王十二年正月，就是尼散月，人在 哈曼 面前抽普珥，普珥即籤，要定何月何日；抽到了十二月，就是亞達月。
ESTH|3|8|哈曼 對 亞哈隨魯 王說：「有一民族散居在王國各省的民族中，與眾不同；他們的律例與萬民的律例不同，也不守王的律例，所以容留他們對王無益。
ESTH|3|9|王若以為好，請下諭旨滅絕他們，我就捐一萬他連得銀子交給管財政的人，納入王的府庫。」
ESTH|3|10|於是王從自己手上摘下戒指給 猶太 人的仇敵， 亞甲 人 哈米大他 的兒子 哈曼 。
ESTH|3|11|王對 哈曼 說：「這銀子賜給你，這民族也交給你，可以照你眼中看為好的待他們。」
ESTH|3|12|正月十三日，王的一些書記受召而來，照著 哈曼 一切所吩咐的，用各省的文字、各族的語言，奉 亞哈隨魯 王的名寫諭旨，又用王的戒指蓋印，傳給王的總督、各省的省長，以及各族的領袖。
ESTH|3|13|詔書由信差傳到王的各省，限令一日之內，就是在十二月，亞達月十三日，把所有的 猶太 人，無論老少婦女孩子，全然剪除，殺戮滅絕，並搶奪他們的財產。
ESTH|3|14|這諭旨的抄本以敕令的方式在各省頒佈，通知各族，預備等候那日。
ESTH|3|15|信差奉王的命令急忙起行，敕令傳遍了 書珊 城堡。王同 哈曼 坐下飲酒， 書珊 城堡卻陷入慌亂中。
ESTH|4|1|末底改 知道所發生的這一切事，就撕裂衣服，披麻蒙灰，在城中行走，痛哭哀號。
ESTH|4|2|他到了朝門前就停住腳步，因為穿麻衣的不可進朝門。
ESTH|4|3|王的諭旨和敕令所到的各省各處， 猶太 人都極其悲哀，禁食哭泣哀號，許多人躺在麻布和爐灰中。
ESTH|4|4|以斯帖 王后的宮女和太監來把這事告訴 以斯帖 ，她非常憂愁，就送衣服給 末底改 穿，要他脫下身上的麻衣，他卻不肯接受。
ESTH|4|5|以斯帖 把王所派伺候她的一個太監 哈他革 召來，吩咐他去見 末底改 ，要知道到底發生了甚麼事，為何如此。
ESTH|4|6|於是 哈他革 出來，到朝門前的廣場見 末底改 。
ESTH|4|7|末底改 把自己遭遇的一切，以及 哈曼 為滅絕 猶太 人答應捐入王庫的銀數都告訴了他；
ESTH|4|8|又把那傳遍 書珊 、要滅絕 猶太 人的諭旨抄本交給 哈他革 ，要他給 以斯帖 看，並向她說明，囑咐她去晉見王，向王懇求，為本族的人在王面前請命。
ESTH|4|9|哈他革 回來，把 末底改 的話告訴 以斯帖 。
ESTH|4|10|以斯帖 吩咐 哈他革 去見 末底改 ，說：
ESTH|4|11|「王所有的臣僕和各省的百姓都知道有一個定例，若未奉召見，擅入內院見王的，無論男女必被處死；除非王向他伸出金杖，不得存活。但我沒有被召進去見王已經有三十天了。」
ESTH|4|12|他們把 以斯帖 的話告訴 末底改 。
ESTH|4|13|末底改 託人回覆 以斯帖 說：「你不要自己以為在王宮裏強過任何 猶太 人，得以倖免。
ESTH|4|14|此時你若閉口不言， 猶太 人必從別處得解脫，蒙拯救；你和你父家必致滅亡。焉知你得了王后的位分不是為現今的機會嗎？」
ESTH|4|15|以斯帖 吩咐人回覆 末底改 說：
ESTH|4|16|「你當去召集 書珊 所有的 猶太 人，為我禁食三晝三夜，不吃不喝；我和我的宮女也要這樣禁食。然後我違例去晉見王，我若死就死吧！」
ESTH|4|17|於是 末底改 照 以斯帖 一切所吩咐的去做。
ESTH|5|1|第三日， 以斯帖 穿上朝服，站立在王宮的內院，對著王宮。王在殿裏坐在寶座上，對著殿的門。
ESTH|5|2|王見 以斯帖 王后站在院內，她在王的眼中得恩寵，王向她伸出手中的金杖。 以斯帖 往前去摸杖頭。
ESTH|5|3|王對她說：「 以斯帖 王后啊，你要甚麼？無論你求甚麼，就是國的一半也必賜給你。」
ESTH|5|4|以斯帖 說：「王若以為好，請王帶著 哈曼 今日赴我為王預備的宴席。」
ESTH|5|5|王說：「叫 哈曼 速速照 以斯帖 的話去做。」於是王帶著 哈曼 赴 以斯帖 所預備的宴席。
ESTH|5|6|在宴席喝酒的時候，王又對 以斯帖 說：「你要甚麼，必賜給你；無論你求甚麼，就是國的一半也必給你。」
ESTH|5|7|以斯帖 回答說：「我所要的、我所求的，嗯......。
ESTH|5|8|我若在王眼前蒙恩，王若願意賜我所要的，准我所求的，就請王和 哈曼 再赴我為你們預備的宴席。明日我必照王的話去做。」
ESTH|5|9|那日 哈曼 心中快樂，歡歡喜喜地出來。但是當他看見 末底改 在朝門不站起來，也不因他動一下，就滿心惱怒 末底改 。
ESTH|5|10|哈曼 忍著氣回家，叫人請他的一些朋友和他妻子 細利斯 來。
ESTH|5|11|哈曼 將他的榮華富貴、眾多的兒女，和王使他尊大、提升他高過官長和臣僕的事，都述說給他們聽。
ESTH|5|12|哈曼 又說：「 以斯帖 王后預備宴席，除了我之外不許別人隨王赴席。明日王后又請我隨王赴席。
ESTH|5|13|只是每當我看見 猶太 人 末底改 坐在朝門，這一切對我就都毫無意義了。」
ESTH|5|14|他的妻子 細利斯 和他所有的朋友對他說：「叫人做一個五十肘高的木架，早晨求王把 末底改 掛在其上，然後你可以歡歡喜喜隨王赴席。」 哈曼 認為這話很好，就叫人做了木架。
ESTH|6|1|那夜王睡不著覺，吩咐人取歷史書，就是史籍，念給他聽，
ESTH|6|2|發現書上寫著：王有兩個守門的太監 辟探 和 提列 ，想要下手害 亞哈隨魯 王， 末底改 告發了這件事。
ESTH|6|3|王說：「 末底改 做了這事，有沒有賜給他甚麼尊榮或高位呢？」伺候王的臣僕說：「沒有賜給他甚麼。」
ESTH|6|4|王說：「誰在院子裏？」那時 哈曼 正進入王宮的外院，要請王把 末底改 掛在他所預備的木架上。
ESTH|6|5|王的臣僕對他說：「看哪， 哈曼 站在院子裏。」王說：「叫他進來。」
ESTH|6|6|哈曼 就進去。王對他說：「王所喜愛要賜尊榮的人，當如何待他呢？」 哈曼 心裏說：「王所喜愛要賜尊榮的人，除了我，還有誰呢？」
ESTH|6|7|哈曼 就對王說：「王所喜愛要賜尊榮的人，
ESTH|6|8|當把王所穿的王袍拿來，牽了戴冠的御馬，
ESTH|6|9|把王袍和御馬都交給王一個極尊貴的大臣，吩咐人把王袍給王所喜愛要賜尊榮的人穿上，領他騎著御馬走遍城裏的廣場，在他面前宣告：『王所喜愛要賜尊榮的人，就是這樣待他。』」
ESTH|6|10|王對 哈曼 說：「你速速把這王袍和御馬，照你所說的，向坐在朝門的 猶太 人 末底改 去做。凡你所說的，一樣都不可缺。」
ESTH|6|11|於是 哈曼 把王袍給 末底改 穿上，領他騎著御馬走遍城裏的廣場，在他面前宣告：「王所喜愛要賜尊榮的人，就是這樣待他。」
ESTH|6|12|末底改 仍回到朝門， 哈曼 卻憂憂悶悶地蒙著頭，急忙回家去了。
ESTH|6|13|哈曼 把所遭遇的一切都說給他妻子 細利斯 和他所有的朋友聽。他的智囊團和他的妻子 細利斯 對他說：「你在 末底改 面前開始敗落；他既是 猶太 人，你必不能勝過他，終必在他面前敗落。」
ESTH|6|14|他們正跟 哈曼 說話的時候，王的幾位太監來了，催 哈曼 快去赴 以斯帖 所預備的宴席。
ESTH|7|1|王帶著 哈曼 來赴 以斯帖 王后的宴席。
ESTH|7|2|第二天在宴席喝酒的時候，王又對 以斯帖 說：「 以斯帖 王后啊，你要甚麼，必賜給你；無論你求甚麼，就是國的一半也必給你。」
ESTH|7|3|以斯帖 王后回答說：「王啊，我若在你眼前蒙恩，王若以為好，我所要的，是王把我的性命賜給我；我所求的，是求我的本族。
ESTH|7|4|因為我和我的本族被出賣了，要被剪除，殺戮，滅絕。我們若被賣為奴為婢，我就閉口不言；但我們的痛苦比起王的損失，算不得甚麼 。」
ESTH|7|5|亞哈隨魯 王問 以斯帖 王后說：「擅敢起意如此行的是誰？這人在哪裏呢？」
ESTH|7|6|以斯帖 說：「仇人敵人就是這惡人 哈曼 ！」 哈曼 在王和王后面前非常驚惶。
ESTH|7|7|王大怒，起來離開酒席往御花園去了。 哈曼 見王定意要加罪於他，就留下來求 以斯帖 王后救他的命。
ESTH|7|8|王從御花園回到酒席廳，見 哈曼 伏在 以斯帖 所靠的榻上；王說：「他竟敢在宮內、在我面前凌辱王后嗎？」這話一出王口， 哈曼 的臉就被蒙住了。
ESTH|7|9|有一個伺候王名叫 哈波拿 的太監說：「看哪， 哈曼 還為那報告給王、救王有功的 末底改 做了一個五十肘高的木架，現今立在 哈曼 的家裏。」王說：「把 哈曼 掛在木架上。」
ESTH|7|10|於是 哈曼 被掛在他為 末底改 所預備的木架上；王的憤怒才平息了。
ESTH|8|1|那日， 亞哈隨魯 王把 猶太 人的仇敵 哈曼 的家產賜給 以斯帖 王后。 末底改 也來到王面前，因為 以斯帖 已經告訴王， 末底改 跟她是甚麼關係。
ESTH|8|2|王摘下自己的戒指，就是從 哈曼 取回的，給了 末底改 。 以斯帖 派 末底改 管理 哈曼 的家產。
ESTH|8|3|以斯帖 又在王面前求情，俯伏在他腳前，流淚哀求他阻止 亞甲 人 哈曼 害 猶太 人的惡謀。
ESTH|8|4|王向 以斯帖 伸出金杖， 以斯帖 就起來，站在王面前，
ESTH|8|5|說：「王若以為好，我若在王面前蒙恩，王若認為合宜，我若在王眼前得喜悅，請王下諭旨，廢除 亞甲 人 哈米大他 的兒子 哈曼 設謀，要殺滅王各省的 猶太 人所頒的詔書。
ESTH|8|6|我何忍見我本族的人受害？何忍見我同宗的人被滅呢？」
ESTH|8|7|亞哈隨魯 王對 以斯帖 王后和 猶太 人 末底改 說：「因為 哈曼 要下手害 猶太 人，看哪，我已把他的家產賜給 以斯帖 ，也把 哈曼 掛在木架上了。
ESTH|8|8|你們可以照你們看為好的，奉王的名寫諭旨給 猶太 人，用王的戒指蓋印；因為奉王的名所寫、用王的戒指蓋印的諭旨是不能廢除的。」
ESTH|8|9|三月，就是西彎月二十三日，當時王的一些書記受召而來，按著 末底改 所吩咐的，用各省的文字、各族的語言，以及 猶太 人的文字語言寫諭旨，傳給那從 印度 直到 古實 一百二十七省的 猶太 人，以及總督、省長和領袖。
ESTH|8|10|末底改 奉 亞哈隨魯 王的名寫諭旨，用王的戒指蓋印，交給信差們騎上御用的王室快馬去頒佈。
ESTH|8|11|王准各城各鎮的 猶太 人在一日之內，在十二月，就是亞達月的十三日聚集，在 亞哈隨魯 王的各省保護自己的性命，剪除，殺戮，滅絕那要攻擊 猶太 人的各省各族所有的軍隊，以及他們的妻子兒女，奪取他們的財產為掠物。
ESTH|8|12|
ESTH|8|13|這諭旨的抄本以敕令的方式在各省頒佈，通知各族，使 猶太 人預備等候那日，好在仇敵身上報仇。
ESTH|8|14|於是騎御用快馬的信差奉王命催促，急忙起行；敕令傳遍了 書珊 城堡。
ESTH|8|15|末底改 穿著藍色白色的朝服，頭戴大金冠冕，又穿紫色細麻布的外袍，從王面前出來； 書珊城 充滿了歡樂的呼聲。
ESTH|8|16|猶太 人有光榮，歡喜快樂，得享尊貴。
ESTH|8|17|王的諭旨和敕令所到的各省各城， 猶太 人都歡喜快樂，擺設宴席，以那日為吉日。國中許多民族的人因懼怕 猶太 人，就自稱為 猶太 人。
ESTH|9|1|十二月，就是亞達月十三日，王的諭旨和敕令要執行的那一日， 猶太 人的仇敵盼望制伏他們，但 猶太 人反倒制伏了恨他們的人。
ESTH|9|2|猶太 人在 亞哈隨魯 王各省的城裏聚集，下手擊殺那些要害他們的人。沒有人能在他們面前站立得住，因為各民族都懼怕他們。
ESTH|9|3|各省的領袖、總督、省長，和辦理王事務的人，因懼怕 末底改 ，就都幫助 猶太 人。
ESTH|9|4|末底改 在朝中為大，名聲傳遍各省； 末底改 這人的權勢日漸擴大。
ESTH|9|5|猶太 人用刀擊殺所有的仇敵，殺滅他們，隨意待那些恨他們的人。
ESTH|9|6|在 書珊 城堡中， 猶太 人殺滅了五百人。
ESTH|9|7|他們殺了 巴珊大他 、 達分 、 亞斯帕他 、
ESTH|9|8|破拉他 、 亞大利雅 、 亞利大他 、
ESTH|9|9|帕瑪斯他 、 亞利賽 、 亞利代 、 瓦耶撒他 ；
ESTH|9|10|這十人都是 哈米大他 的孫子， 猶太 人的仇敵 哈曼 的兒子。 猶太 人卻沒有下手奪取財物。
ESTH|9|11|那日， 書珊 城堡中被殺的人數呈報到王面前。
ESTH|9|12|王對 以斯帖 王后說：「 猶太 人在 書珊 城堡中殺滅了五百人，又殺了 哈曼 的十個兒子，在王其餘的各省不知如何。你要甚麼，必賜給你；你還求甚麼，也必為你成就。」
ESTH|9|13|以斯帖 說：「王若以為好，求你允准 書珊 的 猶太 人，明日也照今日的諭旨去做，並把 哈曼 十個兒子的屍體掛在木架上。」
ESTH|9|14|王允准這麼做。敕令傳遍 書珊 ， 哈曼 十個兒子的屍體被掛了起來。
ESTH|9|15|亞達月十四日，在 書珊 的 猶太 人又聚集，在 書珊 殺了三百人，卻沒有下手奪取財物。
ESTH|9|16|亞達月十三日，在王各省其餘的 猶太 人也都聚集，保護自己的性命，擺脫仇敵得享平安。他們殺了七萬五千個恨他們的人，卻沒有下手奪取財物；十四日他們休息，以這日為設宴歡樂的日子。
ESTH|9|17|
ESTH|9|18|但 書珊 的 猶太 人卻在十三日、十四日聚集；十五日休息，以這日為設宴歡樂的日子。
ESTH|9|19|所以住在無城牆的鄉村的 猶太 人，都以亞達月十四日為設宴歡樂的吉日，彼此餽送禮物。
ESTH|9|20|末底改 記錄這些事，寫信給 亞哈隨魯 王各省遠近所有的 猶太 人，
ESTH|9|21|吩咐他們每年守亞達月十四、十五兩日，
ESTH|9|22|以這兩日為 猶太 人擺脫仇敵得享平安、轉憂為喜、轉悲為樂的吉日，並在這兩日設宴歡樂，彼此餽送禮物，賙濟窮人。
ESTH|9|23|於是， 猶太 人照 末底改 所寫給他們的，把開始所做的作為遵守的定例。
ESTH|9|24|因為 猶太 人的仇敵 亞甲 人 哈米大他 的兒子 哈曼 設謀要殺害 猶太 人，抽普珥，普珥即籤，為要殺盡滅絕他們；
ESTH|9|25|但這陰謀 到了王面前，王卻降旨使 哈曼 謀害 猶太 人的惡事歸到他自己的頭上，他和他的眾子都被掛在木架上。
ESTH|9|26|所以 猶太 人照著普珥這名字稱這兩日為普珥日。他們因這信上一切的話，又因所看見所遇見的事，
ESTH|9|27|就規定自己與後裔，以及歸化他們的人，每年按所寫的、按時守這兩日，永久不廢。
ESTH|9|28|各省各城、世世代代、家家戶戶都記念並守這兩日，使這普珥日在 猶太 人中不可廢掉，在他們後裔中也永不遺忘。
ESTH|9|29|亞比孩 的女兒 以斯帖 王后和 猶太 人 末底改 以全權寫第二封信，堅立這普珥日，
ESTH|9|30|送信給 亞哈隨魯 王國中一百二十七省所有的 猶太 人，祝他們平安和安穩，
ESTH|9|31|勸他們遵照 猶太 人 末底改 和 以斯帖 王后所規定的，按時守這普珥日，並照著 猶太 人為自己與後裔所規定的，禁食與哀求。
ESTH|9|32|以斯帖 規定了守普珥日的條例，這事也記錄在書上。
ESTH|10|1|亞哈隨魯 王向國中和海島的人徵稅。
ESTH|10|2|他以權柄能力所做的一切，以及他使 末底改 尊大、提升他的事，豈不都寫在 瑪代 和 波斯 王的史籍上嗎？
ESTH|10|3|猶太 人 末底改 作 亞哈隨魯 王的宰相，在 猶太 人中為大，得許多弟兄的喜悅，為本族的人爭取福利，為他所有的後代謀求幸福。
JOB|1|1|烏斯 地有一個人名叫 約伯 。這人完全、正直、敬畏上帝、遠離惡事。
JOB|1|2|他生了七個兒子，三個女兒。
JOB|1|3|他的家產有七千隻羊，三千匹駱駝，五百對牛，五百匹母驢，並有許多僕婢。這人在東方人中為至大。
JOB|1|4|他的兒子按著日子各在自己家裏擺設宴席，派人去請他們的三個姊妹來，與他們一同吃喝。
JOB|1|5|宴席的日子過了， 約伯 派人去叫他們自潔。他清早起來，按著他們眾人的數目獻燔祭，因為他說：「恐怕我的兒子犯了罪，心中背棄 上帝。」 約伯 常常這樣行。
JOB|1|6|有一天，上帝的眾使者 來侍立在耶和華面前，撒但也來在其中。
JOB|1|7|耶和華對撒但說：「你從哪裏來？」撒但回答耶和華說：「我從地上走來走去，在那裏往返。」
JOB|1|8|耶和華對撒但說：「你曾用心察看我的僕人 約伯 沒有？地上再沒有人像他那樣完全、正直、敬畏上帝、遠離惡事。」
JOB|1|9|撒但回答耶和華說：「 約伯 敬畏上帝，豈是無故呢？
JOB|1|10|你豈不是四面圈上籬笆圍護他和他的家，以及他一切所有的嗎？他手所做的都蒙你賜福，他的家產也在地上增多。
JOB|1|11|但你若伸手毀他一切所有的，他必當面背棄你。」
JOB|1|12|耶和華對撒但說：「看哪，凡他所有的都在你手中；只是不可伸手加害於他。」於是撒但從耶和華面前退出去。
JOB|1|13|有一天， 約伯 的兒女正在他們長兄的家裏吃飯喝酒，
JOB|1|14|有報信的來見 約伯 ，說：「牛正耕地，母驢在旁邊吃草，
JOB|1|15|示巴 人忽然闖來，把牲畜擄去，並用刀殺了僕人；惟有我一人逃脫，來報信給你。」
JOB|1|16|他還說話的時候，又有人來說：「上帝從天上降下火來，把羊群和僕人都吞滅了；惟有我一人逃脫，來報信給你。」
JOB|1|17|他還說話的時候，又有人來說：「 迦勒底 人分成三隊忽然闖來，把駱駝擄去，並用刀殺了僕人；惟有我一人逃脫，來報信給你。」
JOB|1|18|他還說話的時候，又有人來說：「你的兒女正在他們長兄的家裏吃飯喝酒，
JOB|1|19|看哪，有狂風從曠野颳來，襲擊房屋的四角，房屋倒塌在年輕人身上，他們就都死了；惟有我一人逃脫，來報信給你。」
JOB|1|20|約伯 就起來，撕裂外袍，剃了頭，俯伏在地敬拜，
JOB|1|21|說：「我赤身出於母胎，也必赤身歸回；賞賜的是耶和華，收取的也是耶和華。耶和華的名是應當稱頌的。」
JOB|1|22|在這一切的事上， 約伯 並沒有犯罪，也不以上帝為狂妄。
JOB|2|1|又有一天，上帝的眾使者 來侍立在耶和華面前，撒但也來在其中。
JOB|2|2|耶和華問撒但說：「你從哪裏來？」撒但回答說：「我從地上走來走去，在那裏往返。」
JOB|2|3|耶和華對撒但說：「你曾用心察看我的僕人 約伯 沒有？地上再沒有人像他那樣完全、正直、敬畏上帝、遠離惡事。你雖激起我攻擊他，無故吞滅他，他仍然持守他的純正。」
JOB|2|4|撒但回答耶和華說：「人以皮代皮，情願捨去一切所有的，來保全性命。
JOB|2|5|但你若伸手傷他的骨頭和他的肉，他必當面背棄 你。」
JOB|2|6|耶和華對撒但說：「看哪，他在你手中，只要留下他的性命。」
JOB|2|7|於是撒但從耶和華面前退出去，擊打 約伯 ，使他從腳掌到頭頂長毒瘡。
JOB|2|8|約伯 就坐在灰燼中，拿瓦片刮身體。
JOB|2|9|他的妻子對他說：「你仍然持守你的純正嗎？你背棄上帝，死了吧！」
JOB|2|10|約伯 卻對她說：「你說話，正如愚頑的婦人。唉！難道我們從上帝手裏得福，不也受禍嗎？」在這一切的事上， 約伯 並沒有以口犯罪。
JOB|2|11|約伯 的三個朋友， 提幔 人 以利法 、 書亞 人 比勒達 、 拿瑪 人 瑣法 ，聽說這一切的災禍臨到他身上，各人就從自己的地方相約同來，為他悲傷，安慰他。
JOB|2|12|他們遠遠地舉目觀看，認不出他來，就放聲大哭。各人撕裂外袍，向空中撒塵土，落在自己的頭上。
JOB|2|13|他們同他七天七夜坐在地上，一句話也不對他說，因為他們見到了極大的痛苦。
JOB|3|1|此後， 約伯 開口詛咒自己的生日 。
JOB|3|2|約伯 說：
JOB|3|3|「願我生的那日滅沒， 說『懷了男胎』的那夜也滅沒。
JOB|3|4|願那日變為黑暗， 願上帝不從上面尋找它， 願亮光不照於其上。
JOB|3|5|願黑暗和死蔭索取那日， 願密雲停在其上， 願白天的昏暗 恐嚇它。
JOB|3|6|願那夜被幽暗奪取， 不在一年的日子中喜樂， 也不列入月中的數目。
JOB|3|7|看哪，願那夜沒有生育， 其間也沒有歡樂的聲音。
JOB|3|8|願那些詛咒日子且能惹動 力威亞探 的， 詛咒那夜。
JOB|3|9|願那夜黎明的星宿變為黑暗， 盼亮卻不亮， 也不見晨曦破曉 ；
JOB|3|10|因它沒有把懷我胎的門關閉， 也沒有從我的眼中隱藏患難。
JOB|3|11|「我為何不出母胎而死？ 為何不出母腹就氣絕呢？
JOB|3|12|為何有膝蓋接收我？ 為何有奶哺養我呢？
JOB|3|13|不然，我現在已躺臥安睡， 而且，早已長眠安息；
JOB|3|14|與那些為自己重建荒涼之處， 地上的君王和謀士在一起；
JOB|3|15|或與把銀子裝滿房屋， 擁有金子的王子在一起；
JOB|3|16|我為何不像流產的胎兒被埋藏， 如同未見光的嬰孩？
JOB|3|17|在那裏惡人止息攪擾， 在那裏困乏人得享安息，
JOB|3|18|被囚的人同得安逸， 不再聽見監工的聲音。
JOB|3|19|大的小的都在那裏， 奴僕脫離主人得自由。
JOB|3|20|「遭受患難的人為何有光賜給他呢？ 心中愁苦的人為何有生命賜給他呢？
JOB|3|21|他們等死，卻不得死； 求死，勝於求隱藏的珍寶。
JOB|3|22|他們尋見墳墓， 就歡喜快樂，極其高興。
JOB|3|23|這人的道路遮隱， 上帝又四面圍困他。
JOB|3|24|我吃飯前就發出嘆息， 我的唉哼湧出如水。
JOB|3|25|因我所恐懼的臨到我， 我所懼怕的迎向我；
JOB|3|26|我不得安逸，不得平靜， 也不得安息，卻有患難來到。」
JOB|4|1|提幔 人 以利法 回答說：
JOB|4|2|「人想與你說話，你就厭煩嗎？ 但誰能忍住不發言呢？
JOB|4|3|看哪，你素來教導許多人， 又堅固軟弱的手。
JOB|4|4|你的言語曾扶助跌倒的人； 你使軟弱的膝蓋穩固。
JOB|4|5|但現在禍患臨到 你，你就煩躁了； 它挨近你，你就驚惶。
JOB|4|6|你的倚靠不是在於你敬畏上帝嗎？ 你的盼望不是在於你行事純正嗎？
JOB|4|7|「請你追想：無辜的人有誰滅亡？ 正直的人何處被剪除？
JOB|4|8|按我所見，耕罪孽的， 種毒害的，照樣收割。
JOB|4|9|上帝一噓氣，他們就滅亡； 上帝一發怒，他們就消失。
JOB|4|10|獅子吼叫，猛獅咆哮， 少壯獅子的牙齒被敲斷。
JOB|4|11|公獅因缺獵物而死， 母獅的幼獅都離散。
JOB|4|12|「有話暗中傳遞給我， 耳朵聽其微小的聲音。
JOB|4|13|世人沉睡的時候， 從夜間異象的雜念中，
JOB|4|14|恐懼戰兢臨到我身， 使我百骨戰抖。
JOB|4|15|有靈從我面前經過， 我身上的毫毛豎立。
JOB|4|16|那靈停住， 我卻不能辨其形狀； 有形像在我眼前。 我在靜默中聽見有聲音：
JOB|4|17|『必死的人能比上帝公義嗎？ 壯士能比造他的主純潔嗎？
JOB|4|18|看哪，主不信靠他的僕人， 尚且指他的使者為愚昧，
JOB|4|19|何況那些住在泥屋、 根基在塵土裏、 被蛀蟲所毀壞的人呢？
JOB|4|20|早晚之間，他們就被毀滅， 永歸無有，無人理會。
JOB|4|21|他們帳棚的繩索豈不從中拔出來呢？ 他們死，且是無智慧而死。』」
JOB|5|1|「你呼求吧，有誰回答你呢？ 聖者之中，你轉向哪一位呢？
JOB|5|2|憤怒害死愚妄人， 嫉妒殺死愚蠢的人。
JOB|5|3|我曾見愚妄人扎下根， 但我忽然詛咒他的住處。
JOB|5|4|他的兒女遠離穩妥之地， 在城門口被欺壓，無人搭救。
JOB|5|5|他的莊稼被飢餓的人吃盡了， 就是在荊棘裏的也搶去了； 他的財寶被陷阱 張口吞沒了。
JOB|5|6|因為禍患不是從塵土中出來， 患難也不是從土地裏長出。
JOB|5|7|人生出來必遭遇患難， 如同火花 飛騰。
JOB|5|8|「至於我，我必尋求上帝， 把我的事情交託給他。
JOB|5|9|他行大事不可測度， 行奇事不可勝數。
JOB|5|10|他降雨在地面， 賜水於田野。
JOB|5|11|他將卑微的人安置在高處， 將哀痛的人舉到穩妥之地。
JOB|5|12|他破壞通達人的計謀， 使他們手所做的不得成就。
JOB|5|13|他使有智慧的人中了自己的詭計， 叫狡詐人的計謀速速落空。
JOB|5|14|他們白晝遇見黑暗， 午間摸索如在夜間。
JOB|5|15|上帝拯救貧窮人脫離殘暴人的手， 脫離他們口中的刀。
JOB|5|16|這樣，貧寒人有指望， 不義的人閉口無言。
JOB|5|17|「看哪，上帝所懲治的人是有福的！ 所以你不可輕看全能者的管教。
JOB|5|18|因為他打傷，又包紮； 他擊傷，又親手醫治。
JOB|5|19|你六次遭難，他必救你； 就是七次，災禍也無法害你。
JOB|5|20|在饑荒中，他必救你脫離死亡； 在戰爭中，他必救你脫離刀劍的權勢。
JOB|5|21|你必被隱藏，不受口舌之害； 災害臨到，你也不懼怕。
JOB|5|22|對於災害饑饉，你必譏笑； 至於地上的野獸，你也不懼怕。
JOB|5|23|因為你必與田間的石頭立約， 田裏的野獸也必與你和好。
JOB|5|24|你必知道你的帳棚平安， 你查看你的羊圈，一無所失。
JOB|5|25|你也必知道你的後裔眾多， 你的子孫像地上的青草。
JOB|5|26|你必壽高年邁才歸墳墓， 好像禾捆按時收藏。
JOB|5|27|看哪，這道理我們已經考察，本是如此。 你須要聽，要親自明白。」
JOB|6|1|約伯 回答說：
JOB|6|2|「惟願我的煩惱被秤一秤， 我一切的災害放在天平裏，
JOB|6|3|現今都比海沙更重， 所以我說話急躁。
JOB|6|4|因全能者的箭射中了我， 我的靈喝盡其毒； 上帝的驚嚇擺陣攻擊我。
JOB|6|5|野驢有草豈會叫喚？ 牛有飼料豈會吼叫？
JOB|6|6|食物淡而無鹽豈可吃呢？ 蛋白有甚麼滋味呢？
JOB|6|7|那些可厭的食物， 我心不肯挨近。
JOB|6|8|「惟願我得著所求的， 上帝賞賜我所切望的，
JOB|6|9|願上帝把我壓碎， 伸手將我剪除。
JOB|6|10|我因沒有違棄那聖者的言語， 就仍以此為安慰， 在不止息的痛苦中還可歡躍。
JOB|6|11|我有甚麼氣力使我等候？ 我有甚麼結局使我忍耐？
JOB|6|12|我的氣力豈是石頭的氣力？ 我的肉身豈是銅呢？
JOB|6|13|在我裏面豈不是無助嗎？ 智慧豈不是從我心中被趕逐嗎？
JOB|6|14|「灰心的人，他的朋友當以慈愛待他， 因為他將離棄敬畏全能者的心。
JOB|6|15|我的弟兄詭詐，好像河道， 像溪水流過的河床，
JOB|6|16|因結冰而混濁， 有雪藏在其中，
JOB|6|17|暖和的時候就溶化， 炎熱時便從原處乾涸。
JOB|6|18|商隊偏離道路， 上到荒涼之地而死亡。
JOB|6|19|提瑪 的商隊瞻望， 示巴 的旅客等候。
JOB|6|20|他們因希望落空就抱愧， 來到那裏便蒙羞。
JOB|6|21|現在你們正是這樣 ， 看見驚嚇的事就懼怕。
JOB|6|22|我豈說：『請你們供給我， 從你們的財物中送禮給我』？
JOB|6|23|或說：『請你們拯救我脫離敵人的手， 救贖我脫離殘暴人的手』嗎？
JOB|6|24|「請你們指教我，我就不作聲； 我在何事上有錯，請使我明白。
JOB|6|25|正直言語的力量何其大！ 但你們責備是責備甚麼呢？
JOB|6|26|絕望人的講論既然如風， 你們還計劃批駁言語嗎？
JOB|6|27|你們甚至為孤兒抽籤， 把朋友當貨物。
JOB|6|28|「現在，請你們看著我， 我絕不當面說謊。
JOB|6|29|請你們轉意，不要不公義； 請再轉意，正義在我這裏。
JOB|6|30|我的舌頭豈有不公義嗎？ 我的上膛豈不辨奸惡嗎？」
JOB|7|1|「人在世上豈無勞役呢？ 他的日子不像雇工的日子嗎？
JOB|7|2|像奴僕切慕陰涼， 像雇工等待工錢，
JOB|7|3|我也照樣度過虛空的歲月， 愁煩的夜晚指定給我。
JOB|7|4|我躺臥的時候就說： 『我何時可以起來呢？』漫漫長夜， 我總是翻來覆去，直到天亮。
JOB|7|5|我的肉體以蟲子和塵土為衣， 我的皮膚才收了口又流膿。
JOB|7|6|我的日子比織布的梭更快， 都消耗在沒有指望之中。
JOB|7|7|「你要記得，我的生命不過是一口氣， 我的眼睛必不再看見福樂。
JOB|7|8|觀看我的人，他的眼必不看見我； 你的眼目投向我，我卻不在了。
JOB|7|9|雲彩消散而去； 照樣，人下陰間也不再上來。
JOB|7|10|他不再回自己的家， 他自己的地方也不再認得他。
JOB|7|11|「我甚至不封我的口； 我靈愁苦，要發出言語； 我心苦惱，要吐露哀情。
JOB|7|12|我豈是海洋，豈是大魚， 你竟防守著我呢？
JOB|7|13|我若說：『我的床必安慰我， 我的榻必分擔我的苦情』，
JOB|7|14|你就用夢驚擾我， 用異象恐嚇我。
JOB|7|15|甚至我寧可窒息死亡， 勝似留我這副骨頭。
JOB|7|16|我厭棄生命，不願永遠活著。 你任憑我吧，因我的日子都是虛空。
JOB|7|17|人算甚麼，你竟看他為大， 將他放在心上，
JOB|7|18|每早晨鑒察他， 每時刻考驗他？
JOB|7|19|你到何時才轉眼不看我， 任憑我咽下唾沫呢？
JOB|7|20|鑒察人的主啊，我若有罪，於你何妨？ 為何以我當你的箭靶， 使我成為你的重擔呢？
JOB|7|21|為何不赦免我的過犯， 除掉我的罪孽呢？ 我現今要躺臥在塵土中； 你要切切尋找我，我卻不在了。」
JOB|8|1|書亞 人 比勒達 回答說：
JOB|8|2|「這些話你要說到幾時？ 你口中的言語如狂風要到幾時呢？
JOB|8|3|上帝豈能偏離公平？ 全能者豈能偏離公義？
JOB|8|4|或者你的兒女得罪了他， 他就把他們交在過犯的掌控中。
JOB|8|5|你若切切尋求上帝， 向全能者懇求；
JOB|8|6|你若純潔正直， 他必定為你興起， 使你公義的居所興旺。
JOB|8|7|你起初雖然微小， 日後必非常強盛。
JOB|8|8|「請你詢問上代， 思念他們祖先所查究的。
JOB|8|9|我們不過從昨日才有，一無所知， 因我們在世的日子好像影子。
JOB|8|10|他們豈不指教你，告訴你， 說出發自內心的言語呢？
JOB|8|11|「蒲草沒有泥豈能生長？ 蘆荻沒有水豈能長大？
JOB|8|12|它還青翠，沒有割下的時候， 比百樣的草先枯槁。
JOB|8|13|凡忘記上帝的人，路途也是這樣； 不虔敬人的指望要滅沒。
JOB|8|14|他所仰賴的必折斷， 他所倚靠的是蜘蛛網。
JOB|8|15|他要倚靠房屋，房屋卻站立不住； 他要抓住房屋，房屋卻不能存留。
JOB|8|16|他在日光之下茂盛， 嫩枝在園中蔓延；
JOB|8|17|他的根盤繞石堆， 鑽入石縫 。
JOB|8|18|他若從本地被拔出， 那地就不認識他，說：『我沒有見過你。』
JOB|8|19|看哪，這就是他道路中的喜樂， 以後必另有人從塵土而生。
JOB|8|20|看哪，上帝必不丟棄完全人， 也不扶助邪惡人的手。
JOB|8|21|他還要以喜笑充滿你的口， 以歡呼充滿你的嘴唇。
JOB|8|22|恨惡你的要披戴羞愧， 惡人的帳棚必歸於無有。」
JOB|9|1|約伯 回答說：
JOB|9|2|「我真的知道是這樣， 但人在上帝前怎能成為義呢？
JOB|9|3|人若想要與他爭辯， 千次中也不能回答一次。
JOB|9|4|他心裏有智慧，且大有能力。 誰向上帝剛硬而得平安呢？
JOB|9|5|他把山挪移，山卻不知， 他在怒氣中，把山翻倒。
JOB|9|6|他使地震動，離其本位， 地的柱子就搖撼。
JOB|9|7|他吩咐太陽，太陽就不出來， 又封住眾星。
JOB|9|8|他獨自鋪張諸天， 步行在海浪之上。
JOB|9|9|他造北斗、參星、昴星， 以及南方的星宿 ；
JOB|9|10|他行大事不可測度， 行奇事不可勝數。
JOB|9|11|看哪，他從我旁邊經過，我看不見； 他走過，我沒有察覺他。
JOB|9|12|看哪，他奪去，誰能阻擋他？ 誰敢對他說：『你做甚麼呢？』
JOB|9|13|「上帝必不收回他的怒氣， 扶助 拉哈伯 的，屈身在上帝以下。
JOB|9|14|既是這樣，我怎敢回答他， 怎敢在他之前選擇辯詞呢？
JOB|9|15|我雖有義，也不能回答， 我要向那審判我的懇求。
JOB|9|16|我若呼求，縱然他應允我， 我仍不信他會側耳聽我的聲音。
JOB|9|17|他用暴風 摧折我， 無故加增我的損傷。
JOB|9|18|他不容我喘一口氣， 倒使我飽受苦惱。
JOB|9|19|若論力量，看哪，他真有能力！ 若論審判，『誰能傳我呢？』
JOB|9|20|我雖有義，我的口要定我有罪； 我雖完全，他必證明我為彎曲。
JOB|9|21|我雖完全，不顧自己； 我厭棄我的性命。
JOB|9|22|所以我說，都是一樣； 完全人和惡人，他都滅絕。
JOB|9|23|若災禍忽然帶來死亡， 他必戲笑無辜人的苦難。
JOB|9|24|世界交在惡人手中； 他蒙蔽世界審判官的臉， 若不是他，那麼是誰呢？
JOB|9|25|「我的日子比奔跑者更快， 急速過去，不見福樂。
JOB|9|26|我的日子如蒲草船掠過， 如鷹俯衝抓食。
JOB|9|27|我若說：『我要忘記我的苦情， 強顏歡笑』，
JOB|9|28|我就因一切的愁苦而懼怕； 我知道你必不以我為無辜。
JOB|9|29|我必被定罪， 我何必徒然勞苦呢？
JOB|9|30|我若用雪水洗身， 用鹼潔淨我的手掌，
JOB|9|31|你還要把我扔在坑裏， 我的衣服都憎惡我。
JOB|9|32|他不像我是個人，使我可以回答他， 使我們可以一同受審判。
JOB|9|33|我們中間沒有仲裁者， 可以按手在我們兩造之間。
JOB|9|34|願他使他的杖離開我， 不使他的威嚴恐嚇我，
JOB|9|35|我就說話，不懼怕他； 但對我來說，我卻不是這樣。」
JOB|10|1|「我厭惡自己的性命， 任由我述說自己的苦情； 因心裏苦惱，我要說話。
JOB|10|2|我對上帝說，不要定我有罪， 要指示我，你為何與我爭辯？
JOB|10|3|你手所造的，你又欺壓，又藐視， 卻光照惡人的計謀。 這事你以為美嗎？
JOB|10|4|你的眼豈是肉眼？ 你察看豈像人察看嗎？
JOB|10|5|你的日子豈像人的日子， 你的年歲豈像壯士的年歲，
JOB|10|6|你就追問我的罪孽， 尋察我的罪過嗎？
JOB|10|7|其實，你知道我沒有行惡， 也無人能施行拯救，脫離你的手。
JOB|10|8|你的手塑造我，造了我， 但我整個人卻要一起被你吞滅。
JOB|10|9|求你記得，你製造我如泥土， 你還要使我歸回塵土嗎？
JOB|10|10|你不是倒出我來好像奶， 使我凝結如同奶酪嗎？
JOB|10|11|你以皮和肉給我穿上， 用骨與筋把我聯結起來。
JOB|10|12|你將生命和慈愛賜給我， 你也眷顧保全我的靈。
JOB|10|13|然而，你把這些事藏在你心裏， 我知道這是你的旨意。
JOB|10|14|我若犯罪，你就察看我， 並不赦免我的罪。
JOB|10|15|我若行惡，我就有禍了； 我若行義，也不敢抬頭， 而是飽受羞辱， 看見我的痛苦。
JOB|10|16|你如獅子昂首追捕我 ， 又在我身上顯出奇事。
JOB|10|17|你更新你的見證對付我， 向我加增惱怒， 調遣軍隊攻擊我。
JOB|10|18|「你為何使我出母胎呢？ 甚願我當時氣絕，沒有眼睛看見我。
JOB|10|19|這樣，就如從未有過我， 我一出母胎就被送入墳墓。
JOB|10|20|我的日子不是短少嗎？求你停止， 求你放過我 ，使我可以稍得喜樂，
JOB|10|21|就是在我去而不返， 往黑暗和死蔭之地以先。
JOB|10|22|那是烏黑之地， 猶如幽暗的死蔭， 毫無秩序； 發出的光輝也像幽暗。」
JOB|11|1|拿瑪 人 瑣法 回答說：
JOB|11|2|「這許多的話豈不該回答嗎？ 多嘴多舌的人豈可成為義呢？
JOB|11|3|你誇大的話豈能使人不作聲嗎？ 你戲笑的時候豈沒有人使你受辱嗎？
JOB|11|4|你說：『我的教導純全， 我在你眼前是清潔的。』
JOB|11|5|但是，惟願上帝說話， 願他張開嘴唇攻擊你。
JOB|11|6|願他將智慧的奧祕指示你， 因為健全的知識是兩面的。 你當知道，上帝使你忘記你的一些罪孽。
JOB|11|7|你能尋見上帝的奧祕嗎？ 你能尋見全能者的極限嗎？
JOB|11|8|高如諸天，你能做甚麼？ 比陰間深，你能知道甚麼？
JOB|11|9|其量度比地長， 比海更寬。
JOB|11|10|他若經過，把人拘禁， 召集會眾，誰能阻擋他呢？
JOB|11|11|因為他知道虛妄的人； 當他看見罪惡，豈不留意嗎？
JOB|11|12|空虛的人若獲得知識， 野驢生下的駒子也成了人。
JOB|11|13|「至於你，若堅固己心， 又向主舉手；
JOB|11|14|你若遠遠脫離你手中的罪孽， 不容許不義住在你帳棚之中；
JOB|11|15|這樣，你必仰起臉來，毫無瑕疵； 你也必安穩，無所懼怕。
JOB|11|16|你必忘記你的苦楚， 就是想起來，也如流過的水。
JOB|11|17|你在世要升高，比正午更明， 雖有黑暗，仍像早晨。
JOB|11|18|你因有指望就必穩固， 也必四圍察看 ，安然躺下。
JOB|11|19|你躺臥，無人驚嚇， 並有許多人向你求恩。
JOB|11|20|但惡人的眼睛要失明； 他們無路可逃， 他們的指望就是氣絕身亡。」
JOB|12|1|約伯 回答說：
JOB|12|2|「你們果真是人物啊！ 智慧要與你們一同去死。
JOB|12|3|但我也有聰明，跟你們一樣， 並非不及你們。 這些事，誰不知道呢？
JOB|12|4|我這求告上帝、蒙他應允的人 竟成了朋友所譏笑的； 又公義又完全的人竟遭受譏笑。
JOB|12|5|安逸的人心裏藐視災禍， 這災禍在等待失足滑跌的人。
JOB|12|6|強盜的帳棚安寧， 惹上帝發怒的人穩固， 他們把上帝 握在自己手中 。
JOB|12|7|「你問走獸，走獸必指教你； 你問空中的飛鳥，飛鳥必告訴你；
JOB|12|8|或者你與地說話，地必指教你 ； 海中的魚也必向你說明。
JOB|12|9|在這一切當中， 有誰不知道這是耶和華的手做成的呢？
JOB|12|10|凡動物的生命 和人類的氣息都在他手中。
JOB|12|11|耳朵豈不辨別言語， 正如上膛品嘗食物嗎？
JOB|12|12|年老的有智慧， 壽高的有知識。
JOB|12|13|「在上帝有智慧和能力， 他有謀略和知識。
JOB|12|14|看哪，他拆毀，就不能重建； 他拘禁人，人就不得釋放。
JOB|12|15|看哪，他使水止住，水就乾了； 他把水放出，水就淹沒大地。
JOB|12|16|在他有能力和智慧， 走迷的和使人迷路的都屬他。
JOB|12|17|他把謀士剝衣擄去， 使審判官變為愚妄。
JOB|12|18|他解除君王的權勢 ， 用帶子捆住他們的腰。
JOB|12|19|他把祭司剝衣擄去， 使有權能的人傾覆。
JOB|12|20|他廢去忠信者的言論， 奪去長者的見識。
JOB|12|21|他使貴族蒙羞受辱， 放鬆勇士的腰帶。
JOB|12|22|他從黑暗中彰顯深奧的事， 使死蔭顯出光明。
JOB|12|23|他使邦國興旺而又毀滅， 使邦國擴展又被掠奪。
JOB|12|24|他將地上百姓中領袖的聰明奪去， 使他們迷失在荒涼無路之地。
JOB|12|25|他們在無光的黑暗中摸索； 他使他們搖晃像醉酒的人一樣。」
JOB|13|1|「看哪，這一切，我眼都見過； 我耳都聽過，而且明白。
JOB|13|2|你們所知道的，我也知道， 並非不及你們。
JOB|13|3|然而我要對全能者說話， 我願與上帝理論。
JOB|13|4|但你們是編造謊言的， 全都是無用的醫生。
JOB|13|5|惟願你們全然不作聲， 這就是你們的智慧！
JOB|13|6|請你們聽我的答辯， 留心聽我嘴唇的訴求。
JOB|13|7|你們要為上帝說不義的話嗎？ 要為他說詭詐的言語嗎？
JOB|13|8|你們要看上帝的情面嗎？ 要為他爭辯嗎？
JOB|13|9|他查究你們，這豈是好事嗎？ 人欺騙人，你們也要照樣欺騙他嗎？
JOB|13|10|你們若暗中看人的情面， 他必定要責備你們。
JOB|13|11|他的尊榮豈不叫你們懼怕嗎？ 他豈不使驚嚇臨到你們嗎？
JOB|13|12|你們可記念的諺語是灰燼的箴言； 你們的後盾是泥土的後盾。
JOB|13|13|「你們不要向我作聲， 讓我說話，無論如何我都承當。
JOB|13|14|我為何把我的肉掛在我的牙上， 將我的命放在我的手掌中呢？
JOB|13|15|看哪，他要殺我，我毫無指望 ， 然而我還要在他面前辯明我所行的。
JOB|13|16|這要成為我的拯救， 因為不虔誠的人不可到他面前。
JOB|13|17|你們要細聽我的言語， 讓我的申辯入你們耳中。
JOB|13|18|看哪，我已陳明我的案， 知道自己有義。
JOB|13|19|還有誰要和我爭辯， 我現在就緘默不言，氣絕而死。
JOB|13|20|惟有兩件事不要向我施行， 我就不躲開你的面：
JOB|13|21|就是把你的手縮回，遠離我身； 又不使你的威嚴恐嚇我。
JOB|13|22|這樣，你呼叫，我就回答； 或是讓我說話，你回答我。
JOB|13|23|我的罪孽和我的罪有多少呢？ 求你叫我知道我的過犯與我的罪。
JOB|13|24|你為何轉臉， 拿我當仇敵呢？
JOB|13|25|你要驚動被風吹的葉子嗎？ 要追趕枯乾的碎秸嗎？
JOB|13|26|你寫下苦楚對付我， 又使我擔當幼年的罪孽。
JOB|13|27|你把我的腳鎖上木枷， 察看我一切的道路， 為我的腳掌劃定界限。
JOB|13|28|人像滅絕的爛物， 像蟲蛀的衣裳。」
JOB|14|1|「人為婦人所生， 日子短少，多有患難。
JOB|14|2|他出來如花，凋謝而去； 他飛逝如影，不能存留。
JOB|14|3|這樣的人你豈會睜眼看他， 又叫我 來，在你那裏受審嗎？
JOB|14|4|誰能使潔淨出於污穢呢？ 誰也不能！
JOB|14|5|既然人的日子限定， 他的月數在於你， 你劃定他的界限，他不能越過；
JOB|14|6|求你轉眼不看他，使他得歇息， 直到他像雇工享受他的一天。
JOB|14|7|「因樹有指望， 若被砍下，還可發芽， 嫩枝生長不息。
JOB|14|8|樹根若衰老在地裏， 樹幹也死在土中，
JOB|14|9|及至得了水氣，還會發芽， 長出枝條，像新栽的樹一樣。
JOB|14|10|但壯士一死就消逝了； 人一氣絕，他在何處呢？
JOB|14|11|海中的水枯竭， 江河消散乾涸。
JOB|14|12|人一躺下就不再起來， 等到諸天沒有了 ，仍不復醒， 也不能從睡中喚醒。
JOB|14|13|惟願你把我藏在陰間， 把我隱藏，直到你的憤怒過去； 願你為我定下期限，並記得我。
JOB|14|14|壯士若死了能再活嗎？ 我在一切服役的日子中等待， 直到我退伍的時候來到。
JOB|14|15|你呼叫，我就回答你； 你手所做的，你必期待。
JOB|14|16|但如今你數點我的腳步， 不察看我的罪。
JOB|14|17|我的過犯被你密封在囊中， 你遮掩了我的罪孽。
JOB|14|18|「然而，山崩變為無有， 磐石從原處挪移。
JOB|14|19|流水沖蝕石頭， 急流洗去地上的塵土； 你也照樣滅絕人的指望。
JOB|14|20|你終必勝過人，使他消逝； 你改變他的容貌，把他送走。
JOB|14|21|他的兒子得尊榮，他不知道； 他們降為卑，他也不曉得。
JOB|14|22|他只覺得身上疼痛， 心中為自己悲哀。」
JOB|15|1|提幔 人 以利法 回答說：
JOB|15|2|「智慧人豈可用虛空的知識回答， 用東風充滿自己的肚腹呢？
JOB|15|3|他豈可用無益的話， 用無濟於事的言語理論呢？
JOB|15|4|你誠然廢棄敬畏， 不在上帝面前默想。
JOB|15|5|你的罪孽指教你的口； 你選用詭詐人的舌頭。
JOB|15|6|你自己的口定你有罪，並非是我； 你自己的嘴唇見證你的不是。
JOB|15|7|「你是頭一個生下來的人嗎？ 你受造在諸山之先嗎？
JOB|15|8|你曾聽見上帝的密旨嗎？ 你要獨自得盡智慧嗎？
JOB|15|9|甚麼是你知道，我們不知道的呢？ 甚麼是你明白，我們不明白的呢？
JOB|15|10|我們這裏有白髮的和年老的， 比你父親還年長。
JOB|15|11|上帝的安慰和對你溫和的話， 你以為太小嗎？
JOB|15|12|你的心為何失控， 你的眼為何冒火，
JOB|15|13|以致你的靈反對上帝， 你的口說出這樣的言語呢？
JOB|15|14|人是甚麼，竟算為潔淨呢？ 婦人所生的是甚麼，竟算為義呢？
JOB|15|15|看哪，上帝不信任他的眾聖者； 在他眼前，天也不潔淨，
JOB|15|16|何況那污穢可憎， 喝罪孽如水的世人呢！
JOB|15|17|「我指示你，你要聽我； 我要陳述我所看見的，
JOB|15|18|就是智慧人從列祖所受， 傳講而不隱瞞的事。
JOB|15|19|這地惟獨賜給他們， 並沒有外人從他們中間經過。
JOB|15|20|惡人一生的日子絞痛難熬， 殘暴人存留的年數也是如此。
JOB|15|21|驚嚇的聲音常在他耳中； 在平安時，毀滅者必臨到他。
JOB|15|22|他不信自己能從黑暗中轉回； 他被刀劍看守。
JOB|15|23|他飄流在外求食：『哪裏有食物呢？』 他知道黑暗的日子在他手邊預備好了。
JOB|15|24|急難困苦叫他害怕， 而且勝過他，好像君王預備上陣。
JOB|15|25|因他伸手攻擊上帝， 逞強對抗全能者，
JOB|15|26|挺著頸項， 用盾牌堅厚的凸面向全能者直闖；
JOB|15|27|又因他的臉蒙上油脂， 腰上積滿肥肉。
JOB|15|28|他住在荒涼的城鎮， 房屋無人居住， 將成為廢墟。
JOB|15|29|他不得富足， 財物不得常存， 產業在地上也不加增。
JOB|15|30|他不得脫離黑暗， 火焰要把他的嫩枝燒乾； 因上帝口中的氣，他要離去。
JOB|15|31|不要讓他倚靠虛假，欺騙自己， 因虛假必成為他的報應。
JOB|15|32|他的日期未到之先，這事必實現； 他的枝子不得青綠。
JOB|15|33|他必像葡萄樹，葡萄未熟就掉落； 又像橄欖樹，一開花就凋謝。
JOB|15|34|因不敬虔之輩必不能生育， 受賄賂之人的帳棚必被火吞滅。
JOB|15|35|他們所懷的是毒害，所生的是罪孽， 肚腹裏所預備的是詭詐。」
JOB|16|1|約伯 回答說：
JOB|16|2|「這樣的話我聽了許多； 你們全都是使人愁煩的安慰者。
JOB|16|3|如風的言語有窮盡嗎？ 或者甚麼惹動你回答呢？
JOB|16|4|我也能說你們那樣的話， 你們若處在我的景況， 我也可以堆砌言詞攻擊你們， 又可以向你們搖頭。
JOB|16|5|但我必用口堅固你們， 顫動的嘴唇帶來舒解。
JOB|16|6|「我若說話，痛苦仍不得緩解； 我若停止，痛苦就離開我嗎？
JOB|16|7|但現在上帝使我困倦， 你使所有的親友遠離我，
JOB|16|8|你抓住我 ，成為見證起來攻擊我； 我的枯瘦也當著我的面作證。
JOB|16|9|上帝發怒撕裂我，逼迫我， 向我咬牙切齒； 我的敵人怒目瞪我。
JOB|16|10|他們向我大大張口， 打我的耳光羞辱我， 聚在一起攻擊我。
JOB|16|11|上帝把我交給不敬虔的人， 把我扔到惡人的手中。
JOB|16|12|我本是安逸，他折斷我， 掐住我的頸項，把我摔碎， 又立我作他的箭靶。
JOB|16|13|他的弓箭手圍繞我。 他刺破我的腎臟，並不留情， 把我的膽汁傾倒在地上。
JOB|16|14|他使我破裂，破裂又破裂， 如同勇士向我直闖。
JOB|16|15|「我把麻布縫在我的皮膚上， 把我的角放在塵土中。
JOB|16|16|我的臉因哭泣變紅， 我的眼皮上有死蔭。
JOB|16|17|我的手中卻沒有暴力， 我的祈禱也是純潔的。
JOB|16|18|「地啊，不要遮蓋我的血！ 不要讓我的哀求有藏匿之處！
JOB|16|19|現今，看哪，在天有我的見證， 在上有我的保人。
JOB|16|20|我的朋友譏誚我， 我卻向上帝眼淚汪汪。
JOB|16|21|願人可與上帝理論， 如同人與朋友一樣；
JOB|16|22|因為再過幾年， 我必走那往而不返之路。」
JOB|17|1|「我的靈耗盡，我的日子消逝； 墳墓為我預備好了。
JOB|17|2|戲笑的人果真陪伴著我， 我的眼睛盯住他們的悖逆。
JOB|17|3|「願你親自為我付押擔保。 誰還會與我擊掌呢？
JOB|17|4|因你蒙蔽他們的心，使不明理， 所以你必不高舉他們。
JOB|17|5|控告 朋友為了分享產業的， 他兒女的眼睛要失明。
JOB|17|6|「上帝使我成為人群中的笑談， 他們吐唾沫在我臉上。
JOB|17|7|我的眼睛因憂愁昏花， 我的肢體全像影兒。
JOB|17|8|正直人因此必驚奇； 無辜的人要興起攻擊不敬虔之輩。
JOB|17|9|然而，義人要持守所行的道， 手潔的人要力上加力。
JOB|17|10|至於你們眾人，再回來吧！ 你們中間，我找不到一個智慧人。
JOB|17|11|我的日子已經過去了， 我的謀算、我心的願望已經斷絕了。
JOB|17|12|他們以黑夜為白晝， 即使面臨黑暗，以為亮光已近。
JOB|17|13|我若盼望陰間為我的家， 若下榻在黑暗中，
JOB|17|14|若對地府呼叫：『你是我的父親』， 若對蟲呼叫：『你是我的母親、姊妹』，
JOB|17|15|這樣，我的盼望在哪裏呢？ 我所盼望的，誰能看見呢？
JOB|17|16|這盼望要下到陰間的門閂嗎 ？ 要一起在塵土中安息嗎 ？」
JOB|18|1|書亞 人 比勒達 回答說：
JOB|18|2|「你們尋索言語要到幾時呢 ？ 你們要明白，然後我們才說話。
JOB|18|3|我們為何被視為畜生， 在你們眼中看為愚笨 呢？
JOB|18|4|在怒氣中將自己撕裂的人哪， 難道大地要因你見棄、 磐石要挪開原處嗎？
JOB|18|5|「惡人的亮光必要熄滅， 他的火焰必不照耀。
JOB|18|6|他帳棚中的亮光要變黑暗， 他上面的燈也必熄滅。
JOB|18|7|他強橫的腳步必遭阻礙， 他的計謀必將自己絆倒。
JOB|18|8|他因自己的腳陷入網中， 走在纏人的網子上。
JOB|18|9|羅網必抓住他的腳跟， 陷阱必擒獲他。
JOB|18|10|繩索為他藏在土裏， 羈絆為他藏在路上。
JOB|18|11|四面的驚嚇使他害怕， 在他腳跟後面追趕他。
JOB|18|12|他的力量必因飢餓衰敗， 禍患要在他的旁邊等候，
JOB|18|13|侵蝕他肢體的皮膚； 死亡的長子吞吃他的肢體。
JOB|18|14|他要從所倚靠的帳棚被拔出來， 帶到使人驚恐的王那裏。
JOB|18|15|不屬他的必住在他的帳棚裏， 硫磺必撒在他所住之處。
JOB|18|16|下邊，他的根要枯乾； 上邊，他的枝子要剪除。
JOB|18|17|他的稱號 從地上消失， 他的名字不在街上存留。
JOB|18|18|他必從光明中被驅逐到黑暗裏， 他必被趕出世界。
JOB|18|19|他在自己百姓中必無子無孫， 在寄居之地也沒有倖存者。
JOB|18|20|以後的人 要因他的日子驚訝， 以前的人 也被驚駭抓住。
JOB|18|21|不義之人的住處總是這樣， 這就是不認識上帝之人的下場。」
JOB|19|1|約伯 回答說：
JOB|19|2|「你們攪擾我的心， 用言語壓碎我要到幾時呢？
JOB|19|3|你們這十次羞辱我， 苦待我也不以為恥。
JOB|19|4|果真我有錯， 這錯是在於我。
JOB|19|5|若你們真要向我誇大， 以我的羞辱來責備我，
JOB|19|6|就該知道是上帝傾覆我， 用羅網圍繞我。
JOB|19|7|看哪，我喊冤叫屈，卻不蒙應允； 我呼求，卻沒有公正。
JOB|19|8|上帝攔住我的道路，使我不得經過； 他使黑暗籠罩我的路徑。
JOB|19|9|他剝去我的榮光， 摘去我頭上的冠冕。
JOB|19|10|他在四圍攻擊我，我就走了； 他將我的指望如樹拔出。
JOB|19|11|他向我發烈怒， 以我為他的敵人。
JOB|19|12|他的軍隊一齊上來， 修築道路攻擊我， 在我帳棚的四圍安營。
JOB|19|13|「他把我的兄弟隔在遠處， 使我認識的人全然與我生疏。
JOB|19|14|我的親戚都離開了我； 我的密友都忘記了我。
JOB|19|15|在我家寄居的和我的使女， 都當我是陌生人； 我在他們眼中被視為外邦人。
JOB|19|16|我呼喚僕人，他卻不回答； 我必須親口求他。
JOB|19|17|我口的氣味令我妻子厭惡， 我的同胞都憎惡我。
JOB|19|18|連小男孩也藐視我； 我起來，他們都嘲笑我。
JOB|19|19|我的知心朋友都憎惡我； 我平日所愛的人向我翻臉。
JOB|19|20|我的皮和肉緊貼骨頭， 我得以逃脫，僅剩牙齒 。
JOB|19|21|我的朋友啊，可憐我！可憐我！ 因為上帝的手攻擊我。
JOB|19|22|你們為甚麼彷彿上帝逼迫我， 吃我的肉還不滿足呢？
JOB|19|23|「惟願我的言語現在就寫上， 都記錄在書上；
JOB|19|24|用鐵筆和鉛， 刻在磐石上，存到永遠。
JOB|19|25|我知道我的救贖主 活著， 末後他必站在塵土上。
JOB|19|26|我這皮肉滅絕之後 ， 我必在肉體之外 得見上帝。
JOB|19|27|我自己要見他， 親眼要看他，並不像陌生人。 我的心腸在我裏面耗盡了！
JOB|19|28|你們若說：『我們怎麼逼迫他呢？ 事情的根源是在於他 』，
JOB|19|29|你們就當懼怕刀劍， 因為憤怒帶來刀劍的刑罰。 這樣，你們就知道有審判。」
JOB|20|1|拿瑪 人 瑣法 回答說：
JOB|20|2|「這樣，我的思念叫我回答， 因為我心中急躁。
JOB|20|3|我聽見那羞辱我的責備； 我悟性的靈回答我。
JOB|20|4|你豈不知道嗎？亙古以來， 自從人被安置在地，
JOB|20|5|惡人歡樂的聲音是暫時的， 不敬虔人的喜樂不過是轉眼之間。
JOB|20|6|他的尊榮雖達到天上， 頭雖頂到雲中，
JOB|20|7|他必永遠滅亡，像自己的糞一樣。 看見他的人要說：『他在哪裏呢？』
JOB|20|8|他必如夢飛去，不再尋見； 他被趕走，如夜間的異象。
JOB|20|9|親眼見過他的，必不再見他； 他自己的地方也不再見到他。
JOB|20|10|他的兒女要向窮人求恩； 他的手要賠還錢財。
JOB|20|11|他的骨頭雖然滿有年輕的活力， 卻要和他一同躺臥在塵土之中。
JOB|20|12|「他口中以惡為甘甜， 把惡藏在舌頭底下，
JOB|20|13|愛戀不捨， 含在口中。
JOB|20|14|他的食物在肚裏卻要翻轉， 在他裏面成為虺蛇的毒液。
JOB|20|15|他吞了財寶，還要吐出； 上帝要從他腹中掏出來。
JOB|20|16|他必吸飲虺蛇的毒汁， 毒蛇的舌頭必殺他。
JOB|20|17|他不再看見溪流， 流奶與蜜之河。
JOB|20|18|他勞碌得來的要賠還，不得吞下； 賺取了財貨，也不得歡樂。
JOB|20|19|他欺壓窮人，棄之不顧， 強取非自己所蓋的房屋 。
JOB|20|20|「他的肚腹不知安逸， 所貪戀的連一樣也不放過，
JOB|20|21|剩餘的沒有一樣他不吞吃， 所以他的福樂不能長久。
JOB|20|22|他在滿足有餘的時候，必有困苦臨到； 凡受苦楚之人的手必加在他身上。
JOB|20|23|他的肚腹正要滿足的時候， 上帝必將猛烈的憤怒降在他身上； 他正在吃飯的時候， 上帝要將這憤怒如雨降在他身上。
JOB|20|24|他要躲避鐵的武器， 銅弓要將他射透。
JOB|20|25|箭一抽，就從他背上出來， 發亮的箭頭從他膽中出來； 有驚惶臨到他身上。
JOB|20|26|他的財寶隱藏在深沉的黑暗裏； 有非人吹起的火要把他吞滅， 把他帳棚中所剩下的燒燬。
JOB|20|27|天要顯明他的罪孽， 地要興起去攻擊他。
JOB|20|28|他家裏出產的必消失， 在上帝憤怒的日子被沖走。
JOB|20|29|這是惡人從上帝所得的份， 是上帝為他所定的產業。」
JOB|21|1|約伯 回答說：
JOB|21|2|「你們要細心聽我的言語， 這就算是你們的安慰。
JOB|21|3|請寬容我，我又要說話； 說了以後，任憑你嗤笑吧！
JOB|21|4|我豈是向人訴苦？ 我為何不是沒有耐心呢？
JOB|21|5|你們要轉向我而驚奇， 要用手摀口。
JOB|21|6|我每逢思想，心就驚惶， 戰兢抓住我身。
JOB|21|7|惡人為何存活， 得享高壽，勢力強盛呢？
JOB|21|8|他們的後裔與他們一起 ，堅立在他們面前， 他們得以眼見自己的子孫。
JOB|21|9|他們的家宅平安無懼， 上帝的杖不加在他們身上。
JOB|21|10|他們的公牛傳種而不斷絕， 母牛生牛犢而不掉胎。
JOB|21|11|他們打發小男孩出去，多如羊群， 他們的孩子踴躍跳舞。
JOB|21|12|他們隨著琴鼓歌唱， 因簫聲歡喜。
JOB|21|13|他們度日諸事亨通， 在平安中下到陰間。
JOB|21|14|他們對上帝說：『離開我們吧！ 我們不想知道你的道路。
JOB|21|15|全能者是誰，我們何必事奉他呢？ 求告他有甚麼益處呢？』
JOB|21|16|看哪，他們亨通不是靠自己的手； 惡人的計謀離我好遠。
JOB|21|17|「惡人的燈何嘗熄滅？ 患難何嘗臨到他們呢？ 上帝何嘗發怒，把災禍分給他們呢？
JOB|21|18|他們何嘗像風前的碎秸， 如暴風颳去的糠秕呢？
JOB|21|19|上帝為惡人的兒女積蓄罪孽， 不如本人遭報，好使他親自知道。
JOB|21|20|願他親眼看見自己敗亡， 親自飲全能者的憤怒。
JOB|21|21|他的歲月既盡， 他身後還顧他的家嗎？
JOB|21|22|誰能將知識教導上帝呢？ 是他審判那些居高位的。
JOB|21|23|有人至死身體強壯， 盡得平順安逸；
JOB|21|24|他的肚腹充滿奶汁 ， 他的骨髓滋潤。
JOB|21|25|有人至死心中痛苦， 從未嘗過福樂的滋味；
JOB|21|26|他們同樣躺臥於塵土， 蟲子覆蓋他們。
JOB|21|27|「看哪，我知道你們的意念， 並殘害我的計謀。
JOB|21|28|你們說：『權貴的房屋在哪裏？ 惡人住過的帳棚在哪裏？』
JOB|21|29|你們沒有詢問那些過路的人嗎？ 你們不承認他們的證據嗎？
JOB|21|30|就是惡人在患難的日子得存留， 在憤怒的日子得逃脫。
JOB|21|31|他所行的，有誰當面給他說明？ 他所做的，有誰報應他呢？
JOB|21|32|然而他要被抬到墳地， 並有人看守墓穴。
JOB|21|33|他要以谷中的土塊為甘甜； 人人要跟在他後面， 在他前面去的無數。
JOB|21|34|你們怎能以空話安慰我呢？ 你們的對答全都錯謬！」
JOB|22|1|提幔 人 以利法 回答說：
JOB|22|2|「人能使上帝有益嗎？ 智慧人能使他有益嗎？
JOB|22|3|你為人公義，豈能叫全能者喜悅呢？ 你行為完全，豈能使他得利呢？
JOB|22|4|他豈是因你敬畏的心就責備你， 審判你嗎？
JOB|22|5|你的罪惡豈不是大嗎？ 你的罪孽不是沒有窮盡嗎？
JOB|22|6|因你無故強取弟兄的抵押， 剝去赤身者的衣服。
JOB|22|7|疲乏的人，你沒有給他水喝； 飢餓的人，你沒有給他食物。
JOB|22|8|有能力的人得土地； 尊貴的人住在其中。
JOB|22|9|你打發寡婦空手回去， 你折斷孤兒的膀臂。
JOB|22|10|因此，有羅網環繞你， 有恐懼忽然使你驚惶；
JOB|22|11|或有黑暗使你看不見 ， 有洪水淹沒你。
JOB|22|12|「上帝豈不是在高天嗎？ 你看星宿的頂點何其高呢！
JOB|22|13|你說：『上帝知道甚麼？ 他豈能透過幽暗施行審判呢？
JOB|22|14|密雲將他遮蓋，使他不能看見； 他周遊穹蒼。』
JOB|22|15|你要依從上古的道嗎？ 這道是惡人行過的。
JOB|22|16|他們未到時候就被抓去 ； 他們的根基被江河沖去。
JOB|22|17|他們向上帝說：『離開我們吧！』 全能者能把他們怎麼樣呢？
JOB|22|18|然而，是上帝以美物充滿他們的房屋； 惡人的計謀離我好遠！
JOB|22|19|義人看見他們的結局 就歡喜； 無辜的人嗤笑他們：
JOB|22|20|『攻擊我們的果然被剪除， 剩餘的都被火吞滅。』
JOB|22|21|「你要與上帝和好，要和平， 這樣，福氣必臨到你。
JOB|22|22|你當領受他口中的教導， 將他的言語存在心裏。
JOB|22|23|你若歸向全能者，就必得建立。 你要從你帳棚中遠離不義，
JOB|22|24|你要將黃金丟到塵土裏， 將 俄斐 的金子丟在溪河石頭之間；
JOB|22|25|全能者就必作你的黃金， 作你成堆的銀子。
JOB|22|26|那時，你要以全能者為喜樂， 向上帝仰臉。
JOB|22|27|你要向他禱告，他就聽你； 你也要還你的願。
JOB|22|28|你定意要做何事，必然為你成就； 亮光也必照耀你的路。
JOB|22|29|當人降卑，你說：是因驕傲； 眼目謙卑的人，上帝必然拯救。
JOB|22|30|不是無辜的人，上帝尚且要搭救他 ； 他必因你手中的清潔得蒙拯救。」
JOB|23|1|約伯 回答說：
JOB|23|2|「如今我的哀告還算為悖逆； 我雖唉哼，他的手仍然重重責罰我 。
JOB|23|3|惟願我知道哪裏可以尋見上帝， 能到他的臺前，
JOB|23|4|我就在他面前陳明我的案件， 滿口辯訴。
JOB|23|5|我必知道他回答我的言語， 明白他向我所要說的。
JOB|23|6|他豈用大能與我爭辯呢？ 不！他必理會我。
JOB|23|7|在那裏正直人可以與他辯論， 我就必永遠脫離那審判我的。
JOB|23|8|「看哪，我往前走，他不在那裏； 往後退，也沒有察覺他。
JOB|23|9|他在左邊行事，我卻看不見他； 他轉向右邊 ，我也見不到他。
JOB|23|10|然而他知道我所走的路； 他試煉我，我就如純金。
JOB|23|11|我的腳緊跟他的步伐； 我謹守他的道，並不偏離。
JOB|23|12|他嘴唇的命令，我未曾背棄； 我看重他口中的言語，過於我需用的飲食 。
JOB|23|13|只是他心志已定，誰能使他轉意呢？ 他心裏所願的，就行出來。
JOB|23|14|因此，為我所定的，他必做成， 這類的事他還有許多。
JOB|23|15|所以我在他面前驚惶； 我思想就懼怕他。
JOB|23|16|上帝使我喪膽， 全能者使我驚惶。
JOB|23|17|但我並非被黑暗剪除， 只是幽暗遮蓋了我的臉。
JOB|24|1|「為何全能者不定下期限？ 為何認識他的人看不到那些日子呢？
JOB|24|2|有人挪移地界， 搶奪群畜去放牧。
JOB|24|3|他們拉走孤兒的驢， 強取寡婦的牛作抵押。
JOB|24|4|他們使貧窮人離開正道； 世上的困苦人盡都隱藏。
JOB|24|5|看哪，他們如同野驢出到曠野，殷勤尋找食物， 在野地給孩童餬口。
JOB|24|6|他們收割別人田間的莊稼， 摘取惡人剩餘的葡萄。
JOB|24|7|他們終夜赤身無衣， 在寒冷中毫無遮蓋。
JOB|24|8|他們在山上被大雨淋濕， 因沒有避身之處就擁抱磐石。
JOB|24|9|又有人從母懷中搶走孤兒， 在困苦人身上強取抵押品 。
JOB|24|10|困苦人赤身無衣，到處流浪， 餓著肚子扛抬禾捆，
JOB|24|11|他們在圍牆內榨油， 踹壓酒池，自己卻口渴。
JOB|24|12|在城內垂死的人呻吟， 受傷的人哀號； 上帝卻不理會狂妄的事。
JOB|24|13|「又有人背棄光明， 不認識光明的道， 不留在光明的路上。
JOB|24|14|殺人者黎明起來， 殺害困苦人和貧窮人， 夜間又作盜賊。
JOB|24|15|姦夫的眼等候黃昏， 說：『沒有眼睛能見我』， 就把臉蒙住。
JOB|24|16|盜賊黑夜挖洞； 他們白日躲藏， 並不認識光明。
JOB|24|17|他們全都看早晨如死蔭， 因為他們熟悉死蔭的驚駭。
JOB|24|18|「惡人在水面上快速飄盪， 他們在地上所得的產業被詛咒； 無人再回到他們的葡萄園。
JOB|24|19|乾旱炎熱融化雪水； 陰間也如此吞沒犯罪的人。
JOB|24|20|懷他的母胎忘記他； 蟲子要吃他，覺得甘甜； 他不再被人記念； 不義的人必如樹折斷。
JOB|24|21|「他與不懷孕不生育的婦人交往 ， 卻不善待寡婦。
JOB|24|22|然而上帝用能力保全有勢力的人； 那性命難保的人仍然興起。
JOB|24|23|上帝使他安穩，他就有所倚靠； 上帝的眼目看顧他們的道路。
JOB|24|24|他們高升，不過片刻就沒有了； 他們降為卑，被除滅，與眾人一樣 ， 又如穀的穗子被割下。
JOB|24|25|若不是這樣，誰能指證我是說謊的， 以我的言語為毫無根據呢？」
JOB|25|1|書亞 人 比勒達 回答說：
JOB|25|2|「上帝有統治之權，威嚴可畏； 他在高處施行和平。
JOB|25|3|他的軍隊豈能數算？ 他的光向誰不會升起呢 ？
JOB|25|4|這樣，在上帝面前人怎能稱義？ 婦人所生的怎能潔淨？
JOB|25|5|看哪，在上帝眼前，月亮無光， 星宿也不皎潔，
JOB|25|6|更何況是如蟲的人， 如蛆的世人呢！
JOB|26|1|約伯 回答說：
JOB|26|2|「無能的人蒙你何等的幫助！ 膀臂無力的人蒙你何等的拯救！
JOB|26|3|無智慧的人蒙你何等的指教！ 你向他顯出豐富的知識。
JOB|26|4|你向誰發出言語？ 誰的靈從你而出？
JOB|26|5|在大水和水族以下， 陰魂戰兢。
JOB|26|6|在上帝面前，陰間顯露； 冥府 也不得遮掩。
JOB|26|7|上帝將北極鋪在空中， 將大地懸在虛空。
JOB|26|8|他將水包在密雲中， 盛水的雲卻不破裂。
JOB|26|9|他遮蔽寶座的正面， 把他的雲彩鋪在其上。
JOB|26|10|他在水面上劃一圓圈， 直到光明與黑暗的交界。
JOB|26|11|天的柱子震動， 因他的斥責驚奇。
JOB|26|12|他以能力攪動 大海 ， 藉知識打傷 拉哈伯 。
JOB|26|13|他藉自己的靈使天空晴朗； 他的手刺殺爬得快的蛇。
JOB|26|14|看哪，這不過是上帝工作的些微； 我們聽見他的話，是何等細微的聲音！ 他大能的雷聲誰能明白呢？」
JOB|27|1|約伯 繼續發表他的言論說：
JOB|27|2|「我指著奪去我公道的永生上帝， 並使我心中愁苦的全能者起誓：
JOB|27|3|只要我的生命尚在我裏面， 上帝所賜的氣息仍在我鼻孔內，
JOB|27|4|我的唇絕不說不義， 我的舌也不說詭詐。
JOB|27|5|我斷不以你們為義； 我至死不放棄自己的純正！
JOB|27|6|我持定我的義，並不放鬆； 在世的日子，我的心不責備我。
JOB|27|7|「願我的仇敵如惡人一樣； 願那起來攻擊我的，如不義之人一般。
JOB|27|8|不敬虔的人有甚麼指望呢？ 上帝要剪除他，取他的性命。
JOB|27|9|患難臨到他， 上帝豈聽他的呼求？
JOB|27|10|他豈以全能者為樂， 隨時求告上帝呢？
JOB|27|11|上帝手所做的，我要指教你們； 全能者所行的，我也不會隱瞞。
JOB|27|12|看哪，你們自己也都見過， 為何全變為這樣虛妄呢？
JOB|27|13|「這是上帝為惡人所定的份， 殘暴人從全能者所得的產業：
JOB|27|14|倘若他的兒女增多，仍被刀所殺； 他的子孫必不得飽食。
JOB|27|15|他遺留的人必死而埋葬， 他的寡婦也不哀哭。
JOB|27|16|他雖積蓄銀子如塵沙， 堆積衣服如泥土，
JOB|27|17|他儘管堆積，義人卻要穿上， 無辜的人卻要分取銀子。
JOB|27|18|他建造房屋如蟲做窩， 又如守望者所搭的棚。
JOB|27|19|他雖富足躺臥，卻不得收殮 ， 他張開眼睛，就不在了。
JOB|27|20|驚恐如洪水將他追上， 暴風在夜間將他颳去。
JOB|27|21|東風把他吹去，他就走了； 風將他颳離原地。
JOB|27|22|風 無情地擊打他， 他試圖逃脫風的手。
JOB|27|23|風要因他拍掌， 並要發叱聲，使他離開原地。」
JOB|28|1|「銀子有礦； 煉金有場。
JOB|28|2|鐵從土裏開採， 銅從礦石鎔出。
JOB|28|3|人探索黑暗的盡頭， 查究礦石直到極處， 那是幽暗和死蔭；
JOB|28|4|他在無人居住之處開鑿礦穴， 在無足跡之地被遺忘 ， 與人遠離，懸空搖擺。
JOB|28|5|地出產糧食， 地底翻騰如火。
JOB|28|6|地的石頭是藍寶石之處， 那裏還有金沙。
JOB|28|7|鷙鳥不知那條路， 鷹眼也未曾見過。
JOB|28|8|狂傲的野獸未曾踩踏， 猛烈的獅子也未曾經過。
JOB|28|9|「人動手鑿開堅石， 翻倒山的根基，
JOB|28|10|在磐石中鑿出水道， 親眼看見各樣寶物。
JOB|28|11|他封閉河川不得涓滴 ， 使隱藏之物顯露出來。
JOB|28|12|「然而，智慧何處可尋？ 聰明之地在哪裏？
JOB|28|13|智慧的價值 無人能知， 活人之地也無處可尋。
JOB|28|14|深淵說：『不在我裏面。』 滄海說：『不在我這裏。』
JOB|28|15|智慧不可用黃金換取， 也不能用白銀秤她的價值。
JOB|28|16|俄斐 的金子和貴重的紅瑪瑙， 以及藍寶石，不足與她比擬；
JOB|28|17|黃金和玻璃不足與她比較； 純金的器皿不足兌換她。
JOB|28|18|珊瑚、水晶都不值得提； 智慧的價值勝過寶石 。
JOB|28|19|古實 的紅璧璽不足與她比較； 純金也不足與她比擬。
JOB|28|20|「智慧從何處來呢？ 聰明之地在哪裏？
JOB|28|21|她隱藏，遠離眾生的眼目， 她掩蔽，遠離空中的飛鳥。
JOB|28|22|毀滅和死亡說： 『我們風聞其名。』
JOB|28|23|「上帝明白智慧的道路， 知道智慧的所在。
JOB|28|24|因為他鑒察直到地極， 遍觀普天之下，
JOB|28|25|要為風定輕重， 又度量諸水，
JOB|28|26|為雨定律例， 為雷電定道路。
JOB|28|27|那時他看見智慧，就談論她， 堅定她，並且查究她。
JOB|28|28|他對人說：『看哪，敬畏主就是智慧； 遠離惡事就是聰明。』」
JOB|29|1|約伯 繼續發表他的言論說：
JOB|29|2|「惟願我如從前的歲月， 如上帝保護我的日子。
JOB|29|3|那時他的燈照在我頭上， 我藉他的光行過黑暗。
JOB|29|4|在我壯年的時候， 上帝親密的情誼臨到我的帳棚中。
JOB|29|5|全能者仍與我同在， 我的兒女都環繞我。
JOB|29|6|我的腳洗在乳酪當中； 磐石為我流出油河。
JOB|29|7|我出到城門， 在廣場安排座位，
JOB|29|8|年輕人見我而迴避， 老年人起身站立。
JOB|29|9|王子都停止說話， 用手摀口；
JOB|29|10|領袖靜默無聲， 舌頭貼住上膛。
JOB|29|11|耳朵聽見了，稱我有福； 眼睛看見了，就稱讚我。
JOB|29|12|因我拯救了哀求的困苦人 和無人幫助的孤兒。
JOB|29|13|將要滅亡的為我祝福， 我使寡婦心中歡呼。
JOB|29|14|我穿上公義，它遮蔽我； 我的公平如外袍和冠冕。
JOB|29|15|我作瞎子的眼， 瘸子的腳。
JOB|29|16|我作貧窮人的父； 我不認識之人的案件，我也去查明。
JOB|29|17|我打破不義之人的大牙， 從他牙齒中奪走他所搶的。
JOB|29|18|我說：『我要增添我的日子如塵沙， 我必死在自己家中 。
JOB|29|19|我的根伸展到水邊， 露水夜宿我的枝上。
JOB|29|20|我的榮耀在我身上更新， 我的弓在我手中日新。』
JOB|29|21|「人聽我說話而等候， 為我的教導而靜默。
JOB|29|22|我說話之後，他們就不再說； 我的言語滴在他們身上。
JOB|29|23|他們等候我如等雨水， 又張口如切慕春雨。
JOB|29|24|我向他們微笑，他們不敢相信； 他們不使我臉上的光失色。
JOB|29|25|我為他們選擇道路，又坐首位； 我如君王在軍隊中居住， 又如人安慰哀傷的人。」
JOB|30|1|「但如今，比我年輕的人譏笑我； 我曾藐視他們的父親， 不放在我的牧羊犬中。
JOB|30|2|他們的精力既已衰敗， 手中的氣力於我何益？
JOB|30|3|他們因窮乏飢餓，沒有生氣， 在荒廢淒涼的幽暗中啃乾燥之地。
JOB|30|4|他們在草叢之中採鹹草， 羅騰 樹的根成為他們的食物。
JOB|30|5|他們從人群中被趕出， 人追喊他們如賊一般，
JOB|30|6|以致他們住在荒谷， 住在地洞和巖穴中。
JOB|30|7|他們在草叢中叫喚， 在荊棘下擠成一團。
JOB|30|8|這都是愚頑卑微人的兒女； 他們被鞭打，趕出境外。
JOB|30|9|「現在這些人以我為歌曲， 以我為笑談。
JOB|30|10|他們厭惡我，躲避我， 不住地吐唾沫在我臉上。
JOB|30|11|上帝鬆開我的弓弦 使我受苦， 他們就在我面前脫去轡頭。
JOB|30|12|這夥人在我右邊起來， 他們推開我的腳， 築災難之路攻擊我。
JOB|30|13|他們毀壞我的道， 加增我的災害； 他們毋須人幫助。
JOB|30|14|他們來，如同闖進大缺口， 在暴風間滾動。
JOB|30|15|驚恐傾倒在我身上， 我的尊榮被逐如風； 我的福祿如雲飄去。
JOB|30|16|「現在我的心極其悲傷， 困苦的日子將我抓住。
JOB|30|17|夜間，我裏面的骨頭刺痛， 啃著我的沒有止息。
JOB|30|18|我的外衣因大力扭皺 ， 內衣的領子把我勒住。
JOB|30|19|上帝把我扔在淤泥之中， 我就像塵土和灰燼一樣。
JOB|30|20|我呼求你，你不應允我； 我站起來，你只是望著我。
JOB|30|21|你對我變得殘忍， 大能的手追逼我。
JOB|30|22|你把我提到風中，使我乘風而去， 使我消失在烈風之中。
JOB|30|23|我知道你要使我歸於死亡， 到那為眾生所定的陰宅。
JOB|30|24|「然而，人在廢墟豈不伸手？ 遇災難時一定呼救。
JOB|30|25|人遭難的日子，我豈不為他哭泣呢？ 人貧窮的時候，我豈不為他憂愁呢？
JOB|30|26|我仰望福氣，災禍就來到； 我等待光明，黑暗便來臨。
JOB|30|27|我內心煩擾不安， 困苦的日子臨到我身。
JOB|30|28|我在陰暗中行走，沒有日光 ， 我在會眾中站立求救。
JOB|30|29|我與野狗為弟兄， 我跟鴕鳥為同伴。
JOB|30|30|我的皮膚變黑脫落， 我的骨頭因熱燒焦。
JOB|30|31|我的琴音變為哀泣； 我的簫聲變為哭聲。」
JOB|31|1|「我與眼睛立約， 怎能凝望少女呢？
JOB|31|2|從至上的上帝所得之分， 從至高全能者所得之業是甚麼呢？
JOB|31|3|豈不是禍患臨到不義的， 災害臨到作惡的嗎？
JOB|31|4|上帝豈不察看我的道路， 數點我所有的腳步嗎？
JOB|31|5|「我若與虛謊同行， 我腳若緊跟詭詐，
JOB|31|6|願上帝用公道的天平秤我， 願他知道我的純正。
JOB|31|7|我的腳步若偏離正路， 我的心若隨從我眼目， 我的手掌若黏有污穢；
JOB|31|8|願我栽種，別人來吃， 我的農作物連根拔出。
JOB|31|9|「我心若因婦人受迷惑， 在鄰舍的門外等候，
JOB|31|10|就願我妻子給別人推磨， 別人與她同寢。
JOB|31|11|因為這是邪惡的事， 審判官裁定的罪孽。
JOB|31|12|這是一場火，直燒到毀滅 ， 必拔除我一切的家產。
JOB|31|13|「我的僕婢與我爭辯， 我若藐視不聽他們的冤情，
JOB|31|14|上帝興起的時候，我怎樣行呢？ 他察問的時候，我怎樣回答他呢？
JOB|31|15|造我在母腹中的，不也是造了他嗎？ 在母胎中使我們成形的，豈不是同一位嗎？
JOB|31|16|「我若不讓貧寒人遂其所願， 或是叫寡婦眼中失望，
JOB|31|17|或獨自吃自己的食物， 孤兒沒有吃其中些許；
JOB|31|18|從我年輕時，孤兒就與我一同長大，我好像他的父親， 我從出母腹就扶助寡婦 ；
JOB|31|19|我若見人因無衣死亡， 或見貧窮人毫無遮蓋；
JOB|31|20|我若不使他真心為我祝福， 不使他因我羊的毛得暖；
JOB|31|21|我若舉手攻擊孤兒， 因為在城門口見有幫助我的；
JOB|31|22|情願我的肩膀從肩胛骨脫落， 我的膀臂從肱骨折斷。
JOB|31|23|因上帝降的災禍使我恐懼 ， 因他的威嚴，我甚麼都不能。
JOB|31|24|「我若以黃金為我的指望， 對純金說：你是我的倚靠；
JOB|31|25|我若因財物豐裕， 因手多得資財而歡喜；
JOB|31|26|我若見太陽發光， 明月運行，
JOB|31|27|心就暗暗被引誘， 口親吻自己的手；
JOB|31|28|這也是審判官裁定的罪孽， 因為我背棄了至上的上帝。
JOB|31|29|「我若見恨我的遇難就歡喜， 見他遭災就高興；
JOB|31|30|其實我沒有容許口犯罪， 以詛咒要他的性命；
JOB|31|31|若我帳棚中的人未曾說： 『誰不以他的肉食吃飽呢？』
JOB|31|32|我未曾讓旅客在街上過夜， 卻開門迎接行路的人；
JOB|31|33|我若像 亞當 遮掩自己的過犯， 將罪孽藏在懷中；
JOB|31|34|我若因大大懼怕眾人， 又因宗族的藐視而恐懼， 以致我緘默不言，閉門不出；
JOB|31|35|惟願有一位肯聽我！ 看哪，我的記號，願全能者回答我！ 願那與我爭訟的寫下狀詞！
JOB|31|36|我必把它帶在肩上， 綁在頭上為冠冕。
JOB|31|37|我必向上帝述說我腳步的數目， 如同王子進到他面前。
JOB|31|38|「若我的田地喊冤告我， 犁溝也一同哭泣；
JOB|31|39|我若吃地的出產不給銀錢， 或叫地的原主喪命；
JOB|31|40|願蒺藜生長代替麥子， 惡臭的草代替大麥。」 約伯 的話說完了。
JOB|32|1|於是這三個人因 約伯 看自己為義就停止，不再回答他。
JOB|32|2|那時 布西 人， 蘭 族 巴拉迦 的兒子 以利戶 發怒了。他向 約伯 發怒，因 約伯 自以為義，不以上帝為義。
JOB|32|3|他又向 約伯 的三個朋友發怒，因為他們想不出回答的話來，仍以 約伯 為有罪。
JOB|32|4|以利戶 因為他們比自己年老，就等候要與 約伯 說話。
JOB|32|5|以利戶 見這三個人口中無話回答，就發怒。
JOB|32|6|布西 人 巴拉迦 的兒子 以利戶 回答說： 「我年輕，你們年長， 因此我退讓，不敢向你們陳述我的意見。
JOB|32|7|我說：『年長的當先說話； 壽高的當以智慧教導人。』
JOB|32|8|其實，是人裏面的靈， 全能者的氣使人有聰明。
JOB|32|9|壽高的不都有智慧， 年老的不都明白公平。
JOB|32|10|因此我說：『你們要聽我， 我也要陳述我的意見。』
JOB|32|11|「看哪，我等候你們的話， 側耳聽你們的高見； 直到你們找到要說的言語。
JOB|32|12|我留心聽你們， 看哪，你們中間無一人能折服 約伯 ， 回答他的話。
JOB|32|13|你們切不可說：『我們尋得智慧； 上帝能勝他 ，人卻不能。』
JOB|32|14|約伯 沒有用言語與我爭辯； 我也不用你們的話回答他。
JOB|32|15|「他們驚惶不再回答， 一言不發。
JOB|32|16|我豈因他們不說話， 因他們站住不再回答，仍舊等候呢？
JOB|32|17|我也要以我的一番話回答， 我也要陳述我的意見。
JOB|32|18|因為我滿懷言語， 我裏面的靈激動我。
JOB|32|19|看哪，我的肚腹如酒囊沒有氣孔， 又如新皮袋 快要破裂。
JOB|32|20|我要說話，使我舒暢； 我要張開嘴唇回答。
JOB|32|21|我必不看人的情面， 也不奉承人。
JOB|32|22|我不懂得奉承； 不然，造我的主必快快除滅我。」
JOB|33|1|「但是， 約伯 啊，請聽我的言語， 側耳聽我一切的話。
JOB|33|2|看哪，我開口， 我的舌在上膛發言。
JOB|33|3|我的言語要表明心中的正直， 我嘴唇所知道的就誠實地說。
JOB|33|4|上帝的靈造了我， 全能者的氣使我得生。
JOB|33|5|你若能夠，就請回答我； 請你站起來，在我面前陳明。
JOB|33|6|看哪，我在上帝面前與你一樣， 也是用泥土造成的。
JOB|33|7|看哪，我不用威嚴恐嚇你， 也不用勢力重壓你。
JOB|33|8|「其實，你向我耳朵說話， 我聽見你言語的聲音：
JOB|33|9|『我是純潔無過的， 我是無辜的，在我裏面沒有罪孽。
JOB|33|10|看哪，上帝找機會攻擊我， 以我為他的仇敵，
JOB|33|11|把我的腳鎖上木枷， 察看我一切的道路。』
JOB|33|12|「看哪，你這話無理，我要回答你， 因上帝比世人更大。
JOB|33|13|你為何與他爭論： 『他任何事都不向人解答』？
JOB|33|14|上帝說一次、兩次， 人卻不理會。
JOB|33|15|世人在床上沉睡安眠時， 在夢中和夜間的異象裏，
JOB|33|16|上帝就開通世人的耳朵， 把警告印在他們心上 ，
JOB|33|17|好叫人轉離自己的行為， 叫壯士遠離驕傲，
JOB|33|18|攔阻人不陷入地府， 不讓他命喪刀下 。
JOB|33|19|「人在床上被疼痛懲治， 骨頭不住地掙扎，
JOB|33|20|以致生命厭棄食物， 心中厭惡美味。
JOB|33|21|他的肉消瘦，難以看見； 先前看不見的骨頭都凸出來。
JOB|33|22|他的性命臨近地府， 他的生命挨近滅命者。
JOB|33|23|一千天使中， 若有一個作傳話的臨到他， 指示人所當行的事，
JOB|33|24|上帝就施恩給他，說： 『要救贖他 免得下入地府， 我已經得了贖價。
JOB|33|25|他的肉要比孩童的肉更嫩； 他就返老還童。』
JOB|33|26|他向上帝禱告，上帝就悅納他； 他必歡呼朝見上帝的面， 因上帝恢復他的義。
JOB|33|27|他在人前歌唱說： 『我犯了罪，顛倒是非， 卻沒有受該得的報應。
JOB|33|28|上帝救贖我的性命免入地府， 我的生命也必見光。』
JOB|33|29|「看哪，上帝兩次、三次 向人行這一切的事，
JOB|33|30|為要從地府救回人的性命， 使他被生命之光照耀。
JOB|33|31|約伯 啊，你當留心聽我； 不要作聲，我要說話。
JOB|33|32|你若有話說，可以回答我； 你只管說，因我願以你為義。
JOB|33|33|若不然，你當聽我； 不要作聲，我要把智慧教導你。」
JOB|34|1|以利戶 繼續說：
JOB|34|2|「你們智慧人要聽我的言語， 有知識的人要側耳聽我。
JOB|34|3|因為耳朵辨別言語， 好像上膛品嘗食物。
JOB|34|4|我們當選擇公理， 彼此知道何為善。
JOB|34|5|約伯 曾說：『我是公義的， 上帝奪去我的公理。
JOB|34|6|我有理，豈能說謊呢？ 我無過，受的箭傷卻不能醫治。』
JOB|34|7|哪一個人像 約伯 ， 喝譏誚如同喝水呢？
JOB|34|8|他與作惡的結伴， 和惡人同行。
JOB|34|9|他說：『人以上帝為樂， 總是無益。』
JOB|34|10|「所以，你們明理的人要聽我， 上帝斷不致行惡， 全能者斷不致不義。
JOB|34|11|他必按人所做的報應人， 使各人照所行的得報。
JOB|34|12|確實地，上帝必不作惡， 全能者必不偏離公平。
JOB|34|13|誰派他治理大地？ 誰安定全世界呢？
JOB|34|14|他若專心為己， 將靈和氣收歸自己，
JOB|34|15|凡血肉之軀必一同死亡； 世人必歸於塵土。
JOB|34|16|「你若明理，當聽這話， 側耳聽我言語的聲音。
JOB|34|17|難道恨惡公平的可以掌權嗎？ 那有公義、有大能的，你豈可定他有罪呢？
JOB|34|18|你會對君王說：『你是卑鄙的』； 對貴族說：『你們是邪惡的』嗎？
JOB|34|19|他待王子不徇情面， 也不看重富足的過於貧寒的， 因為他們都是他手所造的。
JOB|34|20|一瞬間他們就死亡。 百姓在半夜中被震動而去世； 有權力的被奪去，非藉人手。
JOB|34|21|「上帝的眼目觀看人的道路， 察看他每一腳步。
JOB|34|22|沒有黑暗，沒有死蔭， 能給作惡者在那裏藏身。
JOB|34|23|上帝不必再三傳人 到他面前受審判。
JOB|34|24|他毋須調查就粉碎有大能的人， 指定別人代替他們。
JOB|34|25|所以他知道他們的行為， 使他們在夜間傾倒壓碎。
JOB|34|26|他在眾目睽睽下擊打他們， 如同擊打惡人。
JOB|34|27|因為他們轉離不跟從他， 不留心他一切的道，
JOB|34|28|甚至使貧寒人的哀聲達到他那裏； 他也聽了困苦人的哀聲。
JOB|34|29|他安靜，誰能定罪呢？ 他轉臉，誰能見他呢？ 無論一國或一人都是如此。
JOB|34|30|不虔敬的人不得作王， 免得百姓陷入圈套。
JOB|34|31|「有誰對上帝說： 『我受了責罰，必不再犯罪；
JOB|34|32|我所看不明的，求你指教我； 我若行了不義，必不再行』？
JOB|34|33|他因你拒絕不接受， 就隨你的心願施行報應嗎？ 選擇的是你，不是我。 你所知道的，只管說吧！
JOB|34|34|明理的人必對我說， 聽我的智慧人也說：
JOB|34|35|『 約伯 說話沒有知識， 他的言語毫無智慧。』
JOB|34|36|願 約伯 被考驗到底， 因他回答像惡人一樣。
JOB|34|37|他在罪上又加悖逆； 在我們中間引起疑惑 ， 用許多言語輕慢上帝。」
JOB|35|1|以利戶 繼續說：
JOB|35|2|「你以為這話有理， 說：『我在上帝面前是公義的。』
JOB|35|3|你說：『這對你有甚麼益處？ 我不犯罪有甚麼好處呢？』
JOB|35|4|至於我，我要用言語回答你 和跟你一起的朋友。
JOB|35|5|你要向天觀看， 瞻望那高於你的穹蒼。
JOB|35|6|你若犯罪，能使上帝受何害呢？ 你的過犯加增，能使上帝受何損呢？
JOB|35|7|你若是公義，能加增他甚麼呢？ 他從你手裏還接受甚麼呢？
JOB|35|8|你的罪惡只影響像你這類的人； 你的公義也只影響世人。
JOB|35|9|「人因多受欺壓就哀求， 因強權者的膀臂而求救。
JOB|35|10|但無人說：『造我的上帝在哪裏？ 他使人夜間歌唱，
JOB|35|11|教導我們多過地上的走獸， 使我們比空中的飛鳥更聰明。』
JOB|35|12|因為惡人驕傲， 他們在那裏呼求，他卻不回答。
JOB|35|13|虛妄的呼求，上帝必不垂聽； 全能者必不留意。
JOB|35|14|何況你說，你不得見他。 案件就在他面前，你等候他吧。
JOB|35|15|但如今因他未曾發怒降罰， 也一點都不理會狂傲，
JOB|35|16|所以 約伯 開口說虛妄的話， 多多發表無知識的言語。」
JOB|36|1|以利戶 繼續說：
JOB|36|2|「你再給我片時，我就指示你， 因我還有話要為上帝說。
JOB|36|3|我要把我的知識從遠處引來， 我要將公義歸給造我的主。
JOB|36|4|我的言語絕不虛假， 有全備知識的與你同在。
JOB|36|5|「看哪，上帝有大能，並不藐視人； 他的心智能力廣大。
JOB|36|6|他不讓惡人活著， 卻為困苦人伸冤。
JOB|36|7|他的眼目不遠離義人， 卻使他們和君王同坐寶座， 永遠被高舉 。
JOB|36|8|他們若被鎖鏈捆住， 被苦難的繩索纏住，
JOB|36|9|他就向他們指示他們的作為和過犯， 以及他們的狂妄自大。
JOB|36|10|他也開通他們的耳朵來領受教導， 吩咐他們回轉離開罪孽。
JOB|36|11|他們若聽從事奉他， 就必度日亨通， 歷年享福。
JOB|36|12|他們若不聽從，就要被刀殺滅， 無知無識而死。
JOB|36|13|「那心中不敬虔的人積蓄怒氣； 上帝捆綁他們，他們竟不求救。
JOB|36|14|他們必在青年時死亡， 與神廟娼妓一樣喪命。
JOB|36|15|上帝藉著困苦救拔困苦人， 藉所受的欺壓開通他們的耳朵。
JOB|36|16|上帝也必引你脫離患難， 進入寬闊不狹窄之地； 擺在你席上的必滿有肥甘。
JOB|36|17|「但你充滿著惡人的辯辭， 辯辭和審判抓住你。
JOB|36|18|不可讓憤怒觸動你，使你破口謾罵 ； 也不可因贖價大而偏行。
JOB|36|19|你的呼求 和一切的勢力， 果真有用，使你不遭患難嗎？
JOB|36|20|不要切慕黑夜， 就是眾民在本處被除滅的時候。
JOB|36|21|你要謹慎，不可偏向罪孽， 因你選擇罪孽過於苦難。
JOB|36|22|看哪，上帝因他的能力而崇高； 有誰像他那樣作教師呢？
JOB|36|23|誰派定他的道路呢？ 誰能說：『你行了不義』？
JOB|36|24|「你要記得頌讚他的作為， 就是人所歌頌的。
JOB|36|25|他的作為，萬人都看見； 世人也從遠處觀看。
JOB|36|26|看哪，上帝崇高，我們不能知道； 他的年數，不能測度。
JOB|36|27|因他吸取水點， 水點就從雲霧中變成雨；
JOB|36|28|雲彩將雨落下， 沛然降於世人。
JOB|36|29|又有誰能明白密雲如何鋪張， 和上帝行宮的雷聲呢？
JOB|36|30|看哪，他的亮光普照自己的四圍； 他覆蓋海的深處。
JOB|36|31|因他用這些審判 眾民， 又賜豐富的糧食。
JOB|36|32|他以閃電遮手掌， 命令它擊中靶子。
JOB|36|33|所發的雷聲將他顯明， 牲畜也指明要起暴風 。」
JOB|37|1|「因此我心戰兢， 從原處移動。
JOB|37|2|聽啊，聽他轟轟的聲音， 是上帝口中所發的響聲。
JOB|37|3|他發響聲震遍天下， 他的閃電直到地極。
JOB|37|4|隨後，人聽見他的聲音， 是那轟轟的聲音； 他發出威嚴的雷聲， 而不加以遏止。
JOB|37|5|上帝發出奇妙的雷聲； 他行大事，我們不能測透。
JOB|37|6|他對雪說：『要降在地上』； 對大雨和暴雨也是這樣說。
JOB|37|7|他封住各人的手， 叫所造的萬人都知道他的作為。
JOB|37|8|野獸進入穴中， 臥在自己洞內。
JOB|37|9|暴風來自內宮， 寒冷出於狂風。
JOB|37|10|上帝噓氣成冰， 凝結寬闊之水，
JOB|37|11|使密雲盛滿水氣， 烏雲散佈閃電。
JOB|37|12|雲藉著他的指引遊行旋轉， 在世界的地面上行他一切所吩咐的，
JOB|37|13|或為責罰，或為他的地， 或為慈愛，都是他所行的。
JOB|37|14|「 約伯 啊，側耳聽這話， 要站立，思想上帝奇妙的作為。
JOB|37|15|你知道上帝如何安排這些， 如何使雲中的閃電照耀嗎？
JOB|37|16|你知道雲彩如何浮於空中， 知識全備者奇妙的作為嗎？
JOB|37|17|你知道南風使地寂靜， 你的衣服就變為熱嗎？
JOB|37|18|你豈能與上帝同鋪穹蒼， 堅固如同鑄成的鏡子嗎？
JOB|37|19|我們因在黑暗中，不會陳說， 請你指教我們該對他說甚麼。
JOB|37|20|有人告訴他我要說話嗎？ 豈有人說他願被吞滅嗎？
JOB|37|21|「現在，人不得見穹蒼的亮光； 風一吹過，天色晴朗。
JOB|37|22|金色的光輝來自北方， 在上帝那裏有可畏的威嚴。
JOB|37|23|全能者，我們不能測度； 他大有能力，又有公平， 滿有公義，必不苦待人。
JOB|37|24|所以，世人敬畏他； 凡自以為 有智慧的，他都不看顧。」
JOB|38|1|那時，耶和華從旋風中回答 約伯 說：
JOB|38|2|「誰用無知的言語使我的旨意暗昧不明？
JOB|38|3|你要如勇士束腰； 我問你，你可以讓我知道。
JOB|38|4|「我立大地根基的時候，你在哪裏？ 你若明白事理，只管說吧！
JOB|38|5|你知道是誰定地的尺度， 是誰把準繩拉在其上嗎？
JOB|38|6|地的根基安置在何處？ 地的角石是誰安放的？
JOB|38|7|那時，晨星一同歌唱； 上帝的眾使者也都歡呼。
JOB|38|8|「當海水衝出，如出母胎， 誰用門將它關閉呢？
JOB|38|9|是我用雲彩當海的衣服， 用幽暗當包裹它的布，
JOB|38|10|為它定界限， 又安門和閂，
JOB|38|11|說：『你只可到這裏，不可越過； 你狂傲的浪要到此止住。』
JOB|38|12|「你有生以來，曾命定晨光， 曾使黎明知道自己的地位，
JOB|38|13|抓住地的四極， 把惡人從其中驅逐出來嗎？
JOB|38|14|地改變如泥上蓋印， 萬物出現如衣服一樣。
JOB|38|15|亮光不照惡人， 高舉的膀臂也必折斷。
JOB|38|16|「你曾進到海之源， 或在深淵的隱密處行走嗎？
JOB|38|17|死亡的門曾向你顯露嗎？ 死蔭的門你曾見過嗎？
JOB|38|18|地的廣大，你能測透嗎？ 你若全知道，只管說吧！
JOB|38|19|「往光明居所的路在哪裏？ 黑暗的地方在何處？
JOB|38|20|你能將它帶到其領域， 能辨明其居所之路嗎？
JOB|38|21|你知道的，因為那時你已出生， 你活的日子數目也多。
JOB|38|22|「你曾進入雪之庫， 或見過雹的倉嗎？
JOB|38|23|雪雹是我為災難的時候， 為打仗和戰爭的日子所預備。
JOB|38|24|光亮從何路分開？ 東風從何路分散遍地？
JOB|38|25|「誰為大雨分道， 誰為雷電開路，
JOB|38|26|使雨降在無人之地， 在無人居住的曠野，
JOB|38|27|使荒廢淒涼之地得以豐足， 青草得以生長？
JOB|38|28|「雨有父親嗎？ 露珠是誰生的呢？
JOB|38|29|冰出於誰的胎？ 天上的霜是誰生的呢？
JOB|38|30|諸水堅硬如石頭， 深淵之面凝結成冰。
JOB|38|31|「你能為昴星繫結嗎？ 你能為參星解帶嗎？
JOB|38|32|你能按時領出星宿嗎？ 能引導北斗與其眾星嗎？
JOB|38|33|你知道天的定律嗎？ 你能使地歸其權下嗎？
JOB|38|34|「你能向密雲揚起聲來， 使傾盆的雨遮蓋你嗎？
JOB|38|35|你能發出閃電，使它們 行走， 並對你說：『我們在這裏』嗎？
JOB|38|36|誰將智慧放在朱鷺 中？ 誰將聰明賜給雄雞 ？
JOB|38|37|誰能用智慧數算雲彩？ 誰能傾倒天上的瓶呢？
JOB|38|38|那時，塵土聚集成團， 土塊緊緊結連。
JOB|38|39|「你能為母獅抓取獵物， 使少壯的獅子飽足嗎？
JOB|38|40|那時，牠們在洞中蹲伏， 在隱密處埋伏。
JOB|38|41|誰能為烏鴉預備食物呢？ 那時，烏鴉之雛哀求上帝， 因無食物飛來飛去。」
JOB|39|1|「你知道巖石間的野山羊幾時生產嗎？ 你能觀察母鹿下小鹿嗎？
JOB|39|2|你能數算牠們懷胎的月數嗎？ 你知道牠們幾時生產嗎？
JOB|39|3|牠們屈身，生下幼兒， 就解除了陣痛。
JOB|39|4|其子漸漸肥壯，在荒野長大； 牠們出去，不再歸回。
JOB|39|5|「誰放野驢自由？ 誰解開快驢的繩索？
JOB|39|6|我使曠野作牠的住處， 使鹽地當牠的居所。
JOB|39|7|牠嘲笑城內的喧嚷， 不聽趕牲口的喝聲。
JOB|39|8|諸山是牠漫遊的草場， 牠尋找各樣青綠之物。
JOB|39|9|「野牛豈肯服事你？ 豈肯在你的槽旁過夜？
JOB|39|10|你豈能用套繩將野牛繫於犁溝？ 牠豈肯隨你耙鬆山谷之地？
JOB|39|11|你豈可因牠力大就倚靠牠？ 豈可把你的工交給牠做呢？
JOB|39|12|你豈能靠牠把你的穀物運回， 又收聚在你的禾場上嗎？
JOB|39|13|「鴕鳥的翅膀歡然拍動， 但豈是鸛的翎毛和羽毛嗎 ？
JOB|39|14|因牠把蛋留在地上， 使蛋在塵土中得溫暖，
JOB|39|15|卻忘記腳會把蛋踹碎， 野獸會踐踏它。
JOB|39|16|牠粗暴待雛，似乎不是自己生的； 雖徒然勞苦 ，也不懼怕。
JOB|39|17|因為上帝使牠忘記智慧， 也未將悟性分給牠。
JOB|39|18|牠幾時挺身展開翅膀， 就嘲笑馬和騎馬的人。
JOB|39|19|「馬的力量是你所賜的嗎？ 牠頸項上的鬃是你披上的嗎？
JOB|39|20|是你叫牠跳躍像蝗蟲嗎？ 牠噴氣之威嚴使人驚惶。
JOB|39|21|牠用蹄在谷中挖地 ，以能力歡躍； 牠出去迎擊仇敵 。
JOB|39|22|牠嘲笑懼怕，並不驚惶， 也不因刀劍退卻。
JOB|39|23|箭袋在牠身上錚錚有聲， 槍和短槍閃閃發亮。
JOB|39|24|牠震顫激動，將地吞下 ； 一聽角聲就站不住。
JOB|39|25|每逢角聲一響，牠說：『啊哈！』 牠從遠處聞到戰爭的氣息， 聽見軍官如雷的吼聲和吶喊。
JOB|39|26|「鷹展開翅膀向南飛翔， 豈是藉著你的智慧嗎？
JOB|39|27|大鷹上騰在高處搭窩， 豈是聽你的指示嗎？
JOB|39|28|牠住在山巖， 以山峰和堅固之所為家，
JOB|39|29|從那裏窺察食物， 眼睛自遠方瞭望。
JOB|39|30|牠的雛吸血； 被殺的人在哪裏，牠也在哪裏。」
JOB|40|1|耶和華繼續對 約伯 說：
JOB|40|2|「強辯的豈可與全能者爭論？ 與上帝辯駁的可以回答吧！」
JOB|40|3|於是， 約伯 回答耶和華說：
JOB|40|4|「看哪，我是卑賤的！我用甚麼回答你呢？ 我只好用手摀住我的口。
JOB|40|5|我說了一次，就不回答； 說了兩次，不再說了。」
JOB|40|6|於是，耶和華從旋風中回答 約伯 說：
JOB|40|7|「你要如勇士束腰； 我問你，你可以讓我知道。
JOB|40|8|你豈可廢棄我的判斷？ 豈可定我有罪，好顯自己為義嗎？
JOB|40|9|你有上帝那樣的膀臂嗎？ 你能像他那樣發雷聲嗎？
JOB|40|10|「你要以榮耀莊嚴為妝飾， 以尊榮威嚴為衣服。
JOB|40|11|你要發出你滿溢的怒氣， 見一切驕傲的人，使他降卑；
JOB|40|12|你見一切驕傲的人，將他制伏， 把惡人踐踏在原來地方。
JOB|40|13|你將他們一同埋藏在塵土中， 把他們的臉遮蔽在隱密處 。
JOB|40|14|這樣，我也向你承認， 你的右手能救你自己。
JOB|40|15|「看哪，我造河馬， 也造了你； 牠吃草像牛一樣。
JOB|40|16|看哪，牠的力氣在腰間， 能力在肚腹的肌肉上。
JOB|40|17|牠挺直 尾巴如香柏樹， 牠大腿的筋緊密結合。
JOB|40|18|牠的骨頭好像銅管； 牠的肢體彷彿鐵棍。
JOB|40|19|「牠在上帝所造之物中為首， 只有創造牠的能攜刀臨近牠。
JOB|40|20|諸山為牠產出食物， 百獸也在那裏遊玩。
JOB|40|21|牠伏在蓮葉之下， 在蘆葦和沼澤的隱密處。
JOB|40|22|蓮葉的陰影遮蔽牠， 溪旁的柳樹環繞牠。
JOB|40|23|看哪，河水氾濫，牠不慌張； 連 約旦河 漲到牠口邊，牠也安然自若。
JOB|40|24|誰能在牠眼前捉拿牠呢？ 誰能以圈套穿牠鼻子呢？」
JOB|41|1|「你能用魚鉤釣上 力威亞探 嗎？ 能用繩子壓下牠的舌頭嗎？
JOB|41|2|你能用繩索穿牠的鼻子嗎？ 能用鉤子穿牠的腮骨嗎？
JOB|41|3|牠豈向你連連懇求， 向你說溫柔的話嗎？
JOB|41|4|牠豈肯與你立約， 讓你拿牠永遠作奴僕嗎？
JOB|41|5|你豈可拿牠當雀鳥玩耍？ 豈可將牠繫來給你幼女？
JOB|41|6|合夥的魚販豈可拿牠當貨物？ 他們豈可把牠分給商人呢？
JOB|41|7|你能用倒鉤扎滿牠的皮， 能用魚叉叉滿牠的頭嗎？
JOB|41|8|把你的手掌按在牠身上吧！ 想一想與牠搏鬥，你就不再這樣做了！
JOB|41|9|看哪，對牠有指望是徒然的； 一見牠，豈不也喪膽嗎？
JOB|41|10|沒有那麼兇猛的人敢惹牠。 這樣，誰能在我面前站立得住呢？
JOB|41|11|誰能與我對質，使我償還呢？ 天下萬物都是我的。
JOB|41|12|「我不能緘默不提 牠的肢體和力量，以及健美的骨骼。
JOB|41|13|誰能剝牠的外皮？ 誰能進牠的鎧甲之間 呢？
JOB|41|14|誰能開牠的腮頰？ 牠牙齒的四圍是可畏的。
JOB|41|15|牠的背上有一排排的鱗甲 ， 緊緊閉合，封得嚴密。
JOB|41|16|這鱗甲一一相連， 氣不得透入其間，
JOB|41|17|互相連接， 膠結一起，不能分開。
JOB|41|18|牠打噴嚏就發出光來， 牠的眼睛好像晨曦 。
JOB|41|19|從牠口中發出燒著的火把， 有火星飛迸出來；
JOB|41|20|從牠鼻孔冒出煙來， 如燒開的鍋在沸騰 。
JOB|41|21|牠的氣點著煤炭， 有火焰從牠口中發出。
JOB|41|22|牠頸項中存著勁力， 恐懼在牠面前蹦跳。
JOB|41|23|牠的肉塊緊緊結連， 緊貼其身，不能搖動。
JOB|41|24|牠的心結實如石頭， 如下面的磨石那樣結實。
JOB|41|25|牠一起來，神明都恐懼， 因崩潰而驚慌失措。
JOB|41|26|人用刀劍扎牠，是無用的， 槍、標槍、尖槍也一樣。
JOB|41|27|牠以鐵為乾草， 以銅為爛木。
JOB|41|28|箭不能使牠逃走， 牠看彈石如碎秸。
JOB|41|29|牠當棍棒作碎秸， 牠嘲笑短槍的颼颼聲。
JOB|41|30|牠肚腹下面是尖瓦片； 牠如釘耙刮過淤泥。
JOB|41|31|牠使深淵滾沸如鍋， 使海洋如鍋中膏油。
JOB|41|32|牠使走過以後的路發光， 令人覺得深淵如同白髮。
JOB|41|33|塵世上沒有像牠那樣的受造物， 一無所懼。
JOB|41|34|凡高大的，牠盯著看； 牠在一切狂傲的野獸中作王。」
JOB|42|1|約伯 回答耶和華說：
JOB|42|2|「我知道，你萬事都能做； 你的計劃不能攔阻。
JOB|42|3|誰無知使你的旨意隱藏呢？ 因此我說的，我不明白； 這些事太奇妙，是我不知道的。
JOB|42|4|求你聽我，我要說話； 我問你，求你讓我知道。
JOB|42|5|我從前風聞有你， 現在親眼看見你。
JOB|42|6|因此我撤回 ， 在塵土和爐灰中懊悔。」
JOB|42|7|耶和華對 約伯 說話以後，耶和華就對 提幔 人 以利法 說：「我的怒氣向你和你兩個朋友發作，因為你們議論我，不如我的僕人 約伯 說的正確。
JOB|42|8|現在你們要為自己取七頭公牛，七隻公羊，到我的僕人 約伯 那裏去，為自己獻上燔祭，我的僕人 約伯 就為你們祈禱。我必悅納他，不按你們的愚妄處置你們。你們議論我，不如我的僕人 約伯 說的正確。」
JOB|42|9|於是 提幔 人 以利法 、 書亞 人 比勒達 、 拿瑪 人 瑣法 遵照耶和華所吩咐的去做，耶和華就悅納 約伯 。
JOB|42|10|約伯 為他的朋友祈禱。耶和華就使 約伯 從苦境 中轉回，並且耶和華賜給他的比他從前所有的加倍。
JOB|42|11|約伯 的兄弟、姊妹，和以前所認識的人都來到他那裏，在他家裏跟他一同吃飯。他們因耶和華所降於他的一切災禍，都為他悲傷，安慰他。每人送他一塊可錫塔 和一個金環。
JOB|42|12|這樣，耶和華後來賜福給 約伯 比先前更多。他有一萬四千隻羊，六千匹駱駝，一千對牛，一千匹母驢。
JOB|42|13|他也有七個兒子，三個女兒。
JOB|42|14|他給長女起名叫 耶米瑪 ，次女叫 基洗亞 ，三女叫 基連哈樸 。
JOB|42|15|在全地的婦女中找不著像 約伯 的女兒那樣美貌的。她們的父親使她們在兄弟中得產業。
JOB|42|16|此後， 約伯 又活了一百四十年，得見他的四代兒孫。
JOB|42|17|這樣， 約伯 年紀老邁，日子滿足而死。
PS|1|1|不從惡人的計謀， 不站罪人的道路， 不坐傲慢人的座位， 惟喜愛耶和華的律法， 晝夜思想 他的律法； 這人便為有福！
PS|1|2|
PS|1|3|他要像一棵樹栽在溪水旁， 按時候結果子， 葉子也不枯乾。 凡他所做的盡都順利。
PS|1|4|惡人並不是這樣， 卻像糠秕被風吹散。
PS|1|5|因此，當審判的時候惡人必站立不住， 罪人在義人的會眾中也是如此。
PS|1|6|因為耶和華知道義人的道路， 惡人的道路卻必滅亡。
PS|2|1|列國為甚麼爭鬧？ 萬民為甚麼圖謀虛妄？
PS|2|2|世上的君王都站穩， 臣宰一同算計， 要對抗耶和華， 對抗他的受膏者：
PS|2|3|「我們要掙脫他們的捆綁， 脫去他們的繩索。」
PS|2|4|那坐在天上的必譏笑， 主必嗤笑他們。
PS|2|5|那時，他要在怒中責備他們， 在烈怒中驚嚇他們：
PS|2|6|「我已經在 錫安 －我的聖山 膏立了我的君王。」
PS|2|7|我要傳耶和華的聖旨， 他對我說：「你是我的兒子， 我今日生了你。
PS|2|8|你求我，我就將列國賜你為基業， 將地極賜你為田產。
PS|2|9|你必用鐵杖打破他們， 把他們如同陶匠的瓦器摔碎。」
PS|2|10|現在，君王啊，應當謹慎！ 世上的審判官哪，要聽勸戒！
PS|2|11|當存敬畏的心事奉耶和華， 又當戰兢而快樂。
PS|2|12|當親吻兒子，免得他發怒， 你們就在半途中滅亡， 因為他的怒氣快要發作。 凡投靠他的，都是有福的。
PS|3|1|耶和華啊，我的敵人何其增多！ 許多人起來攻擊我。
PS|3|2|許多人議論我： 「他得不到上帝的幫助。」（細拉）
PS|3|3|但你－耶和華是我四圍的盾牌， 是我的榮耀，又是令我抬起頭來的。
PS|3|4|我用我的聲音求告耶和華， 他就從他的聖山上應允我。（細拉）
PS|3|5|我躺下，我睡覺，我醒來， 耶和華都保佑我。
PS|3|6|雖有成萬的百姓周圍攻擊我， 我也不懼怕。
PS|3|7|耶和華啊，求你興起！ 我的上帝啊，求你救我！ 因為你打斷我所有仇敵的腮骨， 敲碎了惡人的牙齒。
PS|3|8|救恩屬於耶和華； 願你賜福給你的百姓。（細拉）
PS|4|1|顯我為義的上帝啊， 我呼求的時候，求你應允我！ 我在困境中，你曾使我寬暢； 求你憐憫我，聽我的禱告！
PS|4|2|你們這些人哪，你們把我的尊榮變為羞辱，要到幾時呢？ 你們喜愛虛妄，尋找虛假，要到幾時呢？ （細拉）
PS|4|3|你們要知道，耶和華已將虔誠人分別出來歸他自己； 我求告耶和華，他必垂聽。
PS|4|4|應當畏懼，不可犯罪； 在床上的時候，要心裏思想，並要安靜。（細拉）
PS|4|5|當獻上公義的祭， 又當倚靠耶和華。
PS|4|6|有許多人說：「誰能指示我們甚麼好處？ 耶和華啊，求你用你臉上的光照耀我們。」
PS|4|7|你使我心裏喜樂， 勝過那豐收五穀新酒的人。
PS|4|8|我必平安地躺下睡覺， 因為獨有你－耶和華使我安然居住。
PS|5|1|耶和華啊，求你側耳聽我的言語， 顧念我的心思！
PS|5|2|我的王，我的上帝啊，求你留心聽我呼求的聲音！ 因為我向你祈禱。
PS|5|3|耶和華啊，早晨你必聽我的聲音； 早晨我要向你陳明我的心思，並要警醒。
PS|5|4|因為你不是喜愛邪惡的上帝， 惡人不能與你同住。
PS|5|5|狂傲的人不能站在你眼前； 凡作惡的，都是你所恨惡的。
PS|5|6|說謊言的，你必滅絕； 好流人血、玩弄詭詐的，都為耶和華所憎惡。
PS|5|7|至於我，我必憑你豐盛的慈愛進入你的居所， 我要存敬畏你的心向你的聖殿下拜。
PS|5|8|耶和華啊，求你因我仇敵的緣故，憑你的公義引領我， 使你的道路在我面前正直。
PS|5|9|因為他們口中沒有誠實， 心裏充滿邪惡， 他們的喉嚨是敞開的墳墓； 他們用舌頭諂媚人。
PS|5|10|上帝啊，求你定他們的罪！ 願他們因自己的計謀跌倒； 求你因他們過犯眾多趕逐他們， 因為他們背叛了你。
PS|5|11|凡投靠你的，願他們喜樂，時常歡呼， 因為你庇護他們； 又願那愛你名的人都靠你歡欣。
PS|5|12|耶和華啊，因為你必賜福給義人， 你必用恩惠如同盾牌四面護衛他。
PS|6|1|耶和華啊，求你不要在怒中責備我， 不要在烈怒中懲罰我！
PS|6|2|耶和華啊，求你憐憫我，因為我軟弱。 耶和華啊，求你醫治我，因為我的骨頭戰抖。
PS|6|3|我的心也大大驚惶。 耶和華啊，你要等到幾時呢？
PS|6|4|耶和華啊，求你轉回搭救我， 因你的慈愛拯救我。
PS|6|5|因為死了的人不會記念你， 在陰間有誰稱謝你？
PS|6|6|我因呻吟而困乏； 我每夜流淚，使床鋪漂起， 把褥子濕透。
PS|6|7|我的眼睛因憂愁而昏花， 因敵人的緣故，我的眼目模糊不清。
PS|6|8|你們所有作惡的人，離開我吧！ 因為耶和華聽了我哀哭的聲音。
PS|6|9|耶和華聽了我的懇求， 耶和華必接納我的禱告。
PS|6|10|我所有的仇敵都必羞愧，大大驚惶； 轉眼之間，他們要羞愧撤退。
PS|7|1|耶和華－我的上帝啊，我投靠你！ 求你救我脫離所有追趕我的人，搭救我出來！
PS|7|2|免得他們像獅子撕裂我， 甚至撕碎，無人搭救。
PS|7|3|耶和華－我的上帝啊，我若行了這事， 若有罪孽在我手裏，
PS|7|4|我若以惡回報我的朋友， 連那無故與我為敵的，我也救了他 ，
PS|7|5|就任憑仇敵追趕我，直到追上， 把我的性命踏在地上， 使我的榮耀歸於灰塵。（細拉）
PS|7|6|耶和華啊，求你在怒中起來， 挺身而立，抵擋我敵人的烈怒！ 求你為我興起！你已經發令施行審判。
PS|7|7|願萬民聚集環繞你！ 願你居高位統治他們！
PS|7|8|耶和華向萬民施行審判； 耶和華啊，求你按我的公義 和我心中的純正判斷我。
PS|7|9|願惡人的惡斷絕！ 願你堅立義人！ 因為公義的上帝察驗人的心腸肺腑。
PS|7|10|上帝是我的盾牌， 他拯救心裏正直的人。
PS|7|11|上帝是公義的審判者， 又是天天向惡人發怒的上帝。
PS|7|12|若有人不回頭，他的刀必磨快， 弓必上弦，預備妥當。
PS|7|13|他也預備了致死的兵器， 他所射的是火箭。
PS|7|14|看哪，惡人懷邪惡， 養毒害，生虛假。
PS|7|15|他掘了坑，挖得太深， 竟掉在自己所挖的陷阱裏。
PS|7|16|他的毒害必回到自己頭上， 他的殘暴必落到自己的腦袋上。
PS|7|17|我要照著耶和華的公義稱謝他， 要歌頌耶和華至高者的名。
PS|8|1|耶和華－我們的主啊， 你的名在全地何其美！ 你將你的榮耀彰顯於天 。
PS|8|2|你因敵人的緣故， 從孩童和吃奶的口中建立了能力， 使仇敵和報仇的閉口無言。
PS|8|3|我觀看你手指所造的天， 並你所陳設的月亮星宿。
PS|8|4|人算甚麼，你竟顧念他！ 世人算甚麼，你竟眷顧他！
PS|8|5|你使他比上帝 微小一點， 賜他榮耀尊貴為冠冕。
PS|8|6|你派他管理你手所造的， 使萬物，就是一切的牛羊、 田野的牲畜、空中的鳥、海裏的魚， 凡游在水裏的，都服在他的腳下。
PS|8|7|
PS|8|8|
PS|8|9|耶和華－我們的主啊， 你的名在全地何其美！
PS|9|1|我要一心稱謝耶和華， 傳揚你一切奇妙的作為。
PS|9|2|我要因你歡喜快樂； 至高者啊，我要歌頌你的名！
PS|9|3|我的仇敵回轉撤退的時候， 他們在你面前跌倒滅亡。
PS|9|4|因你已經為我伸冤，為我辯護； 你坐在寶座上，按公義審判。
PS|9|5|你曾斥責列國，滅絕惡人； 你曾塗去他們的名，直到永永遠遠。
PS|9|6|仇敵到了盡頭； 他們遭毀壞，直到永遠。 你拆毀他們的城鎮， 連他們的名字 也都消滅！
PS|9|7|惟耶和華坐在王位上，直到永遠； 他已經為審判擺設寶座。
PS|9|8|他要按公義審判世界， 按正直判斷萬民。
PS|9|9|耶和華要作受欺壓者的庇護所， 在患難時的庇護所。
PS|9|10|耶和華啊，認識你名的人要倚靠你， 因你沒有離棄尋求你的人。
PS|9|11|應當歌頌居於 錫安 的耶和華， 將他所做的傳揚在萬民中。
PS|9|12|那位追討流人血的， 他記念受屈的人， 不忘記困苦人的哀求。
PS|9|13|耶和華啊，求你憐憫我！ 你是從死門把我提升起來的， 求你看那恨我的人所加給我的苦難，
PS|9|14|好讓我述說你一切的美德。 我要在 錫安 的城門因你的救恩歡樂。
PS|9|15|外邦人陷在自己所掘的坑中， 他們的腳被自己暗設的網羅纏住了。
PS|9|16|耶和華已將自己顯明，他已施行審判； 惡人被自己手所做的纏住了 。（細拉）
PS|9|17|惡人，就是忘記上帝的外邦人， 都必歸到陰間。
PS|9|18|貧窮人必不永久被忘， 困苦人的指望必不永遠落空。
PS|9|19|耶和華啊，求你興起，不容世人得勝！ 願外邦人在你面前受審判！
PS|9|20|耶和華啊，求你使他們恐懼， 願外邦人知道自己不過是人。（細拉）
PS|10|1|耶和華啊，你為甚麼站在遠處？ 在患難的時候為甚麼隱藏？
PS|10|2|惡人驕橫地追逼困苦人； 願他們陷在自己所設的計謀裏。
PS|10|3|因為惡人以自己的心願自誇， 貪財的背棄耶和華，並且輕慢他 。
PS|10|4|惡人面帶驕傲，不尋找耶和華； 他的思想中全無上帝。
PS|10|5|他的路時常亨通， 你的審判不在他眼裏。 至於他所有的敵人，他都向他們發怒氣。
PS|10|6|他心裏說：「我必不動搖， 世世代代不遭災難。」
PS|10|7|他滿口咒罵、詭詐、欺壓， 舌底盡是毒害、奸惡。
PS|10|8|他在村莊埋伏等候， 在隱密處殺害無辜的人， 他的眼睛窺探無倚無靠的人。
PS|10|9|他埋伏在暗地，如獅子蹲在洞中。 他埋伏，要俘擄困苦人； 他拉網，就把困苦人擄去。
PS|10|10|他屈身蹲伏， 無倚無靠的人就倒在他的暴力之下。
PS|10|11|他心裏說：「上帝竟忘記了， 上帝轉臉永不觀看。」
PS|10|12|耶和華啊，求你興起！ 上帝啊，求你舉手！ 不要忘記困苦人！
PS|10|13|惡人為何輕慢上帝， 心裏說「你必不追究」？
PS|10|14|你已經察看， 顧念人的憂患和愁苦， 放在你的手中。 無倚無靠的人把自己交託給你， 你向來是幫助孤兒的。
PS|10|15|求你打斷惡人的膀臂， 至於壞人，求你追究他的惡，直到淨盡。
PS|10|16|耶和華永永遠遠為王， 外邦人從他的地已經滅絕了。
PS|10|17|耶和華啊，困苦人的心願你早已聽見； 你必堅固他們的心，也必側耳聽他們的祈求，
PS|10|18|為要給孤兒和受欺壓的人伸冤， 使世上的人不再威嚇他們。
PS|11|1|我投靠耶和華； 你們怎麼對我說：「你當像鳥逃到你們的山去；
PS|11|2|看哪，惡人彎弓，把箭搭在弦上， 要在暗中射那心裏正直的人。
PS|11|3|根基若毀壞， 義人還能做甚麼呢？」
PS|11|4|耶和華在他的聖殿裏， 耶和華在天上的寶座上； 他的眼睛察看， 他的眼目 察驗世人。
PS|11|5|耶和華考驗義人； 惟有惡人和喜愛暴力的人，他心裏恨惡。
PS|11|6|他要向惡人密佈羅網， 烈火、硫磺、熱風作他們杯中的份。
PS|11|7|因為耶和華是公義的，他喜愛義行， 正直人必得見他的面。
PS|12|1|耶和華啊，求你幫助，因虔誠人斷絕了， 世人中間忠信的人消失了。
PS|12|2|人人向鄰舍說謊； 他們說話嘴唇油滑，心口不一。
PS|12|3|願耶和華剪除一切油滑的嘴唇， 誇大的舌頭。
PS|12|4|他們說：「我們必能以舌頭取勝， 我們的嘴唇是自己的， 誰能作我們的主呢？」
PS|12|5|耶和華說：「因為困苦人的冤屈 和貧窮人的嘆息， 我現在要起來， 把他安置在他所切慕的穩妥之地。」
PS|12|6|耶和華的言語是純淨的言語， 如同銀子在泥做的爐中煉過七次。
PS|12|7|耶和華啊，你必保護他們， 你必保佑他們永遠脫離這世代的人。
PS|12|8|卑鄙的人在世人中高升時， 就有惡人四處橫行。
PS|13|1|耶和華啊，你忘記我要到幾時呢？要到永遠嗎？ 你轉臉不顧我要到幾時呢？
PS|13|2|我心裏籌算，終日愁苦，要到幾時呢？ 我的仇敵升高壓制我，要到幾時呢？
PS|13|3|耶和華－我的上帝啊，求你看顧我，應允我！ 求你使我眼目明亮，免得我沉睡至死；
PS|13|4|免得我的仇敵說「我勝了他」； 免得我的敵人在我動搖的時候喜樂。
PS|13|5|但我倚靠你的慈愛， 我的心因你的救恩快樂。
PS|13|6|我要向耶和華歌唱， 因他厚厚地恩待我。
PS|14|1|愚頑人心裏說：「沒有上帝。」 他們都敗壞，行了可憎惡的事， 沒有一個人行善。
PS|14|2|耶和華從天上垂看世人， 要看有明白的沒有， 有尋求上帝的沒有。
PS|14|3|他們都偏離正路，一同變為污穢， 沒有行善的， 連一個也沒有。
PS|14|4|作惡的都沒有知識嗎？ 他們吞吃我的百姓如同吃飯一樣， 並不求告耶和華。
PS|14|5|他們在那裏大大害怕， 因為上帝在義人的族類中。
PS|14|6|你們叫困苦人的籌算變為羞辱， 然而耶和華是他的避難所。
PS|14|7|但願 以色列 的救恩出自 錫安 。 當耶和華救回他被擄子民的時候， 雅各 要快樂， 以色列 要歡喜。
PS|15|1|耶和華啊，誰能寄居你的帳幕？ 誰能居住你的聖山？
PS|15|2|就是行為正直、做事公義、 心裏說實話的人。
PS|15|3|他不以舌頭讒害人， 不惡待朋友， 也不隨夥毀謗鄰舍。
PS|15|4|他眼中藐視匪類， 卻尊重那敬畏耶和華的人。 他發了誓，雖然自己吃虧也不更改。
PS|15|5|他不放債取利， 不受賄賂以害無辜。 做這些事的人必永不動搖。
PS|16|1|上帝啊，求你保佑我， 因為我投靠你。
PS|16|2|我 曾對耶和華說：「你是我的主， 我的福氣惟獨從你而來。」
PS|16|3|論到世上的聖民，他們是尊貴的人， 是我最喜悅的。
PS|16|4|追逐 別神的， 他們的愁苦必增加； 他們所澆奠的血我不獻上， 我嘴唇也不提別神的名號。
PS|16|5|耶和華是我的產業，是我杯中的福分； 我所得的，你為我持守。
PS|16|6|用繩量給我的地界，坐落在佳美之處； 我的產業實在美好。
PS|16|7|我要稱頌那指引我的耶和華， 在夜間我的心腸也指教我。
PS|16|8|我讓耶和華常在我面前， 因他在我右邊，我就不致動搖。
PS|16|9|因此，我的心歡喜，我的靈 快樂； 我的肉身也要安然居住。
PS|16|10|因為你必不將我的靈魂 撇在陰間， 也不讓你的聖者見地府 。
PS|16|11|你必將生命的道路指示我。 在你面前有滿足的喜樂， 在你右手中有永遠的福樂。
PS|17|1|耶和華啊，求你垂聽公義的呼聲， 留心聽我的呼求！ 求你側耳聽我這沒有詭詐的嘴唇的祈禱！
PS|17|2|願判我公正的話從你面前發出， 願你的眼睛察看正直。
PS|17|3|你已經考驗我的心， 你在夜間鑒察我。 你熬煉我，卻找不到錯失， 我立志叫我口中沒有過失。
PS|17|4|論到人的行為，我謹守你嘴唇的言語， 不走殘暴人的道路。
PS|17|5|我的腳緊緊跟隨你的腳蹤， 我的兩腳未曾滑跌。
PS|17|6|上帝啊，我求告你，因為你必應允我； 求你向我側耳，聽我的言語。
PS|17|7|求你顯出你奇妙的慈愛， 你用右手拯救投靠你的人，脫離那起來攻擊他們的人。
PS|17|8|求你保護我，如同保護眼中的瞳人， 把我隱藏在你翅膀的蔭下，
PS|17|9|使我脫離欺壓我的惡人， 脫離那圍困我要害我命的仇敵。
PS|17|10|他們的心被油脂包裹， 用口說驕傲的話。
PS|17|11|他們追逼我 ，現在他們圍困了我們， 瞪著眼，要把我們推倒在地。
PS|17|12|他像獅子要貪吃獵物， 又像少壯獅子蹲伏在暗處。
PS|17|13|耶和華啊，求你興起，前去迎敵，把他打倒！ 求你用你的刀救我的命脫離惡人。
PS|17|14|耶和華啊，求你用手救我脫離世人， 脫離那只在今生有福分的世人！ 你以財寶充滿他們的肚腹， 他們因有兒女就滿足， 將其餘的財物留給他們的孩子。
PS|17|15|至於我，我必因公正得見你的面； 我醒了的時候，你的形像使我滿足。
PS|18|1|耶和華我的力量啊，我愛你！
PS|18|2|耶和華是我的巖石、我的山寨、我的救主、 我的上帝、我的磐石、我所投靠的。 他是我的盾牌， 是拯救我的角，是我的碉堡。
PS|18|3|我要求告當讚美的耶和華， 我必從仇敵手中被救出來。
PS|18|4|死亡的繩索勒住我， 毀滅的急流驚嚇我，
PS|18|5|陰間的繩索纏繞我， 死亡的圈套臨到我。
PS|18|6|我在急難中求告耶和華， 向我的上帝呼求。 他從殿中聽了我的聲音， 我在他面前的呼求必進入他耳中。
PS|18|7|那時，因他發怒地就震動戰抖， 山的根基也震動挪移。
PS|18|8|他的鼻孔冒煙上騰， 他的口發火焚燒，連煤炭也燒著了。
PS|18|9|他使天垂下，親自降臨， 黑雲在他腳下。
PS|18|10|他乘坐基路伯飛行， 藉著風的翅膀快飛，
PS|18|11|以黑暗為藏身之處， 以水的黑暗、天空的密雲作四圍的行宮。
PS|18|12|因他發出光輝， 冰雹和火炭穿透密雲。
PS|18|13|耶和華在天上打雷， 至高者發出聲音，就有冰雹和火炭 。
PS|18|14|他射出箭來，使仇敵四散； 發出連串的閃電，擊潰他們。
PS|18|15|耶和華啊，你的斥責一發， 你鼻孔的氣一出， 海底就顯現， 大地的根基也暴露。
PS|18|16|他從高天伸手抓住我， 把我從大水中拉上來。
PS|18|17|他救我脫離強敵和那些恨我的人， 因為他們比我強盛。
PS|18|18|我遭遇災難的日子，他們來攻擊我； 但耶和華是我的倚靠。
PS|18|19|他領我到寬闊之處， 他救拔我，因他喜愛我。
PS|18|20|耶和華必按我的公義報答我， 按我手中的清潔賞賜我。
PS|18|21|因為我遵守耶和華的道， 未曾作惡離開我的上帝。
PS|18|22|他的一切典章常在我面前， 他的律例我也未曾丟棄。
PS|18|23|我在他面前作了完全人， 我也保護自己遠離罪孽。
PS|18|24|所以耶和華按我的公義， 在他眼前按我手中的清潔賞賜我。
PS|18|25|慈愛的人，你以慈愛待他； 完全的人，你以完善待他。
PS|18|26|清潔的人，你以清潔待他； 歪曲的人，你以彎曲待他。
PS|18|27|困苦的百姓，你必拯救； 高傲的眼目，你使他降卑。
PS|18|28|你必點亮我的燈； 耶和華－我的上帝必照明我的黑暗。
PS|18|29|我藉著你衝入敵軍， 藉著我的上帝跳過城牆。
PS|18|30|至於上帝，他的道是完全的； 耶和華的話是純淨的。 凡投靠他的，他就作他們的盾牌。
PS|18|31|除了耶和華，誰是上帝呢？ 除了我們的上帝，誰是磐石呢？
PS|18|32|惟有那以力量束我的腰、 使我行為完全的，他是上帝。
PS|18|33|他使我的腳快如母鹿， 使我站穩在高處。
PS|18|34|他教導我的手能爭戰， 我的膀臂能開銅造的弓。
PS|18|35|你賜救恩給我作盾牌， 你的右手扶持我， 你的庇護 使我為大。
PS|18|36|你使我腳步寬闊， 我的腳踝未曾滑跌。
PS|18|37|我要追趕我的仇敵，且要追上他們； 若不將他們滅絕，我總不歸回。
PS|18|38|我要打傷他們，使他們站不起來； 他們必倒在我的腳下。
PS|18|39|你曾以力量束我的腰，使我能爭戰； 也曾使那起來攻擊我的，都服在我以下。
PS|18|40|你又使我的仇敵在我面前轉身逃跑， 使我剪除那恨我的人。
PS|18|41|他們呼求，卻無人拯救； 就是呼求耶和華，他也不應允。
PS|18|42|我搗碎他們，如同風前的灰塵； 傾倒 他們，如同街上的泥土。
PS|18|43|你救我脫離百姓的紛爭， 立我作列國的元首； 我素不認識的百姓必事奉我。
PS|18|44|他們一聽見我的名聲就必順從我， 外邦人要投降我。
PS|18|45|外邦人要喪膽， 戰戰兢兢地出營寨。
PS|18|46|耶和華永遠活著。 願我的磐石被稱頌， 願救我的上帝受尊崇。
PS|18|47|這位上帝為我伸冤， 使萬民服在我以下。
PS|18|48|他拯救我脫離仇敵， 又把我舉起，高過那些起來攻擊我的人， 救我脫離殘暴的人。
PS|18|49|耶和華啊，因此我要在外邦中稱謝你， 歌頌你的名。
PS|18|50|耶和華賜極大的救恩給他所立的王， 施慈愛給他的受膏者， 就是給 大衛 和他的後裔，直到永遠。
PS|19|1|諸天述說上帝的榮耀， 穹蒼傳揚他手的作為。
PS|19|2|這日到那日發出言語， 這夜到那夜傳出知識。
PS|19|3|無言無語， 也無聲音可聽。
PS|19|4|它們的聲浪 傳遍天下， 它們的言語傳到地極。 上帝在其中為太陽安設帳幕，
PS|19|5|太陽如同新郎步出洞房， 又如勇士歡然奔路。
PS|19|6|它從天這邊出來，繞到天那邊， 沒有一物可隱藏得不到它的熱氣。
PS|19|7|耶和華的律法全備，使人甦醒； 耶和華的法度確定，使愚蒙人有智慧。
PS|19|8|耶和華的訓詞正直，使人心快活； 耶和華的命令清潔，使人眼目明亮。
PS|19|9|耶和華的典章真實，全然公義， 敬畏耶和華是純潔的，存到永遠，
PS|19|10|比金子可羨慕，比極多的純金可羨慕； 比蜜甘甜，比蜂房下滴的蜜甘甜。
PS|19|11|因此你的僕人受警戒， 遵守這些有極大的賞賜。
PS|19|12|誰能察覺自己的錯失呢？ 求你赦免我隱藏的過犯。
PS|19|13|求你攔阻僕人不犯任意妄為的罪， 不容這罪轄制我， 我就完全，免犯大罪。
PS|19|14|耶和華－我的磐石，我的救贖主啊， 願我口中的言語，心裏的意念在你面前蒙悅納。
PS|20|1|願耶和華在你患難的日子應允你， 願 雅各 的上帝的名保護你。
PS|20|2|願他從聖所救助你， 從 錫安 堅固你，
PS|20|3|記念你的一切祭物， 悅納你的燔祭，（細拉）
PS|20|4|將你心所願的賜給你， 成就你的一切籌算。
PS|20|5|我們要因你的救恩誇勝， 要奉我們上帝的名豎立旌旗。 願耶和華成就你一切所求的！
PS|20|6|現在我知道耶和華必救護他的受膏者， 從他神聖的天上應允他， 用右手的能力救護他。
PS|20|7|有人靠車，有人靠馬， 但我們要提耶和華－我們上帝的名。
PS|20|8|他們都屈身仆倒， 我們卻起來，堅立不移。
PS|20|9|耶和華啊，求你拯救； 我們呼求的時候，願王應允我們！
PS|21|1|耶和華啊，王必因你的能力歡喜； 因你的救恩，他的快樂何其大！
PS|21|2|他心裏所願的，你已經賜給他； 他嘴唇所求的，你未嘗不應允。（細拉）
PS|21|3|你以美善的福氣迎接他， 把純金的冠冕戴在他頭上。
PS|21|4|他向你祈求長壽，你就賜給他， 就是日子長久，直到永遠。
PS|21|5|他因你的救恩大有榮耀， 你將尊榮威嚴加在他身上。
PS|21|6|你使他有洪福，直到永遠， 又使他在你面前歡喜快樂。
PS|21|7|王倚靠耶和華， 因至高者的慈愛，王必不動搖。
PS|21|8|你的手要搜出所有的仇敵， 你的右手要搜出那些恨你的人。
PS|21|9|你的臉出現的時候，要使他們如在炎熱的火爐中。 耶和華要在他的震怒中吞滅他們， 那火要把他們燒盡。
PS|21|10|你必從世上滅絕他們的幼苗， 從人間滅絕他們的後裔。
PS|21|11|因為他們有意加害於你； 他們想出計謀，卻不能做成。
PS|21|12|你必使他們轉身逃跑， 向著他們的臉搭箭在弦。
PS|21|13|耶和華啊，願你因自己的能力顯為至高！ 這樣，我們就唱詩，歌頌你的大能。
PS|22|1|我的上帝，我的上帝，為甚麼離棄我？ 為甚麼遠離不救我，不聽我的呻吟？
PS|22|2|我的上帝啊，我白日呼求，你不應允； 夜間呼求，也不得安寧。
PS|22|3|但你是神聖的， 用 以色列 的讚美為寶座。
PS|22|4|我們的祖宗倚靠你； 他們倚靠你，你解救他們。
PS|22|5|他們哀求你，就蒙解救； 他們倚靠你，就不羞愧。
PS|22|6|但我是蟲，不是人， 被眾人羞辱，被百姓藐視。
PS|22|7|凡看見我的都嗤笑我； 他們撇嘴搖頭：
PS|22|8|「他把自己交託給耶和華，讓耶和華救他吧！ 耶和華既喜愛他，可以搭救他吧！」
PS|22|9|但你是叫我出母腹的， 我在母懷裏，你就使我有倚靠的心。
PS|22|10|我自出母胎就交在你手裏， 自我出母腹，你就是我的上帝。
PS|22|11|求你不要遠離我！ 因為災難臨頭，無人幫助。
PS|22|12|許多公牛環繞我， 巴珊 大力的公牛四面圍困我。
PS|22|13|牠們向我張口， 好像獵食吼叫的獅子。
PS|22|14|我如水被倒出， 我的骨頭都脫了節， 我的心如蠟，在我裏面熔化。
PS|22|15|我的精力枯乾，如同瓦片， 我的舌頭緊貼上顎。 你將我安置在死灰中。
PS|22|16|犬類圍著我，惡黨環繞我； 他們扎了我的手、我的腳。
PS|22|17|我數遍我的骨頭； 他們瞪著眼看我。
PS|22|18|他們分我的外衣， 為我的內衣抽籤。
PS|22|19|耶和華啊，求你不要遠離我！ 我的救主啊，求你快來幫助我！
PS|22|20|求你救我的性命脫離刀劍， 使我僅有的 脫離犬類，
PS|22|21|求你救我脫離獅子的口； 你已經應允我，使我脫離野牛的角。
PS|22|22|我要將你的名傳給我的弟兄， 在會眾中我要讚美你。
PS|22|23|敬畏耶和華的人哪，要讚美他！ 雅各 的後裔啊，要榮耀他！ 以色列 的後裔啊，要懼怕他！
PS|22|24|因為他沒有藐視、憎惡受苦的人， 也沒有轉臉不顧他們； 那受苦之人呼求的時候，他就垂聽。
PS|22|25|我在大會中讚美你的話是從你而來， 我要在敬畏耶和華的人面前還我的願。
PS|22|26|願困苦的人吃得飽足， 願尋求耶和華的人讚美他。 願你們的心永遠活著！
PS|22|27|地的四極都要想念耶和華，並且歸順他， 列國的萬族都要在你面前敬拜。
PS|22|28|因為國度屬於耶和華， 他是管理列國的。
PS|22|29|地上富足的人都必吃喝而敬拜， 凡下到塵土中不能存活自己性命的人， 都要在他面前下拜 ；
PS|22|30|必有後裔事奉他， 主所做的事必傳給後代。
PS|22|31|他們必來傳他的公義給尚未出生的子民， 這是他的作為。
PS|23|1|耶和華是我的牧者， 我必不致缺乏。
PS|23|2|他使我躺臥在青草地上， 領我在可安歇的水邊。
PS|23|3|他使我的靈魂甦醒 ， 為自己的名引導我走義路。
PS|23|4|我雖然行過死蔭的幽谷， 也不怕遭害， 因為你與我同在； 你的杖、你的竿，都安慰我。
PS|23|5|在我敵人面前，你為我擺設筵席； 你用油膏了我的頭，使我的福杯滿溢。
PS|23|6|我一生一世必有恩惠慈愛隨著我； 我且要住在 耶和華的殿中，直到永遠。
PS|24|1|地和其中所充滿的， 世界和住在其中的，都屬耶和華。
PS|24|2|他把地建立在海上， 安定在江河之上。
PS|24|3|誰能登耶和華的山？ 誰能站在他的聖所？
PS|24|4|就是手潔心清，意念不向虛妄， 起誓不懷詭詐的人。
PS|24|5|他必蒙耶和華賜福， 又蒙救他的上帝使他成義。
PS|24|6|這是尋求耶和華的族類， 是尋求你面的 雅各 。（細拉）
PS|24|7|眾城門哪，要抬起頭來！ 永久的門戶啊，你們要被舉起！ 榮耀的王將要進來！
PS|24|8|這榮耀的王是誰呢？ 就是有力有能的耶和華， 在戰場上大有能力的耶和華！
PS|24|9|眾城門哪，要抬起頭來！ 永久的門戶啊，你們要高舉！ 榮耀的王將要進來！
PS|24|10|這榮耀的王是誰呢？ 萬軍之耶和華是榮耀的王！（細拉）
PS|25|1|耶和華啊，我的心仰望你。
PS|25|2|我的上帝啊，我素來倚靠你； 求你不要叫我羞愧， 不要叫我的仇敵向我誇勝。
PS|25|3|凡等候你的必不羞愧， 惟有那無故行奸詐的必要羞愧。
PS|25|4|耶和華啊，求你將你的道指示我， 將你的路指教我！
PS|25|5|求你指教我，引導我進入你的真理， 因為你是救我的上帝。 我整日等候你。
PS|25|6|耶和華啊，求你記念你的憐憫和慈愛， 因為這是亙古以來所常有的。
PS|25|7|求你不要記得我幼年的罪愆和我的過犯； 耶和華啊，求你因你的良善，按你的慈愛記念我。
PS|25|8|耶和華是良善正直的， 因此，他必教導罪人走正路。
PS|25|9|他要按公平引領謙卑人， 將他的道指教他們。
PS|25|10|凡遵守他的約和他法度的人， 耶和華都以慈愛信實待他。
PS|25|11|耶和華啊，求你因你名的緣故赦免我的罪， 因我的罪重大。
PS|25|12|誰敬畏耶和華， 耶和華必教導他當選擇的道路。
PS|25|13|他要安然居住， 他的後裔必承受土地。
PS|25|14|耶和華與敬畏他的人親密， 他要將自己的約指示他們。
PS|25|15|我的眼目時常仰望耶和華， 因他必將我的腳從網裏拉出來。
PS|25|16|求你轉向我，憐憫我， 因我孤獨困苦。
PS|25|17|我心裏愁苦甚多， 求你救我脫離我的禍患。
PS|25|18|求你看顧我的困苦、我的艱難， 赦免我一切的罪。
PS|25|19|求你察看我的仇敵， 因為他們人數眾多，並且痛恨我。
PS|25|20|求你保護我的性命，搭救我， 使我不致羞愧，因為我投靠你。
PS|25|21|願純全、正直保護我， 因為我等候你。
PS|25|22|上帝啊，求你救贖 以色列 脫離他一切的愁苦。
PS|26|1|耶和華啊，求你為我伸冤， 因我向來行事純正； 我倚靠耶和華，必不動搖。
PS|26|2|耶和華啊，求你察看我，考驗我， 熬煉我的肺腑心腸。
PS|26|3|因為你的慈愛常在我眼前， 我也按你的真理而行。
PS|26|4|我未曾與虛妄的人同坐， 也不與偽善的人來往。
PS|26|5|我痛恨惡人的集會， 必不與惡人同坐。
PS|26|6|耶和華啊，我要洗手表明無辜， 才環繞你的祭壇；
PS|26|7|我好發出稱謝的聲音， 述說你一切奇妙的作為。
PS|26|8|耶和華啊，我喜愛你所住的殿 和你顯榮耀的居所。
PS|26|9|不要把我的性命和罪人一同除掉， 不要把我的生命和好流人血的一同除掉。
PS|26|10|他們的手中有奸惡， 他們的右手滿有賄賂。
PS|26|11|至於我，卻要行事純正； 求你救贖我，憐憫我！
PS|26|12|我的腳站在平坦的地方， 在聚會中我要稱頌耶和華！
PS|27|1|耶和華是我的亮光，是我的拯救， 我還怕誰呢？ 耶和華是我生命的保障， 我還懼誰呢？
PS|27|2|那作惡的就是我的仇敵， 前來吃我肉的時候就絆跌仆倒。
PS|27|3|雖有軍隊安營攻擊我，我的心也不害怕； 雖然興起戰爭攻擊我，我仍舊安穩。
PS|27|4|有一件事，我曾求耶和華，我仍要尋求， 就是一生一世住在耶和華的殿中， 瞻仰他的榮美，在他的殿宇裏求問。
PS|27|5|因為我遭遇患難，他必將我隱藏在他的帳棚裏， 把我藏在他帳幕的隱密處， 將我高舉在磐石上。
PS|27|6|現在我得以昂首，高過四面的仇敵。 我要在他的帳幕裏歡然獻祭， 我要唱詩歌頌耶和華。
PS|27|7|耶和華啊，我呼求的時候，求你垂聽我的聲音； 求你憐憫我，應允我。
PS|27|8|你說：「你們當尋求我的面。」 那時我的心向你說： 「耶和華啊，你的面我正要尋求。」
PS|27|9|求你不要轉臉不顧我， 不要發怒趕逐你的僕人， 你向來是幫助我的。 救我的上帝啊，不要離開我， 也不要撇棄我。
PS|27|10|即使我的父母撇棄我， 耶和華終必收留我。
PS|27|11|耶和華啊，求你將你的道指教我， 因我仇敵的緣故引導我走平坦的路。
PS|27|12|求你不要把我交給敵人，遂其所願； 因為妄作見證的和口吐凶言的都起來攻擊我。
PS|27|13|我深信在活人之地 必得見耶和華的恩惠。
PS|27|14|要等候耶和華， 當壯膽，堅固你的心， 要等候耶和華！
PS|28|1|耶和華啊，我要求告你！ 我的磐石啊，求你不要向我緘默！ 倘若你向我閉口， 我就如下入地府的人一樣。
PS|28|2|我呼求你，向你至聖所舉手的時候， 求你垂聽我懇求的聲音！
PS|28|3|不要把我和壞人並作惡的一同除掉； 他們跟鄰舍說平安，心裏卻是奸惡。
PS|28|4|求你按著他們所做的， 按他們的惡行對待他們； 求你照著他們手所做的對待他們， 將他們應得的報應加給他們。
PS|28|5|他們既然不尊重耶和華的作為， 也不尊重他手所做的， 耶和華就必毀壞他們，不建立他們。
PS|28|6|耶和華是應當稱頌的， 因為他聽了我懇求的聲音。
PS|28|7|耶和華是我的力量，是我的盾牌， 我心裏倚靠他就得幫助。 我心中歡樂， 我要用詩歌稱謝他。
PS|28|8|耶和華是他百姓的力量， 又是他受膏者得救的保障。
PS|28|9|求你拯救你的百姓，賜福給你的產業； 求你牧養他們，扶持他們，直到永遠。
PS|29|1|上帝的子民 哪，你們要將榮耀、能力歸給耶和華， 都歸給耶和華！
PS|29|2|要將耶和華的名的榮耀歸給他， 要敬拜神聖榮耀的耶和華 。
PS|29|3|耶和華的聲音在眾水上， 榮耀的上帝打雷； 耶和華打雷在大水之上。
PS|29|4|耶和華的聲音大有能力， 耶和華的聲音滿有威嚴。
PS|29|5|耶和華的聲音震碎香柏樹， 耶和華震碎 黎巴嫩 的香柏樹。
PS|29|6|他使 黎巴嫩 跳躍如牛犢， 使 西連 跳躍如野牛犢。
PS|29|7|耶和華的聲音使火焰分岔。
PS|29|8|耶和華的聲音震動曠野， 耶和華震動 加低斯 的曠野。
PS|29|9|耶和華的聲音驚動母鹿落胎， 樹林也脫落淨光。 凡在他殿中的，都述說他的榮耀。
PS|29|10|耶和華坐在洪水之上為王； 耶和華坐著為王，直到永遠。
PS|29|11|耶和華必賜力量給他的百姓， 耶和華必賜平安的福給他的百姓。
PS|30|1|耶和華啊，我要尊崇你， 因為你救了我，不讓仇敵向我誇耀。
PS|30|2|耶和華－我的上帝啊， 我呼求你，你醫治了我。
PS|30|3|耶和華啊，你救我的性命脫離陰間， 使我存活，不至於下入地府。
PS|30|4|耶和華的聖民哪，你們要歌頌他， 要頌揚他神聖的名字 。
PS|30|5|因為，他的怒氣不過是轉眼之間； 他的恩典乃是一生之久。 一宿雖然有哭泣， 早晨便必歡呼。
PS|30|6|至於我，我凡事順利，就說： 「我永不動搖。」
PS|30|7|耶和華啊，你曾施恩，使我穩固如山； 你轉臉不顧，我就驚惶。
PS|30|8|耶和華啊，我曾求告你； 我向耶和華懇求：
PS|30|9|「我被害流血，下到地府，有何益處呢？ 塵土豈能稱謝你、傳揚你的信實嗎？
PS|30|10|耶和華啊，求你應允我，憐憫我！ 耶和華啊，求你幫助我！」
PS|30|11|你將我的哀哭變為跳舞， 脫去我的麻衣，為我披上喜樂，
PS|30|12|使我的靈 歌頌你，不致緘默。 耶和華－我的上帝啊，我要稱謝你，直到永遠！
PS|31|1|耶和華啊，我投靠你， 求你使我永不羞愧， 憑你的公義搭救我！
PS|31|2|求你側耳聽我， 快快救我！ 求你作我堅固的磐石， 拯救我的保障！
PS|31|3|你真是我的巖石、我的山寨， 求你為你名的緣故引導我，指教我。
PS|31|4|求你救我脫離人為我暗設的網羅， 因為你是我的保障。
PS|31|5|我將我的靈交在你手裏； 耶和華─信實的上帝啊，你救贖了我。
PS|31|6|我 恨惡那信奉虛無神明 的人； 我卻倚靠耶和華。
PS|31|7|我要因你的慈愛歡喜快樂， 因為你見過我的困苦， 知道我心中的艱難。
PS|31|8|你未曾把我交在仇敵手裏， 你使我的腳站在寬闊的地方。
PS|31|9|耶和華啊，求你憐憫我， 因為我在急難之中； 我的眼睛因憂愁而昏花， 我的身心也已耗盡。
PS|31|10|我的生命為愁苦所消耗， 我的年歲為嘆息所荒廢； 我的力量因我的罪孽 衰敗， 我的骨頭也枯乾。
PS|31|11|我因所有的敵人成了羞辱， 在我鄰舍跟前更加羞辱； 那認識我的都懼怕我， 在街上看見我的都躲避我。
PS|31|12|我被遺忘，如同死人，無人記念； 我好像破碎的器皿。
PS|31|13|我聽見許多人的毀謗， 四圍盡是驚嚇； 他們一同商議攻擊我， 圖謀害我的性命。
PS|31|14|耶和華啊，我仍要倚靠你； 我說：「你是我的上帝。」
PS|31|15|我終生的事在你手中， 求你救我脫離仇敵的手和那些迫害我的人。
PS|31|16|求你使你的臉向僕人發光， 憑你的慈愛拯救我。
PS|31|17|耶和華啊，求你叫我不致羞愧， 因為我曾呼求你； 求你使惡人羞愧， 使他們在陰間緘默無聲。
PS|31|18|那撒謊的人逞驕傲輕慢， 出狂妄的話攻擊義人， 願他的嘴啞而無言。
PS|31|19|在世人眼前， 你為敬畏你的人所積存的， 為投靠你的人所施行的， 是何等大的恩惠啊！
PS|31|20|你必將他們藏在你面前的隱密處， 免得遭人暗算； 你要隱藏他們在棚子裏， 免受口舌的爭鬧。
PS|31|21|耶和華是應當稱頌的， 因為我在圍城裏，他向我施展奇妙的慈愛。
PS|31|22|至於我，我曾驚惶地說： 「我從你眼前被隔絕。」 然而，我呼求你的時候， 你仍聽我懇求的聲音。
PS|31|23|耶和華的聖民哪，你們都要愛他！ 耶和華保護誠實可靠的人， 卻加倍報應行事驕傲的人。
PS|31|24|凡仰望耶和華的人， 你們都要壯膽，堅固你們的心！
PS|32|1|過犯得赦免， 罪惡蒙遮蓋的人有福了！
PS|32|2|耶和華不算為有罪， 內心沒有詭詐的人有福了！
PS|32|3|我閉口不認罪的時候， 因終日呻吟而骨頭枯乾。
PS|32|4|黑夜白日，你的手壓在我身上沉重； 我的精力耗盡 ，如同夏天的乾旱。（細拉）
PS|32|5|我向你陳明我的罪， 不隱瞞我的惡。 我說：「我要向耶和華承認我的過犯」； 你就赦免我的罪惡。（細拉）
PS|32|6|為此，凡虔誠人都當趁你可尋找 的時候向你禱告； 大水氾濫的時候，必不臨到他。
PS|32|7|你是我藏身之處， 你必保佑我脫離苦難， 以得救的歡呼 四面環繞我。（細拉）
PS|32|8|我要教導你，指示你當行的路， 我要定睛在你身上勸戒你。
PS|32|9|你不可像那無知的騾馬， 須用嚼環韁繩勒住， 不然，牠就不會靠近你。
PS|32|10|惡人必多受苦楚； 惟獨倚靠耶和華的，必有慈愛四面環繞他。
PS|32|11|義人哪，你們應當靠耶和華歡喜快樂， 心裏正直的人哪，你們都當歡呼。
PS|33|1|義人哪，你們當因耶和華歡呼， 正直人理當讚美耶和華。
PS|33|2|你們要彈琴稱謝耶和華， 用十弦瑟歌頌他。
PS|33|3|應當向他唱新歌， 彈得巧妙，聲音洪亮。
PS|33|4|因為耶和華的言語正直， 他的作為盡都信實。
PS|33|5|他喜愛公義和公平， 遍地滿了耶和華的慈愛。
PS|33|6|諸天藉耶和華的話而造， 萬象藉他口中的氣而成。
PS|33|7|他聚集海水如壘， 收藏深洋在倉庫。
PS|33|8|願全地都敬畏耶和華！ 願世上的居民都懼怕他！
PS|33|9|因為他說有，就有， 命立，就立。
PS|33|10|耶和華使列國的籌算歸於無有， 使萬民的計謀全無功效。
PS|33|11|耶和華的籌算永遠立定， 他心中的計劃萬代長存。
PS|33|12|以耶和華為上帝的，那國有福了！ 耶和華揀選為自己產業的，那民有福了！
PS|33|13|耶和華從天上觀看， 看見所有的人，
PS|33|14|從他的居所察看地上每一個居民，
PS|33|15|他塑造他們的心， 洞察他們一切的作為。
PS|33|16|君王不能因兵多得勝， 勇士不能因力大得救。
PS|33|17|靠馬得救是枉然的， 馬也不能因力大救人。
PS|33|18|看哪，耶和華的眼目看顧敬畏他的人 和仰望他慈愛的人，
PS|33|19|要救他們的性命脫離死亡， 使他們在饑荒中存活。
PS|33|20|我們的心向來等候耶和華； 他是我們的幫助，是我們的盾牌。
PS|33|21|我們的心必靠他歡喜， 因為我們向來倚靠他的聖名。
PS|33|22|耶和華啊，求你照著我們所仰望你的， 向我們施行慈愛！
PS|34|1|我要時時稱頌耶和華， 讚美他的話常在我口中。
PS|34|2|我的心必因耶和華誇耀， 謙卑的人聽見就喜樂。
PS|34|3|你們要和我一同尊耶和華為大， 讓我們一同高舉他的名。
PS|34|4|我曾尋求耶和華，他就應允我， 救我脫離一切的恐懼。
PS|34|5|仰望他的人，就有光榮； 他們 的臉必不蒙羞。
PS|34|6|這困苦人呼求，耶和華就垂聽， 救他脫離一切的患難。
PS|34|7|耶和華的使者在敬畏他的人四圍安營， 要搭救他們。
PS|34|8|你們要嘗嘗主恩的滋味，便知道他是美善； 投靠他的人有福了！
PS|34|9|耶和華的聖民哪，你們當敬畏他， 因敬畏他的一無所缺。
PS|34|10|少壯獅子尚且缺食忍餓， 但尋求耶和華的甚麼好處都不缺。
PS|34|11|孩子們哪，來聽我！ 我要將敬畏耶和華的道教導你們。
PS|34|12|有誰喜愛生命， 愛慕長壽，得享美福？
PS|34|13|你要禁止舌頭不出惡言， 嘴唇不說詭詐的話。
PS|34|14|要棄惡行善， 尋求和睦，一心追求。
PS|34|15|耶和華的眼目看顧義人， 他的耳朵聽他們的呼求。
PS|34|16|耶和華向行惡的人變臉， 要從地上除滅他們的名字 。
PS|34|17|義人呼求，耶和華聽見了， 就拯救他們脫離一切患難。
PS|34|18|耶和華靠近傷心的人， 拯救心靈痛悔的人。
PS|34|19|義人多有苦難， 但耶和華救他脫離這一切，
PS|34|20|又保護他全身的骨頭， 連一根也不折斷。
PS|34|21|惡必害死惡人， 恨惡義人的，必被定罪。
PS|34|22|耶和華救贖他僕人的性命， 凡投靠他的，必不致定罪。
PS|35|1|耶和華啊，與我相爭的，求你與他們相爭！ 與我爭戰的，求你與他們爭戰！
PS|35|2|求你拿著大小盾牌， 起來幫助我；
PS|35|3|舉起槍來，抵擋那追趕我的。 求你對我說：「我是拯救你的。」
PS|35|4|願那尋索我命的，蒙羞受辱！ 願那謀害我的，退後羞愧！
PS|35|5|願他們像風前的糠秕， 有耶和華的使者趕逐他們。
PS|35|6|願他們的道路又暗又滑， 有耶和華的使者追趕他們。
PS|35|7|因他們無故為我暗設網羅， 無故挖坑，要害我的命。
PS|35|8|願災禍忽然臨到他身上！ 願他暗設的網羅纏住自己！ 願他落在其中遭災禍！
PS|35|9|我的心必靠耶和華快樂， 靠他的救恩歡喜。
PS|35|10|我全身的骨頭要說： 「耶和華啊，誰能像你 救護困苦人脫離那比他強壯的， 救護困苦貧窮人脫離那搶奪他的？」
PS|35|11|兇惡的見證人起來， 盤問我所不知道的事。
PS|35|12|他們向我以惡報善， 使我喪失兒子。
PS|35|13|至於我，他們有病的時候， 我穿麻衣，禁食，刻苦己心； 我所求的都歸到自己身上。
PS|35|14|我如此行，好像他是我的朋友，我的兄弟； 我屈身悲哀，如同哀悼自己的母親。
PS|35|15|我在患難中，他們卻歡喜，大家聚集， 我所不認識的卑賤人 聚集攻擊我， 他們不住地撕裂我。
PS|35|16|他們試探我，不斷嘲笑我 ， 向我咬牙切齒。
PS|35|17|主啊，你看著不理要到幾時呢？ 求你救我的性命脫離他們的殘害， 救我僅有的 脫離少壯獅子！
PS|35|18|我在大會中要稱謝你， 在許多百姓中要讚美你。
PS|35|19|求你不容那無理與我為仇的向我誇耀！ 不容那無故恨我的向我瞪眼！
PS|35|20|因為他們不說平安， 倒想出詭詐的言語擾害地上安靜的人。
PS|35|21|他們大大張口攻擊我，說： 「啊哈，啊哈，我們已經親眼看見了！」
PS|35|22|耶和華啊，你已經看見了，求你不要沉默！ 主啊，求你不要遠離我！
PS|35|23|我的上帝─我的主啊，求你醒來，求你奮起， 還我公正，伸明我冤！
PS|35|24|耶和華－我的上帝啊，求你按你的公義判斷我， 不容他們向我誇耀！
PS|35|25|不容他們心裏說：「啊哈，遂我們的心願了！」 不容他們說：「我們已經把他吞了！」
PS|35|26|願那喜歡我遭難的一同抱愧蒙羞！ 願那向我妄自尊大的披戴慚愧，蒙受羞辱！
PS|35|27|願那喜悅我被判為義 的歡呼快樂； 願他們常說：「當尊耶和華為大！ 耶和華喜悅他的僕人平安。」
PS|35|28|我的舌頭要論說你的公義， 要常常讚美你。
PS|36|1|過犯在惡人的心底向他說話 ， 他的眼中不怕上帝。
PS|36|2|他自誇自媚， 以致罪孽無法察覺，不被恨惡。
PS|36|3|他口中的言語盡是罪孽詭詐， 他不再有智慧，也不再行善。
PS|36|4|他在床上圖謀罪孽， 定意行不善的道，不憎惡惡事。
PS|36|5|耶和華啊，你的慈愛上及諸天， 你的信實達到穹蒼，
PS|36|6|你的公義好像高山， 你的判斷如同深淵； 耶和華啊，人民、牲畜，你都救護。
PS|36|7|上帝啊，你的慈愛何其寶貴！ 世人投靠在你翅膀的蔭下。
PS|36|8|他們必因你殿裏的豐盛得以飽足， 你也必叫他們喝你那喜樂的泉水。
PS|36|9|因為在你那裏有生命的泉源， 在你的光中，我們必得見光。
PS|36|10|願你常施慈愛給認識你的人， 常以公義待心裏正直的人。
PS|36|11|不容驕傲人的腳踐踏我， 不容兇惡人的手趕逐我。
PS|36|12|在那裏，作惡的人已經仆倒； 他們被推倒，不能再起來。
PS|37|1|不要為作惡的心懷不平， 也不要嫉妒那行不義的人。
PS|37|2|因為他們如草快被割下， 又如綠色的嫩草快要枯乾。
PS|37|3|你當倚靠耶和華而行善， 安居地上，以他的信實為糧；
PS|37|4|又當以耶和華為樂， 他就將你心裏所求的賜給你。
PS|37|5|當將你的道路交託耶和華， 並倚靠他，他就必成全。
PS|37|6|他要使你的公義如光發出， 使你的公平明如正午。
PS|37|7|你當安心倚靠耶和華，耐性等候他， 不要因那道路通達的和那惡謀成就的心懷不平。
PS|37|8|當止住怒氣，離棄憤怒； 不要心懷不平，以致作惡。
PS|37|9|因為作惡的必被剪除； 惟有等候耶和華的必承受土地。
PS|37|10|還有片時，惡人要歸於無有； 你就是細察他的住處，也不存在。
PS|37|11|但謙卑的人必承受土地， 以豐盛的平安為樂。
PS|37|12|惡人設謀要害義人， 向他咬牙。
PS|37|13|但主必笑他， 因見他受罰的日子將要來到。
PS|37|14|惡人刀已出鞘，弓已上弦， 要砍倒困苦貧窮的人， 要殺害行為正直的人。
PS|37|15|他們的刀必刺入自己的心， 他們的弓必折斷。
PS|37|16|一個義人所有的雖少， 強過許多惡人的富餘。
PS|37|17|因為惡人的膀臂必折斷； 但耶和華扶持義人。
PS|37|18|耶和華知道完全人的日子， 他們的產業要存到永遠。
PS|37|19|他們在患難的時候必不致羞愧， 在饑荒的日子必得飽足。
PS|37|20|惡人卻要滅亡。 耶和華的仇敵要像草地的華美 ； 他們要毀滅，在煙中消失 。
PS|37|21|惡人借貸卻不償還； 義人恩待人，並且施捨。
PS|37|22|蒙耶和華賜福的必承受土地； 他所詛咒的必被剪除。
PS|37|23|義人的腳步為耶和華所穩定； 他的道路，耶和華也喜愛。
PS|37|24|他雖失腳也不致全身仆倒， 因為耶和華攙扶他的手。
PS|37|25|我從前年幼，現在年老， 卻未見過義人被棄， 也未見過他的後裔求乞。
PS|37|26|他常常恩待人，借貸給人， 他的後裔也必蒙福。
PS|37|27|你當離惡行善， 就可永遠安居。
PS|37|28|因為耶和華喜愛公平， 不撇棄他的聖民， 他們永蒙保佑； 但惡人的後裔必被剪除。
PS|37|29|義人必承受土地， 永居其上。
PS|37|30|義人的口發出智慧， 他的舌頭講說公平。
PS|37|31|上帝的律法在他心裏， 他的步伐總不搖動。
PS|37|32|惡人窺探義人， 想要殺他。
PS|37|33|耶和華必不把他交在惡人手中， 當審判的時候，也不定他的罪。
PS|37|34|你當等候耶和華，遵守他的道， 他就抬舉你，使你承受土地； 你必看到惡人被剪除。
PS|37|35|我見過惡人大有勢力， 高聳如本地青翠的樹木。
PS|37|36|有人 從那裏經過，看哪，他已不存在， 我尋找他，卻尋不著了。
PS|37|37|你要細察那完全人，觀看那正直人， 因為和平的人有好結局。
PS|37|38|至於罪人，必一同滅絕， 惡人的結局必被剪除。
PS|37|39|義人得救是出於耶和華， 在患難時耶和華作他們的避難所。
PS|37|40|耶和華幫助他們，解救他們； 他解救他們脫離惡人，把他們救出來， 因為他們投靠他。
PS|38|1|耶和華啊，求你不要在怒中責備我， 不要在烈怒中懲罰我！
PS|38|2|因為你的箭射入我身， 你的手壓住我。
PS|38|3|因你的惱怒，我的肉無一完全； 因我的罪過，我的骨頭也不安寧。
PS|38|4|我的罪孽高過我的頭， 如同重擔叫我擔當不起。
PS|38|5|因我的愚昧， 我的傷發臭流膿。
PS|38|6|我疼痛，大大蜷曲， 整日哀痛。
PS|38|7|我滿腰灼熱， 我的肉無一完全。
PS|38|8|我被壓碎，身心虛弱； 因心裏痛苦，我就呻吟。
PS|38|9|主啊，我的心願都在你面前， 我的嘆息不向你隱瞞。
PS|38|10|我心顫慄，體力衰微， 眼中無光。
PS|38|11|我遭遇災病，良朋密友都袖手旁觀， 我的親戚本家也遠遠站立。
PS|38|12|那尋索我命的設下羅網， 那想要害我的口出惡言， 整日思想詭計。
PS|38|13|但我如聾子聽不見， 像啞巴不能開口。
PS|38|14|我如聽不見的人， 無法用口答辯。
PS|38|15|耶和華啊，我仰望你！ 主－我的上帝啊，你必應允我！
PS|38|16|我曾說：「恐怕他們向我誇耀， 我失腳的時候，他們向我誇口。」
PS|38|17|我就要跌倒， 我的痛苦常在我面前。
PS|38|18|我要承認我的罪孽， 要因我的罪憂愁。
PS|38|19|但我的仇敵又活潑又強壯， 無理恨我的增多了。
PS|38|20|以惡報善的與我作對， 但我追求良善。
PS|38|21|耶和華啊，求你不要撇棄我！ 我的上帝啊，求你不要遠離我！
PS|38|22|拯救我的主啊， 求你快快幫助我！
PS|39|1|我曾說：「我要謹慎我的言行， 免得我的舌頭犯罪； 惡人在我面前的時候， 我要用嚼環勒住我的口。」
PS|39|2|我默然無聲，連好話也不出口， 我的愁苦就更加深。
PS|39|3|我的心在我裏面發熱； 我默想的時候，火就燒起， 我用舌頭說話：
PS|39|4|「耶和華啊，求你讓我曉得我的結局， 我的壽數幾何， 使我知道我的生命何等短暫！
PS|39|5|看哪，你使我的年日窄如手掌， 我一生的年數，在你面前如同無有； 各人最穩妥的時候，真是全然虛幻。（細拉）
PS|39|6|世人行動實係幻影， 他們忙亂，真是枉然， 積蓄財寶，不知將來有誰收取。
PS|39|7|「主啊，如今我等甚麼呢？ 我的指望在乎你！
PS|39|8|求你救我脫離一切的過犯， 不要使我受愚頑人的羞辱。
PS|39|9|我保持沉默，閉口不言， 因為這一切都是你所做的。
PS|39|10|求你從我身上免去你的責罰； 因你手的責打，我就消滅。
PS|39|11|因人的罪惡你懲罰管教他的時候， 如蛀蟲一般，吃掉他所喜愛的。 世人真是虛幻！（細拉）
PS|39|12|「耶和華啊，求你聽我的禱告， 側耳聽我的呼求！ 我流淚，求你不要靜默無聲！ 因為在你面前我是客旅， 是寄居的，像我列祖一般。
PS|39|13|求你寬容我， 使我在去而不返之先可以喜樂。」
PS|40|1|我曾耐性等候耶和華， 他垂聽我的呼求。
PS|40|2|他從泥坑裏， 從淤泥中，把我拉上來， 使我的腳立在磐石上， 使我腳步穩健。
PS|40|3|他使我口唱新歌， 就是讚美我們上帝的話。 許多人必看見而懼怕， 並要倚靠耶和華。
PS|40|4|那倚靠耶和華、 不理會狂傲和偏向虛假的， 這人有福了！
PS|40|5|耶和華－我的上帝啊，你所行的奇事 和你為我們設想的計劃，多到無法盡述； 若要述說陳明，不可勝數。
PS|40|6|祭物和禮物，你不喜愛， 你已經開通我的耳朵； 燔祭和贖罪祭非你所要。
PS|40|7|那時我說：「看哪，我來了！ 我的事在經卷上已經記載了。
PS|40|8|我的上帝啊，我樂意照你的旨意行， 你的律法在我心裏。」
PS|40|9|我在大會中傳講公義的佳音， 看哪，必不制止我的嘴唇； 耶和華啊，這一切你都知道。
PS|40|10|我未曾把你的公義藏在心裏， 我已陳明你的信實和你的救恩； 在大會中我未曾隱瞞你的慈愛和信實。
PS|40|11|耶和華啊，求你不要向我止住你的憐憫！ 願你的慈愛和信實常常保佑我！
PS|40|12|因有無數的禍患圍困我， 我的罪孽追上了我，使我不能看見， 這罪孽比我的頭髮還多， 我的膽量喪失了。
PS|40|13|耶和華啊，求你開恩搭救我！ 耶和華啊，求你速速幫助我！
PS|40|14|願那些尋找我、要滅我命的，一同抱愧蒙羞！ 願那些喜悅我遭害的，退後受辱！
PS|40|15|願那些對我說「啊哈、啊哈」的， 因羞愧而敗亡！
PS|40|16|願一切尋求你的，因你歡喜快樂！ 願那些喜愛你救恩的，常說：「當尊耶和華為大！」
PS|40|17|我本是困苦貧窮的，主卻顧念我。 你是幫助我的，搭救我的； 我的上帝啊，求你不要耽延！
PS|41|1|眷顧貧寒人的有福了 ！ 在患難的日子，耶和華必搭救他。
PS|41|2|耶和華必保全他，使他存活， 他要在地上享福。 求你不要把他交給仇敵，遂其所願。
PS|41|3|他病重在榻，耶和華必扶持他； 他在病中，你必使他離開病床。
PS|41|4|我曾說：「耶和華啊，求你憐憫我， 醫治我，因為我得罪了你。」
PS|41|5|我的仇敵用惡言議論我： 「他幾時才會死，他的名幾時才會消滅呢？」
PS|41|6|當他來看我的時候，說的是假話； 他心存奸惡，走到外邊才說出來。
PS|41|7|所有恨我的，都一同交頭接耳議論我， 他們設計要害我。
PS|41|8|他們說：「他有怪病纏身， 他已躺下，必不能再起來。」
PS|41|9|連我知己的朋友， 我所信賴、吃我飯的人也用腳踢我。
PS|41|10|耶和華啊，求你憐憫我， 使我起來，好報復他們！
PS|41|11|我因此就知道你喜愛我， 我的仇敵不得向我誇勝。
PS|41|12|你因我純正就扶持我， 使我永遠站立在你面前。
PS|41|13|耶和華－ 以色列 的上帝是應當稱頌的， 從亙古直到永遠。阿們！阿們！ 可拉後裔的詩。交給聖詠團長。
PS|42|1|上帝啊，我的心切慕你， 如鹿切慕溪水。
PS|42|2|我的心渴想上帝，就是永生上帝， 我幾時得朝見上帝呢？
PS|42|3|我晝夜以眼淚當食物， 人不住地對我說：「你的上帝在哪裏呢？」
PS|42|4|我從前與眾人同往， 領他們到上帝的殿裏， 大家用歡呼稱頌的聲音守節； 我追想這些事， 我的心極其悲傷。
PS|42|5|我的心哪，你為何憂悶？ 為何在我裏面煩躁？ 應當仰望上帝， 因我還要稱謝他，我當面的拯救，
PS|42|6|我的上帝。我的心在我裏面憂悶， 所以我從 約旦 地， 從 黑門嶺 ，從 米薩山 記念你。
PS|42|7|你的瀑布發聲，深淵就與深淵響應， 你的波浪洪濤漫過我身。
PS|42|8|白晝，耶和華必施慈愛； 黑夜，我要歌頌祈禱賜我生命的上帝。
PS|42|9|我要對上帝－我的磐石說： 「你為何忘記我呢？ 我為何因仇敵的欺壓時常哀痛呢？」
PS|42|10|我的敵人辱罵我， 好像敲碎我的骨頭， 他們不住地對我說： 「你的上帝在哪裏呢？」
PS|42|11|我的心哪，你為何憂悶？ 為何在我裏面煩躁？ 應當仰望上帝， 因我還要稱謝他，我當面的拯救，我的上帝。
PS|43|1|上帝啊，求你為我伸冤， 向不虔誠的國為我辯護； 求你救我脫離詭詐不義的人。
PS|43|2|你是作我保障 的上帝，為何丟棄我呢？ 我為何因仇敵的欺壓時常哀痛呢？
PS|43|3|求你發出你的亮光和信實，好引導我， 帶我到你的聖山，到你的居所！
PS|43|4|我就走到上帝的祭壇， 到賜我喜樂的上帝那裏。 上帝，我的上帝啊， 我要彈琴稱謝你！
PS|43|5|我的心哪，你為何憂悶？ 為何在我裏面煩躁？ 應當仰望上帝， 我還要稱謝他，我當面的拯救，我的上帝。
PS|44|1|上帝啊，你在古時， 我們列祖的日子所做的事， 我們親耳聽見了， 我們的列祖曾為我們述說。
PS|44|2|你曾用手趕出外邦人， 卻栽培了我們的列祖； 你苦待萬民， 卻叫我們的列祖發達。
PS|44|3|因為他們不是靠自己的刀劍承受土地， 也不是靠自己的膀臂得勝， 而是靠你的右手、你的膀臂， 和你臉上的亮光， 因為你喜愛他們。
PS|44|4|上帝啊，你是我的君王， 求你發命令使 雅各 得勝。
PS|44|5|靠你，我們要推倒我們的敵人； 靠你的名，我們要踐踏那興起攻擊我們的人。
PS|44|6|因為我必不倚靠我的弓， 我的刀也不能使我得勝。
PS|44|7|惟有你拯救我們脫離敵人， 使恨我們的人羞愧。
PS|44|8|我們要常常因上帝誇耀， 要永遠頌揚你的名。（細拉）
PS|44|9|但如今你丟棄了我們，使我們受辱， 不和我們的軍隊同去。
PS|44|10|你使我們在敵人前轉身撤退， 使那恨我們的人任意搶奪。
PS|44|11|你使我們如羊當作食物， 把我們分散在列國中。
PS|44|12|你賣了你的子民也不獲利， 所得的並未加添你的資財。
PS|44|13|你使我們受鄰國的羞辱， 被四圍的人嗤笑譏諷。
PS|44|14|你使我們在列國中成了笑柄， 在萬民中使人搖頭。
PS|44|15|因辱罵者和毀謗者的聲音， 因仇敵和報仇者的緣故， 我的凌辱常常在我面前， 我臉上的羞愧將我遮蔽，
PS|44|16|
PS|44|17|這些事都臨到我們身上， 我們卻沒有忘記你， 也沒有違背你的約；
PS|44|18|我們的心並未退縮， 我們的腳也沒有偏離你的路。
PS|44|19|你在野狗出沒之處壓傷我們， 以死蔭籠罩我們。
PS|44|20|倘若我們忘記上帝的名， 或向外邦神明舉手，
PS|44|21|上帝豈不鑒察這事嗎？ 因為他曉得人心裏的隱祕。
PS|44|22|我們為你的緣故終日被殺， 人看我們如將宰的羊。
PS|44|23|主啊，求你睡醒，為何儘睡呢？ 求你醒來，不要永遠丟棄我們！
PS|44|24|你為何轉臉， 不顧我們所遭的苦難和所受的欺壓呢？
PS|44|25|我們俯伏在塵土上， 我們的肚腹緊貼地面。
PS|44|26|求你興起幫助我們！ 因你的慈愛救贖我們！
PS|45|1|我心裏湧出美辭， 我為王朗誦我的詩章， 我的舌頭是敏捷文士的手筆。
PS|45|2|你比世人更美， 你嘴裏滿有恩惠； 所以上帝賜福給你，直到永遠。
PS|45|3|勇士啊，願你腰間佩刀， 大展榮耀和威嚴，
PS|45|4|為真理、謙卑、公義威嚴地駕車前進，無不得勝； 願你的右手顯明可畏的事。
PS|45|5|你的箭鋒快，射中王的仇敵的心， 萬民仆倒在你之下。
PS|45|6|上帝啊，你的寶座是永永遠遠的， 你國度的權杖是正直的權杖。
PS|45|7|你喜愛公義，恨惡罪惡， 所以上帝，就是你的上帝，用喜樂油膏你， 勝過膏你的同伴。
PS|45|8|你的衣服散發沒藥、沉香、肉桂的香氣， 象牙宮中絲弦樂器的聲音使你歡喜。
PS|45|9|你的妃嬪之中有列王的女兒， 王后佩戴 俄斐 金飾站立在你右邊。
PS|45|10|女子啊，要傾聽，要思想，要側耳而聽！ 不要記念你本族和你父家，
PS|45|11|王就羨慕你的美貌； 因為他是你的主，你當向他下拜。
PS|45|12|推羅 必來送禮， 百姓中富足的人也必向你求恩。
PS|45|13|君王的女兒在宮裏極其榮華， 她的衣服是金線繡的；
PS|45|14|她穿錦繡的衣服，引到王面前， 陪伴她的童女隨從她，也被帶到你面前。
PS|45|15|她們要歡喜快樂， 被引導進入王宮。
PS|45|16|你的子孫要接續你列祖， 你要立他們在各地作王。
PS|45|17|我必使萬代記念你的名， 萬民要永永遠遠稱謝你。
PS|46|1|上帝是我們的避難所，是我們的力量， 是我們在患難中隨時的幫助。
PS|46|2|所以，地雖改變， 山雖搖動到海心，
PS|46|3|其中的水雖澎湃翻騰， 山雖因海漲而戰抖， 我們也不害怕。（細拉）
PS|46|4|有一道河，這河的分汊使上帝的城歡喜， 這城就是至高者居住的聖所。
PS|46|5|上帝在其中，城必不動搖； 到天一亮，上帝必幫助這城。
PS|46|6|萬邦喧嚷，國度動搖； 上帝出聲，地就熔化。
PS|46|7|萬軍之耶和華與我們同在， 雅各 的上帝是我們的避難所！（細拉）
PS|46|8|你們來看耶和華的作為， 看他使地怎樣荒涼。
PS|46|9|他止息戰爭，直到地極； 他折弓、斷槍，把戰車焚燒在火中。
PS|46|10|你們要休息，要知道我是上帝！ 我必在列國中受尊崇，在全地也受尊崇。
PS|46|11|萬軍之耶和華與我們同在， 雅各 的上帝是我們的避難所！
PS|47|1|萬民哪，你們都要鼓掌！ 用歡呼的聲音向上帝呼喊！
PS|47|2|因為耶和華至高者是可畏的， 他是治理全地的大君王。
PS|47|3|他使萬民服在我們以下， 又使萬族服在我們腳下。
PS|47|4|他為我們選擇產業， 就是他所愛之 雅各 的榮耀。（細拉）
PS|47|5|上帝上升，有喊聲相送； 耶和華上升，有角聲相送。
PS|47|6|你們要向上帝歌頌，歌頌！ 向我們的王歌頌，歌頌！
PS|47|7|因為上帝是全地的王， 你們要用聖詩歌頌！
PS|47|8|上帝作王治理列國， 上帝坐在他的聖寶座上。
PS|47|9|萬民的君王聚集， 要作 亞伯拉罕 的上帝的子民， 因為地上的盾牌是屬上帝的， 他為至高！
PS|48|1|耶和華本為大！ 在我們上帝的城中， 在他的聖山上， 當受大讚美。
PS|48|2|錫安山 －大君王的城， 在北面居高華美， 為全地所喜悅。
PS|48|3|上帝在城的宮殿中， 自顯為避難所。
PS|48|4|看哪，諸王會合， 一同經過。
PS|48|5|他們見了這城就驚奇喪膽， 急忙逃跑。
PS|48|6|戰兢在那裏抓住他們， 他們好像臨產的婦人一樣陣痛。
PS|48|7|上帝啊，你用東風擊破 他施 的船隻。
PS|48|8|我們在萬軍之耶和華的城裏， 就是我們上帝的城裏， 所看見的正如我們所聽見的。 上帝必堅立這城，直到永遠。（細拉）
PS|48|9|上帝啊，我們在你的殿中 想念你的慈愛。
PS|48|10|上帝啊，你受的讚美正與你的名相稱，直到地極！ 你的右手滿了公義。
PS|48|11|因你的判斷， 錫安山 應當歡喜， 猶大 的城鎮 應當快樂。
PS|48|12|你們當周遊 錫安 ， 四圍環繞，數點城樓，
PS|48|13|細看它的城郭， 察看它的宮殿， 為要傳揚給後代。
PS|48|14|因為這上帝永永遠遠為我們的上帝， 他必作我們引路的，直到死時 。
PS|49|1|萬民哪，你們都當聽這話！ 世上所有的居民， 無論貴賤貧富， 都當側耳而聽！
PS|49|2|
PS|49|3|我口要說智慧的言語， 我心思想通達的道理。
PS|49|4|我要側耳聽比喻， 用琴解謎語。
PS|49|5|在患難的日子，追逼我的人的奸惡 環繞我， 我何必懼怕？
PS|49|6|他們那些倚靠財貨， 自誇錢財多的人，
PS|49|7|沒有一個能贖自己的弟兄 ， 能將贖價給上帝，
PS|49|8|讓他長遠活著，不見地府 ； 因為贖生命的價值極貴， 只可永遠罷休。
PS|49|9|
PS|49|10|他要見智慧人死， 愚昧人和畜牲一般的人一同滅亡， 把他們的財貨留給別人。
PS|49|11|他們雖以自己的名叫自己的地， 墳墓卻作他們永遠的家， 作他們世世代代的居所。
PS|49|12|人居尊貴中不能長久， 如同死亡的畜類一樣。
PS|49|13|他們所行之道本為自己的愚昧， 後來的人卻還佩服他們的話語。（細拉）
PS|49|14|他們如同羊群註定要下陰間， 死亡必作他們的牧者； 到了早晨，正直人必管轄他們。 他們的形像必被陰間所滅，無處可容身。
PS|49|15|然而上帝必救贖我的命脫離陰間的掌控， 因他必收納我。（細拉）
PS|49|16|見人發財、家室日益顯赫的時候， 你不要懼怕；
PS|49|17|因為他死的時候甚麼也不能帶去， 他的榮耀不能隨他下去。
PS|49|18|他活著的時候，雖然自誇為有福 ─你若自己行得好，人必誇獎你─
PS|49|19|他仍必與歷代的祖宗一樣同歸死亡， 永不見光。
PS|49|20|人在尊貴中而不醒悟， 就如死亡的畜類一樣。
PS|50|1|大能者上帝－耶和華已經發言呼召天下， 從日出之地到日落之處。
PS|50|2|從全然美麗的 錫安 中， 上帝已經發光了。
PS|50|3|我們的上帝要來，絕不閉口； 有烈火在他面前吞滅， 有暴風在他四圍颳起。
PS|50|4|他呼召上天下地， 為要審判他的子民：
PS|50|5|「召集我的聖民， 就是那些用祭物與我立約的人，到我這裏來。」
PS|50|6|諸天必表明他的公義， 因為上帝是施行審判的。（細拉）
PS|50|7|「聽啊，我的子民，我要說話！ 以色列 啊，我要審問你； 我是上帝，是你的上帝！
PS|50|8|我並不因你的祭物責備你； 你的燔祭常在我面前。
PS|50|9|我不從你家中取公牛， 也不從你圈內取公山羊；
PS|50|10|因為，林中的百獸是我的， 千山的牲畜也是我的。
PS|50|11|山中 的飛鳥，我都知道， 田野的走獸也都屬我。
PS|50|12|「我若是飢餓，不用告訴你， 因為世界和其中所充滿的都是我的。
PS|50|13|我豈吃公牛的肉呢？ 我豈喝公山羊的血呢？
PS|50|14|你們要以感謝為祭獻給上帝， 又要向至高者還你的願，
PS|50|15|並要在患難之日求告我， 我必搭救你，你也要榮耀我。」
PS|50|16|但上帝對惡人說：「你怎敢傳講我的律例， 口中提到我的約呢？
PS|50|17|其實你恨惡管教， 將我的言語拋在腦後。
PS|50|18|你見了盜賊就樂意與他同夥， 又和行姦淫的人同流合污。
PS|50|19|「你的口出惡言， 你的舌編造詭詐。
PS|50|20|你坐著，毀謗你的兄弟， 讒害你親母的兒子。
PS|50|21|你做了這些事，我閉口不言， 你想我正如你一樣； 其實我要責備你，將這些事擺在你眼前。
PS|50|22|「你們忘記上帝的，要思想這事， 免得我把你們撕碎，無人搭救。
PS|50|23|凡以感謝獻祭的就是榮耀我； 那按正路而行的，我必使他得著上帝的救恩。」
PS|51|1|上帝啊，求你按你的慈愛恩待我！ 按你豐盛的憐憫塗去我的過犯！
PS|51|2|求你將我的罪孽洗滌淨盡， 潔除我的罪！
PS|51|3|因為我知道我的過犯； 我的罪常在我面前。
PS|51|4|我向你犯罪，惟獨得罪了你， 在你眼前行了這惡， 以致你責備的時候顯為公義， 判斷的時候顯為清白。
PS|51|5|看哪，我是在罪孽裏生的， 在我母親懷胎的時候就有了罪。
PS|51|6|你所喜愛的是內心的誠實； 求你在我隱密處使我得智慧。
PS|51|7|求你用牛膝草潔淨我，我就乾淨； 求你洗滌我，我就比雪更白。
PS|51|8|求你使我得聽歡喜快樂的聲音， 使你所壓傷的骨頭可以踴躍。
PS|51|9|求你轉臉不看我的罪， 塗去我一切的罪孽。
PS|51|10|上帝啊，求你為我造清潔的心， 使我裏面重新有正直 的靈。
PS|51|11|不要丟棄我，使我離開你的面； 不要從我收回你的聖靈。
PS|51|12|求你使我重得救恩之樂， 以樂意的靈來扶持我，
PS|51|13|我就把你的道指教有過犯的人， 罪人必歸順你。
PS|51|14|上帝啊，你是拯救我的上帝； 求你救我脫離流人血的罪！ 我的舌頭就高唱你的公義。
PS|51|15|主啊，求你使我嘴唇張開， 我的口就傳揚讚美你的話！
PS|51|16|你本不喜愛祭物，若喜愛，我就獻上； 燔祭你也不喜悅。
PS|51|17|上帝所要的祭就是憂傷的靈； 上帝啊，憂傷痛悔的心，你必不輕看。
PS|51|18|求你隨你的美意善待 錫安 ， 建造 耶路撒冷 的城牆。
PS|51|19|那時，你必喜愛公義的祭 和燔祭，全牲的燔祭； 那時，人必將公牛獻在你壇上。
PS|52|1|勇士啊，你為何作惡自誇？ 上帝的慈愛是常存的。
PS|52|2|你這行詭詐的人哪， 你的舌頭像快利的剃刀，圖謀毀滅。
PS|52|3|你愛惡勝似愛善， 又愛說謊，勝於愛說公義。（細拉）
PS|52|4|詭詐的舌頭啊， 你愛說一切毀滅的話！
PS|52|5|上帝也要毀滅你，直到永遠。 他要抓住你，從帳棚中拉你出來， 從活人之地將你拔除。（細拉）
PS|52|6|義人要看見而懼怕， 並要笑他。
PS|52|7|看哪，這就是那不以上帝為保障的人， 他只倚靠豐富的財物，在邪惡上堅立自己。
PS|52|8|至於我，就像上帝殿中的青橄欖樹， 我永永遠遠倚靠上帝的慈愛。
PS|52|9|我要稱謝你，直到永遠， 因為你做了這事。 我也要在你聖民面前仰望你的名， 這名本為美好。
PS|53|1|愚頑人心裏說：「沒有上帝。」 他們都敗壞，行了可憎惡的罪孽， 沒有一個人行善。
PS|53|2|上帝從天上垂看世人， 要看有明白的沒有， 有尋求上帝的沒有。
PS|53|3|他們全都退後，一同變為污穢， 沒有行善的， 連一個也沒有。
PS|53|4|作惡的都沒有知識嗎？ 他們吞吃我的百姓如同吃飯一樣， 並不求告上帝。
PS|53|5|他們在無可懼怕之處就大大害怕， 因為上帝使那安營攻擊你之人的骨頭散開了。 你使他們蒙羞，因為上帝棄絕了他們。
PS|53|6|但願 以色列 的救恩出自 錫安 。 當上帝救回他被擄子民的時候， 雅各 要快樂， 以色列 要歡喜。
PS|54|1|上帝啊，求你因你的名拯救我， 憑你的大能為我伸冤。
PS|54|2|上帝啊，求你聽我的禱告， 側耳聽我口中的言語。
PS|54|3|因為陌生人興起攻擊我， 強橫的人尋索我的性命； 他們眼中沒有上帝。（細拉）
PS|54|4|看哪，上帝是幫助我的， 主是扶持我性命的，
PS|54|5|他要報應我仇敵所作的惡； 求你憑你的信實滅絕他們。
PS|54|6|我要把甘心祭獻給你； 耶和華啊，我要頌揚你的名，這名本為美好。
PS|54|7|他從一切的急難中把我救出來， 我的眼睛也看見了我的仇敵遭報。
PS|55|1|上帝啊，求你側耳聽我的禱告， 不要隱藏不聽我的懇求！
PS|55|2|求你留心聽我，應允我。 我哀嘆不安，發出呻吟，
PS|55|3|都因仇敵的聲音，惡人的欺壓； 他們將罪孽加在我身上，發怒氣加害我。
PS|55|4|我的心在我裏面陣痛， 死亡的恐怖落在我身。
PS|55|5|恐懼戰兢臨到了我， 驚恐籠罩我。
PS|55|6|我說：「但願我有翅膀像鴿子， 我就飛去，得享安息。
PS|55|7|看哪，我要遠走高飛， 宿在曠野。（細拉）
PS|55|8|我要速速逃到避難之所， 脫離狂風暴雨。」
PS|55|9|主啊，求你吞滅他們，變亂他們的言語！ 因為我在城中見了兇暴爭吵的事。
PS|55|10|他們晝夜在城牆上繞行， 城內也有罪孽和奸惡。
PS|55|11|邪惡在其中， 欺壓和詭詐不離街市。
PS|55|12|原來，不是仇敵辱罵我， 若是仇敵，還可忍受； 也不是恨我的人向我狂妄自大， 若是恨我的人，我必躲避他。
PS|55|13|不料是你；你原與我同等， 是我的朋友，是我的知己！
PS|55|14|我們素常彼此交談，以為甘甜； 我們結伴在上帝的殿中同行。
PS|55|15|願死亡忽然臨到他們！ 願他們活生生地下入陰間！ 因為他們的住處都是邪惡， 他們的內心充滿奸惡。
PS|55|16|至於我，我要求告上帝， 耶和華必拯救我。
PS|55|17|晚上、早晨、中午我要哀聲悲嘆， 他就垂聽我的聲音。
PS|55|18|他救贖我的命脫離攻擊我的人， 使我得享平安， 因為與我相爭的人很多。
PS|55|19|那不願改變、不敬畏上帝的人， 從太古常存的上帝必聽見而使他受苦。（細拉）
PS|55|20|他背了約， 伸手攻擊與他和好的人。
PS|55|21|他的口如奶油光滑， 他的心卻懷著敵意； 他的話比油柔和， 其實是拔出的刀。
PS|55|22|你要把你的重擔卸給耶和華， 他必扶持你， 他永不叫義人動搖。
PS|55|23|上帝啊，你必使惡人墜入滅亡的坑； 那好流人血、行詭詐的人必活不過半生， 但我要倚靠你。
PS|56|1|上帝啊，求你憐憫我，因為有人踐踏我， 終日攻擊欺壓我。
PS|56|2|我的仇敵終日踐踏我， 逞驕傲攻擊我的人很多。
PS|56|3|我懼怕的時候要倚靠你。
PS|56|4|我倚靠上帝，我要讚美他的話語； 我倚靠上帝，必不懼怕。 血肉之軀能把我怎麼樣呢？
PS|56|5|他們終日扭曲我的話， 千方百計加害於我。
PS|56|6|他們聚集，埋伏，窺探我的腳蹤， 等候要害我的命。
PS|56|7|他們豈能脫罪呢 ？ 上帝啊，求你在怒中使萬民敗落！
PS|56|8|我幾次流離，你都數算； 求你把我的眼淚裝在你的皮袋裏。 這一切不都記在你的冊子上嗎？
PS|56|9|我呼求的日子，仇敵都要轉身撤退。 上帝幫助我，這是我所知道的。
PS|56|10|我倚靠上帝，我要讚美他的話語； 我倚靠耶和華，我要讚美他的話語。
PS|56|11|我倚靠上帝，必不懼怕。 人能把我怎麼樣呢？
PS|56|12|上帝啊，我要向你還所許的願， 我要以感謝祭回報你；
PS|56|13|因為你救我的命脫離死亡。 你保護我的腳不跌倒， 使我在生命的光中行在上帝面前。
PS|57|1|上帝啊，求你憐憫我，憐憫我， 因為我的心投靠你。 我要投靠在你翅膀蔭下， 直等到災害過去。
PS|57|2|我要求告至高的上帝， 就是為我成全萬事的上帝。
PS|57|3|那踐踏我的人辱罵我的時候， 上帝必從天上施恩救我，(細拉) 他必向我施行慈愛和信實。
PS|57|4|至於我的性命， 我好像躺臥在吞噬人的獅子當中； 他們的牙齒是槍、箭， 他們的舌頭是快刀。
PS|57|5|上帝啊，願你崇高過於諸天！ 願你的榮耀高過全地！
PS|57|6|他們為我的腳設下網羅，壓迫我； 他們在我面前掘了坑，自己反掉在其中。（細拉）
PS|57|7|上帝啊，我心堅定，我心堅定； 我要唱詩，我要歌頌！
PS|57|8|我的靈 啊，你當醒起！ 琴瑟啊，當醒起！ 我自己要極早醒起！
PS|57|9|主啊，我要在萬民中稱謝你， 在萬族中歌頌你！
PS|57|10|因為你的慈愛高及諸天， 你的信實達到穹蒼。
PS|57|11|上帝啊，願你崇高過於諸天！ 願你的榮耀高過全地！
PS|58|1|你們緘默不語，真合公義嗎？ 你們審判世人，豈按正直嗎？
PS|58|2|不然！你們心中作惡， 量出你們在地上手中的殘暴。
PS|58|3|惡人一出母胎就與上帝疏遠， 一離母腹就走錯路，說謊話。
PS|58|4|他們的毒氣好像蛇的毒氣， 他們好像聾的毒蛇塞住耳朵，
PS|58|5|聽不見弄蛇者的聲音， 也聽不見魔術師的咒語。
PS|58|6|上帝啊，求你敲碎他們口中的牙！ 耶和華啊，求你敲掉少壯獅子的大牙！
PS|58|7|願他們消滅，如急流的水一般； 他們瞄準射箭的時候，箭頭彷彿折斷。
PS|58|8|願他們像蝸牛腐爛消失， 又像婦人流掉的胎兒，未見天日。
PS|58|9|你們用荊棘燒火，鍋還未熱， 上帝就用旋風把未燒著的和已燒著的一齊颳去。
PS|58|10|義人見仇敵遭報就歡喜， 他要在惡人的血中洗腳。
PS|58|11|因此，人必說：「義人誠然有善報， 在地上果然有施行審判的上帝！」
PS|59|1|我的上帝啊，求你救我脫離仇敵， 把我安置在高處，脫離那些起來攻擊我的人。
PS|59|2|求你救我脫離作惡的人， 救我脫離好流人血的人！
PS|59|3|因為他們埋伏要害我命， 強悍的人聚集攻擊我， 耶和華啊，不是為我的過犯， 也不是為我的罪愆。
PS|59|4|我雖然無過，他們急忙擺陣攻擊我。 求你興起，來幫助我，來鑒察！
PS|59|5|萬軍之耶和華上帝－ 以色列 的上帝啊， 求你醒起，懲治萬國！ 不要憐憫行詭詐的惡人！（細拉）
PS|59|6|他們晚上轉回， 叫號如狗，圍城繞行。
PS|59|7|看哪，他們口中噴吐惡言， 嘴裏有刀： 「有誰聽見呢？」
PS|59|8|但你－耶和華必譏笑他們， 你要嗤笑萬國。
PS|59|9|我 的力量啊，我要等候你， 因為上帝是我的庇護所。
PS|59|10|我的上帝要以慈愛 迎接我， 上帝要叫我看見我的仇敵遭報。
PS|59|11|主，我們的盾牌啊， 不要殺他們，免得我的子民遺忘； 求你用你的能力使他們四散， 使他們降為卑。
PS|59|12|願他們因口中的罪和嘴唇的言語， 被自己的驕傲抓住， 他們所說的盡是咒罵和謊話。
PS|59|13|求你發怒，使他們消滅， 求你使他們消滅，歸於無有， 使他們知道上帝在 雅各 中間掌權， 直到地極。（細拉）
PS|59|14|他們晚上轉回， 叫號如狗，圍城繞行。
PS|59|15|他們到處走動覓食， 若不飽足就咆哮不已。
PS|59|16|但我要歌頌你的能力， 早晨要高唱你的慈愛； 因為你是我的庇護所， 在急難的日子作過我的避難所。
PS|59|17|我的力量啊，我要歌頌你； 因為上帝是我的庇護所， 是賜恩給我的上帝。
PS|60|1|上帝啊，你丟棄了我們，破壞了我們； 你曾發怒，求你使我們復興！
PS|60|2|你使地震動，崩裂； 求你將裂口補好，因為地在搖動。
PS|60|3|你讓你的子民遇見艱難， 使我們喝那令人東倒西歪的酒。
PS|60|4|你把旌旗賜給敬畏你的人， 可以躲避弓箭 。（細拉）
PS|60|5|求你應允我們 ，用右手施行拯救， 好讓你所親愛的人得救。
PS|60|6|上帝在他的聖所 說： 「我要歡樂； 要劃分 示劍 ， 丈量 疏割谷 。
PS|60|7|基列 是我的， 瑪拿西 是我的。 以法蓮 是護衛我頭的， 猶大 是我的權杖。
PS|60|8|摩押 是我的沐浴盆， 我要向 以東 扔鞋。 非利士 啊，你還能因我歡呼嗎？」
PS|60|9|誰能領我進堅固城？ 誰能引我到 以東 地？
PS|60|10|上帝啊，你真的丟棄了我們嗎？ 上帝啊，你不和我們的軍隊同去嗎？
PS|60|11|求你幫助我們攻擊敵人， 因為人的幫助是枉然的。
PS|60|12|我們倚靠上帝才得施展大能， 因為踐踏我們敵人的就是他。
PS|61|1|上帝啊，求你聽我的呼求， 留心聽我的禱告！
PS|61|2|我心裏發昏的時候， 要從地極求告你。 求你領我到那比我更高的磐石，
PS|61|3|因為你是我的避難所， 是我的堅固臺，使我脫離仇敵。
PS|61|4|我要永遠住在你的帳幕裏！ 我要投靠在你翅膀下的隱密處！（細拉）
PS|61|5|上帝啊，你聽了我所許的願； 你將產業賜給敬畏你名的人。
PS|61|6|求你加添王的壽數， 使他的年歲存到世世代代。
PS|61|7|願他在上帝面前永遠坐在王位上， 求你預備慈愛和信實保佑他！
PS|61|8|這樣，我要歌頌你的名，直到永遠， 天天還我所許的願。
PS|62|1|我的心默默無聲，專等候上帝， 我的救恩從他而來。
PS|62|2|惟獨他是我的磐石，我的拯救； 他是我的庇護所，我必不大大動搖。
PS|62|3|你們大家攻擊一人，使他被殺， 如歪斜的牆、將倒的壁，要到幾時呢？
PS|62|4|他們彼此商議，要把他從高位上拉下來； 他們喜愛謊話，口雖祝福，心卻詛咒。（細拉）
PS|62|5|我的心哪，你當默默無聲，專等候上帝， 因為我的盼望是從他而來。
PS|62|6|惟獨他是我的磐石，我的拯救； 他是我的庇護所，我必不動搖。
PS|62|7|我的拯救、我的榮耀都在於上帝； 我力量的磐石、我的避難所都在於上帝。
PS|62|8|百姓啊，要時時倚靠他， 在他面前傾心吐意； 上帝是我們的避難所。（細拉）
PS|62|9|人真是虛空， 人真是虛假； 放在天平裏就必浮起， 他們一共比空氣還輕。
PS|62|10|不要仗勢欺人， 也不要因搶奪而驕傲； 若財寶加增，不要放在心上。
PS|62|11|上帝說了一次、兩次，我都聽見了， 就是能力屬乎上帝。
PS|62|12|主啊，慈愛也是屬乎你， 因為你照著各人所做的報應他。
PS|63|1|上帝啊，你是我的上帝， 我要切切尋求你； 在乾旱疲乏無水之地， 我的心靈渴想你，我的肉身切慕你。
PS|63|2|我在聖所中曾如此瞻仰你， 為要見你的能力和你的榮耀。
PS|63|3|因你的慈愛比生命更好， 我的嘴唇要頌讚你。
PS|63|4|我還活著的時候要這樣稱頌你， 我要奉你的名舉手。
PS|63|5|我在床上記念你， 在夜更的時候思念你； 我的心像吃飽了骨髓肥油， 我也要以歡樂的嘴唇讚美你。
PS|63|6|
PS|63|7|因為你曾幫助了我， 我要在你翅膀的蔭下歡呼。
PS|63|8|我的心緊緊跟隨你； 你的右手扶持了我。
PS|63|9|但那些尋索要滅我命的人 必往地底下去；
PS|63|10|他們必被刀劍所殺， 成為野狗的食物。
PS|63|11|但是王必因上帝歡喜， 凡指著他發誓的都要誇耀， 因為說謊之人的口必被塞住。
PS|64|1|上帝啊，我哀嘆的時候，求你聽我的聲音！ 求你保護我的性命，不受仇敵的驚嚇！
PS|64|2|求你把我隱藏， 使我脫離作惡之人的暗謀， 脫離作孽之人的擾亂。
PS|64|3|他們磨舌如刀， 發出苦毒的言語，好像瞄準了的箭，
PS|64|4|要在暗地裏射完全人； 他們忽然射他，並不懼怕。
PS|64|5|他們彼此勉勵，設下惡計； 他們商量，暗設圈套， 說：「誰能看見呢？」
PS|64|6|他們圖謀奸惡： 「我們完成了精密的策劃。」 各人的意念心思是深沉的。
PS|64|7|但上帝要用箭射他們， 他們忽然受了傷。
PS|64|8|他們必然絆跌，被自己的舌頭所害； 凡看見他們的都必搖頭。
PS|64|9|眾人都要害怕， 要傳揚上帝的工作， 並且明白他的作為。
PS|64|10|義人必因耶和華歡喜，並要投靠他； 凡心裏正直的人都必誇耀。
PS|65|1|上帝啊，在 錫安 ，人都等候讚美你， 也要向你還所許的願。
PS|65|2|聽禱告的主啊， 凡有血肉之軀的都要來就你。
PS|65|3|罪孽勝了我； 至於我們的過犯，你都要赦免。
PS|65|4|你所揀選、使他親近你、住在你院中的， 這人有福了！ 我們要因你居所、你聖殿的美福知足。
PS|65|5|拯救我們的上帝啊，你必以威嚴秉公義應允我們； 地極和海角遠方的人都倚靠你。
PS|65|6|你既以大能束腰， 就用力量安定諸山，
PS|65|7|使諸海的響聲和其中波浪的響聲， 並萬民的喧嘩，都平靜了。
PS|65|8|住在地極的人因你的神蹟懼怕， 你使日出日落之地都歡呼。
PS|65|9|你眷顧地， 降雨使地大大肥沃。 上帝的河滿了水； 你這樣澆灌了地， 好為人預備五穀。
PS|65|10|你澆透地的犁溝，潤澤犁脊， 降甘霖，使地鬆軟； 其中生長的，蒙你賜福。
PS|65|11|你以恩惠為年歲的冠冕， 你的路徑都滴下油脂，
PS|65|12|滴在曠野的草場上。 小山以歡樂束腰，
PS|65|13|草場以羊群為衣， 谷中也長滿了五穀； 這一切都歡呼歌唱。
PS|66|1|全地都當向上帝歡呼！
PS|66|2|當歌頌他名的榮耀， 使讚美他的話大有榮耀！
PS|66|3|當對上帝說：「你的作為何等可畏！ 因你的大能，仇敵要向你投降。
PS|66|4|全地要敬拜你，歌頌你， 要歌頌你的名。」（細拉）
PS|66|5|你們來看上帝所做的， 他向世人所做之事是可畏的。
PS|66|6|他將海變成乾地，使百姓步行過河； 我們在那裏要因他歡喜。
PS|66|7|他用權能治理，直到永遠。 他的眼睛鑒察萬民； 悖逆的人不可自高。（細拉）
PS|66|8|萬民哪，你們當稱頌我們的上帝， 使人得聽讚美他的聲音。
PS|66|9|他使我們的性命存活， 不叫我們的腳搖動。
PS|66|10|上帝啊，你曾考驗我們， 你熬煉我們，如煉銀子一樣。
PS|66|11|你使我們進入羅網， 把重擔放在我們身上。
PS|66|12|你使人坐車軋我們的頭； 我們經過水火， 你卻使我們到豐富之地。
PS|66|13|我要帶著燔祭進你的殿， 向你還我的願，
PS|66|14|就是在急難時我嘴唇所發的、 口中所許的。
PS|66|15|我要將肥牛的燔祭 和公羊的香祭獻給你， 又要把公牛和公山羊獻上。（細拉）
PS|66|16|敬畏上帝的人哪，你們都來聽！ 我要述說他為我所做的事。
PS|66|17|我曾用口求告他， 我的舌頭也稱他為高。
PS|66|18|我若心裏注重罪孽， 主必不聽。
PS|66|19|但上帝實在聽見了， 他留心聽了我禱告的聲音。
PS|66|20|上帝是應當稱頌的！ 他沒有推卻我的禱告， 也沒有使他的慈愛離開我。
PS|67|1|願上帝憐憫我們，賜福給我們， 使他的臉向我們發光，（細拉）
PS|67|2|好讓全地得知你的道路， 萬國得知你的救恩。
PS|67|3|上帝啊，願萬民稱謝你！ 願萬民都稱謝你！
PS|67|4|願萬族都快樂歡呼； 因為你必按公正審判萬民， 引導地上的萬族。（細拉）
PS|67|5|上帝啊，願萬民稱謝你！ 願萬民都稱謝你！
PS|67|6|地已經出了土產， 上帝，我們的上帝，要賜福給我們。
PS|67|7|上帝要賜福給我們， 地的四極都要敬畏他！
PS|68|1|願上帝興起，使他的仇敵四散， 使那恨他的人從他面前逃跑。
PS|68|2|你驅逐他們 ，如煙被吹散； 惡人見上帝的面就消滅，如蠟被火熔化。
PS|68|3|惟有義人必然歡喜， 在上帝面前快樂， 他們要在喜樂中歡欣。
PS|68|4|你們當向上帝唱詩，歌頌他的名； 為那駕車經過曠野的修平道路 。 他的名是耶和華， 你們要在他面前歡樂！
PS|68|5|上帝在他的聖所作孤兒的父， 作寡婦的伸冤者。
PS|68|6|上帝使孤獨的有家， 使被囚的出來享福； 惟有悖逆的要住在乾旱之地。
PS|68|7|上帝啊，當你走在百姓前頭， 在曠野行進，（細拉）
PS|68|8|地見上帝的面就震動，天也降雨； 西奈山 見 以色列 上帝的面也震動。
PS|68|9|上帝啊，你降下大雨； 你的產業 以色列 疲乏的時候，你使他堅固。
PS|68|10|你的會眾住在境內； 上帝啊，你在恩惠中為困苦人預備所需的。
PS|68|11|主發命令， 傳好信息的婦女成了大群：
PS|68|12|「統領大軍的君王逃跑了，逃跑了！」 在家等候的婦女也分得了掠物。
PS|68|13|你們躺臥在羊圈， 好像鴿子的翅膀鍍銀，翎毛鍍金一般。
PS|68|14|全能者在境內趕散列王的時候， 勢如飄雪在 撒們 。
PS|68|15|巴珊山 是極其宏偉 的山， 巴珊山 是多峰多嶺的山。
PS|68|16|你們多峰多嶺的山哪， 為何以妒忌的眼光看上帝所願居住的山？ 耶和華必住這山，直到永遠！
PS|68|17|上帝的車輦累萬盈千； 主在其中，好像在 西奈 聖山一樣。
PS|68|18|你已經升上高天，擄掠了俘虜； 你在人間，就是在悖逆的人中，受了供獻， 使耶和華上帝可以與他們同住。
PS|68|19|天天背負我們重擔的主， 就是拯救我們的上帝， 是應當稱頌的！（細拉）
PS|68|20|上帝是為我們施行拯救的上帝； 人能脫離死亡是在乎主─耶和華。
PS|68|21|但上帝要打破他仇敵的頭， 就是那常犯罪之人的頭顱。
PS|68|22|主說：「我要使百姓從 巴珊 歸來， 使他們從深海轉回，
PS|68|23|好叫你打碎仇敵，使你的腳踹在血中， 使你狗的舌頭也有份。」
PS|68|24|上帝啊，你是我的上帝，我的王； 人已經看見你行走，進入聖所。
PS|68|25|歌唱的行在前，作樂的隨在後， 都在擊鼓的童女中間：
PS|68|26|「從 以色列 源頭而來的啊， 你們當在各會中稱頌上帝─耶和華！」
PS|68|27|在那裏，有統管他們的小 便雅憫 ， 有 猶大 的領袖和他們的一群人， 有 西布倫 的領袖， 有 拿弗他利 的領袖。
PS|68|28|你的上帝已賜給你力量 ； 上帝啊，求你堅固你為我們所成全的事！
PS|68|29|因你 耶路撒冷 的殿， 列王必帶貢物獻給你。
PS|68|30|求你斥責蘆葦中的野獸和公牛群， 並萬民中的牛犢。 直到他們帶著銀塊來朝貢 ； 上帝已經趕散好戰的萬民 。
PS|68|31|埃及 的使臣要出來， 古實 人要急忙向上帝伸出手來。
PS|68|32|地上的國度啊， 你們要向上帝歌唱， 要歌頌主，（細拉）
PS|68|33|就是那駕行在亙古的諸天之上的主！ 聽啊，他發出聲音，是極大的聲音。
PS|68|34|你們要將能力歸給上帝； 他的威榮在 以色列 之上， 他的能力顯在天上。
PS|68|35|上帝啊，你從聖所顯為可畏， 以色列 的上帝是那將力量權能賜給他百姓的。 上帝是應當稱頌的！
PS|69|1|上帝啊，求你救我！ 因為眾水就要淹沒我。
PS|69|2|我深陷在淤泥中，沒有立腳之地； 我到了深水之中，波濤漫過我身。
PS|69|3|我因呼求困乏，喉嚨發乾； 我因等候上帝，眼睛失明。
PS|69|4|無故恨我的，比我的頭髮還多； 無理與我為仇、要把我剪除的，甚為強盛。 我沒有搶奪，他們竟然要我償還！
PS|69|5|上帝啊，我的愚昧，你原知道， 我的罪愆不能向你隱瞞。
PS|69|6|萬軍之主耶和華啊， 求你不要讓那等候你的因我蒙羞！ 以色列 的上帝啊， 求你不要讓那尋求你的因我受辱！
PS|69|7|因我為你的緣故受了辱罵， 滿面羞愧。
PS|69|8|我的兄弟把我當陌生人， 我母親的兒子把我當外邦人。
PS|69|9|因我為你的殿心裏焦急，如同火燒， 並且辱罵你的人的辱罵都落在我身上。
PS|69|10|我哭泣，以禁食刻苦我心； 這倒成了我的羞辱。
PS|69|11|我拿麻布當衣裳， 卻成了他們的笑柄。
PS|69|12|坐在城門口的談論我， 酒徒也以我為歌曲。
PS|69|13|至於我，耶和華啊，在悅納的時候我向你祈禱。 上帝啊，求你按你豐盛的慈愛， 憑你拯救的信實應允我！
PS|69|14|求你搭救我脫離淤泥， 不叫我陷在其中； 求你使我脫離那些恨我的人， 使我脫離深水。
PS|69|15|求你不容波濤漫過我， 不容深淵吞滅我， 不容深坑在我以上合口。
PS|69|16|耶和華啊，求你應允我！ 因為你的慈愛本為美好； 求你按你豐盛的憐憫轉回眷顧我！
PS|69|17|不要轉臉不顧你的僕人； 我在急難之中，求你速速應允我！
PS|69|18|求你親近我，救贖我！ 求你因我仇敵的緣故將我贖回！
PS|69|19|你知道我所受的辱罵、欺凌、羞辱； 我的敵人都在你面前。
PS|69|20|辱罵刺傷我的心， 使我憂愁。 我指望有人體恤，卻沒有一個； 指望有人安慰，卻找不著一個。
PS|69|21|他們拿苦膽給我當食物； 我渴了，他們拿醋給我喝。
PS|69|22|願他們的筵席在他們面前變為羅網， 在他們平安的時候 變為圈套。
PS|69|23|願他們的眼睛昏花，看不見； 求你使他們的腰常常戰抖。
PS|69|24|求你將你的惱恨倒在他們身上， 使你的烈怒追上他們。
PS|69|25|願他們的住處變為廢墟， 他們的帳棚無人居住。
PS|69|26|因為你所擊打的，他們就迫害； 你所擊傷的，他們述說 他的愁苦。
PS|69|27|求你使他們罪上加罪， 不容他們在你面前稱義。
PS|69|28|願他們從生命冊上被塗去， 不得名列在義人之中。
PS|69|29|但我困苦憂傷； 上帝啊，願你的救恩將我安置在高處。
PS|69|30|我要以詩歌讚美上帝的名， 以感謝尊他為大！
PS|69|31|這就讓耶和華喜悅，勝似獻牛， 獻有角有蹄的公牛。
PS|69|32|謙卑的人看見了就喜樂； 尋求上帝的人，願你們的心甦醒。
PS|69|33|因為耶和華聽了窮乏的人， 不藐視被囚的人。
PS|69|34|願天和地、 海洋和其中一切的動物都讚美他！
PS|69|35|因為上帝要拯救 錫安 ，建造 猶大 的城鎮； 他的子民要在那裏居住，得地為業。
PS|69|36|他僕人的後裔要承受這地， 愛他名的人要住在其中。
PS|70|1|上帝啊，求你快快搭救我！ 耶和華啊，求你速速幫助我！
PS|70|2|願那些尋索我命的，抱愧蒙羞； 願那些喜悅我遭害的，退後受辱。
PS|70|3|願那些對我說「啊哈、啊哈」的， 因羞愧退後。
PS|70|4|願所有尋求你的，因你歡喜快樂； 願那些喜愛你救恩的，常說：「當尊上帝為大！」
PS|70|5|但我是困苦貧窮的； 上帝啊，求你速速到我這裏來！ 你是幫助我的，搭救我的； 耶和華啊，求你不要耽延！
PS|71|1|耶和華啊，我投靠你， 求你叫我永不羞愧！
PS|71|2|求你憑你的公義搭救我，救拔我； 側耳聽我，拯救我！
PS|71|3|求你作我常來棲身 的磐石， 你已經吩咐要救我， 因為你是我的巖石、我的山寨。
PS|71|4|我的上帝啊，求你救我脫離惡人的手， 脫離不義和殘暴之人的手。
PS|71|5|主耶和華啊，你是我所盼望的； 自我年幼，你是我所倚靠的。
PS|71|6|我自出母胎被你扶持， 使我出母腹的是你。 我要常常讚美你！
PS|71|7|許多人看我為異類， 但你是我堅固的避難所。
PS|71|8|我要滿口述說讚美你的話 終日榮耀你。
PS|71|9|我年老的時候，求你不要丟棄我！ 我體力衰弱時，求你不要離棄我！
PS|71|10|我的仇敵議論我， 那些窺探要害我命的一同商議，
PS|71|11|說：「上帝已經離棄他； 你們去追趕他，捉拿他吧！ 因為沒有人搭救。」
PS|71|12|上帝啊，求你不要遠離我！ 我的上帝啊，求你速速幫助我！
PS|71|13|願那與我為敵的，羞愧滅亡； 願那謀害我的，受辱蒙羞。
PS|71|14|我卻要常常仰望， 並要越發讚美你。
PS|71|15|我的口要終日述說你的公義和你的救恩， 因我無從計算其數。
PS|71|16|我要述說主耶和華的大能， 我單要提說你的公義。
PS|71|17|上帝啊，自我年幼，你就教導我； 直到如今，我傳揚你奇妙的作為。
PS|71|18|上帝啊，我年老髮白的時候， 求你不要離棄我！ 等我宣揚你的能力給下一代， 宣揚你的大能給後世的人。
PS|71|19|上帝啊，你的公義極高； 行過大事的上帝啊，誰能像你？
PS|71|20|你是叫我多經歷重大急難的， 必使我再活過來， 從地的深處救我上來。
PS|71|21|你必使我越發昌大， 又轉來安慰我。
PS|71|22|我的上帝啊，我要鼓瑟稱謝你， 稱謝你的信實！ 以色列 的聖者啊，我要彈琴歌頌你！
PS|71|23|我歌頌你的時候，我的嘴唇要歡呼； 我的性命，就是你所救贖的，也要歡呼。
PS|71|24|我的舌頭也必終日講論你的公義， 因為那些謀害我的人已經蒙羞受辱了。
PS|72|1|上帝啊，求你將你的公平賜給王， 將你的公義賜給王的兒子。
PS|72|2|使他按公義審判你的子民， 按公平審判你的困苦人。
PS|72|3|大山小山都要因公義 使百姓得享平安。
PS|72|4|他必為百姓中困苦的人伸冤， 拯救貧窮之輩， 壓碎那欺壓人的人。
PS|72|5|太陽還存，月亮猶在， 人要敬畏你 ，直到萬代！
PS|72|6|他必降臨，像雨降在已割的草地上， 如甘霖滋潤田地。
PS|72|7|在他的日子，公義 要興旺， 大有平安，除非月亮不在。
PS|72|8|他要執掌權柄，從這海直到那海， 從 大河 直到地極。
PS|72|9|住在曠野的必在他面前下拜， 他的仇敵必要舔土。
PS|72|10|他施 和海島的王要進貢， 示巴 和 西巴 的王要獻禮物。
PS|72|11|眾王都要叩拜他， 萬國都要事奉他。
PS|72|12|貧窮人呼求，他要搭救， 無人幫助的困苦人，他也搭救。
PS|72|13|他要憐憫貧寒和貧窮的人， 拯救貧窮人的性命。
PS|72|14|他要救贖他們脫離欺壓和殘暴， 他們的血在他眼中看為寶貴。
PS|72|15|願他永遠活著， 示巴 的金子要獻給他； 願人常常為他禱告，終日祝福他。
PS|72|16|在地的山頂上，願五穀茂盛， 所結的穀實響動，如 黎巴嫩 的樹林； 願城裏的人興旺，如地上的草。
PS|72|17|願他的名存到永遠， 他的名如太陽之長久 ； 願人因他蒙福， 萬國稱他為有福。
PS|72|18|惟獨耶和華－ 以色列 的上帝能行奇事， 他是應當稱頌的！
PS|72|19|他榮耀的名也當稱頌，直到永遠。 願他的榮耀充滿全地！ 阿們！阿們！
PS|72|20|耶西 的兒子－ 大衛 的祈禱完畢。 亞薩的詩。
PS|73|1|上帝實在恩待 以色列 那些清心的人！
PS|73|2|至於我，我的腳幾乎失閃， 我的步伐險些走偏；
PS|73|3|因為我嫉妒狂傲的人， 我看見惡人享平安。
PS|73|4|他們的力氣強壯， 他們死的時候也沒有疼痛。
PS|73|5|他們不像別人受苦， 也不像別人遭災。
PS|73|6|所以，驕傲如鏈子戴在他們項上， 殘暴像衣裳覆蓋在他們身上。
PS|73|7|他們的眼睛 因體胖而凸出， 他們的內心放任不羈 。
PS|73|8|他們譏笑人，憑惡意說欺壓人的話。 他們說話自高；
PS|73|9|他們的口褻瀆上天， 他們的舌毀謗全地。
PS|73|10|所以他的百姓歸到這裏， 享受滿杯的水 。
PS|73|11|他們說：「上帝怎能曉得？ 至高者哪會知道呢？」
PS|73|12|看哪，這就是惡人， 他們常享安逸，財寶增多。
PS|73|13|我實在徒然潔淨了我的心， 徒然洗手表明我的無辜，
PS|73|14|因為我終日遭災難， 每日早晨受懲治。
PS|73|15|我若說「我要這樣講」， 就是愧對這世代的眾兒女了。
PS|73|16|我思索要明白這事， 眼看實係為難，
PS|73|17|直到我進了上帝的聖所， 思想他們的結局。
PS|73|18|你實在把他們安放在滑地， 使他們跌倒滅亡；
PS|73|19|他們轉眼之間成了何等荒涼！ 他們被驚恐滅盡了。
PS|73|20|人睡醒了，怎樣看夢， 主啊，你醒了也必照樣輕看他們的影像。
PS|73|21|因此，我心裏苦惱， 肺腑被刺。
PS|73|22|我這樣愚昧無知， 在你面前如同畜牲。
PS|73|23|然而，我常與你同在； 你攙扶我的右手。
PS|73|24|你要以你的訓言引導我， 以後你必接我到榮耀裏。
PS|73|25|除你以外，在天上我有誰呢？ 除你以外，在地上我也沒有所愛慕的。
PS|73|26|我的肉體和我的心腸衰殘； 但上帝是我心裏的力量， 又是我的福分，直到永遠。
PS|73|27|看哪，遠離你的，必要死亡； 凡離棄你行淫的，你都滅絕了。
PS|73|28|但我親近上帝是於我有益； 我以主耶和華為我的避難所， 好叫我述說你一切的作為。
PS|74|1|上帝啊，你為何永遠丟棄我們呢？ 為何向你草場的羊發怒，如煙冒出呢？
PS|74|2|求你記念你古時得來的會眾， 就是你所贖、作你產業支派的， 並記念你向來居住的 錫安山 。
PS|74|3|求你舉步去看那日久荒涼之地， 看仇敵在聖所中所做的一切惡事。
PS|74|4|你的敵人在你會中吼叫， 他們豎起自己的標幟為記號，
PS|74|5|好像人揚起斧子 對著林中的樹，
PS|74|6|現在將聖所中的雕刻 ， 全都用斧子錘子打壞。
PS|74|7|他們用火焚燒你的聖所， 褻瀆你名的居所於地。
PS|74|8|他們心裏說「我們要盡行毀滅」； 就在遍地燒燬敬拜上帝聚會的所在。
PS|74|9|我們看不見自己的標幟，不再有先知， 我們當中也無人知道這災禍要到幾時。
PS|74|10|上帝啊，敵人辱罵要到幾時呢？ 仇敵藐視你的名要到永遠嗎？
PS|74|11|你為甚麼縮回你的右手？ 求你從懷中伸出手來，毀滅他們。
PS|74|12|上帝自古以來是我的王， 在這地上施行拯救。
PS|74|13|你曾用能力將海分開， 你打破水裏大魚的頭。
PS|74|14|你曾壓碎 力威亞探 的頭， 把牠給曠野的禽獸作食物。
PS|74|15|你曾分裂泉源和溪流； 使長流的江河枯乾。
PS|74|16|白晝屬你，黑夜也屬你； 亮光和太陽是你預備的。
PS|74|17|地的一切疆界是你立的， 夏天和冬天是你定的。
PS|74|18|耶和華啊，仇敵辱罵，愚頑之輩藐視你的名； 求你記念這事。
PS|74|19|不要將屬你的斑鳩 交給野獸， 不要永遠忘記你困苦人的性命。
PS|74|20|求你顧念所立的約， 因為地上黑暗之處遍滿了兇暴。
PS|74|21|不要讓受欺壓的人蒙羞回去； 要使困苦貧窮的人讚美你的名。
PS|74|22|上帝啊，求你起來為自己辯護！ 求你記念愚頑人怎樣終日辱罵你。
PS|74|23|不要忘記你敵人的喧鬧， 就是那時常上升、起來對抗你之人的喧嘩。
PS|75|1|上帝啊，我們稱謝你，我們稱謝你！ 你的名臨近，人 都述說你奇妙的作為。
PS|75|2|我選定了日期， 必按正直施行審判。
PS|75|3|地和其上的居民都熔化了； 我親自堅立地的柱子。（細拉）
PS|75|4|我對狂傲的人說：「不要狂傲！」 對兇惡的人說：「不要舉角！」
PS|75|5|不要把你們的角高舉， 不要挺著頸項 說話。
PS|75|6|因為高舉非從東，非從西， 也非從南而來。
PS|75|7|惟有上帝斷定， 他使這人降卑，使那人升高。
PS|75|8|耶和華的手裏有杯， 杯內滿了調和起沫的酒； 他倒出來， 地上的惡人都必喝，直到喝盡它的渣滓。
PS|75|9|但我要宣揚，直到永遠！ 我要歌頌 雅各 的上帝！
PS|75|10|惡人一切的角，我要砍斷； 惟有義人的角必被高舉。
PS|76|1|在 猶大 ，上帝為人所認識； 在 以色列 ，他的名為大。
PS|76|2|在 撒冷 有他的住處， 在 錫安 有他的居所。
PS|76|3|他在那裏折斷弓上的火箭、 盾牌、刀劍和戰爭的兵器。（細拉）
PS|76|4|你是光榮的， 比獵物 之山更威嚴。
PS|76|5|心中勇敢的人都被掠奪； 他們睡了長覺，沒有一個英雄能措手。
PS|76|6|雅各 的上帝啊，你的斥責一發， 戰車和戰馬都沉睡了。
PS|76|7|你，惟獨你是可畏的！ 你的怒氣一發，誰能在你面前站得住呢？
PS|76|8|你從天上使人聽判斷。 上帝起來施行審判， 要救地上所有困苦的人； 那時地就懼怕而靜默。（細拉）
PS|76|9|
PS|76|10|人的憤怒終必稱謝你， 你要以人的餘怒束腰。
PS|76|11|你們當向耶和華－你們的上帝許願，還願； 在他四圍的人都當拿貢物獻給那可畏的主。
PS|76|12|他要挫折王子的驕氣， 向地上的君王顯為可畏。
PS|77|1|我要向上帝發聲呼求； 我向上帝發聲，他必側耳聽我。
PS|77|2|我在患難之日尋求主， 在夜間不住地舉手禱告 ， 我的心不肯受安慰。
PS|77|3|我想念上帝，就煩躁不安； 我沉思默想，心靈發昏。（細拉）
PS|77|4|你使我不能閉眼； 我心煩亂，甚至不能說話。
PS|77|5|我追想古時之日， 上古之年。
PS|77|6|夜間我想起我的歌曲 ， 我的心默想，我的靈仔細省察：
PS|77|7|「難道主要永遠丟棄我， 不再施恩嗎？
PS|77|8|難道他的慈愛永遠窮盡， 他的應許世世廢棄嗎？
PS|77|9|難道上帝忘記施恩， 因發怒就止住他的憐憫嗎？」（細拉）
PS|77|10|我說，至高者右手的能力已改變， 這是我的悲哀。
PS|77|11|我要記念耶和華所做的， 要記念你古時的奇事；
PS|77|12|我要思想你所做的， 默念你的作為。
PS|77|13|上帝啊，你的道是神聖的； 有何神明大如上帝呢？
PS|77|14|你是行奇事的上帝， 你曾在萬民中彰顯能力。
PS|77|15|你曾用膀臂贖了你的子民， 就是 雅各 和 約瑟 的子孫。（細拉）
PS|77|16|上帝啊，眾水見你， 眾水一見你就都驚惶， 深淵也都戰抖。
PS|77|17|密雲倒出水來， 天空發出響聲， 你的箭也飛行四方。
PS|77|18|你的雷聲在旋風之中， 閃電照亮世界， 大地戰抖震動。
PS|77|19|你的道在海中， 你的路在大水之中， 你的腳蹤無人知道。
PS|77|20|你曾藉 摩西 和 亞倫 的手引導你的百姓， 好像領羊群一般。
PS|78|1|我的子民哪，要側耳聽我的訓誨， 豎起耳朵聽我口中的言語。
PS|78|2|我要開口說比喻， 我要解開古時的謎語，
PS|78|3|是我們所聽見、所知道， 我們的祖宗告訴我們的。
PS|78|4|我們不要向子孫隱瞞這些事， 而要將耶和華的美德和他的能力， 並他所行的奇事，述說給後代聽。
PS|78|5|他在 雅各 中立法度， 在 以色列 中設律法； 他吩咐我們的祖宗要傳給子孫，
PS|78|6|使將要生的後代子孫可以曉得。 他們也要起來告訴他們的子孫，
PS|78|7|好讓他們仰望上帝， 不忘記上帝的作為， 惟遵守他的命令；
PS|78|8|不要像他們的祖宗， 是頑梗悖逆、心不堅定， 向上帝心不忠實之輩。
PS|78|9|以法蓮 人帶著兵器，拿著弓， 臨陣之日轉身退後。
PS|78|10|他們不遵守上帝的約， 不肯照他的律法行；
PS|78|11|又忘記他的作為 和他所彰顯的奇事。
PS|78|12|他在 埃及 地，在 瑣安 田， 在他們祖宗眼前施行奇事。
PS|78|13|他把海分開，使他們過去， 又叫水立起如壘。
PS|78|14|他白日用雲彩， 終夜用火光引導他們。
PS|78|15|他在曠野使磐石裂開， 多多地給他們水喝，如從深淵而出。
PS|78|16|他使水從磐石湧出， 叫水如江河下流。
PS|78|17|他們卻仍舊得罪他， 在乾旱之地悖逆至高者。
PS|78|18|他們心中試探上帝， 隨自己所欲的求食物，
PS|78|19|並且妄論上帝說： 「上帝豈能在曠野擺設筵席嗎？
PS|78|20|他雖曾擊打磐石，使水湧出，如江河氾濫； 他還能賜糧食嗎？ 還能為他的百姓預備吃的肉嗎？」
PS|78|21|所以，耶和華聽見就發怒， 有烈火向 雅各 點燃， 有怒氣向 以色列 上騰；
PS|78|22|因為他們不信服上帝， 不倚賴他的拯救。
PS|78|23|然而他卻吩咐天空， 又敞開天上的門，
PS|78|24|降嗎哪像雨，給他們吃， 將天上的糧食賜給他們。
PS|78|25|各人就吃大能者的食物； 他賜下糧食，使他們飽足。
PS|78|26|他令東風吹在天空， 用能力引來南風。
PS|78|27|他降肉像雨，多如塵土， 降飛鳥，多如海沙，
PS|78|28|落在他自己的營中， 在他帳幕的四周圍。
PS|78|29|他們吃了，而且飽足； 這樣就隨了他們所欲的。
PS|78|30|但在他們滿足食慾以前， 食物還在他們口中的時候，
PS|78|31|上帝的怒氣就向他們上騰， 殺了他們當中肥壯的人， 打倒 以色列 的青年。
PS|78|32|雖是這樣，他們仍舊犯罪， 不信他奇妙的作為。
PS|78|33|因此，他使他們的日子全歸虛空， 叫他們的年歲盡屬驚恐。
PS|78|34|他殺他們的時候，他們才求問他， 回心轉意，切切尋求上帝。
PS|78|35|他們追念上帝是他們的磐石， 至高的上帝是他們的救贖主。
PS|78|36|他們卻用口諂媚他， 用舌向他說謊。
PS|78|37|他們的心向他不堅定， 不忠於他的約。
PS|78|38|但他有憐憫， 赦免他們的罪孽， 沒有滅絕他們， 而且屢次撤銷他的怒氣， 不發盡他的憤怒。
PS|78|39|他想念他們不過是血肉之軀， 是一陣去而不返的風。
PS|78|40|他們在曠野悖逆他， 在荒地令他擔憂，何其多呢！
PS|78|41|他們再三試探上帝， 惹動 以色列 的聖者。
PS|78|42|他們不追念他手的能力， 和他救贖他們脫離敵人的日子；
PS|78|43|他怎樣在 埃及 顯神蹟， 在 瑣安 田顯奇事，
PS|78|44|把江河並河汊的水都變為血， 使他們不能喝。
PS|78|45|他使蒼蠅成群落在他們當中，吃盡他們， 又叫青蛙滅了他們，
PS|78|46|將他們的果實交給螞蚱， 把他們勞碌得來的交給蝗蟲。
PS|78|47|他降冰雹打壞他們的葡萄樹， 下寒霜打壞他們的桑樹，
PS|78|48|將他們的牲畜交給冰雹， 把他們的群畜交給閃電。
PS|78|49|他使猛烈的怒氣和憤怒、惱恨、苦難， 成了一群降災的使者，臨到他們。
PS|78|50|他為自己的怒氣修平了路， 將他們的性命交給瘟疫， 使他們死亡，
PS|78|51|在 埃及 擊殺所有的長子， 在 含 的帳棚中擊殺他們壯年時頭生的。
PS|78|52|他卻領出自己的子民如羊， 在曠野引導他們如羊群。
PS|78|53|他領他們穩穩妥妥地，使他們不致害怕； 海卻淹沒他們的仇敵。
PS|78|54|他帶他們到自己聖地的邊界， 到他右手所得的這山地。
PS|78|55|他在他們面前趕出外邦人， 用繩子抽籤量地給他們為業， 讓 以色列 支派的人住在自己的帳棚裏。
PS|78|56|他們仍舊試探，悖逆至高的上帝， 不遵守他的法度，
PS|78|57|反倒退後，行詭詐，像他們的祖宗一樣， 他們翻轉，如同鬆弛的弓，
PS|78|58|以丘壇惹他發怒， 以雕刻的偶像使他忌恨。
PS|78|59|上帝聽見就發怒， 全然棄絕了 以色列 ，
PS|78|60|甚至離棄 示羅 的帳幕， 就是他在人間所搭的帳棚；
PS|78|61|又將他有能力的約櫃 交給人擄去， 將他的榮耀交在敵人手中；
PS|78|62|並將他的百姓交給刀劍， 向他的產業發怒。
PS|78|63|壯丁被火燒滅， 童女也無婚禮頌歌。
PS|78|64|祭司倒在刀下， 寡婦卻不哀哭。
PS|78|65|那時，主像睡覺的人醒來， 如勇士飲酒呼喊。
PS|78|66|他擊退敵人， 叫他們永蒙羞辱。
PS|78|67|他撇棄 約瑟 的帳棚， 不揀選 以法蓮 支派，
PS|78|68|卻揀選 猶大 支派， 揀選他所喜愛的 錫安山 ；
PS|78|69|建造他的聖所如同高峰， 又像他所建立的永存之地。
PS|78|70|他揀選他的僕人 大衛 ， 從羊圈中將他召來，
PS|78|71|叫他不再牧放那些母羊， 為要牧養自己的百姓 雅各 和自己的產業 以色列 。
PS|78|72|於是，他以純正的心牧養他們， 用巧妙的手引導他們。
PS|79|1|上帝啊，外邦人侵犯你的產業， 玷污你的聖殿，使 耶路撒冷 變成廢墟，
PS|79|2|將你僕人的屍首交給天空的飛鳥為食， 把你聖民的肉交給地上的走獸，
PS|79|3|耶路撒冷 的周圍流出他們的血如水， 無人埋葬。
PS|79|4|我們成為鄰國羞辱的對象， 被四圍的人嗤笑譏刺。
PS|79|5|耶和華啊，你發怒要到幾時呢？ 要到永遠嗎？ 你的忌恨要如火焚燒嗎？
PS|79|6|求你將你的憤怒傾倒在那不認識你的萬邦 和那不求告你名的國度。
PS|79|7|因為他們吞了 雅各 ， 將他的住處變為廢墟。
PS|79|8|求你不要記得我們先前世代的罪孽； 願你的憐憫速速臨到我們， 因為我們落到極卑微的地步。
PS|79|9|拯救我們的上帝啊，求你因你名的榮耀幫助我們！ 為你名的緣故搭救我們，赦免我們的罪。
PS|79|10|為何讓列國說「他們的上帝在哪裏」呢？ 求你讓列國知道， 你在我們眼前伸你僕人流血的冤。
PS|79|11|願被囚之人的嘆息達到你面前， 求你以強大的膀臂存留那些將死的人。
PS|79|12|主啊，求你將我們鄰邦所加給你的羞辱 七倍歸到他們身上。
PS|79|13|這樣，你的子民，你草場的羊， 要稱謝你，直到永遠； 要述說讚美你的話，直到萬代。
PS|80|1|領 約瑟 如領羊群的 以色列 牧者啊，求你側耳而聽！ 在基路伯之上坐寶座的啊，求你發出光來！
PS|80|2|在 以法蓮 、 便雅憫 、 瑪拿西 面前 求你施展你的大能，拯救我們。
PS|80|3|上帝啊，求你使我們回轉 ， 使你的臉發光，我們就會得救！
PS|80|4|耶和華─萬軍之上帝啊， 你因你百姓的禱告發怒，要到幾時呢？
PS|80|5|你以眼淚當食物給他們吃， 量出滿碗的眼淚給他們喝。
PS|80|6|你使鄰邦因我們紛爭， 我們的仇敵彼此戲笑。
PS|80|7|萬軍之上帝啊，求你使我們回轉， 使你的臉發光，我們就會得救！
PS|80|8|你從 埃及 拔出一棵葡萄樹， 趕出外邦人，把這樹栽上。
PS|80|9|你在它面前清除雜物， 它就深深扎根，蔓延滿地。
PS|80|10|它的影子遮蔽群山， 枝子好像高大的香柏樹。
PS|80|11|它長出枝子，直到大海， 伸展嫩枝，延到 大河 。
PS|80|12|你為何拆毀這樹的籬笆， 任憑路人摘取？
PS|80|13|林中的野豬踐踏它， 田裏的走獸吞吃它。
PS|80|14|萬軍之上帝啊，求你轉回， 從天上垂看觀察，眷顧這葡萄樹；
PS|80|15|保護你右手所栽的根， 你為自己所堅固的幼苗。
PS|80|16|這樹已經被火焚燒，被刀砍伐， 因你臉上的怒容就滅亡了。
PS|80|17|願你的手扶持你右邊的人， 你為自己所堅固的人子。
PS|80|18|這樣，我們就不背離你； 求你救活我們，讓我們得以求告你的名。
PS|80|19|耶和華─萬軍之上帝啊，求你使我們回轉， 使你的臉發光，我們就會得救！
PS|81|1|你們當向上帝－我們的力量大聲歌唱， 向 雅各 的上帝歡呼！
PS|81|2|高唱詩歌，擊打手鼓， 彈奏悅耳的琴瑟。
PS|81|3|當在新月和滿月－ 我們過節的日期吹角，
PS|81|4|因這是為 以色列 所定的律例， 是 雅各 上帝的典章。
PS|81|5|他攻擊 埃及 地的時候， 曾立此為 約瑟 的法度。 我聽見我所不明白的語言：
PS|81|6|「我使你 的肩頭得脫重擔， 使你的手放下筐子。
PS|81|7|你在急難中呼求，我就搭救你， 在雷的隱密處應允你， 在 米利巴 水那裏考驗你。（細拉）
PS|81|8|聽啊，我的子民，我要勸戒你； 以色列 啊，我真願你肯聽從我。
PS|81|9|在你當中，不可有外族的神明； 外邦的神明，你也不可下拜。
PS|81|10|我是耶和華－你的上帝， 曾將你從 埃及 地領上來； 你要大大張口，我就使你滿足。
PS|81|11|「無奈，我的子民不聽我的聲音， 以色列 不肯聽從我。
PS|81|12|我就任憑他們心裏頑梗， 隨自己的計謀而行。
PS|81|13|我的子民若肯聽從我， 以色列 肯行我的道，
PS|81|14|我就速速制伏他們的仇敵， 反手攻擊他們的敵人。
PS|81|15|恨耶和華的人必來投降， 願他們的厄運直到永遠。
PS|81|16|他必拿上好的麥子給 以色列 吃， 又拿磐石出的蜂蜜使你飽足。 」
PS|82|1|上帝站立在神聖的會中， 在諸神中施行審判。
PS|82|2|你們審判不秉公義， 抬舉惡人的臉面，要到幾時呢？（細拉）
PS|82|3|當為貧寒的人和孤兒伸冤， 為困苦和窮乏的人施行公義。
PS|82|4|當保護貧寒和貧窮的人， 救他們脫離惡人的手。
PS|82|5|他們愚昧，他們無知， 在黑暗中走來走去； 地的根基都搖動了。
PS|82|6|我曾說：「你們是諸神， 都是至高者的兒子。
PS|82|7|然而，你們要死去，與世人一樣， 要仆倒，像任何一位王子一般。」
PS|82|8|上帝啊，求你起來審判全地， 因為你必得萬國為業。
PS|83|1|上帝啊，求你不要靜默！ 上帝啊，求你不要閉口，不要不作聲！
PS|83|2|因為你的仇敵喧嚷， 恨你的抬起頭來。
PS|83|3|他們同謀奸詐要害你的百姓， 彼此商議要害你所保護的人。
PS|83|4|他們說：「來吧，我們將他們除滅， 使他們不再成國！ 使 以色列 的名不再被人記念！」
PS|83|5|他們同心商議， 彼此結盟，要抵擋你；
PS|83|6|他們就是住帳棚的 以東 和 以實瑪利 人， 摩押 和 夏甲 人，
PS|83|7|迦巴勒 、 亞捫 、 亞瑪力 、 非利士 和 推羅 的居民。
PS|83|8|亞述 也與他們聯合， 作 羅得 子孫的幫手。（細拉）
PS|83|9|求你待他們，如待 米甸 ， 如在 基順河 待 西西拉 和 耶賓 一樣。
PS|83|10|他們在 隱‧多珥 滅亡， 成了地上的糞土。
PS|83|11|求你使他們的貴族像 俄立 和 西伊伯 ， 使他們的王子都像 西巴 和 撒慕拿 。
PS|83|12|因為他們說：「我們要得上帝的住處， 作自己的產業。」
PS|83|13|我的上帝啊，求你使他們像旋風中的塵土， 如風前的碎秸。
PS|83|14|火怎樣焚燒樹林， 火焰怎樣燒著山嶺，
PS|83|15|求你也照樣用狂風追趕他們， 用暴雨恐嚇他們。
PS|83|16|耶和華啊，求你使他們滿面羞恥， 好叫他們尋求你的名！
PS|83|17|願他們永遠羞愧驚惶！ 願他們慚愧滅亡！
PS|83|18|願他們認識你的名是耶和華， 惟獨你是掌管全地的至高者！
PS|84|1|萬軍之耶和華啊， 你的居所何等可愛！
PS|84|2|我羨慕渴想耶和華的院宇， 我的內心，我的肉體向永生上帝歡呼。
PS|84|3|萬軍之耶和華－我的王，我的上帝啊， 在你祭壇那裏，麻雀為自己找到了家， 燕子為自己找著菢雛之窩。
PS|84|4|如此住在你殿中的有福了！ 他們不斷地讚美你。（細拉）
PS|84|5|靠你有力量、心中嚮往 錫安 大道的， 這人有福了！
PS|84|6|他們經過「流淚谷」 ，叫這谷變為泉源之地； 且有秋雨之福蓋滿了全谷。
PS|84|7|他們行走，力上加力， 各人到 錫安 朝見上帝。
PS|84|8|萬軍之耶和華上帝啊，求你聽我的禱告！ 雅各 的上帝啊，求你側耳而聽！（細拉）
PS|84|9|上帝啊，我們的盾牌，求你觀看， 求你垂顧你受膏者的面！
PS|84|10|在你的院宇一日， 勝似千日； 寧可在我上帝的殿中看門， 不願住在惡人的帳棚裏。
PS|84|11|因為耶和華上帝是太陽，是盾牌， 耶和華要賜下恩惠和榮耀。 他未嘗留下福氣不給那些行動正直的人。
PS|84|12|萬軍之耶和華啊， 倚靠你的人有福了！
PS|85|1|耶和華啊，你已經向你的地施恩， 救回被擄的 雅各 。
PS|85|2|你赦免了你百姓的罪孽， 遮蓋了他們一切的過犯。（細拉）
PS|85|3|你收回所發的憤怒， 撤銷你猛烈的怒氣。
PS|85|4|拯救我們的上帝啊，求你使我們回轉， 使你向我們所發的憤怒止息。
PS|85|5|你要向我們發怒到永遠嗎？ 要將你的怒氣延留到萬代嗎？
PS|85|6|你不再將我們救活， 使你的百姓因你歡喜嗎？
PS|85|7|耶和華啊，求你使我們得見你的慈愛， 又將你的救恩賜給我們。
PS|85|8|我要聽上帝－耶和華所說的話， 因為他必應許賜平安給他的百姓，就是他的聖民； 他們卻不可再轉向愚昧 。
PS|85|9|他的救恩誠然與敬畏他的人相近， 使榮耀住在我們的地上。
PS|85|10|慈愛和誠實彼此相遇， 公義與和平彼此相親。
PS|85|11|誠實從地而生， 公義從天而現。
PS|85|12|耶和華必賜福氣給我們； 我們的地也要出土產。
PS|85|13|公義要行在他面前， 使他的腳蹤有可走之路。
PS|86|1|耶和華啊，求你側耳應允我， 因我是困苦貧窮的。
PS|86|2|求你保住我的性命，因我是虔誠的人。 我的上帝啊，求你拯救我這倚靠你的僕人！
PS|86|3|主啊，求你憐憫我， 因我終日求告你。
PS|86|4|主啊，求你使你的僕人心裏歡喜， 因為我的心仰望你。
PS|86|5|主啊，你本為良善，樂於饒恕人， 以豐盛的慈愛對待凡求告你的人。
PS|86|6|耶和華啊，求你側耳聽我的禱告， 留心聽我懇求的聲音。
PS|86|7|我在患難之日要求告你， 因為你必應允我。
PS|86|8|主啊，諸神之中沒有可與你相比的， 你的作為也無以為比。
PS|86|9|主啊，你所造的萬民都要來敬拜你， 他們要榮耀你的名。
PS|86|10|因你本為大，且行奇妙的事， 惟獨你是上帝。
PS|86|11|耶和華啊，求你將你的道指教我， 我要照你的真理而行； 求你使我專心敬畏你的名！
PS|86|12|主－我的上帝啊，我要一心稱謝你； 我要榮耀你的名，直到永遠。
PS|86|13|因為你的慈愛在我身上浩大， 你救了我的性命免入陰間的深處。
PS|86|14|上帝啊，驕傲的人起來攻擊我， 又有一群強橫的人尋索我的命； 他們沒有將你放在眼裏。
PS|86|15|主啊，你是有憐憫，有恩惠的上帝， 不輕易發怒，並有豐盛的慈愛和信實。
PS|86|16|求你轉向我，憐憫我， 將你的力量賜給僕人，拯救你使女的兒子。
PS|86|17|求你向我顯出恩待我的憑據， 使恨我的人看見就羞愧， 因為你－耶和華幫助我，安慰了我。
PS|87|1|耶和華所立的根基在聖山上。
PS|87|2|耶和華愛 錫安 的門， 勝於愛 雅各 一切的住處。
PS|87|3|上帝的城啊， 有榮耀的事是指著你說的。（細拉）
PS|87|4|我要提起 拉哈伯 和 巴比倫 人， 是在認識我之中的； 看哪， 非利士 、 推羅 和 古實 人， 個個生在那裏。
PS|87|5|論到 錫安 ，必有話說： 「這一個、那一個都生在其中」； 而且至高者必親自堅立這城。
PS|87|6|當耶和華記錄萬民的時候， 他要寫出人的出生地。（細拉）
PS|87|7|歌唱的、跳舞的，都要說： 「我的泉源都在你裏面。」
PS|88|1|耶和華－拯救我的上帝啊， 我晝夜在你面前呼求；
PS|88|2|願我的禱告達到你面前， 求你側耳聽我的懇求！
PS|88|3|因為我心裏滿了患難， 我的性命臨近陰間；
PS|88|4|我與下到地府的人同列， 如同無人幫助的人一樣。
PS|88|5|我被丟在死人中， 好像被殺的人躺在墳墓裏， 不再被你記得， 與你的手隔絕了。
PS|88|6|你把我放在極深的地府裏， 在黑暗地，在深處。
PS|88|7|你的憤怒重壓我身， 你用一切的波浪困住我。（細拉）
PS|88|8|你把我所認識的人隔在遠處， 使我為他們所憎惡； 我被拘禁，不能出來。
PS|88|9|我的眼睛因困苦而昏花； 耶和華啊，我天天求告你，向你舉手。
PS|88|10|你豈要行奇事給死人看嗎？ 陰魂還能起來稱謝你嗎？（細拉）
PS|88|11|你的慈愛豈能在墳墓裏被人述說嗎？ 你的信實豈能在冥府 被人傳揚嗎？
PS|88|12|你的奇事豈能在幽暗裏為人所知嗎？ 你的公義豈能在遺忘之地為人所識嗎？
PS|88|13|耶和華啊，至於我，我要呼求你； 每早晨，我的禱告要達到你面前。
PS|88|14|耶和華啊，你為何丟棄我？ 為何轉臉不顧我？
PS|88|15|我自幼受苦，幾乎死亡； 你使我驚恐，煩亂不安。
PS|88|16|你的烈怒漫過我身， 你用驚嚇把我除滅。
PS|88|17|這些如水終日環繞我， 一起圍困我。
PS|88|18|你把我的良朋密友隔在遠處， 使我所認識的人都在黑暗裏 。
PS|89|1|我要歌唱耶和華的慈愛，直到永遠， 我要用口將你的信實傳到萬代。
PS|89|2|因我曾說：「你的慈愛必建立到永遠， 你的信實必堅立在天上。」
PS|89|3|「我與我所揀選的人立了約， 向我的僕人 大衛 起了誓：
PS|89|4|『我要堅立你的後裔，直到永遠， 要建立你的寶座，直到萬代。』」（細拉）
PS|89|5|耶和華啊，諸天要稱謝你的奇事； 在聖者的會中，要稱謝你的信實。
PS|89|6|因在天空誰能比耶和華呢？ 諸神之中，誰能像耶和華呢？
PS|89|7|在聖者的會中，他是大有威嚴的上帝， 比在他四圍所有的更可畏懼。
PS|89|8|耶和華－萬軍之上帝啊， 哪一個大能者像耶和華？ 你的信實在你四圍。
PS|89|9|你管轄海的狂傲； 波浪翻騰，你使它平靜了。
PS|89|10|你打碎了 拉哈伯 ，使牠如遭刺殺的人； 你用大能的膀臂打散了你的仇敵。
PS|89|11|天屬你，地也屬你； 世界和其中所充滿的都為你所建立。
PS|89|12|南北為你所創造； 他泊 和 黑門 都因你的名歡呼。
PS|89|13|你有大能的膀臂， 你的手有力，你的右手也高舉。
PS|89|14|公義和公平是你寶座的根基， 慈愛和信實行在你前面。
PS|89|15|知道向你歡呼的，那民有福了！ 耶和華啊，他們要行走在你臉的光中。
PS|89|16|他們因你的名終日歡樂， 因你的公義得以高舉。
PS|89|17|你是他們力量的榮耀。 我們的角必被高舉，因為你喜愛我們。
PS|89|18|我們的盾牌是耶和華， 我們的王是 以色列 的聖者。
PS|89|19|當時，你在異象中吩咐你的聖民，說： 「我已把救助之力加在壯士身上， 高舉了那從百姓中所揀選的人。
PS|89|20|我尋得我的僕人 大衛 ， 用我的聖膏膏他。
PS|89|21|我的手必使他堅立， 我的膀臂也必堅固他。
PS|89|22|仇敵必不勒索他， 兇惡之子也不苦害他。
PS|89|23|我要在他面前打碎他的敵人， 擊殺那些恨他的人。
PS|89|24|我的信實和我的慈愛要與他同在； 因我的名，他的角必被高舉。
PS|89|25|我要使他的手伸到海上， 右手伸到河上。
PS|89|26|他要稱呼我說：『你是我的父， 是我的上帝，是拯救我的磐石。』
PS|89|27|我也要立他為長子， 為世上最高的君王。
PS|89|28|我要為他存留我的慈愛，直到永遠， 我與他所立的約必堅定不移。
PS|89|29|我也要使他的後裔存到永遠， 使他的寶座如天之久。
PS|89|30|「倘若他的子孫離棄我的律法， 不照我的典章行，
PS|89|31|背棄我的律例， 不遵守我的誡命，
PS|89|32|我就要用杖責罰他們的過犯， 用鞭責罰他們的罪孽。
PS|89|33|只是我不將我的慈愛全然收回， 也不叫我的信實廢除。
PS|89|34|我必不毀損我的約， 也不改變我口中所出的話。
PS|89|35|我僅此一次指著自己的神聖起誓， 我絕不向 大衛 說謊！
PS|89|36|他的後裔要存到永遠， 他的寶座在我面前如太陽，
PS|89|37|又如月亮永遠堅立； 天上的見證是確實的。」（細拉）
PS|89|38|但你惱怒你的受膏者， 拒絕他，離棄了他。
PS|89|39|你厭惡與你僕人所立的約， 將他的冠冕踐踏於地。
PS|89|40|你拆毀了他一切的圍牆， 使他的堡壘變為廢墟。
PS|89|41|過路的人都搶奪他， 他成了鄰邦羞辱的對象。
PS|89|42|你高舉了他敵人的右手， 使他所有的仇敵歡喜。
PS|89|43|你叫他的刀劍捲刃， 使他在戰爭中站立不住。
PS|89|44|你使他的光輝止息， 將他的寶座推倒於地。
PS|89|45|你減少他年輕的日子， 又使他蒙羞。（細拉）
PS|89|46|耶和華啊，這要到幾時呢？ 你要隱藏自己到永遠嗎？ 你的憤怒如火焚燒要到幾時呢？
PS|89|47|求你想念我的生命是何等短暫。 你創造世人，要使他們歸於何等的虛空呢？
PS|89|48|誰能常活不見死亡、 救自己脫離陰間的掌控呢？（細拉）
PS|89|49|主啊，你從前憑你的信實 向 大衛 起誓要施行的慈愛在哪裏呢？
PS|89|50|主啊，求你記念僕人們所受的羞辱， 記念我怎樣將萬族所加的羞辱都放在我的胸懷。
PS|89|51|耶和華啊，這是你仇敵所加的羞辱， 羞辱了你受膏者的腳蹤。
PS|89|52|耶和華是應當稱頌的，直到永遠。 阿們！阿們！ 神人摩西的祈禱。
PS|90|1|主啊，你世世代代作我們的居所。
PS|90|2|諸山未曾生出， 地與世界你未曾造成， 從亙古到永遠，你是上帝。
PS|90|3|你使人歸於塵土，說： 「世人哪，你們要歸回。」
PS|90|4|在你看來，千年如已過的昨日， 又如夜間的一更。
PS|90|5|你叫他們如水沖去， 他們如睡一覺。 早晨，他們如生長的草；
PS|90|6|早晨發芽生長， 晚上割下枯乾。
PS|90|7|我們因你的怒氣而消滅， 因你的憤怒而驚惶。
PS|90|8|你將我們的罪孽擺在你面前， 將我們的隱惡擺在你面光之中。
PS|90|9|我們經過的日子，都在你震怒之下， 我們度盡的年歲，好像一聲嘆息。
PS|90|10|我們一生的年日是七十歲， 若是強壯可到八十歲； 但其中所矜誇的不過是勞苦愁煩， 轉眼即逝，我們便如飛而去。
PS|90|11|誰曉得你怒氣的權勢？ 誰因著敬畏你而曉得你的憤怒呢？
PS|90|12|求你指教我們怎樣數算自己的日子， 好叫我們得著智慧的心。
PS|90|13|耶和華啊，我們要等到幾時呢？ 求你轉回，憐憫你的僕人們。
PS|90|14|求你使我們早早飽得你的慈愛， 好叫我們一生一世歡呼喜樂。
PS|90|15|求你照著你使我們受苦的日子， 和我們遭難的年歲，使我們喜樂。
PS|90|16|願你的作為向你僕人們顯現， 願你的榮耀向他們子孫顯明。
PS|90|17|願主－我們上帝的恩寵歸於我們身上。 願你堅立我們手所做的工， 我們手所做的工，願你堅立。
PS|91|1|住在至高者隱密處的， 必住在全能者的蔭下。
PS|91|2|我要向耶和華說： 「我的避難所、我的山寨、 我的上帝，你是我所倚靠的。」
PS|91|3|他必救你脫離捕鳥者的羅網 和毀滅人的瘟疫。
PS|91|4|他必用自己的翎毛遮蔽你； 你要投靠在他翅膀底下， 他的信實是大小的盾牌。
PS|91|5|你必不怕黑夜的驚駭， 或是白日飛的箭，
PS|91|6|也不怕黑夜流行的瘟疫， 或是午間滅人的災害。
PS|91|7|雖有千人仆倒在你旁邊， 萬人仆倒在你右邊， 這災卻不得臨近你。
PS|91|8|你惟親眼觀看， 見惡人遭報。
PS|91|9|因為耶和華是我的避難所， 你以至高者為居所，
PS|91|10|禍患必不臨到你， 災害也不挨近你的帳棚。
PS|91|11|因他要為你命令他的使者， 在你所行的一切道路上保護你。
PS|91|12|他們要用手托住你， 免得你的腳碰在石頭上。
PS|91|13|你要踹踏獅子和毒蛇， 踐踏少壯獅子和大蛇。
PS|91|14|「因為他專心愛我，我要搭救他； 因為他認識我的名，我要把他安置在高處。
PS|91|15|他若求告我，我就應允他； 他在急難中，我與他同在； 我要搭救他，使他尊貴。
PS|91|16|我要使他享足長壽， 將我的救恩顯明給他。」
PS|92|1|這是多麼好啊！ 稱謝耶和華， 歌頌你至高者的名，
PS|92|2|早晨傳揚你的慈愛， 每夜傳揚你的信實。
PS|92|3|用十弦的樂器和瑟， 用琴優雅的聲音；
PS|92|4|因你－耶和華藉著你的作為使我高興， 我要因你手的工作歡呼。
PS|92|5|耶和華啊，你的工作何其大！ 你的心思極其深！
PS|92|6|畜牲一般的人不曉得， 愚昧人也不明白。
PS|92|7|惡人雖茂盛如草， 作惡的人雖全都興旺， 他們卻要滅亡， 直到永遠。
PS|92|8|耶和華啊，惟有你是至高， 直到永遠。
PS|92|9|耶和華啊，看哪，你的仇敵， 看哪，你的仇敵都要滅亡； 作惡的全都要離散。
PS|92|10|你卻高舉了我的角，如野牛的角； 我是被新油膏抹的。
PS|92|11|我的眼睛看見我的仇敵遭報， 我的耳朵聽見那些起來攻擊我的惡人受罰。
PS|92|12|義人要興旺如棕樹， 生長如 黎巴嫩 的香柏樹。
PS|92|13|他們栽於耶和華的殿中， 發旺在我們上帝的院裏。
PS|92|14|他們髮白的時候仍結果子， 而且鮮美多汁，
PS|92|15|好顯明耶和華是正直的； 他是我的磐石，在他毫無不義。
PS|93|1|耶和華作王！ 他以威嚴為衣穿上； 耶和華以能力為衣，以能力束腰， 世界就堅定，不得動搖。
PS|93|2|你的寶座從太初立定， 你從亙古就有。
PS|93|3|耶和華啊，大水揚起， 大水發聲，大水澎湃。
PS|93|4|耶和華在高處大有威力， 勝過諸水的響聲，洋海的大浪。
PS|93|5|耶和華啊，你的法度最為確定； 你的殿宜稱為聖，直到永遠。
PS|94|1|耶和華啊，你是伸冤的上帝； 伸冤的上帝啊，求你發出光來！
PS|94|2|審判世界的主啊，求你挺身而立， 使驕傲的人受應得的報應！
PS|94|3|耶和華啊，惡人誇勝要到幾時呢？ 要到幾時呢？
PS|94|4|他們咆哮，說狂妄的話， 作惡的人全都誇耀自己。
PS|94|5|耶和華啊，他們強壓你的百姓， 苦害你的產業。
PS|94|6|他們殺死寡婦和寄居的人， 又殺害孤兒。
PS|94|7|他們說：「耶和華必不看見， 雅各 的上帝必不留意。」
PS|94|8|百姓中像畜牲一般的人當思想， 你們愚昧人要到幾時才有智慧呢？
PS|94|9|造耳朵的，難道自己聽不見嗎？ 造眼睛的，難道自己看不見嗎？
PS|94|10|管教列國的，就是叫人得知識的， 難道自己不懲治人嗎？
PS|94|11|耶和華知道人的意念是虛妄的。
PS|94|12|耶和華啊，你所管教、 用律法教導的人有福了！
PS|94|13|你使他在遭難的日子仍得平安， 直到為惡人挖好了坑。
PS|94|14|因為耶和華必不丟棄他的百姓， 也不離棄他的產業。
PS|94|15|審判要回復公義， 心裏正直的，都必跟隨它。
PS|94|16|誰肯為我起來攻擊邪惡的？ 誰肯為我站起抵擋作惡的？
PS|94|17|若不是耶和華幫助我， 我早就住在寂靜 之中了。
PS|94|18|我若說：「我失了腳！」 耶和華啊，你的慈愛必扶持我。
PS|94|19|我心裏多憂多疑， 你的安慰使我歡樂。
PS|94|20|那藉著律例玩弄奸惡、 以權位肆行殘害的，豈能與你交往呢？
PS|94|21|他們大家聚集攻擊義人， 將無辜的人定了死罪。
PS|94|22|但耶和華向來作我的碉堡， 我的上帝作了我投靠的磐石。
PS|94|23|他叫他們的罪孽歸到自己身上， 要因他們的邪惡剪除他們； 耶和華－我們的上帝要把他們剪除。
PS|95|1|來啊，我們要向耶和華歌唱， 向拯救我們的磐石歡呼！
PS|95|2|我們要以感謝來到他面前， 用詩歌向他歡呼！
PS|95|3|因耶和華是偉大的上帝， 是超越萬神的大君王。
PS|95|4|地的深處在他手中； 山的高峰也屬他。
PS|95|5|海洋屬他，是他造的； 旱地也是他手造成的。
PS|95|6|來啊，我們要俯伏敬拜， 在造我們的耶和華面前跪拜。
PS|95|7|因為他是我們的上帝； 我們是他草場的百姓，是他手中的羊。 惟願你們今天聽他的話！
PS|95|8|你們不可硬著心，像在 米利巴 ， 就是在曠野 瑪撒 的日子。
PS|95|9|那時，你們的祖宗試我，探我， 並且觀看我的作為。
PS|95|10|四十年之久，我厭煩那世代，說： 「這是心裏迷糊的百姓， 竟不知道我的道路！」
PS|95|11|所以，我在怒中起誓： 「他們斷不可進入我的安息！」
PS|96|1|你們要向耶和華唱新歌！ 全地都要向耶和華歌唱！
PS|96|2|要向耶和華歌唱，稱頌他的名！ 天天傳揚他的救恩！
PS|96|3|在列國中述說他的榮耀！ 在萬民中述說他的奇事！
PS|96|4|因耶和華本為大，當受極大的讚美； 他在萬神之上，當受敬畏。
PS|96|5|因萬民的神明都屬虛無； 惟獨耶和華創造諸天。
PS|96|6|有尊榮和威嚴在他面前， 有能力與華美在他聖所。
PS|96|7|民中的萬族啊，要將榮耀、能力歸給耶和華， 都歸給耶和華！
PS|96|8|要將耶和華的名所當得的榮耀歸給他， 拿供物來進入他的院宇。
PS|96|9|當敬拜神聖榮耀的耶和華 ， 全地都要在他面前戰抖！
PS|96|10|要在列國中說：「耶和華作王了！ 世界堅定，不得動搖； 他要按公正審判萬民。」
PS|96|11|願天歡喜，願地快樂！ 願海和其中所充滿的澎湃！
PS|96|12|願田和其中所有的都歡樂！ 那時，林中的樹木都要在耶和華面前歡呼。
PS|96|13|因為他來了，他來要審判全地。 他要按公義審判世界， 按信實審判萬民。
PS|97|1|耶和華作王！願地快樂！ 願眾海島歡喜！
PS|97|2|密雲和幽暗在他四圍， 公義和公平是他寶座的根基。
PS|97|3|烈火在他前頭行， 燒滅他四圍的敵人。
PS|97|4|他的閃電光照世界， 大地看見就震動。
PS|97|5|諸山見耶和華的面， 就是全地之主的面，就如蠟熔化。
PS|97|6|諸天表明他的公義， 萬民看見他的榮耀。
PS|97|7|願所有事奉雕刻偶像、 靠虛無神明自誇的，都蒙羞愧。 萬神哪，你們都當拜他。
PS|97|8|耶和華啊，因你的判斷， 錫安 聽見就歡喜； 猶大 的城鎮 也都快樂。
PS|97|9|因為你－耶和華至高，超乎全地； 受尊崇，遠超萬神之上。
PS|97|10|你們愛耶和華的，都當恨惡罪惡； 他保護聖民的性命， 搭救他們脫離惡人的手。
PS|97|11|散播亮光是為義人 ， 喜樂歸於心裏正直的人。
PS|97|12|義人哪，你們當靠耶和華歡喜， 當頌揚他神聖的名字 。
PS|98|1|你們要向耶和華唱新歌！ 因為他行過奇妙的事， 他的右手和聖臂施行救恩。
PS|98|2|耶和華顯明了他的救恩， 在列國眼前顯出公義；
PS|98|3|記念他對 以色列 家的慈愛和信實。 地的四極都看見我們上帝的救恩。
PS|98|4|全地都要向耶和華歡呼， 要揚聲，歡唱，歌頌！
PS|98|5|用琴歌頌耶和華， 用琴和詩歌的聲音歌頌他！
PS|98|6|用號筒和角聲， 在大君王耶和華面前歡呼！
PS|98|7|願海和其中所充滿的澎湃， 願世界和住在其間的發聲。
PS|98|8|願大水拍掌， 願諸山在耶和華面前一同歡呼；
PS|98|9|因為他來要審判全地。 他要按公義審判世界， 按公正審判萬民。
PS|99|1|耶和華作王，萬民當戰抖！ 他坐在基路伯的寶座上，地當動搖。
PS|99|2|耶和華在 錫安 為大， 他超越萬民之上。
PS|99|3|願他們頌揚他大而可畏的名， 他本為聖！
PS|99|4|喜愛公平、大能的王啊，你堅立公正， 在 雅各 中施行公平和公義。
PS|99|5|當尊崇耶和華－我們的上帝， 在他腳凳前下拜。 他本為聖！
PS|99|6|在他的祭司中有 摩西 和 亞倫 ， 在求告他名的人中有 撒母耳 。 他們求告耶和華，他就應允他們。
PS|99|7|他在雲柱中向他們說話， 他們遵守他的法度和他所賜給他們的律例。
PS|99|8|耶和華－我們的上帝啊，你應允了他們； 你是赦免他們的上帝， 卻按他們所做的報應他們。
PS|99|9|當尊崇耶和華－我們的上帝， 在他的聖山下拜， 因為耶和華－我們的上帝本為聖！
PS|100|1|普天下當向耶和華歡呼！
PS|100|2|當樂意事奉耶和華， 當歡唱來到他面前！
PS|100|3|當認識耶和華是上帝！ 我們是他造的，也是屬他的； 我們是他的民，是他草場的羊。
PS|100|4|當稱謝進入他的門， 當讚美進入他的院。 當感謝他，稱頌他的名！
PS|100|5|因為耶和華本為善； 他的慈愛存到永遠， 他的信實直到萬代。
PS|101|1|我要歌唱慈愛和公平， 耶和華啊，我要向你歌頌！
PS|101|2|我要用智慧行完全的道。 你幾時到我這裏來呢？ 我要以純正的心行在我家中。
PS|101|3|邪僻的事，我都不擺在我眼前； 悖逆的人所做的事，我甚恨惡， 不容沾在我身上。
PS|101|4|歪曲的心思，我必遠離； 邪惡的事情，我不知道。
PS|101|5|暗中讒害他鄰居的，我必將他滅絕； 眼目高傲、心裏驕縱的，我必不容忍。
PS|101|6|我眼要看顧地上誠實可靠的人，使他們與我同住； 行正直路的，他要侍候我。
PS|101|7|行詭詐的，必不得住在我家裏； 說謊言的，必不得立在我眼前。
PS|101|8|我每日早晨要滅絕地上所有的惡人， 把作惡的從耶和華的城裏全都剪除。
PS|102|1|耶和華啊，求你聽我的禱告， 願我的呼求達到你面前！
PS|102|2|我急難的日子，求你不要轉臉不顧我！ 我呼求的日子，求你向我側耳，快快應允我！
PS|102|3|因為我的年日在煙中消失 ， 我的骨頭如火把燒著。
PS|102|4|我的心如草被踩碎而枯乾， 甚至我忘記吃飯。
PS|102|5|因我嘆息的聲音， 我的肉緊貼骨頭。
PS|102|6|我如同曠野的鵜鶘， 好像荒地的貓頭鷹。
PS|102|7|我清醒難以入眠， 如同房頂上孤單的麻雀。
PS|102|8|我的仇敵整日辱罵我， 向我叫號的人指著我賭咒。
PS|102|9|我吃灰燼如同吃飯， 我喝的有眼淚攙雜。
PS|102|10|這都因你的惱恨和憤怒， 你把我舉起，又把我摔下。
PS|102|11|我的年日如夕陽， 我也如草枯乾。
PS|102|12|惟你－耶和華必永遠坐在寶座上， 你的名 存到萬代。
PS|102|13|你必起來憐憫 錫安 ； 因現在是可憐它的時候， 因所定的日期已經到了。
PS|102|14|你的僕人們喜愛 錫安 的石頭， 憐憫它的塵土。
PS|102|15|列國要敬畏耶和華的名， 地上眾王都要敬畏你的榮耀。
PS|102|16|因為耶和華建造了 錫安 ， 在他的榮耀裏顯現。
PS|102|17|他垂聽窮乏人的禱告， 不藐視他們的祈求。
PS|102|18|這必為後代的人記下， 將來受造的百姓要讚美耶和華。
PS|102|19|因為他從至高的聖所垂看； 耶和華從天向地觀看，
PS|102|20|要垂聽被囚之人的嘆息， 要釋放將死的人，
PS|102|21|使人在 錫安 傳揚耶和華的名， 在 耶路撒冷 傳揚讚美他的話，
PS|102|22|就是在萬民和列國 聚集事奉耶和華的時候。
PS|102|23|他使我的力量半途衰弱， 使我的年日短少。
PS|102|24|我說：「我的上帝啊， 不要使我中年去世。 你的年數世世無窮！」
PS|102|25|你起初立了地的根基， 天也是你手所造的。
PS|102|26|天地都會消滅，你卻長存； 天地都會像外衣漸漸舊了。 你要將天地如內衣更換， 天地就都改變了。
PS|102|27|惟有你永不改變， 你的年數沒有窮盡。
PS|102|28|你僕人的子孫要安然居住， 他們的後裔要堅立在你面前。
PS|103|1|我的心哪，你要稱頌耶和華！ 凡在我裏面的，都要稱頌他的聖名！
PS|103|2|我的心哪，你要稱頌耶和華！ 不可忘記他一切的恩惠！
PS|103|3|他赦免你一切的罪孽， 醫治你一切的疾病。
PS|103|4|他救贖你的命脫離地府， 以仁愛和憐憫為你的冠冕。
PS|103|5|他用美物使你的生命 得以滿足， 以致你如鷹返老還童。
PS|103|6|耶和華施行公義， 為所有受欺壓的人伸冤。
PS|103|7|他使 摩西 知道他的法則， 使 以色列 人曉得他的作為。
PS|103|8|耶和華有憐憫，有恩惠， 不輕易發怒，且有豐盛的慈愛。
PS|103|9|他不長久責備， 也不永遠懷怒。
PS|103|10|他沒有按我們的罪待我們， 也沒有照我們的罪孽報應我們。
PS|103|11|天離地何等的高， 他的慈愛向敬畏他的人也是何等的大！
PS|103|12|東離西有多遠， 他叫我們的過犯離我們也有多遠！
PS|103|13|父親怎樣憐憫他的兒女， 耶和華也怎樣憐憫敬畏他的人！
PS|103|14|因為他知道我們的本體， 思念我們不過是塵土。
PS|103|15|至於世人，他的年日如草一樣。 他興旺如野地的花，
PS|103|16|經風一吹，就歸無有， 它的原處也不再認識它。
PS|103|17|但耶和華的慈愛歸於敬畏他的人， 從亙古到永遠； 他的公義也歸於子子孫孫，
PS|103|18|就是那些遵守他的約、 記念他的訓詞而遵行的人。
PS|103|19|耶和華在天上立定寶座， 他的國統管萬有。
PS|103|20|聽從他命令、成全他旨意、 有大能的天使啊，你們都要稱頌耶和華！
PS|103|21|你們行他所喜悅的， 作他諸軍，作他僕役的啊，都要稱頌耶和華！
PS|103|22|你們一切被他造的， 在他所治理的各處， 都要稱頌耶和華！ 我的心哪，你要稱頌耶和華！
PS|104|1|我的心哪，你要稱頌耶和華！ 耶和華－我的上帝啊，你為至大！ 你以尊榮威嚴為衣，
PS|104|2|披上亮光，如披外袍， 鋪張穹蒼，如鋪幔子，
PS|104|3|在水中立樓閣的棟梁， 用雲彩為車輦， 藉著風的翅膀而行，
PS|104|4|以風為使者， 以火焰為僕役，
PS|104|5|將地立在根基上， 使地永不動搖。
PS|104|6|你用深水遮蓋地面，猶如衣裳； 諸水高過山嶺。
PS|104|7|你的斥責一發，水就奔逃； 你的雷聲一發，水就奔流。
PS|104|8|諸山上升，諸谷下沉， 歸你為它所立定之地。
PS|104|9|你定了界限，使水不能超越， 不再轉回淹沒大地。
PS|104|10|耶和華使泉源湧在山谷， 流在山間，
PS|104|11|使野地的走獸有水喝， 野驢得解其渴。
PS|104|12|天上的飛鳥在水旁住宿， 在枝幹間啼叫。
PS|104|13|他從樓閣中澆灌山嶺； 因他作為的功效，地就豐足。
PS|104|14|他使草生長，給牲畜吃， 使菜蔬生長，供給人用 ， 使人從地裏得食物，
PS|104|15|得酒能悅人心， 得油能潤人面， 得糧能養人心。
PS|104|16|佳美的樹木， 就是耶和華所栽種的 黎巴嫩 的香柏樹， 都滿了汁漿。
PS|104|17|雀鳥在其上搭窩， 鸛以松樹 為家。
PS|104|18|高山為野山羊的居所， 巖石為石獾的藏身處。
PS|104|19|你安置月亮以定季節， 太陽自知沉落。
PS|104|20|你造黑暗為夜， 林中的百獸就都爬出來。
PS|104|21|少壯獅子吼叫覓食， 向上帝尋求食物。
PS|104|22|太陽一出，獸就躲避， 躺臥在洞裏。
PS|104|23|人出去做工， 勞碌直到晚上。
PS|104|24|耶和華啊，你所造的何其多！ 都是你用智慧造成的， 全地遍滿了你所造之物。
PS|104|25|那裏有海，又大又廣， 其中有無數的動物， 大小活物都有。
PS|104|26|那裏有船行走， 有你所造的 力威亞探 悠游在其中。
PS|104|27|這些都仰望你按時給牠們食物。
PS|104|28|你給牠們，牠們就拾起來； 你張手，牠們就飽得美食。
PS|104|29|你轉臉，牠們就驚惶； 你收回牠們的氣，牠們就死亡，歸於塵土。
PS|104|30|你差遣你的靈，牠們就受造； 你使地面更換為新。
PS|104|31|願耶和華的榮耀存到永遠！ 願耶和華喜愛自己所造的！
PS|104|32|他看地，地便震動； 他摸山，山就冒煙。
PS|104|33|我一生要向耶和華唱詩！ 我還活的時候，要向我的上帝歌頌！
PS|104|34|願他悅納我的默念！ 我要因耶和華歡喜！
PS|104|35|願罪人從世上消滅！ 願惡人歸於無有！ 我的心哪，你要稱頌耶和華！ 哈利路亞 ！
PS|105|1|你們要稱謝耶和華，求告他的名， 在萬民中傳揚他的作為！
PS|105|2|要向他唱詩，向他歌頌， 述說他一切奇妙的作為！
PS|105|3|要誇耀他的聖名！ 願尋求耶和華的人心中歡喜！
PS|105|4|要尋求耶和華與他的能力， 時常尋求他的面。
PS|105|5|他僕人 亞伯拉罕 的後裔， 他所揀選 雅各 的子孫哪， 要記念他奇妙的作為和他的奇事， 並他口中的判語。
PS|105|6|
PS|105|7|他是耶和華－我們的上帝， 全地都有他的判斷。
PS|105|8|他記念他的約，直到永遠； 記念他吩咐的話，直到千代，
PS|105|9|就是與 亞伯拉罕 所立的約， 向 以撒 所起的誓。
PS|105|10|他將這約向 雅各 定為律例， 向 以色列 定為永遠的約，
PS|105|11|說：「我必將 迦南 地賜給你， 作你們應得的產業。」
PS|105|12|當時，他們人丁有限， 數目稀少，在那地寄居。
PS|105|13|他們從這邦遊到那邦， 從這國去到另一民族。
PS|105|14|他不容人欺負他們， 為他們的緣故責備君王：
PS|105|15|「不可傷害我的受膏者， 也不可惡待我的先知。」
PS|105|16|他命饑荒降在那地， 斷絕日用的糧食 ，
PS|105|17|在他們以先差遣一個人前往， 約瑟 被賣為奴。
PS|105|18|人用腳鐐傷他的腳， 他被鐵的項鏈捆鎖。
PS|105|19|耶和華的話試煉他， 直等所說的應驗了。
PS|105|20|王差人將他解開， 治理萬民的把他釋放，
PS|105|21|立他為王家之主， 掌管他一切所有的，
PS|105|22|使他隨意捆綁他的臣宰， 將智慧教導他的長老。
PS|105|23|以色列 也到了 埃及 ， 雅各 在 含 地寄居。
PS|105|24|耶和華使他的百姓生養眾多， 使他們比敵人強盛，
PS|105|25|他使敵人的心轉去恨他的百姓， 用詭計待他的僕人。
PS|105|26|他差遣他的僕人 摩西 和他所揀選的 亞倫 ，
PS|105|27|在敵人中間顯他的神蹟， 在 含 地顯他的奇事。
PS|105|28|他差遣黑暗，就有黑暗； 他們沒有違背他的話。
PS|105|29|他使 埃及 的水變為血， 令他們的魚死了。
PS|105|30|在他們的地上，青蛙多多滋生， 王宮的內室也是如此。
PS|105|31|他一吩咐，蒼蠅就成群飛來， 並有蚊子進入他們四境。
PS|105|32|他給他們降下冰雹為雨， 在他們的地上降下火焰。
PS|105|33|他擊打他們的葡萄樹和無花果樹， 毀壞他們境內的樹木。
PS|105|34|他一吩咐，就有蝗蟲蝻子上來， 不計其數，
PS|105|35|吃光他們地上各樣的菜蔬， 吞盡他們田地的出產。
PS|105|36|他又擊殺他們國內 所有的長子， 就是他們強壯時頭生的。
PS|105|37|他卻帶領自己的百姓帶著金子銀子出來， 他支派中沒有一個走不動的。
PS|105|38|他們出來的時候， 埃及 人就歡喜； 因為 埃及 人懼怕他們。
PS|105|39|他鋪張雲彩當遮蔽， 夜間使火光照。
PS|105|40|他們祈求，他就使鵪鶉飛來， 並用天上的糧食使他們飽足。
PS|105|41|他敲開磐石，水就湧出； 在乾旱之處，水流成河。
PS|105|42|這都因他記念他的聖言 和他的僕人 亞伯拉罕 。
PS|105|43|他帶領自己的百姓歡樂而出， 帶領自己的選民歡呼前往。
PS|105|44|他把列國的地賜給他們， 他們就承受萬民勞碌得來的，
PS|105|45|好讓他們遵他的律例， 守他的律法。 哈利路亞！
PS|106|1|哈利路亞！ 你們要稱謝耶和華，因他本為善， 他的慈愛永遠長存！
PS|106|2|誰能傳揚耶和華的大能？ 誰能表明他一切的美德？
PS|106|3|凡遵守公平、常行公義的， 這人有福了！
PS|106|4|耶和華啊，你恩待你百姓的時候，求你記念我； 你拯救他們的時候，求你眷顧我，
PS|106|5|好使我經歷你選民的福分， 享受你國民的喜樂， 與你的產業一同誇耀。
PS|106|6|我們與我們的祖宗一同犯罪， 偏邪行惡。
PS|106|7|我們的祖宗在 埃及 不明白你的奇事， 不記念你豐盛的慈愛， 反倒在 紅海 行了悖逆。
PS|106|8|然而，他因自己的名拯救他們， 為要彰顯他的大能。
PS|106|9|他斥責 紅海 ，海就乾了， 帶領他們走過深海，如走曠野。
PS|106|10|他拯救他們脫離恨他們之人的手， 從仇敵手中救贖他們。
PS|106|11|水淹沒他們的敵人， 沒有一個存留。
PS|106|12|那時，他們才信他的話， 歌唱讚美他。
PS|106|13|很快地，他們就忘了他的作為， 不仰望他的指引，
PS|106|14|反倒在曠野起了貪婪之心， 在荒地試探上帝。
PS|106|15|他將他們所求的賜給他們， 卻使他們心靈軟弱。
PS|106|16|他們在營中嫉妒 摩西 和耶和華的聖者 亞倫 。
PS|106|17|地就裂開，吞下 大坍 ， 掩蓋 亞比蘭 一夥的人。
PS|106|18|有火在他們黨中點燃， 有火焰燒燬了惡人。
PS|106|19|他們在 何烈山 造了牛犢， 叩拜鑄成的像，
PS|106|20|將他們榮耀的主 換為吃草之牛的像，
PS|106|21|忘了上帝－他們的救主， 就是曾在 埃及 行大事，
PS|106|22|在 含 地行奇事， 在 紅海 行可畏之事的那位。
PS|106|23|因此，他說要滅絕他們； 若非他所揀選的 摩西 在他面前站在破裂之處， 使他的憤怒轉消， 恐怕他就滅絕他們了。
PS|106|24|他們又藐視那美地， 不信他的話，
PS|106|25|在自己帳棚內發怨言， 不聽耶和華的聲音。
PS|106|26|所以他向他們起誓， 必叫他們倒在曠野，
PS|106|27|叫他們的後裔倒在列國之中， 分散在各地。
PS|106|28|他們又與 巴力‧毗珥 連合， 吃了祭死人的物。
PS|106|29|他們這樣行，惹耶和華發怒， 就有瘟疫流行在他們中間。
PS|106|30|那時， 非尼哈 起而干預， 瘟疫這才止息。
PS|106|31|那就算他為義， 世世代代，直到永遠。
PS|106|32|他們在 米利巴 水又惹耶和華發怒， 甚至 摩西 也因他們的緣故受虧損，
PS|106|33|是因他們觸怒了他的靈， 摩西就用嘴說了急躁的話。
PS|106|34|他們不照耶和華所吩咐的 滅絕外邦人，
PS|106|35|反倒與列國相交， 學習他們的行為，
PS|106|36|事奉他們的偶像， 這就成了自己的圈套。
PS|106|37|他們把自己的兒女祭祀鬼魔，
PS|106|38|流無辜人的血， 就是自己兒女的血， 用他們祭祀 迦南 的偶像， 那地就被血玷污了。
PS|106|39|這樣，他們被自己所做的玷污了， 在行為上犯了淫亂。
PS|106|40|耶和華的怒氣向他的百姓發作， 他憎惡自己的產業，
PS|106|41|將他們交在外邦人手裏， 恨他們的人就轄制他們。
PS|106|42|他們的仇敵欺壓他們， 他們伏在敵人手下。
PS|106|43|他屢次搭救他們， 他們卻圖謀悖逆， 就因自己的罪孽降為卑下。
PS|106|44|然而，他聽見他們哀告的時候， 就眷顧他們的急難，
PS|106|45|為了他們，他記念自己的約， 照他豐盛的慈愛改變心意，
PS|106|46|使他們在凡擄掠他們的人面前蒙憐憫。
PS|106|47|耶和華－我們的上帝啊，求你拯救我們， 從列國中召集我們， 我們好頌揚你的聖名， 以讚美你為誇勝。
PS|106|48|耶和華－ 以色列 的上帝是應當稱頌的， 從亙古直到永遠。 願全體百姓都說：「阿們！」 哈利路亞！
PS|107|1|你們要稱謝耶和華，因他本為善， 他的慈愛永遠長存！
PS|107|2|願耶和華救贖的百姓說這話， 就是他從敵人手中所救贖，
PS|107|3|從各地，從東從西， 從北從海那邊召集來的。
PS|107|4|他們在曠野、在荒地飄流， 找不到可居住的城，
PS|107|5|又飢又渴， 心裏發昏。
PS|107|6|於是他們在急難中哀求耶和華， 他就搭救他們脫離禍患，
PS|107|7|又領他們行走直路， 前往可居住的城。
PS|107|8|但願人因耶和華的慈愛 和他向人所做的奇事都稱謝他；
PS|107|9|因他使心裏渴慕的人得以滿足， 使飢餓的人得飽美食。
PS|107|10|那些坐在黑暗中、死蔭裏的人， 被困苦和鐵鏈捆鎖，
PS|107|11|是因他們違背上帝的言語， 藐視至高者的旨意。
PS|107|12|所以，他用勞苦制伏他們的心； 他們仆倒，無人扶助。
PS|107|13|於是他們在急難中哀求耶和華， 他就拯救他們脫離禍患。
PS|107|14|他從黑暗中、從死蔭裏領他們出來， 扯斷他們的捆綁。
PS|107|15|但願人因耶和華的慈愛 和他向人所做的奇事都稱謝他；
PS|107|16|因為他打破了銅門， 砍斷了鐵閂。
PS|107|17|愚妄人因自己叛逆的行徑 和自己的罪孽受苦楚。
PS|107|18|他們心裏厭惡各樣的食物， 就臨近死亡之門。
PS|107|19|於是他們在急難中哀求耶和華， 他就拯救他們脫離禍患。
PS|107|20|他發出自己的話語醫治他們， 救他們脫離陰府。
PS|107|21|但願人因耶和華的慈愛 和他向人所做的奇事都稱謝他。
PS|107|22|願他們以感謝為祭獻給他， 歡呼述說他的作為！
PS|107|23|那些搭船出海， 在大水中做生意的，
PS|107|24|他們看見耶和華的作為， 並他在深海中的奇事。
PS|107|25|他一出令，狂風捲起， 波浪翻騰。
PS|107|26|他們上到天空，下到海底， 他們的心因患難而消沉。
PS|107|27|他們搖搖晃晃，東倒西歪，好像醉酒的人， 他們的智慧無法可施。
PS|107|28|於是他們在急難中哀求耶和華， 他就領他們脫離禍患。
PS|107|29|他使狂風止息， 波浪平靜，
PS|107|30|既平靜了，他們就歡喜， 他就領他們到想要去的海港。
PS|107|31|但願人因耶和華的慈愛 和他向人所做的奇事都稱謝他。
PS|107|32|願他們在百姓的會中尊崇他， 在長老的座位上讚美他！
PS|107|33|他使江河變為曠野， 叫水泉變為乾涸之地，
PS|107|34|使肥沃之地變為荒蕪的鹽地， 都因當地居民的邪惡。
PS|107|35|他使曠野變為水潭， 叫旱地變為水泉，
PS|107|36|使飢餓的人住在那裏， 建造可居住的城，
PS|107|37|又種田地，栽葡萄園， 得享所出產的果實。
PS|107|38|他賜福給他們，使他們生養眾多， 也不叫他們的牲畜減少。
PS|107|39|但他們因欺壓、患難、愁苦， 人口減少而且卑微。
PS|107|40|他使貴族蒙羞受辱， 使他們迷失在荒涼無路之地；
PS|107|41|卻將窮乏人安置在高處，脫離苦難， 使他的家屬多如羊群。
PS|107|42|正直的人看見就歡喜， 罪孽之輩卻要啞口無言。
PS|107|43|凡有智慧的必在這些事上留心， 他必思想耶和華的慈愛。
PS|108|1|上帝啊，我心堅定； 我口 要唱詩歌頌！
PS|108|2|琴瑟啊，當醒起！ 我要喚起曙光！
PS|108|3|耶和華啊，我要在萬民中稱謝你， 在萬族中歌頌你！
PS|108|4|因為你的慈愛大過諸天， 你的信實達到穹蒼。
PS|108|5|上帝啊，願你崇高過於諸天！ 願你的榮耀高過全地！
PS|108|6|求你應允我，用右手施行拯救， 好讓你所親愛的人得救。
PS|108|7|上帝在他的聖所 說： 「我要歡樂； 要劃分 示劍 ， 丈量 疏割谷 。
PS|108|8|基列 是我的， 瑪拿西 是我的， 以法蓮 是護衛我頭的， 猶大 是我的權杖。
PS|108|9|摩押 是我的沐浴盆， 我要向 以東 扔鞋， 我必因勝 非利士 而歡呼。」
PS|108|10|誰能領我進堅固城？ 誰能引我到 以東 地？
PS|108|11|上帝啊，你真的丟棄了我們嗎？ 上帝啊，你不和我們的軍隊同去嗎？
PS|108|12|求你幫助我們攻擊敵人， 因為人的幫助是枉然的。
PS|108|13|我們倚靠上帝才得施展大能， 因為踐踏我們敵人的就是他。
PS|109|1|我所讚美的上帝啊， 求你不要閉口不言。
PS|109|2|因為惡人的嘴和詭詐人的口張開攻擊我， 他們用撒謊的舌頭對我說話。
PS|109|3|他們圍繞我，說怨恨的話， 又無故地攻打我。
PS|109|4|他們與我作對回報我的愛， 但我專心祈禱。
PS|109|5|他們向我以惡報善， 以恨報愛。
PS|109|6|求你派惡人轄制他， 派對頭站在他右邊！
PS|109|7|他受審判的時候， 願他背負罪名而出！ 願他的祈禱反成為罪！
PS|109|8|願他的年歲短少！ 願別人得他的職分！
PS|109|9|願他的兒女成為孤兒， 他的妻子成為寡婦！
PS|109|10|願他的兒女飄流討飯， 從荒涼之處出來求乞 ！
PS|109|11|願債主牢籠他一切所有的！ 願陌生人搶走他勞碌得來的！
PS|109|12|願無人向他佈施恩惠， 無人恩待他的孤兒！
PS|109|13|願他的後人斷絕， 名字被塗去，不傳於下代！
PS|109|14|願耶和華記得他祖宗的罪孽， 不塗去他母親的罪過！
PS|109|15|願這些罪常在耶和華面前！ 願他們的名字 從地上除滅！
PS|109|16|因為他從未想過要施恩， 卻迫害困苦貧窮的和傷心的人， 把他們處死。
PS|109|17|他愛咒罵，咒罵就臨到他； 他不喜愛祝福，祝福就遠離他！
PS|109|18|他拿咒罵當衣服穿上； 這咒罵就如水進到他裏面， 如油進入他骨頭。
PS|109|19|願這咒罵當他遮身的衣服， 作他經常束腰的帶子！
PS|109|20|這就是那些與我作對、用惡言議論我的人 從耶和華所受的報應。
PS|109|21|但是你，主－耶和華啊， 求你因你的名採取行動； 因你的慈愛美好，求你搭救我！
PS|109|22|因為我困苦貧窮， 內心受傷。
PS|109|23|我如日影偏斜而去， 如蝗蟲被抖出來。
PS|109|24|我因禁食，膝蓋軟弱； 我身體消瘦，不再豐潤。
PS|109|25|我受他們的羞辱， 他們看見我就搖頭。
PS|109|26|耶和華－我的上帝啊，求你幫助我， 照你的慈愛拯救我，
PS|109|27|好讓他們知道這是你的手， 是你－耶和華所做的事。
PS|109|28|任憑他們咒罵，你卻要賜福； 他們幾時起來就必蒙羞， 你的僕人卻要歡喜。
PS|109|29|願與我作對的人披戴羞辱！ 願他們以自己的羞愧作外袍遮身！
PS|109|30|我要用口極力稱謝耶和華， 我要在眾人中間讚美他；
PS|109|31|因為他必站在貧窮人的右邊， 救他脫離定他死罪的人。
PS|110|1|耶和華對我主說： 「你坐在我的右邊， 等我使你仇敵作你的腳凳。」
PS|110|2|耶和華必使你從 錫安 伸出你能力的權杖； 你務要在仇敵中掌權。
PS|110|3|你在聖山上 掌權的日子， 你的子民必甘心跟隨 ； 從晨曦初現， 你就有清晨 的甘露。
PS|110|4|耶和華起了誓，絕不改變： 「你是照著 麥基洗德 的體系永遠為祭司。」
PS|110|5|在你右邊的主， 當他發怒的日子，必打傷列王。
PS|110|6|他要審判列國， 屍首就佈滿各處； 他要痛擊遍地的領袖。
PS|110|7|他要喝路旁的河水， 因此必抬起頭來。
PS|111|1|哈利路亞！ 我要在正直人的大會和會眾中 一心稱謝耶和華。
PS|111|2|耶和華的作為本為大， 被所有喜愛的人所探尋。
PS|111|3|他所做的是尊榮和威嚴， 他的公義存到永遠。
PS|111|4|他行了奇事，使人記念； 耶和華有恩惠，有憐憫。
PS|111|5|他賜糧食給敬畏他的人， 他必永遠記念他的約。
PS|111|6|他向百姓顯出大能的作為， 將列國賜給他們為業。
PS|111|7|他手所做的信實公平， 他的訓詞全然可靠，
PS|111|8|是永永遠遠堅定的， 是按信實正直設立的。
PS|111|9|他向百姓施行救贖， 頒佈他的約，直到永遠； 他的名聖而可畏。
PS|111|10|敬畏耶和華是智慧的開端， 凡遵行他命令的有美好的見識。 耶和華是永遠當讚美的！
PS|112|1|哈利路亞！ 敬畏耶和華，甚喜愛他命令的， 這人有福了！
PS|112|2|他的後裔在世必強盛， 正直人的後代必蒙福。
PS|112|3|他的家中有金銀財寶， 他的義行存到永遠。
PS|112|4|正直人在黑暗中有光向他照耀， 他有恩惠，有憐憫，有公義。
PS|112|5|施恩與人、借貸與人、秉公處事的人 必享美福，
PS|112|6|他永不動搖。 義人被記念，直到永遠。
PS|112|7|他不懼怕兇惡的信息， 他的心堅定，倚靠耶和華。
PS|112|8|他的心確定，總不懼怕， 直到他看見敵人遭報。
PS|112|9|他施捨，賙濟貧窮， 他的義行存到永遠， 他的角必被高舉，大有榮耀。
PS|112|10|惡人看見就憤怒，必咬牙而消亡， 惡人的心願要歸於幻滅。
PS|113|1|哈利路亞！ 耶和華的僕人哪，你們要讚美， 讚美耶和華的名！
PS|113|2|耶和華的名是應當稱頌的， 從今時直到永遠！
PS|113|3|從日出之地到日落之處， 耶和華的名是應當讚美的！
PS|113|4|耶和華超乎萬國之上， 他的榮耀高過諸天。
PS|113|5|誰像耶和華－我們的上帝呢？ 他坐在至高之處，
PS|113|6|自己謙卑， 觀看天上地下的事。
PS|113|7|他從灰塵裏抬舉貧寒的人， 從糞堆中提拔貧窮的人，
PS|113|8|使他們與貴族同坐， 與本國的貴族同坐。
PS|113|9|他使不孕的婦女安居家中， 成為快樂的母親，兒女成群。 哈利路亞！
PS|114|1|以色列 出 埃及 ， 雅各 家離開說陌生語言之民時，
PS|114|2|猶大 作主的聖所， 以色列 為他所治理的國。
PS|114|3|滄海看見就奔逃， 約旦河 也倒流。
PS|114|4|大山踴躍如公羊， 小山跳舞如羔羊。
PS|114|5|滄海啊，你為何奔逃？ 約旦 哪，你為何倒流？
PS|114|6|大山哪，你為何踴躍如公羊？ 小山哪，你為何跳舞如羔羊？
PS|114|7|大地啊，在主的面前， 在 雅各 的上帝的面前，震動吧！
PS|114|8|他叫磐石變為水池， 使堅石變為泉源。
PS|115|1|耶和華啊，榮耀不要歸與我們， 不要歸與我們； 要因你的慈愛和信實歸在你的名下！
PS|115|2|為何讓列國說 「他們的上帝在哪裏」呢？
PS|115|3|但是，我們的上帝在天上， 萬事都隨自己的旨意而行。
PS|115|4|他們的偶像是金的，是銀的， 是人手所造的，
PS|115|5|有口卻不能言， 有眼卻不能看，
PS|115|6|有耳卻不能聽， 有鼻卻不能聞，
PS|115|7|有手卻不能摸， 有腳卻不能走， 有喉卻不能說話。
PS|115|8|造它們的要像它們一樣， 凡靠它們的也必如此。
PS|115|9|以色列 啊，要倚靠耶和華！ 他是人的幫助和盾牌。
PS|115|10|亞倫 家啊，要倚靠耶和華！ 他是人的幫助和盾牌。
PS|115|11|敬畏耶和華的人哪，要倚靠耶和華！ 他是人的幫助和盾牌。
PS|115|12|耶和華向來眷念我們， 他還要賜福， 賜福給 以色列 家， 賜福給 亞倫 家。
PS|115|13|凡敬畏耶和華的，無論大小， 主必賜福給他。
PS|115|14|願耶和華使你們 和你們的子孫日見增加。
PS|115|15|你們蒙了耶和華的福， 他是創造天地的主宰。
PS|115|16|天，是耶和華的天； 地，他卻給了世人。
PS|115|17|死人不能讚美耶和華， 下到寂靜 中的也都不能。
PS|115|18|但我們要稱頌耶和華， 從今時直到永遠。 哈利路亞！
PS|116|1|我愛耶和華， 因為他聽了我的聲音和我的懇求。
PS|116|2|他既向我側耳， 我一生要求告他。
PS|116|3|死亡的繩索勒住我， 陰間的痛苦抓住我， 我遭遇患難愁苦。
PS|116|4|那時，我求告耶和華的名： 「耶和華啊，求你救我！」
PS|116|5|耶和華有恩惠，有公義， 我們的上帝有憐憫。
PS|116|6|耶和華保護愚蒙的人； 我落到卑微的地步，他救了我。
PS|116|7|我的心哪！你要復歸安寧， 因為耶和華用厚恩待你。
PS|116|8|主啊，你救我的命脫離死亡， 使我的眼不再流淚， 使我的腳不致跌倒。
PS|116|9|我行在耶和華面前， 走在活人之地。
PS|116|10|我信，儘管我說： 「我受了極大的困苦。」
PS|116|11|我曾驚惶地說： 「人都是說謊的！」
PS|116|12|耶和華向我賞賜一切厚恩， 我拿甚麼來報答他呢？
PS|116|13|我要舉起救恩的杯， 稱揚耶和華的名。
PS|116|14|我要在他的全體百姓面前 向耶和華還我所許的願。
PS|116|15|在耶和華眼中， 聖民之死極為寶貴。
PS|116|16|耶和華啊，哦，我是你的僕人； 我是你的僕人，是你使女的兒子。 你已經解開我的捆索。
PS|116|17|我要以感謝為祭獻給你， 又要求告耶和華的名。
PS|116|18|我要在 耶路撒冷 當中， 在耶和華殿的院內， 在他的全體百姓面前， 向耶和華還我所許的願。 哈利路亞！
PS|116|19|
PS|117|1|萬國啊，你們要讚美耶和華！ 萬族啊，你們都要頌讚他！
PS|117|2|因為他向我們大施慈愛， 耶和華的信實存到永遠。 哈利路亞！
PS|118|1|你們要稱謝耶和華，因他本為善； 他的慈愛永遠長存！
PS|118|2|願 以色列 說： 「他的慈愛永遠長存！」
PS|118|3|願 亞倫 家說： 「他的慈愛永遠長存！」
PS|118|4|願敬畏耶和華的人說： 「他的慈愛永遠長存！」
PS|118|5|我在急難中求告耶和華， 耶和華就應允我，把我安置在寬闊之地。
PS|118|6|耶和華在我這邊 ，我必不懼怕， 人能把我怎麼樣呢？
PS|118|7|在那幫助我的人中，有耶和華幫助我， 所以我要看見那些恨我的人遭報。
PS|118|8|投靠耶和華， 強似倚賴人；
PS|118|9|投靠耶和華， 強似倚賴權貴。
PS|118|10|列邦圍繞我， 我靠耶和華的名必剿滅他們。
PS|118|11|他們圍繞我，圍困我， 我靠耶和華的名必剿滅他們。
PS|118|12|他們如同蜜蜂一般地圍繞我， 他們熄滅，好像燒荊棘的火； 我靠耶和華的名，必剿滅他們。
PS|118|13|你用力推我，要叫我跌倒， 但耶和華幫助了我。
PS|118|14|耶和華是我的力量，是我的詩歌， 他也成了我的拯救。
PS|118|15|在義人的帳棚裏，有歡呼拯救的聲音， 耶和華的右手施展大能。
PS|118|16|耶和華的右手高舉， 耶和華的右手施展大能。
PS|118|17|我不至於死，仍要存活， 並要傳揚耶和華的作為。
PS|118|18|耶和華雖嚴嚴地懲治我， 卻未曾將我交於死亡。
PS|118|19|給我敞開義門， 我要進去稱謝耶和華！
PS|118|20|這是耶和華的門， 義人要進去！
PS|118|21|我要稱謝你，因為你已經應允我， 又成了我的拯救！
PS|118|22|匠人所丟棄的石頭 已成了房角的頭塊石頭。
PS|118|23|這是耶和華所做的， 在我們眼中看為奇妙。
PS|118|24|這是耶和華所定的日子， 我們在其中要高興歡喜！
PS|118|25|耶和華啊，求你拯救 ！ 耶和華啊，求你使我們順利！
PS|118|26|奉耶和華的名來的是應當稱頌的！ 我們從耶和華的殿中為你們祝福！
PS|118|27|耶和華是上帝， 他光照了我們。 你們要用繩索把祭牲拴住， 直牽到壇角。
PS|118|28|你是我的上帝，我要稱謝你！ 我的上帝啊，我要尊崇你 ！
PS|118|29|你們要稱謝耶和華，因他本為善； 他的慈愛永遠長存！
PS|119|1|行為正直、遵行耶和華律法的， 這人有福了！
PS|119|2|遵守他的法度、一心尋求他的， 這人有福了！
PS|119|3|他們不做不義的事， 但遵行他的道。
PS|119|4|耶和華啊，你曾將你的訓詞吩咐我們， 為要我們切實遵守。
PS|119|5|但願我行事堅定， 得以遵守你的律例。
PS|119|6|我看重你的一切命令， 就不致羞愧。
PS|119|7|我學習你公義的典章， 要以正直的心稱謝你。
PS|119|8|我必遵守你的律例， 求你不要把我全然棄絕！
PS|119|9|青年要如何保持純潔呢？ 是要遵行你的話！
PS|119|10|我曾一心尋求你， 求你不要使我偏離你的命令。
PS|119|11|我將你的話藏在心裏， 免得我得罪你。
PS|119|12|耶和華啊，你是應當稱頌的！ 求你將你的律例教導我！
PS|119|13|我用嘴唇傳揚 你口中一切的典章。
PS|119|14|我喜愛你的法度， 如同喜愛一切的財物。
PS|119|15|我要默想你的訓詞， 看重你的道路。
PS|119|16|我要以你的律例為樂， 我不忘記你的話。
PS|119|17|求你用厚恩待你的僕人，使我存活， 我就遵守你的話。
PS|119|18|求你開我的眼睛， 使我看出你律法中的奇妙。
PS|119|19|我在地上是寄居的人， 求你不要向我隱藏你的命令！
PS|119|20|我時常切慕你的典章， 耗盡心力。
PS|119|21|受詛咒、偏離你命令的驕傲人， 你已經責備他們。
PS|119|22|求你除掉我所受的羞辱和藐視， 因我遵守你的法度。
PS|119|23|雖有掌權者坐著妄論我， 你僕人卻思想你的律例。
PS|119|24|你的法度也是我的喜樂， 我的導師 。
PS|119|25|我的性命幾乎歸於塵土， 求你照你的話將我救活！
PS|119|26|我述說我所做的，你應允了我； 求你將你的律例教導我！
PS|119|27|求你使我明白你的訓詞， 我要默想你的奇事。
PS|119|28|我因愁苦身心耗盡， 求你照你的話使我堅立！
PS|119|29|求你使我離開奸詐的道路， 開恩將你的律法賜給我！
PS|119|30|我選擇了忠信的道路， 將你的典章擺在我面前。
PS|119|31|我持守你的法度； 耶和華啊，求你不要叫我羞愧！
PS|119|32|你使我心胸開闊的時候， 我就往你命令的道路直奔。
PS|119|33|耶和華啊，求你將你的律例指教我， 我必遵守到底！
PS|119|34|求你賜我悟性，我就遵守你的律法， 且要一心遵守。
PS|119|35|求你叫我遵行你的命令， 因為這是我所喜愛的。
PS|119|36|求你使我的心趨向你的法度， 不趨向不義之財。
PS|119|37|求你叫我轉眼不看虛假， 使我活在你的道路 中。
PS|119|38|求你向敬畏你的僕人 堅守你的話！
PS|119|39|求你使我所懼怕的羞辱遠離我， 因你的典章本為美。
PS|119|40|看哪，我切慕你的訓詞， 求你因你的公義賜我生命 ！
PS|119|41|耶和華啊，求你使你的慈愛臨到我， 照你的話使你的救恩臨到我，
PS|119|42|我就有話回答那羞辱我的， 因我倚靠你的話。
PS|119|43|求你叫真理的話總不離開我的口， 因我仰望你的典章。
PS|119|44|我要常守你的律法， 直到永永遠遠。
PS|119|45|我要自由而行 ， 因我尋求了你的訓詞。
PS|119|46|我要在列王面前宣講你的法度， 也不致羞愧。
PS|119|47|我以你的命令為樂， 這命令是我所喜愛的。
PS|119|48|我向我所愛的，就是你的命令高舉雙手 ， 我也要默想你的律例。
PS|119|49|求你記念你向僕人所說的話， 這話使我有盼望。
PS|119|50|你的話將我救活了； 這是我在患難中的安慰。
PS|119|51|驕傲的人極度地侮慢我， 我卻未曾偏離你的律法。
PS|119|52|耶和華啊，我記念你從古以來的典章， 就得了安慰。
PS|119|53|我因惡人離棄你的律法， 怒火中燒。
PS|119|54|我在世寄居， 以你的律例為詩歌。
PS|119|55|耶和華啊，我夜間記念你的名， 我也要遵守你的律法。
PS|119|56|這臨到我， 是因我謹守你的訓詞。
PS|119|57|耶和華是我的福分； 我曾說，我要遵守你的話。
PS|119|58|我一心懇求你的面， 求你照你的話憐憫我！
PS|119|59|我思想自己所行的道路， 我的腳步就轉向你的法度。
PS|119|60|我速速遵守你的命令， 並不遲延。
PS|119|61|惡人的繩索纏繞我， 我卻沒有忘記你的律法。
PS|119|62|我因你公義的典章， 夜半起來稱謝你。
PS|119|63|凡敬畏你、守你訓詞的人， 我都與他作伴。
PS|119|64|耶和華啊，遍地滿了你的慈愛； 求你將你的律例教導我！
PS|119|65|耶和華啊，你照你的話， 善待你的僕人。
PS|119|66|求你教我明辨和知識， 因我信靠你的命令。
PS|119|67|我未受苦以先曾經迷失， 現在卻遵守你的話。
PS|119|68|你本為善，所行的也善； 求你將你的律例教導我！
PS|119|69|驕傲的人編造謊言攻擊我， 我卻要一心遵守你的訓詞。
PS|119|70|他們的心蒙昧如蒙油脂， 我卻喜愛你的律法。
PS|119|71|我受苦是與我有益， 為要使我學習你的律例。
PS|119|72|你口中的律法與我有益， 勝於千萬金銀。
PS|119|73|你的手造了我，塑造我； 求你賜我悟性學習你的命令！
PS|119|74|敬畏你的人看見我就歡喜， 因我仰望你的話。
PS|119|75|耶和華啊，我知道你的典章是公義的； 你使我受苦是以信實待我。
PS|119|76|求你照著你向僕人所說的話， 以慈愛安慰我。
PS|119|77|求你的憐憫臨到我，使我存活， 因你的律法是我的喜樂。
PS|119|78|願驕傲的人蒙羞，因為他們無理傾覆我； 但我要默想你的訓詞。
PS|119|79|願敬畏你的人和知道你法度的人 都歸向我。
PS|119|80|願我的心在你的律例上完全， 使我不致蒙羞。
PS|119|81|我渴想你的救恩身心耗盡， 我仰望你的話。
PS|119|82|我因渴望你的話眼睛失明，說： 「你何時安慰我呢？」
PS|119|83|我雖像煙薰的皮囊， 卻不忘記你的律例。
PS|119|84|你僕人的年日有多少呢？ 你幾時向迫害我的人施行審判呢？
PS|119|85|不順從你律法的驕傲人 為我掘了坑。
PS|119|86|你的命令盡都信實； 他們無理迫害我，求你幫助我！
PS|119|87|他們幾乎把我從世上除滅； 但我沒有離棄你的訓詞。
PS|119|88|求你照你的慈愛將我救活， 我就遵守你口中的法度。
PS|119|89|耶和華啊，你的話安定在天， 直到永遠。
PS|119|90|你的信實存到萬代； 你堅立了地，地就長存。
PS|119|91|天地照你的典章存到今日； 萬物都是你的僕役。
PS|119|92|我若不以你的律法為樂， 早就在苦難中滅絕了！
PS|119|93|我永不忘記你的訓詞， 因你用這訓詞將我救活。
PS|119|94|我是屬你的，求你救我， 因我尋求了你的訓詞。
PS|119|95|惡人等著要滅絕我， 我卻要揣摩你的法度。
PS|119|96|我看萬事盡都有限， 惟有你的命令極其寬廣。
PS|119|97|我何等愛慕你的律法， 終日不住地思想。
PS|119|98|你的命令常存在我心裏， 使我比仇敵有智慧。
PS|119|99|我比我的教師更通達， 因我思想你的法度。
PS|119|100|我比年老的更明白， 因我謹守你的訓詞。
PS|119|101|我阻止我的腳走一切邪路， 為要遵守你的話。
PS|119|102|我沒有偏離你的典章， 因為你教導了我。
PS|119|103|你的言語在我上膛何等甘美， 在我口中比蜜更甜！
PS|119|104|我藉著你的訓詞得以明白， 因此，我恨惡一切虛假的行徑。
PS|119|105|你的話是我腳前的燈， 是我路上的光。
PS|119|106|你公義的典章，我曾起誓遵守， 我必按著誓言而行。
PS|119|107|我極其痛苦； 耶和華啊，求你照你的話將我救活！
PS|119|108|耶和華啊，求你悅納我口中的讚美為甘心祭， 又將你的典章教導我！
PS|119|109|我的性命常在我手掌中 ， 我卻不忘記你的律法。
PS|119|110|惡人為我設下羅網， 我卻沒有偏離你的訓詞。
PS|119|111|我以你的法度為永遠的產業， 因這是我心中所喜愛的。
PS|119|112|我的心傾向你的律例， 謹守到底，直到永遠。
PS|119|113|心懷二意的人為我所恨； 但你的律法為我所愛。
PS|119|114|你是我藏身之處，是我的盾牌； 我仰望你的話。
PS|119|115|作惡的人哪，你們離開我吧！ 我要遵守我上帝的命令。
PS|119|116|求你照你的話扶持我，使我存活， 不要叫我因失望而蒙羞。
PS|119|117|求你扶持我，使我得救， 時常看重你的律例。
PS|119|118|凡偏離你律例的人，你都輕看他們， 因為他們的詭詐必歸虛空。
PS|119|119|你除掉地上所有的惡人，好像除掉渣滓 ； 因此我喜愛你的法度。
PS|119|120|我因懼怕你，肉體戰慄； 我害怕你的典章。
PS|119|121|我行公平和公義， 求你不要撇下我，交給欺壓我的人！
PS|119|122|求你保證你的僕人得福， 不容驕傲的人欺壓我！
PS|119|123|我因盼望你的救恩 和你公義的言語眼睛失明。
PS|119|124|求你照你的慈愛待僕人， 將你的律例教導我。
PS|119|125|我是你的僕人，求你賜我悟性， 得以認識你的法度。
PS|119|126|這是耶和華採取行動的時候， 因人廢棄了你的律法。
PS|119|127|所以，我喜愛你的命令勝於金子， 更勝於純金。
PS|119|128|你的一切訓詞，在萬事上我都以為正直； 我恨惡一切虛假的行徑。
PS|119|129|你的法度奇妙， 所以我一心謹守。
PS|119|130|你的話一開啟就發出亮光， 使愚蒙人通達。
PS|119|131|我大大張口，呼吸急促， 因我切慕你的命令。
PS|119|132|求你轉向我，憐憫我， 就像你待那些喜愛你名的人。
PS|119|133|求你用你的言語使我腳步穩健， 不容罪孽轄制我。
PS|119|134|求你救我脫離人的欺壓， 我要遵守你的訓詞。
PS|119|135|求你使你的臉向僕人發光， 又將你的律例教導我。
PS|119|136|我的眼睛流淚成河， 因為他們不守你的律法。
PS|119|137|耶和華啊，你是公義的； 你的典章正直！
PS|119|138|你所頒佈的法度是公義的， 極其可靠。
PS|119|139|我的狂熱把我燒滅， 因我敵人忘記你的話。
PS|119|140|你的言語極其精煉， 令你僕人喜愛。
PS|119|141|我渺小，被人藐視， 卻不忘記你的訓詞。
PS|119|142|你的公義永遠公義， 你的律法是確實的。
PS|119|143|我遭遇患難愁苦， 你的命令是我的喜樂。
PS|119|144|你的法度永遠公義； 求你賜我悟性，使我存活。
PS|119|145|耶和華啊，我一心呼求你，求你應允我！ 我必謹守你的律例。
PS|119|146|我向你呼求，求你救我！ 我要遵守你的法度。
PS|119|147|天尚未亮我呼喊求救， 我仰望你的話。
PS|119|148|我終夜雙眼睜開， 為要思想你的言語。
PS|119|149|求你按你的慈愛聽我的聲音， 耶和華啊，求你照你的典章將我救活！
PS|119|150|追逐奸惡的人 迫近了， 他們遠離你的律法。
PS|119|151|耶和華啊，你就在我身邊， 你一切的命令是確實的！
PS|119|152|我從你的法度早已知道， 這法度是你永遠立定的。
PS|119|153|求你看顧我的苦難，搭救我， 因我不忘記你的律法。
PS|119|154|求你為我的冤屈辯護，救贖我， 照你的言語將我救活。
PS|119|155|救恩遠離惡人， 因為他們不尋求你的律例。
PS|119|156|耶和華啊，你的憐憫本為大； 求你照你的典章將我救活。
PS|119|157|迫害我的、抵擋我的甚多， 我卻沒有偏離你的法度。
PS|119|158|我看見奸惡的人就憎惡， 因為他們不遵守你的言語。
PS|119|159|你看我何等喜愛你的訓詞！ 耶和華啊，求你按你的慈愛將我救活！
PS|119|160|你話語的精髓是真實的， 你一切公義的典章永遠長存。
PS|119|161|掌權者無故迫害我， 然而我的心畏懼你的話。
PS|119|162|我喜愛你的言語， 好像人得到許多戰利品。
PS|119|163|我恨惡，憎惡虛假； 惟喜愛你的律法。
PS|119|164|我因你公義的典章 一天七次讚美你。
PS|119|165|喜愛你律法的人大有平安， 任何事都不能使他們跌倒。
PS|119|166|耶和華啊，我仰望你的救恩， 遵行你的命令。
PS|119|167|我心謹守你的法度， 這法度我極其喜愛。
PS|119|168|我遵守你的訓詞和法度， 因我所行的道路都在你的面前。
PS|119|169|耶和華啊，願我的呼求達到你面前， 求你照你的話賜我悟性。
PS|119|170|願我的懇求達到你面前， 求你照你的言語搭救我。
PS|119|171|願我的嘴唇發出讚美， 因為你將律例教導我。
PS|119|172|願我的舌頭歌唱你的言語， 因你一切的命令盡都公義。
PS|119|173|求你用你的手幫助我， 因我選擇你的訓詞。
PS|119|174|耶和華啊，我切慕你的救恩！ 你的律法是我的喜樂。
PS|119|175|願我的性命存活，得以讚美你！ 願你的典章幫助我！
PS|119|176|我走迷了路如同失喪的羊，求你尋找你的僕人， 因我不忘記你的命令。
PS|120|1|我在急難中求告耶和華， 他就應允我。
PS|120|2|耶和華啊，求你救我脫離 說謊的嘴唇和詭詐的舌頭！
PS|120|3|詭詐的舌頭啊，他會給你甚麼呢？ 會加給你甚麼呢？
PS|120|4|就是勇士的利箭、 羅騰木 的炭火。
PS|120|5|禍哉！我寄居在 米設 ， 住在 基達 帳棚之中。
PS|120|6|我與那恨惡和平的人 許久同住。
PS|120|7|我願和平， 當我發言，他們卻要戰爭。
PS|121|1|我要向山舉目， 我的幫助從何而來？
PS|121|2|我的幫助 從造天地的耶和華而來。
PS|121|3|他不叫你的腳搖動， 保護你的必不打盹！
PS|121|4|保護 以色列 的 必不打盹，也不睡覺。
PS|121|5|保護你的是耶和華， 耶和華在你右邊蔭庇你。
PS|121|6|白日，太陽必不傷你； 夜間，月亮也不害你。
PS|121|7|耶和華要保護你，免受一切的災害， 他要保護你的性命。
PS|121|8|你出你入，耶和華要保護你， 從今時直到永遠。
PS|122|1|我喜樂， 因人對我說：「我們到耶和華的殿去。」
PS|122|2|耶路撒冷 啊， 我們的腳站在你門內。
PS|122|3|耶路撒冷 被建造， 如同連結整齊的一座城。
PS|122|4|眾支派就是耶和華的支派，上那裏去， 按 以色列 的法度頌揚耶和華的名。
PS|122|5|他們在那裏設立審判的寶座， 就是 大衛 家的寶座。
PS|122|6|你們要為 耶路撒冷 求平安： 「願愛你的人興旺！
PS|122|7|願你城中有平安！ 願你宮內得平靜！」
PS|122|8|為我弟兄和同伴的緣故，我要說： 「願你平安！」
PS|122|9|為耶和華－我們上帝殿的緣故， 我要為你求福！
PS|123|1|坐在天上的主啊， 我向你舉目。
PS|123|2|看哪，僕人的眼睛怎樣仰望主人的手， 婢女的眼睛怎樣仰望女主人的手， 我們的眼睛也照樣仰望耶和華－我們的上帝， 直到他憐憫我們。
PS|123|3|耶和華啊，求你憐憫我們，憐憫我們！ 因為我們受盡了藐視。
PS|123|4|我們受盡了安逸人的譏誚 和驕傲人的藐視。
PS|124|1|說吧， 以色列 ： 「若不是耶和華幫助我們，
PS|124|2|若不是耶和華幫助我們， 當人起來攻擊我們，
PS|124|3|那時，人向我們發怒， 就把我們活活吞了；
PS|124|4|那時，波濤必漫過我們， 河水必淹沒我們；
PS|124|5|那時，狂傲的水 必淹沒我們。」
PS|124|6|耶和華是應當稱頌的！ 他沒有把我們交給他們，作牙齒的獵物。
PS|124|7|我們好像雀鳥，從捕鳥人的羅網裏逃脫， 羅網破裂，我們就逃脫了。
PS|124|8|我們得幫助， 是因造天地之耶和華的名。
PS|125|1|倚靠耶和華的人好像 錫安山 ， 安穩坐鎮，永不動搖。
PS|125|2|眾山怎樣圍繞 耶路撒冷 ， 耶和華也照樣圍繞他的百姓，從今時直到永遠。
PS|125|3|惡人的杖必不在義人的土地上停留， 免得義人伸手作惡。
PS|125|4|耶和華啊，求你善待 行善和心裏正直的人。
PS|125|5|至於那偏行彎曲道路的人， 耶和華必將他們和作惡的人一同驅逐出去。 願平安歸於 以色列 ！
PS|126|1|當耶和華使 錫安 被擄的人歸回的時候， 我們好像做夢的人。
PS|126|2|那時，我們滿口喜笑、 滿舌歡呼； 那時，列國中就有人說： 「耶和華為他們行了大事！」
PS|126|3|耶和華果然為我們行了大事， 我們就歡喜。
PS|126|4|耶和華啊，求你使我們這些被擄的人歸回， 好像 尼革夫 的河水復流。
PS|126|5|流淚撒種的， 必歡呼收割！
PS|126|6|那帶種流淚出去的， 必歡呼地帶禾捆回來！
PS|127|1|若不是耶和華建造房屋， 建造的人就枉然勞力； 若不是耶和華看守城池， 看守的人就枉然警醒。
PS|127|2|你們清晨早起，夜晚安歇， 吃勞碌得來的飯，本是枉然； 惟有耶和華所親愛的， 必叫他安然睡覺。
PS|127|3|看哪，兒女是耶和華所賜的產業， 所懷的胎是他所給的賞賜。
PS|127|4|人在年輕時生的兒女 好像勇士手中的箭。
PS|127|5|箭袋充滿的人有福了！ 他們在城門口和仇敵爭論時必不蒙羞。
PS|128|1|凡敬畏耶和華、 遵行他道的人有福了！
PS|128|2|你要吃勞碌得來的； 你要享福，凡事順利。
PS|128|3|你妻子在你內室，好像多結果子的葡萄樹； 你兒女圍繞你的桌子，如同橄欖樹苗。
PS|128|4|看哪，敬畏耶和華的人 必要這樣蒙福！
PS|128|5|願耶和華從 錫安 賜福給你！ 願你一生一世看見 耶路撒冷 興旺！
PS|128|6|願你看見 你的子子孫孫！ 願平安歸於 以色列 ！
PS|129|1|說吧， 以色列 ： 「從我幼年以來，人屢次苦害我；
PS|129|2|從我幼年以來，人屢次苦害我， 卻沒有勝過我。
PS|129|3|扶犁的人在我背上扶犁而耕， 耕的犁溝很長。」
PS|129|4|耶和華是公義的， 他砍斷了惡人的繩索。
PS|129|5|願恨惡 錫安 的 都蒙羞退後！
PS|129|6|願他們像房頂上的草， 一發芽就枯乾，
PS|129|7|收割的不夠用手抓一把， 捆禾的也不夠抱滿懷。
PS|129|8|過路的也不說：「願耶和華所賜的福歸與你們！ 我們奉耶和華的名給你們祝福！」
PS|130|1|耶和華啊， 我從深處求告你！
PS|130|2|主啊，求你聽我的聲音！ 求你側耳聽我懇求的聲音！
PS|130|3|耶和華啊，你若究察罪孽， 主啊，誰能站得住呢？
PS|130|4|但在你有赦免之恩， 要叫人敬畏你。
PS|130|5|我等候耶和華，我的心等候； 我也仰望他的話。
PS|130|6|我的心等候主，勝於守夜的等候天亮， 勝於守夜的等候天亮。
PS|130|7|以色列 啊，你當仰望耶和華， 因耶和華有慈愛，有豐盛的救恩。
PS|130|8|他必救贖 以色列 脫離一切的罪孽。
PS|131|1|耶和華啊，我的心不狂妄， 我的眼不高傲； 重大和測不透的事， 我也不敢行。
PS|131|2|我使我心安穩平靜，好像母親懷中斷奶的孩子； 我的心在我裏面如同斷過奶的孩子。
PS|131|3|以色列 啊，你當仰望耶和華， 從今時直到永遠！
PS|132|1|耶和華啊，求你記念 大衛 ， 記念他所受的一切苦難！
PS|132|2|他怎樣向耶和華起誓， 向 雅各 的大能者許願：
PS|132|3|「我必不進我的帳幕， 也不上我的床鋪；
PS|132|4|我不容我的眼睛睡覺， 也不容我的眼皮打盹；
PS|132|5|直等到我為耶和華尋得所在， 為 雅各 的大能者尋得居所。」
PS|132|6|我們聽說約櫃在 以法他 ， 我們在 雅珥 的田野尋見它。
PS|132|7|「我們要進他的居所， 在他腳凳前下拜。」
PS|132|8|耶和華啊，求你興起， 與你有能力的約櫃同入安歇之所！
PS|132|9|願你的祭司披上公義！ 願你的聖民歡呼！
PS|132|10|求你因你僕人 大衛 的緣故， 不要厭棄你的受膏者！
PS|132|11|耶和華憑信實向 大衛 起了誓，絕不改變： 「我要立你身所生的 坐在你的寶座上。
PS|132|12|你的眾子若謹守我的約和我所教導他們的法度， 他們的子孫必永遠坐在你的寶座上。」
PS|132|13|因為耶和華揀選了 錫安 ， 願意當作自己的居所：
PS|132|14|「這是我永遠安歇之所； 我要住在這地方，因為我願意在這裏。
PS|132|15|我要賜福使糧食豐足， 使其中的貧窮人飽享食物。
PS|132|16|我要使祭司披上救恩， 聖民就要大聲歡呼！
PS|132|17|在那裏我要使 大衛 的角茁壯， 為我的受膏者預備明燈。
PS|132|18|我要使他的仇敵披上羞恥； 但他的冠冕要在他頭上發光。」
PS|133|1|看哪，弟兄和睦同住 是何等的善，何等的美！
PS|133|2|這好比那貴重的油澆在 亞倫 的頭上， 流到鬍鬚，又流到他的衣襟；
PS|133|3|又好比 黑門 的甘露降在 錫安山 ； 因為在那裏有耶和華所命定的福，就是永遠的生命。
PS|134|1|來，稱頌耶和華！ 夜間侍立在耶和華殿中，耶和華的僕人，
PS|134|2|當向聖所舉手， 稱頌耶和華！
PS|134|3|願造天地的耶和華 從 錫安 賜福給你們！
PS|135|1|哈利路亞！ 你們要讚美耶和華的名！ 侍立在耶和華殿中，耶和華的僕人， 侍立在我們上帝殿院中的，要讚美他！
PS|135|2|
PS|135|3|你們要讚美耶和華， 因耶和華本為善； 要歌頌他的名， 因為這是美好的。
PS|135|4|耶和華揀選 雅各 歸自己， 揀選 以色列 作他寶貴的產業。
PS|135|5|我知道耶和華本為大， 也知道我們的主超乎萬神之上。
PS|135|6|在天，在地，在海洋，在各深淵， 耶和華都隨自己的旨意而行。
PS|135|7|他使雲霧從地極上騰， 造電隨雨而閃， 從倉庫中吹出風來。
PS|135|8|他將 埃及 頭生的， 連人帶牲畜都擊殺了。
PS|135|9|埃及 啊，他施行神蹟奇事， 在你們中間，在法老和他所有臣僕身上。
PS|135|10|他擊打許多國家， 殺戮大能的君王，
PS|135|11|就是 亞摩利 王 西宏 、 巴珊 王 噩 ， 和 迦南 一切的國度，
PS|135|12|他賞賜他們的地為業， 作為自己百姓 以色列 的產業。
PS|135|13|耶和華啊，你的名字存到永遠！ 耶和華啊，你的稱號 存到萬代！
PS|135|14|耶和華要為自己的百姓伸冤， 為自己的僕人發憐憫。
PS|135|15|外邦的偶像是金的，是銀的， 是人手所造的，
PS|135|16|有口卻不能言， 有眼卻不能看，
PS|135|17|有耳卻不能聽， 口中也沒有氣息。
PS|135|18|造它們的要像它們一樣， 凡靠它們的也必如此。
PS|135|19|以色列 家啊，要稱頌耶和華！ 亞倫 家啊，要稱頌耶和華！
PS|135|20|利未 家啊，要稱頌耶和華！ 你們敬畏耶和華的，要稱頌耶和華！
PS|135|21|住在 耶路撒冷 的、 錫安 的耶和華， 是應當稱頌的。 哈利路亞！
PS|136|1|你們要稱謝耶和華，因他本為善； 他的慈愛永遠長存。
PS|136|2|你們要稱謝萬神之神， 因他的慈愛永遠長存。
PS|136|3|你們要稱謝萬主之主， 因他的慈愛永遠長存。
PS|136|4|稱謝那惟一能行大 奇事的， 因他的慈愛永遠長存。
PS|136|5|稱謝那用智慧造天的， 因他的慈愛永遠長存。
PS|136|6|稱謝那鋪地在水以上的， 因他的慈愛永遠長存。
PS|136|7|稱謝那造成大光的， 因他的慈愛永遠長存。
PS|136|8|他造太陽管白晝， 因他的慈愛永遠長存。
PS|136|9|他造月亮星宿管黑夜， 因他的慈愛永遠長存。
PS|136|10|稱謝那擊殺 埃及 凡是頭生的， 因他的慈愛永遠長存。
PS|136|11|他以大能的手和伸出來的膀臂， 因他的慈愛永遠長存。 領 以色列 人從 埃及 人中出來， 因他的慈愛永遠長存。
PS|136|12|
PS|136|13|稱謝那分裂 紅海 的， 因他的慈愛永遠長存。
PS|136|14|他領 以色列 從其中經過， 因他的慈愛永遠長存；
PS|136|15|卻把法老和他的軍隊推落 紅海 裏， 因他的慈愛永遠長存。
PS|136|16|稱謝那引導自己子民行走曠野的， 因他的慈愛永遠長存。
PS|136|17|稱謝那擊殺大君王的， 因他的慈愛永遠長存。
PS|136|18|他殺戮威武的君王， 因他的慈愛永遠長存；
PS|136|19|殺戮 亞摩利 王 西宏 ， 因他的慈愛永遠長存；
PS|136|20|殺戮 巴珊 王 噩 ， 因他的慈愛永遠長存。
PS|136|21|他賞賜他們的地為業， 因他的慈愛永遠長存；
PS|136|22|作為他僕人 以色列 的產業， 因他的慈愛永遠長存。
PS|136|23|我們身處卑微，他顧念我們， 因他的慈愛永遠長存。
PS|136|24|他搭救我們脫離敵人， 因他的慈愛永遠長存。
PS|136|25|凡有血有肉的，他賜糧食， 因他的慈愛永遠長存。
PS|136|26|你們要稱謝天上的上帝， 因他的慈愛永遠長存。
PS|137|1|我們在 巴比倫 河邊， 坐在那裏，追想 錫安 ，就哭了。
PS|137|2|在一排柳樹中， 我們掛上我們的豎琴。
PS|137|3|擄掠我們的在那裏 要我們唱歌； 搶奪我們的要我們為他們作樂： 「給我們唱一首 錫安 的歌吧！」
PS|137|4|我們怎能在外邦之土 唱耶和華的歌呢？
PS|137|5|耶路撒冷 啊，我若忘記你， 寧願我的右手枯萎；
PS|137|6|我若不記得你，不看你過於我最喜樂的， 寧願我的舌頭貼於上膛！
PS|137|7|耶路撒冷 攻破的日子， 以東 人說：「拆毀！拆毀！ 直拆到根基！」 耶和華啊，求你記得！
PS|137|8|將要被滅的 巴比倫 哪， 用你待我們的惡行報復你的，那人有福了。
PS|137|9|抓起你的嬰孩摔在磐石上的， 那人有福了。
PS|138|1|我要一心稱謝你 ， 在諸神面前歌頌你。
PS|138|2|我要向你的聖殿下拜， 我要因你的慈愛和信實頌揚你的名； 因你使你的名和你的言語顯為大， 超乎一切 。
PS|138|3|我呼求的日子，你應允我， 使我壯膽，心裏有能力。
PS|138|4|耶和華啊，地上的君王都要稱謝你， 因他們聽見了你口中的言語。
PS|138|5|他們要歌頌耶和華的作為， 因耶和華大有榮耀。
PS|138|6|耶和華雖崇高，卻看顧卑微的人； 驕傲的人，他從遠處即能認出。
PS|138|7|我雖困在患難中，你必將我救活； 我的仇敵發怒，你必伸手抵擋他們， 你的右手也必拯救我。
PS|138|8|耶和華必成全他在我身上的旨意； 耶和華啊，你的慈愛永遠長存！ 求你不要離棄你手所造的。
PS|139|1|耶和華啊，你已經鑒察我， 認識我。
PS|139|2|我坐下，我起來，你都曉得； 你從遠處知道我的意念。
PS|139|3|我行路，我躺臥，你都細察； 你也深知我一切所行的。
PS|139|4|耶和華啊，我舌頭上的話， 你沒有一句不知道的。
PS|139|5|你前後環繞我， 按手在我身上。
PS|139|6|這樣的知識奇妙，是我不能測的； 至高，是我不能及的。
PS|139|7|我往哪裏去，躲避你的靈？ 我往哪裏逃，躲避你的面？
PS|139|8|我若升到天上，你在那裏； 我若躺在陰間，你也在那裏。
PS|139|9|我若展開清晨的翅膀， 飛到海極居住，
PS|139|10|就是在那裏，你的手必引導我， 你的右手也必扶持我。
PS|139|11|我若說「黑暗必定壓碎我， 我周圍的亮光必成為黑夜」，
PS|139|12|黑暗對你不再是黑暗， 黑夜卻如白晝發亮。 黑暗和光明， 在你看來都是一樣。
PS|139|13|我的肺腑是你所造的， 我在母腹中，你已編織 我。
PS|139|14|我要稱謝你，因我受造奇妙可畏， 你的作為奇妙，這是我心深知道的。
PS|139|15|我在暗中受造，在地的深處被塑造； 那時，我的形體並不向你隱藏。
PS|139|16|我未成形的體質， 你的眼早已看見了； 你所定的日子，我尚未度一日， 都在你的冊子寫上了。
PS|139|17|上帝啊，你的意念向我何等寶貴！ 其數何等眾多！
PS|139|18|我若數點，比海沙更多； 我睡醒的時候，仍和你同在。
PS|139|19|上帝啊，惟願你殺戮惡人； 你們好流人血的，離開我去吧！
PS|139|20|他們說惡言頂撞你， 你的仇敵妄稱你的名 。
PS|139|21|耶和華啊，恨惡你的，我豈不恨惡他們嗎？ 攻擊你的，我豈不憎惡他們嗎？
PS|139|22|我恨惡他們到極點， 以他們為我的仇敵。
PS|139|23|上帝啊，求你鑒察我，知道我的心思， 試煉我，知道我的意念；
PS|139|24|看在我裏面有甚麼惡行沒有， 引導我走永生的道路。
PS|140|1|耶和華啊，求你救我脫離邪惡的人， 保護我脫離殘暴的人！
PS|140|2|他們心中圖謀奸惡， 日日不停挑起戰爭。
PS|140|3|他們的舌頭銳利如蛇， 嘴唇裏有毒蛇的毒液。（細拉）
PS|140|4|耶和華啊，求你庇護我脫離惡人的手， 保護我脫離殘暴的人，他們想要推倒我。
PS|140|5|驕傲的人為我暗設羅網和繩索； 他們在路旁張開網，為我設下圈套。（細拉）
PS|140|6|我曾對耶和華說：「你是我的上帝。」 耶和華啊，求你側耳聽我懇求的聲音！
PS|140|7|主－耶和華、我救恩的力量啊， 在戰爭的日子，你遮蔽了我的頭。
PS|140|8|耶和華啊，求你不要遂惡人的心願； 不要成就他們的計謀，免得他們自高。（細拉）
PS|140|9|至於那些昂首圍困我的人， 願他們嘴唇的奸惡陷害 自己！
PS|140|10|願他們被丟在火中，火炭落在他們身上； 願他們被拋在深坑裏，不能再起來！
PS|140|11|願說惡言的人在地上站立不住； 願禍患獵取殘暴的人，把他打倒。
PS|140|12|我知道耶和華必為困苦人伸冤， 為貧窮人辯護。
PS|140|13|義人必頌揚你的名， 正直人要在你面前居住。
PS|141|1|耶和華啊，我曾求告你， 求你快快臨到我這裏！ 我求告你的時候， 求你側耳聽我的聲音！
PS|141|2|願我的禱告如香呈到你面前！ 願我的手舉起 ，如獻晚祭！
PS|141|3|耶和華啊，求你看守我的口， 把守我的嘴唇！
PS|141|4|不要使我的心偏向邪惡的事， 以致我和作惡的人一同行惡； 也不叫我吃他們的美食。
PS|141|5|任憑義人擊打我，這算為仁慈； 任憑他責備我，這算為頭上的膏油； 我的頭不躲閃。 人正行惡的時候，我仍要祈禱。
PS|141|6|他們的審判官被扔在巖下， 他們就要聽我的話，因為這話甘甜。
PS|141|7|我們的 骨頭散落在陰間的口， 就像人耕田刨地 一樣。
PS|141|8|主－耶和華啊，我的眼目仰望你； 我投靠你，求你不要使我的性命陷入危險！
PS|141|9|求你保護我脫離惡人為我設的羅網 和作惡之人的圈套！
PS|141|10|願惡人落在自己的網中， 我卻得以逃脫。
PS|142|1|我出聲哀告耶和華， 出聲懇求耶和華。
PS|142|2|我在他面前傾訴我的苦情， 在他面前陳說我的患難。
PS|142|3|我的靈在我裏面發昏的時候， 你知道我的道路。 在我所行的路上， 人為我暗設羅網。
PS|142|4|求你留意向我右邊觀看， 無人認識我； 我無避難之處， 也無人眷顧我。
PS|142|5|耶和華啊，我曾向你哀求。 我說：「你是我的避難所， 在活人之地，你是我的福分。」
PS|142|6|求你留心聽我的呼求， 因我落到極卑微之地； 求你救我脫離迫害我的人， 因為他們比我強盛。
PS|142|7|求你從被囚之地領我出來， 我好頌揚你的名。 義人必環繞我， 因為你用厚恩待我。
PS|143|1|耶和華啊，求你聽我的禱告， 側耳聽我的懇求，憑你的信實和公義應允我。
PS|143|2|求你不要審問僕人， 因為在你面前，凡活著的人沒有一個是義的。
PS|143|3|因為仇敵迫害我， 將我打倒在地， 使我住在幽暗之處， 像死了許久的人一樣。
PS|143|4|我的靈在我裏面發昏， 我的心在我裏面顫慄。
PS|143|5|我追想古時之日，思想你的一切作為， 默念你手的工作。
PS|143|6|我向你舉手， 我的心渴想你，如乾旱之地盼雨一樣。（細拉）
PS|143|7|耶和華啊，求你速速應允我！ 我的心神耗盡！ 求你不要轉臉不顧我， 免得我像那些下入地府的人一樣。
PS|143|8|求你使我清晨得聽你慈愛的聲音， 因我倚靠你； 求你使我知道當走的路， 因我的心仰望你。
PS|143|9|耶和華啊，求你救我脫離我的仇敵！ 我往你那裏藏身。
PS|143|10|求你指教我遵行你的旨意， 因你是我的上帝； 願你至善的靈 引我到平坦之地。
PS|143|11|耶和華啊，求你為你名的緣故將我救活， 憑你的公義，將我從患難中領出來，
PS|143|12|憑你的慈愛剪除我的仇敵， 滅絕所有苦待我的人，因我是你的僕人。
PS|144|1|耶和華─我的磐石是應當稱頌的！ 他教導我的手爭戰， 教導我的指頭打仗。
PS|144|2|他是我慈愛的主、我的山寨、 我的碉堡、我的救主、 我的盾牌，是我所投靠的。 他使我的百姓 服在我以下。
PS|144|3|耶和華啊，人算甚麼，你竟認識他！ 世人算甚麼，你竟顧念他！
PS|144|4|人不過像一口氣， 他的年日如影消逝。
PS|144|5|耶和華啊，求你使天下垂，親自降臨； 求你摸山，使山冒煙。
PS|144|6|求你發出閃電，使仇敵四散， 射出你的箭，使他們混亂。
PS|144|7|求你從高處伸手救拔我， 救我脫離大水，脫離外邦人的手。
PS|144|8|他們的口說謊話， 他們的右手起假誓。
PS|144|9|上帝啊，我要向你唱新歌， 用十弦瑟向你歌頌。
PS|144|10|你是那拯救君王的， 你是那救僕人 大衛 脫離害命之刀的。
PS|144|11|求你救拔我， 救我脫離外邦人的手。 他們的口說謊話， 他們的右手起假誓。
PS|144|12|我們的兒子從幼年好像樹苗長大， 我們的女兒如同房角石，按照建宮殿的樣式鑿成。
PS|144|13|我們的倉盈滿，能供應各種糧食； 我們的羊在田野孳生千萬。
PS|144|14|我們的牲口馱滿貨物， 沒有人闖進來搶奪， 也沒有人出去爭戰； 我們的街市上也沒有哭號的聲音。
PS|144|15|這樣情況的百姓有福了！ 以耶和華為他們上帝的百姓有福了！
PS|145|1|我的上帝、我的王啊、我要尊崇你！ 我要永永遠遠稱頌你的名！
PS|145|2|我要天天稱頌你， 也要永永遠遠讚美你的名！
PS|145|3|耶和華本為大，該受大讚美， 其大無法測度。
PS|145|4|這一代要對那一代頌讚你的作為， 他們要傳揚你的大能。
PS|145|5|他們要述說你威嚴榮耀的尊榮， 我要默念你奇妙的作為 。
PS|145|6|人要傳講你可畏的能力， 我也要傳揚你的偉大。
PS|145|7|他們要將你可記念的大恩傳開， 並要高唱你的公義。
PS|145|8|耶和華有恩惠，有憐憫， 不輕易發怒，大有慈愛。
PS|145|9|耶和華善待萬有， 他的憐憫覆庇他一切所造的。
PS|145|10|耶和華啊，你一切所造的都要稱謝你， 你的聖民也要稱頌你。
PS|145|11|他們要傳講你國度的榮耀， 談論你的大能，
PS|145|12|好讓世人知道你大能的作為 和你國度威嚴的榮耀。
PS|145|13|你的國是永遠的國！ 你執掌的權柄存到萬代！ 耶和華一切的話信實可靠， 他一切的作為都有慈愛 。
PS|145|14|耶和華扶起所有跌倒的， 扶起所有被壓下的。
PS|145|15|萬有的眼目都仰望你， 你按時給他們食物。
PS|145|16|你張手， 使一切有生命的都隨願飽足。
PS|145|17|耶和華一切所行的，無不公義， 一切所做的，都有慈愛。
PS|145|18|耶和華臨近凡求告他的， 臨近所有誠心求告他的人。
PS|145|19|敬畏他的，他必成就他們的心願， 也必聽他們的呼求，拯救他們。
PS|145|20|耶和華保護凡愛他的人， 卻要滅絕所有的惡人。
PS|145|21|我的口要述說讚美耶和華的話； 惟願有血肉之軀的都永永遠遠稱頌他的聖名。
PS|146|1|哈利路亞！ 我的心哪，你要讚美耶和華！
PS|146|2|我一生要讚美耶和華！ 我還活著的時候要歌頌我的上帝！
PS|146|3|你們不要倚靠君王，不要倚靠世人， 他一點也不能幫助。
PS|146|4|他的氣一斷，就歸回塵土， 他所打算的，當日就消滅了。
PS|146|5|以 雅各 的上帝為幫助、 仰望耶和華－他上帝的，這人有福了！
PS|146|6|耶和華造天、地、海和其中的萬物， 他守信實，直到永遠。
PS|146|7|他為受欺壓的伸冤， 賜食物給飢餓的人。 耶和華釋放被囚的，
PS|146|8|耶和華開了盲人的眼睛， 耶和華扶起被壓下的人， 耶和華喜愛義人。
PS|146|9|耶和華保護寄居的，扶持孤兒和寡婦， 卻使惡人的道路彎曲。
PS|146|10|耶和華要作王，直到永遠！ 錫安 哪，你的上帝要作王，直到萬代！ 哈利路亞！
PS|147|1|哈利路亞！ 歌頌我們的上帝是美善的， 因為他是美好的，讚美他是合宜的。
PS|147|2|耶和華建造 耶路撒冷 ， 聚集 以色列 中被趕散的人。
PS|147|3|他醫好傷心的人， 包紮他們的傷處。
PS|147|4|他數點星宿的數目， 一一稱它們的名。
PS|147|5|我們的主本為大，大有能力， 他的智慧無法測度。
PS|147|6|耶和華扶持謙卑的人， 將惡人傾覆於地。
PS|147|7|你們要以感謝向耶和華歌唱， 用琴向我們的上帝歌頌。
PS|147|8|他用密雲遮天，為地預備雨水， 使草生長在山上。
PS|147|9|他賜食物給走獸 和啼叫的小烏鴉。
PS|147|10|他不喜悅馬的力大， 不喜愛人的腿快。
PS|147|11|耶和華喜愛敬畏他 和盼望他慈愛的人。
PS|147|12|耶路撒冷 啊，要頌讚耶和華！ 錫安 哪，要讚美你的上帝！
PS|147|13|因為他堅固了你的門閂， 賜福給你中間的兒女。
PS|147|14|他使你境內平安， 用上好的麥子使你滿足。
PS|147|15|他向大地發出命令， 他的話速速頒行。
PS|147|16|他降雪如羊毛， 撒霜如灰燼。
PS|147|17|他擲下冰雹如碎渣， 他發出寒冷，誰能當得起呢？
PS|147|18|他一出令，這些就都融化， 他使風颳起，水便流動。
PS|147|19|他將他的道指示 雅各 ， 將他的律例典章指示 以色列 。
PS|147|20|他未曾這樣對待別國， 至於他的典章，他們向來都不知道 。 哈利路亞！
PS|148|1|哈利路亞！ 你們要從天上讚美耶和華， 在高處讚美他！
PS|148|2|他的眾使者啊，要讚美他！ 他的諸軍啊，都要讚美他！
PS|148|3|太陽月亮啊，要讚美他！ 放光的星宿啊，都要讚美他！
PS|148|4|天上的天和天上的水啊， 你們都要讚美他！
PS|148|5|願這些都讚美耶和華的名！ 因他一吩咐就都造成。
PS|148|6|他將這些設定，直到永永遠遠； 他訂了律例，不能廢去。
PS|148|7|你們哪，都當讚美耶和華： 地上一切所有的，大魚和深洋，
PS|148|8|火和冰雹，雪和霧氣， 成就他命令的狂風，
PS|148|9|大山和小山， 結果子的樹木和一切香柏樹，
PS|148|10|野獸和一切牲畜， 昆蟲和飛鳥，
PS|148|11|世上的君王和萬民， 領袖和世上所有的審判官，
PS|148|12|少年和少女， 老人和孩童，
PS|148|13|願這些都讚美耶和華的名！ 因為獨有他的名被尊崇，他的榮耀在天地之上。
PS|148|14|他高舉自己百姓的角， 使他的聖民 以色列 人，就是與他相近的百姓得榮耀 。 哈利路亞！
PS|149|1|哈利路亞！ 你們要向耶和華唱新歌， 在聖民的會中讚美他！
PS|149|2|願 以色列 因造他的主歡喜！ 願 錫安 的民因他們的王快樂！
PS|149|3|願他們跳舞讚美他的名， 擊鼓彈琴歌頌他！
PS|149|4|因為耶和華喜愛自己的百姓， 他要用救恩當作謙卑人的妝飾。
PS|149|5|願聖民因所得的榮耀歡樂！ 願他們在床上也歡呼！
PS|149|6|願他們口中稱頌上帝為至高， 手裏有兩刃的劍，
PS|149|7|為要報復列國， 懲罰萬民。
PS|149|8|要用鏈子捆他們的君王， 用鐵鐐鎖他們的貴族，
PS|149|9|要在他們身上施行所記錄的審判。 他的聖民都享榮耀。 哈利路亞！
PS|150|1|哈利路亞！ 你們要在上帝的聖所讚美他！ 在他顯能力的穹蒼讚美他！
PS|150|2|要因他大能的作為讚美他， 因他極其偉大讚美他！
PS|150|3|要用角聲讚美他， 鼓瑟彈琴讚美他！
PS|150|4|擊鼓跳舞讚美他！ 用絲弦的樂器和簫的聲音讚美他！
PS|150|5|用大響的鈸讚美他！ 用高聲的鈸讚美他！
PS|150|6|凡有生命的都要讚美耶和華！ 哈利路亞！
PROV|1|1|大衛 的兒子， 以色列 王 所羅門 的箴言：
PROV|1|2|要使人懂得智慧和訓誨， 明白通達的言語，
PROV|1|3|使人領受明智的訓誨， 就是公義、公平和正直，
PROV|1|4|使愚蒙人靈巧， 使年輕人有知識，有智謀。
PROV|1|5|智慧人聽見，增長學問， 聰明人得著智謀，
PROV|1|6|明白箴言和譬喻， 懂得智慧人的言詞和謎語。
PROV|1|7|敬畏耶和華是知識的開端； 愚妄人藐視智慧和訓誨。
PROV|1|8|我兒啊，要聽你父親的訓誨， 不可離棄你母親的教誨；
PROV|1|9|因為這要作你頭上恩惠的華冠， 作你頸上的項鏈。
PROV|1|10|我兒啊，罪人若引誘你， 你不可隨從。
PROV|1|11|他們若說：「你與我們同去， 我們要埋伏殺人流血， 無故地潛藏，殺害無辜；
PROV|1|12|我們好像陰間，把他們活活吞下， 囫圇吞下，如吞下那下到地府的人；
PROV|1|13|我們必得各樣寶物， 將所奪來的裝滿房屋；
PROV|1|14|你來與我們同夥， 共用一個錢囊。」
PROV|1|15|我兒啊，不要與他們走同一道路， 禁止你的腳走他們的路徑。
PROV|1|16|因為他們的腳奔跑行惡， 他們急速殺人流血。
PROV|1|17|在飛鳥眼前張設網羅， 一定會徒勞無功；
PROV|1|18|同樣，他們埋伏，是自流己血， 他們潛藏，是自害己命。
PROV|1|19|凡靠暴力歛財的，所行之路都是如此， 這種念頭必奪去自己的生命。
PROV|1|20|智慧 在街市上呼喊， 在廣場上高聲吶喊，
PROV|1|21|在熱鬧街頭呼叫， 在城門口，在城中，發出言語，說：
PROV|1|22|「你們無知的人喜愛無知， 傲慢人喜歡傲慢， 愚昧人恨惡知識， 要到幾時呢？
PROV|1|23|你們當因我的責備回轉， 我要將我的靈澆灌你們， 將我的話指示你們。
PROV|1|24|因為我呼喚，你們不聽， 我招手，無人理會。
PROV|1|25|你們忽視我一切的勸戒， 拒聽我的責備。
PROV|1|26|你們遭難，我就發笑； 驚恐臨到你們， 驚恐如狂風來臨， 災難好像暴風來到， 急難痛苦臨到你們身上， 我必嗤笑。
PROV|1|27|
PROV|1|28|那時，他們就會呼求我，我卻不回答， 懇切尋求我，卻尋不見。
PROV|1|29|因為他們恨惡知識， 選擇不敬畏耶和華，
PROV|1|30|不聽我的勸戒， 藐視我一切的責備，
PROV|1|31|所以他們要自食其果， 飽脹在自己的計謀中。
PROV|1|32|愚蒙人背道，害死自己， 愚昧人安逸，自取滅亡。
PROV|1|33|惟聽從我的，必安然居住， 得享寧靜，不怕災禍。」
PROV|2|1|我兒啊，你若領受我的言語， 珍藏我的命令，
PROV|2|2|留心聽智慧， 專心求聰明；
PROV|2|3|你若呼求明理， 揚聲求聰明，
PROV|2|4|尋找她，如尋找銀子， 搜尋她，如搜尋寶藏，
PROV|2|5|你就懂得敬畏耶和華， 得以認識上帝。
PROV|2|6|因為耶和華賞賜智慧， 知識和聰明都由他口而出。
PROV|2|7|他為正直人珍藏健全的知識， 給行為純正的人作盾牌，
PROV|2|8|為要保護公正的路， 庇護虔誠人的道。
PROV|2|9|那時，你就明白公義、公平、 正直，和一切完善的道路。
PROV|2|10|因為智慧要進入你的心， 知識要使你內心歡愉。
PROV|2|11|智謀要庇護你， 聰明必保護你，
PROV|2|12|救你脫離惡人的道， 脫離言談乖謬的人。
PROV|2|13|他們離棄正直的路， 行走黑暗的道，
PROV|2|14|喜歡作惡， 喜愛惡人的錯謬。
PROV|2|15|他們的路歪曲， 他們偏離中道。
PROV|2|16|智慧要救你遠離陌生女子， 遠離那油嘴滑舌的外邦女子。
PROV|2|17|她離棄年輕時的配偶， 忘了自己神聖的盟約。
PROV|2|18|她的家陷入死亡， 她的路偏向陰魂。
PROV|2|19|凡到她那裏去的，不得回轉， 也得不到生命的路。
PROV|2|20|智慧使你行善人的道， 守義人的路。
PROV|2|21|正直人必在地上居住， 完全人必在其上存留；
PROV|2|22|惟惡人要從地上剪除， 奸詐人要被拔出。
PROV|3|1|我兒啊，不要忘記我的教誨， 你的心要謹守我的命令，
PROV|3|2|因為它們 必加給你長久的日子， 生命的年數與平安。
PROV|3|3|不可使慈愛和誠信離開你， 要繫在你頸項上，刻在你心版上。
PROV|3|4|這樣，你必在上帝和世人眼前 蒙恩惠，有美好的見識。
PROV|3|5|你要專心仰賴耶和華， 不可倚靠自己的聰明，
PROV|3|6|在你一切所行的路上都要認定他， 他必使你的道路平直。
PROV|3|7|不要自以為有智慧； 要敬畏耶和華，遠離惡事。
PROV|3|8|這便醫治你的肉體 ， 滋潤你的百骨。
PROV|3|9|你要以財物 和一切初熟的土產尊崇耶和華，
PROV|3|10|這樣，你的倉庫必充滿有餘， 你的酒池有新酒盈溢。
PROV|3|11|我兒啊，不可輕看耶和華的管教， 也不可厭煩他的責備，
PROV|3|12|因為耶和華所愛的，他必責備， 正如父親責備所喜愛的兒子。
PROV|3|13|得智慧，得聰明的， 這人有福了。
PROV|3|14|因為智慧的獲利勝過銀子， 所得的盈餘強如金子，
PROV|3|15|比寶石 更寶貴， 你一切所喜愛的，都不足與其比較。
PROV|3|16|她的右手有長壽， 左手有富貴。
PROV|3|17|她的道是安樂， 她的路全是平安。
PROV|3|18|她給持守她的人作生命樹， 謹守她的必定蒙福。
PROV|3|19|耶和華以智慧奠立地基， 以聰明鋪設諸天，
PROV|3|20|以知識使深淵裂開， 使天空滴下甘露。
PROV|3|21|我兒啊，要謹守健全的知識和智謀， 不可使它們偏離你的眼目。
PROV|3|22|這樣，它們必使你的生命有活力， 又作你頸項的美飾。
PROV|3|23|那時，你就坦然行路， 不致跌倒。
PROV|3|24|你躺下，必不懼怕； 你躺臥，睡得香甜。
PROV|3|25|忽然來的驚恐，你不要害怕； 惡人遭毀滅，也不要恐懼，
PROV|3|26|因為耶和華是你的倚靠， 他必保護你的腳不陷入羅網。
PROV|3|27|你的手若有行善的力量， 不可推辭，要施與那應得的人。
PROV|3|28|你若手頭方便， 不可對鄰舍說： 「去吧，明天再來，我必給你。」
PROV|3|29|你的鄰舍既在你附近安居， 不可設計害他。
PROV|3|30|人若未曾加害你， 不可無故與他相爭。
PROV|3|31|不可嫉妒殘暴的人， 不可選擇他的任何道路。
PROV|3|32|因為走偏方向的人是耶和華所憎惡的； 正直人為他所親密。
PROV|3|33|耶和華詛咒惡人的家； 義人的居所他卻賜福。
PROV|3|34|他譏誚那愛譏誚的人； 但賜恩給謙卑的人。
PROV|3|35|智慧人必承受尊榮； 愚昧人高升卻是羞辱。
PROV|4|1|孩子們，要聽父親的訓誨， 留心明白道理。
PROV|4|2|因我給你們好的教導， 不可離棄我的教誨。
PROV|4|3|當我在父親面前還是小孩， 是母親獨一嬌兒的時候，
PROV|4|4|他教導我說：「你的心要持守我的話， 遵守我的命令，你就會存活。
PROV|4|5|要獲得智慧，要獲得聰明， 不可忘記， 也不可偏離我口中的言語。
PROV|4|6|不可離棄智慧，智慧就庇護你， 要愛她，她就保護你。
PROV|4|7|智慧為首，所以要獲得智慧， 要用你一切所有的換取聰明。
PROV|4|8|高舉智慧，她就使你升高， 擁抱智慧，她就使你尊榮。
PROV|4|9|她必將恩惠的華冠加在你頭上， 把榮冕賜給你。」
PROV|4|10|我兒啊，要聽，要領受我的言語， 你就必延年益壽。
PROV|4|11|我已指教你走智慧的道， 引導你行正直的路。
PROV|4|12|你行走，腳步沒有阻礙； 你奔跑，也不致跌倒。
PROV|4|13|要持定訓誨，不可放鬆； 要謹守它，因為它是你的生命。
PROV|4|14|不可行惡人的路， 不要走壞人的道；
PROV|4|15|要躲避，不可經過， 要轉離而去。
PROV|4|16|他們若不行惡，難以成眠， 不使人跌倒，就睡臥不安；
PROV|4|17|因為他們以邪惡當餅吃， 以暴力當酒喝。
PROV|4|18|但義人的路好像黎明的光， 越照越明，直到正午。
PROV|4|19|惡人的道幽暗， 自己不知因何跌倒。
PROV|4|20|我兒啊，要留心聽我的話， 側耳聽我的言語，
PROV|4|21|不可使它們偏離你的眼目， 要存記在你心中。
PROV|4|22|因為找到它們的，就找到生命， 得到全身的醫治。
PROV|4|23|你要保守你心，勝過保守一切， 因為生命的泉源由心發出。
PROV|4|24|要離開歪曲的口， 轉離偏邪的嘴唇。
PROV|4|25|你的兩眼要向前看， 你的雙目 直視前方。
PROV|4|26|要修平 你腳下的路， 你一切的道就必穩固。
PROV|4|27|不可偏左偏右， 你的腳要離開邪惡。
PROV|5|1|我兒啊，要留心聽我的智慧， 側耳聽我的聰明，
PROV|5|2|為要使你謹守智謀， 嘴唇保護知識。
PROV|5|3|因為陌生女子的嘴唇滴下蜂蜜， 她的口比油更滑，
PROV|5|4|後來卻苦似茵蔯， 銳利如兩刃的劍。
PROV|5|5|她的腳墜落死亡， 她的腳步踏入陰間，
PROV|5|6|她無法找到生命的道路， 她的路變遷不定，自己卻不知道。
PROV|5|7|孩子們，現在要聽從我， 不可離棄我口中的言語。
PROV|5|8|你所行的道要遠離她， 不可靠近她家的門口，
PROV|5|9|免得將你的尊榮給別人， 將你的歲月給殘忍的人；
PROV|5|10|免得陌生人滿得你的財富， 你勞苦所得的歸入外邦人的家。
PROV|5|11|在你人生終結，你皮肉和身體衰殘時， 你必唉聲嘆氣，
PROV|5|12|說：「我為何恨惡管教， 心裏輕看責備呢？
PROV|5|13|我不聽從教師的話， 也沒有側耳聽那教導我的。
PROV|5|14|在聚集的會眾中， 我幾乎墜入深淵。」
PROV|5|15|你要喝自己池中的水， 飲自己井裏的活水。
PROV|5|16|你的泉源豈可溢流在外？ 你的河水豈可流到街上？
PROV|5|17|讓它們惟獨歸你， 不可與陌生人同享。
PROV|5|18|要使你的泉源蒙福， 要喜愛你年輕時的妻子。
PROV|5|19|她如可愛的母鹿，如優美的母羊， 願她的胸懷使你時時滿足， 願你常常迷戀她的愛情。
PROV|5|20|我兒啊，你為何迷戀陌生女子？ 為何擁抱外邦女子的胸懷？
PROV|5|21|因為人所行的道都在耶和華眼前， 他察驗 人一切的路。
PROV|5|22|惡人被自己的罪孽抓住， 被自己罪惡的繩索纏繞。
PROV|5|23|他因不受管教而死亡， 因極度愚昧而走迷。
PROV|6|1|我兒啊，你若為朋友擔保， 替陌生人擊掌，
PROV|6|2|你就被口中的言語套住， 被嘴裏的言語抓住。
PROV|6|3|我兒啊，你既落在朋友手中，當這樣行才可救自己： 你要謙卑自己，去懇求你的朋友。
PROV|6|4|不要讓你的眼睛睡覺， 不可容你的眼皮打盹。
PROV|6|5|要救自己，如羚羊脫離獵人的手， 如鳥脫離捕鳥人的手。
PROV|6|6|懶惰人哪， 你去察看螞蟻的動作，就可得智慧。
PROV|6|7|螞蟻沒有領袖， 沒有官長，沒有君王，
PROV|6|8|尚且在夏天預備食物， 在收割時儲存糧食。
PROV|6|9|懶惰人哪，你要睡到幾時呢？ 你甚麼時候才睡醒呢？
PROV|6|10|再睡片時，打盹片時， 抱著雙臂躺臥片時，
PROV|6|11|你的貧窮就如盜賊來到， 你的貧乏彷彿拿盾牌的人來臨。
PROV|6|12|無賴的惡徒 行事全憑歪曲的口，
PROV|6|13|他眨眼傳神， 以腳示意，用指點劃，
PROV|6|14|存心乖謬， 常設惡謀，散播紛爭。
PROV|6|15|所以，災難必突然臨到他， 他必頃刻被毀，無從醫治。
PROV|6|16|耶和華所恨惡的有六樣， 他心所憎惡的共有七樣：
PROV|6|17|就是高傲的眼，撒謊的舌， 殺害無辜的手，
PROV|6|18|圖謀惡計的心， 飛奔行惡的腳，
PROV|6|19|口吐謊言的假證人， 並在弟兄間散播紛爭的人。
PROV|6|20|我兒啊，要遵守你父親的命令， 不可離棄你母親的教誨。
PROV|6|21|要常掛在你心上， 繫在你頸項上。
PROV|6|22|你行走，她必引導你， 你躺臥，她必保護你， 你睡醒，她必與你談論。
PROV|6|23|因為誡命是燈，教誨是光， 管教的責備是生命的道，
PROV|6|24|要保護你遠離邪惡的婦女， 遠離外邦女子諂媚的舌頭。
PROV|6|25|你不要因她的美色而動心， 也不要被她的眼皮勾引。
PROV|6|26|因為連最後一塊餅都會被妓女拿走 ； 有夫之婦會獵取寶貴的生命。
PROV|6|27|人若兜火在懷中， 他的衣服豈能不燒著呢？
PROV|6|28|人若走在火炭上， 他的腳豈能不燙傷呢？
PROV|6|29|與鄰舍之妻同寢的，也是如此， 凡親近她的，難免受罰。
PROV|6|30|賊因飢餓偷竊充飢， 人不藐視他，
PROV|6|31|但若被抓到，要賠償七倍， 他必賠上家中一切財物。
PROV|6|32|與婦人行姦淫的，便是無知， 做這事的，必毀了自己。
PROV|6|33|他必受損傷和羞辱， 他的羞恥不得消除。
PROV|6|34|丈夫因嫉恨發怒， 報仇的時候絕不留情。
PROV|6|35|他不接受任何賠償， 你送許多禮物，他也不肯和解。
PROV|7|1|我兒啊，要遵守我的言語， 存記我的命令。
PROV|7|2|遵守我的命令就得存活， 謹守我的教誨，好像保護眼中的瞳人。
PROV|7|3|要繫在你指頭上， 刻在你心版上。
PROV|7|4|對智慧說「你是我的姊妹」， 稱呼聰明為親人，
PROV|7|5|她就保護你遠離陌生女子， 遠離油嘴滑舌的外邦女子。
PROV|7|6|我曾在我房屋的窗戶內， 透過窗格子往外觀看，
PROV|7|7|看見在愚蒙人中， 注意到孩兒中有一個無知的青年，
PROV|7|8|從街上經過，靠近她的巷口， 直往她家的路去，
PROV|7|9|在黃昏，在傍晚， 在半夜，黑暗之中。
PROV|7|10|看哪，有一個女子來迎接他， 是妓女的打扮，有詭詐的心思。
PROV|7|11|她喧嚷，不守約束， 她的腳在家裏留不住，
PROV|7|12|有時在街市，有時在廣場， 或在各巷口等候。
PROV|7|13|她拉住那青年吻他， 厚著臉皮對他說：
PROV|7|14|「我已獻了平安祭， 今日我還了所許的願。
PROV|7|15|因此，我出來迎接你， 渴望見你的面，我總算找到你了！
PROV|7|16|我已在床上鋪好被單， 是 埃及 麻織的花紋布，
PROV|7|17|又用沒藥、沉香、桂皮 薰了我的床。
PROV|7|18|你來，讓我們飽享愛情，直到早晨， 讓我們彼此親愛歡樂。
PROV|7|19|因為我丈夫不在家， 出門遠行，
PROV|7|20|他手帶錢囊， 要到月圓才回家。」
PROV|7|21|這女子用許多巧言引誘他， 用諂媚的嘴唇催逼他。
PROV|7|22|青年立刻跟隨她，好像牛去被宰殺， 又像愚妄人帶著腳鐐去受刑，
PROV|7|23|直到箭穿進他的肝，如同雀鳥急投羅網， 卻不知會賠上自己的生命。
PROV|7|24|孩子們，現在要聽從我， 要留心聽我口中的言語。
PROV|7|25|你的心不可偏向她的道， 不要誤入她的迷途。
PROV|7|26|因為她擊倒許多人， 無數的人被她殺戮 。
PROV|7|27|她的家是在陰間之路， 下到死亡之宮。
PROV|8|1|智慧豈不呼喚？ 聰明豈不揚聲？
PROV|8|2|她站立在十字路口， 在道路旁高處的頂上，
PROV|8|3|在城門旁，城門口， 入口處，她呼喊：
PROV|8|4|「人哪，我呼喚你們， 我向世人揚聲。
PROV|8|5|愚蒙人哪，你們要學習靈巧， 愚昧人哪，你們的心要明辨。
PROV|8|6|你們當聽，因我要說尊貴的事， 我要張開嘴唇講正直的事。
PROV|8|7|我的口要發出真理， 我的嘴唇憎惡邪惡。
PROV|8|8|我口中的言語都是公義， 並無奸詐和歪曲。
PROV|8|9|聰明人看為正確， 有知識的，都以為正直。
PROV|8|10|你們當領受我的訓誨，勝過領受銀子， 寧得知識，強如得上選的金子。
PROV|8|11|「因為智慧比寶石更美， 一切可喜愛的都不足與其比較。
PROV|8|12|我－智慧以靈巧為居所， 又尋得知識和智謀。
PROV|8|13|敬畏耶和華就是恨惡邪惡； 我恨惡驕傲、狂妄、惡道，和乖謬的口。
PROV|8|14|我有策略和健全的知識， 我聰明，又有能力。
PROV|8|15|君王藉我治國， 王子藉我定公平，
PROV|8|16|王公貴族，所有公義的審判官， 都藉我掌權 。
PROV|8|17|愛我的，我也愛他， 懇切尋求我的，必尋見。
PROV|8|18|財富和尊榮在我， 恆久的財寶和繁榮 也在我。
PROV|8|19|我的果實勝過金子，強如純金， 我的出產超乎上選的銀子。
PROV|8|20|我在公義的道上走， 在公平的路中行，
PROV|8|21|使愛我的承受財產， 充滿他們的庫房。
PROV|8|22|「耶和華在造化的起頭， 在太初創造萬物之先，就有 了我。
PROV|8|23|從亙古，從太初， 未有大地以前，我已被立。
PROV|8|24|沒有深淵， 沒有大水的泉源，我已出生。
PROV|8|25|大山未曾奠定， 小山未有之先，我已出生。
PROV|8|26|那時，他還沒有創造大地和田野， 並世上頭一撮塵土。
PROV|8|27|他立高天，我在那裏， 他在淵面的周圍劃出圓圈，
PROV|8|28|上使穹蒼堅硬， 下使淵源穩固，
PROV|8|29|為滄海定出範圍，使水不越過界限， 奠定大地的根基。
PROV|8|30|那時，我在他旁邊為工程師， 天天充滿喜樂，時時在他面前歡笑，
PROV|8|31|在他的全地歡笑， 喜愛住在人世間。
PROV|8|32|「孩子們，現在要聽從我， 謹守我道的有福了。
PROV|8|33|要聽訓誨，得智慧， 不可棄絕。
PROV|8|34|聽從我，天天在我門口守望， 在我門框旁等候的，那人有福了。
PROV|8|35|因為尋得我的，就尋得生命， 他必蒙耶和華的恩惠。
PROV|8|36|得罪我的，害了自己的生命， 凡恨惡我的，喜愛死亡。」
PROV|9|1|智慧建造房屋， 鑿成七根柱子，
PROV|9|2|宰殺牲畜，調好美酒， 又擺設筵席，
PROV|9|3|派遣女僕出去， 自己在城中至高處呼喚：
PROV|9|4|「誰是愚蒙的人，讓他轉到這裏來！」 又對那無知的人說：
PROV|9|5|「你們來，吃我的餅， 喝我調的酒。
PROV|9|6|你們要離棄愚蒙，就得存活， 並要走明智的道路。」
PROV|9|7|糾正傲慢人的，必招羞辱， 責備惡人的，必被侮辱。
PROV|9|8|不要責備傲慢人，免得他恨你； 要責備智慧人，他必愛你。
PROV|9|9|教導智慧人，他就越有智慧， 指示義人，他就增長學問。
PROV|9|10|敬畏耶和華是智慧的開端， 認識至聖者便是聰明。
PROV|9|11|藉著我，你的日子必增多， 你生命的年數也必加添。
PROV|9|12|你若有智慧，是自己有智慧； 你若傲慢，就自己承擔。
PROV|9|13|愚昧的女子喧嚷， 她是愚蒙，一無所知。
PROV|9|14|她坐在自己家門口， 在城中高處的座位上，
PROV|9|15|呼喚過路的， 向那些在路上直走的人說：
PROV|9|16|「誰是愚蒙的人，讓他轉到這裏來！」 又對那無知的人說：
PROV|9|17|「偷來的水是甜的， 暗藏的餅是美的。」
PROV|9|18|人卻不知有陰魂在她那裏， 她召喚的人是在陰間的深處。
PROV|10|1|所羅門的箴言： 智慧之子使父親喜樂； 愚昧之子使母親擔憂。
PROV|10|2|不義之財毫無益處； 惟有公義能救人脫離死亡。
PROV|10|3|耶和華不使義人捱餓； 惡人所欲的，耶和華必拒絕。
PROV|10|4|手懶的，必致窮乏； 手勤的，卻要富足。
PROV|10|5|夏天儲存的，是智慧之子； 收割時沉睡的，是蒙羞之子。
PROV|10|6|福祉臨到義人頭上； 惡人的口藏匿殘暴。
PROV|10|7|義人的稱號帶來祝福； 惡人的名字必然敗壞。
PROV|10|8|智慧的心，領受誡命； 愚妄的嘴唇，必致傾倒。
PROV|10|9|行正直路的，步步安穩； 走彎曲道的，必致敗露。
PROV|10|10|擠眉弄眼的，使人憂患； 愚妄的嘴唇，必致傾倒。
PROV|10|11|義人的口是生命的泉源； 惡人的口藏匿殘暴。
PROV|10|12|恨能挑啟爭端； 愛能遮掩一切過錯。
PROV|10|13|聰明人嘴裏有智慧； 無知的人背上受刑杖。
PROV|10|14|智慧人積存知識； 愚妄人的口速致敗壞。
PROV|10|15|有錢人的財物是他堅固的城； 貧寒人的貧乏使他敗壞。
PROV|10|16|義人的報酬帶來生命； 惡人的所得用來犯罪。
PROV|10|17|遵守訓誨的，行在生命道上； 離棄責備的，走迷了路。
PROV|10|18|隱藏怨恨的，有說謊的嘴唇； 口出毀謗的，是愚昧人。
PROV|10|19|多言多語難免有過； 節制嘴唇是有智慧。
PROV|10|20|義人的舌如上選的銀子； 惡人的心所值無幾。
PROV|10|21|義人的嘴唇牧養多人； 愚妄人因無知而死亡。
PROV|10|22|耶和華所賜的福使人富足， 並不加上憂慮。
PROV|10|23|愚昧人以行惡為樂； 聰明人以智慧為樂。
PROV|10|24|惡人所怕的，必臨到他； 義人的心願，必蒙應允。
PROV|10|25|暴風一過，惡人歸於無有； 義人卻有永久的根基。
PROV|10|26|懶惰人使那差他的人， 如醋倒牙，如煙薰目。
PROV|10|27|敬畏耶和華使人長壽； 惡人的年歲必減少。
PROV|10|28|義人的盼望帶來喜樂； 惡人的指望必致滅沒。
PROV|10|29|耶和華的道是正直人的保障； 卻成了作惡人的敗壞。
PROV|10|30|義人永不動搖； 惡人不得住在地上。
PROV|10|31|義人的口結出智慧； 乖謬的舌必被割斷。
PROV|10|32|義人的嘴唇懂得令人喜悅； 惡人的口只知乖謬。
PROV|11|1|詭詐的天平為耶和華所憎惡； 公平的法碼為他所喜悅。
PROV|11|2|驕傲來，羞恥也來； 謙遜人卻有智慧。
PROV|11|3|正直人的純正必引導自己； 奸詐人的邪惡必毀滅自己。
PROV|11|4|遭怒的日子錢財無益； 惟有公義能救人脫離死亡。
PROV|11|5|完全人的義修平自己的路； 但惡人必因自己的惡跌倒。
PROV|11|6|正直人的義必拯救自己； 奸詐人必被自己的慾望纏住。
PROV|11|7|惡人一死，他的指望就滅絕； 罪人的盼望也必滅絕。
PROV|11|8|義人得脫離患難， 有惡人來代替他。
PROV|11|9|不虔敬的人用口敗壞鄰舍； 義人卻因知識得救。
PROV|11|10|義人享福，全城喜樂； 惡人滅亡，人人歡呼。
PROV|11|11|因正直人的祝福，城必升高； 因邪惡人的口，它必傾覆。
PROV|11|12|藐視鄰舍的，便是無知； 聰明人卻靜默不言。
PROV|11|13|到處傳話的，洩漏機密； 內心老實的，保守祕密。
PROV|11|14|無智謀，民就敗落； 謀士多，就必得勝。
PROV|11|15|為陌生人擔保的，必受虧損； 恨惡擊掌的，卻得安穩。
PROV|11|16|恩慈的婦女得尊榮； 強壯的男子得財富。
PROV|11|17|仁慈的人善待自己； 殘忍的人擾害己身。
PROV|11|18|惡人做事，得虛幻的報酬； 撒公義種子的，得實在的報償。
PROV|11|19|真正行義的，必得生命； 追求邪惡的，必致死亡。
PROV|11|20|心中歪曲的，為耶和華所憎惡； 行為正直的，為他所喜悅。
PROV|11|21|擊掌保證，惡人難免受罰； 義人的後裔必得拯救。
PROV|11|22|婦女美貌而無見識， 如同金環戴在豬鼻上。
PROV|11|23|義人的心願盡是好的； 惡人的指望卻帶來憤怒。
PROV|11|24|有施捨的，錢財增添； 吝惜過度，反致窮乏。
PROV|11|25|慷慨待人，必然豐裕； 滋潤人的，連自己也得滋潤。
PROV|11|26|屯糧不賣的，百姓必詛咒他； 願意出售的，祝福臨到頭上。
PROV|11|27|懇切求善的，就求得恩寵； 但那求惡的，惡必臨到他。
PROV|11|28|倚靠財富的，自己必跌倒； 義人必興旺如綠葉。
PROV|11|29|擾害己家的，必承受虛空 ； 愚妄人作心中有智慧者的僕人。
PROV|11|30|義人的果實是生命樹； 智慧人必能得人。
PROV|11|31|看哪，義人在地上尚且受報， 何況惡人和罪人呢？
PROV|12|1|喜愛管教的，就是喜愛知識； 恨惡責備的，卻像畜牲。
PROV|12|2|善人蒙耶和華的恩寵； 設詭計的，耶和華必定罪。
PROV|12|3|人靠惡行不能堅立； 義人的根必不動搖。
PROV|12|4|才德的妻子是丈夫的冠冕； 蒙羞的婦人使丈夫骨頭朽爛。
PROV|12|5|義人的思念是公平； 惡人的計謀是詭詐。
PROV|12|6|惡人的言論埋伏流人的血； 正直人的口卻拯救人。
PROV|12|7|惡人傾覆，歸於無有； 義人的家卻屹立不倒。
PROV|12|8|人按自己的智慧得稱讚； 心中偏邪的，必被藐視。
PROV|12|9|被人藐視，但有自己僕人 的， 勝過妄自尊大，卻缺乏食物。
PROV|12|10|義人顧惜他牲畜的命； 惡人的憐憫也是殘忍。
PROV|12|11|耕種自己田地的，必得飽食； 追求虛浮的，卻是無知。
PROV|12|12|惡人想得壞人的獵物； 義人的根結出果實。
PROV|12|13|嘴唇的過錯是惡人的圈套； 但義人必脫離患難。
PROV|12|14|人因口所結的果實，必飽得美福； 人手所做的，必歸到自己身上。
PROV|12|15|愚妄人所行的，在自己眼中看為正直； 惟智慧人從善如流。
PROV|12|16|愚妄人的惱怒立時顯露； 通達人卻能忍辱。
PROV|12|17|說出真話的，顯明公義； 作假見證的，顯出詭詐。
PROV|12|18|說話浮躁，猶如刺刀； 智慧人的舌頭卻能醫治。
PROV|12|19|誠實的嘴唇永遠堅立； 說謊的舌頭只存片時。
PROV|12|20|圖謀惡事的，心存詭詐； 勸人和睦的，便得喜樂。
PROV|12|21|義人不遭災害； 惡人滿受禍患。
PROV|12|22|說謊的嘴唇，為耶和華所憎惡； 行事誠實，為他所喜悅。
PROV|12|23|通達人隱藏知識； 愚昧人的心彰顯愚昧。
PROV|12|24|殷勤人的手必掌權； 懶惰的人必服苦役。
PROV|12|25|人心憂慮，就必沉重； 一句良言，使心歡樂。
PROV|12|26|義人引導他的鄰舍 ； 惡人的道叫人迷失。
PROV|12|27|懶惰的人不烤獵物； 殷勤的人卻得寶貴的財物。
PROV|12|28|在公義的路上有生命； 在其道上並無死亡。
PROV|13|1|智慧之子聽父親的訓誨； 傲慢人不聽責備。
PROV|13|2|人因口所結的果實，必享美福； 奸詐人卻意圖殘暴。
PROV|13|3|謹慎守口的，得保生命； 大張嘴唇的，必致敗亡。
PROV|13|4|懶惰的人奢求，卻無所得； 殷勤的人必然豐裕。
PROV|13|5|義人恨惡謊言； 惡人可憎可恥。
PROV|13|6|行為純正的，有公義保護； 犯罪的，被罪惡傾覆。
PROV|13|7|假冒富足的，一無所有； 裝作窮乏的，多有財物。
PROV|13|8|財富可作人的生命贖價； 窮乏人卻聽不見威嚇的話。
PROV|13|9|義人的光使人歡喜 ； 惡人的燈要熄滅。
PROV|13|10|驕傲挑啟紛爭； 聽勸言卻有智慧。
PROV|13|11|不勞而獲之財 必減少； 逐漸積蓄的必增多。
PROV|13|12|盼望遲延，令人心憂； 願望實現，就是得到生命樹。
PROV|13|13|藐視訓言的，自取滅亡； 敬畏誡命的，必得善報。
PROV|13|14|智慧人的教誨是生命的泉源， 使人避開死亡的圈套。
PROV|13|15|美好的見識使人得寵； 奸詐人的道路恆久奸詐 。
PROV|13|16|通達人都憑知識行事； 愚昧人張揚自己的愚昧。
PROV|13|17|邪惡的使者必陷入禍患； 忠信的使臣帶來醫治。
PROV|13|18|棄絕管教的，必貧窮受辱； 領受責備的，必享尊榮。
PROV|13|19|願望實現，心覺甘甜； 遠離惡事，為愚昧人所憎惡。
PROV|13|20|與智慧人同行的，必得智慧； 和愚昧人作伴的，必受虧損。
PROV|13|21|禍患追趕罪人； 義人卻得善報。
PROV|13|22|善人給子孫遺留產業； 罪人積財卻歸義人。
PROV|13|23|窮乏人開墾的地雖多產糧食， 卻因不公而被奪走。
PROV|13|24|不忍用杖打兒子的，是恨惡他； 疼愛兒子的，勤加管教。
PROV|13|25|義人吃喝食慾滿足； 惡人肚腹卻是缺乏。
PROV|14|1|婦人的智慧建立家室； 愚昧卻親手拆毀它 。
PROV|14|2|行事正直的，敬畏耶和華； 偏離正路的，卻藐視他。
PROV|14|3|在愚妄人的口中有驕傲的杖； 智慧人的嘴唇必保護自己。
PROV|14|4|沒有牛，槽就空空； 土產豐盛卻憑牛的力氣。
PROV|14|5|誠實的證人不說謊； 虛假的證人口吐謊言。
PROV|14|6|傲慢人枉尋智慧； 聰明人易得知識。
PROV|14|7|不要到愚昧人面前， 你無法從他嘴唇裏知道知識。
PROV|14|8|通達人的智慧使他認清自己的道路； 愚昧人的愚昧卻是自欺。
PROV|14|9|愚妄人嘲笑贖愆祭 ； 但正直人蒙悅納。
PROV|14|10|心中的苦楚，只有自己知道； 心裏的喜樂，陌生人無法分享。
PROV|14|11|惡人的房屋必倒塌； 正直人的帳棚必興旺。
PROV|14|12|有一條路，人以為正， 至終成為死亡之路。
PROV|14|13|人在喜笑中，心也會憂愁； 快樂的終點就是愁苦。
PROV|14|14|心中背道的，必滿嘗其果； 善人必從自己的行為得到回報。
PROV|14|15|無知的人甚麼話都信； 通達人謹慎自己的腳步。
PROV|14|16|智慧人有所懼怕，就遠離惡事； 愚昧人卻狂傲自恃。
PROV|14|17|輕易發怒的，行事愚昧； 擅長詭計的，被人恨惡。
PROV|14|18|愚蒙人承受愚昧為產業； 通達人得知識為冠冕。
PROV|14|19|壞人在善人面前俯伏； 惡人在義人門口也是如此。
PROV|14|20|窮乏人，連鄰舍也恨他； 有錢人，愛他的人眾多。
PROV|14|21|藐視鄰舍的，這人有罪； 施恩給困苦人的，這人有福。
PROV|14|22|謀惡的，豈非走入迷途？ 謀善的，有慈愛和誠實。
PROV|14|23|任何勤勞總有收穫； 僅耍嘴皮必致窮乏。
PROV|14|24|智慧人的冠冕是富有智慧； 愚昧人的愚昧終究是愚昧。
PROV|14|25|誠實作證，救人性命； 口吐謊言是詭詐。
PROV|14|26|敬畏耶和華的，大有倚靠； 他的兒女也有避難所。
PROV|14|27|敬畏耶和華是生命的泉源， 使人離開死亡的圈套。
PROV|14|28|君王的榮耀在乎民多； 沒有百姓，王就衰敗。
PROV|14|29|不輕易發怒的，大有聰明； 性情暴躁的，大顯愚昧。
PROV|14|30|平靜的心使肉體有生氣； 嫉妒使骨頭朽爛。
PROV|14|31|欺壓貧寒人的，是蔑視造他的主； 憐憫貧窮人的，是尊敬主。
PROV|14|32|惡人因所行的惡必被推倒； 義人臨死 ，有所投靠。
PROV|14|33|智慧安居在聰明人的心中， 在愚昧人的心中卻不認識 。
PROV|14|34|公義使邦國高舉； 罪惡是百姓的羞辱。
PROV|14|35|君王的恩寵臨到智慧的臣僕； 但其憤怒臨到蒙羞的臣僕。
PROV|15|1|回答柔和，使怒消退； 言語粗暴，觸動怒氣。
PROV|15|2|智慧人的舌善發知識； 愚昧人的口吐出愚昧。
PROV|15|3|耶和華的眼目無處不在， 惡人善人，他都鑒察。
PROV|15|4|溫良的舌是生命樹； 邪惡的舌使人心碎。
PROV|15|5|愚妄人藐視父親的管教； 領受責備，使人精明。
PROV|15|6|義人家中多有財富； 惡人獲利反受擾害。
PROV|15|7|智慧人的嘴傳揚知識； 愚昧人的心並非如此。
PROV|15|8|惡人獻祭，為耶和華所憎惡； 正直人祈禱，為他所喜悅。
PROV|15|9|惡人的道路，為耶和華所憎惡； 追求公義的，為他所喜愛。
PROV|15|10|背棄正路的，必受嚴刑； 恨惡責備的，必致死亡。
PROV|15|11|陰間和冥府 尚且在耶和華面前， 何況世人的心呢？
PROV|15|12|傲慢人不愛受責備， 也不去接近智慧人。
PROV|15|13|心中喜樂，面有喜色； 心裏憂愁，靈就憂傷。
PROV|15|14|聰明人的心追求知識； 愚昧人的口吞吃愚昧。
PROV|15|15|困苦人的日子都是愁苦； 心中歡暢的，常享宴席。
PROV|15|16|財寶稀少，敬畏耶和華， 強如財寶眾多，煩亂不安。
PROV|15|17|有愛，吃素菜， 強如相恨，吃肥牛。
PROV|15|18|暴怒的人挑啟爭端； 忍怒的人止息紛爭。
PROV|15|19|懶惰人的道像荊棘的籬笆； 正直人的路是平坦大道。
PROV|15|20|智慧之子使父親喜樂； 愚昧的人藐視母親。
PROV|15|21|無知的人以愚昧為樂； 聰明的人按正直而行。
PROV|15|22|不先商議，所謀無效； 謀士眾多，所謀得成。
PROV|15|23|口善應對，自覺喜樂； 話合其時，何等美好。
PROV|15|24|生命之道使智慧人上升， 使他遠離底下的陰間。
PROV|15|25|耶和華必拆毀驕傲人的家， 卻要立定寡婦的地界。
PROV|15|26|惡謀為耶和華所憎惡； 良言卻是純淨的。
PROV|15|27|暴力歛財的，擾害己家； 恨惡賄賂的，必得存活。
PROV|15|28|義人的心思量應答； 惡人的口吐出惡言。
PROV|15|29|耶和華遠離惡人， 卻聽義人的祈禱。
PROV|15|30|眼睛發光，使心喜樂； 好的信息，滋潤骨頭。
PROV|15|31|耳聽使人得生命的責備， 必居住在智慧人之中。
PROV|15|32|棄絕管教的，輕看自己的生命； 領受責備的，卻得智慧的心。
PROV|15|33|敬畏耶和華是智慧的訓誨； 要得尊榮，先有謙卑。
PROV|16|1|心中的籌謀在乎人， 舌頭的應對出於耶和華。
PROV|16|2|人一切所行的，在自己眼中看為純潔， 惟有耶和華衡量人的內心。
PROV|16|3|你所做的，要交託耶和華， 你所謀的，就必堅立。
PROV|16|4|耶和華造萬物各適其用， 就是惡人也為禍患的日子所造。
PROV|16|5|凡心裏驕傲的，為耶和華所憎惡； 擊掌保證，他難免受罰。
PROV|16|6|因慈愛和信實，罪孽得贖； 敬畏耶和華的，遠離惡事。
PROV|16|7|人所行的若蒙耶和華喜悅， 耶和華也使仇敵與他和好。
PROV|16|8|少獲利，行事公義， 強如多獲利，行事不義。
PROV|16|9|人心籌算自己的道路； 惟耶和華指引他的腳步。
PROV|16|10|王的嘴唇有聖言， 審判之時，他的口必不差錯。
PROV|16|11|公道的秤和天平屬耶和華， 囊中一切的法碼是他所定。
PROV|16|12|作惡，為王所憎惡， 因國位是靠公義堅立。
PROV|16|13|公義的嘴唇，王喜悅， 說正直話的，他喜愛。
PROV|16|14|王的震怒是死亡的使者， 但智慧人能平息王怒。
PROV|16|15|王臉上的光使人有生命， 他的恩惠好像雲帶來的春雨。
PROV|16|16|得智慧勝過得金子， 選聰明強如選銀子。
PROV|16|17|正直人的道遠離惡事， 謹守己路的，保全性命。
PROV|16|18|驕傲在敗壞以先， 內心高傲在跌倒之前。
PROV|16|19|心裏謙卑與困苦人來往， 強如與驕傲人同分戰利品。
PROV|16|20|留心訓言的 ，必得福樂； 倚靠耶和華的，這人有福。
PROV|16|21|心中有智慧的，必稱為聰明人； 嘴唇的甜言，增長人的學問。
PROV|16|22|人有智慧就有生命的泉源； 愚妄人必受愚妄的懲戒。
PROV|16|23|智慧人的心使他的口謹慎， 又使他的嘴唇增長學問。
PROV|16|24|良言如同蜂巢， 使心甘甜，使骨得醫治。
PROV|16|25|有一條路，人以為正， 至終卻成為死亡之路。
PROV|16|26|勞力的人為自己勞力， 因為他的口腹催逼他。
PROV|16|27|匪徒圖謀奸惡， 嘴唇上的言語彷彿燒焦的火。
PROV|16|28|乖謬的人散播紛爭， 造謠的離間密友。
PROV|16|29|殘暴的人引誘鄰舍， 領他走不好的道路。
PROV|16|30|緊閉雙目的，圖謀乖謬； 緊咬嘴唇的，成就惡事。
PROV|16|31|白髮是榮耀的冠冕， 行在公義道上的，必能得著。
PROV|16|32|不輕易發怒的，勝過勇士； 控制自己脾氣的，強如取城。
PROV|16|33|人雖可擲籤在膝上， 定事卻由耶和華。
PROV|17|1|一塊乾餅，大家相安； 勝過宴席滿屋，大家相爭。
PROV|17|2|明智的僕人必管轄蒙羞的兒子， 並在兄弟中同分產業。
PROV|17|3|鼎為煉銀，爐為煉金， 惟有耶和華熬煉人心。
PROV|17|4|行惡的，留心聽惡毒的嘴唇； 說謊的，側耳聽邪惡的舌頭。
PROV|17|5|譏笑窮乏人的，是蔑視造他的主； 幸災樂禍的，難免受罰。
PROV|17|6|子孫為老人的冠冕； 父母是兒女的榮耀。
PROV|17|7|愚頑人說美言並不相宜， 君子說謊言也不合宜。
PROV|17|8|賄賂在餽贈者的眼中看為玉石， 隨處運轉都得順利。
PROV|17|9|包容過錯的，尋求友愛； 喋喋不休的，離間密友。
PROV|17|10|一句責備的話深入聰明人的心， 強如打愚昧人一百下。
PROV|17|11|惡人只尋求背叛， 殘忍的使者必奉差攻擊他。
PROV|17|12|寧可遇見失喪小熊的母熊， 也不願遇見正行愚昧的愚昧人。
PROV|17|13|以惡報善的， 禍患必不離他的家。
PROV|17|14|紛爭掀起，如同缺口的水； 因此，爭端尚未爆發就當制止。
PROV|17|15|定惡人為義的，定義人為有罪的， 都為耶和華所憎惡。
PROV|17|16|愚昧人既無知， 為何手拿銀錢去買智慧呢？
PROV|17|17|朋友時常親愛， 弟兄為患難而生。
PROV|17|18|在鄰舍面前擊掌擔保的， 是無知的人。
PROV|17|19|喜愛爭吵的，是喜愛過犯； 門蓋得高的，自取敗壞。
PROV|17|20|心中歪曲的，得不著福樂； 舌頭顛倒是非的，陷在禍患中。
PROV|17|21|生愚昧之子的，自己必愁苦； 愚頑人的父親毫無喜樂。
PROV|17|22|喜樂的心能治好疾病； 憂傷的靈使骨頭枯乾。
PROV|17|23|惡人暗中受賄賂， 以致彎曲公正的路。
PROV|17|24|聰明人面前有智慧； 愚昧人眼望地的盡頭。
PROV|17|25|愚昧的兒子使父親愁煩， 使那生他的母親憂苦。
PROV|17|26|刑罰義人實為不善， 責打正直的君子也不宜。
PROV|17|27|節制言語的，有見識； 性情溫良的人，有聰明。
PROV|17|28|愚妄人若靜默不言，可算為智慧， 閉上嘴唇也可算為聰明。
PROV|18|1|孤僻的人只顧自己的心願 ， 他鄙視一切健全的知識。
PROV|18|2|愚昧人不喜愛聰明， 只喜愛表達自己的心意。
PROV|18|3|邪惡來，藐視跟著來； 羞恥到，辱罵同時到。
PROV|18|4|人的口所講的話如同深水， 智慧之泉如湧流的河水。
PROV|18|5|偏袒惡人的情面，是不好的。 審判時使義人受屈，也是不善。
PROV|18|6|愚昧人的嘴唇挑起爭端， 一開口就招鞭打。
PROV|18|7|愚昧人的口自取敗壞， 他的嘴唇是自己生命的圈套。
PROV|18|8|造謠者的話如同美食， 深入人的肚腹。
PROV|18|9|做工懈怠的， 是破壞者的兄弟。
PROV|18|10|耶和華的名是堅固臺， 義人奔入就得安穩。
PROV|18|11|有錢人的財物是他堅固的城， 在他幻想中，猶如高牆。
PROV|18|12|敗壞之先，人心驕傲； 要得尊榮，先有謙卑。
PROV|18|13|未聽完就回話的， 就是他的愚昧和羞辱。
PROV|18|14|人的心靈忍耐疾病； 心靈憂傷，誰能承當呢？
PROV|18|15|聰明人的心得知識； 智慧人的耳求知識。
PROV|18|16|人的禮物為他開路， 引他到高位的人面前。
PROV|18|17|先訴情由的，似乎有理； 另一人來到，就察出實情。
PROV|18|18|掣籤能止息紛爭， 也能化解雙方激烈的爭辯。
PROV|18|19|被冒犯的弟兄 強如難以攻下的堅城； 紛爭如同城堡的門閂。
PROV|18|20|人的肚腹必因口所結的果實飽足； 他必因嘴唇所出的感到滿足。
PROV|18|21|生死在舌頭的掌握之下， 喜愛弄舌的，必吃它所結的果實。
PROV|18|22|得著妻子的，得著好處， 他是蒙了耶和華的恩惠。
PROV|18|23|窮乏人說哀求的話； 有錢人卻用威嚇的話回答。
PROV|18|24|朋友太多的人，必受損害 ； 但有一知己比兄弟更親密。
PROV|19|1|行為純正的窮乏人 勝過嘴唇歪曲的愚昧人。
PROV|19|2|熱心而無見識，實為不善； 腳步急快的，易入歧途。
PROV|19|3|人因愚昧自毀前途， 他的心卻埋怨耶和華。
PROV|19|4|財富使朋友增多； 貧寒人連僅有的朋友也離棄他。
PROV|19|5|作假見證的，難免受罰； 口吐謊言的，不能逃脫。
PROV|19|6|有權貴的，許多人求他賞臉； 愛送禮的，人都作他的朋友。
PROV|19|7|窮乏人連兄弟都恨他， 何況朋友，更是遠離他！ 他用言語追隨，他們卻不在。
PROV|19|8|得著智慧的，愛惜生命； 持守聰明的，尋得好處。
PROV|19|9|作假見證的，難免受罰； 口吐謊言的，必定滅亡。
PROV|19|10|愚昧人奢華度日並不相宜， 僕人管轄王子，也不應該。
PROV|19|11|人有見識就不輕易發怒， 寬恕人的過失便是自己的榮耀。
PROV|19|12|王的憤怒好像獅子吼叫； 他的恩惠卻如草上的甘露。
PROV|19|13|愚昧的兒子是父親的禍患， 妻子的爭吵如雨連連滴漏。
PROV|19|14|房屋錢財是祖宗所遺留的； 惟有賢慧的妻是耶和華所賜的。
PROV|19|15|懶惰使人沉睡， 懈怠的人必捱餓。
PROV|19|16|遵守誡命的，保全生命； 輕忽己路的，必致死亡。
PROV|19|17|憐憫貧寒人的，就是借給耶和華， 他的報償，耶和華必歸還他。
PROV|19|18|趁還有指望，管教你的兒子， 不可執意摧毀他。
PROV|19|19|暴怒的人必受懲罰， 你若救他，必須再救。
PROV|19|20|要聽勸言，接受訓誨， 使你終久有智慧。
PROV|19|21|人心多有計謀； 惟有耶和華的籌算才能成就。
PROV|19|22|仁慈的人令人喜愛 ， 窮乏人強如說謊言的。
PROV|19|23|敬畏耶和華的，得著生命， 他必飽足安居，不遭禍患。
PROV|19|24|懶惰人把手埋入盤裏， 連縮回送進口中也不肯。
PROV|19|25|責打傲慢人，能使無知的人變精明； 責備聰明人，他就明白知識。
PROV|19|26|虐待父親、驅逐母親的， 是蒙羞致辱之子。
PROV|19|27|我兒啊，停止聽 那叫你偏離知識言語的教導 。
PROV|19|28|卑劣的見證嘲笑公平， 惡人的口吞下罪孽。
PROV|19|29|刑罰是為傲慢人預備的， 鞭打則是為愚昧人的背預備的。
PROV|20|1|酒能使人傲慢，烈酒使人喧嚷， 凡沉溺其中的，都無智慧。
PROV|20|2|王的威嚇如獅子吼叫， 激怒他的是自害己命。
PROV|20|3|止息紛爭是人的尊榮， 愚妄人爭鬧不休。
PROV|20|4|懶惰人因冬寒不去耕種， 到收割時，他去尋找，一無所得。
PROV|20|5|人心中的籌算如同深水， 惟聰明人才能汲引出來。
PROV|20|6|很多人聲稱自己忠信， 但誠信的人誰能遇著呢？
PROV|20|7|義人行為純正， 他後代的子孫有福了！
PROV|20|8|王坐在審判的位上， 以眼目驅散一切邪惡。
PROV|20|9|誰能說：「我已經潔淨了我的心， 脫淨了我的罪？」
PROV|20|10|兩樣的法碼和兩樣的伊法 ， 都為耶和華所憎惡。
PROV|20|11|孩童的行動或純潔，或正直， 都以行為顯明自己。
PROV|20|12|能聽的耳，能看的眼， 二者都為耶和華所造。
PROV|20|13|不要貪睡，免致貧窮； 眼要睜開，就可吃飽。
PROV|20|14|買東西的說：「不好，不好！」 及至離去，他卻自誇。
PROV|20|15|有金子和許多寶石， 惟知識的嘴唇是貴重的珍寶。
PROV|20|16|誰為陌生人擔保，就拿誰的衣服； 誰為外邦人作保，誰就要承當。
PROV|20|17|靠謊言而得的食物，令人愉悅； 到後來，他的口必充滿碎石。
PROV|20|18|計謀憑籌算立定， 打仗要憑智謀。
PROV|20|19|到處傳話的，洩漏機密； 口無遮攔的，不可與他結交。
PROV|20|20|咒罵父母的， 他的燈必熄滅，在漆黑中。
PROV|20|21|起初很快得來的產業， 終久卻不是福。
PROV|20|22|你不要說：「我要以惡報惡」； 要等候耶和華，他必拯救你。
PROV|20|23|兩樣的法碼為耶和華所憎惡， 詭詐的天平也為不善。
PROV|20|24|人的腳步為耶和華所定， 人豈能明白自己的道路呢？
PROV|20|25|人冒失地聲稱：「這是神聖的！」 許願之後才細想，就是自陷圈套。
PROV|20|26|智慧的王驅散惡人， 用輪子滾過他們。
PROV|20|27|人的靈是耶和華的燈， 鑒察人的內心深處。
PROV|20|28|慈愛和誠實庇護君王， 他的王位因慈愛而立穩。
PROV|20|29|強壯是青年的榮耀； 白髮為老人的尊榮。
PROV|20|30|鞭傷除淨邪惡， 責打可潔淨人心深處。
PROV|21|1|王的心在耶和華手中像河水， 他能使它隨意流轉。
PROV|21|2|人一切所行的，在自己眼中看為正直， 惟有耶和華衡量人心。
PROV|21|3|行公義和公平 比獻祭更蒙耶和華悅納。
PROV|21|4|眼高心傲，就是惡人的燈， 都是罪。
PROV|21|5|殷勤籌劃的，足致豐裕； 行事急躁的，必致缺乏。
PROV|21|6|用詭詐之舌所得的財富 如被吹散的霧氣，趨向滅亡 。
PROV|21|7|惡人的殘暴必掃去自己， 因他們不肯按公平行事。
PROV|21|8|有罪的人其路彎曲； 純潔的人行為正直。
PROV|21|9|寧可住在房頂的一角， 也不與好爭吵的婦人同住。
PROV|21|10|惡人的心渴想邪惡， 他的眼並不憐憫鄰舍。
PROV|21|11|傲慢人受懲罰，愚蒙人可得智慧； 智慧人受訓誨，便得知識。
PROV|21|12|公義的上帝 鑒察惡人的家， 他傾覆惡人，以致滅亡。
PROV|21|13|塞耳不聽貧寒人哀求的， 他自己呼求，也不蒙應允。
PROV|21|14|暗中送的禮物挽回怒氣， 懷裏的賄賂能止息暴怒。
PROV|21|15|秉公行義使義人喜樂， 卻使作惡的人敗壞。
PROV|21|16|人偏離智慧的路， 必與陰魂為伍 。
PROV|21|17|愛宴樂的，必致窮乏； 貪愛酒和油的，必不富足。
PROV|21|18|惡人作義人的贖價， 奸詐人代替正直人。
PROV|21|19|寧可住在曠野之地， 也不與爭吵易怒的婦人同住。
PROV|21|20|智慧人的居所積蓄寶物與膏油 ； 愚昧人卻揮霍一空。
PROV|21|21|追求公義慈愛的， 就尋得生命、公義 和尊榮。
PROV|21|22|智慧人爬上勇士的城牆， 摧毀他所倚靠的堡壘。
PROV|21|23|謹守口和舌的， 就保護自己免受災難。
PROV|21|24|心驕氣傲的人名叫傲慢， 他行事出於狂妄驕傲。
PROV|21|25|懶惰人的慾望害死自己， 因為他的手不肯做工；
PROV|21|26|有人終日貪得無饜， 義人卻施捨而不吝惜。
PROV|21|27|惡人獻的祭是可憎的， 何況他存惡意來獻呢？
PROV|21|28|不實的見證必消滅； 惟聆聽真情的，他的證詞有力。
PROV|21|29|惡人臉無羞恥； 正直人行事堅定 。
PROV|21|30|沒有人能以智慧、聰明、 謀略抵擋耶和華。
PROV|21|31|馬是為打仗之日預備的； 得勝卻在於耶和華。
PROV|22|1|美名勝過大財， 宏恩強如金銀。
PROV|22|2|有錢人與窮乏人相遇 ， 他們都為耶和華所造。
PROV|22|3|通達人見禍就藏躲； 愚蒙人卻前往受害。
PROV|22|4|敬畏耶和華心存謙卑， 就得財富、尊榮、生命為賞賜。
PROV|22|5|歪曲的人路上有荊棘和羅網， 保護自己生命的，必要遠離。
PROV|22|6|教養孩童走當行的道， 就是到老他也不偏離。
PROV|22|7|有錢人管轄窮乏人， 欠債的是債主的僕人。
PROV|22|8|撒不義種子的必收割災禍， 他逞怒的杖也必廢掉。
PROV|22|9|眼目仁慈的必蒙福， 因他將食物分給貧寒人。
PROV|22|10|趕出傲慢人，爭端就消除， 紛爭和羞辱也必止息。
PROV|22|11|喜愛清心，嘴唇有恩言的， 王必與他為友。
PROV|22|12|耶和華的眼目保護知識， 卻毀壞奸詐人的言語。
PROV|22|13|懶惰人說：「外面有獅子， 我在街上必被殺害。」
PROV|22|14|陌生女子的口是深坑， 耶和華所憎惡的，必陷在其中。
PROV|22|15|愚昧迷住孩童的心， 用管教的杖可以遠遠趕除。
PROV|22|16|欺壓貧寒人為要利己的， 並送禮給有錢人的，都必缺乏。
PROV|22|17|你要側耳聽智慧人的言語 ， 留心領會我的知識。
PROV|22|18|你若心中存記， 嘴唇也準備就緒，這是美的。
PROV|22|19|我今日特地指教你， 為要使你倚靠耶和華。
PROV|22|20|謀略和知識的美事 ， 我豈沒有寫給你嗎？
PROV|22|21|要使你明白真情實理， 好將實情回覆那差你來的人。
PROV|22|22|不可因人貧寒就搶奪他， 也不可在城門口欺壓困苦人，
PROV|22|23|因耶和華必為他們辯護， 也必奪取那搶奪者的命。
PROV|22|24|不可結交好生氣的人， 也不可與暴怒的人來往，
PROV|22|25|恐怕你效法他的行為， 自己就陷在圈套裏。
PROV|22|26|不要為人擊掌擔保， 也不要為債務作保。
PROV|22|27|你若沒有甚麼可償還， 何必使人奪去你睡臥的床呢？
PROV|22|28|祖先所立的地界， 你不可挪移。
PROV|22|29|你看見辦事殷勤的人嗎？ 他必侍立在君王面前， 不在平庸的人面前。
PROV|23|1|你若與長官坐席， 要留意在你面前的是誰。
PROV|23|2|你若是胃口大的人， 就當拿刀放在喉嚨上。
PROV|23|3|不可貪戀長官的美食， 因為那是欺哄人的食物。
PROV|23|4|不要勞碌求富， 要有聰明來節制。
PROV|23|5|你定睛在財富，它就消失， 因為它必長翅膀，如鷹向天飛去。
PROV|23|6|守財奴 的飯，你不要吃， 也不要貪戀他的美味；
PROV|23|7|因為他的心怎樣算計 ， 他為人就是這樣。 他雖對你說：請吃，請喝， 他的心卻與你相背。
PROV|23|8|你所吃的那點食物必吐出來， 你恭維的話語也必落空。
PROV|23|9|不要說話給愚昧人聽， 因他必藐視你智慧的言語。
PROV|23|10|不可挪移古時的地界， 也不可侵佔孤兒的田地，
PROV|23|11|因他們的救贖者 大有能力， 他必向你為他們辯護。
PROV|23|12|你要留心領受訓誨， 側耳聽從知識的言語。
PROV|23|13|不可不管教孩童， 因為你用杖打他，他不會死。
PROV|23|14|你用杖打他， 就可以救他的性命免下陰間。
PROV|23|15|我兒啊，你若心存智慧， 我的心就甚歡喜。
PROV|23|16|你的嘴唇若說正直話， 我的心腸也必快樂。
PROV|23|17|你的心不要羨慕罪人， 卻要羨慕常常敬畏耶和華的人，
PROV|23|18|因為你必有前途， 你的指望也不致斷絕。
PROV|23|19|我兒啊，你當聽，當存智慧， 好在正道上引導你的心。
PROV|23|20|不可與好飲酒的人在一起， 也不要跟貪吃肉的人來往，
PROV|23|21|因為貪食好酒的，必致貧窮， 愛睡覺的，必穿破爛衣服。
PROV|23|22|你要聽從生你的父親； 不可因母親年老而輕看她。
PROV|23|23|你當獲得真理，不可出賣， 智慧、訓誨和聰明也是一樣。
PROV|23|24|義人的父親必大大快樂， 生智慧兒子的，必因他歡喜。
PROV|23|25|願你的父母歡喜， 願那生你的母親快樂。
PROV|23|26|我兒啊，要將你的心歸我， 你的眼目也要喜愛 我的道路。
PROV|23|27|妓女是深坑， 外邦女子是窄井。
PROV|23|28|她像強盜埋伏， 她使奸詐的人增多。
PROV|23|29|誰有禍患？誰有災難？ 誰有紛爭？誰有焦慮？ 誰無故受傷？誰的眼目紅赤？
PROV|23|30|就是那流連飲酒的人， 常去尋找調和的酒。
PROV|23|31|酒發紅，在杯中閃爍時， 你不可觀看； 雖下咽舒暢， 終究它必咬你如蛇，刺你如毒蛇。
PROV|23|32|
PROV|23|33|你的眼睛必看見怪異的事， 你的心必發出乖謬的話。
PROV|23|34|你必像躺在深海中， 或臥在桅杆頂上，
PROV|23|35|說：「人擊打我，但我未受傷， 重擊我，我不覺得。 我幾時清醒， 還要再去尋酒。」
PROV|24|1|你不要嫉妒惡人， 也不要渴望與他們相處，
PROV|24|2|因為他們的心圖謀暴行， 他們的嘴唇談論奸惡。
PROV|24|3|房屋因智慧建造， 因聰明立穩；
PROV|24|4|又因知識， 屋內充滿各樣美好寶貴的財物。
PROV|24|5|有智慧的勇士大有能力， 有知識的人力上加力。
PROV|24|6|你去打仗，要憑智謀； 謀士眾多，就必得勝。
PROV|24|7|對愚妄人，智慧高不可及， 所以他在城門不敢開口。
PROV|24|8|圖謀行惡的， 必稱為奸詐人。
PROV|24|9|愚妄人的籌劃盡是罪惡， 傲慢者為人所憎惡。
PROV|24|10|在患難時你若灰心， 你的力量就微小。
PROV|24|11|人被拉到死亡，你要解救； 人將被殺，你須攔阻。
PROV|24|12|你若說：「看哪，這事我們不知道」， 那衡量人心的豈不明白嗎？ 保護你性命的豈不知道嗎？ 他豈不按各人所做的報應各人嗎？
PROV|24|13|我兒啊，你要吃蜜，因為它是美好的， 要讓甘甜的蜜滴入你的口。
PROV|24|14|你要知道，智慧對你的生命正像如此。 你若找著，必有前途， 你的指望也不致斷絕。
PROV|24|15|你這惡人，不可埋伏攻擊義人的家， 也不可毀壞他安居之所。
PROV|24|16|因為義人雖七次跌倒，仍必興起； 惡人卻被禍患傾倒。
PROV|24|17|你的仇敵跌倒，你不要歡喜， 他傾倒，你的心不要快樂；
PROV|24|18|恐怕耶和華看見就不喜悅， 將怒氣從仇敵身上轉過來。
PROV|24|19|不要為作惡的心懷不平， 也不要嫉妒惡人，
PROV|24|20|因為壞人沒有前途， 惡人的燈也必熄滅。
PROV|24|21|我兒啊，你要敬畏耶和華與君王， 不可結交反覆無常的人，
PROV|24|22|因為他們的災難必忽然興起。 誰能知道耶和華與君王所施行的毀滅呢？
PROV|24|23|以下也是智慧人的箴言： 審判時看人情面是不好的。
PROV|24|24|對惡人說「你是義人」的， 萬民必詛咒，萬族必惱恨。
PROV|24|25|責備惡人的，必得喜悅， 美好的福分也必臨到他。
PROV|24|26|應對合宜的， 猶如與人親吻。
PROV|24|27|你要在外面預備材料， 在田間為自己準備齊全， 然後才建造你的房屋。
PROV|24|28|不可無故作證反對鄰舍， 也不可用嘴唇欺騙人。
PROV|24|29|不可說：「人怎樣待我，我也怎樣待他， 我必照他所做的報復他。」
PROV|24|30|我經過懶惰人的田地， 走過無知人的葡萄園，
PROV|24|31|看哪，它長滿了荊棘， 蕁麻蓋地面， 石牆也坍塌了。
PROV|24|32|我看見就留心思想， 我看著就領受訓誨。
PROV|24|33|再睡片時，打盹片時， 抱著雙臂躺臥片時，
PROV|24|34|你的貧窮就如盜賊來到， 你的貧乏彷彿拿盾牌的人來臨。
PROV|25|1|以下也是 所羅門 的箴言，是 猶大 王 希西家 的人所謄錄的。
PROV|25|2|隱藏事情是上帝的榮耀； 查明事情乃君王的榮耀。
PROV|25|3|天之高，地之深， 君王之心測不透。
PROV|25|4|除去銀子的渣滓， 銀匠就做出器皿來。
PROV|25|5|除去王面前的惡人， 國位就靠公義堅立。
PROV|25|6|不可在君王面前妄自尊大， 也不要站在大人的位上。
PROV|25|7|寧可讓人家說「請你上到這裏來」， 強如在你覲見的貴人面前令你退下。
PROV|25|8|不要冒失出去與人爭訟 ， 免得你的鄰舍羞辱你， 最後你就不知怎麼做。
PROV|25|9|要與鄰舍爭辯你的案情， 不可洩漏他人的隱密，
PROV|25|10|恐怕聽見的人責罵你， 你就難以擺脫臭名。
PROV|25|11|一句話說得合宜， 就如金蘋果在銀網子裏
PROV|25|12|智慧人的勸戒在順從的人耳中， 好像金環和金首飾。
PROV|25|13|忠信的使者對那差他的人， 就如收割時有冰雪的涼氣， 使主人的心舒暢。
PROV|25|14|人空誇禮物而不肯贈送， 就好像有風有雲卻無雨。
PROV|25|15|恆常的忍耐可以勸服君王， 柔和的舌頭能折斷骨頭。
PROV|25|16|你得了蜜，吃夠就好， 免得過飽就吐出來。
PROV|25|17|你的腳要少進鄰舍的家， 免得他厭煩你，恨惡你。
PROV|25|18|作假見證陷害鄰舍的， 就是大錘，是利刀，是快箭。
PROV|25|19|患難時倚靠奸詐的人， 好像牙齒斷裂，又如腳脫臼。
PROV|25|20|對傷心的人唱歌， 就如冷天脫他的衣服， 又如在鹼上倒醋 。
PROV|25|21|你的仇敵若餓了，就給他飯吃， 若渴了，就給他水喝；
PROV|25|22|因為你這樣做，就是把炭火堆在他的頭上， 耶和華必回報你。
PROV|25|23|正如北風生雨， 毀謗的舌頭也生怒容。
PROV|25|24|寧可住在房頂的一角， 也不與好爭吵的婦人同住。
PROV|25|25|有好消息從遙遠的地方來， 就如涼水滋潤口渴的人。
PROV|25|26|義人在惡人面前退縮， 好像攪渾之泉，污染之井。
PROV|25|27|吃蜜過多是不好的， 自求榮耀也是一樣。
PROV|25|28|人不克制自己的心， 就像毀壞的城沒有牆。
PROV|26|1|愚昧人得尊榮不相宜， 正如夏天落雪，收割時下雨。
PROV|26|2|詛咒不會無故臨到 ， 正如麻雀掠過，燕子翻飛。
PROV|26|3|鞭子是為打馬，轡頭是為勒驢， 刑杖正是為打愚昧人的背。
PROV|26|4|不要照愚昧人的愚昧話回答他， 免得你與他一樣。
PROV|26|5|要照愚昧人的愚昧話回答他， 免得他自以為有智慧。
PROV|26|6|藉愚昧人的手寄信的， 就像砍斷雙腳，喝下殘暴。
PROV|26|7|箴言在愚昧人的口中， 正如瘸子的腳懸空無用。
PROV|26|8|將尊榮給愚昧人的， 就像石頭綁在彈弓上。
PROV|26|9|箴言在愚昧人的口中， 好像荊棘刺入醉漢的手。
PROV|26|10|雇愚昧人的，與雇過路人的， 就像弓箭手射傷任何人。
PROV|26|11|愚昧人重複做愚昧之事， 就如狗轉過來吃自己所吐的。
PROV|26|12|你看見自以為有智慧的人嗎？ 愚昧人比他更有指望。
PROV|26|13|懶惰人說：「道路有猛獅， 街上有壯獅。」
PROV|26|14|懶惰人在床上， 就像門在軸心上轉動一樣。
PROV|26|15|懶惰人把手埋入盤裏， 就是送進口中也覺得累。
PROV|26|16|懶惰人眼看自己 比七個善於應對的人更有智慧。
PROV|26|17|過路時捲入與己無關的紛爭， 好像人揪住狗耳一般。
PROV|26|18|人欺騙鄰舍，卻說 「我只是開玩笑而已」， 他就像瘋狂的人拋擲致死的火把和利箭。
PROV|26|19|
PROV|26|20|火缺了柴就必熄滅； 無人造謠，紛爭就止息。
PROV|26|21|好爭吵的人煽動爭端， 就如餘火加炭，火上加柴一樣。
PROV|26|22|造謠者的話如同美食， 深入人的肚腹。
PROV|26|23|火熱的 嘴唇，邪惡的心， 好像銀渣包在瓦器上。
PROV|26|24|仇敵用嘴唇掩飾， 心裏卻藏著詭詐；
PROV|26|25|他用甜言蜜語，你不能相信他， 因為他心中有七樣可憎惡的事。
PROV|26|26|他雖用詭詐掩飾怨恨， 他的邪惡必在集會中顯露。
PROV|26|27|挖陷坑的，自己必陷在其中； 滾石頭的，石頭反滾在他身上。
PROV|26|28|虛謊的舌憎恨他所壓傷的人； 諂媚的口敗壞人的事。
PROV|27|1|不要為明天自誇， 因為你不知道每天會發生何事。
PROV|27|2|要讓陌生人誇獎你，不可用口自誇； 讓外邦人稱讚你，不可用嘴唇稱讚自己。
PROV|27|3|石頭沉，沙土重， 愚妄人的惱怒比這兩樣更沉重。
PROV|27|4|憤怒為殘忍，怒氣像狂瀾， 惟有嫉妒，誰能擋得住呢？
PROV|27|5|當面的責備 勝過隱藏的愛情。
PROV|27|6|朋友加的傷痕出於忠誠； 敵人的親吻卻是多餘。
PROV|27|7|人吃飽了，厭惡蜂房的蜜； 人飢餓了，一切苦物都覺甘甜。
PROV|27|8|人離故鄉漂泊， 就像雀鳥離窩四處飛翔。
PROV|27|9|膏油與香料使人心喜悅， 朋友誠心的勸勉也是如此甘美。
PROV|27|10|你的朋友和父親的朋友， 你都不可離棄。 你遭難時，不要上兄弟的家去； 相近的鄰舍強如遠方的兄弟。
PROV|27|11|我兒啊，你要做智慧人，好叫我的心歡喜， 使我可以回答那辱罵我的人。
PROV|27|12|通達人見禍就藏躲； 愚蒙人卻前往受害。
PROV|27|13|誰為陌生人擔保，就拿誰的衣服； 誰為外邦女子作保，誰就要承當。
PROV|27|14|清晨起來大聲給朋友祝福的， 就算是詛咒他。
PROV|27|15|下雨天連連滴漏， 好爭吵的婦人就像這樣；
PROV|27|16|攔阻她的，就是攔阻風， 又像用右手抓油。
PROV|27|17|以鐵磨鐵，越磨越利， 朋友當面琢磨，也是如此。
PROV|27|18|看守無花果樹的，必吃樹上的果子； 敬奉主人的，必得尊榮。
PROV|27|19|水中照臉，彼此相符； 人心相映，也是如此。
PROV|27|20|陰間和冥府 永不滿足， 人的眼目也是如此。
PROV|27|21|鼎為煉銀，爐為煉金， 口中的稱讚也試煉人。
PROV|27|22|用杵把愚妄人與穀粒一同搗在臼中， 他的愚昧還是離不了他。
PROV|27|23|你要詳細知道你羊群的景況， 留心照顧你的牛群，
PROV|27|24|因為財富不能永留， 冠冕豈能存到萬代？
PROV|27|25|青草除去，嫩草長出， 山上的菜蔬也被採收。
PROV|27|26|綿羊可以做衣服， 公山羊可作田地的價值，
PROV|27|27|並有母山羊奶夠你吃， 夠你養家和女僕的生活。
PROV|28|1|惡人雖無人追趕也逃跑； 義人卻膽壯像獅子。
PROV|28|2|地上因有罪過，君王就多更換； 因聰明和有見識的人，國必長存。
PROV|28|3|窮乏人欺壓貧寒人， 好像暴雨掃過，不留糧食。
PROV|28|4|離棄律法的，誇獎惡人； 遵守律法的，卻與惡人相爭。
PROV|28|5|惡人不明白公義； 惟有尋求耶和華的，無不明白。
PROV|28|6|行為純正的窮乏人 勝過行事歪曲的有錢人。
PROV|28|7|謹守教誨的，是聰明之子； 與貪食者為伍的，卻羞辱其父。
PROV|28|8|人以厚利增加財富， 是給那憐憫貧寒人的積財。
PROV|28|9|轉耳不聽教誨的， 他的祈禱也可憎。
PROV|28|10|誘惑正直人行惡道的，必掉在自己的坑裏； 惟有完全人必承受福分。
PROV|28|11|有錢人自以為有智慧， 但聰明的貧寒人能看穿他。
PROV|28|12|義人高升，有大榮耀； 惡人興起，人就躲藏。
PROV|28|13|遮掩自己過犯的，必不順利； 承認且離棄過犯的，必蒙憐憫。
PROV|28|14|常存敬畏的，這人有福了； 心裏剛硬的，必陷在禍患裏。
PROV|28|15|邪惡的君王壓制貧民， 好像吼叫的獅子，又如覓食的熊。
PROV|28|16|無知的君王多行暴虐； 恨惡非分之財的，必年長日久。
PROV|28|17|背負流人血之罪的，必逃跑直到地府； 願無人幫助他！
PROV|28|18|行為正直的，必蒙拯救； 行事彎曲的，立時跌倒。
PROV|28|19|耕種自己田地的，糧食充足； 追求虛浮的，窮困潦倒。
PROV|28|20|誠實人必多得福； 想要急速發財的，難免受罰。
PROV|28|21|看人情面是不好的； 卻有人因一塊餅而犯法。
PROV|28|22|守財奴 想要急速發財， 卻不知窮乏必臨到他身上。
PROV|28|23|責備人的，後來蒙人喜悅， 多於那用舌頭諂媚人的。
PROV|28|24|搶奪父母竟說「這不是罪過」， 此人與毀滅者同類。
PROV|28|25|心中貪婪的，挑起爭端； 倚靠耶和華的，必得豐裕。
PROV|28|26|心中自以為是的，就是愚昧人； 憑智慧行事的，必蒙拯救。
PROV|28|27|賙濟窮乏人的，不致缺乏； 遮眼不看的，多受詛咒。
PROV|28|28|惡人興起，人就躲藏； 惡人敗亡，義人必增多。
PROV|29|1|人屢次受責罰，仍然硬著頸項， 他必頃刻被毀，無從醫治。
PROV|29|2|義人增多，民就喜樂； 惡人掌權，民就嘆息。
PROV|29|3|愛慕智慧的，使父親喜樂； 結交妓女的，卻浪費錢財。
PROV|29|4|王藉公平，使國堅定； 強索貢物的，使它毀壞。
PROV|29|5|諂媚鄰舍的， 就是設網羅絆他的腳。
PROV|29|6|惡人犯罪，自陷圈套； 惟獨義人歡呼喜樂。
PROV|29|7|義人關注貧寒人的案情； 惡人不明瞭這種知識。
PROV|29|8|傲慢人煽動全城； 智慧人止息眾怒。
PROV|29|9|智慧人與愚妄人有爭訟， 或怒或笑，總不得安寧。
PROV|29|10|好流人血的，恨惡完全人， 正直人卻顧惜 他的性命。
PROV|29|11|愚昧人怒氣全發； 智慧人自我平息。
PROV|29|12|君王若聽謊言， 他一切臣僕都是奸惡。
PROV|29|13|窮乏人和欺壓者相遇 ， 耶和華使他們的眼目明亮。
PROV|29|14|君王憑誠信判斷貧寒人， 他的國位必永遠堅立。
PROV|29|15|杖打和責備能增加智慧； 任性的少年使母親羞愧。
PROV|29|16|惡人多，過犯也加多， 義人必看見他們敗亡。
PROV|29|17|管教你的兒子，他就使你得安寧， 也使你心裏喜樂。
PROV|29|18|沒有異象 ，民就放肆； 惟遵守律法的，便為有福。
PROV|29|19|僕人不能靠言語受教； 他即使明白，也不回應。
PROV|29|20|你見過言語急躁的人嗎？ 愚昧人比他更有指望。
PROV|29|21|人將僕人從小嬌養， 至終必帶來憂傷 。
PROV|29|22|好生氣的人挑起爭端， 暴怒的人多多犯錯。
PROV|29|23|人的高傲使自己蒙羞； 心裏謙遜的，必得尊榮。
PROV|29|24|與盜賊分贓的，是恨惡自己的性命； 他雖聽見發誓的聲音，也不告訴人。
PROV|29|25|懼怕人的，陷入圈套； 惟有倚靠耶和華的，必得安穩。
PROV|29|26|求王恩的人多； 人獲公正來自耶和華。
PROV|29|27|不義之人，義人憎惡； 行事正直的，惡人憎惡。
PROV|30|1|雅基 的兒子、 瑪撒 人 亞古珥 的言語 ，是這人對 以鐵 和 烏甲 說的。
PROV|30|2|我比眾人更像畜牲， 也沒有人的聰明。
PROV|30|3|我沒有學好智慧， 也不認識至聖者。
PROV|30|4|誰升天又降下來？ 誰聚風在手掌中？ 誰包水在衣服裏？ 誰立定地的四極？ 他名叫甚麼？ 他兒子名叫甚麼？ 你知道嗎？
PROV|30|5|上帝的言語句句都是煉淨的， 投靠他的，他便作他們的盾牌。
PROV|30|6|你不可加添他的言語， 恐怕他責備你，你就顯為說謊的。
PROV|30|7|我求你兩件事， 在我未死之先，不要拒絕我：
PROV|30|8|求你使虛假和謊言遠離我， 使我不貧窮也不富足， 賜給我需用的飲食。
PROV|30|9|免得我飽足了，就不認你，說： 「耶和華是誰呢？」 又恐怕我貧窮就偷竊， 以致褻瀆我上帝的名。
PROV|30|10|不要向主人讒害他的僕人， 恐怕他詛咒你，你便算為有罪。
PROV|30|11|有一類人，詛咒父親， 不給母親祝福。
PROV|30|12|有一類人，自以為純潔， 卻沒有洗淨自己的污穢。
PROV|30|13|有一類人，眼目何其高傲， 眼皮也是高舉。
PROV|30|14|有一類人，牙如劍，齒如刀， 要吞滅地上的困苦人和世間的貧窮人。
PROV|30|15|水蛭有兩個女兒： 「給呀，給呀。」 有三樣不知足的， 不說「夠了」的有四樣：
PROV|30|16|陰間和不生育的子宮， 吸水不足的地，還有不說「夠了」的火。
PROV|30|17|嘲笑父親、藐視而不聽從母親的， 谷中的烏鴉必啄他的眼睛，小鷹也必吃它。
PROV|30|18|我所測不透的奇妙有三樣， 我所不知道的有四樣：
PROV|30|19|就是鷹在空中飛的道， 蛇在磐石上爬的道， 船在海中行的道， 男與女交合的道。
PROV|30|20|淫婦的道是這樣， 她吃了，把嘴一擦就說： 「我沒有行惡。」
PROV|30|21|使地震動的有三樣， 地承擔不起的有四樣：
PROV|30|22|就是僕人作王， 愚頑人吃得飽足，
PROV|30|23|令人憎惡的女子出嫁， 婢女取代她的女主人。
PROV|30|24|地上有四樣東西雖小，卻甚聰明：
PROV|30|25|螞蟻是無力之類， 卻在夏天預備糧食。
PROV|30|26|石獾並非強壯之類， 卻在巖石中造房子。
PROV|30|27|蝗蟲沒有君王， 卻分隊而出。
PROV|30|28|壁虎你用手就可抓住， 牠卻住在王宮。
PROV|30|29|腳步威武的有三樣， 行走威武的有四樣：
PROV|30|30|獅子－百獸中最勇猛的、 無論遇見甚麼絕不退縮，
PROV|30|31|獵狗，公山羊， 和有整排士兵的君王。
PROV|30|32|你若行事愚頑，自高自傲， 或是設計惡謀，就當用手摀口。
PROV|30|33|攪動牛奶必成乳酪， 扭鼻子必出血， 照樣，激發烈怒必挑起爭端。
PROV|31|1|瑪撒 王 利慕伊勒 的言語，就是他母親教導他的 。
PROV|31|2|我兒，怎麼了？ 我腹中生的兒，怎麼了？ 我許願而得的兒，怎麼了？
PROV|31|3|不要將你的精力給婦女， 也不要有敗壞君王的行為。
PROV|31|4|利慕伊勒 啊，君王不宜，君王不宜喝酒， 王子尋找烈酒也不相宜；
PROV|31|5|恐怕喝了就忘記所頒的法令， 顛倒所有困苦人的是非。
PROV|31|6|可以把烈酒給將亡的人喝， 把酒給心裏愁苦的人喝，
PROV|31|7|讓他喝了，就忘記他的貧窮， 不再記得他的苦楚。
PROV|31|8|你當為不能自辯的人 開口， 為所有孤獨無助者伸冤。
PROV|31|9|你當開口按公義判斷， 當為困苦和貧窮的人辯護。
PROV|31|10|才德的婦人誰能得著呢？ 她的價值遠勝過寶石。
PROV|31|11|她丈夫心裏信賴她， 必不缺少利益；
PROV|31|12|她終其一生， 使丈夫有益無損。
PROV|31|13|她尋找羊毛和麻， 歡喜用手做工。
PROV|31|14|她好像商船， 從遠方運來糧食，
PROV|31|15|未到黎明她就起來， 把食物分給家中的人， 將當做的工分派女僕。
PROV|31|16|她想得田地，就去買來， 用手中的成果栽葡萄園。
PROV|31|17|她以能力束腰， 使膀臂有力。
PROV|31|18|她覺得自己獲利不錯， 她的燈終夜不滅。
PROV|31|19|她伸手拿捲線桿， 她的手掌把住紡車。
PROV|31|20|她張手賙濟困苦人， 伸手幫助貧窮人。
PROV|31|21|她不因下雪為家裏的人擔心， 因為全家都穿上朱紅衣服。
PROV|31|22|她為自己製作被單， 她的衣服是細麻和紫色布做的。
PROV|31|23|她丈夫在城門口與本地的長老同坐， 為人所認識。
PROV|31|24|她做細麻布衣裳來賣， 又將腰帶賣給商家。
PROV|31|25|能力和威儀是她的衣服， 她想到日後的景況就喜笑。
PROV|31|26|她開口就發智慧， 她舌上有仁慈的教誨。
PROV|31|27|她管理家務， 並不吃閒飯。
PROV|31|28|她的兒女起來稱她有福， 她的丈夫也稱讚她：
PROV|31|29|「才德的女子很多， 惟獨你超過一切。」
PROV|31|30|魅力是虛假的，美貌是虛浮的； 惟敬畏耶和華的婦女必得稱讚。
PROV|31|31|她手中的成果你們要賞給她， 願她的工作在城門口榮耀她。
ECCL|1|1|在 耶路撒冷 作王、 大衛 的兒子、傳道者的言語。
ECCL|1|2|傳道者說：虛空的虛空， 虛空的虛空，全是虛空。
ECCL|1|3|人一切的勞碌， 就是他在日光之下的勞碌，有甚麼益處呢？
ECCL|1|4|一代過去，一代又來， 地卻永遠長存。
ECCL|1|5|太陽上升，太陽下落， 急歸所出之地。
ECCL|1|6|風往南颳，又向北轉， 不停旋轉，繞回原路。
ECCL|1|7|江河都往海裏流，海卻不滿； 江河從何處流，仍歸回原處。
ECCL|1|8|萬事令人厭倦， 人不能說盡。 眼看，看不飽； 耳聽，聽不足。
ECCL|1|9|已有的事，後必再有； 已行的事，後必再行。 日光之下並無新事。
ECCL|1|10|有一件事人指著說：「看，這是新的！」 它在我們以前的世代早已有了。
ECCL|1|11|已過的事，無人記念； 將來的事，後來的人也不記念。
ECCL|1|12|我傳道者在 耶路撒冷 作過 以色列 的王。
ECCL|1|13|我用智慧專心探尋、考察天下所發生的一切事：上帝給世人何等沉重的擔子，使他們在其中勞苦！
ECCL|1|14|我見日光之下所發生的一切事，看哪，全是虛空，全是捕風。
ECCL|1|15|彎曲的，不能變直； 缺乏的，不計其數。
ECCL|1|16|我心裏說：「看哪，我大有智慧，勝過在我以前所有統治 耶路撒冷 的人；我的心也多經歷智慧和知識的事。」
ECCL|1|17|我專心想要明白智慧，想要明白狂妄與愚昧，方知這也是捕風。
ECCL|1|18|因為多有智慧，就多有愁煩； 增加知識，就增加憂傷。
ECCL|2|1|我心裏說：「來吧，讓我用喜樂試試你，使你享福！」看哪，這也是虛空。
ECCL|2|2|論嬉笑，我說：「這是狂妄。」論享樂，「這有甚麼用呢？」
ECCL|2|3|我心以智慧引導我，我心裏探究，如何用酒使身體舒暢，如何抓住愚昧，直等我看明世人在天下短暫一生中，當行何事為美。
ECCL|2|4|我大興土木，為自己建造房屋，栽葡萄園，
ECCL|2|5|修造庭園和公園，在其中栽種各樣果樹，
ECCL|2|6|挖造水池，用以灌溉林中的幼樹。
ECCL|2|7|我買了僕婢，也有生在家中的僕婢；又有許多牛群羊群，勝過我以前所有在 耶路撒冷 的人。
ECCL|2|8|我為自己積蓄金銀，搜集各君王、各省份的財寶；又為自己得男女歌手和世人所喜愛的物，以及一個又一個的妃嬪。
ECCL|2|9|這樣，我就日漸昌盛，勝過我以前所有在 耶路撒冷 的人。我的智慧仍然存留。
ECCL|2|10|凡我眼所求的，我沒有克制它；我心所樂的，我沒有不享受。因我的心要為一切的勞碌快樂，這是我從一切勞碌中所得的報償 。
ECCL|2|11|後來，我回顧我手所經營的一切和我勞碌所做的工。看哪，全是虛空，全是捕風；在日光之下毫無益處。
ECCL|2|12|我轉而回顧智慧、狂妄和愚昧。在王以後來的人又如何呢？不過做先前所做的就是了。
ECCL|2|13|於是我看出智慧勝過愚昧，如同光明勝過黑暗。
ECCL|2|14|智慧人的眼目光明 ，愚昧人卻在黑暗裏行。但我知道他們都有相同的遭遇。
ECCL|2|15|我心裏就說：「愚昧人所遇見的，我也一樣遇見，那麼我何必更有智慧呢？」我心裏說：「這也是虛空。」
ECCL|2|16|智慧人和愚昧人一樣，不會長久被人記念，因為日後都被遺忘。可嘆！智慧人和愚昧人都一樣會死亡。
ECCL|2|17|於是我恨惡生命，因為在日光之下所發生的事我都以為煩惱，全是虛空，全是捕風。
ECCL|2|18|我恨惡一切的勞碌，就是我在日光之下所勞碌的，因為我所得的必須留給我以後的人。
ECCL|2|19|那人是智慧是愚昧，誰能知道呢？他竟要掌管我在日光之下用智慧勞碌所得的。這也是虛空。
ECCL|2|20|我轉想我在日光之下所勞碌的一切工作，心就絕望。
ECCL|2|21|因為有人用智慧、知識、靈巧勞碌工作，所得來的卻要遺留給未曾勞碌的人作產業。這也是虛空，大大不幸。
ECCL|2|22|人一切的勞碌操心，就是他在日光之下所勞碌的，又得著了甚麼呢？
ECCL|2|23|他日日憂慮，他的勞苦成為愁煩，連夜間心也不得休息。這也是虛空。
ECCL|2|24|難道一個人有吃有喝，且在勞碌中享福，不是福氣嗎？我看這也是出於上帝的手。
ECCL|2|25|論到吃用、享福，誰能勝過我呢？
ECCL|2|26|上帝喜愛誰，就給誰智慧、知識和喜樂；惟有罪人，上帝使他勞苦，將他所儲藏、所堆積的歸給上帝所喜愛的人。這也是虛空，也是捕風。
ECCL|3|1|凡事都有定期， 天下每一事務都有定時。
ECCL|3|2|生有時，死有時； 栽種有時，拔出 有時；
ECCL|3|3|殺戮有時，醫治有時； 拆毀有時，建造有時；
ECCL|3|4|哭有時，笑有時； 哀慟有時，跳舞有時；
ECCL|3|5|丟石頭有時，撿石頭有時； 懷抱有時，不抱有時；
ECCL|3|6|尋找有時，失落有時； 保存有時，拋棄有時；
ECCL|3|7|撕裂有時，縫補有時； 沉默有時，說話有時；
ECCL|3|8|喜愛有時，恨惡有時； 戰爭有時，和平有時。
ECCL|3|9|這樣，做事的人在他所勞碌的事上得到甚麼益處呢？
ECCL|3|10|我觀看上帝給世人的擔子，使他們在其中勞苦：
ECCL|3|11|上帝造萬物，各按其時成為美好，又將永恆安放在世人心裏；然而上帝從始至終的作為，人不能測透。
ECCL|3|12|我知道，人除了終身喜樂納福，沒有一件幸福的事。
ECCL|3|13|並且人人吃喝，在他的一切勞碌中享福，這也是上帝的賞賜。
ECCL|3|14|我知道上帝所做的都必存到永遠；無所增添，無所減少。上帝這樣做，是要人在他面前存敬畏的心。
ECCL|3|15|現今的事以前就有了，將來的事也早已有了，並且上帝使已過的事重新再來 。
ECCL|3|16|我又見日光之下，應有公平之處有奸惡，應有公義之處也有奸惡。
ECCL|3|17|我心裏說：「上帝必審判義人和惡人，因為在那裏，各樣事務，一切工作，都有定時。」
ECCL|3|18|我心裏說：「為世人的緣故，上帝考驗他們，讓他們看見自己不過像走獸一樣。」
ECCL|3|19|因為世人遭遇的，走獸也遭遇，所遭遇的都一樣：這個怎樣死，那個也怎樣死，他們都有一樣的氣息。人不能強於走獸，全是虛空；
ECCL|3|20|都歸一處，都是出於塵土，也都歸於塵土。
ECCL|3|21|誰知道人的氣息是往上升，走獸的氣息是下入地呢？
ECCL|3|22|總而言之，人能夠在他經營的事上喜樂，是最好不過了，因為這是他應得的報償。他身後的事誰能領他回來看呢？
ECCL|4|1|我轉而觀看日光之下所發生的一切欺壓之事。看哪，受欺壓的流淚，無人安慰；欺壓他們的有權勢，也無人安慰。
ECCL|4|2|因此，我讚歎那已死的死人，勝過那還活著的活人。
ECCL|4|3|但那尚未出生，就是未曾見過日光之下所發生之惡事的，比這兩種人更幸福。
ECCL|4|4|我見人因彼此嫉妒而有一切的勞碌和各樣工作的成就，這也是虛空，也是捕風。
ECCL|4|5|愚昧人抱著雙臂， 自食其肉。
ECCL|4|6|一掌滿滿而得享安靜， 勝過兩掌滿滿而勞碌捕風。
ECCL|4|7|我轉而觀看日光之下有一件虛空的事：
ECCL|4|8|有人孤單無雙，無子無兄弟，竟勞碌不息，眼目也不以財富為滿足。他說：「我勞碌，自己卻不享福，到底是為了誰呢？」這也是虛空，是極沉重的擔子。
ECCL|4|9|兩個人總比一個人好，他們勞碌同得美好的報償。
ECCL|4|10|若是跌倒，這人可以扶起他的同伴；倘若孤身跌倒，沒有別人扶起他來，這人就有禍了。
ECCL|4|11|再者，二人同睡就都暖和，一人獨睡怎能暖和呢？
ECCL|4|12|若遇敵攻擊，孤身難擋，二人就能抵擋他；三股合成的繩子不易折斷。
ECCL|4|13|貧窮而有智慧的年輕人，勝過年老不再納諫的愚昧王，
ECCL|4|14|那人從監牢裏出來作王，在國中原是出身貧寒。
ECCL|4|15|我見日光之下所有行走的活人，都跟隨那年輕人，就是接續作王的那位。
ECCL|4|16|他的百姓，就是他所治理的眾人，多得無數；但後來的人還是不喜歡他。這也是虛空，也是捕風。
ECCL|5|1|你到上帝的殿要謹慎你的腳步；近前聽，勝過愚昧人獻祭，他們不知道自己在作惡。
ECCL|5|2|在上帝面前你不可冒失開口，也不可心急發言；因為上帝在天上，你在地上，所以你的話語要少。
ECCL|5|3|事務多，令人做夢；話語多，顯出愚昧。
ECCL|5|4|你向上帝許願，還願不可遲延，因他不喜歡愚昧人，你許的願應當償還。
ECCL|5|5|你許願不還，不如不許。
ECCL|5|6|不可放任你的口使肉體犯罪，也不可在使者 面前說是錯許了。為何使上帝因你的聲音發怒，敗壞你手所做的呢？
ECCL|5|7|多夢多言，其中多有虛空，你只要敬畏上帝。
ECCL|5|8|你若在一個地區看見窮人受欺壓，公義公平被掠奪，不要因此驚奇；有一位高過居高位的在鑒察，在他們之上還有更高的。
ECCL|5|9|況且地的益處歸眾人，就是君王也受田地的供應。
ECCL|5|10|喜愛銀子的，不因得銀子滿足；喜愛財富的，也不因得利益知足。這也是虛空。
ECCL|5|11|貨物增添，吃的人也增添，物主得甚麼益處呢？不過眼看而已！
ECCL|5|12|勞碌的人不拘吃多吃少，睡得香甜；富人的豐足卻不容他睡覺。
ECCL|5|13|我見日光之下有一件令人憂傷的禍患，就是財主積存財富，反害自己。
ECCL|5|14|他因遭遇不幸 ，財產盡失；他生了兒子，手裏卻一無所有。
ECCL|5|15|他怎樣從母胎赤身而來，也必照樣赤身而去；他所勞碌得來的，手中分毫不能帶去。
ECCL|5|16|這是一件令人憂傷的禍患。他來的時候怎樣，去的時候也必怎樣。他為風勞碌有甚麼益處呢？
ECCL|5|17|並且他終身在黑暗中吃喝 ，多有煩惱、病痛和怒氣。
ECCL|5|18|看哪，我所見為善為美的，就是人在上帝賜他一生的日子吃喝，享受日光之下勞碌得來的好處，因為這是他應得的報償。
ECCL|5|19|而且，一個人蒙上帝賞賜財富與資產，又使他能享用，能獲取自己當有的報償 ，在他的勞碌中喜樂，這是上帝的賞賜。
ECCL|5|20|他不多思念自己一生的日子，因為上帝使他的心充滿喜樂。
ECCL|6|1|我見日光之下有一件禍患重壓在人身上，
ECCL|6|2|就是人蒙上帝賜他財富、資產和尊榮，以致他心裏所願的一樣都不缺，只是上帝使他不能享用，反被外人享用。這是虛空，也是禍患。
ECCL|6|3|人若生一百個兒子，活許多歲數；他即使壽命很長，心裏卻不因福樂而滿足，又不得埋葬；我說，那流掉的胎比他倒好。
ECCL|6|4|因為這胎虛虛而來，暗暗而去，名字被黑暗遮蔽，
ECCL|6|5|而且沒有見過天日，甚麼都不知道，這胎比那人倒享安息。
ECCL|6|6|那人雖然活千年，再活千年，卻不能享福；眾人豈不都歸同一個地方去嗎？
ECCL|6|7|人的勞碌都為口腹，心裏卻不知足。
ECCL|6|8|智慧人比愚昧人有甚麼益處呢？困苦人在眾人面前知道如何行，有甚麼益處呢？
ECCL|6|9|眼睛所看的比心裏妄想的倒好。這也是虛空，也是捕風。
ECCL|6|10|先前所有的，早已起了名，人早知道人是如何的，不能與比自己強壯的相爭。
ECCL|6|11|話語多，虛空也增多，這對人有甚麼益處呢？
ECCL|6|12|人一生虛度的日子，如影兒經過，誰知道甚麼才是對他有益呢？誰能告訴他身後在日光之下會發生甚麼事呢？
ECCL|7|1|名譽強如美好的膏油， 人死去的日子勝過他出生的日子。
ECCL|7|2|往喪家去， 強如往宴樂的家， 因為死是眾人的結局， 活人必將這事放在心上。
ECCL|7|3|憂愁強如喜笑， 因為面帶愁容，終必使心喜樂。
ECCL|7|4|智慧人的心在遭喪之家； 愚昧人的心在快樂之家。
ECCL|7|5|聽智慧人的責備， 強如聽愚昧人歌唱；
ECCL|7|6|因為愚昧人的笑聲， 好像鍋子下面燒荊棘的爆聲， 這也是虛空。
ECCL|7|7|勒索使智慧人變為愚妄， 賄賂能敗壞人的心。
ECCL|7|8|事情的終局強如它的起頭； 存心忍耐的，勝過居心驕傲的。
ECCL|7|9|你的心不要急躁惱怒， 因為惱怒存在愚昧人的懷中。
ECCL|7|10|不要說： 為甚麼先前的日子強過現今的日子呢？ 你這樣問不是出於智慧。
ECCL|7|11|智慧加上產業是美好的， 對見天日的人都有益處。
ECCL|7|12|因為智慧庇護人， 好像金錢庇護人一樣； 智慧能保全智慧者的生命， 這就是知識的益處。
ECCL|7|13|你要觀看上帝的作為， 誰能使他所彎曲的變直呢？
ECCL|7|14|順利時要喜樂；患難時當思考。上帝使這兩樣都發生，因此，人不知將會發生甚麼事。
ECCL|7|15|在虛度的日子裏，我見過各樣的事情，義人在他的義中滅亡，惡人在他的惡中倒享長壽。
ECCL|7|16|不要行義過分，也不要過於自逞智慧，何必自取敗亡呢？
ECCL|7|17|不要行惡過分，也不要為人愚昧，何必未到期而死呢？
ECCL|7|18|你持守這個，那個也不要鬆手才好。敬畏上帝的人，這一切都能兼得。
ECCL|7|19|智慧使擁有智慧的人比城中十個官長更有能力。
ECCL|7|20|其實世上沒有行善而不犯罪的義人。
ECCL|7|21|人所說的話，你不要都放在心上，免得聽見你的僕人詛咒你。
ECCL|7|22|因為你心裏知道，自己也曾屢次詛咒別人。
ECCL|7|23|我曾用智慧試驗這一切事，我說：「要得智慧。」智慧卻離我遠。
ECCL|7|24|萬事之理遙不可及，太深奧，誰能測透呢？
ECCL|7|25|我轉念，一心要知道，要考察，要尋求智慧和萬事的來由，要知道邪惡為愚昧，愚昧為狂妄。
ECCL|7|26|我發現有一種婦人比死還苦毒：她本身是陷阱，她的心是羅網，手是鎖鏈。凡蒙上帝喜愛的人必能躲開她；有罪的人卻被她纏住了。
ECCL|7|27|傳道者說：「你看，我考察一件又一件，為要尋求萬事的來由，這是我所尋得的：
ECCL|7|28|我繼續尋找，卻未找到；一千當中，我找到一個男的，但在這一切當中，卻找不到一個女的。
ECCL|7|29|你看，我所找到的只有一件，就是上帝造的人是正直的，但他們卻尋出許多詭計。」
ECCL|8|1|誰如 智慧人呢？ 誰知道事情的解釋呢？ 人的智慧使他的臉發光， 改變他臉上的暴戾之氣 。
ECCL|8|2|我勸你 因上帝誓言的緣故，當遵守王的命令。
ECCL|8|3|不要急躁離開王的面前，不要固執行惡，因為他凡事都隨自己心意而行。
ECCL|8|4|王的話本有權力，誰能對他說：「你在做甚麼？」
ECCL|8|5|凡遵守命令的，必不經歷禍患；智慧人的心知道適當的時機和必經的過程。
ECCL|8|6|各樣事務都有時機和過程，但人有苦難重壓在身。
ECCL|8|7|他不知道將來的事，其實將來如何，誰能告訴他呢？
ECCL|8|8|沒有人能掌握生命，將生命留住；也沒有人有權力掌管死期。這場爭戰無人能免；邪惡也不能救那行邪惡的人。
ECCL|8|9|這一切我都見過，我專心考察日光之下所發生的一切事，有時這人管轄那人，令他受害。
ECCL|8|10|我見惡人埋葬；從前他們進出聖地，他們在城中的作為被人忘記。這也是虛空。
ECCL|8|11|判罪之後不立刻執行，所以世人滿懷作惡的心思。
ECCL|8|12|罪人雖然作惡百次，倒享長壽；然而我也知道，福樂必臨到敬畏上帝的人，就是在他面前心存敬畏的人。
ECCL|8|13|惡人卻不得福樂，他的日子好像影兒不得長久，因為他不敬畏上帝。
ECCL|8|14|世上有一件虛空的事，就是義人所遭遇的，反而照惡人所做的；惡人所遭遇的，反而照義人所做的。我說，這也是虛空。
ECCL|8|15|我就稱讚快樂，原來人在日光之下，最大的福氣莫過於吃喝快樂；他在日光之下，上帝賜他一生的日子，要從勞碌中享受所得。
ECCL|8|16|我專心想要明白智慧，要觀看世上所發生的事。有人晝夜不得闔眼睡覺。
ECCL|8|17|我觀看上帝一切的作為，知道人不能探求日光之下所發生的事；任憑他費多少力探索，都找不出來，智慧人雖說他明白，仍不能找出來。
ECCL|9|1|我將這一切事放在心上，詳細研究這些，就知道義人和智慧人，並他們的作為都在上帝手中；或是愛，或是恨，都在他們面前，但人不能知道。
ECCL|9|2|凡臨到眾人的際遇都一樣：義人和惡人，好人 ，潔淨的人和不潔淨的人，獻祭的和不獻祭的，都一樣。好人如何，罪人也如何；起誓的如何，怕起誓的也如何。
ECCL|9|3|在日光之下發生的一切事中有一件禍患，就是眾人的際遇都一樣，並且世人的心充滿了惡；活著的時候心裏狂妄，後來就歸死人那裏去了。
ECCL|9|4|與一切活人相連的，那人還有指望，因為活著的狗勝過死了的獅子。
ECCL|9|5|活著的人知道必死；死了的人毫無所知，也不再得賞賜，因為他們的名 已被遺忘。
ECCL|9|6|他們的愛，他們的恨，他們的嫉妒，早就消滅了。在日光之下所發生的一切事，他們永不再有份了。
ECCL|9|7|你只管歡歡喜喜吃你的飯，心中快樂喝你的酒，因為上帝已經悅納你的作為。
ECCL|9|8|你的衣服要時時潔白，你頭上也不要缺少膏油。
ECCL|9|9|在你一生虛空的日子，就是上帝賜你在日光之下虛空 的日子，當與你所愛的妻快活度日，因為那是你一生中在日光之下勞碌所得的報償。
ECCL|9|10|凡你手所當做的事，要盡力去做；因為在你所必須去的陰間沒有工作，沒有謀算，沒有知識，也沒有智慧。
ECCL|9|11|我轉而回顧日光之下，快跑的未必能贏，強壯的未必戰勝，智慧的未必得糧食，聰明的未必得財富，有學問的未必得人喜悅，全在乎各人遇上的時候和機會。
ECCL|9|12|人不知道自己的定期。魚被險惡的網圈住，鳥被羅網捉住，禍患的時刻忽然臨到，世人陷在其中也是如此。
ECCL|9|13|我見日光之下有一樣智慧，在我看來是偉大的，
ECCL|9|14|就是有一人口稀少的小城，遇大君王前來攻擊，修築營壘，將城圍困。
ECCL|9|15|城中有一個貧窮的智慧人，他用智慧救了那城，卻沒有人記念那窮人。
ECCL|9|16|我就說，智慧勝過勇力；然而那貧窮人的智慧被人藐視，他的話也無人聽從。
ECCL|9|17|寧可聽智慧人安靜的話語，不聽掌權者在愚昧人中的喊聲。
ECCL|9|18|智慧勝過打仗的兵器；但一個罪人能敗壞許多善事。
ECCL|10|1|死蒼蠅使做香的膏油散發臭氣； 同樣，一點愚昧也能壓倒智慧和尊榮。
ECCL|10|2|智慧人的心居右； 愚昧人的心居左。
ECCL|10|3|愚昧人的行徑顯出無知， 對眾人說，他是愚昧人。
ECCL|10|4|掌權者的怒氣若向你發作， 不要離開你的本位， 因為鎮定能平息大過。
ECCL|10|5|我見日光之下有一件禍患， 似乎出於統治者的錯誤，
ECCL|10|6|就是愚昧人立在高位； 有錢人卻坐在低位。
ECCL|10|7|我見僕人騎馬， 王子像僕人在地上步行。
ECCL|10|8|挖陷坑的，自己必陷在其中； 拆城牆的，自己必被蛇咬。
ECCL|10|9|開鑿石頭的，會受損傷； 劈開木頭的，必遭危險。
ECCL|10|10|鐵器鈍了，若不將刃磨快，就必多費力氣； 但智慧的益處在於使人成功。
ECCL|10|11|尚未行法術，蛇若咬人， 行法術的人就得不到甚麼好處了。
ECCL|10|12|智慧人的口說出恩言； 愚昧人的嘴吞滅自己，
ECCL|10|13|他口中的話語起頭是愚昧， 終局是邪惡的狂妄。
ECCL|10|14|愚昧人多有話語。 人不知將來會發生甚麼事， 他身後的事誰能告訴他呢？
ECCL|10|15|愚昧人的勞碌使自己困乏， 連進城的路他也不知道。
ECCL|10|16|邦國啊，你的君王若年少， 你的群臣早晨宴樂， 你就有禍了！
ECCL|10|17|邦國啊，你的君王若是貴族之子， 你的群臣按時吃喝， 是為強身，不為酒醉， 你就有福了！
ECCL|10|18|因人懶惰，房頂塌下； 因人手懶，房屋滴漏。
ECCL|10|19|擺設宴席是為歡樂。 酒能使人快活， 錢能叫萬事應心。
ECCL|10|20|不可詛咒君王， 連起意也不可， 在臥室裏也不可詛咒富人； 因為空中的飛鳥必傳揚這聲音， 有翅膀的必述說這事。
ECCL|11|1|當將你的糧食撒在水面上， 因為日子久了，你必能得著它。
ECCL|11|2|將你所擁有的分給七人，或八人， 因為你不知道會有甚麼災禍臨到地上。
ECCL|11|3|雲若滿了雨，就必傾倒在地上。 樹向南倒，或向北倒， 樹倒在何處，就留在何處。
ECCL|11|4|看風的，必不撒種； 望雲的，必不收割。
ECCL|11|5|你不知道氣息如何進入孕婦的骨頭裏 ；照樣，造萬物之上帝的作為，你也無從得知。
ECCL|11|6|早晨要撒種，晚上也不要歇手，因為你不知道哪一樣發旺；前者或後者，或兩者都一樣好。
ECCL|11|7|光是甜美的，眼見日光是多麼好啊！
ECCL|11|8|人活多少年，就當快樂多少年，然而也當想到黑暗的日子；因為這樣的日子必多，所要來臨的全是虛空。
ECCL|11|9|年輕人哪，你在年少時當快樂；在年輕時使你的心歡暢，做你心所願做的，看你眼所愛看的；卻要知道，為這一切，上帝必審問你。
ECCL|11|10|所以，當從心中除掉愁煩，從肉體除去痛苦；因為年少和年輕之時，全是虛空。
ECCL|12|1|你趁著年輕、衰老的日子尚未來到，就是你所說，我毫無喜悅的那些歲月來臨之前，當記念造你的主。
ECCL|12|2|不要等到太陽、光明、月亮、星宿變為黑暗，雨後雲又返回；
ECCL|12|3|看守房屋的發顫，強壯的屈身，推磨的婦女因人少而停工，從窗戶往外看的眼光變為昏暗；
ECCL|12|4|街門關閉，推磨的聲音微小，鳥一叫，就驚醒，唱歌女子的聲音也都微弱；
ECCL|12|5|人怕高處，路上有驚慌；杏樹開花，蚱蜢成為重擔，慾望不再挑起；因為人歸他永遠的家，弔喪的在街上往來。
ECCL|12|6|不要等到銀鏈折斷 ，金罐破裂，瓶子在泉旁損壞，水輪在井口斷裂，
ECCL|12|7|塵土仍歸於地，像原來一樣，氣息仍歸於賜氣息的上帝。
ECCL|12|8|傳道者說：「虛空的虛空，全是虛空。」
ECCL|12|9|再者，傳道者因有智慧，將知識教導眾人；他思量，考察，並列舉出許多箴言。
ECCL|12|10|傳道者專心尋求可喜悅的言語，是憑正直寫的誠實話。
ECCL|12|11|智慧人的話語如同刺棒；這些嘉言好像釘穩的釘子，都是一個牧者所賜的。
ECCL|12|12|我兒，還有一點，你當受勸戒：著書多，沒有窮盡；讀書多，身體疲倦。
ECCL|12|13|這些事都已聽見了，結論就是：敬畏上帝，謹守他的誡命，這是人當盡的本分。
ECCL|12|14|因為人所做的事，連一切隱藏的事，無論是善是惡，上帝都必審問。
SONG|1|1|所羅門 的雅歌 。
SONG|1|2|願他用口與我親吻。 你的愛情比酒更美，
SONG|1|3|你的膏油馨香， 你的名如傾瀉而出的香膏， 所以童女都愛你。
SONG|1|4|願你吸引我跟隨你；讓我們快跑吧！ 王領我進入他的內室。 我們必因你歡喜快樂， 我們要思念你的愛情， 勝似思念美酒。 她們愛你是理所當然的。
SONG|1|5|耶路撒冷 的女子啊， 我雖然黑，卻是秀美， 如同 基達 的帳棚， 好像 所羅門 的幔子，
SONG|1|6|不要因太陽把我曬黑了就瞪著我。 我母親的兒子向我發怒， 他們使我看守葡萄園； 我自己的葡萄園我卻沒有看守。
SONG|1|7|我心所愛的啊，請告訴我， 你在何處牧羊？ 正午在何處使羊歇臥？ 我何必像蒙著臉的女子 在你同伴的羊群旁邊呢？
SONG|1|8|你這女子中最美麗的， 你若不知道， 只管跟隨羊群的腳蹤行， 在牧人的帳棚邊，牧放你的小山羊。
SONG|1|9|我的佳偶， 你好比法老戰車上的駿馬。
SONG|1|10|你的兩頰因髮辮而秀美， 你的頸項因珠串而華麗。
SONG|1|11|我們要為你編上金鏈，鑲上銀飾。
SONG|1|12|王正坐席的時候， 我的哪噠香膏散發香味。
SONG|1|13|我的良人好像一袋沒藥， 在我胸懷中。
SONG|1|14|我的良人好像一束鳳仙花， 在 隱‧基底 的葡萄園中。
SONG|1|15|看哪，我的佳偶，你真美麗！ 看哪，你真美麗！你的眼睛是鴿子。
SONG|1|16|看哪，我的良人，你多英俊可愛！ 讓我們以青草為床榻，
SONG|1|17|以香柏樹為房子的棟梁， 以松樹作屋頂的椽木。
SONG|2|1|我是 沙崙 的玫瑰花， 是谷中的百合花。
SONG|2|2|我的佳偶在女子中， 好像荊棘裏的百合花。
SONG|2|3|我的良人在男子中， 如同蘋果樹在樹林裏。 我歡歡喜喜坐在他的蔭下， 嘗他果子的滋味，覺得甘甜。
SONG|2|4|他領我進入宴會廳， 為我插上愛的旗幟。
SONG|2|5|請你們用葡萄餅增補我力， 以蘋果暢快我的心， 因我為愛而生病。
SONG|2|6|他的左手在我頭下， 他的右手將我環抱。
SONG|2|7|耶路撒冷 的女子啊， 我指著羚羊或田野的母鹿囑咐你們， 不要喚醒，不要挑動愛情，等它自發。
SONG|2|8|聽啊！我良人的聲音， 看哪！他穿山越嶺而來。
SONG|2|9|我的良人像羚羊，像小鹿。 看哪，他站在我們的牆壁邊， 從窗戶往裏觀看， 從窗格子往裏窺探。
SONG|2|10|我的良人對我說： 「我的佳偶，起來！ 我的美人，與我同去！
SONG|2|11|看哪，因為冬天已逝， 雨水止住，已經過去了。
SONG|2|12|地上百花開放， 歌唱的時候到了， 斑鳩的聲音在我們境內也聽見了。
SONG|2|13|無花果樹的果子漸漸成熟， 葡萄樹開花，散發香氣。 我的佳偶，起來！ 我的美人，與我同去！
SONG|2|14|我的鴿子啊，你在磐石穴中， 在陡巖的隱密處。 求你容我得見你的面貌， 求你容我得聽你的聲音； 因你的聲音悅耳， 你的容貌秀美。
SONG|2|15|請為我們擒拿狐狸， 就是毀壞葡萄園的小狐狸， 我們的葡萄正在開花。」
SONG|2|16|我的良人屬我，我也屬他， 他在百合花中放牧。
SONG|2|17|我的良人哪， 等到天起涼風、 日影飛去的時候， 願你歸回，像羚羊， 像小鹿，在崎嶇的山 上。
SONG|3|1|我夜間躺臥在床上， 尋找我心所愛的； 我尋找他，卻尋不著。
SONG|3|2|「我要起來，繞行城中， 在街市上，在廣場上， 尋找我心所愛的。」 我尋找他，卻尋不著。
SONG|3|3|城中巡邏的守衛遇見我， 「你們看見我心所愛的沒有？」
SONG|3|4|我剛離開他們，就遇見我心所愛的。 我拉住他，不放他走， 領他進入我母親的家， 到懷我者的內室。
SONG|3|5|耶路撒冷 的女子啊， 我指著羚羊或田野的母鹿囑咐你們， 不要喚醒，不要挑動愛情，等它自發。
SONG|3|6|那如煙柱從曠野上來， 薰了沒藥、乳香，撲上商人各樣香粉的是誰呢？
SONG|3|7|看哪，是 所羅門 的轎， 周圍有六十個勇士， 都是 以色列 中的勇士。
SONG|3|8|他們的手都持刀，善於爭戰， 各人腰間佩刀，防備夜間恐怖的攻擊。
SONG|3|9|所羅門 王用 黎巴嫩 木 為自己製作轎子。
SONG|3|10|轎柱是用銀做的， 轎底是用金做的， 坐墊是紫色的， 其中所鋪的是 耶路撒冷 女子的愛情。
SONG|3|11|錫安的女子啊， 你們要出去觀看 所羅門 王！ 他頭戴冠冕，就是在他結婚當天 心中喜樂的時候，他母親給他戴上的。
SONG|4|1|看哪，我的佳偶，你真美麗！看哪，你真美麗！ 你的眼睛在面紗後好像鴿子。 你的頭髮如同一群山羊，從 基列山 下來。
SONG|4|2|你的牙齒如新剪毛的一群母羊，洗淨之後走上來， 它們成對，沒有一顆是單獨的。
SONG|4|3|你的唇好像一條朱紅線， 你的嘴秀美。 你的鬢角在面紗後， 如同迸開的石榴。
SONG|4|4|你的頸項猶如 大衛 為收藏軍器而造的高塔， 其上懸掛一千個盾牌， 都是勇士的盾牌。
SONG|4|5|你的兩乳好像百合花中吃草的一對小鹿， 是母鹿雙生的。
SONG|4|6|我要往沒藥山和乳香岡去， 直到天起涼風、 日影飛去的時候。
SONG|4|7|我的佳偶，你全然美麗， 毫無瑕疵！
SONG|4|8|我的新娘，請你與我一同離開 黎巴嫩 ， 與我一同離開 黎巴嫩 。 從 亞瑪拿 山巔， 從 示尼珥 ，就是 黑門山 頂， 從獅子的洞， 從豹子的山往下觀看。
SONG|4|9|我的妹子，我的新娘， 你奪了我的心。 你明眸一瞥， 你頸項的鏈子， 奪了我的心！
SONG|4|10|我的妹子，我的新娘， 你的愛情 何其美！ 你的愛情比酒甜美！ 你膏油的馨香勝過一切香料！
SONG|4|11|我的新娘，你的唇滴下蜂蜜， 你的舌下有蜜，有奶。 你衣服的香氣宛如 黎巴嫩 的芬芳。
SONG|4|12|我的妹子，我的新娘 是上鎖的園子， 是禁閉的園子 ， 是封閉的泉源。
SONG|4|13|你園內所種的結了石榴， 有佳美的果子， 並鳳仙花與哪噠樹。
SONG|4|14|有哪噠和番紅花， 香菖蒲和桂樹， 並各樣乳香木、沒藥、沉香， 與一切上等的香料。
SONG|4|15|你是園中的泉，活水的井， 是從 黎巴嫩 湧流而下的溪水。
SONG|4|16|北風啊，興起！ 南風啊，吹來！ 吹在我的園內， 使其中的香氣散發出來。 願我的良人進入自己園裏， 吃他佳美的果子。
SONG|5|1|我的妹子，我的新娘， 我進入我的園中， 採了我的沒藥和香料， 吃了我的蜂房和蜂蜜， 喝了我的酒和奶。 我的朋友，請吃！ 我親愛的，請喝，多多地喝！
SONG|5|2|我身躺臥，我心卻醒。 這是我良人的聲音； 他敲門： 「我的妹子，我的佳偶， 我的鴿子，我完美的人兒， 請你為我開門； 因我的頭沾滿露水， 我的髮被夜露滴濕。」
SONG|5|3|我脫了衣裳，怎能再穿上呢？ 我洗了腳，怎可再弄髒呢？
SONG|5|4|我的良人從門縫裏伸進他的手， 我便因他動了心。
SONG|5|5|我起來，要為我的良人開門。 我的兩手滴下沒藥， 我的指頭有沒藥汁滴在門閂上。
SONG|5|6|我為我的良人開了門， 我的良人卻已轉身走了。 他說話的時候，我魂不守舍。 我尋找他，竟尋不著， 我呼叫他，他卻不回答。
SONG|5|7|城中巡邏的守衛遇見我， 打了我，傷了我， 看守城牆的人奪去我的披肩。
SONG|5|8|耶路撒冷 的女子啊，我囑咐你們： 若遇見我的良人， 要告訴他，我為愛而生病。
SONG|5|9|你這女子中最美麗的， 你的良人有甚麼勝過別的良人呢？ 你的良人有甚麼勝過別的良人， 使你這樣囑咐我們？
SONG|5|10|我的良人紅潤發亮， 超乎萬人之上。
SONG|5|11|他的頭像千足的純金， 他的髮綹卷曲，黑如烏鴉。
SONG|5|12|他的眼如溪水旁的鴿子， 沐浴在奶中，安得合式 。
SONG|5|13|他的兩頰如香花園， 如香草臺 ； 他的嘴唇像百合花， 滴下沒藥汁。
SONG|5|14|他的雙手宛如金條， 鑲嵌水蒼玉； 他的身體如同雕刻的象牙， 周圍鑲嵌藍寶石。
SONG|5|15|他的腿好比白玉石柱， 安在精金座上； 他的容貌如 黎巴嫩 ， 佳美如香柏樹。
SONG|5|16|他的口甘甜， 他全然可愛。 耶路撒冷 的女子啊， 這是我的良人， 這是我的朋友。
SONG|6|1|你這女子中最美麗的， 你的良人往何處去？ 你的良人轉向何處去了？ 我們好與你同去尋找他。
SONG|6|2|我的良人進入自己園中， 到香花園， 在園內放牧， 採百合花。
SONG|6|3|我屬我的良人， 我的良人屬我； 他在百合花中放牧。
SONG|6|4|我的佳偶啊，你美麗如 得撒 ， 秀美如 耶路撒冷 ， 威武如展開旌旗的軍隊。
SONG|6|5|求你轉開眼睛不要看我， 因你的眼睛使我慌亂。 你的頭髮如同一群山羊，從 基列山 下來。
SONG|6|6|你的牙齒如一群母羊，洗淨之後走上來， 它們成對，沒有一顆是單獨的。
SONG|6|7|你的鬢角在面紗後， 如同迸開的石榴。
SONG|6|8|雖有六十王后、八十妃嬪， 並有無數的童女。
SONG|6|9|她是我獨一的鴿子、我完美的人兒， 是她母親獨生的， 是生養她的所寵愛的。 女子見了都稱她有福， 王后妃嬪見了也讚美她。
SONG|6|10|那俯視如晨曦、 美麗如月亮、皎潔如太陽、 威武如展開旌旗軍隊的是誰呢？
SONG|6|11|我下到堅果園， 要看谷中青翠的植物， 要看葡萄可曾發芽， 石榴可曾放蕊；
SONG|6|12|不知不覺， 我彷彿坐在我百姓高官 的戰車中。
SONG|6|13|回來，回來， 書拉密 的女子； 回來，回來，我們要看你。 你們為何要觀看 書拉密 的女子， 像觀看兩隊人馬在跳舞 呢？
SONG|7|1|尊貴的女子啊，你的腳在鞋中何等秀美！ 你的大腿圓潤，好像美玉， 是巧匠的手做成的。
SONG|7|2|你的肚臍如圓杯， 不缺調和的酒。 你的肚子如一堆麥子， 周圍有百合花。
SONG|7|3|你的兩乳好像一對小鹿， 是母鹿雙生的。
SONG|7|4|你的頸項如象牙塔， 你的眼睛像 希實本 、 巴特‧拉併 門旁的水池， 你的鼻子彷彿朝向 大馬士革 的 黎巴嫩 塔。
SONG|7|5|你的頭在你身上好像 迦密山 ， 你頭上的髮呈紫色， 王被這髮綹繫住了。
SONG|7|6|我親愛的，喜樂的女子啊， 你何等美麗！何等令人喜悅！
SONG|7|7|你的身材好像棕樹， 你的兩乳如同纍纍的果實。
SONG|7|8|我說：我要爬上棕樹，抓住枝子。 願你的兩乳好像葡萄纍纍， 願你鼻子的香氣如蘋果；
SONG|7|9|你的上顎如美酒， 直流入我良人的口裏， 流入沉睡者的口中 。
SONG|7|10|我屬我的良人， 他也戀慕我。
SONG|7|11|來吧！我的良人， 讓我們往田間去， 在村莊住宿。
SONG|7|12|早晨讓我們起來往葡萄園去， 看葡萄樹發芽沒有， 花開了沒有， 石榴放蕊沒有， 在那裏我要將我的愛情給你。
SONG|7|13|曼陀羅草 散發香味， 在我們的門內有各樣新陳佳美的果子； 我的良人，這都是我為你保存的。
SONG|8|1|惟願你像我的兄弟， 像吃我母親奶的兄弟。 我在外頭遇見你就與你親吻， 誰也不輕看我。
SONG|8|2|我必引導你， 領你進入我母親的家， 她必教導我， 我必使你喝石榴汁釀的香酒。
SONG|8|3|他的左手在我頭下， 他的右手將我環抱。
SONG|8|4|耶路撒冷 的女子啊， 我囑咐你們， 不要喚醒、不要挑動愛情，等它自發。
SONG|8|5|那靠著良人從曠野上來的是誰呢？ 在蘋果樹下，我叫醒了你； 在那裏，你母親曾為了生你而陣痛， 在那裏，生你的為你陣痛。
SONG|8|6|求你將我放在你心上如印記， 帶在你臂上如戳記。 因為愛情如死之堅強， 熱戀如陰間之牢固， 所發的光是火焰的光， 是極其猛烈的火焰 。
SONG|8|7|愛情，眾水不能熄滅， 江河也不能淹沒。 若有人拿家中所有的財寶要換愛情， 就全被藐視。
SONG|8|8|我們有一小妹， 她還沒有乳房， 人來提親的日子， 我們當為她怎麼辦呢？
SONG|8|9|她若是牆， 我們要在其上建造銀塔； 她若是門， 我們要用香柏木板圍護她。
SONG|8|10|我是牆， 我的兩乳像塔。 那時，我在他眼中是找到平安的人。
SONG|8|11|所羅門 在 巴力‧哈們 有一葡萄園， 他將這葡萄園租給看守的人， 每人為其中的果子要交一千銀子。
SONG|8|12|我有屬自己的葡萄園。 所羅門 哪，一千歸你， 兩百歸看守果子的人。
SONG|8|13|你這住在園中的， 同伴都要聽你的聲音， 求你使我也得以聽見。
SONG|8|14|我的良人哪，求你快來！ 像羚羊，像小鹿，在香草山上。
ISA|1|1|當 烏西雅 、 約坦 、 亞哈斯 、 希西家 作 猶大 王的時候， 亞摩斯 的兒子 以賽亞 見異象，論到 猶大 和 耶路撒冷 。
ISA|1|2|天哪，要聽！地啊，側耳而聽！ 因為耶和華說： 「我養育兒女，將他們養大， 他們竟悖逆我。
ISA|1|3|牛認識主人， 驢認識主人的槽； 以色列 卻不認識， 我的民卻不明白。」
ISA|1|4|禍哉！犯罪的國民， 擔著罪孽的百姓， 行惡的族類， 敗壞的兒女！ 他們離棄耶和華， 藐視 以色列 的聖者， 背向他，與他疏遠。
ISA|1|5|你們為甚麼屢次悖逆，繼續受責打呢？ 你們已經滿頭疼痛， 全心發昏；
ISA|1|6|從腳掌到頭頂， 沒有一處是完好的， 盡是創傷、瘀青，與流血的傷口， 未曾擠淨，未曾包紮， 也沒有用膏滋潤。
ISA|1|7|你們的土地荒蕪， 城鎮被火燒燬； 你們的田地在你們眼前被陌生人侵吞， 既被陌生人傾覆，就成為荒蕪 。
ISA|1|8|僅存的 錫安 ， 好似葡萄園的草棚， 如瓜田中的茅屋， 又如被圍困的城。
ISA|1|9|若不是萬軍之耶和華為我們留下一些倖存者， 我們早已變成 所多瑪 ，像 蛾摩拉 一樣了。
ISA|1|10|所多瑪 的官長啊， 你們要聽耶和華的言語！ 蛾摩拉 的百姓啊， 要側耳聽我們上帝的教誨！
ISA|1|11|耶和華說： 「你們許多的祭物於我何益呢？ 公綿羊的燔祭和肥畜的油脂， 我已經膩煩了； 公牛、羔羊、公山羊的血， 我都不喜悅。
ISA|1|12|「你們來朝見我， 誰向你們的手要求這些， 使你們踐踏我的院宇呢？
ISA|1|13|不要再獻無謂的供物了， 香是我所憎惡的。 我不能容忍行惡又守嚴肅會： 初一、安息日和召集的大會。
ISA|1|14|你們的初一和節期，我心裏恨惡， 它們成了我的重擔， 擔當這些，令我厭煩。
ISA|1|15|你們舉手禱告，我必遮眼不看， 就算你們多多祈禱，我也不聽； 你們的手沾滿了血。
ISA|1|16|你們要洗滌、自潔， 從我眼前除掉惡行； 要停止作惡，
ISA|1|17|學習行善， 尋求公平， 幫助受欺壓的 ， 替孤兒伸冤， 為寡婦辯護。」
ISA|1|18|耶和華說： 「來吧，我們彼此辯論。 你們的罪雖像硃紅，必變成雪白； 雖紅如丹顏，必白如羊毛。
ISA|1|19|你們若甘心聽從， 必吃地上的美物；
ISA|1|20|若不聽從，反倒悖逆， 必被刀劍吞滅； 這是耶和華親口說的。」
ISA|1|21|忠信的城竟然變為妓女！ 從前充滿了公平， 公義居在其中， 現今卻有兇手居住。
ISA|1|22|你的銀子變為渣滓， 你的酒用水沖淡。
ISA|1|23|你的官長悖逆， 與盜賊為伍， 全都喜愛賄賂， 追求贓物； 他們不為孤兒伸冤， 寡婦的案件也呈不到他們面前。
ISA|1|24|因此，主－萬軍之耶和華、 以色列 的大能者說： 「唉！我要向我的對頭雪恨， 向我的敵人報仇。
ISA|1|25|我必反手對付你， 如鹼煉淨你的渣滓， 除盡你的雜質。
ISA|1|26|我必回復你的審判官，像起初一樣， 回復你的謀士，如起先一般。 然後，你必稱為公義之城， 忠信之邑。」
ISA|1|27|錫安 必因公平得蒙救贖， 其中歸正的人必因公義得蒙救贖。
ISA|1|28|但悖逆的和犯罪的必一同敗亡， 離棄耶和華的必致消滅。
ISA|1|29|那等人必因所喜愛的聖樹抱愧； 你們必因所選擇的園子 蒙羞，
ISA|1|30|因為你們必如葉子枯乾的橡樹， 如無水的園子。
ISA|1|31|有權勢的必如麻線， 他的作為好像火花， 都要一同焚燒，無人撲滅。
ISA|2|1|亞摩斯 的兒子 以賽亞 所見，有關 猶大 和 耶路撒冷 的事。
ISA|2|2|末後的日子，耶和華殿的山必堅立， 超乎諸山，高舉過於萬嶺； 萬國都要流歸這山。
ISA|2|3|必有許多民族前往，說： 「來吧，我們登耶和華的山， 到 雅各 上帝的殿。 他必將他的道教導我們， 我們也要行他的路。」 因為教誨必出於 錫安 ， 耶和華的言語必出於 耶路撒冷 。
ISA|2|4|他必在萬國中施行審判， 為許多民族斷定是非。 他們要將刀打成犁頭， 把槍打成鐮刀； 這國不舉刀攻擊那國， 他們也不再學習戰事。
ISA|2|5|雅各 家啊， 來吧！讓我們在耶和華的光明中行走。
ISA|2|6|你離棄了你的百姓 雅各 家， 因為他們充滿了東方的習俗 ， 又像 非利士 人一樣觀星象， 並與外邦人擊掌。
ISA|2|7|他們的國滿了金銀， 財寶也無窮； 他們的地滿了馬匹， 戰車也無數。
ISA|2|8|他們的地滿了偶像； 他們跪拜自己手所造的， 就是自己手指所做的。
ISA|2|9|有人屈膝， 有人下跪； 所以，不要饒恕他們。
ISA|2|10|當進入磐石，藏在土中， 躲避耶和華的驚嚇和他威嚴的榮光。
ISA|2|11|到那日，眼目高傲的必降卑， 狂妄的人必屈膝； 惟獨耶和華被尊崇。
ISA|2|12|因萬軍之耶和華的一個日子 要臨到所有驕傲狂妄的， 臨到一切自高的， 使他們降為卑；
ISA|2|13|臨到 黎巴嫩 高大的香柏樹、 巴珊 的橡樹，
ISA|2|14|臨到一切高山、 一切峻嶺，
ISA|2|15|臨到一切碉堡、 一切堅固的城牆，
ISA|2|16|臨到 他施 一切的船隻、 一切華麗的船艇。
ISA|2|17|人的驕傲必屈膝， 人的狂妄必降卑； 在那日，惟獨耶和華被尊崇，
ISA|2|18|偶像必全然廢棄。
ISA|2|19|耶和華興起使地大震動的時候， 人就進入石洞和土穴裏， 躲避耶和華的驚嚇和他威嚴的榮光。
ISA|2|20|到那日，人必將造來敬拜的金偶像、銀偶像 拋給田鼠和蝙蝠。
ISA|2|21|耶和華興起使地大震動的時候， 人就進入磐縫和巖隙裏， 躲避耶和華的驚嚇和他威嚴的榮光。
ISA|2|22|你們不要倚靠世人， 他只不過鼻孔裏有氣息， 算得了甚麼呢？
ISA|3|1|看哪，主－萬軍之耶和華要從 耶路撒冷 和 猶大 除掉眾人所倚靠的，所仰賴的， 就是所倚靠的糧，所仰賴的水；
ISA|3|2|除掉勇士和戰士， 審判官和先知， 占卜的和長老，
ISA|3|3|除掉五十夫長和顯要、 謀士和巧匠， 以及擅長法術的人。
ISA|3|4|我必使孩童作他們的領袖， 幼兒管轄他們。
ISA|3|5|百姓要彼此欺壓， 各人欺壓鄰舍； 青年要侮慢老人， 卑賤的要侮慢尊貴的。
ISA|3|6|人在父家拉住自己的兄弟： 「你有外衣，來作我們的官長， 讓這些敗壞的事歸於你的手下吧！」
ISA|3|7|那時，他必揚聲說： 「我不作醫治你們的人； 我家裏沒有糧食，也沒有衣服， 你們不可立我作百姓的官長。」
ISA|3|8|耶路撒冷 敗落， 猶大 傾倒； 因為他們的舌頭和行為與耶和華相悖， 無視於他榮光的眼目。
ISA|3|9|他們的臉色證明自己不正， 他們述說自己像 所多瑪 一樣的罪惡，毫不隱瞞。 他們有禍了！因為作惡自害。
ISA|3|10|你們要對義人說，他是有福的， 因為他必吃自己行為所結的果實。
ISA|3|11|惡人有禍了！他必遭災難！ 因為他要按自己手所做的受報應。
ISA|3|12|至於我的百姓， 統治者剝削你們， 放高利貸的人管轄你們 。 我的百姓啊，引導你的使你走錯， 並毀壞你所行的道路。
ISA|3|13|耶和華興起訴訟， 站著審判萬民。
ISA|3|14|耶和華必審問他國中的長老和領袖： 「你們，你們摧毀葡萄園， 搶奪困苦人，囤積在你們家中。
ISA|3|15|你們為何壓碎我的百姓， 碾磨困苦人的臉呢？」 這是萬軍之主耶和華說的。
ISA|3|16|耶和華說： 因為 錫安 狂傲， 行走挺項，賣弄眼目， 俏步徐行，腳下玎璫，
ISA|3|17|主必使 錫安 頭頂長瘡， 耶和華又暴露其下體。
ISA|3|18|到那日，主必除掉華美的足飾、額帶、月牙圈、
ISA|3|19|耳環、手鐲、面紗、
ISA|3|20|頭巾、足鏈、華帶、香盒、符囊、
ISA|3|21|戒指、鼻環、
ISA|3|22|禮服、外套、披肩、皮包、
ISA|3|23|手鏡、細麻衣、頭飾、紗巾。
ISA|3|24|必有腐爛代替馨香， 繩子代替腰帶， 光禿代替美髮， 麻衣繫腰代替華服， 烙痕代替美貌。
ISA|3|25|你的男丁必倒在刀下， 你的勇士必死在陣上。
ISA|3|26|錫安 的城門必悲傷、哀號； 它必荒涼，坐在地上。
ISA|4|1|在那日，七個女人必拉住一個男人，說：「我們吃自己的食物，穿自己的衣服，但求你允許我們歸你名下，除掉我們的羞恥。」
ISA|4|2|在那日，耶和華的苗必華美尊榮，地的出產必成為倖存的 以色列 民的驕傲和光榮。
ISA|4|3|主以公平的靈和焚燒的靈洗淨 錫安 居民 的污穢，又除淨在 耶路撒冷 流人血的罪。那時，剩在 錫安 、留在 耶路撒冷 的，就是一切住 耶路撒冷 、在生命冊上記名的，必稱為聖。
ISA|4|4|
ISA|4|5|耶和華必在整座 錫安山 ，在會眾之上，白天造雲，黑夜發出煙和火焰的光，因為在一切榮耀之上必有華蓋；
ISA|4|6|這要作為棚子，白天可以遮蔭避暑，暴風雨侵襲時，可作藏身處和避難所。
ISA|5|1|我要為我親愛的唱歌， 我所愛的、他的葡萄園之歌。 我親愛的有葡萄園 在肥沃的山岡上。
ISA|5|2|他刨挖園子，清除石頭， 栽種上等的葡萄樹， 在園中蓋了一座樓， 又鑿出酒池； 指望它結葡萄， 反倒結了野葡萄。
ISA|5|3|耶路撒冷 的居民和 猶大 人哪， 現在，請你們在我與我的葡萄園之間斷定是非。
ISA|5|4|我為我葡萄園所做的之外， 還有甚麼可做的呢？ 我指望它結葡萄， 怎麼倒結了野葡萄呢？
ISA|5|5|現在我告訴你們， 我要向我的葡萄園怎麼做。 我必撤去籬笆，使它被燒燬； 拆毀圍牆，使它被踐踏。
ISA|5|6|我必使它荒廢，不再修剪， 不再鋤草，任荊棘蒺藜生長； 我也必吩咐密雲， 不再降雨在其上。
ISA|5|7|萬軍之耶和華的葡萄園就是 以色列 家； 他所喜愛的樹就是 猶大 人。 他指望公平， 看哪，卻有流血； 指望公義， 看哪，卻有冤聲。
ISA|5|8|禍哉！你們以房接房， 以地連地， 以致不留餘地， 只顧自己獨居境內。
ISA|5|9|我耳聞萬軍之耶和華說： 「許多房屋必然荒廢； 宏偉華麗，無人居住。
ISA|5|10|十畝 的葡萄園只釀出一罷特的酒， 一賀梅珥的穀種只結一伊法糧食。」
ISA|5|11|禍哉！那些清晨早起，追尋烈酒， 因酒狂熱，流連到深夜的人，
ISA|5|12|他們在宴席上 彈琴，鼓瑟，擊鼓，吹笛，飲酒， 卻不留意耶和華的作為， 也不留心他手所做的。
ISA|5|13|所以，我的百姓因無知就被擄去； 尊貴的人甚是飢餓， 平民也極其乾渴。
ISA|5|14|因此，陰間胃口 大開， 張開無限量的口； 令 耶路撒冷 的貴族與平民、狂歡的與作樂的人 都掉落其中。
ISA|5|15|人為之屈膝， 人就降為卑； 高傲的眼目也降為卑。
ISA|5|16|惟有萬軍之耶和華因公平顯為崇高， 神聖的上帝因公義顯為聖。
ISA|5|17|羔羊必來吃草，如同在自己的草場； 在富有人的廢墟，流浪的牲畜也來吃 。
ISA|5|18|禍哉！那些以虛假的繩子牽引罪孽， 以套車的繩索緊拉罪惡的人。
ISA|5|19|他們說： 「任 以色列 的聖者急速前行，快快成就他的作為， 好讓我們看看； 任他的籌算臨近成就， 好使我們知道。」
ISA|5|20|禍哉！那些稱惡為善，稱善為惡， 以暗為光，以光為暗， 以苦為甜，以甜為苦的人。
ISA|5|21|禍哉！那些在自己眼中有智慧， 在自己面前有通達的人。
ISA|5|22|禍哉！那些以飲酒稱雄， 以調烈酒稱霸的人。
ISA|5|23|他們因受賄賂，就稱惡人為義， 將義人的義奪去。
ISA|5|24|火苗怎樣吞滅碎秸， 乾草怎樣落在火焰之中， 照樣，他們的根必然腐朽， 他們的花像灰塵揚起； 因為他們厭棄萬軍之耶和華的教誨， 藐視 以色列 聖者的言語。
ISA|5|25|因此，耶和華的怒氣向他的百姓發作。 他伸手攻擊他們，山嶺就震動； 他們的屍首在街市上好像糞土。 雖然如此，他的怒氣並未轉消， 他的手依然伸出。
ISA|5|26|他必豎立大旗，召集遠方的國民， 把他們從地極叫來。 看哪，他們必急速奔來，
ISA|5|27|其中沒有疲倦的，絆跌的； 沒有打盹的，睡覺的； 腰帶並不放鬆， 鞋帶也不拉斷。
ISA|5|28|他們的箭銳利， 弓也上了弦； 馬蹄如堅石， 車輪像旋風。
ISA|5|29|他們要吼叫，像母獅， 咆哮，像少壯獅子； 他們要咆哮，抓取獵物， 穩穩叼走，無人能救回。
ISA|5|30|那日，他們要向 以色列 人咆哮， 像海浪澎湃； 人若望地，看哪，只有黑暗與禍患， 光明因密雲而變黑暗。
ISA|6|1|當 烏西雅 王崩的那年，我看見主坐在高高的寶座上。他的衣裳下襬遮滿聖殿。
ISA|6|2|上有撒拉弗侍立，各有六個翅膀：兩個翅膀遮臉，兩個翅膀遮腳，兩個翅膀飛翔，
ISA|6|3|彼此呼喊說： 「聖哉！聖哉！聖哉！萬軍之耶和華； 他的榮光遍滿全地！」
ISA|6|4|因呼喊者的聲音，門檻的根基震動，殿裏充滿了煙雲。
ISA|6|5|那時我說：「禍哉！我滅亡了！因為我是嘴唇不潔的人，住在嘴唇不潔的民中，又因我親眼看見大君王－萬軍之耶和華。」
ISA|6|6|有一撒拉弗向我飛來，手裏拿著燒紅的炭，是用火鉗從壇上取下來的，
ISA|6|7|用炭沾我的口，說：「看哪，這炭沾了你的嘴唇，你的罪孽便除掉，你的罪惡就赦免了。」
ISA|6|8|我聽見主的聲音說：「我可以差遣誰呢？誰肯為我們去呢？」我說：「我在這裏，請差遣我！」
ISA|6|9|他說：「你去告訴這百姓說： 『你們聽了又聽，卻不明白； 看了又看，卻不曉得。』
ISA|6|10|要使這百姓心蒙油脂， 耳朵發沉， 眼睛昏花； 恐怕他們眼睛看見， 耳朵聽見， 心裏明白， 回轉過來，就得醫治。」
ISA|6|11|我就說：「主啊，這到幾時為止呢？」他說： 「直到城鎮荒涼，無人居住， 房屋空無一人，土地極其荒蕪；
ISA|6|12|耶和華將人遷到遠方， 國內被撇棄的土地很多。
ISA|6|13|國內剩下的人若還有十分之一， 也必被吞滅。 然而如同大樹與橡樹，雖被砍伐， 殘幹卻仍存留， 聖潔的苗裔是它的殘幹。」
ISA|7|1|烏西雅 的孫子， 約坦 的兒子， 猶大 王 亞哈斯 在位的時候， 亞蘭 王 利汛 和 利瑪利 的兒子 以色列 王 比加 上來攻打 耶路撒冷 ，卻不能攻取。
ISA|7|2|有人告訴 大衛 家說：「 亞蘭 與 以法蓮 已經結盟。」王的心和百姓的心就都顫動，好像林中的樹被風吹動一樣。
ISA|7|3|耶和華對 以賽亞 說：「你和你的兒子 施亞‧雅述 要出去，到 上池 的水溝盡頭，往漂布地的大路上，迎見 亞哈斯 ，
ISA|7|4|對他說：『你要謹慎，要鎮定，不要害怕，不要因 利汛 和 亞蘭 ，以及 利瑪利 的兒子這兩個冒煙火把的頭所發的烈怒而心裏膽怯。
ISA|7|5|因為 亞蘭 、 以法蓮 ，和 利瑪利 的兒子設惡謀要害你，說：
ISA|7|6|我們要上去攻擊 猶大 ，擾亂它，攻破它來歸我們，在其中立 他比勒 的兒子為王。
ISA|7|7|主耶和華如此說： 這事必站立不住， 也不得成就。
ISA|7|8|因為 亞蘭 的首都是 大馬士革 ， 大馬士革 的領袖是 利汛 ； 六十五年之內， 以法蓮 必然國破族亡，
ISA|7|9|以法蓮 的首都是 撒瑪利亞 ； 撒瑪利亞 的領袖是 利瑪利 的兒子。 你們若是不信， 必站立不穩。』」
ISA|7|10|耶和華又吩咐 亞哈斯 ：
ISA|7|11|「你向耶和華－你的上帝求一個預兆：在陰間的深淵，或往上的高處。」
ISA|7|12|但 亞哈斯 說：「我不求；我不試探耶和華。」
ISA|7|13|以賽亞 說：「聽啊， 大衛 家！你們使人厭煩豈算小事，還要使我的上帝厭煩嗎？
ISA|7|14|因此，主自己要給你們一個預兆，看哪，必有童女懷孕生子，給他起名叫 以馬內利 。
ISA|7|15|到他曉得棄惡擇善的時候，他必吃乳酪與蜂蜜。
ISA|7|16|因為在這孩子還不曉得棄惡擇善之先，你所憎惡的那兩個王的土地必被撇棄。
ISA|7|17|耶和華必使 亞述 王臨到你和你的百姓，並你的父家，自從 以法蓮 脫離 猶大 的時候，未曾有過這樣的日子。
ISA|7|18|「那時，耶和華要呼叫，召來 埃及 江河源頭的蒼蠅和 亞述 地的蜂；
ISA|7|19|牠們都必飛來，停在陡峭的谷中、巖石縫裏、一切荊棘叢中和片片草場上。
ISA|7|20|「那時，主必用 大河 外雇來的剃刀，就是 亞述 王，剃去你的頭髮和腳毛，並要剃淨你的鬍鬚。
ISA|7|21|「那時，每一個人要養活一頭母牛犢和兩隻母羊；
ISA|7|22|因為奶量充足，他就有乳酪可吃，國內剩餘的人也都能吃乳酪與蜂蜜。
ISA|7|23|「那時，凡種一千棵葡萄樹、價值一千銀子的地方，必長出荊棘和蒺藜。
ISA|7|24|人到那裏去，必帶弓箭，因為遍地長滿了荊棘和蒺藜。
ISA|7|25|所有鋤頭刨過的山地，你因懼怕荊棘和蒺藜，不敢到那裏去；只能作放牛之處，羊群踐踏之地。」
ISA|8|1|耶和華對我說：「你取一塊大板子，拿人的筆 ，寫上『瑪黑珥‧沙拉勒‧哈施‧罷斯』 。
ISA|8|2|我 要用可靠的證人， 烏利亞 祭司和 耶比利家 的兒子 撒迦利亞 為我作證。」
ISA|8|3|我親近女先知 ；她就懷孕生子，耶和華對我說：「給他起名叫 瑪黑珥‧沙拉勒‧哈施‧罷斯 ；
ISA|8|4|因為在這孩子還不曉得叫爸爸媽媽以前， 大馬士革 的財寶和 撒瑪利亞 的擄物必被 亞述 王掠奪一空。」
ISA|8|5|耶和華又吩咐我：
ISA|8|6|「這百姓既厭棄 西羅亞 緩流的水，喜歡 利汛 以及 利瑪利 的兒子，
ISA|8|7|因此，看哪，主必使 亞述 王和他的威勢如 大河 翻騰洶湧的水上漲，蓋過他們，必上漲超過一切水道，漲過兩岸，
ISA|8|8|必沖入 猶大 ，漲溢氾濫，直到頸項。他展開翅膀，遮蔽你的全地。 以馬內利 啊！」
ISA|8|9|萬民哪，任憑你們行惡 ，終必毀滅； 遠方的眾人哪，當側耳而聽！ 任憑你們束腰，終必毀滅； 你們束起腰來，終必毀滅。
ISA|8|10|任憑你們籌算甚麼，終必無效； 不管你們講定甚麼，總不成立； 因為上帝與我們同在。
ISA|8|11|耶和華以大能的手訓誡我不可行 這百姓所行的道，對我這樣說：
ISA|8|12|「這百姓說同謀背叛的，你們不要說同謀背叛。他們所怕的，你們不要怕，也不要畏懼；
ISA|8|13|但要尊萬軍之耶和華為聖，他才是你們所當怕的，所當畏懼的。
ISA|8|14|他必作為聖所，卻向 以色列 的兩家成為絆腳的石頭，使人跌倒的磐石；作 耶路撒冷 居民的羅網和圈套。
ISA|8|15|許多人在其上絆倒，他們跌倒，甚至跌傷，並且落入陷阱，被抓住了。」
ISA|8|16|你要捲起律法書，在我門徒中間封住教誨。
ISA|8|17|我要等候那轉臉不顧 雅各 家的耶和華，也要仰望他。
ISA|8|18|看哪，我與耶和華所賜給我的兒女成了 以色列 的預兆和奇蹟，這是從住在 錫安山 萬軍之耶和華來的。
ISA|8|19|有人對你們說：「當求問招魂的與行巫術的，他們唧唧喳喳，念念有詞。」然而，百姓不當求問自己的上帝嗎？豈可為活人求問死人呢？
ISA|8|20|當以教誨和律法書為準；人所說的若不與此相符，必沒有黎明。
ISA|8|21|他必經過這地，遇艱難，受飢餓；飢餓的時候，心中焦躁，咒罵自己的君王和上帝。他仰觀上天，
ISA|8|22|俯察下地，看哪，盡是艱難、黑暗和駭人的昏暗。他必被趕入幽暗中去。
ISA|9|1|但那受過痛苦的必不再見幽暗。 從前上帝使 西布倫 地和 拿弗他利 地被藐視，末後卻使這沿海的路， 約旦河 東，外邦人居住的 加利利 地得榮耀。
ISA|9|2|在黑暗中行走的百姓看見了大光； 住在死蔭之地的人有光照耀他們。
ISA|9|3|你使這國民眾多 ， 使他們喜樂大增； 他們在你面前歡喜， 好像收割時的歡喜， 又像人分戰利品那樣的快樂。
ISA|9|4|因為他們所負的重軛 和肩頭上的杖， 並欺壓者的棍， 你都已經折斷， 如同在 米甸 的日子一般。
ISA|9|5|戰士在戰亂中所穿的靴子， 以及那滾在血中的衣服， 都必當作柴火燃燒。
ISA|9|6|因有一嬰孩為我們而生； 有一子賜給我們。 政權必擔在他的肩頭上； 他名稱為「奇妙策士、全能的上帝、永在的父、和平的君」。
ISA|9|7|他的政權與平安必加增無窮。 他必在 大衛 的寶座上治理他的國， 以公平公義使國堅定穩固， 從今直到永遠。 萬軍之耶和華的熱心必成就這事。
ISA|9|8|主向 雅各 家發出言語， 主的話臨到 以色列 家。
ISA|9|9|眾百姓，就是 以法蓮 和 撒瑪利亞 的居民， 都將知道； 他們憑驕傲自大的心說：
ISA|9|10|「磚塊掉落了，我們要鑿石頭重建； 桑樹砍了，我們要改種香柏樹。」
ISA|9|11|因此，耶和華興起 利汛 的敵人 前來攻擊 以色列 ， 要激起它的仇敵，
ISA|9|12|東有 亞蘭 人，西有 非利士 人； 他們張口吞吃 以色列 。 雖然如此，耶和華的怒氣並未轉消； 他的手依然伸出。
ISA|9|13|這百姓還沒有歸向擊打他們的主， 也沒有尋求萬軍之耶和華。
ISA|9|14|耶和華在一日之間 從 以色列 中剪除了頭與尾－ 棕樹枝與蘆葦－
ISA|9|15|長老和顯要就是頭， 以謊言教人的先知就是尾。
ISA|9|16|因為引導這百姓的使他們走入迷途， 被引導的都必被吞滅。
ISA|9|17|所以，主不喜愛 他們的青年， 也不憐憫他們的孤兒和寡婦； 因為他們都是褻瀆的，行惡的， 並且各人的口都說愚妄的話。 雖然如此，耶和華的怒氣並未轉消； 他的手依然伸出。
ISA|9|18|邪惡如火焚燒， 吞滅荊棘和蒺藜， 在稠密的樹林中點燃， 成為煙柱，旋轉上騰。
ISA|9|19|因萬軍之耶和華的烈怒，地都燒遍了； 百姓成為柴火， 無人憐惜弟兄。
ISA|9|20|有人右邊搶奪，猶受飢餓； 左邊吞吃，仍不飽足， 各人吃自己膀臂上的肉。
ISA|9|21|瑪拿西 吞吃 以法蓮 ， 以法蓮 吞吃 瑪拿西 ， 他們又一同攻擊 猶大 。 雖然如此，耶和華的怒氣並未轉消； 他的手依然伸出。
ISA|10|1|禍哉！那些設立不義之律例的， 和記錄奸詐之判詞的，
ISA|10|2|為要扭曲貧寒人的案件， 奪去我民中困苦人的理， 以寡婦當作擄物， 以孤兒當作掠物。
ISA|10|3|到降罰的日子，災禍從遠方臨到， 那時，你們要怎麼辦呢？ 你們要向誰逃奔求救呢？ 你們的財寶要存放何處呢？
ISA|10|4|他們只得屈身在被擄的人之下， 仆倒在被殺的人中間 。 雖然如此，耶和華的怒氣並未轉消； 他的手依然伸出。
ISA|10|5|禍哉！ 亞述 ，我怒氣的棍！ 他們手中的杖是我的惱恨。
ISA|10|6|我要差遣他攻擊褻瀆的國， 吩咐他對付我所惱怒的民， 搶走擄物，奪取掠物， 將他們踐踏，如同街上的泥土一般。
ISA|10|7|然而，這並非他的意念， 他的心不是這樣打算； 他的心要摧毀， 要剪除不少的國家。
ISA|10|8|他說：「我的官長豈不都是君王嗎？
ISA|10|9|迦勒挪 豈不像 迦基米施 嗎？ 哈馬 豈不像 亞珥拔 嗎？ 撒瑪利亞 豈不像 大馬士革 嗎？
ISA|10|10|既然我的手已伸到了這些有偶像的國， 他們所雕刻的偶像 過於 耶路撒冷 和 撒瑪利亞 的偶像，
ISA|10|11|我豈不照樣待 耶路撒冷 和其中的偶像， 如同我待 撒瑪利亞 和其中的偶像嗎？」
ISA|10|12|主在 錫安山 和 耶路撒冷 成就他一切工作的時候，說：「我必懲罰 亞述 王自大的心和他高傲尊貴的眼目。」
ISA|10|13|因為他說： 「我所成就的事是靠我手的能力 和我的智慧， 因為我本有聰明。 我挪移列國的地界， 搶奪他們所積蓄的財寶， 並且像勇士，使坐寶座的降為卑。
ISA|10|14|我的手奪取列國的財寶， 好像人奪取鳥窩； 我得了全地， 好像人拾起被棄的鳥蛋； 沒有振動翅膀的， 沒有張嘴的，也沒有鳴叫的。」
ISA|10|15|斧豈可向用斧砍伐的自誇呢？ 鋸豈可向拉鋸的自大呢？ 這好比棍揮動那舉棍的， 好比杖舉起那不是木頭的人。
ISA|10|16|因此，主－萬軍之耶和華 必使 亞述 王的壯士變為瘦弱， 在他的榮華之下必有火點燃， 如同火在燃燒一般。
ISA|10|17|以色列 的光必變成火， 它的聖者必成為火焰； 一日之間，將 亞述 王的荊棘和蒺藜焚燒淨盡，
ISA|10|18|又毀滅樹林和田園的榮華， 連魂帶體，好像病重的人消逝 一樣。
ISA|10|19|他林中只剩下稀少的樹木， 連孩童也能寫其數目。
ISA|10|20|到那日， 以色列 所剩下的和 雅各 家所逃脫的，必不再倚靠那擊打他們的，卻要誠心仰賴耶和華－ 以色列 的聖者。
ISA|10|21|所剩下的，就是 雅各 家的餘民，必歸回全能的上帝。
ISA|10|22|以色列 啊，你的百姓雖多如海沙，惟有剩下的歸回。滅絕之事已成定局，公義必如水漲溢。
ISA|10|23|因為萬軍之主耶和華在全地必成就所定的滅絕之事。
ISA|10|24|所以，萬軍之主耶和華如此說：「住 錫安 我的百姓啊， 亞述 王雖然用棍擊打你，又如 埃及 舉杖攻擊你，你不要怕他。
ISA|10|25|因為還有一點點時候，我向你們發的憤怒就要結束，我的怒氣要使他們滅亡。
ISA|10|26|萬軍之耶和華要舉起鞭子來攻擊他，好像在 俄立 磐石那裏擊打 米甸 人一樣。他的杖向海伸出，他必把杖舉起，如在 埃及 一般。
ISA|10|27|到那日， 亞述 王的重擔必離開你的肩頭，他的軛必離開你的頸項；那軛必因肥壯而撐斷 。」
ISA|10|28|亞述 王來到 亞葉 ， 經過 米磯崙 ， 在 密抹 安放輜重。
ISA|10|29|他們過了隘口， 要在 迦巴 住宿。 拉瑪 戰兢， 掃羅 的 基比亞 逃命。
ISA|10|30|迦琳 哪，要高聲呼喊！ 注意聽， 萊煞 啊！ 困苦的 亞拿突 啊 ！
ISA|10|31|瑪得米那 躲避， 基柄 的居民逃遁。
ISA|10|32|當那日， 亞述 王要在 挪伯 停留， 揮手攻擊 錫安 的山， 就是 耶路撒冷 的山。
ISA|10|33|看哪，主－萬軍之耶和華 以猛撞削斷樹枝； 巨木必被砍下， 高大的樹必降為低。
ISA|10|34|稠密的樹林，他要用鐵器砍下， 黎巴嫩 必被大能者伐倒 。
ISA|11|1|從 耶西 的殘幹必長出嫩枝， 他的根所抽的枝子必結果實。
ISA|11|2|耶和華的靈必住在他身上， 就是智慧和聰明的靈， 謀略和能力的靈， 知識和敬畏耶和華的靈。
ISA|11|3|他必以敬畏耶和華為樂； 行審判不憑眼見， 斷是非也不憑耳聞；
ISA|11|4|卻要以公義審判貧寒人， 以正直判斷地上的困苦人， 以口中的棍擊打全地， 以嘴裏的氣殺戮惡人。
ISA|11|5|公義必當他的腰帶， 信實必作他脅下的帶子。
ISA|11|6|野狼必與小綿羊同住， 豹子與小山羊同臥； 少壯獅子、牛犢和肥畜同群 ； 孩童要牽引牠們。
ISA|11|7|牛必與熊同食， 牛犢與小熊同臥； 獅子與牛一樣吃草。
ISA|11|8|吃奶的嬰孩在虺蛇的洞口玩耍， 斷奶的幼兒必按手在毒蛇的穴上。
ISA|11|9|在我聖山各處， 牠們都不傷人，不害物； 因為認識耶和華的知識要遍滿全地， 好像水充滿海洋一般。
ISA|11|10|到那日， 耶西 的根立作萬民的大旗；列國的人必尋求他，他安歇之所大有榮耀。
ISA|11|11|當那日，主必再度伸手救回自己百姓中所剩餘的，就是在 亞述 、 埃及 、 巴特羅 、 古實 、 以攔 、 示拿 、 哈馬 ，並眾海島所剩下的。
ISA|11|12|他要向列國豎立大旗， 召集 以色列 被趕散的人， 又從地極四方聚集分散的 猶大 人。
ISA|11|13|以法蓮 的嫉妒必消散， 苦待 猶大 的也被剪除； 以法蓮 必不嫉妒 猶大 ， 猶大 也不苦待 以法蓮 。
ISA|11|14|他們要飛向西方， 撲在 非利士 人的肩頭上， 他們要一同擄掠東方人， 他們的手伸到 以東 和 摩押 ； 亞捫 人也必順服他們。
ISA|11|15|耶和華必使 埃及 的海灣全然毀壞 ， 他舉手在 大河 之上颳起了暴熱的風， 擊打它，使它分成七條溪流， 人穿鞋便可渡過。
ISA|11|16|必有一條大道， 為百姓中從 亞述 逃脫生還的餘民而開， 如當日為 以色列 從 埃及 上來一樣。
ISA|12|1|在那日，你要說： 「耶和華啊，我要稱謝你！ 因為你雖然向我發怒， 你的怒氣卻已轉消； 你又安慰了我。
ISA|12|2|「看哪！上帝是我的拯救； 我要倚靠他，並不懼怕。 因為主耶和華是我的力量， 是我的詩歌， 他也成了我的拯救。」
ISA|12|3|你們必從救恩的泉源歡然取水。
ISA|12|4|在那日，你們要說： 「當稱謝耶和華，求告他的名； 在萬民中傳揚他的作為， 宣告他的名已被尊崇。
ISA|12|5|「你們要向耶和華唱歌， 因他所做的十分宏偉； 但願這事遍傳全地。
ISA|12|6|錫安 的居民哪，當揚聲歡呼， 因為在你們當中的 以色列 聖者最為偉大。」
ISA|13|1|亞摩斯 的兒子 以賽亞 所見，有關 巴比倫 的默示。
ISA|13|2|你們要在荒涼的山上豎立大旗， 向他們揚聲， 揮手招呼他們進入貴族之門。
ISA|13|3|我吩咐我所分別為聖的人， 召喚我的勇士， 就是我那狂喜高傲的人， 為要執行我的怒氣。
ISA|13|4|聽啊，山間有喧鬧的聲音， 好像有許多百姓聚集， 聽啊，多國之民聚集鬧鬨的聲音； 這是萬軍之耶和華召集作戰的軍隊。
ISA|13|5|他們從遠方來， 從天邊來， 耶和華和他惱恨的兵器 要毀滅全地。
ISA|13|6|你們要哀號， 因為耶和華的日子臨近了！ 這日來到，好像毀滅從全能者來到。
ISA|13|7|因此，人的手都變軟弱， 人的心都必惶惶。
ISA|13|8|他們必驚恐， 悲痛和愁苦將他們抓住。 他們陣痛，好像臨產的婦人一樣， 彼此驚奇對看，臉如火焰。
ISA|13|9|看哪！耶和華的日子臨到， 必有殘忍、憤恨、烈怒， 使這地荒蕪， 除滅其中的罪人。
ISA|13|10|天上的星宿都不發光， 太陽一升起就變黑暗， 月亮也不放光。
ISA|13|11|我必因邪惡懲罰世界， 因罪孽懲罰惡人， 我要止息驕傲人的狂妄， 制伏殘暴者的傲慢。
ISA|13|12|我要使人比純金更少， 比 俄斐 的赤金還少。
ISA|13|13|我，萬軍之耶和華狂怒，就是發烈怒的日子， 要令天震動， 地必搖撼，離其本位。
ISA|13|14|人如被追趕的羚羊， 像無人聚集的羊群， 各自歸回本族， 逃到本地。
ISA|13|15|凡被追上的必被刺死， 凡被捉拿的必倒在刀下。
ISA|13|16|他們的嬰孩必在他們眼前被摔死， 他們的房屋被搶劫， 他們的妻子被污辱。
ISA|13|17|看哪，我必激起 瑪代 人攻擊他們， 瑪代 人並不看重銀子， 也不喜愛金子。
ISA|13|18|他們必用弓擊潰青年， 不憐憫婦人所生的； 眼也不顧惜孩子。
ISA|13|19|巴比倫 為列國的榮耀， 為 迦勒底 人所誇耀的華美， 必像上帝所傾覆的 所多瑪 、 蛾摩拉 一樣；
ISA|13|20|國中必永無人煙， 世世代代無人居住； 阿拉伯 人不在那裏支搭帳棚， 牧羊的人也不使羊群躺臥在那裏。
ISA|13|21|曠野的走獸躺臥在那裏， 咆哮的動物擠滿棲身之所； 鴕鳥住在那裏， 山羊鬼魔也在那裏跳舞。
ISA|13|22|土狼必在它的宮殿 呼號， 野狗在華美的殿裏吼叫。 巴比倫 的時辰臨近了， 它的日子必不長久。
ISA|14|1|耶和華要憐憫 雅各 ，再度揀選 以色列 ，將他們安頓在本地。寄居的必與他們聯合，加入 雅各 家。
ISA|14|2|外邦人要將他們帶回本地。 以色列 家必在耶和華的地上得外邦人為僕婢，也要擄掠先前擄掠他們的，轄制先前欺壓他們的。
ISA|14|3|當耶和華使你得享安息，脫離愁苦、煩惱，和被迫做苦工的日子，
ISA|14|4|你必唱這詩歌嘲諷 巴比倫 王說： 「欺壓人的竟然滅亡！ 他的兇暴 竟然止息！
ISA|14|5|耶和華折斷惡人的杖， 打斷統治者的權杖；
ISA|14|6|他們在憤怒中連連攻擊萬民， 在怒氣中轄制列國， 逼迫他們，毫不留情。
ISA|14|7|現在全地得安息，享平靜， 人都出聲歡呼。
ISA|14|8|松樹和 黎巴嫩 的香柏樹 都因你歡樂： 自從你仆倒， 再也無人上來砍伐我們。
ISA|14|9|下面的陰間因你震動， 迎接你的到來； 在世曾為領袖的陰魂為你驚動， 那曾為列國君王的，都從寶座起立。
ISA|14|10|他們都要發言，對你說： 『你也變為軟弱，像我們一樣嗎？ 你也成了我們的樣子嗎？』
ISA|14|11|你的威嚴和琴瑟的聲音都下到陰間。 你下面鋪的是蟲，上面蓋的是蛆。
ISA|14|12|「明亮之星，早晨之子啊， 你竟然從天墜落！ 你這攻敗列國的，竟然被砍倒在地上！
ISA|14|13|你心裏曾說： 『我要升到天上， 我要高舉我的寶座在上帝的眾星之上， 我要坐在會眾聚集的山上，在極北的地方。
ISA|14|14|我要升到高雲之上， 我要與至高者同等。』
ISA|14|15|然而，你必墜落陰間， 到地府極深之處。
ISA|14|16|凡看見你的都要定睛望你， 留意看你，說： 『就是這個人嗎？ 他使大地顫抖， 使列國震動，
ISA|14|17|使世界如同荒野， 使城鎮傾覆； 是他，不釋放被擄的人歸家。』
ISA|14|18|列國的君王各自在自己的墳墓中， 在尊榮裏長眠。
ISA|14|19|惟獨你被拋棄在你的墳墓之外， 有如被厭惡的枝子 ， 被許多用刀刺透殺死的人覆蓋著， 一同墜落地府的石頭那裏， 像被踐踏的屍首。
ISA|14|20|你不得與君王同葬， 因為你毀壞你的國，殺戮你的民。 「惡人的後裔永不留名。
ISA|14|21|為了祖先的罪孽， 要預備他子孫的屠宰場， 免得他們興起，奪得全地， 使城市遍滿地面。」
ISA|14|22|萬軍之耶和華說： 「我必起來攻擊他們， 將 巴比倫 的名號和剩餘的人， 連子帶孫一併剪除； 這是耶和華說的。
ISA|14|23|「我必使 巴比倫 為豪豬佔據， 成為泥沼之地； 我要用滅命的掃帚掃淨它； 這是萬軍之耶和華說的。」
ISA|14|24|萬軍之耶和華起誓說： 「我怎樣思想，必照樣成就； 我怎樣定意，必照樣堅立，
ISA|14|25|要在我的地上擊破 亞述 ， 在我的山上將它踐踏。 它的軛必離開受壓制的人， 它的重擔必離開他們的肩頭。」
ISA|14|26|這是向全地所定的旨意， 向萬國所伸出的手。
ISA|14|27|萬軍之耶和華既然定意，誰能阻撓呢？ 他的手已經伸出，誰能使它縮回呢？
ISA|14|28|亞哈斯 王崩的那年，有默示如下：
ISA|14|29|「全 非利士 啊， 不要因擊打你的杖折斷就喜樂。 因為蛇必生出毒蛇， 牠所生的是會飛的火蛇。
ISA|14|30|貧寒人的長子必有得吃； 貧窮人必安然躺臥。 我必以饑荒滅絕你的根， 牠 必殺盡你所剩餘的人。
ISA|14|31|門哪，哀號吧！ 城啊，呼喊吧！ 全 非利士 都熔化了！ 因為有煙從北方而來， 在它的行伍中沒有掉隊的。」
ISA|14|32|當如何回答外邦的使者呢？ 「耶和華建立了 錫安 ， 在其中他困苦的百姓必有倚靠。」
ISA|15|1|論 摩押 的默示。 一夜之間， 摩押 的 亞珥 變為荒廢， 歸於無有； 一夜之間， 摩押 的 基珥 變為荒廢， 歸於無有。
ISA|15|2|摩押 上到神廟和 底本 的丘壇去哭泣； 它因 尼波 和 米底巴 哀號， 各人頭上光禿，鬍鬚剃淨。
ISA|15|3|他們在街市上腰束麻布， 都在房頂和廣場上哀號， 淚流不停。
ISA|15|4|希實本 和 以利亞利 呼喊， 他們的聲音達到 雅雜 ， 所以 摩押 的士兵高聲喊叫， 他們的心戰兢。
ISA|15|5|我的心 為 摩押 哀號； 它的難民逃到 瑣珥 ， 逃到 伊基拉‧施利施亞 。 他們上 魯希坡 ，隨走隨哭， 在 何羅念 的路上，因毀滅發出哀聲。
ISA|15|6|寧林 的水乾涸， 青草枯乾，嫩草死光， 青綠之物，一無所有。
ISA|15|7|因此， 摩押 人所得的財物和積蓄 都要運過 柳樹河 。
ISA|15|8|哀聲遍傳 摩押 四境， 哀號的聲音達到 以基蓮 ， 哀號的聲音遠及 比珥‧以琳 。
ISA|15|9|底們 的水充滿了血， 然而我還要加添 底們 的災難， 讓獅子追上 摩押 的難民 和那地 剩餘的人。
ISA|16|1|你們當將 羔羊奉送給那地的掌權者， 從 西拉 往曠野，送到 錫安 的山。
ISA|16|2|摩押 的居民 來到 亞嫩 渡口， 如逃遁的飛鳥，被趕離鳥巢 。
ISA|16|3|求你賜謀略，行公平， 使你的影子在正午如黑夜， 掩護逃亡的人，不洩露逃難者的行蹤。
ISA|16|4|願我 摩押 逃亡的人 寄居在你那裏， 你作他們的避難所，躲避滅命者的面。 勒索的人消失， 毀滅的事止息， 欺壓者從國中除滅，
ISA|16|5|在 大衛 帳幕中必有寶座因慈愛堅立， 必有一位君王憑信實坐在其上， 施行審判，尋求公平，迅速行公義。
ISA|16|6|我們聽聞 摩押 的驕傲， 極其驕傲； 它狂妄、驕傲、自大， 它誇大的言詞都是空的。
ISA|16|7|因此， 摩押 人必為 摩押 哀號， 人人都要哀號。 你們要為 吉珥‧哈列設 的葡萄餅哀嘆， 極其憂傷。
ISA|16|8|因為 希實本 的田地 和 西比瑪 的葡萄樹都衰殘了， 列國的君主折斷它的枝幹， 這枝子曾長到 雅謝 ，延伸到曠野， 嫩枝向外伸出，直伸過海；
ISA|16|9|所以，我要為 西比瑪 的葡萄樹哀哭， 像 雅謝 人一樣哀哭。 希實本 、 以利亞利 啊， 我要以眼淚澆灌你， 你因夏天果子和收割的莊稼， 歡呼聲已經止息了。
ISA|16|10|田園中不再有歡喜快樂， 葡萄園裏必無人歌唱，無人歡呼， 在壓酒池中踹酒的不再踹酒了， 我使歡呼的聲音止息了 。
ISA|16|11|因此，我的心腸為 摩押 哀鳴如琴， 我的內心為 吉珥‧哈列設 哀哭。
ISA|16|12|當 摩押 人出現在丘壇，筋疲力盡時，雖然到自己的聖所祈禱，卻仍無濟於事。
ISA|16|13|這是耶和華曾論到 摩押 的話。
ISA|16|14|但現在，耶和華說：「三年之內，按照雇工年數的算法， 摩押 的榮華必變為羞辱，人口雖曾眾多，剩餘的又少又弱。」
ISA|17|1|論 大馬士革 的默示。 看哪， 大馬士革 不再為城市， 變為廢墟。
ISA|17|2|亞羅珥 的城鎮被撇棄 ， 將成為牧羊之處， 羊群在那裏躺臥， 無人使牠們驚嚇。
ISA|17|3|以法蓮 不再有堡壘， 大馬士革 失去其王國， 亞蘭 的百姓所剩無幾， 如 以色列 人的榮美消失一般； 這是萬軍之耶和華說的。
ISA|17|4|到那日， 雅各 的榮美必失色， 它肥胖的身軀漸漸消瘦；
ISA|17|5|像人收割成熟的禾稼， 用手臂割取麥穗， 又像人在 利乏音谷 拾取穗子；
ISA|17|6|其間所剩不多，好像人打橄欖樹， 在最高的樹梢上只剩兩、三顆橄欖， 在多結果子的旁枝上只剩四、五顆； 這是耶和華－ 以色列 的上帝說的。
ISA|17|7|當那日，人必仰望造他們的主，眼目看著 以色列 的聖者。
ISA|17|8|他們必不仰望自己手所築的祭壇，也不理會自己指頭所造的 亞舍拉 和香壇。
ISA|17|9|當那日，他們堅固的城必因 以色列 人的緣故，如同樹林中和山頂上所撇棄的地方 。這樣，地就荒蕪了。
ISA|17|10|因你忘記拯救你的上帝， 忘記那保護你的磐石； 所以，你雖栽上佳美的樹苗， 插上別樣的枝子，
ISA|17|11|栽種的日子，你使它生長， 栽種的早晨，你使它開花， 但在愁苦、極其傷痛的日子， 所收割的都歸無有。
ISA|17|12|唉！萬民鬧鬨，好像海浪澎湃， 列邦喧鬧，如同洪水滔滔，
ISA|17|13|列邦喧鬧，如同大水滔滔； 但上帝一斥責，他們就遠遠躲避， 他們被追趕，如同山上風前的糠秕， 又如暴風前的碎秸；
ISA|17|14|看哪，晚上有驚嚇，未到早晨它就消失無蹤。 這是擄掠我們之人的厄運，是搶奪我們之人的報應。
ISA|18|1|禍哉！ 古實河 的那一邊、翅膀刷刷作響之地，
ISA|18|2|差遣使者在水面上， 坐蒲草船過海。 你們這些疾行的使者， 要到高大光滑的民那裏去； 那民遠近都畏懼， 是強大好征服的國， 土地有河流穿過。
ISA|18|3|世上所有的居民，住在地上的人哪， 山上大旗豎起時，你們要看， 號角吹響時，你們要聽。
ISA|18|4|耶和華對我如此說： 「我要安靜，從我的居所觀看， 如同日光下閃爍的熱氣， 又如收割時 露水蒸發的雲霧。」
ISA|18|5|收割之前，花蕾先謝， 花成了將熟的葡萄； 他必用刀削去嫩枝， 砍掉蔓延的枝條，
ISA|18|6|一起丟給山間的鷙鳥和地上的野獸； 鷙鳥要在其上避暑， 地上一切的野獸都在那裏過冬。
ISA|18|7|到那時，這高大光滑的民， 遠近都畏懼的民、 強大好征服之國、 土地有河流穿過； 他們必被當作 禮物獻給萬軍之耶和華， 獻到 錫安山 － 萬軍之耶和華立他名的地方。
ISA|19|1|論 埃及 的默示。 看哪，耶和華乘駕快雲， 臨到 埃及 ； 埃及 的偶像在他面前戰兢， 埃及 人的心在裏面消溶。
ISA|19|2|我要激起 埃及 人攻擊 埃及 人， 弟兄攻擊弟兄， 鄰舍攻擊鄰舍， 這城攻擊那城， 這國攻擊那國。
ISA|19|3|埃及 人的心神在裏面耗盡， 我要破壞他們的計謀。 他們必求問偶像和念咒的， 求問招魂的與行巫術的人。
ISA|19|4|我要將 埃及 人交在嚴厲的主人手中， 殘暴的君王必管轄他們； 這是主－萬軍之耶和華說的。
ISA|19|5|海水枯竭， 河流乾涸，
ISA|19|6|江河發臭， 埃及 的河水必然減少而枯乾。 蘆葦和蘆荻枯萎，
ISA|19|7|尼羅河 旁的植物 ，在 尼羅河 的沿岸， 並 尼羅河 旁所種的一切 全都枯焦，被風吹去，歸於無有。
ISA|19|8|打魚的哀哭， 所有在 尼羅河 釣魚的都必悲傷， 在水上撒網的也都衰殘。
ISA|19|9|以細緻的麻編織的必羞愧， 織布的必變蒼白 ；
ISA|19|10|織布的心情沮喪 ， 所有的傭工心都愁煩。
ISA|19|11|瑣安 的官長極其愚昧， 法老智慧的謀士籌劃愚謀； 你們怎敢對法老說： 「我是智慧人的子孫， 是古代國王的後裔？」
ISA|19|12|你的智慧人在哪裏？ 萬軍之耶和華向 埃及 所定的旨意， 他們既然知道，就讓他們告訴你吧！
ISA|19|13|瑣安 的官長愚昧， 挪弗 的官長受蒙蔽； 作 埃及 支派棟梁的， 帶領 埃及 走錯了路。
ISA|19|14|耶和華使歪曲的靈滲入 埃及 中間， 讓他們使 埃及 一切所做的都出差錯， 好像醉酒之人嘔吐時東倒西歪一樣。
ISA|19|15|在 埃及 ，無論是頭是尾， 棕樹枝與蘆葦，所做的事都不得成就。
ISA|19|16|到那日， 埃及 必像婦人一樣，因萬軍之耶和華揮手攻擊而戰兢懼怕。
ISA|19|17|猶大 地必使 埃及 驚恐，不論向誰提起，他都懼怕。這是因萬軍之耶和華向 埃及 所定的旨意。
ISA|19|18|當那日， 埃及 地必有五個城市的人說 迦南 的語言，又指著萬軍之耶和華起誓。有一城必稱為「太陽城」 。
ISA|19|19|在那日，在 埃及 地將有獻給耶和華的一座壇，邊界上必有為耶和華立的一根柱子。
ISA|19|20|這都要在 埃及 地為萬軍之耶和華作記號和證據。 埃及 人因受欺壓哀求耶和華，他就差遣一位救主作護衛者，拯救他們，
ISA|19|21|耶和華就被 埃及 所認識。在那日， 埃及 人要認識耶和華，獻牲祭和素祭敬拜他，並向耶和華許願還願。
ISA|19|22|耶和華必擊打 埃及 ，又擊打又醫治， 埃及 人就歸向耶和華。他必應允他們的禱告，醫治他們。
ISA|19|23|在那日，必有從 埃及 通往 亞述 的大道。 亞述 人要進入 埃及 ， 埃及 人也要進入 亞述 ； 埃及 人要與 亞述 人一同敬拜。
ISA|19|24|在那日， 以色列 將與 埃及 、 亞述 三國一起，使地上的人得福。
ISA|19|25|萬軍之耶和華必賜福給他們，說：「 埃及 －我的百姓， 亞述 －我手的工作， 以色列 －我的產業，都有福了！」
ISA|20|1|亞述 元帥 受 亞述 王 撒珥根 派遣往 亞實突 的那年，他攻打 亞實突 ，將城攻取。
ISA|20|2|那時，耶和華吩咐 亞摩斯 的兒子 以賽亞 說：「你去解掉你腰間的麻布，脫下你腳上的鞋。」 以賽亞 就這樣做，赤身赤腳行走。
ISA|20|3|耶和華說：「我僕人 以賽亞 怎樣赤身赤腳行走三年，作為關於 埃及 和 古實 的預兆奇蹟，
ISA|20|4|照樣， 亞述 王必擄去 埃及 人，掠去 古實 人，無論老少，都赤身赤腳，露出下體，使 埃及 蒙羞。
ISA|20|5|以色列 人必驚惶羞愧，因為他們仰望 古實 ，以 埃及 為榮。
ISA|20|6|「那時，沿海一帶的居民必說：『看哪，我們素來所仰望的，就是為躲避 亞述 王所逃往 求救的，不過如此！我們怎能逃脫呢？』」
ISA|21|1|論海邊曠野的默示。 它像 尼革夫 的旋風掃過， 從曠野，從可怕之地而來。
ISA|21|2|有悽慘的異象向我揭示： 「詭詐的在行詭詐，毀滅的在行毀滅。 以攔 哪，前進吧！ 瑪代 啊，圍攻吧！ 我使它一切的嘆息停止了。」
ISA|21|3|為此，我腰部滿是疼痛， 痛苦將我抓住， 好像臨產的婦人一樣的痛。 我疼痛甚至不能聽， 我驚惶甚至不能看 。
ISA|21|4|我心慌亂，驚恐威嚇我。 我所渴望的黃昏，反成為我的恐懼。
ISA|21|5|有人擺設筵席， 鋪上地毯，又吃又喝。 「官長啊，起來， 抹亮盾牌。」
ISA|21|6|主對我如此說： 「你去設立守望者， 讓他報告他所看見的。
ISA|21|7|他會看見一對一對騎著馬的軍隊， 又看見驢隊，駱駝隊， 他要留心聽，仔細地聽。」
ISA|21|8|他如獅子般吼叫 ： 「主啊，我白天常站在暸望樓， 徹夜立在我的暸望臺。」
ISA|21|9|看哪，有一對一對騎著馬的軍隊前來。 他就回應說：「 巴比倫 傾倒了！傾倒了！ 他把 巴比倫 神明的一切雕刻偶像都打碎在地上了。」
ISA|21|10|我被打的禾稼，我禾場上的穀物啊， 我從萬軍之耶和華－ 以色列 的上帝那裏所聽見的，都告訴你們了。
ISA|21|11|論 度瑪 的默示。 有人聲從 西珥 呼喊： 「守望的啊，夜裏如何？ 守望的啊，夜裏如何？」
ISA|21|12|守望者說： 「早晨來到，黑夜將臨。 你們若要問，問吧， 也可以回頭再來。」
ISA|21|13|論 阿拉伯 的默示。 底但 的旅行商隊啊， 你們在 阿拉伯 的樹林中住宿。
ISA|21|14|提瑪 地的居民哪， 提水來迎接口渴的人， 帶餅來迎接難民。
ISA|21|15|他們躲避刀劍和出了鞘的刀， 躲避上了弦的弓與戰爭的重災。
ISA|21|16|主對我這樣說：「一年之內，按照雇工年數的算法， 基達 一切的繁華必歸無有。
ISA|21|17|基達 人中強壯弓箭手剩下的數目甚為稀少，這是耶和華－ 以色列 的上帝說的。」
ISA|22|1|論異象谷的默示。 甚麼事使你們上去， 全都上到屋頂呢？
ISA|22|2|你這四處吶喊、大聲喧嘩的城、 歡樂的邑啊， 你被殺的並非被刀所殺， 也不是因打仗陣亡。
ISA|22|3|你所有的官長一同奔逃， 不用弓箭就被捆綁 ； 你們即使逃往遠方， 也要被找到，一同被捆綁。
ISA|22|4|因此我說： 「不要看我， 讓我痛哭吧！ 不要因我百姓 的毀滅竭力安慰我。」
ISA|22|5|因為這是萬軍之主耶和華使異象谷 混亂、踐踏、煩擾的日子； 城牆被攻破， 哀聲達到山上。
ISA|22|6|以攔 提著箭袋， 有戰車、士兵、騎兵； 吉珥 亮出盾牌，
ISA|22|7|你佳美的山谷遍佈戰車， 騎兵排列在城門前。
ISA|22|8|他除掉 猶大 的防禦。 那時，你指望森林庫裏的兵器。
ISA|22|9|你們看見 大衛城 缺口很多，就匯集 下池 的水；
ISA|22|10|你們數點 耶路撒冷 的房屋，拆毀房屋，用以修補城牆，
ISA|22|11|又在兩道城牆中間挖水池，用以盛舊池的水，卻不仰望成就這事的主，也不顧念從古時定這事的主。
ISA|22|12|當那日，萬軍之主耶和華使人哭泣哀號， 頭上光禿，身披麻布。
ISA|22|13|看哪，人卻歡喜快樂， 宰牛殺羊，吃肉喝酒： 「讓我們吃吃喝喝吧！因為明天要死了。」
ISA|22|14|萬軍之耶和華開啟我的耳朵： 「這罪孽直到你們死，斷不得赦免！」 這是萬軍之主耶和華說的。
ISA|22|15|萬軍之主耶和華如此說：「你到 舍伯那 宮廷總管那裏去，說：
ISA|22|16|『你在這裏憑甚麼？你在這裏靠誰？竟敢在這裏為自己鑿墳墓，在高處為自己鑿墳墓，在巖石中為自己挖安身之所！
ISA|22|17|你這偉大的人，看哪，耶和華必將你用力拋出，將你緊緊纏裹。
ISA|22|18|他必將你捲成一團，好像拋球一樣拋向寬闊之地。你這主人家的羞辱啊，你必死在那裏，你引以為榮的戰車也毀在那裏。
ISA|22|19|我要革除你的官職，你必從原位被逐 。』
ISA|22|20|「到那日，我要召 希勒家 的兒子─我的僕人 以利亞敬 來，
ISA|22|21|將你的外袍給他穿上，將你的腰帶給他繫緊，將你的政權交在他手中。他必作 耶路撒冷 居民和 猶大 家的父。
ISA|22|22|我要將 大衛 家的鑰匙放在他肩頭上。他開了，無人能關；他關了，無人能開。
ISA|22|23|我要使他立穩，像釘子釘在堅固的地方；他必成為他父家榮耀的寶座。
ISA|22|24|他父家所有的榮耀，連兒女帶子孫，有如杯碗、瓶罐的小器皿，都掛在他身上。
ISA|22|25|當那日，萬軍之耶和華說，釘在堅固處的釘子必挪移，被砍斷落地，掛在上面的各樣重擔都被切斷。這是耶和華說的。」
ISA|23|1|論 推羅 的默示。 哀號吧， 他施 的船隻！ 因為 推羅 已成廢墟，沒有房屋存留， 他們從 基提 地來的時候，得到這個消息 。
ISA|23|2|沿海的居民， 西頓 的商家啊， 當靜默無聲。 你差人航海 ，
ISA|23|3|在大水之上， 西曷河 的糧食、 尼羅河 的莊稼是 推羅 的進項， 它就成為列國的商埠。
ISA|23|4|西頓 ，你這海洋中的堡壘啊，應當羞愧， 因為大海說 ： 「我未經歷產痛，也沒有生產， 未曾養育男孩，也沒有撫養女孩。」
ISA|23|5|推羅 的風聲傳到 埃及 時， 他們為這風聲極其疼痛。
ISA|23|6|你們當渡到 他施 去， 哀號吧，沿海的居民！
ISA|23|7|這就是你們那古老歡樂的城市嗎？ 它的腳曾帶人到遠方居住。
ISA|23|8|誰定意 推羅 有這樣的遭遇呢？ 它本是賜冠冕的， 它的商家是王子， 生意人是世上尊貴的人。
ISA|23|9|這是萬軍之耶和華所定的， 為要貶抑一切榮耀的狂傲， 使地上一切尊貴的人被藐視。
ISA|23|10|他施 啊， 你要像 尼羅河 一樣在你的地氾濫， 不再有腰帶的束縛了。
ISA|23|11|耶和華已經向海伸手， 震動列國； 他出令對付 迦南 ， 要拆毀其中的堡壘。
ISA|23|12|他說：「受欺壓的少女 西頓 哪， 你必不再歡樂。 起來！渡到 基提 去， 就是在那裏也不得安歇。
ISA|23|13|看哪， 迦勒底 人之地，這國民如今已不復存在。 亞述 人使它 成為住曠野者的居所。他們建築自己的瞭望樓，拆毀它的宮殿，使它成為荒涼。
ISA|23|14|哀號吧， 他施 的船隻！ 因你們的堡壘已成廢墟。
ISA|23|15|到那時， 推羅 必被忘記七十年，就是一位君王的年數。七十年後， 推羅 的景況必如妓女之歌：
ISA|23|16|「你這被遺忘的妓女啊， 帶著琴周遊城內， 彈得美妙，唱許多歌， 好讓人記得你。」
ISA|23|17|七十年後，耶和華必巡視 推羅 ，使它再度獲利 ，與地面上的世界各國貿易 。
ISA|23|18|它的收益和獲利都要歸耶和華為聖，不再私自屯積存留；因為它的收益必歸給住在耶和華面前的人，使他們吃飽，穿華麗的衣服。
ISA|24|1|看哪，耶和華使地空虛，變為荒蕪， 地面扭曲，居民四散。
ISA|24|2|那時，百姓如何，祭司也如何； 僕人如何，主人也如何； 婢女如何，主母也如何； 買主如何，賣主也如何； 放債的如何，借貸的也如何； 債主如何，欠債的也如何。
ISA|24|3|地必全然空虛，盡都荒蕪， 因為這話是耶和華說的。
ISA|24|4|大地悲哀凋零， 世界敗落衰殘， 地上居高位的人也沒落了。
ISA|24|5|地被其上的居民所污穢， 因為他們犯了律法， 廢了律例，背了永約。
ISA|24|6|所以，詛咒吞滅大地， 住在其上的都有罪； 地上的居民被火焚燒， 剩下的人稀少。
ISA|24|7|新酒悲哀，葡萄樹凋殘， 心中歡樂的都嘆息。
ISA|24|8|擊鼓之樂停止， 狂歡者的喧嘩止住， 彈琴之樂也停止了。
ISA|24|9|人不再飲酒唱歌， 喝烈酒的，必以為苦。
ISA|24|10|荒涼的城拆毀了， 各家關閉，無法進入。
ISA|24|11|有人在街上嚷著要酒喝， 一切的喜樂變為昏暗， 地上的歡樂全都消失。
ISA|24|12|城裏盡是荒涼， 城門全都摧毀。
ISA|24|13|地上的萬民正像打過的橄欖樹， 又如葡萄釀酒以後再去摘取，所剩無幾。
ISA|24|14|他們要高聲歡呼， 從海那邊揚聲讚美耶和華的威嚴。
ISA|24|15|因此，你們要在日出之地榮耀耶和華， 在眾海島榮耀耶和華－ 以色列 上帝的名。
ISA|24|16|我們聽見從地極有人歌唱： 「榮耀歸於公義的那一位！」 我卻說：「我滅亡了！ 我滅亡了，我有禍了！ 詭詐的還在行詭詐， 詭詐的還在大行詭詐。」
ISA|24|17|地上的居民哪， 驚嚇、陷阱、羅網都臨到你；
ISA|24|18|躲過驚嚇之聲的墜入陷阱， 逃離陷阱的又被羅網纏住， 因為天上的窗戶都打開， 地的根基也震動。
ISA|24|19|地必全然破壞，盡都崩裂， 劇烈震動。
ISA|24|20|地要搖搖晃晃，好像醉酒的人， 又如小屋子搖來搖去； 罪過重壓其上， 它就塌陷，不能復起。
ISA|24|21|到那日，耶和華在天上必懲罰天上的軍隊， 在地上必懲罰地上的列王。
ISA|24|22|他們必被聚集， 像囚犯困在牢裏， 他們被關在監獄， 多日之後便受懲罰。
ISA|24|23|那時，月亮要蒙羞，太陽要慚愧， 因為萬軍之耶和華必在 錫安山 ， 在 耶路撒冷 作王， 在他眾長老面前彰顯榮耀。
ISA|25|1|耶和華啊，你是我的上帝， 我要尊崇你，稱頌你的名。 因為你以信實忠信 行遠古所定奇妙的事。
ISA|25|2|你使城市變為廢墟， 使堅固的城荒涼， 使外邦人的城堡不再為城， 永遠不再重建。
ISA|25|3|所以，強大的民必尊敬你， 殘暴之國的城必敬畏你。
ISA|25|4|因為你是貧寒人的保障， 貧窮人急難中的保障， 暴風雨之避難所， 炎熱地之陰涼處。 當殘暴者盛氣凌人的時候， 如暴風直吹牆壁，
ISA|25|5|如乾旱地的熱氣， 你要制止外邦人的喧嚷， 殘暴者的歌要停止， 好像熱氣因雲的陰影而消失。
ISA|25|6|在這山上，萬軍之耶和華必為萬民擺設宴席，有肥甘與美酒，就是滿有骨髓的肥甘與精釀的美酒。
ISA|25|7|在這山上，他必吞滅纏裹萬民的面紗和那遮蓋列國的遮蔽物。
ISA|25|8|他已吞滅死亡直到永遠。主耶和華必擦乾各人臉上的眼淚，在全地除去他百姓的羞辱；這是耶和華說的。
ISA|25|9|到那日，人必說：「看哪，這是我們的上帝，我們向來等候他，他必拯救我們。這是耶和華，我們向來等候他，我們必因他的救恩歡喜快樂。」
ISA|25|10|耶和華的手必按住這山， 摩押 人要被踐踏在他底下，好像乾草被踐踏在糞池 裏。
ISA|25|11|他們要在其中伸展雙手，好像游泳的人伸手游泳。他們的手雖靈巧，耶和華卻使他們的驕傲降為卑下。
ISA|25|12|他使你城牆上堅固的碉堡傾倒，夷為平地，化為塵土。
ISA|26|1|當那日，在 猶大 地，人必唱這歌： 「我們有堅固的城， 耶和華賜救恩為城牆，為城郭。
ISA|26|2|你們要敞開城門， 使守信的公義之民得以進入。
ISA|26|3|堅心倚賴你的，你必保守他十分平安， 因為他倚靠你。
ISA|26|4|你們當倚靠耶和華，直到永遠， 因為耶和華，耶和華是永遠的磐石。
ISA|26|5|他使居住高處的與高處的城市一同降為卑下， 將城拆毀，夷為平地，化為塵土，
ISA|26|6|使它被腳踐踏， 就是被困苦人和貧寒人的腳踐踏。」
ISA|26|7|義人的道是正直的， 正直的主啊，你修平義人的路。
ISA|26|8|耶和華啊，我們在你行審判的路上等候你 ， 我們心裏所渴慕的，就是你的名和你的稱號 。
ISA|26|9|夜間，我的心渴想你， 我裏面的靈切切尋求你。 因為你在地上行審判的時候， 世上的居民就學習公義。
ISA|26|10|惡人雖然領受恩惠， 仍未學到公義。 在正直之地，他行不義， 也不看耶和華的威嚴。
ISA|26|11|耶和華啊，你的手高舉，他們不觀看； 願他們觀看你為百姓發的熱心而羞愧， 願火吞滅你的敵人。
ISA|26|12|耶和華啊，你必賞賜我們平安， 因為我們所做的一切，都是你為我們成就的。
ISA|26|13|耶和華－我們的上帝啊， 在你以外曾有別的主管轄我們， 但我們惟獨稱揚你的名。
ISA|26|14|死去的不能再復活， 陰魂不能再興起； 你懲罰他們，使他們毀滅， 他們的名號 就全然消滅。
ISA|26|15|耶和華啊，你增添國民， 你增添國民，得了榮耀， 又拓展國土的疆界。
ISA|26|16|耶和華啊，他們在急難中尋求你。 你的管教臨到他們身上時， 他們傾吐低聲的禱告。
ISA|26|17|婦人懷孕，臨產疼痛， 在痛苦之中喊叫； 耶和華啊，我們在你面前也是如此。
ISA|26|18|我們曾懷孕，曾疼痛， 所生產的竟像風一樣， 並未帶給地上任何拯救； 世上也未曾有居民生下來 。
ISA|26|19|你的死人要復活， 我的屍首要起來。 睡在塵土裏的啊，要醒起歌唱！ 你的甘露好像晨曦 的甘露， 地要交出陰魂。
ISA|26|20|我的百姓啊，要進入內室， 關上你的門，躲避片刻， 等到憤怒過去。
ISA|26|21|因為，看哪，耶和華從他的居所出來， 要懲罰地上居民的罪孽。 地必露出其中的血， 不再掩蓋被殺的人。
ISA|27|1|到那日，耶和華必用他堅硬銳利的大刀懲罰 力威亞探 ，就是那爬得快的蛇，懲罰 力威亞探 ，就是那彎彎曲曲的蛇，並殺死海裏的大魚。
ISA|27|2|當那日，你們要唱這美好 葡萄園的歌：
ISA|27|3|「我－耶和華看守葡萄園，按時灌溉， 晝夜看守，免得有人損害。
ISA|27|4|我心中不存憤怒。 惟願在戰爭中我有荊棘和蒺藜， 我就起步攻擊他， 把他一同焚燒；
ISA|27|5|或者讓他緊靠我，以我為避難所， 與我和好， 與我和好。」
ISA|27|6|將來 雅各 要扎根， 以色列 要發芽開花， 果實遍滿地面。
ISA|27|7|耶和華擊打 以色列 ， 豈像擊打那些擊打他們的人嗎？ 以色列 被殺戮， 豈像其他人所遭遇的殺戮嗎？
ISA|27|8|你驅趕他們，放逐他們， 與他們相爭。 在颳東風的日子， 他以暴風趕逐他們。
ISA|27|9|所以， 雅各 的罪孽藉此得赦免， 除罪的效果盡在乎此； 他使祭壇的石頭變為粉碎的石灰， 使 亞舍拉 和香壇不再立起。
ISA|27|10|因為堅固的城變為荒涼， 成了被撇棄的居所，像曠野一樣； 牛犢在那裏吃草， 在那裏躺臥，吃盡其中的樹枝。
ISA|27|11|它的枝條一枯乾，就被折斷， 婦女用以點火燃燒。 因為這百姓蒙昧無知， 所以，造他們的必不憐憫他們， 造成他們的也不施恩給他們。
ISA|27|12|到那日， 以色列 人哪，耶和華必像人打樹拾果一般，從 大河 的支流，直到 埃及 的溪谷，將你們一一收集。
ISA|27|13|當那日，號角大響；在 亞述 地將亡的，與被趕散至 埃及 地的，都要前來，在 耶路撒冷 聖山上敬拜耶和華。
ISA|28|1|禍哉！ 以法蓮 酒徒高傲的冠冕， 其榮美竟如花凋殘； 他們在肥沃的山谷頂上， 被酒擊敗。
ISA|28|2|看哪，主有一位大能大力者， 如強烈的冰雹， 如毀滅的暴風雨， 如漲溢的洪水， 他必親手將他們摔落在地。
ISA|28|3|以法蓮 酒徒高傲的冠冕， 必被腳踐踏；
ISA|28|4|那如凋殘之花的榮美， 在肥沃的山谷頂上， 必如夏令前初熟的無花果， 讓看見的人注意， 摘到手裏，隨即吞吃。
ISA|28|5|到那日，萬軍之耶和華 必成為他餘民的榮冠華冕，
ISA|28|6|成為在位審判者的公平之靈， 和城門口制敵的力量。
ISA|28|7|這些人也因酒搖晃， 因烈酒東倒西歪。 祭司和先知因烈酒搖晃， 被酒所困， 因烈酒東倒西歪。 他們錯解默示， 審判時不分是非。
ISA|28|8|筵席上都滿了嘔吐的污穢， 沒有一處乾淨。
ISA|28|9|「他要將知識指教誰呢？ 要向誰闡明信息呢？ 是向那些剛斷奶的， 離開母親胸懷的嗎？
ISA|28|10|因為他咕噥咕噥，咕噥咕噥， 嘮嘮叨叨，嘮嘮叨叨， 這裏一點，那裏一點。」
ISA|28|11|耶和華要藉嘲弄的嘴唇和外邦人的舌頭， 向這百姓說話。
ISA|28|12|他曾對他們說： 「這是安歇之所， 你們要使疲乏的人得安歇， 這是歇息之處。」 他們卻不肯聽。
ISA|28|13|耶和華的話對他們而言是 「咕噥咕噥，咕噥咕噥， 嘮嘮叨叨， 嘮嘮叨叨， 這裏一點，那裏一點」； 以致他們往前行， 卻後仰跌倒，甚至跌傷， 落入陷阱，被抓住了。
ISA|28|14|因此，你們這些傲慢的人， 就是管轄住 耶路撒冷 這百姓的， 要聽耶和華的話。
ISA|28|15|你們曾說： 「我們已與死亡立約， 與陰間結盟， 不可擋的鞭子揮過時， 必不臨到我們； 因我們以謊言為避難所， 靠虛假來藏身」；
ISA|28|16|所以，主耶和華如此說： 「看哪，我在 錫安 放一塊石頭作為根基， 是衡量的石頭， 是寶貴的房角石，穩固的根基； 信靠他的人必不致驚恐。
ISA|28|17|我以公平為準繩， 以公義為鉛垂線； 冰雹必沖去謊言的避難所， 大水必漫過藏身之處。
ISA|28|18|你們與死亡所立的約必廢除， 與陰間所結的盟不得堅立； 不可擋的鞭子揮過時， 你們必被踐踏。
ISA|28|19|每逢它揮來，必將你們擄去； 每早晨它必揮過， 白晝黑夜都是如此。 明白這信息的都必驚恐。」
ISA|28|20|床榻短，人不能伸展； 被子窄，人無從裹身。
ISA|28|21|耶和華必興起，像在 毗拉心山 ， 他必發怒，如在 基遍谷 ； 為要做成他的工，就是非常的工， 成就他的事，就是奇異的事。
ISA|28|22|現在你們不可傲慢， 免得捆綁你們的繩索更結實， 因為我從萬軍之主耶和華那裏聽見， 在全地施行滅絕的事已定。
ISA|28|23|你們當側耳聽我的聲音， 留心聽我的言語。
ISA|28|24|那為撒種而耕地的 會不停地耕地，鬆土，耙地嗎？
ISA|28|25|他剷平了地面， 豈不就種小茴香， 播種大茴香， 按行列種小麥， 在定處種大麥， 在田邊種粗麥嗎？
ISA|28|26|他的上帝教導他， 指導他合宜的方法。
ISA|28|27|原來打小茴香，不用尖利的器具， 軋大茴香，也不是用車輪； 卻要用杖打小茴香， 用棍打大茴香。
ISA|28|28|穀要打， 但不能持續地搗， 用車輪和馬軋， 卻不軋碎它。
ISA|28|29|這也是出於萬軍之耶和華， 他的謀略奇妙， 他的智慧廣大。
ISA|29|1|禍哉！ 亞利伊勒 ， 亞利伊勒 ， 大衛 安營的城， 任憑你年復一年， 節期照常循環，
ISA|29|2|我卻要使 亞利伊勒 遭難； 它必悲傷哀號， 它對我是 亞利伊勒 。
ISA|29|3|我必四圍安營攻擊你， 築臺圍困你， 堆壘攻擊你。
ISA|29|4|你必敗落，從地裏說話， 你的言語細微出於塵埃。 你的聲音必像那招魂者的聲音出於地， 你的言語呢喃出於塵埃。
ISA|29|5|你那成群的陌生人 要像細塵， 暴民要像吹起的糠秕； 這事必頃刻之間忽然臨到。
ISA|29|6|萬軍之耶和華必使雷轟、地震、巨響、旋風、暴風， 並吞滅的火焰臨到它。
ISA|29|7|那時，攻擊 亞利伊勒 列國的軍隊， 與一切攻擊 亞利伊勒 和它城堡， 並帶給它患難的， 必如夢，如夜間的異象；
ISA|29|8|又像飢餓的人在夢中吃飯， 醒了仍覺飢腸轆轆； 或像口渴的人在夢中喝水， 醒了仍覺發昏，心裏想喝。 攻擊 錫安山 列國的軍隊也必如此。
ISA|29|9|你們等候驚奇吧！ 你們沉迷宴樂吧！ 他們醉了，卻非因酒； 東倒西歪，卻非因烈酒。
ISA|29|10|因為耶和華將沉睡的靈澆灌你們， 遮住你們的眼， 眼就是先知， 覆蓋你們的頭， 頭就是先見。
ISA|29|11|所有的默示，在你們看來都如封住的書卷，人將這書卷交給識字的人，說：「請念吧！」他說：「我不能念，因為它封住了。」
ISA|29|12|又將這書卷交給不識字的人，說：「請念吧！」他說：「我不識字。」
ISA|29|13|主說：「因這百姓以口親近我， 用嘴唇尊敬我， 心卻遠離我； 他們敬畏我， 不過是領受前人的命令。
ISA|29|14|所以，看哪，我要在這百姓中行奇妙的事， 就是奇妙又奇妙的事。 他們智慧人的智慧必然消滅， 聰明人的聰明必然消失。」
ISA|29|15|禍哉！那些向耶和華深藏謀略的， 他們在暗中行事，說： 「有誰看見我們呢？ 誰會注意我們呢？」
ISA|29|16|你們把事情顛倒了， 豈可看陶匠如陶土呢？ 受造物豈可論創造者說， 「他並沒有造我」？ 製成物豈可論製作者說， 「他根本不懂」？
ISA|29|17|黎巴嫩 變為田園， 田園看似森林， 不是只需要一些時間嗎？
ISA|29|18|那時，聾子必聽見這書上的話； 盲人的眼必從迷矇黑暗中看見。
ISA|29|19|困苦的人必因耶和華增添歡喜， 人間貧窮的必因 以色列 的聖者快樂。
ISA|29|20|因為殘暴的人歸於無有， 傲慢的人已經滅絕， 一切存心作惡的都被剪除。
ISA|29|21|他們憑一句話定一個人有罪， 為在城門口斷是非的設下羅網， 又用虛無的事屈枉義人。
ISA|29|22|所以，救贖 亞伯拉罕 的耶和華 論到 雅各 家時如此說： 「 雅各 必不再羞愧， 面容也不再變色。
ISA|29|23|當他的兒女看見 我的手在他們當中所成就的事情 ， 他們就必尊我的名為聖， 尊 雅各 的聖者為聖， 他們必敬畏 以色列 的上帝。
ISA|29|24|心中迷糊的必明白， 發怨言的必領受訓誨。」
ISA|30|1|耶和華說： 「禍哉！這悖逆的兒女。 他們同謀，卻不出於我， 結盟，卻不出於我的靈， 以致罪上加罪。
ISA|30|2|他們沒有尋求我的指示，就起身下 埃及 去， 要倚靠法老的庇護堅固自己， 並投在 埃及 的蔭下。
ISA|30|3|但法老的庇護反成為你們的羞辱； 你們投在 埃及 蔭下，反使你們慚愧。
ISA|30|4|他們的領袖已在 瑣安 ， 他們的使臣到了 哈內斯 。
ISA|30|5|他們必因那無益於他們的民蒙羞； 那民並非幫助，也非有益， 只帶來羞恥和凌辱。」
ISA|30|6|論 尼革夫 牲畜的默示。 他們將財物馱在驢背上， 將寶物馱在駱駝的背脊， 經過艱難困苦之地， 就是母獅、公獅、毒蛇、飛蛇之地， 往那無益於他們的民那裏去。
ISA|30|7|埃及 的幫助是徒然的， 因此，我稱它為「毫不中用的 拉哈伯 」 。
ISA|30|8|現在你要去， 在他們面前將這話刻在版上， 寫在書上， 以便流傳後世，直到永永遠遠 。
ISA|30|9|因為他們是悖逆的百姓、說謊的兒女， 是不肯聽從耶和華訓誨的兒女。
ISA|30|10|他們對先見說：「不要再看了」； 對先知說：「不要向我們預言正直的事； 要對我們說好聽的話， 預言虛幻的事。
ISA|30|11|要離開這道，偏離這路， 不要在我們面前再提說 以色列 的聖者。」
ISA|30|12|所以， 以色列 的聖者如此說： 「因你們藐視這話， 倚賴欺壓和詭詐，以此為可靠，
ISA|30|13|因此，這罪孽在你們身上， 好像高牆裏有凸起的裂縫， 頃刻之間忽然坍下來了；
ISA|30|14|它被砸碎，好像把陶匠的瓦器摔碎， 毫不顧惜， 甚至在碎塊中找不到一片 可用以從爐內取火，或從池中舀水。
ISA|30|15|主耶和華－ 以色列 的聖者如此說： 「你們得救在乎歸回安息， 得力在乎平靜安穩。」 你們卻是不肯，
ISA|30|16|你們說：「不然，我們要騎馬奔走」， 所以你們必然奔走。 你們又說：「我們要騎快馬」， 所以追趕你們的，也必飛快。
ISA|30|17|一人叱喝，令千人逃跑， 五人叱喝，你們都逃跑； 以致剩下的如山頂的旗杆， 如山岡上的大旗。
ISA|30|18|耶和華必然等候，要施恩給你們； 必然興起，好憐憫你們。 因為耶和華是公平的上帝； 凡等候他的都是有福的！
ISA|30|19|住在 錫安 、居於 耶路撒冷 的百姓啊，你必不再哭泣。主必因你哀求的聲音施恩給你，他聽見的時候就必應允你。
ISA|30|20|主雖然以艱難給你當餅，以困苦給你當水，你的教師卻不再隱藏，你的眼睛必看見你的教師。
ISA|30|21|你或向左或向右，必聽見後邊有聲音說：「這是正路，要行在其間。」
ISA|30|22|你要玷污那雕刻偶像所包的銀子和鑄造偶像所鍍的金子。你要拋棄它們，如拋棄污穢之物；對偶像說：「去吧！」
ISA|30|23|你撒種在地裏，主必降雨在其上，使地所出的糧食肥美豐盛。那時，你的牲畜必在遼闊的草場吃草。
ISA|30|24|耕地的牛和驢必吃加鹽的飼料，是用鏟子和杈子揚淨的。
ISA|30|25|在大行殺戮的日子，城樓倒塌的時候，高山峻嶺必有川河湧流。
ISA|30|26|當耶和華包紮他百姓的傷口，醫治他所擊打傷痕的日子，月光必像日光，日光必加七倍，像七日的光一樣。
ISA|30|27|看哪，耶和華的名從遠方來， 他的怒氣燒起，濃煙上騰。 他的嘴唇滿有憤恨， 他的舌頭像吞滅的火。
ISA|30|28|他的氣息如漲溢的河水，直漲到頸項， 要用毀滅的篩網篩淨列國， 並在眾民口中安放導錯方向的嚼環。
ISA|30|29|你們必唱歌，像守聖節的夜間一樣；並且心中喜樂，像人吹笛，來到耶和華的山，到 以色列 的磐石那裏。
ISA|30|30|耶和華必使人聽見他威嚴的聲音，又以極大的憤怒、吞滅的火焰、雷雨、暴風和像石塊的冰雹，使人看見他降罰的膀臂。
ISA|30|31|亞述 必因耶和華的聲音驚惶，耶和華必用杖擊打它。
ISA|30|32|耶和華必將定規要打 的杖加在它身上；每打一下，都必配合擊鼓彈琴的節奏。打仗時，耶和華必振臂與它交戰。
ISA|30|33|原來 陀斐特 早已預備好了，是為君王預備的；又深又寬，堆滿了火和木柴；耶和華的氣息猶如一股硫磺使它燃起。
ISA|31|1|禍哉！那些下 埃及 求幫助的， 他們仰賴馬匹，倚靠甚多的戰車， 並倚靠強壯的騎兵， 卻不仰望 以色列 的聖者， 也不求問耶和華。
ISA|31|2|其實，耶和華有智慧， 他降災禍， 並不撤回自己的話， 卻要興起攻擊作惡之家， 攻擊那幫助人作惡的。
ISA|31|3|埃及 人不過是人，並非上帝， 他們的馬不過是血肉，並不是靈。 耶和華一伸手， 那幫助人的必絆跌，受幫助的也必跌倒， 都一同滅亡。
ISA|31|4|耶和華對我如此說， 獅子和少壯獅子為獵物而咆哮， 許多牧人被召來攻擊牠， 牠總不因他們的聲音驚惶， 也不因他們的喧嚷退縮； 萬軍之耶和華也必如此 降臨在 錫安 的大小山岡上爭戰。
ISA|31|5|雀鳥盤旋護衛， 萬軍之耶和華也必照樣保護 耶路撒冷 ； 他必保護拯救， 必逾越而搭救。
ISA|31|6|以色列 人哪，要歸向你們嚴重悖逆的那一位！
ISA|31|7|到那日，你們各人要拋棄親手所造、陷自己於罪中的金偶像和銀偶像。
ISA|31|8|亞述 必倒在刀下，並非人的刀； 有刀要將它吞滅，並非人的刀。 它要逃避這刀， 它的年輕人必做苦工。
ISA|31|9|它的磐石必因驚嚇而消失， 它的領袖必因大旗驚惶； 這是那有火在 錫安 、 有爐在 耶路撒冷 的耶和華說的。
ISA|32|1|看哪，必有一位君王憑公義執政， 必有王子藉公平掌權。
ISA|32|2|必有一人如避風港， 如暴風雨的藏身處； 如乾旱地的溪流， 又如乾燥地巨石的陰影。
ISA|32|3|看的人眼睛不再昏花， 聽的人耳朵必留心聽。
ISA|32|4|性急的人懂得分辨， 口吃的人說話流暢。
ISA|32|5|愚頑人不再稱為君子， 流氓不再稱為紳士。
ISA|32|6|因為愚頑人必說愚妄的話， 他的心作惡 ， 行褻瀆的事， 傳播惡言攻擊耶和華， 使飢餓的人仍然飢餓， 口渴的人無水可喝。
ISA|32|7|流氓的手段邪惡， 他圖謀惡計， 用謊言毀滅困苦人； 貧窮人講求公理時， 他也是如此行。
ISA|32|8|君子卻圖謀高尚的事， 他必因高尚的事站立得穩。
ISA|32|9|安逸的婦女啊，起來聽我的聲音！ 無慮的女子啊，側耳聽我的言語！
ISA|32|10|無慮的女子啊，再過一年，你們必顫慄， 因為無葡萄可摘， 也無果實可收。
ISA|32|11|安逸的婦女啊，要戰兢； 無慮的女子啊，要顫慄， 要脫去衣服，赤著身體， 腰束麻布。
ISA|32|12|你們要為美好的田地 和多結果子的葡萄樹捶胸哀哭。
ISA|32|13|刺草和荊棘要長在我百姓的田地上， 長在歡樂城中一切快樂家園上。
ISA|32|14|宮殿必被撇下， 繁華的城必被拋棄， 堡壘和瞭望樓永為洞穴， 成為野驢的樂土， 羊群的草場。
ISA|32|15|等到聖靈從高處澆灌我們， 曠野將變為田園， 田園看似森林。
ISA|32|16|公平要居住在曠野， 公義要安歇在田園。
ISA|32|17|公義的果實是平安， 公義的效果是平靜和安穩，直到永遠。
ISA|32|18|我的百姓要住在平安的居所， 安穩的住處，寧靜的安歇之地。
ISA|32|19|雖有冰雹擊倒樹林， 城也夷為平地；
ISA|32|20|然而你們在水邊撒種， 牧放牛驢的有福了！
ISA|33|1|禍哉！你這未遭毀滅而毀滅人的人， 人未以詭詐待你而你以詭詐待人的人！ 等你行完了毀滅， 自己必被毀滅； 你行完了詭詐， 人必以詭詐待你。
ISA|33|2|耶和華啊，求你施恩給我們， 我們等候你。 求你每早晨作我們的膀臂， 遭難時作我們的拯救。
ISA|33|3|轟然之聲一發出，萬民就奔逃； 你一興起 ，列國就四散。
ISA|33|4|你們的擄物必被斂盡， 有如螞蚱斂盡禾稼； 人為擄物奔走，宛如蝗蟲蹦跳。
ISA|33|5|耶和華受尊崇，居高處， 使公平和公義充滿 錫安 。
ISA|33|6|他是你這世代安定的力量， 豐盛的救恩、 智慧和知識； 敬畏耶和華是 錫安 的至寶。
ISA|33|7|看哪，他們的英雄在外面哀號 ， 求和的使臣在痛哭。
ISA|33|8|大路荒涼，行人止息； 盟約撕毀，見證 被棄， 人也不受尊重。
ISA|33|9|大地悲哀衰殘， 黎巴嫩 羞愧且枯乾， 沙崙 好像曠野， 巴珊 和 迦密 必凋殘。
ISA|33|10|耶和華說： 「現在我要興起， 要高升， 要受尊崇。
ISA|33|11|你們懷的是糠秕，生的是碎秸； 你們的氣息如火吞滅自己。
ISA|33|12|萬民必像燒著的石灰， 又如斬斷的荊棘，在火裏燃燒。」
ISA|33|13|你們遠方的人，當聽我所做的事； 你們近處的人，當承認我的大能。
ISA|33|14|錫安 的罪人都懼怕， 戰兢抓住不敬虔的人。 我們中間有誰能與吞噬的火同住？ 我們中間有誰能與不滅的火共存呢？
ISA|33|15|那行事公義、說話正直、 憎惡欺壓所得之財、 搖手不受賄賂、 掩耳不聽流血的計謀、 閉眼不看邪惡之事的，
ISA|33|16|這人必居高處， 他的保障是磐石的堡壘， 必有糧食賜給他， 飲水也不致斷絕。
ISA|33|17|你必親眼看見君王的榮美， 看見遼闊之地。
ISA|33|18|你的心必回想那些恐怖的事： 「那數算的人在哪裏？ 秤重的人在哪裏？ 數點城樓的又在哪裏呢？」
ISA|33|19|你必不再看見那兇暴的民， 他們嘴唇說艱澀的言語，難以理解； 舌頭結巴，說無意義的話。
ISA|33|20|你要注視 錫安 ，我們守聖節的城！ 你必親眼看見 耶路撒冷 成為安靜的居所， 成為不挪移的帳幕， 橛子永不拔出， 繩索一根也不折斷。
ISA|33|21|在那裏，威嚴的耶和華對我們是寬闊的江河， 其中必沒有搖槳的小船來往， 也沒有巨大的船舶經過。
ISA|33|22|耶和華是審判我們的， 耶和華為我們設立律法； 耶和華是我們的君王， 他必拯救我們。
ISA|33|23|船上的繩索鬆開， 不能穩住桅杆， 也無法揚起船帆。 那時許多擄物被瓜分， 連瘸腿的也能奪走掠物。
ISA|33|24|城內的居民無人說：「我病了」； 城裏居住的百姓，罪孽都蒙赦免。
ISA|34|1|列國啊，要近前來聽！ 萬民哪，要側耳而聽！ 全地和其上所充滿的， 世界和其中所出的，都應當聽！
ISA|34|2|因為耶和華向列國發怒， 向他們的全軍發烈怒， 要將他們滅盡，任人殺戮。
ISA|34|3|被殺的人必被拋棄， 屍首臭氣上騰， 諸山為他們的血所融化。
ISA|34|4|天上萬象都要朽壞， 天被捲起，有如書卷， 其上的萬象盡都衰殘； 如葡萄樹的葉子凋落， 又如無花果樹枯萎一樣。
ISA|34|5|因為我的刀在天上將要顯現 ； 看哪，這刀臨到 以東 和我所詛咒的民， 要施行審判。
ISA|34|6|耶和華的刀沾滿了血， 是用油脂和羔羊、公山羊的血， 並公綿羊腎上的油脂滋潤的； 因為在 波斯拉 有祭物獻給耶和華， 在 以東 地有大屠殺。
ISA|34|7|野牛與他們一起倒下， 牛犢和壯牛也一同倒下。 他們的地被血染遍， 他們的塵土因油脂肥潤。
ISA|34|8|這是耶和華報仇之日， 為 錫安 伸冤的報應之年。
ISA|34|9|它的河水要變為柏油， 塵埃變為硫磺， 大地成為燃燒的柏油，
ISA|34|10|晝夜總不熄滅， 它的煙永遠上騰， 必世世代代成為荒廢， 永永遠遠無人經過。
ISA|34|11|鵜鶘、豪豬要得它為業， 貓頭鷹、烏鴉要住在其間。 耶和華必將空虛的準繩、 混沌的石垂線，拉在 以東 之上。
ISA|34|12|人必宣稱那裏沒有王國， 它的貴族和所有領袖都歸於無有。
ISA|34|13|以東 的宮殿要長出荊棘， 城堡要生長蒺藜和刺草； 成為野狗的住處， 鴕鳥的居所。
ISA|34|14|野獸要和土狼相遇， 山羊鬼魔要與同伴對唱， 莉莉絲 必在那裏棲身， 為自己尋找安歇之處。
ISA|34|15|箭頭蛇要在那裏做窩， 下蛋，孵蛋，並招聚幼蛇在其保護之下； 鷂鷹也與伴侶聚集在那裏。
ISA|34|16|你們要查考並誦讀耶和華的書； 這些現象必然存在， 沒有一樣動物缺少伴侶。 因為是他，藉著我的口 吩咐， 他的靈將牠們聚集。
ISA|34|17|他為牠們抽籤， 親手用準繩為牠們分地； 直到牠們永遠得地為業， 世世代代住在其間。
ISA|35|1|曠野和乾旱之地必然歡喜， 沙漠也必快樂； 又如玫瑰綻放，
ISA|35|2|朵朵繁茂， 其樂融融，而且歡呼。 黎巴嫩 的榮耀， 並 迦密 與 沙崙 的華美，必賜給它。 人要看見耶和華的榮耀， 看見我們上帝的榮美。
ISA|35|3|你們要使軟弱的手強壯， 使無力的膝蓋穩固；
ISA|35|4|對心裏焦急的人說： 「要剛強，不要懼怕。 看哪，你們的上帝要來施報， 要施行極大的報應， 他必來拯救你們。」
ISA|35|5|那時，盲人的眼必睜開， 聾子的耳必開通。
ISA|35|6|那時，瘸子必跳躍如鹿， 啞巴的舌頭必歡呼。 在曠野有水噴出， 在沙漠有江河湧流。
ISA|35|7|火熱之地要變為水池， 乾渴之地要變為泉源。 野狗躺臥休息之處 必長出青草、蘆葦和蒲草。
ISA|35|8|在那裏必有一條大道， 就是一條路 ，稱為聖路。 污穢的人不得經過， 是專為走路的人 預備的， 愚昧的人也不會迷路。
ISA|35|9|在那裏沒有獅子， 猛獸也不經過； 在那裏牠們未現蹤跡， 只有救贖的民在那裏行走。
ISA|35|10|耶和華救贖的民必歸回， 歌唱來到 錫安 ； 永遠的快樂必歸到他們頭上， 他們必得著歡喜快樂， 憂傷嘆息盡都逃避。
ISA|36|1|希西家 王十四年， 亞述 王 西拿基立 上來攻擊 猶大 的一切堅固的城，將城攻取。
ISA|36|2|亞述 王從 拉吉 差遣將軍 率領大軍前往 耶路撒冷 ，到 希西家 王那裏去。將軍站在 上池 的水溝旁，在往漂布地的大路上。
ISA|36|3|希勒家 的兒子 以利亞敬 宮廷總管、 舍伯那 書記和 亞薩 的兒子 約亞 史官，出來見他。
ISA|36|4|將軍對他們說：「你們去告訴 希西家 ，大王 亞述 王如此說：『你倚靠甚麼，讓你如此自信滿滿？
ISA|36|5|我說 ，你有打仗的計謀和能力，我看不過是空話。你到底倚靠誰，竟敢背叛我呢？
ISA|36|6|看哪，你所倚靠的 埃及 是那斷裂的葦杖，人若倚靠這杖，它就刺進他的手，穿透它。 埃及 王法老向所有倚靠他的人都是這樣。
ISA|36|7|你若對我說：我們倚靠耶和華－我們的上帝， 希西家 豈不是將上帝的丘壇和祭壇廢去，並且吩咐 猶大 和 耶路撒冷 的人說：你們只當在這一個壇前敬拜嗎？
ISA|36|8|現在你與我主 亞述 王打賭，我給你兩千匹馬，看你能否派得出騎士來騎牠們。
ISA|36|9|若不然，怎能使我主臣僕中最小的一個軍官轉臉而逃呢？你難道要倚靠 埃及 的戰車和騎兵嗎？
ISA|36|10|現在我上來攻擊毀滅這地，豈不是出於耶和華嗎？耶和華吩咐我說，你上去攻擊這地，毀滅它吧！』」
ISA|36|11|以利亞敬 、 舍伯那 、 約亞 對將軍說：「求你用 亞蘭 話對僕人說，因為我們聽得懂；不要用 猶大 話對我們說，免得傳到城牆上百姓的耳中。」
ISA|36|12|將軍說：「我主差遣我來，豈是單對你和你的主人說這些話嗎？不也是對這些坐在城牆上，要與你們一同吃自己糞、喝自己尿的人說的嗎？」
ISA|36|13|於是 亞述 將軍站著，用 猶大 話大聲喊著說：「你們當聽大王 亞述 王的話，
ISA|36|14|王如此說：『你們不要被 希西家 欺哄了，因他不能拯救你們。
ISA|36|15|不要聽憑 希西家 說服你們倚靠耶和華，他說，耶和華必要拯救我們，這城必不交在 亞述 王的手中。』
ISA|36|16|你們不要聽 希西家 的話！因 亞述 王如此說：『你們要與我講和，出來投降，各人就可以吃自己葡萄樹和無花果樹的果子，喝自己井裏的水，
ISA|36|17|等我來領你們到一個地方，與你們本地一樣，就是有五穀和新酒之地，有糧食和葡萄園之地。
ISA|36|18|恐怕 希西家 誤導你們說，耶和華必拯救我們。列國的神明有哪一個曾救它本國脫離 亞述 王的手呢？
ISA|36|19|哈馬 和 亞珥拔 的神明在哪裏呢？ 西法瓦音 的神明在哪裏呢？它們曾救 撒瑪利亞 脫離我的手嗎？
ISA|36|20|這些國的神明有誰曾救自己的國家脫離我的手呢？難道耶和華能救 耶路撒冷 脫離我的手嗎？』」
ISA|36|21|百姓靜默不言，一句不答，因為 希西家 王曾吩咐說：「不要回答他。」
ISA|36|22|當下 希勒家 的兒子 以利亞敬 宮廷總管、 舍伯那 書記，和 亞薩 的兒子 約亞 史官都撕裂衣服，來到 希西家 那裏，將 亞述 將軍的話告訴他。
ISA|37|1|希西家 王聽見了，就撕裂衣服，披上麻布，進了耶和華的殿。
ISA|37|2|他差遣 以利亞敬 宮廷總管和 舍伯那 書記，並祭司中年長的，都披上麻布，到 亞摩斯 的兒子 以賽亞 先知那裏去。
ISA|37|3|他們對他說：「 希西家 如此說：『今日是急難、懲罰、凌辱的日子，就如嬰孩快要出生，卻沒有力氣生產。
ISA|37|4|或許耶和華－你的上帝聽見 亞述 將軍的話，就是他主人 亞述 王差他來辱罵永生上帝的話，耶和華－你的上帝就斥責所聽見的這些話。求你為倖存的餘民揚聲禱告。』」
ISA|37|5|希西家 王的臣僕就來到 以賽亞 那裏。
ISA|37|6|以賽亞 對他們說：「要對你們的主人這樣說，耶和華如此說：『你聽見 亞述 王的僕人褻瀆我的話，不要懼怕。
ISA|37|7|看哪，因為我必驚動他的心 ，他要聽見風聲就歸回本地，在那裏我必使他倒在刀下。』」
ISA|37|8|亞述 將軍聽見 亞述 王已拔營離開 拉吉 ，就啟程返回，正遇見 亞述 王去攻打 立拿 。
ISA|37|9|亞述 王聽見有人談論 古實 王 特哈加 說：「他出來要與你爭戰。」 亞述 王一聽見，就差使者去見 希西家 ，說：
ISA|37|10|「你們要對 猶大 王 希西家 如此說：『不要聽你所倚靠的上帝欺哄你說： 耶路撒冷 必不交在 亞述 王的手中。
ISA|37|11|看哪，你總聽說 亞述 諸王向列國所行的是盡行滅絕，難道你能倖免嗎？
ISA|37|12|我祖先所毀滅的，就是 歌散 、 哈蘭 、 利色 和 提‧拉撒 的 伊甸 人；這些國的神明何曾拯救他們呢？
ISA|37|13|哈馬 的王， 亞珥拔 的王， 西法瓦音城 的王， 希拿 和 以瓦 的王，都在哪裏呢？』」
ISA|37|14|希西家 從使者手裏接過書信，看完了，就上耶和華的殿，在耶和華面前展開書信。
ISA|37|15|希西家 向耶和華禱告說：
ISA|37|16|「坐在基路伯之上萬軍之耶和華－ 以色列 的上帝啊，你，惟有你是地上萬國的上帝，你創造了天和地。
ISA|37|17|耶和華啊，求你側耳而聽；耶和華啊，求你睜眼而看，聽 西拿基立 差遣使者辱罵永生上帝的一切話。
ISA|37|18|耶和華啊， 亞述 諸王果然使列國和列國之地變為荒蕪，
ISA|37|19|將列國的神明扔在火裏，因為它們不是神明，是人手所造的，是木頭、石頭，所以被滅絕了。
ISA|37|20|耶和華－我們的上帝啊，現在求你救我們脫離 亞述 王的手，使地上萬國都知道惟有你是耶和華。」
ISA|37|21|亞摩斯 的兒子 以賽亞 就差人去見 希西家 ，說：「耶和華－ 以色列 的上帝如此說，你因 亞述 王 西拿基立 的事向我祈求，
ISA|37|22|所以耶和華論他這樣說： 『少女 錫安 藐視你，嘲笑你； 耶路撒冷 向你搖頭。
ISA|37|23|「『你辱罵誰，褻瀆誰， 揚起聲來，高舉眼目攻擊誰呢？ 你攻擊的是 以色列 的聖者。
ISA|37|24|你藉臣僕辱罵主說： 我率領許多戰車登上高山， 到 黎巴嫩 的頂端； 我要砍伐其中高大的香柏樹 和上好的松樹。 我必上到極高之處， 進入茂盛的森林裏。
ISA|37|25|我已經挖井喝水 我必用腳掌踏乾 埃及 一切的河流。
ISA|37|26|「『你豈沒有聽見 我早先所定、古時所立、現今實現的事嗎？ 就是讓你去毀壞堅固的城鎮，使它們變為廢墟；
ISA|37|27|城裏居民的力量甚小， 他們驚惶羞愧； 像野草，像青菜， 如房頂上的草， 被東風颳散 。
ISA|37|28|「『你站起，你坐下，你出去，你進來， 你向我發烈怒，我都知道。
ISA|37|29|因你向我發烈怒， 你的狂傲上達我耳中， 我要用鉤子鉤住你的鼻子， 將嚼環放在你口裏， 使你從原路轉回去。』
ISA|37|30|「我賜給你的預兆：你們今年要吃野生的，明年也要吃自長的；後年，你們就要耕種收割，栽葡萄園，吃其中的果子。
ISA|37|31|猶大 家所逃脫剩餘的，仍要往下扎根，向上結果。
ISA|37|32|必有剩餘的民從 耶路撒冷 而出；有逃脫的人從 錫安山 而來。萬軍之耶和華的熱心必成就這事。
ISA|37|33|「所以耶和華論 亞述 王如此說：他必不得來到這城，也不在這裏射箭，不得拿盾牌到城前，也不能建土堆攻城。
ISA|37|34|他從哪條路來，必從那條路回去，必不得來到這城。這是耶和華說的。
ISA|37|35|因我為自己的緣故，又為我僕人 大衛 的緣故，必保護拯救這城。」
ISA|37|36|耶和華的使者出去，在 亞述 營中殺了十八萬五千人。清早有人起來，看哪，都是死屍。
ISA|37|37|亞述 王 西拿基立 就拔營回去，住在 尼尼微 。
ISA|37|38|一日，他在他的神明 尼斯洛 廟裏叩拜，他兒子 亞得米勒 和 沙利色 用刀殺了他，然後逃到 亞拉臘 地；他兒子 以撒．哈頓 接續他作王。
ISA|38|1|那些日子， 希西家 病得要死， 亞摩斯 的兒子 以賽亞 先知來見他，對他說：「耶和華如此說：『你當留遺囑給你的家，因為你必死，不能活了。』」
ISA|38|2|希西家 就轉臉朝牆，向耶和華禱告，
ISA|38|3|說：「耶和華啊，求你記念我在你面前怎樣存完全的心，按誠實行事，又做你眼中看為善的事。」 希西家 就痛哭。
ISA|38|4|耶和華的話臨到 以賽亞 說：
ISA|38|5|「你去告訴 希西家 說，耶和華－你祖先 大衛 的上帝如此說：『我聽見了你的禱告，看見了你的眼淚。看哪，我必加添你十五年的壽數；
ISA|38|6|我要救你和這城脫離 亞述 王的手，也要保護這城。』
ISA|38|7|「耶和華必成就他所說的這話。這是耶和華給你的預兆：
ISA|38|8|看哪，我要使 亞哈斯 日晷上隨太陽前進的影子，往後退十度。」於是，在日晷上照下來的日影果然往後退了十度。
ISA|38|9|猶大 王 希西家 患病痊癒後的詩：
ISA|38|10|我說，在如日中天的時候我就走了， 將剩餘的年歲交給陰間的門。
ISA|38|11|我說，我必不得見耶和華，不得在活人之地見耶和華， 也不再看見世人，就是短暫世界 中的居民。
ISA|38|12|我的住處好像牧人的帳棚， 遭人掀起，離我而去； 我將性命捲起， 像織布的捲布一樣。 他從織布機頭那裏將我剪斷， 你使我命喪於旦夕。
ISA|38|13|我令自己安靜 直到天亮； 他像獅子折斷我所有的骨頭， 你使我命喪於旦夕。
ISA|38|14|我像燕子呢喃， 像白鶴鳴叫， 又如鴿子哀鳴； 我因仰望，眼睛困倦。 主啊，我受欺壓， 求你為我作保。
ISA|38|15|我還有甚麼可說的呢？ 他應許我的 ，他已成就了。 我因心裏的苦楚， 在一生的年日必謙卑而行 。
ISA|38|16|主啊，人得存活是在乎此， 我的靈存活也全在乎此 ； 求你使我痊癒，仍然存活。
ISA|38|17|看哪，我受大苦是為使我得平安； 你愛我，救我的性命脫離敗壞的地府， 將我一切的罪扔在你背後。
ISA|38|18|原來，陰間不能稱謝你， 死亡不能頌揚你， 下到地府的人也不能盼望你的信實。
ISA|38|19|只有活人，活人必稱謝你， 像我今日稱謝你一樣。 為父的，必使兒女知道你的信實。
ISA|38|20|耶和華肯救我， 所以，我們要一生一世 在耶和華殿中 彈奏我弦樂的歌。
ISA|38|21|以賽亞 說：「拿一塊無花果餅來，貼在瘡上，王必痊癒。」
ISA|38|22|希西家 說：「我能上耶和華的殿，有甚麼預兆呢？」
ISA|39|1|那時， 巴拉但 的兒子， 巴比倫 王 米羅達‧巴拉但 聽見 希西家 病得痊癒，就送書信和禮物給他。
ISA|39|2|希西家 歡喜見使者，就將自己寶庫裏的金子、銀子、香料、貴重的膏油和他軍械庫裏一切的兵器，以及他所有的財寶，都給他們看；在他家中和全國之內， 希西家 沒有一樣不給他們看的。
ISA|39|3|於是 以賽亞 先知到 希西家 王那裏去，對他說：「這些人說了些甚麼？他們從哪裏來見你？」 希西家 說：「他們從遠方的 巴比倫 來見我。」
ISA|39|4|以賽亞 說：「他們在你家裏看見了甚麼？」 希西家 說：「凡我家中所有的，他們都看見了；我財寶中沒有一樣東西不給他們看的。」
ISA|39|5|以賽亞 對 希西家 說：「你要聽萬軍之耶和華的話，
ISA|39|6|耶和華說：『看哪，日子將到，凡你家裏所有的，並你祖先積蓄到如今的一切，都要被擄到 巴比倫 去，不留下一樣；
ISA|39|7|從你本身所生的孩子，其中必有被擄到 巴比倫 王宮當太監的。』」
ISA|39|8|希西家 對 以賽亞 說：「你所說耶和華的話甚好。」因為他想：「在我有生之年必有太平和安穩。」
ISA|40|1|你們的上帝說： 「要安慰，安慰我的百姓。
ISA|40|2|要對 耶路撒冷 說安慰的話， 向它宣告， 它的戰爭已結束， 它的罪孽已赦免； 它為自己一切的罪， 已從耶和華手中加倍受罰。」
ISA|40|3|有聲音呼喊著： 「要在曠野為耶和華預備道路， 在沙漠為我們的上帝修直大道。
ISA|40|4|一切山窪都要填滿， 大小山岡都要削平； 陡峭的要變為平坦， 崎嶇的必成為平原。
ISA|40|5|耶和華的榮耀必然顯現， 凡有血肉之軀的都一同看見， 因為這是耶和華親口說的。」
ISA|40|6|有聲音說：「你喊叫吧！」 我 說：「我喊叫甚麼呢？」 凡有血肉之軀的盡都如草， 他的一切榮美像野地的花。
ISA|40|7|耶和華吹一口氣， 草就枯乾，花也凋謝。 百姓誠然是草；
ISA|40|8|草必枯乾，花必凋謝， 惟有我們上帝的話永遠立定。
ISA|40|9|報好信息的 錫安 哪， 要登高山； 報好信息的 耶路撒冷 啊， 要極力揚聲。 揚聲不要懼怕， 對 猶大 的城鎮說： 「看哪，你們的上帝！」
ISA|40|10|看哪，主耶和華必以大能臨到， 他的膀臂必為他掌權； 看哪，他的賞賜在他那裏， 他的報應在他面前。
ISA|40|11|他要像牧人牧養自己的羊群， 用膀臂聚集羔羊，抱在胸懷， 慢慢引導那乳養小羊的。
ISA|40|12|誰曾用手心量諸水， 用手虎口量蒼天， 用升斗盛大地的塵土， 用秤稱山嶺， 用天平稱岡陵呢？
ISA|40|13|誰曾測度耶和華的靈， 或作他的謀士指教他呢？
ISA|40|14|他與誰商議， 誰教導他， 以公平的路指示他， 將知識傳授與他， 又將通達的道指教他呢？
ISA|40|15|看哪，列國都像水桶裏的一滴， 又如天平上的微塵； 看哪，他舉起眾海島，好像舉起極微小之物。
ISA|40|16|黎巴嫩 不夠當柴燒， 其中的走獸也不夠作燔祭。
ISA|40|17|列國在他面前如同不存在， 在他看來微不足道，只是虛空。
ISA|40|18|你們究竟將誰比上帝， 用甚麼形像與他相較呢？
ISA|40|19|至於偶像，匠人鑄造它， 銀匠用金子包裹它， 又為它鑄造銀鏈。
ISA|40|20|沒有能力捐獻的人， 就挑選不易朽壞的木頭， 為自己尋找巧匠， 豎立不會倒的偶像。
ISA|40|21|你們豈不知道嗎？ 豈未曾聽見嗎？ 難道沒有人從起頭就告訴你們嗎？ 自從地的根基立定， 你們豈不明白嗎？
ISA|40|22|上帝坐在地的穹窿之上， 地上的居民有如蚱蜢。 他鋪張穹蒼如幔子， 展開諸天如可住的帳棚。
ISA|40|23|他使君王歸於虛無， 使地上的審判官成為虛空。
ISA|40|24|他們剛栽上， 剛種好， 根也剛扎在地裏， 經他一吹，就都枯乾； 旋風將他們吹去，像碎秸一樣。
ISA|40|25|那聖者說：「你們將誰與我相比， 與我相等呢？」
ISA|40|26|你們要向上舉目， 看是誰創造這萬象， 按數目領出它們， 一一稱其名， 以他的權能 和他的大能大力， 使它們一個都不缺。
ISA|40|27|雅各 啊，你為何說， 以色列 啊，你為何言， 「我的道路向耶和華隱藏， 我的冤屈上帝並不查問」？
ISA|40|28|你豈不曾知道嗎？ 你豈未曾聽見嗎？ 永在的上帝耶和華，創造地極的主， 他不疲乏，也不困倦； 他的智慧無法測度。
ISA|40|29|疲乏的，他賜能力； 軟弱的，他加力量。
ISA|40|30|就是年輕人也要疲乏困倦， 強壯的也必全然跌倒。
ISA|40|31|但那等候耶和華的必重新得力。 他們必如鷹展翅上騰； 他們奔跑卻不困倦， 行走卻不疲乏。
ISA|41|1|眾海島啊，在我面前靜默； 萬民要重新得力， 讓他們近前來陳述， 我們可以彼此辯論。
ISA|41|2|誰從東方興起一人， 憑公義召他來到腳前？ 誰將列國交給他， 使他管轄列王， 把他們如灰塵交與他的刀， 如風吹的碎秸交與他的弓？
ISA|41|3|他追趕君王， 安然走過， 快速地腳不落地 。
ISA|41|4|誰做成這事， 從起初宣召歷代呢？ 就是我－耶和華！ 我是首先的， 也與末後的同在。
ISA|41|5|眾海島看見就都害怕， 地極也都戰兢， 他們近前來；
ISA|41|6|各人互相幫助， 對弟兄說：「壯膽吧！」
ISA|41|7|木匠鼓勵銀匠， 用鎚子打光的鼓勵打砧的， 對銲工說：「銲得好！」 又用釘子釘穩，免得它倒下。
ISA|41|8|惟你 以色列 ，我的僕人， 雅各 ，我所揀選的， 我朋友 亞伯拉罕 的後裔，
ISA|41|9|你是我從地極領來， 從地角召來的， 我對你說：「你是我的僕人； 我揀選你，並不棄絕你。」
ISA|41|10|你不要害怕，因為我與你同在； 不要驚惶，因為我是你的上帝。 我必堅固你，幫助你， 用我公義的右手扶持你。
ISA|41|11|看哪，凡向你發怒的都抱愧蒙羞， 與你相爭的必如無有，並要滅亡。
ISA|41|12|與你爭鬥的，你要尋找他們，卻遍尋不著； 與你爭戰的必如無有，成為虛無。
ISA|41|13|因為我耶和華－你的上帝 必攙扶你的右手， 對你說：「不要害怕！ 我必幫助你。」
ISA|41|14|蟲子 雅各 ， 以色列 人哪， 不要害怕！ 我必幫助你； 救贖你的是 以色列 的聖者。 這是耶和華說的。
ISA|41|15|看哪，我使你成為 全新的打穀機，齒輪銳利； 你要把山嶺打得粉碎， 使岡陵如同糠秕。
ISA|41|16|你要簸揚它們，風要將它們吹去； 旋風要颳散它們。 你卻要以耶和華為喜樂， 因 以色列 的聖者誇耀。
ISA|41|17|困苦貧窮人尋找水，卻尋不著； 他們因口渴，舌頭乾燥。 我－耶和華必應允他們， 我─ 以色列 的上帝必不離棄他們。
ISA|41|18|我要在光禿的高地開江河， 在谷中開泉源； 我要使沙漠變為水池， 使乾地變為湧泉。
ISA|41|19|我要在曠野栽植香柏樹、 皂莢樹、番石榴樹，和野橄欖樹。 在沙漠一同栽上松樹、杉樹， 和黃楊樹，
ISA|41|20|好叫人看見，知道， 思想，明白； 這是耶和華親手做的， 是 以色列 的聖者所造的。
ISA|41|21|耶和華說： 「你們要呈上你們的案件。」 雅各 的君王說： 「你們要提出你們的理由。」
ISA|41|22|讓它們近前來，告訴我們將來要發生甚麼事！ 你們要說明先前發生的事，好讓我們思索； 或者告訴我們將來的事，使我們得知事情的結局。
ISA|41|23|你們要指明未來的事， 使我們知道你們是神明！ 你們或降福，或降禍， 好使我們驚奇，一同觀看。
ISA|41|24|看哪，你們屬乎虛無， 你們的作為也屬虛空； 那選擇你們的是可憎惡的。
ISA|41|25|我從北方興起一人， 他從日出之地而來， 是求告我名的； 他必踩踏 掌權者，如踩踏泥土， 又如陶匠踹泥一般。
ISA|41|26|有誰從起初宣佈這事，使我們知道呢？ 有誰從先前指明，使我們說「他是對的」呢？ 沒有人宣佈， 沒有人指明， 也沒有人聽見你們的話。
ISA|41|27|我首先對 錫安 說，看哪，他們在此！ 我要將一位報好信息的賜給 耶路撒冷 。
ISA|41|28|然而我觀看，並無一人； 我詢問的時候， 他們中間也沒有謀士可回答。
ISA|41|29|看哪，他們盡是麻煩 ， 所做的工都屬虛無； 所鑄的偶像是風，是虛空。
ISA|42|1|看哪，我的僕人， 我所扶持、所揀選、心所喜悅的！ 我已將我的靈賜給他， 他必將公理傳給萬邦。
ISA|42|2|他不喧嚷，不揚聲， 也不使街上聽見他的聲音。
ISA|42|3|壓傷的蘆葦，他不折斷； 將殘的燈火，他不吹滅。 他憑信實將公理傳開。
ISA|42|4|他不灰心，也不喪膽， 直到他在地上設立公理； 眾海島都等候他的訓誨。
ISA|42|5|那創造諸天，鋪張穹蒼， 鋪開地與地的出產， 賜氣息給地上眾人， 賜生命給行走其上之人的 上帝耶和華如此說：
ISA|42|6|「我－耶和華憑公義召你， 要攙扶你的手，保護你， 要藉著你與百姓立約， 使你成為萬邦之光，
ISA|42|7|開盲人的眼， 領囚犯出監獄， 領坐在黑暗中的出地牢。
ISA|42|8|我是耶和華，這是我的名； 我必不將我的榮耀歸給別神 ， 也不將我所得的頌讚歸給雕刻的偶像。
ISA|42|9|看哪，先前的事已經成就， 現在我要指明新事， 告訴你們尚未發生的事。
ISA|42|10|航海的人和海中一切所有的， 眾海島和其中的居民， 都當向耶和華唱新歌， 從地極讚美他。
ISA|42|11|曠野和其中的城鎮， 並 基達 人居住的村莊都當揚聲 ； 西拉 的居民當歡呼， 在山頂上大聲呼喊。
ISA|42|12|願他們將榮耀歸給耶和華， 在海島中傳揚頌讚他的話。
ISA|42|13|耶和華必如勇士出征， 如戰士激起憤恨， 他要喊叫，大聲吶喊， 擊敗他的敵人。
ISA|42|14|我許久閉口不言，沉默不語； 現在我要像臨產的婦人，大聲喊叫， 呼吸急促而喘氣。
ISA|42|15|我要使大小山岡變為荒蕪， 使其上的花草都枯乾； 我要使江河變為沙洲， 使水池盡都乾涸。
ISA|42|16|我要引導盲人行他們所不認識的道， 引領他們走他們未曾走過的路； 我在他們面前使黑暗變為光明， 使彎曲變為平直。 這些事我都要做， 並不離棄他們。
ISA|42|17|但那倚靠雕刻的偶像， 對鑄造的偶像說： 「你是我們的神明」； 這種人要退後，大大蒙羞。
ISA|42|18|你們這耳聾的，聽吧！ 你們這眼瞎的，看吧， 使你們得以看見！
ISA|42|19|誰比我的僕人眼瞎呢？ 誰比我所差遣的使者耳聾呢？ 誰瞎眼像那獻身給我的人？ 誰瞎眼 像耶和華的僕人呢？
ISA|42|20|看見許多事卻不領會， 耳朵開通卻聽不見。
ISA|42|21|耶和華因自己的公義， 樂意使律法為大為尊。
ISA|42|22|但這百姓是被搶被奪的， 全都陷在洞穴中，關在監牢裏； 他們成了掠物，無人拯救， 成了擄物，無人索還。
ISA|42|23|你們中間誰肯側耳聽這話， 誰肯留心聽，以防將來呢？
ISA|42|24|誰將 雅各 交出作為擄物， 將 以色列 交給搶奪者呢？ 豈不是耶和華 ─我們所得罪的那位嗎？ 他們不肯遵行他的道， 也不聽從他的訓誨。
ISA|42|25|所以，他將猛烈的怒氣和戰爭的威力 傾倒在 以色列 身上； 在他周圍如火燃起，他竟然不知， 燒著了，他也不在意。
ISA|43|1|雅各 啊，創造你的耶和華， 以色列 啊，造成你的那位， 現在如此說： 「你不要害怕，因為我救贖了你； 我曾提你的名召你，你是屬我的。
ISA|43|2|你從水中經過，我必與你同在， 你渡過江河，水必不漫過你； 你在火中行走，也不被燒傷， 火焰必不燒著你身。
ISA|43|3|因為我是耶和華－你的上帝， 是 以色列 的聖者－你的救主； 我使 埃及 作你的贖價， 使 古實 和 西巴 代替你。
ISA|43|4|因我看你為寶貝為尊貴； 又因我愛你， 所以使人代替你， 使萬民替換你的生命。
ISA|43|5|你不要害怕，因我與你同在； 我必領你的後裔從東方來， 又從西方召集你。
ISA|43|6|我要對北方說，交出來！ 對南方說，不可扣留！ 要將我的兒子從遠方帶來， 將我的女兒從地極領回，
ISA|43|7|就是凡稱為我名下的人， 是我為自己的榮耀創造的， 是我所塑造，所做成的。」
ISA|43|8|你要將有眼卻瞎、 有耳卻聾的民都帶出來！
ISA|43|9|任憑萬國聚集， 任憑萬民會合。 他們當中誰能說明， 並將先前的事指示我們呢？ 讓他們帶來見證，顯明他們有理， 看是否聽見的人會說：「果然是真的。」
ISA|43|10|你們是我的見證， 是我所揀選的僕人， 為了要使你們知道，且信服我， 又明白我就是耶和華。 在我以前沒有任何被造的真神， 在我以後也必沒有。 這是耶和華說的。
ISA|43|11|我，惟有我是耶和華； 除我以外沒有救主。
ISA|43|12|我曾指示，我曾拯救，我曾說明， 並沒有外族的神明 在你們中間。 你們是我的見證， 我是上帝。 這是耶和華說的。
ISA|43|13|自有日子以來，我就是上帝， 誰也不能救人脫離我的手。 我要行事，誰能逆轉呢？
ISA|43|14|耶和華─你們的救贖主、 以色列 的聖者如此說： 「因你們的緣故， 我已派遣人到 巴比倫 去； 要使 迦勒底 人都如難民， 坐自己素來宴樂的船下來。
ISA|43|15|我是耶和華－你們的聖者， 是創造 以色列 的，是你們的君王。」
ISA|43|16|那在滄海中開道， 在大水中開路， 使戰車、馬匹、軍兵、勇士一同出來， 使他們仆倒，不再起來， 使他們滅沒，好像熄滅之燈火的耶和華如此說：
ISA|43|17|
ISA|43|18|「你們不要追念從前的事， 也不要思想古時的事。
ISA|43|19|看哪，我要行一件新事， 如今就要顯明，你們豈不知道嗎？ 我必在曠野開道路， 在沙漠開江河 。
ISA|43|20|野地的走獸要尊敬我， 野狗和鴕鳥也必尊敬我。 因我使曠野有水， 使沙漠有河， 好賜給我的百姓、我的選民喝。
ISA|43|21|這百姓是我為自己造的， 為要述說我的美德。」
ISA|43|22|「 雅各 啊，你並沒有求告我； 以色列 啊，你倒厭煩我。
ISA|43|23|你並沒有將你的羊帶來獻給我做燔祭， 也沒有用牲祭尊敬我； 我未曾因素祭使你操勞， 也沒有因乳香使你厭煩。
ISA|43|24|你沒有用銀子為我買香菖蒲， 也沒有用祭物的油脂使我飽足； 倒使我因你的罪惡操勞， 使我因你的罪孽厭煩。
ISA|43|25|我，惟有我為自己的緣故塗去你的過犯， 我也不再記得你的罪惡。
ISA|43|26|你儘管提醒我，讓我們來辯論； 儘管陳述，自顯為義。
ISA|43|27|你的始祖犯罪， 你的師傅違背我；
ISA|43|28|因此，我要凌辱聖所的領袖 ， 使 雅各 遭毀滅， 使 以色列 受辱罵。」
ISA|44|1|「我的僕人 雅各 ， 我所揀選的 以色列 啊， 現在你當聽。
ISA|44|2|那位造你，使你在母腹中成形， 並要幫助你的耶和華如此說： 我的僕人 雅各 ， 我所揀選的 耶書崙 哪， 不要害怕！
ISA|44|3|因為我要把水澆灌乾渴的地方， 使水湧流在乾旱之地。 我要將我的靈澆灌你的後裔， 使我的福臨到你的子孫。
ISA|44|4|他們要在草叢中生長 ， 如溪水旁的柳樹。
ISA|44|5|這個要說：『我是屬耶和華的』， 那個要以 雅各 的名自稱， 又有一個在手上寫著：『歸耶和華』， 並自稱為 以色列 。」
ISA|44|6|耶和華－ 以色列 的君王， 以色列 的救贖主－萬軍之耶和華如此說： 「我是首先的，也是末後的； 除我以外再沒有上帝。
ISA|44|7|自從古時我設立了人， 誰能像我宣告，指明，又為自己陳說呢？ 讓他指明未來的事和必成的事吧！
ISA|44|8|你們不要恐懼，也不要害怕。 我豈不是從上古就告訴並指示你們了嗎？ 你們是我的見證人！ 除我以外，豈有上帝呢？ 誠然沒有磐石，就我所知，一個也沒有！」
ISA|44|9|製造偶像的人盡都虛空，他們所喜悅的全無益處；偶像的見證人毫無所見，毫無所知，以致他們羞愧。
ISA|44|10|誰製造神像，鑄造偶像？這些都是無益的。
ISA|44|11|看哪，他的同夥都必羞愧。工匠不過是人，任他們聚集，任他們站立吧！他們都必懼怕，一同羞愧。
ISA|44|12|鐵匠用工具在火炭上工作 ，用鎚打出形狀，用他有力的膀臂來錘。他因飢餓而無力氣；因未喝水而疲倦。
ISA|44|13|木匠拉線，用筆劃出樣子，用鉋子鉋成形狀，又用圓規劃了模樣。他仿照人的體態，做出美妙的人形，放在廟裏。
ISA|44|14|他砍伐香柏樹，又取杉樹和橡樹，在樹林中讓它茁壯；或栽種松樹，得雨水滋潤長大。
ISA|44|15|這樹，人可用以生火；他拿一些來取暖，又搧火烤餅，而且做神像供跪拜，做雕刻的偶像向它叩拜。
ISA|44|16|他將一半的木頭燒在火中，用它烤肉來吃；吃飽了，就自己取暖說：「啊哈，我暖和了，我看到火了！」
ISA|44|17|然後又用剩下的一半做了一個神明，就是雕刻的偶像，向這偶像俯伏叩拜，向它禱告說：「求你拯救我，因你是我的神明。」
ISA|44|18|他們既無知，又不思想；因為耶和華蒙蔽他們的眼，使他們看不見，塞住他們的心，使他們不明白。
ISA|44|19|沒有一個心裏醒悟，有知識，有聰明，能說：「我曾拿一部分用火燃燒，在炭火上烤餅，也烤肉來吃。這剩下的，我豈要做可憎之像嗎？我豈可向木頭叩拜呢？」
ISA|44|20|他以灰塵為食，心裏迷糊，以致偏邪，不能自救，也不能說：「我右手中豈不是有虛謊嗎？」
ISA|44|21|雅各 啊，要思念這些事； 以色列 啊，你是我的僕人。 我造了你，你是我的僕人， 以色列 啊，我必不忘記你 。
ISA|44|22|我塗去你的過犯，像厚雲消散； 塗去你的罪惡，如薄霧消失。 你當歸向我，因我救贖了你。
ISA|44|23|諸天哪，應當歌唱， 因為耶和華成就這事。 地的深處啊，應當歡呼； 眾山哪，要出聲歌唱； 樹林和其中所有的樹木啊，你們都當歌唱！ 因為耶和華救贖了 雅各 ， 並要因 以色列 榮耀自己。
ISA|44|24|從你在母腹中就造了你，你的救贖主－耶和華如此說： 「我－耶和華創造萬物， 獨自鋪張諸天，親自展開大地 ；
ISA|44|25|我使虛謊的預兆失效， 愚弄占卜的人， 使智慧人退後， 使他的知識變為愚拙；
ISA|44|26|卻使我僕人的話站得住， 成就我使者的籌算。 我論 耶路撒冷 說：『必有人居住』； 論 猶大 的城鎮說：『必被建造， 我必重建其中的廢墟。』
ISA|44|27|我對深淵說：『乾了吧！ 我要使你的江河乾涸』；
ISA|44|28|論 居魯士 說：『他是我的牧人， 他要成就我所喜悅的， 下令建造 耶路撒冷 ， 發命令立穩聖殿的根基。』」
ISA|45|1|耶和華對所膏的 居魯士 如此說， 他的右手我曾攙扶， 使列國降服在他面前， 列王的腰帶我曾鬆開， 使城門在他面前敞開， 不得關閉：
ISA|45|2|「我要在你前面行， 修平崎嶇之地。 我必打破銅門， 砍斷鐵閂。
ISA|45|3|我要將暗中的寶物和隱藏的財富賜給你， 使你知道提名召你的 就是我－耶和華， 以色列 的上帝。
ISA|45|4|因我的僕人 雅各 ， 我所揀選的 以色列 ， 我提名召你； 你雖不認識我， 我也加給你名號。
ISA|45|5|我是耶和華，再沒有別的了； 除了我以外再沒有上帝。 你雖不認識我， 我必給你束腰。
ISA|45|6|從日出之地到日落之處使人都知道 除我以外，沒有別的。 我是耶和華，再沒有別的了。
ISA|45|7|我造光，又造暗； 施平安，又降災禍； 做成這一切的是我－耶和華。
ISA|45|8|「諸天哪，要如雨傾盆而降， 雲要降下公義， 地要裂開，救恩湧出 ， 使公義也一同滋長； 這都是我－耶和華造的。」
ISA|45|9|「那與造他的主爭論的人有禍了！ 他不過是地上瓦塊中的一片 。 泥土豈可對塑造它的說：『你做的是甚麼？ 你所做的物怎麼沒有把手呢？ 』
ISA|45|10|有人對父親說， 『你生的是甚麼』， 對母親 說， 『你生產的是甚麼』； 這人有禍了！」
ISA|45|11|耶和華－ 以色列 的聖者， 就是造 以色列 的如此說： 「難道我孩子的未來，你們能質問我， 我手的工作，你們可以吩咐我嗎？
ISA|45|12|我造大地，又創造人在地上。 我親手鋪張諸天， 天上萬象也是我所任命的。
ISA|45|13|我憑公義興起 居魯士 ， 又要修直他一切的道路。 他必建造我的城， 釋放我被擄的民， 不為工價，也不為獎賞。」 這是萬軍之耶和華說的。
ISA|45|14|耶和華如此說： 「 埃及 的出產和 古實 的貨物必歸你； 身量高大的 西巴 人，他們必過來歸你，為你所有。 他們必帶著鎖鏈過來跟隨你， 向你下拜，祈求你說： 『上帝真是在你中間，再沒有別的， 沒有別的上帝。』」
ISA|45|15|救主－ 以色列 的上帝啊， 你誠然是隱藏自己的上帝。
ISA|45|16|製造偶像的都要抱愧蒙羞， 他們要一同歸於慚愧。
ISA|45|17|惟有 以色列 必蒙耶和華拯救， 得永遠的救恩。 你們必不蒙羞，也不抱愧， 直到永世無盡。
ISA|45|18|耶和華如此說， 他創造諸天，他是上帝； 他造了地，形成它，堅固它， 並非創造它為荒涼， 而是要給人居住： 「我是耶和華，再沒有別的。
ISA|45|19|我不在隱密黑暗之地說話， 也沒有對 雅各 的後裔說， 『你們尋求我是徒然的』， 我－耶和華所講的是公義， 所說的是正直。」
ISA|45|20|「你們從列國逃脫的人， 要一同聚集前來。 那些抬著雕刻的木偶、 祈求不能救人之神明的， 毫無知識。
ISA|45|21|你們要近前來說明， 讓他們彼此商議。 誰從古時指明這事？ 誰從上古述說它？ 不是我－耶和華嗎？ 除了我以外，再沒有上帝； 我是公義的上帝，又是救主； 除了我以外，再沒有別的了。
ISA|45|22|「地的四極都當轉向我， 就必得救； 因為我是上帝，再沒有別的。
ISA|45|23|我指著自己起誓， 公義從我的口發出，這話並不返回： 『萬膝必向我跪拜， 萬口必憑我起誓。』
ISA|45|24|人論我說 ， 「公義、能力，惟獨在乎耶和華。 人必歸向他， 凡向他發怒的都必蒙羞。
ISA|45|25|以色列 的後裔必因耶和華得稱為義， 並要彼此誇耀。」
ISA|46|1|彼勒 叩拜， 尼波 屈身； 巴比倫 的偶像馱在走獸和牲畜背上。 你們所抬的成了重馱， 使牲畜疲乏。
ISA|46|2|這些神明一同屈身叩拜， 不能救自己 ， 反倒遭人擄去。
ISA|46|3|雅各 家， 以色列 家所有的餘民哪， 你們自從生下就蒙我抱， 自出母胎便由我來背， 你們都要聽從我。
ISA|46|4|直到你們年老，我不改變； 直到你們髮白，我仍扶持。 我已造你，就必背你； 我必抱你，也必拯救。
ISA|46|5|你們將誰與我相比，與我相等， 將誰與我相較，使我們相似呢？
ISA|46|6|他們從錢囊中倒出金子， 用天平秤出銀子， 雇銀匠造成神像， 他們又俯伏，又叩拜。
ISA|46|7|他們抬起神像，扛在肩上， 安置在定處，使它站立， 不離本位； 人呼求它，它卻不回答， 也無法救人脫離災難。
ISA|46|8|你們當記得這事，立定心意 。 叛逆的人哪，要留心思想。
ISA|46|9|要追念上古的事， 因為我是上帝，並無別的； 我是上帝，沒有能與我相比的。
ISA|46|10|我從起初就指明末後的事， 從古時便言明未成的事， 說：「我的籌算必立定； 凡我所喜悅的，我必成就。」
ISA|46|11|我召鷙鳥從東方來， 召那成就我籌算的人從遠方來。 我已說出，就必成就； 我已謀定，也必做成。
ISA|46|12|你們這些心中頑固、 遠離公義的人，要聽從我。
ISA|46|13|我使我的公義臨近，它已不遠。 我的救恩必不遲延。 我要為 以色列 －我的榮耀 在 錫安 施行救恩。
ISA|47|1|少女 巴比倫 哪， 下來坐在塵埃； 迦勒底 啊， 沒有寶座，要坐在地上； 你不再稱為柔弱嬌嫩。
ISA|47|2|要用磨磨麵， 揭去面紗， 脫去長裙， 露腿渡河。
ISA|47|3|你的下體必被露出； 你的羞辱必被看見。 我要報復， 誰也不寬容 。
ISA|47|4|我們的救贖主是 以色列 的聖者， 他的名為萬軍之耶和華。
ISA|47|5|迦勒底 啊， 你要靜坐，進入黑暗中， 因你不再稱為萬國之后。
ISA|47|6|我向我的百姓發怒， 使我的產業受凌辱， 將他們交在你手中； 然而你毫不憐憫他們， 連老年人你也加極重的軛。
ISA|47|7|你說：「我必永遠為后。」 你不將這事放在心上， 也不思想事情的結局。
ISA|47|8|你這專好宴樂、以為地位穩固的， 現在當聽這話。 你心中說： 「惟有我，除我以外再沒有別的。 我必不致寡居， 也不經歷喪子之痛。」
ISA|47|9|哪知，喪子、寡居這兩件事 一日之間忽然臨到你； 你雖多行邪術、廣施魔咒， 這兩件事必全然臨到你身上。
ISA|47|10|你倚靠自己的惡行，說： 「無人看見我。」 你的智慧聰明使你走偏， 你心裏說： 「惟有我，除我以外再沒有別的了。」
ISA|47|11|但災禍臨到你， 你不知如何驅除； 災害落在你身上， 你也無法除掉， 你所不知道的毀滅必忽然臨到你身上。
ISA|47|12|儘管使用從幼年就施行的魔符和眾多的邪術吧！ 或許有些幫助， 或許可以致勝。
ISA|47|13|你籌劃太多，以致疲倦。 讓那些觀天象，看星宿， 在初一說預言的都起來， 救你脫離所要臨到你的事！
ISA|47|14|看哪，他們要像碎秸被火焚燒， 無法救自己脫離火焰的魔掌； 沒有炭火可以取暖 ， 你也不能坐在火旁。
ISA|47|15|你所操勞的事都像這樣； 從你幼年以來與你交易的都各奔己路， 沒有一人來救你。
ISA|48|1|雅各 家，稱為 以色列 名下， 從 猶大 的源頭而出的啊， 你們指著耶和華的名起誓， 提說 以色列 的上帝， 卻不憑誠信，也不憑公義； 你們自稱為聖城之民， 倚靠名為萬軍之耶和華－ 以色列 的上帝； 現在，當聽我言：
ISA|48|2|
ISA|48|3|「先前的事，我自古已說明， 已從我口而出， 是我所指示的； 我瞬間行事，事便成就。
ISA|48|4|因為我知道你是頑梗的； 你的頸項是鐵的， 你的額頭是銅的。
ISA|48|5|所以，我自古就給你說明， 在事未成以先指示你， 免得你說：『這些事是我的偶像所行的， 是我雕刻的偶像和鑄造的神像所命定的。』
ISA|48|6|「你既已聽見，現在要察看這一切； 你們不是要說明嗎？ 從今以後，我要指示你新事， 就是你所不知道的隱密事。
ISA|48|7|這事是現今造的，並非自古就有， 在今日以先，你未曾聽見； 免得你說：『看哪，這事我早已知道了。』
ISA|48|8|誠然你未曾聽見，也未曾知道； 你的耳朵從來未曾開通。 我原知道你行事極其詭詐， 你自從出母胎以來， 就稱為悖逆的。
ISA|48|9|「我為我的名暫且忍怒， 為了我的榮耀向你容忍， 不將你剪除。
ISA|48|10|看哪，我熬煉你，卻不像熬煉銀子； 你在苦難的火爐中，我試煉 你。
ISA|48|11|我為自己的緣故必做這事， 我豈能被褻瀆？ 我必不將我的榮耀歸給別神 。
ISA|48|12|雅各 －我所選召的 以色列 啊， 當聽從我： 我是耶和華， 「我是首先的，也是末後的。
ISA|48|13|我親手立了地的根基， 以右手鋪張諸天； 我一召喚，天地就都立定。
ISA|48|14|你們都當聚集而聽， 偶像 之中誰曾說明這些事？ 耶和華愛他，他必向 巴比倫 成就耶和華的旨意， 耶和華的膀臂也要加在 迦勒底 人身上 。
ISA|48|15|我，惟有我曾說過， 我選召他，領他來， 他的道路必亨通。
ISA|48|16|你們要接近我來聽這話， 我從起初就未曾在隱密之處說話， 萬事之始，我就在那裏。」 現在，主耶和華差遣了我， 帶著他的靈而來 。
ISA|48|17|耶和華－你的救贖主， 以色列 的聖者如此說： 「我是耶和華－你的上帝， 我教導你，使你得益處， 指引你當走的路。
ISA|48|18|甚願你聽從我的命令， 你的平安就會如河水， 你的公義如海浪，
ISA|48|19|你的後裔必多如海沙， 你腹中所生的必多如沙粒。 他的名絕不從我面前剪除， 也不滅絕。」
ISA|48|20|你們要從 巴比倫 出來， 從 迦勒底 人中逃脫， 以歡呼的聲音宣告， 將這事傳揚到地極，說： 耶和華救贖了他的僕人 雅各 ！
ISA|48|21|他引導他們經過沙漠， 他們卻未嘗乾渴； 他為他們使水從磐石流出， 磐石裂開，水就湧出。
ISA|48|22|耶和華說： 「惡人必不得平安！」
ISA|49|1|眾海島啊，當聽從我！ 遠方的眾民哪，要留心聽！ 自出母胎，耶和華就選召我； 自出母腹，他就稱呼我的名。
ISA|49|2|他使我的口如快刀， 把我藏在他手蔭之下； 又使我成為磨利的箭， 把我藏在他箭袋之中；
ISA|49|3|對我說：「你是我的僕人 以色列 ； 我必因你得榮耀。」
ISA|49|4|我卻說：「我勞碌是徒然， 我盡力是虛無虛空。 耶和華誠然以公平待我， 我的賞賜在我的上帝那裏。」
ISA|49|5|現在耶和華說話，他從我出母胎，就造我作他的僕人， 要使 雅各 歸向他， 使 以色列 聚集在他那裏。 耶和華看我為尊貴， 我的上帝是我的力量。
ISA|49|6|他說：「你作我的僕人， 使 雅各 眾支派復興， 使 以色列 中蒙保存的人歸回； 然而此事尚小， 我還要使你作萬邦之光， 使你施行我的救恩，直到地極。」
ISA|49|7|救贖主－ 以色列 的聖者耶和華 對那被人藐視、本國憎惡、 統治者奴役的如此說： 「君王看見就站起來， 領袖也要下拜； 這都是因信實的耶和華， 因揀選你的 以色列 的聖者。」
ISA|49|8|耶和華如此說： 「在悅納的時候，我應允了你； 在拯救的日子，我幫助了你。 我要保護你， 要藉著你與百姓立約， 為了復興遍地， 使人承受荒蕪之地為業；
ISA|49|9|對那被捆綁的人說：『出來吧！』 對在黑暗裏的人說：『顯現吧！』 他們在路上必得飲食， 在光禿的高地必有食物。
ISA|49|10|他們不飢不渴， 炎熱和烈日必不傷害他們； 因為憐憫他們的必引導他們， 領他們到水泉旁邊。
ISA|49|11|我必在眾山開闢路徑， 大道也要填高。
ISA|49|12|看哪，他們從遠方來； 有些從北方來，有些從西方來， 有些從 色弗尼 地來。」
ISA|49|13|諸天哪，應當歡呼！ 大地啊，應當快樂！ 眾山哪，應當揚聲歌唱！ 因為耶和華已經安慰他的百姓， 他要憐憫他的困苦之民。
ISA|49|14|錫安 說：「耶和華離棄了我， 主忘記了我。」
ISA|49|15|婦人焉能忘記她吃奶的嬰孩， 不憐憫她所生的兒子？ 即或有忘記的， 我卻不忘記你。
ISA|49|16|看哪，我將你銘刻在我掌上， 你的城牆常在我眼前。
ISA|49|17|建立你的勝過毀壞你的， 使你荒廢的必都離你而去。
ISA|49|18|你舉目向四圍觀看， 他們都聚集來到你這裏。 我指著我的永生起誓， 你定要以他們為妝飾佩戴， 帶著他們，像新娘一樣。 這是耶和華說的。
ISA|49|19|至於你荒廢淒涼之處， 並你被毀壞之地， 如今居民必嫌太窄， 吞滅你的必離你遙遠。
ISA|49|20|你要再聽見喪失子女後所生的兒女說： 「這地方我居住太窄， 請你給我地方居住。」
ISA|49|21|那時你心裏必說：「我既喪子不育， 被擄，飄流在外 ， 誰給我生了這些？ 誰將他們養大呢？ 看哪，我被撇下獨自一人時， 他們都在哪裏呢？」
ISA|49|22|主耶和華如此說： 「看哪，我必向列國舉手， 向萬民豎立大旗； 他們必將你的兒子抱在懷中帶來， 將你的女兒背在肩上扛來。
ISA|49|23|列王必作你的養父， 王后必作你的乳母。 他們必以臉伏地，向你下拜， 並舔你腳上的塵土。 你就知道我是耶和華， 等候我的必不致羞愧。」
ISA|49|24|勇士搶去的豈能奪回？ 被殘暴者擄掠的豈能得解救呢？
ISA|49|25|但耶和華如此說： 「就是勇士所擄掠的，也可以奪回； 殘暴者所搶的，也可以得解救。 與你相爭的，我必與他相爭， 我也要拯救你的兒女。
ISA|49|26|我必使那欺壓你的吃自己的肉， 飲自己的血，如喝甜酒喝醉一樣。 凡有血肉之軀的都必知道我－耶和華是你的救主， 是你的救贖主，是 雅各 的大能者。」
ISA|50|1|耶和華如此說： 「我休了你們的母親， 她的休書在哪裏呢？ 我將你們賣給了我哪一個債主呢？ 看哪，你們被賣是因你們的罪孽； 你們的母親被休，是因你們的過犯。
ISA|50|2|我來的時候，為何沒有人呢？ 我呼喚的時候，為何無人回應呢？ 我的膀臂豈是過短、不能救贖嗎？ 我豈無拯救之力嗎？ 看哪，我一斥責，海就乾了； 我使江河變為曠野， 其中的魚因無水腥臭，乾渴而死。
ISA|50|3|我使諸天以黑暗為衣， 以麻布為遮蓋。」
ISA|50|4|主耶和華賜我受教者的舌頭， 使我知道怎樣用言語扶助疲乏的人。 主每天早晨喚醒，喚醒我的耳朵， 使我能聽，像受教者一樣。
ISA|50|5|主耶和華開啟我的耳朵， 我並未違背，也未退後。
ISA|50|6|人打我的背，我任他打； 人拔我兩頰的鬍鬚，我由他拔； 人侮辱我，向我吐唾沫，我並不掩面。
ISA|50|7|主耶和華必幫助我， 所以我不抱愧。 我硬著臉面好像堅石， 也知道我必不致蒙羞。
ISA|50|8|稱我為義的與我相近； 誰與我爭論， 讓我們來對質； 誰與我作對， 讓他近前來吧！
ISA|50|9|看哪，主耶和華必幫助我， 誰能定我有罪呢？ 看哪，他們都要像衣服漸漸破舊， 被蛀蟲蛀光。
ISA|50|10|你們當中有誰是敬畏耶和華， 聽從他僕人的話語， 卻行在黑暗中，沒有亮光的， 當倚靠耶和華的名， 仰賴自己的上帝。
ISA|50|11|看哪，你們當中所有點火、以火把圍繞自己的人， 當行走在你們的火焰 裏， 並你們所點的火把中。 這是我親手為你們定的： 你們必躺臥在悲慘之中。
ISA|51|1|追求公義、 尋求耶和華的人哪， 當聽從我！ 你們要追想自己是從哪塊磐石鑿出， 從哪個巖穴挖掘而來；
ISA|51|2|要追想你們的祖宗 亞伯拉罕 和生你們的 撒拉 ； 因為我選召 亞伯拉罕 時，他只有一個人， 但我賜福給他， 使他增多。
ISA|51|3|耶和華已經安慰 錫安 ， 安慰了 錫安 一切的廢墟， 使曠野如 伊甸 ， 使沙漠像耶和華的園子； 其中必有歡喜、快樂、感謝， 和歌唱的聲音。
ISA|51|4|我的民哪，要留心聽我， 我的國啊，要向我側耳； 因為訓誨必從我而出， 我必使我的公理成為萬民之光。
ISA|51|5|我的公義臨近， 我的救恩發出。 我的膀臂要審判萬民， 眾海島都要等候我，倚賴我的膀臂。
ISA|51|6|你們要向天舉目， 觀看下面的地； 天必像煙雲消散， 地必如衣服漸漸破舊； 其上的居民也要如此 死亡。 惟有我的救恩永遠長存， 我的公義也不廢掉。
ISA|51|7|知道公義、將我的訓誨存在心中的人哪， 當聽從我！ 不要怕人的辱罵， 也不要因人的毀謗驚惶。
ISA|51|8|因為他們必像衣服被蛀蟲蛀； 像羊毛被蟲子咬。 惟有我的公義永遠長存， 我的救恩直到萬代。
ISA|51|9|耶和華的膀臂啊，興起，興起！ 以能力為衣穿上， 像古時的年日，像上古的世代一樣興起！ 從前砍碎 拉哈伯 、 刺透大魚的，不是你嗎？
ISA|51|10|使海與深淵的水乾涸， 在海的深處開路， 使救贖的民走過的，不是你嗎？
ISA|51|11|耶和華救贖的民必歸回， 歌唱來到 錫安 ； 永恆的喜樂必歸到他們頭上。 他們必得著歡喜快樂， 憂傷嘆息盡都逃避。
ISA|51|12|我，惟有我是安慰你們的。 你是誰，竟怕那必死的人， 怕那生命如草的世人，
ISA|51|13|卻忘記鋪張諸天、立定地基、 造你的耶和華？ 你因欺壓者圖謀毀滅所發的暴怒， 終日害怕， 其實那欺壓者的暴怒在哪裏呢？
ISA|51|14|被擄的即將得釋放， 不至於死而下入地府， 也不致缺乏食物。
ISA|51|15|我是耶和華－你的上帝， 我攪動大海，使海中的波浪澎湃， 萬軍之耶和華是我的名。
ISA|51|16|我已將我的話放在你口中， 用我的手影遮蔽你， 為要安定諸天，立定地基， 並對 錫安 說：「你是我的百姓。」
ISA|51|17|耶路撒冷 啊，興起，興起！ 站起來！ 你從耶和華手中喝了他憤怒的杯， 那使人東倒西歪的杯，直到喝盡。
ISA|51|18|她所生育的孩子中，沒有一個攙她的； 她所撫養的孩子中，沒有一個扶她的。
ISA|51|19|這雙重的災難臨到你， 有誰憐憫你呢？ 破壞和毀滅，饑荒和戰爭臨到， 我如何能安慰你呢 ？
ISA|51|20|你的孩子發昏， 在各街頭躺臥， 如同網羅裏的羚羊， 滿了耶和華的憤怒， 滿了你上帝的斥責。
ISA|51|21|因此，你這困苦卻非因酒而醉的， 當聽這話，
ISA|51|22|你的主，耶和華， 就是為他百姓辯護的上帝如此說： 「看哪，我已從你手中接過 那使人東倒西歪的杯， 就是我憤怒的杯， 你必不再喝。
ISA|51|23|我必將這杯遞在苦待你的人 手中。 他們曾對你說：『你屈身， 任我們踐踏過去吧！』 你就以背為地， 又如街道，任人走過。
ISA|52|1|錫安 哪，興起！興起！ 穿上你的能力！ 聖城 耶路撒冷 啊，穿上你華美的衣服！ 因為從今以後， 未受割禮、不潔淨的必不再進入你中間。
ISA|52|2|耶路撒冷 啊，抖去塵埃， 起來坐在王位上！ 被擄的 錫安 哪， 解開你頸上的鎖鏈！
ISA|52|3|耶和華如此說：「你們白白地被賣，也必不用銀子贖回。」
ISA|52|4|主耶和華如此說：「先前我的百姓下到 埃及 ，在那裏寄居，末後又有 亞述 人欺壓他們。」
ISA|52|5|我的百姓既是白白地被擄，如今我在這裏做甚麼呢？這是耶和華說的。轄制他們的人歡呼 ，我的名終日不斷受褻瀆，這是耶和華說的。
ISA|52|6|因此，我的百姓必認識我的名；在那日，他們必知道說這話的就是我。看哪，是我！」
ISA|52|7|在山上報佳音，傳平安， 報好信息，傳揚救恩， 那人的腳蹤何等佳美啊！ 他對 錫安 說：「你的上帝作王了！」
ISA|52|8|聽啊，你守望之人的聲音， 他們揚聲一同歡唱； 因為他們必親眼看見耶和華返回 錫安 。
ISA|52|9|耶路撒冷 的廢墟啊， 要出聲一同歡唱； 因為耶和華安慰了他的百姓， 救贖了 耶路撒冷 。
ISA|52|10|耶和華在萬國眼前露出聖臂， 地的四極都要看見我們上帝的救恩。
ISA|52|11|離開吧！離開吧！ 你們要從 巴比倫 出來。 你們扛抬耶和華器皿的人哪， 不要沾不潔淨的東西， 離去時務要保持潔淨。
ISA|52|12|你們出來必不致匆忙， 也不致奔逃； 因為耶和華要在你們前頭行， 以色列 的上帝必作你們的後盾。
ISA|52|13|看哪，我的僕人行事必有智慧， 他必被高升，高舉， 升到至高之處。
ISA|52|14|許多人因他 驚奇 ─他的面貌比別人憔悴， 他的外表比世人枯槁─
ISA|52|15|同樣，他也必使許多國家驚奇 ， 君王要向他閉口。 未曾傳給他們的，他們必看見； 未曾聽見過的事，他們要明白。
ISA|53|1|我們所傳的有誰信呢？ 耶和華的膀臂向誰顯露呢？
ISA|53|2|他在耶和華面前生長如嫩芽， 像根出於乾地。 他無佳形美容使我們注視他， 也無美貌使我們仰慕他。
ISA|53|3|他被藐視，被人厭棄； 多受痛苦，常經憂患。 他被藐視， 好像被人掩面不看的一樣， 我們也不尊重他。
ISA|53|4|他誠然擔當我們的憂患， 背負我們的痛苦； 我們卻以為他受責罰， 是被上帝擊打苦待。
ISA|53|5|他為我們的過犯受害， 為我們的罪孽被壓傷。 因他受的懲罰，我們得平安； 因他受的鞭傷，我們得醫治。
ISA|53|6|我們都如羊走迷， 各人偏行己路； 耶和華使我們眾人的罪孽都歸在他身上。
ISA|53|7|他被欺壓受苦， 卻不開口； 他像羔羊被牽去宰殺， 又像羊在剪毛的人手下無聲， 他也是這樣不開口。
ISA|53|8|因受欺壓和審判，他被奪去， 誰能想到他的世代呢？ 因為他從活人之地被剪除， 為我百姓 的罪過他被帶到死裏 。
ISA|53|9|他雖然未行殘暴， 口中也沒有詭詐， 人還使他與惡人同穴， 與財主同墓 。
ISA|53|10|耶和華的旨意要壓傷他， 使他受苦。 當他的生命作為贖罪祭時 ， 他必看見後裔，他的年日必然長久。 耶和華所喜悅的事，必在他手中亨通。
ISA|53|11|因自己的勞苦，他必看見光 就心滿意足。 因自己的認識，我的義僕使許多人得稱為義， 他要擔當他們的罪孽。
ISA|53|12|因此，我要使他與位大的同份， 與強盛的均分擄物。 因為他傾倒自己的生命，以致於死， 也列在罪犯之中。 他卻擔當多人的罪， 為他們的過犯代求 。
ISA|54|1|你這不懷孕、不生育的，要歡呼； 你這未曾經過產難的，要歡呼，揚聲呼喊； 因為被遺棄的婦人， 比有丈夫的人兒女更多； 這是耶和華說的。
ISA|54|2|要擴張你帳幕之地， 伸展你居所的幔子，不要縮回； 要放長你的繩子， 堅固你的橛子。
ISA|54|3|因為你要向左向右開展， 你的後裔必得列國為業， 又使荒廢的城鎮有人居住。
ISA|54|4|不要懼怕，因你必不致蒙羞； 不要抱愧，因你必不致受辱。 你必忘記年輕時的羞愧， 不再記得守寡的恥辱。
ISA|54|5|因為造你的是你的丈夫， 萬軍之耶和華是他的名； 救贖你的是 以色列 的聖者， 他必稱為全地之上帝。
ISA|54|6|耶和華召你， 如同召回心中憂傷遭遺棄的婦人， 就是年輕時所娶被遺棄的妻子； 這是你的上帝說的。
ISA|54|7|我離棄你不過片時， 卻要大施憐憫將你尋回。
ISA|54|8|我因漲溢的怒氣， 一時向你轉臉， 但我要以永遠的慈愛憐憫你； 這是耶和華－你的救贖主說的。
ISA|54|9|這事於我有如 挪亞 的洪水； 我怎樣起誓不再使 挪亞 的洪水淹沒全地， 也照樣起誓不再向你發怒， 且不斥責你。
ISA|54|10|大山可以挪開， 小山可以遷移， 但我的慈愛必不離開你， 我平安的約也不遷移； 這是憐憫你的耶和華說的。
ISA|54|11|你這受困苦、被暴風捲走、不得憐憫的城， 看哪，我必以灰泥來做你的石頭， 以藍寶石立你的根基，
ISA|54|12|又以紅寶石造你的女牆， 以晶瑩的珠玉造你的城門， 以珍貴的寶石造你四圍的邊界。
ISA|54|13|你的兒女都要領受耶和華的教導， 你的兒女必大享平安。
ISA|54|14|你必因公義得堅立， 必遠離欺壓，毫不懼怕； 你必遠離驚嚇，驚嚇必不臨近你。
ISA|54|15|若有人攻擊你，這非出於我； 凡攻擊你的，必因你仆倒。
ISA|54|16|看哪，我造了那吹炭火、打造合用兵器的鐵匠； 我也造了那殘害人、行毀滅的人。
ISA|54|17|凡為攻擊你而造的兵器必無效用； 在審判時興起用口舌攻擊你的， 你必駁倒他。 這是耶和華僕人的產業， 是他們從我所得的義； 這是耶和華說的。
ISA|55|1|來！你們所有乾渴的，都當來到水邊； 沒有銀錢的也可以來。 你們都來，買了吃； 不用銀錢，不付代價， 就可買酒和奶。
ISA|55|2|你們為何花錢買那不是食物的東西， 用勞碌得來的買那無法使人飽足的呢？ 你們要留意聽從我的話，就能吃那美物， 得享肥甘，心中喜樂。
ISA|55|3|當側耳而聽，來到我這裏； 要聽，就必存活。 我要與你們立永約， 就是應許給 大衛 那可靠的慈愛。
ISA|55|4|看哪，我已立他作萬民的見證， 立他作萬民的君王和發令者。
ISA|55|5|看哪，你要召集素不認識的國民， 素不認識的國民要奔向你； 這都因耶和華─你的上帝， 因 以色列 的聖者已經榮耀了你。
ISA|55|6|當趁耶和華可尋找的時候尋找他， 在他接近的時候求告他。
ISA|55|7|惡人當離棄自己的道路， 不義的人應除掉自己的意念。 歸向耶和華，耶和華就必憐憫他； 當歸向我們的上帝，因為他必廣行赦免。
ISA|55|8|我的意念非同你們的意念， 我的道路非同你們的道路。 這是耶和華說的。
ISA|55|9|天怎樣高過地， 照樣，我的道路高過你們的道路， 我的意念高過你們的意念。
ISA|55|10|雨雪從天而降，並不返回， 卻要滋潤土地，使地面發芽結實， 使撒種的有種，使要吃的有糧。
ISA|55|11|我口所出的話也必如此， 絕不徒然返回， 卻要成就我的旨意， 達成我差它的目的。
ISA|55|12|你們必歡歡喜喜出來， 平平安安蒙引導。 大山小山必在你們面前歡呼， 田野的樹木也都拍掌。
ISA|55|13|松樹長出，代替荊棘； 番石榴長出，代替蒺藜。 這要為耶和華留名， 作為永不磨滅的證據。
ISA|56|1|耶和華如此說： 「你們當守公平，行公義； 因我的救恩臨近， 我的公義將要顯現。
ISA|56|2|謹守安息日不予干犯， 禁止己手不作惡， 如此行、如此持守的人有福了！」
ISA|56|3|與耶和華聯合的外邦人不要說： 「耶和華將我和他的子民分別出來。」 太監也不要說：「看哪，我是枯樹。」
ISA|56|4|因為耶和華如此說： 「那些謹守我的安息日， 選擇我旨意， 持守我約的太監，
ISA|56|5|我必使他們在我殿中，在我牆內， 有紀念碑，有名號， 勝過有兒有女； 我必賜他們永遠的名，不能剪除。
ISA|56|6|「那些與耶和華聯合， 事奉他，愛他名， 作他僕人的外邦人， 凡謹守安息日不予干犯， 又持守我約的人，
ISA|56|7|我必領他們到我的聖山， 使他們在我的禱告的殿中喜樂。 他們的燔祭和祭物， 在我壇上必蒙悅納， 因我的殿必稱為萬民禱告的殿。
ISA|56|8|我還要召集更多的人 歸併到這些被召集的人中。 這是召集被趕散的 以色列 人的 主耶和華說的。」
ISA|56|9|野地的走獸，你們都來吞吃吧！ 林中的野獸，你們也來吞吃！
ISA|56|10|以色列 的守望者都瞎了眼， 沒有知識； 都是啞狗，不會吠叫， 只知做夢，躺臥，貪睡，
ISA|56|11|這些狗貪食，不知飽足。 這些牧人不知明辨， 他們都偏行己路， 人人追求自己的利益。
ISA|56|12|他們說：「來吧！我去拿酒， 讓我們暢飲烈酒吧！ 明天必和今天一樣， 甚至更好！」
ISA|57|1|義人死亡， 無人放在心上； 虔誠的人被接去， 無人理解； 義人被接去，以免禍患。
ISA|57|2|行為正直的人進入平安， 得以在床上安歇 。
ISA|57|3|到這裏來吧！ 你們這些巫婆的兒子， 姦夫和妓女的後代；
ISA|57|4|你們向誰戲笑？ 向誰張口吐舌呢？ 你們豈不是叛逆所生的兒女， 虛謊所生的後代嗎？
ISA|57|5|你們在橡樹 中間，在各青翠的樹下慾火攻心； 在山谷間，在巖隙下殺了兒女；
ISA|57|6|去拜谷中光滑的石頭有你們的份， 這些就是你們的命運。 你向它們獻澆酒祭，獻供物， 這事我豈能容忍嗎？
ISA|57|7|你在高而又高的山上安設床舖， 上那裏去獻祭。
ISA|57|8|你在門後，在門框後， 立起你的牌來； 你離棄了我，赤露己身， 又爬上自己所鋪寬闊的床鋪， 與它們立約； 你喜愛它們的床，看著它們的赤體 。
ISA|57|9|你帶了油到 摩洛 那裏， 加上許多香水。 你派遣使者往遠方去， 甚至降到陰間，
ISA|57|10|因路途遙遠，你就疲倦， 卻不說，這是枉然， 以為能找到復興之力， 所以不覺疲憊。
ISA|57|11|你怕誰，因誰恐懼， 竟說謊，不記得我， 不將這事放在心上。 是否因我許久閉口不言， 你就不怕我了呢？
ISA|57|12|我可以宣告你的公義和你的作為， 但它們與你無益。
ISA|57|13|你哀求的時候， 讓你所搜集的神像 拯救你吧！ 風要把它們全都颳散， 吹一口氣就都吹走。 但那投靠我的必得地產， 承受我的聖山為業。
ISA|57|14|耶和華說： 「你們要修築，修築，要預備道路， 除掉我百姓路中的絆腳石。」
ISA|57|15|那至高無上、永遠長存、 名為聖者的如此說： 「我住在至高至聖的所在， 卻與心靈痛悔的謙卑人同住； 要使謙卑的人心靈甦醒， 使痛悔的人內心復甦。
ISA|57|16|我必不長久控訴，也不永遠懷怒， 因為我雖使靈性發昏，我也造了人的氣息。
ISA|57|17|我因人貪婪的罪孽，發怒擊打他； 我轉臉向他發怒， 他卻仍隨意背道而行。
ISA|57|18|我看見他的行為， 要醫治他，引導他 ， 使他和與他一同哀傷的人都得安慰。
ISA|57|19|我要醫治他， 他要結出嘴唇的果實。 平安，平安，歸給遠處和近處的人！ 這是耶和華說的。」
ISA|57|20|但是惡人好像翻騰的海， 不得平靜； 其中的水常湧出污穢和淤泥。
ISA|57|21|我的上帝說：「惡人必不得平安！」
ISA|58|1|你要大聲喊叫，不要停止； 要揚聲，好像吹角； 向我的百姓宣告他們的過犯， 向 雅各 家陳述他們的罪惡。
ISA|58|2|他們天天尋求我， 樂意明白我的道， 好像行義的國家， 未離棄它的上帝的典章； 他們向我求問公義的判詞， 喜悅親近上帝。
ISA|58|3|「我們禁食，你為何不看呢？ 我們刻苦己心，你為何不理會呢？」 看哪，你們禁食的時候仍追求私利， 剝削為你們做苦工的人。
ISA|58|4|看哪，你們禁食，卻起紛爭興訟， 以兇惡的拳頭打人。 你們今日這種禁食 無法使你們的聲音聽聞於高處。
ISA|58|5|這豈是我所要的禁食， 為人所用以刻苦己心的日子嗎？ 我難道只是叫人如蘆葦般低頭， 鋪上麻布和灰燼嗎？ 你能稱此為禁食， 為耶和華所悅納的日子嗎？
ISA|58|6|我所要的禁食，豈不是要你鬆開兇惡的繩， 解開軛上的索， 使被欺壓的得自由， 折斷一切的軛嗎？
ISA|58|7|豈不是要你把食物分給飢餓的人， 將流浪的窮人接到家中， 見赤身的給他衣服遮體， 而不隱藏自己避開你的骨肉嗎？
ISA|58|8|這樣，必有光如晨光破曉照耀你， 你也要快快得到醫治； 你的公義在你前面行， 耶和華的榮光必作你的後盾。
ISA|58|9|那時你求告，耶和華必應允； 你呼求，他必說：「我在這裏。」 你若從你中間除掉重軛 和指摘人的指頭，並發惡言的事，
ISA|58|10|向飢餓的人施憐憫， 使困苦的人得滿足； 你在黑暗中就必得著光明， 你的幽暗必變如正午。
ISA|58|11|耶和華必時常引導你， 在乾旱之地使你心滿意足， 又使你骨頭強壯。 你必如有水澆灌的園子， 又像水流不絕的泉源。
ISA|58|12|你們中間必有人起來修造久已荒廢之處， 立起代代相承的根基。 你必稱為修補裂痕的， 和重修路徑給人居住的。
ISA|58|13|你若禁止自己的腳踐踏安息日， 不在我的聖日做自己高興的事， 稱安息日為「可喜樂的」， 稱耶和華的聖日為「可尊重的」， 尊敬這日， 不走自己的道路， 不求自己的喜悅， 也不隨意說話；
ISA|58|14|那麼，你就會以耶和華為樂。 耶和華要使你乘駕於地的高處， 又要以你祖先 雅各 的產業養育你； 這是耶和華親口說的。
ISA|59|1|看哪，耶和華的膀臂並非過短，不能拯救， 耳朵並非發沉，不能聽見，
ISA|59|2|但你們的罪孽使你們與上帝隔絕， 你們的罪惡使他轉臉不聽你們。
ISA|59|3|因你們的手掌被血沾染， 你們的指頭被罪玷污， 你們的嘴唇說謊言， 你們的舌頭出惡語。
ISA|59|4|無人按公義控訴， 也無人憑誠實辯白； 卻倚靠虛妄，口說謊言， 懷毒害，生罪孽。
ISA|59|5|他們孵毒蛇蛋， 結蜘蛛網。 凡吃這蛋的必死， 蛋一打破，就孵出蛇來。
ISA|59|6|所結的網不能當衣服， 無法掩蓋自己所作所為。 他們的行為全是邪惡， 手所做的盡都殘暴。
ISA|59|7|他們的腳奔跑行惡， 急速流無辜者的血； 他們的思想全是惡念， 走過的路盡是破壞與毀滅。
ISA|59|8|平安的路，他們不知道， 所行的事無一公平。 他們為自己修築彎曲的路， 凡走這路的都不得平安。
ISA|59|9|因此，公平離我們甚遠， 公義追不上我們。 我們指望光亮，看哪，卻只有黑暗， 指望光明，卻行在幽暗中。
ISA|59|10|我們用手摸牆，好像盲人， 四處摸索，如同失明的人； 中午時我們絆倒，如在黃昏一樣， 在強壯的人中，我們好像死人一般。
ISA|59|11|我們全都咆哮如熊， 哀鳴如鴿子； 指望公平，卻得不著； 指望救恩，它卻遠離。
ISA|59|12|我們的過犯在你面前增加， 罪惡作證控告我們； 過犯與我們同在。 至於我們的罪孽，我們都知道：
ISA|59|13|就是悖逆，否認耶和華， 轉去不跟從我們的上帝， 口說欺壓和叛逆的話， 心懷謊言，隨即說出；
ISA|59|14|公平轉而退後， 公義站在遠處， 誠實仆倒在廣場上， 正直不得進入；
ISA|59|15|誠實少見， 離棄邪惡的人反成掠物。 那時，耶和華見沒有公平， 就不喜悅。
ISA|59|16|他見無人， 竟無一人代求，甚為詫異， 就用自己的膀臂拯救他， 以公義扶持他。
ISA|59|17|他穿上公義為鎧甲， 戴上救恩為頭盔， 穿上報復為衣服， 披戴熱心為外袍。
ISA|59|18|他必按人的行為報應， 惱怒他的敵人， 報復他的仇敵， 向眾海島施行報應。
ISA|59|19|在日落之處，人必敬畏耶和華的名； 在日出之地，人必敬畏他的榮耀。 他必如湍急的河流沖來， 耶和華的靈催逼他自己。
ISA|59|20|必有一位救贖主來到 錫安 ， 來到 雅各 族中離棄過犯的人那裏； 這是耶和華說的。
ISA|59|21|耶和華說：「這就是我與他們所立的約：我加給你的靈，傳給你的話，必不離你的口，也不離你後裔與你後裔之後裔的口，從今直到永遠；這是耶和華說的。」
ISA|60|1|興起，發光！因為你的光已來到！ 耶和華的榮光發出照耀著你。
ISA|60|2|看哪，黑暗籠罩大地， 幽暗遮蓋萬民， 耶和華卻要升起照耀你， 他的榮光要顯在你身上。
ISA|60|3|列國要來就你的光， 列王要來就你發出的光輝。
ISA|60|4|你舉目向四圍觀看， 眾人都聚集到你這裏。 你的兒子從遠方來， 你的女兒也被抱著帶來。
ISA|60|5|那時，你看見就有光榮， 你的心興奮歡暢 ； 因為大海那邊的財富必歸你， 列國的財寶也來歸你。
ISA|60|6|成群的駱駝， 並 米甸 和 以法 的獨峰駝遮滿你； 示巴 的眾人都必來到， 要奉上黃金和乳香， 又要傳揚讚美耶和華的話。
ISA|60|7|基達 的羊群都聚集到你這裏， 尼拜約 的公羊供你使用， 獻在我壇上蒙悅納； 我必榮耀我那榮耀的殿。
ISA|60|8|那些飛來如雲、 又像鴿子飛向窗戶的是誰呢？
ISA|60|9|眾海島必等候我 ， 他施 的船隻領先， 將你的兒女，連同他們的金銀從遠方帶來， 這都因 以色列 的聖者、耶和華－你上帝的名， 因為他已經榮耀了你。
ISA|60|10|外邦人要建造你的城牆， 他們的君王必服事你。 我曾發怒擊打你， 如今卻施恩憐憫你。
ISA|60|11|你的城門必時常開放， 晝夜不關， 使人將列國的財物帶來歸你， 他們的君王也被牽引而來。
ISA|60|12|不事奉你的那邦、那國要滅亡， 那些國家必全然荒廢。
ISA|60|13|黎巴嫩 的榮耀， 就是松樹、杉樹、黃楊樹， 都必一同歸你， 用以裝飾我聖所坐落之處； 我也要使我腳所踏之地得榮耀。
ISA|60|14|壓制你的，他的子孫必來向你屈身； 藐視你的，都要在你腳前下拜。 人要稱你為「耶和華的城」， 為「 以色列 聖者的 錫安 」。
ISA|60|15|你雖曾被拋棄，被恨惡， 甚至無人經過， 我卻使你有永遠的榮華， 成為世世代代的喜樂。
ISA|60|16|你要吃列國的奶， 吃列王的乳。 你就知道我－耶和華是你的救主， 是你的救贖主，是 雅各 的大能者。
ISA|60|17|我要賞賜金子代替銅， 賞賜銀子代替鐵， 銅代替木頭， 鐵代替石頭。 我要以和平為你的官長， 以公義為你的監督。
ISA|60|18|你的地不再聽聞殘暴的事， 境內不再聽見破壞與毀滅。 你必稱你的牆為「拯救」， 稱你的門為「讚美」。
ISA|60|19|白晝太陽不再作你的光， 月亮 也不再發光照耀你； 耶和華卻要作你永遠的光， 你的上帝要成為你的榮耀。
ISA|60|20|你的太陽不再落下， 月亮也不消失； 因為耶和華必作你永遠的光。 你悲哀的日子定要結束。
ISA|60|21|你的居民全是義人， 永遠得地為業； 他們是我栽的苗，是我手的工作， 為了彰顯我的榮耀。
ISA|60|22|稀少的要成為大族， 弱小的要變為強國。 我－耶和華到了時候必速速成就這事。
ISA|61|1|主耶和華的靈在我身上， 因為耶和華用膏膏我， 叫我報好信息給貧窮的人， 差遣我醫好傷心的人， 報告被擄的得釋放， 被捆綁的得自由；
ISA|61|2|宣告耶和華的恩年 和我們的上帝報仇的日子； 安慰所有悲哀的人，
ISA|61|3|為 錫安 悲哀的人，賜華冠代替灰燼， 喜樂的油代替悲哀， 讚美為衣代替憂傷的靈； 稱他們為「公義樹」， 是耶和華所栽植的，為要彰顯他的榮耀。
ISA|61|4|他們必修造久已荒涼的廢墟， 建立先前淒涼之處， 重修歷代荒涼之城。
ISA|61|5|那時，陌生人要伺候、牧放你們的羊群； 外邦人必為你們耕種田地， 修整你們的葡萄園。
ISA|61|6|但你們要稱為「耶和華的祭司」， 稱作「我們上帝的僕人」。 你們必享用列國的財物， 必承受他們的財富 。
ISA|61|7|因為他們所受雙倍的羞辱， 凌辱被稱為他們的命運， 因此，他們在境內必得雙倍的產業， 永遠之樂必歸給他們。
ISA|61|8|因為我－耶和華喜愛公平， 恨惡搶奪與惡行 ； 我要憑誠實施行報償， 與我的百姓立永約。
ISA|61|9|他們的後裔必在列國中為人所知， 他們的子孫在萬民中為人所識； 凡看見他們的必承認他們是耶和華所賜福的後裔。
ISA|61|10|我因耶和華大大歡喜， 我的心因上帝喜樂； 因他以拯救為衣給我穿上， 以公義為外袍給我披上， 好像新郎戴上華冠， 又如新娘佩戴首飾。
ISA|61|11|地怎樣使芽長出， 園子怎樣使所栽種的生長， 主耶和華也必照樣 使公義和讚美在萬國中發出。
ISA|62|1|我因 錫安 必不靜默， 為 耶路撒冷 必不安寧， 直到它的公義如光輝發出， 它的救恩如火把燃燒。
ISA|62|2|列國要看見你的公義， 列王要看見你的榮耀。 你必得新的名字， 是耶和華親口起的。
ISA|62|3|你在耶和華的手中成為華冠， 在你上帝的掌上成為冠冕。
ISA|62|4|你不再稱為「被撇棄的」， 你的地也不再稱為「荒蕪的」； 你要稱為「我所喜悅的」， 你的地要稱為「有歸屬的」。 因為耶和華喜悅你， 你的地必歸屬於他。
ISA|62|5|年輕人怎樣娶童女， 你的百姓也要照樣娶你； 新郎怎樣因新娘而喜樂， 你的上帝也要如此以你為樂。
ISA|62|6|耶路撒冷 啊， 我在你城牆上設立守望者， 他們晝夜不停地呼喊。 呼求耶和華的啊，你們不要歇息，
ISA|62|7|也不要使他歇息， 直等他建立 耶路撒冷 ， 使 耶路撒冷 在地上為人所讚美。
ISA|62|8|耶和華指著自己的右手和大能的膀臂起誓說： 「我必不再將你的五穀給仇敵作食物， 外邦人也必不再喝你勞碌得來的新酒。
ISA|62|9|惟有那收割的要吃，並讚美耶和華； 那儲藏葡萄的要在我聖所院內喝。」
ISA|62|10|你們當從門經過，經過， 預備百姓的路。 你們要修築，修築大道， 清除石頭， 為萬民豎立大旗。
ISA|62|11|看哪，耶和華曾宣告到地極， 你們要對 錫安 說： 「看哪，你的拯救者已來到。 看哪，他的賞賜在他那裏， 他的報償在他面前。」
ISA|62|12|人稱他們為「聖民」，為「耶和華救贖的民」， 你也必稱為「受眷顧的」，為「不被撇棄的城」。
ISA|63|1|這從 以東 的 波斯拉 來， 穿紅衣服， 裝扮華美， 能力廣大， 大步向前邁進的是誰呢？ 就是我， 憑公義說話， 以大能施行拯救的。
ISA|63|2|你為何以紅色裝扮？ 你的衣服為何像踹醡酒池的人呢？
ISA|63|3|我獨自踹醡酒池， 萬民中並無一人與我同在。 我發怒，將他們踹下， 發烈怒將他們踐踏。 他們的血濺在我的衣服上， 玷污了我一切的衣裳。
ISA|63|4|因為報仇之日在我心中， 救贖我民之年已經來到。
ISA|63|5|我仰望，見無人幫助； 我詫異，竟無人扶持。 因此，我的膀臂為我施行拯救； 我的烈怒將我扶持。
ISA|63|6|我發怒，踹下眾民； 發烈怒，使他們喝醉， 又將他們的血倒在地上。
ISA|63|7|我要照耶和華一切所賜給我們的， 並他憑憐憫與豐盛的慈愛 所賜給 以色列 家的大恩， 述說他的慈愛和美德。
ISA|63|8|他說：「他們誠然是我的百姓， 未行虛假的子民。」 這樣，他就作了他們的救主。
ISA|63|9|他們在一切苦難當中， 他也同受苦難， 並且他面前的使者拯救他們 。 他以慈愛和憐憫救贖他們， 在古時的日子時常抱他們，背他們。
ISA|63|10|他們竟然悖逆，使他的聖靈憂傷。 他就轉變，成為他們的仇敵， 親自攻擊他們。
ISA|63|11|那時，他的百姓想起古時 摩西 的日子： 「那將百姓和牧養群羊的人 從海裏領上來的在哪裏呢？ 那將聖靈降在他們中間，
ISA|63|12|以榮耀的膀臂在 摩西 右邊行動， 在百姓面前將水分開， 為要建立自己永遠的名，
ISA|63|13|又帶領他們經過深處的在哪裏呢？」 他們如馬行走曠野，不致絆跌；
ISA|63|14|又如牲畜下到山谷， 耶和華的靈使他們得安息； 照樣，你也引導你的百姓， 為要建立自己榮耀的名。
ISA|63|15|求你從天上， 從你神聖榮耀的居所垂顧觀看。 你的熱心和你大能的作為在哪裏呢？ 你內心的關懷和你的憐憫向我們停止了。
ISA|63|16|亞伯拉罕 雖然不承認我們， 以色列 也不承認我們， 你卻是我們的父。 耶和華啊，你是我們的父； 自古以來，你的名是「我們的救贖主」。
ISA|63|17|耶和華啊，你為何使我們偏離你的道， 使我們心裏剛硬、不敬畏你呢？ 求你為你的僕人， 為你產業的支派而回轉。
ISA|63|18|你的聖民暫時得你的聖所， 但我們的敵人踐踏了它。
ISA|63|19|我們就成了你未曾治理的人， 成了未曾稱為你名下的人。
ISA|64|1|願你破天而降， 願山在你面前震動，
ISA|64|2|好像火燒乾柴， 又如火將水燒開， 使你敵人知道你的名， 列國必在你面前發顫！
ISA|64|3|你曾做我們不能逆料可畏的事； 那時你降臨，山嶺在你面前震動。
ISA|64|4|自古以來，人未曾聽見，未曾耳聞，未曾眼見， 除你以外，還有上帝能為等候他的人行事。
ISA|64|5|你迎見那歡喜行義、記念你道的人； 看哪，你曾發怒，因我們犯了罪； 這景況已久，我們還能得救嗎？
ISA|64|6|我們都如不潔淨的人， 所行的義都像污穢的衣服。 我們如葉子漸漸枯乾， 罪孽像風把我們吹走。
ISA|64|7|無人求告你的名， 無人奮力抓住你。 你轉臉不顧我們， 你使我們因罪孽而融化 。
ISA|64|8|但耶和華啊，現在你仍是我們的父！ 我們是泥，你是陶匠； 我們都是你親手所造的。
ISA|64|9|耶和華啊，求你不要大發震怒， 也不要永遠記得罪孽； 看哪，求你垂顧我們， 因我們都是你的百姓。
ISA|64|10|你的聖城已變為曠野； 錫安 變為曠野， 耶路撒冷 成為廢墟。
ISA|64|11|我們那神聖華美的殿， 就是我們祖先讚美你的地方，已被火焚燒； 我們所羨慕的美地盡都荒蕪。
ISA|64|12|耶和華啊，有這些事，你還能忍受嗎？ 你還靜默，使我們大受苦難嗎？
ISA|65|1|沒有求問我的，我要讓他們找到； 沒有尋找我的，我要讓他們尋見； 我對沒有呼求我名的國 說： 「我在這裏！我在這裏！」
ISA|65|2|我整天向那悖逆的百姓招手， 他們隨自己的意念行不善之道。
ISA|65|3|這百姓時常當面惹我發怒， 在園中獻祭， 在磚上燒香，
ISA|65|4|在墳墓間停留， 在隱密處過夜， 吃豬肉， 器皿中有不潔淨之肉熬的湯；
ISA|65|5|且對人說：「你站開吧！ 不要挨近我，因為我對你來說太神聖了 。」 這些人惹我鼻中冒煙， 如終日燃燒的火。
ISA|65|6|看哪，這些都寫在我面前。 我必不靜默，卻要施行報應， 將你們和你們祖先的罪孽 全都報應在後人身上； 因為他們在山上燒香， 在岡上褻瀆我， 我要按他們先前所行的，報應在他們身上 ； 這是耶和華說的。
ISA|65|7|
ISA|65|8|耶和華如此說： 「人在葡萄中尋得新酒時會說： 『不要毀壞它，因為它還有用處』； 同樣，我必因我僕人的緣故， 不將他們全然毀滅。
ISA|65|9|我必從 雅各 中領出後裔， 從 猶大 中領出那要繼承我眾山的； 我的選民要繼承它， 我的僕人要在那裏居住。
ISA|65|10|沙崙 必成為羊群的圈， 亞割谷 成為牛群躺臥之處， 都為尋求我的民所得。
ISA|65|11|但你們這些離棄耶和華， 就是忘記我的聖山、 為『幸運之神』擺設筵席、 為『命運之神』裝滿調和酒的，
ISA|65|12|我命定你們歸於刀下， 你們都要屈身被殺； 因為我呼喚，你們不回應； 我說話，你們不聽從； 反倒做我眼中看為惡的事， 選擇我所不喜悅的事。」
ISA|65|13|所以，主耶和華如此說： 「看哪，我的僕人必得吃，你們卻飢餓； 看哪，我的僕人必得喝，你們卻乾渴； 看哪，我的僕人必歡喜，你們卻蒙羞。
ISA|65|14|看哪，我的僕人因心中喜樂而歡呼， 你們卻因心裏悲痛而哀哭， 因靈裏憂傷而哀號。
ISA|65|15|你們必留下自己的名 給我選民指著賭咒： 主耶和華必殺你們， 另起別名稱呼他的僕人。
ISA|65|16|在地上為自己求福的， 必憑真實的上帝求福； 在地上起誓的， 必指著真實的上帝起誓。 因為從前的患難已被遺忘， 從我眼前消逝。」
ISA|65|17|「看哪，我造新天新地！ 從前的事不再被記念，也不被人放在心上；
ISA|65|18|當因我所造的歡喜快樂，直到永遠； 看哪，因為我造 耶路撒冷 為人所喜， 造其中的居民為人所樂。
ISA|65|19|我必因 耶路撒冷 歡喜， 因我的百姓快樂， 那裏不再聽見哭泣和哀號的聲音。
ISA|65|20|那裏沒有數日夭折的嬰孩， 也沒有壽數不滿的老人； 因為百歲死的仍算孩童， 未達百歲而亡的 算是被詛咒的。
ISA|65|21|他們建造房屋，居住其中， 栽葡萄園，吃園中的果子；
ISA|65|22|並非造了給別人居住， 也非栽種給別人享用； 因為我百姓的日子必長久如樹木， 我的選民必享受親手勞碌得來的。
ISA|65|23|他們必不徒然勞碌， 所生產的，也不遭災害， 因為他們和他們的子孫 都是蒙耶和華賜福的後裔。
ISA|65|24|他們尚未求告，我就應允； 正說話的時候，我就垂聽。
ISA|65|25|野狼必與羔羊同食， 獅子必吃草，與牛一樣， 蛇必以塵土為食物； 在我聖山的遍處， 牠們都不傷人，也不害物； 這是耶和華說的。」
ISA|66|1|耶和華如此說： 「天是我的座位； 地是我的腳凳。 你們能為我造怎樣的殿宇呢？ 哪裏是我安歇的地方呢？
ISA|66|2|這一切是我手所造的， 這一切就都存在了。 我所看顧的是困苦、靈裏痛悔、 因我言語而戰兢的人。 這是耶和華說的。
ISA|66|3|「至於那些宰牛，殺人， 獻羔羊，打斷狗頸項， 獻豬血為供物， 燒乳香，稱頌偶像的， 他們選擇自己的道路， 心裏喜愛可憎惡的事；
ISA|66|4|我也必選擇苦待他們， 使他們所懼怕的臨到他們； 因為我呼喚，無人回應； 我說話，他們不聽從； 反倒做我眼中看為惡的事， 選擇我所不喜悅的事。」
ISA|66|5|你們因耶和華言語而戰兢的人哪，當聽他的話： 「你們的弟兄，就是恨惡你們， 因我名趕出你們的，曾說： 『願耶和華彰顯榮耀 ， 好讓我們看見你們的喜樂。』 但蒙羞的終究是他們！
ISA|66|6|「有喧嘩的聲音出自城中！ 有聲音來自殿裏！ 是耶和華向仇敵施行報應的聲音！
ISA|66|7|「 錫安 未曾陣痛就生產， 疼痛尚未來到，就生出男孩。
ISA|66|8|國豈能一日而生？ 民豈能一時而產？ 但 錫安 一陣痛就生下兒女， 這樣的事有誰聽見， 有誰看見呢？
ISA|66|9|耶和華說：我使人臨產， 豈不讓她 生產呢？ 你的上帝說：我使人生產， 難道還讓她關閉 不生嗎？
ISA|66|10|「你們所有愛慕 耶路撒冷 的啊， 要與她一同歡喜，為她高興； 你們所有為她悲哀的啊， 都要與她一同樂上加樂；
ISA|66|11|使你們在她安慰的懷中吃奶得飽， 盡情吸取她豐盛的榮耀，滿心喜樂。」
ISA|66|12|耶和華如此說： 「看哪，我要使平安臨到她，好像江河； 使列國的榮耀及於她，如同漲溢的溪流。 你們要盡情吸吮； 你們必被抱在身旁 ，搖弄在膝上。
ISA|66|13|我要安慰你們，如同母親安慰兒女； 你們也必在 耶路撒冷 得安慰。
ISA|66|14|你們看見，心裏就喜樂， 你們的骨頭必如草生長； 耶和華的手在他僕人身上彰顯， 他卻要向他的仇敵發怒。」
ISA|66|15|看哪，耶和華必在火中降臨， 他的戰車宛如暴風， 以烈怒施行報應， 以火焰施行責罰；
ISA|66|16|耶和華必以火與刀審判凡有血肉之軀的， 被耶和華所殺的很多。
ISA|66|17|那些潔淨自己獻給偶像，進入園內，跟隨其中一個人去吃豬肉和鼠肉，並可憎之物的，他們必一同滅絕。這是耶和華說的。
ISA|66|18|我知道他們的行為和他們的意念。聚集萬國萬族 的時候到了 ，他們要來瞻仰我的榮耀；
ISA|66|19|我要在他們中間顯神蹟，差遣他們當中的倖存者到列國去，就是到 他施 、 普勒 、以善射聞名的 路德 、 土巴 、 雅完 ，和未曾聽見我名聲，未曾看見我榮耀的遙遠海島那裏去；他們必在列國中傳揚我的榮耀。
ISA|66|20|他們要將你們的弟兄從列國中帶回，或騎馬，或坐車，或乘蓬車，或騎騾子，或騎獨峰駝，到我的聖山 耶路撒冷 ，作為供物獻給耶和華。這是耶和華說的。正如 以色列 人用潔淨的器皿盛供物奉到耶和華的殿中，
ISA|66|21|我也必從他們中間立人作祭司，作 利未 人。這是耶和華說的。
ISA|66|22|「我所造的新天新地在我面前長存， 你們的後裔和你們的名號也必照樣長存。 這是耶和華說的。
ISA|66|23|每逢初一、安息日， 凡有血肉之軀的必前來，在我面前下拜； 這是耶和華說的。
ISA|66|24|「他們要出去觀看那些違背我的人的屍首， 他們的蟲是不死的， 他們的火是不滅的， 凡有血肉之軀的都必憎惡他們。」
JER|1|1|這些是 便雅憫 地 亞拿突城 的祭司， 希勒家 的兒子 耶利米 的話。
JER|1|2|亞們 的兒子 猶大 王 約西亞 在位第十三年，耶和華的話臨到 耶利米 。
JER|1|3|從 約西亞 的兒子 猶大 王 約雅敬 在位的時候，直到 約西亞 的兒子 猶大 王 西底家 在位的末年，就是第十一年五月間 耶路撒冷 被擄時，耶和華的話也常臨到 耶利米 。
JER|1|4|耶利米 說，耶和華的話臨到我，說：
JER|1|5|「我尚未將你造在母腹中，就已認識你； 你未出母胎，我已將你分別為聖， 派你作列國的先知。」
JER|1|6|我就說：「唉，主耶和華！看哪，我不知道怎麼說，因為我年輕。」
JER|1|7|耶和華對我說： 「不要說：『我年輕』， 因為我差遣你到誰那裏去，你都要去； 我吩咐你說甚麼話，你都要說。
JER|1|8|你不要怕他們， 因為我與你同在，要拯救你。 這是耶和華說的。」
JER|1|9|於是耶和華伸手按住我的口， 對我說： 「看哪，我已將我的話放在你口中。
JER|1|10|我今日立你在列邦列國之上， 為要拔出，拆毀，毀壞，傾覆， 又要建立，栽植。」
JER|1|11|耶和華的話臨到我，說：「 耶利米 ，你看見甚麼？」我說：「我看見一根杏樹枝。」
JER|1|12|耶和華對我說：「你看得不錯；因為我要看守 我的話，使它實現。」
JER|1|13|耶和華的話第二次臨到我，說：「你看見甚麼？」我說：「我看見一個水燒開的鍋，從北而傾。」
JER|1|14|耶和華對我說：「必有災禍從北方發出，臨到這地所有的居民。
JER|1|15|看哪，我要召北方列國的萬族。這是耶和華說的。他們要來，各安寶座在 耶路撒冷 的城門口，周圍攻擊城牆，又要攻擊 猶大 的一切城鎮。
JER|1|16|這百姓離棄我，向別神燒香，跪拜自己手所造的，我要針對這一切惡行，向他們宣讀我的判決。
JER|1|17|所以你當束腰，起來，將我所吩咐你的一切話都告訴他們；不要因他們驚惶，免得我使你在他們面前驚惶。
JER|1|18|看哪，我今日使你成為堅城、鐵柱、銅牆，對抗全地和 猶大 的君王、官長、祭司，並這地的百姓。
JER|1|19|他們要攻擊你，卻不能勝過你，因為我與你同在，要拯救你。這是耶和華說的。」
JER|2|1|耶和華的話臨到我，說：
JER|2|2|「你去向 耶路撒冷 居民的耳朵呼喊說，耶和華如此說： 『你年輕時的恩愛， 新婚時的愛情， 你怎樣在曠野， 在未耕種之地跟隨我， 我都記得。
JER|2|3|那時 以色列 歸耶和華為聖， 作為他初熟的土產； 凡吞吃它的必算為有罪， 災禍必臨到他們。 這是耶和華說的。』」
JER|2|4|雅各 家， 以色列 家的各族啊，當聽耶和華的話，
JER|2|5|耶和華如此說： 「你們的祖先看我有甚麼錯處， 竟遠離我，隨從那虛無的神明 ， 自己成為虛無呢？
JER|2|6|他們並不問： 『那領我們從 埃及 地上來， 引導我們走過曠野、沙漠有坑洞之地， 走過乾旱死蔭、無人經過、 無人居住之地的耶和華在哪裏呢？』
JER|2|7|我領你們進入肥沃之地， 使你們得吃其中的果子和美物； 你們進入時，卻使我的地玷污， 使我的產業成為可憎惡的。
JER|2|8|祭司從來不問：『耶和華在哪裏呢？』 傳講律法的不認識我， 官長違背我， 先知藉 巴力 說預言， 隨從無益的東西。」
JER|2|9|「我因此必與你們爭辯， 也與你們的子孫爭辯。 這是耶和華說的。
JER|2|10|你們且渡到 基提 海島察看， 派人往 基達 去留心查考， 看可曾有過這樣的事。
JER|2|11|豈有一國換了它的神明嗎？ 其實那不是神明！ 但我的百姓將他們的榮耀換了那無益的東西。
JER|2|12|諸天哪，要因此震驚， 顫慄，極其淒涼！ 這是耶和華說的。
JER|2|13|因為我的百姓做了兩件惡事： 離棄我這活水的泉源； 又為自己鑿出水池， 卻是破裂不能儲水的池子。」
JER|2|14|「 以色列 是僕人嗎？ 是家中生的奴僕嗎？ 為何成為掠物呢？
JER|2|15|少壯獅子向它咆哮，大聲吼叫， 使它的地荒蕪； 城鎮燒燬，無人居住。
JER|2|16|挪弗 人和 答比匿 人打破你的頭顱。
JER|2|17|這不是你自己招惹的嗎？ 不是因耶和華－你上帝引導你行路時， 你離棄了他嗎？
JER|2|18|現今你為何在 埃及 路上喝 西曷河 的水呢？ 為何在 亞述 路上喝 大河 的水呢？
JER|2|19|你自己的惡必懲治你， 你背道的事必責罰你。 由此可知可見，你離棄耶和華－你的上帝， 不存敬畏我的心， 實為惡事，為苦事； 這是萬軍之主耶和華說的。」
JER|2|20|「你 在古時折斷你的軛，解開你的繩索， 說：『我必不事奉耶和華 。』 你在各高岡上、各青翠的樹下屈身行淫。
JER|2|21|然而，我栽種你為上等的葡萄樹， 全用純正的種子； 你怎麼向我變為外邦葡萄樹的壞枝子呢？
JER|2|22|你雖用鹼、多用皂莢清洗， 你罪孽的痕跡仍顯在我面前。 這是主耶和華說的。
JER|2|23|你怎能說： 『我沒有玷污，沒有隨從 巴力 』？ 看看你在谷中所做的，思想你自己的所作所為； 你是快行的獨峰駝，狂奔亂闖。
JER|2|24|你是野驢，習慣曠野， 慾心發動時就呼吸急促， 發情時誰能使牠轉回呢？ 凡尋找牠的必不費力， 在牠的季節必能尋見牠。
JER|2|25|你不要弄到赤足而行， 喉嚨乾渴。 你卻說：『沒有用的， 我喜愛陌生人， 我必隨從他們。』」
JER|2|26|「賊被捉拿，怎樣羞愧， 以色列 家和他們的君王、官長、 祭司、先知也都照樣羞愧。
JER|2|27|他們向木頭說：『你是我的父』； 向石頭說：『你是生我的。』 他們以背向我， 不肯以面向我； 及至遭遇患難時卻說： 『起來拯救我們吧！』
JER|2|28|你為自己做的神明在哪裏呢？ 你遭遇患難的時候， 讓它們起來拯救你吧！ 猶大 啊，你神明的數目與你城的數目相等。
JER|2|29|「你們為何與我爭辯呢？ 你們都違背了我。 這是耶和華說的。
JER|2|30|我責打你們的兒女是徒然的， 他們不受管教。 你們自己的刀吞滅你們的先知， 好像殘害人的獅子。
JER|2|31|這世代的人哪， 你們要留意耶和華的話。 我向 以色列 豈是曠野， 或幽暗之地呢？ 我的百姓為何說： 『我們脫離約束，不再歸向你了』？
JER|2|32|少女豈能忘記她的妝飾呢？ 新娘豈能忘記她的美衣呢？ 我的百姓卻在無數的日子裏忘記了我！
JER|2|33|「你竟然如此精於求愛之道， 可把你的門徑教邪惡的女人！
JER|2|34|你衣服的邊上有無辜貧窮人的血， 其實你並未發現他們挖洞進屋偷竊 。 雖有這一切的事 ，
JER|2|35|你還說：『我無辜； 耶和華的怒氣必定轉離我了。』 看哪，我必審問你； 因你自己說：『我沒有犯罪。』
JER|2|36|你為何東奔西跑改變你的道路呢？ 你必因 埃及 蒙羞， 像從前因 亞述 蒙羞一樣。
JER|2|37|你也必兩手抱頭離開這裏； 因為耶和華已經棄絕你所倚靠的， 你不能因他們而得順利。」
JER|3|1|耶和華說 ：「人若休妻， 妻離他而去，做了別人的妻子， 前夫豈能再回到她那裏呢？ 那地豈不是大大污穢了嗎？ 但你和許多情郎行淫， 還是可以回到我這裏。 這是耶和華說的。
JER|3|2|你舉目向光禿的高地觀看， 何處沒有你的淫行呢？ 你坐在道路旁等候， 好像 阿拉伯 人在曠野埋伏， 你的淫行和邪惡使全地污穢了。
JER|3|3|因此甘霖停止， 春雨不降。 你還是一副娼妓之臉， 不顧羞恥。
JER|3|4|你不是才向我呼叫說： 『我父啊，你是我年輕時的密友，
JER|3|5|人豈永遠懷恨，長久存怒嗎？』 看哪，你雖這樣說，還是竭盡所能去行惡。」
JER|3|6|約西亞 王在位的時候，耶和華對我說：「你看見背道的 以色列 所做的嗎？她上到各高山，在各青翠的樹下行淫。
JER|3|7|我說：『她行這些事以後會回轉歸向我』，她卻不回轉。她奸詐的妹妹 猶大 也看見了。
JER|3|8|我看見背道的 以色列 行淫，我為這緣故給她休書休了她，她奸詐的妹妹 猶大 還不懼怕，也去行淫。
JER|3|9|因 以色列 輕忽了她的淫亂，與石頭和木頭行姦淫 ，她和這地就都污穢了 。
JER|3|10|雖有這一切的事，她奸詐的妹妹 猶大 還不一心歸向我，不過是假意歸我。這是耶和華說的。」
JER|3|11|耶和華對我說：「背道的 以色列 比奸詐的 猶大 還顯為義。
JER|3|12|你去向北方宣告這些話，說： 『背道的 以色列 啊，回來吧！ 這是耶和華說的。 我必不怒目看你們， 因為我是慈愛的， 這是耶和華說的。 我必不永遠懷怒；
JER|3|13|只要你承認你的罪孽， 就是違背耶和華－你的上帝， 在各青翠的樹下追逐外族的神明 ， 沒有聽從我的話。 這是耶和華說的。
JER|3|14|背道的兒女啊，回來吧！ 這是耶和華說的。 因為我作你們的丈夫， 要將你們從一城取一人， 從一族取兩人，帶到 錫安 。
JER|3|15|「『我必將合我心意的牧者賞賜給你們，他們要以知識和智慧牧養你們。
JER|3|16|你們在國中生養眾多的時候，那些日子，人必不再提說耶和華的約櫃，不追想，不記念，不覺缺少，也不再製造。這是耶和華說的。
JER|3|17|那時，人必稱 耶路撒冷 為耶和華的寶座；萬國聚集在那裏，為耶和華的名來到 耶路撒冷 ，他們必不再隨從自己頑梗的惡心行事。
JER|3|18|當那些日子， 猶大 家要和 以色列 家同行，從北方之地一同來到我所賜給你們祖先為業之地。』」
JER|3|19|我說，我多麼樂意把你列在兒女之中， 賜給你美地， 就是萬國中最美的產業。 我說，你會以「我父啊」稱呼我， 不再轉離而跟從我。
JER|3|20|以色列 家啊，你們向我行詭詐， 真像妻子行詭詐離開丈夫。 這是耶和華說的。
JER|3|21|有聲音從光禿的高地傳來， 就是 以色列 人哭泣懇求的聲音， 因為他們走彎曲之道， 忘記耶和華－他們的上帝。
JER|3|22|「你們這背道的兒女啊，回來吧！ 我要醫治你們背道的病。」 「看哪，我們來到你這裏， 因你是耶和華－我們的上帝。
JER|3|23|從小山來的真是枉然， 大山的喧嚷也是枉然 。 以色列 得救，誠然在乎耶和華－我們的上帝。
JER|3|24|「從我們幼年以來，那可恥之物 吞吃了我們祖先勞碌得來的，就是他們的羊群、牛群和他們的兒女。
JER|3|25|我們在羞恥中躺臥吧！願慚愧將我們遮蓋！因為從我們幼年以來，我們和我們的祖先都得罪了耶和華－我們的上帝，沒有聽從耶和華－我們上帝的話。」
JER|4|1|耶和華說：「 以色列 啊， 你若回轉，回轉歸向我， 若從我眼前除掉你可憎的偶像， 不再猶疑不定，
JER|4|2|憑誠實、公平、公義 指著永生的耶和華起誓； 列國就必因他蒙福， 也必因他誇耀。」
JER|4|3|耶和華對 猶大 人和 耶路撒冷 人如此說： 「你們要為自己開墾荒地， 不要撒種在荊棘裏。
JER|4|4|猶大 人和 耶路撒冷 的居民哪， 你們當自行割禮，歸耶和華， 將你們心裏的污穢 除掉； 免得我的憤怒因你們的惡行發作， 如火燃起， 甚至無人能熄滅！」
JER|4|5|你們要在 猶大 傳揚， 在 耶路撒冷 宣告，說： 「當在國中吹角，高聲呼叫說： 『你們當聚集！ 我們好進入堅固城！』
JER|4|6|應當向 錫安 豎立大旗。 逃吧，不要遲延， 因我必使災禍與大毀滅從北方來到。
JER|4|7|有獅子從密林中上來， 是毀壞列國的。 牠已動身出離本處， 要使你的地荒涼， 使你的城鎮變為廢墟，無人居住。
JER|4|8|因此，你們當腰束麻布，哭泣哀號， 因為耶和華的烈怒並未轉離我們。」
JER|4|9|耶和華說：「到那時，君王和領袖的心要失喪，祭司都要驚奇，先知都要詫異。」
JER|4|10|我說：「哀哉！主耶和華啊，你真是大大欺哄這百姓和 耶路撒冷 ，說：『你們必得平安。』其實刀劍已經抵住喉嚨了！」
JER|4|11|那時，必有話對這百姓和 耶路撒冷 說：「來自曠野光禿高地的熱風吹向我的百姓 ，不是為簸揚，也不是為揚淨。
JER|4|12|又有一陣比這更大的風向我颳來；現在，我要向他們宣讀我的判決。」
JER|4|13|看哪，他必如雲湧上； 他的戰車如旋風， 他的馬比鷹更快。 我們有禍了！ 我們敗落了！
JER|4|14|耶路撒冷 啊，你當洗去心中的惡， 使你可以得救。 惡念在你裏面要存到幾時呢？
JER|4|15|有聲音從 但 傳出， 有災禍從 以法蓮山 傳來。
JER|4|16|你們當傳給列國， 看哪，要向 耶路撒冷 報告： 「有圍攻的人從遠方來到， 向 猶大 的城鎮大聲喊叫。
JER|4|17|他們包圍 耶路撒冷 ， 好像看守田園的， 因為它背叛了我。 這是耶和華說的。
JER|4|18|你的作風和行為招惹這事； 這是你罪惡的結果， 實在是苦， 刺透了你的心！」
JER|4|19|我的肺腑啊，我的肺腑啊，我心疼痛！ 我的心在我裏面煩躁不安。 我不能靜默不言， 因我已聽見角聲和打仗的喊聲。
JER|4|20|毀壞的信息不斷傳來， 因為全地荒廢。 我的帳棚忽然毀壞， 我的幔子頃刻破裂。
JER|4|21|我看見大旗，聽見角聲， 要到幾時呢？
JER|4|22|「我的百姓愚頑，不認識我； 他們是愚昧無知的兒女， 有智慧行惡，沒有知識行善。」
JER|4|23|我觀看地， 看哪，地是空虛混沌； 我觀看天，天也無光。
JER|4|24|我觀看大山，看哪，盡都震動， 小山也都搖來搖去。
JER|4|25|我觀看，看哪，無人； 空中的飛鳥也都躲避。
JER|4|26|我觀看，看哪，肥田變為荒地； 所有城鎮在耶和華面前， 因他的烈怒都被拆毀。
JER|4|27|耶和華如此說：「全地必然荒涼， 我卻不毀滅淨盡。
JER|4|28|因此，地要悲哀， 天上也必黑暗； 因為我言已出，我意已定， 必不改變，也不由此轉回。」
JER|4|29|各城的人因騎兵和弓箭手的響聲就都逃跑， 進入密林，爬上磐石； 城鎮都被拋棄， 無人住在其中。
JER|4|30|你這被毀滅的啊， 你要做甚麼呢？ 你穿上朱紅衣服， 佩戴黃金飾物， 用眼影修飾眼睛， 徒然美化你自己。 戀慕你的卻藐視你， 尋索你的性命。
JER|4|31|我聽見彷彿婦人臨產的聲音， 好像生頭胎疼痛的聲音， 原來是 錫安 的聲音； 她喘著氣，伸開手： 「我有禍了！ 在殺人者跟前，我的心靈發昏。」
JER|5|1|你們要走遍 耶路撒冷 的街市， 在廣場尋找， 看是否有人行公平、求誠實； 若有，我就赦免這城。
JER|5|2|雖然他們說「我對永生的耶和華發誓」， 所起的誓實在是假的。
JER|5|3|耶和華啊，你的眼目不是在尋找誠實嗎？ 你擊打他們，他們卻不傷慟； 你摧毀他們，他們仍不領受管教。 他們使臉剛硬過於磐石， 不肯回頭。
JER|5|4|我說：「這些人實在是貧寒的， 他們是愚昧的， 因為不知道耶和華的作為， 也不知道他們上帝的法則。
JER|5|5|我要去見尊貴的人，向他們說話， 他們應該知道耶和華的作為， 知道他們上帝的法則。」 然而，這些人卻齊心將軛折斷， 掙開繩索。
JER|5|6|因此，林中的獅子必害死他們， 野地的狼必滅絕他們， 豹子在城外窺伺。 凡出城的必被撕碎， 因為他們的罪過極多， 背道的事也增加。
JER|5|7|我怎能赦免你呢？ 你的兒女離棄我， 又指著那不是上帝的起誓。 我使他們飽足， 他們就行姦淫， 居住 在娼妓家裏。
JER|5|8|他們如餵飽的馬，精力旺盛， 各向鄰舍的妻子吹哨。
JER|5|9|我豈不因這些事施行懲罰嗎？ 像這樣的國家，我豈能不報復呢？ 這是耶和華說的。
JER|5|10|你們要上去毀壞它的葡萄園， 但不可毀壞淨盡， 只可除掉其枝子， 因為不屬耶和華。
JER|5|11|以色列 家和 猶大 家向我大行詭詐。 這是耶和華說的。
JER|5|12|關乎耶和華他們說了虛謊的話： 「他不會的， 災禍必不臨到我們， 我們也不會遇見刀劍和饑荒。
JER|5|13|先知不過是一陣風， 道也不在他們裏面； 這災禍必臨到他們身上。」
JER|5|14|所以耶和華－萬軍之上帝如此說： 「因為他們說這話， 看哪，我必使我的話在你口中為火， 使這百姓為柴， 火便將他們燒滅。
JER|5|15|以色列 家啊， 看哪，我必使一國從遠方來攻擊你， 是強盛的國， 是古老的國； 他們的言語你不知道， 所說的話你不明白。 這是耶和華說的。
JER|5|16|他們的箭袋有如敞開的墳墓， 他們全都是勇士。
JER|5|17|他們必吃盡你的莊稼和糧食， 是你兒女該吃的 ； 必吃盡你的牛羊， 吃盡你的葡萄和無花果； 又必用刀劍毀壞你所倚靠的堅固城。
JER|5|18|「就是在那些日子，我也不會將你們毀滅淨盡。這是耶和華說的。
JER|5|19|百姓若說：『耶和華－我們的上帝為甚麼向我們行這一切事呢？』你就對他們說：『你們怎樣離棄我，在你們的地上事奉外邦神明，也必照樣在不屬你們的地上事奉外族人。』」
JER|5|20|當在 雅各 家傳揚， 在 猶大 宣告，說：
JER|5|21|「愚昧無知的百姓啊， 你們有眼不看， 有耳不聽， 現在當聽這話。
JER|5|22|你們難道不懼怕我嗎？ 在我面前還不戰兢嗎？ 這是耶和華說的。 我以沙為海的界限， 作永遠的條例，使它不得越過。 波浪洶湧，卻不能勝過； 怒濤澎湃，仍無法越過。
JER|5|23|但這百姓有背叛忤逆的心， 他們轉離而去。
JER|5|24|他們心裏並不說： 『我們應當敬畏耶和華－我們的上帝； 他按時賜雨，就是秋雨和春雨， 又為我們定收割的季節。』
JER|5|25|你們的罪孽使這些轉離你們， 你們的罪惡使你們不能得福。
JER|5|26|在我百姓當中有惡人， 他們埋伏，好像捕鳥的人在窺探 ； 他們設羅網陷害人。
JER|5|27|籠子怎樣裝滿雀鳥， 他們的屋裏也照樣充滿詭詐； 他們因此得以強大富足。
JER|5|28|他們肥胖光潤，作惡過甚， 不為人伸冤， 不為孤兒伸冤，使他們勝訴， 也不為貧窮人辯護。
JER|5|29|我豈不因這些事施行懲罰嗎？ 像這樣的國家，我豈能不報復呢？ 這是耶和華說的。
JER|5|30|「國中有令人驚駭、 恐怖的事發生，
JER|5|31|先知說假預言， 祭司把權柄抓在自己手上， 我的百姓也喜愛這樣， 到了結局你們要怎麼辦呢？」
JER|6|1|便雅憫 人哪，當逃離 耶路撒冷 ， 在 提哥亞 吹號角， 在 伯‧哈基琳 升信號， 因為有災禍與大毀滅從北方逼近。
JER|6|2|那秀美嬌嫩的 錫安 ， 我必剪除。
JER|6|3|牧人必引領羊群到它那裏， 在它周圍支搭帳棚， 各在自己的地方放牧。
JER|6|4|「你們要準備攻擊它。 起來吧，我們要趁正午上去。」 「哀哉！日已漸斜， 黃昏的影子拖長了。」
JER|6|5|「起來吧，我們要在夜間上去， 毀壞它的宮殿。」
JER|6|6|萬軍之耶和華如此說： 「你們要砍伐樹木， 建土堆攻打 耶路撒冷 ， 就是那該受罰的城 ， 其中盡是欺壓。
JER|6|7|井怎樣湧出水來， 這城也照樣湧出惡來； 其中常聽聞殘暴毀滅的事， 病痛損傷也常在我面前。
JER|6|8|耶路撒冷 啊，當受管教， 免得我心與你生疏， 免得我使你荒涼， 成為無人居住之地。」
JER|6|9|萬軍之耶和華如此說： 「他們洗劫 以色列 剩下的民， 如摘淨葡萄一樣； 現你的手如採收葡萄的人，在樹枝上採了又採 。」
JER|6|10|現在我可以向誰說話，警告誰，使他們聽呢？ 看哪，他們的耳朵未受割禮，不能聽見。 看哪，他們以耶和華的話為羞辱， 不以為喜悅。
JER|6|11|因此我被耶和華的憤怒充滿，難以忍受。 「你要把它倒在街上孩童 和成群的年輕人身上， 他們連夫帶妻， 年長者與高齡的人都必被擒拿。
JER|6|12|他們的房屋、田地， 和妻子都要一起轉歸別人， 我要伸手攻擊這地的居民。」 這是耶和華說的。
JER|6|13|「因為他們從最小的到最大的都貪圖不義之財， 從先知到祭司全都行事虛假。
JER|6|14|他們輕忽地醫治我百姓的損傷， 說：『平安了！平安了！』 其實沒有平安。
JER|6|15|他們行可憎之事，應當羞愧； 然而他們卻一點也不覺得羞愧， 也不知羞恥。 因此，他們必與仆倒的人一同仆倒， 我懲罰他們的時候， 他們必跌倒。」 這是耶和華說的。
JER|6|16|耶和華如此說： 「你們當站在路邊察看， 尋訪古老的路， 哪裏是完善的道路，就行走在其上； 這樣，你們自己必找到安息。 他們卻說：『我們不走。』
JER|6|17|我為你們設立守望的人， 要留心聽角聲。 他們卻說：『我們不聽。』
JER|6|18|因此，列國啊，當聽！ 會眾啊，要知道他們必遭遇的事。
JER|6|19|地啊，當聽！ 看哪，我必使災禍臨到這百姓， 是他們計謀所結的果子； 因為他們不肯留心聽我的話， 至於我的律法，他們也厭棄。
JER|6|20|從 示巴 來的乳香， 從遠方出的香菖蒲， 奉來給我有何用呢？ 你們的燔祭不蒙悅納； 你們的祭物，我也不喜悅。」
JER|6|21|所以耶和華如此說： 「看哪，我要將絆腳石放在這百姓面前； 父親和兒子要一同跌在其上， 鄰舍與朋友也都滅亡。」
JER|6|22|耶和華如此說： 「看哪，有一民族從北方而來； 有一大國被激起，從地極來到。
JER|6|23|他們拿弓和槍， 性情殘忍，不施憐憫； 他們的聲音如海浪澎湃。 錫安 哪， 他們都騎馬， 如上戰場的人擺陣攻擊你。」
JER|6|24|我們聽見這樣的風聲，手就發軟； 痛苦將我們抓住， 疼痛彷彿臨產的婦人。
JER|6|25|你們不要出到田野去， 也不要行走在路上， 因四圍有仇敵的刀劍和驚嚇。
JER|6|26|我的百姓 啊，應當腰束麻布，滾在灰中。 要悲傷，如喪獨子般痛痛哭號， 因為滅命的忽然臨到我們。
JER|6|27|我使你作我百姓的測試者 和考驗者 ， 使你知道並考驗他們的行為。
JER|6|28|他們極其悖逆， 到處毀謗人， 他們是銅是鐵， 全都敗壞了。
JER|6|29|風箱吹火，鉛被燒燬， 煉而又煉，終是徒然， 因為惡劣的還未除掉。
JER|6|30|人必稱他們為被拋棄的銀子， 因為耶和華已經拋棄了他們。
JER|7|1|耶和華的話臨到 耶利米 ，說：
JER|7|2|「你當站在耶和華殿的門口，在那裏宣講這話說：所有從這些門進來敬拜耶和華的 猶大 人哪，當聽耶和華的話。
JER|7|3|萬軍之耶和華－ 以色列 的上帝如此說：你們要改正你們的所作所為，我就使你們仍然居住這地 。
JER|7|4|不要倚靠虛謊的話，說：『這是耶和華的殿，是耶和華的殿，是耶和華的殿！』
JER|7|5|「你們若實在改正你們的所作所為，彼此誠然施行公平，
JER|7|6|不欺壓寄居的和孤兒寡婦，不在這地方流無辜人的血，也不隨從別神陷害自己，
JER|7|7|我就使你們仍然居住這地 ，就是我從古時所賜給你們祖先的地，從永遠到永遠。
JER|7|8|「看哪，你們倚靠虛謊無益的話語。
JER|7|9|你們豈可偷盜，殺害，姦淫，起假誓，向 巴力 燒香，隨從素不認識的別神，
JER|7|10|又來到這稱為我名下的殿，在我面前敬拜，說『我們平安無事』，為了要行這一切可憎的事呢？
JER|7|11|這稱為我名下的殿在你們眼中豈可看為賊窩呢？看哪，我真的都看見了。這是耶和華說的。
JER|7|12|你們到我的地方 示羅 去，就是我先前在那裏立為我名的居所，察看我因這百姓 以色列 的罪惡向那地方所行的事。
JER|7|13|現在，因你們行了這一切的事，我一再警戒你們，你們卻不聽從；我呼喚你們，你們也不回應。這是耶和華說的。
JER|7|14|所以我要向這稱為我名下、你們所倚靠的殿，與我所賜給你們和你們祖先的地這樣行，正如我從前向 示羅 所行的。
JER|7|15|我必將你們從我眼前趕出，正如趕出你們的眾弟兄，就是所有 以法蓮 的後裔。」
JER|7|16|「所以，你不要為這百姓祈禱；不要為他們呼求禱告，也不要為他們向我祈求，因我不聽你。
JER|7|17|他們在 猶大 城鎮和 耶路撒冷 街上所做的，你難道沒有看見嗎？
JER|7|18|孩子撿柴，父親燒火，婦女揉麵做餅，獻給天后，又向別神獻澆酒祭，惹我發怒。
JER|7|19|他們豈是惹我發怒呢？不是自己惹禍，以致臉上慚愧嗎？這是耶和華說的。
JER|7|20|所以主耶和華如此說：看哪，我必將我的怒氣和憤怒傾倒在這地方的人和牲畜身上、田野的樹木和地裏的出產上，它必燃燒，不會熄滅。」
JER|7|21|萬軍之耶和華－ 以色列 的上帝如此說：「你們要將燔祭加在你們的祭物上，又要吃肉；
JER|7|22|因為我將你們祖先從 埃及 地領出來的那日，燔祭和祭物的事我並沒有提說，也沒有吩咐他們。
JER|7|23|我只吩咐他們這一件事說：『你們當聽從我的話，我就作你們的上帝，你們也作我的子民。你們行走我所吩咐的一切道路，就可以得福。』
JER|7|24|他們卻不聽從，也不側耳而聽，竟隨從自己的計謀和頑梗的惡心去行，不進反退。
JER|7|25|自從你們祖先出 埃及 地的那日，直到今日，我每日一再差遣我的僕人眾先知到你們那裏去。
JER|7|26|你們卻不聽我，不側耳而聽，竟硬著頸項行惡，比你們的祖先更甚。
JER|7|27|「你要將這一切的話告訴他們，他們卻不聽你；呼喚他們，他們卻不回應。
JER|7|28|你要對他們說：『這就是不聽從耶和華－他們上帝的話、不領受訓誨的國民；誠信已從他們口中消失殆盡了。
JER|7|29|耶路撒冷 啊，要剪頭髮，扔掉它， 在光禿的高地唱哀歌， 因為耶和華棄絕、離棄了惹他發怒的世代。』」
JER|7|30|「 猶大 人行我眼中看為惡的事，將可憎之偶像立在稱為我名下的殿裏，玷污這殿。這是耶和華說的。
JER|7|31|他們在 欣嫩子谷 建造 陀斐特 的丘壇，要在火中焚燒自己的兒女。這並不是我所吩咐的，我心裏也從來沒有想過。
JER|7|32|因此，看哪，日子將到，這地方不再稱為 陀斐特 和 欣嫩子谷 ，反倒稱為 殺戮谷 。他們要在 陀斐特 埋葬屍首，甚至無處可葬。這是耶和華說的。
JER|7|33|並且這百姓的屍首要給空中的飛鳥和地上的走獸作食物，無人嚇走牠們。
JER|7|34|那時，我必止息 猶大 城鎮和 耶路撒冷 街上歡喜和快樂的聲音、新郎和新娘的聲音，因為這地必然荒蕪。」
JER|8|1|耶和華說：「那時，人必將 猶大 諸王和領袖的骸骨、祭司和先知的骸骨，以及 耶路撒冷 居民的骸骨，都從墳墓中取出來，
JER|8|2|散佈在太陽、月亮和天上眾星之下，就是他們從前所喜愛、所事奉、所隨從、所求問、所敬拜的。這些骸骨不被收殮，不被埋葬，必在地面上成為糞土。
JER|8|3|這邪惡家族所倖存的餘民，就是在我趕他們到的各處所剩下的 ，全都寧可選死不選活。這是萬軍之耶和華說的。」
JER|8|4|「你要對他們說，耶和華如此說： 人跌倒，不再起來嗎？ 人轉去，不再轉回來嗎？
JER|8|5|這 耶路撒冷 的百姓為何永久背道呢？ 他們抓住詭詐，不肯回頭。
JER|8|6|我留心聽，聽見他們說不誠實的話。 無人懊悔自己的惡行，說： 『我做的是甚麼呢？』 他們全都轉奔己路， 如馬直闖戰場。
JER|8|7|空中的鸛鳥知道自己的季節， 斑鳩、燕子與白鶴也守候當來的時令； 我的百姓卻不知道耶和華的法則。
JER|8|8|「你們怎麼說：『我們有智慧， 耶和華的律法在我們這裏』？ 看哪，其實文士的假筆舞弄虛假。
JER|8|9|智慧人慚愧，驚惶，被擒拿； 看哪，他們背棄耶和華的話， 還會有甚麼智慧呢？
JER|8|10|因此，我必將他們的妻子給別人， 將他們的田地給別人為業； 因為他們從最小的到最大的都貪圖不義之財， 從先知到祭司全都行事虛假。
JER|8|11|他們輕忽地醫治我百姓的損傷，說： 『平安了！平安了！』 其實沒有平安。
JER|8|12|他們行可憎之事，應當羞愧； 然而他們卻一點也不覺得羞愧， 又不知羞恥。 因此，他們必與仆倒的人一樣仆倒； 我懲罰他們的時候， 他們必跌倒。 這是耶和華說的。
JER|8|13|我必使他們全然滅絕； 葡萄樹上必沒有葡萄 ， 無花果樹上沒有果子， 葉子也必枯乾。 我所賜給他們的， 必離他們而去。 這是耶和華說的。」
JER|8|14|我們為何靜坐不動呢？ 我們當聚集，進入堅固城， 在那裏靜默不言； 因為耶和華－我們的上帝使我們靜默不言， 又將苦水給我們喝， 都因我們得罪了耶和華。
JER|8|15|我們指望平安， 卻得不著福氣； 指望痊癒的時刻， 看哪，受了驚惶。
JER|8|16|「從 但 那裏傳來敵人的馬噴氣的聲音， 壯馬發出嘶聲， 全地就都震動； 因為他們來吞滅這地和其上所有的， 吞滅這城與其中的居民。
JER|8|17|看哪，我必派蛇進到你們中間， 就是法術無法驅除的毒蛇， 牠們必咬你們。 這是耶和華說的。」
JER|8|18|憂愁時我尋找安慰 ， 我心在我裏面發昏。
JER|8|19|聽啊，是我百姓呼救的聲音從遠地傳來： 「耶和華不是在 錫安 嗎？ 錫安 的王不是在其中嗎？」 「他們為甚麼以自己雕刻的偶像 和外邦虛無的神明 惹我發怒呢？」
JER|8|20|「秋收已過，夏季已完， 我們還未得救！」
JER|8|21|因我百姓的損傷， 我也受了損傷。 我哀慟，驚惶將我抓住。
JER|8|22|在 基列 豈沒有乳香呢？ 在那裏豈沒有醫生呢？ 我百姓 為何得不著醫治呢？
JER|9|1|但願我的頭為水， 我的眼為淚水的泉源， 我好為我百姓 中被殺的人晝夜哭泣。
JER|9|2|惟願在曠野有旅客的客棧， 我好離開我的百姓而去； 因他們全都行姦淫， 是行詭詐的一黨。
JER|9|3|他們彎起舌頭像弓， 為要說謊話； 他們在國中增長勢力， 不是為誠信。 他們惡上加惡， 並不認識我。 這是耶和華說的。
JER|9|4|你們各人當謹防鄰舍， 不可信賴弟兄； 因為弟兄盡行欺騙， 鄰舍也都往來毀謗人。
JER|9|5|他們互相欺騙， 不說真話， 訓練自己的舌頭說謊， 竭盡所能地作惡。
JER|9|6|你居住在詭詐的人中； 他們因行詭詐 ，不願意認識我。 這是耶和華說的。
JER|9|7|所以萬軍之耶和華如此說： 「看哪，我要熬煉他們，考驗他們； 不然，為了我的百姓 ，我該如何行呢？
JER|9|8|他們的舌頭是毒箭，說話詭詐， 跟鄰舍口說平安， 心卻謀害他。
JER|9|9|我豈不因這些事向他們施行懲罰嗎？ 像這樣的國家，我豈能不報復呢？ 這是耶和華說的。」
JER|9|10|我要為山嶺哭泣悲哀， 為曠野的草場揚聲哀號； 因為都已枯焦，甚至無人經過。 牲畜的鳴叫聽不見， 空中的飛鳥和地上的走獸也都逃離。
JER|9|11|我必使 耶路撒冷 成為廢墟，為野狗的住處， 也必使 猶大 的城鎮荒廢，無人居住。
JER|9|12|誰是智慧人，可以明白這事？耶和華的口可向誰述說，使他傳講呢？這地為何毀滅，枯焦如曠野，無人經過呢？
JER|9|13|耶和華說：「因為這百姓離棄我在他們面前所設立的律法，不聽從我的話，不肯遵行，
JER|9|14|反隨從自己頑梗的心行事，照他們祖先所教訓的隨從諸 巴力 。」
JER|9|15|所以萬軍之耶和華－ 以色列 的上帝如此說：「看哪，我必將茵蔯給這百姓吃，又用苦水給他們喝。
JER|9|16|我要把他們分散在他們和他們祖宗所不認識的列國；我也要使刀劍追殺他們，直到將他們滅盡。」
JER|9|17|萬軍之耶和華如此說： 「你們要考慮， 將唱哀歌的婦女召來， 差人召善哭的婦女前來，
JER|9|18|叫她們速速為我們舉哀， 使我們淚眼汪汪， 使我們的眼皮湧出淚水。
JER|9|19|因為有哀聲從 錫安 傳來： 『我們竟然敗落！ 我們何等慚愧！ 我們撇下土地， 人拆毀了我們的房屋。』」
JER|9|20|婦女們哪，當聽耶和華的話， 領受他口中的言語； 當教導你們的女兒舉哀， 各人教導女伴唱哀歌。
JER|9|21|因為死亡從窗戶進來， 進入我們的宮殿， 從外邊剪除孩童， 從街上剪除少年。
JER|9|22|你當說，耶和華如此說： 人的屍首必倒在田野像糞土， 又像收割的人身後遺落的禾稼， 無人拾取。
JER|9|23|耶和華如此說：「智慧人不要因他的智慧誇口，勇士不要因他的力氣誇口，財主也不要因他的財富誇口；
JER|9|24|誇口的卻要誇自己有聰明，認識我是耶和華，知道我喜悅在世上施行慈愛、公平和公義。這是耶和華說的。
JER|9|25|「看哪，日子將到，這是耶和華說的，我要懲罰只在肉身受割禮的人，
JER|9|26|就是 埃及 、 猶大 、 以東 、 亞捫 人、 摩押 人，和住曠野所有剃鬢髮的人；因為列國都未受割禮， 以色列 全家心中也未受割禮。」
JER|10|1|以色列 家啊，要聽耶和華對你們所說的話，
JER|10|2|耶和華如此說： 「不要效法列國的行為， 任憑列國因天象驚惶， 你們不要驚惶。
JER|10|3|萬民的習俗是虛空的； 偶像 不過是從樹林中砍來的木頭， 是匠人用斧頭做成的手工。
JER|10|4|人用金銀妝飾它， 用釘子和錘子釘穩， 使它不動搖。
JER|10|5|偶像好像瓜田裏的稻草人， 不能說話，不能行走， 必須有人抬著。 不要怕它們， 因它們不能降禍， 也無力降福。」
JER|10|6|耶和華啊，沒有誰能與你相比！ 你本為大，你的名也大有能力。
JER|10|7|萬國的王啊，誰不敬畏你？ 敬畏你本是合宜的； 列國所有的智慧人中， 在他們一切的國度裏， 都沒有能與你相比的。
JER|10|8|他們如同畜牲，盡都愚昧。 偶像的訓誨算甚麼呢？ 偶像不過是木頭，
JER|10|9|錘煉的銀片是從 他施 來的， 金子則從 烏法 而來， 都是匠人和銀匠的手工； 又有藍色和紫色的衣服， 全都是巧匠的作品。
JER|10|10|惟耶和華是真上帝， 是活的上帝，是永遠的王。 他一發怒，大地震動； 他一惱恨，列國擔當不起。
JER|10|11|你們要對他們這樣說：「那些不是創造天地的神明，必從地上、從天下被除滅！」
JER|10|12|耶和華以能力創造大地， 以智慧建立世界， 以聰明鋪張穹蒼。
JER|10|13|他一出聲，天上就有眾水澎湃； 他使雲霧從地極上騰， 造電隨雨而閃， 從倉庫中吹出風來。
JER|10|14|人人都如同畜牲，毫無知識； 銀匠都因偶像羞愧， 他所鑄的偶像本是虛假， 它們裏面並無氣息。
JER|10|15|偶像都是虛無的， 是迷惑人的作品， 到受罰的時刻必被除滅。
JER|10|16|雅各 所得的福分不是這樣， 因主 是那創造萬有的， 以色列 是他產業的支派， 萬軍之耶和華是他的名。
JER|10|17|受圍困的居民哪，當收拾你的行囊， 離開這地。
JER|10|18|因為耶和華如此說： 「看哪，這一次，我必將此地的居民拋出去， 又必加害他們， 使他們覺悟 。」
JER|10|19|禍哉！我受損傷， 我的傷痕極其重大。 我卻說：「這真的是我必須忍受的痛苦。」
JER|10|20|我的帳棚毀壞， 我的繩索折斷， 我的兒女都離我而去，不在了。 再無人來支搭我的帳棚，掛起我的幔子。
JER|10|21|因為牧人如同畜牲， 沒有尋求耶和華， 所以不得順利； 他們的羊群也都分散了。
JER|10|22|有風聲！看哪，來了！ 有大擾亂從北方而來， 要使 猶大 的城鎮變為廢墟， 成為野狗的住處。
JER|10|23|耶和華啊，我知道人的道路不由自己， 行路的人也不能定自己的腳步。
JER|10|24|耶和華啊，求你按公平管教我， 不要在你的怒中懲治我， 免得你使我歸於無有。
JER|10|25|求你將憤怒傾倒在不認識你的列國中， 傾倒在不求告你名的各族上； 因為他們吞了 雅各 ，不但吞吃，而且滅絕， 使他的住處變為荒涼。
JER|11|1|耶和華的話臨到 耶利米 ，說：
JER|11|2|「當聽這約的話，告訴 猶大 人和 耶路撒冷 的居民，
JER|11|3|對他們說，耶和華－ 以色列 的上帝如此說：『不聽從這約之話的人必受詛咒。
JER|11|4|這約是我將你們祖先從 埃及 地領出來，脫離鐵爐的那日所吩咐他們的，說：你們要聽從我的話，照我所吩咐的一切去做。這樣，你們作我的子民，我也作你們的上帝，
JER|11|5|我好堅定我向你們列祖所起的誓，賞賜他們流奶與蜜之地，正如今日一樣。』」我就回應說：「耶和華啊，阿們！」
JER|11|6|耶和華對我說：「你要在 猶大 城鎮和 耶路撒冷 街市宣告這一切話，說：『當聽從遵行這約的話，
JER|11|7|因為我將你們祖先從 埃及 地領出來的那日，直到今日，都一再切切告誡他們說：當聽從我的話。
JER|11|8|他們卻不聽從，也不側耳而聽，竟隨從自己頑梗的惡心去行。我就使這約中一切詛咒的話臨到他們身上；這約是我吩咐他們遵行的，他們卻不遵行。』」
JER|11|9|耶和華對我說：「在 猶大 人和 耶路撒冷 居民中有同謀背叛的事。
JER|11|10|他們轉去效法他們祖先的惡行，不肯聽我的話，竟隨從別神，事奉它們。 以色列 家和 猶大 家違背了我與他們列祖所立的約。
JER|11|11|所以耶和華如此說：看哪，我必使災禍臨到他們，是他們不能逃脫的。他們向我哀求，我卻不聽。
JER|11|12|那時， 猶大 城鎮的人和 耶路撒冷 的居民要哀求他們燒香所供奉的神明；只是遭難的時候，這些神明一點也不能拯救他們。
JER|11|13|猶大 啊，你神明的數目與你城鎮的數目相等；你所築可恥的壇，就是向 巴力 燒香的壇 ，也與 耶路撒冷 街道的數目相等。
JER|11|14|「所以你不要為這百姓祈禱，也不要為他們呼求禱告，因為他們遭難向我哀求的時候，我必不應允。
JER|11|15|我所親愛的既多設惡謀，還能在我殿中做甚麼呢？你因作惡就喜樂，聖肉要離開你。
JER|11|16|從前耶和華給你起名叫青橄欖樹，又華美又結好果子；如今他用一聲巨響點火在其上，枝子就折斷了。
JER|11|17|「原來栽培你的萬軍之耶和華已經說要降禍給你，是因 以色列 家和 猶大 家行惡。他們向 巴力 燒香，惹我發怒，是自作自受。」
JER|11|18|耶和華指示我，我才知道； 你將他們所做的給我指明。
JER|11|19|我像柔順的羔羊被牽去宰殺， 並不知道他們設計謀害我： 「我們把樹連果子都滅了吧！ 把他從活人之地剪除， 使他的名不再被記得。」
JER|11|20|按公義判斷、察驗人肺腑心腸的萬軍之耶和華啊， 求你使我得見你在他們身上報仇， 因我已將我的案件向你稟明了。
JER|11|21|所以，耶和華論到尋索你命的 亞拿突 人如此說：「他們說：你不要奉耶和華的名說預言，免得你死在我們手中。
JER|11|22|所以萬軍之耶和華如此說：看哪，我必懲罰他們；他們的壯丁必被刀劍殺死，他們的兒女必因饑荒而死，
JER|11|23|他們當中必無任何倖存者；因為在他們受罰之年，我必使災禍臨到 亞拿突 人。」
JER|12|1|耶和華啊，我與你爭辯的時候， 你總是顯為義； 但有一件，我還要與你理論： 惡人的道路為何亨通呢？ 大行詭詐的為何得安逸呢？
JER|12|2|你栽培了他們， 他們也扎了根， 長大，而且結果。 他們的口與你相近， 心卻與你遠離。
JER|12|3|耶和華啊，你認識我，看見我， 你察驗我向你的心如何。 求你將他們拉出來， 如將宰的羊， 為殺戮的日子分別出來。
JER|12|4|這地悲哀， 一切田野的青草枯乾要到幾時呢？ 因其上居民的惡行， 牲畜和飛鳥都滅絕了。 因為他們說：「他看不見 我們的結局 。」
JER|12|5|「你與步行的人同跑， 尚且覺得累， 怎能與馬賽跑呢？ 你在安全之地尚且會跌倒 ， 在 約旦河 邊的叢林要怎麼辦呢？
JER|12|6|因為連你兄弟和你父家都以詭詐待你， 甚至在你後邊大聲喊叫。 雖然他們向你說好話， 你也不要相信他們。」
JER|12|7|我離棄了我的殿宇， 撇棄了我的產業， 將我心裏所親愛的交在她 仇敵手中。
JER|12|8|我的產業向我如林中的獅子， 出聲攻擊我， 因此我恨惡她。
JER|12|9|我的產業向我如斑點的鷙鳥， 有鷙鳥在四圍攻擊她。 你們去聚集田野的百獸， 叫牠們來吞吃吧！
JER|12|10|許多牧人毀壞我的葡萄園， 踐踏我的地產， 使我美好的地產變為荒涼的曠野。
JER|12|11|他們使地荒涼； 地既荒涼，就向我哀哭。 全地荒涼，卻無人在意。
JER|12|12|滅命的來到曠野中一切光禿的高地； 耶和華的刀從地這邊直到地那邊，盡行殺滅， 凡血肉之軀都不得平安。
JER|12|13|他們種的是麥子， 收的卻是荊棘； 辛辛苦苦卻無收穫。 因耶和華的烈怒， 你們必為自己的收成感到羞愧。
JER|12|14|耶和華如此說：「看哪，我要將所有的惡鄰拔出本地，他們曾佔據了我賜給 以色列 百姓所承受的產業；我也要將 猶大 家從他們中間拔出來。
JER|12|15|我拔出他們以後，必回轉過來憐憫他們，使他們歸回，各歸本業，各歸故土。
JER|12|16|他們若殷勤學習我百姓的道，指著我的名起誓：『我指著永生的耶和華起誓』，正如他們從前教我百姓指著 巴力 起誓，他們必在我百姓中得以建立。
JER|12|17|他們若是不聽，我必拔出那國，不但拔出，還要毀滅。這是耶和華說的。」
JER|13|1|耶和華對我如此說：「你去買一條麻布帶子，束在你腰上，不可把它泡在水裏。」
JER|13|2|我就照耶和華的話，買了一條帶子，束在我的腰上。
JER|13|3|耶和華的話第二次臨到我，說：
JER|13|4|「要拿你所買、在你腰上的帶子，起來往 幼發拉底河 去，把腰帶藏在那裏的磐石穴中。」
JER|13|5|我就去，照著耶和華命令我的，把腰帶藏在 幼發拉底河 邊。
JER|13|6|過了多日，耶和華對我說：「你起來往 幼發拉底河 去，把我命令你藏在那裏的腰帶取出來。」
JER|13|7|我就往 幼發拉底河 去，把那腰帶從我所藏的地方挖出來。看哪，腰帶已經破爛，毫無用處了。
JER|13|8|耶和華的話臨到我，說：
JER|13|9|「耶和華如此說：我要照樣敗壞 猶大 的驕傲和 耶路撒冷 的狂傲。
JER|13|10|這惡民不肯聽我的話，按自己頑梗的心而行，隨從別神，事奉敬拜它們；這惡民必像這腰帶，毫無用處。
JER|13|11|腰帶怎樣緊貼人的腰，照樣，我也曾使 以色列 全家和 猶大 全家緊貼著我，歸我為子民，使我得名聲，得頌讚，得榮耀；他們卻不肯聽從。這是耶和華說的。」
JER|13|12|「所以你要對他們說：『耶和華－ 以色列 的上帝如此說：各罈都要裝滿酒。』他們必對你說：『我們豈不知道各罈都要裝滿酒嗎？』
JER|13|13|你就對他們說：『耶和華如此說：看哪，我必使這地所有的居民，就是坐 大衛 寶座的君王、祭司和先知，並 耶路撒冷 所有的居民，都酩酊大醉。
JER|13|14|我要使他們彼此衝突，連父與子也互相衝突；我必不可憐，不顧惜，不憐憫，以致將他們滅絕。這是耶和華說的。』」
JER|13|15|你們當聽，當側耳而聽； 不可驕傲，因為耶和華已經吩咐了。
JER|13|16|當耶和華－你們的上帝 尚未使黑暗來臨， 在昏暗的山上 你們的腳未絆跌以前， 要將榮耀歸給他。 你們盼望光明， 他卻使光明變為死蔭， 成為幽暗。
JER|13|17|你們若不聽這話， 我的心必因你們的驕傲暗自哭泣； 我的眼必痛哭流淚， 因為耶和華的羊群被擄去了。
JER|13|18|你要對君王和太后說： 「你們當自卑，坐下； 因你們的王冠， 就是你們華美的冠冕已經掉落了 。」
JER|13|19|尼革夫 的城鎮都被關閉， 無人打開； 猶大 全被擄掠， 擄掠淨盡。
JER|13|20|你們要舉目觀看從北方來的人。 先前賜給你的羊群， 就是你所引以為榮的羊， 現今在哪裏呢？
JER|13|21|耶和華立你自己所教導的盟友， 立他們為頭來轄制你， 你還有甚麼話可說呢？ 痛苦豈不將你抓住像臨產的婦人嗎？
JER|13|22|你若心裏說：「這一切的事為何臨到我呢？」 是因你罪孽甚多。 你的下襬揭起， 你的腳跟受傷。
JER|13|23|古實 人豈能改變皮膚呢？ 豹豈能改變斑點呢？ 若能，你們這善於行惡的便能行善了。
JER|13|24|我必吹散他們， 如碎秸隨曠野的風飄動。
JER|13|25|這是你所當得的， 是我量給你的報應 ； 因為你忘記了我， 倚靠虛假 。 這是耶和華說的。
JER|13|26|我要揭起你的下襬， 蒙在你臉上， 顯露你的羞恥。
JER|13|27|你在田野的山上行姦淫， 發嘶聲，謀淫亂， 這些可憎之事我都看見了。 耶路撒冷 啊，你有禍了！ 你不肯潔淨 還要等到幾時呢？
JER|14|1|耶和華的話臨到 耶利米 ，論到旱災的事：
JER|14|2|「 猶大 悲哀，城門衰敗； 眾人坐在地上哀慟， 耶路撒冷 的哀聲上達。
JER|14|3|他們的貴族打發童僕去打水； 他們來到水池， 找不到水，就拿著空器皿， 蒙羞慚愧，抱頭而回。
JER|14|4|因為無雨降在地上，土地就乾裂， 農夫為此蒙羞抱頭。
JER|14|5|田野的母鹿因為無草 也撇棄才生的小鹿。
JER|14|6|野驢站在光禿的高地喘氣，好像野狗； 牠們的眼目因無草而失明。」
JER|14|7|耶和華啊，雖然我們的罪孽控告我們， 求你為你名的緣故行動吧！ 我們本是多次背道，得罪了你。
JER|14|8|以色列 所盼望，在患難時作他救主的啊， 你在這地為何像寄居的， 又如旅行的只住一夜呢？
JER|14|9|你為何像受驚嚇的人， 像不能救人的勇士呢？ 耶和華啊，你在我們中間， 我們是稱為你名下的人， 求你不要離開我們。
JER|14|10|耶和華論到這百姓如此說： 「這百姓喜愛遊蕩， 不約束自己的腳步， 所以耶和華不悅納他們。 現今他要記起他們的罪孽， 懲罰他們的罪惡。」
JER|14|11|耶和華又對我說：「不要為這百姓求福。
JER|14|12|他們禁食的時候，我不聽他們的呼求；他們獻燔祭和素祭，我也不悅納。我卻要用刀劍、饑荒、瘟疫滅絕他們。」
JER|14|13|我就說：「唉！主耶和華，看哪，那些先知常對他們說：『你們必不見刀劍，也不遭饑荒；耶和華要在這地方賞賜你們真正的平安。』」
JER|14|14|耶和華對我說：「那些先知託我的名說假預言，我並未差遣他們，沒有吩咐他們，也沒有對他們說話；他們向你們預言的是虛假的異象、占卜、虛無，以及心中的詭詐。
JER|14|15|所以耶和華如此說：『論到託我名說預言的那些先知，我並未差遣他們；他們說這地不會有刀劍、饑荒，其實那些先知自己必被刀劍、饑荒滅絕。
JER|14|16|聽他們說預言的百姓必因饑荒、刀劍被扔在 耶路撒冷 的街道上，無人埋葬。他們連妻子帶兒女，都是如此。我必將他們的惡倒在他們身上。』」
JER|14|17|你要向他們說這些話： 願我眼淚汪汪， 晝夜不息， 因為少女─我百姓 受了重大的打擊， 傷口極其嚴重。
JER|14|18|我若出到田間， 看哪，有被刀殺的； 我若進入城內， 看哪，有因饑荒患病的； 先知和祭司也在各地往來經商， 不知如何是好。
JER|14|19|你全然棄絕 猶大 嗎？ 你的心厭惡 錫安 嗎？ 你為何擊打我們，使我們無法得醫治呢？ 我們指望平安，卻得不著福氣； 指望痊癒，看哪，受了驚惶。
JER|14|20|耶和華啊，我們承認自己的罪惡 和我們祖先的罪孽， 因我們得罪了你。
JER|14|21|求你為你名的緣故， 不厭惡，不輕視你榮耀的寶座。 求你記念， 不要違背你與我們所立的約。
JER|14|22|外邦虛無的神明 中有能降雨的嗎？ 天能自降甘霖嗎？ 耶和華－我們的上帝啊，不是你嗎？ 我們要等候你， 因為這一切都是你所造的。
JER|15|1|耶和華對我說：「雖有 摩西 和 撒母耳 站在我面前，我的心也不顧惜這百姓。你把他們從我眼前趕出，叫他們出去吧！
JER|15|2|他們若問你說：『我們往哪裏去呢？』你就告訴他們，耶和華如此說： 『定為死亡的，必致死亡； 定為刀殺的，必被刀殺； 定為饑荒的，必遭饑荒； 定為擄掠的，必被擄掠。』」
JER|15|3|「我命定四樣災害臨到他們，就是刀劍殺戮、群狗拖拉、空中的飛鳥和地上的走獸吞吃毀滅。這是耶和華說的。
JER|15|4|我必使地上萬國因他們而驚駭，都因 希西家 的兒子 猶大 王 瑪拿西 在 耶路撒冷 所做的事。」
JER|15|5|耶路撒冷 啊，有誰同情你呢？ 有誰為你悲傷呢？ 有誰轉身問你安呢？
JER|15|6|你棄絕了我， 轉身退後； 因此我伸手攻擊你，毀滅你， 我已憐憫到厭煩了。 這是耶和華說的。
JER|15|7|我在境內各關口 用簸箕篩我的百姓， 使他們喪掉兒女， 又毀滅他們， 他們仍不轉離所行的道。
JER|15|8|他們的寡婦在我面前比海沙更多； 我使滅命者在正午來到， 攻擊年輕人的母親， 使痛苦驚嚇忽然臨到她身上。
JER|15|9|生過七個孩子的婦人衰弱； 尚在白晝，太陽忽然落下， 她就抱愧蒙羞。 我必當著敵人的面， 將他們當中的倖存者交給刀劍。 這是耶和華說的。
JER|15|10|我的母親哪，我有禍了！因你生我作全地爭相指控的人。我素來沒有借貸給人，人也沒有借貸給我，人人卻都咒罵我。
JER|15|11|耶和華說：「我必定釋放 你，使你得福氣。災禍苦難來臨時，我必使仇敵央求你。
JER|15|12|人豈能將銅與鐵，就是北方的鐵折斷呢？
JER|15|13|「我必因你在四境之內所犯的一切罪，將你的貨物財寶當掠物，白白地交出來 。
JER|15|14|我要使你的仇敵過去，到你所不認識的地方 ，因為你們要被我怒中所起的火焚燒。」
JER|15|15|耶和華啊，你是知道的； 求你記念我，眷顧我， 向迫害我的人為我報仇； 不要把我取去，因你不輕易發怒， 要知道我為你的緣故受了凌辱。
JER|15|16|耶和華－萬軍之上帝啊， 我得著你的話就把它們吃了， 你的話是我心中的歡喜快樂； 因我是稱為你名下的人。
JER|15|17|我並未坐在享樂人的會中歡樂； 因你的手，我就獨自靜坐， 你使我滿心憤慨。
JER|15|18|我的痛苦為何長久不止呢？ 我的傷痕為何無法可醫，不能痊癒呢？ 難道你以詭詐待我，像流乾的河道嗎？
JER|15|19|所以耶和華如此說：「你若回轉， 我就使你歸回， 站在我面前。 你若能將寶物和無用之物分別出來， 你就可以當作我的口。 他們必歸向你， 你卻不可歸向他們。
JER|15|20|我必使你向這百姓成為堅固的銅牆。 他們必攻擊你，卻不能勝過你； 因我與你同在，要拯救你，搭救你。 這是耶和華說的。
JER|15|21|我必搭救你脫離惡人的手， 救贖你脫離殘暴之人的手。」
JER|16|1|耶和華的話又臨到我，說：
JER|16|2|「你不可在這地方娶妻，為自己生兒育女。
JER|16|3|因為論到在這地方所生的兒女，又論到在這國中生他們的父母，耶和華如此說：
JER|16|4|他們必死於致命的疾病，無人哀哭，不得埋葬，在地上如糞土，因刀劍和饑荒而滅絕；他們的屍首必給空中的飛鳥和地上的走獸作食物。
JER|16|5|「耶和華如此說：不要進入喪家，不要去哀哭，也不要為他們悲傷，因我已使我的平安、慈愛、憐憫離開這百姓。這是耶和華說的。
JER|16|6|他們連大帶小，都必在這地死亡，不得埋葬。人必不為他們哀哭，不為他們割劃自己，也不剃光頭。
JER|16|7|有喪事，人不為他們擘餅 ，也不因死人安慰他們；他們喪父喪母，人也不給他們一杯酒安慰他們。
JER|16|8|你不可進入宴樂的家，與人同坐又吃又喝，
JER|16|9|因為萬軍之耶和華－ 以色列 的上帝如此說：看哪，你們還活著的日子，我必在你們眼前止息這地方歡喜和快樂的聲音、新郎和新娘的聲音。
JER|16|10|「你將這一切的話指示這百姓，他們若問你說：『耶和華為甚麼說，要降這大災禍攻擊我們呢？我們有甚麼罪孽呢？我們向耶和華－我們的上帝犯了甚麼罪呢？』
JER|16|11|你就對他們說：『因為你們祖先離棄了我，隨從別神，事奉敬拜它們，卻離棄我，不遵守我的律法。這是耶和華說的。
JER|16|12|你們行惡比你們祖先更甚，看哪，各人隨從自己頑梗的惡心行事，不聽從我。
JER|16|13|所以我必將你們從這地趕出，直趕到你們和你們祖先素不認識之地。你們在那裏晝夜必事奉別神，因為我必不再向你們施恩。』」
JER|16|14|「看哪，日子將到，人必不再指著那領 以色列 人從 埃及 地上來的永生耶和華起誓。這是耶和華說的。
JER|16|15|人卻要指著那領 以色列 人離開北方之地，離開他們被趕到的各國之永生的耶和華起誓；並且我要領他們歸回我從前賜給他們祖先之地。」
JER|16|16|「看哪，我要差派許多打魚的捕獲他們；以後，我也要派許多打獵的，從各山上、各岡上、各石穴中獵取他們。這是耶和華說的。
JER|16|17|因我的眼目察看他們一切的行為；他們不能在我面前遮掩，他們的罪孽也不能在我眼前隱藏。
JER|16|18|我要先加倍報應他們的罪孽和罪惡，因為他們以可憎之偶像的屍首使我的地玷污，使我的產業充斥可厭之物。」
JER|16|19|耶和華啊，你是我的力量， 是我的保障， 在患難之日是我的避難所。 列國的人必從地極來到你這裏，說： 「我們祖先所承受的， 不過是虛假，是虛空無益之物。
JER|16|20|人豈可為自己製造神明呢？ 其實它們不是神明。」
JER|16|21|「所以，看哪，我要使他們知道，就是這一次使他們知道我的手和我的能力。他們就知道我的名是耶和華了。」
JER|17|1|猶大 的罪是用鐵筆、用金剛石記錄的，銘刻在他們的心版和祭壇角上。
JER|17|2|他們的兒女思念他們在高岡上、青翠樹旁的祭壇和 亞舍拉 。
JER|17|3|我田野的山哪，因你在全境內的丘壇所犯的罪，我必使你的財富和一切的財寶成為掠物。
JER|17|4|因自己所做的 ，你必失去我所賜給你的產業。我也必使你在你所不認識的地服侍你的仇敵；因你們激起了我的怒火，直燒到永遠。
JER|17|5|耶和華如此說： 「倚靠人，以血肉為膀臂， 心中離棄耶和華的， 那人該受詛咒！
JER|17|6|他必像沙漠裏的矮樹， 不見福樂來到； 他要住在曠野乾旱之處， 無人居住的鹽地。
JER|17|7|倚靠耶和華、以耶和華為他所仰賴的， 那人有福了！
JER|17|8|他必像樹栽於水旁， 在河邊扎根， 炎熱來到，毫不察覺 ， 葉子仍必青翠； 在乾旱之年，一無掛慮， 並且結果不止。
JER|17|9|「人心比萬物都詭詐， 壞到極處， 誰能識透呢？
JER|17|10|我－耶和華是鑒察人心，考驗人肺腑的， 要按各人所行的和他做事的結果報應他。」
JER|17|11|那不按正道得財富的， 好像鷓鴣孵不是自己生的； 到了中年，財富必離開他， 終久他必成為愚頑人。
JER|17|12|我們的聖所是榮耀的寶座， 從太初就在高處。
JER|17|13|耶和華－ 以色列 的盼望啊， 凡離棄你的必蒙羞。 離我而去的， 他們必被寫在地裏， 因為他們離棄耶和華，這活水的泉源。
JER|17|14|耶和華啊，求你醫治我，我就痊癒， 拯救我，我便得救； 因你是我所讚美的。
JER|17|15|看哪，他們對我說： 「耶和華的話在哪裏呢？ 讓它應驗吧！」
JER|17|16|至於我，我並沒有逃避作牧人跟隨你 ， 也沒有想望那災殃的日子； 這是你所知道的。 我嘴唇所出的都在你面前。
JER|17|17|不要使我因你驚恐； 災禍來臨時，你是我的避難所。
JER|17|18|願那些迫害我的蒙羞， 卻不要使我蒙羞； 使他們驚惶， 卻不要使我驚惶； 願災禍的日子臨到他們， 以加倍的毀壞毀壞他們。
JER|17|19|耶和華對我如此說：「你去站在 猶大 君王出入的 平民門 ，和 耶路撒冷 的各城門口，
JER|17|20|對他們說：『你們這 猶大 君王、 猶大 眾人和 耶路撒冷 所有的居民，凡從這些城門進入的，都當聽耶和華的話。
JER|17|21|耶和華如此說：你們要謹慎，不可在安息日挑甚麼擔子進入 耶路撒冷 的城門，
JER|17|22|也不可在安息日從家中挑擔子出去。無論何工都不可做，只要以安息日為聖日，正如我所吩咐你們祖先的。』
JER|17|23|他們卻不聽從，也不側耳而聽，竟硬著頸項不聽，不肯領受訓誨。
JER|17|24|「你們若留意聽從我，在安息日不挑甚麼擔子進入這城的各門，只以安息日為聖日，在那日不做任何工作，這是耶和華說的，
JER|17|25|就必有坐 大衛 寶座的君王和領袖，與 猶大 人，並 耶路撒冷 的居民，或坐車，或騎馬，進入這城的各門，而且這城必存到永遠。
JER|17|26|也必有人從 猶大 城鎮和 耶路撒冷 四圍的各處，從 便雅憫 地、 謝非拉 、山區，並 尼革夫 而來，都帶燔祭和祭物，素祭和乳香，並感謝祭，到耶和華的殿去。
JER|17|27|你們若不聽從我，不以安息日為聖日，仍在安息日挑擔子進入 耶路撒冷 的各城門，我必在城門中點火；這火必燒燬 耶路撒冷 的宮殿，不會熄滅。」
JER|18|1|耶和華的話臨到 耶利米 ，說：
JER|18|2|「你起來，下到陶匠的家裏去，在那裏我要使你聽見我的話。」
JER|18|3|我就下到陶匠的家裏去，看哪，他在轉盤上做器皿。
JER|18|4|陶匠用泥做的器皿在他手中做壞了，他就用它另做別的器皿，照他看為好的去做。
JER|18|5|耶和華的話臨到我，說：
JER|18|6|「 以色列 家啊，我待你們豈不能像這陶匠弄泥嗎？ 以色列 家，看哪，泥在陶匠的手中怎樣，你們在我的手中也怎樣。這是耶和華說的。
JER|18|7|我何時論到一邦或一國說，要拔出、拆毀、毀壞；
JER|18|8|我所說的那一邦若回轉離開他們的惡，我就改變心意，不將我想要施行的災禍降與他們。
JER|18|9|我何時論到一邦或一國說，要建立、栽植；
JER|18|10|他們若行我眼中看為惡的事，不聽從我的話，我就改變心意，不將我所說的福氣賜給他們。
JER|18|11|現在你要對 猶大 人和 耶路撒冷 的居民說：『耶和華如此說：看哪，我捏塑災禍降給你們，定意懲罰你們。你們各人當回轉離開所行的惡道，改正你們的所作所為。』
JER|18|12|「他們卻說：『沒有用的，我們要照自己的計謀去行，各人要隨自己頑梗的惡心行事。』」
JER|18|13|「所以，耶和華如此說： 你們且往各國訪問， 有誰聽見這樣的事？ 少女 以色列 行了一件極恐怖的事。
JER|18|14|黎巴嫩 的雪豈能從田野 的磐石上融化呢？ 從遠處 流下的涼水豈能乾涸呢？
JER|18|15|我的百姓竟忘記我， 向那虛無的神明 燒香， 它們使百姓在所行的路上、在古道上絆跌， 去行未修築的斜路，
JER|18|16|他們的地就變為荒涼， 長久被人嘲笑； 凡經過這地的必驚駭搖頭。
JER|18|17|在仇敵面前，我必如東風颳散他們， 遭難的日子，我要以背向他們， 不以臉看他們。」
JER|18|18|他們說：「來吧！讓我們設計謀害 耶利米 ；因為我們有祭司講律法，有智慧人設謀略，有先知說預言，都未曾斷絕。來吧！讓我們用舌頭攻擊他，不要理他一切的話。」
JER|18|19|耶和華啊，求你留心聽我， 且聽那些指控我的人的話。
JER|18|20|人豈可以惡報善呢？ 他們竟挖坑要害我的性命！ 求你記念我站在你面前為他們說好話， 要使你的憤怒轉離他們。
JER|18|21|因此，願他們的兒女忍受饑荒， 願他們死於刀劍之手； 願他們的妻無子，且作寡婦， 願他們的男人被死亡所滅， 他們的壯丁在陣上被刀擊殺。
JER|18|22|你使敵軍忽然臨到他們的時候， 願人聽見哀聲從他們的屋內發出； 因他們挖坑要捉拿我， 暗設羅網要絆我的腳。
JER|18|23|耶和華啊，他們要殺我的那一切計謀， 你都知道。 求你不要赦免他們的罪孽， 也不要從你面前塗去他們的罪惡。 願他們在你面前跌倒， 願你在發怒的時候對付他們。
JER|19|1|耶和華如此說：「你去買陶匠的瓷瓶 ，你和 百姓中的長老、位尊的祭司
JER|19|2|出去到 欣嫩子谷 、 哈珥西 的門口，在那裏宣告我所吩咐你的話，
JER|19|3|說：『 猶大 君王和 耶路撒冷 的居民哪，當聽耶和華的話。萬軍之耶和華－ 以色列 的上帝如此說：看哪，我必使災禍臨到這地方，凡聽見的人都必耳鳴；
JER|19|4|因為他們和他們祖先，並 猶大 君王都離棄我，使這地方與我疏遠 ，在這裏向素不認識的別神燒香，又使這地方遍滿無辜人的血。
JER|19|5|他們建造 巴力 的丘壇，要在火中焚燒自己的兒女，作為燔祭獻給 巴力 。這不是我命令的，不是我吩咐的，我心裏也從來沒有想過。
JER|19|6|因此，看哪，日子將到，這地方不再稱為 陀斐特 和 欣嫩子谷 ，反倒稱為 殺戮谷 。這是耶和華說的。
JER|19|7|我要在這地方使 猶大 和 耶路撒冷 的計謀落空，也必使他們在仇敵面前倒在刀下，倒在尋索其命的人手下。我要把他們的屍首給空中的飛鳥和地上的走獸作食物。
JER|19|8|我必使這城令人驚駭嘲笑；凡路過的，必因這城所遭的災難驚駭嘲笑。
JER|19|9|仇敵和尋索其命的人追逼他們，使他們落在圍困窘迫之中，我必使他們各人吃自己兒女的肉和朋友的肉。』
JER|19|10|「你要在跟你同去的人眼前打碎那瓶，
JER|19|11|對他們說：『萬軍之耶和華如此說：我要打碎這百姓和這城，正如人打碎陶匠的器皿，不能再使其完整。他們要在 陀斐特 埋葬，甚至無處可葬。
JER|19|12|我必向這地方和其中的居民如此行，使這城與 陀斐特 一樣。這是耶和華說的。
JER|19|13|耶路撒冷 的房屋和 猶大 君王的宮殿，就是他們在其上向天上的萬象燒香、向別神獻澆酒祭的宮殿房屋，都必被玷污，和 陀斐特 一樣。』」
JER|19|14|耶利米 從耶和華差他去說預言的 陀斐特 回來，站在耶和華殿的院中對眾百姓說：
JER|19|15|「萬軍之耶和華－ 以色列 的上帝如此說：『看哪，我必使我所說的一切災禍臨到這城和屬它的城鎮，因為他們硬著頸項不聽我的話。』」
JER|20|1|音麥 的兒子 巴施戶珥 祭司作耶和華殿的總管，聽見 耶利米 預言這些事，
JER|20|2|就打 耶利米 先知，用耶和華殿裏 上便雅憫門 內的枷鎖，把他鎖在那裏。
JER|20|3|次日， 巴施戶珥 開枷釋放 耶利米 。於是 耶利米 對他說：「耶和華不叫你的名為 巴施戶珥 ，而叫你 瑪歌珥‧米撒畢 ，
JER|20|4|因耶和華如此說：『看哪，我要使你和你的眾朋友驚嚇；你們要親眼看見他們倒在仇敵的刀下。我必將 猶大 人全都交在 巴比倫 王的手中，他要把他們擄到 巴比倫 去，用刀殺他們。
JER|20|5|我要將這城中一切的貨財和勞碌得來的，並一切的珍寶，以及 猶大 君王所有的寶物，都交在仇敵手中。仇敵要搶奪他們，抓住他們，把他們帶到 巴比倫 去。
JER|20|6|你， 巴施戶珥 ，和所有住在你家中的人都必被擄；你和你的朋友，就是你向他們說假預言的，都要到 巴比倫 去，死在那裏，葬在那裏。』」
JER|20|7|耶和華啊，你欺哄了我， 我也被你欺哄了。 你比我強，並且得勝。 我終日成為笑柄， 人人都戲弄我。
JER|20|8|我每逢講話的時候，就哀嘆， 我喊叫：「有暴力和毀滅！」 因為耶和華的話終日成了我的凌辱和譏刺。
JER|20|9|我若說：「我不再提耶和華， 也不再奉他的名講論」， 我心裏便覺得 似乎有燒著的火悶在我骨中， 我忍受不住，不能自禁。
JER|20|10|我聽見許多的毀謗， 四圍都是驚嚇； 連我知己朋友都看著我跌倒： 「告他吧，我們要告他！ 或者他被引誘， 我們就能勝他， 在他身上報仇。」
JER|20|11|然而，耶和華與我同在， 好像可怕的勇士。 因此，迫害我的都絆跌， 不能得勝； 他們大大蒙羞， 由於行事沒有智慧， 必永遠受那不能忘懷的羞辱。
JER|20|12|考驗義人、察看人肺腑心腸的萬軍之耶和華啊， 求你使我得見你在他們身上報仇， 因我已將我的案件向你稟明了。
JER|20|13|你們要向耶和華唱歌！ 要讚美耶和華！ 因他救了窮人的性命 脫離惡人的手。
JER|20|14|願我出生的那日受詛咒！ 願我母親生我的那天不蒙福！
JER|20|15|報信給我父親說 「你得了兒子」， 使我父親甚歡喜的， 願那人受詛咒。
JER|20|16|願那人像耶和華所傾覆而不憐惜的城鎮； 願他早晨聽見哀聲， 中午聽見吶喊；
JER|20|17|因他沒有在我未出胎就把我殺了， 以致我母親成為我的墳墓， 她卻一直懷著胎 。
JER|20|18|我為何出胎見勞碌愁苦， 在羞愧中度盡我的年日呢？
JER|21|1|耶和華的話臨到 耶利米 。那時， 西底家 王差派 瑪基雅 的兒子 巴施戶珥 和 瑪西雅 的兒子 西番雅 祭司到他那裏去，說：
JER|21|2|「請你為我們求問耶和華，因為 巴比倫 王 尼布甲尼撒 前來攻擊我們；或者耶和華照他一切奇妙的作為待我們，使 巴比倫 王離開我們而去。」
JER|21|3|耶利米 對他們說：「你們當對 西底家 這樣說：
JER|21|4|『耶和華－ 以色列 的上帝如此說：看哪，我要使你們手中的兵器，就是你們與城外圍困你們的 巴比倫 王和 迦勒底 人打仗所用的兵器轉回來，把它們聚集在這城中。
JER|21|5|我要在怒氣、憤怒和大惱怒中，用伸出來的手和大能的膀臂，親自攻擊你們；
JER|21|6|又要擊打這城的居民，他們連人帶牲畜都必遭遇大瘟疫而死亡。
JER|21|7|以後，我要將 猶大 王 西底家 和他的臣僕百姓，就是在城內，從瘟疫、刀劍、饑荒中倖存的人，都交在 巴比倫 王 尼布甲尼撒 手中，交在仇敵和尋索其命的人手中。 巴比倫 王必用刀擊殺他們，不顧惜，不同情，不憐憫。這是耶和華說的。』
JER|21|8|「你要對這百姓說：『耶和華如此說：看哪，我將生命的路和死亡的路擺在你們面前。
JER|21|9|住在這城裏的必遭刀劍、饑荒、瘟疫而死；但出去投降圍困你們之 迦勒底 人的必得存活，保全自己的性命。
JER|21|10|我向這城板臉，降禍不降福；這城必交在 巴比倫 王的手中，他必用火焚燒。這是耶和華說的。』」
JER|21|11|「至於 猶大 王的家，你們當聽耶和華的話。
JER|21|12|大衛 家啊，耶和華如此說： 『每早晨你們要施行公平， 拯救被搶奪的脫離欺壓者的手， 免得我的憤怒因你們的惡行發作， 如火燃起，無人能熄滅。』
JER|21|13|住在山谷和平原磐石上的居民啊， 看哪，我與你們為敵， 因為你們說：『誰能下來攻擊我們？ 誰能進入我們的住處呢？』 這是耶和華說的。
JER|21|14|我必按你們行事的結果懲罰你們， 也必使火在 耶路撒冷 的林中燃起， 將四圍所有的盡行燒滅。 這是耶和華說的。」
JER|22|1|耶和華如此說：「你要下到 猶大 王的宮中，在那裏說這話，
JER|22|2|你要說：『坐 大衛 寶座的 猶大 王啊，你和你的臣僕，並進入這些城門的百姓，都當聽耶和華的話。
JER|22|3|耶和華如此說：你們要施行公平和公義，拯救被搶奪的脫離欺壓者的手，不可虧負寄居的和孤兒寡婦，不可用殘暴對待他們，也不可在這地方流無辜人的血。
JER|22|4|你們若切實遵行這話，就必有坐 大衛 寶座的君王和他的臣僕百姓，或坐車或騎馬，從這王宮的各門進入。
JER|22|5|你們若不聽這些話，我指著自己起誓，這王宮必變為廢墟。這是耶和華說的。』
JER|22|6|耶和華論到 猶大 王的家如此說： 「我看你如 基列 ， 如 黎巴嫩 的山頂； 然而，我必使你變為曠野， 成為無人居住的城鎮。
JER|22|7|我要預備施行毀滅的人， 各人佩帶兵器攻擊你； 他們要砍伐你佳美的香柏樹， 扔在火中。
JER|22|8|「許多國的百姓經過這城，就彼此談論說：『耶和華為何向這大城這樣做呢？』
JER|22|9|必有人回答說：『是因他們離棄了耶和華－他們上帝的約，事奉敬拜別神。』」
JER|22|10|不要為已死的人哀哭， 也不要為他悲傷， 卻要為離家外出的人大大哀哭； 因為他不再回來見自己的出生地。
JER|22|11|因為論到離開這地方的 約西亞 之子 猶大 王 沙龍 ，就是接續他父親 約西亞 作王的，耶和華這樣說：「他必不再回到這裏來，
JER|22|12|卻要死在被擄去的地方，必不得再見這地。」
JER|22|13|禍哉！那以不公義蓋房，以不公平造樓， 白白使鄰舍做工，卻不給工錢的人，
JER|22|14|他說：「我要為自己蓋寬敞的房，蓋高大的樓。」 他為它開窗戶， 以香柏木為牆板， 漆上丹紅色。
JER|22|15|難道你作王就是要蓋香柏木樓房爭勝的嗎？ 你的父親豈不是也吃也喝， 也施行公平和公義嗎？ 那時他得了福樂。
JER|22|16|他為困苦和貧窮的人伸冤， 那時就得了福樂。 認識我不就在此嗎？ 這是耶和華說的。
JER|22|17|你的眼和你的心卻專顧不義之財， 流無辜人的血， 行欺壓和殘暴。
JER|22|18|所以，耶和華論到 約西亞 的兒子 猶大 王 約雅敬 如此說： 人必不為他舉哀： 「哀哉，我的哥哥！ 哀哉，我的姊姊！」 也不為他舉哀： 「哀哉，我的主！ 哀哉，我主的榮華！」
JER|22|19|他被埋葬好像埋驢子一樣， 被拖出去，扔在 耶路撒冷 城門外。
JER|22|20|你要上 黎巴嫩 哀號， 在 巴珊 揚聲， 從 亞巴琳 哀號， 因為你所親愛的都毀滅了。
JER|22|21|你興盛的時候，我對你說話； 你卻說：「我不聽。」 你從年輕時就是這樣， 不肯聽我的話。
JER|22|22|你的牧人要被風吞吃， 你所親愛的必被擄去； 那時你必因你一切的惡行抱愧蒙羞。
JER|22|23|你這住 黎巴嫩 、在香柏樹上搭窩的， 有痛苦臨到你， 如疼痛臨到臨產的婦人， 那時你何等可憐 ！
JER|22|24|耶和華說：「 約雅敬 的兒子 猶大 王 哥尼雅 ，雖是我右手上帶印的戒指，我憑我的永生起誓，我必將你從其上摘下來。
JER|22|25|我要將你交在尋索你命的人和你所懼怕的人手中，就是 巴比倫 王 尼布甲尼撒 和 迦勒底 人手中。
JER|22|26|我也要將你和生你的母親趕到別國，不是你們出生的地方；你們必死在那裏，
JER|22|27|心中雖然很想歸回那地，卻不得歸回。」
JER|22|28|哥尼雅 這人是被輕看、遭毀壞的罐子， 是無人喜愛的器皿嗎？ 他和他的後裔為何被趕到素不認識之地呢？
JER|22|29|地啊，地啊，地啊，當聽耶和華的話！
JER|22|30|耶和華如此說： 「要把這人登記為無子， 是平生不得亨通的人； 因為他後裔中再無一人得亨通， 能坐在 大衛 的寶座上治理 猶大 。」
JER|23|1|耶和華說：「禍哉！那些殘害、趕散我草場之羊的牧人！」
JER|23|2|耶和華－ 以色列 的上帝論到那些牧養他百姓的牧人如此說：「你們趕散我的羊群，並未看顧他們；看哪，我必懲罰你們的惡行。這是耶和華說的。
JER|23|3|我要從我趕他們到的各國召集我羊群中剩餘的，領他們歸回本處；他們必生養眾多。
JER|23|4|我必設立牧人照管他們，牧養他們。他們不再懼怕，不再驚惶，沒有一個失喪的。這是耶和華說的。
JER|23|5|「看哪，日子將到，我要為 大衛 興起公義的苗裔； 他必掌王權，行事有智慧，在地上施行公平和公義。這是耶和華說的。
JER|23|6|在他的日子， 猶大 必得救， 以色列 也安然居住。他的名必稱為『耶和華－我們的義』。
JER|23|7|「看哪，日子將到，人必不再指著那領 以色列 人從 埃及 地上來的永生耶和華起誓。這是耶和華說的。
JER|23|8|人卻要指著那領 以色列 家的後裔離開北方之地、離開我趕他們到的各國的永生耶和華起誓。他們必住在本地。」
JER|23|9|論到那些先知， 我心在我裏面憂傷， 我的骨頭全都發顫； 因耶和華和他的聖言， 我像醉酒的人， 像被酒所勝的人。
JER|23|10|全地滿了犯姦淫的人！ 因妄自賭咒，地就悲哀， 曠野的草場都枯乾了。 他們所行的道是惡的； 他們的權力用得不對。
JER|23|11|連先知帶祭司都是褻瀆的， 就是在我殿中，我也看見他們的惡行。 這是耶和華說的。
JER|23|12|因此，他們的道路必像黑暗中的滑地， 他們必被追趕，仆倒在其上； 因為在他們受罰之年， 我必使災禍臨到他們。 這是耶和華說的。
JER|23|13|我在 撒瑪利亞 的先知中曾見狂妄的事； 他們藉 巴力 說預言， 使我的百姓 以色列 走迷了路。
JER|23|14|我在 耶路撒冷 的先知中曾見恐怖的事； 他們犯姦淫，行虛謊， 又堅固惡人的手， 無人回轉離開自己的惡行。 他們在我面前都像 所多瑪 ， 耶路撒冷 的居民都像 蛾摩拉 。
JER|23|15|因此，萬軍之耶和華論到先知如此說： 「看哪，我必使他們吃茵蔯， 喝苦水； 因為褻瀆的事出於 耶路撒冷 的先知，遍及各地。」
JER|23|16|萬軍之耶和華如此說：「你們不要聽這些先知向你們所說的預言。他們使你們成為虛無，所說的異象是出於自己的心，不是出於耶和華的口。
JER|23|17|他們常對藐視我的人說：『耶和華說：你們必享平安。』 又對一切按自己頑梗之心而行的人說：『災禍必不臨到你們。』」
JER|23|18|有誰站在耶和華的會中 察看並聽見他的話呢？ 有誰留心聽他的話呢？
JER|23|19|看哪！耶和華的暴風 在震怒中發出， 是旋轉的暴風， 必轉到惡人頭上。
JER|23|20|耶和華的怒氣必不轉消， 直到他心中所定的成就了，實現了。 末後的日子，你們要全然明白。
JER|23|21|我並未差遣那些先知， 他們竟自奔跑； 我沒有對他們說話， 他們竟自預言。
JER|23|22|他們若站在我的會中， 必使我的百姓聽我的話， 又使他們回轉離開惡道， 離開他們所行的惡。
JER|23|23|我是靠近你們的上帝，不是遙遠的上帝，不是嗎？ 這是耶和華說的。
JER|23|24|人豈能在隱密處藏身，使我看不見他呢？這是耶和華說的。我豈不遍滿天和地嗎？這是耶和華說的。
JER|23|25|我已聽見那些先知所說的，他們託我的名說假預言：「我做了夢！我做了夢！」
JER|23|26|所言虛假、心存詭詐的先知，他們這樣存心要到幾時呢？
JER|23|27|他們彼此述說所做的夢，想要使我的百姓忘記我的名，正如他們祖先因 巴力 忘記我的名一樣。
JER|23|28|得夢的先知可以述說那夢；領受我話的人可以誠實講我的話。糠秕怎能與麥子比較呢？這是耶和華說的。
JER|23|29|我的話豈不像火，又像能打碎磐石的大錘嗎？這是耶和華說的。
JER|23|30|看哪，那些先知各從鄰舍偷竊我的話，因此我必與他們為敵。這是耶和華說的。
JER|23|31|那些先知用自己的舌頭說是耶和華說的；看哪，我必與他們為敵。這是耶和華說的。
JER|23|32|那些以假夢為預言，又述說這夢，以謊言和魯莽使我百姓走迷了路的，看哪，我必與他們為敵。這是耶和華說的。我並未差遣他們，也沒有吩咐他們。他們對這百姓毫無益處。這是耶和華說的。
JER|23|33|無論是這百姓、是先知、是祭司，問你說：「耶和華有甚麼默示呢？」你就對他們說：「甚麼默示啊？ 我已撇棄你們了。這是耶和華說的。」
JER|23|34|凡說「耶和華的默示」的，無論是先知、是祭司、是百姓，我必懲罰那人和他的家。
JER|23|35|你們各人要對鄰舍、對弟兄如此說：「耶和華回答了甚麼？耶和華說了甚麼呢？」
JER|23|36|你們不可再提「耶和華的默示」，因為各人所說的話必成為自己的重擔 ；你們錯用了永生上帝、萬軍之耶和華－我們上帝的話。
JER|23|37|你們要對先知如此說：「耶和華回答了你甚麼？耶和華說了甚麼呢？」
JER|23|38|你們若說「耶和華的默示」，耶和華就必如此說：「我曾差人到你們那裏去，告訴你們不可說『耶和華的默示』這幾個字，你們卻說『耶和華的默示』；
JER|23|39|所以，看哪，我必忘記你們 ，將你們和我所賜給你們並你們祖先的城都撇棄了；
JER|23|40|又必使永遠的凌辱和長久的羞恥臨到你們，是不能忘記的。」
JER|24|1|巴比倫 王 尼布甲尼撒 將 約雅敬 的兒子 猶大 王 耶哥尼雅 和 猶大 的領袖，並工匠、鐵匠從 耶路撒冷 擄去，帶到 巴比倫 。這事以後，耶和華指給我看，看哪，有兩筐無花果放在耶和華殿前。
JER|24|2|一筐是極好的無花果，像是初熟的；一筐是極壞的無花果，壞得不能吃。
JER|24|3|耶和華對我說：「 耶利米 ，你看見甚麼？」我說：「我看見無花果，好的極好，壞的極壞，壞得不能吃。」
JER|24|4|於是耶和華的話臨到我，說：
JER|24|5|「耶和華－ 以色列 的上帝如此說：『被擄去的 猶大 人，就是我所打發離開這地到 迦勒底 人之地去的，我必看顧他們如這好的無花果，使他們得福樂。
JER|24|6|我要眷顧他們，使他們得福樂，領他們歸回這地。我也要建立他們，必不拆毀；栽植他們，必不拔出。
JER|24|7|我要賜給他們認識我的心，認識我是耶和華。他們要作我的子民，我要作他們的上帝，他們要一心歸向我。』」
JER|24|8|耶和華如此說：「我必將 猶大 王 西底家 和他的眾領袖，以及留在這地 耶路撒冷 剩餘的人，並住在 埃及 地的 猶大 人都交出來，好像那極壞、壞得不能吃的無花果。
JER|24|9|我必使他們在地上萬國中成為恐懼，成為災禍，在我趕逐他們到的各處成為凌辱、笑柄、譏笑、詛咒的對象。
JER|24|10|我必使刀劍、饑荒、瘟疫臨到他們，直到他們從我所賜給他們和他們祖先之地滅絕。」
JER|25|1|約西亞 的兒子 猶大 王 約雅敬 第四年，就是 巴比倫 王 尼布甲尼撒 的元年，耶和華論 猶大 眾百姓的話臨到 耶利米 。
JER|25|2|耶利米 先知就將這些話對 猶大 眾百姓和 耶路撒冷 所有的居民說：
JER|25|3|「從 亞們 的兒子 猶大 王 約西亞 十三年直到今日，在這二十三年中，常有耶和華的話臨到我；我也一再對你們傳講，只是你們不聽從。
JER|25|4|耶和華也曾一再差遣他的僕人眾先知到你們這裏來，只是你們不聽從，也不側耳而聽，
JER|25|5|說：『你們各人當回轉離開惡道和惡行，就可居住耶和華從古時所賜給你們和你們祖先之地，直到永遠。
JER|25|6|不可隨從別神，事奉敬拜它們，以你們手所做的惹我發怒；這樣，我就不會降災禍給你們。
JER|25|7|然而你們不聽從我，竟以手所做的惹我發怒，害了自己。這是耶和華說的。』」
JER|25|8|所以萬軍之耶和華如此說：「因為你們不聽我的話，
JER|25|9|看哪，我必召北方的眾族和我僕人 巴比倫 王 尼布甲尼撒 前來攻擊這地和這地的居民，並四圍所有的國民。我要將他們盡行滅絕，以致他們令人驚駭、嗤笑，並且永久荒涼 。這是耶和華說的。
JER|25|10|我又要止息他們歡喜和快樂的聲音、新郎和新娘的聲音、推磨的聲音和燈的亮光。
JER|25|11|這全地必然荒涼，令人驚駭。這些國家要服事 巴比倫 王七十年。
JER|25|12|七十年滿了以後，我必懲罰 巴比倫 王和那國，並 迦勒底 人之地，因他們的罪孽使那地永遠荒涼。這是耶和華說的。
JER|25|13|我也必使我向那地所說的話，就是所有記在這書上， 耶利米 向這些國家說的預言，都臨到那地。
JER|25|14|因為必有許多國家和大君王使 迦勒底 人作奴僕；我也必照他們的行為，按他們手所做的報應他們。」
JER|25|15|耶和華－ 以色列 的上帝對我如此說：「你從我手中拿這杯憤怒的酒，給我所差遣你去的各國的百姓喝。
JER|25|16|他們喝了就要東倒西歪，並要發狂，因我使刀劍臨到他們中間。」
JER|25|17|我就從耶和華的手中拿了這杯，給耶和華所差遣我去的各國的百姓喝，
JER|25|18|其中有 耶路撒冷 和 猶大 的城鎮，並 耶路撒冷 的君王與領袖；因此這城鎮荒涼，令人驚駭、嗤笑、詛咒，正如今日一樣。
JER|25|19|又有 埃及 王法老和他的臣僕、官長，以及他的眾百姓，
JER|25|20|並混居的各族和 烏斯 地的諸王，與 非利士 人之地的諸王，包括 亞實基倫 、 迦薩 、 以革倫 ，以及 亞實突 剩下的人，
JER|25|21|還有 以東 、 摩押 、 亞捫 人，
JER|25|22|推羅 的諸王、 西頓 的諸王、海的那邊沿海地區的諸王，
JER|25|23|底但 、 提瑪 、 布斯 ，和所有剃鬢髮的人，
JER|25|24|阿拉伯 的諸王、住曠野混居各族的諸王、
JER|25|25|心利 的諸王、 以攔 的諸王、 瑪代 的諸王、
JER|25|26|北方遠近的諸王，以及天下、地面上的萬國也一個一個都喝了，以後 示沙克 王也要喝。
JER|25|27|「你要對他們說：『萬軍之耶和華－ 以色列 的上帝如此說：你們要喝，且要喝醉，要嘔吐，且要跌倒，不再起來，都因我使刀劍臨到你們中間。』
JER|25|28|「他們若不肯從你手中拿這杯來喝，你就要對他們說：『萬軍之耶和華如此說：你們一定要喝！
JER|25|29|看哪，我既從稱為我名下的城起首施行災禍，你們能免去懲罰嗎？你們必不能免，因為我要命刀劍臨到地上所有的居民。這是萬軍之耶和華說的。』
JER|25|30|「所以你要向他們預言這一切的話，對他們說： 『耶和華從高天吼叫， 從聖所發出聲音， 向自己的羊群大聲吼叫； 他要向地上所有的居民吶喊， 像踹葡萄的人一樣。
JER|25|31|必有響聲達到地極， 因為耶和華與列國爭辯。 凡有血肉之軀的，他必審問； 至於惡人，他必交給刀劍。 這是耶和華說的。』
JER|25|32|「萬軍之耶和華如此說： 看哪，必有災禍發出，從這國到那國， 並有大暴風從地極颳起。
JER|25|33|「到那日，從地這邊到地那邊，都有耶和華所殺戮的人。必無人哀哭，不得收殮，不得埋葬，必在地面上成為糞土。
JER|25|34|「牧人哪，你們當哀號，呼喊； 羊群的領導者啊，你們要在灰中翻滾； 因為你們被宰殺、被分散 的日子已經來到。 你們要仆倒，好像珍貴的器皿打碎一樣。
JER|25|35|牧人無路可逃， 羊群的領導者也無法逃脫。
JER|25|36|聽啊，有牧人呼喊， 有羊群領導者哀號的聲音， 因為耶和華摧毀他們的草場。
JER|25|37|因耶和華猛烈的怒氣， 平安的羊圈都被肅清。
JER|25|38|他像獅子離開洞穴， 他們的地因兇猛的怒氣 和他強烈的怒氣，都變為荒涼。」
JER|26|1|約西亞 的兒子 猶大 王 約雅敬 登基時，有這話從耶和華臨到 耶利米 ，說：
JER|26|2|「耶和華如此說：你要站在耶和華殿的院內，對 猶大 所有城鎮的人，就是到耶和華的殿來禮拜的，傳講我所吩咐你的一切話，一字也不可刪減。
JER|26|3|或者他們肯聽從，各人回轉離開惡道，我就改變心意，不將我因他們所行的惡、想要施行的災禍降與他們。
JER|26|4|你要對他們說，耶和華如此說：『你們若不聽從我，不遵行我在你們面前所設立的律法，
JER|26|5|不聽從我一再差遣我僕人眾先知到你們那裏去所說的話，你們果然沒有聽從，
JER|26|6|我就必使這殿如 示羅 ，使這城成為地上萬國所詛咒的。』」
JER|26|7|耶利米 在耶和華殿中所說的這些話，祭司、先知與眾百姓都聽見了。
JER|26|8|耶利米 說完了耶和華吩咐他對眾百姓說的一切話，祭司、先知與眾百姓都來抓住他，說：「你該死！
JER|26|9|你為何假借耶和華的名預言，說這殿必如 示羅 ，這城必荒廢無人居住呢？」於是眾百姓都聚集在耶和華的殿中圍住 耶利米 。
JER|26|10|猶大 的官長們聽見這些事，就從王宮上到耶和華的殿，坐在耶和華殿 新門 的入口。
JER|26|11|祭司、先知對官長和眾百姓說：「這人該死，因為他說預言攻擊這城，正如你們親耳聽見的。」
JER|26|12|耶利米 就對官長和眾百姓說：「耶和華差遣我預言攻擊這殿和這城，傳講你們所聽見的這一切話。
JER|26|13|現在，要改正你們的所作所為，聽從耶和華－你們上帝的話，他就必改變心意，不把所說的災禍降與你們。
JER|26|14|至於我，看哪，我在你們手中，你們眼裏看甚麼是好的，是正確的，就那樣待我吧！
JER|26|15|但你們要確實知道，你們若把我處死，就使流無辜人血的罪歸給你們和這城，以及城裏的居民了；因為耶和華確實差遣我到你們這裏來，將這一切話傳到你們耳中。」
JER|26|16|官長和眾百姓對祭司和先知說：「這人是不該死的，因為他奉耶和華－我們上帝的名向我們說話。」
JER|26|17|國中的長老就有幾個人起來，對聚集的眾百姓說：
JER|26|18|「當 猶大 王 希西家 的日子，有 摩利沙 人 彌迦 對 猶大 眾百姓預言說： 『萬軍之耶和華如此說： 錫安 要被耕種像一塊田地， 耶路撒冷 要變為廢墟， 這殿的山必像叢林的高處。』
JER|26|19|「 猶大 王 希西家 和 猶大 人豈是把他處死呢？ 希西家 豈不是敬畏耶和華，懇求耶和華施恩嗎？耶和華就改變心意，不把所說的災禍降與他們。若處死這人，我們就做了大惡，害死自己了。」
JER|26|20|有一個人，就是 示瑪雅 的兒子 基列‧耶琳 人 烏利亞 ，也奉耶和華的名說預言；他說預言攻擊這城和這地，和 耶利米 所說的完全一樣。
JER|26|21|約雅敬 王和他所有的勇士、官長聽見了 烏利亞 的話，王想要把他處死。 烏利亞 聽見就懼怕，逃往 埃及 去了。
JER|26|22|約雅敬 王差 亞革波 的兒子 以利拿單 ，帶領幾個人前往 埃及 。
JER|26|23|他們將 烏利亞 從 埃及 帶出來，解送到 約雅敬 王那裏；王用刀殺了他，把他的屍首拋在平民的墳地中。
JER|26|24|然而， 沙番 的兒子 亞希甘 保護 耶利米 ，不將他交在百姓手中，以免他們把他處死。
JER|27|1|約西亞 的兒子 猶大 王 約雅敬 登基時，有這話從耶和華臨到 耶利米 ，說：
JER|27|2|「耶和華對我如此說：你要為自己做皮帶和木軛，套在你的頸項上，
JER|27|3|然後託那些來到 耶路撒冷 ，到 猶大 王 西底家 那裏的使節，把皮帶和木軛送到 以東 王、 摩押 王、 亞捫 王、 推羅 王、 西頓 王那裏，
JER|27|4|且囑咐他們轉達他們的主人。萬軍之耶和華－ 以色列 的上帝如此說，你們要對你們的主人這樣說：
JER|27|5|我用大能和伸出來的膀臂創造大地和地上的人民、牲畜。我看給誰合適，就把地給誰。
JER|27|6|現在我將全地都交在我僕人 巴比倫 王 尼布甲尼撒 手中，也把野地的走獸給他使用。
JER|27|7|列國都要服事他和他的子孫，直到他本國遭報的日期來到；那時，許多國家和大君王要使他作奴隸。
JER|27|8|「無論哪一邦、哪一國，不肯服事 巴比倫 王 尼布甲尼撒 ，不把頸項放在他的軛下，我必用刀劍、饑荒、瘟疫懲罰那邦，直到我藉 巴比倫 王的手毀滅他們。這是耶和華說的。
JER|27|9|至於你們，不可聽從你們的先知和占卜的、做夢的 、觀星象的，以及行邪術的；他們對你們說：『你們必不致服事 巴比倫 王。』
JER|27|10|他們向你們傳的是假預言，要叫你們遠離本地，以致我將你們趕出去，使你們滅亡。
JER|27|11|但哪一邦肯把頸項放在 巴比倫 王的軛下服事他，我必使那邦仍在本地存留，在那裏耕種居住。這是耶和華說的。」
JER|27|12|我就照這一切話對猶大王 西底家 說：「你們要把頸項放在 巴比倫 王的軛下，服事他和他的百姓，就得存活。
JER|27|13|你和你的百姓何必因刀劍、饑荒、瘟疫而死亡，像耶和華所論不肯服事 巴比倫 王的國家呢？
JER|27|14|不可聽那些先知對你們所說的話，他們說：『你們必不致服事 巴比倫 王』，其實他們向你們傳的是假預言。
JER|27|15|耶和華說：『我並未差遣他們，他們卻託我的名傳假預言，使我將你們和向你們說預言的那些先知趕出去，一同滅亡。』」
JER|27|16|我又對祭司和這眾百姓說：「耶和華如此說：你們不可聽那先知對你們所說的預言，他們說：『看哪，耶和華殿中的器皿快要從 巴比倫 帶回來』；其實他們向你們傳的是假預言。
JER|27|17|不可聽從他們，只管服事 巴比倫 王，就得存活。何必使這城變為廢墟呢？
JER|27|18|他們若真是先知，有耶和華的話臨到他們，讓他們祈求萬軍之耶和華，使耶和華殿中和 猶大 王宮內，並 耶路撒冷 剩下的器皿，不致被帶到 巴比倫 去。
JER|27|19|萬軍之耶和華這樣論柱子、銅海、盆座，並留在這城裏剩下的器皿，
JER|27|20|就是 巴比倫 王 尼布甲尼撒 擄掠 約雅敬 的兒子 猶大 王 耶哥尼雅 ，並 猶大 、 耶路撒冷 所有貴族時，沒有從 耶路撒冷 掠去 巴比倫 的器皿。
JER|27|21|論到那在耶和華殿中和 猶大 王宮內，並 耶路撒冷 剩下的器皿，萬軍之耶和華－ 以色列 的上帝如此說：
JER|27|22|它們必被帶到 巴比倫 ，存放在那裏，直到我眷顧 以色列 人，將這些器皿帶回歸還此地的日子。這是耶和華說的。」
JER|28|1|當年，就是 猶大 王 西底家 登基第四年五月， 押朔 的兒子 基遍 人 哈拿尼雅 先知，在耶和華的殿中當著祭司和眾百姓的面對我說：
JER|28|2|「萬軍之耶和華－ 以色列 的上帝如此說：我已經折斷 巴比倫 王的軛。
JER|28|3|二年之內，我要將 巴比倫 王 尼布甲尼撒 從這地擄掠到 巴比倫 的器皿，就是耶和華殿中的一切器皿，都帶回此地。
JER|28|4|我又要將 約雅敬 的兒子 猶大 王 耶哥尼雅 和被擄到 巴比倫 所有的 猶大 人帶回此地，因為我要折斷 巴比倫 王的軛。這是耶和華說的。」
JER|28|5|耶利米 先知當著祭司和站在耶和華殿裏眾百姓的面，對 哈拿尼雅 先知說：
JER|28|6|「阿們！願耶和華如此行，願耶和華實現你所預言的話，將耶和華殿中的器皿和所有被擄去的人從 巴比倫 帶回此地。
JER|28|7|然而我在你和眾百姓耳中所要說的話，你應當聽。
JER|28|8|從古以來，在你我以前的眾先知，向多國和大邦說預言，論到戰爭、災禍 、瘟疫的事。
JER|28|9|至於那預言平安的先知，到先知的話應驗的時候，人就知道他真是耶和華所差來的。」
JER|28|10|哈拿尼雅 先知就取下 耶利米 先知頸項上的軛，把它折斷。
JER|28|11|哈拿尼雅 又當著眾百姓的面說：「耶和華如此說：二年之內我必照樣從列國的頸項上折斷 巴比倫 王 尼布甲尼撒 的軛。」 耶利米 先知就離開了。
JER|28|12|哈拿尼雅 先知折斷 耶利米 先知頸項上的軛以後，耶和華的話臨到 耶利米 ，說：
JER|28|13|「你去告訴 哈拿尼雅 說，耶和華如此說：你折斷木軛，卻換來鐵軛！
JER|28|14|萬軍之耶和華－ 以色列 的上帝如此說：我已將鐵軛加在這些國的頸項上，使他們服事 巴比倫 王 尼布甲尼撒 。他們總要服事他，我也把野地的走獸給了他。」
JER|28|15|於是 耶利米 先知對 哈拿尼雅 先知說：「 哈拿尼雅 啊，你應當聽！耶和華並沒有差遣你，你竟使這百姓倚靠謊言。
JER|28|16|所以耶和華如此說：看哪，我要把你從地面上除掉，你今年必死，因為你向耶和華說了叛逆的話。」
JER|28|17|這樣， 哈拿尼雅 先知當年七月間就死了。
JER|29|1|耶利米 先知從 耶路撒冷 送信給被擄倖存的長老，以及祭司、先知，和 尼布甲尼撒 從 耶路撒冷 擄到 巴比倫 去的眾百姓。
JER|29|2|這是在 耶哥尼雅 王和太后、官員，並 猶大 和 耶路撒冷 的領袖，以及工匠、鐵匠都離開 耶路撒冷 之後。
JER|29|3|他藉 沙番 的兒子 以利亞薩 和 希勒家 的兒子 基瑪利 的手送去；他們二人是 猶大 王 西底家 差往 巴比倫 去見 巴比倫 王 尼布甲尼撒 的。
JER|29|4|信上說：「萬軍之耶和華－ 以色列 的上帝對所有被擄的，就是我使他們從 耶路撒冷 被擄到 巴比倫 去的人如此說：
JER|29|5|你們要建造房屋，住在其中；要開墾田園，吃園中所出產的；
JER|29|6|要娶妻生兒養女，為你們的兒子娶妻，使你們的女兒嫁人，生兒養女。你們要在那裏生養眾多，不可減少。
JER|29|7|我使你們被擄到的那城，你們要為那城求平安，為那城向耶和華祈求，因為那城得平安，你們也隨著得平安。
JER|29|8|萬軍之耶和華－ 以色列 的上帝如此說：不要被你們中間的先知和占卜的所誘惑，也不要聽信你們 所做的夢，
JER|29|9|因為他們託我的名對你們說假預言，我並未差遣他們。這是耶和華說的。
JER|29|10|「耶和華如此說：為 巴比倫 所定的七十年滿了以後，我要眷顧你們，向你們實現我的恩言，使你們歸回此地。
JER|29|11|我知道我向你們所懷的意念是賜平安的意念，不是降災禍的意念，要叫你們末後有指望。這是耶和華說的。
JER|29|12|你們呼求我，向我禱告，我就應允你們。
JER|29|13|你們尋求我，若專心尋求我，就必尋見。
JER|29|14|我必被你們尋見，也必使你們被擄的人歸回。這是耶和華說的。我必將你們從各國和我趕你們到的各處召集過來，又將你們帶回我使你們被擄離開的地方。這是耶和華說的。
JER|29|15|「你們說：『耶和華已在 巴比倫 為我們興起先知。』
JER|29|16|所以耶和華如此論坐 大衛 寶座的君王和住在這城裏所有的百姓，就是未曾與你們一同被擄的弟兄，
JER|29|17|萬軍之耶和華如此說：『看哪，我必使刀劍、饑荒、瘟疫臨到他們，使他們像極壞的無花果，壞得不能吃。
JER|29|18|我必用刀劍、饑荒、瘟疫追趕他們，使地上萬國因他們而驚駭；在我趕他們到的各國，令人詛咒、驚駭、嗤笑、羞辱。
JER|29|19|這是因為他們不聽從我先前一再差遣我僕人眾先知說的話。這是耶和華說的。你們 也一樣不聽。這是耶和華說的。』
JER|29|20|所以你們所有被擄去的，就是我從 耶路撒冷 放逐到 巴比倫 去的，當聽耶和華的話。
JER|29|21|萬軍之耶和華－ 以色列 的上帝論 哥賴雅 的兒子 亞哈 和 瑪西雅 的兒子 西底家 如此說：『他們託我的名向你們說假預言，看哪，我必把他們交在 巴比倫 王 尼布甲尼撒 的手中，他要在你們眼前殺害他們。
JER|29|22|在 巴比倫 所有被擄的 猶大 人必藉這二人賭咒說：願耶和華使你像 巴比倫 王在火中焚燒的 西底家 和 亞哈 一樣。
JER|29|23|這二人在 以色列 中做了醜事，與鄰舍的妻行淫，又假託我的名說我未曾吩咐他們的話。我知道這一切，也作見證。這是耶和華說的。』」
JER|29|24|「你要對 尼希蘭 人 示瑪雅 說：
JER|29|25|萬軍之耶和華－ 以色列 的上帝如此說：你曾用自己的名送信給 耶路撒冷 的眾百姓和 瑪西雅 的兒子 西番雅 祭司，並眾祭司，說：
JER|29|26|『耶和華已經立你 西番雅 為祭司，代替 耶何耶大 祭司，使耶和華的殿中有總管，好把所有狂妄自稱先知的人用枷枷住，用鎖鎖住。
JER|29|27|現在 亞拿突 人 耶利米 向你們自稱先知，你為甚麼不責備他呢？
JER|29|28|他送信給我們在 巴比倫 的人說：被擄的事必長久，你們要建造房屋，住在其中；要開墾田園，吃園中所出產的。』」
JER|29|29|西番雅 祭司就把這信念給 耶利米 先知聽。
JER|29|30|於是耶和華的話臨到 耶利米 ，說：
JER|29|31|「你當送信給所有被擄的人，說：『耶和華論到 尼希蘭 人 示瑪雅 說：因為 示瑪雅 向你們說預言，使你們倚靠謊言，而我並沒有差遣他，
JER|29|32|所以耶和華如此說：看哪，我必懲罰 尼希蘭 人 示瑪雅 和他的後裔，他必無一人存留住在這民中，也看不見我所要賞賜給我百姓的福樂，因為他向耶和華說了叛逆的話。這是耶和華說的。』」
JER|30|1|耶和華的話臨到 耶利米 ，說：
JER|30|2|「耶和華－ 以色列 的上帝如此說：你要將我對你說過的一切話都寫在書上。
JER|30|3|看哪，日子將到，我要使我的百姓 以色列 和 猶大 被擄的人歸回。這是耶和華說的。耶和華說：我要使他們回到我所賜給他們祖先之地，他們就得這地為業。」
JER|30|4|以下是耶和華論到 以色列 和 猶大 所說的話：
JER|30|5|耶和華如此說： 「我們聽見顫抖的聲音， 令人懼怕，沒有平安。
JER|30|6|你們且訪查看看， 男人會生孩子嗎？ 我怎麼看見人人都用手撐腰， 像臨產的婦人， 臉都發白了呢？
JER|30|7|哀哉！ 那日為大， 無日可比； 這是 雅各 遭難的時刻， 但他必從患難中得拯救。」
JER|30|8|萬軍之耶和華說：「到那日，我必折斷你頸項上仇敵的軛，拉斷你的皮帶。陌生人必不再使他作奴隸。
JER|30|9|他們卻要事奉耶和華－他們的上帝，事奉我為他們所興起的 大衛 王。」
JER|30|10|我的僕人 雅各 啊，不要懼怕； 以色列 啊，不要驚惶； 因我從遠方拯救你， 從被擄之地拯救你的後裔； 雅各 必回來得享平靜安逸， 無人能使他害怕。 這是耶和華說的。
JER|30|11|因我與你同在，要拯救你， 也要將那些國滅絕淨盡， 就是我趕你去的那些國； 卻不將你滅絕淨盡， 倒要從寬懲治你， 但絕不能不罰你。 這是耶和華說的。
JER|30|12|耶和華如此說： 「你的損傷無法醫治， 你的傷痕極其重大。
JER|30|13|無人為你的傷痛辯護， 也沒有可醫治你的良藥。
JER|30|14|你所親愛的都忘記你， 不來探望你。 我因你罪孽甚大，罪惡眾多， 曾藉仇敵加的傷害傷害你， 藉殘忍者懲治你。
JER|30|15|你為何因所受的損傷哀號呢？ 你的痛苦無法醫治。 我因你罪孽甚大，罪惡眾多， 曾將這些加在你身上。
JER|30|16|因此，凡吞吃你的必被吞吃， 你的敵人個個都被擄去； 擄掠你的必成為擄物， 我使搶奪你的成為掠物。
JER|30|17|我必使你痊癒， 醫好你的傷痕， 都因人稱你為被趕散的， 這是 錫安 ，是無人來探望的！ 這是耶和華說的。」
JER|30|18|耶和華如此說： 「看哪，我必使 雅各 被擄去的帳棚歸回， 也必顧惜他的住處。 城必建造在原有的廢墟上， 宮殿也必照樣有人居住。
JER|30|19|必有感謝和歡樂的聲音從其中發出， 我使他們增多，不致減少； 使他們尊榮，不致卑微。
JER|30|20|他們的兒女必如往昔； 他們的會眾堅立在我面前； 凡欺壓他們的，我必懲罰。
JER|30|21|他們的君王是他們自己的人， 掌權的必出自他們。 我要使他接近我， 他也要親近我； 不然，誰敢放膽親近我呢？ 這是耶和華說的。
JER|30|22|你們要作我的子民， 我要作你們的上帝。」
JER|30|23|看哪，耶和華的憤怒 如暴風已經發出； 是掃滅的暴風， 必轉到惡人的頭上。
JER|30|24|耶和華的烈怒必不轉消， 直到他心中所定的成就了，實現了； 末後的日子你們就會明白。
JER|31|1|耶和華說：「那時，我必作 以色列 各家的上帝，他們必作我的子民。」
JER|31|2|耶和華如此說： 「從刀劍生還的百姓 在曠野蒙恩； 以色列 尋找安歇之處。」
JER|31|3|耶和華從遠方向我顯現： 「我以永遠的愛愛你， 因此，我以慈愛吸引你。」
JER|31|4|少女 以色列 啊， 我要再建立你，你就得以建立； 你必再拿起手鼓， 隨著歡樂的舞者而出。
JER|31|5|你必在 撒瑪利亞 的山上栽葡萄園， 栽種的人栽種，而且享用。
JER|31|6|日子將到，守望的人必在 以法蓮 山上呼叫： 「起來吧！我們要上 錫安 ， 到耶和華－我們的上帝那裏去。」
JER|31|7|耶和華如此說： 「你們當為 雅各 歡樂歌唱， 為萬國中為首的歡呼。 當傳揚，頌讚說： 『耶和華啊， 求你拯救你的百姓 ， 拯救 以色列 的餘民。』
JER|31|8|看哪，我必將他們從北方之地領來， 從地極召集而來； 同他們來的有盲人、瘸子、孕婦、產婦； 他們必成群結隊回到這裏。
JER|31|9|他們要哭泣而來。 我要照他們懇求的引導他們， 使他們在河水旁行走正直的路， 他們在其上必不致絆跌； 因為我是 以色列 的父， 以法蓮 是我的長子。
JER|31|10|列國啊，要聽耶和華的話， 要在遠方的海島傳揚，說： 「趕散 以色列 的必召集他， 看守他，如牧人看守羊群。」
JER|31|11|因為耶和華救贖了 雅各 ， 救贖他脫離比他更強之人的手。
JER|31|12|他們來到 錫安 的高處歌唱， 因耶和華的宏恩而喜樂洋溢， 就是五穀、新酒和新的油， 並羔羊和牛犢。 他們必像有水澆灌的園子， 一點也不再有愁煩。
JER|31|13|那時，少女必歡樂跳舞； 年輕的、年老的，都一同歡樂； 因為我要使他們的悲哀變為歡喜， 並要安慰他們，使他們的愁煩轉為喜樂。
JER|31|14|我必以肥油使祭司的心滿足， 我的百姓也要因我的恩惠知足。 這是耶和華說的。
JER|31|15|耶和華如此說： 「在 拉瑪 聽見號咷痛哭的聲音， 是 拉結 哭她兒女，不肯因她兒女受安慰， 因為他們都不在了。」
JER|31|16|耶和華如此說： 「不要出聲哀哭， 你的眼目也不要流淚； 因你的辛勞必有報償， 他們必從仇敵之地歸回。 這是耶和華說的。
JER|31|17|你末後必有指望， 你的兒女必回到自己的疆土。 這是耶和華說的。
JER|31|18|我聽見 以法蓮 為自己悲嘆說： 『你管教我，我便受管教， 我如未馴服的牛犢。 求你使我回轉，我便回轉， 因為你是耶和華－我的上帝。
JER|31|19|我背離以後就懊悔， 受教以後就捶胸 ； 我因擔當年輕時的凌辱就抱愧蒙羞。』
JER|31|20|以法蓮 是我的愛子嗎？ 是我喜歡的孩子嗎？ 我每逢責備他，仍深顧念他。 因此，我的心腸牽掛著他， 我必要憐憫他。 這是耶和華說的。
JER|31|21|少女 以色列 啊， 當為自己設立路標， 為自己豎起指路牌。 要留心向著大道， 就是你曾走過的路； 你當回轉，回到你自己的城鎮。
JER|31|22|背道的女子啊， 你翻來覆去要到幾時呢？ 耶和華在地上造了一件新事， 就是女子護衛男子。」
JER|31|23|萬軍之耶和華－ 以色列 的上帝如此說：「我使被擄之人歸回的時候，他們在 猶大 地和其中的城鎮必再這樣說： 公義的居所啊，聖山哪， 願耶和華賜福給你。
JER|31|24|猶大 和 猶大 城鎮的人，耕地的和帶著群畜遊牧的人，都要一同住在其中。
JER|31|25|疲乏的人，我使他振作；愁煩的人，我使他滿足。」
JER|31|26|於是我醒了，我看到我睡得香甜。
JER|31|27|「看哪，日子將到，我要使人的後代和牲畜的種，在 以色列 家和 猶大 家繁衍。這是耶和華說的。
JER|31|28|我先前怎樣看守他們，為要拔出、拆毀、毀壞、傾覆、苦害，也必照樣看守他們，為要建立、栽植。這是耶和華說的。
JER|31|29|當那些日子，人不再說： 『父親吃了酸葡萄， 兒子牙齒就酸倒。』
JER|31|30|但各人要因自己的罪死亡；凡吃酸葡萄的，自己的牙必酸倒。
JER|31|31|「看哪，日子將到，我要與 以色列 家和 猶大 家另立新的約。這是耶和華說的。
JER|31|32|這約不像我拉著他們祖宗的手，領他們出 埃及 地的時候與他們所立的約。我雖作他們的丈夫，他們卻背了我的約。這是耶和華說的。
JER|31|33|那些日子以後，我與 以色列 家所立的約是這樣：我要將我的律法放在他們裏面，寫在他們心上。我要作他們的上帝，他們要作我的子民。這是耶和華說的。
JER|31|34|他們各人不再教導自己的鄰舍和弟兄說：『你該認識耶和華』，因為他們從最小的到最大的都必認識我。我要赦免他們的罪孽，不再記得他們的罪惡。這是耶和華說的。」
JER|31|35|耶和華使太陽白晝發光， 按定例使月亮和星辰照耀黑夜， 又攪動大海，使海中波浪澎湃， 萬軍之耶和華是他的名， 他如此說：
JER|31|36|「這些定例若能在我面前廢掉， 以色列 的後裔才會在我面前斷絕， 永遠不再成國。 這是耶和華說的。」
JER|31|37|耶和華如此說： 「若有人能測量上面的天， 探索下面地的根基， 我才會因 以色列 後裔所做的一切棄絕他們。 這是耶和華說的。」
JER|31|38|看哪，日子將到，這城必為耶和華而造，從 哈楠業樓 直到 角門 。這是耶和華說的。
JER|31|39|丈量的繩子要往外拉出，直到 迦立山 ，又轉到 歌亞 ；
JER|31|40|拋屍的全谷和倒灰之處，並一切田地，直到 汲淪溪 ，又到東邊 馬門 的角落，都要歸耶和華為聖；不再拔出，不再傾覆，直到永遠。
JER|32|1|猶大 王 西底家 第十年，就是 尼布甲尼撒 十八年，耶和華的話臨到 耶利米 。
JER|32|2|那時 巴比倫 王的軍隊圍困 耶路撒冷 ， 耶利米 先知被囚在 猶大 王宮中護衛兵的院內；
JER|32|3|因為 猶大 王 西底家 囚禁他，說：「你為甚麼預言耶和華如此說：『看哪，我要把這城交在 巴比倫 王的手中，他必攻下這城。
JER|32|4|猶大 王 西底家 必不能逃脫 迦勒底 人的手，定要交在 巴比倫 王手中，他要親眼看到 巴比倫 王，親口跟他說話。
JER|32|5|巴比倫 王要將 西底家 帶到 巴比倫 ； 西底家 必住在那裏，直到我懲罰 他的時候。你們雖與 迦勒底 人爭戰，卻不順利。這是耶和華說的。』」
JER|32|6|耶利米 說：「耶和華的話臨到我，說：
JER|32|7|『看哪，你叔父 沙龍 的兒子 哈拿篾 必到你這裏來，說：請你買我在 亞拿突 的那塊地，因為你有代贖的責任。』
JER|32|8|我叔父的兒子 哈拿篾 果然照耶和華的話來到護衛兵的院內，對我說：『請你買我在 便雅憫 境內、 亞拿突 的那塊地；因為它應該由你來承受，而且你也有代贖的責任。請你買下它吧！』我就知道這確是耶和華的話。
JER|32|9|「我便向我叔父的兒子 哈拿篾 買了 亞拿突 的那塊地，秤了十七舍客勒銀子給他。
JER|32|10|我在契上簽字，將契封緘，又請證人來，用天平把銀子秤給他。
JER|32|11|我又將按照法定條例所立的買契，就是封緘的那一張和敞開的那一張，
JER|32|12|在我叔父的兒子 哈拿篾 和簽字作證的人，並坐在護衛兵院內所有 猶大 人眼前，交給 瑪西雅 的孫子 尼利亞 的兒子 巴錄 。
JER|32|13|我在眾人眼前囑咐 巴錄 說：
JER|32|14|『萬軍之耶和華－ 以色列 的上帝如此說：你拿著這文件，就是封緘的和敞開的買契，把它們放在瓦器裏，以便長久保存。
JER|32|15|因為萬軍之耶和華－ 以色列 的上帝如此說：將來在這地必有人再購置房屋、田地和葡萄園。』」
JER|32|16|「我將買契交給 尼利亞 的兒子 巴錄 以後，就向耶和華禱告說：
JER|32|17|『唉！主耶和華，看哪，你曾用大能和伸出來的膀臂創造天和地，在你沒有難成的事。
JER|32|18|你施慈愛給千萬人，又將祖先的罪孽報應在他後世子孫身上。至大全能的上帝啊，萬軍之耶和華是你的名，
JER|32|19|你謀事有大略，行事有大能，注目觀看世人一切的舉動，為要照各人所做的和他做事的結果報應他。
JER|32|20|你在 埃及 地顯神蹟奇事，直到今日在 以色列 和世人中間也是如此，建立了自己的名聲，正如今日一樣。
JER|32|21|你用神蹟奇事、大能的手、伸出來的膀臂和大可畏的事，領你的百姓 以色列 出了 埃及 ，
JER|32|22|把這地賞賜給他們，就是你向他們列祖起誓應許要賜給他們的流奶與蜜之地。
JER|32|23|他們進入並取得這地，卻不聽從你的話，也不遵行你的律法。你吩咐他們所當行的，他們都不去行，因此你使這一切的災禍臨到他們。
JER|32|24|看哪，敵人已經來到，用土堆攻取這城；這城也因刀劍、饑荒、瘟疫被交在攻城的 迦勒底 人手中。你所說的話都應驗了，看哪，你也看見了。
JER|32|25|主耶和華啊，你卻對我說，要用銀子為自己買那塊地，又請人作證；其實這城已交在 迦勒底 人的手中了。』」
JER|32|26|耶和華的話臨到 耶利米 ，說：
JER|32|27|「看哪，我是耶和華，是凡有血肉之軀者的上帝，在我豈有難成的事嗎？
JER|32|28|耶和華如此說：看哪，我必將這城交給 迦勒底 人的手和 巴比倫 王 尼布甲尼撒 的手，他必攻取這城。
JER|32|29|攻城的 迦勒底 人必來放火焚燒這城和城裏的房屋；人曾在這房頂上向 巴力 燒香，向別神獻澆酒祭，惹我發怒。
JER|32|30|以色列 人和 猶大 人從年輕時，就專做我眼中看為惡的事。 以色列 人盡以手所做的惹我發怒。這是耶和華說的。
JER|32|31|這城自從建造的那日直到今日，常惹我的怒氣和憤怒，以致我將這城從我面前除掉；
JER|32|32|這是因 以色列 人和 猶大 人一切的邪惡，就是他們和他們的君王、官長、祭司、先知，並 猶大 人，以及 耶路撒冷 居民所做的，惹我發怒。
JER|32|33|他們以背向我，不以面向我；我雖然一再教導他們，他們卻不聽從，不領受訓誨，
JER|32|34|竟把可憎之偶像設立在稱為我名下的殿中，玷污了這殿。
JER|32|35|他們在 欣嫩子谷 建造 巴力 的丘壇，把自己的兒女經火獻給 摩洛 ；他們行這可憎的事，使 猶大 陷在罪裏，這並不是我吩咐的，我心裏也從來沒有想過。」
JER|32|36|現在論到這城，就是你們所說，已經因刀劍、饑荒、瘟疫被交在 巴比倫 王手中的，耶和華－ 以色列 的上帝如此說：
JER|32|37|「看哪，我曾在怒氣、憤怒和大惱怒中，將 以色列 人趕到各國；我必從那裏將他們召集出來，領他們回到此地，使他們安然居住。
JER|32|38|他們要作我的子民，我要作他們的上帝。
JER|32|39|我要使他們彼此同心同道，好叫他們永遠敬畏我，使他們和他們後世的子孫得享福樂。
JER|32|40|我要跟他們立永遠的約，要施恩給他們，絕不轉離；又要把敬畏我的心放在他們心裏，不離棄我。
JER|32|41|我必歡喜施恩給他們，盡心盡意、真誠地將他們栽於此地。
JER|32|42|「因為耶和華如此說：我怎樣使這一切大災禍臨到這百姓，也要照樣使我所應許他們的一切福樂都臨到他們。
JER|32|43|你們所說荒涼、無人、無牲畜，已交給 迦勒底 人手的這地，必有人購置田地。
JER|32|44|在 便雅憫 地、 耶路撒冷 四圍的各處、 猶大 的城鎮、山區的城鎮、 謝非拉 的城鎮，並 尼革夫 的城鎮，人必用銀子買田地，在契上簽字，將契封緘，找人作證，因為我必使被擄的人歸回。這是耶和華說的。」
JER|33|1|耶利米 還囚在護衛兵的院內，耶和華的話第二次臨到他，說：
JER|33|2|「成事的耶和華，塑造它為要建立它的耶和華，名為耶和華的那位如此說：
JER|33|3|『你求告我，我就應允你，並將你所不知道、又大又隱密的事指示你。
JER|33|4|論到這城中的房屋和 猶大 君王的宮殿，就是拆毀來擋圍城工事和刀劍的，耶和華－ 以色列 的上帝如此說：
JER|33|5|他們與 迦勒底 人爭戰，用我在怒氣和憤怒中所殺之人的屍首塞滿這房屋；我因他們一切的惡，轉臉不顧這城。
JER|33|6|看哪，我要使這城得以痊癒安舒，我要醫治他們，將豐盛的平安與信實顯明給他們。
JER|33|7|我也要使 猶大 被擄的和 以色列 被擄的人歸回，並要建立他們，如起初一樣。
JER|33|8|我要洗淨他們干犯我的一切罪，赦免他們干犯我、違背我的一切罪。
JER|33|9|這城在地上萬國面前要因我的緣故，以喜樂得名，得頌讚，得榮耀，因為他們聽見我所賞賜的一切福樂。他們因我向這城所施的一切福樂平安，就懼怕戰兢。」
JER|33|10|耶和華如此說：「你們論這地方，說是荒廢、無人、無牲畜之地，但在這荒涼、無人、無居民、無牲畜的 猶大 城鎮和 耶路撒冷 街上，必再聽見
JER|33|11|歡喜和快樂的聲音、新郎和新娘的聲音，並聽見有人說： 你們要稱謝萬軍之耶和華， 因耶和華本為善， 他的慈愛永遠長存！ 他們奉感謝祭到耶和華的殿中；因為我必使這地被擄的人歸回，如起初一樣。這是耶和華說的。」
JER|33|12|萬軍之耶和華如此說：「在這荒廢、無人、無牲畜之地，並其中所有的城鎮，必再有牧人的草場，可讓羊群躺臥在那裏。
JER|33|13|在山區的城鎮、 謝非拉 的城鎮、 尼革夫 的城鎮、 便雅憫 地、 耶路撒冷 四圍的各處和 猶大 的城鎮，必再有羊群從數點的人手下經過。這是耶和華說的。
JER|33|14|「看哪，日子將到，我應許 以色列 家和 猶大 家的恩言必然實現。這是耶和華說的。
JER|33|15|在那些日子、那時候，我必使 大衛 公義的苗裔長起來；他必在地上施行公平和公義。
JER|33|16|在那些日子， 猶大 必得救， 耶路撒冷 必安然居住，他的名必稱為『耶和華－我們的義』。
JER|33|17|「因為耶和華如此說： 大衛 家必永遠不斷有人坐在 以色列 家的寶座上；
JER|33|18|利未 家的祭司也不斷有人在我面前獻燔祭、燒素祭，時常辦理獻祭的事。」
JER|33|19|耶和華的話臨到 耶利米 ，說：
JER|33|20|「耶和華如此說：你們若能廢棄我所立白日黑夜的約，使白日黑夜不按時輪轉，
JER|33|21|就能廢棄我與我僕人 大衛 所立的約，使他沒有後裔在他的寶座上作王，並能廢棄我與事奉我的 利未 家的祭司所立的約。
JER|33|22|正如天上的萬象不能數算，海邊的塵沙不能斗量，我必照樣使我僕人 大衛 的後裔和事奉我的 利未 人多起來。」
JER|33|23|耶和華的話臨到 耶利米 ，說：
JER|33|24|「你沒有留意這百姓所說的話嗎？他們說：『耶和華所揀選的二族，他已經棄絕了。』他們這樣藐視我的百姓，不把他們當作國來看待。
JER|33|25|耶和華如此說：除非我沒有立白日黑夜之約，也未曾安排天和地的定例，
JER|33|26|否則我不會棄絕 雅各 的後裔和我僕人 大衛 的後裔，使 大衛 的後裔不再治理 亞伯拉罕 、 以撒 、 雅各 的後裔。我必使他們被擄的人歸回，也必憐憫他們。」
JER|34|1|巴比倫 王 尼布甲尼撒 率領他的全軍和地上他管轄的各國各邦，攻打 耶路撒冷 和 耶路撒冷 所有的城鎮。那時，耶和華的話臨到 耶利米 ，說：
JER|34|2|「耶和華－ 以色列 的上帝說，你去告訴 猶大 王 西底家 ，耶和華如此說：看哪，我要把這城交在 巴比倫 王的手中，他必用火焚燒。
JER|34|3|你必不能逃脫他的手，定被拿住，交在他手中。你要親眼看到 巴比倫 王，他要親口跟你說話，你也必到 巴比倫 去。
JER|34|4|猶大 王 西底家 啊，你一定要聽耶和華的話。耶和華論到你如此說：你必不死於刀下；
JER|34|5|必平安而終，人要為你焚燒，好像為你祖先，就是在你以前早先的王焚燒一樣。人要為你舉哀說：『哀哉！我主啊。』這話是我說的。這是耶和華說的。」
JER|34|6|於是， 耶利米 先知在 耶路撒冷 把這一切話告訴 猶大 王 西底家 。
JER|34|7|那時， 巴比倫 王的軍隊正攻打 耶路撒冷 ，又攻打 猶大 僅存的城鎮，就是 拉吉 和 亞西加 ；原來 猶大 的堅固城只剩下這兩座。
JER|34|8|西底家 王與 耶路撒冷 的眾百姓立約，要他們宣告自由，叫各人釋放自己的僕人和婢女，使 希伯來 的男人和女人得自由，誰也不可使他的 猶大 弟兄作奴僕。這事以後，耶和華的話臨到 耶利米 。
JER|34|9|
JER|34|10|所有前來立約的領袖和眾百姓都順從，各人釋放自己的僕人和婢女，使他們得自由，不再叫他們作奴僕。大家都順從，將僕婢釋放了。
JER|34|11|但後來他們又反悔，叫被釋放得自由的僕人婢女回來，強迫他們仍為僕婢。
JER|34|12|因此耶和華的話臨到 耶利米 ，說：
JER|34|13|「耶和華－ 以色列 的上帝如此說：我將你們祖先從 埃及 地為奴之家領出時，與他們立約說：
JER|34|14|『你的一個 希伯來 弟兄若賣給你，服事你六年，到第七年你們各人就要釋放他自由出去。』只是你們祖先不聽我，不側耳而聽。
JER|34|15|如今你們回轉，行我眼中看為正的事，各人向鄰舍宣告自由，並且在我面前、在稱為我名下的殿中立約。
JER|34|16|你們卻反悔，褻瀆我的名，各人叫所釋放得自由的僕人婢女回來，強迫他們仍為僕婢。
JER|34|17|所以耶和華如此說：你們不聽從我，各人不向弟兄鄰舍宣告自由。看哪！我要向你們宣告自由，把你們自由地交給刀劍、饑荒、瘟疫，並且使地上萬國因你們而驚駭。這是耶和華說的。
JER|34|18|那些違背我約的人，就是不遵守在我面前立約之話的，我要使他們成了那劈成兩半的牛犢，使人從切塊中經過：
JER|34|19|猶大 的領袖、 耶路撒冷 的領袖、官員、祭司，和從牛犢切塊中經過的這地的眾百姓，
JER|34|20|我必將他們交在仇敵和尋索其命的人手中；他們的屍首必給空中的飛鳥和地上的走獸作食物。
JER|34|21|我必將 猶大 王 西底家 和他的眾領袖交在仇敵和尋索其命的人手中，與那暫時離你們而去的 巴比倫 王軍隊的手中。
JER|34|22|看哪，我要吩咐他們回到這城，攻打這城，將城攻取，用火焚燒；我也要使 猶大 的城鎮變為廢墟，無人居住。這是耶和華說的。」
JER|35|1|當 約西亞 的兒子 約雅敬 作 猶大 王的時候，耶和華的話臨到 耶利米 ，說：
JER|35|2|「你去見 利甲 族的人，吩咐他們，領他們進入耶和華殿的一個房間，給他們酒喝。」
JER|35|3|我就帶 哈巴洗尼雅 的孫子 雅利米雅 的兒子 雅撒尼亞 ，和他的兄弟，並他所有的兒子，以及 利甲 全族的人，
JER|35|4|領他們到耶和華的殿，進入 伊基大利 的兒子神人 哈難 兒子們的房間；那房間靠近官長的房間，在 沙龍 之子門口的守衛 瑪西雅 的房間上面。
JER|35|5|於是我在 利甲 族的人面前擺設盛滿了酒的碗和杯，對他們說：「請喝酒。」
JER|35|6|他們卻說：「我們不喝酒，因為我們祖先 利甲 的兒子 約拿達 曾吩咐我們說：『你們與你們的子孫永不可喝酒，
JER|35|7|不可蓋房子，不可撒種，也不可栽葡萄園，連擁有都不可；但一生的年日要住帳棚，使你們的日子在寄居的地面上得以長久。』
JER|35|8|凡我們祖先 利甲 的兒子 約拿達 所吩咐我們的話，我們都聽從了。我們和我們的妻子兒女一生的年日都不喝酒，
JER|35|9|不蓋房子居住，我們也沒有葡萄園、田地和種子；
JER|35|10|但住在帳棚裏，聽從並遵行我們祖先 約拿達 所吩咐我們的一切話。
JER|35|11|巴比倫 王 尼布甲尼撒 上來攻打這地的時候，我們說：『來吧，我們到 耶路撒冷 去，躲避 迦勒底 的軍隊和 亞蘭 的軍隊。』這樣，我們才住在 耶路撒冷 。」
JER|35|12|耶和華的話臨到 耶利米 ，說：
JER|35|13|「萬軍之耶和華－ 以色列 的上帝如此說：你去對 猶大 人和 耶路撒冷 的居民說，你們不肯領受訓誨，聽從我的話嗎？這是耶和華說的。
JER|35|14|利甲 的兒子 約拿達 所吩咐他子孫不可喝酒的話，他們已經遵守了；他們因為聽從祖先的吩咐，直到今日都不喝酒。至於我，我一再警戒你們，你們卻不肯聽從我。
JER|35|15|我一再差遣我的僕人眾先知到你們那裏去，說：『你們各人當回頭離開惡道，改正行為，不再隨從事奉別神，如此，就必住在我所賜給你們和你們祖先的地上。』只是你們不側耳而聽，也不聽我。
JER|35|16|利甲 的兒子 約拿達 的子孫能遵守祖先所吩咐他們的命令，這百姓卻不肯聽從我！
JER|35|17|因此，耶和華－萬軍之上帝、 以色列 的上帝如此說：看哪，我要使我所說的一切災禍臨到 猶大 人和 耶路撒冷 所有的居民。因為我向他們說話，他們不聽從；我呼喚他們，他們也沒有回應。」
JER|35|18|耶利米 對 利甲 族的人說：「萬軍之耶和華－ 以色列 的上帝如此說：因你們聽從你們祖先 約拿達 的吩咐，謹守他的一切命令，照他所吩咐的去做，
JER|35|19|所以萬軍之耶和華－ 以色列 的上帝如此說： 利甲 的兒子 約拿達 必永遠不斷有人侍立在我面前。」
JER|36|1|約西亞 的兒子 猶大 王 約雅敬 第四年，有這話從耶和華臨到 耶利米 ，說：
JER|36|2|「你要取一書卷，把我對你所說攻擊 以色列 和 猶大 ，並各國的一切話，從我對你說話的那日，就是從 約西亞 的日子起直到今日，都寫在其上；
JER|36|3|或者 猶大 家聽見我想要降給他們的一切災禍，各人就回轉離開惡道，我就赦免他們的罪孽和罪惡。」
JER|36|4|耶利米 召了 尼利亞 的兒子 巴錄 來； 巴錄 就從 耶利米 口中，把耶和華對 耶利米 所說的一切話寫在書卷上。
JER|36|5|耶利米 吩咐 巴錄 說：「我被禁止，不能進耶和華的殿。
JER|36|6|所以你要趁禁食的日子進入耶和華的殿中，把耶和華的話，就是你從我口中寫在書卷上的話，念給百姓和所有從各城鎮前來的 猶大 人親耳聽；
JER|36|7|或者他們的懇求達到耶和華面前，各人回轉離開惡道，因為耶和華向這百姓所說要發的怒氣和憤怒實在很大。」
JER|36|8|尼利亞 的兒子 巴錄 就照 耶利米 先知所吩咐的一切去做，在耶和華殿中宣讀書卷上耶和華的話。
JER|36|9|約西亞 的兒子 猶大 王 約雅敬 第五年九月， 耶路撒冷 的眾百姓和那從 猶大 城鎮前來 耶路撒冷 的眾百姓，在耶和華面前宣告禁食，
JER|36|10|巴錄 就在耶和華殿的上院，靠近耶和華殿的 新門 口， 沙番 的兒子 基瑪利雅 文士的房間裏，宣讀書卷上 耶利米 的話給眾百姓親耳聽。
JER|36|11|沙番 的孫子 基瑪利雅 的兒子 米該亞 聽見書卷上耶和華的一切話，
JER|36|12|就下到王宮，進入書記的房間。看哪，所有的官長都坐在那裏，包括 以利沙瑪 文士、 示瑪雅 的兒子 第萊雅 、 亞革波 的兒子 以利拿單 、 沙番 的兒子 基瑪利雅 、 哈拿尼雅 的兒子 西底家 和其餘的官長。
JER|36|13|米該亞 向他們述說他所聽見的一切話，就是當 巴錄 向眾百姓宣讀那書卷時親耳聽見的。
JER|36|14|官長們就派 猶底 ，就是 古示 的曾孫， 示利米雅 的孫子， 尼探雅 的兒子到 巴錄 那裏，對他說：「你把你所念給百姓聽的書卷拿在手裏，到我們這裏來。」 尼利亞 的兒子 巴錄 就手拿書卷到他們那裏來。
JER|36|15|他們對他說：「請坐下，念給我們親耳聽。」 巴錄 就念給他們親耳聽。
JER|36|16|他們聽見這一切話就害怕，面面相覷，對 巴錄 說：「我們必須將這一切話稟告王。」
JER|36|17|他們問 巴錄 說：「請你告訴我們，你怎樣從他口中寫下這一切話呢？」
JER|36|18|巴錄 回答說：「他向我口述這一切話，我就用筆墨把它寫在書卷上。」
JER|36|19|眾官長對 巴錄 說：「你和 耶利米 要去躲起來，不可叫人知道你們躲在哪裏。」
JER|36|20|眾官長把書卷留在 以利沙瑪 文士的房間裏，然後進院見王，把這一切話說給王聽。
JER|36|21|王就派 猶底 去拿這書卷來；他就從 以利沙瑪 文士的房間內取來，念給王和侍立在王左右的眾官長親耳聽。
JER|36|22|那時正是九月，王坐在過冬的房屋裏，王前面有燃燒的火盆 。
JER|36|23|猶底 念了三、四段 ，王就用文士的刀把書卷割破，丟在火盆裏，直到全卷在火中燒盡了。
JER|36|24|王和聽見這一切話的臣僕都不懼怕，也不撕裂衣服。
JER|36|25|以利拿單 和 第萊雅 ，並 基瑪利雅 懇求王不要燒這書卷，王卻不聽。
JER|36|26|王吩咐王 的兒子 耶拉篾 、 亞斯列 的兒子 西萊雅 和 亞伯疊 的兒子 示利米雅 ，去捉拿 巴錄 文士和 耶利米 先知；耶和華卻將他們隱藏起來。
JER|36|27|王燒了有 巴錄 從 耶利米 口中所寫之話的書卷以後，耶和華的話臨到 耶利米 ，說：
JER|36|28|「你再取一書卷，將 猶大 王 約雅敬 所燒前一卷書上原有的一切話寫在上面。
JER|36|29|論到 猶大 王 約雅敬 你要說，耶和華如此說：你燒了這書卷，說：『你為甚麼在上面寫著， 巴比倫 王必要來毀滅這地，使這地絕了人民和牲畜呢？』
JER|36|30|所以耶和華論到 猶大 王 約雅敬 說：他後裔中必沒有人坐在 大衛 的寶座上；他的屍首必被拋棄，白天受炎熱，黑夜受寒霜。
JER|36|31|我必因他和他後裔，並他臣僕的罪孽懲罰他們。我要使我所說的一切災禍臨到他們和 耶路撒冷 的居民，並 猶大 人；只是他們不肯聽從。」
JER|36|32|於是， 耶利米 又取一書卷交給 尼利亞 的兒子 巴錄 文士，他就從 耶利米 的口中寫了 猶大 王 約雅敬 在火中所燒書卷上的一切話，另外又添了許多相仿的話。
JER|37|1|約西亞 的兒子 西底家 接續 約雅敬 的兒子 哥尼雅 作王，因為 巴比倫 王 尼布甲尼撒 立他在 猶大 地作王。
JER|37|2|但 西底家 、他的臣僕和這地的百姓都不聽從耶和華藉 耶利米 先知所說的話。
JER|37|3|西底家 王派 示利米雅 的兒子 猶甲 和 瑪西雅 的兒子 西番雅 祭司，去見 耶利米 先知，說：「求你為我們祈求耶和華－我們的上帝。」
JER|37|4|那時 耶利米 仍在百姓中進出，因為他們還沒有把他囚在監裏。
JER|37|5|法老的軍隊已經從 埃及 出來，那圍困 耶路撒冷 的 迦勒底 人聽見這風聲，就拔營離開 耶路撒冷 去了。
JER|37|6|耶和華的話臨到 耶利米 先知，說：
JER|37|7|「耶和華－ 以色列 的上帝如此說：你們要對派你們來求問我的 猶大 王如此說：『看哪，那出來幫助你們的法老軍隊必回 埃及 本國去。
JER|37|8|迦勒底 人必再來攻打這城，並要攻下，用火焚燒。
JER|37|9|耶和華如此說：你們不要自欺說「 迦勒底 人必定離開我們」，因為他們必不離開。
JER|37|10|你們即使擊敗與你們爭戰的 迦勒底 全軍，他們當中剩下受傷的人也必各自從帳棚裏起來，用火焚燒這城。』」
JER|37|11|迦勒底 的軍隊因躲避法老的軍隊，拔營離開 耶路撒冷 的時候，
JER|37|12|耶利米 離開 耶路撒冷 ，往 便雅憫 地去，要在那裏從百姓當中取得自己的地產。
JER|37|13|他到了 便雅憫門 ，那裏的守門官名叫 伊利雅 ，是 哈拿尼亞 的孫子， 示利米雅 的兒子，他逮捕 耶利米 先知，說：「你是去投降 迦勒底 人的！」
JER|37|14|耶利米 說：「你這是謊話，我並不是去投降 迦勒底 人。」 伊利雅 不聽 耶利米 的話，就逮捕他，把他帶到官長那裏。
JER|37|15|官長們惱怒 耶利米 ，打了他，把他囚在 約拿單 文士的房屋中，因為他們把這屋子當作監牢。
JER|37|16|耶利米 來到地牢，進入牢房，在那裏拘留多日。
JER|37|17|西底家 王差人提他出來，在自己的宮內私下問他說：「有甚麼話從耶和華臨到沒有？」 耶利米 說：「有！」又說：「你必被交在 巴比倫 王手中。」
JER|37|18|耶利米 又對 西底家 王說：「我在甚麼事上得罪你，或你的臣僕，或這百姓，你們竟將我囚在監裏呢？
JER|37|19|對你們預言『 巴比倫 王必不來攻擊你們和這地』的先知在哪裏呢？
JER|37|20|主－我的王啊，現在求你垂聽，允准我在你面前的懇求：不要把我送回 約拿單 文士的房屋中，免得我死在那裏。」
JER|37|21|於是 西底家 王下令，他們就把 耶利米 交在護衛兵的院中，每天從餅店街取一個餅給他，直到城中所有的餅都用盡了。這樣， 耶利米 仍拘留在護衛兵的院中。
JER|38|1|瑪坦 的兒子 示法提雅 、 巴施戶珥 的兒子 基大利 、 示利米雅 的兒子 猶甲 、 瑪基雅 的兒子 巴示戶珥 聽見 耶利米 對眾百姓所說的話，說：
JER|38|2|「耶和華如此說：留在這城裏的必遭刀劍、饑荒、瘟疫而死，但歸向 迦勒底 人的必得存活；至少能保全自己的性命，得以存活。
JER|38|3|耶和華如此說：這城必要交在 巴比倫 王軍隊的手中，他必攻下這城。」
JER|38|4|於是官長們對王說：「求你把這人處死，因他向城裏剩下的士兵和眾人說這樣的話，使他們的手發軟。這人不是為這百姓求平安，而是叫他們受災禍。」
JER|38|5|西底家 王說：「看哪，他在你們手中，王不能反對你們所做的事。」
JER|38|6|他們就拿住 耶利米 ，把他丟在王 的兒子 瑪基雅 的井裏；那口井在護衛兵的院中。他們用繩子把 耶利米 縋下去，井裏沒有水，只有淤泥， 耶利米 就陷在淤泥中。
JER|38|7|在王宮裏的太監 古實 人 以伯‧米勒 ，聽見他們把 耶利米 丟進井裏，那時王坐在 便雅憫門 前。
JER|38|8|以伯‧米勒 從王宮裏出來，對王說：
JER|38|9|「主－我的王啊，這些人向 耶利米 先知一味地行惡，把他丟在井裏；他在那裏必因飢餓而死，因為城裏不再有糧食了。」
JER|38|10|王就吩咐 古實 人 以伯‧米勒 說：「你從這裏帶領三十人，趁 耶利米 先知還沒死，把他從井裏拉上來。」
JER|38|11|於是 以伯‧米勒 帶領這些人同去，進入王宮，到庫房以下 ，從那裏取了些碎布和破衣服，用繩子縋下去，到井裏 耶利米 那裏。
JER|38|12|古實 人 以伯‧米勒 對 耶利米 說：「你用這些碎布和破衣服放在繩子上，墊你的腋下。」 耶利米 就照樣做。
JER|38|13|這樣，他們用繩子將 耶利米 從井裏拉上來。 耶利米 仍在護衛兵的院中。
JER|38|14|西底家 王差人將 耶利米 先知帶進耶和華殿的第三個門，到王那裏去。王對 耶利米 說：「我要問你一件事，你一點都不可向我隱瞞。」
JER|38|15|耶利米 對 西底家 說：「我若告訴你，你豈不是一定要把我處死嗎？我若勸你，你必不聽我。」
JER|38|16|西底家 王就私下對 耶利米 說：「我指著那造我們生命之永生的耶和華起誓：我必不把你處死，也不將你交在尋索你命的人手中。」
JER|38|17|耶利米 對 西底家 說：「耶和華－萬軍之上帝、 以色列 的上帝如此說：你若歸順 巴比倫 王的官長，你的命就必存活，這城也不致被火焚燒，你和你的全家都必存活。
JER|38|18|你若不歸順 巴比倫 王的官長，這城必交在 迦勒底 人手中。他們必用火焚燒，你也不得脫離他們的手。」
JER|38|19|西底家 王對 耶利米 說：「我怕那些投降 迦勒底 人的 猶大 人，恐怕 迦勒底 人把我交在他們手中，他們就戲弄我。」
JER|38|20|耶利米 說：「 迦勒底 人必不把你交出。求你聽從我對你所說耶和華的話，這樣對你有好處，你的命也必存活。
JER|38|21|你若不肯歸順，耶和華指示我的話是這樣：
JER|38|22|看哪， 猶大 王宮裏所留下來的婦女必被帶到 巴比倫 王的官長那裏。這些婦女要說： 你知己的朋友引誘你， 他們勝過你； 你的腳陷入淤泥， 他們卻離棄你。
JER|38|23|「人必將你的后妃和你的兒女帶到 迦勒底 人那裏；你也不得脫離他們的手，必被 巴比倫 王的手捉住，這城也必被火焚燒 。」
JER|38|24|西底家 對 耶利米 說：「不要讓人知道這些對話，你就不至於死。
JER|38|25|官長們若聽見我跟你說話，到你那裏對你說：『告訴我們，你對王說了甚麼話，王又向你說了甚麼；不可向我們隱瞞，否則我們就要殺你。』
JER|38|26|你就對他們說：『我在王面前懇求不要把我送回 約拿單 的房屋，免得我死在那裏。』」
JER|38|27|隨後官長們到 耶利米 那裏，問他，他就照王所吩咐的一切話回答他們。他們就不再問他，因為事情沒有洩漏。
JER|38|28|於是 耶利米 仍在護衛兵的院中，直到 耶路撒冷 被攻下的日子。當 耶路撒冷 被攻下時，他仍在那裏。
JER|39|1|猶大 王 西底家 第九年十月， 巴比倫 王 尼布甲尼撒 率領全軍前來圍困 耶路撒冷 。
JER|39|2|西底家 十一年四月初九日，城被攻破。
JER|39|3|耶路撒冷 被攻下的時候， 巴比倫 王的眾官長， 尼甲‧沙利薛 、 三甲‧尼波 、 撒西金 將軍 、 尼甲‧沙利薛 將軍 ，並 巴比倫 王其餘的官長都來坐在 中門 。
JER|39|4|猶大 王 西底家 和所有士兵看見他們，就在夜間從靠近王的花園、兩城牆中間的門逃跑出城，往 亞拉巴 逃去。
JER|39|5|迦勒底 的軍隊追趕他們，在 耶利哥 的平原追上 西底家 ，將他逮住，帶到 哈馬 地的 利比拉 、 巴比倫 王 尼布甲尼撒 那裏； 尼布甲尼撒 就判他的罪。
JER|39|6|在 利比拉 ， 巴比倫 王在 西底家 眼前殺了他的兒女； 巴比倫 王又殺了 猶大 所有的貴族，
JER|39|7|並且挖了 西底家 的眼睛，用銅鏈鎖住他，要帶到 巴比倫 去。
JER|39|8|迦勒底 人用火焚燒王宮和百姓的房屋，又拆毀 耶路撒冷 的城牆。
JER|39|9|那時， 尼布撒拉旦 護衛長把城裏所剩下的百姓和投降他的降民，以及其餘的百姓都擄到 巴比倫 去了。
JER|39|10|尼布撒拉旦 護衛長卻把百姓中一無所有的窮人留在 猶大 地，當時就賞給他們葡萄園和田地 。
JER|39|11|巴比倫 王 尼布甲尼撒 為了 耶利米 ，囑咐 尼布撒拉旦 護衛長：
JER|39|12|「你領他去，好好地看待他，切不可害他；他對你怎麼說，你就向他怎樣做。」
JER|39|13|尼布撒拉旦 護衛長和 尼布沙斯班 將軍 、 尼甲‧沙利薛 將軍 ，並 巴比倫 王眾官長，
JER|39|14|派人把 耶利米 從護衛兵的院中提出來，交給 沙番 的孫子， 亞希甘 的兒子 基大利 ，讓他自由進出屋子；於是 耶利米 住在百姓中間。
JER|39|15|耶利米 還囚在護衛兵院中的時候，耶和華的話臨到他，說：
JER|39|16|「你去告訴 古實 人 以伯‧米勒 說，萬軍之耶和華－ 以色列 的上帝如此說：看哪，我說降禍不降福的話必臨到這城，到那時必在你面前實現。
JER|39|17|到那日我必拯救你，你必不致交在你所怕的人手中。這是耶和華說的。
JER|39|18|我定要搭救你，你必不致倒在刀下，卻要保全自己的性命，因你倚靠我。這是耶和華說的。」
JER|40|1|耶利米 被鏈子鎖在 耶路撒冷 和 猶大 被擄到 巴比倫 的人中， 尼布撒拉旦 護衛長把他從 拉瑪 提出來，釋放他以後，耶和華的話臨到 耶利米 。
JER|40|2|護衛長提 耶利米 來，對他說：「耶和華－你的上帝曾說要降這災禍給此地。
JER|40|3|耶和華照他所說的做了，已使這災禍臨到；因你們得罪耶和華，不聽從他的話，所以這事臨到你們。
JER|40|4|看哪，現在我解開你手上的鏈子，你若看與我同往 巴比倫 去好，就可以去，我必厚待你；你若看與我同往 巴比倫 去不好，就不必去。看哪，全地在你面前，你以為哪裏美好，哪裏合宜，只管去吧
JER|40|5|─ 耶利米 尚未回去 ─你可以回到 巴比倫 王所立管理 猶大 城鎮的 沙番 的孫子， 亞希甘 的兒子 基大利 那裏去，在他那裏住在百姓當中。不然，你看哪裏合宜就可以去。」於是護衛長送他糧食和禮物，釋放了他。
JER|40|6|耶利米 就來到 米斯巴 ， 亞希甘 的兒子 基大利 那裏去，與他同住，住在留於境內的百姓當中。
JER|40|7|在鄉間所有的軍官和屬他們的人，聽見 巴比倫 王立了 亞希甘 的兒子 基大利 作當地的省長，並將沒有擄到 巴比倫 的男人、婦女、孩童和當地極窮的人全交給他，
JER|40|8|於是 尼探雅 的兒子 以實瑪利 ， 加利亞 的兩個兒子 約哈難 和 約拿單 ， 單戶篾 的兒子 西萊雅 ，並 尼陀法 人 以斐 的眾子， 瑪迦 人的兒子 耶撒尼亞 ，和屬他們的人，都來到 米斯巴 的 基大利 那裏。
JER|40|9|沙番 的孫子， 亞希甘 的兒子 基大利 向他們和屬他們的人起誓說：「不要怕服事 迦勒底 人，只管住在這地，服事 巴比倫 王，就可以得福。
JER|40|10|至於我，我要住在 米斯巴 ，侍候那些到我們這裏來的 迦勒底 人；只是你們當積蓄酒、油和夏天的果子，收藏在器皿裏，並住在你們所佔的城鎮中。」
JER|40|11|在 摩押 地和 亞捫 人當中，在 以東 地和各國，所有的 猶大 人聽見 巴比倫 王留下一些 猶大 人，並立 沙番 的孫子、 亞希甘 的兒子 基大利 管理他們，
JER|40|12|所有的 猶大 人就從被趕到的各處回來，到 猶大 地 米斯巴 的 基大利 那裏。他們積蓄了許多的酒，並夏天的果子。
JER|40|13|加利亞 的兒子 約哈難 和在鄉間的軍官來到 米斯巴 的 基大利 那裏，
JER|40|14|對他說：「 亞捫 人的王 巴利斯 派 尼探雅 的兒子 以實瑪利 來謀害你的命，你知道嗎？」 亞希甘 的兒子 基大利 卻不相信他們的話。
JER|40|15|加利亞 的兒子 約哈難 在 米斯巴 私下對 基大利 說：「求你容我去殺 尼探雅 的兒子 以實瑪利 ，必無人知道。何必讓他害你的命，使聚集到你這裏來的 猶大 人都分散，以致 猶大 剩餘的人都滅亡呢？」
JER|40|16|亞希甘 的兒子 基大利 對 加利亞 的兒子 約哈難 說：「你不可做這事，你所論 以實瑪利 的話是假的。」
JER|41|1|七月中，王的大臣，就是王室後裔 以利沙瑪 的孫子、 尼探雅 的兒子 以實瑪利 帶著十個人，來到 米斯巴 ， 亞希甘 的兒子 基大利 那裏；他們在 米斯巴 一同吃飯。
JER|41|2|尼探雅 的兒子 以實瑪利 和同他來的那十個人起來，用刀擊殺 沙番 的孫子， 亞希甘 的兒子 基大利 ，就是 巴比倫 王所立為當地省長的，把他殺死。
JER|41|3|以實瑪利 把所有在 米斯巴 與 基大利 一起的 猶大 人，以及他們在那裏所遇見的 迦勒底 人和士兵都殺了。
JER|41|4|他殺了 基大利 的第二天，還沒有人知道的時候，
JER|41|5|有八十人從 示劍 、 示羅 和 撒瑪利亞 前來，鬍鬚剃去，衣服撕裂，身體劃破，手拿素祭和乳香，要奉到耶和華的殿。
JER|41|6|尼探雅 的兒子 以實瑪利 從 米斯巴 出來迎接他們，隨走隨哭，遇見了他們，就對他們說：「你們可以到 亞希甘 的兒子 基大利 那裏。」
JER|41|7|他們到了城中， 尼探雅 的兒子 以實瑪利 和與他一起的人就把他們殺了，丟在坑裏。
JER|41|8|只是他們中間有十個人對 以實瑪利 說：「不要殺我們，因為我們有許多大麥、小麥、油和蜜藏在田間。」於是他住手，沒有在弟兄中間殺他們。
JER|41|9|以實瑪利 把那些因 基大利 事件所殺之人的屍首都丟在坑裏；這坑是從前 亞撒 王因怕 以色列 王 巴沙 所挖的。 尼探雅 的兒子 以實瑪利 把那些被殺的人填滿了坑。
JER|41|10|以實瑪利 把 米斯巴 剩下的人，就是眾公主和仍住在 米斯巴 所有的百姓都擄去，他們原是 尼布撒拉旦 護衛長交給 亞希甘 的兒子 基大利 的。 尼探雅 的兒子 以實瑪利 擄了他們，要到 亞捫 人那裏去。
JER|41|11|加利亞 的兒子 約哈難 和與他一起的軍官，聽見 尼探雅 的兒子 以實瑪利 所做的一切惡事，
JER|41|12|就帶領眾人前往，要和 尼探雅 的兒子 以實瑪利 爭戰，他們在 基遍 的大水池 旁遇見他。
JER|41|13|在 以實瑪利 那裏的眾人看見 加利亞 的兒子 約哈難 和與他一起的軍官，就都歡喜。
JER|41|14|這樣， 以實瑪利 從 米斯巴 所擄去的眾人都轉而歸向 加利亞 的兒子 約哈難 。
JER|41|15|尼探雅 的兒子 以實瑪利 和八個人脫離 約哈難 的手，逃到 亞捫 人那裏去。
JER|41|16|尼探雅 的兒子 以實瑪利 殺了 亞希甘 的兒子 基大利 ，從 米斯巴 把所有倖存的百姓、士兵、婦女、孩童、太監擄到 基遍 之後， 加利亞 的兒子 約哈難 和與他一起的軍官把他們都搶回來，
JER|41|17|帶到靠近 伯利恆 的 基羅特金罕 住下，要到 埃及 去，
JER|41|18|躲避 迦勒底 人。他們懼怕 迦勒底 人，因為 尼探雅 的兒子 以實瑪利 殺了 巴比倫 王所立管理那地的 亞希甘 的兒子 基大利 。
JER|42|1|眾軍官和 加利亞 的兒子 約哈難 ，並 何沙雅 的兒子 耶撒尼亞 以及眾百姓，從最小的到最大的都進前來，
JER|42|2|對 耶利米 先知說：「請你准我們在你面前祈求，為我們這倖存的人向耶和華－你的上帝禱告。我們本來眾多，現在剩下的極少，這是你親眼看見的。
JER|42|3|願耶和華－你的上帝指示我們當走的路，當做的事。」
JER|42|4|耶利米 先知對他們說：「我已經聽見了，看哪，我必照你們的話向耶和華－你們的上帝禱告。耶和華無論回答甚麼，我都必告訴你們，絕不隱瞞。」
JER|42|5|於是他們對 耶利米 說：「我們若不照耶和華－你上帝差遣你說的一切話去做，願耶和華在我們中間作真實可靠的見證。
JER|42|6|我們請你到耶和華－我們的上帝面前，他說的無論是好是歹，我們都必聽從；因為我們聽從耶和華－我們上帝的話，就可以得福。」
JER|42|7|過了十天，耶和華的話臨到 耶利米 。
JER|42|8|他就將 加利亞 的兒子 約哈難 和與他一起所有的軍官和百姓，從最小的到最大的都召來，
JER|42|9|對他們說：「你們請我到耶和華－ 以色列 的上帝面前為你們祈求，他如此說：
JER|42|10|『你們若仍留在這地，我就建立你們，必不拆毀；栽植你們，必不拔出；因我為所降與你們的災禍感到遺憾。
JER|42|11|不要怕你們所懼怕的 巴比倫 王。不要怕他！因為我與你們同在，要拯救你們脫離他的手。這是耶和華說的。
JER|42|12|我要向你們施憐憫，他 就憐憫你們，使你們歸回本地。』
JER|42|13|倘若你們說：『我們不留在這地』，不聽從耶和華－你們上帝的話，
JER|42|14|說：『我們不留在這地，卻要進入 埃及 地，在那裏我們看不見戰爭，聽不見角聲，也不致缺食挨餓；我們要住在那裏。』
JER|42|15|倖存的 猶大 人哪，你們現在要聽耶和華的話；萬軍之耶和華－ 以色列 的上帝如此說：『你們若定意進入 埃及 ，在那裏寄居，
JER|42|16|你們所懼怕的刀劍在 埃及 地必追上你們，你們所懼怕的饑荒在 埃及 要緊緊跟隨你們，你們必死在那裏。
JER|42|17|凡定意進入 埃及 在那裏寄居的，必遭刀劍、饑荒、瘟疫而死，無一人存留，得以逃脫我所降與他們的災禍。』
JER|42|18|「萬軍之耶和華－ 以色列 的上帝如此說：『我怎樣將我的怒氣和憤怒傾倒在 耶路撒冷 的居民身上，你們進入 埃及 的時候，我也必照樣將我的憤怒傾倒在你們身上，以致你們受辱罵、驚駭、詛咒、羞辱，並且不得再看見這地方。』
JER|42|19|倖存的 猶大 人哪，耶和華論到你們說：『不要進入 埃及 。』你們要確實知道，我今日已警戒你們了。
JER|42|20|你們行詭詐害自己；因為你們請我到耶和華－你們上帝那裏，說：『請你為我們向耶和華－我們的上帝禱告，你把耶和華－我們上帝所說的一切告訴我們，我們就必遵行。』
JER|42|21|我今日把這話告訴你們，你們卻不聽耶和華－你們上帝為這一切事差我到你們那裏所說的話。
JER|42|22|現在你們要確實知道，你們在所要去的寄居之地必遭刀劍、饑荒、瘟疫而死。」
JER|43|1|耶利米 向眾百姓說完了耶和華－他們上帝一切的話，就是耶和華－他們上帝差他去說的這一切話，
JER|43|2|何沙雅 的兒子 亞撒利雅 和 加利亞 的兒子 約哈難 ，以及所有狂傲的人，就對 耶利米 說：「你說謊！耶和華－我們的上帝並沒有差遣你說：『你們不可進入 埃及 ，在那裏寄居。』
JER|43|3|這是 尼利亞 的兒子 巴錄 挑唆你害我們，要把我們交在 迦勒底 人手中，使我們被殺或被擄到 巴比倫 去。」
JER|43|4|加利亞 的兒子 約哈難 和所有的軍官、百姓，都不肯聽從耶和華的話留在 猶大 地。
JER|43|5|加利亞 的兒子 約哈難 和所有的軍官卻將倖存的 猶大 人，就是從被趕到的各國回來，在 猶大 地寄居的男人、婦女、孩童和眾公主，並 尼布撒拉旦 護衛長留在 沙番 的孫子， 亞希甘 的兒子 基大利 那裏的眾人，與 耶利米 先知，以及 尼利亞 的兒子 巴錄 ，
JER|43|6|
JER|43|7|都帶入 埃及 地，到了 答比匿 ；這是因他們不肯聽從耶和華的話。
JER|43|8|在 答比匿 ，耶和華的話臨到 耶利米 ，說：
JER|43|9|「你要在 猶大 人眼前用手拿幾塊大石頭，藏在 答比匿 法老的宮門砌磚的石墩上，
JER|43|10|對他們說：『萬軍之耶和華－ 以色列 的上帝如此說：看哪，我必召我的僕人 巴比倫 王 尼布甲尼撒 前來，安置他的寶座在所藏的這些石頭上；他要在其上支搭華麗的帳幕。
JER|43|11|他要來攻擊 埃及 地： 定為死亡的，必致死亡； 定為擄掠的，必遭擄掠； 定為刀殺的，必被刀殺。
JER|43|12|我要用火點燃 埃及 眾神明的廟宇， 巴比倫 王要焚燒廟宇，擄去神像；他要圍住 埃及 地，好像牧人披上外衣，從那裏安然而去。
JER|43|13|他必打碎 埃及 地 伯‧示麥 的柱像，用火焚燒 埃及 眾神明的廟宇。』」
JER|44|1|有話臨到 耶利米 ，論到住 埃及 地所有的 猶大 人，就是住在 密奪 、 答比匿 、 挪弗 、 巴特羅 境內的 猶大 人，說：
JER|44|2|「萬軍之耶和華－ 以色列 的上帝如此說：我所降與 耶路撒冷 和 猶大 各城的一切災禍，你們都看見了。看哪，那些城鎮今日荒涼，無人居住；
JER|44|3|這是因居民所行的惡，去燒香事奉別神，就是他們和你們，以及你們列祖所不認識的神明，惹我發怒。
JER|44|4|我一再差遣我的僕人眾先知去，說：你們切不可行我所厭惡這可憎之事。
JER|44|5|他們卻不聽從，不側耳而聽，也不轉離惡事，仍向別神燒香。
JER|44|6|因此，我的怒氣和憤怒都傾倒出來，在 猶大 城鎮和 耶路撒冷 街市上燃起，以致它們都荒廢淒涼，正如今日一樣。
JER|44|7|現在耶和華－萬軍之上帝、 以色列 的上帝如此說：你們為何做這大惡自害己命，使你們的男人、婦女、孩童和吃奶的都從 猶大 剪除，不留一人呢？
JER|44|8|你們以手所做的，在寄居的 埃及 地向別神燒香，惹我發怒，使你們被剪除，在天下萬國中受詛咒羞辱。
JER|44|9|你們祖先的惡行， 猶大 諸王和后妃的惡行，你們自己和你們妻子的惡行，就是在 猶大 地和 耶路撒冷 街市上所做的，你們都忘了嗎？
JER|44|10|到如今你們還不懊悔，不懼怕，不肯遵行我在你們和你們祖先面前所設立的法度律例。
JER|44|11|「所以萬軍之耶和華－ 以色列 的上帝如此說：看哪，我必向你們變臉降災，剪除 猶大 眾人。
JER|44|12|我必使那定意進入 埃及 地、在那裏寄居的，就是倖存的 猶大 人，盡都滅絕。他們必在 埃及 地仆倒，因刀劍饑荒滅絕，從最小的到最大的都必遭刀劍饑荒而死，甚至受辱罵、驚駭、詛咒、羞辱。
JER|44|13|我怎樣用刀劍、饑荒、瘟疫懲罰 耶路撒冷 ，也必照樣懲罰那些住在 埃及 地的 猶大 人。
JER|44|14|那進入 埃及 地、在那裏寄居的，就是倖存的 猶大 人，都不得逃脫，也不得歸回 猶大 地。他們心中很想歸回，居住在那裏；但除了少數逃脫的以外，都不得歸回。」
JER|44|15|那些知道自己妻子向別神燒香的男人，與站在那裏的一大群婦女，就是住 埃及 地 巴特羅 所有的百姓，回答 耶利米 說：
JER|44|16|「論到你奉耶和華的名向我們所說的話，我們必不聽從。
JER|44|17|我們定要照我們口中所說的一切話去做，向天后燒香，獻澆酒祭，按著我們與我們祖先、君王、官長在 猶大 城鎮和 耶路撒冷 街市上素常所做的一樣；因為那時我們得以吃飽、享福樂，並未遇見災禍。
JER|44|18|自從我們停止向天后燒香，獻澆酒祭，我們倒缺乏這一切，又因刀劍饑荒滅絕。」
JER|44|19|婦女們說 ：「我們向天后燒香，獻澆酒祭，做天后像的餅供奉它，向它獻澆酒祭，難道我們的丈夫沒有參與嗎？」
JER|44|20|耶利米 對這樣回答他的男人和婦女說：
JER|44|21|「你們與你們祖先、君王、官長，以及這地的百姓，在 猶大 城鎮和 耶路撒冷 街市上所燒的香，耶和華豈不記得，放在他心上嗎？
JER|44|22|耶和華因你們所行的惡、所做可憎的事，不能再容忍，所以使你們的地荒涼，受驚駭詛咒，無人居住，正如今日一樣。
JER|44|23|你們燒香，得罪耶和華，不聽耶和華的話，不遵行他的律法、條例、法度，所以你們遭遇這災禍，正如今日一樣。」
JER|44|24|耶利米 又對眾百姓和婦女說：「所有在 埃及 地的 猶大 人哪，當聽耶和華的話。
JER|44|25|萬軍之耶和華－ 以色列 的上帝如此說：你們和你們的妻子口中說過、手裏做到，說：『我們定要向天后還願，向它燒香，獻澆酒祭。』現在你們儘管堅定所許的願，去還願吧！
JER|44|26|所有住 埃及 地的 猶大 人哪，當聽耶和華的話。耶和華說：看哪，我指著我至大的名起誓，在 埃及 全地，我的名必不再被 猶大 任何人的口呼喊：『我指著主－永生的耶和華起誓。』
JER|44|27|看哪，我看守他們，為要降禍不降福；在 埃及 地的 猶大 人必因刀劍、饑荒而滅亡，直到滅絕。
JER|44|28|從 埃及 地能脫離刀劍、歸回 猶大 地的人數很少。那進入 埃及 地、在那裏寄居的，就是倖存的 猶大 人，必知道是誰的話站得住，是我的話呢，還是他們的話。
JER|44|29|我在這地方懲罰你們，必有預兆，使你們知道我降禍給你們的話必站得住。這是耶和華說的。
JER|44|30|耶和華如此說：看哪，我必將 埃及 王 合弗拉 法老交在他仇敵和尋索其命的人手中，像我將 猶大 王 西底家 交在他仇敵和尋索其命的 巴比倫 王 尼布甲尼撒 手中一樣。」
JER|45|1|約西亞 的兒子 猶大 王 約雅敬 第四年， 尼利亞 的兒子 巴錄 把 耶利米 先知口中所說的話寫在書上； 耶利米 對 巴錄 說：
JER|45|2|「 巴錄 啊，耶和華－ 以色列 的上帝說：
JER|45|3|你曾說：『哀哉！耶和華使我愁上加愁，我因呻吟而困乏，不得安歇。』
JER|45|4|你要這樣告訴他，耶和華如此說：看哪，我所建立的，我必拆毀；我所栽植的，我必拔出；在全地我都如此行。
JER|45|5|你為自己圖謀大事嗎？不要圖謀！看哪，我必使災禍臨到凡有血肉之軀的。但你無論往哪裏去，我要保全你的性命。這是耶和華說的。」
JER|46|1|耶和華論列國的話臨到 耶利米 先知。
JER|46|2|論到 埃及 ，關於 埃及 王 尼哥 法老的軍隊，這軍隊安營在 幼發拉底河 邊的 迦基米施 ，是 巴比倫 王 尼布甲尼撒 在 約西亞 的兒子 猶大 王 約雅敬 第四年所打敗的。
JER|46|3|你們要預備大小盾牌， 往前上陣，
JER|46|4|套上車， 騎上馬！ 頂盔站立， 磨槍披甲！
JER|46|5|我為何看見他們驚惶， 轉身退後呢？ 他們的勇士打敗仗， 急忙逃跑，並不回頭； 四圍都有驚嚇！ 這是耶和華說的。
JER|46|6|不要容快跑的逃避， 也不要容勇士逃脫 ； 在北方 幼發拉底河 邊， 他們絆跌仆倒。
JER|46|7|這是誰，像 尼羅河 漲溢， 如江河的水翻騰呢？
JER|46|8|埃及 像 尼羅河 漲溢， 如江河的水翻騰。 它說：「我要漲溢遮蓋全地； 我要毀滅城鎮和其中的居民。
JER|46|9|馬匹啊，上去吧！ 戰車啊，要疾行！ 手拿盾牌的 古實 和 弗 的勇士， 擅長拉弓的 路德 人，前進吧！」
JER|46|10|那日是萬軍之主耶和華報仇的日子， 要向敵人報仇。 刀劍必吞吃飽足， 飲血滿足； 因為在北方 幼發拉底河 邊， 有祭物獻給萬軍之主耶和華。
JER|46|11|少女 埃及 啊， 要上 基列 去取乳香； 你雖服用許多藥， 還是徒然，不得治好。
JER|46|12|列國聽見你的羞辱， 遍地滿了你的哀聲； 勇士與勇士彼此相撞， 二人一起跌倒。
JER|46|13|以下是耶和華對 耶利米 先知說的話，論到 巴比倫 王 尼布甲尼撒 要來攻擊 埃及 地。
JER|46|14|你們要在 埃及 傳揚，在 密奪 報告， 在 挪弗 、 答比匿 宣告說： 「要擺好陣勢，預備作戰， 因為刀劍在你四圍施行吞滅。」
JER|46|15|你的壯士為何被掃除呢？ 他們站立不住， 因為耶和華驅逐他們；
JER|46|16|他使多人絆跌，彼此撞倒。 他們說：「起來，讓我們回到自己的同胞、 回到自己的出生地去， 好躲避欺壓的刀劍。」
JER|46|17|他們在那裏稱 埃及 王法老 為 「錯失良機的誇大者」。
JER|46|18|名為萬軍之耶和華的君王說： 我指著我的永生起誓： 「 尼布甲尼撒 來的時候， 必像眾山之中的 他泊 ， 像海邊的 迦密 。」
JER|46|19|住在 埃及 的啊， 要預備被擄時需用的物品； 因為 挪弗 必成為廢墟， 被燒燬，無人居住。
JER|46|20|埃及 是肥美的母牛犢； 但來自北方的牛虻來到了！來到了！
JER|46|21|它的傭兵好像圈裏的肥牛犢， 他們轉身退後， 一齊逃跑，站立不住； 因為他們遭難的日子、 受罰的時刻已經來臨。
JER|46|22|它的聲音好像蛇在滑行。 敵人要成隊而來，如砍伐樹木的人， 手拿斧頭攻擊它。
JER|46|23|雖然它的樹林不易穿過， 敵人卻要砍伐， 因敵人比蝗蟲還多，不可勝數。 這是耶和華說的。
JER|46|24|埃及 必然蒙羞， 被交在北方人的手中。
JER|46|25|萬軍之耶和華－ 以色列 的上帝說：「看哪，我要懲罰 挪 的 亞捫 和法老、 埃及 和它的神明，以及君王，也要懲罰法老和倚靠他的人。
JER|46|26|我要將他們交給尋索其命之人的手和 巴比倫 王 尼布甲尼撒 與他臣僕的手。但 埃及 日後必再有人居住，與從前一樣。這是耶和華說的。」
JER|46|27|我的僕人 雅各 啊，不要懼怕！ 以色列 啊，不要驚惶！ 因我要從遠方拯救你， 從被擄之地拯救你的後裔。 雅各 必回來，得享平靜安逸， 無人令他害怕。
JER|46|28|我的僕人 雅各 啊，不要懼怕！ 因我與你同在。 我要將那些國滅絕淨盡， 就是我趕你去的那些國； 卻不將你滅絕淨盡， 倒要從寬懲治你， 但絕不能不罰你。 這是耶和華說的。
JER|47|1|在法老攻擊 迦薩 之前，耶和華論 非利士 人的話臨到 耶利米 先知。
JER|47|2|耶和華如此說： 看哪，有水從北方漲起，成為漲溢的河， 要淹沒全地和其中所充滿的， 淹沒城和城裏的居民。 人必呼喊， 境內的居民都必哀號。
JER|47|3|一聽見敵人壯馬蹄踏的響聲、 戰車隆隆、車輪轟轟， 為父的手就發軟， 不能回頭看顧兒女。
JER|47|4|因為日子將到， 耶和華必毀滅所有 非利士 人， 剪除 推羅 、 西頓 僅存的幫助者； 他要毀滅 非利士 人、 迦斐託 海島剩餘的人。
JER|47|5|迦薩 成了光禿， 亞實基倫 歸於無有。 平原 中所剩的啊， 你割劃自己，要到幾時呢？
JER|47|6|耶和華的刀劍哪，你要到幾時才止息呢？ 要入鞘，安靜不動。
JER|47|7|耶和華吩咐它攻擊 亞實基倫 和海邊之地， 既已派定它，你 怎能靜止不動呢？
JER|48|1|論 摩押 。 萬軍之耶和華－ 以色列 的上帝如此說： 禍哉， 尼波 ！它要變為廢墟。 基列亭 蒙羞被攻取， 米斯迦 蒙羞被毀壞，
JER|48|2|摩押 不再被稱讚。 有人在 希實本 設計謀害它： 「來吧！我們將它剪除，使它不再成國。」 瑪得緬 哪，你也必靜默無聲； 刀劍必追趕你。
JER|48|3|從 何羅念 有哀號聲： 「荒涼！大毀滅！」
JER|48|4|「 摩押 毀滅了！」 它的孩童哀號，使人聽見。
JER|48|5|人上 魯希坡 隨走隨哭， 因為在 何羅念 的下坡聽見毀滅的哀聲。
JER|48|6|你們要奔逃，自救己命， 使你們的性命如曠野裏的矮樹 。
JER|48|7|你因倚靠自己所做的 和自己的財寶，必被攻取。 基抹 和屬它的祭司、官長也要一同被擄去。
JER|48|8|那行毀滅的要來到各城， 並無一城倖免。 山谷必敗落， 平原必毀壞， 正如耶和華所說的。
JER|48|9|你們要將翅膀給 摩押 ， 使它可以飛去 。 它的城鎮必荒涼， 無人居住。
JER|48|10|懶惰不肯為耶和華做事的，必受詛咒；禁止刀劍不見血的，必受詛咒。
JER|48|11|摩押 自幼年以來常享安逸， 如沉澱未被攪動的酒 ， 沒有從這器皿倒在那器皿， 也未曾被擄掠過。 因此，它的原味尚存， 香氣未變。
JER|48|12|看哪，日子將到，我必差倒酒的到它那裏去，將它倒出來；他們要倒空器皿，打碎罈子。這是耶和華說的。
JER|48|13|摩押 必因 基抹 羞愧，像 以色列 家因倚靠 伯特利 羞愧一樣。
JER|48|14|你們怎麼說： 「我們是勇士，是會打仗的壯士」呢？
JER|48|15|摩押 變為廢墟， 敵人上去佔它的城鎮。 它精良的壯丁都下去遭殺戮； 這是名為萬軍之耶和華的君王說的。
JER|48|16|摩押 的災殃臨近， 災難速速來到。
JER|48|17|凡在它四圍的和認識它名的， 都要為它悲傷，說： 那結實的杖和美好的棍， 竟然折斷了！
JER|48|18|底本 的居民哪， 要從你榮耀的座位上下來， 坐著忍受乾渴； 因毀滅 摩押 的人上來攻擊你， 毀壞了你的堡壘。
JER|48|19|住 亞羅珥 的啊， 要站在道路的邊上觀望， 問逃跑的男人和逃脫的女人說： 「發生了甚麼事呢」？
JER|48|20|摩押 因毀壞蒙羞； 你們要哀號呼喊， 要在 亞嫩 報告： 「 摩押 已成廢墟！」
JER|48|21|審判臨到平原之地的 何倫 、 雅雜 、 米法押 、
JER|48|22|底本 、 尼波 、 伯‧低比拉太音 、
JER|48|23|基列亭 、 伯‧迦末 、 伯‧米恩 、
JER|48|24|加略 、 波斯拉 和 摩押 地遠近所有的城鎮。
JER|48|25|摩押 的角砍斷了，膀臂折斷了。這是耶和華說的。
JER|48|26|你們要使 摩押 沉醉，因它向耶和華誇大。它要在自己所吐之物中打滾，又要被人嗤笑。
JER|48|27|以色列 不是你的笑柄嗎？它難道是在賊中被逮到，使你每逢提到它就搖頭的嗎？
JER|48|28|摩押 的居民哪， 要離開城鎮，住在山崖裏， 像鴿子在峽谷口上搭窩。
JER|48|29|我們聽聞 摩押 人的驕傲， 極其驕傲； 他們自高、自傲、 自我狂妄、居心自大。
JER|48|30|我知道他們的憤怒是虛空的， 他們誇大的話一無所成。 這是耶和華說的。
JER|48|31|因此，我要為 摩押 哀號， 為 摩押 全地呼喊； 人必為 吉珥‧哈列設 人嘆息。
JER|48|32|西比瑪 的葡萄樹啊，我為你哀哭， 甚於 雅謝 人的哀哭。 你的枝子蔓延過海， 直伸到 雅謝海 。 那行毀滅的已經臨到你夏天的果子和葡萄。
JER|48|33|肥田和 摩押 地的歡喜快樂都被奪去， 我使酒池不再流出酒來， 無人踹酒歡呼； 呼喊的聲音不再是歡呼。
JER|48|34|有哀聲從 希實本 達到 以利亞利 ，他們發的哀聲達到 雅雜 ；從 瑣珥 達到 何羅念 ，達到 伊基拉‧施利施亞 ，因為 寧林 的水必然乾涸。
JER|48|35|我必在 摩押 地使那在丘壇獻祭的，和那向他的神明燒香的都滅絕了。這是耶和華說的。
JER|48|36|因此，我的心為 摩押 哀鳴如簫，我的心為 吉珥‧哈列設 人哀哭； 摩押 人所得的財物都毀滅了。
JER|48|37|各人頭上光禿，鬍鬚剪短，手有劃傷，腰束麻布。
JER|48|38|在 摩押 的各房頂上和街市上到處有人哀哭，因我打碎 摩押 ，好像打碎無人喜愛的器皿。這是耶和華說的。
JER|48|39|打得粉碎了！他們要哀號了！ 摩押 要羞愧轉背了！這樣， 摩押 必受四圍的人嗤笑驚駭。
JER|48|40|耶和華如此說： 看哪，仇敵必如鷹展翅快飛， 攻擊 摩押 。
JER|48|41|加略 被攻取，堡壘也被佔據。 到那日， 摩押 的勇士心中疼痛如臨產的婦人。
JER|48|42|摩押 必被毀滅，不再成國， 因它向耶和華誇大。
JER|48|43|摩押 的居民哪， 驚嚇、陷阱、羅網都臨近你。 這是耶和華說的。
JER|48|44|躲過驚嚇的必墜入陷阱， 逃離陷阱的又被羅網纏住， 因我必使懲罰之年臨到 摩押 。 這是耶和華說的。
JER|48|45|逃難的人站在 希實本 的蔭下，筋疲力盡， 因為有火從 希實本 發出， 有火焰出自 西宏 ， 燒盡 摩押 的鬢角和鬧鬨人的頭頂。
JER|48|46|摩押 啊，你有禍了！ 屬 基抹 的百姓滅亡了！ 因你的兒子都被擄去， 你的女兒也被擄去。
JER|48|47|到末後，我卻要使 摩押 被擄的人歸回。 摩押 受審判的話到此為止。 這是耶和華說的。
JER|49|1|論 亞捫 人。 耶和華如此說： 以色列 沒有兒子嗎？ 沒有後嗣嗎？ 米勒公 為何承受 迦得 為業呢？ 屬它的百姓為何住其中的城鎮呢？
JER|49|2|看哪，日子將到，我必使人聽見打仗的喊聲， 攻擊 亞捫 人所住的 拉巴 的喊聲。 拉巴 要成為廢墟， 屬它的鄉鎮 要被火焚燒。 這是耶和華說的。 先前承受 以色列 為業的， 此時 以色列 倒要承受他們為業。 這是耶和華說的。
JER|49|3|希實本 哪，要哀號， 因為 愛 地已成荒地。 拉巴 的鄉鎮哪，要呼喊， 以麻布束腰； 要哭號，在籬笆中往來奔跑； 因 米勒公 和它的祭司、 官長要一同被擄去。
JER|49|4|背道的民 哪， 你為何因有山谷， 因有水流的山谷誇耀呢？ 為何倚靠自己的財寶，說： 「誰能來到我們這裏呢？」
JER|49|5|萬軍之主耶和華說： 看哪，我要使驚嚇從四圍的鄰邦臨到你們； 你們必被趕出， 各人一直往前， 無人收容難民。
JER|49|6|但後來，我卻要使被擄的 亞捫 人歸回。這是耶和華說的。
JER|49|7|論 以東 。 萬軍之耶和華如此說： 提幔 不再有智慧了嗎？ 聰明人的謀略都用盡了嗎？ 他們的智慧盡歸無有了嗎？
JER|49|8|底但 的居民哪，要轉身逃跑， 住在深密處； 因為我懲罰 以掃 的時候， 必使災殃臨到他。
JER|49|9|摘葡萄的若來到你那裏， 豈不留下幾串嗎？ 賊若夜間來到， 豈不是只毀壞他們要毀壞的嗎？
JER|49|10|我卻使 以掃 赤裸， 暴露他的藏身處； 他不能隱藏自己。 他的後裔、弟兄、鄰舍全都滅絕， 他也歸於無有。
JER|49|11|你撇下孤兒，我必保全他們的性命； 你的寡婦可以倚靠我。
JER|49|12|耶和華如此說：「看哪，既然原不該喝那杯的一定要喝，你能免去懲罰嗎？必不能免，一定要喝！
JER|49|13|我指著自己起誓， 波斯拉 必令人驚駭、受羞辱、被詛咒，並且全然荒廢。它所有的城鎮都要永遠成為廢墟。這是耶和華說的。」
JER|49|14|我從耶和華那裏聽見消息， 有使者被差往列國去，說： 「你們要聚集前來攻擊 以東 ， 要起來爭戰。」
JER|49|15|看哪，我使你在列國中為最小， 在世人中被藐視。
JER|49|16|住在山穴中盤據山頂的啊， 你被自己的聲勢與心中的狂傲所蒙蔽； 你雖如大鷹高高搭窩， 我卻要從那裏拉你下來。 這是耶和華說的。
JER|49|17|以東 必令人驚駭；凡經過的人都驚駭，又因它一切的災禍嗤笑。
JER|49|18|耶和華說：它要像 所多瑪 、 蛾摩拉 和鄰近的城鎮一樣傾覆，必無人住在那裏，也無人在其中寄居。
JER|49|19|看哪，就像獅子從 約旦河 邊的叢林上來，攻擊堅固的居所，我要在轉眼之間使 以東 人逃跑，離開這地。我揀選誰，就派誰治理這地。誰能像我呢？誰能召我出庭呢？ 有哪一個牧人能在我面前站得住呢？
JER|49|20|你們要聽耶和華攻擊 以東 所定的計劃和他攻擊 提幔 居民所定的旨意。他們羊群當中微弱的定要被拖走，他們的草場定要變為荒涼。
JER|49|21|因他們仆倒的聲音，地就震動，哀號的聲音傳到 紅海 那裏。
JER|49|22|看哪，仇敵必如大鷹飛起，展開翅膀攻擊 波斯拉 。到那日， 以東 的勇士心中疼痛如臨產的婦人。
JER|49|23|論 大馬士革 。 哈馬 和 亞珥拔 蒙羞， 因為他們聽見兇惡的消息就融化； 焦慮像海浪洶湧，不得平靜。
JER|49|24|大馬士革 發軟，轉身逃跑； 戰兢將它捉住， 痛苦憂愁將它抓住， 如臨產的婦人一樣。
JER|49|25|我所喜樂受稱讚的城， 怎能被撇棄 呢？
JER|49|26|它的壯丁必仆倒在街上， 當那日，戰士全都靜默無聲。 這是萬軍之耶和華說的。
JER|49|27|我必用火點燃 大馬士革 的城牆， 燒滅 便‧哈達 的宮殿。
JER|49|28|論 巴比倫 王 尼布甲尼撒 所攻打的 基達 和 夏瑣 諸國。 耶和華如此說： 迦勒底 人哪，起來上 基達 去， 毀滅東方人。
JER|49|29|人要奪去他們的帳棚和羊群， 人要帶走他們的幔子、一切器皿，和駱駝，佔為己有。 人向他們喊著說： 四圍都有驚嚇。
JER|49|30|夏瑣 的居民哪，要逃奔遠方， 住在深遠之處； 因為 巴比倫 王 尼布甲尼撒 設計謀害你們， 起意攻擊你們。 這是耶和華說的。
JER|49|31|迦勒底 人哪，起來！ 上到安逸無慮的國民那裏去， 他們是無門無閂、單獨居住的。 這是耶和華說的。
JER|49|32|他們的駱駝必成為掠物， 他們眾多的牲畜必成為擄物。 我要將剃鬢髮的人分散四方 ， 使災殃從四圍臨到他們。 這是耶和華說的。
JER|49|33|夏瑣 必成為野狗的住處， 永遠荒廢； 無人住在那裏， 也無人在其中寄居。
JER|49|34|猶大 王 西底家 登基的時候，耶和華論 以攔 的話臨到 耶利米 先知，說：
JER|49|35|「萬軍之耶和華如此說：看哪，我必折斷 以攔 人的弓，那是他們戰鬥的主力。
JER|49|36|我要使風從天的四方颳來，臨到 以攔 ，將他們分散四方。 以攔 被趕散的人沒有一國不到的。
JER|49|37|我必使 以攔 人在仇敵和尋索其命的人面前驚惶；我也必使災禍，就是我的烈怒臨到他們，又必使刀劍追殺他們，直到將他們滅盡。這是耶和華說的。
JER|49|38|我要在 以攔 設立我的寶座，在那裏除滅君王和官長。這是耶和華說的。
JER|49|39|「到末後，我卻要使被擄的 以攔 人歸回。這是耶和華說的。」
JER|50|1|以下是耶和華藉 耶利米 先知論 巴比倫 和 迦勒底 人之地所說的話。
JER|50|2|你們要在萬國中傳揚，宣告， 豎立大旗； 要宣告，不可隱瞞，說： 「 巴比倫 被攻取， 彼勒 蒙羞， 米羅達 驚惶。 巴比倫 的神像都蒙羞， 它的偶像都驚惶。」
JER|50|3|因有一國從北方上來攻擊它，使它的地荒涼，無人居住，連人帶牲畜都逃走了。
JER|50|4|在那日、在那時， 以色列 人要和 猶大 人同來，隨走隨哭，尋求耶和華－他們的上帝。這是耶和華說的。
JER|50|5|他們要問到 錫安 之路，又面向那裏，說：「來吧，他們要 在永不被遺忘的約中與耶和華聯合。」
JER|50|6|我的百姓成了失喪的羊，牧人使他們走迷了路，轉入叢山之間。他們從大山走到小山，竟忘了自己安歇之處。
JER|50|7|凡遇見他們的，就把他們吞滅。敵人說：「我們不算有罪；因他們得罪了那可作真正 居所的耶和華，就是他們祖先所仰望的耶和華。」
JER|50|8|「你們要逃離 巴比倫 ，要離開 迦勒底 人之地，像走在羊群前面的公山羊。
JER|50|9|看哪，因我必激起大國聯盟，帶領他們從北方來攻擊 巴比倫 ，他們要擺陣攻擊它，它必在那裏被攻取。他們的箭好像善射 勇士的箭，絕不徒然返回。
JER|50|10|迦勒底 要成為掠物，凡擄掠它的都必心滿意足。這是耶和華說的。」
JER|50|11|搶奪我產業的啊， 你們因歡喜快樂， 像踹穀 嬉戲的母牛犢， 又像發嘶聲的壯馬。
JER|50|12|你們的母親極其抱愧， 生你們的必然蒙羞。 看哪，她要列在諸國之末， 成為曠野、旱地、沙漠；
JER|50|13|因耶和華的憤怒， 巴比倫 必無人居住， 全然荒涼， 凡經過的都要受驚駭， 又因它所遭的災殃嗤笑。
JER|50|14|所有拉弓的啊，要在 巴比倫 的四圍擺陣， 射箭攻擊它， 不用愛惜箭枝， 因為它得罪了耶和華。
JER|50|15|要在它四圍吶喊： 「它已經投降， 堡壘坍塌了， 城牆拆毀了！」 這是耶和華所報的仇。 你們要向它報仇； 它怎樣待人，你們也要怎樣待它。
JER|50|16|你們要將 巴比倫 撒種的 和收割時拿鐮刀的全都剪除。 他們各人因躲避欺壓的刀劍， 必歸回本族，逃到本土。
JER|50|17|以色列 是打散的羊，被獅子趕散。首先是 亞述 王將他吞滅，末後是 巴比倫 王 尼布甲尼撒 折斷他的骨頭。
JER|50|18|所以萬軍之耶和華－ 以色列 的上帝如此說：「看哪，我必懲罰 巴比倫 王和他的地，像我從前懲罰 亞述 王一樣。
JER|50|19|我必領 以色列 回他自己的草場，他要在 迦密 和 巴珊 吃草，又在 以法蓮 山上和 基列 境內得以飽足。
JER|50|20|在那日、在那時，你尋找 以色列 的罪孽，一無所有；尋找 猶大 的罪惡，也無所得；因為我所留下的人，我必赦免。這是耶和華說的。」
JER|50|21|你要上去攻擊 米拉大翁 之地， 又攻擊 比割 的居民。 將他們追殺滅盡， 照我所吩咐你的一切去做。 這是耶和華說的。
JER|50|22|境內有打仗和大毀滅的響聲。
JER|50|23|全地的大錘竟然砍斷破壞！ 巴比倫 在列國中竟然荒涼！
JER|50|24|巴比倫 哪，我為你設下羅網， 你被纏住，竟不自覺。 你被尋著，也被捉住， 因為你對抗耶和華。
JER|50|25|耶和華已經打開軍械庫， 拿出他惱恨的兵器； 這是萬軍之主耶和華 在 迦勒底 人之地要做的事。
JER|50|26|你們要從極遠的邊界前來攻擊它 ， 要開它的倉廩， 將它堆起如高堆， 毀滅淨盡，絲毫不留。
JER|50|27|要殺它一切的牛犢， 使牠們下去遭殺戮。 他們有禍了， 因為他們的日子，就是他們受罰的時刻已經來到。
JER|50|28|從 巴比倫 之地逃出來的難民，在 錫安 揚聲宣告耶和華－我們的上帝要報仇，為他的聖殿報仇。
JER|50|29|你們要招集一切弓箭手來攻擊 巴比倫 ，在 巴比倫 四圍安營，不容一人逃脫。要照著它所做的報應它；它怎樣待人，你們也要怎樣待它，因為它向耶和華－ 以色列 的聖者狂傲。
JER|50|30|所以它的壯丁必仆倒在街上。當那日，它的士兵全都靜默無聲。這是耶和華說的。
JER|50|31|「看哪，你這狂傲的啊，我與你為敵， 因為你的日子， 我懲罰你的時刻已經來到。 這是萬軍之主耶和華說的。
JER|50|32|狂傲的必絆跌仆倒，無人扶起。 我必用火點燃他的城鎮， 將他四圍所有的盡行燒滅。」
JER|50|33|萬軍之耶和華如此說：「 以色列 人和 猶大 人一同受欺壓；凡擄掠他們的都緊緊抓住他們，不肯釋放。
JER|50|34|他們的救贖主大有能力，萬軍之耶和華是他的名。他必定為他們伸冤，使全地得享平靜；他卻要攪擾 巴比倫 的居民。」
JER|50|35|有刀劍臨到 迦勒底 人和 巴比倫 的居民， 臨到它的領袖與智慧人。 這是耶和華說的。
JER|50|36|有刀劍臨到矜誇的人， 他們就變為愚昧； 有刀劍臨到它的勇士， 他們就驚惶。
JER|50|37|有刀劍臨到它的馬匹、戰車， 和其中混居的各族， 他們變成與婦女一樣； 有刀劍臨到它的寶物， 寶物就被搶奪。
JER|50|38|有乾旱 臨到它的眾水， 它們就必乾涸； 因為這是雕刻偶像之地， 人因偶像顛狂 。
JER|50|39|所以野獸和土狼必住在那裏，鴕鳥也住在其中，永遠無人居住，世世代代無人定居。
JER|50|40|巴比倫 要像上帝所傾覆的 所多瑪 、 蛾摩拉 和鄰近的城鎮一樣，必無人住在那裏，也無人在其中寄居。這是耶和華說的。
JER|50|41|看哪，有一民族從北方而來， 有一大國和許多君王被激起，從地極來到。
JER|50|42|他們拿弓和槍， 性情殘忍，毫不留情； 他們的聲音像海浪澎湃。 巴比倫 啊， 他們騎著馬， 如上戰場的人擺列隊伍， 要攻擊你。
JER|50|43|巴比倫 王聽見他們的風聲， 手就發軟， 痛苦將他抓住， 彷彿臨產的婦人疼痛一般。
JER|50|44|「看哪，就像獅子從 約旦河 邊的叢林上來，攻擊堅固的居所，我要在轉眼之間使 迦勒底 人逃跑，離開這地。我揀選誰，就派誰治理這地。誰能像我呢？誰能召我出庭呢？有哪一個牧人能在我面前站得住呢？
JER|50|45|你們要聽耶和華攻擊 巴比倫 所定的計劃和他攻擊 迦勒底 人之地所定的旨意。他們羊群當中微弱的定要被拖走，他們的草場定要變為荒涼。
JER|50|46|因 巴比倫 被攻下的聲音，地就震動，人在列國都聽見呼喊的聲音。」
JER|51|1|耶和華如此說： 看哪，我必颳起毀滅的風， 攻擊 巴比倫 和住在 立加米 的人。
JER|51|2|我要差陌生人 來到 巴比倫 ， 他們要簸揚它，使它的地空無一物。 在它遭禍的日子， 他們要四圍攻擊它。
JER|51|3|不要叫拉弓的拉弓， 不要叫他佩戴盔甲 ； 不要憐惜 巴比倫 的壯丁， 要滅盡它的全軍。
JER|51|4|他們必在 迦勒底 人之地被殺仆倒， 在 巴比倫 的街市上被刺透。
JER|51|5|以色列 和 猶大 境內雖然充滿違背 以色列 聖者的罪， 卻沒有被他的上帝－萬軍之耶和華所遺棄。
JER|51|6|你們要奔逃，離開 巴比倫 ， 各救自己的性命！ 不要陷在它的罪孽中一同滅亡， 因為這是耶和華報仇的時刻， 他必向 巴比倫 施行報應。
JER|51|7|巴比倫 素來是耶和華手中的金杯， 使全地沉醉， 列國喝了它的酒就顛狂。
JER|51|8|巴比倫 忽然傾覆毀壞； 要為它哀號， 拿乳香來止它的疼痛， 或者可以治好。
JER|51|9|我們想醫治 巴比倫 ， 它卻未獲痊癒。 離開它吧！讓我們各人歸回本國， 因為它受的審判通於上天，達到穹蒼。
JER|51|10|耶和華已經彰顯出我們的義。 來吧！我們要在 錫安 傳揚耶和華－我們上帝的作為。
JER|51|11|你們要磨尖箭頭， 抓住盾牌。 論到 巴比倫 ，耶和華定意要毀滅它，所以激起 瑪代 君王的心；這是耶和華報仇，為他的聖殿報仇。
JER|51|12|你們要豎立大旗， 攻擊 巴比倫 的城牆； 要堅固瞭望臺， 派定守望的設下埋伏； 因為耶和華指著 巴比倫 居民所說的， 他不但這樣定意，也已成就。
JER|51|13|住在眾水之上多有財寶的啊， 你的結局已到！ 你貪婪之量已滿盈 ！
JER|51|14|萬軍之耶和華指著自己起誓說： 我必使人遍滿各處像蝗蟲一樣， 他們必吶喊攻擊你。
JER|51|15|耶和華以能力創造大地， 以智慧建立世界， 以聰明鋪張穹蒼。
JER|51|16|他一出聲，天上就有眾水澎湃； 他使雲霧從地極上騰， 造電隨雨而閃， 從倉庫中吹出風來。
JER|51|17|人人都如同畜牲，毫無知識； 銀匠都因偶像羞愧， 他所鑄的偶像本為虛假， 它們裏面並無氣息。
JER|51|18|它們都是虛無的， 是迷惑人的東西， 到它們受罰的時刻必被除滅。
JER|51|19|雅各 所得的福分不是這樣， 因主 是那創造萬有的， 以色列 是他產業的支派， 萬軍之耶和華是他的名。
JER|51|20|你是我爭戰的斧子和打仗的兵器。 我要用你打碎列邦， 毀滅列國；
JER|51|21|用你打碎馬和騎馬的， 打碎戰車和坐在其上的；
JER|51|22|用你打碎男人和女人， 打碎老人和少年， 打碎壯丁和少女；
JER|51|23|用你打碎牧人和他的羊群， 打碎農夫和他的一對耕牛， 打碎省長和官員。
JER|51|24|我必在你們眼前報復 巴比倫 人和 迦勒底 居民在 錫安 所做的一切惡事。這是耶和華說的。
JER|51|25|行毀滅的山，看哪，我與你為敵， 你毀滅全地， 我必伸手攻擊你， 將你從山巖滾下去， 使你成為燒燬了的山。 這是耶和華說的。
JER|51|26|人必不從你那裏取石頭為房角石， 也不取石頭來作根基， 因為你必永遠荒廢。 這是耶和華說的。
JER|51|27|你們要在境內豎立大旗， 在列邦中吹角， 使列邦預備攻擊 巴比倫 。 要招集 亞拉臘 、 米尼 、 亞實基拿 各國前來攻擊它， 派將軍攻擊它， 使馬匹上來如粗暴的蝗蟲；
JER|51|28|使列邦和 瑪代 君王，省長和官員， 他們所管的全地，都預備攻擊它。
JER|51|29|地必震動而移轉； 因耶和華向 巴比倫 旨意已確定， 要使 巴比倫 土地荒涼，無人居住。
JER|51|30|巴比倫 的勇士停止爭戰， 躲在堡壘之中。 他們的力氣耗盡， 他們變成與婦女一樣。 巴比倫 的住處焚燒， 門閂都折斷了。
JER|51|31|通報的彼此相遇， 送信的彼此相遇， 報告 巴比倫 王， 城的四方都被攻下了，
JER|51|32|渡口被佔據了， 蘆葦被火焚燒， 戰士都驚慌。
JER|51|33|萬軍之耶和華－ 以色列 的上帝如此說： 巴比倫 好像踹穀的禾場； 再過片時，它收割的時候就到了。
JER|51|34|巴比倫 王 尼布甲尼撒 吞滅我，壓碎我， 使我成為空器皿。 他如大魚將我吞下， 以我的美物充滿他的肚腹， 又把我趕出去。
JER|51|35|錫安 的居民要說： 願我和我骨肉之親所受的殘暴 歸給 巴比倫 。 耶路撒冷 人要說： 願我們所流的血 歸給 迦勒底 的居民。
JER|51|36|所以，耶和華如此說： 看哪，我必為你伸冤，為你報仇； 我必使 巴比倫 的海枯竭， 使它的泉源乾涸。
JER|51|37|巴比倫 必成為廢墟， 為野狗的住處， 令人驚駭、嗤笑， 並且無人居住。
JER|51|38|他們要像少壯獅子一同咆哮， 像小獅子吼叫。
JER|51|39|他們食慾一來的時候， 我必為他們擺設酒席， 使他們沉醉，好叫他們快樂； 他們睡了長覺，永不醒起。 這是耶和華說的。
JER|51|40|我必使他們像羔羊、 像公綿羊和公山羊被牽去宰殺。
JER|51|41|示沙克 竟然被攻取！ 全地所稱讚的被佔據！ 巴比倫 在列國中竟然變為荒涼！
JER|51|42|海水漲起，漫過 巴比倫 ； 澎湃的海浪遮蓋了它。
JER|51|43|它的城鎮變廢墟， 地變乾旱，成為沙漠， 成為無人居住、 無人經過之地。
JER|51|44|我要懲罰 巴比倫 的 彼勒 ， 使它吐出所吞之物。 列國必不再流歸到它那裏， 巴比倫 的城牆也必坍塌。
JER|51|45|我的子民哪，你們要離開 巴比倫 ！ 各人逃命，躲避耶和華的烈怒。
JER|51|46|不要因境內所聽見的風聲 心驚膽怯或懼怕； 因為這年有風聲傳來， 那年也有風聲傳來； 境內有殘暴的事， 官長攻擊官長。
JER|51|47|所以，看哪，日子將到， 我必懲罰 巴比倫 雕刻的偶像。 它的全地必然抱愧， 它被殺的人必仆倒在其上。
JER|51|48|那時，天地和其中所有的， 必因 巴比倫 歡呼， 因為行毀滅的要從北方來到它那裏。 這是耶和華說的。
JER|51|49|巴比倫 要因 以色列 被殺的人而仆倒， 正如全地被刺殺的人是因 巴比倫 仆倒一般。
JER|51|50|你們躲避刀劍的要快走， 不要站住！ 要在遠方懷念耶和華， 心中追想 耶路撒冷 。
JER|51|51|我們聽見辱罵就蒙羞，滿面慚愧， 因為外邦人進入耶和華殿的聖所。
JER|51|52|所以，看哪，日子將到， 我必懲罰 巴比倫 雕刻的偶像， 在全境內到處都有刺傷的人在呻吟。 這是耶和華說的。
JER|51|53|巴比倫 雖升到天上， 雖使它堅固的高處更堅固， 我也要差毀滅者到它那裏。 這是耶和華說的。
JER|51|54|有哀號的聲音從 巴比倫 出來， 有大毀滅從 迦勒底 人之地而來。
JER|51|55|耶和華使 巴比倫 變為廢墟， 使其中喧嘩的大聲滅絕。 仇敵彷彿眾水， 波浪澎湃，發出響聲；
JER|51|56|這是行毀滅的臨到 巴比倫 。 巴比倫 的勇士被捉住， 他們的弓折斷了； 因為耶和華是施行報應的上帝， 他必施行報應。
JER|51|57|我必使 巴比倫 的領袖、 智慧人、省長、官員和勇士都喝醉， 使他們永遠沉睡，不再醒起。 這是名為萬軍之耶和華的君王說的。
JER|51|58|萬軍之耶和華如此說： 巴比倫 寬闊的城牆要夷為平地， 它高大的城門必被火焚燒。 萬民所勞碌的必致虛空， 萬族所勞碌的被火焚燒， 他們都必困乏。
JER|51|59|猶大 王 西底家 在位第四年， 瑪西雅 的孫子， 尼利亞 的兒子 西萊雅 與王同去 巴比倫 ， 西萊雅 是王宮的大臣， 耶利米 先知有話吩咐他。
JER|51|60|耶利米 把一切要臨到 巴比倫 的災禍，就是論到 巴比倫 的這一切話，寫在一書卷上。
JER|51|61|耶利米 對 西萊雅 說：「你到了 巴比倫 ，務要宣讀這一切話，
JER|51|62|說：『耶和華啊，你曾論到這地方說：要剪除它，不再有人與牲畜居住此地，必永遠荒涼。』
JER|51|63|你讀完這書卷，就要把一塊石頭拴在其上，投入 幼發拉底河 中，
JER|51|64|說：『 巴比倫 因耶和華所要降與它的災禍，必如此沉下去，不再浮起來，百姓也必困乏。』」 耶利米 的話到此為止。
JER|52|1|西底家 登基的時候年二十一歲，在 耶路撒冷 作王十一年。他母親名叫 哈慕她 ，是 立拿 人 耶利米 的女兒。
JER|52|2|西底家 行耶和華眼中看為惡的事，像 約雅敬 所做的一切。
JER|52|3|因此，耶和華向 耶路撒冷 和 猶大 發怒，以致把他們從自己面前趕出去。 西底家 背叛 巴比倫 王，
JER|52|4|他作王第九年十月初十， 巴比倫 王 尼布甲尼撒 率領全軍前來攻擊 耶路撒冷 ，對著城安營，四圍築堡壘攻城，
JER|52|5|城被圍困，直到 西底家 王十一年。
JER|52|6|四月初九，城裏的饑荒非常嚴重，當地的百姓都沒有糧食。
JER|52|7|城被攻破，士兵全都在夜間從靠近王園兩城牆中間的門逃跑出城； 迦勒底 人正在四圍攻城，他們就往 亞拉巴 逃去。
JER|52|8|迦勒底 的軍隊追趕 西底家 王，在 耶利哥 的平原追上他。他的全軍都離開他潰散了。
JER|52|9|迦勒底 人就拿住王，帶他到 哈馬 地 利比拉 的 巴比倫 王那裏； 巴比倫 王就判他的罪。
JER|52|10|巴比倫 王在 西底家 眼前殺了他的兒女，又在 利比拉 殺了 猶大 全體的官長，
JER|52|11|並且挖了 西底家 的眼睛，用銅鏈鎖著他，帶到 巴比倫 去，將他囚在監裏，直到他死的日子。
JER|52|12|巴比倫 王 尼布甲尼撒 十九年五月初十，在 巴比倫 王面前侍立的 尼布撒拉旦 護衛長進入 耶路撒冷 ，
JER|52|13|他焚燒了耶和華的殿、王宮和 耶路撒冷 的房屋；用火焚燒所有大戶人家的房屋。
JER|52|14|跟隨護衛長的 迦勒底 全軍拆毀了 耶路撒冷 四圍的城牆。
JER|52|15|那時 尼布撒拉旦 護衛長將百姓中最窮的和城裏所剩下的百姓，並那些投降 巴比倫 王的人，以及剩下的工匠，都擄去了。
JER|52|16|但 尼布撒拉旦 護衛長留下一些當地最窮的人，叫他們修整葡萄園，耕種田地。
JER|52|17|耶和華殿的銅柱並殿內的盆座和銅海， 迦勒底 人都打碎了，把那些銅運到 巴比倫 去；
JER|52|18|他們又帶走鍋、鏟子、鉗子、盤子、勺子，和供奉用的一切銅器；
JER|52|19|杯、火盆、碗、鍋、燈臺、勺子、酒杯，無論金的銀的，護衛長都帶走了；
JER|52|20|還有 所羅門 為耶和華殿所造的兩根柱子、一面銅海，並座下的十二隻銅牛，這些器皿的銅多得無法可秤。
JER|52|21|至於柱子，這一根柱子高十八肘，厚四指，周圍十二肘，中間是空的；
JER|52|22|柱上有銅頂，每個銅頂高五肘；銅頂的周圍有網子和石榴，也都是銅的。另一根柱子與此相同，也有石榴。
JER|52|23|柱子四面有九十六個石榴，在網子周圍，總共有一百個石榴。
JER|52|24|護衛長拿住 西萊雅 大祭司、 西番亞 副祭司和門口的三個守衛，
JER|52|25|又從城中拿住一個管理士兵的官 ，並在城裏找到王面前的七個親信，和召募當地百姓之將軍的書記官，以及在城中找到的六十個當地百姓。
JER|52|26|尼布撒拉旦 護衛長把這些人帶到 利比拉 的 巴比倫 王那裏。
JER|52|27|巴比倫 王擊殺他們，在 哈馬 地的 利比拉 把他們處死。這樣， 猶大 人就被擄去離開本地。
JER|52|28|這是 尼布甲尼撒 所擄百姓的數目：他在位第七年擄去 猶大 人三千零二十三人；
JER|52|29|尼布甲尼撒 十八年從 耶路撒冷 擄去八百三十二人；
JER|52|30|尼布甲尼撒 二十三年， 尼布撒拉旦 護衛長擄去 猶大 人七百四十五人；共有四千六百人。
JER|52|31|巴比倫 王 以未‧米羅達 作王的元年，就是 猶大 王 約雅斤 被擄後三十七年十二月二十五日，他使 猶大 王 約雅斤 抬起頭來，提他出監，
JER|52|32|對他說好話，使他的位高過與他一同被擄、在 巴比倫 眾王的位；
JER|52|33|又給他脫了囚服，使他終身常在 巴比倫 王面前吃飯。
JER|52|34|巴比倫 王賜給他日常需用的食物，日日一份，終身都是這樣，直到他死的日子。
LAM|1|1|唉！先前人口稠密的城市， 現在為何獨坐！ 先前在列國中為大的， 現在竟如寡婦！ 先前在各省中為王后的， 現在竟成為服苦役的人！
LAM|1|2|她 夜間痛哭，淚流滿頰， 在所有親愛的人中，找不到一個安慰她的。 她的朋友都以詭詐待她， 成為她的仇敵。
LAM|1|3|猶大 被擄， 遭遇苦難，多服勞役。 她住在列國中，得不著安息； 追逼她的在狹窄之地追上她。
LAM|1|4|錫安 的道路因無人前來過節就哀傷， 她的城門荒涼， 祭司嘆息， 少女悲傷； 她自己充滿痛苦。
LAM|1|5|她的敵人作主， 她的仇敵亨通； 耶和華因她過犯多而使她受苦， 她的孩童在敵人面前去作俘虜。
LAM|1|6|錫安 的威榮全都失去。 她的領袖如找不著草場的鹿， 在追趕的人面前無力行走。
LAM|1|7|耶路撒冷 在困苦窘迫之時， 就追想古時一切的榮華。 她的百姓落在敵人手中，無人幫助； 敵人看見，就因她的毀滅嗤笑。
LAM|1|8|耶路撒冷 犯了大罪， 因此成為不潔淨； 素來尊敬她的，見她裸露就都藐視她， 她自己也嘆息退後。
LAM|1|9|她的污穢是在下襬上； 她未曾思想自己的結局， 她的敗落令人驚詫， 無人安慰她。 「耶和華啊，求你看顧我的苦難， 因為仇敵強大。」
LAM|1|10|敵人伸手奪取她的一切貴重物品； 她眼見列國侵入她的聖所， 你曾吩咐他們不可進入你的集會。
LAM|1|11|她的百姓都嘆息，尋求食物； 他們用貴重物品換取糧食，要救性命。 「耶和華啊，求你觀看， 留意我多麼卑微。」
LAM|1|12|所有過路的人哪，願這事不要發生在你們身上 。 你們要留意觀看， 有像這樣臨到我的痛苦沒有？ 耶和華在他發烈怒的日子使我受苦。
LAM|1|13|他從高處降火進入我的骨頭， 剋制了我； 他張開網，絆我的腳， 使我退後， 又令我終日淒涼發昏。
LAM|1|14|他用手綁我罪過的軛， 捲繞著加在我頸項上； 他使我力量衰敗。 主將我交在我不能抵擋的人手中。
LAM|1|15|主棄絕我們當中所有的勇士， 聚集會眾攻擊我， 要壓碎我的年輕人。 主踹下少女 猶大 ， 在醡酒池中。
LAM|1|16|我因這些事哭泣， 眼淚汪汪； 因為那安慰我、使我重新得力的， 離我甚遠。 我的兒女孤苦， 因為仇敵得勝了。
LAM|1|17|錫安 伸出雙手，卻無人安慰。 論到 雅各 ，耶和華已經出令， 使四圍的人作他的仇敵； 耶路撒冷 在他們中間成為不潔淨。
LAM|1|18|耶和華是公義的！ 我違背了他的命令。 萬民哪，請聽， 來看我的痛苦； 我的少女和壯丁都被擄去。
LAM|1|19|我招呼我所親愛的， 他們卻欺騙了我。 我的祭司和長老尋找食物，要救性命的時候， 就在城中斷了氣。
LAM|1|20|耶和華啊，求你觀看， 因為我在急難中； 我的心腸煩亂， 我心在我裏面翻轉， 因我大大背逆。 在外，刀劍使人喪亡； 在家，猶如死亡。
LAM|1|21|有人聽見我嘆息 ， 卻無人安慰我！ 我所有的仇敵聽見我的患難就喜樂， 因這是你所做的。 你使你所宣告的日子來臨， 願他們像我一樣。
LAM|1|22|願他們的惡行都呈現在你面前； 你怎樣因我一切的罪過待我， 求你也照樣待他們； 因我嘆息甚多，心中發昏。
LAM|2|1|唉！主竟發怒，使黑雲遮蔽 錫安 ！ 他將 以色列 的華美從天扔在地上， 在他發怒的日子並不顧念自己的腳凳。
LAM|2|2|主吞滅 雅各 一切的住處，並不顧惜。 他發怒傾覆 猶大 的堡壘， 將它們夷為平地， 凌辱這國與她的領袖。
LAM|2|3|他發烈怒，砍斷 以色列 一切的角， 在仇敵面前收回右手。 他將 雅各 燒燬，如火焰四圍吞滅。
LAM|2|4|他張弓好像仇敵， 他站立舉起右手， 如同敵人殺戮我們眼目所喜愛的。 他在 錫安 的帳棚 傾倒憤怒，如火一般。
LAM|2|5|主如仇敵吞滅 以色列 ， 吞滅它一切的宮殿， 毀壞境內的堡壘； 在 猶大 加添悲傷和哭號。
LAM|2|6|他摧毀自己的帳幕如摧毀園子， 毀壞自己的會幕。 耶和華使節慶和安息日在 錫安 盡被遺忘， 又在極其憤怒中厭棄君王與祭司。
LAM|2|7|耶和華撇棄自己的祭壇， 憎惡自己的聖所， 把宮殿的牆交給仇敵。 他們在耶和華的殿中喧嚷， 如在節慶之日一樣。
LAM|2|8|耶和華定意拆毀 錫安 的城牆； 他拉了準繩， 不將手收回，定要毀滅。 他使城郭和城牆都悲哀， 一同衰敗。
LAM|2|9|錫安 的門陷入地裏， 主毀壞，折斷她的門閂。 她的君王和官長都置身列國中，沒有律法； 她的先知也不再從耶和華領受異象。
LAM|2|10|錫安 的長老坐在地上，默默無聲； 他們揚起塵土落在頭上，腰束麻布； 耶路撒冷 的少女垂頭至地。
LAM|2|11|我的眼睛流淚，以致失明； 我的心腸煩亂，肝膽落地， 都因我的百姓 遭毀滅， 又因孩童和吃奶的在城內的廣場上昏厥。
LAM|2|12|他們如受傷的人在城內廣場上昏厥， 在母親的懷裏將要喪命時， 就對母親說：「餅和酒在哪裏呢？」
LAM|2|13|耶路撒冷 啊，我可用甚麼向你證明 呢？ 我可用甚麼與你相比呢？ 少女 錫安 哪，我拿甚麼和你比較，好安慰你呢？ 因你的裂傷大如海； 誰能醫治你呢？
LAM|2|14|你的先知為你看見虛假和粉飾的異象， 並未揭露你的罪孽， 使你被擄的歸回； 卻傳給你虛假與誤導人的默示。
LAM|2|15|凡過路的都向你拍掌。 他們向 耶路撒冷 嗤笑，搖頭： 「這就是人稱為全美的、 稱為全地所喜悅的城嗎？」
LAM|2|16|你所有的仇敵 張口來攻擊你； 他們嗤笑，切齒，說： 「我們把她吞滅了， 這是我們所盼望的日子！ 我們終於等到了，親眼看見了！」
LAM|2|17|耶和華成就了他所定的， 應驗了他古時所命定的。 他傾覆，並不顧惜， 他使仇敵向你誇耀， 使你敵人的角高舉。
LAM|2|18|他們的心哀求主。 錫安 的城牆啊， 願你日夜淚流如河，不讓自己休息， 你眼中的瞳人也不歇息。
LAM|2|19|夜間每逢時辰開始，要起來呼喊， 在主面前傾心吐意如水。 你的孩童在街頭上挨餓昏厥， 你要為他們的性命向主舉手。
LAM|2|20|耶和華啊，求你觀看， 留意你向誰這樣行。 婦人豈可吃自己所生、所撫育的嬰孩嗎？ 祭司和先知豈可在主的聖所中被殺嗎？
LAM|2|21|年輕人和老年人躺臥在街上， 我的少女和壯丁都倒在刀下。 你在發怒的日子殺了他們， 你殺戮，並不顧惜。
LAM|2|22|你從四圍招聚使我驚嚇的人， 像在節慶的日子一樣。 耶和華發怒的日子， 無人逃脫，無人生還。 我所撫育養大的， 仇敵都殺盡了。
LAM|3|1|因耶和華憤怒的杖， 我是遭遇困苦的人。
LAM|3|2|他驅趕我走入黑暗， 沒有光明。
LAM|3|3|他反手攻擊我， 終日不停。
LAM|3|4|他使我皮肉枯乾， 折斷我的骨頭。
LAM|3|5|他築壘攻擊我， 以苦楚和艱難圍困我；
LAM|3|6|使我住在幽暗之處， 像死了許久的人一樣。
LAM|3|7|他圍住我，使我無法脫身； 他使我的銅鏈沉重。
LAM|3|8|儘管我哀號求救， 他仍攔阻我的禱告。
LAM|3|9|他用鑿過的石頭擋住我的道路， 使我的路徑彎曲。
LAM|3|10|他向我如埋伏的熊， 如在隱密處的獅子。
LAM|3|11|他使我轉離正路， 把我撕碎 ，使我淒涼。
LAM|3|12|他拉弓，命我站立， 作為箭靶；
LAM|3|13|把箭袋中的箭 射入我的肺腑。
LAM|3|14|我成了全體百姓的笑柄， 成了他們終日的歌曲。
LAM|3|15|他使我受盡苦楚， 飽食茵蔯；
LAM|3|16|用沙石磨斷我的牙， 以灰塵覆蓋我。
LAM|3|17|你使我遠離平安， 我忘了何為福樂。
LAM|3|18|於是我說：「我的力量衰敗， 在耶和華那裏我毫無指望！」
LAM|3|19|求你記得我的困苦和流離， 它如茵蔯和苦膽一般；
LAM|3|20|我心想念這些， 就在我裏面憂悶 。
LAM|3|21|但我的心回轉過來， 因此就有指望；
LAM|3|22|因耶和華的慈愛，我們不致滅絕 ， 因他的憐憫永不斷絕，
LAM|3|23|每早晨，這些都是新的； 你的信實極其廣大！
LAM|3|24|我心裏說：「耶和華是我的福分， 因此，我要仰望他。」
LAM|3|25|凡等候耶和華，心裏尋求他的， 耶和華必施恩給他。
LAM|3|26|人仰望耶和華， 安靜等候他的救恩， 這是好的。
LAM|3|27|人在年輕時負軛， 這是好的。
LAM|3|28|他當安靜獨坐， 因為這是耶和華加在他身上的。
LAM|3|29|讓他臉伏於地 吧！ 或者還會有指望。
LAM|3|30|讓人打他耳光， 使他飽受凌辱吧！
LAM|3|31|主必不永遠撇棄，
LAM|3|32|他雖使人憂愁， 還要照他豐盛的慈愛施憐憫；
LAM|3|33|他並不存心要人受苦， 令世人憂愁。
LAM|3|34|把世上所有的囚犯 踹在腳下，
LAM|3|35|在至高者面前 扭曲人的公正，
LAM|3|36|在人的訴訟上 顛倒是非， 這都是主看不中的。
LAM|3|37|若非主發命令， 誰能說了就成呢？
LAM|3|38|是禍，是福， 不都出於至高者的口嗎？
LAM|3|39|人都有自己的罪， 活人有甚麼好發怨言的呢？
LAM|3|40|讓我們省察，檢討自己的行為， 歸向耶和華吧！
LAM|3|41|讓我們獻上我們的心， 向天上的上帝舉手！
LAM|3|42|我們犯罪悖逆， 你並未赦免。
LAM|3|43|你渾身是怒氣，追趕我們； 你施行殺戮，並不顧惜。
LAM|3|44|你以密雲圍著自己， 禱告不能穿透。
LAM|3|45|你使我們在萬民中 成為污物和垃圾。
LAM|3|46|我們所有的仇敵 張口來攻擊我們；
LAM|3|47|驚嚇和陷阱臨到我們， 殘害和毀滅也臨到我們。
LAM|3|48|因我百姓 遭毀滅， 我的眼睛淚流成河。
LAM|3|49|我的眼睛流淚不停， 流淚不止，
LAM|3|50|直等到耶和華垂顧， 從天上觀看。
LAM|3|51|為我城中的百姓 ， 我眼所見的使我心痛。
LAM|3|52|無故與我為敵的追逼我， 像追捕雀鳥一樣。
LAM|3|53|他們要在坑中了結我的性命， 丟石頭在我身上。
LAM|3|54|眾水淹沒我的頭， 我說：「我沒命了！」
LAM|3|55|耶和華啊， 在極深的地府裏，我求告你的名。
LAM|3|56|我的聲音你聽見了， 求你不要掩耳不聽 我的呼聲，我的求救。
LAM|3|57|我求告你的時候， 你臨近我，說：「不要懼怕！」
LAM|3|58|主啊，你為我伸冤， 你救贖了我的命。
LAM|3|59|耶和華啊，你已看見我的委屈， 求你為我主持正義。
LAM|3|60|他們要報復，謀害我， 你都看見了。
LAM|3|61|耶和華啊，你聽見他們的辱罵， 他們害我的一切計謀，
LAM|3|62|那些起來攻擊我的人嘴唇所說的話 和他們終日攻擊我的計謀。
LAM|3|63|求你留意！ 他們無論坐下或起來， 我都是他們的笑柄。
LAM|3|64|耶和華啊，求你照他們手所做的 向他們施行報應。
LAM|3|65|求你使他們心裏剛硬， 使你的詛咒臨到他們。
LAM|3|66|求你發怒追趕他們， 從耶和華的地上 除滅他們。
LAM|4|1|唉！黃金竟然無光！ 純金竟然變色！ 聖所的石頭散落在街上。
LAM|4|2|錫安 寶貝的孩子雖然好比精金， 現在竟當作陶匠手所做的瓦瓶！
LAM|4|3|野狗尚且哺乳其子， 我百姓 的婦人反倒殘忍， 如曠野的鴕鳥一般；
LAM|4|4|吃奶孩子的舌頭因乾渴貼住上膛， 孩童求餅，卻無人擘給他們。
LAM|4|5|素來吃美好食物的， 如今遭遺棄在街上； 素來穿著朱紅衣裳長大的， 如今卻擁抱糞堆。
LAM|4|6|我百姓的罪孽比 所多瑪 的罪還大； 所多瑪 雖無人伸手攻擊， 轉眼之間就被傾覆。
LAM|4|7|錫安 的拿細耳人 比雪純淨， 比奶更白； 他們的身體比寶石更紅， 身軀之美如藍寶石一般。
LAM|4|8|但如今他們的面貌比煤炭更黑， 在街上無人認識； 他們的皮膚緊貼骨頭， 枯乾形同槁木。
LAM|4|9|被刀劍刺殺的 勝過因飢餓而死 的； 飢餓者由於缺乏田裏的出產 就消瘦而亡 。
LAM|4|10|當我百姓遭毀滅的時候， 慈心的婦人親手烹煮自己的兒女為食物。
LAM|4|11|耶和華發盡他的憤怒， 傾倒他的烈怒， 用火焚燒 錫安 ， 燒燬 錫安 的根基。
LAM|4|12|地上的君王和世上的居民都不信 敵人和仇敵竟能進入 耶路撒冷 的城門。
LAM|4|13|這都因她先知的罪惡和祭司的罪孽， 他們在城中流了義人的血。
LAM|4|14|他們如盲人在街上徘徊， 又被血玷污， 以致人不敢摸他們的衣服。
LAM|4|15|人向他們喊著： 「你這不潔淨的，走開！ 走開！走開！不要摸我！」 他們逃走流浪的時候， 列國中有人說： 「他們不可再寄居此地。」
LAM|4|16|耶和華親自趕散他們， 不再眷顧他們； 不看重祭司，也不厚待長老。
LAM|4|17|我們的眼目徒然仰望幫助，以致失明， 我們從瞭望臺所守望的，竟是一個不能救人的國！
LAM|4|18|仇敵追逐我們的腳蹤， 使我們不敢在自己的街上行走。 我們的結局臨近， 日子已滿， 我們的結局已經來到。
LAM|4|19|追趕我們的比空中的鷹更快； 他們在山上追逼我們， 在曠野埋伏，等候我們。
LAM|4|20|耶和華的受膏者是我們鼻中的氣， 被抓到他們的坑裏， 論到他，我們曾說： 「我們必在他蔭下， 在列國中存活。」
LAM|4|21|住 烏斯 地的 以東 啊，儘管歡喜快樂， 苦杯必傳到你那裏； 你要喝醉，裸露自己。
LAM|4|22|錫安 哪，你罪孽的懲罰已經結束， 耶和華必不再使你被擄去。 以東 啊，耶和華必懲罰你的罪孽， 揭露你的罪惡。
LAM|5|1|耶和華啊，求你顧念我們所遭遇的， 留意看我們所受的凌辱。
LAM|5|2|我們的產業歸陌生人， 我們的房屋歸外邦人。
LAM|5|3|我們是無父的孤兒， 我們的母親如同寡婦。
LAM|5|4|我們出銀錢才得水喝， 我們的柴也是用錢買來的。
LAM|5|5|我們被追趕，迫及頸項， 疲乏卻不得歇息。
LAM|5|6|我們束手投降 埃及 和 亞述 ， 為要得糧吃飽。
LAM|5|7|我們的祖先犯罪，而今他們不在了， 我們卻擔當他們的罪孽。
LAM|5|8|奴僕轄制我們， 無人救我們脫離他們的手。
LAM|5|9|因曠野有刀劍， 我們冒生命的危險才能得糧食。
LAM|5|10|因饑荒的乾熱， 我們的皮膚熱如火爐。
LAM|5|11|他們在 錫安 玷污婦人， 在 猶大 城鎮污辱少女。
LAM|5|12|他們吊起領袖的手， 使長老臉上無光。
LAM|5|13|年輕人扛磨石， 孩童背木柴而跌倒。
LAM|5|14|城門口不再有老年人， 年輕人也不再奏樂。
LAM|5|15|我們心中的快樂止息， 跳舞轉為悲哀。
LAM|5|16|冠冕從我們的頭上掉落； 我們有禍了，因為犯了罪。
LAM|5|17|因這些事我們心裏發昏， 眼睛昏花。
LAM|5|18|錫安山 荒涼， 狐狸行在其上。
LAM|5|19|耶和華啊，你治理直到永遠， 你的寶座萬代長存。
LAM|5|20|你為何全然忘記我們？ 為何長久離棄我們？
LAM|5|21|耶和華啊，求你使我們回轉歸向你， 我們就得以回轉。 求你更新我們的年日，像古時一樣，
LAM|5|22|難道你全然棄絕了我們， 向我們大發烈怒？
EZEK|1|1|在三十年四月初五，我在 迦巴魯河 邊被擄的人當中，那時天開了，我看見上帝的異象。
EZEK|1|2|正是 約雅斤 王被擄的第五年四月初五，
EZEK|1|3|在 迦勒底 人之地的 迦巴魯河 邊，耶和華的話特地臨到 布西 的兒子 以西結 祭司，耶和華的手按在他身上。
EZEK|1|4|我觀看，看哪，狂風從北方颳來，有一朵大雲閃爍著火，周圍有光輝，其中的火好像閃耀的金屬；
EZEK|1|5|又從其中顯出四個活物的形像。他們的形狀是這樣：有人的形像，
EZEK|1|6|各有四張臉，四個翅膀。
EZEK|1|7|他們的腿是直的，腳掌好像牛犢的蹄，燦爛如磨亮的銅。
EZEK|1|8|在四面的翅膀以下有人的手。這四個活物的臉和翅膀是這樣：
EZEK|1|9|翅膀彼此相接，行走時並不轉彎，各自往前直行。
EZEK|1|10|至於臉的形像：四個活物各有人的臉，右面有獅子的臉，左面有牛的臉，也有鷹的臉；
EZEK|1|11|這就是他們的臉 。他們的翅膀向上張開，各有兩個翅膀彼此相接，用另外兩個翅膀遮體。
EZEK|1|12|他們各自往前直行。靈往哪裏去，他們就往哪裏去，行走時並不轉彎。
EZEK|1|13|至於四活物的形像，就如燒著火炭的形狀，又如火把的形狀。有火在四活物中間來回移動，這火有光輝，從火中發出閃電。
EZEK|1|14|這些活物往來奔走，好像電光一閃。
EZEK|1|15|我觀看活物，看哪，有四張臉的活物旁邊各有一個輪子在地上。
EZEK|1|16|輪子的形狀結構 好像耀眼的水蒼玉。四輪都是一個樣式，形狀 結構好像輪中套輪。
EZEK|1|17|輪子行走的時候，向四方直行，行走時並不轉彎。
EZEK|1|18|至於輪圈，高而可畏；四個輪圈周圍佈滿眼睛。
EZEK|1|19|活物行走，輪子也在旁邊行走；活物離地上升，輪子也上升。
EZEK|1|20|靈往哪裏去，活物就往哪裏去；輪子在活物旁邊上升，因為活物的靈在輪中。
EZEK|1|21|活物行走，輪子也行走；活物站住，輪子也站住；活物離地上升，輪子也在旁邊上升，因為活物的靈在輪中。
EZEK|1|22|活物的頭上面有穹蒼的形像，像耀眼驚人的水晶，鋪張在活物的頭頂上。
EZEK|1|23|穹蒼之下，活物的翅膀伸直，彼此相對，每個活物用兩個翅膀遮住自己；每個活物用兩個翅膀遮住自己 ，就是自己的身體。
EZEK|1|24|活物行走的時候，我聽見翅膀的響聲，像大水的聲音，像全能者的聲音，又像軍隊鬧鬨的聲音。活物站住的時候，翅膀垂下。
EZEK|1|25|在他們頭上的穹蒼之上有聲音。他們站住的時候，翅膀垂下。
EZEK|1|26|在他們頭上的穹蒼之上有寶座的形像，彷彿藍寶石的樣子；寶座的形像上方有彷彿人的樣子的形像。
EZEK|1|27|我見他的腰以上有彷彿閃耀的金屬，周圍有彷彿火的形狀，又見他的腰以下有彷彿火的形狀，周圍也有光輝。
EZEK|1|28|下雨的日子，雲中彩虹的形狀怎樣，周圍光輝的形狀也是怎樣。 這就是耶和華榮耀形像的樣式，我一看見就臉伏於地。我又聽見一位說話者的聲音。
EZEK|2|1|他對我說：「人子啊，你站起來，我要和你說話。」
EZEK|2|2|他對我說話的時候，靈進入我裏面，使我站起來，我就聽見他對我說話。
EZEK|2|3|他對我說：「人子啊，我差你往悖逆我的國家， 以色列 人那裏去，他們是悖逆我的。他們和他們的祖先違背我，直到今日。
EZEK|2|4|這些人厚著臉皮，心裏剛硬。我差你到他們那裏去，你要對他們說：『主耶和華如此說。』
EZEK|2|5|他們是悖逆之家，他們或聽，或不聽，必知道在他們中間有了先知。
EZEK|2|6|你，人子啊，雖有荊棘和蒺藜在你那裏，你又住在蠍子中間，總不要怕他們，也不要怕他們的話；他們雖是悖逆之家，但你不要怕他們的話，也不要因他們的臉色驚惶。
EZEK|2|7|他們或聽，或不聽，你只管將我的話告訴他們；他們是極其悖逆的。
EZEK|2|8|「但是你，人子啊，要聽我對你說的話，不要像那悖逆之家一樣悖逆，要開口吃我所賜給你的。」
EZEK|2|9|我觀看，看哪，有一隻手向我伸來；看哪，手中有一書卷。
EZEK|2|10|他在我面前展開書卷，它內外都寫著字，上面所寫的有哀號、嘆息、悲痛的話。
EZEK|3|1|他對我說：「人子啊，要吃你所得到的，吃下這書卷；然後要去，對 以色列 家宣講。」
EZEK|3|2|於是我張開了口，他就使我吃這書卷。
EZEK|3|3|他對我說：「人子啊，要吃我所賜給你的這書卷，塞滿你的肚腹。」我就吃了，口中覺得其甜如蜜。
EZEK|3|4|他對我說：「人子啊，你要到 以色列 家那裏去，對他們傳講我的話。
EZEK|3|5|你奉差遣不是往那說話艱澀、言語難懂的民那裏，而是往 以色列 家去；
EZEK|3|6|你不是往那說話艱澀、言語難懂的許多民族那裏去，他們的話你不懂。然而，我若差你往他們那裏去，他們會聽從你。
EZEK|3|7|以色列 家卻不肯聽從你，因為他們不肯聽從我；原來 以色列 全家是額頭堅硬、心裏剛愎的人。
EZEK|3|8|看哪，我使你的臉堅硬，對抗他們的臉；使你的額頭堅硬，對抗他們的額頭。
EZEK|3|9|我使你的額頭像金剛石，比火石更堅硬。他們雖是悖逆之家，但你不要怕他們，也不要因他們的臉色而驚惶。」
EZEK|3|10|他又對我說：「人子啊，我對你說的一切話，你心裏要領會，耳朵要聽。
EZEK|3|11|要到被擄的人，到你本國百姓那裏去，他們或聽，或不聽，你要對他們宣講，告訴他們這是主耶和華說的。」
EZEK|3|12|那時，靈將我舉起，我就聽見在我身後有極大震動的聲音：「耶和華的榮耀，從他所在之處，是應當稱頌的！」
EZEK|3|13|有活物的翅膀相碰的聲音，也有活物旁邊輪子的聲音，是極大震動的聲音。
EZEK|3|14|於是靈將我舉起，帶著我走。我就去了，十分苦惱，我的靈火熱；耶和華的手重重地按在我身上。
EZEK|3|15|我就來到 提勒‧亞畢 那些住在 迦巴魯河 邊被擄的人那裏，到他們住的地方 ，在他們中間驚愕地坐了七日。
EZEK|3|16|過了七日，耶和華的話臨到我，說：
EZEK|3|17|「人子啊，我立你作 以色列 家的守望者，所以你要聽我口中的話，替我警戒他們。
EZEK|3|18|我何時指著惡人說：『他必要死』；你若不警戒他，也不勸告他，使他離開惡行，拯救他的性命，這惡人必死在罪孽之中；我卻要從你手裏討他的血債。
EZEK|3|19|倘若你警戒惡人，他仍不轉離罪惡，也不離開惡行，他必死在罪孽之中，你卻救了自己的命。
EZEK|3|20|但是義人若轉離他的義而作惡，我要把絆腳石放在他面前，他必死亡；因你沒有警戒他，他必死在罪中，他素來所行的義不被記念；我卻要從你手裏討他的血債。
EZEK|3|21|倘若你警戒義人，使他不犯罪，他就不犯罪；他因領受警戒就必存活，你也救了自己的命。」
EZEK|3|22|在那裏耶和華的手按在我身上。他對我說：「起來，到平原去，我要在那裏和你說話。」
EZEK|3|23|於是我起來，到平原去，看哪，耶和華的榮耀停在那裏，正如我在 迦巴魯河 邊所見到的一樣，我就臉伏於地。
EZEK|3|24|靈進入我裏面，使我站起來。耶和華對我說：「你進屋裏去，把門關上。
EZEK|3|25|你，人子，看哪，人要用繩索捆綁你，使你不能出去到他們中間。
EZEK|3|26|我必使你的舌頭貼住上膛，以致你啞口，不能作責備他們的人；他們原是悖逆之家。
EZEK|3|27|但我對你說話的時候，必使你開口，你就要對他們說：『主耶和華如此說。』聽的，讓他聽；不聽的，任他不聽，因為他們是悖逆之家。」
EZEK|4|1|「你，人子啊，拿一塊磚，擺在你面前，將一座城 耶路撒冷 畫在上面。
EZEK|4|2|你要圍攻這城，築堡壘，建土堆，安營攻擊，周圍設撞城槌攻城，
EZEK|4|3|又要拿一個鐵盤放在你和城的中間，作為鐵牆。你要把你的臉對著這城，使城被困。你要圍攻這城，這要成為 以色列 家的預兆。
EZEK|4|4|「你要向左側臥，承擔 以色列 家的罪孽；按你向左側臥的日數，擔當他們的罪孽。
EZEK|4|5|我已將他們作惡的年數定了日期，就是三百九十天，你要如此擔當 以色列 家的罪孽。
EZEK|4|6|這些日子結束之後，你還要向右側臥，擔當 猶大 家的罪孽。我為你定了四十天，一天頂一年。
EZEK|4|7|你要把你的臉對著被困的 耶路撒冷 ，露出膀臂，說預言攻擊這城。
EZEK|4|8|看哪，我用繩索捆綁你，使你不能從這邊翻到那邊，直等到你圍困的日子結束。
EZEK|4|9|「你要取小麥、大麥、豆子、紅豆、小米、粗麥，裝在一個器皿裏，為自己做餅；在你側臥的三百九十天吃這餅。
EZEK|4|10|你所吃食物的量是每天二十舍客勒，要按時吃。
EZEK|4|11|你喝水的量是每天六分之一欣，要按時喝。
EZEK|4|12|你要吃這餅像大麥餅一樣，在眾人眼前用人的糞烤它。」
EZEK|4|13|耶和華說：「 以色列 人在我趕他們到的列國中，也必這樣吃不潔淨的食物。」
EZEK|4|14|我說：「唉！主耶和華，看哪，我從來未曾被玷污，從幼年到如今沒有吃過自然死的，或被野獸撕裂的，那不潔淨的肉也未曾入我的口。」
EZEK|4|15|於是他對我說：「看，我給你牛糞代替人糞，你要在上面烤你的餅。」
EZEK|4|16|他又對我說：「人子，看哪，我必斷絕 耶路撒冷 糧食的供應 。他們要帶著憂慮限量吃餅；帶著驚惶限量喝水。
EZEK|4|17|他們因缺糧缺水，彼此驚惶，在自己的罪孽中消滅。」
EZEK|5|1|「你，人子啊，拿一把快刀當作剃刀，用這刀剃你的頭髮和鬍鬚，然後用天平將鬚髮分成幾份。
EZEK|5|2|圍困的日子滿了，你要把三分之一放在城中用火焚燒；三分之一放在城的四圍用刀砍碎；三分之一任風吹散，我要拔刀追趕它們。
EZEK|5|3|你要從其中取幾根鬚髮，用衣服的邊包起來，
EZEK|5|4|再從其中取一些扔在火裏，在火中焚燒；必有火從其中出來燒盡 以色列 全家。
EZEK|5|5|主耶和華如此說：這就是 耶路撒冷 。我曾將它安置在列國中，列邦都在它的四圍。
EZEK|5|6|耶路撒冷 行惡，違背我的典章，過於列國；干犯我的律例，過於四圍的列邦。它棄絕我的典章，也沒有遵行我的律例。
EZEK|5|7|所以主耶和華如此說：因為你們混亂，過於四圍的列國，不遵行我的律例，不順從我的典章，甚至也不順從四圍列國的規條 ，
EZEK|5|8|所以主耶和華如此說：看哪，我，我必與你為敵，必在列國眼前，在你中間施行審判；
EZEK|5|9|並且因你一切可憎的事，我要在你中間行未曾行過，將來也不會行的事。
EZEK|5|10|在你中間，父親要吃兒子，兒子要吃父親。我必向你施行審判，將你剩下的人分散四方 。
EZEK|5|11|主耶和華說：我指著我的永生起誓，因你用一切可憎之物、可厭的事玷污我的聖所，所以，我要把你剃光 ，我的眼必不顧惜你，也不可憐你。
EZEK|5|12|你的百姓三分之一必遭瘟疫而死，因饑荒在你們中間而消滅；三分之一必在你四圍倒在刀下；我必將三分之一分散四方，要拔刀追趕他們。
EZEK|5|13|「我要這樣發盡我的怒氣；我向他們發的憤怒停止以後，自己就得到平息。當我向他們發盡我的憤怒時，他們就知道我─耶和華所說的是出於妒忌。
EZEK|5|14|在四圍的列國中，我要使你成為荒涼，在所有過路人的眼前看為羞辱。
EZEK|5|15|這樣，我必以怒氣、憤怒和烈怒的責備，向你施行審判。那時，它 就在四圍的列國中成為羞辱、譏刺、警戒、驚駭；這是我─耶和華說的。
EZEK|5|16|我向滅亡的人射出饑荒的惡箭，將它們射出，毀滅你們；那時，我要加重你們的饑荒，斷絕你們糧食的供應。
EZEK|5|17|我要令饑荒和惡獸臨到你，使你喪失兒女。瘟疫和流血的事必在你那裏盛行，我也要使刀劍臨到你。這是我─耶和華說的。」
EZEK|6|1|耶和華的話臨到我，說：
EZEK|6|2|「人子啊，你要面向 以色列 的眾山說預言。
EZEK|6|3|你要說： 以色列 的眾山哪，要聽主耶和華的話。主耶和華對大山、小岡、水溝、山谷如此說：看哪，我要使刀劍臨到你們，也必毀壞你們的丘壇。
EZEK|6|4|你們的祭壇要荒廢，香壇必打碎。我要使你們當中被殺的人仆倒在你們的偶像面前，
EZEK|6|5|將 以色列 人的屍首放在他們的偶像面前，把你們的骸骨拋散在祭壇的四周圍。
EZEK|6|6|無論你們住在何處，城鎮要變為廢墟，丘壇也必毀壞，以至於你們的祭壇荒廢，被定罪 ，偶像打碎消除，香壇砍倒；你們所做的被塗去。
EZEK|6|7|被殺的人必仆倒在你們中間，你們就知道我是耶和華。
EZEK|6|8|「我必留下一些人，你們中有人得以在列國中脫離刀劍，分散在列邦。
EZEK|6|9|那些逃脫的人，必在被擄所到的各國中記得我，我心裏何等傷痛，因他們起淫心，離棄我，淫蕩的眼追隨偶像。他們因所做一切可憎的惡事，必厭惡自己。
EZEK|6|10|他們必知道我是耶和華；我說過要使這災禍臨到他們身上，並非空話。
EZEK|6|11|「主耶和華如此說：你當擊掌頓足，說：哀哉！ 以色列 家做了這一切可憎的惡事，必仆倒在刀劍、饑荒、瘟疫之下。
EZEK|6|12|在遠方的，必遭瘟疫而死；在近處的，必倒在刀劍之下；那存留被圍困的，必因饑荒而死；我要在他們身上發盡我的憤怒。
EZEK|6|13|被殺的要仆倒在祭壇四圍的偶像中，在各高岡、各山頂、各青翠的樹下，和各茂密的橡樹下，就是他們獻馨香的祭給一切偶像的地方。那時，他們就知道我是耶和華。
EZEK|6|14|我必伸手攻擊他們，使他們的地荒廢，從 第伯拉他 的曠野起 ，一切的住處都荒涼。他們就知道我是耶和華。」
EZEK|7|1|耶和華的話又臨到我，說：
EZEK|7|2|「你，人子啊，主耶和華對 以色列 地如此說：結局，結局臨到了地的四境！
EZEK|7|3|現在你的結局已經來臨；我要使我的怒氣臨到你，也要按你的行為審判你，照你所做一切可憎的事懲罰你。
EZEK|7|4|我的眼必不顧惜你，也不可憐你，卻要按你所做的報應你，照你們中間可憎的事懲罰你；你就知道我是耶和華。
EZEK|7|5|「主耶和華如此說：災難，惟一的災難 ，看哪，臨近了！
EZEK|7|6|結局到了，結局到了，它要醒起來攻擊你。看哪，它已來到！
EZEK|7|7|境內的居民哪，厄運臨到你；時候到了，日子近了，有鬧鬨，但不是山上歡呼的聲音。
EZEK|7|8|我快要將我的憤怒傾倒在你身上，向你發盡我的怒氣，按你的行為審判你，照你所做一切可憎的事懲罰你。
EZEK|7|9|我的眼必不顧惜你，也不可憐你，必按你所做的報應你，照你中間可憎的事懲罰你；你就知道擊打你的是我─耶和華。
EZEK|7|10|「看哪，那日子！看哪，已來到！厄運已經發生！杖已開花，驕傲已發芽。
EZEK|7|11|殘暴興起，成了罰惡的杖。他們將一無所有，他們的富足 、他們的財寶 都不復存在；他們中間也不再有尊榮。
EZEK|7|12|時候到了，日子近了，買主不可歡喜，賣主也不用愁煩，因為烈怒已經臨到他們眾人身上。
EZEK|7|13|賣主即使存活，也不能討回所賣的，因為這異象關乎他們眾人；誰都不能討回，也沒有人能在罪孽中使自己的生命剛強。」
EZEK|7|14|「他們吹了角，預備齊全，卻無一人出戰，因為我的烈怒臨到他們眾人身上。
EZEK|7|15|外有刀劍，內有瘟疫、饑荒。在田野的，必因刀劍而死；在城中的，必遭饑荒、瘟疫吞滅。
EZEK|7|16|其中倖存的要逃脫，各人因自己的罪孽在山上發出悲聲，如谷中的鴿子哀鳴；
EZEK|7|17|雙手發軟，膝蓋軟弱如水，
EZEK|7|18|腰束麻布，戰慄籠罩他們；各人臉上羞愧，頭上光禿。
EZEK|7|19|他們要把銀子拋棄在街上，看金子如污穢之物。正當耶和華發怒的日子，金銀不能拯救他們，不能滿足食慾，也不能使肚腹飽滿，反倒成了自己罪孽的絆腳石。
EZEK|7|20|他們用所誇耀華美的妝飾製造可憎可厭的偶像，所以我使他們看它如污穢之物。
EZEK|7|21|我必將它交給外邦人為掠物，交給地上的惡人為擄物；他們要褻瀆它。
EZEK|7|22|他們褻瀆我寶貴之所 ，強盜也進去褻瀆它。我必轉臉不顧 以色列 人 。
EZEK|7|23|「要製造鎖鏈；因為遍地都有流血的罪，滿城都是殘暴的事。
EZEK|7|24|所以，我要使列國中最兇惡的人前來佔據他們的房屋；我要止息殘暴人的驕傲，他們的聖所也要被褻瀆。
EZEK|7|25|毀滅來到；他們求平安，卻沒有平安。
EZEK|7|26|災害加上災害，風聲接連風聲；他們要向先知尋求異象，但祭司的教誨、長老的謀略都必斷絕。
EZEK|7|27|君王要悲哀，官長要披絕望為衣，這地百姓的手都發顫。我必照他們所做的待他們，按他們所應得的審判他們，他們就知道我是耶和華。」
EZEK|8|1|第六年六月初五，我坐在家中； 猶大 的眾長老坐在我面前。在那裏主耶和華的手降在我身上。
EZEK|8|2|我觀看，看哪，有形像彷彿火 的形狀，從他腰部以下形狀是火，從他腰部以上有光輝的形狀，好像閃耀的金屬。
EZEK|8|3|他伸出一隻手的樣式，抓住我的一綹頭髮，靈就將我舉到天地中間；在上帝的異象中，他帶我到 耶路撒冷 朝北的內院門口，在那裏有惹動妒忌的偶像的座位，它惹動了妒忌。
EZEK|8|4|看哪，在那裏有 以色列 上帝的榮耀，形狀與我在平原所見的一樣。
EZEK|8|5|上帝對我說：「人子啊，你舉目向北觀看。」我就舉目向北觀看，看哪，祭壇門北邊的門口有那惹動妒忌的偶像。
EZEK|8|6|他又對我說：「人子啊，你看見 以色列 家所做的嗎？他們在這裏做了極其可憎的事，使我遠離我的聖所。你還要看見另有極其可憎的事。」
EZEK|8|7|他領我到院子門口。我觀看，看哪，牆上有一個洞。
EZEK|8|8|他對我說：「人子啊，你要挖牆。」我就挖牆。看哪，有一扇門。
EZEK|8|9|他說：「你進去，看他們在這裏所做可憎的惡事。」
EZEK|8|10|於是我進去看。看哪，四面牆上刻著各樣爬行的動物、可憎的走獸和 以色列 家各樣的偶像。
EZEK|8|11|以色列 家的七十個長老站在這些像前， 沙番 的兒子 雅撒尼亞 也站在其中，各人手拿他的香爐，煙雲的香氣上騰。
EZEK|8|12|他對我說：「人子啊，你看見 以色列 家的長老，暗中在自己偶像的房間裏所做的嗎？因為他們說：『耶和華看不見我們；耶和華已經離棄這地。』」
EZEK|8|13|他又說：「你還要看見他們所做另外極其可憎的事。」
EZEK|8|14|他領我到耶和華殿朝北的門口。看哪，在那裏有婦女們坐著，為 搭模斯 哭泣。
EZEK|8|15|他對我說：「人子啊，你看見了嗎？你還要看見比這更可憎的事。」
EZEK|8|16|然後他領我到耶和華殿的內院。看哪，在耶和華殿門口、走廊和祭壇中間，約有二十五個人背向耶和華的殿，面向東方，向東拜太陽。
EZEK|8|17|他對我說：「人子啊，你看見了嗎？ 猶大 家在這裏行可憎的事還算為小嗎？他們遍地行殘暴，再三惹我發怒。看哪，他們手拿枝條舉向鼻前 ！
EZEK|8|18|因此，我也要以憤怒行事。我的眼必不顧惜，也不可憐他們；他們雖在我耳邊大聲呼求，我還是不聽。」
EZEK|9|1|他在我耳邊大聲喊叫，說：「上前來啊，懲罰這城的人，手中要各拿毀滅的兵器。」
EZEK|9|2|看哪，有六個人從朝北的 上門 而來，各人手裏拿著致命的兵器；他們當中有一人身穿細麻衣，腰間繫著文士用的墨盒。他們進來，站在銅的祭壇旁。
EZEK|9|3|在基路伯之上， 以色列 上帝的榮耀從那裏上升，到殿的入口處。上帝召那身穿細麻衣、腰間繫著墨盒的人前來。
EZEK|9|4|耶和華對他說：「你去走遍 耶路撒冷 全城，那些為城中所做可憎之事嘆息哀哭的人，你要在他們額上做記號。」
EZEK|9|5|我耳中聽見耶和華對其餘的人說：「要跟隨他走遍全城去擊殺。你們的眼不要顧惜，也不要可憐他們。
EZEK|9|6|要將年老的、年輕的、少女、孩童和婦女，從我的聖所開始全都殺盡，只是不可挨近凡有記號的人。」於是他們從殿前的長老殺起。
EZEK|9|7|他對他們說：「要使這殿污穢，使院中遍滿被殺的人。你們出去吧！」他們就出去，在城中擊殺。
EZEK|9|8|他們擊殺的時候，只剩我一人，我就臉伏在地上，呼喊說：「唉！主耶和華啊，你將憤怒傾倒在 耶路撒冷 ，豈要把 以色列 所剩餘的人都滅絕嗎？」
EZEK|9|9|他對我說：「 以色列 家和 猶大 家的罪孽極其重大。遍地都有流血的事，滿城有冤屈，因為他們說：『耶和華已經離棄這地，他看不見我們。』
EZEK|9|10|因此，我的眼必不顧惜，也不可憐他們，要照他們所做的報應在他們頭上。」
EZEK|9|11|看哪，那身穿細麻衣、腰間繫著墨盒的人回覆這事說：「我已經照你所吩咐的做了。」
EZEK|10|1|我觀看，看哪，在穹蒼之中，也就是基路伯的頭上，有藍寶石的形狀，彷彿寶座的形像顯在他們上面。
EZEK|10|2|耶和華對那身穿細麻衣的人說：「你進到基路伯下面旋轉的輪子中，從基路伯之間取出火炭裝滿兩手掌，撒在城上。」 我親眼看見他進去。
EZEK|10|3|那人進去的時候，基路伯站在殿的南邊，雲彩充滿了內院。
EZEK|10|4|耶和華的榮耀從基路伯那裏上升，到殿的入口處；殿內滿佈雲彩，院子也充滿了耶和華榮耀的光輝。
EZEK|10|5|基路伯翅膀的響聲傳到外院，好像全能上帝說話的聲音。
EZEK|10|6|耶和華吩咐那身穿細麻衣的人說：「要從基路伯之間旋轉的輪子中取火。」那人就進去站在一個輪子旁邊。
EZEK|10|7|基路伯中的一個基路伯伸手到基路伯中間的火那裏，取一些放在那身穿細麻衣人的手掌中，那人拿了就出去。
EZEK|10|8|在基路伯翅膀以下，顯出有人手的樣式。
EZEK|10|9|我又觀看，看哪，這些基路伯的旁邊有四個輪子。一個基路伯旁有一個輪子，另一個基路伯旁也有一個輪子；輪子的形狀好像水蒼玉石。
EZEK|10|10|至於四輪的形狀，都是一個樣式，好像輪中套輪。
EZEK|10|11|輪子行走的時候，向四方都能直行，行走時並不轉彎。頭轉向何方，它們也隨著向何方行走，行走時並不轉彎。
EZEK|10|12|基路伯的全身，連背帶手和翅膀，並輪子周圍都佈滿眼睛。他們四個的輪子都是如此。
EZEK|10|13|我耳中聽見這些輪子稱為「旋轉的輪」。
EZEK|10|14|基路伯各有四張臉：第一是基路伯的臉，第二是人的臉，第三是獅子的臉，第四是鷹的臉。
EZEK|10|15|基路伯升上去了；這就是我在 迦巴魯河 邊所看見的活物。
EZEK|10|16|基路伯行走，輪子也在旁邊行走。基路伯展開翅膀，離地上升，輪子也不轉離他們的旁邊。
EZEK|10|17|基路伯站住，輪子也站住；基路伯上升，輪子也跟著上升，因為活物的靈在輪中。
EZEK|10|18|耶和華的榮耀離開殿的入口處，停在基路伯之上。
EZEK|10|19|基路伯展開翅膀，在我眼前離地上升；他們離去的時候，輪子在旁邊，都停在耶和華殿的東門口。在他們上面有 以色列 上帝的榮耀。
EZEK|10|20|這是我在 迦巴魯河 邊所見的活物，他們在 以色列 上帝之下；因此我知道他們是基路伯。
EZEK|10|21|他們各有四張臉、四個翅膀，翅膀以下有人手的樣式。
EZEK|10|22|至於他們臉的模樣，以及身體的形像 ，正是我從前在 迦巴魯河 邊所看見的。他們各自往前直行。
EZEK|11|1|靈將我舉起，帶我到耶和華聖殿面向東方的東門。看哪，門口有二十五個人。我見其中有百姓的領袖 押朔 的兒子 雅撒尼亞 和 比拿雅 的兒子 毗拉提 。
EZEK|11|2|耶和華對我說：「人子啊，他們就是圖謀罪孽，在這城中設計惡謀的人。
EZEK|11|3|他們說：『蓋房屋的時候尚未臨近；這城是鍋，我們是肉。』
EZEK|11|4|人子啊，因此你當說預言，說預言攻擊他們。」
EZEK|11|5|耶和華的靈降在我身上，對我說：「你當說，耶和華如此說： 以色列 家啊，你們所說的，你們心裏所想的，我都知道。
EZEK|11|6|你們在這城裏大行屠殺，被殺的人遍滿街道。
EZEK|11|7|所以主耶和華如此說：你們在城中殺的人是肉，這城是鍋；你們卻要從其中被帶出去。
EZEK|11|8|你們怕刀劍，我卻要使刀劍臨到你們。這是主耶和華說的。
EZEK|11|9|我要把你們從這城中帶出去，交在外邦人的手裏，且要在你們中間施行審判。
EZEK|11|10|你們要仆倒在刀下；我必在 以色列 的邊界審判你們，你們就知道我是耶和華。
EZEK|11|11|這城必不作你們的鍋，你們也不作鍋中的肉。我要在 以色列 的邊界審判你們，
EZEK|11|12|你們就知道我是耶和華；因為你們不遵行我的律例，也不順從我的典章，卻隨從你們四圍列國的規條。」
EZEK|11|13|我正說預言的時候， 比拿雅 的兒子 毗拉提 死了。於是我臉伏在地，大聲呼叫說：「唉！主耶和華啊，你要把 以色列 剩餘的人都滅絕淨盡嗎？」
EZEK|11|14|耶和華的話臨到我，說：
EZEK|11|15|「人子啊， 耶路撒冷 的居民對你的兄弟、你的本家、你的親屬、 以色列 全家所有的人說：『你們遠離耶和華吧！這地是賜給我們為業的。』
EZEK|11|16|所以你當說：『主耶和華如此說：我雖將 以色列 全家遠遠流放到列國，使他們分散在列邦，我卻要在他們所到的列邦，暫時作他們的聖所。』
EZEK|11|17|你當說：『主耶和華如此說：我必從萬民中召集你們，從分散的列邦中聚集你們，又將 以色列 地賜給你們。』
EZEK|11|18|他們到了那裏，必從其中除掉一切可憎之物、可厭的事。
EZEK|11|19|我要使他們有合一的心，也要將新靈放在你們 裏面，又從他們的肉體中除掉石心，賜給他們肉心，
EZEK|11|20|使他們順從我的律例，謹守遵行我的典章。他們要作我的子民，我要作他們的上帝。
EZEK|11|21|至於那些心中隨從可憎之物、可厭的事的人，我必照他們所做的報應在他們頭上。這是主耶和華說的。」
EZEK|11|22|於是，基路伯展開翅膀，輪子都在他們旁邊；在他們上面有 以色列 上帝的榮耀。
EZEK|11|23|耶和華的榮耀從城中上升，停在城東的那座山上。
EZEK|11|24|靈將我舉起，在異象中上帝的靈將我帶回 迦勒底 地，到被擄的人那裏；之後我所見的異象就離我上升去了。
EZEK|11|25|我就把耶和華指示我的一切事都說給被擄的人聽。
EZEK|12|1|耶和華的話臨到我，說：
EZEK|12|2|「人子啊，你住在悖逆之家中；他們有眼可看卻看不見，有耳可聽卻聽不到，因為他們是悖逆之家。
EZEK|12|3|所以人子啊，你要收拾被擄時需用的物件，白天在他們眼前離去，在他們眼前離開你所住的地方，移到別處去；他們雖是悖逆之家，或者可以領悟。
EZEK|12|4|你要白天在他們眼前拿出你被擄時需用的物件。到了晚上，要在他們眼前離去，像被擄的人離去一樣。
EZEK|12|5|你要在他們眼前挖通牆壁，從其中將物件帶出去 。
EZEK|12|6|到天黑時，在他們眼前背在肩上帶走 ，並要蒙住臉看不見地，因為我要使你成為 以色列 家的預兆。」
EZEK|12|7|我就照著所吩咐的去做，白天拿出被擄時需用的物件。到了晚上，用手挖通牆壁；天黑的時候，在他們眼前背在肩上帶走。
EZEK|12|8|次日早晨，耶和華的話臨到我，說：
EZEK|12|9|「人子啊， 以色列 家，就是那悖逆之家，豈不是問你說：『你在做甚麼呢？』
EZEK|12|10|你要對他們說：『主耶和華如此說：這是關乎 耶路撒冷 君王和其中 以色列 全家的默示。』
EZEK|12|11|你要說：『我是你們的預兆：我怎樣做，他們所遭遇的也必這樣，他們必被擄去，作俘虜。』
EZEK|12|12|他們中間的君王也必在天黑時把物件背在肩上帶走。他們要挖通牆壁，從其中帶出去 。他必蒙住臉，眼看不見地。
EZEK|12|13|我要把我的網撒在他身上，他就被我的羅網纏住。我要帶他到 迦勒底 人之地的 巴比倫 ；他沒有看見那地，就死在那裏。
EZEK|12|14|我要把四圍幫助他的和他所有的軍隊分散到四方 ，也要拔刀追趕他們。
EZEK|12|15|我把他們驅逐到列國，分散在列邦的時候，他們就知道我是耶和華。
EZEK|12|16|我卻要留下他們當中幾個人得免刀劍、饑荒、瘟疫，使他們在所到的列國述說自己所做一切可憎的事；他們就知道我是耶和華。」
EZEK|12|17|耶和華的話臨到我，說：
EZEK|12|18|「人子啊，你吃飯時必戰抖，喝水時必驚惶憂慮。
EZEK|12|19|你要對這地的百姓說：主耶和華論 以色列 地的 耶路撒冷 居民如此說，他們吃飯時必憂慮，喝水時必驚惶，因其中居民所行殘暴的事，這地必然荒廢，一無所存。
EZEK|12|20|有人居住的城鎮必變為廢墟，地必荒涼；你們就知道我是耶和華。」
EZEK|12|21|耶和華的話臨到我，說：
EZEK|12|22|「人子啊，在 以色列 地你們怎麼有這俗語說：『日子延長，一切異象卻落了空』呢？
EZEK|12|23|你要告訴他們說：『主耶和華如此說：我必令這俗語止息， 以色列 中不再有人引用這俗語。』你卻要對他們說：『日子臨近，一切的異象都必應驗。』
EZEK|12|24|從此以後， 以色列 家不再有虛假的異象和奉承的占卜。
EZEK|12|25|我─耶和華說話，所說的必定實現，不再耽延。你們這悖逆之家啊，你們在世的日子，我所說的話必定實現。這是主耶和華說的。」
EZEK|12|26|耶和華的話臨到我，說：
EZEK|12|27|「人子，看哪， 以色列 家的人說：『他所見的異象是許多日子以後的事，所說的預言是指著遙遠的時候。』
EZEK|12|28|所以你要對他們說：『主耶和華如此說：我的話不再有一句耽延，我所說的話必定實現。』這是主耶和華說的。」
EZEK|13|1|耶和華的話臨到我，說：
EZEK|13|2|「人子啊，你要說預言，攻擊 以色列 中說預言的先知，對那些隨心說預言的人說：『你們當聽耶和華的話。』」
EZEK|13|3|主耶和華如此說：「禍哉！那些愚頑的先知，隨從自己的心意，卻一無所見
EZEK|13|4|以色列 啊，你的先知好像廢墟中的狐狸，
EZEK|13|5|沒有上去堵住缺口，也沒有為 以色列 家重修城牆，使它在耶和華的日子來臨時，可以在戰爭中站得住。
EZEK|13|6|他們看見的是虛假，是謊詐的占卜，說是耶和華說的；其實耶和華並沒有差遣他們，他們卻指望那話必站立得住。
EZEK|13|7|你們豈不是見了虛假的異象嗎？豈不是說了謊詐的占卜嗎？你們說，這是耶和華說的，其實我沒有說過。」
EZEK|13|8|所以主耶和華如此說：「因你們說的是虛假，見的是謊詐，所以，看哪，我要敵對你們。這是主耶和華說的。
EZEK|13|9|我的手必攻擊那見虛假異象、用謊詐占卜的先知，他們必不列在我百姓的會中，不錄在 以色列 家的名冊上，也不能進入 以色列 地；你們就知道我是主耶和華。
EZEK|13|10|他們誘惑我的百姓，說：『平安！』其實沒有平安，就像有人築牆壁，看哪，他們倒去粉刷它。
EZEK|13|11|所以你要對那些粉刷的人說：『牆要倒塌，暴雨漫過。你們大冰雹啊，要降下 ，狂風要吹裂這牆。』
EZEK|13|12|看哪，這牆倒塌，人豈不是要問你們說：『你們所粉刷的在哪裏呢？』」
EZEK|13|13|所以主耶和華如此說：「我要發怒，使狂風吹裂它，在怒中令暴雨漫過，又發怒降下大冰雹，毀壞它。
EZEK|13|14|我要這樣拆毀你們那粉飾的牆，把它夷為平地，以致根基露出；牆一倒塌，你們也要在其中滅亡。你們就知道我是耶和華。
EZEK|13|15|我要對牆和粉刷它的人發盡我的憤怒，我 要對你們說：『牆沒有了！粉刷它的人也沒有了！』
EZEK|13|16|這就是 以色列 的先知，他們指著 耶路撒冷 說預言，見到這城平安的異象，其實沒有平安。這是主耶和華說的。」
EZEK|13|17|「你，人子啊，要面向你百姓中隨心說預言的婦女們，說預言攻擊她們，
EZEK|13|18|說，主耶和華如此說：『這些婦女有禍了！她們為眾人的手腕縫驅邪帶，替身材高矮不同的人做頭巾，為要獵取人的性命。難道你們要獵取我百姓的性命，使自己存活嗎？
EZEK|13|19|你們為幾把大麥、幾塊餅，在我的百姓中褻瀆我，對那肯聽謊言的百姓說謊言，讓不該死的人死，讓不該活的人活。』」
EZEK|13|20|所以主耶和華如此說：「看哪，我要對付你們那用以獵取人，如獵飛鳥般的驅邪帶。我要把驅邪帶從你們的手腕扯去，釋放那些如飛鳥被你們獵取的人。
EZEK|13|21|我也必撕裂你們的頭巾，救我百姓脫離你們的手，使他們不再被獵取，落在你們手中；你們就知道我是耶和華。
EZEK|13|22|我未曾使義人傷心，你們卻以謊話使他傷心，且又堅固惡人的手，不使他回轉離開惡道得以存活。
EZEK|13|23|所以，你們必不再看見虛假的異象，也不再行占卜的事；我要救我的百姓脫離你們的手；你們就知道我是耶和華。」
EZEK|14|1|有幾個 以色列 的長老到我這裏來，坐在我面前。
EZEK|14|2|耶和華的話臨到我，說：
EZEK|14|3|「人子啊，這些人在心中設立偶像，把陷自己於罪的絆腳石放在面前，我真的能讓他們求問嗎？
EZEK|14|4|所以你要告訴他們，對他們說：『主耶和華如此說： 以色列 家的人，凡在心中設立偶像，把陷自己於罪的絆腳石放在面前，卻來到先知那裏的，我─耶和華在他所求的事上，必因他拜許多偶像向他施行報應 ，
EZEK|14|5|為要奪回 以色列 家的心，他們全都拜偶像，與我疏遠了。』
EZEK|14|6|「所以你要對 以色列 家說：『主耶和華如此說：回轉吧！回轉離開你們的偶像，轉臉離開一切可憎的事。』
EZEK|14|7|因為 以色列 家的人，或在 以色列 中寄居的外人，凡與我隔絕，在心中設立偶像，把陷自己於罪的絆腳石放在面前，卻來到先知那裏，要為自己的事求問我的，我─耶和華必親自報應他。
EZEK|14|8|我要向那人變臉，使他成為警戒和笑柄，並且我要把他從我民中剪除；你們就知道我是耶和華。
EZEK|14|9|先知若被騙說了一句預言，是我─耶和華騙了那先知，我要伸手攻擊他，把他從我百姓 以色列 中除滅。
EZEK|14|10|他們必擔當自己的罪孽。先知的罪孽和求問之人的罪孽都一樣，
EZEK|14|11|使 以色列 家不再走迷離開我，也不再因各樣的罪過玷污自己，卻要作我的子民，我也作他們的上帝。這是主耶和華說的。」
EZEK|14|12|耶和華的話臨到我，說：
EZEK|14|13|「人子啊，若有一國犯罪干犯我，我也伸手攻擊它，斷絕他們糧食的供應，使饑荒臨到那地，將人與牲畜從其中剪除；
EZEK|14|14|雖有 挪亞 、 但以理 、 約伯 這三人在那裏，他們只能因自己的義救自己的命。這是主耶和華說的。
EZEK|14|15|我若使惡獸經過那地，大肆蹂躪，使地荒涼，以致因這些獸，人都不得經過；
EZEK|14|16|雖有這三人在其中，主耶和華說：我指著我的永生起誓，他們不能救兒子女兒，只有他們自己可以得救，那地仍然荒涼。
EZEK|14|17|或者我使刀劍臨到那地，說：『讓刀劍穿越那地』，以致我把人與牲畜從其中剪除；
EZEK|14|18|雖有這三人在其中，主耶和華說：我指著我的永生起誓，他們不能救兒子女兒，只有他們自己可以得救。
EZEK|14|19|或者我叫瘟疫流行那地，把我的憤怒帶著血傾在其中，好使人與牲畜從其中剪除；
EZEK|14|20|雖有 挪亞 、 但以理 、 約伯 在那裏，主耶和華說：我指著我的永生起誓，他們不能救兒子女兒，只能因自己的義救自己的命。
EZEK|14|21|「主耶和華如此說：我若將這四樣大災，就是刀劍、饑荒、惡獸、瘟疫降在 耶路撒冷 ，將人與牲畜從其中剪除，豈不是更嚴重嗎？
EZEK|14|22|看哪，在那裏必有倖免於難的人帶著兒子女兒；看哪，他們來到你們這裏；你們看見他們的所作所為，就會因我降給 耶路撒冷 的災禍，因我降給它的一切，得到安慰。
EZEK|14|23|你們因看見他們的所作所為，得到安慰，就會知道我在 耶路撒冷 所做的並非毫無緣故。這是主耶和華說的。」
EZEK|15|1|耶和華的話臨到我，說：
EZEK|15|2|「人子啊，葡萄樹比一切其他的樹，就是樹林裏眾樹木的樹枝，有甚麼長處呢？
EZEK|15|3|可以從其中取木料來做工嗎？人可以拿來做釘子，掛東西在上面嗎？
EZEK|15|4|看哪，它已經拋在火中當柴燒，火既燒了兩頭，中間也燒焦了，它還有甚麼用處呢？
EZEK|15|5|看哪，它完整的時候尚且不能拿來做工，何況被火燒焦了，還能拿來做工嗎？
EZEK|15|6|所以，主耶和華如此說：我怎樣使林中樹裏的葡萄樹在火中當柴燒，我也必照樣對待 耶路撒冷 的居民。
EZEK|15|7|我必向他們變臉；他們雖從火中逃出來，火仍要燒滅他們。我向他們變臉的時候，你們就知道我是耶和華。
EZEK|15|8|我必使這地荒涼，因為他們做了背叛的事。這是主耶和華說的。」
EZEK|16|1|耶和華的話臨到我，說：
EZEK|16|2|「人子啊，你要使 耶路撒冷 知道它那些可憎的事。
EZEK|16|3|你要說，主耶和華對 耶路撒冷 如此說：你的根源，你的出身，是在 迦南 地；你的父親是 亞摩利 人，母親是 赫 人。
EZEK|16|4|論到你出世的景況，在你出生的日子沒有人為你斷臍帶，也沒有用水清洗，使你潔淨；沒有人撒鹽在你身上，也沒有人用布包你。
EZEK|16|5|沒有人顧惜你，為你做一件這樣的事來可憐你。你卻被扔在田野上面，因你出生的日子就被厭惡。
EZEK|16|6|「我從你旁邊經過，見你在血中打滾，就對你說：『你雖在血中，卻要活下去！』我又說：『你雖在血中，卻要活下去！』
EZEK|16|7|我使你成長如田間所生長的；你就漸長，美而又美 ，兩乳成形，頭髮秀長，但你仍然赤身露體。
EZEK|16|8|「我從你旁邊經過看見你，看哪，正是你渴慕愛情的時候，我就用我衣服的邊搭在你身上，遮蓋你的赤體；又向你起誓，與你立約，你就歸我。這是主耶和華說的。
EZEK|16|9|那時我用水洗你，洗淨你身上的血，又用油抹你。
EZEK|16|10|我使你身穿錦繡衣裳，腳穿海狗皮鞋，用細麻布裹著你，精緻衣料披在你身上。
EZEK|16|11|我用首飾打扮你：我把手鐲戴在你手上，項鏈在你頸上，
EZEK|16|12|我也把環子戴在你鼻上，耳環在你耳上，華冠在你頭上。
EZEK|16|13|這樣，你就有金銀的首飾，穿的是細麻衣和精緻衣料，以及錦繡衣裳；吃的是細麵、蜂蜜和油。你也極其美貌，配登王后之位。
EZEK|16|14|你美貌的名聲傳到列國，因我加給你榮華，使你完美。這是主耶和華說的。
EZEK|16|15|「只是你仗著自己美貌，又憑著你的名聲行淫。你向路人縱情淫亂，你的美貌就屬於他的了 。
EZEK|16|16|你拿你的衣服為自己做成彩色丘壇，在其上行淫。這樣的事本不該有，以後也不該發生。
EZEK|16|17|你拿我所賜給你的那些美麗的金銀寶物，為自己製造男性的偶像，與它們行淫；
EZEK|16|18|你拿你的錦繡衣裳為它們披上，把我的膏油和香料擺在它們面前；
EZEK|16|19|你把我賜給你的食物，就是我賜給你享用的細麵、油和蜂蜜，都擺在它們面前作為馨香的供物。事情就是這樣。這是主耶和華說的。
EZEK|16|20|你拿你為我所生的兒女獻給它們吞噬。你的淫亂豈是小事？
EZEK|16|21|你竟把我的兒女殺了，使他們經火獻給它們！
EZEK|16|22|你做這一切可憎和淫亂的事，並未追念你幼年的日子，那時你赤身露體，在血中打滾。」
EZEK|16|23|「你有禍了！你有禍了！這是主耶和華說的。你做這一切惡事之後，
EZEK|16|24|又為自己建造土墩，在各廣場上築起高臺。
EZEK|16|25|你在各個街頭建造高臺，使你的美貌變為可憎；又向所有過路的人招手 ，多行淫亂。
EZEK|16|26|你也和你那放縱情慾的鄰邦 埃及 人行淫，增添你的淫亂，惹我發怒。
EZEK|16|27|看哪，我伸手攻擊你，減少你的福分，卻將你交給恨惡你的 非利士 人 ，讓他們任意待你。他們為你的淫行也感到羞恥。
EZEK|16|28|你尚且不滿意，又與 亞述 人行淫，但與他們行淫之後，仍不滿足；
EZEK|16|29|於是你與那稱為貿易之地的 迦勒底 多行淫亂，即使這樣，你仍不滿足。
EZEK|16|30|「你的心何等脆弱！這是主耶和華說的。你做這一切事，都是不知羞恥的妓女所做的，
EZEK|16|31|在各個街頭建造土墩，在各廣場上築高臺；但你藐視行淫的賞金，又不像妓女。
EZEK|16|32|你這行淫的妻子啊，竟然接外人，替代丈夫。
EZEK|16|33|凡妓女都是得人贈禮，你反倒餽贈你所愛的人，倒貼他們，使他們從四圍來與你行淫。
EZEK|16|34|你的淫行與其他婦女相反，不是人要求與你行淫；是你給人賞金，不是人給你賞金；你是相反的。」
EZEK|16|35|「你這妓女啊，要聽耶和華的話。
EZEK|16|36|主耶和華如此說：因你放縱情慾，露出下體，與你所愛的行淫，因你敬拜一切可憎的偶像，就像 自己兒女的血獻給它們，
EZEK|16|37|所以，看哪，我要聚集所有與你交歡的情人，不論是你所愛的或你所恨的，聚集他們從四圍到你那裏來；我要在他們面前暴露你的下體，使他們看盡你的下體。
EZEK|16|38|我也要審判你，如審判淫婦和流人血的婦女一樣。我要在憤怒和妒忌中使流血的罪歸到你身上。
EZEK|16|39|我要把你交在他們手中；他們必拆毀你的土墩，毀壞你的高臺，剝去你的衣服，奪取你美麗的寶物，留下你赤身露體。
EZEK|16|40|他們必聚集眾人攻擊你，用石頭打死你，用刀劍刺透你，
EZEK|16|41|用火焚燒你的房屋，在許多婦女眼前審判你。我必使你不再行淫，你也不再給賞金。
EZEK|16|42|我止息了向你所發的憤怒，我的妒忌也離開了你；這樣，我就平靜，不再惱怒。
EZEK|16|43|因你不追念幼年的日子，反而在這一切的事上惹我發烈怒，所以，看哪，我必照你所做的報應在你頭上。在你一切可憎的事上，你不是還行了淫亂嗎？這是主耶和華說的。」
EZEK|16|44|「看哪，凡說俗語的必用這俗語攻擊你，說：『有其母必有其女。』
EZEK|16|45|你實在是你母親的女兒，厭棄丈夫和兒女；你也是你姊妹的姊妹，厭棄丈夫和兒女。你的母親是 赫 人，父親是 亞摩利 人。
EZEK|16|46|你的姊姊是 撒瑪利亞 ，她和她的女兒們住在你北邊；你的妹妹是 所多瑪 ，她和她的女兒們住在你南邊。
EZEK|16|47|你不只效法她們的行為，照她們可憎的事去做，不消多時 ，你所做的一切就比她們更惡。
EZEK|16|48|主耶和華說：我指著我的永生起誓，你的妹妹 所多瑪 與她的女兒們並未做你和你女兒們所做的事。
EZEK|16|49|看哪，你的妹妹 所多瑪 的罪孽是這樣：她和她的女兒們都驕傲，糧源充足，大享安逸，卻不扶持困苦和貧窮人的手。
EZEK|16|50|她們狂傲，在我面前做可憎的事，我看見了就把她們除掉。
EZEK|16|51|撒瑪利亞 所犯的罪不及你的一半，你所做可憎的事比她更多；比起你所做這一切可憎的事，你的姊妹倒顯為義。
EZEK|16|52|你既為你的姊妹辯護，就要擔當自己的羞辱。因你所犯的罪比她們更可憎，她們比你倒顯為義；你既使你的姊妹顯為義，就要抱愧，擔當自己的羞辱。」
EZEK|16|53|「我必使她們被擄的歸回，使 所多瑪 和她的女兒們、 撒瑪利亞 和她的女兒們，並與你一起被擄的都歸回；
EZEK|16|54|好使你擔當自己的羞辱，為所做的一切抱愧，讓她們得到安慰。
EZEK|16|55|你的妹妹 所多瑪 和她的女兒們必回復原狀； 撒瑪利亞 和她的女兒們必回復原狀；你和你的女兒們也必回復原狀。
EZEK|16|56|在你驕傲的日子，你的妹妹 所多瑪 豈不是你口中的笑柄嗎？
EZEK|16|57|在你的惡行顯露以前，那受了凌辱的 亞蘭 女兒們和 亞蘭 四圍 非利士 的女兒們，都在四圍藐視你。
EZEK|16|58|耶和華說：你的淫蕩和可憎之事，你自己要擔當。」
EZEK|16|59|「主耶和華如此說：你這輕看誓言而背約的，我必照你所做的報應你。
EZEK|16|60|然而我要追念在你幼年時我與你所立的約，也要與你立定永約。
EZEK|16|61|當你接納你的姊姊和妹妹時，你要追念你所行的，自覺慚愧；並且我要將她們賞給你做女兒，卻不是按著我與你所立的約。
EZEK|16|62|我要堅定與你所立的約，你就知道我是耶和華，
EZEK|16|63|使你在我赦免你一切惡行時，心中追念，自覺慚愧，又因羞辱就不再開口。這是主耶和華說的。」
EZEK|17|1|耶和華的話臨到我，說：
EZEK|17|2|「人子啊，你要向 以色列 家出謎語，設比喻，
EZEK|17|3|說，主耶和華如此說：有一隻大鷹，翅膀大，翎毛長，羽毛豐滿，色彩繽紛；牠飛到 黎巴嫩 ，啄去香柏樹梢，
EZEK|17|4|啄斷它頂端的嫩枝，叼到貿易之地，放在商業城中。
EZEK|17|5|牠又從這地取了一些種子，種在肥沃的田裏，栽於豐沛的水源旁，如種植柳樹。
EZEK|17|6|它漸漸生長，成為低矮蔓生的葡萄樹；樹枝伸向那鷹，根部在牠下面。這樣，它就長成了一棵葡萄樹，生出枝子，長出枝幹。
EZEK|17|7|「有一隻 大鷹，翅膀大，羽毛多。看哪，葡萄樹從栽種它的苗圃向這鷹伸出根來，長出枝子，期盼從牠得到澆灌。
EZEK|17|8|這棵樹栽於肥田豐沛的水源旁，原是為了生枝、結果，成為佳美的葡萄樹。
EZEK|17|9|你要說，主耶和華如此說：這棵葡萄樹豈能發旺呢？鷹豈不拔出它的根來，摘光它的果子，使它枯乾，連長出的嫩葉都枯萎了嗎？要把它連根拔除，並不需要費大力或動用許多人。
EZEK|17|10|看哪，葡萄樹雖然栽種了，豈能發旺呢？一經東風擊打，豈不全然枯乾了嗎？它必在生長的苗圃中枯乾了。」
EZEK|17|11|耶和華的話臨到我，說：
EZEK|17|12|「你要對那悖逆之家說：你們不知道這些事是甚麼意思嗎？你要這樣說，看哪， 巴比倫 王曾到 耶路撒冷 ，把其中的君王和官長帶到 巴比倫 去，
EZEK|17|13|又從 以色列 王室後裔中選取一人，與他立約，令他發誓，又擄走國中有勢力的人，
EZEK|17|14|使王國衰弱，不再強盛，只能靠守盟約方得生存。
EZEK|17|15|他卻背叛 巴比倫 王，差派使者前往 埃及 ，要求 埃及 人給他馬匹和許多人。他豈能亨通呢？這樣做的人豈能逃脫呢？他背了約豈能逃脫呢？
EZEK|17|16|主耶和華說：我指著我的永生起誓，他定要死在 巴比倫 ，就是 巴比倫 王所在之處；因為 巴比倫 王立他為王，他竟輕看向王所起的誓，背棄王與他所立的約。
EZEK|17|17|當敵人建土堆，築堡壘，要殲滅許多人時，法老雖有強大軍隊和大批人馬，在戰場上還是不能幫助他。
EZEK|17|18|他輕看誓言，背棄盟約，看哪，雖已投降 ，卻又做這一切的事，他必不能逃脫。
EZEK|17|19|所以主耶和華如此說：我指著我的永生起誓，他既輕看我的誓言，背棄我的約，我必使這罪歸到他頭上。
EZEK|17|20|我要把我的網撒在他身上，他就被我的羅網纏住。我要帶他到 巴比倫 ，在那裏因他背叛我的罪懲罰他。
EZEK|17|21|所有逃跑的 軍隊必倒在刀下；剩餘的也必分散四方 。你們就知道說這話的是我─耶和華。」
EZEK|17|22|主耶和華如此說：「我要從香柏樹高高的樹梢摘取並栽上，從頂端的嫩枝中折下一嫩枝，栽於極高的山上，
EZEK|17|23|栽在 以色列 高處的山上。它就生枝、結果，成為高大的香柏樹，各類飛禽中的鳥都來宿在其下，宿在枝子的蔭下 。
EZEK|17|24|田野的樹木因此就知道是我─耶和華使高樹矮小，使矮樹高大，使綠樹枯乾，使枯樹發旺。我─耶和華說了這話，就必成就。」
EZEK|18|1|耶和華的話又臨到我，說：
EZEK|18|2|「你們在 以色列 地何以有這俗語，『父親吃了酸葡萄，兒子牙齒就酸倒』呢？
EZEK|18|3|主耶和華說：我指著我的永生起誓，你們在 以色列 必不再引用這俗語。
EZEK|18|4|看哪，所有的生命都是屬我的；父親的生命怎樣屬我，兒子的生命也照樣屬我；然而犯罪的，他必定死。
EZEK|18|5|「人若是公義，行公平公義的事：
EZEK|18|6|未曾在山上吃祭物，未曾向 以色列 家的偶像舉目；未曾污辱鄰舍的妻，也未曾在婦人的經期間親近她；
EZEK|18|7|未曾虧負人，而是將欠債之人的抵押品還給他；未曾搶奪人的物件，卻把食物給飢餓的人吃，把衣服給赤身的人穿；
EZEK|18|8|未曾向人取利息，也未曾索取高利，反倒縮手不作惡，在人與人之間施行誠實的判斷；
EZEK|18|9|遵行我的律例，謹守我的典章，按誠實行事 ；這人是公義的，必要存活。這是主耶和華說的。
EZEK|18|10|「他若生了兒子，兒子作強盜，流人的血，作父親的 雖然未犯此過，兒子卻對弟兄 行了以上所說的惡，在山上吃祭物，污辱鄰舍的妻；
EZEK|18|11|
EZEK|18|12|虧負困苦和貧窮的人，搶奪別人的物件，不歸還抵押品，卻向偶像舉目，做可憎的事；
EZEK|18|13|向人取利息，索取高利，這人豈能存活呢？他不能存活。他因做這一切可憎的事，必要死亡，他的血要歸到自己身上。
EZEK|18|14|「看哪，他若生了兒子，兒子見父親所犯的一切罪，他見了，卻不照樣去做；
EZEK|18|15|他未曾在山上吃祭物，未曾向 以色列 家的偶像舉目，未曾污辱鄰舍的妻；
EZEK|18|16|也未曾虧負人，未曾取人的抵押品，未曾搶奪人的物件，卻把食物給飢餓的人吃，把衣服給赤身的人穿，
EZEK|18|17|縮手不害困苦人，未曾向人索取利息或高利；反倒順從我的典章，遵行我的律例；如此，他必不因父親的罪孽死亡，定要存活。
EZEK|18|18|至於他父親，因為施行欺壓，搶奪弟兄，在百姓中行不善，看哪，他必因自己的罪孽死亡。
EZEK|18|19|「你們還說：『兒子為甚麼不擔當父親的罪孽呢？』兒子若行公平公義的事，謹守遵行我一切的律例，他必要存活。
EZEK|18|20|惟有犯罪的，卻必死亡。兒子不擔當父親的罪孽，父親也不擔當兒子的罪孽。義人的善果要歸自己，惡人的惡報也要歸自己。
EZEK|18|21|「惡人若回轉離開所做的一切罪惡，謹守我的一切律例，行公平公義的事，他必要存活，不致死亡。
EZEK|18|22|他所犯的一切罪過都不被記念；他因所行的義，必要存活。
EZEK|18|23|惡人死亡，豈是我所喜悅的呢？我豈不是喜悅他回轉離開所行的道而存活嗎？這是主耶和華說的。
EZEK|18|24|至於義人，他若轉離義行而作惡，照著惡人所做一切可憎的事去做，豈能存活呢？他所行的一切義都不被記念；反而因所行的惡、所犯的罪死亡。
EZEK|18|25|「你們卻說：『主的道不公平！』 以色列 家啊，你們要聽，我的道不公平嗎？你們的道不是不公平嗎？
EZEK|18|26|義人若轉離義行而作惡，他就因這些惡而死亡。他要死在他所作的惡中。
EZEK|18|27|惡人若回轉離開所行的惡，行公平公義的事，他必救自己的命；
EZEK|18|28|因為他省察，回轉離開所犯的一切罪過，他必要存活，不致死亡。
EZEK|18|29|以色列 家還說：『主的道不公平！』 以色列 家啊，我的道不公平嗎？你們的道不是不公平嗎？
EZEK|18|30|所以， 以色列 家啊，我必按你們各人所做的審判你們。當回轉，回轉離開你們一切的罪過，免得罪孽成為你們的絆腳石。這是主耶和華說的。
EZEK|18|31|你們要把所犯的一切罪過盡行拋棄，為自己造一個新的心和新的靈。 以色列 家啊，你們為甚麼要死呢？
EZEK|18|32|我不喜歡有任何人死亡，所以你們當回轉，要存活！這是主耶和華說的。」
EZEK|19|1|你當為 以色列 的領袖們唱哀歌，
EZEK|19|2|說： 你的母親在獅子中 是怎樣的母獅呢？ 牠蹲伏在少壯獅子中， 養育小獅子。
EZEK|19|3|牠養大了其中一隻小獅子， 成了少壯獅子， 學會抓食， 牠就吃人。
EZEK|19|4|列國聽見了就把牠逮住在他們的坑裏， 用鉤子拉牠到 埃及 地去。
EZEK|19|5|母獅見自己等候， 期望落空， 就從小獅子中取一隻 ， 養為少壯獅子；
EZEK|19|6|牠在眾獅子中徜徉， 長大成為少壯獅子， 學會抓食， 牠就吃人。
EZEK|19|7|牠拆毀他們的宮殿 ， 使他們的城鎮變為廢墟； 因牠咆哮的聲音， 遍地和其中所充滿的都荒廢了。
EZEK|19|8|於是四圍列國 從各省前來攻擊牠， 把網撒在牠身上， 把牠逮住在他們的坑裏。
EZEK|19|9|他們又用鉤子鉤住牠，把牠放入籠中， 帶到 巴比倫 王那裏， 把牠押進城堡， 以色列 山上就不再聽見牠的聲音。
EZEK|19|10|你的母親如葡萄樹， 在葡萄園中 ， 栽於水邊，因為水多， 就多結果子，多生枝子；
EZEK|19|11|它長出堅固的枝幹， 可作統治者的權杖。 這枝幹高舉在茂密的樹枝中， 可見樹身高大，枝子繁多。
EZEK|19|12|但在烈怒中它被拔出，摔在地上； 東風吹乾其果子， 那堅固的枝幹因折斷而枯乾， 被火燒燬；
EZEK|19|13|如今這葡萄樹移植於曠野， 在乾旱無水之地，
EZEK|19|14|火從枝幹中發出， 燒滅它的枝條和它的果子 ， 以致不再有堅固的枝幹， 可作統治者的權杖。 這是哀傷之歌，成為一首哀歌。
EZEK|20|1|第七年五月初十，有 以色列 的幾個長老前來求問耶和華，坐在我面前。
EZEK|20|2|耶和華的話臨到我，說：
EZEK|20|3|「人子啊，你要告訴 以色列 的長老，對他們說，主耶和華如此說：你們來是為求問我嗎？主耶和華說：我指著我的永生起誓，我必不讓你們求問。
EZEK|20|4|人子啊，你要審問他們嗎？你要審問嗎？你當使他們知道他們祖先那些可憎的事；
EZEK|20|5|你要對他們說，主耶和華如此說：當日我揀選 以色列 ，對 雅各 家的後裔起誓，在 埃及 地向他們顯現，起誓說：我是耶和華─你們的上帝；
EZEK|20|6|那日我向他們起誓，要領他們出 埃及 地，到我為他們所找到的流奶與蜜之地，就是全地中最美好之地。
EZEK|20|7|我對他們說，你們各人要拋棄眼中所喜愛的可憎之物，不可用 埃及 的偶像玷污自己。我是耶和華─你們的上帝。
EZEK|20|8|他們卻悖逆我，不肯聽從我，不拋棄他們眼中所喜愛的可憎之物，離棄 埃及 的偶像。 「我就說，在 埃及 地，我要把我的憤怒傾倒在他們身上，向他們發盡我的怒氣。
EZEK|20|9|我這麼做是為了我名的緣故，免得我的名在他們所居住之列國眼中被褻瀆；我曾在這些列國眼前向他們顯現，領他們出了 埃及 地。
EZEK|20|10|我領他們出 埃及 地，帶他們到曠野。
EZEK|20|11|我將我的律例賜給他們，將我的典章指示他們；人若遵行就必因此存活。
EZEK|20|12|我將我的安息日賜給他們，在我與他們中間作記號，讓他們知道我─耶和華是使他們分別為聖的。
EZEK|20|13|以色列 家卻在曠野中悖逆我，不順從我的律例，厭棄我的典章；人若遵行就必因此存活。他們卻大大干犯我的安息日。 「因此我說，我要在曠野把我的憤怒傾倒在他們身上，滅絕他們。
EZEK|20|14|我這麼做是為了我名的緣故，免得我的名在列國眼中被褻瀆，因為在這些列國眼前我領了他們出來。
EZEK|20|15|並且我在曠野向他們起誓，必不領他們進入我所賜的流奶與蜜之地，就是全地中最美好之地；
EZEK|20|16|因為他們厭棄我的典章，不順從我的律例，干犯我的安息日，他們的心隨從自己的偶像。
EZEK|20|17|雖然如此，我的眼仍顧惜他們，不毀滅他們，不在曠野把他們滅絕淨盡。
EZEK|20|18|「我在曠野對他們的兒女說：『不要遵行你們祖先的律例，不要謹守他們的規條，也不要用他們的偶像玷污自己。
EZEK|20|19|我是耶和華─你們的上帝，你們要順從我的律例，謹守遵行我的典章，
EZEK|20|20|且以我的安息日為聖。這日必在我與你們中間作記號，使你們知道我是耶和華─你們的上帝。』
EZEK|20|21|只是他們的兒女悖逆我，不順從我的律例，也不謹守遵行我的典章；人若遵行就必因此存活。他們卻干犯我的安息日。 「因此我說，我要在曠野把我的憤怒傾倒在他們身上，向他們發盡我的怒氣。
EZEK|20|22|但我卻縮手而未如此行；我這麼做是為了我名的緣故，免得我的名在列國眼中被褻瀆，因為在這些列國眼前我領了他們出來。
EZEK|20|23|並且我在曠野向他們起誓，要把他們驅散到列國，分散在列邦；
EZEK|20|24|因為他們不遵行我的典章，厭棄我的律例，干犯我的安息日，眼目向著他們祖先的偶像。
EZEK|20|25|我也任他們遵行那無益的律例，隨從那不能使人存活的規條。
EZEK|20|26|他們使所有頭生的經火，我就任憑他們在這供物上玷污自己；我令他們驚恐，他們就知道我是耶和華。
EZEK|20|27|「人子啊，你要告訴 以色列 家，對他們說，主耶和華如此說：你們的祖先在背叛我的事上再次褻瀆了我；
EZEK|20|28|我領他們到我起誓應許賜給他們的地，他們看見各高岡、各茂密的樹，就在那裏獻祭，獻上惹我發怒的供物，也在那裏焚燒馨香的祭，獻澆酒祭。
EZEK|20|29|我就對他們說：你們去的那丘壇叫甚麼呢？它名叫 巴麻 ，直到今日。
EZEK|20|30|所以你要對 以色列 家說，主耶和華如此說：你們仍要照你們祖先所做的玷污自己嗎？還要照他們可憎的事行淫嗎？
EZEK|20|31|當你們獻上供物，使你們兒子經火的時候，你們仍用各樣的偶像玷污自己，直到今日。 以色列 家啊，我豈能讓你們求問呢？主耶和華說：我指著我的永生起誓，我必不讓你們求問。
EZEK|20|32|「你們說：『我們要像列國和列邦的宗族一樣，去事奉木頭與石頭。』你們所起的心意萬不能成就。」
EZEK|20|33|「主耶和華說：我指著我的永生起誓，我要作王，用大能的手和伸出的膀臂，並傾倒出來的憤怒治理你們。
EZEK|20|34|我必用大能的手和伸出的膀臂，並傾倒出來的憤怒，把你們從萬民中領出來，從被趕散到的列邦聚集你們。
EZEK|20|35|我必帶你們到萬民的曠野，在那裏當面審判你們。
EZEK|20|36|我怎樣在 埃及 地的曠野審判你們的祖先，也必照樣審判你們。這是主耶和華說的。
EZEK|20|37|我要使你們從杖下經過，按著約的拘束 帶領你們。
EZEK|20|38|我必從你們中間除盡叛逆和得罪我的人；我將他們從所寄居的地方領出來，他們卻不得進入 以色列 地，你們就知道我是耶和華。
EZEK|20|39|「你們， 以色列 家啊，主耶和華如此說：你們若不聽從我，從今以後就讓各人去事奉他的偶像吧，只是不可再以你們的供物和偶像褻瀆我的聖名。
EZEK|20|40|「在我的聖山，就是 以色列 高處的山， 以色列 全家，那地所有的人，都要在那裏事奉我。在那裏我悅納他們，並要你們獻供物和初熟的土產，以及一切的聖物。這是主耶和華說的。
EZEK|20|41|我把你們從萬民中領出來，從被趕散到的列邦聚集你們，那時我必悅納你們如同悅納馨香之祭，我要在列國眼前，在你們中間顯為聖。
EZEK|20|42|我領你們進入 以色列 地，就是我起誓應許賜給你們列祖之地，那時你們就知道我是耶和華。
EZEK|20|43|你們在那裏要追念那玷污自己的所作所為，又要因所行的一切惡事厭惡自己。
EZEK|20|44|以色列 家啊，我為我名的緣故，沒有照著你們的惡行和你們的敗壞對待你們；你們就知道我是耶和華。這是主耶和華說的。」
EZEK|20|45|耶和華的話臨到我，說：
EZEK|20|46|「人子啊，你要面向南方，向南方傳講 ，向 尼革夫 田野的樹林說預言。
EZEK|20|47|你要對 尼革夫 的樹林說，要聽耶和華的話。主耶和華如此說：看哪，我要在你那裏點火，燒滅你們中間所有的綠樹和枯樹，猛烈的火焰必不熄滅；從南到北，人的臉都被燒焦。
EZEK|20|48|凡血肉之軀都知道是我─耶和華點了火，這火必不熄滅。」
EZEK|20|49|於是我說：「唉！主耶和華啊，人都指著我說：他不是說比喻的人嗎？」
EZEK|21|1|耶和華的話臨到我，說：
EZEK|21|2|「人子啊，把你的臉正對著 耶路撒冷 ，對著聖所 傳講 ，向 以色列 地說預言。
EZEK|21|3|你要向 以色列 地說，耶和華如此說：看哪，我與你為敵，拔刀出鞘，把義人和惡人從你中間剪除。
EZEK|21|4|因為我要剪除你當中的義人和惡人，所以我的刀要出鞘，從南到北攻擊所有的血肉之軀；
EZEK|21|5|凡血肉之軀都知道我─耶和華已拔刀出鞘，刀必不再入鞘。
EZEK|21|6|你，人子啊，要嘆息，在他們眼前斷了腰，愁苦地嘆息。
EZEK|21|7|若有人對你說：『你為甚麼嘆息呢？』你就說：『因為有風聲傳來，人心惶惶，雙手發軟，精神衰敗，膝弱如水。看哪，它臨近了，一定會發生。』這是主耶和華說的。」
EZEK|21|8|耶和華的話臨到我，說：
EZEK|21|9|「人子啊，你要預言說，耶和華如此吩咐，你要說： 有刀，刀已磨快， 又擦亮了；
EZEK|21|10|磨快為要大大殺戮， 擦亮為要像閃電。 我們豈能快樂呢？ 它藐視我兒的權杖和一切的木頭 。
EZEK|21|11|它已經交給人擦亮，可以掌握使用；這刀已經磨快擦亮，好交在行殺戮的人手中。
EZEK|21|12|人子啊，你要呼喊哀號，因為這刀將臨到我的百姓，臨到 以色列 所有的領袖身上。他們和我的百姓都要交在刀下，所以你要捶胸 。
EZEK|21|13|因為這是一個考驗，若它藐視權杖，也不算一回事，又怎麼樣呢？這是主耶和華說的。」
EZEK|21|14|「人子啊，你要拍掌預言，使這刀三番兩次臨到；這是致人死傷的刀，就是包圍人，使人大受死傷的刀。
EZEK|21|15|我設立這恐嚇 的刀，攻擊他們一切的城門，為要使他們的心驚慌害怕，許多人因而跌倒。唉！它 造得像閃電，磨得尖利 ，要行殺戮。
EZEK|21|16|刀啊，要行動一致 ，向右邊，或指向左邊；面向哪方，就向哪方。
EZEK|21|17|我也要拍掌，使我的憤怒平息。這是我─耶和華說的。」
EZEK|21|18|耶和華的話臨到我，說：
EZEK|21|19|「人子啊，你要畫定兩條路線，使 巴比倫 王的刀過來，這兩條路必從同一地分出來；要在通往城裏的路口畫手作指標。
EZEK|21|20|你要劃定一條路，使刀來到 亞捫 人的 拉巴 ，來到 猶大 ，在堅固城 耶路撒冷 。
EZEK|21|21|因為 巴比倫 王站在岔路上，在兩條路口占卜。他搖籤 求問神像，察看肝臟；
EZEK|21|22|右手是 耶路撒冷 的占卜，以便安設撞城槌，張口喊殺 ，揚聲呼叫，建土堆，築堡壘，以撞城槌攻打城門。
EZEK|21|23|在那些曾鄭重起誓的 猶大 人眼中，這是虛假的占卜；但 巴比倫 王要使他們想起自己的罪孽，以便俘擄他們。」
EZEK|21|24|於是，主耶和華如此說：「因你們的過犯顯露，你們的罪孽被記得，以致你們的罪惡在你們一切的行為上都彰顯出來；你們既被記得，就被擄在掌中。
EZEK|21|25|你這褻瀆行惡的 以色列 王啊，你的日子，最後懲罰的時刻已來臨。
EZEK|21|26|主耶和華如此說：當除掉榮冕，摘下華冠，景況已不復從前；要使卑者升為高，使高者降為卑。
EZEK|21|27|我要將這國傾覆，傾覆，再傾覆；這國必不存在，直等到那應得的人來到，我就將國賜給他。」
EZEK|21|28|「人子啊，你要說預言；你要說，論到 亞捫 人和他們的凌辱，主耶和華吩咐我如此說：有刀，拔出來的刀，已經擦亮，為了行殺戮；它亮如閃電以行吞滅。
EZEK|21|29|他們為你見虛假的異象，行謊詐的占卜，使你倒在褻瀆之惡人的頸項上；他們的日子，最後懲罰的時刻已來臨。
EZEK|21|30|你收刀入鞘吧！我要在你受造之處、生長之地懲罰你。
EZEK|21|31|我要把我的憤怒傾倒在你身上，把我烈怒的火噴在你身上；又將你交在善於殺滅、畜牲一般的人手中。
EZEK|21|32|你要成為火中之柴，你的血必在地裏；你必不再被記得，因為這是我─耶和華說的。」
EZEK|22|1|耶和華的話臨到我，說：
EZEK|22|2|「你，人子啊，你要審問，審問這流人血的城嗎？要使它知道它一切可憎的事。
EZEK|22|3|你要說，主耶和華如此說：那在其中流人血的城啊，它的時刻已到，它製造偶像玷污了自己。
EZEK|22|4|你因流了人的血，算為有罪；因所製造的偶像，玷污自己；你使你的日子臨近，你的年數已來到 。所以我使你承受列國的凌辱和列邦的譏誚。
EZEK|22|5|你這惡名昭彰、混亂的城啊，離你或遠或近的國家都必譏誚你。
EZEK|22|6|「看哪， 以色列 的領袖在你那裏，為了流人的血各逞其能。
EZEK|22|7|你那裏有輕慢父母的，在你當中有欺壓寄居者的，你那裏也有虧負孤兒寡婦的。
EZEK|22|8|你藐視我的聖物，干犯我的安息日。
EZEK|22|9|你那裏有為流人血而毀謗人的，你那裏有在山上吃祭物的，在你當中也有行淫亂的，
EZEK|22|10|有露父親下體的 ，有玷辱經期中不潔淨之婦人的。
EZEK|22|11|這人與鄰舍的妻子行可憎的事，那人行淫污辱媳婦，在你那裏還有人污辱他的姊妹，父親的女兒。
EZEK|22|12|你那裏有收取報酬而流人血的。你取利息，又索取高利；欺壓鄰舍，奪取財物；你竟然忘了我。這是主耶和華說的。
EZEK|22|13|「看哪，我因你所得不義之財和你們中間所流的血，就擊打手掌。
EZEK|22|14|到了我對付你的日子，你的心豈能忍受呢？你的手還能有力嗎？我─耶和華說了這話，就必成就。
EZEK|22|15|我要把你驅散到列國，分散在列邦。我也必除掉你們中間的污穢。
EZEK|22|16|你在列國眼前因自己所做的被侮辱 ，你就知道我是耶和華。」
EZEK|22|17|耶和華的話臨到我，說：
EZEK|22|18|「人子啊，我看 以色列 家為渣滓。他們是爐中的銅、錫、鐵、鉛，是煉銀的渣滓 。
EZEK|22|19|所以主耶和華如此說：因你們全都成為渣滓，所以，看哪，我必將你們聚集在 耶路撒冷 中。
EZEK|22|20|人怎樣把銀、銅、鐵、鉛、錫聚在爐中，吹火使它鎔化；照樣，我也要在我的怒氣和憤怒中聚集你們，把你們安置在城中，使你們鎔化。
EZEK|22|21|我必聚集你們，把我烈怒的火吹在你們身上，你們就在其中鎔化。
EZEK|22|22|銀子怎樣在爐中鎔化，你們也必照樣在城中鎔化，因此就知道是我─耶和華把憤怒傾倒在你們身上。」
EZEK|22|23|耶和華的話臨到我，說：
EZEK|22|24|「人子啊，你要向這地說：你是未被潔淨 之地，在我盛怒的日子，沒有雨水在其上。
EZEK|22|25|其中的先知同謀背叛 ，如咆哮的獅子抓撕掠物。他們吞滅人命，搶奪財寶，使這地寡婦增多。
EZEK|22|26|其中的祭司曲解我的律法，褻瀆我的聖物，不分別聖與俗，也不使人分辨潔淨和不潔淨，又遮眼不顧我的安息日；在他們中間連我也被褻慢了。
EZEK|22|27|其中的領袖彷彿野狼抓撕掠物，流人的血，傷害人命，為得不義之財。
EZEK|22|28|其中的先知為他們粉刷，見虛假的異象，行謊詐的占卜，說：『主耶和華如此說』，其實耶和華並沒有說。
EZEK|22|29|這地的百姓慣行欺壓搶奪之事，虧負困苦和貧窮的人，欺壓寄居者，沒有公平。
EZEK|22|30|我在他們中間尋找一人重修城牆，在我面前為這地站在缺口上，使我不致滅絕它，卻連一個也找不著。
EZEK|22|31|所以我把憤怒傾倒在他們身上，用烈怒之火消滅他們，照他們所做的報應在他們頭上。這是主耶和華說的。」
EZEK|23|1|耶和華的話臨到我，說：
EZEK|23|2|「人子啊，有兩個女子，是一母所生，
EZEK|23|3|她們在 埃及 行淫，年少時就開始行淫；在那裏任人擁抱胸懷，撫弄她們少女的乳房。
EZEK|23|4|她們的名字，大的叫 阿荷拉 ，妹妹叫 阿荷利巴 。她們都歸於我，生了兒女。論到她們的名字， 阿荷拉 是 撒瑪利亞 ， 阿荷利巴 是 耶路撒冷 。
EZEK|23|5|「 阿荷拉 歸我之後卻仍行淫，戀慕所愛的人，就是 亞述 人，都是戰士 ，
EZEK|23|6|穿著藍衣，作省長、副省長，全都是俊美的年輕人，騎著馬的騎士。
EZEK|23|7|阿荷拉 與 亞述 人中所有的美男子放縱淫行，她因拜所戀慕之人的一切偶像，玷污了自己。
EZEK|23|8|她從 埃及 的時候，就沒有離開過淫亂；因為她年輕時，有人與她同寢，撫弄她少女的乳房，和她縱慾行淫。
EZEK|23|9|因此，我把她交在她所愛的人手中，就是她所戀慕的 亞述 人手中。
EZEK|23|10|他們暴露她的下體，擄掠她的兒女，用刀殺了她；他們向她施行審判，使她在婦女中留下臭名。
EZEK|23|11|「她妹妹 阿荷利巴 雖然看見了，卻還是縱慾，比姊姊更加腐敗，行淫亂比姊姊更甚。
EZEK|23|12|她戀慕 亞述 人，就是省長和副省長，披掛整齊的戰士，騎著馬的騎士，全都是俊美的年輕人。
EZEK|23|13|我看見她被污辱，姊妹二人同行一路。
EZEK|23|14|阿荷利巴 又加增淫行，她看見牆上刻有人像，就是鮮紅色的 迦勒底 人雕刻的像。
EZEK|23|15|它們腰間繫著帶子，頭上有飄揚的裹頭巾，都是將軍的樣子， 巴比倫 人的形像； 迦勒底 是他們的出生地。
EZEK|23|16|阿荷利巴 一看見就戀慕他們，派遣使者往 迦勒底 他們那裏去。
EZEK|23|17|巴比倫 人來到她那裏，上了她愛情的床，與她行淫污辱她。她被污辱，隨後她的心卻與他們生疏。
EZEK|23|18|這樣，她既暴露淫行，暴露下體；我的心就與她生疏，像先前與她的姊姊生疏一樣。
EZEK|23|19|她仍繼續增添淫行，追念她年輕時在 埃及 地行淫的日子，
EZEK|23|20|戀慕情人的身壯精足，如驢似馬。
EZEK|23|21|這樣，你就渴望年輕時的淫蕩；那時， 埃及 人因你年輕時的胸懷，撫弄你的乳房 。」
EZEK|23|22|阿荷利巴 啊，主耶和華如此說：「看哪，我要激起先前你喜愛，而後生疏的人前來攻擊你。我必使他們前來，在你四圍攻擊你；
EZEK|23|23|有 巴比倫 人、 迦勒底 眾人、 比割 人、 書亞 人、 哥亞 人，還有 亞述 眾人與他們一起，都是俊美的年輕人。他們是省長、副省長、將軍、有名聲的，全都騎著馬。
EZEK|23|24|他們用兵器、 戰車、輜重車，率領大軍前來攻擊你。他們要拿大小盾牌，戴著頭盔，在你四圍擺陣攻擊你。我要把審判交給他們，他們必按著自己的規條審判你。
EZEK|23|25|我要向你傾洩我的妒忌，使他們以憤怒對待你。他們必割去你的鼻子和耳朵，你剩餘的人必倒在刀下。他們必擄去你的兒女，你所剩餘的必被火焚燒。
EZEK|23|26|他們必剝去你的衣服，奪取你美麗的寶物。
EZEK|23|27|這樣，我必止息你的淫行和你從 埃及 地就開始犯的淫亂，使你不再仰望 亞述 ，也不再追念 埃及 。
EZEK|23|28|主耶和華如此說：看哪，我必把你交在你所恨惡的人手中，就是你心與他生疏的人手中。
EZEK|23|29|他們要以恨惡對待你，奪取你勞碌得來的一切，留下你赤身露體。你淫亂的下體，連你的淫行和淫蕩，都必顯露。
EZEK|23|30|人必向你行這些事；因為你隨從外邦人行淫，用他們的偶像玷污自己。
EZEK|23|31|你走了你姊姊的路，所以我必把她的杯交在你的手中。」
EZEK|23|32|主耶和華如此說： 「你必喝你姊姊的杯， 那杯又深又廣， 盛得很多， 使你遭受嗤笑譏刺。
EZEK|23|33|你必酩酊大醉， 滿有愁苦。 你姊姊 撒瑪利亞 的杯， 驚駭和淒涼的杯，
EZEK|23|34|你必喝它，並且喝乾。 甚至咀嚼杯片， 撕裂自己的胸脯； 因為我曾說過。 這是主耶和華說的。」
EZEK|23|35|主耶和華如此說：「因你忘記我，將我丟在背後，所以你要擔當你的淫行和淫蕩。」
EZEK|23|36|耶和華對我說：「人子啊，你要審問 阿荷拉 與 阿荷利巴 嗎？要指出她們所做可憎的事。
EZEK|23|37|她們行姦淫，手中有血。她們與偶像行姦淫，使她們為我所生的兒女經火，給它們當食物。
EZEK|23|38|此外，她們還向我這樣做：同一天又玷污我的聖所，干犯我的安息日。
EZEK|23|39|她們殺了兒女獻給偶像，當天又進入我的聖所，褻瀆了它。看哪，這就是她們在我殿中所做的。
EZEK|23|40|「況且你們兩姊妹派人從遠方召人來。使者到了他們那裏，看哪，他們就來了。為了他們，你們沐浴，畫眼影，佩戴首飾，
EZEK|23|41|坐在華美的床上，前面擺設桌子，把我的香料和膏油放在其上。
EZEK|23|42|在那裏有一群人歡樂的聲音；有許多的平民，從曠野來的醉漢 ，把鐲子戴在她們手上，把華冠戴在她們頭上。
EZEK|23|43|「我論到這久行姦淫而色衰的婦人說：現在人們還要與她行淫，她也要與人行淫。
EZEK|23|44|人去到 阿荷拉 和 阿荷利巴 二淫婦那裏 ，好像與妓女行淫。
EZEK|23|45|義人必按照審判淫婦和流人血之婦人的規條，審判她們；因為她們是淫婦，她們的手中有血。」
EZEK|23|46|主耶和華如此說：「我要讓軍隊上來攻擊她們，使她們驚駭，成為擄物。
EZEK|23|47|這軍隊必用石頭打死她們，用刀劍殺害她們，又殺戮她們的兒女，用火焚燒她們的房屋。
EZEK|23|48|我必使這地不再有淫行，所有的婦女都受警戒，不再效法你們的淫行 。
EZEK|23|49|人必因你們的淫行報應你們；你們要擔當拜偶像的罪，因此你們就知道我是主耶和華。」
EZEK|24|1|第九年十月初十，耶和華的話臨到我，說：
EZEK|24|2|「人子啊，你要記錄這一天的名稱，這特別的一天， 巴比倫 王圍困 耶路撒冷 ，就在這特別的一天。
EZEK|24|3|你要向這悖逆之家設比喻，對他們說，主耶和華如此說： 把鍋放在火上， 放好了，倒水在其中；
EZEK|24|4|要將肉塊，一切肥美的肉塊， 腿和肩都放在鍋裏， 要裝滿上等的骨頭；
EZEK|24|5|要取羊群中最好的， 把柴 堆在下面， 把它煮開， 骨頭煮在其中。
EZEK|24|6|「主耶和華如此說：禍哉！這流人血的城，就是長銹的鍋。它的銹未曾除掉，要將肉塊從其中一一取出，不必抽籤。
EZEK|24|7|這城所流的血還在城中，血倒在光滑的磐石上，沒有倒在地上，用土掩蓋；
EZEK|24|8|是我使這城所流的血倒在光滑的磐石上，不得掩蓋，為要惹動憤怒，施行報應。
EZEK|24|9|所以主耶和華如此說：禍哉！這流人血的城，我必親自加大柴堆。
EZEK|24|10|你要添上木柴，使火著旺，將肉煮爛，加上香料 ，烤焦骨頭；
EZEK|24|11|你要把空鍋放在炭火上，將鍋燒熱，把銅燒紅，鎔化其中的污穢，除淨其上的銹。
EZEK|24|12|然而這一切勞碌無效 ，它厚厚的銹，即使用火也除不掉。
EZEK|24|13|雖然我想潔淨你污穢的淫行，你卻不潔淨，你的污穢再也不能潔淨，直等我止息了向你發的憤怒。
EZEK|24|14|我─耶和華說了這話，時候到了，就必成就；必不退縮，不顧惜，也不憐憫。人必照你的所作所為審判你。這是主耶和華說的。」
EZEK|24|15|耶和華的話臨到我，說：
EZEK|24|16|「人子，看哪，我要以災病奪取你眼中所喜愛的，你卻不可悲哀哭泣，也不可流淚，
EZEK|24|17|只可嘆息，不可出聲，不可辦理喪事；裹上頭巾，腳上穿鞋，不可摀著鬍鬚，也不可吃一般人的食物 。」
EZEK|24|18|到了早晨我把這事告訴百姓，晚上我的妻子就死了。次日早晨我就遵命而行。
EZEK|24|19|百姓對我說：「你這樣做跟我們有甚麼關係，你不告訴我們嗎？」
EZEK|24|20|我對他們說：「耶和華的話臨到我，說：
EZEK|24|21|『你告訴 以色列 家，主耶和華如此說：我要使我的聖所被褻瀆，就是你們憑勢力所誇耀、眼裏所喜愛、心中所愛惜的；並且你們所遺留的兒女必倒在刀下。
EZEK|24|22|那時，你們要照我所做的去做。你們不可摀著鬍鬚，也不可吃一般人的食物。
EZEK|24|23|你們頭要裹上頭巾，腳要穿上鞋；不可悲哀哭泣。你們必因自己的罪孽衰殘，相對嘆息。
EZEK|24|24|以西結 必這樣成為你們的預兆；凡他所做的，你們也必照樣做。那事來到，你們就知道我是主耶和華。』」
EZEK|24|25|「你，人子啊，那日當我除掉他們所倚靠的保障、所歡喜的榮耀，並眼中所喜愛的，心裏所重看的兒女時，
EZEK|24|26|逃脫的人豈不來到你這裏，使你耳聞這事嗎？
EZEK|24|27|那日你要向逃脫的人開口說話，不再啞口無言。你必這樣成為他們的預兆，他們就知道我是耶和華。」
EZEK|25|1|耶和華的話臨到我，說：
EZEK|25|2|「人子啊，你要面向 亞捫 人說預言，攻擊他們。
EZEK|25|3|你要對 亞捫 人說，當聽主耶和華的話。主耶和華如此說：我的聖所遭褻瀆， 以色列 地變荒涼， 猶大 家被擄掠；那時，你因這些事說『啊哈』，
EZEK|25|4|所以，看哪，我要把你交給東方人為業；他們必在你中間安營居住，設立居所，吃你的果子，喝你的奶。
EZEK|25|5|我必使 拉巴 成為牧放駱駝之地，使 亞捫 成為羊群躺臥之處，你們就知道我是耶和華。
EZEK|25|6|主耶和華如此說：因你們拍手頓足，幸災樂禍，藐視 以色列 地，
EZEK|25|7|所以，看哪，我要伸手攻擊你，把你交給列國作為擄物。我必從萬民中剪除你，從列邦中消滅你。我必除滅你，你就知道我是耶和華。」
EZEK|25|8|「主耶和華如此說：因 摩押 和 西珥 人說『看哪， 猶大 家與列國無異』，
EZEK|25|9|所以，看哪，我要破開 摩押 邊界的城鎮，就是 摩押 人所誇耀的城鎮， 伯‧耶施末 、 巴力‧免 、 基列亭 ，
EZEK|25|10|令東方人前來攻擊 亞捫 人。我必將 亞捫 交給他們為業，使 亞捫 人在列國中不再被記念。
EZEK|25|11|我也必向 摩押 施行審判，他們就知道我是耶和華。」
EZEK|25|12|「主耶和華如此說：因為 以東 向 猶大 家報仇，因向他們報仇而大大顯為有罪，
EZEK|25|13|所以主耶和華如此說：我要伸手攻擊 以東 ，將人與牲畜剪除，使 以東 從 提幔 起，直到 底但 ，地變荒涼，人也都倒在刀下。
EZEK|25|14|我要藉我子民 以色列 的手報復 以東 ；他們必照我的怒氣，按我的憤怒對待 以東 ， 以東 人就知道施報的是我。這是主耶和華說的。」
EZEK|25|15|「主耶和華如此說：因 非利士 人報仇，就是心存輕蔑報仇；他們永懷仇恨，意圖毀滅，
EZEK|25|16|所以主耶和華如此說：看哪，我要伸手攻擊 非利士 人，剪除 基利提 人，滅絕沿海剩餘的居民。
EZEK|25|17|我要大大報復他們，發怒斥責他們。我報復他們的時候，他們就知道我是耶和華。」
EZEK|26|1|第十一年某月初一，耶和華的話臨到我，說：
EZEK|26|2|「人子啊，因 推羅 向 耶路撒冷 說：『啊哈！那眾民之門已經破壞，向我敞開；它既變為廢墟，我必豐盛。』
EZEK|26|3|所以，主耶和華如此說： 推羅 ，看哪，我與你為敵，使許多國家湧上攻擊你，如同海洋使波浪湧上一樣。
EZEK|26|4|他們要破壞 推羅 的城牆，拆毀它的城樓。我也要刮淨它的塵土，使它成為光滑的磐石。
EZEK|26|5|推羅 必成為海中的曬網場，因為我曾說過， 這是主耶和華說的。它必成為列國的擄物，
EZEK|26|6|推羅 鄉間鄰近的城鎮 必遭刀劍滅絕，他們就知道我是耶和華。」
EZEK|26|7|主耶和華如此說：「看哪，我必使諸王之王，就是 巴比倫 王 尼布甲尼撒 ，率領馬匹、戰車、騎兵、軍隊和許多人從北方來攻擊 推羅 。
EZEK|26|8|他必用刀劍殺滅你鄉間鄰近的城鎮，也必築堡壘，建土堆，舉盾牌攻擊你。
EZEK|26|9|他要安設撞城槌攻破你的城牆，以刀劍拆毀你的城樓。
EZEK|26|10|因他馬匹眾多，塵土必揚起遮蔽你。他進入你的城門，如同進入已有缺口之城。那時，你的城牆必因騎兵、車輪和戰車的響聲震動。
EZEK|26|11|他的馬蹄必踐踏你所有的街道；他必用刀劍殺戮你的居民。你堅固的柱子 必倒在地上。
EZEK|26|12|人必擄獲你的財寶，掠奪你的貨財；他們要破壞你的城牆，拆毀你華美的房屋，將你的石頭、木頭、塵土都拋在水中。
EZEK|26|13|我要使你唱歌的聲音止息；人不再聽見你彈琴的聲音。
EZEK|26|14|我必使你成為光滑的磐石，作曬網的場所。你不得再被建造，因為我─耶和華已這樣說了。這是主耶和華說的。」
EZEK|26|15|主耶和華對 推羅 如此說：「在你中間行殺戮，受傷的人唉哼時，海島豈不都因你傾倒的響聲震動嗎？
EZEK|26|16|那時沿海的君王都要從寶座下來，除去朝服，脫下錦衣，披上戰兢，坐在地上，不停發抖，為你而驚駭。
EZEK|26|17|他們必為你作哀歌，向你說： 『你這聞名之城， 航海之人居住， 海上最為堅固的， 你和居民使所有住在沿海的人 無不驚恐， 現在竟然毀滅了！
EZEK|26|18|如今在你傾覆的日子， 海島都要戰兢； 海中的群島見你歸於無有 就都驚惶。』」
EZEK|26|19|主耶和華如此說：「 推羅 啊 ，我要使你變為荒涼，如無人居住的城鎮；又使深水漫過你，大水淹沒你。
EZEK|26|20|那時，我要使你和下到地府的人同去，到古時候的人那裏；我要使你和下到地府的人一同住在地的深處，在久已荒廢的地方，使你那裏不再有人居住；我要在活人之地顯榮耀 。
EZEK|26|21|我必叫你令人驚恐，使你不再存留於世；人雖尋找你，卻永不尋見。這是主耶和華說的。」
EZEK|27|1|耶和華的話臨到我，說：
EZEK|27|2|「人子啊，要為 推羅 作哀歌。
EZEK|27|3|你要對位於海口，跟許多海島的百姓做生意的 推羅 說，主耶和華如此說： 推羅 啊，你曾說： 『我全然美麗。』
EZEK|27|4|你的疆界在海的中心， 造你的使你全然美麗。
EZEK|27|5|他們用 示尼珥 的松樹作你的甲板， 用 黎巴嫩 的香柏樹作桅杆，
EZEK|27|6|用 巴珊 的橡樹作你的槳， 用鑲嵌象牙的 基提 海島黃楊木 為艙板。
EZEK|27|7|你的帆是用 埃及 繡花細麻布做的， 可作你的大旗； 你的篷是用 以利沙島 的藍色和紫色布做的。
EZEK|27|8|西頓 和 亞發 的居民為你划槳； 推羅 啊，你們中間的智慧人為你掌舵。
EZEK|27|9|迦巴勒 的長者和智者 在你中間修補裂縫； 海上一切的船隻和水手 都在你那裏進行貨物交易。
EZEK|27|10|「 波斯 人、 路德 人、 弗 人在你的軍營中作戰士；他們在你們中間懸掛盾牌和頭盔，彰顯你的尊榮。
EZEK|27|11|亞發 人和你的軍隊都駐守在四圍的城牆上，你的城樓上也有勇士；他們懸掛盾牌，成全你的美麗。
EZEK|27|12|「 他施 因你多有財物，就作你的客商，他們帶著銀、鐵、錫、鉛前來換你的商品。
EZEK|27|13|雅完 、 土巴 、 米設 都與你交易，以人口和銅器換你的貨物。
EZEK|27|14|陀迦瑪 族用馬匹、戰馬和騾子換你的商品。
EZEK|27|15|底但 人與你交易，許多海島成為你的碼頭；他們拿象牙、黑檀木與你交換。
EZEK|27|16|亞蘭 因你貨品充裕，就作你的客商；他們用綠寶石、紫色布、刺繡、細麻布、珊瑚、紅寶石換你的商品。
EZEK|27|17|猶大 和 以色列 地都與你交易；他們用 米匿 的小麥、餅、蜜、油、乳香換你的貨物。
EZEK|27|18|大馬士革 也因你貨品充裕，多有各類財物，就帶來 黑本 酒和白羊毛與你交易。
EZEK|27|19|威但 和從 烏薩 來的 雅完 人 為了你的貨物，以加工的鐵、桂皮、香菖蒲換你的商品。
EZEK|27|20|底但 以騎馬用的座墊毯子與你交換。
EZEK|27|21|阿拉伯 和 基達 所有的領袖都作你的客商，用羔羊、公綿羊、公山羊與你交換。
EZEK|27|22|示巴 和 拉瑪 的商人也來與你交易，他們用各類上好的香料、各類的寶石和黃金換你的商品。
EZEK|27|23|哈蘭 、 干尼 、 伊甸 、 示巴 商人、 亞述 和 基抹 都與你交易。
EZEK|27|24|這些商人將美好的貨物包在藍色的繡花包袱內，又將華麗的衣服裝在香柏木的箱子裏，用繩索捆著，以此與你交易 。
EZEK|27|25|他施 的船隻為你運貨， 你在海中滿載貨物，極其沉重。
EZEK|27|26|划槳的把你划到水深之處， 東風在海中將你擊破。
EZEK|27|27|你的財寶、商品、貨物、 水手、掌舵的、 修補船縫的、進行貨物交易的， 並你那裏所有的戰士 和你中間所有的軍隊， 在你傾覆的日子都必沉在海底。
EZEK|27|28|因掌舵者的呼聲， 郊野就必震動。
EZEK|27|29|所有划槳的 都從他們的船下來； 水手和所有在海上掌舵的， 都要登岸。
EZEK|27|30|他們必為你放聲痛哭， 撒塵土於頭上， 在灰中打滾；
EZEK|27|31|又為你使頭光禿， 用麻布束腰， 號咷痛哭， 痛苦至極。
EZEK|27|32|他們哀號的時候， 為你作哀歌， 為你痛哭： 有何城如 推羅 ， 在海中沉寂呢？
EZEK|27|33|你由海上運出商品， 使許多民族充裕； 你以許多財寶貨物 令地上的君王豐富。
EZEK|27|34|在深水中被海浪打破的時候， 你的貨物和你中間所有的軍隊都下沉。
EZEK|27|35|海島所有的居民為你驚奇， 他們的君王都甚恐慌，面帶愁容。
EZEK|27|36|萬民中的商人向你發噓聲； 你令人驚恐， 不再存留於世，直到永遠。」
EZEK|28|1|耶和華的話臨到我，說：
EZEK|28|2|「人子啊，你要對 推羅 的君王說，主耶和華如此說： 你心裏高傲，說：『我是神明； 我在海中坐諸神之位。』 雖然你把你的心比作神明的心， 你卻不過是人，並不是神明！
EZEK|28|3|看哪，你比 但以理 更有智慧， 任何祕密都不能向你隱藏。
EZEK|28|4|你靠自己的智慧聰明得了財寶， 把金銀收入庫房；
EZEK|28|5|你靠自己的大智慧以貿易增添財寶， 又因你的財寶心裏高傲；
EZEK|28|6|所以主耶和華如此說： 因你把你的心比作神明的心，
EZEK|28|7|所以，看哪，我必使外國人， 就是列國中兇暴的人臨到你這裏； 他們要拔刀摧毀你用智慧得來的美物， 污損你的榮光。
EZEK|28|8|他們必使你墜入地府； 你要像被刺殺之人的死，死在海中。
EZEK|28|9|在殺你的人面前， 你還能說『我是神明』嗎？ 在殺害你的人手中， 你不過是人，並不是神明。
EZEK|28|10|你要死在陌生人手中， 像未受割禮之人的死， 因為我曾說過， 這是主耶和華說的。」
EZEK|28|11|耶和華的話臨到我，說：
EZEK|28|12|「人子啊，要為 推羅 王作哀歌，對他說，主耶和華如此說： 你曾是完美的典範， 智慧充足，全然美麗。
EZEK|28|13|你在 伊甸 ─上帝的園中， 佩戴各樣寶石， 就是紅寶石、紅璧璽、金剛石、 水蒼玉、紅瑪瑙、碧玉、 藍寶石、綠寶石、紅玉； 你的寶石有黃金的底座，手工精巧 ， 都是在你受造之日預備的。
EZEK|28|14|我指定你為受膏的基路伯， 看守保護； 你在上帝的聖山上； 往來在如火的寶石中。
EZEK|28|15|你從受造之日起行為正直， 直到後來查出你的不義。
EZEK|28|16|你因貿易發達， 暴力充斥其中，以致犯罪， 所以我污辱你，使你離開上帝的山。 守護者基路伯啊， 我已將你從如火的寶石中殲滅。
EZEK|28|17|你因美麗心中高傲， 因榮光而敗壞智慧， 我已將你拋棄在地， 把你擺在君王面前， 好叫他們目睹眼見。
EZEK|28|18|你因罪孽眾多，貿易不公， 褻瀆了你的聖所； 因此我使火從你中間發出， 燒滅了你， 使你在所有觀看的人眼前 變為地上的灰燼。
EZEK|28|19|萬民中凡認識你的 都必為你驚奇。 你令人驚恐， 不再存留於世，直到永遠。」
EZEK|28|20|耶和華的話臨到我，說：
EZEK|28|21|「人子啊，你要面向 西頓 ，向它說預言。
EZEK|28|22|你要說，主耶和華如此說： 『 西頓 ，看哪，我與你為敵， 我要在你中間得榮耀。』 我在它中間施行審判、顯為聖的時候， 人就知道我是耶和華。
EZEK|28|23|我必令瘟疫進入 西頓 ， 使血流在街上。 刀劍從四圍臨到它， 被殺的要仆倒在其中； 人就知道我是耶和華。」
EZEK|28|24|「四圍恨惡 以色列 家的人，對他們必不再如刺人的荊棘，傷人的蒺藜；他們就知道我是主耶和華。」
EZEK|28|25|主耶和華如此說：「我將分散在萬民中的 以色列 家召集回來，在列國眼前向他們顯為聖的時候，他們仍可在我所賜給我僕人 雅各 之地居住。
EZEK|28|26|他們要在這地上安然居住。我向四圍恨惡他們的眾人施行審判之後，他們要建造房屋，栽葡萄園，安然居住，他們就知道我是耶和華─他們的上帝。」
EZEK|29|1|第十年十月十二日，耶和華的話臨到我，說：
EZEK|29|2|「人子啊，你要面向 埃及 王法老，向他和 埃及 全地說預言。
EZEK|29|3|你要說，主耶和華如此說： 埃及 王法老， 你這臥在自己江河中的海怪， 看哪，我與你為敵。 你曾說：『我的 尼羅河 是我的， 是我為自己造的。』
EZEK|29|4|我必用鉤子鉤住你的腮頰， 令江河中的魚貼住你的鱗甲； 我要把你和所有貼著鱗甲的魚 從你的江河中拉上來。
EZEK|29|5|我要把你和江河中的魚全都拋棄在曠野； 你必仆倒在田間， 無人收殮，無人掩埋。 我已將你給了地上的走獸、空中的飛鳥作食物。
EZEK|29|6|「 埃及 所有的居民必定知道我是耶和華。因為你已成為 以色列 家蘆葦的杖；
EZEK|29|7|他們用手掌一握，你就斷裂，傷了他們的肩；他們靠著你，你卻折斷，閃了他們的腰 。
EZEK|29|8|所以主耶和華如此說：我必使刀劍臨到你，把人與牲畜從你中間剪除。
EZEK|29|9|埃及 地必荒蕪廢棄，他們就知道我是耶和華。 「因為法老說『 尼羅河 是我的，是我所造的』，
EZEK|29|10|所以，看哪，我必與你和你的江河為敵，使 埃及 地，從 密奪 到 色弗尼 ，直到 古實 邊界，全然廢棄荒蕪。
EZEK|29|11|人的腳不經過，獸的蹄也不經過，四十年之久無人居住。
EZEK|29|12|我要使 埃及 地成為荒蕪中最荒蕪的地，使它的城鎮變為荒廢中最荒廢的城鎮，共四十年之久。我必將 埃及 人分散到列國，四散在列邦。
EZEK|29|13|「主耶和華如此說：滿了四十年後，我必招聚分散在萬民中的 埃及 人。
EZEK|29|14|我要令 埃及 被擄的人歸回，使他們回到本地 巴特羅 。在那裏，他們必成為弱小的國家，
EZEK|29|15|成為列國中最低微的，不再自高於列邦之上。我必使他們變為小國，不再轄制列邦。
EZEK|29|16|埃及 必不再作 以色列 家的倚靠，卻使 以色列 家想起他們仰賴 埃及 的罪。他們就知道我是主耶和華。」
EZEK|29|17|第二十七年正月初一，耶和華的話臨到我，說：
EZEK|29|18|「人子啊， 巴比倫 王 尼布甲尼撒 令他的軍兵大力攻打 推羅 ，以致頭都光禿，肩都磨破；然而他和軍兵雖然為攻打 推羅 花這麼多力氣，卻沒有從那裏得到甚麼犒賞。
EZEK|29|19|所以主耶和華如此說：我要將 埃及 地賜給 巴比倫 王 尼布甲尼撒 ；他必擄掠 埃及 的財富，搶奪它的擄物，擄掠它的掠物，用以犒賞他的軍兵。
EZEK|29|20|我將 埃及 地賜給他，犒賞他，因他們為我效勞。這是主耶和華說的。
EZEK|29|21|「當那日，我必使 以色列 家壯大 ，又必使你─ 以西結 在他們中間開口；他們就知道我是耶和華。」
EZEK|30|1|耶和華的話臨到我，說：
EZEK|30|2|「人子啊，你要說預言；你要說，主耶和華如此說： 哀哉這日！你們應當哭號，
EZEK|30|3|因為日子近了， 耶和華的日子臨近了； 那是密雲之日， 是列國受罰 之期。
EZEK|30|4|必有刀劍臨到 埃及 ； 被殺的人仆倒在 埃及 時， 古實 人顫驚不已。 埃及 的財富遭擄掠， 根基被拆毀。
EZEK|30|5|古實 人、 弗 人、 路德 人、混居的各族和 古伯 人，以及盟國的人都要與 埃及 人一同倒在刀下。」
EZEK|30|6|耶和華如此說： 扶助 埃及 的必傾倒， 埃及 驕傲的權勢必降為卑， 從 密奪 到 色弗尼 ，人必倒在刀下。 這是主耶和華說的。
EZEK|30|7|埃及 成為荒涼中最荒涼的國， 它的城鎮變為荒廢中最荒廢的城鎮。
EZEK|30|8|我在 埃及 放火， 幫助 埃及 的，都遭滅絕； 那時，他們就知道我是耶和華。
EZEK|30|9|「到那日，必有使者從我面前乘船出去，使安逸無慮的 古實 人驚懼；當 埃及 遭難的日子，痛苦也必臨到他們。看哪，這事臨近了！
EZEK|30|10|主耶和華如此說： 我要藉 巴比倫 王 尼布甲尼撒 的手 除滅 埃及 的軍隊。
EZEK|30|11|他和隨從他的人， 就是列國中兇暴的人， 要前來毀滅這地， 拔刀攻擊 埃及 ， 使遍地佈滿被殺的人。
EZEK|30|12|我要使江河乾涸， 將這地賣在惡人手中； 我要藉外國人的手， 使這地和其中所充滿的變為荒蕪； 這是我─耶和華說的。
EZEK|30|13|「主耶和華如此說： 我要毀滅偶像， 從 挪弗 除掉神像； 不再有君王出自 埃及 地， 我要使 埃及 地的人懼怕。
EZEK|30|14|我必令 巴特羅 荒涼， 在 瑣安 放火， 向 挪 施行審判。
EZEK|30|15|我要將我的憤怒傾倒在 訓 ， 埃及 的堡壘上， 要剪除 挪 的眾民。
EZEK|30|16|我必在 埃及 放火， 訓 必大大痛苦， 挪 被攻破， 挪弗 終日遭敵侵襲。
EZEK|30|17|亞文 和 比‧伯實 的年輕人必倒在刀下， 這些城鎮將被擄掠。
EZEK|30|18|我在 答比匿 折斷 埃及 的軛 ， 使它驕傲的權勢止息。 那時，日光必退去； 至於這城，必有密雲遮蔽， 鄰近的城鎮 也遭擄掠。
EZEK|30|19|我要如此向 埃及 施行審判， 他們就知道我是耶和華。」
EZEK|30|20|第十一年正月初七，耶和華的話臨到我，說：
EZEK|30|21|「人子啊，我已折斷 埃及 王法老的一隻膀臂；看哪，無人為他敷藥，也無人為他包紮繃帶，使他有力持刀。
EZEK|30|22|因此，主耶和華如此說：看哪，我與 埃及 王法老為敵，要折斷他的膀臂，折斷強壯的和已受傷的，使刀從他手中掉落。
EZEK|30|23|我必將 埃及 人分散到列國，四散在列邦。
EZEK|30|24|我要使 巴比倫 王的膀臂有力，把我的刀交在他手中；卻要折斷法老的膀臂，使他在 巴比倫 王面前呻吟，如同被殺的人一樣。
EZEK|30|25|我要使 巴比倫 王的膀臂強壯，法老的膀臂卻要下垂；當我把我的刀交在 巴比倫 王手中時，他要舉刀攻擊 埃及 地，他們就知道我是耶和華。
EZEK|30|26|我必將 埃及 人分散到列國，四散在列邦；他們就知道我是耶和華。」
EZEK|31|1|第十一年三月初一，耶和華的話臨到我，說：
EZEK|31|2|「人子啊，你要對 埃及 王法老和他的軍隊說： 論到你的強盛，誰能與你相比呢？
EZEK|31|3|看哪， 亞述 是 黎巴嫩 的香柏樹， 枝條榮美，蔭密如林， 極其高大，樹頂高聳入雲。
EZEK|31|4|眾水使它生長， 深水使它長高； 所栽之地有江河環繞， 汊出的水道流至田野的樹木。
EZEK|31|5|所以它高大超過田野的樹木； 生長時因水源豐沛， 枝子繁多，枝條增長。
EZEK|31|6|空中所有的飛鳥在枝子上搭窩， 野地所有的走獸在枝條下生子， 所有的大國也在它的蔭下居住。
EZEK|31|7|它樹大枝長，極為榮美， 因它的根在眾水之旁。
EZEK|31|8|上帝園中的香柏樹不能遮蔽它； 松樹不及它的枝子， 楓樹不及它的枝條， 上帝園中的樹都沒有它榮美。
EZEK|31|9|我使它枝條繁多， 極為榮美； 在上帝的園中， 伊甸 所有的樹都嫉妒它。」
EZEK|31|10|所以主耶和華如此說：「因它 高大，樹頂高聳入雲，心高氣傲，
EZEK|31|11|我要把它交給 列國中強人的手裏，他們必定按它的罪惡懲治它。我已經驅逐它。
EZEK|31|12|外國人，就是列國中兇暴的人，已把它砍斷拋棄。它的枝條掉落山間和一切谷中，枝子折斷，落在地上一切河道。地上的萬民都離開它的遮蔭，拋棄了它。
EZEK|31|13|空中的飛鳥都棲身在掉落的樹幹上，野地的走獸也都躺臥在它的枝條中。
EZEK|31|14|為了要使水邊的樹木枝幹不再長高，樹頂也不再高聳入雲；那些得水滋潤的，不再屹立於其中。因為它們和下到地府的人一起，都被交與死亡，到了地底下。」
EZEK|31|15|主耶和華如此說：「它墜落陰間的那日，我為它遮蓋深淵，攔住江河，使眾水停流，以表哀悼。我使 黎巴嫩 為它悲哀，田野的樹木都因它枯萎。
EZEK|31|16|我把它扔到陰間，與下到地府的人一同墜落。那時，列國聽見墜落的響聲就震驚； 伊甸 一切的樹木，就是 黎巴嫩 中得水滋潤、最佳最美的樹，在地底下都得了安慰。
EZEK|31|17|這些樹也要與它同下陰間，到被刀所殺的人那裏；它們曾作它的膀臂 ，在列國中曾居住在它的蔭下。
EZEK|31|18|在這樣的榮耀與威勢中， 伊甸 樹木有誰能與你相比呢？然而你要與 伊甸 的樹木一同到地底下；在未受割禮的人中，與被刀所殺的人一同躺下。 「法老和他的軍隊正是如此。這是主耶和華說的。」
EZEK|32|1|第十二年十二月初一，耶和華的話臨到我，說：
EZEK|32|2|「人子啊，你要為 埃及 王法老作哀歌，說： 你在列國中，如同少壯獅子， 卻像海裏的海怪， 衝出江河， 以爪攪動諸水， 使江河渾濁。
EZEK|32|3|主耶和華如此說： 許多民族聚集時， 我要將我的網撒在你身上， 他們要把你拉上來。
EZEK|32|4|我要把你丟在地上， 拋在田野， 使空中的飛鳥落在你身上， 遍地的野獸因你得以飽足。
EZEK|32|5|我要將你的肉丟在山間， 用你巨大的屍首 填滿山谷。
EZEK|32|6|我要以你所流的血 浸透大地， 漫過山頂， 溢滿河道。
EZEK|32|7|我毀滅你時， 要遮蔽諸天， 使眾星昏暗； 我必以密雲遮掩太陽， 月亮也不放光。
EZEK|32|8|我要使天上發亮的光體 在你上面變為昏暗， 使你的地也變為黑暗。 這是主耶和華說的。
EZEK|32|9|「我使你在列國，在你所不認識的列邦中滅亡 。那時，我必使許多民族的心因你愁煩。
EZEK|32|10|當我在他們面前舉起我的刀，我要使許多民族因你驚恐，他們的君王也必因你極其恐慌。在你仆倒的日子，他們各人為自己的性命時時戰兢。
EZEK|32|11|主耶和華如此說： 巴比倫 王的刀必臨到你。
EZEK|32|12|我必藉勇士的刀使你的軍隊仆倒；這些勇士都是列國中兇暴的人。 他們必使 埃及 的驕傲歸於無有， 埃及 的軍隊必被滅絕。
EZEK|32|13|我要除滅眾水旁一切的走獸， 人的腳必不再攪渾這水， 獸的蹄也不攪渾這水。
EZEK|32|14|那時，我必使他們的水澄清， 使他們的江河像油緩流。 這是主耶和華說的。
EZEK|32|15|我使 埃及 地荒廢， 使這地空無一物， 又擊殺其中所有的居民； 那時，他們就知道我是耶和華。
EZEK|32|16|「這是一首為人所吟唱的哀歌；列國的女子要唱這哀歌，她們要為 埃及 和它的軍隊唱這哀歌。這是主耶和華說的。」
EZEK|32|17|第十二年某月 十五日，耶和華的話臨到我，說：
EZEK|32|18|「人子啊，你要為 埃及 的軍隊哀號，把他們和強盛之國 一同扔到地底下，與那些下到地府的人在一起。
EZEK|32|19|『你的美麗勝過誰呢？ 墜落吧，與未受割禮的人躺在一起！』
EZEK|32|20|他們要仆倒在被刀所殺的人當中。 埃及 被交給刀劍，人要把它和它的軍隊拉走。
EZEK|32|21|強壯的勇士要在陰間對 埃及 王和他的盟友說話；他們未受割禮，被刀劍所殺，已經墜落躺下。
EZEK|32|22|「 亞述 和它的全軍在那裏，四圍都是墳墓；他們全都是被殺倒在刀下的人。
EZEK|32|23|他們的墳墓在地府極深之處，它的眾軍環繞它的墳墓，他們全都是被殺倒在刀下的人，曾在活人之地使人驚恐。
EZEK|32|24|「 以攔 在那裏，它的全軍環繞它的墳墓；他們全都是被殺倒在刀下、未受割禮而到地底下的，曾在活人之地使人驚恐；他們與下到地府的人一同擔當羞辱。
EZEK|32|25|人為它和它的軍隊在被殺的人中設立床榻，四圍都是墳墓；他們都是未受割禮被刀所殺的，曾在活人之地使人驚恐；他們與下到地府的人一同擔當羞辱。 以攔 已列在被殺的人中。
EZEK|32|26|「 米設 、 土巴 和他們的全軍都在那裏，四圍都是墳墓；他們都是未受割禮被刀所殺的，曾在活人之地使人驚恐。
EZEK|32|27|他們不得與那未受割禮 仆倒的勇士躺在一起；這些勇士帶著兵器下到陰間，頭枕著刀劍，骨頭帶著本身的罪孽，曾在活人之地使人驚恐。
EZEK|32|28|法老啊，你必與未受割禮的人一起毀滅，與被刀所殺的人躺在一起。
EZEK|32|29|「 以東 在那裏，它的君王和所有官長雖然英勇，還是與被刀所殺的人同列；他們必與未受割禮的和下到地府的人躺在一起。
EZEK|32|30|「在那裏有北方的眾王子和所有的 西頓 人，全都與被殺的人一同下去。他們雖然英勇，使人驚恐，還是蒙羞。他們未受割禮，和被刀所殺的人躺在一起，與下到地府的人一同擔當羞辱。
EZEK|32|31|「法老看見他們，就為他的軍兵，就是被刀所殺屬法老的人和他的全軍感到安慰。這是主耶和華說的。
EZEK|32|32|我任憑法老在活人之地使人驚恐，法老和他的軍兵必躺在未受割禮和被刀所殺的人中。這是主耶和華說的。」
EZEK|33|1|耶和華的話臨到我，說：
EZEK|33|2|「人子啊，你要吩咐本國的百姓，對他們說：我使刀劍臨到哪一國，哪一國的百姓從他們中間選立一人，作為守望者。
EZEK|33|3|守望者見刀劍臨到那地，若吹角警戒百姓，
EZEK|33|4|有人聽見角聲卻不受警戒，刀劍來除滅了他，這人的血必歸到自己頭上。
EZEK|33|5|他聽見角聲，不受警戒，他的血必歸到自己身上；他若受警戒，就救了自己的命。
EZEK|33|6|倘若守望者見刀劍臨到，卻不吹角，以致百姓未受警戒，刀劍來殺了他們中間的一個人，這人雖然因自己的罪孽而死，我卻要從守望者的手裏討他的血債。
EZEK|33|7|「人子啊，我照樣立你作 以色列 家的守望者；你要聽我口中的話，替我警戒他們。
EZEK|33|8|我對惡人說：『惡人哪，你必要死！』你若不開口警戒惡人，使他離開所行的道，這惡人必因自己的罪孽而死，我卻要從你手裏討他的血債。
EZEK|33|9|但是你，你若警戒惡人，叫他離棄所行的道，他仍不轉離，他必因自己的罪孽而死，你卻救了自己的命。」
EZEK|33|10|「人子啊，你要對 以色列 家說：你們曾這樣說：『我們的過犯罪惡在自己身上，我們必因此消滅，怎能存活呢？』
EZEK|33|11|你要對他們說，主耶和華說：我指著我的永生起誓，我斷不喜悅惡人死亡，惟喜悅惡人轉離他所行的道而存活。 以色列 家啊，你們回轉，回轉離開惡道吧！何必死亡呢？
EZEK|33|12|人子啊，你要對本國的百姓說：義人的義，在他犯罪之日不能救他；至於惡人的惡，在他轉離惡行之日不會使他傾倒；義人在他犯罪之日不能因自己的義存活。
EZEK|33|13|我對義人說：『你必存活！』他若倚靠自己的義作惡，所行的義就不被記念；他必因所作的惡死亡。
EZEK|33|14|我對惡人說：『你必死亡！』他若轉離他的罪惡，行公平公義的事；
EZEK|33|15|惡人若歸還抵押品，歸回所搶奪的東西，遵行生命的律例，不再作惡；他必存活，不致死亡。
EZEK|33|16|他所犯的一切罪必不被記念；他行了公平公義的事，必要存活。
EZEK|33|17|「你本國的百姓說：『主的道不公平。』其實他們，他們的道才是不公平。
EZEK|33|18|義人轉離自己的義作惡，他必因此而死亡。
EZEK|33|19|惡人轉離他的惡，行公平公義的事，他必因此而存活。
EZEK|33|20|你們還說：『主的道不公平。』 以色列 家啊，我必按你們各人所行的審判你們。」
EZEK|33|21|我們被擄後第十二年的十月初五，有人從 耶路撒冷 逃到我這裏，說：「城已被攻破。」
EZEK|33|22|逃來的人到的前一天晚上，耶和華的手按在我身上，開我的口。第二天早晨，等那人來到我這裏，我的口就開了，不再說不出話來。
EZEK|33|23|耶和華的話臨到我，說：
EZEK|33|24|「人子啊，住在 以色列 荒廢之地的人說：『 亞伯拉罕 一人能得這地為業，我們人數眾多，這地更是給我們為業的。』
EZEK|33|25|所以你要對他們說，主耶和華如此說：你們吃帶血的食物，向偶像舉目，並且流人的血，你們還能得這地為業嗎？
EZEK|33|26|你們倚靠自己的刀劍行可憎的事，人人污辱鄰舍的妻，你們還能得這地為業嗎？
EZEK|33|27|你要對他們這樣說，主耶和華如此說：我指著我的永生起誓，在廢墟的，必倒在刀下；在田野的，必交給野獸吞吃；在堡壘和洞中的，必遭瘟疫而死。
EZEK|33|28|我必使這地荒廢荒涼，它驕傲的權勢也必止息； 以色列 的山都必荒廢，無人經過。
EZEK|33|29|我因他們所做一切可憎的事，使地荒廢荒涼；那時，他們就知道我是耶和華。」
EZEK|33|30|「你，人子啊，你本國的百姓在城牆旁邊、在房屋門口談論你。弟兄對弟兄彼此說：『來吧！聽聽有甚麼話從耶和華而出。』
EZEK|33|31|他們如同百姓前來，來到你這裏，坐在你面前彷彿是我的子民。他們聽了你的話，卻不實行；因為他們口裏說愛，心卻追隨財利。
EZEK|33|32|看哪，他們看你如同一個唱情歌的人 ，聲音優雅、善於奏樂；他們聽了你的話，卻不實行。
EZEK|33|33|看哪，這話就要應驗；應驗時，他們就知道在他們中間有了先知。」
EZEK|34|1|耶和華的話臨到我，說：
EZEK|34|2|「人子啊，你要向 以色列 的牧人說預言，對他們說，主耶和華如此說：禍哉！ 以色列 的牧人只知牧養自己。牧人豈不當牧養群羊嗎？
EZEK|34|3|你們吃肥油 、穿羊毛、宰殺肥羊，卻不牧養群羊。
EZEK|34|4|瘦弱的，你們不調養；有病的，你們不醫治；受傷的，你們未包紮；被逐的，你們不去領回；失喪的，你們不尋找；卻用暴力嚴嚴地轄制牠們 。
EZEK|34|5|牠們因無牧人就分散；既分散，就成為一切野獸的食物。
EZEK|34|6|我的羊流落眾山之間和各高岡上，分散在全地，無人去尋，無人去找。
EZEK|34|7|「所以，你們這些牧人要聽耶和華的話。
EZEK|34|8|主耶和華說：我指著我的永生起誓，我的羊因無牧人就成為掠物，也作了一切野獸的食物。我的牧人不尋找我的羊；這些牧人只知餵養自己，並不餵養我的羊。
EZEK|34|9|所以你們這些牧人要聽耶和華的話。
EZEK|34|10|主耶和華如此說：看哪，我必與牧人為敵，從他們手裏討回我的羊，使他們不再牧放群羊；牧人也不再餵養自己。我必救我的羊脫離他們的口，不再作他們的食物。」
EZEK|34|11|「主耶和華如此說：『看哪，我必親自尋找我的羊，將牠們尋見。
EZEK|34|12|牧人在羊群四散的日子怎樣尋找他的羊，我必照樣尋找我的羊。這些羊在密雲黑暗的日子散在各處，我要從那裏救回牠們。
EZEK|34|13|我要從萬民中領出牠們，從各國聚集牠們，引領牠們歸回故土。我要在 以色列 山上，在一切溪水旁邊，在境內所有可居住的地牧養牠們。
EZEK|34|14|我要在肥美的草場牧養牠們。牠們的圈必在 以色列 高處的山上，牠們必躺臥在佳美的圈內，在 以色列 山肥美的草場上吃草。
EZEK|34|15|我要親自牧養我的群羊，使牠們得以躺臥。這是主耶和華說的。
EZEK|34|16|失喪的，我必尋找；被逐的，我必領回；受傷的，我必包紮；有病的，我必醫治；只是肥的壯的，我要除滅 ；我必秉公牧養牠們。』
EZEK|34|17|「我的羊群哪，論到你們，主耶和華如此說：看哪，我要在羊與羊中間、公綿羊與公山羊中間施行審判。
EZEK|34|18|你們在肥美的草場上吃草還以為是小事嗎？竟用你們的腳踐踏剩下的草；你們喝了清水，竟用你們的腳攪渾剩下的水。
EZEK|34|19|至於我的羊，只能吃你們所踐踏的，喝你們所攪渾的。
EZEK|34|20|「所以，主耶和華對牠們如此說：看哪，我要親自在肥羊和瘦羊中間施行審判。
EZEK|34|21|因為你們用側邊用肩推擠一切瘦弱的羊，又用角牴撞，使牠們四散在外；
EZEK|34|22|所以，我要拯救我的群羊，牠們必不再作掠物；我也要在羊和羊中間施行審判。
EZEK|34|23|我必在他們之上立一牧人 ，就是我的僕人 大衛 ，牧養牠們；他必牧養他們，作他們的牧人。
EZEK|34|24|我─耶和華必作他們的上帝，我的僕人 大衛 要在他們中間作王。這是我─耶和華說的。
EZEK|34|25|「我要與他們立平安的約，使惡獸從境內斷絕；他們在曠野也能安然居住，在樹林也能躺臥。
EZEK|34|26|我要使他們和我山岡的四圍蒙福；我也必叫時雨落下，使福如甘霖降下。
EZEK|34|27|田野的樹木必結果子，地也必有出產；他們要在自己的土地安然居住。我折斷他們所負的軛，救他們脫離奴役他們之人的手；那時，他們就知道我是耶和華。
EZEK|34|28|他們必不再作外邦人的掠物，地上的野獸也不再吞吃他們；他們卻要安然居住，無人使他們驚嚇。
EZEK|34|29|我必為他們建立聞名的 栽種之地；他們在境內就不再為饑荒所滅，也不再受列國的羞辱。
EZEK|34|30|他們必知道我─耶和華他們的上帝與他們同在，並知道他們， 以色列 家，是我的子民。這是主耶和華說的。
EZEK|34|31|你們這些人，你們是我的羊，我草場上的羊；我是你們的上帝。這是主耶和華說的。」
EZEK|35|1|耶和華的話臨到我，說：
EZEK|35|2|「人子啊，你要面向 西珥山 ，向它說預言，
EZEK|35|3|對它說，主耶和華如此說： 西珥山 ，看哪，我與你為敵，必伸手攻擊你，使你荒涼荒廢。
EZEK|35|4|我必使你的城鎮變為廢墟，使你成為荒涼；你就知道我是耶和華。
EZEK|35|5|因為你永懷仇恨，在 以色列 人遭遇災難、罪孽到了盡頭時，把他們交給刀劍，
EZEK|35|6|所以主耶和華說：我指著我的永生起誓，我必使你遭遇血的報應，血必追趕你；你既不恨惡血，血必追趕你。
EZEK|35|7|我要使 西珥山 荒涼荒廢，把來往經過的人從它那裏剪除。
EZEK|35|8|我要使 西珥山 佈滿被殺的人。被刀殺的要倒在小山和山谷，並一切的溪水中。
EZEK|35|9|我必使你永遠荒涼，使你的城鎮無人居住，你們就知道我是耶和華。
EZEK|35|10|「因為你曾說『這二國、這二邦必歸我，我們必得為業』，其實耶和華仍在那裏；
EZEK|35|11|所以主耶和華說：我指著我的永生起誓，我必照你因仇恨向他們發的怒氣和嫉妒對待你；我審判你的時候，要在他們中間顯明自己。
EZEK|35|12|你必知道我─耶和華已聽見你一切凌辱的話，是針對 以色列 群山說的：『這些山荒涼了，它們是給我們作食物的。』
EZEK|35|13|你們用口向我說誇大的話，增多與我敵對的話，我都聽見了。
EZEK|35|14|主耶和華如此說：全地歡樂的時候，我必使你荒涼。
EZEK|35|15|你怎樣因 以色列 家的地業荒涼而喜樂，我也要照你所做的對待你。 西珥山 哪，你和 以東 全地都必荒涼；人就知道 我是耶和華。」
EZEK|36|1|「人子啊，你要對 以色列 群山說預言： 以色列 群山哪，要聽耶和華的話。
EZEK|36|2|主耶和華如此說，因仇敵說：『啊哈！這古老的丘壇都歸我們為業了！』
EZEK|36|3|所以你要預言，說：主耶和華如此說：因為敵人使你荒涼，四圍踐踏你，要叫你歸其餘的列國為業，使你們成為各族的話柄與百姓的笑談；
EZEK|36|4|因此， 以色列 群山哪，要聽主耶和華的話。對那遭四圍其餘列國佔據、譏刺的大山小岡、水溝山谷、荒廢之地、被棄之城，主耶和華如此說；
EZEK|36|5|所以，主耶和華如此說：我因妒火中燒，就責備其餘的列國和 以東 的眾人。他們快樂滿懷，心存恨惡，將我的地佔為己有，視為被拋棄的掠物。
EZEK|36|6|所以，你要指著 以色列 地說預言，對大山小岡、水溝山谷說，主耶和華如此說：看哪，我在妒忌和憤怒中宣佈：因你們曾受列國的羞辱，
EZEK|36|7|所以我起誓說，你們四圍的列國要擔當自己的羞辱。這是主耶和華說的。
EZEK|36|8|「 以色列 群山哪，要長出枝條，為我子民 以色列 結出果子，因為他們即將來到。
EZEK|36|9|看哪，我是幫助你們的，我要轉向你們，使你們得以耕作栽種。
EZEK|36|10|我要使 以色列 全家在你們那裏人數增多，城鎮有人居住，廢墟重新建造。
EZEK|36|11|我要使人丁和牲畜在你們那裏加增，他們必生養眾多。我要使你們那裏像以前一樣有人居住，並要賜福，比先前更多；你們就知道我是耶和華。
EZEK|36|12|我要使我的子民 以色列 在你們那裏行走，他們必得你為業；你就成為他們的產業，不再使他們喪失兒女。
EZEK|36|13|主耶和華如此說，因為人對你們說『你是吞吃人的，又使國民喪失兒女』，
EZEK|36|14|所以你必不再吞吃人，也不再使國民喪失兒女。這是主耶和華說的。
EZEK|36|15|我使你不再聽見列國的羞辱；你必不再受萬民的辱罵，也不再使國民絆跌。這是主耶和華說的。」
EZEK|36|16|耶和華的話臨到我，說：
EZEK|36|17|「人子啊， 以色列 家住本地的時候，所作所為使那地玷污。他們的行為在我面前，好像婦人在經期中那樣污穢。
EZEK|36|18|所以我因他們在那地流人的血，且以偶像使那地玷污，就把我的憤怒傾倒在他們身上。
EZEK|36|19|我將他們分散到列國，四散在列邦，按他們的所作所為懲罰他們。
EZEK|36|20|他們到了 所去的列國，使我的聖名被褻瀆；因為人談論他們說，這是耶和華的子民，卻從耶和華的地出來。
EZEK|36|21|但我顧惜我的聖名，就是 以色列 家在所到的列國中褻瀆的。
EZEK|36|22|「所以，你要對 以色列 家說，主耶和華如此說： 以色列 家啊，我做這事不是為你們，而是為了我的聖名，就是你們在所到的列國中褻瀆的。
EZEK|36|23|我要使我至大的名顯為聖；這名在列國中已遭褻瀆，是你們在他們中間褻瀆的。我在他們眼前，在你們身上顯為聖的時候，他們就知道我是耶和華。這是主耶和華說的。
EZEK|36|24|我必從列國帶領你們，從列邦聚集你們，領你們回到本地。
EZEK|36|25|我必灑清水在你們身上，你們就潔淨了。我要潔淨你們，使你們脫離一切的污穢，棄絕一切的偶像。
EZEK|36|26|我也要賜給你們一顆新心，將新靈放在你們裏面，又從你們的肉體中除掉石心，賜給你們肉心。
EZEK|36|27|我必將我的靈放在你們裏面，使你們順從我的律例，謹守遵行我的典章。
EZEK|36|28|你們必住在我所賜給你們祖先之地；你們要作我的子民，我要作你們的上帝。
EZEK|36|29|我要救你們脫離一切的污穢，也要令五穀豐登，使你們不再遭遇饑荒。
EZEK|36|30|我要使樹木多結果子，田地多出土產，好叫你們不再因饑荒被列國凌辱。
EZEK|36|31|那時，你們必追念自己的惡行和不好的作為，就因你們的罪孽和可憎的事厭惡自己。
EZEK|36|32|你們要知道，我這樣做不是為你們。 以色列 家啊，你們當為自己的行為抱愧蒙羞。這是主耶和華說的。
EZEK|36|33|「主耶和華如此說：我潔淨你們，使你們脫離一切罪孽的日子，必使城鎮有人居住，廢墟重新建造。
EZEK|36|34|這荒蕪的土地，曾被過路的人看為荒蕪，現今卻得以耕種。
EZEK|36|35|他們必說：『這荒蕪之地，現在成了像 伊甸園 一樣；這荒涼、荒廢、毀壞的城鎮，現今堅固，有人居住。』
EZEK|36|36|那時，在你們四圍其餘的列國必知道，我─耶和華修造那毀壞之處，開墾那荒蕪之地。我─耶和華說了這話，就必成就。
EZEK|36|37|「主耶和華如此說：我要回應 以色列 家的求問，成全他們，增添他們的人數，使他們多如羊群。
EZEK|36|38|在 耶路撒冷 守節時，作為祭物所獻的羊群有多少，照樣，荒涼的城鎮必為人群所充滿；他們就知道我是耶和華。」
EZEK|37|1|耶和華的手按在我身上。耶和華藉著他的靈帶我出去，把我放在平原中，平原遍滿骸骨。
EZEK|37|2|他使我從骸骨的四圍經過，看哪，平原上面的骸骨甚多，看哪，極其枯乾。
EZEK|37|3|他對我說：「人子啊，這些骸骨能活過來嗎？」我說：「主耶和華啊，你是知道的。」
EZEK|37|4|他又對我說：「你要向這些骸骨說預言，對它們說：枯乾的骸骨啊，要聽耶和華的話。
EZEK|37|5|主耶和華對這些骸骨如此說：『看哪，我必使氣息 進入你們裏面，你們就要活過來。
EZEK|37|6|我要給你們加上筋，長出肉，又給你們包上皮，使氣息進入你們裏面，你們就要活過來；你們就知道我是耶和華。』」
EZEK|37|7|於是，我遵命說預言。正說預言的時候，有響聲，看哪，有地震；骨與骨彼此接連。
EZEK|37|8|我觀看，看哪，骸骨上面有筋，長了肉，又包上皮，只是裏面還沒有氣息。
EZEK|37|9|耶和華對我說：「人子啊，你要說預言，向風 說預言。你要說，耶和華如此說：氣息啊，要從四方 而來，吹在這些被殺的人身上，使他們活過來。」
EZEK|37|10|於是我遵命說預言，氣息就進入骸骨，骸骨就活過來，並且用腳站起來，成為極大的軍隊。
EZEK|37|11|他對我說：「人子啊，這些骸骨就是 以色列 全家。他們說：『看哪，我們的骨頭枯乾了，我們的指望失去了，我們滅絕淨盡了！』
EZEK|37|12|所以你要說預言，對他們說，主耶和華如此說：我的子民，看哪，我要打開你們的墳墓，把你們帶出墳墓，領你們進入 以色列 地。
EZEK|37|13|我的子民哪，我打開你們的墳墓，把你們帶出墳墓時，你們就知道我是耶和華。
EZEK|37|14|我必將我的靈放在你們裏面，你們就要活過來。我把你們安置在本地，你們就知道我─耶和華說了這話，就必成就。這是耶和華說的。」
EZEK|37|15|耶和華的話臨到我，說：
EZEK|37|16|「人子啊，你要取一根木杖，在其上寫『為 猶大 和他的盟友 以色列 人』；又取一根 木杖，在其上寫『為 約瑟 ，就是 以法蓮 的杖，和他的盟友 以色列 全家』。
EZEK|37|17|你要將這兩根木杖彼此相接，連成一根，使它們在你手中合而為一。
EZEK|37|18|當你本國的子民對你說：『你這是甚麼意思，你不指示我們嗎？』
EZEK|37|19|你就對他們說，主耶和華如此說：看哪，我要將 約瑟 和他的盟友 以色列 支派的杖，就是在 以法蓮 手中的那根，與 猶大 的杖接連成為一根，在我手中合而為一。
EZEK|37|20|你要在他們眼前，把寫了字的那兩根杖拿在手中，
EZEK|37|21|對他們說，主耶和華如此說：看哪，我要從 以色列 人所到的列國帶領他們，從四圍聚集他們，領他們回到本地。
EZEK|37|22|我要使他們在這地，在 以色列 群山上成為一國，必有一王作他們全體的王。他們不再成為二國，絕不再分為二國。
EZEK|37|23|他們不再因偶像和可憎的物，並一切的罪過玷污自己。我卻要救他們離開一切犯罪所住的地方 ；我要潔淨他們，如此，他們要作我的子民，我要作他們的上帝。』
EZEK|37|24|「我的僕人 大衛 要作他們的王；他們全體必歸一個牧人。他們必順從我的典章，謹守遵行我的律例。
EZEK|37|25|他們要住在我賜給我僕人 雅各 的地上，就是你們列祖所住之地。他們和他們的子孫，並子孫的子孫，都永遠住在那裏。我的僕人 大衛 要作他們的王，直到永遠；
EZEK|37|26|並且我要與他們立平安的約，作為永約。我要安頓他們，使他們人數增多，又在他們中間設立我的聖所，直到永遠。
EZEK|37|27|我的居所必在他們中間；我要作他們的上帝，他們要作我的子民。
EZEK|37|28|我的聖所在 以色列 人中間直到永遠，列國就知道是我─耶和華使 以色列 分別為聖。」
EZEK|38|1|耶和華的話臨到我，說：
EZEK|38|2|「人子啊，你要面向 瑪各 地的 歌革 ，就是 米設 和 土巴 的大王，向他說預言。
EZEK|38|3|你要說，主耶和華如此說： 米設 和 土巴 的大王 歌革 ，看哪，我與你為敵。
EZEK|38|4|我要把你掉轉過來，用鉤子鉤住你的腮頰，把你和你的軍兵、馬匹、騎兵都帶走。他們全都披掛整齊，成為大軍，佩帶大小盾牌，各人拿著刀劍；
EZEK|38|5|他們當中有 波斯 人、 古實 人和 弗 人，都帶著盾牌和頭盔；
EZEK|38|6|還有 歌篾 人和他的軍隊，北方極遠的 陀迦瑪 族和他的軍隊，這許多民族都跟著你。
EZEK|38|7|「你和聚集到你那裏的軍隊都要預備，預備妥當，你要作他們的守衛。
EZEK|38|8|過了多日，你必被差派；到末後之年，你要來到那脫離刀劍、從列國召集回來的人所住之地，來到 以色列 常久荒涼的山上；他們都從列國中被領出，在那裏安然居住。
EZEK|38|9|你和你的全軍，並跟隨你的許多民族都要上來，如暴風刮來，如密雲遮蓋地面。
EZEK|38|10|「主耶和華如此說：那時，你的心必起意念，圖謀惡計，
EZEK|38|11|說：『我要上那無牆的鄉村之地，到那安靜的居民那裏，他們無牆，無門、無閂，安然居住。
EZEK|38|12|我去那裏要搶財為擄物，奪貨為掠物，反手攻擊那從前荒涼、現在有人居住之地，又攻擊那從列國招聚出來、得了牲畜財貨、住在地的高處的百姓。』
EZEK|38|13|示巴 人、 底但 人、 他施 的商人和他們的少壯獅子都對你說：『你來是要搶財為擄物嗎？你聚集軍隊是要奪貨為掠物，奪取金銀，擄去牲畜、財貨，搶奪許多財寶為擄物嗎？』
EZEK|38|14|「人子啊，你要因此說預言，對 歌革 說，主耶和華如此說：我的子民 以色列 安然居住時，你是知道的。
EZEK|38|15|你從你的地方，從北方極遠處率領許多民族前來，他們都騎著馬，是一隊強而多的軍兵。
EZEK|38|16|歌革 啊，你必上來攻擊我的子民 以色列 ，如密雲遮蓋地面。末後的日子，我必領你來攻擊我的地，我藉你在列國眼前顯為聖的時候，他們就要認識我。
EZEK|38|17|主耶和華如此說：我在古時藉我僕人 以色列 眾先知所說的，不就是你嗎？ 他們在那些日子，多年說預言，我必領你來攻擊 以色列 人。」
EZEK|38|18|「主耶和華說： 歌革 上來攻擊 以色列 地的時候，我的怒氣要從鼻孔裏發出。
EZEK|38|19|我在妒忌和如火的烈怒中說：那日在 以色列 地必有大震動，
EZEK|38|20|甚至海中的魚、天空的鳥、野地的獸，和地上爬的各種爬行動物，並地面上的眾人，因見我的面就都震動；山嶺崩裂，陡巖塌陷，一切的牆都必坍塌。
EZEK|38|21|我必令刀劍在我的眾山攻擊 歌革 ；人要用刀劍殺害弟兄。這是主耶和華說的。
EZEK|38|22|我要用瘟疫和血懲罰他。我也必降暴雨、大冰雹、火及硫磺在他和他的軍隊，並跟隨他的許多民族身上。
EZEK|38|23|我必顯為大，顯為聖，在許多國家眼前顯明自己；他們就知道我是耶和華。」
EZEK|39|1|「你，人子啊，要向 歌革 說預言。你要說，主耶和華如此說： 米設 和 土巴 的大王 歌革 ，看哪，我與你為敵。
EZEK|39|2|我要把你調轉過來，帶領你，從北方極遠的地方上來，帶你到 以色列 的群山上。
EZEK|39|3|我要打落你左手的弓，打掉你右手的箭。
EZEK|39|4|你和你的全軍，並跟隨你的列國的人，都必倒在 以色列 的群山上。我要將你給各類攫食的飛鳥和野地的走獸作食物。
EZEK|39|5|你必倒在田野，因為我曾說過，這是主耶和華說的。
EZEK|39|6|我要降火在 瑪各 和海島安然居住的人身上，他們就知道我是耶和華。
EZEK|39|7|「我要在我的子民 以色列 中彰顯我的聖名，不容我的聖名再被褻瀆，列國就知道我─耶和華是 以色列 中的聖者。
EZEK|39|8|看哪，時候到了，必然成就，這就是我曾說過的日子。這是主耶和華說的。
EZEK|39|9|「住 以色列 城鎮的人要出去生火，用軍器燃燒，就是大小盾牌、弓箭、棍棒、槍矛；用它們來燒火，直燒了七年。
EZEK|39|10|他們不必從田野撿柴，也不必從森林伐木，因為他們要用這些軍器燒火。他們要搶奪那搶奪他們的人，擄掠那擄掠他們的人。這是主耶和華說的。」
EZEK|39|11|「當那日，我要把 以色列 境內、海東邊的 旅人谷 給 歌革 在那裏作墳地 ，阻擋了旅行的人 。在那裏，人要埋葬 歌革 和他的軍兵，稱那地為 哈們‧歌革谷 。
EZEK|39|12|以色列 家的人要用七個月埋葬他們，好使那地潔淨。
EZEK|39|13|那地所有的百姓都來埋葬他們。當我得榮耀的日子，這事必叫百姓得名聲。這是主耶和華說的。
EZEK|39|14|他們要分派人專職巡查遍地，埋葬那遺留在地面上入侵者的屍首，好潔淨全地。過了七個月，他們還要再巡查。
EZEK|39|15|巡查的人要遍行全地，見有人的骸骨，就在旁邊立一標記，等埋葬的人來將骸骨葬在 哈們‧歌革谷 ，
EZEK|39|16|且有一城要取名為 哈摩那 。他們必這樣潔淨那地。
EZEK|39|17|「你，人子啊，主耶和華如此說：你要向各類的飛鳥和野地的走獸說：你們要聚集，來吧，從四方聚集來吃我為你們準備的祭物，就是在 以色列 的群山上豐盛的祭物，叫你們吃肉、喝血。
EZEK|39|18|你們要吃勇士的肉，喝地上領袖的血，如吃公綿羊、羔羊、公山羊、公牛；他們全都是 巴珊 的肥畜。
EZEK|39|19|你們吃我為你們準備的祭物，必吃油脂直到飽了，喝血直到醉了。
EZEK|39|20|你們要因我席上的馬匹、騎兵、勇士和所有的戰士而飽足。這是主耶和華說的。」
EZEK|39|21|「我要在列國中彰顯我的榮耀，萬國就必看見我怎樣把手加在他們身上，施行審判。
EZEK|39|22|從那日以後， 以色列 家就知道我是耶和華─他們的上帝，
EZEK|39|23|列國也必知道， 以色列 家被擄掠是因他們的罪孽。他們得罪我，我就轉臉不顧他們，將他們交在敵人手中，使他們全都倒在刀下。
EZEK|39|24|我照他們的污穢和罪過待他們，轉臉不顧他們。
EZEK|39|25|「所以主耶和華如此說：現在，我要使 雅各 被擄的人歸回，要憐憫 以色列 全家，又為我的聖名發熱心。
EZEK|39|26|我將他們從萬民中領回，從仇敵之地召來，在許多國家的眼前，在他們身上顯為聖，他們在本地安然居住，無人使他們驚嚇，那時，他們要擔當 自己的羞辱和干犯我的一切罪。
EZEK|39|27|
EZEK|39|28|我使他們被擄到列國，後又聚集他們回到本地，不再留一人在那裏，那時他們就知道我是耶和華─他們的上帝。
EZEK|39|29|我不再轉臉不顧他們，因我已將我的靈澆灌 以色列 家。這是主耶和華說的。」
EZEK|40|1|我們被擄的第二十五年， 耶路撒冷城 攻破後十四年，正在年初，某月初十，就在那一天，耶和華的手按在我身上，把我帶到那裏。
EZEK|40|2|在上帝的異象中，他帶我到 以色列 地，把我安置在一座極高的山上；在山的南邊有彷彿一座城的建築物。
EZEK|40|3|他帶我到那裏，看哪，有一人面貌 如銅，手拿麻繩和丈量的蘆葦竿，站在門口。
EZEK|40|4|那人對我說：「人子啊，凡我所指示你的，你都要用眼看，用耳聽，並要放在心上。我帶你到這裏來，為要指示你；凡你所見的，都要告訴 以色列 家。」
EZEK|40|5|看哪，殿外四圍有牆。那人手拿丈量的蘆葦竿，長六肘，每肘再加一掌。他量圍牆，寬一竿，高一竿。
EZEK|40|6|他到了朝東的門，就上臺階，量這門的門檻，寬一竿；這門檻寬一竿。
EZEK|40|7|又有守衛房，每間長一竿，寬一竿，守衛房之間相隔五肘。挨著通往殿之門走廊的門檻，一竿。
EZEK|40|8|他量通往殿之門的走廊，一竿。
EZEK|40|9|他量門的走廊，八肘；牆柱，二肘；門的走廊通往殿那裏。
EZEK|40|10|往東的門有守衛房：這旁三間，那旁三間，大小都一樣；這邊和那邊的牆柱，大小也一樣。
EZEK|40|11|他量門的入口，寬十肘，門長十三肘。
EZEK|40|12|守衛房前有矮牆，一肘，那邊的矮牆也是一肘；守衛房這邊六肘，那邊也是六肘。
EZEK|40|13|他量門，從守衛房這邊的房頂到那邊的房頂，寬二十五肘；入口與入口相對。
EZEK|40|14|他量牆柱，六十肘，院子的四周圍有挨著牆柱的門。
EZEK|40|15|從大門入口到裏面門的走廊，五十肘。
EZEK|40|16|守衛房和四圍挨著牆柱的門，都有嵌壁式的窗戶，廊子也有；裏面到處都有窗戶，牆柱上雕刻著棕樹。
EZEK|40|17|他帶我到外院，看哪，院子的四圍有房間，有石板地；石板地上有三十個房間。
EZEK|40|18|沿著門側邊的石板地，就是下面的石板地，與門的長度相同。
EZEK|40|19|他量寬度，從下門的前面到內院外的前面，東向北向一百肘。
EZEK|40|20|他量外院朝北的門的長和寬。
EZEK|40|21|門的守衛房，這旁三間，那旁三間；牆柱和廊子，與第一個門的大小一樣。長五十肘，寬二十五肘。
EZEK|40|22|其窗戶和廊子，並雕刻的棕樹，與朝東的門大小一樣。要登七個臺階才能上到這門，前面 有廊子。
EZEK|40|23|內院有門與這門相對，北面東面都是如此。他從這門量到那門，共一百肘。
EZEK|40|24|他帶我往南去，看哪，朝南有門，他量門的牆柱 和廊子，大小與先前一樣。
EZEK|40|25|門兩旁與廊子的周圍都有窗戶，和先前量的窗戶一樣。門長五十肘，寬二十五肘。
EZEK|40|26|要登七個臺階才能上到這門，前面 有廊子；牆柱上雕刻著棕樹，這邊一棵，那邊一棵。
EZEK|40|27|內院朝南也有門，從這門量到朝南的那門，共一百肘。
EZEK|40|28|他帶我從南門到內院，他量南門，大小與先前一樣。
EZEK|40|29|守衛房和牆柱、廊子，大小與先前一樣。門兩旁與廊子的周圍都有窗戶。門長五十肘，寬二十五肘。
EZEK|40|30|周圍有廊子，長二十五肘，寬五肘。
EZEK|40|31|廊子朝著外院，牆柱上雕刻著棕樹。要登八個臺階才能上到這門。
EZEK|40|32|他帶我到內院的東邊，他量那門，大小與先前一樣。
EZEK|40|33|守衛房和牆柱、廊子，大小與先前一樣。門兩旁與廊子的周圍都有窗戶。長五十肘，寬二十五肘。
EZEK|40|34|廊子朝著外院。牆柱兩邊都雕刻著棕樹。要登八個臺階才能上到這門。
EZEK|40|35|他帶我到北門，他量了，大小與先前一樣，
EZEK|40|36|就是量守衛房和牆柱、廊子。門的周圍都有窗戶；門長五十肘，寬二十五肘。
EZEK|40|37|牆柱 朝著外院。牆柱兩邊都雕刻著棕樹。要登八個臺階才能上到這門。
EZEK|40|38|有房間和它的入口在門的牆柱 旁，那裏是洗燔祭牲的地方。
EZEK|40|39|在門的走廊內，這邊有兩張桌子，那邊也有兩張桌子，其上可宰殺燔祭牲、贖罪祭牲和贖愆祭牲。
EZEK|40|40|上到北門的入口，朝向外面的這邊有兩張桌子，門的走廊那邊也有兩張桌子。
EZEK|40|41|門這邊有四張桌子，那邊也有四張桌子，共八張，在其上宰殺祭牲。
EZEK|40|42|為燔祭牲的四張桌子是用石頭鑿成的，長一肘半，寬一肘半，高一肘。宰殺燔祭牲和其他祭牲所用的器皿可放在其上。
EZEK|40|43|有鉤子，寬一掌，掛在廊內的四周圍。桌子上可放祭牲的肉。
EZEK|40|44|從外面進到內門，內院裏有房間，為歌唱的人而設 ；一間在北門旁，朝南，又有一間在南 門旁，朝北。
EZEK|40|45|他對我說：「這朝南的房間是為了聖殿供職的祭司，
EZEK|40|46|那朝北的房間是為了祭壇前供職的祭司；這些祭司是 利未 人中 撒督 的子孫，近前來事奉耶和華的。」
EZEK|40|47|他又量內院，長一百肘，寬一百肘，是正方的。祭壇就在殿前。
EZEK|40|48|於是他帶我到殿前的走廊，量走廊的牆柱。這面寬五肘，那面寬五肘。 門的兩旁，這邊三肘，那邊三肘。
EZEK|40|49|走廊長二十肘，寬十一肘 。要登臺階 才能上到走廊。靠近牆柱又有柱子，這邊一根，那邊一根。
EZEK|41|1|他帶我到殿那裏，他量牆柱：這面寬六肘，那面寬六肘，寬窄與會幕相同 。
EZEK|41|2|門口寬十肘。門的兩旁，這邊五肘，那邊五肘。他又量了殿，長四十肘，寬二十肘。
EZEK|41|3|他到內殿量門的牆柱，二肘，門口六肘，門的兩旁各寬七肘。
EZEK|41|4|他量內殿，長二十肘，寬二十肘。他對我說：「這是至聖所。」
EZEK|41|5|他又量殿的牆，六肘；圍著殿有廂房，各寬四肘。
EZEK|41|6|廂房有三層，層疊而上，每層排列三十間。殿的牆四周有凸出的牆支撐廂房，廂房就不必以殿的牆為支柱。
EZEK|41|7|這圍繞著殿的廂房越高越寬；廂房圍著殿懸疊而上，所以越上面越寬，從下一層，到中一層，到上一層。
EZEK|41|8|我又見有高臺圍繞著殿，作為廂房的根基，高足足有一竿，就是六大肘。
EZEK|41|9|廂房的外牆寬五肘。殿的廂房和那邊的房間中間還有空地，寬二十肘，圍繞著殿。
EZEK|41|10|
EZEK|41|11|廂房的門口向著空地：一門向北，一門向南。周圍的空地寬五肘。
EZEK|41|12|在西邊空地之後有房子，寬七十肘，長九十肘，牆四圍厚五肘。
EZEK|41|13|這樣，他量了殿，長一百肘，又量空地和那房子並牆，共長一百肘。
EZEK|41|14|殿的前面和東邊的空地，寬一百肘。
EZEK|41|15|他量了空地後面的那房子，並兩旁的樓廊，共長一百肘。 內殿、院的走廊、
EZEK|41|16|門檻 、嵌壁式的窗戶，並對著門檻的三層樓廊，周圍都鑲上木板；地板到窗戶，窗戶都關著，
EZEK|41|17|直到門以上，就是到內殿和外殿內外四圍牆壁，都這樣測量。
EZEK|41|18|牆上雕刻基路伯和棕樹，基路伯和基路伯之間有一棵棕樹，每基路伯有兩張臉；
EZEK|41|19|人的臉向著這邊的棕樹，獅子的臉向著那邊的棕樹，殿內四周圍都是如此。
EZEK|41|20|從地板到門的上面，都有基路伯和棕樹。殿的牆就是這樣。
EZEK|41|21|殿的門柱是方的。至聖所的前面有個東西形狀像
EZEK|41|22|木頭做的壇，高三肘，長二肘 。壇角和底座 ，並四面，都是木頭做的。他對我說：「這是耶和華面前的供桌。」
EZEK|41|23|殿和聖所各有一個雙層門。
EZEK|41|24|每個門有兩扇，每扇又有兩個摺疊頁；這一扇有兩頁，另一扇也有兩頁。
EZEK|41|25|殿的門扇上雕刻著基路伯和棕樹，與刻在牆上的一樣。在外面門的走廊前有木頭做的飛簷。
EZEK|41|26|門的走廊這邊和那邊都有嵌壁式的窗戶和棕樹；殿的廂房和飛簷也是這樣。
EZEK|42|1|他帶我出來往北，到外院，又帶我進入一個房間，一面對著空地，一面對著北邊的房子。
EZEK|42|2|前面長一百肘，寬五十肘，有門向北；
EZEK|42|3|對著內院那二十肘 ，又對著外院的石板地，在第三層樓有樓廊對著樓廊。
EZEK|42|4|那些房間前有一條走道，寬十肘，往裏面有寬一肘的通道 。房門都向北。
EZEK|42|5|房間因為樓廊佔掉一些地方，所以房子的上層比中下兩層窄。
EZEK|42|6|房間分三層，卻不像外院的屋子用柱子支撐，而是從地面往上，所以一層比一層更窄。
EZEK|42|7|外面有一道牆，長五十肘，在房間前面，與朝外院的房間平行。
EZEK|42|8|靠著外院的房間長五十肘，看哪，朝聖殿的長一百肘。
EZEK|42|9|這些房間下面的東邊有一個入口，從外院可由此進入；
EZEK|42|10|其寬如院牆。朝東 也有房間，一面對著空地，一面對著房子。
EZEK|42|11|這些房間前的通道與北邊房間的通道一樣；長、寬、出口、樣式和入口都相同。
EZEK|42|12|在東邊通道的開端，正對著那道牆有門可以進入，與向南邊房間的門一樣。
EZEK|42|13|他對我說：「面對空地南邊的房間和北邊的房間，都是聖的房間；親近耶和華的祭司當在那裏吃至聖的東西，也當在那裏存放至聖的東西，就是素祭、贖罪祭和贖愆祭，因此處為聖。
EZEK|42|14|祭司進聖所，出來的時候，不可直接到外院，要在那裏放下他們供職的衣服，因為這是聖衣；要穿上別的衣服才可以到百姓所在之處。」
EZEK|42|15|他量完了內殿的大小，就帶我出朝東的門，去量院的四周圍。
EZEK|42|16|他用丈量的蘆葦竿量東面，五百竿 ；又轉去
EZEK|42|17|用丈量的蘆葦竿量北面，五百竿；又轉去
EZEK|42|18|用丈量的蘆葦竿量南面，五百竿。
EZEK|42|19|他又轉到西面，用丈量的蘆葦竿去量，五百竿。
EZEK|42|20|他量四面，長五百，寬五百，四周圍有牆，為要分別聖與俗。
EZEK|43|1|以後，他帶我到一座門，就是朝東的門。
EZEK|43|2|看哪， 以色列 上帝的榮光從東而來，他的聲音如同眾水的響聲，地因他的榮耀發光。
EZEK|43|3|我所見的異象如同從前我 來滅城的時候所見的異象，又如我在 迦巴魯河 邊所見的異象，我就臉伏於地。
EZEK|43|4|耶和華的榮光從朝東的門照入殿中。
EZEK|43|5|靈將我舉起，帶入內院，看哪，耶和華的榮光充滿了殿。
EZEK|43|6|我聽見有一位從殿中向我說話，有一人站在我旁邊。
EZEK|43|7|他對我說：「人子啊，這是我寶座之地，是我腳掌所踏之地。我要住在這裏，住在 以色列 人中間直到永遠。 以色列 家和他們的君王不可再以淫行，或在高處以君王的屍首 玷污我的聖名。
EZEK|43|8|因他們使自己的門檻挨近我的門檻，使自己的門框挨近我的門框，又使他們與我之間僅隔一牆，並且行可憎的事，玷污我的聖名，所以我發怒滅絕他們。
EZEK|43|9|現在，他們當從我面前遠離淫行和君王的屍首，我就要住在他們中間，直到永遠。
EZEK|43|10|「你，人子啊，要將這殿指示 以色列 家，讓他們量殿的大小 ，使他們因自己的罪孽羞愧。
EZEK|43|11|他們若因自己所做的一切感到羞愧，你就要將殿的規模、樣式、出口、入口，以及有關整體規模的條例、禮儀、律法指示他們 ，在他們眼前寫下，使他們遵照殿整體的規模和條例去做。
EZEK|43|12|這是殿的律法：山頂上四周圍的全地界都稱為至聖；看哪，這就是殿的律法 。」
EZEK|43|13|這些是祭壇的大小，以肘來量，這肘是一肘一掌。底座高一肘，邊寬一肘，四周圍有邊，高一虎口；這是祭壇的座 。
EZEK|43|14|從底座到下層的臺座，二肘，邊寬一肘。從小臺座到大臺座，四肘，邊寬一肘。
EZEK|43|15|壇上的爐臺，高四肘，從爐臺向上突起四個角。
EZEK|43|16|這爐臺長十二肘，寬十二肘，四面見方。
EZEK|43|17|臺座長十四肘，寬十四肘，四面見方。四周圍有邊，高半肘，底座四圍的邊寬一肘。有臺階朝東。
EZEK|43|18|他對我說：「人子啊，主耶和華如此說：這些是建造祭壇，為要在其上獻燔祭，把血灑在上面的條例：
EZEK|43|19|你要將一頭公牛犢作為贖罪祭，交給那近前來事奉我的 利未 家的祭司 撒督 的後裔；這是主耶和華說的。
EZEK|43|20|你要取那公牛犢的一些血，抹在壇的四角和臺座的四角，並周圍的邊上。你要這樣潔淨壇，為壇贖罪。
EZEK|43|21|你又要將那作贖罪祭的公牛燒在聖所外面，殿的預定之處。
EZEK|43|22|次日，要將無殘疾的公山羊獻為贖罪祭；要潔淨壇，像用公牛潔淨一樣。
EZEK|43|23|你潔淨了壇，就要將一頭無殘疾的公牛犢和羊群中一隻無殘疾的公綿羊
EZEK|43|24|奉到耶和華面前。祭司要撒鹽在其上，獻給耶和華為燔祭。
EZEK|43|25|七日內，你要每日獻一隻公山羊為贖罪祭，也要獻一頭公牛犢和羊群中的一隻公綿羊，都要沒有殘疾的。
EZEK|43|26|七日內祭司要為壇贖罪，使它潔淨，把它分別為聖。
EZEK|43|27|滿了七日，自八日以後，祭司要在壇上獻你們的燔祭和平安祭；我必悅納你們。這是主耶和華說的。」
EZEK|44|1|他又帶我回到聖所朝東的外門，那門關閉了。
EZEK|44|2|耶和華對我說：「這門必須關閉，不可敞開，誰也不可由其中進入；因為耶和華─ 以色列 的上帝已經由其中進入，所以必須關閉。
EZEK|44|3|至於君王，他必按君王的位分坐在其內，在耶和華面前吃餅。他必由這門的走廊而入，也必由此而出。」
EZEK|44|4|他又帶我由北門來到殿前。我觀看，看哪，耶和華的榮光充滿耶和華的殿，我就臉伏於地。
EZEK|44|5|耶和華對我說：「人子啊，我對你所說耶和華殿中一切的條例和律法，你要留心，用眼看，用耳聽，要留心殿的入口和聖所一切的出口。
EZEK|44|6|你要對那悖逆的 以色列 家說，主耶和華如此說： 以色列 家啊，你們行這一切可憎的事，夠了吧！
EZEK|44|7|你們把我的食物，就是脂肪和血獻上的時候，竟把心和肉體未受割禮的外邦人領進我的聖所，玷污我的殿；你們行這一切可憎的事，違背了我的約。
EZEK|44|8|你們未盡看守我聖物的職責，竟派別人在我的聖所替你們盡看守之責。
EZEK|44|9|「主耶和華如此說：所有心和肉體未受割禮的外邦人，就是住在 以色列 中間的任何外邦人，都不可進入我的聖所。」
EZEK|44|10|「 以色列 人走迷的時候， 利未 人遠離我，隨從他們的偶像走迷離開我，他們必擔當自己的罪孽。
EZEK|44|11|他們必在我的聖所當僕役，照管殿門，在殿裏伺候；他們要為百姓宰殺燔祭牲和其他祭牲，站在百姓面前伺候他們。
EZEK|44|12|因為這些 利未 人曾在偶像前伺候他們，成了 以色列 家罪孽的絆腳石，所以我向他們起誓：他們必擔當自己的罪孽。這是主耶和華說的。
EZEK|44|13|他們不可親近我，作事奉我的祭司，也不可挨近我任何一件聖物，就是至聖的物；他們卻要擔當自己的羞辱和所行可憎之事的報應。
EZEK|44|14|我要指派他們在殿裏看守，辦理殿中一切事務，做一切當做的工。」
EZEK|44|15|「 以色列 人走迷離開我的時候， 利未 家的祭司 撒督 的子孫仍然盡看守我聖所的職責；因此他們必親近我，事奉我，並且侍立在我面前，把脂肪與血獻給我。這是主耶和華說的。
EZEK|44|16|只有他們可以進我的聖所，來到我的桌前事奉我，守我吩咐的職責。
EZEK|44|17|他們進內院的門要穿細麻衣，在內院門和殿內供職時不可穿羊毛衣服。
EZEK|44|18|他們要頭戴細麻布的頭巾，腰穿細麻布的褲子；不可穿容易出汗的衣服。
EZEK|44|19|他們出到外院，到外院 百姓那裏，要脫下供職所穿的衣服，放在聖的房間內，換上別的衣服，免得因他們的衣服使百姓成為聖。
EZEK|44|20|他們不可剃頭，也不可留長髮，頭髮一定要修剪。
EZEK|44|21|祭司進內院時不可喝酒。
EZEK|44|22|他們不可娶寡婦或被休的婦人為妻，只可娶 以色列 後裔中的處女，或祭司的寡婦。
EZEK|44|23|他們要教導我的子民分辨聖與俗，使他們知道潔淨和不潔淨的分別。
EZEK|44|24|有爭訟的事，他們應當審判，按我的典章審判。他們要在我的節期守我的律法和條例，也當以我的安息日為聖日。
EZEK|44|25|祭司不可挨近死屍使自己不潔淨，只可為父親、母親、兒子、女兒、兄弟和未出嫁的姊妹使自己不潔淨。
EZEK|44|26|他潔淨之後，他們必須再為他計算七天。
EZEK|44|27|當他進內院，入聖所，在聖所中事奉的日子，要為自己獻上贖罪祭。這是主耶和華說的。
EZEK|44|28|「祭司必有產業，我就是他們的產業。不可在 以色列 中給他們基業，我就是他們的基業。
EZEK|44|29|素祭、贖罪祭和贖愆祭他們都可以吃， 以色列 中一切永獻的祭物都歸他們。
EZEK|44|30|各樣上好的初熟之物和所獻的供物，都要歸祭司。你們也要將最先的麵團給祭司；這樣，福氣就必臨到你們的家。
EZEK|44|31|無論是鳥是獸，凡自然死去的，或是被撕裂的，祭司都不可吃。」
EZEK|45|1|你們抽籤分地為業，要獻上一份作為獻給耶和華的聖地，長二萬五千肘 ，寬二萬 肘。整個地區都作為聖地。
EZEK|45|2|再從其中劃出一塊作為聖所，長五百肘，寬五百肘，四面見方；四圍再加五十肘的空地。
EZEK|45|3|從這整個範圍要劃出長二萬五千肘，寬一萬肘的地，其中要有聖所，是至聖的。
EZEK|45|4|這是地上的一塊聖地，要歸給在聖所供職、親近事奉耶和華的祭司，作為他們房屋用地與聖所的聖地。
EZEK|45|5|其餘長二萬五千肘，寬一萬肘，要歸給在殿中供職的 利未 人，作為他們二十間房屋 的地業。
EZEK|45|6|在那塊獻上的聖地旁邊，你們要劃分造城的地業，寬五千肘，長二萬五千肘，歸 以色列 全家。
EZEK|45|7|劃歸君王的地要在獻上的聖地和城用地的兩旁，面對著聖地，又面對城的用地，西至西邊的疆界，東至東邊的疆界，從西到東，長度與每支派所分得的一樣。
EZEK|45|8|這地要在 以色列 中歸君王為業。我所立的君王必不再欺壓我的子民，卻要按支派把地分給 以色列 家。
EZEK|45|9|主耶和華如此說：「 以色列 的王啊，你們夠了吧！要除掉殘暴和搶奪的事，行公平和公義，不可再勒索我的百姓。這是主耶和華說的。
EZEK|45|10|「你們要用公道的天平、公道的伊法、公道的罷特。
EZEK|45|11|伊法要與罷特等量；一罷特為賀梅珥的十分之一，一伊法也是賀梅珥的十分之一，都以賀梅珥為計算單位。
EZEK|45|12|一舍客勒是二十季拉；二十舍客勒，二十五舍客勒，十五舍客勒，合起來為你們的一彌那。
EZEK|45|13|「你們當獻的供物是這樣：一賀梅珥麥子要獻六分之一伊法，一賀梅珥大麥也要獻六分之一伊法。
EZEK|45|14|獻油的條例是這樣，按油的罷特：每一歌珥油，即十罷特或一賀梅珥，要獻十分之一罷特，原來十罷特等於一賀梅珥。
EZEK|45|15|從 以色列 水源豐沛的草場上，每二百隻羊中要獻一隻羔羊。這都可作素祭、燔祭、平安祭，來為民贖罪。這是主耶和華說的。
EZEK|45|16|這地所有的百姓都要帶這些供物到 以色列 王那裏。
EZEK|45|17|王的本分是在節期、初一、安息日，就是 以色列 家一切的盛會，奉上燔祭、素祭、澆酒祭。他要獻上贖罪祭、素祭、燔祭和平安祭，為 以色列 家贖罪。」
EZEK|45|18|主耶和華如此說：「正月初一，你要取無殘疾的公牛犢，潔淨聖所。
EZEK|45|19|祭司要取一些贖罪祭牲的血，抹在殿的門柱上和祭壇臺座的四角上，並內院的門框上。
EZEK|45|20|本月初七，你也要為誤犯罪的和因無知而犯罪的這樣做；你們要為聖殿贖罪。
EZEK|45|21|「正月十四日，你們要守逾越節，七天的節期都要吃無酵餅。
EZEK|45|22|當日，王要為自己和全國百姓預備一頭公牛作贖罪祭。
EZEK|45|23|節期的七天內，每天他要預備無殘疾的七頭公牛、七隻公綿羊，給耶和華為燔祭；每天又要預備一隻公山羊為贖罪祭。
EZEK|45|24|他也要預備素祭，為一頭公牛同獻一伊法細麵，為一隻公綿羊同獻一伊法細麵，每一伊法加一欣油。
EZEK|45|25|七月十五日守節的時候，七天他都要像這樣預備贖罪祭、燔祭、素祭和油。」
EZEK|46|1|主耶和華如此說：「內院朝東的門，在六個工作的日子必須關閉；惟有安息日和初一要敞開。
EZEK|46|2|王從外面要由門的走廊進入，站在門框旁邊；祭司要為他預備燔祭和平安祭，王要在門的門檻那裏敬拜，然後退出。這門直到晚上不可關閉。
EZEK|46|3|安息日和初一，這地的百姓要在這門口，在耶和華面前敬拜。
EZEK|46|4|安息日，王要用六隻無殘疾的羔羊、一隻無殘疾的公綿羊，獻給耶和華為燔祭；
EZEK|46|5|同獻的素祭，要為公綿羊獻一伊法細麵，為羔羊則按照他的力量獻，一伊法要加一欣油。
EZEK|46|6|初一，他要獻一頭無殘疾的公牛犢、六隻羔羊、一隻公綿羊，全都要用無殘疾的。
EZEK|46|7|他也要預備素祭，為公牛獻一伊法細麵，為公綿羊獻一伊法細麵，為羔羊則按照他的力量獻，一伊法要加一欣油。
EZEK|46|8|王進入的時候要由這門的走廊而入，也要從原路出去。
EZEK|46|9|「在各節期，這地的百姓朝見耶和華的時候，從北門進入敬拜的，要由南門而出；從南門進入的，要由北門而出。不可從進入的門出去，要往前直行，從對面的門出去。
EZEK|46|10|他們進入時，王也跟他們一同進入；他們出去，他也要出去。
EZEK|46|11|「在節期和盛會的日子同獻的素祭，要為一頭公牛獻一伊法細麵，為一隻公綿羊獻一伊法細麵，為羔羊則按照各人的力量獻，一伊法要加一欣油。
EZEK|46|12|王奉獻甘心祭，就是向耶和華甘心獻的燔祭或平安祭時，當有人為他開朝東的門。他就獻上燔祭和平安祭，與安息日所獻的一樣，然後退出。他出去之後，當有人將門關閉。」
EZEK|46|13|「每日，你要取一隻無殘疾一歲的羔羊獻給耶和華為燔祭；要每天早晨獻上。
EZEK|46|14|每天早晨你也要預備同獻的素祭，六分之一伊法細麵，並三分之一欣油，調和細麵。這素祭要經常獻給耶和華，作為永遠的定例。
EZEK|46|15|每天早晨要這樣獻上羔羊、素祭和油，為經常獻的燔祭。」
EZEK|46|16|主耶和華如此說：「王若將禮物賜給他的任何一個兒子，這就成為兒子的產業，可留給子孫，是他們所承受的地業。
EZEK|46|17|倘若王將他產業的一份賜給他的一個臣僕，這就成為他臣僕的產業，直到自由之年，然後地要歸還王；王的產業終究要歸自己的兒子。
EZEK|46|18|王不可奪取百姓的產業，以致趕逐他們離開自己的地業；他應該從自己的地業中將產業賜給子孫，免得我的子民離開自己的地業，四散各處。」
EZEK|46|19|他帶領我從大門旁邊的入口，進到朝北為祭司所預備聖的房間，看哪，西邊盡頭有一塊土地。
EZEK|46|20|他對我說：「這是祭司煮贖愆祭牲、贖罪祭牲，烤素祭的地方，免得帶出外院，使百姓成為聖。」
EZEK|46|21|他又帶我出到外院，使我經過院子的四個角落，看哪，院子的每個角落都有一個小院子。
EZEK|46|22|院子四個角落有小院子，周圍有牆，每個小院子長四十肘 ，寬三十肘；四個角落的小院子大小都一樣，
EZEK|46|23|小院子周圍各有一排石牆，每排石牆下面有爐灶。
EZEK|46|24|他對我說：「這些是煮肉用的屋子，殿內的僕役要在這裏煮百姓的祭物。」
EZEK|47|1|他帶我回到殿門，看哪，有水從殿的門檻下面往東流出，因為這殿是朝東的。水從殿的側面，就是右邊，從祭壇的南邊往下流。
EZEK|47|2|他帶我出北門，又領我從外邊轉到朝東的外門，看哪，水從右邊流出。
EZEK|47|3|他手拿繩子往東出去，量了一千肘，使我涉水而過，水到腳踝。
EZEK|47|4|他又量了一千，使我涉水而過，水就到膝；再量了一千，使我過去，水就到腰；
EZEK|47|5|又量了一千，水已成河，無法過去；因為水勢高漲成河，只能游泳，無法走過。
EZEK|47|6|他對我說：「人子啊，你看見了嗎？」 他帶我回到河邊。
EZEK|47|7|我回到河邊時，看哪，河這邊與那邊的岸上有極多的樹木。
EZEK|47|8|他對我說：「這水往東方流，下到 亞拉巴 ，直到海。所流出來的水，一入海 就使水變淡 。
EZEK|47|9|這兩條河 所到之處，凡滋生的動物都必存活；這水流到那裏，使那裏的水變淡，因此裏面有極多的魚。這河水所到之處，百物都必存活。
EZEK|47|10|必有漁夫站在河邊，從 隱‧基底 直到 隱‧以革蓮 ，全都成了曬 網的場所。那裏的魚各從其類，好像大海的魚甚多。
EZEK|47|11|但是沼澤與池塘的水無法變淡，只能作產鹽之用。
EZEK|47|12|河這邊與那邊的岸上必生長各類樹木，可作食物；葉子不枯乾，果子不斷絕。每月必結新果子，因為這水是從聖所流出來的。樹上的果子必作食物，葉子可以治病。」
EZEK|47|13|主耶和華如此說：「這是你們按 以色列 十二支派分地為業的地界， 約瑟 要得兩份。
EZEK|47|14|你們承受這地為業，要彼此均分；我曾起誓應許將這地賜給你們的列祖，這地必歸你們為業。
EZEK|47|15|「這地的疆界如下：北界從 大海 往 希特倫 ，直到 西達達 口；
EZEK|47|16|又往 哈馬 、 比羅他 、 西伯蓮 ( 西伯蓮 在 大馬士革 的邊界與 哈馬 的邊界中間)，到 浩蘭 邊界的 哈撒‧哈提干 。
EZEK|47|17|這樣，疆界是從 大海 往 大馬士革 地界上的 哈薩‧以難 ，北邊以 哈馬 為界。這是北界。
EZEK|47|18|「東界在 浩蘭 和 大馬士革 中間， 基列 和 以色列 地的中間，以 約旦河 為界。你們要量疆界直到東海 。這是東界。
EZEK|47|19|「南界是從 他瑪 到 加低斯 的 米利巴 水，經 埃及 溪谷 ，直到 大海 。這是南界。
EZEK|47|20|「西界就是 大海 ，從南界直到 哈馬口 對面。這是西界。
EZEK|47|21|「你們要為自己按 以色列 的支派分這地。
EZEK|47|22|要抽籤分這地為業，歸自己和那在你們中間寄居，生兒育女的外人。你們要看他們如本地出生的 以色列 人，他們要在 以色列 支派中與你們同得地業。
EZEK|47|23|外人寄居在哪個支派，你們就在哪裏將地業分給他們。這是主耶和華說的。」
EZEK|48|1|眾支派的名字如下：從北邊盡頭，由 希特倫 往 哈馬 口，到 大馬士革 地界上的 哈薩‧以難 。北邊靠著 哈馬 地，從東到西是 但 的一份。
EZEK|48|2|靠著 但 的地界，從東到西，是 亞設 的一份。
EZEK|48|3|靠著 亞設 的地界，從東到西，是 拿弗他利 的一份。
EZEK|48|4|靠著 拿弗他利 的地界，從東到西，是 瑪拿西 的一份。
EZEK|48|5|靠著 瑪拿西 的地界，從東到西，是 以法蓮 的一份。
EZEK|48|6|靠著 以法蓮 的地界，從東到西，是 呂便 的一份。
EZEK|48|7|靠著 呂便 的地界，從東到西，是 猶大 的一份。
EZEK|48|8|靠著 猶大 的地界，從東到西，必有你們所當獻的聖地，寬二萬五千肘 ；長短與各族從東到西所分的地相同，聖所當在其中。
EZEK|48|9|你們獻給耶和華的聖地要長二萬五千肘，寬一萬肘。
EZEK|48|10|這聖地要歸祭司，北長二萬五千肘，西寬一萬肘，東寬一萬肘，南長二萬五千肘。耶和華的聖所當在其中。
EZEK|48|11|這地要歸 撒督 的子孫中成為聖的祭司，他們謹守我所吩咐的；當 以色列 人走迷的時候，他們不像那些 利未 人走迷了。
EZEK|48|12|在聖地中要特別保留一份歸他們，為至聖，緊鄰著 利未 人的地界。
EZEK|48|13|利未 人所得的地長二萬五千肘，寬一萬肘，與祭司的地界相等，都長二萬五千肘，寬一萬肘。
EZEK|48|14|這地不可賣，不可換；這上好的部分不可轉讓給別人，因為它歸耶和華為聖。
EZEK|48|15|剩下的地長二萬五千肘、寬五千肘，要作公用，為造城、蓋房、空地之用；城要在中間。
EZEK|48|16|以下是城的大小：北面四千五百肘，南面四千五百肘，東面四千五百肘，西面四千五百肘。
EZEK|48|17|城要有空地，向北二百五十肘，向南二百五十肘，向東二百五十肘，向西二百五十肘。
EZEK|48|18|靠著聖地並排剩餘的，東長一萬肘，西長一萬肘；它與聖地並排，其中所出產的要作城內工人的食物。
EZEK|48|19|以色列 支派中所有在城內做工的，都要耕種這地。
EZEK|48|20|你們要將整塊四方的聖地，長二萬五千肘，寬二萬五千肘，連同城的用地都獻作聖地。
EZEK|48|21|聖地和城的用地兩邊剩餘的要歸給王。地的東邊，南北二萬五千肘，東至東界；西邊，南北二萬五千肘，西至西界；靠著各支派所分的地，都要歸給王。聖地和殿的聖所要在其中。
EZEK|48|22|利未 人的地與城的用地都在王的地中間， 猶大 邊界和 便雅憫 邊界之間，要歸給王。
EZEK|48|23|論到其餘的支派，從東到西，是 便雅憫 的一份。
EZEK|48|24|靠著 便雅憫 的地界，從東到西，是 西緬 的一份。
EZEK|48|25|靠著 西緬 的地界，從東到西，是 以薩迦 的一份。
EZEK|48|26|靠著 以薩迦 的地界，從東到西，是 西布倫 的一份。
EZEK|48|27|靠著 西布倫 的地界，從東到西，是 迦得 的一份。
EZEK|48|28|靠著 迦得 南邊的地界，界限從 他瑪 到 加低斯 的 米利巴 水，經 埃及 溪谷 ，直到 大海 。
EZEK|48|29|這就是你們要抽籤分給 以色列 支派為業之地，是他們各支派所得的份。這是主耶和華說的。
EZEK|48|30|以下是城的出口：北面四千五百肘，
EZEK|48|31|城的各門要按 以色列 的支派命名。北面有三個門，一為 呂便 門，一為 猶大 門，一為 利未 門。
EZEK|48|32|東面四千五百肘，有三個門，一為 約瑟 門，一為 便雅憫 門，一為 但 門。
EZEK|48|33|南面四千五百肘，有三個門，一為 西緬 門，一為 以薩迦 門，一為 西布倫 門。
EZEK|48|34|西面四千五百肘，有三個門，一為 迦得 門，一為 亞設 門，一為 拿弗他利 門。
EZEK|48|35|城的周圍共一萬八千肘。從此以後，這城的名字必稱為「耶和華的所在」。
DAN|1|1|猶大 王 約雅敬 在位第三年， 巴比倫 王 尼布甲尼撒 來到 耶路撒冷 ，將城圍困。
DAN|1|2|主將 猶大 王 約雅敬 和上帝殿中的一些器皿交在他的手中。他就把他們帶到 示拿 地他神明的廟裏，將器皿收入他神明的庫房中。
DAN|1|3|王吩咐太監長 亞施毗拿 ，從 以色列 人的王室後裔和貴族中帶進幾個人來，
DAN|1|4|就是沒有殘疾、相貌俊美、通達各樣學問 、知識聰明俱備、足能在王宮侍立的少年，要教他們 迦勒底 的文字和語言。
DAN|1|5|王從自己所用的膳和所飲的酒中，派給他們每日的分量，養育他們三年，好叫他們期滿以後侍立在王面前。
DAN|1|6|他們中間有 猶大 人 但以理 、 哈拿尼雅 、 米沙利 和 亞撒利雅 。
DAN|1|7|太監長給他們另外起名，稱 但以理 為 伯提沙撒 ，稱 哈拿尼雅 為 沙得拉 ，稱 米沙利 為 米煞 ，稱 亞撒利雅 為 亞伯尼歌 。
DAN|1|8|但以理 卻立志，不以王的膳和王所飲的酒玷污自己，於是懇求太監長容他不使自己玷污。
DAN|1|9|上帝使 但以理 在太監長眼前蒙恩，得憐憫。
DAN|1|10|太監長對 但以理 說：「我懼怕我主我王，他已經派給你們飲食，何必讓他見你們的面貌比你們同年齡的少年憔悴呢？這樣，你們就使我的頭在王那裏不保了。」
DAN|1|11|但以理 對太監長所派監管 但以理 、 哈拿尼雅 、 米沙利 、 亞撒利雅 的管理者說：
DAN|1|12|「請你考驗僕人們十天，給我們素菜吃，清水喝，
DAN|1|13|然後你親自觀察我們的面貌和那用王膳的少年的面貌；就照你所觀察的待你的僕人吧！」
DAN|1|14|管理者准許他們這件事，考驗他們十天。
DAN|1|15|過了十天，他們的身材看來比所有享用王膳的少年更加俊美健壯，
DAN|1|16|於是管理者撤去王派給他們用的膳和所飲的酒，只給他們素菜。
DAN|1|17|這四個少年，上帝在各樣文字學問上賜給他們知識和聰明； 但以理 又明白各樣異象和夢兆。
DAN|1|18|王吩咐帶他們進宮的日子到了，太監長就把他們帶到 尼布甲尼撒 面前。
DAN|1|19|王與他們談論，在所有少年中找不到人能與 但以理 、 哈拿尼雅 、 米沙利 、 亞撒利雅 相比，於是他們就在王面前侍立。
DAN|1|20|王考問他們一切智慧和聰明的事，發現他們比全國所有的術士和巫師勝過十倍。
DAN|1|21|到 居魯士 王元年， 但以理 還健在。
DAN|2|1|尼布甲尼撒 在位第二年，他做了很多夢，心裏煩亂，不能睡覺。
DAN|2|2|王吩咐人將術士、巫師、行邪術的和 迦勒底 人召來，要他們把王的夢告訴王；他們就來，站在王面前。
DAN|2|3|王對他們說：「我做了一個夢，心裏煩亂，想要知道這是甚麼夢。」
DAN|2|4|迦勒底 人用 亞蘭 話對王說：「願王萬歲！請將夢告訴僕人，我們就可以講解。」
DAN|2|5|王回答 迦勒底 人說：「這事我已決定，你們若不把夢和夢的解釋告訴我，就必被凌遲，你們的房屋必成糞堆；
DAN|2|6|但你們若能說出這個夢和夢的解釋，就必從我得到禮物、賞賜和殊榮。現在，你們要把夢和夢的解釋告訴我。」
DAN|2|7|他們再一次回答說：「請王將夢告訴僕人，我們就可以講解。」
DAN|2|8|王回答說：「我確實知道你們是故意拖延，因為你們知道這事我已決定。
DAN|2|9|你們若不將夢告訴我，只有一個辦法對待你們；因為你們彼此串通，向我胡言亂語，要等候情勢改變。現在，你們要將夢告訴我，讓我知道你們真能為我解夢。」
DAN|2|10|迦勒底 人回答王說：「世上沒有人能解釋王的事情；從來沒有君王、大臣、掌權者向術士、巫師，或 迦勒底 人問過這樣的事。
DAN|2|11|王所問的事很難，除了不與血肉之軀同住的上帝，沒有人能在王面前解釋。」
DAN|2|12|王因這事生氣，大大震怒，吩咐滅絕 巴比倫 所有的智慧人。
DAN|2|13|命令發出，智慧人將要被殺，人就尋找 但以理 和他的同伴，要殺他們。
DAN|2|14|王的護衛長 亞略 奉命去殺 巴比倫 的智慧人， 但以理 用婉言和智慧回應，
DAN|2|15|向王的大臣 亞略 說：「王的命令為何這樣緊急呢？」 亞略 就把事情告訴 但以理 。
DAN|2|16|於是 但以理 進去求王寬限，好為王解夢。
DAN|2|17|但以理 回到他的居所，把這事告訴他的同伴 哈拿尼雅 、 米沙利 、 亞撒利雅 ，
DAN|2|18|要他們祈求天上的上帝施憐憫，將這奧祕指明，免得 但以理 和他的同伴與 巴比倫 其餘的智慧人一同滅亡。
DAN|2|19|這奧祕就在夜間異象中顯明給 但以理 ， 但以理 就稱頌天上的上帝。
DAN|2|20|但以理 說： 「上帝的名是應當稱頌的，從亙古直到永遠！ 因為智慧和能力都屬乎他。
DAN|2|21|他改變時間、季節， 他廢王，立王； 將智慧賜給智慧人， 將知識賜給聰明人。
DAN|2|22|他顯明深奧隱祕的事， 洞悉幽暗中的一切， 光明也與他同住。
DAN|2|23|我列祖的上帝啊，我感謝你，讚美你， 因你將智慧才能賜給我， 我們所求問的現在你已指明給我， 把王的事給我們指明。」
DAN|2|24|於是， 但以理 進到王所派滅絕 巴比倫 智慧人的 亞略 那裏去，對他這樣說：「不要滅絕 巴比倫 的智慧人，求你領我到王面前，我可以為王解夢。」
DAN|2|25|亞略 就急忙領 但以理 到王面前，對王這樣說：「我在被擄的 猶大 人中找到一人，能將夢的解釋告訴王。」
DAN|2|26|王對那稱為 伯提沙撒 的 但以理 說：「你能將我所做的夢和夢的解釋告訴我嗎？」
DAN|2|27|但以理 回答王說：「王所問的那奧祕，智慧人、巫師、術士、觀兆的都不能告訴王，
DAN|2|28|只有那在天上的上帝能顯明奧祕。他已把日後將要發生的事指示 尼布甲尼撒 王。你在床上做的夢和你腦中的異象是這樣：
DAN|2|29|你，王啊，你在床上所思想的是關乎日後的事，那顯明奧祕的主已把將來要發生的事指示你。
DAN|2|30|至於我，那奧祕顯明給我，並非因我智慧勝過一切活著的人，而是為了讓王知道夢的解釋，知道你心裏的意念。
DAN|2|31|「你，王啊，你正觀看，看哪，有一個很大的像，這像甚高，極其光耀，立在你面前，形狀非常可怕。
DAN|2|32|這像的頭是純金的，胸膛和膀臂是銀的，腹部和腰是銅的，
DAN|2|33|腿是鐵的，腳是半鐵半泥的。
DAN|2|34|你正觀看，見有一塊非人手鑿出來的石頭打在它半鐵半泥的腳上，把腳砸碎；
DAN|2|35|於是鐵、泥、銅、銀、金都一同砸得粉碎，如夏天禾場上的糠秕，被風吹散，無處可尋。打碎這像的石頭成了一座大山，覆蓋全地。
DAN|2|36|「這就是那夢；我們要在王面前講解那夢。
DAN|2|37|你，王啊，你是諸王之王。天上的上帝已將國度、權勢、能力、尊榮都賜給你。
DAN|2|38|世人和走獸，並天空的飛鳥，不論居住何處，他都交在你的手中，令你掌管這一切。你就是那金的頭。
DAN|2|39|在你以後必興起另一國，不及於你；又有第三國如銅，必掌管全地。
DAN|2|40|第四國必堅壯如鐵，就像鐵能打碎砸碎一切；鐵怎樣壓碎一切，那國也必照樣打碎壓碎。
DAN|2|41|你既看見像的腳和腳趾頭，一半是陶匠的泥，一半是鐵，那國將來也必分裂。你既看見鐵和泥攙雜，那國也必有鐵的力量。
DAN|2|42|那腳趾頭既是半鐵半泥，那國也必半強半弱。
DAN|2|43|你既看見鐵和泥攙雜，他們必有混雜的後裔，卻不能彼此相合，正如鐵和泥不能相合。
DAN|2|44|當諸王在位的時候，天上的上帝必另立一個永不敗壞的國度，這國度必不歸給其他百姓，卻要打碎滅絕所有的國度，存立到永遠。
DAN|2|45|你既看見非人手鑿出來的一塊石頭從山而出，打碎鐵、銅、泥、銀、金，那就是至大的上帝把將來要發生的事給王指明。這夢是確實的，這解釋也是準確的。」
DAN|2|46|當時， 尼布甲尼撒 王臉伏於地，向 但以理 下拜，並且吩咐人給他奉上供物和香。
DAN|2|47|王對 但以理 說：「你既能講明這奧祕，你們的上帝誠然是萬神之神、萬王之主，是奧祕的啟示者。」
DAN|2|48|於是王使 但以理 高升，賞賜他極多的禮物，派他管理 巴比倫 全省，又立他為總理，掌管 巴比倫 所有的智慧人。
DAN|2|49|但以理 求王，王就派 沙得拉 、 米煞 、 亞伯尼歌 管理 巴比倫 省的事務，只是 但以理 仍在朝中侍立。
DAN|3|1|尼布甲尼撒 王造了一個金像，高六十肘，寬六肘，立在 巴比倫 省的 杜拉 平原。
DAN|3|2|尼布甲尼撒 王差人將總督、欽差、省長、參謀、財務、法官、地方官和各省的官員都召了來，為 尼布甲尼撒 王所立的像行開光禮。
DAN|3|3|於是總督、欽差、省長、參謀、財務、法官、地方官和各省的官員都聚集，站在 尼布甲尼撒 所立的像前，要為 尼布甲尼撒 王所立的像行開光禮。
DAN|3|4|那時傳令的大聲呼叫說：「各方、各國、各族 的人哪，有命令傳給你們：
DAN|3|5|你們一聽見角、號、琴、瑟、三角琴、鼓和各樣樂器的聲音，就當俯伏，拜 尼布甲尼撒 王所立的金像。
DAN|3|6|凡不俯伏下拜的，必立刻扔在烈火的窯中。」
DAN|3|7|因此百姓一聽見角、號、琴、瑟、三角琴 和各樣樂器的聲音，各方、各國、各族的人就都俯伏，拜 尼布甲尼撒 王所立的金像。
DAN|3|8|在那時，有幾個 迦勒底 人進前來控告 猶大 人。
DAN|3|9|他們對 尼布甲尼撒 王說：「願王萬歲！
DAN|3|10|你，王啊，你曾降旨，凡聽見角、號、琴、瑟、三角琴、鼓和各樣樂器聲音的，都當俯伏拜這金像。
DAN|3|11|凡不俯伏下拜的，必扔在烈火的窯中。
DAN|3|12|現在有幾個 猶大 人，就是王所派管理 巴比倫 省事務的 沙得拉 、 米煞 、 亞伯尼歌 ；王啊，這些人不理你的諭旨，不事奉你的神明，也不拜你所立的金像。」
DAN|3|13|當時， 尼布甲尼撒 大發烈怒，命令把 沙得拉 、 米煞 、 亞伯尼歌 帶過來；他們就把這幾個人帶到王面前。
DAN|3|14|尼布甲尼撒 對他們說：「 沙得拉 、 米煞 、 亞伯尼歌 ，你們不事奉我的神明，不拜我所立的金像，是真的嗎？
DAN|3|15|現在，你們若準備好，一聽見角、號、琴、瑟、三角琴、鼓和各樣樂器的聲音，就俯伏拜我所造的像；若不下拜，必立刻扔在烈火的窯中，有哪一個神明能救你們脫離我的手呢？」
DAN|3|16|沙得拉 、 米煞 、 亞伯尼歌 對王說：「 尼布甲尼撒 啊，這件事我們不必回答你，
DAN|3|17|即便如此，我們所事奉的上帝能將我們從烈火的窯中救出來。王啊，他必救我們脫離你的手；
DAN|3|18|即或不然，王啊，你當知道，我們絕不事奉你的神明，也不拜你所立的金像。」
DAN|3|19|當時， 尼布甲尼撒 怒氣填胸，向 沙得拉 、 米煞 、 亞伯尼歌 變了臉色，命令把窯燒熱，比平常熱七倍；
DAN|3|20|又命令他軍中的幾個壯士，把 沙得拉 、 米煞 、 亞伯尼歌 捆起來，扔在烈火的窯中。
DAN|3|21|這三人穿著內袍、外衣、頭巾和其他的衣服，被捆起來扔在烈火的窯中。
DAN|3|22|因為王的命令緊急，窯又非常熱，那抬 沙得拉 、 米煞 、 亞伯尼歌 的人都被火焰燒死。
DAN|3|23|但是這三個人， 沙得拉 、 米煞 、 亞伯尼歌 被捆綁著，掉進烈火的窯中。
DAN|3|24|那時， 尼布甲尼撒 王驚奇，急忙站起來，對謀士說：「我們捆起來扔在火裏的不是三個人嗎？」他們回答王說：「王啊，是的。」
DAN|3|25|王說：「看哪，我看見有四個人，並沒有捆綁，在火中行走，也沒有受傷；那第四個的相貌好像神明的兒子。」
DAN|3|26|於是 尼布甲尼撒 靠近烈火窯門，說：「至高上帝的僕人 沙得拉 、 米煞 、 亞伯尼歌 ，出來，來吧！」 沙得拉 、 米煞 、 亞伯尼歌 就從火中出來。
DAN|3|27|那些總督、欽差、省長和王的謀士一同聚集來看這三個人，見火不能傷他們的身體，頭髮沒有燒焦，衣裳也沒有變色，都沒有火燒過的氣味。
DAN|3|28|尼布甲尼撒 說：「 沙得拉 、 米煞 、 亞伯尼歌 的上帝是應當稱頌的！他差遣使者救護倚靠他的僕人，他們不遵王的命令，甚至捨身，在他們上帝以外不肯事奉敬拜別神。
DAN|3|29|現在我降旨，無論何方、何國、何族，凡有人毀謗 沙得拉 、 米煞 、 亞伯尼歌 的上帝，他必被凌遲，他的房屋必成糞堆，因為沒有別神能像這樣施行拯救。」
DAN|3|30|那時王在 巴比倫 省使 沙得拉 、 米煞 、 亞伯尼歌 高升。
DAN|4|1|尼布甲尼撒 王對住在全地各方、各國、各族的人說：「願你們大享平安！
DAN|4|2|我樂意宣揚至高上帝向我所行的神蹟奇事。
DAN|4|3|他的神蹟何其大！ 他的奇事何其盛！ 他的國度存到永遠； 他的權柄存到萬代！
DAN|4|4|「我－ 尼布甲尼撒 安居在家中，在宮裏享受榮華。
DAN|4|5|我做了一個夢，使我懼怕。我在床上的意念和腦中的異象，使我驚惶。
DAN|4|6|因此我降旨召 巴比倫 的智慧人全都到我面前，要他們將夢的解釋告訴我。
DAN|4|7|於是那些術士、巫師、 迦勒底 人、觀兆的都進來，我將那夢告訴他們，他們卻不能把夢的解釋告訴我。
DAN|4|8|最後， 但以理 ，就是按照我神明的名字稱為 伯提沙撒 的，來到我面前，他裏頭有神聖神明的靈，我將夢告訴他：
DAN|4|9|『術士的領袖 伯提沙撒 啊，我知道你裏頭有神聖神明的靈，甚麼奧祕都不能為難你。現在你要把我夢中所見的異象和夢的解釋告訴我 。』
DAN|4|10|「我在床上腦中的異象是這樣：我觀看，看哪，大地中間有一棵樹，極其高大。
DAN|4|11|那樹漸長，而且茁壯，高得頂天，從地極都能看見，
DAN|4|12|葉子華美，果子甚多，可作所有動物的食物；野地的走獸臥在蔭下，天空的飛鳥宿在枝上，凡有血肉的都從這樹得食物。
DAN|4|13|「我觀看，我在床上腦中的異象是這樣，看哪，有守望者，就是神聖的一位，從天而降，
DAN|4|14|大聲呼叫說：『砍倒這樹！砍下枝子！拔掉葉子！拋散果子！使走獸逃離樹下，飛鳥躲開樹枝。
DAN|4|15|樹的殘幹卻要留在地裏，在田野的青草中用鐵圈和銅圈套住。任他讓天上的露水滴濕，和地上的走獸一同吃草，
DAN|4|16|使他的心改變，不再是人的心，而給他一個獸心，使他經過七個時期 。
DAN|4|17|這是眾守望者所發的命令，是眾聖者所作的決定，好叫世人知道至高者在人的國中掌權，要將國賜給誰就賜給誰，並且立極卑微的人執掌國權。』
DAN|4|18|「這是我－ 尼布甲尼撒 王所做的夢。 伯提沙撒 啊，你要說明這夢的解釋；我國中所有的智慧人都不能把夢的解釋告訴我，惟獨你能，因你裏頭有神聖神明的靈。」
DAN|4|19|於是稱為 伯提沙撒 的 但以理 驚駭片時，心意驚惶。王說：「 伯提沙撒 啊，不要因夢和夢的解釋驚惶。」 伯提沙撒 回答說：「我主啊，願這夢歸給恨惡你的人，這夢的解釋歸給你的敵人。
DAN|4|20|你所見的樹漸長，而且茁壯，高得頂天，全地都能看見，
DAN|4|21|葉子華美，果子甚多，可作所有動物的食物；野地的走獸住在其下，天空的飛鳥宿在枝上。
DAN|4|22|「王啊，這成長又茁壯的樹就是你。你的威勢成長及於天，你的權柄達到地極。
DAN|4|23|王既看見一位神聖的守望者從天而降，說：『將這樹砍倒毀壞，樹的殘幹卻要留在地裏，在田野的青草中用鐵圈和銅圈套住。任他讓天上的露水滴濕，與野地的走獸一同吃草，直到經過七個時期。』
DAN|4|24|「王啊，夢的解釋就是這樣：臨到我主我王的事是出於至高者的命令。
DAN|4|25|你必被趕出離開世人，與野地的走獸同住，吃草如牛，讓天上的露水滴濕，且要經過七個時期，直等到你知道至高者在人的國中掌權，要將國賜給誰就賜給誰。
DAN|4|26|這使樹的殘幹存留的命令，是要等你知道天在掌權，你的國必定歸你。
DAN|4|27|王啊，求你悅納我的諫言，以施行公義除去罪過，以憐憫窮人除掉罪惡，或者你的平安可以延長。」
DAN|4|28|這些事都臨到 尼布甲尼撒 王。
DAN|4|29|過了十二個月，他在 巴比倫 王宮頂上散步。
DAN|4|30|王說：「這大 巴比倫 豈不是我用大能大力建為首都，要顯示我威嚴的榮耀嗎？」
DAN|4|31|這話還在王口中的時候，有聲音從天降下，說：「 尼布甲尼撒 王啊，有話對你說，你的國離開你了。
DAN|4|32|你必被趕出離開世人，與野地的走獸同住，吃草如牛，且要經過七個時期；等你知道至高者在人的國中掌權，要將國賜給誰就賜給誰。」
DAN|4|33|當時這話就應驗在 尼布甲尼撒 身上，他被趕出離開世人，吃草如牛，身體被天上的露水滴濕，頭髮長得像鷹的羽毛，指甲長得像鳥爪。
DAN|4|34|「時候到了，我－ 尼布甲尼撒 舉目望天，我的知識復歸於我，我就稱頌至高者，讚美尊敬活到永遠的上帝。 他的權柄存到永遠， 他的國度存到萬代。
DAN|4|35|地上所有的居民都算為虛無； 在天上萬軍和地上居民中， 他都憑自己的旨意行事。 無人能攔住他的手， 或問他說，你在做甚麼呢？
DAN|4|36|「那時，我的知識復歸於我，威嚴和光榮也復歸於我，使我的國度得榮耀，我的謀士和大臣也來朝見我。我又重建我的國度，更大的權勢加添在我身上。
DAN|4|37|現在我－ 尼布甲尼撒 讚美、尊崇、恭敬天上的王，因為他所行的全都信實，他所做的盡都公平。那行事驕傲的，他能降為卑。」
DAN|5|1|伯沙撒 王為他的一千大臣擺設盛筵，與這一千人飲酒。
DAN|5|2|伯沙撒 在歡飲之間，吩咐人將他父 尼布甲尼撒 從 耶路撒冷 聖殿所擄掠的金銀器皿拿來，好使王與大臣、王后、妃嬪用這器皿飲酒。
DAN|5|3|於是他們把聖殿，就是 耶路撒冷 上帝殿中所擄掠的金器皿拿來，王和大臣、王后、妃嬪就用這器皿飲酒。
DAN|5|4|他們飲酒，讚美金、銀、銅、鐵、木、石造的神明。
DAN|5|5|當時，忽然有人的指頭出現，在燈臺對面王宮粉刷的牆上寫字。王看見寫字的指頭，
DAN|5|6|就變了臉色，心意驚惶，腰骨好像脫節，雙膝彼此相碰，
DAN|5|7|大聲吩咐將巫師、 迦勒底 人和觀兆的領進來。王對 巴比倫 的智慧人說：「誰能讀這文字，並且向我講解它的意思，他必身穿紫袍，項帶金鏈，在我國中位列第三。」
DAN|5|8|於是王所有的智慧人都進前來，他們卻不能讀那文字，也不能為王講解它的意思。
DAN|5|9|伯沙撒 王就甚驚惶，臉色改變，他的大臣也都困惑。
DAN|5|10|太后 因王和他大臣所說的話，就進入宴會廳，說：「願王萬歲！你的心不要驚惶，臉不要變色。
DAN|5|11|在你國中有一人，他裏頭有神聖神明的靈，你父在世的日子，這人心中光明，又有聰明智慧，好像神明的智慧。你父 尼布甲尼撒 王，就是王的父，曾立他為術士、巫師、 迦勒底 人和觀兆者的領袖，
DAN|5|12|都因他有美好的靈性，又有知識聰明，能解夢，釋謎語，解疑惑。這人名叫 但以理 ， 尼布甲尼撒 王又稱他為 伯提沙撒 ，現在可以召他來，他必解明這意思。」
DAN|5|13|於是 但以理 被領到王面前。王問 但以理 說：「你就是我父王從 猶大 帶來、被擄的 猶大 人 但以理 嗎？
DAN|5|14|我聽說你裏頭有神明的靈，心中有光，又有聰明和高超的智慧。
DAN|5|15|現在智慧人和巫師都被帶到我面前，要叫他們讀這文字，為我講解它的意思；無奈他們都不能講解它的意思。
DAN|5|16|我聽說你能講解，能解疑惑；現在你若能讀這文字，為我講解它的意思，就必身穿紫袍，項戴金鏈，在我國中位列第三。」
DAN|5|17|但以理 回答王說：「你的禮物可以歸你自己，你的賞賜可以歸給別人；我卻要為王讀這文字，講解它的意思。
DAN|5|18|你，王啊，至高的上帝曾將國度、大權、榮耀、威嚴賜給你父 尼布甲尼撒 ；
DAN|5|19|因上帝所賜給他的大權，各方、各國、各族的人都在他面前恐懼戰兢，因他要殺就殺，要人活就活，要升就升，要降就降。
DAN|5|20|但他的心高傲，靈也剛愎，以致行事狂傲，就被革去國度的王位，奪走榮耀。
DAN|5|21|他被趕出離開世人，他的心變為獸心，與野驢同住，吃草如牛，身體被天上的露水滴濕，直到他知道，至高的上帝在人的國中掌權，憑自己的旨意立人治國。
DAN|5|22|伯沙撒 啊，你是他的兒子 ，你雖知道這一切，卻不謙卑自己，
DAN|5|23|竟向天上的主自高，差人將他殿中的器皿拿到你面前，你和大臣、王后、妃嬪用這器皿飲酒。你又讚美那不能看、不能聽、無知無識，用金、銀、銅、鐵、木、石造的神明，沒有將榮耀歸與那手中掌管你氣息，管理你一切行動的上帝。
DAN|5|24|於是從他那裏顯出指頭寫這文字。
DAN|5|25|「所寫的文字是：『彌尼，彌尼，提客勒，烏法珥新 。』
DAN|5|26|解釋是這樣：彌尼就是上帝數算你國的年日到此完畢。
DAN|5|27|提客勒就是你被秤在天平上，秤出你的虧欠來。
DAN|5|28|毗勒斯 就是你的國要分裂，歸給 瑪代 人和 波斯 人。」
DAN|5|29|於是 伯沙撒 下令，人就把紫袍給 但以理 穿上，把金鏈給他戴在頸項上，又傳令使他在國中位列第三。
DAN|5|30|當夜， 迦勒底 王 伯沙撒 被殺。
DAN|5|31|瑪代 人 大流士 年六十二歲，取了 迦勒底 國。
DAN|6|1|大流士 隨心所願，立了一百二十個總督，治理全國，
DAN|6|2|又在他們以上立總長三人， 但以理 也在其中；使總督在他們三人面前呈報，免得王受虧損。
DAN|6|3|這 但以理 因有卓越的靈性，超乎其餘的總長和總督，王想立他治理全國。
DAN|6|4|那時，總長和總督在治國的事務上尋找 但以理 的把柄，為要控告他；只是找不到任何的把柄和過失，因他忠心辦事，毫無錯誤過失。
DAN|6|5|那些人就說：「我們要找 但以理 的把柄，若不從他上帝的律法中下手，就尋不著。」
DAN|6|6|於是，總長和總督紛紛聚集來見王，說：「 大流士 王萬歲！
DAN|6|7|國中的總長、欽差、總督、謀士和省長彼此商議，求王下旨，立一條禁令，三十天之內，不拘何人，若在王以外，或向神明或向人求甚麼，就必扔在獅子坑中。
DAN|6|8|王啊，現在求你立這禁令，在這文件上簽署，使它不能更改；照 瑪代 人和 波斯 人的例，絕不更動。」
DAN|6|9|於是 大流士 王在這禁令的文件上簽署。
DAN|6|10|但以理 知道這文件已經簽署，就進自己的家，他家樓上的窗戶開向 耶路撒冷 。他一天三次，雙膝跪著，在他的上帝面前禱告感謝，像平常一樣。
DAN|6|11|於是，那些人紛紛聚集，發現 但以理 在他上帝面前祈禱懇求。
DAN|6|12|他們就進到王面前，向王提及禁令，說：「三十天之內不拘何人，若在王以外，或向神明或向人求甚麼，必被扔在獅子坑中，王不是在這禁令上簽署了嗎？」王回答說：「確有這事，照 瑪代 人和 波斯 人的例是不可更改的。」
DAN|6|13|他們對王說：「王啊，那被擄的 猶大 人 但以理 不理會你，也不遵守你簽署的禁令，竟一天三次祈禱。」
DAN|6|14|王聽見這話，就甚愁煩，一心要救 但以理 ，直到日落的時候，他還在籌劃解救他。
DAN|6|15|那些人就紛紛聚集到王那裏，對王說：「王啊，當知道 瑪代 人和 波斯 人有例，凡王所立的禁令和律例都不可更改。」
DAN|6|16|於是王下令，人就把 但以理 帶來，扔在獅子坑中。王對 但以理 說：「你經常事奉的上帝，他必拯救你。」
DAN|6|17|有人搬來一塊石頭放在坑口，王用自己的璽和大臣的印，封閉那坑，使懲辦 但以理 的事絕不更改。
DAN|6|18|王回到宮裏，終夜禁食，不讓人帶樂器 到他面前，他也失眠了。
DAN|6|19|次日黎明，王起來，急忙往獅子坑那裏去，
DAN|6|20|臨近坑邊，哀聲呼叫 但以理 。王對 但以理 說：「永生上帝的僕人 但以理 啊，你經常事奉的上帝能救你脫離獅子嗎？」
DAN|6|21|但以理 對王說：「願王萬歲！
DAN|6|22|我的上帝差遣使者封住獅子的口，叫獅子不傷我，因我在上帝面前無辜。王啊，在你面前我也沒有做過任何虧損的事。」
DAN|6|23|王因此就甚喜樂，吩咐把 但以理 從坑裏拉上來。於是 但以理 從坑裏被拉上來，身上毫無損傷，因為他信靠他的上帝。
DAN|6|24|王下令，把那些控告 但以理 的人和他們的妻子兒女都帶來，扔在獅子坑中。他們還沒有到坑底，獅子就制伏他們，咬碎他們的骨頭。
DAN|6|25|於是， 大流士 王傳旨給住在全地各方、各國、各族的人說：「願你們大享平安！
DAN|6|26|現在我降旨，我所統轄全國的人民，都要在 但以理 的上帝面前戰兢畏懼。 因為他是活的上帝， 永遠長存， 他的國度永不敗壞， 他的權柄永存無極！
DAN|6|27|他庇護，搭救， 在天上地下施行神蹟奇事， 救了 但以理 脫離獅子的口。」
DAN|6|28|如此，這 但以理 ，當 大流士 在位的時候和 波斯 的 居魯士 在位的時候，大享亨通。
DAN|7|1|巴比倫 王 伯沙撒 元年， 但以理 在床上做夢，腦中看見異象，就記錄這夢，述說其中的大意。
DAN|7|2|但以理 說： 我在夜間的異象中觀看，看哪，天上有四風，突然颳在大海之上。
DAN|7|3|有四隻巨獸從海裏上來，牠們各不相同：
DAN|7|4|頭一個像獅子，有鷹的翅膀；我正觀看的時候，牠的翅膀被拔去，牠從地上被扶起來，用兩腳站立，像人一樣，還給了牠人的心。
DAN|7|5|看哪，另有一獸如熊，就是第二獸，半身側立，口裏的牙齒中有三根獠牙 。有人吩咐這獸說：「起來，吞吃許多的肉。」
DAN|7|6|其後，我觀看，看哪，另有一獸如豹，背上有四個鳥的翅膀；這獸有四個頭，還給了牠權柄。
DAN|7|7|其後，我在夜間的異象中觀看，看哪，第四獸可怕可懼，極其強壯，有大鐵牙，吞吃嚼碎，剩下的用腳踐踏。這獸與前面所有的獸不同，牠有十隻角。
DAN|7|8|我正思考這些角的時候，看哪，其中又長出另一隻小角；先前的角中有三隻角在它面前連根被拔出。看哪，這角有眼，像人的眼，有口說誇大的話。
DAN|7|9|我正觀看的時候， 有寶座設立， 上面坐著亙古常在者。 他的衣服潔白如雪， 頭髮如純淨的羊毛。 寶座是火焰， 其輪為烈火。
DAN|7|10|有火如河湧出， 從他面前流出來； 事奉他的有千千， 在他面前侍立的有萬萬； 他坐著要行審判 ， 案卷都展開了。
DAN|7|11|於是我觀看，因這角說誇大的話，我正觀看的時候，那獸被殺，身體被毀，扔在火中焚燒。
DAN|7|12|其餘的獸，權柄都被奪去，生命卻得以延續，直到所定的時候和日期。
DAN|7|13|我在夜間的異象中觀看， 看哪，有一位像人子的， 駕著天上的雲而來， 被領到亙古常在者面前。
DAN|7|14|他得了權柄、榮耀、國度， 使各方、各國、各族的人都事奉他。 他的權柄是永遠的，不能廢去， 他的國度必不敗壞。
DAN|7|15|至於我－ 但以理 ，我的靈在我裏面憂傷，我腦中的異象使我驚惶。
DAN|7|16|我走近其中一位侍立者，問他這一切的實情。他就告訴我，使我知道這事的解釋：
DAN|7|17|這四隻巨獸就是將要在世上興起的四個王 。
DAN|7|18|然而，至高者的眾聖者必要得到這國度，並且擁有它，直到永遠，永永遠遠。
DAN|7|19|於是我想要更清楚知道第四獸的實情，牠與一切的獸不同，甚是可怕，有鐵牙銅爪，吞吃嚼碎，剩下的用腳踐踏；
DAN|7|20|頭上有十隻角和那另長出的一角，三隻角在這角面前掉落；這角有眼，有口說誇大的話，形狀比牠的同類更強。
DAN|7|21|我觀看，這角與眾聖者爭戰，勝了他們，
DAN|7|22|直到亙古常在者來到，為至高者的眾聖者伸冤，眾聖者得到國度的時候就到了。
DAN|7|23|那侍立者這樣說： 第四獸就是世上要興起的第四國， 與其他各國不同， 它要併吞全地， 並且踐踏嚼碎。
DAN|7|24|至於那十隻角，就是從這國中興起的十個王； 後來又興起另一王， 與先前的不相同， 他要制伏三個王。
DAN|7|25|他說話抵擋至高者， 折磨至高者的眾聖者， 又改變節期和律法。 眾聖者要交在他手中一年 、兩年、又半年。
DAN|7|26|然而，他坐著要行審判； 他的權柄要被奪去， 毀壞，滅絕，一直到底。
DAN|7|27|國度、權柄和天下諸國的大權 必賜給至高者的眾聖民。 他的國是永遠的國， 所有掌權的都必事奉他，順從他。
DAN|7|28|這事到此結束。我－ 但以理 因這些念頭甚是驚惶，臉色也變了，卻將這事記在心裏。
DAN|8|1|伯沙撒 王在位第三年，有異象向我－ 但以理 顯現，是在先前所見的異象之後。
DAN|8|2|我在異象中觀看，見自己在 以攔 省 書珊 的城堡中；我在異象中又見自己在 烏萊河 邊。
DAN|8|3|我舉目觀看，看哪，有一隻公綿羊站在河邊，牠有兩隻角，這兩角都高，一角高過另一角，後長出來的比較高。
DAN|8|4|我見那公綿羊向西、向北、向南牴撞，沒有任何獸在牠面前站立得住，沒有能逃脫牠手的；牠任意而行，自高自大。
DAN|8|5|我正思想的時候，看哪，有一隻公山羊從西而來，遍行全地，腳不著地。這山羊兩眼當中有一隻顯眼的角。
DAN|8|6|牠往我先前所見、站在河邊、有雙角的公綿羊那裏，以猛烈的怒氣向牠直闖。
DAN|8|7|我見公山羊靠近公綿羊，向牠發怒，攻擊牠，折斷牠的兩角。公綿羊在公山羊面前站立不住；牠把公綿羊撞倒在地，用腳踐踏，沒有能救公綿羊脫離牠手的。
DAN|8|8|這公山羊長得極其高大，正強壯的時候，那大角折斷了，從角的下面向天的四方 長出四隻顯眼的角來。
DAN|8|9|從四角中的一角又長出另一隻小角，向南、向東、向佳美之地，日漸壯大。
DAN|8|10|牠漸壯大，高及諸天萬象，把一些天象和星辰摔落在地，用腳踐踏。
DAN|8|11|牠自高自大 ，自以為高及萬象之君，牠除掉經常獻給君的祭，毀壞君的聖所。
DAN|8|12|因罪過的緣故，有軍隊和經常獻的祭交給牠。牠把真理拋在地上，任意而行 ，無往不利。
DAN|8|13|我聽見有一位聖者說話，又有一位聖者向那說話的聖者說：「這經常獻的祭、帶來荒涼的罪過、聖所與軍隊被踐踏的異象，要持續到幾時呢？」
DAN|8|14|他對我 說：「要到二千三百日，聖所就必潔淨 。」
DAN|8|15|我－ 但以理 見了這異象，想要明白其中的意思。看哪，有一位形狀像人的站在我面前。
DAN|8|16|我聽見 烏萊河 中有人聲呼叫說：「 加百列 啊，要使這人明白這異象。」
DAN|8|17|他就來到我所站的地方。他一來，我就驚慌，臉伏於地。他對我說：「人子啊，你要明白，因為這是關乎末後時期的異象。」
DAN|8|18|他對我說話的時候，我正沉睡，臉伏於地。他就摸我，扶我站起來。
DAN|8|19|他說：「看哪，我要指示你惱怒結束的時候必成的事，因為這是關乎末後指定的時期。
DAN|8|20|你所看見那有雙角的公綿羊就是 瑪代 王和 波斯 王。
DAN|8|21|那公山羊就是 希臘 王；兩眼當中的大角就是第一個王。
DAN|8|22|至於角折斷了，又從角的下面長出四隻角，意思就是有四個國要從這國興起，只是權勢都不及它。
DAN|8|23|這四國末期，惡貫滿盈的時候，必有一王興起，面貌兇惡，詭計多端。
DAN|8|24|他的權柄極大，卻不是因自己的能力；他要施行驚人的毀滅，無往不利，任意而行，又要毀滅強有力的人和眾聖民。
DAN|8|25|他用權術使手中的詭計成功；他的心自高自大，趁人無備的時候毀滅多人。他又起來攻擊萬君之君，至終卻非因人的手而遭毀滅。
DAN|8|26|所說二千三百日 的異象是真的，但你要將這異象封住，因為它關乎未來許多的日子。」
DAN|8|27|於是我－ 但以理 昏倒，病了數日，然後起來辦理王的事務。我因這異象驚駭不已，但還是不能了解。
DAN|9|1|瑪代 族 亞哈隨魯 的兒子 大流士 被立為王，統治 迦勒底 國元年，
DAN|9|2|就是他在位第一年，我－ 但以理 從書上得知，耶和華的話臨到 耶利米 先知，論 耶路撒冷 荒涼期滿的年數為七十年。
DAN|9|3|我面向主上帝，禁食，披麻蒙灰，懇切禱告祈求。
DAN|9|4|我向耶和華－我的上帝祈禱、認罪，說：「主啊，你是大而可畏的上帝，向愛主、守主誡命的人守約施慈愛。
DAN|9|5|我們犯罪作惡，行惡叛逆，偏離你的誡命典章，
DAN|9|6|沒有聽從你僕人眾先知奉你的名向我們君王、官長、祖先和這地所有百姓所說的話。
DAN|9|7|主啊，你是公義的，但我們 猶大 人和 耶路撒冷 的居民，並你所趕到各國的 以色列 眾人，不論遠近，因為背叛了你，臉上蒙羞，正如今日一樣。
DAN|9|8|耶和華啊，我們和我們的君王、官長、祖先因得罪了你，臉上就都蒙羞。
DAN|9|9|主－我們的上帝是憐憫饒恕人的，我們卻違背了他，
DAN|9|10|沒有聽從耶和華－我們上帝的話，沒有遵行他藉僕人眾先知向我們頒佈的律法。
DAN|9|11|以色列 眾人都犯了你的律法，偏離、不聽從你的話；因此，你僕人 摩西 律法上所寫的詛咒和誓言傾倒在我們身上，因我們得罪了上帝。
DAN|9|12|上帝使大災禍臨到我們，實現了警戒我們和審判我們官長的話；原來 耶路撒冷 所遭遇的災禍是普天之下未曾有過的。
DAN|9|13|這一切災禍臨到我們，是照 摩西 律法上所寫的，我們卻沒有求耶和華－我們上帝的恩惠，使我們回轉離開罪孽，明白你的真理。
DAN|9|14|所以耶和華特意使這災禍臨到我們，耶和華－我們的上帝在他所行的事上都是公義的；我們並沒有聽從他的話。
DAN|9|15|主－我們的上帝啊，你曾用大能的手領你的子民出 埃及 地，使自己得了名聲，正如今日一樣，現在，我們犯了罪，作了惡。
DAN|9|16|主啊，求你按你豐盛的公義，使你的怒氣和憤怒轉離你的城 耶路撒冷 ，就是你的聖山。因我們的罪惡和我們祖先的罪孽， 耶路撒冷 和你的子民被四圍的人羞辱。
DAN|9|17|我們的上帝啊，現在求你垂聽你僕人的祈禱懇求，為你自己的緣故使你的臉向荒涼的聖所發光。
DAN|9|18|我的上帝啊，求你側耳而聽，睜眼而看，眷顧我們那荒涼之地和稱為你名下的城。我們在你面前懇求，不是因自己的義，而是因你豐富的憐憫。
DAN|9|19|主啊，求你垂聽！主啊，求你赦免！主啊，求你側耳，求你實行！為你自己的緣故不要遲延。我的上帝啊，因這城和這民都是稱為你名下的。」
DAN|9|20|我正說話、禱告，承認我的罪和我百姓 以色列 的罪，為我上帝的聖山，在耶和華－我的上帝面前懇求；
DAN|9|21|我正在禱告中說話，先前在異象中所見的那位 加百列 ，約在獻晚祭的時候迅速飛到我這裏來。
DAN|9|22|他指教我說 ：「 但以理 啊，現在我來要使你有智慧，有聰明。
DAN|9|23|你剛開始懇求的時候，就有命令發出。現在我來告訴你，因你是蒙愛的；所以你要思想這事，明白這異象。
DAN|9|24|「為你百姓和你聖城，已經定了七十個七，要止住罪過，除淨罪惡，贖盡罪孽，引進永恆的公義，封住異象和預言，並膏至聖所 。
DAN|9|25|你當知道，當明白，從發出命令恢復並重建 耶路撒冷 ，直到受膏的君出現，必有七個七和六十二個七。 耶路撒冷城 連街帶濠都必在艱難中恢復並重建。
DAN|9|26|過了六十二個七，那受膏者 被剪除，一無所有；必有一王的百姓來毀滅這城和聖所，它的結局 必如洪水沖沒。必有戰爭，一直到末了，荒涼的事已經定了。
DAN|9|27|在一七之期，他必與許多人堅立盟約；一七之半，他必使獻祭與供獻止息。那施行毀滅的可憎之物必立在聖殿裏 ，直到所定的結局傾倒在那行毀滅者的身上。」
DAN|10|1|波斯 王 居魯士 第三年，有話指示那稱為 伯提沙撒 的 但以理 。這話是確實的，指著大戰爭； 但以理 明白這話，明白這異象。
DAN|10|2|那時，我－ 但以理 悲傷了三個七日；
DAN|10|3|美味我沒有吃，酒和肉沒有入我的口，也沒有用油抹我的身，直到滿了三個七日。
DAN|10|4|正月二十四日，我在 大河 ，就是 底格里斯河 邊，
DAN|10|5|舉目觀看，看哪，有一人身穿細麻衣，腰束 烏法 的純金腰帶。
DAN|10|6|他的身體如水蒼玉，面貌如閃電，眼目如火把，手臂和腳如明亮的銅，說話的聲音像眾人的聲音。
DAN|10|7|我－ 但以理 一人看見這異象，跟我一起的人沒有看見，卻有極大的戰兢落在他們身上，他們就逃跑躲避，
DAN|10|8|只剩下我一人。我看見這大異象就渾身無力，面容變色，毫無氣力。
DAN|10|9|我聽見他說話的聲音；一聽見他說話的聲音，我就沉睡，臉伏於地。
DAN|10|10|看哪，有一隻手摸我，使我膝蓋和手掌戰抖。
DAN|10|11|他對我說：「蒙愛的 但以理 啊，要思想我對你所說的話，只管站起來，因為我現在奉差遣來到你這裏。」他對我說這話，我就戰戰兢兢地站起來。
DAN|10|12|他說：「 但以理 啊，不要懼怕！因為自從第一日你立志要明白，又在你上帝面前刻苦自己，你的話已蒙應允；我就是因你的話而來。
DAN|10|13|但 波斯 國的領袖攔阻了我二十一天。看哪，天使長 中的一位 米迦勒 來幫助我，因為我被留在 波斯 諸王那裏。
DAN|10|14|現在我來，要使你明白你百姓日後必遭遇的事，因為這異象關乎未來的日子。」
DAN|10|15|他向我這樣說，我就臉面朝地，啞口無聲。
DAN|10|16|看哪，有一位形狀像人的，摸我的嘴唇，我就開口說話，向那站在我面前的說：「我主啊，因這異象使我感到劇痛，毫無氣力。
DAN|10|17|我主的僕人怎能跟我主說話呢？我現在渾身無力，毫無氣息。」
DAN|10|18|有一位形狀像人的再一次摸我，使我有力量。
DAN|10|19|他說：「蒙愛的人哪，不要懼怕，願你平安！你要剛強！要剛強！ 」他一對我說話，我就覺得有力量，說：「我主請說，因你使我有力量。」
DAN|10|20|他說：「你知道我為甚麼到你這裏來嗎？現在我要回去與 波斯 的領袖爭戰，我去了之後，看哪， 希臘 的領袖必來。
DAN|10|21|但我要將那記錄在真理之書上的話告訴你。除了你們的天使 米迦勒 之外，沒有人幫助我抵擋他們。」
DAN|11|1|「至於我，當 瑪代 的 大流士 元年，我曾起來扶助 米迦勒 ，使他堅強。
DAN|11|2|現在我要指示你確實的事。」 「看哪， 波斯 還有三個王要興起，第四王必富足遠勝諸王。他因富足成為強盛，就煽動各國攻擊 希臘 國。
DAN|11|3|必有一個勇敢的王興起，執掌大權，隨意而行。
DAN|11|4|他正興起的時候，他的國必瓦解，向天的四方 裂開，卻不歸他的後裔，也不如他當年統治的權威；他的國必被拔出，歸給他後裔之外的人。
DAN|11|5|「南方的王必強盛，他的將帥中必有一個比他更強，執掌權柄，權柄甚大。
DAN|11|6|過了幾年，他們必結盟，南方王的女兒必來到北方王那裏，使約生效；但這女子不能保留實力，王的力量 也未能存留。這女子、帶她來的、生她的 和當時扶助她的必被殺害 。
DAN|11|7|但從這女子的本家必另有一子 接續王位，他要率領軍隊進入北方王的堡壘，攻擊他們，而且得勝，
DAN|11|8|把他們的神像和鑄成的偶像，與金銀寶器都擄掠到 埃及 去。數年之內，他不去攻擊北方的王。
DAN|11|9|北方的王必侵入南方王的國土，但卻要撤回本地。
DAN|11|10|「北方王的兒子們必動干戈，招聚許多軍兵。他要前進，如洪水氾濫；要再度爭戰，直搗南方王的堡壘。
DAN|11|11|南方王必發烈怒，出來與北方王爭戰，擺列大軍；北方王的軍兵必敗在南方王的手下。
DAN|11|12|這大軍既被掃蕩，南方王的心就自高；他雖使萬人仆倒，卻不能保持勝利。
DAN|11|13|「北方王要再度擺列大軍，比先前更多。過了幾年，他必率領大軍，帶極多的裝備而來。
DAN|11|14|那時，必有許多人起來攻擊南方王，並且你百姓中的殘暴人要興起，應驗異象，他們卻要敗亡。
DAN|11|15|北方王必來建土堆攻取堅固城，南方的軍兵抵擋不住，就是精選的部隊也無力抵擋；
DAN|11|16|前來攻擊南方王的必任意而行，無人在北方王面前站立得住。他要站在那佳美之地，用手施行毀滅。
DAN|11|17|「他必定意傾全國之力而來，與南方王訂約，把自己的女兒 給南方王為妻，企圖敗壞他的國度。這計謀卻未得逞，自己也得不到好處。
DAN|11|18|其後北方王必轉頭，奪取許多海島。但有一將帥除掉北方王對人的羞辱，並且使羞辱歸到他自己身上。
DAN|11|19|他必轉頭回到本地的堡壘，卻要絆跌仆倒，歸於無有。
DAN|11|20|「那時，有一人興起接續他的王位，他為了王國的榮華，差官員橫征暴斂。這王過不多時就死了，不是因怒氣 ，也不是因戰役。」
DAN|11|21|「後來，有一個卑鄙的人興起接續他的王位，人未曾將國的尊榮給他，他卻趁人無備的時候前來，用詭詐奪取政權。
DAN|11|22|勢如洪水般的軍兵在他面前被沖沒，遭擊潰；立約的領袖也是如此。
DAN|11|23|他與人結盟之後，卻行詭詐。跟隨他的人雖不多，他卻日漸強盛。
DAN|11|24|他趁人無備的時候，來到國中極肥沃之地，做他祖宗和祖宗的祖宗未曾做過的事，瓜分擄物、掠物和財寶，又策劃進攻堡壘；然而這都是暫時的。
DAN|11|25|「他必奮勇向前，率領大軍攻擊南方王；南方王以極強的大軍迎戰，卻抵擋不住，因為有人設計謀害南方王。
DAN|11|26|吃王餉的使王敗壞，王的軍隊必被沖沒，仆倒被殺的甚多。
DAN|11|27|至於這二王，他們心懷惡計，同席吃飯卻彼此說謊，但計謀不成，因為結局要在指定的時期來到。
DAN|11|28|北方王必帶許多財寶回本地，但他的心反對聖約；他恣意橫行，回到本地。
DAN|11|29|「到了指定的時期，他必返回，侵入南方。這一次卻不像前一次，
DAN|11|30|因為 基提 的戰船要來攻擊他，他就喪膽而退。他惱恨聖約，恣意橫行，要回來善待那些背棄聖約的人。
DAN|11|31|他要興兵，這兵必褻瀆聖所，就是堡壘，除掉經常獻的祭，設立那施行毀滅的可憎之物。
DAN|11|32|他必用巧言奉承違背聖約的惡人；惟獨認識上帝的子民必剛強行事。
DAN|11|33|民間的智慧人必訓誨許多人，然而在一段日子裏，他們必因刀劍、火燒、擄掠、搶奪而仆倒。
DAN|11|34|他們仆倒的時候，會得到少許援助，卻有許多人用詭詐加入他們。
DAN|11|35|智慧人中有些人仆倒，為要使他們受熬煉，成為潔淨、潔白，直到末了；因為還有一段日子才到所定的時期。
DAN|11|36|「王必任意而行，自高自大，超過所有的神明，又用荒謬的話攻擊萬神之神。他必行事亨通，直到主的憤怒結束，因為所定的事必然實現。
DAN|11|37|他不顧他祖宗的神明，也不顧婦女所仰慕的神明，任何神明他都不顧；因為他自大，高過一切，
DAN|11|38|以敬奉堡壘的神明取而代之，用金、銀、寶石和珍寶敬奉他祖宗所不認識的神明。
DAN|11|39|他靠外邦神明的幫助，攻破最堅固的堡壘。凡承認他的，他要給他們許多尊榮，使他們管轄許多人，又分封土地作為報償。
DAN|11|40|「到末了，南方王要與北方王交戰。北方王要用戰車、騎兵和許多戰船，勢如暴風來攻擊他，又要侵入列國，如洪水氾濫。
DAN|11|41|他要侵入那佳美之地，許多國就被傾覆 ，但 以東 人、 摩押 人和大半的 亞捫 人必逃離他的手。
DAN|11|42|他要伸手攻擊列國，連 埃及 地也不得逃脫。
DAN|11|43|他要掌管 埃及 的金銀財寶和各樣珍寶， 路比 人和 古實 人都跟從他的腳步。
DAN|11|44|但從東方和北方必有消息傳來擾亂他，他就大發烈怒出去，要將許多人殺滅淨盡。
DAN|11|45|他要在海和榮美的聖山之間搭起王宮的帳幕；然而他的結局到了，無人能幫助他。」
DAN|12|1|「那時，保佑你百姓的天使長 米迦勒 必站起來，並且有大艱難，自從有國以來直到此時，未曾有過這樣的事。那時，你的百姓凡記錄在冊上的，必得拯救。
DAN|12|2|睡在地裏塵埃中的必有多人醒過來；其中有得永生的，有受羞辱永遠被憎惡的。
DAN|12|3|智慧人要發光，如同天上的光；那領許多人歸於義的必發光如星，直到永永遠遠。
DAN|12|4|但以理 啊，你要隱藏這話，封閉這書，直到末時。必有許多人往來奔跑 ，知識 就必增長。」
DAN|12|5|我－ 但以理 觀看，看哪，另有兩個人站立：一個在河這邊，一個在河那邊。
DAN|12|6|其中一個對那在河水之上、穿細麻衣的說：「這奇異的事要到幾時才應驗呢？」
DAN|12|7|我聽見那在河水之上、穿細麻衣的，向天舉起左右手，指著那活到永遠的起誓說：「要到一年 、兩年，又半年，粉碎聖民力量結束的時候，這一切的事就要應驗。」
DAN|12|8|我聽了卻不明白，就說：「我主啊，這些事的結局是怎樣呢？」
DAN|12|9|他說：「 但以理 ，去吧！因為這話已經隱藏封閉，直到末時。
DAN|12|10|必有許多人使自己潔淨、潔白，且受熬煉；但惡人仍必行惡，沒有一個惡人明白，惟獨智慧人能明白。
DAN|12|11|從除掉經常獻的祭，設立那施行毀滅的可憎之物的時候起，必有一千二百九十日。
DAN|12|12|那等候，直到一千三百三十五日的有福了。
DAN|12|13|「至於你，你要去等候結局。你必安息，到了末期，你必起來，享受你的福分。」
HOS|1|1|當 烏西雅 、 約坦 、 亞哈斯 、 希西家 作 猶大 王， 約阿施 的兒子 耶羅波安 作 以色列 王的時候，耶和華的話臨到 備利 的兒子 何西阿 。
HOS|1|2|耶和華初次向 何西阿 說話。耶和華對他說：「你去娶一個淫蕩的女子為妻，收那從淫亂所生的兒女；因為這地行大淫亂，離棄耶和華。」
HOS|1|3|於是， 何西阿 去娶了 滴拉音 的女兒 歌篾 。她就懷孕，為 何西阿 生了一個兒子。
HOS|1|4|耶和華對 何西阿 說：「給他起名叫 耶斯列 ；因為再過片時，我要懲罰 耶戶 家在 耶斯列 流人血的罪，也必終結 以色列 家的王朝。
HOS|1|5|到那日，我必在 耶斯列 平原折斷 以色列 的弓。」
HOS|1|6|歌篾 又懷孕，生了一個女兒，耶和華對 何西阿 說：「給她起名叫 羅‧路哈瑪 ；因為我必不再憐憫 以色列 家，絕不赦免他們。
HOS|1|7|我卻要憐憫 猶大 家，使他們靠耶和華－他們的上帝得救；我必不讓他們靠弓、刀、戰爭、馬匹與騎兵得救。」
HOS|1|8|歌篾 在 羅‧路哈瑪 斷奶以後，又懷孕生了一個兒子。
HOS|1|9|耶和華說：「給他起名叫 羅‧阿米 ；因為你們不是我的子民，我也不是你們的上帝 。」
HOS|1|10|然而， 以色列 的人數必多如海沙，不可量，不可數。從前在甚麼地方對他們說「你們不是我的子民」，將來就在那裏稱他們為「永生上帝的兒子」。
HOS|1|11|猶大 人和 以色列 人要一同聚集，為自己設立一個「頭」，從這地上來，因為 耶斯列 的日子必為大日。
HOS|2|1|你們要稱你們的眾弟兄 為 阿米 ，稱你們的眾姊妹 為 路哈瑪 。
HOS|2|2|要跟你們的母親理論，理論， ─因為她不是我的妻子， 我也不是她的丈夫─ 叫她除掉臉上的淫相 和胸間的淫態，
HOS|2|3|免得我剝光她，使她赤身， 如剛出生的時候一樣， 使她如曠野，如乾旱之地， 乾渴而死。
HOS|2|4|我必不憐憫她的兒女， 因為他們是從淫亂生的兒女。
HOS|2|5|他們的母親行了淫亂， 懷他們的做了可羞恥的事； 因為她說：「我要跟隨我所愛的， 我的餅、水、羊毛、麻、油、酒， 都是他們給的。」
HOS|2|6|因此，看哪，我要用荊棘堵塞她 的道， 築牆擋住她， 使她找不著路；
HOS|2|7|以致她追隨所愛的人，卻追不上， 尋找他們，卻尋不著， 就說：「我要回到前夫那裏去， 因我那時比現在還好。」
HOS|2|8|她不知道是我給她五穀、新酒和新的油， 又加添她的金銀； 他們卻用來供奉 巴力 。
HOS|2|9|因此，我要在收割的日子收回我的五穀， 在當令的季節收回我的新酒， 我要奪回她用以遮體的羊毛和麻。
HOS|2|10|如今我必在她所愛的人眼前顯露她的羞恥 ， 無人能救她脫離我的手。
HOS|2|11|我必使她的宴樂、節期、初一、安息日， 她一切的盛會都止息。
HOS|2|12|我要毀壞她的葡萄樹和無花果樹， 就是她所說「我所愛的給我為賞賜」的； 我要使它們變為荒林， 為野地的走獸所吞吃。
HOS|2|13|我要懲罰她素日給諸 巴力 燒香的罪； 那時她佩戴耳環和珠寶， 跟隨她所愛的，卻忘記我。 這是耶和華說的。
HOS|2|14|因此，看哪，我要誘導她，領她到曠野， 我要說動她的心。
HOS|2|15|在那裏，我必賜她葡萄園， 又賜她 亞割谷 作為指望的門。 她必在那裏回應， 像在年輕時從 埃及 地上來的時候一樣。
HOS|2|16|那日你必稱呼我 伊施 ，不再稱呼我 巴力 。這是耶和華說的。
HOS|2|17|因為我必從她口中除掉諸 巴力 的名號，不再有人提這名號。
HOS|2|18|當那日，我必為我的百姓，與野地的走獸、天空的飛鳥和地上爬行的動物立約；又要在國中折斷弓和刀，止息戰爭，使他們安然躺臥。
HOS|2|19|我必聘你永遠歸我為妻，以公義、公平、慈愛、憐憫聘你歸我；
HOS|2|20|又以信實聘你歸我，你就必認識耶和華。
HOS|2|21|耶和華說：那日我必應允， 我必應允天，天必應允地，
HOS|2|22|地必應允五穀、新酒和新的油； 這些都必應允在 耶斯列 身上。
HOS|2|23|我為自己必將她種在這地。 我必憐憫 羅‧路哈瑪 ； 對 羅‧阿米 說： 「你是我的子民」； 他必說：「我的上帝。」
HOS|3|1|耶和華又對我說：「你去愛那情人所愛卻犯姦淫的婦人，正如耶和華愛那偏向別神、喜愛葡萄餅 的 以色列 人。」
HOS|3|2|於是我用十五舍客勒銀子和一賀梅珥半大麥買她歸我。
HOS|3|3|我對她說：「你當多日與我同住，不可行淫，不可歸與別人，我對你也一樣。」
HOS|3|4|因為 以色列 人必多日過著無君王，無領袖，無祭祀，無柱像，無以弗得，無家中神像的生活。
HOS|3|5|後來 以色列 人必歸回 ，尋求耶和華─他們的上帝和他們的王 大衛 。在末後的日子，他們必敬畏耶和華，領受他的恩惠。
HOS|4|1|以色列 人哪，當聽耶和華的話。 耶和華指控這地的居民， 因為在這地上無誠信， 無慈愛，無人認識上帝；
HOS|4|2|惟起誓、欺騙、殺害、 偷盜、姦淫、殘暴、 流血又流血。
HOS|4|3|因此，這地悲哀， 其上的居民、野地的走獸、 天空的飛鳥都日趨衰微， 海中的魚也必消滅。
HOS|4|4|然而，人都不必爭辯，也不必指責。 你的百姓與抗拒祭司的人一樣。
HOS|4|5|日間你必跌倒， 夜間先知也要與你一同跌倒； 我要滅絕你的母親。
HOS|4|6|我的百姓因無知識而滅亡。 你拋棄知識， 我也必拋棄你， 使你不再作我的祭司。 你既忘了你上帝的律法， 我也必忘記你的兒女。
HOS|4|7|祭司越發增多，就越發得罪我； 我必使他們的榮耀變為羞辱。
HOS|4|8|他們吞吃我百姓的贖罪祭 ， 滿心願意我的子民犯罪。
HOS|4|9|將來百姓所受的， 祭司也必承受； 我必因他們所行的懲罰他們， 照他們所做的報應他們。
HOS|4|10|他們吃，卻不得飽足； 行淫，卻不繁衍； 因為他們離棄耶和華， 常行
HOS|4|11|淫亂。 酒和新酒奪去人的心。
HOS|4|12|我的百姓求問木頭， 以為木杖能指示他們； 淫亂的心使他們失迷， 以致行淫離棄他們的上帝，
HOS|4|13|在各山頂獻祭，在各高岡上燒香， 在橡樹、楊樹、大樹之下， 因為那裏樹影美好。 所以，你們的女兒行淫， 你們的媳婦 犯姦淫。
HOS|4|14|我不因你們的女兒行淫 或你們的媳婦犯姦淫懲罰她們； 因為人自己轉去與娼妓同居， 與神廟娼妓一同獻祭。 這無知的百姓必致傾倒。
HOS|4|15|以色列 啊，你雖然行淫， 猶大 卻不可犯罪； 不要往 吉甲 去， 不要上到 伯‧亞文 ， 也不要指著永生的耶和華起誓。
HOS|4|16|以色列 倔強， 猶如倔強的母牛； 現在耶和華能牧放他們， 如在寬闊之地牧放羔羊嗎？
HOS|4|17|以法蓮 親近偶像， 任憑他吧！
HOS|4|18|他們喝完了酒， 荒淫無度， 他們的官長甚愛羞恥的事。
HOS|4|19|風把他們捲在翅膀裏， 他們必因所獻的祭 蒙羞。
HOS|5|1|眾祭司啊，要聽這話！ 以色列 家啊，要留心聽！ 王室啊，要側耳而聽！ 審判將臨到你們， 因你們在 米斯巴 如羅網， 在 他泊山 如張開的網。
HOS|5|2|這些悖逆的人大行殺戮， 我要斥責他們眾人。
HOS|5|3|至於我，我認識 以法蓮 ， 以色列 不能向我隱藏。 以法蓮 哪，現在你竟然行淫 ， 以色列 竟然被污辱。
HOS|5|4|他們所做的使他們不能歸向上帝， 因有淫亂的心在他們裏面； 他們不認識耶和華。
HOS|5|5|以色列 的驕傲使自己臉面無光 ； 以色列 和 以法蓮 必因自己的罪孽跌倒， 猶大 也必與他們一同跌倒。
HOS|5|6|他們牽著牛羊去尋求耶和華， 卻尋不著； 因他已轉去離開他們。
HOS|5|7|他們不忠於耶和華， 生了私生子。 現在新月必吞滅他們和他們的地業。
HOS|5|8|你們當在 基比亞 吹角， 在 拉瑪 吹號， 在 伯‧亞文 發出警報； 便雅憫 哪，留意你的背後！
HOS|5|9|到了懲罰的日子， 以法蓮 必變為廢墟； 我在 以色列 眾支派中，已指示將來必成的事。
HOS|5|10|猶大 的領袖如同挪移地界的人， 我必把我的憤怒如水傾倒在他們身上。
HOS|5|11|以法蓮 因喜愛遵從荒謬的命令 就受欺壓，在審判中被壓碎。
HOS|5|12|我對 以法蓮 竟如蛀蟲， 向 猶大 家竟如朽爛。
HOS|5|13|以法蓮 見自己有病， 猶大 見自己有傷， 以法蓮 就前往 亞述 ， 差遣人去見大王 ； 他卻不能醫治你們， 不能治好你們的傷。
HOS|5|14|我必向 以法蓮 如獅子， 向 猶大 家如少壯獅子。 我要撕裂，並且離去， 我必奪去，無人搭救。
HOS|5|15|我要去，我要回到原處， 等他們自覺有罪，尋求我的面； 急難時他們必切切尋求我。
HOS|6|1|來，我們歸向耶和華吧！ 他撕裂我們，也必醫治； 打傷我們，也必包紮。
HOS|6|2|過兩天他必使我們甦醒， 第三天他必使我們興起， 我們就在他面前得以存活。
HOS|6|3|我們要認識，要追求認識耶和華。 他如黎明必然出現， 他必臨到我們像甘霖， 像滋潤土地的春雨。
HOS|6|4|以法蓮 哪，我可以向你怎樣行呢？ 猶大 啊，我可以向你怎樣做呢？ 因為你們的慈愛如同早晨的雲霧， 又如速散的露水。
HOS|6|5|因此，我藉先知砍伐他們， 以我口中的話殺戮他們； 對你的審判 如光發出。
HOS|6|6|我喜愛慈愛 ，不喜愛祭物； 喜愛人認識上帝，勝於燔祭。
HOS|6|7|他們卻如 亞當 背約， 在那裏向我行詭詐。
HOS|6|8|基列 是作惡之人的城， 被血沾染。
HOS|6|9|成群的祭司如強盜埋伏等候， 在 示劍 的路上殺戮， 行了邪惡。
HOS|6|10|在 以色列 家我看見可憎的事， 在 以法蓮 那裏有淫行， 以色列 被污辱了。
HOS|6|11|猶大 啊，我使被擄之民歸回的時候， 必有為你所預備的豐收。
HOS|7|1|我正要醫治 以色列 的時候， 以法蓮 的罪孽 和 撒瑪利亞 的邪惡就顯露出來。 他們行事虛謊， 內有賊人入侵， 外有群盜劫掠。
HOS|7|2|他們以為我不在意他們一切的惡行； 現在，他們所做的在我面前纏繞他們。
HOS|7|3|他們行惡使君王歡喜， 說謊使官長快樂。
HOS|7|4|他們全都犯姦淫， 如同烤熱的火爐， 師傅在揉麵到發麵時 暫時停止煽火。
HOS|7|5|在我們君王宴樂的日子， 官長因酒的烈性而生病 ， 王與褻慢的人握手。
HOS|7|6|他們臨近，心裏如火爐一般， 他們等待，如烤餅的整夜睡覺， 到了早晨卻如火焰熊熊。
HOS|7|7|他們全都熱如火爐， 吞滅他們的審判官。 他們的君王都仆倒， 他們中間無一人求告我。
HOS|7|8|以法蓮 混居在萬民中 ， 以法蓮 是沒有翻過的餅。
HOS|7|9|外邦人消耗他的力量，他卻不知道； 頭髮斑白，他也不覺得。
HOS|7|10|以色列 的驕傲使自己臉面無光。 他們雖遭遇這一切， 仍不歸向耶和華－他們的上帝， 也不尋求他。
HOS|7|11|以法蓮 好像鴿子愚蠢無知， 他們求告 埃及 ，投奔 亞述 。
HOS|7|12|他們去的時候，我要把我的網撒在他們身上； 我要捕獲他們如同空中的鳥。 我必按他們會眾所聽到的 懲罰他們。
HOS|7|13|他們因離棄我，必定有禍； 因違背我，必遭毀滅。 我雖想要救贖他們，他們卻向我說謊。
HOS|7|14|他們在床上呼號， 卻不誠心哀求我； 他們為求五穀新酒而聚集 ， 卻背叛我。
HOS|7|15|我雖管教他們，堅固他們的膀臂， 他們卻圖謀邪惡抗拒我。
HOS|7|16|他們歸向，但不是歸向至上者 ； 終究必如鬆弛的弓。 他們的領袖必因舌頭的狂傲倒在刀下， 這在 埃及 地必成為人的笑柄。
HOS|8|1|你用口吹角吧！ 敵人如鷹攻打耶和華的家； 因為他們違背了我的約， 干犯了我的律法。
HOS|8|2|他們必呼求我： 「我的上帝啊，我們 以色列 認識你了 。」
HOS|8|3|以色列 丟棄良善 ； 仇敵必追逼他。
HOS|8|4|他們立君王，並非出於我； 立官長，我卻不知道。 他們用金銀為自己製造偶像， 以致被剪除。
HOS|8|5|撒瑪利亞 啊，耶和華已拋棄你的牛犢； 我的怒氣向拜牛犢的人發作。 他們要到幾時方能無罪呢？
HOS|8|6|因這牛犢是出於 以色列 ， 是匠人所造的， 並不是上帝。 撒瑪利亞 的牛犢必被打碎。
HOS|8|7|他們所栽種的是風， 所收割的是暴風； 禾稼不長穗， 無以製成麵粉； 即便製成， 外邦人也必吞吃它。
HOS|8|8|以色列 被吞吃， 如今在列國中像人所不喜愛的器皿。
HOS|8|9|他們投奔 亞述 如獨行的野驢。 以法蓮 雇用情人，
HOS|8|10|他們雇用列國； 如今我要聚集他們， 他們必因君王和官長所加的重擔開始衰微 。
HOS|8|11|以法蓮 為贖罪增添許多祭壇， 這些祭壇卻使他犯罪。
HOS|8|12|我為他寫了許多條 律法， 他卻以為與他毫無關係。
HOS|8|13|他們獻祭物作為給我的供物， 卻自食其肉， 耶和華並不悅納他們。 現在他必記起他們的罪孽， 懲罰他們的罪惡； 他們必返回 埃及 。
HOS|8|14|以色列 忘記造他的主，建造宮殿， 猶大 增添許多堅固的城； 我卻要降火在他的城鎮， 吞滅其堡壘。
HOS|9|1|以色列 啊，不要歡喜， 像 萬民一樣快樂； 因為你行淫離棄你的上帝， 喜愛各禾場上賣淫所得的賞金。
HOS|9|2|禾場和壓酒池都不足以餵養他們， 它的新酒也必缺乏。
HOS|9|3|他們必不得住耶和華的地； 以法蓮 卻要返回 埃及 ， 在 亞述 吃不潔淨的食物。
HOS|9|4|他們必不得向耶和華獻澆酒祭， 所獻的祭也不蒙悅納。 他們的祭物如居喪者的食物， 凡吃的必使自己玷污； 因為他們的食物只為自己的口腹， 必不得入耶和華的殿。
HOS|9|5|到盛會的日子，在耶和華的節期， 你們要怎樣行呢？
HOS|9|6|看哪，他們要逃避災難； 埃及 人要收殮他們， 摩弗 人要埋葬他們。 蒺藜盤踞他們貴重的銀器， 荊棘必佔據他們的帳棚。
HOS|9|7|降罰的日子近了， 報應的時候已經來到。 以色列 必知道， 先知愚昧， 受靈感動的人狂妄， 皆因你多多作惡，大懷怨恨。
HOS|9|8|以法蓮 替我的上帝守望； 至於先知，他所到之處都有捕鳥人的羅網， 在他上帝的家中也遭人懷恨。
HOS|9|9|他們深深敗壞， 如在 基比亞 的日子一樣。 耶和華必記起他們的罪孽， 懲罰他們的罪惡。
HOS|9|10|我發現 以色列 ， 如在曠野的葡萄； 我看見你們的祖先， 如春季無花果樹上初熟的果子。 他們卻來到 巴力‧毗珥 ， 獻上自己做羞恥的事， 成為可憎惡的， 與他們所愛的一樣。
HOS|9|11|以法蓮 ，他們的榮耀如鳥飛去， 必不生產，不懷胎，不成孕；
HOS|9|12|他們縱然將兒女養大， 我卻要使他們喪子，一個也不留。 我離棄他們， 他們就有禍了。
HOS|9|13|我看 以法蓮 如 推羅 栽於美地。 以法蓮 卻要將自己的兒女帶出來， 交給行殺戮的人。
HOS|9|14|耶和華啊，求你加給他們， 加給他們甚麼呢？ 要使他們懷孕流產， 乳房枯乾。
HOS|9|15|因他們在 吉甲 的一切惡事， 我在那裏憎惡他們。 因他們所行的惡， 我必把他們趕出我的殿， 不再愛他們； 他們的領袖都是悖逆的。
HOS|9|16|以法蓮 受擊打， 其根枯乾，不能結果， 即或生產， 我也要殺他們所生的愛子。
HOS|9|17|我的上帝必棄絕他們， 因為他們不聽從他； 他們必飄流在列國中。
HOS|10|1|以色列 是茂盛的葡萄樹， 結果繁多。 果子越多， 就越增添祭壇； 土地越肥美， 就越建造美麗的柱像。
HOS|10|2|他們心懷二意， 現今要定為有罪。 耶和華必拆毀他們的祭壇， 粉碎他們的柱像。
HOS|10|3|現在他們要說： 「我們沒有王； 因為我們不敬畏耶和華， 王又能為我們做甚麼呢？」
HOS|10|4|他們講空話， 以假誓立約； 因此，懲罰如苦菜滋生 在田間的犁溝中。
HOS|10|5|撒瑪利亞 的居民必因 伯‧亞文 的牛犢驚恐； 它的百姓為它悲哀， 它的祭司為它戰兢， 因為榮耀已經離開它。
HOS|10|6|人必將牛犢帶到 亞述 ， 當作禮物獻給大王。 以法蓮 必蒙羞， 以色列 必因自己的計謀慚愧。
HOS|10|7|撒瑪利亞 的王要滅亡， 如水面上的泡沫一般。
HOS|10|8|亞文 的丘壇， 以色列 犯罪的地方必毀壞， 荊棘和蒺藜必長在他們的祭壇上。 他們要向大山說：遮蓋我們！ 向小山說：倒在我們身上！
HOS|10|9|以色列 啊， 你從 基比亞 的日子以來就時常犯罪， 他們仍停留在那裏。 攻擊罪孽之輩的戰事豈不會臨到 基比亞 嗎？
HOS|10|10|我必隨己意懲罰他們， 他們為雙重的罪所纏； 萬民必聚集攻擊他們。
HOS|10|11|以法蓮 是馴良的母牛犢，喜愛踹穀， 我要將軛套在牠肥美的頸項上， 我要使 以法蓮 被套住； 猶大 必耕田， 雅各 必耙地。
HOS|10|12|你們要為自己栽種公義， 收割慈愛。 你們要開墾荒地， 現今正是尋求耶和華的時候； 等他臨到，公義必如雨降給你們。
HOS|10|13|你們耕種奸惡， 收割罪孽， 吃的是謊言的果實。 因你倚靠自己的行為， 仰賴你眾多的勇士，
HOS|10|14|所以在你百姓中必掀起鬧鬨， 你一切的堡壘必被拆毀， 就如 沙勒幔 在爭戰的日子拆毀 伯‧亞比勒 ， 將城中的母子一同摔死。
HOS|10|15|伯特利 啊，因你們的大惡， 你們必遭遇如此。 黎明來臨， 以色列 的王必全然滅絕。
HOS|11|1|以色列 年幼的時候，我愛他， 就從 埃及 召我的兒子出來。
HOS|11|2|先知 越是呼喚他們， 他們越是遠離 ， 向諸 巴力 獻祭， 為雕刻的偶像燒香。
HOS|11|3|我曾教導 以法蓮 行走， 我用膀臂 抱起他們， 他們卻不知道是我醫治他們。
HOS|11|4|我用慈繩愛索牽引他們； 我待他們如人鬆開牛兩腮旁邊的軛， 彎下身來餵養他們。
HOS|11|5|他們必不返回 埃及 地； 然而 亞述 人要作他們的王， 因他們不肯歸向我。
HOS|11|6|刀劍必臨到他們的城鎮， 毀壞門閂，吞滅眾人， 都因他們自己的計謀。
HOS|11|7|我的百姓偏要背離我， 他們雖向至高者呼求， 他卻不抬舉他們 。
HOS|11|8|以法蓮 哪，我怎能捨棄你？ 以色列 啊，我怎能棄絕你？ 我怎能使你如 押瑪 ？ 怎能使你如 洗扁 ？ 我回心轉意， 我的憐憫燃了起來。
HOS|11|9|我必不發猛烈的怒氣， 也不再毀滅 以法蓮 。 因我是上帝，並非世人， 是你們中間的聖者； 我必不在怒中臨到你們。
HOS|11|10|耶和華如獅子吼叫， 他的兒女必跟隨他。 他一吼叫， 他們就從西方戰兢而來。
HOS|11|11|他們必如雀鳥從 埃及 戰兢而來， 又如鴿子從 亞述 地來到。 我必使他們住自己的房屋； 這是耶和華說的。
HOS|11|12|以法蓮 用謊言圍繞我， 以色列 家用詭計環繞我； 猶大 卻仍與上帝同行 ， 向聖者忠心。
HOS|12|1|以法蓮 以風為食物， 終日追逐東風， 增添虛謊和殘暴， 與 亞述 立約， 也把油送到 埃及 。
HOS|12|2|耶和華指控 猶大 ， 要照 雅各 所行的懲罰他， 按他所做的報應他。
HOS|12|3|他在腹中抓住哥哥的腳跟， 壯年的時候與上帝角力，
HOS|12|4|他與天使角力，並且得勝。 他曾哀哭，懇求施恩。 在 伯特利 遇見耶和華， 耶和華在那裏吩咐我們 ，
HOS|12|5|耶和華是萬軍之上帝， 耶和華是他可記念的名。
HOS|12|6|所以你當歸向你的上帝， 謹守慈愛和公平， 常常等候你的上帝。
HOS|12|7|商人 手持詭詐的天平， 喜愛欺壓。
HOS|12|8|以法蓮 說： 我果然富有，得了財寶； 我所勞碌得來的一切 人必找不到我有甚麼可算為有罪的惡。
HOS|12|9|自從你出 埃及 地以來， 我就是耶和華－你的上帝； 我必使你再住帳棚， 如同節期的日子一樣。
HOS|12|10|我已吩咐眾先知， 又增加異象， 藉先知設比喻。
HOS|12|11|基列 沒有罪孽嗎？ 他們誠然是虛假的， 在 吉甲 獻牛犢為祭； 他們的祭壇如同田間犁溝中的亂堆。
HOS|12|12|從前 雅各 逃到 亞蘭 地， 以色列 為娶妻子工作， 為娶妻子而牧放。
HOS|12|13|後來耶和華藉先知領 以色列 從 埃及 上來， 也藉先知看顧他們。
HOS|12|14|然而 以法蓮 大大惹動主怒， 他所流的血必歸到他身上。 主必使他的羞辱歸還給他。
HOS|13|1|從前 以法蓮 說話，人都戰兢， 他在 以色列 中居處高位； 但他因 巴力 犯罪就死了。
HOS|13|2|如今他們罪上加罪， 為自己鑄造偶像， 憑自己的聰明用銀子造偶像， 全都是匠人所製的。 論到它，有話說： 獻祭的人都要親吻牛犢。
HOS|13|3|因此，他們必如早晨的雲霧， 又如速散的露水， 如被狂風吹離禾場的糠秕， 又如煙囪冒出的煙。
HOS|13|4|自從你出 埃及 地以來， 我就是耶和華－你的上帝； 除了我上帝以外，你不認識別的， 在我以外，並沒有救主。
HOS|13|5|我曾在曠野， 就是那乾旱之地認識你。
HOS|13|6|他們得到餵養，就飽足； 既得飽足，就心高氣傲， 因而忘記了我。
HOS|13|7|因此我向他們如同獅子， 又如豹伏在道旁。
HOS|13|8|我如失去小熊的母熊，攻擊他們， 撕裂他們的胸膛。 在那裏我必如母獅吞吃他們， 如野獸撕開他們。
HOS|13|9|以色列 啊，你自取滅亡了 ， 因為我才是你的幫助。
HOS|13|10|現在，你的王在哪裏呢？ 讓他在你的各城中拯救你吧！ 你曾說「給我立君王和官長」， 那些治理你的又在哪裏呢？
HOS|13|11|我在怒氣中將王賜給你， 又在烈怒中將王廢去。
HOS|13|12|以法蓮 的罪孽被捲起來， 他的罪惡被收藏起來。
HOS|13|13|產婦的疼痛必臨到他身上； 他是無智慧之子， 如同臨盆時未出現的胎兒。
HOS|13|14|我必救贖他們脫離陰間， 救贖他們脫離死亡。 死亡啊，你的災害在哪裏？ 陰間哪，你的毀滅在哪裏？ 憐憫必從我眼前消逝。
HOS|13|15|他在弟兄中雖然旺盛， 卻有東風颳來， 就是耶和華的風從曠野上來。 他的泉源必乾涸， 他的源頭必枯竭， 這風必奪走他所積蓄的一切寶物。
HOS|13|16|撒瑪利亞 要擔當罪孽， 因為背叛自己的上帝。 他們必倒在刀下， 嬰孩必被摔死， 孕婦必被剖開。
HOS|14|1|以色列 啊，你要歸向耶和華－你的上帝， 你因自己的罪孽跌倒了。
HOS|14|2|當歸向耶和華， 用言語向他說： 「求你除盡罪孽，悅納善行， 我們就用嘴唇的祭代替牛犢獻上。
HOS|14|3|亞述 不能救我們， 我們不再騎馬， 也不再對我們手所造的偶像說： 『你是我們的上帝』； 孤兒在你那裏得蒙憐憫。」
HOS|14|4|我必醫治他們背道的病， 甘心愛他們， 因為我向他們所發的怒氣已轉消。
HOS|14|5|我必向 以色列 如甘露； 他必如百合花開放， 如 黎巴嫩 的樹扎根。
HOS|14|6|他的嫩枝必延伸， 他的榮華如橄欖樹， 香氣如 黎巴嫩 的香柏樹。
HOS|14|7|曾住在他蔭下的必歸回，使五穀生長 ， 他們要發旺如葡萄樹， 他的名氣 如 黎巴嫩 的酒。
HOS|14|8|以法蓮 說： 「我與偶像有何相干？」 我應允他，顧念他： 我如青翠的松樹， 你的果實從我而來。
HOS|14|9|智慧人必明白這些事， 聰明人必知道這一切。 耶和華的道是正直的， 義人行在其中， 罪人卻在其上跌倒。
JOEL|1|1|耶和華的話臨到 毗土珥 的兒子 約珥 。
JOEL|1|2|老年人哪，當聽這話； 這地所有的居民哪，要側耳而聽。 在你們的日子， 或你們祖先的日子， 曾發生過這樣的事嗎？
JOEL|1|3|你們要將這事傳與子， 子傳與孫， 孫傳與後代。
JOEL|1|4|剪蟲吃剩的，蝗蟲來吃； 蝗蟲吃剩的，蝻子來吃； 蝻子吃剩的，螞蚱 來吃。
JOEL|1|5|醉酒的人哪，要清醒，要哭泣； 好酒的人哪，都要為甜酒哀號， 因為酒從你們的口中斷絕了。
JOEL|1|6|有一隊蝗蟲 ，強盛且不可數， 上來侵犯我的地； 牠的牙齒如獅子的牙齒， 如母獅的大牙。
JOEL|1|7|牠毀壞我的葡萄樹， 撕裂我的無花果樹， 剝光又丟棄，使枝條露白。
JOEL|1|8|你要像童女腰束麻布， 為她年少時的丈夫哀號。
JOEL|1|9|耶和華的殿中斷絕素祭和澆酒祭， 事奉耶和華的祭司都悲哀。
JOEL|1|10|田荒涼，地悲哀； 因為五穀毀壞， 新酒枯竭， 新的油也缺乏。
JOEL|1|11|農夫啊，要慚愧； 修整葡萄園的啊，你們要哀號； 因為大麥、小麥與田間的莊稼全都毀了。
JOEL|1|12|葡萄樹枯乾， 無花果樹衰殘， 石榴樹、棕樹、蘋果樹， 田野一切的樹木都枯乾； 眾人的喜樂盡都消逝。
JOEL|1|13|祭司啊，當束上麻布痛哭； 事奉祭壇的啊，要哀號； 事奉我上帝的啊，你們要來，披上麻布過夜， 因為在你們上帝的殿中不再有素祭和澆酒祭了。
JOEL|1|14|你們要使禁食的日子分別為聖， 宣告嚴肅會， 召集長老和這地所有的居民 來到耶和華－你們上帝的殿， 向耶和華哀求。
JOEL|1|15|哀哉，這日子！ 因為耶和華的日子臨近， 好像毀滅從全能者來到。
JOEL|1|16|糧食不是在我們眼前斷絕了嗎？ 歡喜快樂不是從我們上帝的殿中止息了嗎？
JOEL|1|17|種子在土塊下朽爛， 倉荒涼，廩破壞， 因為五穀枯乾了。
JOEL|1|18|牲畜哀鳴， 牛群混亂，因無草場， 羊群也受苦。
JOEL|1|19|耶和華啊，我向你求告， 因為有火吞噬野地的草場， 火焰燒盡田野的樹木。
JOEL|1|20|田野的走獸切慕你， 因為溪水乾涸， 火吞噬了野地的草場。
JOEL|2|1|你們要在 錫安 吹角， 在我的聖山發出警報。 這地所有的居民要發顫， 因為耶和華的日子快到， 已經臨近了。
JOEL|2|2|那是黑暗、陰森的日子， 是密雲、烏黑的日子， 如同黎明籠罩山嶺。 有一隊蝗蟲，又大又強， 自古以來沒有像這樣的， 以後直到萬代也必沒有。
JOEL|2|3|牠們前面有火吞噬， 後面有火焰燒盡。 牠們未到以前，地如 伊甸園 ， 過去以後，卻成了荒涼的曠野， 沒有一樣能躲避牠們。
JOEL|2|4|牠們形狀如馬， 奔跑如戰馬。
JOEL|2|5|響聲如戰車在山頂上跳動， 如火焰吞噬碎秸， 好像強大的軍隊擺陣備戰。
JOEL|2|6|在牠們面前，萬民傷慟， 臉都變色。
JOEL|2|7|牠們如勇士奔跑， 如戰士攀登城牆， 各行於自己的道路， 不亂隊伍；
JOEL|2|8|牠們並不彼此推擠， 各行於自己的大道， 衝過防禦 ， 並不停止。
JOEL|2|9|牠們蹦上城， 跳上牆， 爬上房屋， 從窗戶進來，如同盜賊。
JOEL|2|10|在牠們面前， 地動天搖， 日月昏暗， 星宿無光。
JOEL|2|11|耶和華在他的軍旅前出聲， 他的隊伍龐大， 遵行他命令的強盛。 耶和華的日子大而可畏， 誰能當得起呢？
JOEL|2|12|然而你們現在要禁食，哭泣，哀號， 一心歸向我。 這是耶和華說的。
JOEL|2|13|你們要撕裂心腸， 不要撕裂衣服。 歸向耶和華－你們的上帝， 因為他有恩惠，有憐憫， 不輕易發怒， 有豐盛的慈愛， 並且會改變心意， 不降那災難。
JOEL|2|14|誰知道他也許會回心轉意，留下餘福， 就是獻給耶和華－你們上帝的素祭和澆酒祭。
JOEL|2|15|你們要在 錫安 吹角， 使禁食的日子分別為聖， 宣告嚴肅會。
JOEL|2|16|聚集百姓，使會眾自潔； 召集老年人， 聚集孩童和在母懷吃奶的； 使新郎出內室， 新娘離開洞房。
JOEL|2|17|事奉耶和華的祭司 要在走廊和祭壇間哭泣，說： 「耶和華啊，求你顧惜你的百姓， 不要使你的產業受羞辱， 在列國中成為笑柄。 為何讓人在萬民中說 『他們的上帝在哪裏』呢？」
JOEL|2|18|耶和華為自己的地發熱心， 憐憫他的百姓。
JOEL|2|19|耶和華應允他的百姓說： 「看哪，我要賞賜你們五穀、新酒和新的油， 使你們飽足， 我必不再使你們受列國的羞辱。
JOEL|2|20|我要使北方來的隊伍遠離你們， 將他們趕到乾旱荒蕪之地： 前隊趕入東海， 後隊趕入西海； 臭氣上升，惡臭騰空。 耶和華果然行了大事！
JOEL|2|21|「土地啊，不要懼怕， 要歡喜快樂， 因為耶和華行了大事。
JOEL|2|22|田野的走獸啊，不要懼怕， 因為曠野的草已生長， 樹木結果， 無花果樹、葡萄樹也都效力 。
JOEL|2|23|「 錫安 的民哪，你們要歡喜， 要因耶和華－你們的上帝快樂； 因他賞賜你們合宜的秋雨 ， 為你們降下甘霖， 秋雨和春雨，和先前一樣。
JOEL|2|24|「禾場充滿五穀， 池中漫溢新酒和新的油。
JOEL|2|25|我差遣到你們中間的大軍隊， 就是蝗蟲、蝻子、螞蚱、剪蟲， 那些年間所吃的，我要補還給你們。
JOEL|2|26|「你們必吃得飽足， 讚美耶和華－你們上帝的名， 他為你們行了奇妙的事。 我的百姓不致羞愧，直到永遠。
JOEL|2|27|你們必知道我是在 以色列 中， 又知道我是耶和華－你們的上帝，沒有別的。 我的百姓不致羞愧，直到永遠。」
JOEL|2|28|「以後，我要將我的靈澆灌凡有血肉之軀的。 你們的兒女要說預言， 你們的老人要做異夢， 你們的少年要見異象。
JOEL|2|29|在那些日子， 我要將我的靈澆灌我的僕人和婢女。
JOEL|2|30|「我要在天上地下顯出奇事，有血，有火，有煙柱。
JOEL|2|31|太陽要變為黑暗，月亮要變為血，這都在耶和華大而可畏的日子未到以前。
JOEL|2|32|那時，凡求告耶和華名的就必得救；因為照耶和華所說的，在 錫安山 ，在 耶路撒冷 將有逃脫的人。凡耶和華所召的 ，都在餘民之列。」
JOEL|3|1|「看哪，在那些日子，到那個時候，我使 猶大 和 耶路撒冷 被擄之人歸回的時候，
JOEL|3|2|我要聚集萬民，帶他們下到 約沙法谷 去，在那裏我要為我百姓，我產業 以色列 的緣故，向萬民施行審判；因為他們把我的百姓分散到列國，瓜分了我的土地，
JOEL|3|3|為我的百姓抽籤，以男孩換取妓女，為喝酒賣掉女孩。
JOEL|3|4|「 推羅 、 西頓 和 非利士 四境的人哪，你們與我何干？你們要報復我嗎？若要報復我，我必使報應速速歸到你們頭上。
JOEL|3|5|你們奪取我的金銀，把我珍貴的寶物帶入你們的廟宇 ，
JOEL|3|6|並將 猶大 人和 耶路撒冷 人賣給 希臘 人 ，使他們遠離自己的疆土。
JOEL|3|7|看哪，我必激發他們離開你們把他們賣去的地方，又必使報應歸到你們頭上。
JOEL|3|8|我要將你們的兒女賣到 猶大 人手中，他們必轉賣給遠方的國家 示巴 人。這是耶和華說的。」
JOEL|3|9|當在列國中宣告： 預備打仗， 激發勇士， 使所有戰士上前來。
JOEL|3|10|要將犁頭打成刀劍， 鐮刀打成戈矛； 弱者要說：「我是勇士。」
JOEL|3|11|四圍的列國啊， 要速速前來， 一同聚集。 耶和華啊， 求你使你的勇士降臨。
JOEL|3|12|列國都當興起， 上到 約沙法谷 ； 因為我必坐在那裏， 審判四圍的列國。
JOEL|3|13|揮鐮刀吧！因為莊稼熟了； 來踩踏吧！因為醡酒池滿了。 酒池已經滿溢， 因為他們的罪惡甚大。
JOEL|3|14|在 斷定谷 有許多許多的人， 因為耶和華的日子臨近 斷定谷 了。
JOEL|3|15|日月昏暗， 星宿無光。
JOEL|3|16|耶和華必從 錫安 吼叫， 從 耶路撒冷 出聲， 天地就震動。 耶和華卻要作他百姓的避難所， 作 以色列 人的保障。
JOEL|3|17|你們就知道我是耶和華－你們的上帝， 我住在 錫安 －我的聖山。 耶路撒冷 必成為聖； 陌生人不再從其中經過。
JOEL|3|18|在那日，大山要滴甜酒， 小山要流奶， 猶大 的溪河都有水流出； 必有泉源從耶和華的殿中流出， 滋潤 什亭谷 。
JOEL|3|19|埃及 必定荒涼， 以東 成為荒涼的曠野， 因為他們向 猶大 人行殘暴， 又因他們在本地流無辜人的血。
JOEL|3|20|但 猶大 必存到永遠， 耶路撒冷 必存到萬代。
JOEL|3|21|我要免除 流人血的罪， 是先前未曾免除的， 耶和華居住在 錫安 。
AMOS|1|1|這是 猶大 王 烏西雅 在位與 約阿施 的兒子 以色列 王 耶羅波安 在位的時候，大地震前二年，從 提哥亞 來的牧人 阿摩司 所見的─他的話論到 以色列 。
AMOS|1|2|他說：「耶和華必從 錫安 吼叫， 從 耶路撒冷 出聲； 牧人的草場哀傷， 迦密 的山頂枯乾。」
AMOS|1|3|耶和華如此說： 「 大馬士革 三番四次犯罪， 以鐵的打穀機擊打 基列 ， 我必不撤銷對它的懲罰。
AMOS|1|4|我要降火在 哈薛 的王宮， 吞滅 便‧哈達 的宮殿；
AMOS|1|5|我要折斷 大馬士革 的門閂， 剪除 亞文 平原的居民 和 伯‧伊甸 的掌權者， 亞蘭 人必被擄到 吉珥 。」 這是耶和華說的。
AMOS|1|6|耶和華如此說： 「 迦薩 三番四次犯罪， 擄掠全體百姓交給 以東 ， 我必不撤銷對它的懲罰。
AMOS|1|7|我要降火在 迦薩 城內， 吞滅它的宮殿；
AMOS|1|8|我要剪除 亞實突 的居民 和 亞實基倫 的掌權者， 反手攻擊 以革倫 ， 剩餘的 非利士 人都必滅亡。」 這是主耶和華說的。
AMOS|1|9|耶和華如此說： 「 推羅 三番四次犯罪， 將全體百姓交給 以東 ， 不顧念弟兄的盟約， 我必不撤銷對它的懲罰，
AMOS|1|10|我要降火在 推羅 城內， 吞滅它的宮殿。」
AMOS|1|11|耶和華如此說： 「 以東 三番四次犯罪， 怒氣不停發作，永遠懷著憤怒， 拿刀追趕兄弟，絲毫不存憐憫， 我必不撤銷對它的懲罰。
AMOS|1|12|我要降火在 提幔 ， 吞滅 波斯拉 的宮殿。」
AMOS|1|13|耶和華如此說： 「 亞捫 人三番四次犯罪， 剖開 基列 的孕婦， 擴張自己的疆界， 我必不撤銷對它的懲罰。
AMOS|1|14|我要在戰爭吶喊的日子， 在旋風狂吹時， 在 拉巴 城內放火， 吞滅它的宮殿；
AMOS|1|15|他們的君王和官長必一同被擄。」 這是耶和華說的。
AMOS|2|1|耶和華如此說： 「 摩押 三番四次犯罪， 把 以東 王的骸骨焚燒成灰， 我必不撤銷對它的懲罰。
AMOS|2|2|我要降火在 摩押 ， 吞滅 加略 的宮殿， 摩押 必在鬧鬨、吶喊、吹角聲中滅亡；
AMOS|2|3|我要剪除 摩押 的領袖， 把所有的官長和他一同殺戮。」 這是耶和華說的。
AMOS|2|4|耶和華如此說： 「 猶大 三番四次犯罪， 厭棄耶和華的訓誨， 不遵守他的律例； 他們祖先所隨從虛假的偶像 使他們走迷了， 我必不撤銷對它的懲罰。
AMOS|2|5|我要降火在 猶大 ， 吞滅 耶路撒冷 的宮殿。」
AMOS|2|6|耶和華如此說： 「 以色列 三番四次犯罪， 為銀子賣了義人， 為一雙鞋賣了窮人， 我必不撤銷對它的懲罰。
AMOS|2|7|他們把貧寒人的頭踐踏在地的塵土上 ， 又阻礙困苦人的道路。 父子與同一個女子行淫， 以致褻瀆我的聖名。
AMOS|2|8|他們在各祭壇旁邊， 躺臥在人所典當的衣服上， 又在他們上帝的殿裏 喝受罰之人的酒。
AMOS|2|9|「我從他們面前除滅 亞摩利 人； 他雖高大如香柏樹，強壯如橡樹， 我卻上滅其果，下絕其根。
AMOS|2|10|我曾將你們從 埃及 地領上來， 在曠野裏引導你們四十年， 使你們得 亞摩利 人之地為業；
AMOS|2|11|我從你們子孫中興起先知， 又從你們少年中興起拿細耳人。 以色列 人哪，不是這樣嗎？」 這是耶和華說的。
AMOS|2|12|「你們卻把酒給拿細耳人喝， 囑咐先知說：『不要說預言。』
AMOS|2|13|「看哪，我要把你們壓下去， 如同裝滿禾捆的車壓過一樣。
AMOS|2|14|快跑的無從避難， 壯士無法使力， 勇士也不能自救；
AMOS|2|15|拿弓的站立不住， 腿快的不能逃脫， 騎馬的也不能自救。
AMOS|2|16|到那日，勇士中最有膽量的， 必赤身逃跑。」 這是耶和華說的。
AMOS|3|1|以色列 人哪，當聽耶和華責備你們的話，責備我從 埃及 地領上來的全家，說：
AMOS|3|2|「在地上萬族中，我只認識你們； 因此，我必懲罰你們一切的罪孽。」
AMOS|3|3|二人若不同心， 豈能同行呢？
AMOS|3|4|獅子若無獵物， 豈會在林中咆哮呢？ 少壯獅子若無所得， 豈會從洞裏吼叫呢？
AMOS|3|5|若未設圈套， 雀鳥豈能陷入地上的羅網呢？ 羅網若無所得， 豈會從地上翻起呢？
AMOS|3|6|城中若吹角， 百姓豈不戰兢嗎？ 災禍若臨到一城， 豈非耶和華所降的嗎？
AMOS|3|7|主耶和華不會做任何事情， 除非先將奧祕指示他的僕人眾先知。
AMOS|3|8|獅子吼叫，誰不懼怕呢？ 主耶和華既已說了，誰能不說預言呢？
AMOS|3|9|你們要在 亞實突 的宮殿 和 埃及 地的宮殿傳揚，說： 「要聚集在 撒瑪利亞 的山上， 看城裏有何等大的擾亂與欺壓。」
AMOS|3|10|「他們以暴力搶奪， 堆積在自己的宮殿裏， 卻不懂得行正直的事。」 這是耶和華說的。
AMOS|3|11|所以主耶和華如此說： 「敵人必來圍攻這地， 削弱你的勢力， 搶掠你的宮殿。」
AMOS|3|12|耶和華如此說：「牧人怎樣從獅子口中搶回兩條腿或耳朵的一小片，住 撒瑪利亞 的 以色列 人得救也是如此，不過搶回床的一角和床榻的靠枕 而已。」
AMOS|3|13|主耶和華－萬軍之上帝說： 「當聽這話，警戒 雅各 家。
AMOS|3|14|我懲罰 以色列 罪孽的日子， 也要懲罰 伯特利 的祭壇； 祭壇的角必被砍下，墜落於地。
AMOS|3|15|我要拆毀過冬和避暑的房屋， 象牙的房屋必毀滅， 廣廈豪宅都歸無有。」 這是耶和華說的。
AMOS|4|1|「你們這些 撒瑪利亞山 上的 巴珊 母牛啊， 當聽這話！ 你們欺負貧寒人，壓碎貧窮人， 對主人說：『拿酒來，我們喝吧！』
AMOS|4|2|主耶和華指著自己的神聖起誓說： 『看哪，日子將到，人必用鉤子將你們鉤去， 用魚鉤把你們中最後一個鉤去。
AMOS|4|3|你們必從城牆的缺口 出去， 各人直往前行， 投向 哈門 。』」 這是耶和華說的。
AMOS|4|4|「 以色列 人哪，任你們往 伯特利 去犯罪， 到 吉甲 增加罪過， 每早晨獻上你們的祭物， 每三日納你們的十一奉獻；
AMOS|4|5|任你們獻上有酵的感謝祭， 宣揚你們的甘心祭，使人聽見， 因為這是你們所喜愛的。」 這是主耶和華說的。
AMOS|4|6|「我使你們在每一座城裏牙齒乾淨， 使你們各處的糧食缺乏， 你們仍不歸向我。」 這是耶和華說的。
AMOS|4|7|「在收割的前三個月， 我不降雨在你們那裏， 我降雨在這城， 不降雨在那城； 這塊地有雨， 那塊無雨的地就必枯乾。
AMOS|4|8|兩三城的人擠到一個城去找水喝， 卻喝不足， 你們仍不歸向我。」 這是耶和華說的。
AMOS|4|9|「我以焚風 和霉爛攻擊你們， 你們許多的菜園、葡萄園、 無花果樹、橄欖樹屢屢被剪蟲 所吃， 你們仍不歸向我。」 這是耶和華說的。
AMOS|4|10|「我降瘟疫在你們中間， 如在 埃及 的樣子； 用刀殺戮你們的年輕人 和你們遭擄掠的馬匹， 營中臭氣撲鼻， 你們仍不歸向我。」 這是耶和華說的。
AMOS|4|11|「我傾覆你們， 如同上帝從前傾覆 所多瑪 、 蛾摩拉 一樣； 你們好像從火中搶救出來的一根柴， 你們仍不歸向我。」 這是耶和華說的。
AMOS|4|12|「因此， 以色列 啊，我要如此對待你； 因為我要這樣對待你， 以色列 啊， 你當預備迎見你的上帝。」
AMOS|4|13|看哪，那創山，造風，將其心意指示人， 使晨光變幽暗，踩行在地之高處的， 他的名是耶和華－萬軍之上帝。
AMOS|5|1|以色列 家啊，聽我為你們所作的哀歌：
AMOS|5|2|「 以色列 民 跌倒，不得再起； 躺在地上，無人扶起。」
AMOS|5|3|主耶和華如此說： 「 以色列 家的城派出一千，只剩一百； 派出一百，只剩十個。」
AMOS|5|4|耶和華向 以色列 家如此說： 「你們要尋求我，就必存活。
AMOS|5|5|不要往 伯特利 尋求， 不要進入 吉甲 ， 也不要過到 別是巴 ； 因為 吉甲 必被擄走， 伯特利 必歸無有。」
AMOS|5|6|要尋求耶和華，就必存活， 免得他在 約瑟 家如火發出， 焚燒 伯特利 ，無人撲滅。
AMOS|5|7|你們這使公平變為茵蔯， 將公義丟棄於地的人哪！
AMOS|5|8|那造昴星和參星， 使死蔭變為晨光， 使白晝變為黑夜， 召喚海水、 使其傾倒在地面上的， 耶和華是他的名。
AMOS|5|9|他快速摧毀強壯的人， 毀滅就臨到堡壘。
AMOS|5|10|你們怨恨那在城門口斷是非的， 憎惡那說正直話的。
AMOS|5|11|所以，因你們踐踏貧寒人， 向他們勒索糧稅； 你們雖建造石鑿的房屋， 卻不得住在其內； 雖栽植美好的葡萄園， 卻不得喝其中所出的酒。
AMOS|5|12|我知道你們的罪過何其多， 你們的罪惡何其大； 你們迫害義人，收受賄賂， 在城門口屈枉貧窮人。
AMOS|5|13|所以智慧人在這樣的時候必靜默不言， 因為這是險惡的時候。
AMOS|5|14|你們要尋求良善， 不要尋求邪惡，就必存活。 這樣，耶和華－萬軍之上帝 必照你們所說的與你們同在。
AMOS|5|15|要恨惡邪惡，喜愛良善， 在城門口秉公行義； 或者耶和華－萬軍之上帝 會施恩給 約瑟 的餘民。
AMOS|5|16|因此，主耶和華－萬軍之上帝如此說： 「在一切的廣場上必有哀號的聲音； 在各街市上必有人說： 『哀哉！哀哉！』 他們叫農夫來哭號， 叫善唱哀歌的來舉哀；
AMOS|5|17|各葡萄園都有哀號的聲音， 因為我必從你中間經過。」 這是耶和華說的。
AMOS|5|18|想望耶和華日子的人有禍了！ 為甚麼你們要耶和華的日子呢？ 那是黑暗沒有光明的日子，
AMOS|5|19|好像人躲避獅子卻遇見熊； 進房屋以手靠牆，卻被蛇咬。
AMOS|5|20|耶和華的日子豈不是黑暗沒有光明， 幽暗毫無光輝嗎？
AMOS|5|21|「我厭惡你們的節期， 也不喜悅你們的嚴肅會。
AMOS|5|22|你們雖然向我獻燔祭和素祭， 我卻不悅納， 也不看你們用肥畜獻的平安祭。
AMOS|5|23|要使你們歌唱的聲音遠離我， 因為我不聽你們琴瑟的樂曲。
AMOS|5|24|惟願公平如大水滾滾， 公義如江河滔滔。
AMOS|5|25|「 以色列 家啊，你們在曠野四十年，何嘗將祭物和供物獻給我呢？
AMOS|5|26|你們抬著你們的 撒古特 君王 ，和你們為自己所造之偶像 迦溫 ，你們的神明之星。
AMOS|5|27|所以我要把你們擄到 大馬士革 以外。」這是耶和華說的，他的名為萬軍之上帝。
AMOS|6|1|「那在 錫安 安逸， 在 撒瑪利亞山 安穩， 為列國之首，具有名望， 且為 以色列 家所歸向的，有禍了！
AMOS|6|2|你們要過到 甲尼 察看， 從那裏往 哈馬 大城去， 又下到 非利士 人的 迦特 ， 你們比這些國更好嗎？ 或是他們的疆界比你們的疆界廣大呢？
AMOS|6|3|你們以為降禍的日子尚遠， 卻使殘暴的統治 臨近。
AMOS|6|4|「那些躺臥在象牙床上，舒身在榻上的， 吃群中的羔羊和棚裏的牛犢。
AMOS|6|5|他們以琴瑟逍遙歌唱， 為自己作曲 ，像 大衛 一樣；
AMOS|6|6|以大碗喝酒，用上等油抹身， 卻不為 約瑟 所受的苦難憂傷；
AMOS|6|7|所以，現在這些人必首先被擄， 逍遙的歡宴必消失。」
AMOS|6|8|主耶和華指著自己起誓說： 「我憎惡 雅各 的驕傲，厭棄他的宮殿； 我必將城和其中一切所有的都交給敵人。」 這是耶和華－萬軍之上帝說的 。
AMOS|6|9|那時，若一房之內剩下十個人，也都必死。
AMOS|6|10|死人的叔伯要把屍首抬到屋外焚燒，就問房屋內間的人說：「你那裏還有別人嗎？」他說：「沒有。」又說：「不要作聲，不可提耶和華的名。」
AMOS|6|11|看哪，耶和華發命令， 把大房子拆成碎片， 小屋子裂為小塊。
AMOS|6|12|馬豈能在巖石上奔跑？ 人豈能在那裏 用牛耕種呢？ 你們卻使公平變為苦膽， 使公義的果子變為茵蔯。
AMOS|6|13|你們這些喜愛 羅‧底巴 的，自誇說： 「我們不是憑自己的力量攻佔了 加寧 嗎？」
AMOS|6|14|耶和華─萬軍之上帝說： 「 以色列 家，看哪，我必興起一國攻擊你們； 他們必欺壓你們， 從 哈馬口 直到 亞拉巴 的河。」
AMOS|7|1|主耶和華指示我一件事，在春天作物剛長出時，看哪，主 造了蝗蟲；看哪，這是王收割後長出的春天作物。
AMOS|7|2|蝗蟲吃盡那地青草的時候，我說： 「主耶和華啊，求你赦免； 因為 雅各 弱小， 他怎能站立得住呢？」
AMOS|7|3|耶和華對這事改變心意， 耶和華說：「這災可以免了。」
AMOS|7|4|主耶和華又指示我一件事，看哪，主耶和華命火施行審判，火就吞滅深淵，燒盡產業。
AMOS|7|5|我就說： 「主耶和華啊，求你止息； 因為 雅各 弱小， 他怎能站立得住呢？」
AMOS|7|6|耶和華對這事改變心意， 主耶和華說：「這災也可免了。」
AMOS|7|7|他又指示我一件事，看哪，主手拿鉛垂線，站立在依鉛垂線建好的牆邊。
AMOS|7|8|耶和華對我說：「 阿摩司 ，你看見甚麼？」我說：「鉛垂線。」主說： 「看哪，我要在我子民 以色列 中 吊起鉛垂線， 不再寬恕他們。
AMOS|7|9|以撒 的丘壇必荒涼， 以色列 的聖所必荒廢； 我要起來用刀攻擊 耶羅波安 的家。」
AMOS|7|10|伯特利 的祭司 亞瑪謝 派人到 以色列 王 耶羅波安 那裏，說：「 阿摩司 在 以色列 家中圖謀背叛你，他所說的一切話，這地不能承擔；
AMOS|7|11|因為 阿摩司 這樣說： 『 耶羅波安 必被刀殺， 以色列 百姓必被擄， 離開本地。』」
AMOS|7|12|於是 亞瑪謝 對 阿摩司 說：「你這先見哪，要逃到 猶大 地，在那裏過活 ，在那裏說預言；
AMOS|7|13|卻不要在 伯特利 再說預言，因為這裏有王的聖所，有王的宮殿。」
AMOS|7|14|阿摩司 對 亞瑪謝 說：「我原不是先知，也不是先知的門徒；我是牧人，是修剪桑樹的。
AMOS|7|15|耶和華帶領我，叫我不再牧放羊群，對我說：『你去向我子民 以色列 說預言。』
AMOS|7|16|「現在你要聽耶和華的話。 你說：『不要向 以色列 說預言， 也不要向 以撒 家傳講 。』
AMOS|7|17|所以耶和華如此說： 『你的妻子要在城中作妓女， 你的兒女要倒在刀下； 你的地必有人用繩子量了瓜分， 你自己必死在不潔淨之地； 以色列 百姓必被擄， 離開本地。』」
AMOS|8|1|主耶和華又指示我一件事，看哪，有一筐夏天的果子。
AMOS|8|2|他說：「 阿摩司 ，你看見甚麼？」我說：「一筐夏天的果子。」耶和華對我說： 「我子民 以色列 的結局 到了， 我必不再寬恕他們。
AMOS|8|3|那日，宮殿裏的詩歌要變為哀號 ； 必有許多屍首拋在各處， 安靜無聲。」 這是主耶和華說的。
AMOS|8|4|你們這些踐踏貧窮人、 使這地困苦人衰敗的， 當聽這話！
AMOS|8|5|你們說：「初一幾時過去， 我們好賣糧； 安息日幾時過去， 我們好擺開穀物； 我們要把伊法變小， 把舍客勒變大， 以詭詐的天平欺哄人，
AMOS|8|6|用銀子買貧寒人， 以一雙鞋換貧窮人， 把壞的穀物賣給人。」
AMOS|8|7|耶和華指著 雅各 的驕傲起誓說： 「他們這一切的行為，我必永遠不忘。
AMOS|8|8|地豈不因這事震動？ 其中的居民豈不悲哀嗎？ 全地必如 尼羅河 漲起， 如 埃及 的 尼羅河 湧起退落。
AMOS|8|9|「到那日， 我要使太陽在正午落下， 使這地在白晝黑暗。」 這是主耶和華說的。
AMOS|8|10|「我要使你們的節期變為悲哀， 你們一切的歌曲變為哀歌； 我要使眾人腰束麻布， 頭上光禿； 我要使這悲哀如喪獨子， 其結局如悲痛的日子。
AMOS|8|11|「看哪，日子將到， 我必命饑荒降在地上； 人飢餓非因無餅，乾渴非因無水， 而是因不聽耶和華的話。」 這是主耶和華說的。
AMOS|8|12|他們必飄流，從這海到那海， 從北邊到東邊，往來奔跑， 尋求耶和華的話， 卻尋不著。
AMOS|8|13|「當那日，少年和美貌的少女 必因乾渴而發昏。
AMOS|8|14|那些指著 撒瑪利亞 的罪孽 起誓的，說： 『 但 哪，我們指著你那裏的神明起誓』， 又說：『我們指著通往 別是巴 的路起誓』， 這些人都必仆倒，永不再起。」
AMOS|9|1|我看見主站在祭壇旁，說： 「你要擊打柱頂，使門檻震動， 要剪除眾人當中為首的， 他們中最後的 ，我必用刀殺戮； 無一人能逃避，無一人能逃脫。
AMOS|9|2|「雖然他們挖透陰間， 我的手必從那裏拉出他們； 雖然他們爬到天上， 我必從那裏拿下他們；
AMOS|9|3|雖然藏在 迦密山 頂， 我必在那裏搜尋，擒拿他們； 雖然離開我眼前藏在海底， 我必在那裏命令蛇咬他們；
AMOS|9|4|雖然被仇敵擄去， 我也必在那裏命令刀劍殺戮他們； 我必定睛在他們身上， 降禍不降福。」
AMOS|9|5|萬軍的主耶和華觸摸地，地就融化， 凡住在地上的都必悲哀； 全地必如 尼羅河 漲起， 如同 埃及 的 尼羅河 落下。
AMOS|9|6|那在天上建造樓閣、 在地上奠定穹蒼、 召喚海水、 使其傾倒在地面上的， 耶和華是他的名。
AMOS|9|7|耶和華說：「 以色列 人哪， 我豈不是看你們如 古實 人嗎？ 我豈不是領 以色列 人出 埃及 地， 也領 非利士 人出 迦斐託 ， 領 亞蘭 人出 吉珥 嗎？
AMOS|9|8|看哪，主耶和華的眼目 察看這有罪的國度， 要把它從地面上滅絕， 卻不將 雅各 家滅絕淨盡。」 這是耶和華說的。
AMOS|9|9|「看哪，我發命令， 使 以色列 家在萬國中飄流， 好像人用篩子篩穀， 連一粒也不落在地上。
AMOS|9|10|我子民中所有的罪人， 就是那些說 『災禍必不靠近，必不追上我們』的， 都必死在刀下。」
AMOS|9|11|「在那日，我必重建 大衛 倒塌的帳幕， 修補其中的缺口； 我必建立那遭破壞的， 重新修造，如古時一般，
AMOS|9|12|使 以色列 人接管 以東 所剩餘的 和所有稱為我名下的國。 這是耶和華說的，他要行這事。
AMOS|9|13|「看哪，日子將到， 耕種的必接續收割的， 踹葡萄的必接續撒種的； 大山要滴下甜酒， 小山也被漫過。」 這是耶和華說的。
AMOS|9|14|「我要使 以色列 被擄的子民歸回； 他們要重修荒廢的城鎮， 居住在其中； 栽植葡萄園，喝其中所出的酒， 修造果園，吃其中的果子。
AMOS|9|15|我要將他們栽植於本地， 他們必不再從我所賜給他們的地上被拔出。」 這是耶和華－你的上帝說的。
OBAD|1|1|俄巴底亞 所見的異象。 我們從耶和華那裏得到消息， 有使者被差往列國去： 「起來吧， 我們要起來與 以東 爭戰！」 主耶和華論 以東 如此說：
OBAD|1|2|看哪，我要使你在列國中為最小， 被人大大藐視。
OBAD|1|3|你狂傲的心欺騙了你， 你住在巖穴， 居所在高處， 心裏說： 「誰能把我拉下來到地上呢？」
OBAD|1|4|你雖如鷹高飛， 在星宿之間搭窩， 我必從那裏拉你下來。 這是耶和華說的。
OBAD|1|5|盜賊若來到你那裏， 小偷夜間來到， 豈不是只偷他們所需要的嗎？ 摘葡萄的若來到你那裏， 豈不留下幾串嗎？ 你竟全然滅絕！
OBAD|1|6|以掃 遭到搜查， 他隱藏的寶物竟被尋出！
OBAD|1|7|與你結盟的都驅趕你，直到邊界， 與你和好的欺騙你，勝過你， 吃你飯的人設下圈套陷害你─ 他卻毫無聰明 。
OBAD|1|8|到那日， 我豈不從 以東 除滅智慧人？ 從 以掃山 除滅聰明人？ 這是耶和華說的。
OBAD|1|9|提幔 哪， 你的勇士必驚惶， 以致 以掃山 的人都被殺戮剪除。
OBAD|1|10|因你向兄弟 雅各 施暴， 你必蒙羞， 永被剪除。
OBAD|1|11|當陌生人擄掠 雅各 的財物， 當外邦人進入他的城門， 為 耶路撒冷 抽籤分取財物的日子， 你竟站在一旁，像與他們同夥。
OBAD|1|12|你兄弟遭難的日子， 你不該瞪著眼看； 猶大 人被滅的日子， 你不該幸災樂禍； 他們遭難的日子， 你不該說狂傲的話。
OBAD|1|13|我子民遭災的日子， 你不該進他們的城門； 他們遭災的日子， 你不該瞪著眼看他們受苦； 他們遭災的日子， 你不該伸手搶他們的財物。
OBAD|1|14|他們遭難的日子， 你不該站在岔路口 剪除他們逃脫的人， 你不該交出他們的倖存者。
OBAD|1|15|耶和華的日子臨近萬國； 你所做的，人也必向你照樣做， 你的報應必歸到自己頭上。
OBAD|1|16|你們在我聖山怎樣喝了苦杯， 萬國必照樣不停地喝， 且喝且吞， 他們就必歸於無有。
OBAD|1|17|但在 錫安山 必有逃脫的人， 那山必成為聖； 雅各 家必得原有的產業 。
OBAD|1|18|雅各 家必成為大火， 約瑟 家成為火焰； 以掃 家必如碎秸， 遭燃燒，被吞滅， 以掃 家必無倖存者。 這是耶和華說的。
OBAD|1|19|他們必得 尼革夫 和 以掃山 ， 得 謝非拉 ， 非利士 人之地， 他們必得 以法蓮 地和 撒瑪利亞 地， 得 便雅憫 和 基列 ；
OBAD|1|20|被擄的 以色列 大軍 必得 迦南 人的地，直到 撒勒法 ， 在 西法拉 被擄的 耶路撒冷 人 必得 尼革夫 的城鎮。
OBAD|1|21|必有一些解救者 上到 錫安山 ，審判 以掃山 ， 國度就歸耶和華了。
JONAH|1|1|耶和華的話臨到 亞米太 的兒子 約拿 ，說：
JONAH|1|2|「起來，到 尼尼微 大城去，向其中的居民宣告，因為他們的惡已達到我面前。」
JONAH|1|3|約拿 卻起身，逃往 他施 去躲避耶和華。他下到 約帕 ，遇見一條船要往 他施 去。 約拿 付了船費，就上船，與船上的人同往 他施 ，為要躲避耶和華。
JONAH|1|4|耶和華在海上颳起大風，海就狂風大作，船幾乎破裂。
JONAH|1|5|水手都懼怕，各人哀求自己的神明。他們把船上的貨物拋進海裏，為要減輕載重。 約拿 卻下到艙底，躺臥沉睡。
JONAH|1|6|船長到他那裏，對他說：「你怎麼還在沉睡呢？起來，求告你的神明，或者神明顧念我們，使我們不致滅亡。」
JONAH|1|7|船上的人彼此說：「來吧，我們來抽籤，看看這災難臨到我們是因誰的緣故。」於是他們就抽籤，抽出 約拿 來。
JONAH|1|8|他們對 約拿 說：「請你告訴我們，這災難臨到我們是因誰的緣故呢？你做甚麼行業？你從哪裏來？你是哪一國的人？屬哪一族？」
JONAH|1|9|他說：「我是 希伯來 人，我敬畏耶和華，天上的上帝，他創造了滄海和陸地。」
JONAH|1|10|那些人就大大懼怕，對他說：「你做的是甚麼事呢？」原來他們已經知道他在躲避耶和華，因為他告訴了他們。
JONAH|1|11|海浪越來越洶湧，他們就問他說：「我們當向你做甚麼，才能使海浪平靜呢？」
JONAH|1|12|他對他們說：「你們把我抬起來，拋進海裏，海就會平靜了；我知道你們遭遇這大風浪是因我的緣故。」
JONAH|1|13|然而那些人竭力划槳，想要把船靠回陸地，卻是不能；因風浪愈來愈大，撲向他們。
JONAH|1|14|於是他們求告耶和華說：「耶和華啊，求求你不要因這人的性命使我們滅亡，不要使流無辜人血的罪歸給我們；因為你－耶和華隨自己的旨意行事。」
JONAH|1|15|他們把 約拿 抬起來，拋進海裏，海的狂浪就平息了。
JONAH|1|16|那些人就大大懼怕耶和華，向耶和華獻祭許願。
JONAH|1|17|耶和華安排一條大魚吞下 約拿 ， 約拿 在魚腹中三日三夜。
JONAH|2|1|約拿 在魚腹中向耶和華－他的上帝禱告，
JONAH|2|2|說： 「我在患難中求告耶和華， 他就應允我； 我從陰間的深處呼求， 你就俯聽我的聲音。
JONAH|2|3|你將我投下深淵， 直到海心； 大水環繞我， 你的波浪洪濤漫過我身。
JONAH|2|4|我說：『我從你眼前被驅逐， 然而我仍要仰望你的聖殿。』
JONAH|2|5|眾水環繞我，幾乎淹沒我； 深淵圍住我； 海草纏繞我的頭。
JONAH|2|6|我下沉到山的根基， 地的門閂將我永遠關住。 耶和華－我的上帝啊， 你卻將我的性命從地府裏救出來。
JONAH|2|7|我心靈發昏時， 就想起耶和華。 我的禱告進入你的聖殿， 達到你面前。
JONAH|2|8|那信奉虛無神明 的人， 丟棄自己的慈愛；
JONAH|2|9|但我要以感謝的聲音向你獻祭。 我所許的願，我必償還。 救恩出於耶和華。」
JONAH|2|10|耶和華吩咐那魚，魚就把 約拿 吐在陸地上。
JONAH|3|1|耶和華的話第二次臨到 約拿 ，說：
JONAH|3|2|「起來，到 尼尼微 大城去，把我告訴你的信息向其中的居民宣告。」
JONAH|3|3|約拿 就照耶和華的話起來，到 尼尼微 去。 尼尼微 是一座極大的城，約有三天的路程。
JONAH|3|4|約拿 進城，走了一天，宣告說：「再過四十天， 尼尼微 要傾覆了！」
JONAH|3|5|尼尼微 人就信服上帝，宣告禁食，從最大的到最小的都穿上麻衣。
JONAH|3|6|這消息傳到 尼尼微 王那裏，他就從寶座起來，脫下朝服，披上麻布，坐在灰中。
JONAH|3|7|他叫人通告 尼尼微 全城，說：「王和大臣有令，人、畜、牛、羊都不可嘗任何東西，不可吃，也不可喝水。
JONAH|3|8|人與牲畜都要披上麻布，切切求告上帝。各人要回轉離開惡道，離棄自己掌中的殘暴。
JONAH|3|9|誰知道上帝也許會回心轉意，不發烈怒，使我們不致滅亡。」
JONAH|3|10|上帝察看他們的行為，見他們離開惡道，上帝就改變心意，原先所說要降與他們的災難，他不降了。
JONAH|4|1|這事令 約拿 大大不悅，甚至發怒。
JONAH|4|2|他就向耶和華禱告，說：「耶和華啊，這不就是我仍在本國的時候所說的嗎？我知道你是有恩惠，有憐憫的上帝，不輕易發怒，有豐盛的慈愛，並且會改變心意，不降那災難。我就是因為這樣，才急速逃往 他施 去的呀！
JONAH|4|3|耶和華啊，現在求你取走我的性命吧！因為我死了比活著更好。」
JONAH|4|4|耶和華說：「你這樣發怒，對嗎？」
JONAH|4|5|約拿 出城，坐在城的東邊，在那裏為自己搭了一座棚。他坐在棚子的蔭下，要看看城裏會發生甚麼事。
JONAH|4|6|耶和華上帝安排了一棵蓖麻，使它生長高過 約拿 ，影子遮蓋他的頭，使他免受苦難； 約拿 因這棵蓖麻大大歡喜。
JONAH|4|7|次日黎明，上帝卻安排一條蟲來咬這蓖麻，以致枯乾。
JONAH|4|8|太陽出來的時候，上帝安排炎熱的東風，太陽曝曬 約拿 的頭，使他發昏，他就為自己求死，說：「我死了比活著更好！」
JONAH|4|9|上帝對 約拿 說：「你因這棵蓖麻這樣發怒，對嗎？」他說：「我發怒以至於死，都是對的！」
JONAH|4|10|耶和華說：「這棵蓖麻你沒有為它操勞，也不是你使它長大的；它一夜生長，一夜枯死，你尚且愛惜；
JONAH|4|11|何況這 尼尼微 大城，其中不能分辨左右手的就有十二萬多人，還有許多牲畜，我豈能不愛惜呢？」
MIC|1|1|當 猶大 王 約坦 、 亞哈斯 、 希西家 在位的時候，耶和華的話臨到 摩利沙 人 彌迦 ，他見到有關 撒瑪利亞 和 耶路撒冷 的異象。
MIC|1|2|萬民哪，你們都要聽！ 地和其上所有的，要留心聽！ 主耶和華要從他的聖殿 指證你們的不是。
MIC|1|3|看哪，耶和華從他的居所出來， 降臨步行地之高處。
MIC|1|4|眾山在他底下熔化， 諸谷崩裂， 如蠟熔在火中， 如水沖下山坡。
MIC|1|5|這都是因 雅各 的罪過， 因 以色列 家的罪惡。 雅各 的罪過在哪裏呢？ 豈不是在 撒瑪利亞 嗎？ 猶大 的丘壇在哪裏呢？ 豈不是在 耶路撒冷 嗎？
MIC|1|6|因此，我必使 撒瑪利亞 變為田野的廢墟， 用以栽植葡萄； 我必把它的石頭倒在山谷， 掀開它的地基。
MIC|1|7|城裏一切雕刻的偶像必被打碎， 行淫的賞金全被火燒， 我要毀滅它的一切偶像； 因為從妓女的賞金積聚而來的， 它們仍歸為妓女的賞金。
MIC|1|8|為此我要大聲哀號， 赤身赤腳行走； 我要呼號如野狗， 哀鳴如鴕鳥。
MIC|1|9|因為 撒瑪利亞 的創傷無法醫治， 蔓延到 猶大 ， 到了我百姓的城門， 直達 耶路撒冷 。
MIC|1|10|不要在 迦特 宣揚 這事， 千萬不要哭泣； 要在 伯‧亞弗拉 翻滾於灰塵 中。
MIC|1|11|沙斐 的居民哪，要赤身羞愧地經過， 撒南 的居民不敢出門， 伯‧以薛 哀哭，不再支持你們。
MIC|1|12|瑪律 的居民心甚憂急，切望得著福氣， 因為災禍已從耶和華那裏臨到 耶路撒冷 的城門。
MIC|1|13|拉吉 的居民哪，要用快馬 套車； 錫安 的罪由你而起， 以色列 的罪過在你那裏顯出。
MIC|1|14|因此，你要將送別禮送到 摩利設‧迦特 ； 亞革悉 的眾家族必用詭詐 待 以色列 諸王。
MIC|1|15|瑪利沙 的居民哪， 我必使搶奪者來到你這裏； 以色列 的貴族 必來到 亞杜蘭 。
MIC|1|16|猶大 啊，為了你所喜愛的兒女， 你要剪髮，剃光頭， 要使你的頭光禿，如同禿鷹， 因為他們被擄去離開你了。
MIC|2|1|禍哉，那些在床上圖謀罪孽、籌劃惡事的人！ 天一亮，他們因手中有能力就去行惡。
MIC|2|2|他們看上田地就佔據， 貪圖房屋便奪取； 他們欺壓戶主和他的家庭， 霸佔人和他的產業。
MIC|2|3|所以耶和華如此說： 看哪，我籌劃災禍降與這家族； 這災禍在你們頸項上無法解脫， 你們也不能昂首而行， 因為這是災禍的時刻。
MIC|2|4|到那日，必有人為你們唱詩歌， 用悲哀的哀歌哀號，說： 「我們全然敗落， 我百姓的產業易主了！ 耶和華竟然使它離開我， 我們的田地為悖逆的人所瓜分了！」
MIC|2|5|因此，你必無人能在耶和華的會中 抽籤拉繩 。
MIC|2|6|他們傳講說：「不可傳講； 人都不可傳講這些事， 羞辱不會臨到我們。」
MIC|2|7|雅各 家啊，可這麼說嗎 ？ 耶和華沒有耐心嗎？ 這些事是他所行的嗎？ 我的言語豈不是與行動正直的人有益嗎？
MIC|2|8|然而，近來我的百姓興起如仇敵。 你們剝去那些安然行路、不願打仗之人身上的外衣，
MIC|2|9|把我百姓中的婦人從安樂家中趕出， 又將我的榮耀從她們孩子身上永遠奪去。
MIC|2|10|起來，走吧！ 這裏並非安歇之處； 因為不潔淨帶來毀壞， 且是大大的毀壞。
MIC|2|11|若有人心存虛假，用謊言說 ： 「我向你們傳講可得清酒和烈酒 」， 那人就必作這百姓的傳講者。
MIC|2|12|雅各 家啊，我定要聚集你們， 定要召集 以色列 的餘民， 把他們安置在一處，如 波斯拉 的羊， 又如草場上的羊群， 人數眾多，大大喧嘩。
MIC|2|13|開路的在他們前面上去， 直闖過城門，從城門出去； 他們的王在前面行， 耶和華在他們的前頭。
MIC|3|1|於是我說： 雅各 的領袖， 以色列 家的官長啊， 你們要聽！ 你們豈不知道公平嗎？
MIC|3|2|你們惡善好惡， 剝我百姓 身上的皮， 從他們的骨頭上剔肉，
MIC|3|3|你們吃我百姓的肉， 剝他們的皮， 打斷他們的骨頭， 如切塊 下鍋， 如釜中的肉。
MIC|3|4|到了遭災的時候，這些人要哀求耶和華， 他卻不應允他們。 那時，因他們所行的惡， 他必轉臉離開他們。
MIC|3|5|論到使我百姓走入歧途的先知， 他們牙齒有所嚼，就呼喊說：「平安！」 誰不給他們吃，就揚言攻擊他， 耶和華如此說：
MIC|3|6|你們因此必遭遇黑夜，看不到異象； 遭遇幽暗，無法占卜。 太陽必向先知沉落， 白晝轉為黑暗。
MIC|3|7|先見必抱愧， 占卜的必蒙羞， 他們全都摀著鬍鬚， 因為上帝不應允他們。
MIC|3|8|至於我，我藉耶和華的靈， 滿有能力、公平和勇氣， 可向 雅各 述說他的過犯， 向 以色列 指出他的罪惡。
MIC|3|9|當聽這話， 雅各 家的領袖， 以色列 家的官長啊！ 你們厭棄公平， 在一切事上屈枉正直；
MIC|3|10|以血建立 錫安 ， 以罪孽建造 耶路撒冷 。
MIC|3|11|城裏的領袖為賄賂行審判， 祭司為酬勞施訓誨， 先知為銀錢行占卜； 他們卻倚賴耶和華，說： 「耶和華不是在我們中間嗎？ 災禍必不臨到我們。」
MIC|3|12|因此，為你們的緣故， 錫安 要被耕種像一塊田地， 耶路撒冷 要變為廢墟， 這殿的山必如叢林的高處。
MIC|4|1|末後的日子， 耶和華殿的山必堅立， 超乎諸山，高舉過於萬嶺； 萬民都要流歸這山。
MIC|4|2|必有許多民族前往，說： 「來吧，我們登耶和華的山， 到 雅各 上帝的殿。 他必將他的道指教我們， 我們也要行他的路。」 因為教誨必出於 錫安 ， 耶和華的言語必出於 耶路撒冷 。
MIC|4|3|他必在許多民族中施行審判， 為遠方強盛的國斷定是非。 他們要將刀打成犁頭， 把槍打成鐮刀。 這國不舉刀攻擊那國， 他們也不再學習戰事。
MIC|4|4|人人都要坐在自己的葡萄樹 和無花果樹下， 無人使他們驚嚇； 這是萬軍之耶和華親口說的。
MIC|4|5|萬民都奉自己神明的名行事， 我們卻要奉耶和華－我們上帝的名而行， 直到永永遠遠。
MIC|4|6|耶和華說：在那日， 我必聚集瘸腿的， 召集被趕逐的， 以及我所懲治的人。
MIC|4|7|我要使瘸腿的成為餘民， 使被趕到遠方的成為強盛之國。 耶和華要在 錫安山 作王治理他們， 從今直到永遠。
MIC|4|8|你， 以得臺 ， 錫安 的山岡啊， 先前的權柄必歸給你， 耶路撒冷 的國權必將歸還。
MIC|4|9|現在，你為何大聲呼喊呢？ 你中間沒有君王， 你的謀士滅絕， 以致疼痛抓住你， 如臨產的婦人嗎？
MIC|4|10|錫安 哪，你要疼痛生產， 彷彿臨產的婦人； 因你必從城裏出來，住在田野； 你要到 巴比倫 去， 在那裏，你要蒙解救， 在那裏，耶和華必救贖你 脫離仇敵的手掌。
MIC|4|11|現在，許多國家聚集攻擊你，說： 「讓 錫安 被玷污！ 讓我們親眼看到！」
MIC|4|12|他們卻不知道耶和華的意念， 也不明白他的籌算， 他聚集他們， 像把禾捆聚到禾場。
MIC|4|13|錫安 哪，起來踹穀吧！ 我必使你的角成為鐵， 使你的蹄成為銅。 你必打碎許多民族， 將他們的財寶獻給耶和華， 將他們的財富獻給全地的主。
MIC|5|1|成群的民 哪，現在要聚集成隊； 仇敵前來圍攻我們， 要用杖擊打 以色列 領袖的臉頰。
MIC|5|2|伯利恆 的 以法他 啊， 你在 猶大 諸城中雖小， 將來必有一位從你那裏出來， 在 以色列 中為我作掌權者； 他的根源自亙古，從太初就有。
MIC|5|3|因此，耶和華要將 以色列 人交給敵人， 直到臨產的婦人生下孩子； 那時，他其餘的弟兄 必回到 以色列 人那裏。
MIC|5|4|他必倚靠耶和華的大能， 倚靠耶和華－他上帝之名的威嚴， 站立並牧養， 使他們安然居住； 因為現在他必尊大， 直到地極。
MIC|5|5|這位就是和平 。 當 亞述 侵入我們領土， 踐踏我們宮殿時， 我們就立七個牧者， 八個領袖攻擊它。
MIC|5|6|他們要用刀劍毀壞 亞述 地 和 寧錄 地的關口 。 當 亞述 侵入我們領土， 踐踏我們邊境時， 他必拯救我們。
MIC|5|7|雅各 的餘民 必在許多民族中， 如從耶和華降下的露水， 又如甘霖降在草上； 他們不倚靠人， 也不仰賴世人。
MIC|5|8|雅各 的餘民必在列國中， 在許多民族中， 如林間百獸中的獅子， 又如少壯獅子在羊群中； 他若經過就必踐踏撕裂， 無人搭救。
MIC|5|9|願你的手舉起，高過敵人！ 願你的仇敵都被剪除！
MIC|5|10|耶和華說：到那日， 我必從你中間剪除馬匹， 毀壞戰車；
MIC|5|11|除滅你國中的城鎮， 拆毀你一切的堡壘；
MIC|5|12|除掉你手中的邪術， 你那裏不再有占卜的人。
MIC|5|13|我必從你中間除滅雕刻的偶像和柱像， 你就不再跪拜自己手所造的；
MIC|5|14|我必從你中間拔除 亞舍拉 ， 毀滅你的城鎮；
MIC|5|15|我必在怒氣和憤怒中 報應那不聽從我的列國。
MIC|6|1|當聽耶和華說的話： 起來，向山嶺爭辯， 使岡陵聽見你的聲音。
MIC|6|2|山嶺啊，要聽耶和華的指控！ 大地永久的根基啊，要聽！ 因耶和華控告他的百姓， 與 以色列 爭辯。
MIC|6|3|「我的百姓啊，我向你做了甚麼呢？ 我在甚麼事上使你厭煩？ 你回答我吧！
MIC|6|4|我曾將你從 埃及 地領出來， 從為奴之家救贖你， 我差遣 摩西 、 亞倫 和 米利暗 在你前面帶領。
MIC|6|5|我的百姓啊，當記念從前 摩押 王 巴勒 如何籌算， 比珥 的兒子 巴蘭 如何回應他， 當記念從 什亭 到 吉甲 所發生的事， 好使你們明白耶和華公義的作為。」
MIC|6|6|「我朝見耶和華， 在至高上帝面前跪拜，當獻上甚麼呢？ 難道獻一歲的牛犢為燔祭來朝見他嗎？
MIC|6|7|耶和華豈喜悅千千的公羊， 或是萬萬的油河嗎？ 我豈可為自己的過犯獻我的長子， 為自己的罪惡獻我所親生的嗎？」
MIC|6|8|世人哪，耶和華已指示你何為善。 他向你所要的是甚麼呢？ 只要你行公義，好憐憫， 存謙卑的心與你的上帝同行。
MIC|6|9|耶和華向這城呼叫 ─看重你的名是真智慧 ─ 你們當聽懲罰 和派定懲罰的人 。
MIC|6|10|惡人家中不是仍有不義之財 和惹人生氣的變小了的伊法嗎？
MIC|6|11|我若用不公道的天平 和袋中詭詐的法碼， 豈可算為清白呢？
MIC|6|12|城裏的有錢人遍行殘暴， 其中的居民說謊話， 口中的舌頭盡是詭詐。
MIC|6|13|因此，我也擊打你，使你受傷 ， 因你的罪惡使你受驚駭。
MIC|6|14|你要吃，卻吃不飽， 你的肚子仍是空空。 你必被挪去，不得逃脫； 如有逃脫的，我必交給刀劍。
MIC|6|15|你撒種，卻不得收割； 踹橄欖，卻不得油抹身； 有新酒，卻不得酒喝。
MIC|6|16|因為你遵守 暗利 的規條， 行 亞哈 家一切所行的， 順從他們的計謀； 因此，我必使你荒涼， 使你的居民遭人嗤笑， 你們也必擔當我百姓的羞辱。
MIC|7|1|我有禍了！我好像夏日收割後的果子， 又如收成之後剩餘的葡萄， 沒有一掛可吃的， 也沒有我心所渴想初熟的無花果。
MIC|7|2|地上的虔誠人滅盡了， 人世間已無正直的人； 他們都埋伏，為要流人的血， 用羅網獵取自己的弟兄。
MIC|7|3|他們雙手善於作惡， 君王和審判官都索取賄賂； 位高的人吐出心中的慾望， 彼此勾結 。
MIC|7|4|他們當中最好的，不過像蒺藜； 最正直的，不過如荊棘籬笆。 你守候的日子，懲罰已經來到， 他們必擾亂不安。
MIC|7|5|不可倚賴鄰舍， 不可信靠密友； 甚至對躺在你懷中的妻子 也要守住你的口。
MIC|7|6|因為兒子藐視父親， 女兒抵擋母親， 媳婦抗拒婆婆， 人的仇敵就是自己家裏的人。
MIC|7|7|至於我，我要仰望耶和華， 等候那救我的上帝； 我的上帝必應允我。
MIC|7|8|我的仇敵啊，不要向我誇耀。 我雖跌倒，仍要起來； 雖坐在黑暗裏，耶和華卻作我的光。
MIC|7|9|我要承受耶和華的惱怒， 直到他為我辯護，為我伸冤， 因我得罪了他； 他要領我進入光明， 我必得見他的公義。
MIC|7|10|那時我的仇敵看見這事就羞愧， 他曾對我說：「耶和華－你的上帝在哪裏？」 我必親眼見他遭報， 現在，他必被踐踏，如同街上的泥土。
MIC|7|11|你的城牆重修的日子到了！ 到那日，邊界必擴展。
MIC|7|12|到那日，人必從 亞述 ， 從 埃及 的城鎮， 從 埃及 到 大河 ， 從這海到那海， 從這山到那山， 都歸到你這裏。
MIC|7|13|然而，因居民的緣故， 為了他們行事的結果， 這地必然荒涼。
MIC|7|14|求你在 迦密 的樹林中， 以你的杖牧放你獨居的民， 你產業中的羊群； 願他們像古時一樣， 牧放在 巴珊 和 基列 。
MIC|7|15|我要顯奇事給他們看， 好像出 埃及 地的時候一樣。
MIC|7|16|列國看見，雖大有勢力仍覺慚愧； 他們必用手摀口，掩耳不聽。
MIC|7|17|他們要舔土如蛇， 又如地上爬行的動物， 戰戰兢兢離開他們的營寨； 他們必畏懼耶和華─我們的上帝， 也必因你而害怕。
MIC|7|18|有哪一個神明像你，赦免罪孽， 饒恕他產業中餘民的罪過？ 他不永遠懷怒，喜愛施恩。
MIC|7|19|他 必轉回憐憫我們， 把我們的罪孽踏在腳下。 你必將他們 一切的罪投於深海。
MIC|7|20|你必按古時向我們列祖起誓的話， 以信實待 雅各 ， 向 亞伯拉罕 施慈愛。
NAH|1|1|論 尼尼微 的默示， 伊勒歌斯 人 那鴻 所見異象的書。
NAH|1|2|耶和華是忌邪 、報應的上帝。 耶和華施報應，大有憤怒； 耶和華向他的敵人報應， 向他的仇敵懷怒。
NAH|1|3|耶和華不輕易發怒，大有能力， 但耶和華萬不以有罪的為無罪。 他的道路在旋風和暴風之中， 雲彩為他腳下的塵土。
NAH|1|4|他斥責海，使海枯乾， 使一切江河乾涸。 巴珊 和 迦密 衰殘， 黎巴嫩 的花草也衰殘了。
NAH|1|5|大山因他震動， 小山也都融化； 大地在他面前突起， 世界和住在其間的也都如此。
NAH|1|6|他發憤恨，誰能立得住呢？ 他發烈怒，誰能當得起呢？ 他的憤怒如火傾洩而出， 磐石因他崩裂。
NAH|1|7|耶和華本為善， 在患難的日子為人的保障， 並且認識那些投靠他的人；
NAH|1|8|但他必以漲溢的洪水淹沒其地方 ， 又驅逐仇敵進入黑暗。
NAH|1|9|你們籌劃何種計謀攻擊耶和華呢？ 他必終結一切， 仇敵 不會再度興起。
NAH|1|10|你們像雜亂的荊棘， 像喝醉了的人， 又如枯乾的碎秸，全然燒滅。
NAH|1|11|有一人從你那裏出來， 圖謀邪惡，設惡計攻擊耶和華。
NAH|1|12|耶和華如此說： 「他們雖然勢力強大，人數眾多， 也要被剪除，歸於無有。 我雖曾使你受苦， 卻不再使你受苦。
NAH|1|13|現在，我要從你身上折斷他的軛， 解開捆綁你的繩索。」
NAH|1|14|耶和華已經發命令，指著你說： 「你的名下必不再留後； 我要從你神明的廟中除滅雕刻的偶像和鑄造的偶像， 我必因你的卑賤，為你預備墳墓。」
NAH|1|15|看哪，山上有報佳音、傳平安之人的腳蹤。 猶大 啊，守你的節期， 還你的願吧！ 因為惡人不再侵犯你， 他已滅絕淨盡了。
NAH|2|1|那打碎你的人 上到你面前。 要看守堡壘，把守道路， 要挺起腰來，大大使力。
NAH|2|2|耶和華復興 雅各 的榮華， 像復興 以色列 的榮華； 因為蹂躪者曾經蹂躪他們， 毀壞了他們的葡萄枝。
NAH|2|3|他勇士的盾牌是紅的， 精兵都穿朱紅衣服。 在預備打仗的日子， 戰車上的鐵閃爍如火 ， 柏木的槍桿也已舉起 ；
NAH|2|4|戰車在街上疾行， 在廣場上來往奔馳， 形狀如火把， 飛馳如閃電。
NAH|2|5|他 招聚他的貴族； 他們前行時絆跌， 速上城牆， 預備屏障。
NAH|2|6|河閘開放， 宮殿沖沒。
NAH|2|7|這是命定之事： 王后赤身被擄 ， 宮女搥胸， 哀鳴如鴿子。
NAH|2|8|尼尼微 自古以來 如同聚水的池子； 現在居民都在逃跑 。 「站住！站住！」 卻無人回轉。
NAH|2|9|你們搶奪金子吧！ 你們搶奪銀子吧！ 因為所積蓄的無窮， 華美的寶器無數。
NAH|2|10|荒蕪，荒涼，全然荒廢， 人心害怕，雙膝顫抖， 腰部疼痛，臉都變色。
NAH|2|11|獅子的洞， 幼獅餵養之處在哪裏呢？ 公獅、母獅、小獅出入， 無人使牠們驚嚇之地在哪裏呢？
NAH|2|12|公獅撕碎的足夠給幼獅吃， 又為母獅掐死獵物， 把獵物塞滿牠的洞穴， 把撕碎的裝滿牠的窩。
NAH|2|13|看哪，我與你為敵，將它的戰車 焚燒成煙，刀劍必吞滅你的少壯獅子；我必從地上除滅你的獵物，你使者的聲音必不再聽見。這是萬軍之耶和華說的。
NAH|3|1|禍哉！這流人血的城， 欺詐連連，搶奪充斥， 擄掠的事總不止息。
NAH|3|2|鞭聲響亮，車輪轟轟， 馬匹跳躍，戰車奔騰；
NAH|3|3|騎兵爭先，刀劍發光， 槍矛閃爍，被殺的甚多， 屍首成堆，屍骸無數， 人因屍骸而絆跌，
NAH|3|4|都因那美貌的妓女多有淫行， 慣行邪術， 藉淫行誘惑 列國， 用邪術誘惑萬族。
NAH|3|5|看哪，我與你為敵， 掀開你的下襬，蒙在你臉上， 使列邦看見你的赤體， 使列國觀看你的羞辱。 這是萬軍之耶和華說的。
NAH|3|6|我必將可憎污穢之物拋在你身上， 使你被藐視，為眾人所觀看。
NAH|3|7|凡看見你的，都必逃離你，說： 「 尼尼微 荒涼了！有誰為你悲傷呢？ 我何處找到安慰你的人呢？」
NAH|3|8|你能勝過 挪亞們 嗎？ 它坐落在眾河之間， 周圍有水， 海 作它的城郭， 海 作它的城牆。
NAH|3|9|古實 和 埃及 是它的力量， 沒有窮盡， 弗 人和 路比 人是它的幫手。
NAH|3|10|但它被流放，被人擄去， 它的嬰孩也被摔碎在各街頭； 人為它的貴族抽籤， 它的權貴都被鎖鏈鎖住。
NAH|3|11|你也必喝醉，昏迷錯亂， 並因仇敵的緣故尋求庇護。
NAH|3|12|你一切的堡壘必如無花果樹上初熟的果子， 一經搖動，就落在想吃的人口中。
NAH|3|13|看哪，你中間的士兵是婦女， 你國中的關口向仇敵敞開， 你的門閂被火焚燒。
NAH|3|14|你要打水預備受困； 要加強防禦， 取土踹泥， 做成磚模。
NAH|3|15|在那裏，火要吞滅你， 刀必殺戮你， 如蝻子般吞滅你。 你人數增多如蝻子， 增多如蝗蟲吧！
NAH|3|16|你增添商賈，多過天上的星宿； 如蝻子蛻皮飛去。
NAH|3|17|你的領袖多如蝗蟲， 你的將軍彷彿成群的蝗蟲； 天涼時齊落在籬笆上， 太陽一出就飛去， 人不知道落在何處。
NAH|3|18|亞述 王啊， 你的牧人睡覺， 你的貴族躺臥 ， 你的百姓散在山間， 無人招聚。
NAH|3|19|你的損傷並未減輕， 你的傷痕極其重大。 凡聽見這消息的人都因你拍掌。 有誰沒有時常遭受你的暴行呢？
HAB|1|1|哈巴谷 先知所看見的默示。
HAB|1|2|耶和華啊，我呼求， 你不應允，要到幾時呢？ 我向你呼喊「暴力！」 你還不拯救？
HAB|1|3|你為何使我看見罪孽？ 你為何坐視奸惡呢？ 毀滅和兇暴在我面前， 爭執與紛爭不斷發生。
HAB|1|4|因此律法無效， 公理從未彰顯。 因惡人圍困義人， 所以公理遭受扭曲。
HAB|1|5|你們要向列國觀看 ，注意看， 要驚奇，再驚奇！ 因為在你們的日子，有一件事發生 ， 儘管有人說了，你們還是不信。
HAB|1|6|看哪，我必興起 迦勒底 人， 就是那殘忍暴躁之民，通行遍地， 霸佔不屬自己的住處。
HAB|1|7|他威武可畏， 審判與威權都由他而出。
HAB|1|8|他的馬比豹更快， 比晚上 的野狼更猛。 他的戰馬跳躍， 他的戰馬從遠方而來 ； 他們飛跑，如鷹急速抓食，
HAB|1|9|都為施行殘暴而來， 他們的臉面向東 ， 聚集俘虜，多如塵沙。
HAB|1|10|他譏誚列王， 嘲諷領袖， 嗤笑一切堡壘， 堆土攻取它。
HAB|1|11|那時，他如風猛然掃過， 他背叛，顯為有罪； 他以自己的力量為神明。
HAB|1|12|耶和華－我的上帝，我的聖者啊， 你不是從亙古就有嗎？ 我們必不致死。 耶和華啊，你派他為要行審判； 磐石啊，你立他為要懲治人。
HAB|1|13|你的眼目清潔， 不看邪惡，也不看奸惡， 為何你卻看著人行詭詐呢？ 惡人吞滅比自己公義的人， 為何你保持沉默呢？
HAB|1|14|你為何使人如海中的魚， 又如無人管轄的爬行動物呢？
HAB|1|15|他用鉤子把他們全拉上來， 用羅網捕獲他們， 拉漁網聚集他們。 因此，他歡喜快樂，
HAB|1|16|向羅網獻祭， 向漁網燒香； 因為他藉此得豐盛的收穫 與肥美的食物。
HAB|1|17|但他豈可因此屢屢倒空羅網 ， 時常殺戮列國的人，毫不顧惜呢？
HAB|2|1|我要站在我的瞭望臺， 立在城樓 上觀看， 看耶和華要對我說甚麼， 我可用甚麼話向他訴冤。
HAB|2|2|耶和華回答我，說： 將這默示清楚地寫在看板上， 使人容易朗讀 。
HAB|2|3|因為這默示有一定日期， 論及終局，絕不落空。 它雖然耽延，你要等候； 因為它必臨到，不再遲延。
HAB|2|4|看哪，惡人自高自大，心不正直； 惟義人必因他的信得生 。
HAB|2|5|他因酒詭詐、 狂傲、不安於位； 他張開喉嚨 ，好像陰間， 如死亡不能知足， 他聚集萬國， 招聚萬民全歸自己。
HAB|2|6|這些人豈不都要提起詩歌和俗語，嘲諷他說： 禍哉！你增添不屬自己的財物， 靠押金發財，要到幾時呢？
HAB|2|7|咬傷你的 豈不忽然興起， 擾害你的豈不突然崛起， 你就成為他們的擄物嗎？
HAB|2|8|因你搶奪許多國家， 流人的血，向土地、城鎮和全城的居民施行殘暴， 各國殘存之民都必搶奪你。
HAB|2|9|禍哉！那為本家積蓄不義之財、 在高處搭窩、指望得免災禍的人！
HAB|2|10|你圖謀剪除許多民族，犯了罪， 使自己的家蒙羞，自害己命。
HAB|2|11|牆裏的石頭要呼叫， 屋內的棟梁必應聲。
HAB|2|12|禍哉！那以鮮血建城、 以罪孽造鎮的人！
HAB|2|13|看哪，這不都是 出於萬軍之耶和華嗎？ 萬民勞碌得來的被火焚燒， 萬族辛苦建造的，歸於虛空。
HAB|2|14|全地都必認識耶和華的榮耀， 好像水充滿海洋一般。
HAB|2|15|禍哉！那給鄰舍酒喝，加上毒物 ， 使人喝醉，為要看見他們下體的人！
HAB|2|16|你滿受羞辱，不得榮耀； 你也喝吧，顯明你是未受割禮的 ！ 耶和華右手的杯必傳到你那裏， 你的榮耀就變為羞辱。
HAB|2|17|黎巴嫩 所受的殘暴必淹沒你， 野獸所遭遇的毀滅使你驚嚇 ； 因你流人的血， 向土地、城鎮和全城的居民施行殘暴。
HAB|2|18|偶像有甚麼益處呢？ 製造者雕刻它， 鑄成偶像，作虛假的教師； 製造者倚靠的是自己所做的啞巴偶像。
HAB|2|19|禍哉！那對木頭說「醒起」， 對啞巴石頭說「起來」的人！ 偶像豈能教導人呢？ 看哪，它以金銀包裹，其中並無氣息。
HAB|2|20|惟耶和華在他的聖殿中， 全地都當在他面前肅靜。
HAB|3|1|哈巴谷 先知的禱告，調用流離歌。
HAB|3|2|耶和華啊，我聽見你的名聲； 耶和華啊，我懼怕你的作為。 求你在這些年間 復興你的作為， 在這些年間將它顯明出來 ； 在發怒的時候以憐憫為念。
HAB|3|3|上帝從 提幔 而來， 聖者從 巴蘭山 臨到； 他的榮光遮蔽諸天， 頌讚遍滿全地。
HAB|3|4|他的輝煌如同日光， 從他手裏發出光芒， 那裏 隱藏他的能力。
HAB|3|5|在他前面有瘟疫流行， 在他腳下有熱症發出。
HAB|3|6|他站立，震動 大地， 他觀看，震動列國。 永久的山崩裂， 長存的嶺塌陷， 他的作為與古時一樣。
HAB|3|7|我見 古珊 的帳棚遭難， 米甸 地的幔子動搖。
HAB|3|8|耶和華啊，你豈是向江河發怒， 向江河生氣， 向海洋發烈怒嗎？ 你騎在馬上， 坐在得勝的戰車上，
HAB|3|9|你的弓全然顯露 ， 箭是發誓的言語 ； 你以江河分開大地。
HAB|3|10|山嶺見你，無不戰抖； 大水氾濫而過， 深淵發聲， 洶湧翻騰 。
HAB|3|11|因你的箭射出光芒， 你的槍閃出光耀， 日月都停在原處。
HAB|3|12|你發怒遍行大地， 以怒氣責打列國，如打穀一般。
HAB|3|13|你出來拯救你的百姓， 拯救你的受膏者； 你打破惡人之家的頭， 暴露其根基，直到頸項 。
HAB|3|14|你以其戈矛刺透他戰士的頭； 他們如旋風將我 颳散， 他們喜愛暗中吞吃困苦的人。
HAB|3|15|你騎馬踐踏海， 踐踏洶湧的大水。
HAB|3|16|我聽見這聲音，身體戰兢， 嘴唇發顫， 骨中朽爛， 在所立之處戰兢 ； 但我安靜等候 災難之日臨到那上來侵犯我們的民 。
HAB|3|17|雖然無花果樹不發旺， 葡萄樹不結果， 橄欖樹也不收成， 田地不出糧食， 圈中絕了羊， 棚內也沒有牛；
HAB|3|18|然而，我要因耶和華歡欣， 因救我的上帝喜樂。
HAB|3|19|主耶和華是我的力量， 他使我的腳快如母鹿， 又使我穩行在高處。 這歌交給聖詠團長，用絲弦的樂器。
ZEPH|1|1|當 亞們 的兒子 猶大 王 約西亞 在位的時候，耶和華的話臨到 希西家 的玄孫， 亞瑪利雅 的曾孫， 基大利 的孫子， 古示 的兒子 西番雅 。
ZEPH|1|2|耶和華說： 「我必從地面上徹底除滅萬物。
ZEPH|1|3|我必除滅人與牲畜， 除滅空中的鳥、海裏的魚、 絆腳石和惡人； 我必把人從地面上剪除， 這是耶和華說的。
ZEPH|1|4|我必伸手攻擊 猶大 和 耶路撒冷 所有的居民； 從這地方剪除剩下的 巴力 、 事奉偶像之祭司的名字與祭司；
ZEPH|1|5|還有那些在屋頂拜天上萬象的， 那些敬拜耶和華指著他起誓， 卻又指著 米勒公 起誓的；
ZEPH|1|6|並那些轉去不跟從耶和華， 不尋求耶和華，也不求問他的。」
ZEPH|1|7|在主耶和華面前要靜默無聲， 因為耶和華的日子快到了。 耶和華已經預備祭物， 將召來的人分別為聖。
ZEPH|1|8|「到了獻祭給耶和華的日子， 我要懲罰領袖和王子， 及所有穿外邦衣服的人。
ZEPH|1|9|到那日，我必懲罰所有跳過門檻， 以殘暴和詭詐塞滿主人房屋的人。
ZEPH|1|10|「當那日，從 魚門 必發出悲哀的聲音， 從第二城區發出哀號的聲音， 從山間發出破裂的大響聲。 這是耶和華說的。
ZEPH|1|11|瑪革提施 的居民哪，你們要哀號， 因為所有的商人 都滅亡了， 滿載銀子的人都被剪除。
ZEPH|1|12|那時，我必用燈巡查 耶路撒冷 ， 懲罰那些沉湎在酒渣上的人； 他們心裏說： 『耶和華必不降福，也不降禍。』
ZEPH|1|13|他們的財寶成為掠物， 房屋變為廢墟。 他們建造房屋，卻不得住在其內； 栽葡萄園，卻不得喝其中所出的酒。」
ZEPH|1|14|耶和華的大日臨近， 臨近而且甚快； 那是耶和華日子的風聲， 勇士必在那裏痛痛地哭號。
ZEPH|1|15|那日是憤怒的日子， 急難困苦的日子， 荒廢淒涼的日子， 黑暗幽冥的日子， 烏雲密佈的日子，
ZEPH|1|16|是吹角吶喊的日子， 要攻擊堅固的城， 攻擊高大的城樓。
ZEPH|1|17|我必使災禍臨到人身上， 使他們行走如同盲人， 因為他們得罪了耶和華； 他們的血必倒出如灰塵， 肉身拋棄如糞土。
ZEPH|1|18|當耶和華發怒的日子， 他們的金銀不能救自己； 耶和華妒忌的火必燒滅全地， 要向地上所有的居民施行可怕的毀滅。
ZEPH|2|1|不知羞恥的國民哪， 趁命令尚未發出， 日子流逝如糠秕， 耶和華的烈怒尚未臨到你們， 他發怒的日子未到以先， 你們應當聚集，聚集起來。
ZEPH|2|2|
ZEPH|2|3|世上遵守耶和華典章的謙卑人哪， 你們都當尋求耶和華， 尋求公義，尋求謙卑； 或許在耶和華發怒的日子得以隱藏。
ZEPH|2|4|迦薩 必遭遺棄 ， 亞實基倫 必然荒涼； 亞實突 人必在正午被趕出， 以革倫 也要連根拔除 。
ZEPH|2|5|禍哉，住沿海之地的 基利提 人！ 迦南 、 非利士 人之地啊，耶和華的話攻擊你們： 我必毀滅你，以致無人居住。
ZEPH|2|6|沿海之地要變為草場， 牧人的住處 和羊群的圈。
ZEPH|2|7|這地必為 猶大 家的餘民所得； 他們要在那裏放牧， 晚上躺臥在 亞實基倫 的房屋中； 因為耶和華－他們的上帝必眷顧他們， 使被擄的人歸回。
ZEPH|2|8|我聽見 摩押 毀謗， 亞捫 人辱罵； 他們辱罵我的百姓， 自誇自大，侵犯他們的疆土。」
ZEPH|2|9|萬軍之耶和華－ 以色列 的上帝說： 因此，我指著我的永生起誓： 摩押 必如 所多瑪 ， 亞捫 人必像 蛾摩拉 ， 都變為刺草、鹽坑、永遠荒廢之地。 我百姓中剩餘的必擄掠他們， 我國中的倖存者必得他們的地。
ZEPH|2|10|這事臨到他們是因他們的驕傲， 他們自誇自大， 辱罵萬軍之耶和華的百姓。
ZEPH|2|11|耶和華必向他們顯為可畏， 因他使地上的眾神衰微； 列國的海島各在自己的地方敬拜他。
ZEPH|2|12|你們 古實 人， 也是被我的刀所殺的。
ZEPH|2|13|耶和華要伸手攻擊北方， 毀滅 亞述 ， 使 尼尼微 荒涼， 乾旱如同曠野。
ZEPH|2|14|群畜，就是各類 的走獸必臥在其中， 鵜鶘和豪豬要宿在柱頂； 窗戶有鳴叫的聲音， 門檻毀壞 ， 他要毀壞香柏木板 。
ZEPH|2|15|這素來歡樂、安然居住的城， 心裏說：「惟有我，除我以外再沒有別的」， 現在竟然荒涼，成為野獸躺臥之處！ 凡經過的人都必搖著手嗤笑它。
ZEPH|3|1|禍哉，這欺壓的城！ 悖逆，污穢，
ZEPH|3|2|不聽從命令， 不領受訓誨， 不倚靠耶和華， 不親近它的上帝。
ZEPH|3|3|其中的領袖是咆哮的獅子， 審判官是晚上 的野狼， 不留一點到早晨。
ZEPH|3|4|它的先知是虛浮詭詐的人， 祭司褻瀆聖所，強解律法。
ZEPH|3|5|耶和華在它中間行公義， 斷不做非義的事， 每早晨顯明他的公義，無日不然； 只是不義的人不知羞恥。
ZEPH|3|6|「我已經除滅列國， 使他們的城樓荒廢。 我使他們街道荒涼， 無人經過； 他們的城鎮毀壞， 沒有人，沒有居民。
ZEPH|3|7|我說：『只要你敬畏我， 領受訓誨； 其住處就不會照我原先所定的被剪除 。』 然而，他們從早起來就在各樣事上敗壞自己。
ZEPH|3|8|「你們要等候我， 直到我興起擄掠 的日子； 因為我已定意招聚列邦，聚集列國， 將我的惱怒，我一切的烈怒，都傾倒在它們身上。 我妒忌的火必燒滅全地。 這是耶和華說的。
ZEPH|3|9|「那時，我要改變萬民， 使他們有清潔的嘴唇， 好求告耶和華的名， 同心合意事奉我。
ZEPH|3|10|那些向我祈求的， 我所分散的子民 ， 必從 古實河 的那一邊， 獻供物給我。
ZEPH|3|11|「當那日，你必不再因一切得罪我的事蒙羞， 因為那時我必從你中間除掉狂喜高傲的人， 在我的聖山上你也不再狂傲。
ZEPH|3|12|我卻要在你中間留下困苦貧寒的百姓， 他們必投靠耶和華的名。
ZEPH|3|13|以色列 的餘民必不行惡， 不說謊，口中沒有詭詐的舌頭； 他們吃喝躺臥， 無人使他們驚嚇。」
ZEPH|3|14|錫安 哪，應當歌唱！ 以色列 啊，應當歡呼！ 耶路撒冷 啊，應當滿心歡喜快樂！
ZEPH|3|15|耶和華已經免去對你的審判， 趕出你的仇敵。 以色列 的王－耶和華在你中間； 你必不再懼怕災禍。
ZEPH|3|16|當那日，必有話對 耶路撒冷 說： 「不要懼怕！ 錫安 哪，不要手軟！
ZEPH|3|17|耶和華－你的上帝在你中間 大有能力，施行拯救。 他必因你歡欣喜樂， 他在愛中靜默， 且因你而喜樂歡呼。
ZEPH|3|18|我要聚集那些因無節期而愁煩的人， 他們曾遠離你， 是你的重擔和羞辱 。
ZEPH|3|19|那時，看哪，我必對付所有苦待你的人， 拯救瘸腿的，召集被趕出的； 那些在全地受羞辱的， 我必使他們得稱讚，享名聲。
ZEPH|3|20|那時，我必領你們回來，召集你們； 我使你們被擄之人歸回的時候， 我必使你們在地上的萬民中享名聲，得稱讚； 這是耶和華說的。」
HAG|1|1|大流士 王第二年六月初一，耶和華的話藉 哈該 先知向 撒拉鐵 的兒子 猶大 省長 所羅巴伯 和 約撒答 的兒子 約書亞 大祭司傳講，說：
HAG|1|2|「萬軍之耶和華如此說，這百姓說，建造耶和華殿的時候還沒有到 。」
HAG|1|3|耶和華的話藉 哈該 先知傳講，說：
HAG|1|4|「這殿荒涼，你們自己還住天花板的房屋嗎？
HAG|1|5|現在，萬軍之耶和華如此說，你們要省察自己的行為。
HAG|1|6|你們撒的種多，收的卻少；你們吃，卻不得飽；喝，卻不得足；穿衣服，卻不得暖；領工錢的，領了工錢卻裝入有破洞的袋中。
HAG|1|7|「萬軍之耶和華如此說，你們要省察自己的行為。
HAG|1|8|你們要上山取木料，建造這殿，我就因此喜樂，且得榮耀。這是耶和華說的。
HAG|1|9|你們盼望多得，看哪，所得的卻少；你們收到家中，我就吹去。這是為甚麼呢？因為我的殿荒涼，你們各人卻只為自己的房屋奔走。這是萬軍之耶和華說的。
HAG|1|10|所以，因你們的緣故 ，天不降甘露，地也不出土產。
HAG|1|11|我命令乾旱臨到土地、山岡、五穀、新酒、新油和地上的出產，也臨到人和牲畜，以及一切人手勞碌得來的。」
HAG|1|12|那時， 撒拉鐵 的兒子 所羅巴伯 、 約撒答 的兒子 約書亞 大祭司，和所有倖存的百姓都聽從耶和華－他們上帝的話，就是 哈該 先知奉耶和華－他們上帝差遣所說的話；百姓在耶和華面前存敬畏的心。
HAG|1|13|耶和華的使者 哈該 奉耶和華差遣對百姓說：「我與你們同在。這是耶和華說的。」
HAG|1|14|耶和華激發 撒拉鐵 的兒子 猶大 省長 所羅巴伯 、 約撒答 的兒子 約書亞 大祭司，和所有倖存百姓的心，他們就來為萬軍之耶和華－他們上帝的殿做工。
HAG|1|15|這是在 大流士 王第二年六月二十四日。
HAG|2|1|七月二十一日，耶和華的話藉 哈該 先知傳講，說：
HAG|2|2|「你要曉諭 撒拉鐵 的兒子 猶大 省長 所羅巴伯 、 約撒答 的兒子 約書亞 大祭司，和所有倖存的百姓，說：
HAG|2|3|『你們中間存留的，有誰見過這殿從前的榮耀呢？現在你們看如何？在你們眼中豈不是如同無有嗎？
HAG|2|4|所羅巴伯 啊，現在，你當剛強！這是耶和華說的。 約撒答 的兒子 約書亞 大祭司啊，你當剛強！這是耶和華說的。這地的百姓啊，你們都當剛強做工，因為我與你們同在。這是萬軍之耶和華說的。
HAG|2|5|這是照著你們出 埃及 時我與你們立約的話。我的靈仍要住在你們中間，你們不必懼怕。
HAG|2|6|萬軍之耶和華如此說：過些時候，我必再一次震動天地、滄海與乾地。
HAG|2|7|我必震動萬國，萬國的珍寶都必運來 ，我就使這殿充滿榮耀。這是萬軍之耶和華說的。
HAG|2|8|銀子是我的，金子也是我的。這是萬軍之耶和華說的。
HAG|2|9|這後來的殿的榮耀必大過先前的榮耀。這是萬軍之耶和華說的。在這地方我必賜平安。這是萬軍之耶和華說的。』」
HAG|2|10|大流士 王第二年九月二十四日，耶和華的話臨到 哈該 先知，說：
HAG|2|11|「萬軍之耶和華如此說，你要向祭司請教律法，說：
HAG|2|12|『看哪，若有人用衣服的邊兜聖肉，這衣服的邊接觸了餅，或湯，或酒，或油，或別的食物，這些是否成為聖呢？』」祭司回答說：「不。」
HAG|2|13|哈該 又說：「若有人因摸屍體染了不潔淨，然後接觸任何東西，這東西就變為不潔淨嗎？」祭司回答說：「必不潔淨。」
HAG|2|14|於是 哈該 說：「耶和華說，在我面前這民如此，這國也是如此；他們手裏的各樣工作都是如此；他們在那裏所獻的都不潔淨。」
HAG|2|15|「現在，你們心裏要想一想，從今日起，耶和華的殿還沒有一塊石頭放在石頭上的情況。
HAG|2|16|那時你們怎麼了？ 有人來到二十斗的穀堆那裏，卻只得了十斗；有人來到酒池那裏要取五十桶，卻只得了二十桶。
HAG|2|17|我以焚風 、霉爛、冰雹攻擊你們，和你們手上的各樣工作，你們仍不歸向我。這是耶和華說的。
HAG|2|18|你們心裏要想一想，從今日起，就是從這九月二十四日起，從立耶和華殿根基的日子起，你們心裏想一想：
HAG|2|19|倉裏還有穀種嗎？葡萄樹、無花果樹、石榴樹、橄欖樹雖沒有結果子， 從今日起，我必賜福。」
HAG|2|20|這月二十四日，耶和華的話再次臨到 哈該 ，說：
HAG|2|21|「你要告訴 猶大 省長 所羅巴伯 說，我必震動天地，
HAG|2|22|傾覆列國的寶座，除滅列邦列國的勢力，並傾覆戰車和坐在其上的。馬和騎兵都必跌倒，各人被弟兄的刀所殺。
HAG|2|23|萬軍之耶和華說： 撒拉鐵 的兒子我僕人 所羅巴伯 啊，這是耶和華說的，到那日，我必以你為印，因我揀選了你。這是萬軍之耶和華說的。」
ZECH|1|1|大流士 王第二年八月，耶和華的話臨到 易多 的孫子， 比利家 的兒子 撒迦利亞 先知，說：
ZECH|1|2|「耶和華曾向你們祖先大發烈怒。
ZECH|1|3|你要對 以色列 人說，萬軍之耶和華如此說：你們要轉向我，這是萬軍之耶和華說的，我就轉向你們，這是萬軍之耶和華說的。
ZECH|1|4|不要效法你們的祖先。從前的先知呼叫他們說：『萬軍之耶和華如此說，當回轉離開你們的惡道惡行。』他們卻不聽，也不順從我。這是耶和華說的。
ZECH|1|5|你們的祖先在哪裏呢？那些先知能永遠存活嗎？
ZECH|1|6|然而我的言語和律例，就是我所吩咐我僕人眾先知的，豈不臨到你們的祖先嗎？他們就回轉，說：萬軍之耶和華定意按我們的所作所為對待我們，他也已經照樣行了。」
ZECH|1|7|大流士 第二年十一月，就是細罷特月二十四日，耶和華的話臨到 易多 的孫子， 比利家 的兒子 撒迦利亞 先知，說：
ZECH|1|8|「我夜間觀看，看哪，有一人騎著紅馬，站在窪地的番石榴樹中間。在他身後有紅色、褐色和白色的馬。」
ZECH|1|9|我說：「主啊，這是甚麼意思？」與我說話的天使說：「我要指示你這是甚麼意思。」
ZECH|1|10|那站在番石榴樹中間的人回答說：「這是奉耶和華差遣，在遍地巡邏的。」
ZECH|1|11|他們對站在番石榴樹中間耶和華的使者說：「我們在遍地巡邏，看哪，全地都安息平靜。」
ZECH|1|12|於是，耶和華的使者說：「萬軍之耶和華啊，你惱恨 耶路撒冷 和 猶大 的城鎮已經七十年了，你不施憐憫要到幾時呢？」
ZECH|1|13|耶和華就用美善的話和安慰的話回答那與我說話的天使。
ZECH|1|14|與我說話的天使對我說：「你要宣告，萬軍之耶和華如此說：我為 耶路撒冷 而妒忌，為 錫安 大大妒忌。
ZECH|1|15|我非常惱怒那享安逸的列國，因我從前稍微惱怒，他們就越發加害。
ZECH|1|16|所以耶和華如此說：現在我回到 耶路撒冷 ，仍要施憐憫，我的殿要重建在其中，準繩必拉在 耶路撒冷 之上。這是萬軍之耶和華說的。
ZECH|1|17|你要再宣告，萬軍之耶和華如此說：我的城鎮要再度繁榮發達。耶和華必再安慰 錫安 ，揀選 耶路撒冷 。」
ZECH|1|18|我舉目觀看，看哪，有四隻角。
ZECH|1|19|我問那與我說話的天使：「這是甚麼意思？」他對我說：「這是擊散 猶大 、 以色列 和 耶路撒冷 的角。」
ZECH|1|20|耶和華又把四個匠人指給我看。
ZECH|1|21|我問：「這些人來做甚麼呢？」他說：「那是擊散 猶大 的角，使人不敢抬頭；但這些匠人前來威嚇列國，打掉列國的角，因為他們舉起角來擊散 猶大 地。」
ZECH|2|1|我舉目觀看，看哪，有一人手拿丈量的繩。
ZECH|2|2|我問：「你到哪裏去？」他對我說：「要去丈量 耶路撒冷 ，看有多寬多長。」
ZECH|2|3|看哪，與我說話的天使出去 ，另有一位天使迎著他來，
ZECH|2|4|對他說：「你跑去告訴這個年輕人說， 耶路撒冷 必有人居住，如同無城牆的鄉村，因為其中的人和牲畜很多。
ZECH|2|5|耶和華說：『我要作 耶路撒冷 四圍火的城牆，並要作城中的榮耀。』」
ZECH|2|6|耶和華說：「來，來！你們要從北方之地逃回；因我曾把你們分散到天的四方 。這是耶和華說的。」
ZECH|2|7|來！住 巴比倫 的 錫安 百姓啊，逃吧！
ZECH|2|8|萬軍之耶和華在顯出榮耀之後，差遣我到擄掠你們的列國那裏，他如此說：「碰你們的就是碰他自己 眼中的瞳人。
ZECH|2|9|看哪，我要揮手攻擊他們，他們就必作自己奴僕的擄物。」你們就知道萬軍之耶和華差遣了我。
ZECH|2|10|耶和華說：「 錫安 哪，應當歡樂歌唱，因為，看哪，我要來，要住在你中間。
ZECH|2|11|在那日，必有許多國家歸附耶和華，作我的子民。我要住 在你中間。」你就知道萬軍之耶和華差遣我到你那裏去。
ZECH|2|12|耶和華必收回 猶大 ，作為他聖地的產業，他必再度揀選 耶路撒冷 。
ZECH|2|13|凡血肉之軀都當在耶和華面前靜默無聲，因為他從他的聖所奮起了。
ZECH|3|1|天使 指給我看： 約書亞 大祭司站在耶和華的使者面前，撒但站在 約書亞 的右邊控告他。
ZECH|3|2|耶和華向撒但說：「撒但哪，耶和華責備你！揀選 耶路撒冷 的耶和華責備你！這不是從火中抽出來的一根柴嗎？」
ZECH|3|3|約書亞 穿著污穢的衣服，站在那使者面前。
ZECH|3|4|使者吩咐那些侍立在他面前的說：「脫去他污穢的衣服。」又對 約書亞 說：「你看，我使你的罪孽離開你，要給你穿上華美的衣服。」
ZECH|3|5|我說 ：「要將潔淨的冠冕戴在他頭上。」他們就把潔淨的冠冕戴在他頭上，給他穿上華美的衣服，耶和華的使者在旁邊站立。
ZECH|3|6|耶和華的使者告誡 約書亞 說，
ZECH|3|7|萬軍之耶和華如此說：「你若遵行我的道，謹守我的命令，就可以管理我的家，看守我的院宇；我也要使你在這些侍立的人中間來往。
ZECH|3|8|約書亞 大祭司啊，你和坐在你面前的同伴都當聽，因為他們是作預兆的：看哪，我必使我僕人 大衛 的苗裔 長出。
ZECH|3|9|看哪，這是我在 約書亞 面前所立的石頭，這一塊石頭上有七眼。看哪，我要親自雕刻這石頭，並在一日之間除掉這地的罪孽。這是萬軍之耶和華說的。
ZECH|3|10|在那日，你們各人要請鄰舍坐在葡萄樹和無花果樹下。這是萬軍之耶和華說的。」
ZECH|4|1|那與我說話的天使又來叫醒我，好像人睡覺時被喚醒一樣。
ZECH|4|2|他問我：「你看見甚麼？」我說：「我看見了，看哪，有一個純金的燈臺，頂上有燈座，其上有七盞燈，每盞燈的上頭有七根管子；
ZECH|4|3|旁邊有兩棵橄欖樹，一棵在燈座的右邊，一棵在燈座的左邊。」
ZECH|4|4|我問與我說話的天使說：「主啊，這是甚麼意思？」
ZECH|4|5|與我說話的天使回答，對我說：「你不知道這是甚麼意思嗎？」我說：「主啊，我不知道。」
ZECH|4|6|他回答我說：「這是耶和華指示 所羅巴伯 的話。萬軍之耶和華說：不是倚靠勢力，不是倚靠才能，乃是倚靠我的靈方能成事 。
ZECH|4|7|大山哪，你算甚麼呢？在 所羅巴伯 面前，你必夷為平地。他安放頂上的那塊石頭，人就歡呼：『願恩惠、恩惠歸與這殿！』」
ZECH|4|8|耶和華的話臨到我，說：
ZECH|4|9|「 所羅巴伯 的手立了這殿的根基，他的手也必完成這工，你就知道萬軍之耶和華差遣我到你們這裏。
ZECH|4|10|誰藐視這日的事為小呢？他們見 所羅巴伯 手拿石垂線就歡喜。這七盞燈 是耶和華的眼睛，遍察全地。」
ZECH|4|11|我問天使說：「那麼在燈臺左右的這兩棵橄欖樹是甚麼意思呢？」
ZECH|4|12|我再次問他：「這兩根橄欖樹枝在兩根流出金色油的金嘴旁邊，是甚麼意思呢？」
ZECH|4|13|他對我說：「你不知道這是甚麼意思嗎？」我說：「主啊，我不知道。」
ZECH|4|14|他說：「這是兩位受膏者，侍立在全地之主的旁邊。」
ZECH|5|1|我又舉目觀看，看哪，有一飛行的書卷。
ZECH|5|2|他問我：「你看見甚麼？」我回答：「我看見一飛行的書卷，長二十肘，寬十肘。」
ZECH|5|3|他對我說：「這就是向全地面發出的詛咒。凡偷竊的必按書卷這面的話除滅，凡起假誓的必按書卷那面的話除滅。
ZECH|5|4|萬軍之耶和華說：我要把這書卷送出去，進入偷竊者的家和指著我名起假誓者的家，停留在他家裏，連房屋帶木頭和石頭都毀滅了。」
ZECH|5|5|與我說話的天使前來，對我說：「你要舉目觀看，看那出現的是甚麼。」
ZECH|5|6|我問：「這是甚麼呢？」他說：「這出現的是量器 。」又說：「是他們的眼目，遍行全地 。」
ZECH|5|7|看哪，圓形的鉛蓋被抬起來，有一個婦人坐在量器中。
ZECH|5|8|天使說：「這是罪惡。」他就把婦人推進量器裏，把鉛蓋壓在量器的口上。
ZECH|5|9|於是我舉目觀看，看哪，有兩個婦人前來，她們的翅膀中有風，翅膀如同鸛鳥的翅膀。她們把量器抬起來，懸在天地之間。
ZECH|5|10|我問那與我說話的天使：「她們要把量器抬到哪裏去呢？」
ZECH|5|11|他對我說：「要抬到 示拿 地去，為它建造房屋；等預備妥當，就把它安放在自己的臺座上。」
ZECH|6|1|我又舉目觀看，看哪，有四輛馬車從兩座山的中間出來；那兩座山是銅山。
ZECH|6|2|第一輛車套著紅馬，第二輛車套著黑馬，
ZECH|6|3|第三輛車套著白馬，第四輛車套著帶斑點的馬，都是強壯的 。
ZECH|6|4|我就回應與我說話的天使說：「主啊，這是甚麼意思？」
ZECH|6|5|天使回答，對我說：「這是天的四風，是從全地之主面前出來的。」
ZECH|6|6|套著黑馬的車往北方之地去，白馬跟隨在後；有斑點的馬往南方之地去；
ZECH|6|7|那些壯馬出來，急著要在地上巡邏。天使說：「你們只管在地上巡邏。」牠們就在地上巡邏。
ZECH|6|8|他又呼叫我，告訴我說：「你看，往北方地去的已在北方之地使我放心。」
ZECH|6|9|耶和華的話臨到我，說：
ZECH|6|10|「你要拿從 巴比倫 歸來的被擄之人 黑玳 、 多比雅 、 耶大雅 所獻的，當日就要進到 西番雅 的兒子 約西亞 的家裏，
ZECH|6|11|拿這金銀做冠冕，戴在 約撒答 的兒子 約書亞 大祭司的頭上；
ZECH|6|12|對他說，萬軍之耶和華如此說：『看哪，那名稱為 大衛 苗裔的，要在本處生長，並要建造耶和華的殿。
ZECH|6|13|就是他，要建造耶和華的殿，他要承受尊榮，坐在位上掌王權；又有一位祭司坐在自己的位上，兩職之間籌劃和平。
ZECH|6|14|這冠冕要歸 希連 、 多比雅 、 耶大雅 ，和 西番雅 的兒子 賢 ，放在耶和華的殿裏作為紀念。』」
ZECH|6|15|遠方的人要來建造耶和華的殿，你們因此就知道，萬軍之耶和華差遣我到你們這裏來。你們若留意聽從耶和華－你們上帝的話，這事必然成就。
ZECH|7|1|大流士 王第四年九月，就是基斯流月初四，耶和華的話臨到 撒迦利亞 。
ZECH|7|2|那時 伯特利 人已經差遣 沙利色 和 利堅‧米勒 ，並他們的人，去懇求耶和華的恩，
ZECH|7|3|問萬軍之耶和華殿中的祭司，又問先知：「我當如歷年以來所行，在五月哭泣齋戒嗎？」
ZECH|7|4|萬軍之耶和華的話臨到我，說：
ZECH|7|5|「你要向這地全體百姓和祭司說：『你們這七十年來，在五月、七月禁食悲哀，豈是真的向我禁食嗎？
ZECH|7|6|你們吃喝，不是為自己吃，為自己喝嗎？
ZECH|7|7|當 耶路撒冷 和四圍的城鎮有人居住，享繁榮， 尼革夫 和 謝非拉 也有人居住的時候，耶和華藉從前的先知所宣告的，你們不當聽嗎？』」
ZECH|7|8|耶和華的話臨到 撒迦利亞 ，說：
ZECH|7|9|「萬軍之耶和華如此說：你們要按真正的公平來審判，彼此以慈愛憐憫相待。
ZECH|7|10|不可欺壓寡婦、孤兒、寄居的和困苦的人。誰都不可心裏謀害弟兄。
ZECH|7|11|他們卻不留意；聳肩悖逆，耳朵發沉，不肯聽從。
ZECH|7|12|他們的心堅硬如金剛石，不聽律法和萬軍之耶和華藉著他的靈差遣從前先知所說的話。因此，萬軍之耶和華大發烈怒。
ZECH|7|13|萬軍之耶和華說：我曾呼喚他們，他們不聽；將來他們呼求我，我也不聽！
ZECH|7|14|我必以旋風將他們吹散到素不認識的萬國中。他們離開以後，地就荒涼，無人來往經過；他們使美好之地荒涼了。」
ZECH|8|1|萬軍之耶和華的話臨到我，說：
ZECH|8|2|「萬軍之耶和華如此說：我為 錫安 而妒忌，大大妒忌；我為了它妒忌而大發烈怒。
ZECH|8|3|耶和華如此說：我要回到 錫安 ，住在 耶路撒冷 中間。 耶路撒冷 必稱為忠實的城，萬軍之耶和華的山必稱為聖山。
ZECH|8|4|萬軍之耶和華如此說：將來必有年老的男女坐在 耶路撒冷 的廣場上，各人因年紀老邁而手拿枴杖。
ZECH|8|5|城裏的廣場滿有男孩女孩在玩耍。
ZECH|8|6|萬軍之耶和華如此說：在那些日子，即使這事在這餘民眼中看為奇妙，難道在我眼中也看為奇妙嗎？這是萬軍之耶和華說的。
ZECH|8|7|萬軍之耶和華如此說：看哪，我要從日出之地、從日落之地拯救我的子民。
ZECH|8|8|我要領他們來，使他們住在 耶路撒冷 中間。他們要作我的子民，我要作他們的上帝，都憑信實和公義。
ZECH|8|9|「萬軍之耶和華如此說：你們的手要堅強；這些日子，你們已聽見先知的口，在萬軍之耶和華殿的根基立定、聖殿建造的日子所說的這些話。
ZECH|8|10|那些日子以前，人得不著工價，牲畜也無人雇用；且因敵人的緣故，出入不得平安；因我使人與人互相攻擊。
ZECH|8|11|但如今，我對這餘民必不像先前的日子。這是萬軍之耶和華說的。
ZECH|8|12|因為他們要平安撒種，葡萄樹要結果子，土地必有出產，天也必降甘露。我要使這餘民享受這一切。
ZECH|8|13|猶大 家和 以色列 家啊，你們從前在列國中怎樣成為可詛咒的；照樣，我要拯救你們，使你們得福 。不要懼怕，你們的手要堅強。
ZECH|8|14|「萬軍之耶和華如此說：你們祖先惹我發怒的時候，我怎樣定意降禍，並不改變；萬軍之耶和華說，
ZECH|8|15|這些日子我也定意施恩給 耶路撒冷 和 猶大 家；你們不要懼怕。
ZECH|8|16|你們所當行的是這樣：每個人要與鄰舍說誠實話，在城門口要按真正的公平來審判，使人和睦。
ZECH|8|17|誰都不可心裏謀害鄰舍，也不可喜愛起假誓，因為這些事都為我所恨惡。這是耶和華說的。」
ZECH|8|18|萬軍之耶和華的話臨到我，說：
ZECH|8|19|「萬軍之耶和華如此說：四月的禁食、五月的禁食、七月的禁食和十月的禁食，必成為 猶大 家的歡喜和快樂，以及美好的節期；所以你們要喜愛誠實與和平。
ZECH|8|20|「萬軍之耶和華如此說：將來還有眾百姓和許多城鎮的居民要來。
ZECH|8|21|這城的居民必到那城，說：『我們快去懇求耶和華的恩，尋求萬軍之耶和華；我自己也要去。』
ZECH|8|22|必有許多民族和強盛的國家來到 耶路撒冷 尋求萬軍之耶和華，懇求耶和華的恩。
ZECH|8|23|萬軍之耶和華如此說：在那些日子，列國中說各種語言的人，必有十個人強拉住一個 猶大 人衣服的邊，說：『我們要與你們同去，因為我們聽見上帝與你們同在了。』」
ZECH|9|1|耶和華的默示， 他的話臨到 哈得拉 地、 大馬士革 －因世人和 以色列 各支派的眼目都向著耶和華－
ZECH|9|2|和鄰近的 哈馬 ， 以及 推羅 和 西頓 。 因為它極有智慧，
ZECH|9|3|推羅 為自己建造堅固城 ， 堆起銀子如塵沙， 純金如街上的泥土。
ZECH|9|4|看哪，主必趕出它， 重創它海上的勢力， 它必被火吞滅。
ZECH|9|5|亞實基倫 看見必懼怕， 迦薩 看見甚痛苦， 以革倫 因失了盼望而蒙羞； 迦薩 必不再有君王， 亞實基倫 也不再有人居住，
ZECH|9|6|混血的人要住在 亞實突 ； 我必除滅 非利士 人的驕傲。
ZECH|9|7|我要除去他口中帶血之肉 和牙齒內可憎之物。 他必作餘民歸於我們的上帝， 在 猶大 像族長一樣； 以革倫 必如 耶布斯 人。
ZECH|9|8|我要紮營在我的家， 敵軍不得任意往來， 暴虐的人也不再經過， 因為我親眼看顧。
ZECH|9|9|錫安 哪，應當大大喜樂； 耶路撒冷 啊，應當歡呼。 看哪，你的王來到你這裏！ 他是公義的，並且施行拯救， 謙和地騎著驢， 騎著小驢，驢的駒子。
ZECH|9|10|我必除滅 以法蓮 的戰車 和 耶路撒冷 的戰馬； 戰爭的弓也必剪除。 他要向列國講和平； 他的權柄必從這海管到那海， 從 大河 管到地極。
ZECH|9|11|錫安 哪，我因與你立約的血， 要從無水坑裏釋放你中間被囚的人。
ZECH|9|12|被囚而有指望的人哪，要轉回堡壘； 我今日宣告，我必加倍補償你。
ZECH|9|13|我為自己把 猶大 彎緊， 我使 以法蓮 如滿弓。 錫安 哪，我要喚起你的兒女， 希臘 啊，我要攻擊你的兒女， 使你如勇士的刀。
ZECH|9|14|耶和華要顯現在他們身上， 他的箭要射出如閃電。 主耶和華必吹角， 乘南方的旋風而行。
ZECH|9|15|萬軍之耶和華必保護他們； 他們要吞滅，要踐踏彈弓的石頭 ； 他們吶喊，狂飲 如喝酒， 如盛滿的碗， 又如壇的四角。
ZECH|9|16|當那日，耶和華－他們的上帝 必看他的百姓如羊群，拯救他們； 因為他們如冠冕上的寶石， 在他的地上如旗幟高舉 。
ZECH|9|17|他是何等善！ 他是何其美！ 五穀使少男強壯， 新酒使少女健美。
ZECH|10|1|春雨的季節，你們要向耶和華求雨。 耶和華發出雷電， 為眾人降下大雨， 把田園的菜蔬賜給人。
ZECH|10|2|因為家中神像所言的是虛空， 占卜者所見的是虛假， 他們講說假夢， 徒然安慰人。 所以眾人如羊流離， 因無牧人就受欺壓。
ZECH|10|3|我的怒氣向牧人發作， 我必懲罰那為首的 ； 萬軍之耶和華眷顧他的羊群， 就是 猶大 家， 必使他們如戰場上的駿馬。
ZECH|10|4|房角石從他而出， 橛子從他而出， 戰爭的弓也從他而出， 每一個掌權的都從他而出。
ZECH|10|5|他們必如戰場上的勇士， 踐踏仇敵如街上的泥土。 他們必爭戰，因為耶和華與他們同在， 他們必使騎馬的羞愧。
ZECH|10|6|我要堅固 猶大 家， 拯救 約瑟 家， 我要領他們歸回，因我憐憫他們， 他們必像我未曾棄絕他們一樣； 都因我是耶和華－他們的上帝， 我必應允他們。
ZECH|10|7|以法蓮 人必如勇士， 他們心中暢快如同喝酒； 他們的兒女看見就歡喜， 他們的心必因耶和華喜樂。
ZECH|10|8|我要呼叫，聚集他們， 因我已經救贖他們。 他們的人數必增添， 如從前增添一樣。
ZECH|10|9|我要將他們分散在列國中， 他們必在遠方記得我； 他們與兒女都必存活， 他們要歸回。
ZECH|10|10|我必使他們從 埃及 地歸回， 從 亞述 召集他們， 領他們到 基列 地和 黎巴嫩 ； 這些還不夠他們居住。
ZECH|10|11|耶和華 必經過苦海，擊打海浪。 尼羅河 的深處全都枯乾， 亞述 的驕傲必降卑， 埃及 的權杖必除去。
ZECH|10|12|我要使他們倚靠耶和華，得以堅固， 他們必奉他的名而行 ； 這是耶和華說的。
ZECH|11|1|黎巴嫩 哪，敞開你的門， 任火吞滅你的香柏樹。
ZECH|11|2|哀號吧，松樹！ 因為香柏樹傾倒了，高大的樹毀壞了。 哀號吧， 巴珊 的橡樹！ 因為茂盛的樹林倒下來了。
ZECH|11|3|聽啊，有牧人在哀號， 因他們的榮華敗落了； 聽啊，有少壯獅子咆哮， 因 約旦河 旁的叢林荒廢了。
ZECH|11|4|耶和華－我的上帝如此說：「你要牧養這群將宰的羊。
ZECH|11|5|買羊的宰了他們，卻不認為自己有罪；賣他們的也說：『耶和華是應當稱頌的，因我富足了。』牧養他們的並不憐憫他們。
ZECH|11|6|我不再憐憫這地的居民。看哪，我要將這些人交在各人的鄰舍和君王手中；他們必毀滅這地，我卻不救任何一個脫離他們的手。這是耶和華說的。」
ZECH|11|7|於是，我牧養這群將宰的羊，就是羊群中最困苦的 ；我拿著兩根杖，一根我稱為「恩惠」 ，一根稱為「聯合」。這樣，我就牧養這群羊。
ZECH|11|8|一個月之內，我廢除了三個牧人，因為我的心厭煩他們，他們的心也憎惡我。
ZECH|11|9|我就說：「我不牧養你們。要死的，由他死；滅亡的，由他滅亡；剩餘的，由他們彼此吞食。」
ZECH|11|10|我拿起那根稱為「恩惠」的杖，折斷它，表明我廢棄與萬民所立的約。
ZECH|11|11|當日約就廢了。因此，那些羊群中最困苦的 ，看著我，就知道這真是耶和華的話。
ZECH|11|12|我對他們說：「你們若看為美，就給我工價。不然，就罷了！」於是他們秤了三十塊銀錢作為我的工價。
ZECH|11|13|耶和華對我說：「把它丟給窯戶。那是他們對我所估定的好價錢！」我就取這三十塊銀錢，在耶和華的殿中將它丟給窯戶。
ZECH|11|14|我又折斷第二根杖，就是稱為「聯合」的那根杖，表明我廢棄 猶大 與 以色列 弟兄間的情誼。
ZECH|11|15|耶和華對我說：「你再把愚昧牧人所用的器具拿來，
ZECH|11|16|因為，看哪，我要在這地立一個牧人；他不看顧將亡的，不尋找分散的，不醫治受傷的，也不牧養強壯的；卻要吞吃肥羊的肉，撕裂牠們的蹄。
ZECH|11|17|禍哉！無用的牧人丟棄羊群， 刀必臨到他的膀臂和右眼上； 他的膀臂必全然枯乾， 他的右眼也必昏暗失明。」
ZECH|12|1|耶和華的默示，他的話論到 以色列 。 鋪張諸天、建立地基、造人裏面之靈的耶和華說：
ZECH|12|2|「看哪，我要使 耶路撒冷 成為令四圍列國百姓昏醉的杯； 耶路撒冷 被圍困， 猶大 也一樣受困 。
ZECH|12|3|在那日，我要使 耶路撒冷 成為萬民的一塊沉重石頭，凡舉起它的必受重傷；地上的萬國都聚集攻擊它。
ZECH|12|4|到那日，我必令一切的馬匹驚惶，使騎馬的癲狂。我必張開眼睛看顧 猶大 家，卻使列國一切的馬匹瞎眼。這是耶和華說的。
ZECH|12|5|猶大 的族長心裏要說：『 耶路撒冷 的居民因倚靠萬軍之耶和華－他們的上帝，就成為我的力量 。』
ZECH|12|6|「那日，我必使 猶大 的族長如柴堆中的火盆，又如禾捆裏的火把；他們必左右吞滅四圍列國的百姓。 耶路撒冷 卻仍屹立在本處，仍在 耶路撒冷 ！
ZECH|12|7|「耶和華要先拯救 猶大 的帳棚，免得 大衛 家的榮耀和 耶路撒冷 居民的榮耀勝過 猶大 。
ZECH|12|8|那日，耶和華必保護 耶路撒冷 的居民。他們中間軟弱的在那日必如 大衛 ； 大衛 家必如上帝，如行在他們前面的耶和華的使者。
ZECH|12|9|那日，我必定意滅絕前來攻擊 耶路撒冷 的萬國。」
ZECH|12|10|「我要將那施恩與懇求的靈，澆灌 大衛 家和 耶路撒冷 的居民。他們必仰望我，就是他們所扎的那位。他們必為他悲傷，如喪獨子，又為他哀哭，如喪長子。
ZECH|12|11|那日，在 耶路撒冷 必有大大的哀號，如 米吉多 平原上 哈達‧臨門 的哀號。
ZECH|12|12|這地必哀哭：一家一家地哭， 大衛 家的家族聚在一處，他們的婦女聚在一處； 拿單 家的家族聚在一處，他們的婦女聚在一處。
ZECH|12|13|利未 家的家族聚在一處，他們的婦女聚在一處； 示每 家的家族聚在一處，他們的婦女聚在一處。
ZECH|12|14|其餘的各家，每一家的家族聚在一處，他們的婦女聚在一處。」
ZECH|13|1|「在那日，因罪惡與污穢的緣故，必有一泉源為 大衛 家和 耶路撒冷 的居民而開。」
ZECH|13|2|萬軍之耶和華說：「在那日，我要從地上除滅偶像的名，使它不再被記得；我也必使這地不再有先知，不再有污穢的靈。
ZECH|13|3|若還有人說預言，生他的父母必對他說：『你不得存活，因為你假借耶和華的名說謊話。』生他的父母在他說預言時，要將他刺死。
ZECH|13|4|那日，凡作先知說預言的必因所論的異象羞愧，不再穿毛皮外袍哄騙人。
ZECH|13|5|他要說：『我不是先知，我是耕地的；我從幼年就作人的奴僕。』
ZECH|13|6|有人對他說：『你兩手臂間是甚麼傷呢？』他說：『這是我在親友家中所受的傷。』」
ZECH|13|7|萬軍之耶和華說： 刀劍哪，興起攻擊我的牧人， 攻擊我的同伴吧！ 要擊打牧人，羊就分散了； 我必反手攻擊那微小的。
ZECH|13|8|這全地的人， 三分之二將被剪除而死， 三分之一仍必存留。 這是耶和華說的。
ZECH|13|9|我要使這三分之一經過火， 熬煉他們，如熬煉銀子； 試煉他們，如試煉金子。 他們要求告我的名， 我必應允他們。 我說：「這是我的子民。」 他們要說：「耶和華是我的上帝。」
ZECH|14|1|看哪，耶和華的日子臨近了，你的財物必被搶掠，在你中間被瓜分。
ZECH|14|2|我要招聚萬國與 耶路撒冷 爭戰；城必被攻取，房屋被搶奪，婦女被玷污，城中的一半被擄去；但其餘的百姓不會從城中被剪除。
ZECH|14|3|那時，耶和華要出去與那些國家打仗，如同從前戰爭的日子打仗一樣。
ZECH|14|4|那日，他的腳必站在 橄欖山 上，這山面向 耶路撒冷 的東邊。 橄欖山 必從中間裂開，自東至西成為極大的谷；山的一半向北挪移，一半向南挪移。
ZECH|14|5|你們要從我的山谷中逃跑，因為山谷必延到 亞薩 。你們要逃跑，如在 猶大 王 烏西雅 年間逃避大地震一樣 。耶和華－我的上帝必降臨，所有的聖者與你 同來。
ZECH|14|6|在那日，必沒有光，不會放晴，只有烏雲 。
ZECH|14|7|耶和華所知道的那一日，沒有白天，沒有黑夜，到了晚上仍有亮光。
ZECH|14|8|在那日，必有活水從 耶路撒冷 出來，一半往東海流，一半往西海流；冬夏都是如此。
ZECH|14|9|耶和華要作全地的王。那日，耶和華必為獨一無二，他的名也是獨一無二。
ZECH|14|10|從 迦巴 直到 耶路撒冷 南方的 臨門 ，全地要變為曠野。 耶路撒冷 要矗立於本處，從 便雅憫門 到 舊門 ，又到 角門 ，並從 哈楠業樓 ，直到王的酒池。
ZECH|14|11|人要住在其中，不再有詛咒； 耶路撒冷 必安然屹立。
ZECH|14|12|這是耶和華所降的災殃，要攻擊那些與 耶路撒冷 作戰的萬民；他們兩腳站立時，肉要潰爛，眼在眶中潰爛，舌在口中也潰爛。
ZECH|14|13|那日，耶和華必使他們大大混亂。他們彼此用手揪住，用手互相攻擊。
ZECH|14|14|猶大 也要在 耶路撒冷 打仗 。那時四圍各國的財物，就是許許多多的金銀和衣服，必被收聚。
ZECH|14|15|馬匹、騾子、駱駝、驢和營中一切的牲畜所遭的災殃與那災殃一樣。
ZECH|14|16|上來攻擊 耶路撒冷 的列國中所有剩下的人，要年年上來敬拜大君王－萬軍之耶和華，並守住棚節。
ZECH|14|17|地上萬族中，凡不上 耶路撒冷 敬拜大君王－萬軍之耶和華的，雨必不降在他們的地上。
ZECH|14|18|埃及 族若不上來，雨必不降在他們的地上；凡不上來守住棚節的列國，耶和華必用這災攻擊他們。
ZECH|14|19|這就是 埃及 的懲罰和那些不上來守住棚節之列國的懲罰。
ZECH|14|20|在那日，馬的鈴鐺上要刻上「歸耶和華為聖」。耶和華殿內的鍋必如祭壇前的碗一樣。
ZECH|14|21|耶路撒冷 和 猶大 一切的鍋都必歸萬軍之耶和華為聖。凡獻祭的都必來取這鍋，在其中煮肉。當那日，在萬軍之耶和華的殿中必不再有做買賣的人 。
MAL|1|1|耶和華的話，藉 瑪拉基 傳給 以色列 的默示。
MAL|1|2|耶和華說：「我曾愛你們。」你們卻說：「你在何事上愛我們呢？」耶和華說：「 以掃 不是 雅各 的哥哥嗎？我卻愛 雅各 ，
MAL|1|3|惡 以掃 ，使他的山嶺荒涼，把他的地業交給曠野的野狗。」
MAL|1|4|以東 若說：「我們雖被毀壞，卻要重建荒廢之處。」萬軍之耶和華如此說：「任他們建造，我必拆毀；人必稱他們為『邪惡之境』，為『耶和華永遠惱怒之民』。」
MAL|1|5|你們必親眼看見，你們要說：「耶和華在 以色列 疆界之外必尊為大！」
MAL|1|6|萬軍之耶和華對你們說：「兒子孝敬父親，僕人敬畏主人；我既為父親，孝敬我的在哪裏呢？我既為主人，敬畏我的在哪裏呢？你們這些藐視我名的祭司啊！」你們卻說：「我們在何事上藐視你的名呢？」
MAL|1|7|「你們將不潔淨的食物獻在我的祭壇上，卻說：『我們在何事上使你不潔淨呢？』你們說，耶和華的供桌是可藐視的。
MAL|1|8|你們將瞎眼的獻為祭物，這不算為惡嗎？將瘸腿的、有病的獻上，這不算為惡嗎？那麼，請把這些獻給你的省長，他豈會悅納你 ，豈會抬舉你呢？這是萬軍之耶和華說的。」
MAL|1|9|現在我勸你們要懇求上帝，好讓他施恩給我們。這事既出於你們的手，他豈會抬舉你們任何人呢？這是萬軍之耶和華說的。
MAL|1|10|萬軍之耶和華說：「甚願你們中間有人把殿的門 關上，免得你們徒然在我壇上燒火。我不喜歡你們，也不從你們手中悅納供物。」
MAL|1|11|萬軍之耶和華說：「從日出之地到日落之處，我的名在列國中必尊為大。在各處，人必奉我的名燒香，獻潔淨的供物，因為我的名在列國中必尊為大。
MAL|1|12|你們卻褻瀆我的名，說：『主的供桌是不潔淨的，供桌上的果子和食物是可藐視的。』
MAL|1|13|你們又說：『看哪，這些事何等煩瑣！』並嗤之以鼻 。這是萬軍之耶和華說的。你們把搶來的、瘸腿的、有病的拿來獻上為祭，我豈能從你們手中悅納它呢？這是耶和華說的。
MAL|1|14|行詭詐的人是可詛咒的！他的群畜中雖有公羊，他許了願，卻將有殘疾的獻給主。因我是大君王，我的名在列國中是可畏的。這是萬軍之耶和華說的。」
MAL|2|1|現在，眾祭司啊，這誡命是給你們的。
MAL|2|2|萬軍之耶和華說：「你們若不聽，不放在心上，不將榮耀歸給我的名，我就使詛咒臨到你們，使你們的福分變為詛咒；其實我已經詛咒了你們的福分，因你們不把誡命放在心上。
MAL|2|3|看哪，我要斥責你們的後裔，把糞抹在你們臉上，就是你們祭牲 的糞。人要把你們和糞一起抬出去，
MAL|2|4|你們就知道我頒這誡命給你們，使我與 利未 所立的約可以常存。這是萬軍之耶和華說的。
MAL|2|5|我曾與他立生命和平安的約。我將這兩樣賜給他，使他存敬畏的心；他就敬畏我，懼怕我的名。
MAL|2|6|真實的訓誨在他口中，他的嘴唇中沒有不義。他以平安和正直與我同行，使許多人回轉離開罪孽。
MAL|2|7|祭司的嘴唇當守護知識，人也當從他口中尋求訓誨，因為他是萬軍之耶和華的使者。
MAL|2|8|你們卻偏離正道，使許多人在這訓誨上絆跌。你們破壞了我與 利未 人所立的約。這是萬軍之耶和華說的。
MAL|2|9|所以我使你們被眾百姓藐視，看為卑賤；因你們不遵守我的道，在律法上看人的情面 。」
MAL|2|10|我們豈不都有一位父嗎？豈不是一位上帝創造了我們嗎？為何互相行詭詐，褻瀆了上帝與我們列祖所立的約呢？
MAL|2|11|猶大 行事詭詐，在 以色列 和 耶路撒冷 中行了可憎的事；因為 猶大 人褻瀆耶和華所喜愛的聖殿，娶外邦神明的女子為妻。
MAL|2|12|凡做這事的，無論是清醒的 或回應的，即使獻供物給萬軍之耶和華，耶和華也要將他從 雅各 的帳棚中剪除。
MAL|2|13|你們又再做這樣的事，使哭泣和嘆息的眼淚遮蓋耶和華的祭壇，以致耶和華不再理會那供物，也不喜歡從你們的手中收納。
MAL|2|14|你們還說：「這是為甚麼呢？」因為耶和華在你和你年輕時所娶的妻之間作證。她雖是你的配偶，你誓約 的妻，你卻背棄她。
MAL|2|15|一個人如果還剩下一點靈性，他不會這麼做。這人在尋找甚麼呢？上帝的後裔！ 當謹守你們的靈性，誰也不可背棄年輕時所娶的妻。
MAL|2|16|耶和華－ 以色列 的上帝說：「我恨惡休妻的事和衣服外面披上暴力的人。所以當謹守你們的心，不可行詭詐。這是萬軍之耶和華說的。」
MAL|2|17|你們用言語使耶和華厭煩，卻說：「我們在何事上使他厭煩呢？」因為你們說：「凡行惡的，耶和華看為善，並且喜愛他們；」又說：「公平的上帝在哪裏呢？」
MAL|3|1|萬軍之耶和華說：「看哪，我要差遣我的使者在我前面預備道路。你們所尋求的主必忽然來到他的殿；立約的使者，就是你們所仰慕的，看哪，快要來到。」
MAL|3|2|他來的日子，誰能當得起呢？他顯現的時候，誰能立得住呢？因為他如煉金匠的火，如漂洗者的鹼。
MAL|3|3|他必坐下如煉淨銀子的人，必潔淨 利未 人，熬煉他們像金銀一樣；他們就憑公義獻供物給耶和華。
MAL|3|4|那時， 猶大 和 耶路撒冷 所獻的供物必蒙耶和華悅納，彷彿古時之日、上古之年。
MAL|3|5|萬軍之耶和華說：「我必臨近你們，施行審判。我必速速作見證，警戒那些行邪術的、犯姦淫的、起假誓的、剝削雇工工錢的、欺壓孤兒寡婦的、屈枉寄居者的和不敬畏我的人。」
MAL|3|6|「我－耶和華是不改變的；所以， 雅各 的子孫啊，你們不致滅亡。
MAL|3|7|從你們祖先的日子以來，你們就偏離我的律例而不遵守。現在你們要轉向我，我就轉向你們。這是萬軍之耶和華說的。你們卻說：『我們如何轉向呢？』
MAL|3|8|人豈可搶奪上帝呢？你們竟搶奪我！你們卻說：『我們在何事上搶奪你呢？』其實就是在你們當納的十分之一奉獻和當獻的供物上。
MAL|3|9|因你們全國上下都搶奪我的供物，詛咒就臨到你們身上。
MAL|3|10|你們要將當納的十分之一全然送入倉庫，使我家有糧，以此試試我，是否為你們敞開天上的窗戶，傾福與你們，甚至無處可容。這是萬軍之耶和華說的。
MAL|3|11|我必為你們斥責蝗蟲 ，不容牠毀壞你們的土產。你們田間的葡萄樹，果實未熟以先也不會掉落。這是萬軍之耶和華說的。
MAL|3|12|萬國必稱你們為有福的，因你們必成為喜樂之地。這是萬軍之耶和華說的。」
MAL|3|13|耶和華說：「你們用話頂撞我。」你們卻說：「我們說了甚麼話頂撞你呢？」
MAL|3|14|你們說：「事奉上帝是枉然，我們遵守上帝所吩咐的，在萬軍之耶和華面前哀痛而行，有甚麼益處呢？
MAL|3|15|現在，我們稱狂傲的人為有福，並且行惡的人得以建立；他們雖然試探上帝，卻得以逃脫。」
MAL|3|16|那時，敬畏耶和華的人彼此談論，耶和華側耳而聽，且有紀念冊在他面前，記錄那敬畏耶和華、思念他名的人。
MAL|3|17|萬軍之耶和華說：「在我所定的日子，他們必屬我，是我寶貴的產業。我必憐憫他們，如同人憐憫那服侍他的兒子。
MAL|3|18|那時你們必再一次 看出義人和惡人，事奉上帝和不事奉上帝的人有何差別。」
MAL|4|1|萬軍之耶和華說：「看哪，那日臨近，勢如燒著的火爐，凡狂傲的和行惡的都如碎秸，在那日被燒盡，根與枝條無一存留。
MAL|4|2|但是，對你們敬畏我名的人，必有公義的太陽出現，其光線 有醫治的能力。你們必出來跳躍如圈裏的牛犢。
MAL|4|3|你們必踐踏惡人；在我所定的日子，他們必成為你們腳掌下的灰塵。這是萬軍之耶和華說的。
MAL|4|4|「你們當記念我僕人 摩西 的律法，就是我在 何烈山 為 以色列 眾人所吩咐他的律例典章。
MAL|4|5|「看哪，耶和華大而可畏之日未到以前，我要差遣 以利亞 先知到你們那裏去。
MAL|4|6|他必使父親的心轉向兒女，兒女的心轉向父親，免得我來詛咒這地。」
MATT|1|1|亞伯拉罕 的後裔、 大衛 的子孫 耶穌基督的家譜：
MATT|1|2|亞伯拉罕 生 以撒 ， 以撒 生 雅各 ， 雅各 生 猶大 和他的兄弟，
MATT|1|3|猶大 從 她瑪 氏生 法勒斯 和 謝拉 ， 法勒斯 生 希斯崙 ， 希斯崙 生 亞蘭 ，
MATT|1|4|亞蘭 生 亞米拿達 ， 亞米拿達 生 拿順 ， 拿順 生 撒門 ，
MATT|1|5|撒門 從 喇合 氏生 波阿斯 ， 波阿斯 從 路得 氏生 俄備得 ， 俄備得 生 耶西 ，
MATT|1|6|耶西 生 大衛 王。 大衛 從 烏利亞 的妻子生 所羅門 ，
MATT|1|7|所羅門 生 羅波安 ， 羅波安 生 亞比雅 ， 亞比雅 生 亞撒 ，
MATT|1|8|亞撒 生 約沙法 ， 約沙法 生 約蘭 ， 約蘭 生 烏西雅 ，
MATT|1|9|烏西雅 生 約坦 ， 約坦 生 亞哈斯 ， 亞哈斯 生 希西家 ，
MATT|1|10|希西家 生 瑪拿西 ， 瑪拿西 生 亞們 ， 亞們 生 約西亞 ，
MATT|1|11|百姓被遷到 巴比倫 的時候， 約西亞 生 耶哥尼雅 和他的兄弟。
MATT|1|12|遷到 巴比倫 之後， 耶哥尼雅 生 撒拉鐵 ， 撒拉鐵 生 所羅巴伯 ，
MATT|1|13|所羅巴伯 生 亞比玉 ， 亞比玉 生 以利亞敬 ， 以利亞敬 生 亞所 ，
MATT|1|14|亞所 生 撒督 ， 撒督 生 亞金 ， 亞金 生 以律 ，
MATT|1|15|以律 生 以利亞撒 ， 以利亞撒 生 馬但 ， 馬但 生 雅各 ，
MATT|1|16|雅各 生 約瑟 ，就是 馬利亞 的丈夫；那稱為基督的耶穌是從 馬利亞 生的。
MATT|1|17|這樣，從 亞伯拉罕 到 大衛 共有十四代，從 大衛 到遷至 巴比倫 的時候也有十四代，從遷至 巴比倫 的時候到基督又有十四代。
MATT|1|18|耶穌基督降生的事記在下面：他母親 馬利亞 已經許配給 約瑟 ，還沒有迎娶， 馬利亞 就從聖靈懷了孕。
MATT|1|19|她丈夫 約瑟 是個義人，不願意當眾羞辱她，想要暗地裏把她休了。
MATT|1|20|正考慮這些事的時候，忽然主的使者在 約瑟 夢中向他顯現，說：「 大衛 的子孫 約瑟 ，不要怕，把你的妻子 馬利亞 娶過來，因她所懷的孕是從聖靈來的。
MATT|1|21|她將要生一個兒子，你要給他起名叫耶穌，因他要將自己的百姓從罪惡裏救出來。」
MATT|1|22|這整件事的發生，是要應驗主藉先知所說的話：
MATT|1|23|「必有童女懷孕生子； 人要稱他的名為 以馬內利 。」 （ 以馬內利 翻出來就是「上帝與我們同在」。）
MATT|1|24|約瑟 醒來，就遵照主的使者的吩咐把妻子娶過來；
MATT|1|25|但是沒有和她同房，直到她生了兒子 ，就給他起名叫耶穌。
MATT|2|1|在 希律 作王的時候，耶穌生在 猶太 的 伯利恆 。有幾個博學之士 從東方來到 耶路撒冷 ，說：
MATT|2|2|「那生下來作 猶太 人之王的在哪裏？我們在東方看見他的星，特來拜他。」
MATT|2|3|希律 王聽見了，就心裏不安； 耶路撒冷 全城的人也都不安。
MATT|2|4|他就召集了祭司長和民間的文士，問他們：「基督該生在哪裏？」
MATT|2|5|他們說：「在 猶太 的 伯利恆 。因為有先知記著：
MATT|2|6|『 猶大 地的 伯利恆 啊， 你在 猶大 諸城中並不是最小的； 因為將來有一位統治者要從你那裏出來， 牧養我 以色列 民。』」
MATT|2|7|於是， 希律 暗地裏召了博學之士來，查問那星是甚麼時候出現的，
MATT|2|8|就派他們往 伯利恆 去，說：「你們去仔細尋訪那小孩子，找到了就來報信，我也好去拜他。」
MATT|2|9|他們聽了王的話就去了。忽然，在東方所看到的那顆星在前面引領他們，一直行到小孩子所在地方的上方就停住了。
MATT|2|10|他們看見那星，就非常歡喜；
MATT|2|11|進了房子，看見小孩子和他母親 馬利亞 ，就俯伏拜那小孩子，揭開寶盒，拿出黃金、乳香、沒藥，作為禮物獻給他。
MATT|2|12|因為在夢中得到主的指示，不要回去見 希律 ，他們就從別的路回自己的家鄉去了。
MATT|2|13|他們走後，忽然主的使者在 約瑟 夢中向他顯現，說：「起來！帶著小孩子和他母親逃往 埃及 ，住在那裏，等我的指示；因為 希律 要搜尋那小孩子來殺害他。」
MATT|2|14|約瑟 就起來，連夜帶著小孩子和他母親往 埃及 去，
MATT|2|15|住在那裏，直到 希律 死了。這是要應驗主藉先知所說的話：「我從 埃及 召我的兒子出來。」
MATT|2|16|希律 見自己被博學之士愚弄，極其憤怒，差人將 伯利恆 城裏和四境所有的男孩，根據他向博學之士仔細查問到的時間，凡兩歲以內的，都殺盡了。
MATT|2|17|這就應驗了 耶利米 先知所說的話：
MATT|2|18|「在 拉瑪 聽見號咷大哭的聲音， 是 拉結 哭她兒女； 她不肯受安慰， 因為他們都不在了。」
MATT|2|19|希律 死了以後，在 埃及 ，忽然主的使者在 約瑟 夢中向他顯現，
MATT|2|20|說：「起來，帶著小孩子和他母親回 以色列 地去！因為要殺害這小孩子的人已經死了。」
MATT|2|21|約瑟 就起來，帶著小孩子和他母親進入 以色列 地去。
MATT|2|22|但是他因聽見 亞基老 繼承他父親 希律 作了 猶太 王，怕到那裏去；又在夢中得到主的指示，就往 加利利 境內去了。
MATT|2|23|他們到了一座城，名叫 拿撒勒 ，就住在那裏。這是要應驗先知所說的話：「他將稱為 拿撒勒 人。」
MATT|3|1|在那些日子，施洗的 約翰 出來，在 猶太 的曠野宣講：
MATT|3|2|「你們要悔改！因為天國近了。」
MATT|3|3|這人就是 以賽亞 先知所說的： 「在曠野有聲音呼喊著： 預備主的道， 修直他的路。」
MATT|3|4|這 約翰 身穿駱駝毛的衣服，腰束皮帶，吃的是蝗蟲和野蜜。
MATT|3|5|那時， 耶路撒冷 、全 猶太 和全 約旦河 地區的人，都到 約翰 那裏去，
MATT|3|6|承認他們的罪，在 約旦河 裏受他的洗。
MATT|3|7|約翰 看見許多法利賽人和撒都該人也來受洗，就對他們說：「毒蛇的孽種啊，誰指示你們逃避那將要來的憤怒呢？
MATT|3|8|你們要結出果子來，和悔改的心相稱。
MATT|3|9|不要自己心裏說：『我們有 亞伯拉罕 為祖宗。』我告訴你們，上帝能從這些石頭中給 亞伯拉罕 興起子孫來。
MATT|3|10|現在斧子已經放在樹根上，凡不結好果子的樹就砍下來，丟在火裏。
MATT|3|11|我是用水給你們施洗，叫你們悔改；但那在我以後來的，能力比我更大，我就是給他提鞋子也不配，他要用聖靈與火給你們施洗。
MATT|3|12|他手裏拿著簸箕，要揚淨他的穀物，把麥子收在倉裏，把糠用不滅的火燒盡。」
MATT|3|13|當時，耶穌從 加利利 來到 約旦河 ，到了 約翰 那裏，請 約翰 為他施洗。
MATT|3|14|約翰 想要阻止他，說：「我應該受你的洗，你怎麼到我這裏來呢？」
MATT|3|15|耶穌回答他：「暫且這樣做吧，因為我們理當這樣履行全部的義 。」於是 約翰 就依了他。
MATT|3|16|耶穌受了洗，隨即從水裏上來。天忽然為他 開了，他看見上帝的靈降下，彷彿鴿子落在他身上。
MATT|3|17|這時，天上有聲音說：「這是我的愛子，我所喜愛的。」
MATT|4|1|當時，耶穌被聖靈引到曠野，受魔鬼的試探。
MATT|4|2|他禁食四十晝夜，後來就餓了。
MATT|4|3|那試探者進前來對他說：「你若是上帝的兒子，叫這些石頭變成食物吧。」
MATT|4|4|耶穌卻回答說：「經上記著： 『人活著，不是單靠食物， 乃是靠上帝口裏所出的一切話。』」
MATT|4|5|魔鬼就帶他進了聖城，叫他站在聖殿頂上，
MATT|4|6|對他說：「你若是上帝的兒子，就跳下去！因為經上記著： 『主要為你命令他的使者， 用手托住你， 免得你的腳碰在石頭上。』」
MATT|4|7|耶穌對他說：「經上又記著：『不可試探主—你的上帝。』」
MATT|4|8|魔鬼又帶他上了一座很高的山，將世上的萬國和萬國的榮華都指給他看，
MATT|4|9|對他說：「你若俯伏拜我，我就把這一切賜給你。」
MATT|4|10|耶穌說：「撒但 ，退去！因為經上記著： 『要拜主—你的上帝， 惟獨事奉他。』」
MATT|4|11|於是，魔鬼離開了耶穌，立刻有天使來伺候他。
MATT|4|12|耶穌聽見 約翰 下了監，就退到 加利利 去；
MATT|4|13|後來離開 拿撒勒 ，往 迦百農 去，住在那裏。那地方靠海，在 西布倫 和 拿弗他利 地區。
MATT|4|14|這是要應驗 以賽亞 先知所說的話：
MATT|4|15|「 西布倫 ， 拿弗他利 ， 沿海的路， 約旦河 的東邊， 外邦人的 加利利 —
MATT|4|16|那坐在黑暗裏的百姓 看見了大光； 坐在死蔭之地的人 有光照耀他們。」
MATT|4|17|從那時候，耶穌開始宣講，說：「你們要悔改！因為天國近了。」
MATT|4|18|耶穌沿著 加利利 海邊行走，看見兩兄弟，就是那叫 彼得 的 西門 和他弟弟 安得烈 ，正往海裏撒網；他們本是打魚的。
MATT|4|19|耶穌對他們說：「來跟從我，我要叫你們得人如得魚一樣。」
MATT|4|20|他們立刻捨了網，跟從他。
MATT|4|21|耶穌從那裏往前走，看見另外兩兄弟，就是 西庇太 的兒子 雅各 和他弟弟 約翰 ，同他們的父親 西庇太 在船上補網，耶穌就呼召他們。
MATT|4|22|他們立刻捨了船，辭別父親，跟從了耶穌。
MATT|4|23|耶穌走遍 加利利 ，在各會堂裏教導人，宣講天國的福音，醫治百姓各樣的疾病。
MATT|4|24|他的名聲傳遍了 敘利亞 。那裏的人把一切病人，就是有各樣疾病和疼痛的、被鬼附的、癲癇的、癱瘓的，都帶了來，耶穌就治好了他們。
MATT|4|25|當時，有一大群人從 加利利 、 低加坡里 、 耶路撒冷 、 猶太 、 約旦河 的東邊，來跟從他。
MATT|5|1|耶穌看見這一群人，就上了山，坐下後，門徒到他跟前來，
MATT|5|2|他開口教導他們說：
MATT|5|3|「心靈貧窮的人有福了！ 因為天國是他們的。
MATT|5|4|哀慟的人有福了！ 因為他們必得安慰。
MATT|5|5|謙和的人有福了！ 因為他們必承受土地。
MATT|5|6|飢渴慕義的人有福了！ 因為他們必得飽足。
MATT|5|7|憐憫人的人有福了！ 因為他們必蒙憐憫。
MATT|5|8|清心的人有福了！ 因為他們必得見上帝。
MATT|5|9|締造和平的人有福了！ 因為他們必稱為上帝的兒子。
MATT|5|10|為義受迫害的人有福了！ 因為天國是他們的。
MATT|5|11|「人若因我辱罵你們，迫害你們，捏造各樣壞話毀謗你們 ，你們就有福了！
MATT|5|12|要歡喜快樂，因為你們在天上的賞賜是很多的。在你們以前的先知，人也是這樣迫害他們。」
MATT|5|13|「你們是地上的鹽。鹽若失了味，怎能叫它再鹹呢？它不再有用，只好被丟在外面，任人踐踏。
MATT|5|14|你們是世上的光。城造在山上是不能隱藏的。
MATT|5|15|人點燈，不放在斗底下，而是放在燈臺上，就照亮一家的人。
MATT|5|16|你們的光也要這樣照在人前，叫他們看見你們的好行為，把榮耀歸給你們在天上的父。」
MATT|5|17|「不要以為我來是要廢掉律法和先知。我來不是要廢掉，而是要成全。
MATT|5|18|我實在告訴你們，就是到天地都廢去，律法的一點一畫也不能廢去，直到一切都實現。
MATT|5|19|所以，無論誰廢掉這誡命中最小的一條，又教導人也這樣做，他在天國裏要稱為最小的。但無論誰遵行並如此教導人的，他在天國裏要稱為大。
MATT|5|20|我告訴你們，你們的義若不勝過文士和法利賽人的義，絕不能進天國。」
MATT|5|21|「你們聽過有對古人說：『不可殺人』；『凡殺人的，必須受審判。』
MATT|5|22|但是我告訴你們：凡向弟兄動怒的，必須受審判；凡罵弟兄是廢物的，必須受議會的審判；凡罵弟兄是白痴的，必須遭受地獄的火。
MATT|5|23|所以，你在祭壇上獻祭物的時候，若想起有弟兄對你懷恨，
MATT|5|24|就要把祭物留在壇前，先去跟弟兄和好，然後來獻祭物。
MATT|5|25|你同告你的冤家還在路上，就要趕快與他講和，免得他把你送交給法官，法官交給警衛，你就下在監裏了。
MATT|5|26|我實在告訴你，就是有一個大文錢 還沒有還清，你也絕不能從那裏出來。」
MATT|5|27|「你們聽過有話說：『不可姦淫。』
MATT|5|28|但是我告訴你們：凡看見婦女就動淫念的，這人心裏已經與她犯姦淫了。
MATT|5|29|若是你的右眼使你跌倒，就把它挖出來，丟掉。寧可失去身體中的一部分，也不讓整個身體被扔進地獄。
MATT|5|30|若是你的右手使你跌倒，就把它砍下來，丟掉。寧可失去身體中的一部分，也不讓整個身體下地獄。」
MATT|5|31|「又有話說：『無論誰休妻，都要給她休書。』
MATT|5|32|但是我告訴你們：凡休妻的，除非是因不貞的緣故，否則就是使她犯姦淫了；人若娶被休的婦人，也是犯姦淫了。」
MATT|5|33|「你們又聽過有對古人說：『不可背誓，所起的誓總要向主謹守。』
MATT|5|34|但是我告訴你們：甚麼誓都不可起。不可指著天起誓，因為天是上帝的寶座。
MATT|5|35|不可指著地起誓，因為地是他的腳凳；也不可指著 耶路撒冷 起誓，因為 耶路撒冷 是大君王的京城。
MATT|5|36|又不可指著你的頭起誓，因為你不能使一根頭髮變黑變白。
MATT|5|37|你們的話，是，就說是；不是，就說不是。若再多說，就是出於那惡者。」
MATT|5|38|「你們聽過有話說：『以眼還眼，以牙還牙。』
MATT|5|39|但是我告訴你們：不要與惡人作對。有人打你的右臉，連另一邊也轉過去由他打。
MATT|5|40|有人想要告你，要拿你的裏衣，連外衣也由他拿去。
MATT|5|41|有人強迫你走一里 路，你就跟他走二里。
MATT|5|42|有求你的，就給他；有向你借貸的，不可推辭。」
MATT|5|43|「你們聽過有話說：『要愛你的鄰舍，恨你的仇敵。』
MATT|5|44|但是我告訴你們：要愛你們的仇敵，為那迫害你們的禱告。
MATT|5|45|這樣，你們就可以作天父的兒女了。因為他叫太陽照好人，也照壞人；降雨給義人，也給不義的人。
MATT|5|46|你們若只愛那愛你們的人，有甚麼賞賜呢？就是稅吏不也是這樣做嗎？
MATT|5|47|你們若只請你弟兄的安，有甚麼比別人強呢？就是外邦人不也是這樣做嗎？
MATT|5|48|所以，你們要完全，如同你們的天父是完全的。」
MATT|6|1|「你們要謹慎，不可故意在人面前表現虔誠，叫他們看見，若是這樣，就不能得你們天父的賞賜了。
MATT|6|2|「所以，你施捨的時候，不可叫人在你前面吹號，像那假冒為善的人在會堂裏和街道上所做的，故意要得人的稱讚。我實在告訴你們，他們已經得了他們的賞賜。
MATT|6|3|你施捨的時候，不要讓左手知道右手所做的，
MATT|6|4|好使你隱祕地施捨；你父在隱祕中察看，必然賞賜你。」
MATT|6|5|「你們禱告的時候，不可像那假冒為善的人，愛站在會堂裏和十字路口禱告，故意讓人看見。我實在告訴你們，他們已經得了他們的賞賜。
MATT|6|6|你禱告的時候，要進入內室，關上門，向那在隱祕中的父禱告；你父在隱祕中察看，必將賞賜你。
MATT|6|7|你們禱告，不可像外邦人那樣重複一些空話，他們以為話多了必蒙垂聽。
MATT|6|8|你們不可效法他們。因為在你們祈求以前，你們所需要的，你們的父早已知道了。」
MATT|6|9|「所以，你們要這樣禱告： 『我們在天上的父： 願人都尊你的名為聖。
MATT|6|10|願你的國降臨； 願你的旨意行在地上， 如同行在天上。
MATT|6|11|我們日用的飲食，今日賜給我們。
MATT|6|12|免我們的債， 如同我們免了人的債。
MATT|6|13|不叫我們陷入試探； 救我們脫離那惡者。 因為國度、權柄、榮耀，全是你的， 直到永遠。阿們！ 』
MATT|6|14|「你們若饒恕人的過犯，你們的天父也必饒恕你們；
MATT|6|15|你們若不饒恕人 ，你們的天父也必不饒恕你們的過犯。」
MATT|6|16|「你們禁食的時候，不可像那假冒為善的人，臉上帶著愁容；因為他們蓬頭垢面，故意讓人看出他們在禁食。我實在告訴你們，他們已經得了他們的賞賜。
MATT|6|17|你禁食的時候，要梳頭洗臉，
MATT|6|18|不要讓人看出你在禁食，只讓你隱祕中的父看見；你父在隱祕中察看，必然賞賜你。」
MATT|6|19|「不要為自己在地上積蓄財寶；地上有蟲子咬，能銹壞，也有賊挖洞來偷。
MATT|6|20|要在天上積蓄財寶；天上沒有蟲子咬，不會銹壞，也沒有賊挖洞來偷。
MATT|6|21|因為你的財寶在哪裏，你的心也在哪裏。」
MATT|6|22|「眼睛是身體的燈。你的眼睛若明亮，全身就光明；
MATT|6|23|你的眼睛若昏花，全身就黑暗。你裏面的光若黑暗了，那黑暗是何等大呢！」
MATT|6|24|「一個人不能服侍兩個主；他不是恨這個愛那個，就是重這個輕那個。你們不能又服侍上帝，又服侍 瑪門 。」
MATT|6|25|「所以，我告訴你們，不要為你們的生命憂慮吃甚麼喝甚麼 ，或為你們的身體憂慮穿甚麼。生命不勝於飲食嗎？身體不勝於衣裳嗎？
MATT|6|26|你們看一看那天上的飛鳥，也不種也不收，也不在倉裏存糧，你們的天父尚且養活牠們。你們不比飛鳥貴重得多嗎？
MATT|6|27|你們哪一個能藉著憂慮使壽數多加一刻呢 ？
MATT|6|28|何必為衣裳憂慮呢？你們想一想野地裏的百合花是怎麼長起來的：它也不勞動也不紡線。
MATT|6|29|然而我告訴你們，就是 所羅門 極榮華的時候，他所穿戴的還不如這些花的一朵呢！
MATT|6|30|你們這小信的人哪！野地裏的草今天還在，明天就丟在爐裏，上帝還給它這樣的妝飾，何況你們呢？
MATT|6|31|所以，不要憂慮，說：『我們吃甚麼？喝甚麼？穿甚麼？』
MATT|6|32|這都是外邦人所求的。你們需要這一切東西，你們的天父都知道。
MATT|6|33|你們要先求上帝的國和他的義，這些東西都要加給你們了。
MATT|6|34|所以，不要為明天憂慮，因為明天自有明天的憂慮；一天的難處一天當就夠了。」
MATT|7|1|「你們不要評斷別人，免得你們被審判。
MATT|7|2|因為你們怎樣評斷別人，也必怎樣被審判；你們用甚麼量器量給人，也必用甚麼量器量給你們。
MATT|7|3|為甚麼看見你弟兄眼中有刺，卻不想自己眼中有梁木呢？
MATT|7|4|你自己眼中有梁木，怎能對你弟兄說『讓我去掉你眼中的刺』呢？
MATT|7|5|你這假冒為善的人！先去掉自己眼中的梁木，然後才能看得清楚，好去掉你弟兄眼中的刺。
MATT|7|6|不要把聖物給狗，也不要把你們的珍珠丟在豬面前，恐怕牠們踐踏了珍珠，轉過來咬你們。」
MATT|7|7|「你們祈求，就給你們；尋找，就找到；叩門，就給你們開門。
MATT|7|8|因為凡祈求的，就得著；尋找的，就找到；叩門的，就給他開門。
MATT|7|9|你們中間誰有兒子求餅，反給他石頭呢？
MATT|7|10|求魚，反給他蛇呢？
MATT|7|11|你們雖然不好，尚且知道拿好東西給兒女，何況你們在天上的父，他豈不更要把好東西賜給求他的人嗎？
MATT|7|12|所以，無論何事，你們想要人怎樣待你們，你們也要怎樣待人，因為這就是律法和先知的道理。」
MATT|7|13|「你們要進窄門。因為通往滅亡的門是寬的，路是大的，進去的人也多；
MATT|7|14|通往生命的門是窄的，路是小的，找到的人也少。」
MATT|7|15|「你們要防備假先知。他們到你們這裏來，外面披著羊皮，裏面卻是殘暴的狼。
MATT|7|16|豈能在荊棘上摘葡萄呢？豈能在蒺藜裏摘無花果呢？憑著他們的果子，就可以認出他們來。
MATT|7|17|這樣，凡好樹都結好果子，而壞樹結壞果子。
MATT|7|18|好樹不能結壞果子，壞樹也不能結好果子。
MATT|7|19|凡不結好果子的樹就砍下來，丟在火裏。
MATT|7|20|所以，憑著他們的果子就可以認出他們來。」
MATT|7|21|「不是每一個稱呼我『主啊，主啊』的人都能進天國；惟有遵行我天父旨意的人才能進去。
MATT|7|22|在那日必有許多人對我說：『主啊，主啊，我們不是奉你的名傳道，奉你的名趕鬼，奉你的名行許多異能嗎？』
MATT|7|23|我要向他們宣告：『我從來不認識你們，你們這些作惡的人，給我走開！』」
MATT|7|24|「所以，凡聽了我這些話又去做的，好比一個聰明人把房子蓋在磐石上。
MATT|7|25|風吹，雨打，水沖，撞擊那房子，房子總不倒塌，因為根基立在磐石上。
MATT|7|26|凡聽了我這些話而不去做的，好比一個無知的人把房子蓋在沙土上。
MATT|7|27|風吹，雨打，水沖，撞擊那房子，房子就倒塌了，並且倒塌得很厲害。」
MATT|7|28|耶穌講完了這些話，眾人對他的教導都感到驚奇，
MATT|7|29|因為他教導他們正像有權柄的人，不像他們的文士。
MATT|8|1|耶穌下了山，有一大群人跟著他。
MATT|8|2|這時，一個痲瘋病人前來拜他，說：「主啊，你若肯，你能使我潔淨。」
MATT|8|3|耶穌伸手摸他，說：「我肯，你潔淨了吧！」他的痲瘋病立刻就潔淨了。
MATT|8|4|耶穌對他說：「你要注意，不可告訴任何人，只要去，讓祭司為你檢查，並獻上 摩西 所吩咐的祭物，作為證據給眾人看。」
MATT|8|5|耶穌進了 迦百農 ，有一個百夫長進前來，求他，
MATT|8|6|說：「主啊，我的僮僕癱瘓了，躺在家裏，非常痛苦。」
MATT|8|7|耶穌說：「我去醫治他。」
MATT|8|8|百夫長回答：「主啊，你到舍下來，我不敢當；只要你說一句話，我的僮僕就會痊癒。
MATT|8|9|因為我在人的權下，也有兵在我以下。我對這個說：『去！』他就去；對那個說：『來！』他就來；對我的僕人說：『做這事！』他就去做。」
MATT|8|10|耶穌聽了就很驚訝，對跟從的人說：「我實在告訴你們，這麼大的信心，就是在 以色列 ，我也沒有見過。
MATT|8|11|我又告訴你們，從東從西，將有許多人來，在天國裏與 亞伯拉罕 、 以撒 、 雅各 一同坐席；
MATT|8|12|本國的子民反而被趕到外邊黑暗裏去，在那裏要哀哭切齒了。」
MATT|8|13|耶穌對百夫長說：「你回去吧！照你的信心成全你了。」就在那時，他的僮僕好了。
MATT|8|14|耶穌到了 彼得 家裏，見 彼得 的岳母正發燒躺著。
MATT|8|15|耶穌一摸她的手，燒就退了，於是她起來服事耶穌。
MATT|8|16|傍晚的時候，有人帶著許多被鬼附的來到耶穌跟前，他只用一句話就把邪靈都趕出去，並且治好了一切有病的人。
MATT|8|17|這是要應驗 以賽亞 先知所說的話： 「他代替了我們的軟弱， 擔當了我們的疾病。」
MATT|8|18|耶穌見許多人圍著他，就吩咐渡到對岸去。
MATT|8|19|有一個文士進前來對他說：「老師，你無論往哪裏去，我都要跟從你。」
MATT|8|20|耶穌說：「狐狸有洞，天空的飛鳥有窩，人子卻沒有枕頭的地方。」
MATT|8|21|又有一個門徒對耶穌說：「主啊，容許我先回去埋葬我的父親。」
MATT|8|22|耶穌說：「讓死人埋葬他們的死人。你跟從我吧！」
MATT|8|23|耶穌上了船，門徒跟著他。
MATT|8|24|海裏忽然起了猛烈的風暴，以致船幾乎被波浪淹沒，耶穌卻睡著了。
MATT|8|25|門徒去叫醒他，說：「主啊，救命啊，我們快沒命啦！」
MATT|8|26|耶穌說：「你們這些小信的人哪，為甚麼膽怯呢？」於是他起來，斥責風和海，風和海就大大平靜了。
MATT|8|27|眾人驚訝地說：「這是怎樣的一個人？連風和海都聽從他。」
MATT|8|28|耶穌渡到對岸去，到 加大拉 人 的地區，有兩個被鬼附的人從墳墓迎著他走來。他們極其兇猛，甚至沒有人敢從那條路經過。
MATT|8|29|他們喊著說：「上帝的兒子，你為甚麼干擾我們？時候還沒有到，你就上這裏來叫我們受苦嗎？」
MATT|8|30|離他們很遠，有一大群豬正在吃食。
MATT|8|31|鬼就央求耶穌，說：「若要把我們趕出去，就打發我們進入豬群吧！」
MATT|8|32|耶穌對他們說：「去吧！」鬼就出來，進入豬群。一轉眼，整群豬都闖下山崖，投進海裏，淹死了。
MATT|8|33|放豬的就逃進城去，把這一切事和被鬼附的人所遭遇的都告訴眾人。
MATT|8|34|全城的人都出來迎見耶穌，見了他以後，就央求他離開他們的地區。
MATT|9|1|耶穌上了船，渡過海，來到自己的城裏。
MATT|9|2|有人用褥子抬著一個癱子到耶穌跟前來。耶穌見他們的信心，就對癱子說：「孩子，放心吧，你的罪赦了。」
MATT|9|3|這時，有幾個文士心裏說：「這個人說褻瀆的話了。」
MATT|9|4|耶穌知道他們的心思，就說：「你們心裏為甚麼懷著惡念呢？
MATT|9|5|說『你的罪赦了』，或說『你起來行走』，哪一樣容易呢？
MATT|9|6|但要讓你們知道，人子在地上有赦罪的權柄」，於是對癱子說：「起來！拿你的褥子回家去吧。」
MATT|9|7|那人就起來，回家去了。
MATT|9|8|眾人看見都畏懼，歸榮耀給上帝，因為他把這樣的權柄賜給人。
MATT|9|9|耶穌從那裏往前走，看見一個人名叫 馬太 ，在稅關坐著，就對他說：「來跟從我！」他就起來跟從耶穌。
MATT|9|10|耶穌在屋裏坐席的時候，有好些稅吏和罪人來，與耶穌和他的門徒一同坐席。
MATT|9|11|法利賽人看見，就對耶穌的門徒說：「你們的老師為甚麼與稅吏和罪人一同吃飯呢？」
MATT|9|12|耶穌聽見，就說：「健康的人用不著醫生；有病的人才用得著。
MATT|9|13|經上說：『我喜愛憐憫，不喜愛祭祀。』這句話的意思，你們去揣摩。我不是來召義人，而是召罪人。」
MATT|9|14|那時， 約翰 的門徒來見耶穌，說：「我們和法利賽人常常 禁食，你的門徒卻不禁食，這是為甚麼呢？」
MATT|9|15|耶穌對他們說：「新郎和賓客在一起的時候，賓客怎麼能哀慟呢？但日子將到，新郎要被帶走，那時候他們就要禁食了。
MATT|9|16|沒有人把新布補在舊衣服上；因為所補上的會撕破那衣服，裂口就更大了。
MATT|9|17|也沒有人把新酒裝在舊皮袋裏，若是這樣，皮袋會脹破，酒就漏出來，皮袋也糟蹋了。相反地，把新酒裝在新皮袋裏，兩樣就都保全了。」
MATT|9|18|耶穌說這些話的時候，有一個會堂主管來，向他下跪，說：「我女兒剛死了，求你去按手在她身上，她就會活過來。」
MATT|9|19|耶穌就起來跟他去；門徒也跟了去。
MATT|9|20|這時，有一個女人，患了經血不止的病有十二年，來到耶穌背後，摸他的衣裳繸子；
MATT|9|21|因為她心裏說：「我只要摸他的衣裳，就會痊癒。」
MATT|9|22|耶穌轉過來，看見她，就說：「女兒，放心！你的信救了你。」從那時起，這女人就痊癒了。
MATT|9|23|耶穌到了會堂主管的家裏，看見吹鼓手和亂哄哄的一群人，
MATT|9|24|就說：「退去吧！這女孩不是死了，而是睡著了。」他們就嘲笑他。
MATT|9|25|眾人被趕出後，耶穌就進去，拉著女孩的手，女孩就起來了。
MATT|9|26|於是這消息傳遍了那地方。
MATT|9|27|耶穌從那裏往前走，有兩個盲人跟著他，喊叫說：「 大衛 之子，可憐我們吧！」
MATT|9|28|耶穌進了屋子，盲人就來到他跟前。耶穌說：「你們信我能做這事嗎？」他們說：「主啊，我們信。」
MATT|9|29|耶穌就摸他們的眼睛，說：「照著你們的信心成全你們吧。」
MATT|9|30|他們的眼睛就開了。耶穌嚴嚴地叮囑他們說：「要小心，不可讓人知道。」
MATT|9|31|他們出去，竟把他的名聲傳遍了那地方。
MATT|9|32|他們出去的時候，有人把一個被鬼附的啞巴帶到耶穌跟前來。
MATT|9|33|鬼被趕出去，啞巴就說出話來。眾人都很驚訝，說：「在 以色列 ，從來沒有見過這樣的事。」
MATT|9|34|法利賽人卻說：「他是靠著鬼王趕鬼的。」
MATT|9|35|耶穌走遍各城各鄉，在他們的會堂裏教導人，宣講天國的福音，又醫治各樣的病症。
MATT|9|36|他看見一大群人，就憐憫他們；因為他們困苦無助，如同羊沒有牧人一樣。
MATT|9|37|於是他對門徒說：「要收的莊稼多，做工的人少。
MATT|9|38|所以，你們要求莊稼的主差遣做工的人出去收他的莊稼。」
MATT|10|1|耶穌叫了十二個門徒來，給他們權柄，能驅趕污靈和醫治各樣的疾病。
MATT|10|2|這十二使徒的名字如下：頭一個叫 西門 （又稱 彼得 ），還有他弟弟 安得烈 ， 西庇太 的兒子 雅各 和 雅各 的弟弟 約翰 ，
MATT|10|3|腓力 和 巴多羅買 ， 多馬 和稅吏 馬太 ， 亞勒腓 的兒子 雅各 ，和 達太 ，
MATT|10|4|激進黨的 西門 ，還有出賣耶穌的 加略 人 猶大 。
MATT|10|5|耶穌差遣這十二個人出去，吩咐他們說：「外邦人的路，你們不要走； 撒瑪利亞 人的城，你們不要進；
MATT|10|6|寧可往 以色列 家迷失的羊那裏去。
MATT|10|7|要邊走邊傳，說『天國近了』。
MATT|10|8|要醫治病人，使死人復活，使痲瘋病人潔淨，把鬼趕出去。你們白白地得來，也要白白地給人。
MATT|10|9|腰袋裏不要帶金銀銅錢；
MATT|10|10|途中不要帶行囊，不要帶兩件內衣，也不要帶鞋子和手杖，因為工人得飲食是應當的。
MATT|10|11|你們無論進哪一城、哪一村，要打聽那裏誰是合適的人，就住在他家，直住到離開的時候。
MATT|10|12|進他家時，要向那家請安。
MATT|10|13|那家若配得平安，你們所求的平安就臨到那家；若不配得，你們所求的平安仍歸你們。
MATT|10|14|凡不接待你們，不聽你們話的人，你們離開那家，或是那城的時候，要跺掉你們腳上的塵土。
MATT|10|15|我實在告訴你們，在審判的日子， 所多瑪 和 蛾摩拉 地方所受的，比那城還容易受呢！」
MATT|10|16|「看哪！我差你們出去，如同羊進入狼群，所以你們要機警如蛇，純真如鴿。
MATT|10|17|你們要防備那些人，因為他們要把你們交給議會，也要在會堂裏鞭打你們。
MATT|10|18|你們要為我的緣故被送到統治者和君王面前，對他們和外邦人作見證。
MATT|10|19|當人把你們交出時，不要擔心怎樣說話，或說甚麼話。到那時候，必賜給你們該說的話，
MATT|10|20|因為不是你們自己說的，而是你們父的靈在你們裏面說的。
MATT|10|21|兄弟要把兄弟、父親要把兒女置於死地；兒女要起來與父母為敵，害死他們。
MATT|10|22|而且你們要為我的名被眾人憎恨。但堅忍到底的終必得救。
MATT|10|23|有人在這城迫害你們，就逃到另一城去。 我實在告訴你們， 以色列 的城鎮，你們還沒有走遍，人子就要來臨。
MATT|10|24|「學生不高過老師，僕人不高過主人。
MATT|10|25|學生所遭遇的與老師一樣，僕人所遭遇的與主人一樣，也就夠了。既然有人罵一家的主人是『 別西卜 』 ，更何況他的家人呢？」
MATT|10|26|「所以，不要怕他們，因為掩蓋的事沒有不顯露出來的，隱藏的事也沒有不被知道的。
MATT|10|27|我在暗中告訴你們的，你們要在明處說出來；你們耳中所聽的，要在屋頂上宣揚出來。
MATT|10|28|那殺人身體但不能滅人靈魂的，不要怕他們；惟有那能在地獄裏毀滅身體和靈魂的，才要怕他。
MATT|10|29|兩隻麻雀不是賣一銅錢 嗎？你們的父若不許，一隻也不會掉在地上。
MATT|10|30|就是你們的頭髮也都數過了。
MATT|10|31|所以，不要懼怕，你們比許多的麻雀還貴重！」
MATT|10|32|「所以，凡在人面前認我的，我在我天上的父面前也必認他；
MATT|10|33|凡在人面前不認我的，我在我天上的父面前也必不認他。」
MATT|10|34|「你們不要以為我來是帶給地上和平，我來並不是帶來和平，而是刀劍。
MATT|10|35|因為我來是要叫 『人與父親對立， 女兒與母親對立， 媳婦與婆婆對立。
MATT|10|36|人的仇敵就是自己家裏的人。』
MATT|10|37|愛父母勝過愛我的，不配作我的門徒；愛兒女勝過愛我的，不配作我的門徒。
MATT|10|38|不背自己的十字架跟從我的，不配作我的門徒。
MATT|10|39|得著性命的，要喪失性命；為我喪失性命的，要得著性命。」
MATT|10|40|「接納你們的就是接納我；接納我的就是接納差遣我來的那位。
MATT|10|41|把先知當作先知接納的，必得先知的賞賜；把義人當作義人接納的，必得義人的賞賜。
MATT|10|42|無論誰，只因門徒的名，就算把一杯涼水給這些小子中的一個喝，我實在告訴你們，他一定會得到賞賜。」
MATT|11|1|耶穌吩咐完了十二個門徒，就離開那裏，往各城去傳道，教導人。
MATT|11|2|約翰 在監獄裏聽見基督所做的事，就派他的門徒去，
MATT|11|3|問耶穌：「將要來的那位就是你嗎？還是我們要等候另一位呢？」
MATT|11|4|耶穌回答他們：「你們去，把所聽見、所看見的告訴 約翰 ：
MATT|11|5|就是盲人看見，瘸子行走，痲瘋病人得潔淨，聾子聽見，死人復活，窮人聽到福音。
MATT|11|6|凡不因我跌倒的有福了！」
MATT|11|7|他們一走，耶穌就對眾人談到 約翰 ，說：「你們從前到曠野去，是要看甚麼呢？看風吹動的蘆葦嗎？
MATT|11|8|你們出去到底是要看甚麼？看穿細軟衣服的人嗎？那穿細軟衣服的人是在王宮裏。
MATT|11|9|你們出去究竟是要看甚麼？是先知嗎？是的，我告訴你們，他比先知大多了。
MATT|11|10|這個人就是經上所說的： 『看哪，我要差遣我的使者在你面前， 他要在你前面為你預備道路。』
MATT|11|11|我實在告訴你們，凡女子所生的，沒有一個比施洗 約翰 大；但在天國裏，最小的比他還大。
MATT|11|12|從施洗 約翰 的日子到今天，天國受到強烈的攻擊，強者奪取它 。
MATT|11|13|眾先知和律法，直到 約翰 為止，都說了預言。
MATT|11|14|如果你們願意接受，這人就是那要來的 以利亞 。
MATT|11|15|有耳的，就應當聽！
MATT|11|16|「我該用甚麼來比這世代呢？這正像孩童坐在街市上向同伴呼喊：
MATT|11|17|『我們為你們吹笛，你們不跳舞； 我們唱哀歌，你們不捶胸。』
MATT|11|18|約翰 來了，既不吃也不喝，人們就說他是被鬼附的；
MATT|11|19|人子來了，也吃也喝，他們又說這人貪食好酒，是稅吏和罪人的朋友。而智慧是由它的果子來證實的 。」
MATT|11|20|那時，耶穌在一些城行了許多異能。因為城裏的人不肯悔改，他就責備那些城說：
MATT|11|21|「 哥拉汛 哪，你有禍了！ 伯賽大 啊，你有禍了！因為在你們中間所行的異能若行在 推羅 、 西頓 ，他們早已披麻蒙灰悔改了。
MATT|11|22|但我告訴你們，在審判的日子， 推羅 和 西頓 所受的，比你們還容易受呢！
MATT|11|23|迦百農 啊， 你以為要被舉到天上嗎？ 你要被推下陰間！ 因為在你那裏所行的異能，若行在 所多瑪 ，它還可以存留到今日。
MATT|11|24|但我告訴你們，在審判的日子， 所多瑪 地方所受的，比你們還容易受呢！」
MATT|11|25|那時，耶穌說：「父啊，天地的主，我感謝你！因為你把這些事向聰明智慧的人隱藏起來，而向嬰孩啟示出來。
MATT|11|26|父啊，是的，因為你的美意本是如此。
MATT|11|27|一切都是我父交給我的；除了父，沒有人知道子；除了子和子所願意啟示的人，沒有人知道父。
MATT|11|28|凡勞苦擔重擔的人都到我這裏來，我要使你們得安息。
MATT|11|29|我心裏柔和謙卑，你們當負我的軛，向我學習；這樣，你們的心靈就必得安息。
MATT|11|30|因為我的軛是容易的，我的擔子是輕省的。」
MATT|12|1|那時，耶穌在安息日從麥田經過。他的門徒餓了，就摘麥穗來吃。
MATT|12|2|法利賽人看見，對耶穌說：「看哪，你的門徒在安息日做不合法的事了。」
MATT|12|3|耶穌對他們說：「 大衛 和跟從他的人飢餓時所做的事，你們沒有念過嗎？
MATT|12|4|他怎麼進了上帝的居所，吃了供餅呢？這餅是他和跟從他的人不可以吃的，惟獨祭司才可以吃。
MATT|12|5|再者，律法上所記的，在安息日，祭司在聖殿裏犯了安息日也不算有罪，你們沒有念過嗎？
MATT|12|6|但我告訴你們，比聖殿更大的在這裏。
MATT|12|7|『我喜愛憐憫，不喜愛祭祀。』你們若明白這話的意思，就不將無罪的當作有罪了。
MATT|12|8|因為人子是安息日的主。」
MATT|12|9|耶穌離開那地方，進了 猶太 人的會堂；
MATT|12|10|那裏有個一隻手萎縮了的人。有人為了要控告耶穌，就問他：「安息日治病合不合法？」
MATT|12|11|耶穌對他們說：「你們中間誰有一隻羊在安息日掉在坑裏，不抓住牠，把牠拉上來呢？
MATT|12|12|人比羊貴重得多了！所以，在安息日做善事是合法的。」
MATT|12|13|於是對那人說：「伸出手來！」他把手一伸，手就復原了，和另一隻一樣。
MATT|12|14|法利賽人出去，商議怎樣除掉耶穌。
MATT|12|15|耶穌知道了，就離開那裏，有一大群人跟著他。他把所有的病人都治好了，
MATT|12|16|又囑咐他們不要把他宣揚出去。
MATT|12|17|這是要應驗 以賽亞 先知所說的話：
MATT|12|18|「看哪，我所揀選的僕人， 我所親愛，心所喜悅的； 我要將我的靈賜給他， 他必將公理傳給外邦。
MATT|12|19|他不爭吵，不喧嚷， 街上也沒有人聽見他的聲音。
MATT|12|20|壓傷的蘆葦，他不折斷， 將殘的燈火，他不吹滅， 直到他使公理得勝。
MATT|12|21|外邦人都要仰望他的名。」
MATT|12|22|當時，有人把一個被鬼附，又盲又啞的人帶到耶穌那裏，耶穌醫治他，那啞巴就能說話，又能看見。
MATT|12|23|眾人都驚奇，說：「這不是 大衛 之子嗎？」
MATT|12|24|但法利賽人聽見，就說：「這個人趕鬼，無非是靠著鬼王 別西卜 罷了。」
MATT|12|25|耶穌知道他們的心思，就對他們說：「一國自相紛爭，必定荒蕪；一城一家自相紛爭，必立不住。
MATT|12|26|若撒但趕出撒但，就是自相紛爭，他的國怎能立得住呢？
MATT|12|27|我若靠著 別西卜 趕鬼，你們的子弟趕鬼又靠著誰呢？這樣，他們要作你們的判官。
MATT|12|28|我若靠著上帝的靈趕鬼，那麼，上帝的國就已臨到你們了。
MATT|12|29|人怎能進壯士家裏搶奪他的東西呢？除非先綁住那壯士，否則無法搶奪他的家。
MATT|12|30|不跟我一起的，就是反對我；不與我一起收聚的，就是在拆散。
MATT|12|31|所以我告訴你們，人一切的罪和褻瀆的話都可得赦免，但是褻瀆聖靈，總不得赦免。
MATT|12|32|凡說話干犯人子的，還可得赦免；但是說話干犯聖靈的，今世來世總不得赦免。」
MATT|12|33|「你們知道樹好，果子也好；又知道樹壞，果子也壞；因為看果子就可以知道樹。
MATT|12|34|毒蛇的孽種啊，你們既是惡人，怎能說出好話來呢？因為心裏所充滿的，口裏就說出來。
MATT|12|35|善人從他所存的善發出善來；惡人從他所存的惡發出惡來。
MATT|12|36|我告訴你們，凡是人所說的閒話，在審判的日子，要句句供出來；
MATT|12|37|因為要憑你的話定你為義，也要憑你的話定你有罪。」
MATT|12|38|當時，有幾個文士和法利賽人對耶穌說：「老師，我們想請你顯個神蹟給我們看看。」
MATT|12|39|耶穌回答他們：「邪惡淫亂的世代求看神蹟，除了先知 約拿 的神蹟以外，再沒有神蹟給他們看了。
MATT|12|40|約拿 三日三夜在大魚肚腹中，同樣，人子也要三日三夜在地裏面。
MATT|12|41|在審判的時候， 尼尼微 人要起來定這世代的罪，因為 尼尼微 人聽了 約拿 所傳的就悔改了。看哪，比 約拿 更大的在這裏！
MATT|12|42|在審判的時候，南方的女王要起來定這世代的罪，因為她從地極而來，要聽 所羅門 智慧的話。看哪，比 所羅門 更大的在這裏！」
MATT|12|43|「污靈離了人身，走遍無水之地尋找安歇之處，卻找不到。
MATT|12|44|於是他說：『我要回到我原來的屋裏去。』他到了，看見裏面空著，打掃乾淨，修飾好了，
MATT|12|45|就去另帶了七個比自己更惡的靈來，都進去住在那裏。那人後來的景況比先前更壞了。這邪惡的世代也要如此。」
MATT|12|46|耶穌還在對眾人說話的時候，不料，他母親和他兄弟站在外邊想要跟他說話。
MATT|12|47|有人告訴他：「看哪！你母親和你兄弟站在外邊，想要跟你說話。」
MATT|12|48|他卻回答那對他說話的人，說：「誰是我的母親？誰是我的兄弟？」
MATT|12|49|於是他伸手指著門徒，說：「看哪，我的母親，我的兄弟！
MATT|12|50|凡遵行我天父旨意的人就是我的兄弟、姊妹和母親。」
MATT|13|1|就在那天，耶穌從房子裏出來，坐在海邊。
MATT|13|2|有一大群人到他那裏聚集，他只好上船坐下，眾人都站在岸上。
MATT|13|3|他用比喻對他們講了許多話。他說：「有一個撒種的出去撒種。
MATT|13|4|他撒的時候，有的落在路旁，飛鳥來把它們吃掉了。
MATT|13|5|有的落在土淺的石頭地上，因為土不深，很快就長出苗來，
MATT|13|6|太陽出來一曬，因為沒有根就枯乾了。
MATT|13|7|有的落在荊棘裏，荊棘長起來，把它擠住了。
MATT|13|8|又有的落在好土裏，就結出果實，有一百倍的，有六十倍的，有三十倍的。
MATT|13|9|有耳的，就應當聽！」
MATT|13|10|門徒進前來問耶穌：「對眾人講話，為甚麼用比喻呢？」
MATT|13|11|耶穌回答他們說：「因為天國的奧祕只讓你們知道，不讓他們知道。
MATT|13|12|凡有的，還要給他，讓他有餘；凡沒有的，連他所有的也要奪去。
MATT|13|13|我之所以用比喻對他們講，是因為 他們看卻看不清， 聽卻聽不見，也不明白。
MATT|13|14|在他們身上，正應驗了 以賽亞 的預言： 『你們聽了又聽，卻不明白， 看了又看，卻看不清。
MATT|13|15|因為這百姓的心麻木， 耳朵發沉， 眼睛閉著， 免得眼睛看見， 耳朵聽見， 心裏明白，回轉過來， 我會醫治他們。』
MATT|13|16|但你們的眼睛是有福的，因為看得見；你們的耳朵也是有福的，因為聽得見。
MATT|13|17|我實在告訴你們，從前有許多先知和義人要看你們所看的，卻沒有看見；要聽你們所聽的，卻沒有聽見。」
MATT|13|18|「所以，你們要聽這撒種的比喻。
MATT|13|19|凡聽見天國的道而不明白的，那惡者就來，把撒在他心裏的奪了去；這就是撒在路旁的了。
MATT|13|20|撒在石頭地上的，就是人聽了道，立刻歡喜領受，
MATT|13|21|只因心裏沒有根，不過是暫時的，一旦為道遭受患難或迫害，立刻就跌倒。
MATT|13|22|撒在荊棘裏的，就是人聽了道，後來有世上的憂慮、錢財的迷惑把道擠住了，結不出果實。
MATT|13|23|撒在好土裏的，就是人聽了道，明白了，後來結了果實，有一百倍的，有六十倍的，有三十倍的。」
MATT|13|24|耶穌又設個比喻對他們說：「天國好比人撒好種在田裏，
MATT|13|25|在人睡覺的時候，他的仇敵來，把雜草撒在麥子裏就走了。
MATT|13|26|到長苗吐穗的時候，雜草也顯出來。
MATT|13|27|地主的僕人進前來對他說：『主人，你不是撒好種在田裏嗎？哪裏來的雜草呢？』
MATT|13|28|主人回答他們：『這是仇敵做的。』僕人對他說：『你要我們去拔掉嗎？』
MATT|13|29|主人說：『不必，恐怕拔雜草，也把麥子連根拔出來。
MATT|13|30|讓這兩樣一起長，等到收割。當收割的時候，我會對收割的人說，先把雜草拔出來，捆成捆，留著燒，把麥子收在我的倉裏。』」
MATT|13|31|他又設個比喻對他們說：「天國好比一粒芥菜種，有人拿去種在田裏。
MATT|13|32|它原比所有的種子都小，等到長起來，卻比各樣的菜都大，且成了樹，以致天上的飛鳥來在它的枝上築巢。」
MATT|13|33|他又對他們講另一個比喻：「天國好比麵酵，有婦人拿來放進三斗麵裏，直到全團都發起來。」
MATT|13|34|這都是耶穌用比喻對眾人說的話，不用比喻，他就不對他們說甚麼。
MATT|13|35|這是要應驗先知 所說的話： 「我要開口說比喻， 說出從創世以來所隱藏的事。」
MATT|13|36|當時，耶穌離開眾人，進了屋子。他的門徒進前來，說：「請把田間雜草的比喻講給我們聽。」
MATT|13|37|他回答：「那撒好種的就是人子，
MATT|13|38|田地就是世界，好種就是天國之子，雜草就是那惡者之子，
MATT|13|39|撒雜草的仇敵就是魔鬼，收割的時候就是世代的終結，收割的人就是天使。
MATT|13|40|正如把雜草拔出來用火焚燒，世代的終結也要如此。
MATT|13|41|人子要差遣他的使者，把一切使人跌倒的和作惡的從他國裏挑出來，
MATT|13|42|丟在火爐裏，在那裏要哀哭切齒了。
MATT|13|43|那時，義人要在他們父的國裏發出光來，像太陽一樣。有耳的，就應當聽！」
MATT|13|44|「天國好比寶貝藏在地裏，人發現了就把它藏起來，歡歡喜喜地去變賣一切所有的，買這塊地。
MATT|13|45|「天國又好比商人尋找好的珍珠，
MATT|13|46|發現一顆貴重的珍珠，就去變賣他一切所有的，買下這顆珍珠。」
MATT|13|47|「天國又好比網撒在海裏，聚攏各種魚類，
MATT|13|48|網一滿，人們就把它拉上岸，坐下來，揀好的收在桶裏，不好的丟掉。
MATT|13|49|世代的終結也要這樣：天使要出來，把惡人從義人中分別出來，
MATT|13|50|丟在火爐裏，在那裏要哀哭切齒了。」
MATT|13|51|耶穌說：「這一切的話你們都明白了嗎？」他們對他說：「明白了。」
MATT|13|52|他對他們說：「凡文士學習作天國的門徒，就像一個家的主人從他庫裏拿出新的和舊的東西來。」
MATT|13|53|耶穌說完了這些比喻，就離開那裏，
MATT|13|54|來到自己的家鄉，在會堂裏教導人，以致他們都很驚奇，說：「這人哪來這樣的智慧和異能呢？
MATT|13|55|這不是那木匠的兒子嗎？他母親不是叫 馬利亞 嗎？他兄弟們不是叫 雅各 、 約瑟 、 西門 、 猶大 嗎？
MATT|13|56|他姊妹們不是都在我們這裏嗎？他這一切是從哪裏來的呢？」
MATT|13|57|他們就厭棄他。耶穌對他們說：「先知除了在本鄉和自己的家之外，沒有不被尊敬的。」
MATT|13|58|耶穌因為他們不信，沒有在那裏行很多異能。
MATT|14|1|那時， 希律 分封王聽見耶穌的名聲，
MATT|14|2|就對臣僕說：「這是施洗的 約翰 從死人中復活，因此才有這些異能在他裏面運行。」
MATT|14|3|原來， 希律 為他兄弟 腓力 的妻子 希羅底 的緣故，把 約翰 抓住綁了，關進監獄，
MATT|14|4|因為 約翰 曾對他說：「你佔有這婦人是不合法的。」
MATT|14|5|希律 就想要殺他，可是怕民眾，因為他們認為 約翰 是先知。
MATT|14|6|到了 希律 的生日， 希羅底 的女兒在眾人面前跳舞，使 希律 歡喜，
MATT|14|7|於是 希律 發誓許諾隨她所求的給她。
MATT|14|8|女兒被母親指使，就說：「請把施洗 約翰 的頭放在盤子裏，拿來給我。」
MATT|14|9|王就憂愁，然而因他所發的誓，又因同席的人，就下令給她；
MATT|14|10|於是打發人去，在監獄裏斬了 約翰 ，
MATT|14|11|把頭放在盤子裏，拿來給那女孩，她拿去給她母親。
MATT|14|12|約翰 的門徒來，把屍體領去埋葬了，又去告訴耶穌。
MATT|14|13|耶穌聽到了，就從那裏上船，私下退到荒野的地方去。眾人聽到後，從各城來，步行跟隨他。
MATT|14|14|耶穌出來，見有一大群人，就憐憫他們，治好了他們的病人。
MATT|14|15|傍晚的時候，門徒進前來，說：「這地方偏僻，而且時候已經晚了，請叫眾人散去，他們好進村子，自己買些食物。」
MATT|14|16|耶穌對他們說：「不用他們去，你們給他們吃吧！」
MATT|14|17|門徒說：「我們這裏只有五個餅、兩條魚。」
MATT|14|18|耶穌說：「拿過來給我。」
MATT|14|19|於是他吩咐眾人坐在草地上，就拿著這五個餅和兩條魚，望著天祝福，擘開餅，遞給門徒，門徒又遞給眾人。
MATT|14|20|他們都吃，並且吃飽了。門徒把剩下的碎屑收拾起來，裝滿了十二個籃子。
MATT|14|21|吃的人中，男的約有五千，還不算婦女和孩子。
MATT|14|22|耶穌隨即催門徒上船，先渡到對岸，等他叫眾人散去。
MATT|14|23|疏散了眾人以後，他獨自上山去禱告。到了晚上，只有他一人在那裏。
MATT|14|24|那時船已離岸好幾里 ，因風不順，被浪顛簸。
MATT|14|25|天快亮的時候，耶穌在海面上走，往門徒那裏去。
MATT|14|26|但門徒看見他在海面上走，就驚慌了，說：「是個鬼怪！」他們害怕得喊叫起來。
MATT|14|27|耶穌連忙對他們說：「放心！是我，不要怕！」
MATT|14|28|彼得 回答他說：「主啊，如果是你，請叫我從水面上走到你那裏去。」
MATT|14|29|耶穌說：「你來吧！」 彼得 就從船上下去，在水面上走，往耶穌那裏去；
MATT|14|30|只因見風很強 ，害怕起來，將要沉下去，就喊著說：「主啊，救我！」
MATT|14|31|耶穌立刻伸手拉住他，說：「你這小信的人哪，為甚麼疑惑呢？」
MATT|14|32|他們一上船，風就停了。
MATT|14|33|在船上的人都拜他，說：「你真是上帝的兒子。」
MATT|14|34|他們渡過了海，在 革尼撒勒 上岸。
MATT|14|35|那裏的人認出耶穌，就打發人到整個周圍地區去，把所有的病人帶到他那裏，
MATT|14|36|求耶穌讓他們只摸一摸他的衣裳繸子，摸著的人就都好了。
MATT|15|1|那時，有法利賽人和文士從 耶路撒冷 來見耶穌，說：
MATT|15|2|「你的門徒為甚麼違反古人的傳統？因為他們吃飯的時候不洗手。」
MATT|15|3|耶穌回答他們：「你們為甚麼因你們的傳統而違反上帝的誡命呢？
MATT|15|4|上帝說：『當孝敬父母』；又說：『咒罵父母的，必須處死。』
MATT|15|5|你們倒說：『無論誰對父母說：我所當供奉你的已經作了奉獻，
MATT|15|6|就可以不孝敬他的父親 。』這就是你們藉著傳統，廢了上帝的話。
MATT|15|7|假冒為善的人哪！ 以賽亞 指著你們所預言的說得好：
MATT|15|8|『這百姓用嘴唇尊敬我， 他們的心卻遠離我。
MATT|15|9|他們把人的規條當作教義教導人； 他們拜我也是枉然。』」
MATT|15|10|耶穌叫了眾人來，對他們說：「你們要聽，也要明白。
MATT|15|11|從口裏進去的不玷污人，從口裏出來的才玷污人。」
MATT|15|12|當時，門徒進前來對他說：「法利賽人聽見這話很反感，你知道嗎？」
MATT|15|13|耶穌回答：「一切植物，若不是我天父栽植的，都要連根拔出來。
MATT|15|14|由他們吧！他們是瞎子作瞎子的嚮導 ；若是瞎子領瞎子，兩個人都要掉在坑裏。」
MATT|15|15|彼得 回應他說：「請將這比喻講解給我們聽。」
MATT|15|16|耶穌說：「連你們也還不明白嗎？
MATT|15|17|難道你們不了解，凡進到口裏的，是經過肚子，又排入廁所嗎？
MATT|15|18|然而口裏出來的是出於心裏，這才玷污人。
MATT|15|19|因為出於心裏的有種種惡念，如兇殺、姦淫、淫亂、偷盜、偽證、毀謗。
MATT|15|20|這些才玷污人。至於不洗手吃飯，那並不玷污人。」
MATT|15|21|耶穌離開那裏，退到 推羅 、 西頓 境內。
MATT|15|22|有一個 迦南 婦人從那地方出來，喊著說：「主啊， 大衛 之子，可憐我！我女兒被鬼纏得很苦。」
MATT|15|23|耶穌卻一言不答。門徒進前來，求他說：「這婦人在我們後頭喊叫，請打發她走吧。」
MATT|15|24|耶穌回答：「我奉差遣只到 以色列 家迷失的羊那裏去。」
MATT|15|25|那婦人來拜他，說：「主啊，幫幫我！」
MATT|15|26|他回答：「拿孩子的餅丟給小狗吃是不妥的。」
MATT|15|27|婦人說：「主啊，不錯，可是小狗也吃牠主人桌上掉下來的碎屑。」
MATT|15|28|於是耶穌回答她說：「婦人，你的信心很大！照你所要的成全你吧。」從那時起，她的女兒就好了。
MATT|15|29|耶穌離開那地方，來到靠近 加利利 的海邊，就上山坐下。
MATT|15|30|有一大群人到他那裏，帶著瘸子、盲人、肢殘的、聾啞的，和好些別的病人，都放在他腳前，他就治好了他們。
MATT|15|31|於是眾人都驚訝，因為看見聾啞的說話，肢殘的痊癒，瘸子行走，盲人看見，他們就歸榮耀給 以色列 的上帝。
MATT|15|32|耶穌叫門徒來，說：「我憐憫這群人，因為他們同我在這裏已經三天，沒有吃的東西了。我不願意叫他們餓著回去，恐怕他們在路上餓昏了。」
MATT|15|33|門徒說：「我們在這野地，哪裏有這麼多的餅讓這許多人吃飽呢？」
MATT|15|34|耶穌對他們說：「你們有多少餅？」他們說：「有七個，還有幾條小魚。」
MATT|15|35|他就吩咐眾人坐在地上，
MATT|15|36|拿著這七個餅和幾條魚，祝謝了，擘開，遞給門徒；門徒又遞給眾人。
MATT|15|37|他們都吃，並且吃飽了，收拾剩下的碎屑，裝滿了七個筐子。
MATT|15|38|吃的人中，男的有四千，還不算婦女和孩子。
MATT|15|39|耶穌叫眾人散去，就上船，來到 馬加丹 境內。
MATT|16|1|法利賽人和撒都該人來試探耶穌，請他顯個來自天上的神蹟給他們看。
MATT|16|2|耶穌回答他們：「傍晚天發紅，你們就說：『明日天晴。』
MATT|16|3|早晨天色又紅又暗，你們就說：『今日有風雨。』你們知道分辨天上的氣象，倒不能分辨這個時代的神蹟 。
MATT|16|4|邪惡淫亂的世代求看神蹟，除了 約拿 的神蹟以外，再沒有神蹟給他們看了。」於是耶穌離開他們走了。
MATT|16|5|門徒渡到對岸，忘了帶餅。
MATT|16|6|耶穌對他們說：「你們要謹慎，要防備法利賽人和撒都該人的酵。」
MATT|16|7|門徒彼此議論說：「這是因為我們沒有帶餅吧。」
MATT|16|8|耶穌知道了，就說：「你們這小信的人，為甚麼因為沒有餅就彼此議論呢？
MATT|16|9|你們還不明白嗎？不記得那五個餅分給五千人，你們收拾了多少籃子的碎屑嗎？
MATT|16|10|也不記得那七個餅分給四千人，你們又收拾了多少筐子的碎屑嗎？
MATT|16|11|我對你們說『要防備法利賽人和撒都該人的酵』，這話不是指著餅說的，你們怎麼不明白呢？」
MATT|16|12|門徒這才明白他所說的不是要他們防備餅的酵 ，而是要防備法利賽人和撒都該人的教訓。
MATT|16|13|耶穌到了 凱撒利亞．腓立比 的境內，就問門徒：「人們說人子是誰？」
MATT|16|14|他們說：「有人說是施洗的 約翰 ；有人說是 以利亞 ；又有人說是 耶利米 或是先知中的一位。」
MATT|16|15|耶穌問他們：「你們說我是誰？」
MATT|16|16|西門．彼得 回答說：「你是基督，是永生上帝的兒子。」
MATT|16|17|耶穌回答他說：「 約拿 的兒子 西門 ，你是有福的！因為這不是屬血肉的啟示你的，而是我在天上的父啟示的。
MATT|16|18|我還告訴你，你是 彼得 ，我要把我的教會建造在這磐石上，陰間的權柄不能勝過它。
MATT|16|19|我要把天國的鑰匙給你，凡你在地上所捆綁的，在天上也要捆綁；凡你在地上所釋放的，在天上也要釋放。」
MATT|16|20|當時，耶穌囑咐門徒不可對任何人說他是基督。
MATT|16|21|從那時起，耶穌才向門徒明說，他必須上 耶路撒冷 去，受長老、祭司長和文士許多的苦，並且被殺，第三天復活。
MATT|16|22|彼得 就拉著他，責備他說：「主啊，千萬不可如此！這事絕不可臨到你身上。」
MATT|16|23|耶穌轉過來，對 彼得 說：「撒但，退到我後邊去！你是我的絆腳石，因為你不體會上帝的心意，而是體會人的意思。」
MATT|16|24|於是耶穌對門徒說：「若有人要跟從我，就當捨己，背起自己的十字架來跟從我。
MATT|16|25|因為凡要救自己生命的，要喪失生命；凡為我喪失生命的，要得著生命。
MATT|16|26|人若賺得全世界，賠上自己的生命，有甚麼益處呢？人還能拿甚麼換生命呢？
MATT|16|27|人子要在他父的榮耀裏與他的眾使者一起來臨，那時候，他要照各人的行為報應各人。
MATT|16|28|我實在告訴你們，站在這裏的，有人在沒經歷死亡以前，必定看見人子來到他的國裏。」
MATT|17|1|過了六天，耶穌帶著 彼得 、 雅各 和 雅各 的弟弟 約翰 ，領他們悄悄地上了高山。
MATT|17|2|他在他們面前變了形像，他的臉明亮如太陽，衣裳潔白如光。
MATT|17|3|忽然，有 摩西 和 以利亞 向他們顯現，與耶穌說話。
MATT|17|4|彼得 回應，對耶穌說：「主啊，我們在這裏真好！你若願意，我就在這裏搭三座棚，一座為你，一座為 摩西 ，一座為 以利亞 。」
MATT|17|5|說話之間，忽然有一朵明亮的雲彩遮蓋他們，又有聲音從雲彩裏出來，說：「這是我的愛子，我所喜愛的。你們要聽從他！」
MATT|17|6|門徒聽見，就俯伏在地，極其害怕。
MATT|17|7|耶穌進前來，拍拍他們，說：「起來，不要害怕！」
MATT|17|8|他們舉目，不見一人，只見耶穌獨自一人。
MATT|17|9|下山的時候，耶穌囑咐他們說：「人子還沒有從死人中復活，你們不要把所看到的告訴人。」
MATT|17|10|門徒問耶穌：「那麼，文士為甚麼說 以利亞 必須先來？」
MATT|17|11|耶穌回答：「 以利亞 的確要來，並要復興萬事；
MATT|17|12|可是我告訴你們， 以利亞 已經來了，人不認識他，反倒任意待他。人子也將這樣受他們的苦。」
MATT|17|13|門徒這才明白耶穌所說的是指施洗的 約翰 。
MATT|17|14|耶穌和門徒到了眾人那裏，有一個人來見耶穌，跪下，
MATT|17|15|說：「主啊，可憐我的兒子。他害癲癇病很苦，屢次跌進火裏，屢次跌進水裏。
MATT|17|16|我帶他到你門徒那裏，他們卻不能醫治他。」
MATT|17|17|耶穌回答：「唉！這又不信又悖謬的世代啊，我和你們在一起要到幾時呢？我忍耐你們要到幾時呢？把他帶到我這裏來！」
MATT|17|18|耶穌斥責那鬼，鬼就出來；從那時起，孩子就痊癒了。
MATT|17|19|門徒私下進前來問耶穌：「我們為甚麼不能趕出那鬼呢？」
MATT|17|20|耶穌對他們說：「是因你們的信心小。我實在告訴你們，你們若有信心像一粒芥菜種，就是對這座山說：『你從這邊移到那邊』，它也會移過去，並且你們沒有一件不能做的事了。 」
MATT|17|21|
MATT|17|22|他們聚集在 加利利 的時候，耶穌對門徒說：「人子將要被交在人手裏。
MATT|17|23|他們要殺害他，第三天他要復活。」門徒就非常憂愁。
MATT|17|24|他們到了 迦百農 ，收聖殿稅 的人來見 彼得 ，說：「你們的老師不納聖殿稅嗎？」
MATT|17|25|彼得 說：「納。」他進了屋子，耶穌先對他說：「 西門 ，你的意見如何？世上的君王向誰徵收關稅或丁稅？是向自己的兒子呢？還是向外人呢？」
MATT|17|26|彼得 說：「是向外人。」耶穌對他說：「既然如此，兒子就可以免了。
MATT|17|27|但恐怕觸犯他們，你往海邊去釣魚，把先釣上來的魚拿起來，開了牠的口，會發現一個司塔特 ，可以拿去給他們，作你我的稅錢。」
MATT|18|1|當時，門徒前來問耶穌：「天國裏誰是最大的？」
MATT|18|2|耶穌叫一個小孩子來，讓他站在他們當中，
MATT|18|3|說：「我實在告訴你們，你們若不回轉，變成像小孩子一樣，絕不能進天國。
MATT|18|4|所以，凡自己謙卑像這小孩子的，他在天國裏就是最大的。
MATT|18|5|凡為我的名接納一個像這小孩子的，就是接納我。」
MATT|18|6|「凡使這些信我的小子中的一個跌倒的，倒不如把大磨石拴在這人的頸項上，沉在深海裏。
MATT|18|7|這世界有禍了，因為它使人跌倒；絆倒人的事是免不了的，但那絆倒人的有禍了！
MATT|18|8|如果你一隻手或是一隻腳使你跌倒，就把它砍下來扔掉。你缺一隻手或是一隻腳進入永生，比有兩手兩腳被扔進永火裏還好。
MATT|18|9|如果你一隻眼使你跌倒，就把它挖出來扔掉。你只有一隻眼進入永生，比有兩隻眼被扔進地獄的火裏還好。」
MATT|18|10|「你們要小心，不可輕看這些小子中的一個；我告訴你們，他們的天使在天上，常見我天父的面。
MATT|18|11|
MATT|18|12|「一個人若有一百隻羊，其中一隻走迷了路，你們的意見如何？他豈不留下這九十九隻在山上，去找那隻迷路的羊嗎？
MATT|18|13|若是找到了，我實在告訴你們，他為這一隻羊歡喜，比為那沒有迷路的九十九隻歡喜還大呢！
MATT|18|14|你們 在天上的父也是這樣，不願意失去這些小子中的一個。」
MATT|18|15|「若是你的弟兄得罪你 ，你要去，趁著只有他和你在一起的時候，指出他的錯來。他若聽你，你就贏得了你的弟兄；
MATT|18|16|他若不聽，你就另外帶一個或兩個人同去，因為『任何指控都要憑兩個或三個證人的口述才能成立』。
MATT|18|17|他若是不聽他們，就去告訴教會；若是不聽教會，就把他看作外邦人和稅吏。
MATT|18|18|「我實在告訴你們，凡你們在地上所捆綁的，在天上也要捆綁；凡你們在地上所釋放的，在天上也要釋放。
MATT|18|19|我又實在 告訴你們，若是你們中間有兩個人在地上同心合意地求甚麼事，我在天上的父必為他們成全。
MATT|18|20|因為，哪裏有兩三個人奉我的名聚會，哪裏就有我在他們中間。」
MATT|18|21|那時， 彼得 進前來，對耶穌說：「主啊，我弟兄得罪我，我當饒恕他幾次呢？到七次夠嗎？」
MATT|18|22|耶穌說：「我告訴你，不是到七次，而是到七十個七次。
MATT|18|23|因為天國好像一個王要和他僕人算賬。
MATT|18|24|他開始算的時候，有人帶了一個欠一萬他連得的僕人來。
MATT|18|25|因為他沒有甚麼償還之物，主人下令把他和他妻子兒女，以及一切所有的都賣了來償還。
MATT|18|26|那僕人就俯伏向他叩頭，說：『寬容我吧，我都會還你的。』
MATT|18|27|那僕人的主人就動了慈心，把他釋放了，並且免了他的債。
MATT|18|28|那僕人出來，遇見一個欠他一百個銀幣的同伴，就揪著他，扼住他的喉嚨，說：『把你所欠的還我！』
MATT|18|29|他的同伴就俯伏央求他，說：『寬容我吧，我會還你的。』
MATT|18|30|他不肯，卻把他下在監裏，直到他還了所欠的債。
MATT|18|31|同伴們看見他所做的事就很悲憤，把這一切的事都告訴了主人。
MATT|18|32|於是主人叫了他來，對他說：『你這惡奴才！你央求我，我就把你所欠的都免了；
MATT|18|33|你不應該憐憫你的同伴，像我憐憫你嗎？』
MATT|18|34|主人就大怒，把他交給司刑的，直到他還清了所欠的債。
MATT|18|35|你們各人若不從心裏饒恕你的弟兄，我天父也要這樣待你們。」
MATT|19|1|耶穌說完了這些話，就離開 加利利 ，來到 猶太 的境內、 約旦河 的東邊。
MATT|19|2|有一大群人跟著他，他就在那裏治好了他們。
MATT|19|3|有些法利賽人來試探耶穌說：「無論甚麼緣故，人休妻都合法嗎？」
MATT|19|4|耶穌回答：「那起初造人的，是造男造女，並且說：『因此，人要離開父母，與妻子結合，二人成為一體。』這經文你們沒有念過嗎？
MATT|19|5|
MATT|19|6|既然如此，夫妻不再是兩個人，而是一體的了。所以，上帝配合的，人不可分開。」
MATT|19|7|法利賽人說：「這樣， 摩西 為甚麼吩咐給妻子休書就可以休她呢？」
MATT|19|8|耶穌說：「 摩西 因為你們的心硬，所以准許你們休妻，但起初並不是這樣。
MATT|19|9|我告訴你們，凡休妻另娶的，若不是為不貞的緣故，就是犯姦淫了。 」
MATT|19|10|門徒對耶穌說：「丈夫和妻子的關係既是這樣，倒不如不娶。」
MATT|19|11|耶穌對他們說：「這話不是人人都能領受的，惟獨賜給誰，誰才能領受。
MATT|19|12|因為有人從母腹裏就是不宜結婚的，也有因人為的緣故不宜結婚的，並有為天國的緣故自己不結婚的 。這話誰能領受，就領受吧。」
MATT|19|13|那時，有人帶著小孩子來見耶穌，要他給他們按手禱告，門徒就責備那些人。
MATT|19|14|耶穌說：「讓小孩子到我這裏來，不要阻止他們，因為在天國的正是這樣的人。」
MATT|19|15|耶穌給他們按手，然後離開那地方。
MATT|19|16|有一個人進前來問耶穌：「老師，我該做甚麼善事才能得永生？」
MATT|19|17|耶穌對他說：「你為甚麼問我關於善的事呢？只有一位是善良的。你若要進入永生，就該遵守誡命。」
MATT|19|18|他說：「哪些誡命？」耶穌說：「就是不可殺人；不可姦淫；不可偷盜；不可作假見證；
MATT|19|19|當孝敬父母；又當愛鄰 如己。」
MATT|19|20|那青年說：「這一切我都遵守了，還缺少甚麼呢？」
MATT|19|21|耶穌說：「你若願意作完全人，去變賣你所擁有的，分給窮人，就必有財寶在天上；然後來跟從我。」
MATT|19|22|那青年聽見這話，就憂憂愁愁地走了，因為他的產業很多。
MATT|19|23|耶穌對門徒說：「我實在告訴你們，財主進天國是難的。
MATT|19|24|我再告訴你們，駱駝穿過針眼比財主進上帝的國還容易呢！」
MATT|19|25|門徒聽見這話，就非常驚奇，說：「這樣，誰能得救呢？」
MATT|19|26|耶穌看著他們，說：「在人這是不能，在上帝凡事都能。」
MATT|19|27|於是 彼得 回應，對他說：「看哪，我們已經撇下一切跟從你了，我們會得到甚麼呢？」
MATT|19|28|耶穌對他們說：「我實在告訴你們，你們這些跟從我的人，到了萬物更新、人子坐在他榮耀寶座上的時候，你們也要坐在十二個寶座上，審判 以色列 十二個支派。
MATT|19|29|凡為我的名撇下房屋，或是兄弟、姊妹、父親、母親、 兒女、田地的，將得著百倍，並且承受永生。
MATT|19|30|然而，有許多在前的，將要在後；在後的，將要在前。」
MATT|20|1|「因為天國好比一家的主人清早去雇人進他的葡萄園做工。
MATT|20|2|他和工人講定一天一個銀幣 ，就打發他們進葡萄園去。
MATT|20|3|約在上午九點鐘出去，看見市場上還有閒站的人，
MATT|20|4|就對那些人說：『你們也進葡萄園去，我會給你們合理的工錢。』
MATT|20|5|他們也進去了。約在正午和下午三點鐘又出去，他也是這麼做。
MATT|20|6|約在下午五點鐘出去，他看見還有人站在那裏，就問他們：『你們為甚麼整天在這裏閒站呢？』
MATT|20|7|他們說：『因為沒有人雇我們。』他說：『你們也進葡萄園去。』
MATT|20|8|到了晚上，園主對工頭說：『叫工人都來，給他們工錢，從後來的起，到先來的為止。』
MATT|20|9|約在下午五點鐘雇的人來了，各人領了一個銀幣。
MATT|20|10|那些最先雇的來了，以為可以多領，誰知也是各領一個銀幣。
MATT|20|11|他們領了工錢，就埋怨那家的主人說：
MATT|20|12|『我們整天勞苦受熱，那些後來的只做了一小時，你竟待他們和我們一樣嗎？』
MATT|20|13|主人回答其中的一人說：『朋友，我沒虧待你，你與我講定的不是一個銀幣嗎？
MATT|20|14|拿你的錢走吧！我樂意給那後來的和給你的一樣，
MATT|20|15|難道我的東西不可隨我的意思用嗎？因為我作好人，你就眼紅了嗎？』
MATT|20|16|這樣，那在後的，將要在前；在前的，將要在後了。」
MATT|20|17|耶穌上 耶路撒冷 去的時候，在路上把十二個門徒帶到一邊，對他們說：
MATT|20|18|「看哪，我們上 耶路撒冷 去，人子將被交給祭司長和文士；他們要定他死罪，
MATT|20|19|把他交給外邦人戲弄，鞭打，釘在十字架上；第三天他要復活。」
MATT|20|20|那時， 西庇太 兒子的母親和她兩個兒子上前來，向耶穌叩頭，求他一件事。
MATT|20|21|耶穌問她：「你要甚麼呢？」她對耶穌說：「在你的國裏，請讓我這兩個兒子一個坐在你右邊，一個坐在你左邊。」
MATT|20|22|耶穌回答：「你們不知道所求的是甚麼。我將要喝的杯，你們能喝嗎？」他們對他說：「我們能。」
MATT|20|23|耶穌說：「我所喝的杯，你們要喝。可是坐在我的左右，不是我可以賜的，而是我父為誰預備就賜給誰。」
MATT|20|24|其餘十個門徒聽見，就對他們兄弟二人很生氣。
MATT|20|25|耶穌叫了他們來，說：「你們知道，外邦人有君王作主治理他們，有大臣操權管轄他們。
MATT|20|26|但是在你們中間，不可這樣。你們中間誰願為大，就要作你們的用人；
MATT|20|27|誰願為首，就要作你們的僕人。
MATT|20|28|正如人子來，不是要受人的服事，乃是要服事人，並且要捨命，作多人的贖價。」
MATT|20|29|他們出 耶利哥 的時候，有一大群人跟隨耶穌。
MATT|20|30|有兩個盲人坐在路旁，聽說是耶穌經過，就喊著說：「主啊 ， 大衛 之子，可憐我們吧！」
MATT|20|31|眾人責備他們，不許他們作聲，他們卻越發喊著說：「主啊 ， 大衛 之子，可憐我們吧！」
MATT|20|32|耶穌就站住，叫他們來，說：「你們要我為你們做甚麼？」
MATT|20|33|他們說：「主啊，讓我們的眼睛能看見。」
MATT|20|34|耶穌動了慈心，摸了他們的眼睛，他們立刻看得見，就跟從耶穌。
MATT|21|1|耶穌和門徒快到 耶路撒冷 ，進了 橄欖山 的 伯法其 時，打發兩個門徒，
MATT|21|2|對他們說：「你們往對面村子裏去，會立刻看見一匹驢拴在那裏，還有驢駒同在一處，解開牠們，牽到我這裏來。
MATT|21|3|若有人對你們說甚麼，你們就說：『主要用牠們。』那人會立刻讓你們牽來。」
MATT|21|4|這事發生是要應驗先知所說的話：
MATT|21|5|「要對 錫安 的兒女 說： 看哪，你的王來到你這裏， 謙和地騎著驢， 騎著小驢—驢的駒子。」
MATT|21|6|門徒就照耶穌所吩咐的去做，
MATT|21|7|牽了驢和驢駒來，把他們的衣服搭在上面，耶穌就騎上。
MATT|21|8|許許多多的人把自己的衣服鋪在路上，還有人砍下樹枝來鋪在路上。
MATT|21|9|前呼後擁的人群喊著說： 「和散那 歸於 大衛 之子！ 奉主名來的是應當稱頌的！ 至高無上的，和散那！」
MATT|21|10|耶穌進了 耶路撒冷 ，全城都驚動了，說：「這是誰？」
MATT|21|11|眾人說：「這是從 加利利 的 拿撒勒 來的先知耶穌。」
MATT|21|12|耶穌進了聖殿 ，趕出聖殿裏所有在做買賣的人，推倒兌換銀錢之人的桌子和賣鴿子之人的凳子，
MATT|21|13|對他們說：「經上記著： 『我的殿要稱為禱告的殿， 你們倒使它成為賊窩了。』」
MATT|21|14|在聖殿裏有盲人和瘸子到耶穌跟前，他就治好了他們。
MATT|21|15|祭司長和文士看見耶穌所行的奇事，又見小孩子在聖殿裏喊著說：「和散那歸於 大衛 之子！」就很生氣，
MATT|21|16|對他說：「這些人所喊的，你聽到了嗎？」耶穌對他們說：「聽到了。經上說：『你藉孩童和吃奶的口發出完全的讚美』，你們沒有念過嗎？」
MATT|21|17|於是他離開他們，出城到 伯大尼 去，在那裏過夜。
MATT|21|18|早晨回城的時候，他餓了，
MATT|21|19|看見路旁有一棵無花果樹，就走到跟前，在樹上找不到甚麼，只有葉子，就對樹說：「從今以後，你永不結果子！」那無花果樹立刻枯乾了。
MATT|21|20|門徒看見了，驚訝地說：「無花果樹怎麼立刻枯乾了呢？」
MATT|21|21|耶穌回答他們：「我實在告訴你們，你們若有信心，不疑惑，不但能行我對無花果樹所行的事，就是對這座山說：『離開此地，投在海裏！』也會實現。
MATT|21|22|你們禱告，無論求甚麼，只要信，就必得著。」
MATT|21|23|耶穌進了聖殿，正教導人的時候，祭司長和百姓的長老來問他：「你仗著甚麼權柄做這些事？給你這權柄的是誰呢？」
MATT|21|24|耶穌回答他們說：「我也要問你們一句話，你們若告訴我，我就告訴你們我仗著甚麼權柄做這些事。
MATT|21|25|約翰 的洗禮是從哪裏來的？是從天上來的，還是從人間來的呢？」他們彼此商議說：「我們若說『從天上來的』，他會對我們說：『這樣，你們為甚麼不信他呢？』
MATT|21|26|若說『從人間來的』，我們又怕眾人，因為大家都認為 約翰 是先知。」
MATT|21|27|於是他們回答耶穌：「我們不知道。」耶穌也對他們說：「我也不告訴你們，我仗著甚麼權柄做這些事。」
MATT|21|28|「有一件事，你們的意見如何？一個人有兩個兒子。他來對大兒子說：『孩子，今天到葡萄園裏做工去。』
MATT|21|29|他回答：『我不去』，以後自己懊悔，就去了。
MATT|21|30|他來對小兒子也是這樣說。他回答：『父親大人，我去』，卻不去。
MATT|21|31|這兩個兒子是哪一個照著父親的意願做了呢？」他們說：「大兒子。」耶穌說：「我實在告訴你們，稅吏和娼妓倒比你們先進上帝的國。
MATT|21|32|因為 約翰 到你們這裏來指引你們走義路，你們卻不信他，稅吏和娼妓倒信了他。你們看見了以後，還是不悔悟去信他。」
MATT|21|33|「你們再聽一個比喻：有一個家的主人開墾了一個葡萄園，四周圍上籬笆，裏面挖了一個榨酒池，蓋了一座守望樓，租給園戶，就出外遠行去了。
MATT|21|34|收果子的時候快到了，他打發僕人到園戶那裏去收果子。
MATT|21|35|園戶拿住僕人，打了一個，殺了一個，用石頭打死了一個。
MATT|21|36|主人又打發別的僕人去，比先前更多；園戶還是照樣對待他們。
MATT|21|37|最後他打發自己的兒子到他們那裏去，說：『他們會尊敬我的兒子。』
MATT|21|38|可是，園戶看見他兒子，彼此說：『這是承受產業的。來，我們殺了他，佔他的產業！』
MATT|21|39|於是他們拿住他，把他扔出葡萄園外，殺了。
MATT|21|40|葡萄園的主人來的時候，要怎樣處置那些園戶呢？」
MATT|21|41|他們說：「要狠狠地除滅那些惡人，將葡萄園轉租給那些按時候交果子的園戶。」
MATT|21|42|耶穌對他們說： 「『匠人所丟棄的石頭 已作了房角的頭塊石頭。 這是主所做的， 在我們眼中看為奇妙。』 這段經文你們從來沒有念過嗎？
MATT|21|43|所以我告訴你們，上帝的國必從你們奪去，賜給那能結果子的民。
MATT|21|44|誰跌在這石頭上，一定會跌得粉碎；這石頭掉在誰的身上，就要把誰壓得稀爛。 」
MATT|21|45|祭司長和法利賽人聽見他的比喻，就看出他是指著他們說的。
MATT|21|46|他們想要捉拿他，但是懼怕眾人，因為眾人認為他是先知。
MATT|22|1|耶穌又用比喻對他們說：
MATT|22|2|「天國好比一個王為他兒子擺設娶親的宴席。
MATT|22|3|他打發僕人去，請那些被邀的人來赴宴，他們卻不肯來。
MATT|22|4|王又打發別的僕人，說：『你們去告訴那被邀的人，我的宴席已經預備好了，牛和肥畜已經宰了，各樣都齊備，請你們來赴宴。』
MATT|22|5|那些人不理就走了，一個到自己田裏去，一個做買賣去。
MATT|22|6|其餘的抓住僕人，凌辱他們，把他們殺了。
MATT|22|7|王就大怒，發兵除滅那些兇手，燒燬他們的城。
MATT|22|8|於是王對僕人說：『喜宴已經齊備，只是所邀的人不配。
MATT|22|9|所以你們要往岔路口上去，凡遇見的，都邀來赴宴。』
MATT|22|10|那些僕人就出去，到大路上，凡遇見的，不論善惡都招聚了來，宴席上就坐滿了客人。
MATT|22|11|王進來見賓客，看到那裏有一個沒有穿禮服的，
MATT|22|12|就對他說：『朋友，你到這裏來怎麼不穿禮服呢？』那人無言可答。
MATT|22|13|於是王對侍從說：『捆起他的手腳，把他扔在外邊的黑暗裏；在那裏他要哀哭切齒了。』
MATT|22|14|因為被召的人多，選上的人少。」
MATT|22|15|於是，法利賽人出去商議，怎樣找話柄來陷害耶穌，
MATT|22|16|就打發他們的門徒同 希律 黨人去見耶穌，說：「老師，我們知道你是誠實的，並且誠誠實實傳上帝的道，無論誰你都一視同仁，因為你不看人的面子。
MATT|22|17|請告訴我們，你的意見如何？納稅給凱撒合不合法？」
MATT|22|18|耶穌看出他們的惡意，就說：「假冒為善的人哪，為甚麼試探我？
MATT|22|19|拿一個納稅的錢給我看！」他們就拿一個銀幣來給他。
MATT|22|20|耶穌問他們：「這像和這名號是誰的？」
MATT|22|21|他們說：「是凱撒的。」於是耶穌說：「這樣，凱撒的歸凱撒；上帝的歸上帝。」
MATT|22|22|他們聽了十分驚訝，就離開他走了。
MATT|22|23|那天，撒都該人來見耶穌。他們說沒有復活這回事，於是問耶穌：
MATT|22|24|「老師， 摩西 說：『某人若死了，沒有孩子，他弟弟該娶他的妻子，為哥哥生子立後。』
MATT|22|25|從前，在我們這裏有兄弟七人，第一個娶了妻，死了，沒有孩子，撇下妻子給弟弟。
MATT|22|26|第二、第三，直到第七個，都是如此。
MATT|22|27|後來，那婦人也死了。
MATT|22|28|那麼，在復活的時候，她是七個人中哪一個的妻子呢？因為他們都娶過她。」
MATT|22|29|耶穌回答他們說：「你們錯了，因為不明白聖經，也不知道上帝的大能。
MATT|22|30|在復活的時候，人也不娶也不嫁，而是像天上的天使一樣。
MATT|22|31|論到死人復活，上帝向你們所說的話，你們沒有念過嗎？
MATT|22|32|他說：『我是 亞伯拉罕 的上帝， 以撒 的上帝， 雅各 的上帝。』上帝不是死人的上帝，而是活人的上帝。」
MATT|22|33|眾人聽見這話，對他的教導非常驚訝。
MATT|22|34|法利賽人聽見耶穌堵住了撒都該人的口，他們就聚集在一起。
MATT|22|35|其中有一個人是律法師 ，要試探耶穌，就問他：
MATT|22|36|「老師，律法上的誡命哪一條是最大的呢？」
MATT|22|37|耶穌對他說：「你要盡心、盡性、盡意愛主—你的上帝。
MATT|22|38|這是最大的，且是第一條誡命。
MATT|22|39|第二條也如此，就是要愛鄰 如己。
MATT|22|40|這兩條誡命是一切律法和先知書的總綱。」
MATT|22|41|法利賽人聚集的時候，耶穌問他們：
MATT|22|42|「論到基督，你們的意見如何？他是誰的後裔呢？」他們說：「是 大衛 的。」
MATT|22|43|耶穌說：「這樣， 大衛 被聖靈感動，怎麼還稱他為主，說：
MATT|22|44|『主對我主說： 你坐在我的右邊， 等我把你的仇敵放在你腳下？』
MATT|22|45|大衛 既稱他為主，他怎麼又是 大衛 的後裔呢？」
MATT|22|46|沒有一個人能回答一句話，從那日以後沒有人敢再問他甚麼。
MATT|23|1|那時，耶穌對眾人和門徒講論，
MATT|23|2|說：「文士和法利賽人坐在 摩西 的位上，
MATT|23|3|所以凡他們所吩咐你們的，你們都要謹守遵行。但不要效法他們的行為，因為他們能說不能行。
MATT|23|4|他們把難挑的 重擔捆起來，擱在人的肩上，但自己一個指頭也不肯動。
MATT|23|5|他們所做的一切事都是要讓人看見，所以把佩戴的經匣 加寬了，衣裳的繸子加長了，
MATT|23|6|喜愛宴席上的首座、會堂裏的高位，
MATT|23|7|又喜歡人們在街市上向他們問安，稱呼他們拉比 。
MATT|23|8|但你們不要接受拉比的稱呼，因為只有一位是你們的老師；你們都是弟兄。
MATT|23|9|也不要稱呼地上的人為父，因為只有一位是你們的父，就是在天上的父。
MATT|23|10|不要接受師傅的稱呼，因為只有一位是你們的師傅，就是基督。
MATT|23|11|你們中間誰為大，誰就要作你們的用人。
MATT|23|12|凡自高的，必降為卑；自甘卑微的，必升為高。
MATT|23|13|「你們這假冒為善的文士和法利賽人有禍了！因為你們當著人的面把天國的門關了，自己不進去，要進去的人，你們也不容他們進去。
MATT|23|14|
MATT|23|15|「你們這假冒為善的文士和法利賽人有禍了！因為你們走遍海洋陸地，說服一個人入教，既入了教，卻使他成為比你們加倍壞的地獄之子。
MATT|23|16|「你們這瞎眼的嚮導有禍了！你們說：『凡指著聖所起誓的算不得甚麼；但是凡指著聖所中的金子起誓的，他就該謹守。』
MATT|23|17|你們這無知的瞎子啊，哪個更大呢？是金子，還是使金子成聖的聖所呢？
MATT|23|18|你們又說：『凡指著祭壇起誓的算不得甚麼；但是凡指著壇上祭物起誓的，他就該謹守。』
MATT|23|19|你們這些瞎子啊，哪個更大呢？是祭物，還是使祭物成聖的壇呢？
MATT|23|20|所以，人指著祭壇起誓，就是指著壇和壇上一切所有的起誓；
MATT|23|21|人指著聖所起誓，就是指著聖所和那住在聖所裏的起誓；
MATT|23|22|人指著天起誓，就是指著上帝的寶座和那坐在上面的起誓。
MATT|23|23|「你們這假冒為善的文士和法利賽人有禍了！因為你們將薄荷、大茴香、小茴香獻上十分之一，那律法上更重要的事，就是公義、憐憫、信實，你們反倒不做；這原是你們該做的－至於那些奉獻也不可廢棄。
MATT|23|24|你們這瞎眼的嚮導，蠓蟲你們就濾出來，駱駝你們倒吞下去。
MATT|23|25|「你們這假冒為善的文士和法利賽人有禍了！因為你們洗淨杯盤的外面，裏面卻滿了貪婪和放蕩。
MATT|23|26|你這瞎眼的法利賽人，先洗淨杯子 的裏面，好使外面也乾淨了。
MATT|23|27|「你們這假冒為善的文士和法利賽人有禍了！因為你們好像粉飾了的墳墓，外面好看，裏面卻滿了死人的骨頭和一切的污穢。
MATT|23|28|你們也是如此，外面對人顯出公義，裏面卻滿了虛偽和不法的事。
MATT|23|29|「你們這假冒為善的文士和法利賽人有禍了！因為你們建造先知的墳，裝修義人的墓，
MATT|23|30|說：『若是我們在先祖的時代，必不和他們一同流先知的血。』
MATT|23|31|這樣，你們就證明自己是殺害先知的人的子孫了。
MATT|23|32|你們去充滿你們祖宗的惡貫吧！
MATT|23|33|你們這些蛇啊，毒蛇的孽種啊，怎能逃脫地獄的懲罰呢？
MATT|23|34|所以，我差遣先知、智慧人和文士到你們這裏來，有的你們要殺害，要釘十字架；有的你們要在會堂裏鞭打，從這城追逼到那城，
MATT|23|35|如此，地上所有義人流的血都歸到你們身上，從義人 亞伯 的血起，直到你們在聖所和祭壇中間所殺的 巴拉加 的兒子 撒迦利亞 的血為止。
MATT|23|36|我實在告訴你們，這一切的罪都要歸到這世代了。」
MATT|23|37|「 耶路撒冷 啊， 耶路撒冷 啊，你常殺害先知，又用石頭打死那奉差遣到你這裏來的人。我多少次想聚集你的兒女，好像母雞把小雞聚集在翅膀底下，但是你們不願意。
MATT|23|38|看吧，你們的家要被廢棄成為荒蕪。
MATT|23|39|我告訴你們，從今以後，你們絕不會再見到我，直到你們說：『奉主名來的是應當稱頌的！』」
MATT|24|1|耶穌出了聖殿，正離開的時候，門徒前來，把聖殿的建築指給他看。
MATT|24|2|耶穌回應他們說：「你們不是看見這一切嗎？我實在告訴你們，這裏將沒有一塊石頭會留在另一塊石頭上，而不被拆毀的。」
MATT|24|3|耶穌在 橄欖山 上坐著，門徒私下進前來問他：「請告訴我們，甚麼時候有這些事呢？你來臨和世代的終結有甚麼預兆呢？」
MATT|24|4|耶穌回答他們：「你們要謹慎，免得有人迷惑你們。
MATT|24|5|因為將有好些人冒我的名來，說『我是基督』，並且要迷惑許多人。
MATT|24|6|你們也將聽見打仗和打仗的風聲。注意，不要驚慌！因為這些事必須發生，但這還不是終結。
MATT|24|7|民要攻打民，國要攻打國，多處必有饑荒、地震。
MATT|24|8|這都是災難 的起頭。
MATT|24|9|那時，人要使你們陷在患難裏，也要殺害你們；你們又要為我的名被萬民憎恨。
MATT|24|10|那時，會有許多人跌倒，也會彼此陷害，彼此憎恨；
MATT|24|11|且有好些假先知起來，迷惑許多人。
MATT|24|12|因為不法的事增多，許多人的愛心漸漸冷淡了。
MATT|24|13|但堅忍到底的終必得救。
MATT|24|14|這天國的福音要傳遍天下，對萬民作見證，然後終結才來到。」
MATT|24|15|「當你們看見先知 但以理 所說的那『施行毀滅的褻瀆者』站在聖地（讀這經的人要會意），
MATT|24|16|那時，在 猶太 的，應當逃到山上；
MATT|24|17|在屋頂上的，不要下來拿家裏的東西；
MATT|24|18|在田裏的，不要回去取衣裳。
MATT|24|19|在那些日子，懷孕的和奶孩子的就苦了。
MATT|24|20|你們要祈求，好讓你們逃走的時候，不遇見冬天或安息日。
MATT|24|21|因為那時必有大災難，自從世界的起頭直到如今，從沒有這樣的災難，將來也不會有。
MATT|24|22|若不減少那些日子，凡血肉之軀的，就沒有一個能得救；可是為了選民，那些日子將減少。
MATT|24|23|那時，若有人對你們說：『看哪，基督在這裏！』或『在那裏！』你們不要信。
MATT|24|24|因為假基督和假先知將要起來，顯大神蹟、大奇事，如果可能，要把選民也迷惑了。
MATT|24|25|看哪，我已經預先告訴你們了。
MATT|24|26|若有人對你們說：『看哪，基督在曠野裏！』你們不要出去；或說：『看哪，基督在內室中！』你們不要信。
MATT|24|27|好像閃電從東邊發出，直照到西邊，人子來臨也要這樣。
MATT|24|28|屍首在哪裏，鷹也會聚在哪裏。」
MATT|24|29|「那些日子的災難一過去， 太陽要變黑， 月亮也不放光， 眾星要從天上墜落， 天上的萬象都要震動。
MATT|24|30|那時，人子的預兆要顯在天上，地上的萬族都要哀哭。他們要看見人子帶著能力和大榮耀，駕著天上的雲來臨。
MATT|24|31|他要差遣天使，用大聲的號筒，從四方，從天這邊直到天那邊，召集他的選民。」
MATT|24|32|「你們要從無花果樹學習功課：當樹枝發芽長葉的時候，你們就知道夏天近了。
MATT|24|33|同樣，當你們看見這一切，就知道那時候近了，就在門口了。
MATT|24|34|我實在告訴你們，這世代還沒有過去，這一切都要發生。
MATT|24|35|天地要廢去，我的話卻絕不廢去。」
MATT|24|36|「但那日子，那時辰，沒有人知道，連天上的天使也不知道，子也不知道，惟有父知道。
MATT|24|37|挪亞 的日子怎樣，人子來臨也要怎樣。
MATT|24|38|在洪水以前的那些日子，人照常吃喝嫁娶，直到 挪亞 進方舟的那日，
MATT|24|39|不知不覺洪水來了，把他們全都沖去。人子來臨也要這樣。
MATT|24|40|那時，兩個人在田裏，一個被接去，一個被撇下。
MATT|24|41|兩個女人推磨，一個被接去，一個被撇下。
MATT|24|42|所以，你們要警醒，因為不知道你們的主哪一天來到。
MATT|24|43|你們要知道，一家的主人若知道晚上甚麼時候有賊來，就必警醒，不讓賊挖穿房屋。
MATT|24|44|所以，你們也要預備，因為在你們想不到的時候，人子就來了。」
MATT|24|45|「那麼，誰是那忠心又精明的僕人，主人派他管理自己的家僕、按時分糧給他們的呢？
MATT|24|46|主人來到，看見僕人這樣做，那僕人就有福了。
MATT|24|47|我實在告訴你們，主人要派他管理所有的財產。
MATT|24|48|如果那惡僕心裏說：『我的主人會來得遲』，
MATT|24|49|就動手打他的同伴，又和醉酒的人一同吃喝，
MATT|24|50|在想不到的日子，不知道的時候，那僕人的主人要來，
MATT|24|51|重重地懲罰他 ，定他和假冒為善的人同罪，在那裏他要哀哭切齒了。」
MATT|25|1|「那時，天國好比十個童女拿著燈出去迎接新郎。
MATT|25|2|其中有五個是愚拙的，五個是聰明的。
MATT|25|3|愚拙的拿著燈，卻沒有帶油；
MATT|25|4|聰明的拿著燈，又盛了油在器皿裏。
MATT|25|5|新郎遲延的時候，她們都打盹，睡著了。
MATT|25|6|半夜有人喊：『看，新郎來了，你們出來迎接他。』
MATT|25|7|那些童女就都起來挑亮她們的燈。
MATT|25|8|愚拙的對聰明的說：『請分點油給我們，因為我們的燈要滅了。』
MATT|25|9|聰明的回答：『恐怕不夠你我用的；你們還是自己到賣油的那裏去買吧。』
MATT|25|10|她們去買的時候，新郎到了。那預備好了的，與他進去共赴婚宴，門就關了。
MATT|25|11|其餘的童女隨後也來了，說：『主啊，主啊，給我們開門！』
MATT|25|12|他卻回答：『我實在告訴你們，我不認識你們。』
MATT|25|13|所以，你們要警醒，因為那日子，那時辰，你們不知道。」
MATT|25|14|「天國又好比一個人要出外遠行，就叫了僕人來，把他的家業交給他們。
MATT|25|15|他按著各人的才幹，給他們銀子：一個給了五千 ，一個給了二千 ，一個給了一千 ，就出外遠行去了。
MATT|25|16|那領五千的立刻拿去做買賣，另外賺了五千。
MATT|25|17|那領二千的也照樣另賺了二千。
MATT|25|18|但那領一千的去掘開地，把主人的銀子埋藏了。
MATT|25|19|過了許久，那些僕人的主人來了，和他們算賬。
MATT|25|20|那領五千的又帶著另外的五千來，說：『主啊，你交給我五千。請看，我又賺了五千。』
MATT|25|21|主人說：『好，你這又善良又忠心的僕人，你在少許的事上忠心，我要派你管理許多的事，進來享受你主人的快樂吧！』
MATT|25|22|那領二千的也進前來，說：『主啊，你交給我二千。請看，我又賺了二千。』
MATT|25|23|主人說：『好，你這又善良又忠心的僕人，你在少許的事上忠心，我要派你管理許多的事，進來享受你主人的快樂吧！』
MATT|25|24|那領一千的也進前來，說：『主啊，我知道你，你是個嚴厲的人：沒有種的地方也要收割，沒有播的地方也要收穫，
MATT|25|25|我就害怕，去把你的一千銀子埋藏在地裏。請看，你的銀子在這裏。』
MATT|25|26|他的主人回答他說：『你這又惡又懶的僕人，你既知道我沒有種的地方也要收割，沒有播的地方也要收穫，
MATT|25|27|就該把我的銀子放給兌換銀錢的人，到我來的時候可以連本帶利收回。
MATT|25|28|把他這一千奪過來，給那有一萬 的。
MATT|25|29|因為凡有的，還要加給他，叫他有餘；沒有的，連他所有的也要奪過來。
MATT|25|30|把這無用的僕人丟在外面黑暗裏，在那裏他要哀哭切齒了。』」
MATT|25|31|「當人子在他榮耀裏，同著眾天使來臨的時候，要坐在他榮耀的寶座上。
MATT|25|32|萬民都要聚集在他面前。他要把他們分別出來，好像牧人分別綿羊、山羊一般，
MATT|25|33|把綿羊安置在右邊，山羊在左邊。
MATT|25|34|於是王要向他右邊的說：『你們這蒙我父賜福的，可來承受那創世以來為你們所預備的國。
MATT|25|35|因為我餓了，你們給我吃；渴了，你們給我喝；我流浪在外，你們留我住；
MATT|25|36|我赤身露體，你們給我穿；我病了，你們看顧我；我在監獄裏，你們來看我。』
MATT|25|37|義人就回答：『主啊，我們甚麼時候見你餓了，給你吃；渴了，給你喝？
MATT|25|38|甚麼時候見你流浪在外，留你住；或是赤身露體，給你穿？
MATT|25|39|又甚麼時候見你病了，或是在監獄裏，來看你呢？』
MATT|25|40|王回答他們說：『我實在告訴你們，這些事你們做在我弟兄中一個最小的身上，就是做在我身上了。』
MATT|25|41|「王又要向那左邊的說：『你們這被詛咒的人，離開我！進入那為魔鬼和他的使者所預備的永火裏去！
MATT|25|42|因為我餓了，你們沒有給我吃；渴了，你們沒有給我喝；
MATT|25|43|我流浪在外，你們沒有留我住；我赤身露體，你們沒有給我穿；我病了，我在監獄裏，你們沒有來看顧我。』
MATT|25|44|他們也要回答：『主啊，我們甚麼時候見你餓了，或渴了，或流浪在外，或赤身露體，或病了，或在監獄裏，沒有伺候你呢？』
MATT|25|45|王要回答：『我實在告訴你們，這些事你們沒有做在任何一個最小的弟兄身上，就是沒有做在我身上了。』
MATT|25|46|這些人要往永刑裏去；那些義人要往永生裏去。」
MATT|26|1|耶穌說完了這一切的話，就對門徒說：
MATT|26|2|「你們知道，過兩天是逾越節，人子將要被出賣，釘在十字架上。」
MATT|26|3|那時，祭司長和百姓的長老聚集在那稱為 該亞法 的大祭司的院裏。
MATT|26|4|大家商議要設計捉拿耶穌，把他殺掉。
MATT|26|5|可是他們說：「不可在過節的日子，恐怕百姓生亂。」
MATT|26|6|耶穌在 伯大尼 的痲瘋病人 西門 家裏，
MATT|26|7|有一個女人拿著一玉瓶極貴的香膏來，趁耶穌坐席的時候，澆在他的頭上。
MATT|26|8|門徒看見就很不高興，說：「何必這樣浪費呢！
MATT|26|9|這香膏可以賣許多錢，賙濟窮人。」
MATT|26|10|耶穌看出他們的意思，就說：「為甚麼難為這女人呢？她在我身上做的是一件美事。
MATT|26|11|因為常有窮人和你們在一起，但是你們不常有我。
MATT|26|12|她把這香膏澆在我身上是為我安葬作準備的。
MATT|26|13|我實在告訴你們，普天之下，無論在甚麼地方傳這福音，都要述說這女人所做的，來記念她。」
MATT|26|14|當時，十二使徒中有一個叫 加略 人 猶大 的，去見祭司長，
MATT|26|15|說：「我把他交給你們，你們願意給我多少錢？」他們給了他三十塊銀錢。
MATT|26|16|從那時候起，他就找機會要把耶穌交給他們。
MATT|26|17|除酵節的第一天，門徒來問耶穌：「你要我們在哪裏給你預備吃逾越節的宴席呢？」
MATT|26|18|耶穌說：「你們進城去，到某人那裏，對他說：『老師說：我的時候快到了，我要和我的門徒在你家裏守逾越節。』」
MATT|26|19|門徒遵照耶穌所吩咐的去預備了逾越節的宴席。
MATT|26|20|到了晚上，耶穌和十二使徒坐席。
MATT|26|21|他們吃的時候，耶穌說：「我實在告訴你們，你們中間有一個人要出賣我。」
MATT|26|22|他們就非常憂愁，一個一個地問他：「主，該不是我吧？」
MATT|26|23|耶穌回答說：「同我蘸手在盤子裏的，就是要出賣我的。
MATT|26|24|人子要去了，正如經上所寫有關他的；但出賣人子的人有禍了！那人沒有出生倒好。」
MATT|26|25|出賣耶穌的 猶大 回答他說：「拉比，該不是我吧？」耶穌說：「你自己說了。」
MATT|26|26|他們吃的時候，耶穌拿起餅來，祝福了，就擘開，遞給門徒，說：「你們拿去，吃吧。這是我的身體。」
MATT|26|27|他又拿起杯來，祝謝了，遞給他們，說：「你們都喝這個，
MATT|26|28|因為這是我立約的血，為許多人流出來，使罪得赦。
MATT|26|29|但我告訴你們，從今以後，我不再喝這葡萄汁，直到我在我父的國裏與你們同喝新的那日子。」
MATT|26|30|他們唱了詩，就出來往 橄欖山 去。
MATT|26|31|那時，耶穌對他們說：「今夜，你們為我的緣故都要跌倒。因為經上記著： 『我要擊打牧人， 羊就分散了。』
MATT|26|32|但我復活以後，要在你們之前往 加利利 去。」
MATT|26|33|彼得 回答他說：「即使眾人為你的緣故跌倒，我也絕不跌倒。」
MATT|26|34|耶穌說：「我實在告訴你，今夜雞叫以前，你要三次不認我。」
MATT|26|35|彼得 說：「我就是必須和你同死，也絕不會不認你。」所有的門徒都是這樣說。
MATT|26|36|耶穌和門徒來到一個地方，名叫 客西馬尼 。他對他們說：「你們坐在這裏，我到那邊去禱告。」
MATT|26|37|於是他帶著 彼得 和 西庇太 的兩個兒子同去。他憂愁起來，極其難過，
MATT|26|38|就對他們說：「我心裏非常憂傷，幾乎要死；你們留在這裏，和我一同警醒。」
MATT|26|39|他就稍往前走，俯伏在地，禱告說：「我父啊，如果可能，求你使這杯離開我。然而，不是照我所願的，而是照你所願的。」
MATT|26|40|他回到門徒那裏，見他們睡著了，就對 彼得 說：「怎麼樣？你們不能同我警醒一小時嗎？
MATT|26|41|總要警醒禱告，免得陷入試探。你們心靈固然願意，肉體卻軟弱了。」
MATT|26|42|他第二次又去禱告說：「我父啊，這杯若不能離開我，必須我喝，就願你的旨意成全。」
MATT|26|43|他又來，見他們睡著了，因為他們的眼睛困倦。
MATT|26|44|耶穌又離開他們，第三次去禱告，說的話跟先前一樣。
MATT|26|45|然後他來到門徒那裏，對他們說：「現在你們仍在睡覺安歇嗎？看哪，時候到了，人子被出賣在罪人手裏了。
MATT|26|46|起來，我們走吧！看哪，那出賣我的人快來了。」
MATT|26|47|耶穌還在說話的時候，十二使徒之一的 猶大 來了，還有一大群人帶著刀棒，從祭司長和百姓的長老那裏跟他同來。
MATT|26|48|那出賣耶穌的給了他們一個暗號，說：「我親誰，誰就是。你們把他抓住。」
MATT|26|49|猶大 立刻進前來對耶穌說：「拉比，你好！」就跟他親吻。
MATT|26|50|耶穌對他說：「朋友，你來要做的事，就做吧。 」於是那些人上前，下手抓住耶穌。
MATT|26|51|忽然，有一個和耶穌一起的人伸手拔出刀來，把大祭司的僕人砍了一刀，削掉了他一隻耳朵。
MATT|26|52|耶穌對他說：「收刀入鞘吧！凡動刀的，必死在刀下。
MATT|26|53|你想我不能求我父，現在為我差遣比十二營還多的天使來嗎？
MATT|26|54|若是這樣，經上所說事情必須如此發生的話怎麼應驗呢？」
MATT|26|55|就在那時，耶穌對眾人說：「你們帶著刀棒出來抓我，如同拿強盜嗎？我天天坐在聖殿裏教導人，你們並沒有抓我。
MATT|26|56|但這整件事的發生，是要應驗先知書上的話。」那時，門徒都離開他，逃走了。
MATT|26|57|抓耶穌的人把他帶到大祭司 該亞法 那裏去，文士和長老已經在那裏聚集。
MATT|26|58|彼得 遠遠地跟著耶穌，直到大祭司的院子，進到裏面，就和警衛同坐，要看結局怎樣。
MATT|26|59|祭司長和全議會尋找假見證控告耶穌，要處死他。
MATT|26|60|雖然有好些人來作假見證，總找不到實據。最後有兩個人前來，
MATT|26|61|說：「這個人曾說：『我能拆毀上帝的殿，三日內又建造起來。』」
MATT|26|62|大祭司就站起來，對耶穌說：「這些人作證告你的事，你甚麼都不回答嗎？」
MATT|26|63|耶穌卻不言語。大祭司對他說：「我指著永生上帝命令你起誓告訴我們，你是不是基督—上帝的兒子？」
MATT|26|64|耶穌對他說：「你自己說了。然而，我告訴你們， 此後你們要看見人子 坐在權能者的右邊， 駕著天上的雲來臨。」
MATT|26|65|大祭司就撕裂衣服，說：「他說了褻瀆的話，我們何必再要證人呢？現在你們已經聽見他這褻瀆的話了。
MATT|26|66|你們的意見如何？」他們回答：「他該處死。」
MATT|26|67|他們就吐唾沫在他臉上，用拳頭打他，也有打他耳光的，
MATT|26|68|說：「基督啊，向我們說預言吧！打你的是誰？」
MATT|26|69|彼得 在外面院子裏坐著，有一個使女進前來，說：「你素來也是同那 加利利 人耶穌一起的。」
MATT|26|70|彼得 在眾人面前卻不承認，說：「我不知道你說的是甚麼！」
MATT|26|71|他出去，到了門口，又有一個使女看見他，就對那裏的人說：「這個人是同 拿撒勒 人耶穌一起的。」
MATT|26|72|彼得 又不承認，起誓說：「我不認得那個人。」
MATT|26|73|過了不久，旁邊站著的人前來，對 彼得 說：「你的確是他們一夥的，你的口音把你顯露出來了。」
MATT|26|74|彼得 就賭咒發誓說：「我不認得那個人。」立刻雞就叫了。
MATT|26|75|彼得 想起耶穌所說的話：「雞叫以前，你要三次不認我。」他就出去痛哭。
MATT|27|1|到了早晨，眾祭司長和百姓的長老商議要處死耶穌，
MATT|27|2|就把他綁著，解去，交給 彼拉多 總督。
MATT|27|3|這時，出賣耶穌的 猶大 看見耶穌已經定了罪，就後悔，把那三十塊銀錢拿回來給祭司長和長老，
MATT|27|4|說：「我出賣了無辜人的血有罪了。」他們說：「那跟我們有甚麼相干？你自己承當吧！」
MATT|27|5|猶大 就把那銀錢丟在殿裏，出去吊死了。
MATT|27|6|祭司長拾起銀錢來，說：「這是血價，不可放在聖殿的銀庫裏。」
MATT|27|7|他們商議，就用那銀錢買了窯戶的一塊田，用來埋葬外鄉人。
MATT|27|8|所以，那塊田直到今日還叫做「血田」。
MATT|27|9|這就應驗了先知 耶利米 所說的話：「他們用那三十塊銀錢，就是 以色列 人給那被估定的人所估定的價錢，
MATT|27|10|買了窯戶的一塊田；這是照著主所吩咐我的。」
MATT|27|11|耶穌站在總督面前，總督問他：「你是 猶太 人的王嗎？」耶穌說：「是你說的。」
MATT|27|12|他被祭司長和長老控告的時候，甚麼都不回答。
MATT|27|13|彼拉多 就對他說：「他們作證告你這麼多的事，你沒有聽見嗎？」
MATT|27|14|耶穌仍不回答，連一句話也不說，以致總督覺得非常驚訝。
MATT|27|15|總督有一個常例，每逢這節期，隨眾人的意願釋放一個囚犯給他們。
MATT|27|16|當時有一個出名的囚犯叫 巴拉巴 。
MATT|27|17|眾人聚集的時候， 彼拉多 就對他們說：「你們要我釋放哪一個給你們？是 巴拉巴 呢？是稱為基督的耶穌呢？」
MATT|27|18|總督原知道他們是因為嫉妒才把他解了來。
MATT|27|19|正坐堂的時候，他的夫人打發人來說：「這義人的事，你一點不可管，因為我今天在夢中因他受了許多的苦。」
MATT|27|20|祭司長和長老挑唆眾人，要求釋放 巴拉巴 ，除掉耶穌。
MATT|27|21|總督回答他們說：「這兩個人，你們要我釋放哪一個給你們呢？」他們說：「 巴拉巴 。」
MATT|27|22|彼拉多 說：「這樣，那稱為基督的耶穌我怎麼辦他呢？」他們都說：「把他釘十字架！」
MATT|27|23|總督說：「為甚麼？他做了甚麼惡事呢？」他們更加喊著說：「把他釘十字架！」
MATT|27|24|彼拉多 見說也無濟於事，反要生亂，就拿水在眾人面前洗手，說：「流這人 的血，罪不在我，你們承當吧。」
MATT|27|25|眾人都回答：「他的血歸到我們和我們的子孫身上！」
MATT|27|26|於是 彼拉多 釋放 巴拉巴 給他們，把耶穌鞭打後交給人釘十字架。
MATT|27|27|總督的兵把耶穌帶進總督府，把全營的兵都聚集在耶穌那裏。
MATT|27|28|他們脫了他的衣服，穿上一件朱紅色的袍子，
MATT|27|29|用荊棘編了冠冕，戴在他頭上，拿一根蘆葦稈放在他右手裏，跪在他面前，戲弄他，說：「萬歲， 猶太 人的王！」
MATT|27|30|他們又向他吐唾沫，拿蘆葦稈打他的頭。
MATT|27|31|他們戲弄完了，就給他脫了袍子，又穿上他自己的衣服，帶他出去，要釘十字架。
MATT|27|32|他們出去的時候，遇見一個 古利奈 人，名叫 西門 ，就強迫他同去，好背耶穌的十字架。
MATT|27|33|他們到了一個地方，名叫 各各他 ，就是「髑髏地」。
MATT|27|34|士兵拿苦膽調和的酒給耶穌喝。他嘗了，不肯喝。
MATT|27|35|他們把他釘在十字架上，然後抽籤分了他的衣服，
MATT|27|36|又坐在那裏看守他。
MATT|27|37|他們在他頭上方安了一個罪狀牌，寫著：「這是 猶太 人的王耶穌。」
MATT|27|38|當時，有兩個強盜和他同釘十字架，一個在右邊，一個在左邊。
MATT|27|39|從那裏經過的人譏笑他，搖著頭，
MATT|27|40|說：「你這拆毀殿、三日又建造起來的，救救你自己吧！如果你是上帝的兒子，就從十字架上下來呀！」
MATT|27|41|眾祭司長、文士和長老也同樣嘲笑他，說：
MATT|27|42|「他救了別人，不能救自己。他是 以色列 的王，現在從十字架上下來，我們就信他。
MATT|27|43|他倚靠上帝，上帝若願意，現在就來救他，因為他曾說『我是上帝的兒子』。」
MATT|27|44|和他同釘的強盜也這樣譏諷他。
MATT|27|45|從正午到下午三點鐘，遍地都黑暗了。
MATT|27|46|約在下午三點鐘，耶穌大聲高呼，說：「以利！以利！拉馬撒巴各大尼？」就是說：「我的上帝！我的上帝！為甚麼離棄我？」
MATT|27|47|站在那裏的人，有的聽見就說：「這個人呼叫 以利亞 呢！」
MATT|27|48|其中有一個人立刻跑去，拿海綿蘸滿了醋，綁在蘆葦稈上，送給他喝。
MATT|27|49|其餘的人說：「且等著，看 以利亞 來不來救他。」
MATT|27|50|耶穌又大喊一聲，氣就斷了。
MATT|27|51|忽然，殿的幔子從上到下裂為兩半，地震動，磐石崩裂，
MATT|27|52|墳墓也開了，有許多已睡了的聖徒的身體也復活了。
MATT|27|53|耶穌復活以後，他們從墳墓裏出來，進了聖城，向許多人顯現。
MATT|27|54|百夫長和跟他一同看守耶穌的人看見地震和所經歷的事，非常害怕，說：「他真是上帝的兒子！」
MATT|27|55|有好些婦女在那裏，遠遠地觀看，她們是從 加利利 跟隨耶穌，來服事他的；
MATT|27|56|其中有 抹大拉 的 馬利亞 ，又有 雅各 和 約瑟 的母親 馬利亞 ，並有 西庇太 兩個兒子的母親。
MATT|27|57|到了晚上，有一個財主，名叫 約瑟 ，是 亞利馬太 來的，他也是耶穌的門徒。
MATT|27|58|這人去見 彼拉多 ，請求要耶穌的身體， 彼拉多 就吩咐給他。
MATT|27|59|約瑟 取了身體，用乾淨的細麻布裹好，
MATT|27|60|然後把他安放在自己的新墓穴裏，就是他鑿在巖石裏的。他又把大石頭滾到墓門口，然後離開。
MATT|27|61|有 抹大拉 的 馬利亞 和另一個 馬利亞 在那裏，對著墳墓坐著。
MATT|27|62|次日，就是預備日的第二天，祭司長和法利賽人聚集來見 彼拉多 ，
MATT|27|63|說：「大人，我們記得那迷惑人的還活著的時候曾說：『三天後我要復活。』
MATT|27|64|因此，請吩咐人將墳墓把守妥當，直到第三天，恐怕他的門徒來把他偷了去，就告訴百姓說：『他從死人中復活了。』這樣的話，那後來的迷惑就比先前的更厲害了。」
MATT|27|65|彼拉多 說：「你們有看守的兵，去吧！盡你們所能的把守妥當。」
MATT|27|66|他們就帶著看守的兵同去，封了石頭，將墳墓把守妥當。
MATT|28|1|安息日過後，七日的第一日，天快亮的時候， 抹大拉 的 馬利亞 和另一個 馬利亞 來看墳墓。
MATT|28|2|忽然，地大震動；因為有主的一個使者從天上下來，把石頭滾開，坐在上面。
MATT|28|3|他的相貌如同閃電，衣服潔白如雪。
MATT|28|4|看守的人嚇得渾身顫抖，甚至和死人一樣。
MATT|28|5|天使回應婦女說：「不要害怕！我知道你們是尋找那釘十字架的耶穌。
MATT|28|6|他不在這裏，照他所說的，他已經復活了。你們來！看看安放他的地方。
MATT|28|7|快去告訴他的門徒，說他已從死人中復活了，並且要比你們先到 加利利 去，在那裏你們會看見他。看哪！我已經告訴你們了。」
MATT|28|8|婦女們急忙離開墳墓，又害怕，又大為歡喜，跑去告訴他的門徒。
MATT|28|9|忽然，耶穌迎上她們，說：「平安！」她們就上前抱住他的腳拜他。
MATT|28|10|耶穌對她們說：「不要害怕！你們去告訴我的弟兄，叫他們往 加利利 去，在那裏會見到我。」
MATT|28|11|她們去的時候，看守的兵有幾個進城去，把所發生的事都報告祭司長。
MATT|28|12|祭司長和長老聚集商議，就拿許多銀錢給士兵，
MATT|28|13|說：「你們要這樣說：『夜間我們睡覺的時候，他的門徒來把他偷去了。』
MATT|28|14|若是這話被總督聽見，有我們勸他，保你們無事。」
MATT|28|15|士兵收了銀錢，就照所囑咐他們的去做。這話就在 猶太 人中間流傳，直到今日。
MATT|28|16|十一個門徒往 加利利 去，到了耶穌指定他們去的山上。
MATT|28|17|他們見了耶穌就拜他，然而還有人疑惑。
MATT|28|18|耶穌進前來，對他們說：「天上地下所有的權柄都賜給我了。
MATT|28|19|所以，你們要去，使萬民作我的門徒，奉父、子、聖靈的名給他們施洗 ，
MATT|28|20|凡我所吩咐你們的，都教導他們遵守。看哪，我天天與你們同在，直到世代的終結。」
MARK|1|1|上帝的兒子 ，耶穌基督福音的起頭。
MARK|1|2|正如 以賽亞 先知書上記著： 「看哪，我要差遣我的使者在你面前， 他要為你預備道路。
MARK|1|3|在曠野有聲音呼喊著： 預備主的道， 修直他的路。」
MARK|1|4|照這話，施洗 約翰 來到曠野 ，宣講悔改的洗禮，使罪得赦。
MARK|1|5|猶太 全地和全 耶路撒冷 的人都出去，到 約翰 那裏，承認他們的罪，在 約旦河 裏受他的洗。
MARK|1|6|約翰 穿駱駝毛的衣服，腰束皮帶，吃的是蝗蟲和野蜜。
MARK|1|7|他宣講，說：「有一位在我以後來的，能力比我更大，我就是彎腰給他解鞋帶也不配。
MARK|1|8|我用水給你們施洗，他卻要用聖靈給你們施洗。」
MARK|1|9|那時，耶穌從 加利利 的 拿撒勒 來，在 約旦河 裏受了 約翰 的洗。
MARK|1|10|他從水裏一上來，就看見天裂開了，聖靈彷彿鴿子降在他身上。
MARK|1|11|又有聲音從天上來，說：「你是我的愛子，我喜愛你。」
MARK|1|12|聖靈立刻把耶穌催促到曠野裏去。
MARK|1|13|他在曠野四十天，受撒但的試探，並與野獸同在一起，且有天使來伺候他。
MARK|1|14|約翰 下監以後，耶穌來到 加利利 ，宣講上帝的福音，
MARK|1|15|說：「日期滿了，上帝的國近了。你們要悔改，信福音！」
MARK|1|16|耶穌沿著 加利利 的海邊走，看見 西門 和 西門 的弟弟 安得烈 在海上撒網；他們本是打魚的。
MARK|1|17|耶穌對他們說：「來跟從我，我要叫你們得人如得魚一樣。」
MARK|1|18|他們立刻捨了網，跟從他。
MARK|1|19|耶穌稍往前走，又見 西庇太 的兒子 雅各 和他弟弟 約翰 在船上補網。
MARK|1|20|耶穌隨即呼召他們，他們就把父親 西庇太 和雇工留在船上，跟從了耶穌。
MARK|1|21|他們到了 迦百農 ，耶穌就在安息日進了會堂教導人。
MARK|1|22|他們對他的教導感到很驚奇，因為他教導他們正像有權柄的人，不像文士。
MARK|1|23|當時，會堂裏有一個污靈附身的人，他在喊叫，
MARK|1|24|說：「 拿撒勒 人耶穌，你為甚麼干擾我們？你來消滅我們嗎？我知道你是誰，你是上帝的聖者。」
MARK|1|25|耶穌斥責他說：「不要作聲，從這人身上出來吧！」
MARK|1|26|污靈使那人抽了一陣風，大聲喊叫，就出來了。
MARK|1|27|眾人都驚訝，以致彼此對問：「這是甚麼事？是個新的教導啊！他用權柄命令污靈，連污靈也聽從了他。」
MARK|1|28|於是耶穌的名聲立刻傳遍了全 加利利 周圍地區。
MARK|1|29|他們一出會堂，就同 雅各 和 約翰 進了 西門 和 安得烈 的家。
MARK|1|30|西門 的岳母正發燒躺著，就有人告訴耶穌。
MARK|1|31|耶穌進前拉著她的手，扶她起來，燒就退了，於是她服事他們。
MARK|1|32|傍晚日落的時候，有人帶著一切害病的和被鬼附的，來到耶穌跟前。
MARK|1|33|全城的人都聚集在門前。
MARK|1|34|耶穌治好了許多害各樣病的人，又趕出許多鬼，不許鬼說話，因為鬼認識他。
MARK|1|35|次日早晨，天未亮的時候，耶穌起來，到曠野地方去，在那裏禱告。
MARK|1|36|西門 和同伴出去找他，
MARK|1|37|找到了就對他說：「眾人都在找你！」
MARK|1|38|耶穌對他們說：「讓我們往別處去，到鄰近的鄉村，我也好在那裏傳道，因為我是為這事出來的。」
MARK|1|39|於是他走遍全 加利利 ，在他們的會堂傳道，並且趕鬼。
MARK|1|40|有一個痲瘋病人來求耶穌，向他跪下 ，說：「你若肯，你能使我潔淨。」
MARK|1|41|耶穌動了慈心，就伸手摸他，說：「我肯，你潔淨了吧！」
MARK|1|42|痲瘋病立刻離開他，他就潔淨了。
MARK|1|43|耶穌嚴嚴地叮囑他，立刻打發他走，
MARK|1|44|對他說：「你要注意，千萬不可告訴任何人，只要去，讓祭司為你檢查，又因為你已經潔淨，獻上 摩西 所吩咐的祭物，作為證據給眾人看。」
MARK|1|45|那人出去，倒說許多的話，把這件事傳揚開了，使耶穌不能再公開進城，只好留在外邊曠野地方，人從各處都到他跟前來。
MARK|2|1|過了些日子，耶穌又進了 迦百農 。人聽說他在屋裏，
MARK|2|2|於是許多人聚集，甚至連門前都沒有空地；耶穌就對他們講道。
MARK|2|3|有人帶著一個癱子來見耶穌，是由四個人抬來的；
MARK|2|4|因為人多，無法抬到耶穌跟前，就把他所在那房子的屋頂拆了，既拆通了，就把癱子連所躺臥的褥子都縋下去。
MARK|2|5|耶穌見他們的信心，就對癱子說：「孩子，你的罪赦了。」
MARK|2|6|有幾個文士坐在那裏，心裏議論，說：
MARK|2|7|「這個人為甚麼這樣說呢？他說褻瀆的話了。除了上帝一位之外，誰能赦罪呢？」
MARK|2|8|耶穌心中立刻知道他們心裏這樣議論，就說：「你們心裏為甚麼這樣議論呢？
MARK|2|9|對癱子說『你的罪赦了』，或說『起來！拿你的褥子行走』，哪一樣容易呢？
MARK|2|10|但要讓你們知道，人子在地上有赦罪的權柄。」就對癱子說：
MARK|2|11|「我吩咐你，起來！拿你的褥子回家去吧。」
MARK|2|12|那人就起來，立刻拿著褥子，當著眾人面前出去了，以致眾人都驚奇，歸榮耀給上帝，說：「我們從來沒有見過這樣的事！」
MARK|2|13|耶穌又到海邊去，眾人都到他跟前來，他就教導他們。
MARK|2|14|耶穌往前走，看見 亞勒腓 的兒子 利未 在稅關坐著，就對他說：「來跟從我！」他就起來跟從耶穌。
MARK|2|15|耶穌在 利未 家裏坐席的時候，有好些稅吏和罪人與耶穌和他的門徒一同坐席，因為有很多人也跟隨耶穌。
MARK|2|16|法利賽人中的文士 看見耶穌與罪人和稅吏一同吃飯，就對他的門徒說：「他與稅吏和罪人一同吃飯嗎？」
MARK|2|17|耶穌聽見，就對他們說：「健康的人用不著醫生，有病的人才用得著。我不是來召義人，而是召罪人。」
MARK|2|18|那時， 約翰 的門徒和法利賽人都禁食。他們來問耶穌說：「 約翰 的門徒和法利賽人的門徒禁食，你的門徒卻不禁食，這是為甚麼呢？」
MARK|2|19|耶穌對他們說：「新郎和賓客在一起的時候，賓客怎麼能禁食呢？只要新郎和他們在一起，他們不能禁食。
MARK|2|20|但日子將到，新郎要被帶走，那日他們就要禁食了。
MARK|2|21|「沒有人把新布縫在舊衣服上，若是這樣，所補上的新布會撕破舊衣服，裂口就更大了。
MARK|2|22|也沒有人把新酒裝在舊皮袋裏，若是這樣，酒會脹破皮袋，酒和皮袋都糟蹋了 。相反地，新酒要裝在新皮袋裏 。」
MARK|2|23|有一個安息日，耶穌從麥田經過。他的門徒走路的時候，摘起麥穗來。
MARK|2|24|法利賽人對耶穌說：「看哪！他們為甚麼做安息日不合法的事呢？」
MARK|2|25|耶穌對他們說：「 大衛 和跟從他的人飢餓需要食物時所做的事，你們沒有念過嗎？
MARK|2|26|他在 亞比亞他 作大祭司的時候，怎麼進了上帝的居所，吃了供餅，又給跟從他的人吃呢？這餅除了祭司以外，人都不可以吃。」
MARK|2|27|他又對他們說：「安息日是為人設立的，人不是為安息日設立的。
MARK|2|28|所以，人子也是安息日的主。」
MARK|3|1|耶穌又進了會堂，在那裏有一個人，他的一隻手萎縮了。
MARK|3|2|眾人為了要控告耶穌，就窺探他會不會在安息日醫治那人。
MARK|3|3|耶穌對那手萎縮了的人說：「起來站在當中！」
MARK|3|4|他又問眾人：「在安息日行善行惡，救命害命，哪樣是合法的呢？」他們都不作聲。
MARK|3|5|耶穌怒目環視他們，因他們的心剛硬而憂傷，就對那人說：「伸出手來！」他把手一伸，手就復原了。
MARK|3|6|法利賽人出去，立刻同 希律 一黨的人商議怎樣除掉耶穌。
MARK|3|7|耶穌和門徒退到海邊去，有許多人從 加利利 跟隨他。還有許多人聽見他所做的事，就從 猶太 、 耶路撒冷 、 以土買 、 約旦河 的東邊，以及 推羅 和 西頓 的附近地方來到他那裏。
MARK|3|8|
MARK|3|9|因為人多，他吩咐門徒為他預備一隻小船，免得眾人擁擠他。
MARK|3|10|他治好了許多人，所以凡有疾病的，都擠著要摸他。
MARK|3|11|每當污靈看見他，就俯伏在他面前，喊著說：「你是上帝的兒子。」
MARK|3|12|耶穌再三囑咐他們不要把他宣揚出去。
MARK|3|13|耶穌上了山，把自己所要的人召來，他們就來到他那裏。
MARK|3|14|於是他設立十二個人，又稱他們為使徒 ，要他們常和自己同在，也要差他們去傳道，
MARK|3|15|並給他們權柄趕鬼。
MARK|3|16|他設立的十二個人 有 西門 －耶穌又給他起名叫 彼得 ，
MARK|3|17|還有 西庇太 的兒子 雅各 和 雅各 的弟弟 約翰 —耶穌又給他們起名叫 半尼其 ，就是雷的兒子—
MARK|3|18|又有 安得烈 、 腓力 、 巴多羅買 、 馬太 、 多馬 、 亞勒腓 的兒子 雅各 、 達太 和激進黨的 西門 ，
MARK|3|19|還有出賣耶穌的 加略 人 猶大 。
MARK|3|20|耶穌進了屋子，眾人又聚集，甚至他連飯也顧不得吃。
MARK|3|21|耶穌的家人聽見，就出來要拉住他，因為他們說他癲狂了。
MARK|3|22|從 耶路撒冷 下來的文士說：「他是被 別西卜 附身的」，又說：「他是靠著鬼王趕鬼的。」
MARK|3|23|耶穌叫他們來，用比喻對他們說：「撒但怎能趕出撒但呢？
MARK|3|24|一國若自相紛爭，那國就立不住；
MARK|3|25|一家若自相紛爭，那家就立不住。
MARK|3|26|撒但若自相攻打紛爭，他就立不住，必定滅亡。
MARK|3|27|沒有人能進壯士家裏，搶奪他的東西；除非先綁住那壯士，否則無法搶奪他的家。
MARK|3|28|我實在告訴你們，世人一切的罪和一切褻瀆的話都可以得到赦免；
MARK|3|29|凡褻瀆聖靈的，卻永不得赦免，而要擔當永遠的罪。」
MARK|3|30|因為他們說：「他是被污靈附身的。」
MARK|3|31|那時，耶穌的母親和他兄弟來，站在外邊，打發人去叫他。
MARK|3|32|有許多人在耶穌周圍坐著，他們就告訴他說：「看哪！你母親、你兄弟和你姊妹 在外邊找你。」
MARK|3|33|耶穌回答他們：「誰是我的母親？誰是我的兄弟？」
MARK|3|34|就環視那周圍坐著的人，說：「看哪，我的母親，我的兄弟！
MARK|3|35|凡遵行上帝旨意的人就是我的兄弟姊妹和母親。」
MARK|4|1|耶穌又在海邊教導人。有一大群人到他那裏聚集，他只好上船坐下。船在海裏，眾人都靠近海，站在岸上。
MARK|4|2|耶穌就用許多比喻教導他們。在教導的時候，他對他們說：
MARK|4|3|「你們聽啊，有一個撒種的出去撒種。
MARK|4|4|他撒的時候，有的落在路旁，飛鳥來把它吃掉了。
MARK|4|5|有的落在土淺的石頭地上，因為土不深，很快就長出苗來，
MARK|4|6|太陽出來一曬，因為沒有根就枯乾了。
MARK|4|7|有的落在荊棘裏，荊棘長起來，把它擠住了，就結不出果實。
MARK|4|8|又有的落在好土裏，就發芽長大，結出果實，有三十倍的，有六十倍的，有一百倍的。」
MARK|4|9|耶穌又說：「有耳可聽的，就應當聽！」
MARK|4|10|耶穌獨自一人的時候，跟隨他的人和十二使徒問他這些比喻的意思。
MARK|4|11|耶穌對他們說：「上帝國的奧祕只讓你們知道，若是對外人講，凡事就用比喻，
MARK|4|12|要 他們看了又看，卻看不清， 聽了又聽，卻不明白， 免得他們回轉過來，獲得赦免。」
MARK|4|13|耶穌又對他們說：「你們不明白這比喻嗎？這樣怎能明白一切的比喻呢？
MARK|4|14|撒種的人所撒的就是道。
MARK|4|15|那撒在路旁的種子，就是人聽了道，撒但立刻來，把撒在他們心裏的道奪了去。
MARK|4|16|那撒在石頭地上的，就是人聽了道，立刻歡喜領受，
MARK|4|17|因心裏沒有根，不過是暫時的，一旦為道遭受患難或迫害，立刻就跌倒。
MARK|4|18|還有那撒在荊棘裏的，就是人聽了道，
MARK|4|19|後來有世上的憂慮、錢財的迷惑，和別樣的私慾進來，把道擠住了，結不出果實。
MARK|4|20|那撒在好土裏的，就是人聽了道，領受了，並且結了果實，有三十倍的，有六十倍的，有一百倍的。」
MARK|4|21|耶穌又對他們說：「人拿燈來，難道是要放在斗底下，床底下，而不放在燈臺上嗎？
MARK|4|22|因為掩藏的事沒有不顯出來的，隱瞞的事也沒有不露出來的。
MARK|4|23|有耳可聽的，就應當聽！」
MARK|4|24|他又說：「你們要留心所聽的。你們用甚麼量器來量，也將要用甚麼來量給你們，並且要多給你們。
MARK|4|25|因為有的，還要給他；沒有的，連他所有的也要奪去。」
MARK|4|26|耶穌又說：「上帝的國如同人把種子撒在地上，
MARK|4|27|黑夜睡覺，白日起來，這種子就發芽生長，那人卻不知道如何會這樣。
MARK|4|28|土地自然而然地出產五穀，先發苗，後長穗，然後穗上結成飽滿的穀子。
MARK|4|29|五穀熟了，就用鐮刀去割，因為收成的時候到了。」
MARK|4|30|耶穌又說：「我們可用甚麼來比擬上帝的國呢？可用甚麼比喻來說明呢？
MARK|4|31|它像一粒芥菜種，種在地裏的時候，雖比地上所有的種子都小，
MARK|4|32|但種下去以後，它長起來，比各樣的菜都大，又長出大枝，以致天上的飛鳥可以在它的蔭下築巢。」
MARK|4|33|耶穌用許多這樣的比喻，照他們所能聽的，對他們講道；
MARK|4|34|若不用比喻，他就不對他們講，但私下沒有人的時候，就把一切的道講給門徒聽。
MARK|4|35|那天晚上，耶穌對門徒說：「我們渡到對岸去吧。」
MARK|4|36|門徒離開眾人，耶穌已在船上，他們就請他一同去；也有別的船和他同行。
MARK|4|37|忽然狂風大作，波浪打入船內，以致船灌滿了水。
MARK|4|38|耶穌在船尾上，枕著枕頭睡覺。門徒叫醒他，說：「老師！我們快沒命了，你不管嗎？」
MARK|4|39|耶穌醒了，斥責那風，向海說：「住了吧！靜了吧！」風就止住，大大平靜了。
MARK|4|40|耶穌對他們說：「為甚麼膽怯？你們還沒有信心嗎？」
MARK|4|41|他們就非常懼怕，彼此說：「這到底是誰？連風和海都聽從他。」
MARK|5|1|他們渡到海的對岸，到 格拉森 人 的地區。
MARK|5|2|耶穌一下船，就有一個污靈附身的人從墳墓迎著他走來。
MARK|5|3|那人常住在墳墓裏，沒有人能捆住他，就是用鐵鏈也不能；
MARK|5|4|因為人屢次用腳鐐和鐵鏈捆鎖他，鐵鏈被他掙斷，腳鐐也被他弄碎了，總沒有人能制伏他。
MARK|5|5|他晝夜常在墳墓裏和山中喊叫，又用石頭打自己。
MARK|5|6|他遠遠看見耶穌，就跑過來拜他，
MARK|5|7|大聲呼叫說：「至高上帝的兒子耶穌，你為甚麼干擾我？我指著上帝懇求你，不要叫我受苦！」
MARK|5|8|這是因耶穌曾吩咐他說：「污靈啊，從這人身上出來！」
MARK|5|9|耶穌問他：「你叫甚麼名字？」他說：「我名叫 群 ，因為我們數目眾多。」
MARK|5|10|他就再三求耶穌不要叫他們離開那地方。
MARK|5|11|在山坡那裏，有一大群豬正在吃食；
MARK|5|12|污靈就央求耶穌，說：「求你打發我們進入豬群，好附著牠們。」
MARK|5|13|耶穌准了他們，污靈就出來，進入豬裏，那群豬就闖下山崖，投進海裏，淹死了。豬的數目約有二千。
MARK|5|14|放豬的逃跑了，去告訴城裏和鄉下的人。眾人就來，要看發生了甚麼事。
MARK|5|15|他們來到耶穌那裏，看見那被鬼附的人，就是曾被群鬼所附的，坐著，穿著衣服，神智清醒，他們就害怕。
MARK|5|16|看見這事的人把被鬼附的人所遇見的，和那群豬的事，都告訴了眾人，
MARK|5|17|眾人就央求耶穌離開他們的地區。
MARK|5|18|耶穌上船的時候，那曾被鬼附的人懇求要和耶穌在一起。
MARK|5|19|耶穌不許，卻對他說：「你回家去，到你的親友那裏，將主為你所做多麼大的事和他怎樣憐憫你，都告訴他們。」
MARK|5|20|那人就走了，開始在 低加坡里 傳揚耶穌為他做了多麼大的事，眾人就都驚訝。
MARK|5|21|耶穌又坐船 渡到對岸，有一大群人聚集到他身邊；他正在海邊。
MARK|5|22|有一個會堂主管，名叫 葉魯 ，也來了，一見到耶穌，就俯伏在他腳前，
MARK|5|23|再三求他，說：「我的小女兒快要死了，求你去為她按手，使她痊癒，可以活下去。」
MARK|5|24|耶穌就和他同去。 有一大群人跟隨他，擁擠著他。
MARK|5|25|有一個女人，患了經血不止的病有十二年，
MARK|5|26|在好多醫生手裏受了許多苦，又花盡了她所有的，一點也不見好，反而更重了。
MARK|5|27|她聽見耶穌的事，就夾在眾人中間，從後面來摸耶穌的衣裳，
MARK|5|28|因她想：「我只摸到他的衣裳，就會痊癒。」
MARK|5|29|於是她的流血立刻止住，她覺得身上的疾病好了。
MARK|5|30|耶穌頓時心裏覺得有能力從自己身上出去，就在眾人中間轉過來，說：「誰摸我的衣裳？」
MARK|5|31|門徒對他說：「你看眾人擁擠著你，還說『誰摸我』呢？」
MARK|5|32|耶穌周圍觀看，要見做這事的女人。
MARK|5|33|那女人知道在自己身上所成的事，就恐懼戰兢，來俯伏在耶穌跟前，將實情全告訴他。
MARK|5|34|耶穌對她說：「女兒，你的信救了你，平安地回去吧！你的疾病痊癒了。」
MARK|5|35|耶穌還在說話的時候，有人從會堂主管的家裏來，說：「你的女兒死了，何必還勞駕老師呢？」
MARK|5|36|耶穌不理會他們所說的話，就對會堂主管說：「不要怕，只要信！」
MARK|5|37|於是他帶著 彼得 、 雅各 和 雅各 的弟弟 約翰 同去，不許別人跟著他。
MARK|5|38|他們來到會堂主管的家裏，耶穌看到一片吵鬧，並有人大聲哭泣哀號，
MARK|5|39|就進到裏面，對他們說：「為甚麼大吵大哭呢？孩子不是死了，是睡著了。」
MARK|5|40|他們就嘲笑耶穌。耶穌把他們都趕出去，帶著孩子的父母和跟隨的人進了孩子所在的地方，
MARK|5|41|就拉著孩子的手，對她說：「大利大，古米！」翻出來就是說：「女孩，我吩咐你，起來！」
MARK|5|42|那女孩子立刻起來走動—她已經十二歲了；他們就非常驚奇。
MARK|5|43|耶穌切切地囑咐他們，不要讓人知道這事，又吩咐給她東西吃。
MARK|6|1|耶穌離開那裏，來到自己的家鄉；門徒也跟從他。
MARK|6|2|到了安息日，他在會堂裏教導人。眾人聽見，就很驚奇，說：「這人哪來這本事呢？所賜給他的是甚麼智慧？他手所做的是何等的異能呢？
MARK|6|3|這不是那木匠嗎？不是 馬利亞 的兒子 雅各 、 約西 、 猶大 、 西門 的長兄嗎？他姊妹們不也是在我們這裏嗎？」他們就厭棄他。
MARK|6|4|耶穌對他們說：「先知除了在本鄉、本族和自己的家之外，沒有不被尊敬的。」
MARK|6|5|耶穌在那裏不能行甚麼異能，不過為幾個病人按手，治好他們。
MARK|6|6|他也詫異他們不信。 耶穌走遍周圍鄉村教導人。
MARK|6|7|他叫了十二個使徒來，差遣他們兩個兩個地出去，也賜給他們權柄制伏污靈，
MARK|6|8|並且吩咐他們：途中不要帶食物和行囊，腰袋裏也不要帶錢，除了手杖以外，甚麼都不要帶；
MARK|6|9|只要穿鞋子，也不要穿兩件內衣。
MARK|6|10|他又對他們說：「你們無論到何處，進哪家，就住在哪裏，直到離開那地方。
MARK|6|11|若有甚麼地方的人不接待你們，不聽你們，你們離開那裏的時候，要跺掉你們腳上的塵土，證明他們的不是。」
MARK|6|12|使徒就出去傳道，叫人悔改，
MARK|6|13|又趕出許多鬼，用油抹了許多病人，治好他們。
MARK|6|14|耶穌的名聲傳開了， 希律 王也聽見。有人說：「施洗的 約翰 從死人中復活了，因此才有這些異能在他裏面運行。」
MARK|6|15|但別人說：「他是 以利亞 。」又有人說：「是先知，正如先知中的一位。」
MARK|6|16|希律 聽見卻說：「是我所斬的 約翰 ，他復活了。」
MARK|6|17|原來， 希律 為他兄弟 腓力 的妻子 希羅底 的緣故，派人去抓了 約翰 ，把他綁了在監獄裏，因為 希律 已經娶了那婦人。
MARK|6|18|約翰 曾對 希律 說：「你佔有你兄弟的妻子是不合法的。」
MARK|6|19|於是 希羅底 懷恨他，想要殺他，只是不能。
MARK|6|20|因為 希律 怕 約翰 ，知道他是義人，是聖人，所以就保護他，雖然聽了他的講論十分困惑 ，仍然樂意聽他。
MARK|6|21|有一天，恰巧是 希律 的生日， 希律 擺設宴席，請了大臣、千夫長和 加利利 的領袖。
MARK|6|22|他的女兒 希羅底 進來跳舞，使 希律 和同席的人都很高興。王就對女孩說：「無論你要甚麼，向我求，我都會給你」；
MARK|6|23|又對她多次 起誓說：「無論你向我求甚麼，就是我國家的一半，我也會給你。」
MARK|6|24|她就出去對她母親說：「我該求甚麼呢？」她母親說：「施洗 約翰 的頭。」
MARK|6|25|她就急忙進去見王，求他說：「我願王立刻把施洗 約翰 的頭放在盤子裏給我。」
MARK|6|26|王就很憂愁，然而因他所發的誓，又因同席的人，不願食言，
MARK|6|27|就立刻派一個衛兵，吩咐拿 約翰 的頭來。衛兵就去，在監獄裏斬了 約翰 ，
MARK|6|28|把頭放在盤子裏，拿來給那女孩，她就給她母親。
MARK|6|29|約翰 的門徒聽到了，就來把他的屍體領去，放在墳墓裏。
MARK|6|30|使徒們聚集到耶穌那裏，把一切所做的事、所傳的道全告訴他。
MARK|6|31|他就說：「你們來，同我私下到荒野的地方去歇一歇。」這是因為來往的人多，他們連吃飯的時間也沒有。
MARK|6|32|他們就坐船，私下往荒野的地方去。
MARK|6|33|眾人看見他們走了，有許多認識他們的，就從各城步行，一同跑到那裏，比他們先趕到了。
MARK|6|34|耶穌出來，見有一大群的人，就憐憫他們，因為他們如同羊沒有牧人一般，於是開始教導他們許多事。
MARK|6|35|天已經很晚，門徒進前來，說：「這地方偏僻，而且天已經很晚了，
MARK|6|36|請叫眾人散去，他們好往四面的鄉鎮村莊去，自己買些東西吃。」
MARK|6|37|耶穌回答他們說：「你們給他們吃吧！」門徒對他說：「我們要拿兩百個銀幣去買餅給他們吃嗎？」
MARK|6|38|耶穌說：「你們有多少餅？去看看。」他們知道後就說：「有五個，還有兩條魚。」
MARK|6|39|耶穌吩咐他們，叫眾人一組一組地坐在青草地上。
MARK|6|40|眾人就一群一群地坐下，有一百的，有五十的。
MARK|6|41|耶穌拿著這五個餅和兩條魚，望著天祝福，擘開餅，遞給門徒，擺在眾人面前，也把那兩條魚分給眾人。
MARK|6|42|他們都吃，並且吃飽了。
MARK|6|43|門徒把餅和魚的碎屑收拾起來，裝滿了十二個籃子。
MARK|6|44|吃餅的男人共有五千。
MARK|6|45|耶穌隨即催門徒上船，先渡到對岸，到 伯賽大 去，等他叫眾人散去。
MARK|6|46|他辭別了他們，就往山上去禱告。
MARK|6|47|到了晚上，船在海中，耶穌獨自在岸上。
MARK|6|48|他看見門徒因風不順，搖櫓很苦。天快亮的時候，他在海面上走，往他們那裏去，想要超過他們。
MARK|6|49|但門徒看見他在海面上走，以為是鬼怪，就喊叫起來；
MARK|6|50|因為他們都看見了他，甚為驚慌。耶穌連忙對他們說：「放心！是我，不要怕！」
MARK|6|51|於是他到他們那裏，一上船，風就停了；他們心裏十分驚奇。
MARK|6|52|這是因為他們不明白那分餅的事，心裏還是愚頑。
MARK|6|53|他們渡過了海，在 革尼撒勒 靠岸，泊了船，
MARK|6|54|他們一下來，眾人立刻認出是耶穌，
MARK|6|55|就跑遍那整個地區，聽到他在哪裏，就把有病的人用褥子抬到哪裏。
MARK|6|56|耶穌所到的地方，或村中、或城裏、或鄉間，他們都把病人放在街市上，求耶穌讓他們摸一摸他的衣裳繸子，摸著的人就都好了。
MARK|7|1|有法利賽人和幾個從 耶路撒冷 來的文士聚集到耶穌那裏。
MARK|7|2|他們曾看見他的門徒中有人用不潔淨的手，就是沒有洗的手吃飯。
MARK|7|3|法利賽人和所有的 猶太 人都拘守古人的傳統，若不按規矩洗手就不吃飯；
MARK|7|4|從市場來，若不洗淨也不吃飯；他們還拘守好些別的規矩，如洗杯、罐、銅器、床鋪 等。
MARK|7|5|法利賽人和文士問他說：「你的門徒為甚麼不照古人的傳統，竟然用不潔淨的手吃飯呢？」
MARK|7|6|耶穌對他們說：「 以賽亞 指著你們假冒為善的人所預言的說得好。如經上所記： 『這百姓用嘴唇尊敬我， 他們的心卻遠離我。
MARK|7|7|他們把人的規條當作教義教導人； 他們拜我也是枉然。』
MARK|7|8|你們是離棄上帝的誡命，拘守人的傳統。」
MARK|7|9|耶穌又說：「你們誠然是廢棄上帝的誡命，為要守自己的傳統。
MARK|7|10|摩西 說：『當孝敬父母』；又說：『咒罵父母的，必須處死。』
MARK|7|11|你們倒說：『人若對父母說：我所當供奉你的已經作了各耳板』（各耳板就是奉獻的意思），
MARK|7|12|你們就容許他不必再奉養父母。
MARK|7|13|這就是你們藉著繼承傳統，廢了上帝的話。你們還做許多這樣的事。」
MARK|7|14|耶穌又叫眾人來，對他們說：「你們都要聽我的話，也要明白。
MARK|7|15|從外面進去的不能玷污人，惟有從裏面出來的才玷污人。 」
MARK|7|16|
MARK|7|17|耶穌離開眾人，進了屋子，門徒就問他這比喻的意思。
MARK|7|18|耶穌對他們說：「你們也是這樣不明白嗎？難道你們不了解，凡從外面進去的不能玷污人嗎？
MARK|7|19|因為不是進入他的心，而是進入他的肚子，又排入廁所。」（這是說，各樣的食物都是潔淨的。）
MARK|7|20|耶穌又說：「從人裏面出來的，那才玷污人；
MARK|7|21|因為從人心裏發出種種惡念，如淫亂、偷盜、兇殺、
MARK|7|22|姦淫、貪婪、邪惡、詭詐、淫蕩、嫉妒、毀謗、驕傲、狂妄。
MARK|7|23|這一切的惡都是從裏面出來，且能玷污人。」
MARK|7|24|耶穌從那裏起身，往 推羅 境內去，進了一家，他不願意人知道，卻隱藏不住。
MARK|7|25|立刻有一個婦人，她的小女兒被污靈附著，一聽見耶穌的事，就來俯伏在他腳前。
MARK|7|26|這婦人是 希臘 人，屬 敘利亞 的 腓尼基 族。她求耶穌從她女兒身上趕出那鬼。
MARK|7|27|耶穌對她說：「讓孩子們先吃飽，拿孩子的餅丟給小狗吃是不妥的。」
MARK|7|28|婦人回答：「主啊，桌子底下的小狗也吃小孩子的碎屑呀！」
MARK|7|29|耶穌對她說：「憑著這句話，你回去吧，鬼已經離開你的女兒了。」
MARK|7|30|她就回家去，見小孩子躺在床上，鬼已經出去了。
MARK|7|31|耶穌又離開了 推羅 地區，經過 西頓 ，就從 低加坡里 境內來到 加利利海 。
MARK|7|32|有人帶著一個耳聾舌結的人來見耶穌，求他為他按手。
MARK|7|33|耶穌領他離開眾人，到一邊去，就用指頭探他的耳朵，吐唾沫抹他的舌頭，
MARK|7|34|望天嘆息，對他說：「以法大！」就是說「開了吧！」
MARK|7|35|他的耳朵立刻 開了，舌結也解了，他說話也清楚了。
MARK|7|36|耶穌囑咐他們不要告訴人；但他越囑咐，他們越發傳揚。
MARK|7|37|眾人分外驚奇，說：「他所做的事樣樣都好，他甚至使聾子聽見，啞巴說話。」
MARK|8|1|那時，又有一大群人聚集，沒有甚麼吃的。耶穌叫門徒來，說：
MARK|8|2|「我憐憫這群人，因為他們同我在這裏已經三天，沒有吃的東西了。
MARK|8|3|我若叫他們餓著回家，他們會在路上餓昏，因為其中有從遠處來的。」
MARK|8|4|門徒回答：「在這野地，從哪裏能得餅使這些人吃飽呢？」
MARK|8|5|耶穌問他們：「你們有多少餅？」他們說：「七個。」
MARK|8|6|他吩咐眾人坐在地上，就拿著這七個餅祝謝了，擘開，遞給門徒，叫他們擺開，門徒就擺在眾人面前。
MARK|8|7|他們還有幾條小魚；耶穌祝謝了，就吩咐也擺在眾人面前。
MARK|8|8|他們都吃，並且吃飽了，收拾剩下的碎屑，有七筐子。
MARK|8|9|人數約有四千。耶穌打發他們走了，
MARK|8|10|隨即同門徒上船，來到 大瑪努他 境內。
MARK|8|11|法利賽人出來盤問耶穌，要求他從天上顯個神蹟給他們看，想要試探他。
MARK|8|12|耶穌心裏深深嘆息，說：「這世代為甚麼求神蹟呢？我實在告訴你們，沒有神蹟給這世代看。」
MARK|8|13|他就離開他們，又上船往海的對岸去了。
MARK|8|14|門徒忘了帶餅，在船上除了一個餅，沒有別的食物。
MARK|8|15|耶穌囑咐他們說：「你們要謹慎，要防備法利賽人的酵和 希律 的酵。」
MARK|8|16|他們彼此議論說：「這是因為我們沒有餅吧。」
MARK|8|17|耶穌知道了，就說：「你們為甚麼因為沒有餅就議論呢？你們還不領悟，還不明白嗎？你們的心還是愚頑嗎？
MARK|8|18|你們有眼睛，看不見嗎？有耳朵，聽不到嗎？也不記得嗎？
MARK|8|19|我擘開那五個餅分給五千人，你們收拾的碎屑裝滿了多少個籃子呢？」他們說：「十二個。」
MARK|8|20|「又擘開那七個餅分給四千人，你們收拾的碎屑裝滿了多少個筐子呢？」他們說：「七個。」
MARK|8|21|耶穌說：「你們還不明白嗎？」
MARK|8|22|他們來到 伯賽大 ，有人帶一個盲人來，求耶穌摸他。
MARK|8|23|耶穌拉著盲人的手，領他到村外，就吐唾沫在他眼睛上，為他按手，問他：「你看見甚麼？」
MARK|8|24|他抬頭一看，說：「我看見人，他們好像樹木，並且行走。」
MARK|8|25|隨後耶穌又按手在他眼睛上，他定睛一看，就復原了，樣樣都看得清楚了。
MARK|8|26|耶穌打發他回家，說：「連這村子你也不要進去。」
MARK|8|27|耶穌和門徒出去，往 凱撒利亞．腓立比 附近的村莊去。在路上，他問門徒：「人們說我是誰？」
MARK|8|28|他們對他說：「是施洗的 約翰 ；有人說是 以利亞 ；又有人說是先知中的一位。」
MARK|8|29|他又問他們：「你們說我是誰？」 彼得 回答他：「你是基督。」
MARK|8|30|於是耶穌切切地囑咐他們不可對任何人說起他。
MARK|8|31|從此，他教導他們說：「人子必須受許多的苦，被長老、祭司長和文士棄絕，並且被殺，三天後復活。」
MARK|8|32|耶穌明白地說了這話， 彼得 就拉著他，責備他。
MARK|8|33|耶穌轉過來看著門徒，斥責 彼得 說：「撒但，退到我後邊去！因為你不體會上帝的心意，而是體會人的意思。」
MARK|8|34|於是他叫眾人和門徒來，對他們說：「若有人要跟從我，就當捨己，背起自己的十字架來跟從我。
MARK|8|35|因為凡要救自己生命的，必喪失生命；凡為我和福音喪失生命的，必救自己的生命。
MARK|8|36|人就是賺得全世界，賠上自己的生命，有甚麼益處呢？
MARK|8|37|人還能拿甚麼換生命呢？
MARK|8|38|凡在這淫亂罪惡的世代，把我和我的道當作可恥的，人子在他父的榮耀裏與聖天使一同來臨的時候，也要把那人當作可恥的。」
MARK|9|1|耶穌又對他們說：「我實在告訴你們，站在這裏的，有人在沒經歷死亡以前，必定看見上帝的國帶著能力臨到。」
MARK|9|2|過了六天，耶穌帶著 彼得 、 雅各 、 約翰 ，領他們悄悄地上了高山。他在他們面前變了形像，
MARK|9|3|衣服放光，極其潔白，地上漂布的人沒有一個能漂得那樣白。
MARK|9|4|有 以利亞 和 摩西 向他們顯現，並且與耶穌說話。
MARK|9|5|彼得 對耶穌說：「拉比 ，我們在這裏真好！我們來搭三座棚，一座為你，一座為 摩西 ，一座為 以利亞 。」
MARK|9|6|彼得 不知道說甚麼才好，因為他們很害怕。
MARK|9|7|有一朵雲彩來遮蓋他們，又有聲音從雲彩裏出來，說：「這是我的愛子，你們要聽從他！」
MARK|9|8|門徒連忙向周圍觀看，不再看見任何人，只見耶穌同他們在一起。
MARK|9|9|下山的時候，耶穌囑咐他們說：「人子還沒有從死人中復活，你們不要把所看到的告訴人。」
MARK|9|10|門徒將這話存記在心，彼此議論「從死人中復活」是甚麼意思。
MARK|9|11|他們就問耶穌：「文士為甚麼說 以利亞 必須先來？」
MARK|9|12|耶穌說：「 以利亞 的確先來復興萬事。經上不是指著人子說，他要受許多的苦和被人輕慢嗎？
MARK|9|13|我告訴你們， 以利亞 已經來了，他們任意待他，正如經上指著他說的。」
MARK|9|14|他們到了門徒那裏，看見有一大群人圍著他們，又有文士和他們辯論。
MARK|9|15|眾人一見耶穌，都很驚奇，就跑上去向他問安。
MARK|9|16|耶穌問他們：「你們和他們辯論甚麼？」
MARK|9|17|眾人中的一個回答：「老師，我帶了我的兒子到你這裏來，他被啞巴的靈附著。
MARK|9|18|無論在哪裏，那靈拿住他，把他摔倒，他就口吐白沫，牙關緊鎖，身體僵硬。我請過你的門徒把那靈趕出去，他們卻不能。」
MARK|9|19|耶穌回答：「唉！這不信的世代啊，我和你們在一起要到幾時呢？我忍耐你們要到幾時呢？把他帶到我這裏！」
MARK|9|20|他們就帶了他來。那靈一見耶穌，就使他重重地抽風，倒在地上，翻來覆去，口吐白沫。
MARK|9|21|耶穌問他父親：「他得這病有多久了呢？」父親說：「從小的時候。
MARK|9|22|那靈屢次把他扔在火裏、水裏，要治死他。你若能做甚麼，求你憐憫我們，幫助我們。」
MARK|9|23|耶穌對他說：「『你若能』，在信的人，凡事都能。」
MARK|9|24|孩子的父親立刻喊著說：「我信；求你幫助我的不信！」
MARK|9|25|耶穌看見眾人都跑上來，就斥責那污靈說：「你這聾啞的靈，我命令你從他裏頭出來，再不要進去！」
MARK|9|26|那靈大喊一聲，使孩子猛烈地抽了一陣風，就出來了。孩子好像死了一般，以致眾人多半說：「他死了。」
MARK|9|27|但耶穌拉著他的手，扶他起來，他就站起來了。
MARK|9|28|耶穌進了屋子，門徒就私下問他：「我們為甚麼不能趕出那靈呢？」
MARK|9|29|耶穌對他們說：「非用禱告 ，這一類的邪靈總趕不出來。」
MARK|9|30|他們離開那地方，經過 加利利 ；耶穌不願意人知道，
MARK|9|31|因為他正教導門徒說：「人子將要被交在人手裏，他們要殺害他；被殺以後，三天後他要復活。」
MARK|9|32|門徒卻不明白這話，又不敢問他。
MARK|9|33|他們來到 迦百農 。耶穌在屋裏問門徒說：「你們在路上議論的是甚麼？」
MARK|9|34|門徒不作聲，因為他們在路上彼此爭論誰最大。
MARK|9|35|耶穌坐下，叫十二個使徒來，說：「若有人願意為首，他要作眾人之後，作眾人的用人。」
MARK|9|36|於是耶穌領一個小孩過來，讓他站在門徒當中，又抱起他來，對他們說：
MARK|9|37|「凡為我的名接納一個像這小孩子的，就是接納我；凡接納我的，不是接納我，而是接納那差我來的。」
MARK|9|38|約翰 對耶穌說：「老師，我們看見一個人奉你的名趕鬼，我們就阻止他，因為他不跟從我們。」
MARK|9|39|耶穌說：「不要阻止他，因為沒有人奉我的名行異能，反倒輕易毀謗我。
MARK|9|40|不抵擋我們的，就是幫助我們的。
MARK|9|41|凡因你們是屬基督，給你們一杯水喝的，我實在告訴你們，他一定會得到賞賜。」
MARK|9|42|「凡使這些信我的小子 中的一個跌倒的，倒不如把大磨石拴在這人的頸項上，扔在海裏。
MARK|9|43|如果你一隻手使你跌倒，就把它砍下來；你缺一隻手進入永生，比有兩隻手落到地獄，入那不滅的火裏去還好。
MARK|9|44|
MARK|9|45|如果你一隻腳使你跌倒，就把它砍下來；你瘸腿進入永生，比有兩隻腳被扔進地獄裏還好。
MARK|9|46|
MARK|9|47|如果你一隻眼使你跌倒，就去掉它；你只有一隻眼進入上帝的國，比有兩隻眼被扔進地獄裏還好。
MARK|9|48|在那裏，蟲是不死的，火是不滅的。
MARK|9|49|因為每個人必被火像鹽一般醃起來。
MARK|9|50|鹽本是好的，若失了鹹味，你們怎能用它調味呢？你們中間要有鹽，彼此和睦。」
MARK|10|1|耶穌從那裏起身，來到 猶太 的境內， 約旦河 的東邊。眾人又聚集到他那裏，他又照常教導他們。
MARK|10|2|有法利賽人來問他說：「男人休妻合不合法？」意思是要試探他。
MARK|10|3|耶穌回答他們說：「 摩西 吩咐你們的是甚麼？」
MARK|10|4|他們說：「 摩西 准許寫了休書就可以休妻。」
MARK|10|5|耶穌對他們說：「 摩西 因為你們的心硬，所以寫這誡命給你們。
MARK|10|6|但從起初創造的時候，上帝造人是造男造女。
MARK|10|7|因此，人要離開他的父母，與妻子結合 ，
MARK|10|8|二人成為一體。既然如此，夫妻不再是兩個人，而是一體的了。
MARK|10|9|所以，上帝配合的，人不可分開。」
MARK|10|10|他們到了屋裏，門徒又問他這事。
MARK|10|11|耶穌對他們說：「凡休妻另娶的，就是犯姦淫，辜負他的妻子；
MARK|10|12|妻子若離棄丈夫另嫁，也是犯姦淫了。」
MARK|10|13|有人帶著小孩子來見耶穌，要他摸他們，門徒就責備那些人。
MARK|10|14|耶穌看見就很生氣，對門徒說：「讓小孩到我這裏來，不要阻止他們，因為在上帝國的正是這樣的人。
MARK|10|15|我實在告訴你們，凡要接受上帝國的，若不像小孩子，絕不能進去。」
MARK|10|16|於是他抱著小孩子，給他們按手，為他們祝福。
MARK|10|17|耶穌剛上路的時候，有一個人跑來，跪在他面前，問他：「善良的老師，我該做甚麼事才能承受永生？」
MARK|10|18|耶穌對他說：「你為甚麼稱我是善良的？除了上帝一位之外，再沒有善良的。
MARK|10|19|誡命你是知道的：『不可殺人；不可姦淫；不可偷盜；不可作假見證；不可虧負人；當孝敬父母。』」
MARK|10|20|他對耶穌說：「老師，這一切我從小都遵守了。」
MARK|10|21|耶穌看著他，就愛他，對他說：「你還缺少一件：去變賣你所有的，分給窮人，就必有財寶在天上；然後來跟從我。」
MARK|10|22|他聽見這話，臉就變了色，憂憂愁愁地走了，因為他的產業很多。
MARK|10|23|耶穌看了看周圍，對門徒說：「有錢財的人進上帝的國是何等的難哪！」
MARK|10|24|門徒對他的話非常驚奇。耶穌又對他們說：「孩子們， 要進上帝的國是何等的難哪！
MARK|10|25|駱駝穿過針眼比財主進上帝的國還容易呢！」
MARK|10|26|門徒就更為驚訝，彼此對問：「這樣，誰能得救呢？」
MARK|10|27|耶穌看著他們，說：「在人不能，在上帝卻不然，因為在上帝凡事都能。」
MARK|10|28|彼得 就對他說：「看哪，我們已經撇下一切跟從你了。」
MARK|10|29|耶穌說：「我實在告訴你們，凡為我和福音撇下房屋，或是兄弟、姊妹、父親、母親、兒女、田地，
MARK|10|30|沒有不在今世得百倍的，就是房屋、兄弟、姊妹、母親、兒女、田地，並且要受迫害，在來世得永生。
MARK|10|31|然而，有許多在前的，將要在後；在後的，將要在前。」
MARK|10|32|他們行路上 耶路撒冷 去。耶穌在前頭走，他們很驚訝，跟從的人也害怕。耶穌又叫十二使徒來，把自己將要遭遇的事告訴他們，
MARK|10|33|說：「看哪，我們上 耶路撒冷 去，人子將被交給祭司長和文士；他們要定他死罪，又交給外邦人。
MARK|10|34|他們要戲弄他，向他吐唾沫，鞭打他，殺害他；三天後，他要復活。」
MARK|10|35|西庇太 的兒子 雅各 和 約翰 進前來，對耶穌說：「老師，我們無論求你甚麼，願你為我們做。」
MARK|10|36|耶穌對他們說：「要我為你們做甚麼？」
MARK|10|37|他們對他說：「在你的榮耀裏，請賜我們一個坐在你右邊，一個坐在你左邊。」
MARK|10|38|耶穌對他們說：「你們不知道所求的是甚麼。我所喝的杯，你們能喝嗎？我所受的洗，你們能受嗎？」
MARK|10|39|他們對他說：「我們能。」耶穌對他們說：「我所喝的杯，你們要喝；我所受的洗，你們也要受。
MARK|10|40|可是坐在我的左右，不是我可以賜的，而是為誰預備就賜給誰。」
MARK|10|41|其餘十個門徒聽見，就對 雅各 和 約翰 很生氣。
MARK|10|42|耶穌叫了他們來，對他們說：「你們知道，外邦人有君王作主治理他們，有大臣操權管轄他們。
MARK|10|43|但是在你們中間，不可這樣。你們中間誰願為大，就要作你們的用人；
MARK|10|44|在你們中間誰願為首，就要作眾人的僕人。
MARK|10|45|因為人子來，並不是要受人的服事，乃是要服事人，並且要捨命作多人的贖價。」
MARK|10|46|他們到了 耶利哥 。耶穌同門徒並許多人離開 耶利哥 的時候，有一個討飯的盲人，是 底買 的兒子 巴底買 ，坐在路旁。
MARK|10|47|他聽見是 拿撒勒 的耶穌，就喊了起來，說：「 大衛 之子耶穌啊，可憐我吧！」
MARK|10|48|有許多人責備他，不許他作聲，他卻越發喊著：「 大衛 之子啊，可憐我吧！」
MARK|10|49|耶穌就站住，說：「叫他過來。」他們就叫那盲人，對他說：「放心，起來！他在叫你啦。」
MARK|10|50|盲人就丟下衣服，跳起來，走到耶穌那裏。
MARK|10|51|耶穌回答他說：「你要我為你做甚麼？」盲人對他說：「拉波尼 ，我要能看見。」
MARK|10|52|耶穌對他說：「你去吧！你的信救了你。」盲人立刻看得見，就在路上跟隨耶穌。
MARK|11|1|耶穌和門徒快到 耶路撒冷 ，來到 伯法其 和 伯大尼 ，在 橄欖山 那裏。耶穌打發兩個門徒，
MARK|11|2|對他們說：「你們往對面村子裏去，一進去的時候會看見一匹驢駒拴在那裏，是從來沒有人騎過的，把牠解開，牽來。
MARK|11|3|若有人對你們說：『為甚麼做這事？』你們就說：『主要用牠，但會立刻把牠牽回到這裏來。』」
MARK|11|4|他們去了，看見一匹驢駒拴在門外街道上，就把牠解開。
MARK|11|5|在那裏站著的人，有幾個說：「你們解開驢駒做甚麼？」
MARK|11|6|門徒照著耶穌的話說，那些人就任憑他們牽去了。
MARK|11|7|他們把驢駒牽到耶穌那裏，把自己的衣服搭在上面，耶穌就騎上。
MARK|11|8|有許多人把衣服鋪在路上，還有人把田間的樹枝砍下來鋪上。
MARK|11|9|前呼後擁的人都喊著說： 「和散那 ！ 奉主名來的是應當稱頌的！
MARK|11|10|那將要來的我祖 大衛 之國是應當稱頌的！ 至高無上的，和散那！」
MARK|11|11|耶穌到了 耶路撒冷 ，進入聖殿，看了周圍的一切。天色已晚，他就和十二使徒出城，往 伯大尼 去。
MARK|11|12|第二天，他們從 伯大尼 出來，耶穌餓了。
MARK|11|13|他遠遠地看見一棵無花果樹，樹上有葉子，就過去，看是不是在樹上可以找到甚麼。他到了樹下，竟找不到甚麼，只有葉子，因為不是無花果的季節。
MARK|11|14|耶穌就對樹說：「從今以後，永沒有人吃你的果子。」他的門徒都聽到了。
MARK|11|15|他們來到 耶路撒冷 。耶穌一進聖殿，就趕出在聖殿裏做買賣的人，推倒兌換銀錢之人的桌子和賣鴿子之人的凳子；
MARK|11|16|也不許人拿著器具從聖殿裏經過。
MARK|11|17|他教導他們說：「經上不是記著： 『我的殿要稱為萬國禱告的殿嗎？ 你們倒使它成為賊窩了。』」
MARK|11|18|祭司長和文士聽見這話，就想法子要除掉耶穌，卻又怕他，因為眾人都對他的教導感到驚奇。
MARK|11|19|每天晚上，他們 都到城外去。
MARK|11|20|早晨，他們從那裏經過，看見無花果樹連根都枯乾了。
MARK|11|21|彼得 想起耶穌的話來，就對他說：「拉比，你看！你所詛咒的無花果樹已經枯乾了。」
MARK|11|22|耶穌回答：「你們對上帝要有信心。
MARK|11|23|我實在告訴你們，無論何人對這座山說：『離開此地，投在海裏！』他心裏若不疑惑，只信所說的必成，就為他實現。
MARK|11|24|所以我告訴你們，凡你們禱告祈求的，無論是甚麼，只要信你們已經得著了，就為你們實現。
MARK|11|25|你們站著禱告的時候，若想起有人得罪你們，就該饒恕他，好讓你們在天上的父也饒恕你們的過犯。 」
MARK|11|26|
MARK|11|27|他們又來到 耶路撒冷 。耶穌在聖殿裏行走的時候，祭司長、文士和長老進前來，
MARK|11|28|問他說：「你仗著甚麼權柄做這些事？給你權柄做這些事的是誰呢？」
MARK|11|29|耶穌對他們說：「我要問你們一句話，你們回答我，我就告訴你們我仗著甚麼權柄做這些事。
MARK|11|30|約翰 的洗禮是從天上來的，還是從人間來的呢？你們回答我吧。」
MARK|11|31|他們彼此商議說：「我們若說『從天上來的』，他會說：『這樣，你們為甚麼不信他呢？』
MARK|11|32|但若說『從人間來的』，卻又怕眾人，因為大家認為 約翰 確是先知。」
MARK|11|33|於是他們回答耶穌：「我們不知道。」耶穌說：「我也不告訴你們，我仗著甚麼權柄做這些事。」
MARK|12|1|耶穌就用比喻對他們說：「有人開墾了一個葡萄園，四周圍上籬笆，挖了一個榨酒池，蓋了一座守望樓，租給園戶，就出外遠行去了。
MARK|12|2|到了時候，他打發一個僕人到園戶那裏，要向他們收葡萄園的果子。
MARK|12|3|他們拿住他，打了他，叫他空手回去。
MARK|12|4|園主再打發一個僕人到他們那裏。他們打傷他的頭，並且侮辱他。
MARK|12|5|園主又打發一個僕人去，他們就殺了他。以後又打發好些僕人去，有的被他們打了，有的被他們殺了。
MARK|12|6|園主還有一位，是他的愛子，最後又打發他去，說：『他們會尊敬我的兒子。』
MARK|12|7|那些園戶卻彼此說：『這是承受產業的。來，我們殺了他，產業就歸我們了！』
MARK|12|8|於是他們拿住他，殺了他，把他扔出葡萄園。
MARK|12|9|這樣，葡萄園主要怎麼做呢？他要來除滅那些園戶，將葡萄園轉給別人。
MARK|12|10|『匠人所丟棄的石頭 已作了房角的頭塊石頭。 這是主所做的， 在我們眼中看為奇妙。』 這經文你們沒有念過嗎？」
MARK|12|11|
MARK|12|12|他們看出這比喻是指著他們說的，就想要捉拿他，但是懼怕眾人，於是離開他走了。
MARK|12|13|後來，他們打發幾個法利賽人和 希律 黨人到耶穌那裏，要用他自己的話陷害他。
MARK|12|14|他們來了，就對他說：「老師，我們知道你是誠實的，無論誰你都一視同仁；因為你不看人的面子，而是誠誠實實傳上帝的道。納稅給凱撒合不合法？
MARK|12|15|我們該不該納？」耶穌知道他們的虛偽，就對他們說：「你們為甚麼試探我？拿一個銀幣來給我看。」
MARK|12|16|他們就拿了來。耶穌問他們：「這像和這名號是誰的？」他們對他說：「是凱撒的。」
MARK|12|17|耶穌對他們說：「凱撒的歸凱撒；上帝的歸上帝。」他們對他非常驚訝。
MARK|12|18|撒都該人來見耶穌。他們說沒有復活這回事，於是問耶穌：
MARK|12|19|「老師， 摩西 為我們寫下這話：『某人的哥哥若死了，撇下妻子，沒有孩子，他該娶哥哥的妻子，為哥哥生子立後。』
MARK|12|20|那麼，有兄弟七人，第一個娶了妻，死了，沒有留下孩子。
MARK|12|21|第二個娶了她，也死了，沒有留下孩子。第三個也是這樣。
MARK|12|22|那七個人都沒有留下孩子。最後，那婦人也死了。
MARK|12|23|在復活的時候， 她是哪一個的妻子呢？因為他們七個人都娶過她。」
MARK|12|24|耶穌說：「你們錯了，不正是因為不明白聖經，也不知道上帝的大能嗎？
MARK|12|25|當人從死人中復活後，也不娶也不嫁，而是像天上的天使一樣。
MARK|12|26|論到死人復活，你們沒有念過 摩西 書中《荊棘篇》上所記載的嗎？上帝對 摩西 說：『我是 亞伯拉罕 的上帝， 以撒 的上帝， 雅各 的上帝。』
MARK|12|27|上帝不是死人的上帝，而是活人的上帝。你們是大錯了。」
MARK|12|28|有一個文士來，聽見他們的辯論，知道耶穌回答得好，就問他說：「誡命中哪一條是第一呢？」
MARK|12|29|耶穌回答：「第一是：『 以色列 啊，你要聽，主—我們的上帝是獨一的主。
MARK|12|30|你要盡心、盡性、盡意、盡力愛主—你的上帝。』
MARK|12|31|第二是：『要愛鄰 如己。』再沒有比這兩條誡命更大的了。」
MARK|12|32|那文士對耶穌說：「好，老師，你說得對，上帝是一位，除了他以外，再沒有別的了；
MARK|12|33|並且盡心、盡智、盡力愛他，又愛鄰如己，要比一切燔祭和祭祀好得多。」
MARK|12|34|耶穌見他回答得有智慧，就對他說：「你離上帝的國不遠了。」從此以後，沒有人敢再問他甚麼。
MARK|12|35|耶穌在聖殿裏教導人，問他們說：「文士怎麼說基督是 大衛 的後裔呢？
MARK|12|36|大衛 被聖靈感動，說： 『主對我主說： 你坐在我的右邊， 等我把你的仇敵放在你腳下 。』
MARK|12|37|大衛 親自稱他為主，他怎麼又是 大衛 的後裔呢？」一大群的人都喜歡聽他。
MARK|12|38|他在教導的時候，說：「你們要防備文士。他們好穿長袍走來走去，喜歡人們在街市上向他們問安，
MARK|12|39|又喜愛會堂裏的高位，宴席上的首座。
MARK|12|40|他們侵吞寡婦的家產，假意作很長的禱告。這些人要受更重的懲罰！」
MARK|12|41|耶穌面向聖殿銀庫坐著，看眾人怎樣把錢投入銀庫。有好些財主投了許多錢。
MARK|12|42|有一個窮寡婦來，投了兩個小文錢 ，就是一個大文錢 。
MARK|12|43|耶穌叫門徒來，對他們說：「我實在告訴你們，這窮寡婦投入銀庫裏的比眾人所投的更多。
MARK|12|44|因為，眾人都是拿有餘的捐獻，但這寡婦，雖然自己不足，卻把她一生所有的全都投進去了。」
MARK|13|1|耶穌從聖殿裏出來的時候，有一個門徒對他說：「老師，請看，這是多麼了不起的石頭！多麼了不起的建築！」
MARK|13|2|耶穌對他說：「你看見這些宏偉的建築嗎？這裏將沒有一塊石頭會留在另一塊石頭上而不被拆毀的。」
MARK|13|3|耶穌在 橄欖山 上，面向聖殿坐著； 彼得 、 雅各 、 約翰 和 安得烈 私下問他說：
MARK|13|4|「請告訴我們，甚麼時候有這些事呢？這一切事將成的時候有甚麼預兆呢？」
MARK|13|5|耶穌說：「你們要謹慎，免得有人迷惑你們。
MARK|13|6|將有好些人冒我的名來，說『我是基督』，並且要迷惑許多人。
MARK|13|7|當你們聽見打仗和打仗的風聲，不要驚慌；這些事必須發生，但這還不是終結。
MARK|13|8|民要攻打民，國要攻打國，多處必有地震、饑荒。這都是災難 的起頭。
MARK|13|9|但你們自己要謹慎；因為有人要把你們交給議會，並且你們在會堂裏要受鞭打，又為我的緣故站在統治者和君王面前，對他們作見證。
MARK|13|10|然而，福音必須先傳給萬民。
MARK|13|11|有人把你們解送去受審的時候，不要事先擔心說甚麼；到那時候，賜給你們甚麼話，你們就說甚麼；因為說話的不是你們，而是聖靈。
MARK|13|12|兄弟要把兄弟、父親要把兒女置於死地；兒女要起來與父母為敵，害死他們；
MARK|13|13|而且你們要為我的名被眾人憎恨。但堅忍到底的終必得救。」
MARK|13|14|「當你們看見那『施行毀滅的褻瀆者』站在不當站的地方（讀這經的人要會意），那時，在 猶太 的，應當逃到山上；
MARK|13|15|在屋頂上的，不要下來，也不要進家裏去拿東西；
MARK|13|16|在田裏的，不要回去取衣裳。
MARK|13|17|在那些日子，懷孕的和奶孩子的就苦了。
MARK|13|18|你們要祈求，叫這事不在冬天發生。
MARK|13|19|因為，在那些日子必有災難，自從上帝創造萬物直到如今，從沒有這樣的災難，將來也不會有。
MARK|13|20|若不是主減少那些日子，凡血肉之軀的，就沒有一個能得救；但是為了他所揀選的選民，他將那些日子減少了。
MARK|13|21|那時，若有人對你們說：『看哪，基督在這裏！看哪，在那裏！』你們不要信。
MARK|13|22|因為假基督和假先知將要起來，顯神蹟奇事，如果可能，連選民也迷惑了。
MARK|13|23|你們要謹慎！凡事我都預先告訴你們了。」
MARK|13|24|「在那些日子、那災難以後， 太陽要變黑，月亮也不放光，
MARK|13|25|眾星要從天上墜落， 天上的萬象都要震動。
MARK|13|26|那時，他們要看見人子帶著大能力和榮耀駕雲來臨。
MARK|13|27|他要差遣天使，從四方，從地極直到天邊，召集他的選民。」
MARK|13|28|「你們要從無花果樹學習功課：當樹枝發芽長葉的時候，你們就知道夏天近了。
MARK|13|29|同樣，當你們看見這些事發生，就知道那時候近了，就在門口了。
MARK|13|30|我實在告訴你們，這世代還沒有過去，這一切都要發生。
MARK|13|31|天地要廢去，我的話卻絕不廢去。」
MARK|13|32|「但那日子，那時辰，沒有人知道，連天上的天使也不知道，子也不知道，惟有父知道。
MARK|13|33|你們要謹慎，要警醒 ，因為你們不知道那時刻幾時來到。
MARK|13|34|這事正如一個人離家遠行，授權給僕人們，分派各人的工作，又吩咐看門的警醒。
MARK|13|35|所以，你們要警醒，因為你們不知道這家的主人甚麼時候來，是晚上，或半夜，或雞叫時，或早晨，
MARK|13|36|免得他忽然來到，看見你們睡著了。
MARK|13|37|我對你們所說的話，也是對眾人說的：要警醒！」
MARK|14|1|過兩天是逾越節，又是除酵節，祭司長和文士在想法子怎樣設計捉拿耶穌，把他殺掉。
MARK|14|2|他們說：「不可在過節的日子，恐怕百姓生亂。」
MARK|14|3|耶穌在 伯大尼 痲瘋病人 西門 家裏坐席的時候，有一個女人拿著一玉瓶極貴的純哪噠 香膏來，打破玉瓶，把膏澆在耶穌的頭上。
MARK|14|4|有幾個人心中很不高興，說：「何必這樣浪費香膏呢？
MARK|14|5|這香膏可以賣三百多個銀幣賙濟窮人。」他們就對那女人生氣。
MARK|14|6|耶穌說：「由她吧！為甚麼難為她呢？她在我身上做的是一件美事。
MARK|14|7|因為常有窮人和你們在一起，要向他們行善，隨時都可以，但是你們不常有我。
MARK|14|8|她所做的是盡她所能的；她是為了我的安葬，把香膏預先澆在我身上。
MARK|14|9|我實在告訴你們，普天之下，無論在甚麼地方傳這福音，都要述說這女人所做的，來記念她。」
MARK|14|10|十二使徒中有一個 加略 人 猶大 ，去見祭司長，要把耶穌交給他們。
MARK|14|11|他們聽見就很高興，又應許給他銀子；他就想怎樣找機會把耶穌交給他們。
MARK|14|12|除酵節的第一天，就是宰逾越節羔羊的那一天，門徒對耶穌說：「你要我們到哪裏去預備你吃逾越節的宴席呢？」
MARK|14|13|耶穌就打發兩個門徒，對他們說：「你們進城去，會有人拿著一罐水迎面而來，你們就跟著他。
MARK|14|14|無論他進哪一家，你們就對那家的主人說：『老師問：我的客房在哪裏？我和我的門徒要在那裏吃逾越節的宴席。』
MARK|14|15|他會帶你們看一間擺設齊全、準備妥當的樓上大廳，你們就在那裏為我們預備。」
MARK|14|16|門徒出去，進了城，所看到的正如耶穌所說的。他們就預備了逾越節的宴席。
MARK|14|17|到了晚上，耶穌和十二使徒都來了。
MARK|14|18|他們坐席，正吃的時候，耶穌說：「我實在告訴你們，你們中間有一個與我同吃的人要出賣我了。」
MARK|14|19|他們就憂愁起來，一個個地問他：「不是我吧？」
MARK|14|20|耶穌對他們說：「是十二人中的一個，就是同我蘸餅在盤子裏的那個人。
MARK|14|21|人子要去了，正如經上所寫有關他的；但出賣人子的人有禍了！那人沒有出生倒好。」
MARK|14|22|他們吃的時候，耶穌拿起餅來，祝福了，就擘開，遞給他們，說：「你們拿去，這是我的身體。」
MARK|14|23|他又拿起杯來，祝謝了，遞給他們；他們都喝了。
MARK|14|24|耶穌對他們說：「這是我立約的血，為許多人流出來的。
MARK|14|25|我實在告訴你們，我不再喝這葡萄汁，直到我在上帝的國裏喝新的那日子。」
MARK|14|26|他們唱了詩，就出來往 橄欖山 去。
MARK|14|27|耶穌對他們說：「你們都要跌倒，因為經上記著： 『我要擊打牧人， 羊就分散了。』，　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　
MARK|14|28|但我復活以後，要在你們之前往 加利利 去。」
MARK|14|29|彼得 說：「雖然眾人跌倒，但我不會。」
MARK|14|30|耶穌對他說：「我實在告訴你，今天夜裏，雞叫兩遍 以前，你要三次不認我。」
MARK|14|31|彼得 卻極力地說：「我就是必須和你同死，也絕不會不認你。」所有的門徒 都是這樣說。
MARK|14|32|他們來到一個地方，名叫 客西馬尼 。耶穌對門徒說：「你們坐在這裏，我去禱告。」
MARK|14|33|於是他帶著 彼得 、 雅各 和 約翰 同去。他驚恐起來，極其難過，
MARK|14|34|對他們說：「我心裏非常憂傷，幾乎要死；你們留在這裏，要警醒。」
MARK|14|35|他就稍往前走，俯伏在地，禱告說，如果可能，就叫那時候離開他。
MARK|14|36|他說：「阿爸，父啊！在你凡事都能；求你將這杯撤去。然而，不是照我所願的，而是照你所願的。」
MARK|14|37|耶穌回來，見他們睡著了，就對 彼得 說：「 西門 ，你睡著了嗎？不能警醒一小時嗎？
MARK|14|38|總要警醒禱告，免得陷入試探。你們心靈固然願意，肉體卻軟弱了。」
MARK|14|39|耶穌又去禱告，說的話跟先前一樣。
MARK|14|40|他又來，見他們睡著了，因為他們的眼睛很困倦；他們也不知道怎麼回答他。
MARK|14|41|他第三次來對他們說：「現在你們仍在睡覺安歇嗎？夠了，時候到了。看哪，人子被出賣在罪人手裏了。
MARK|14|42|起來，我們走吧！看哪，那出賣我的人快來了。」
MARK|14|43|耶穌還在說話的時候，忽然十二使徒之一的 猶大 來了，還有一群人帶著刀棒，從祭司長、文士和長老那裏跟他同來。
MARK|14|44|那出賣耶穌的人曾給他們一個暗號，說：「我親誰，誰就是。你們把他抓住，穩妥地帶走。」
MARK|14|45|猶大 來了，隨即到耶穌跟前，說：「拉比」，就跟他親吻。
MARK|14|46|他們就下手抓住他。
MARK|14|47|旁邊站著的人，有一個拔出刀來，把大祭司的僕人砍了一刀，削掉了他一隻耳朵。
MARK|14|48|耶穌回應他們說：「你們帶著刀棒出來拿我，如同拿強盜嗎？
MARK|14|49|我天天教導人，同你們在殿裏，你們並沒有抓我。但這是要應驗經上的話。」
MARK|14|50|門徒都離開他，逃走了。
MARK|14|51|有一個青年光著身子，只披一塊麻布，跟隨耶穌，眾人就抓住他。
MARK|14|52|他卻丟下麻布，赤身逃走了。
MARK|14|53|他們把耶穌帶到大祭司那裏，又有眾祭司長、長老和文士都來一同聚集。
MARK|14|54|彼得 遠遠地跟著耶穌，直到進了大祭司的院子，和警衛一同坐在火邊取暖。
MARK|14|55|祭司長和全議會尋找見證控告耶穌，要處死他，卻找不到實據。
MARK|14|56|因為有好些人作假見證告他，他們的見證又各不相符。
MARK|14|57|又有幾個人站起來，作假見證告他說：
MARK|14|58|「我們聽見他說：『我要拆毀這人手所造的殿，三日內另造一座不是人手所造的。』」
MARK|14|59|就是這樣，他們的見證還是不相符。
MARK|14|60|大祭司起來站在中間，問耶穌說：「這些人作證告你的事，你甚麼都不回答嗎？」
MARK|14|61|耶穌卻不言語，一句也不回答。大祭司又問他：「你是不是基督，那當稱頌者的兒子？」
MARK|14|62|耶穌說：「我是。 你們要看見人子 坐在那權能者的右邊， 駕著天上的雲來臨。」
MARK|14|63|大祭司就撕裂衣服，說：「我們何必再要證人呢？
MARK|14|64|你們已經聽見他這褻瀆的話了。你們的決定如何？」他們都判定他該處死。
MARK|14|65|於是有人開始向他吐唾沫，又蒙著他的臉，用拳頭打他，對他說：「你說預言吧！」警衛把他拉過來，打他耳光。
MARK|14|66|彼得 在下邊院子裏，大祭司的一個使女來了，
MARK|14|67|見 彼得 取暖，就看著他，說：「你素來也是同 拿撒勒 人耶穌一起的。」
MARK|14|68|彼得 卻不承認，說：「我不知道，也不明白你說的是甚麼！」於是他出來，到了前院，雞就叫了 。
MARK|14|69|那使女看見他，又對旁邊站著的人說：「這個人也是他們一夥的。」
MARK|14|70|彼得 又不承認。過了不久，旁邊站著的人又對 彼得 說：「你真是他們一夥的，因為你也是 加利利 人。」
MARK|14|71|彼得 就賭咒發誓說：「我不認得你們說的這個人。」
MARK|14|72|立刻，雞叫了第二遍。 彼得 想起耶穌對他所說的話：「雞叫兩遍以前，你要三次不認我。」他就忍不住哭了。
MARK|15|1|一到早晨，眾祭司長、長老、文士，和全議會的人大家商議，就把耶穌綁著，解去，交給 彼拉多 。
MARK|15|2|彼拉多 問他：「你是 猶太 人的王嗎？」耶穌回答：「是你說的。」
MARK|15|3|祭司長們告他許多的事。
MARK|15|4|彼拉多 又問他：「你看，他們告你這麼多的事，你甚麼都不回答嗎？」
MARK|15|5|耶穌仍不回答，以致 彼拉多 覺得驚訝。
MARK|15|6|每逢這節期， 彼拉多 照眾人所求的，釋放一個囚犯給他們。
MARK|15|7|有一個人名叫 巴拉巴 ，和作亂的人監禁在一起。他們作亂的時候曾殺過人。
MARK|15|8|眾人上去求 彼拉多 照常例給他們辦理。
MARK|15|9|彼拉多 說：「你們要我釋放 猶太 人的王給你們嗎？」
MARK|15|10|他原知道祭司長們是因嫉妒才把耶穌解了來。
MARK|15|11|但是祭司長們煽動眾人，寧可要他釋放 巴拉巴 給他們。
MARK|15|12|彼拉多 又說：「那麼，你們稱為 猶太 人的王的 ，要 我怎麼辦他呢？」
MARK|15|13|他們又再喊著：「把他釘十字架！」
MARK|15|14|彼拉多 說：「為甚麼？他做了甚麼惡事呢？」他們更加喊著：「把他釘十字架！」
MARK|15|15|彼拉多 要討好眾人，就釋放 巴拉巴 給他們，把耶穌鞭打後交給人釘十字架。
MARK|15|16|士兵把耶穌帶進總督府的庭院裏，叫齊了全營的兵。
MARK|15|17|他們給他穿上紫袍，又用荊棘編了冠冕給他戴上，
MARK|15|18|然後向他致敬，說：「萬歲， 猶太 人的王！」
MARK|15|19|他們又拿一根蘆葦稈打他的頭，向他吐唾沫，屈膝拜他。
MARK|15|20|他們戲弄完了，就給他脫了紫袍，又穿上他自己的衣服，帶他出去，要把他釘十字架。
MARK|15|21|有一個 古利奈 人 西門 ，就是 亞歷山大 和 魯孚 的父親，從鄉下來，經過那地方，他們就強迫他同去，好背耶穌的十字架。
MARK|15|22|他們帶耶穌到了一個地方叫 各各他 （翻出來就是「髑髏地」），
MARK|15|23|拿沒藥調和的酒給耶穌，他卻不受。
MARK|15|24|於是他們把他釘在十字架上，抽籤分他的衣服，看誰得甚麼。
MARK|15|25|他們把他釘十字架的時候是上午九點鐘。
MARK|15|26|罪狀牌上寫的是：「 猶太 人的王。」
MARK|15|27|他們又把兩個強盜和他同釘十字架，一個在右邊，一個在左邊。
MARK|15|28|
MARK|15|29|從那裏經過的人譏笑他，搖著頭，說：「哼！你這拆毀殿、三日又建造起來的，
MARK|15|30|救救你自己，從十字架上下來呀！」
MARK|15|31|眾祭司長和文士也這樣嘲笑他，彼此說：「他救了別人，不能救自己。
MARK|15|32|以色列 的王基督，現在從十字架上下來，好讓我們看見就信了呀！」那和他同釘的人也譏諷他。
MARK|15|33|到了正午，全地都黑暗了，直到下午三點鐘。
MARK|15|34|下午三點鐘的時候，耶穌大聲呼喊：「以羅伊！以羅伊！拉馬撒巴各大尼？」（翻出來就是：我的上帝！我的上帝！為甚麼離棄我？）
MARK|15|35|旁邊站著的人，有的聽見就說：「看哪，他叫 以利亞 呢！」
MARK|15|36|有一個人跑去，把海綿蘸滿了醋，綁在蘆葦稈上，送給他喝，說：「且等著，看 以利亞 會不會來把他放下來。」
MARK|15|37|耶穌大喊一聲，氣就斷了。
MARK|15|38|殿的幔子從上到下裂為兩半。
MARK|15|39|對面站著的百夫長看見耶穌這樣斷氣 ，就說：「這人真是上帝的兒子！」
MARK|15|40|還有些婦女遠遠地觀看，其中有 抹大拉 的 馬利亞 ，又有小 雅各 和 約西 的母親 馬利亞 ，並有 撒羅米 ，
MARK|15|41|就是耶穌在 加利利 的時候，跟隨他、服事他的那些人，還有同耶穌上 耶路撒冷 的好些婦女。
MARK|15|42|到了晚上，因為這是預備日，就是安息日的前一日，
MARK|15|43|有 亞利馬太 的 約瑟 前來，他是尊貴的議員，也是盼望著上帝國的，他放膽進去見 彼拉多 ，請求要耶穌的身體。
MARK|15|44|彼拉多 詫異耶穌已經死了，就叫百夫長來，問他耶穌是不是死了很久；
MARK|15|45|既從百夫長得知實情，就把耶穌的身體賜給 約瑟 。
MARK|15|46|約瑟 買了細麻布，把耶穌取下來，用細麻布裹好，安放在巖石中鑿出來的墓穴裏，又滾來一塊石頭擋住墓門。
MARK|15|47|抹大拉 的 馬利亞 和 約西 的母親 馬利亞 都看見安放他的地方。
MARK|16|1|過了安息日， 抹大拉 的 馬利亞 、 雅各 的母親 馬利亞 ，和 撒羅米 ，買了香料，要去膏耶穌的身體。
MARK|16|2|七日的第一日清早，太陽出來後，她們來到墳墓那裏，
MARK|16|3|彼此說：「誰要替我們把石頭從墓門滾開呢？」
MARK|16|4|她們抬頭一看，看見石頭已經滾開了，原來那石頭很大。
MARK|16|5|她們進了墳墓，看見一個年輕人坐在右邊，穿著白袍，就很驚奇。
MARK|16|6|那年輕人對她們說：「不要驚慌！你們尋找那釘十字架的 拿撒勒 人耶穌，他已經復活了，不在這裏。來看安放他的地方。
MARK|16|7|你們去，對他的門徒和 彼得 說：『他要比你們先到 加利利 去，在那裏你們會看見他，正如他從前所告訴你們的。』」
MARK|16|8|於是她們出來，從墳墓那裏逃走，又發抖又驚訝，甚麼也沒有告訴人，因為她們害怕。 〔
MARK|16|9|凡耶穌所吩咐的，她們簡潔地告訴 彼得 和他周圍的人。這些事以後，耶穌親自藉著他的門徒，從東到西，把那神聖、不朽、永遠拯救的福音傳出去。阿們！〕 〔 在七日的第一日清早，耶穌復活了，先向 抹大拉 的 馬利亞 顯現；耶穌曾從她身上趕出七個鬼。
MARK|16|10|她去告訴那向來跟隨耶穌的人；那時他們正哀慟哭泣。
MARK|16|11|他們聽見耶穌活了，被 馬利亞 看見，可是不信。〕 〔
MARK|16|12|這些事以後，門徒中有兩個人往鄉下去；正走著的時候，耶穌以另一種形像向他們顯現。
MARK|16|13|他們去告訴其餘的門徒，那些門徒還是不信。〕 〔
MARK|16|14|後來十一使徒坐席的時候，耶穌向他們顯現，責備他們不信，心裏剛硬，因為他們不信那些在他復活以後看見他的人。
MARK|16|15|他又對他們說：「你們往普天下去，傳福音給萬民 聽。
MARK|16|16|信而受洗的必然得救，不信的必被定罪。
MARK|16|17|信的人將有神蹟隨著他們：就是奉我的名趕鬼；說新方言；
MARK|16|18|手 能拿蛇；若喝了甚麼毒物，也不會受害；手按病人，病人就好了。」〕 〔
MARK|16|19|主耶穌 和他們說完了話以後，被接到天上，坐在上帝的右邊。
MARK|16|20|門徒出去，到處傳福音。主和他們同工，藉著伴隨的神蹟證實所傳的道。 〕
LUKE|1|1|提阿非羅 大人哪，有好些人提筆作書，述說在我們中間所實現的事，是照傳道的人從起初親眼看見又傳給我們的。這些事我從起頭都詳細考察了，我也想按著次序寫給你，
LUKE|1|2|
LUKE|1|3|
LUKE|1|4|要讓你知道所學的道都是確實的。
LUKE|1|5|在 希律 作 猶太 王的時候， 亞比雅 班裏有一個祭司，名叫 撒迦利亞 ；他妻子是 亞倫 的後代，名叫 伊利莎白 。
LUKE|1|6|他們兩人在上帝面前都是義人，遵行主的一切誡命和條例，沒有可指責的。
LUKE|1|7|只是他們沒有孩子，因為 伊利莎白 不生育，兩個人又年紀老邁了。
LUKE|1|8|撒迦利亞 按班次在上帝面前執行祭司的職務，
LUKE|1|9|照祭司的規矩抽籤，進到主的殿裏燒香。
LUKE|1|10|燒香的時候，眾百姓在外面禱告。
LUKE|1|11|有主的一個使者站在香壇的右邊，向他顯現。
LUKE|1|12|撒迦利亞 看見，就驚慌害怕。
LUKE|1|13|天使對他說：「 撒迦利亞 ，不要害怕，因為你的祈禱已經被聽見了。你的妻子 伊利莎白 要給你生一個兒子，你要給他起名叫 約翰 。
LUKE|1|14|你必歡喜快樂；有許多人因他出世也必喜樂。
LUKE|1|15|他在主面前將要為大，淡酒烈酒都不喝，從母腹裏就被聖靈充滿。
LUKE|1|16|他要使許多 以色列 人回轉，歸於主—他們的上帝。
LUKE|1|17|他將有 以利亞 的精神和能力，走在主的前面，叫父親的心轉向兒女，叫悖逆的人轉向義人的智慧，又為主預備迎接他的百姓。」
LUKE|1|18|撒迦利亞 對天使說：「我怎麼能知道這事呢？我已經老了，我的妻子也年紀老邁了。」
LUKE|1|19|天使回答他說：「我是站在上帝面前的 加百列 ，奉差遣來對你說話，把這好信息報給你。
LUKE|1|20|到了時候，這些話必然應驗；只因你不信我的話，你會成為啞巴，不能說話，直到這些事實現的日子。」
LUKE|1|21|百姓等候 撒迦利亞 ，詫異他在聖所裏遲延那麼久。
LUKE|1|22|到他出來，卻不能和他們說話，他們就知道他在聖所裏見了異象；他直向他們打手勢，因為他成了啞巴。
LUKE|1|23|他供職的日子一滿，就回家去了。
LUKE|1|24|這些日子以後，他的妻子 伊利莎白 就懷孕，隱藏了五個月；
LUKE|1|25|她說：「主在眷顧我的日子，這樣看顧我，要除掉我在人前的羞恥。」
LUKE|1|26|到了第六個月，天使 加百列 奉上帝的差遣往 加利利 的一座城去，這城名叫 拿撒勒 ，
LUKE|1|27|到一個童女那裏，她已經許配 大衛 家的一個人，名叫 約瑟 ；童女的名字叫 馬利亞 。
LUKE|1|28|天使進去，對她說：「蒙大恩的女子，你好，主和你同在！」
LUKE|1|29|馬利亞 因這話就很驚慌，又反覆思考這樣問候是甚麼意思。
LUKE|1|30|天使對她說： 「 馬利亞 ，不要怕，你在上帝面前已經蒙恩了。
LUKE|1|31|你要懷孕生子，要給他起名叫耶穌。
LUKE|1|32|他將要為大，稱為至高者的兒子； 主上帝要把他祖先 大衛 的王位給他。
LUKE|1|33|他要作 雅各 家的王，直到永遠； 他的國沒有窮盡。」
LUKE|1|34|馬利亞 對天使說：「我沒有出嫁，怎麼會有這事呢？」
LUKE|1|35|天使回答她說： 「聖靈要臨到你身上； 至高者的能力要庇蔭你， 因此，那要出生的聖者要稱為上帝的兒子 。
LUKE|1|36|況且，你的親戚 伊利莎白 ，就是那素來稱為不生育的，在年老的時候也懷了男胎，現在懷孕六個月了。
LUKE|1|37|因為，出於上帝的話，沒有一句不帶能力的。」
LUKE|1|38|馬利亞 說：「我是主的使女，願意照你的話實現在我身上。」於是天使離開她去了。
LUKE|1|39|在那些日子， 馬利亞 起身，急忙前往山區，來到 猶大 的一座城，
LUKE|1|40|進了 撒迦利亞 的家，向 伊利莎白 問安。
LUKE|1|41|伊利莎白 一聽到 馬利亞 問安，所懷的胎就在腹裏跳動。 伊利莎白 被聖靈充滿，
LUKE|1|42|高聲喊著說： 「你在婦女中是有福的！ 你所懷的胎也是有福的！
LUKE|1|43|我主的母親到我這裏來，為何這事臨到我呢？
LUKE|1|44|因為你問安的聲音一入我耳，我腹裏的胎就歡喜跳動。
LUKE|1|45|這相信的女子是有福的！因為主對她所說的話都要應驗。」
LUKE|1|46|馬利亞 說： 「我心尊主為大；
LUKE|1|47|我靈以上帝我的救主為樂；
LUKE|1|48|因為他顧念他使女的卑微； 從今以後，萬代要稱我有福。
LUKE|1|49|因為那有權能的為我做了大事； 他的名是聖的。
LUKE|1|50|他憐憫敬畏他的人， 直到世世代代。
LUKE|1|51|他用膀臂施展大能； 他趕散心裏妄想的狂傲人。
LUKE|1|52|他叫有權柄的失位， 叫卑賤的升高。
LUKE|1|53|他叫飢餓的飽餐美食， 叫富足的空手回去。
LUKE|1|54|他扶助了他的僕人 以色列 ，不忘記施憐憫，
LUKE|1|55|正如他對我們的列祖說過， 『憐憫 亞伯拉罕 和他的後裔，直到永遠。』」
LUKE|1|56|馬利亞 和 伊利莎白 同住，約有三個月，然後回家去了。
LUKE|1|57|伊利莎白 的產期到了，生了一個兒子。
LUKE|1|58|鄰里親屬聽見主向她大施憐憫，就和她一同歡樂。
LUKE|1|59|到了第八日，他們來給孩子行割禮，並要照他父親的名字叫他 撒迦利亞 。
LUKE|1|60|他母親回應說：「不！要叫他 約翰 。」
LUKE|1|61|他們對她說：「你親族中沒有叫這名字的。」
LUKE|1|62|他們就向他父親打手勢，問他這孩子要叫甚麼名字。
LUKE|1|63|他要了一塊寫字的板，寫上：「他的名字是 約翰 。」他們就都驚訝。
LUKE|1|64|撒迦利亞 的口立刻開了，舌頭也鬆了，就開始說話稱頌上帝。
LUKE|1|65|周圍居住的人都懼怕；這一切的事就傳遍了 猶太 山區。
LUKE|1|66|凡聽見的人都把這事放在心裏，他們說：「這個孩子將來會怎麼樣呢？」因為有主的手與他同在。
LUKE|1|67|他父親 撒迦利亞 被聖靈充滿，就預言說：
LUKE|1|68|「主— 以色列 的上帝是應當稱頌的！ 因他眷顧他的百姓，為他們施行救贖，
LUKE|1|69|在他僕人 大衛 家中， 為我們興起了拯救的角，
LUKE|1|70|正如主藉著古時候聖先知的口所說的，
LUKE|1|71|『他拯救我們脫離仇敵， 脫離一切恨我們之人的手。
LUKE|1|72|他向我們列祖施憐憫， 記得他的聖約，
LUKE|1|73|就是他對我們祖宗 亞伯拉罕 所起的誓，
LUKE|1|74|叫我們既從仇敵手中被救出來， 就可以終身在他面前， 無所懼怕地用聖潔和公義事奉他。
LUKE|1|75|
LUKE|1|76|孩子啊，你要稱為至高者的先知； 因為你要走在主的前面，為他預備道路，
LUKE|1|77|叫他的百姓因罪得赦， 認識救恩；
LUKE|1|78|因我們上帝憐憫的心腸， 叫清晨的日光從高天臨到我們，
LUKE|1|79|要照亮坐在黑暗中死蔭裏的人， 把我們的腳引到和平的路上。』」
LUKE|1|80|這孩子漸漸長大，心靈堅強，住在曠野，直到他在 以色列 人面前公開出現的日子。
LUKE|2|1|在那些日子，凱撒 奧古斯都 降旨，叫全國人民都登記戶籍。
LUKE|2|2|這第一次登記戶籍是在 居里扭 作 敘利亞 總督的時候行的。
LUKE|2|3|眾人各歸各城，辦理登記。
LUKE|2|4|約瑟 也從 加利利 的 拿撒勒城 上 猶太 去，到了 大衛 的城名叫 伯利恆 ，因為他是 大衛 家族的人，
LUKE|2|5|要和他所聘之妻 馬利亞 一同登記戶籍。那時 馬利亞 已經懷孕。
LUKE|2|6|他們在那裏的時候， 馬利亞 的產期到了，
LUKE|2|7|就生了頭胎的兒子，用布包起來，放在馬槽裏，因為客店裏沒有地方。
LUKE|2|8|在 伯利恆 的野外有牧羊人，夜間值班看守羊群。
LUKE|2|9|有主的一個使者站在他們旁邊，主的榮光四面照著他們，牧羊人就很懼怕。
LUKE|2|10|那天使對他們說：「不要懼怕！看哪！因為我報給你們大喜的信息，是關乎萬民的：
LUKE|2|11|因今天在 大衛 的城裏，為你們生了救主，就是主基督。
LUKE|2|12|你們要看見一個嬰孩，包著布，臥在馬槽裏，那就是給你們的記號。」
LUKE|2|13|忽然，有一大隊天兵同那天使讚美上帝說：
LUKE|2|14|「在至高之處榮耀歸與上帝！ 在地上平安歸與他所喜悅的人！」
LUKE|2|15|眾天使離開他們，升天去了。牧羊人彼此說：「我們往 伯利恆 去，看看所成的事，就是主所告訴我們的。」
LUKE|2|16|他們急忙去了，找到 馬利亞 和 約瑟 ，還有那嬰孩臥在馬槽裏。
LUKE|2|17|他們看見，就把天使論這孩子的話傳開了。
LUKE|2|18|聽見的人都詫異牧羊人對他們所說的話。
LUKE|2|19|馬利亞 卻把這一切的事存在心裏，反覆思考。
LUKE|2|20|牧羊人回去了，因所聽見所看見的一切事，正如天使向他們所說的，就歸榮耀於上帝，讚美他。
LUKE|2|21|滿了八天，他們就給孩子行割禮，又給他起名叫耶穌；這是他還沒有在母腹裏成胎以前天使所起的名。
LUKE|2|22|按 摩西 律法滿了潔淨的日子，他們就帶著孩子上 耶路撒冷 去，要把他獻給主。
LUKE|2|23|正如主的律法上所記：「凡頭生的男子必歸主為聖」；
LUKE|2|24|又要照主的律法上所說，用一對斑鳩，或用兩隻雛鴿獻祭。
LUKE|2|25|那時，在 耶路撒冷 有一個人，名叫 西面 ；這人又公義又虔誠，素常盼望 以色列 的安慰者來到，又有聖靈在他身上。
LUKE|2|26|他得了聖靈的啟示，知道自己未死以前必看見主所立的基督。
LUKE|2|27|他受了聖靈的感動，進入聖殿，正遇見耶穌的父母抱著孩子進來，要照律法的規矩而行。
LUKE|2|28|西面 就把他抱過來，稱頌上帝說：
LUKE|2|29|「主啊，如今可以照你的話， 容你的僕人安然去世；
LUKE|2|30|因為我的眼睛已經看見你的救恩，
LUKE|2|31|就是你在萬民面前所預備的：
LUKE|2|32|是啟示外邦人的光， 是你民 以色列 的榮耀。」
LUKE|2|33|孩子的父母因論耶穌的這些話就驚訝。
LUKE|2|34|西面 給他們祝福，又對孩子的母親 馬利亞 說：「這孩子被立，是要叫 以色列 中許多人跌倒，許多人興起；又要成為毀謗的對象，
LUKE|2|35|叫許多人心裏的意念顯露出來；你自己的心也要被劍刺透。」
LUKE|2|36|又有位女先知，名叫 亞拿 ，是 亞設 支派 法內力 的女兒，年紀已經老邁，從童女出嫁，同丈夫住了七年，
LUKE|2|37|就寡居了，現在已經八十四歲 。她不離開聖殿，禁食祈求，晝夜事奉上帝。
LUKE|2|38|正當那時，她進前來感謝上帝，對一切盼望 耶路撒冷 得救贖的人講論這孩子的事。
LUKE|2|39|約瑟 和 馬利亞 照主的律法辦完了一切的事，就回 加利利 ，到自己的城 拿撒勒 去了。
LUKE|2|40|孩子漸漸長大，強健起來，充滿智慧，又有上帝的恩典在他身上。
LUKE|2|41|每年逾越節，他父母都上 耶路撒冷 去。
LUKE|2|42|當他十二歲的時候，他們按著過節的規矩上去。
LUKE|2|43|守滿了節期，他們回去，孩童耶穌仍舊在 耶路撒冷 。他的父母並不知道，
LUKE|2|44|以為他在同行的人中間，走了一天的路程才在親屬和熟悉的人中找他，
LUKE|2|45|既找不著，就回 耶路撒冷 去找他。
LUKE|2|46|過了三天，他們發現他在聖殿裏，坐在教師中間，一面聽，一面問。
LUKE|2|47|凡聽見他的人都對他的聰明和應對感到驚奇。
LUKE|2|48|他父母看見就很驚奇。他母親對他說：「我兒啊，為甚麼對我們這樣做呢？看哪，你父親和我很焦急，到處找你！」
LUKE|2|49|耶穌對他們說：「為甚麼找我呢？難道你們不知道我應當在我父的家裏嗎？ 」
LUKE|2|50|他所說的這話，他們不明白。
LUKE|2|51|他就同他們下去，回到 拿撒勒 ，並且順從他們。他母親把這一切的事都存在心裏。
LUKE|2|52|耶穌的智慧和身量 ，並上帝和人喜愛他的心，都一齊增長。
LUKE|3|1|凱撒 提庇留 在位第十五年， 本丟．彼拉多 作 猶太 總督， 希律 作 加利利 分封的王，他兄弟 腓力 作 以土利亞 和 特拉可尼 地區分封的王， 呂撒聶 作 亞比利尼 分封的王，
LUKE|3|2|亞那 和 該亞法 作大祭司。那時， 撒迦利亞 的兒子 約翰 在曠野裏，上帝的話臨到他。
LUKE|3|3|他就走遍 約旦河 一帶地方，宣講悔改的洗禮，使罪得赦。
LUKE|3|4|正如 以賽亞 先知書上所記的話： 「在曠野有聲音呼喊著： 預備主的道， 修直他的路！
LUKE|3|5|一切山窪都要填滿； 大小山岡都要削平！ 彎彎曲曲的地方要改為筆直； 高高低低的道路要改為平坦！
LUKE|3|6|凡血肉之軀的，都要看見上帝的救恩！」
LUKE|3|7|約翰 對那出來要受他洗的眾人說：「毒蛇的孽種啊，誰指示你們逃避那將要來的憤怒呢？
LUKE|3|8|你們要結出果子來，和悔改的心相稱。不要自己心裏說：『我們有 亞伯拉罕 為祖宗。』我告訴你們，上帝能從這些石頭中給 亞伯拉罕 興起子孫來。
LUKE|3|9|現在斧子已經放在樹根上，凡不結好果子的樹就砍下來，丟在火裏。」
LUKE|3|10|眾人問他：「這樣，我們該做甚麼呢？」
LUKE|3|11|約翰 回答：「有兩件衣裳的，就分給那沒有的；有食物的，也該這樣做。」
LUKE|3|12|也有稅吏來要受洗，對他說：「老師，我們該做甚麼呢？」
LUKE|3|13|約翰 對他們說：「除了規定的數目，不要多收。」
LUKE|3|14|也有士兵問他說：「我們該做甚麼呢？」 約翰 說：「不要勒索任何人，也不要敲詐人；自己有糧餉就該知足。」
LUKE|3|15|百姓期待基督的來臨；他們心裏猜測，或許 約翰 是基督。
LUKE|3|16|約翰 對眾人說：「我是用水給你們施洗，但有一位能力比我更大的要來，我就是給他解鞋帶也不配。他要用聖靈與火給你們施洗。
LUKE|3|17|他手裏拿著簸箕，要揚淨他的穀物，把麥子收在倉裏，把糠用不滅的火燒盡。」
LUKE|3|18|約翰 又用許多別的話勸百姓，向他們傳福音。
LUKE|3|19|希律 分封王，因他兄弟之妻 希羅底 的緣故，並因他所做的一切惡事，受了 約翰 的責備。
LUKE|3|20|希律 在一切事上又添了這一件，就是把 約翰 收在監裏。
LUKE|3|21|眾百姓都受了洗，耶穌也受了洗。他正禱告的時候，天開了，
LUKE|3|22|聖靈降在他身上，形狀彷彿鴿子；又有聲音從天上來，說：「你是我的愛子，我喜愛你。」
LUKE|3|23|耶穌開始傳道，年紀約有三十歲。依人看來，他是 約瑟 的兒子， 約瑟 是 希里 的兒子，
LUKE|3|24|希里 是 瑪塔 的兒子， 瑪塔 是 利未 的兒子， 利未 是 麥基 的兒子， 麥基 是 雅拿 的兒子， 雅拿 是 約瑟 的兒子，
LUKE|3|25|約瑟 是 瑪他提亞 的兒子， 瑪他提亞 是 亞摩斯 的兒子， 亞摩斯 是 拿鴻 的兒子， 拿鴻 是 以斯利 的兒子， 以斯利 是 拿該 的兒子，
LUKE|3|26|拿該 是 瑪押 的兒子， 瑪押 是 瑪他提亞 的兒子， 瑪他提亞 是 西美 的兒子， 西美 是 約瑟 的兒子， 約瑟 是 猶大 的兒子， 猶大 是 約亞拿 的兒子，
LUKE|3|27|約亞拿 是 利撒 的兒子， 利撒 是 所羅巴伯 的兒子， 所羅巴伯 是 撒拉鐵 的兒子， 撒拉鐵 是 尼利 的兒子， 尼利 是 麥基 的兒子，
LUKE|3|28|麥基 是 亞底 的兒子， 亞底 是 哥桑 的兒子， 哥桑 是 以摩當 的兒子， 以摩當 是 珥 的兒子， 珥 是 約細 的兒子，
LUKE|3|29|約細 是 以利以謝 的兒子， 以利以謝 是 約令 的兒子， 約令 是 瑪塔 的兒子， 瑪塔 是 利未 的兒子，
LUKE|3|30|利未 是 西緬 的兒子， 西緬 是 猶大 的兒子， 猶大 是 約瑟 的兒子， 約瑟 是 約南 的兒子， 約南 是 以利亞敬 的兒子，
LUKE|3|31|以利亞敬 是 米利亞 的兒子， 米利亞 是 買南 的兒子， 買南 是 瑪達他 的兒子， 瑪達他 是 拿單 的兒子， 拿單 是 大衛 的兒子，
LUKE|3|32|大衛 是 耶西 的兒子， 耶西 是 俄備得 的兒子， 俄備得 是 波阿斯 的兒子， 波阿斯 是 沙拉 的兒子， 沙拉 是 拿順 的兒子 ，
LUKE|3|33|拿順 是 亞米拿達 的兒子， 亞米拿達 是 亞民 的兒子， 亞民 是 亞尼 的兒子， 亞尼 是 希斯崙 的兒子 ， 希斯崙 是 法勒斯 的兒子， 法勒斯 是 猶大 的兒子，
LUKE|3|34|猶大 是 雅各 的兒子， 雅各 是 以撒 的兒子， 以撒 是 亞伯拉罕 的兒子， 亞伯拉罕 是 他拉 的兒子， 他拉 是 拿鶴 的兒子，
LUKE|3|35|拿鶴 是 西鹿 的兒子， 西鹿 是 拉吳 的兒子， 拉吳 是 法勒 的兒子， 法勒 是 希伯 的兒子， 希伯 是 沙拉 的兒子，
LUKE|3|36|沙拉 是 該南 的兒子， 該南 是 亞法撒 的兒子， 亞法撒 是 閃 的兒子， 閃 是 挪亞 的兒子， 挪亞 是 拉麥 的兒子，
LUKE|3|37|拉麥 是 瑪土撒拉 的兒子， 瑪土撒拉 是 以諾 的兒子， 以諾 是 雅列 的兒子， 雅列 是 瑪勒列 的兒子， 瑪勒列 是 該南 的兒子， 該南 是 以挪士 的兒子，
LUKE|3|38|以挪士 是 塞特 的兒子， 塞特 是 亞當 的兒子， 亞當 是上帝的兒子。
LUKE|4|1|耶穌滿有聖靈，從 約旦河 回來，聖靈把他引到曠野，
LUKE|4|2|四十天受魔鬼的試探。在那些日子，他沒有吃甚麼，日子滿了，他餓了。
LUKE|4|3|魔鬼對他說：「你若是上帝的兒子，叫這塊石頭變成食物吧。」
LUKE|4|4|耶穌回答：「經上記著： 『人活著，不是單靠食物。 』」
LUKE|4|5|魔鬼又領他上了高山，霎時間把天下萬國都指給他看，
LUKE|4|6|對他說：「這一切權柄和榮華我都要給你，因為這原是交給我的，我願意給誰就給誰。
LUKE|4|7|你若在我面前下拜，這一切都歸你。」
LUKE|4|8|耶穌回答他說：「經上記著： 『要拜主—你的上帝， 惟獨事奉他。』」
LUKE|4|9|魔鬼又領他到 耶路撒冷 去，叫他站在聖殿頂上，對他說：「你若是上帝的兒子，從這裏跳下去！
LUKE|4|10|因為經上記著： 『主要為你命令他的使者保護你；
LUKE|4|11|他們要用手托住你， 免得你的腳碰在石頭上。』」
LUKE|4|12|耶穌回答他說：「經上說：『不可試探主—你的上帝。』」
LUKE|4|13|魔鬼用完了各樣的試探，就離開耶穌，再等時機。
LUKE|4|14|耶穌帶著聖靈的能力回到 加利利 ，他的名聲傳遍了四方。
LUKE|4|15|他在各會堂裏教導人，眾人都稱讚他。
LUKE|4|16|耶穌來到 拿撒勒 ，就是他長大的地方。在安息日，照他素常的規矩進了會堂，站起來要念聖經。
LUKE|4|17|有人把 以賽亞 先知的書交給他，他就打開，找到一處寫著：
LUKE|4|18|「主的靈在我身上， 因為他用膏膏我， 叫我傳福音給貧窮的人； 差遣我宣告： 被擄的得釋放， 失明的得看見， 受壓迫的得自由，
LUKE|4|19|宣告上帝悅納人的禧年。」
LUKE|4|20|於是他把書捲起來，交還給管理人，就坐下。會堂裏的人都定睛看他。
LUKE|4|21|耶穌對他們說：「你們聽見的這段經文，今天已經應驗了。」
LUKE|4|22|眾人都稱讚他，並對他口中所出的恩言感到驚訝；他們說：「這不是 約瑟 的兒子嗎？」
LUKE|4|23|耶穌對他們說：「你們一定會用這俗語向我說：『醫生，你醫治自己吧！我們聽見你在 迦百農 所做的事，也該在你自己的家鄉做吧。』」
LUKE|4|24|他又說：「我實在告訴你們，沒有先知在自己家鄉被人接納的。
LUKE|4|25|我對你們說實話，在 以利亞 的時候，天閉塞了三年六個月，遍地有大饑荒，那時， 以色列 中有許多寡婦，
LUKE|4|26|以利亞 並沒有奉差往她們中任何一個人那裏去，只奉差往 西頓 的 撒勒法 一個寡婦那裏去。
LUKE|4|27|在 以利沙 先知的時候， 以色列 中有許多痲瘋病人，但除了 敘利亞 的 乃縵 ，沒有一個得潔淨的。」
LUKE|4|28|會堂裏的人聽見這些話，都怒氣填胸，
LUKE|4|29|就起來趕他出城。他們的城造在山上；他們帶他到山崖，要把他推下去。
LUKE|4|30|他卻從他們中間穿過去，走了。
LUKE|4|31|耶穌下到 迦百農 ，就是 加利利 的一座城，在安息日教導眾人。
LUKE|4|32|他們對他的教導感到很驚奇，因為他的話裏有權柄。
LUKE|4|33|在會堂裏有一個人，被污鬼的靈附著，大聲喊叫說：
LUKE|4|34|「唉！ 拿撒勒 人耶穌，你為甚麼干擾我們？你來消滅我們嗎？我知道你是誰，你是上帝的聖者。」
LUKE|4|35|耶穌斥責他說：「不要作聲，從這人身上出來吧！」鬼把那人摔倒在眾人中間，就出來了，卻沒有傷害他。
LUKE|4|36|眾人都驚訝，彼此對問：「這是甚麼道理呢？因為他用權柄能力命令污靈，污靈就出來。」
LUKE|4|37|於是耶穌的名聲傳遍了周圍各地。
LUKE|4|38|耶穌出了會堂，進了 西門 的家。 西門 的岳母在發高燒，有些人為她求耶穌。
LUKE|4|39|耶穌站在她旁邊，斥責那高燒，燒就退了。她立刻起來服事他們。
LUKE|4|40|日落的時候，凡有病人的，不論害甚麼病，都帶到耶穌那裏。耶穌給他們每一個人按手，治好他們。
LUKE|4|41|又有鬼從好些人身上出來，喊著說：「你是上帝的兒子！」耶穌斥責他們，不許他們說話，因為他們知道他是基督。
LUKE|4|42|天亮的時候，耶穌出來，走到荒野的地方。眾人去找他，到了他那裏，要留住他，不讓他離開他們。
LUKE|4|43|但耶穌對他們說：「我也必須在別的城傳上帝國的福音，因我奉差原是為此。」
LUKE|4|44|於是耶穌在 猶太 的各會堂傳道。
LUKE|5|1|耶穌站在 革尼撒勒 湖邊，眾人擁擠他，要聽上帝的道。
LUKE|5|2|他見有兩隻船靠在湖邊，打魚的人卻離開船，洗網去了。
LUKE|5|3|有一隻船是 西門 的，耶穌就上去，請他把船撐開，稍微離岸，就坐下，在船上教導眾人。
LUKE|5|4|他講完了，對 西門 說：「把船開到水深的地方下網打魚。」
LUKE|5|5|西門 說：「老師，我們整夜勞累，並沒有打著甚麼。但依從你的話，我就下網。」
LUKE|5|6|他們下了網，圈住許多魚，網險些裂開，
LUKE|5|7|就招手叫另一隻船上的同伴來幫助。他們就來，把魚裝滿了兩隻船，船甚至要沉下去。
LUKE|5|8|西門．彼得 看見，就俯伏在耶穌膝前，說：「主啊，離開我，我是個罪人。」
LUKE|5|9|他和一切跟他一起的人對打到了這一網的魚都很驚訝。
LUKE|5|10|他的夥伴 西庇太 的兒子 雅各 、 約翰 ，也是這樣。耶穌對 西門 說：「不要怕！從今以後，你要得人了。」
LUKE|5|11|他們把兩隻船靠了岸，就撇下所有的，跟從了耶穌。
LUKE|5|12|有一回，耶穌在一個城裏，有人滿身長了痲瘋，看見他，就俯伏在地，求他說：「主啊，你若肯，你能使我潔淨。」
LUKE|5|13|耶穌伸手摸他，說：「我肯，你潔淨了吧！」痲瘋病立刻離開了他。
LUKE|5|14|耶穌吩咐他：「你不可告訴任何人，只要去，把自己給祭司察看，又因為你已經潔淨，要照 摩西 所吩咐的獻上祭物，作為證據給眾人看。」
LUKE|5|15|但耶穌的名聲越發傳揚出去。有一大群人聚集來聽道，也希望耶穌醫治他們的病。
LUKE|5|16|耶穌卻退到曠野去禱告。
LUKE|5|17|有一天，耶穌教導人，有法利賽人和律法教師在旁邊坐著；他們是從 加利利 各鄉村、 猶太 和 耶路撒冷 來的。主的能力與耶穌同在，使他能治好病人。
LUKE|5|18|這時，有些人用褥子抬著一個癱子，要把他抬進去放在耶穌面前，
LUKE|5|19|卻因人多，找不出法子抬進去，就上了房頂，從瓦間把他連褥子縋到當中，在耶穌面前。
LUKE|5|20|耶穌見他們的信心，就說：「朋友，你的罪赦了。」
LUKE|5|21|文士和法利賽人就開始議論說：「這個人是誰，竟說褻瀆的話？除了上帝一位之外，誰能赦罪呢？」
LUKE|5|22|耶穌知道他們所議論的，就回答他們說：「你們心裏為甚麼議論呢？
LUKE|5|23|說『你的罪赦了』，或說『你起來行走』，哪一樣容易呢？
LUKE|5|24|但要讓你們知道，人子在地上有赦罪的權柄。」他就對癱子說：「我吩咐你，起來！拿你的褥子回家去吧。」
LUKE|5|25|那人當著眾人面前立刻起來，拿了他所躺臥的褥子回家去，歸榮耀給上帝。
LUKE|5|26|眾人都驚奇，也歸榮耀給上帝，並且滿心懼怕，說：「我們今日看見不尋常的事了！」
LUKE|5|27|這些事以後，耶穌出去，看見一個稅吏，名叫 利未 ，在稅關坐著，就對他說：「來跟從我！」
LUKE|5|28|他就撇下所有的，起來跟從耶穌。
LUKE|5|29|利未 在自己家裏為耶穌大擺宴席，有一大群稅吏和別的人與他們一同坐席。
LUKE|5|30|法利賽人和文士就向耶穌的門徒發怨言說：「你們為甚麼跟稅吏和罪人一同吃喝呢？」
LUKE|5|31|耶穌回答他們：「健康的人用不著醫生；有病的人才用得著。
LUKE|5|32|我不是來召義人悔改，而是召罪人悔改。」
LUKE|5|33|他們對耶穌說：「 約翰 的門徒常常禁食祈禱，法利賽人的門徒也是這樣，惟獨跟你在一起的又吃又喝。」
LUKE|5|34|耶穌對他們說：「新郎和賓客在一起的時候，你們怎麼能叫賓客禁食呢？
LUKE|5|35|但日子將到，新郎要被帶走，那些日子他們就要禁食了。」
LUKE|5|36|耶穌又講一個比喻，對他們說：「沒有人把新衣服撕下一塊來補在舊衣服上，若是這樣，會把新的撕裂了，並且所撕下來的那塊新的和舊的也不相稱。
LUKE|5|37|也沒有人把新酒裝在舊皮袋裏；若是這樣，新酒會脹破皮袋，酒就漏出來，皮袋也糟蹋了。
LUKE|5|38|相反地，新酒必須裝在新皮袋裏。
LUKE|5|39|沒有人喝了陳酒又想喝新的；他總說陳的好。」
LUKE|6|1|有一個安息日 ，耶穌從麥田經過。他的門徒摘了麥穗，用手搓著吃。
LUKE|6|2|有幾個法利賽人說：「你們為甚麼做安息日不合法的事呢？」
LUKE|6|3|耶穌回答他們：「 大衛 和跟從他的人飢餓時所做的事，你們沒有念過嗎？
LUKE|6|4|他怎麼進了上帝的居所，拿供餅吃，又給跟從的人吃呢？這餅惟獨祭司可以吃，別人都不可以吃。」
LUKE|6|5|他又對他們說：「人子是安息日的主。」
LUKE|6|6|又有一個安息日，耶穌進了會堂教導人，在那裏有一個人，他的右手萎縮了。
LUKE|6|7|文士和法利賽人窺探耶穌會不會在安息日治病，為要找把柄告他。
LUKE|6|8|耶穌卻知道他們的意念，就對那萎縮了手的人說：「起來，站在當中！」那人就起來，站著。
LUKE|6|9|耶穌對他們說：「我問你們，在安息日行善行惡，救命害命，哪樣是合法的呢？」
LUKE|6|10|他就環視眾人，對那人說：「伸出手來！」他照著做，他的手就復原了。
LUKE|6|11|他們怒氣填胸，彼此商議怎樣對付耶穌。
LUKE|6|12|在那些日子，耶穌出去，上山祈禱，整夜向上帝禱告。
LUKE|6|13|到了天亮，他叫門徒來，就從他們中間挑選十二個人，稱他們為使徒。
LUKE|6|14|這十二個人有 西門 （耶穌又給他起名叫 彼得 ），還有他弟弟 安得烈 ，又有 雅各 和 約翰 ， 腓力 和 巴多羅買 ，
LUKE|6|15|馬太 和 多馬 ， 亞勒腓 的兒子 雅各 和激進黨的 西門 ，
LUKE|6|16|雅各 的兒子 猶大 和後來成為出賣者的 加略 人 猶大 。
LUKE|6|17|耶穌和他們下了山，站在一塊平地上；在一起的有許多門徒，又有許多百姓從全 猶太 和 耶路撒冷 ，並 推羅 、 西頓 的海邊來，
LUKE|6|18|都要聽他講道，又希望耶穌醫治他們的病；還有被污靈纏磨的，也得了醫治。
LUKE|6|19|眾人都想要摸他，因為有能力從他身上發出來，治好了他們。
LUKE|6|20|耶穌舉目看著門徒，說： 「貧窮的人有福了！ 因為上帝的國是你們的。
LUKE|6|21|現在飢餓的人有福了！ 因為你們將得飽足。 現在哭泣的人有福了！ 因為你們將要歡笑。
LUKE|6|22|人為人子的緣故憎恨你們，拒絕你們，辱罵你們，把你們當惡人除掉你們的名，你們就有福了！
LUKE|6|23|在那日，你們要歡欣雀躍，因為你們在天上的賞賜是很多的；他們的祖宗也是這樣待先知的。
LUKE|6|24|但你們富足的人有禍了！ 因為你們已經受過安慰。
LUKE|6|25|你們現在飽足的人有禍了！ 因為你們將要飢餓。 你們現在歡笑的人有禍了！ 因為你們將要哀慟哭泣。
LUKE|6|26|人都說你們好的時候，你們有禍了！因為他們的祖宗也是這樣待假先知的。」
LUKE|6|27|「可是我告訴你們這些聽的人，要愛你們的仇敵！要善待恨你們的人！
LUKE|6|28|要祝福詛咒你們的人！要為凌辱你們的人禱告！
LUKE|6|29|有人打你的臉，連另一邊也由他打。有人拿你的外衣，連內衣也由他拿去。
LUKE|6|30|凡求你的，就給他；有人拿走你的東西，不要討回來。
LUKE|6|31|「你們想要人怎樣待你們，你們也要怎樣待人。
LUKE|6|32|你們若只愛那愛你們的人，有甚麼可感謝的呢？就是罪人也愛那愛他們的人。
LUKE|6|33|你們若善待那善待你們的人，有甚麼可感謝的呢？就是罪人也是這樣做。
LUKE|6|34|你們若借給人，希望從他收回，有甚麼可感謝的呢？就是罪人也借給罪人，再如數收回。
LUKE|6|35|你們倒要愛仇敵，要善待他們，並要借給人不指望償還，你們的賞賜就很多了，你們必作至高者的兒子，因為他恩待那忘恩的和作惡的。
LUKE|6|36|你們要仁慈，像你們的父是仁慈的。」
LUKE|6|37|「你們不要評斷別人，就不被審判；你們不要定人的罪，就不被定罪；你們要饒恕人，就必蒙饒恕。
LUKE|6|38|你們要給人，就必有給你們的，並且用十足的升斗，連搖帶按，上尖下流地倒在你們懷裏；因為你們用甚麼量器量給人，也必用甚麼量器量給你們。」
LUKE|6|39|耶穌又用比喻對他們說：「瞎子豈能領瞎子，兩個人不是都要掉在坑裏嗎？
LUKE|6|40|學生不高過老師，凡學成了的會和老師一樣。
LUKE|6|41|為甚麼看見你弟兄眼中有刺，卻不想自己眼中有梁木呢？
LUKE|6|42|你不見自己眼中有梁木，怎能對你弟兄說：『讓我去掉你眼中的刺』呢？你這假冒為善的人！先去掉自己眼中的梁木，然後才能看得清楚，好去掉你弟兄眼中的刺。」
LUKE|6|43|「沒有好樹結壞果子，也沒有壞樹結好果子。
LUKE|6|44|每一種樹木可以從其果子看出來。人不是從荊棘上摘無花果的，也不是從蒺藜裏摘葡萄的。
LUKE|6|45|善人從他心裏所存的善發出善來，惡人從他所存的惡發出惡來；因為心裏所充滿的，口裏就說出來。」
LUKE|6|46|「你們為甚麼稱呼我『主啊，主啊』，卻不照我的話做呢？
LUKE|6|47|凡到我這裏來，聽了我的話又去做的，我要告訴你們他像甚麼人：
LUKE|6|48|他像一個人蓋房子，把地挖深，將根基立在磐石上，到發大水的時候，水沖那房子，房子總不動搖，因為蓋造得好。
LUKE|6|49|但聽了不去做的，就像一個人在土地上蓋房子，沒有根基，水一沖，立刻倒塌了，並且那房子損壞得很厲害。」
LUKE|7|1|耶穌對百姓講完了這一切的話，就進了 迦百農 。
LUKE|7|2|有一個百夫長所器重的僕人害病，快要死了。
LUKE|7|3|百夫長風聞耶穌的事，就託 猶太 人的幾個長老去求耶穌來救他的僕人。
LUKE|7|4|他們到了耶穌那裏，切切地求他說：「你為他做這事是他配得的；
LUKE|7|5|因為他愛我們的民族，為我們建造會堂。」
LUKE|7|6|耶穌就和他們同去。離那家不遠，百夫長託幾個朋友去見耶穌，對他說：「主啊，不必勞駕，因你到舍下來，我不敢當。
LUKE|7|7|我也自以為不配去見你，只要你說一句話，就會讓我的僮僕得痊癒。
LUKE|7|8|因為我被派在人的權下，也有兵在我之下。我對這個說：『去！』他就去；對那個說：『來！』他就來；對我的僕人說：『做這事！』他就去做。」
LUKE|7|9|耶穌聽到這些話，就很驚訝，轉身對跟隨的眾人說：「我告訴你們，這麼大的信心，就是在 以色列 ，我也沒有見過。」
LUKE|7|10|那差來的人回到百夫長家裏，發現僕人已經好了。
LUKE|7|11|過了不久 ，耶穌往一座城去，這城名叫 拿因 ，他的門徒和一大群人與他同行。
LUKE|7|12|當他走近城門時，有一個死人被抬出來。這人是他母親獨生的兒子，而他母親又是寡婦。城裏的許多人與她一同送殯。
LUKE|7|13|主看見那寡婦就憐憫她，對她說：「不要哭。」
LUKE|7|14|於是耶穌進前來，按著槓，抬的人就站住了。耶穌說：「年輕人，我吩咐你，起來！」
LUKE|7|15|那死人就坐了起來，開始說話，耶穌就把他交給他的母親。
LUKE|7|16|眾人都驚奇，歸榮耀給上帝，說：「有大先知在我們當中興起了！」又說：「上帝眷顧了他的百姓！」
LUKE|7|17|關於耶穌的這事就傳遍了 猶太 和周圍地區。
LUKE|7|18|約翰 的門徒把這些事都告訴 約翰 。於是 約翰 叫了兩個門徒來，
LUKE|7|19|差他們到主 那裏去，說：「將要來的那位就是你嗎？還是我們要等候別人呢？」
LUKE|7|20|那兩個人來到耶穌那裏，說：「施洗的 約翰 差我們來問你：『將要來的那位就是你嗎？還是我們要等候別人呢？』」
LUKE|7|21|就在那時，耶穌治好了許多患疾病的，得瘟疫的，被邪靈附身的，又開恩使好些盲人能看見。
LUKE|7|22|耶穌回答他們：「你們去，把所看見、所聽見的告訴 約翰 ：就是盲人看見，瘸子行走，痲瘋病人得潔淨，聾子聽見，死人復活，窮人聽到福音。
LUKE|7|23|凡不因我跌倒的有福了！」
LUKE|7|24|約翰 所差來的人一走，耶穌就對眾人談到 約翰 ，說：「你們從前到曠野去，是要看甚麼呢？被吹動的蘆葦嗎？
LUKE|7|25|你們出去到底是要看甚麼？穿細軟衣服的人嗎？看哪，那穿華麗衣服、宴樂度日的人是在王宮裏。
LUKE|7|26|你們出去究竟是要看甚麼？是先知嗎？是的，我告訴你們，他比先知大多了。
LUKE|7|27|這個人就是經上所說的： 『看哪，我要差遣我的使者在你面前， 他要在你前面為你預備道路。』
LUKE|7|28|我告訴你們，凡女子所生的，沒有比 約翰 大的；但在上帝國裏，最小的比他還大。」
LUKE|7|29|眾百姓和稅吏已受過 約翰 的洗，聽見這話，就以上帝為義；
LUKE|7|30|但法利賽人和律法師沒有受過 約翰 的洗，竟廢棄了上帝為他們所定的旨意。
LUKE|7|31|主又說：「這樣，我該用甚麼來比這世代的人呢？他們好像甚麼呢？
LUKE|7|32|這正像孩童坐在街市上，彼此喊叫： 『我們為你們吹笛，你們不跳舞； 我們唱哀歌，你們不啼哭。』
LUKE|7|33|施洗的 約翰 來，不吃餅，不喝酒，你們說他是被鬼附的。
LUKE|7|34|人子來，也吃也喝，你們又說這人貪食好酒，是稅吏和罪人的朋友。
LUKE|7|35|而智慧是由所有智慧的人來證實的。」
LUKE|7|36|有一個法利賽人請耶穌和他吃飯，耶穌就到那法利賽人家裏去坐席。
LUKE|7|37|那城裏有一個女人，是個罪人，知道耶穌在法利賽人家裏坐席，就拿著盛滿香膏的玉瓶，
LUKE|7|38|站在耶穌背後，挨著他的腳哭，眼淚滴濕了耶穌的腳，就用自己的頭髮擦乾，又用嘴連連親他的腳，把香膏抹上。
LUKE|7|39|請耶穌的法利賽人看見這事，心裏說：「這人若是先知，一定知道摸他的是誰，是個怎樣的女人；她是個罪人哪！」
LUKE|7|40|耶穌回應他說：「 西門 ，我有話要對你說。」 西門 說：「老師，請說。」
LUKE|7|41|耶穌說：「有兩個人欠了某一個債主的錢，一個欠五百個銀幣，一個欠五十個銀幣。
LUKE|7|42|因為他們無力償還，債主就開恩赦免了他們兩個人的債。那麼，這兩個人哪一個更愛他呢？」
LUKE|7|43|西門 回答：「我想是那多得赦免的人。」耶穌對他說：「你的判斷不錯。」
LUKE|7|44|於是他轉過來向著那女人，對 西門 說：「你看見這女人嗎？我進了你的家，你沒有給我水洗腳，但這女人用眼淚滴濕了我的腳，又用頭髮擦乾。
LUKE|7|45|你沒有親我，但這女人從我進來就不住地親我的腳。
LUKE|7|46|你沒有用油抹我的頭，但這女人用香膏抹我的腳。
LUKE|7|47|所以我告訴你，她許多的罪都赦免了，因為她愛的多；而那少得赦免的，愛的就少。」
LUKE|7|48|於是耶穌對那女人說：「你的罪都赦免了。」
LUKE|7|49|同席的人心裏說：「這是甚麼人，竟赦免人的罪呢？」
LUKE|7|50|耶穌對那女人說：「你的信救了你，平安地回去吧！」
LUKE|8|1|過了不久，耶穌周遊各城各鄉傳道，宣講上帝國的福音。和他同去的有十二個使徒，
LUKE|8|2|還有曾被邪靈所附，被疾病所纏，而已經治好的幾個婦女，其中有稱為 抹大拉 的 馬利亞 ，曾有七個鬼從她身上趕出來，
LUKE|8|3|又有 希律 的管家 苦撒 的妻子 約亞拿 ，和 蘇撒拿 以及好些別的婦女，她們都是用自己的財物供給耶穌和使徒。
LUKE|8|4|當一大群人聚集，又有人從各城裏出來見耶穌的時候，耶穌用比喻說：
LUKE|8|5|「有一個撒種的出去撒種。他撒的時候，有的落在路旁，被人踐踏，天上的飛鳥又來把它吃掉了。
LUKE|8|6|有的落在磐石上，一出來就枯乾了，因為得不著滋潤。
LUKE|8|7|有的落在荊棘裏，荊棘跟它一同生長，把它擠住了。
LUKE|8|8|又有的落在好土裏，生長起來，結實百倍。」耶穌說完這些話，大聲說：「有耳可聽的，就應當聽！」
LUKE|8|9|門徒問耶穌這比喻是甚麼意思。
LUKE|8|10|他說：「上帝國的奧祕只讓你們知道，至於別人，就用比喻，要 他們看也看不見， 聽也不明白。」
LUKE|8|11|「這比喻是這樣的：種子就是上帝的道。
LUKE|8|12|那些在路旁的，就是人聽了道，隨後魔鬼來，從他們心裏把道奪去，以免他們信了得救。
LUKE|8|13|那些在磐石上的，就是人聽道，歡喜領受，但沒有根，不過暫時相信，等到碰上試煉就退後了。
LUKE|8|14|那落在荊棘裏的，就是人聽了道，走開以後，被今生的憂慮、錢財、宴樂擠住了，結不出成熟的子粒來。
LUKE|8|15|那落在好土裏的，就是人聽了道，並用純真善良的心持守它，耐心等候結果實。」
LUKE|8|16|「沒有人點燈用器皿蓋上，或放在床底下，而是放在燈臺上，讓進來的人看見亮光。
LUKE|8|17|因為掩藏的事沒有不顯出來的，隱瞞的事也沒有不露出來被人知道的。
LUKE|8|18|所以，你們應當小心怎樣聽。因為凡有的，還要給他；凡沒有的，連他自以為有的也要奪去。」
LUKE|8|19|耶穌的母親和他兄弟來看他，因為人多，不能到他跟前。
LUKE|8|20|有人告訴他說：「你母親和你兄弟站在外邊，要見你。」
LUKE|8|21|耶穌回答他們：「聽了上帝的道而遵行的人，就是我的母親，我的兄弟了。」
LUKE|8|22|有一天，耶穌和門徒上了船，他對門徒說：「我們渡到湖的對岸去吧。」他們就開了船。
LUKE|8|23|船行的時候，耶穌睡著了。湖上忽然起了狂風，船將灌滿了水，很危險。
LUKE|8|24|門徒去叫醒他，說：「老師！老師！我們快沒命啦！」耶穌醒了，斥責那狂風大浪，風浪就止住，平靜了。
LUKE|8|25|耶穌對他們說：「你們的信心在哪裏呢？」他們又懼怕又驚訝，彼此說：「這到底是誰？他吩咐風和水，連風和水都聽從他。」
LUKE|8|26|他們到了 格拉森 人的地區，就在 加利利 的對面。
LUKE|8|27|耶穌上了岸，就有城裏一個被鬼附的人迎著他走來。這個人好久不穿衣服，不住在屋子裏，而住在墳墓裏。
LUKE|8|28|他看見耶穌，就喊叫著俯伏在他面前，大聲說：「至高上帝的兒子耶穌，你為甚麼干擾我？我求你，不要叫我受苦！」
LUKE|8|29|這是因耶穌曾吩咐污靈從這人身上出來。原來這污靈屢次抓住他；他常被人看守，又被鐵鏈和腳鐐捆鎖，他竟把鎖鏈掙斷，被鬼趕到曠野去。
LUKE|8|30|耶穌問他：「你的名字叫甚麼？」他說：「 群 」；這是因為附著他的鬼多。
LUKE|8|31|鬼就央求耶穌不要命令他們到無底坑裏去。
LUKE|8|32|那裏有一大群豬正在山坡上吃食，鬼央求耶穌准他們進入豬裏；耶穌准了他們。
LUKE|8|33|於是鬼從那人出來，進入豬裏，那群豬就闖下山崖，投進湖裏，淹死了。
LUKE|8|34|放豬的看見這事就逃跑了，去告訴城裏和鄉下的人。
LUKE|8|35|眾人出來，要看發生了甚麼事；到了耶穌那裏，發現那人坐在耶穌腳前，鬼已離開了他，穿著衣服，神智清醒，他們就害怕。
LUKE|8|36|看見這事的人把被鬼附的人怎麼得醫治的事告訴他們。
LUKE|8|37|格拉森 周圍地區的人，因為害怕得很，都求耶穌離開他們；耶穌就上船回去了。
LUKE|8|38|鬼已從身上出去的那人懇求要和耶穌在一起，耶穌卻打發他回去，說：
LUKE|8|39|「你回家去，傳講上帝為你做了多麼大的事。」他就走遍全城，傳揚耶穌為他做了多麼大的事。
LUKE|8|40|耶穌回來的時候，眾人迎接他，因為他們都等候著他。
LUKE|8|41|有一個會堂主管，名叫 葉魯 ，來俯伏在耶穌腳前，求耶穌到他家裏去，
LUKE|8|42|因為他有一個獨生女，約十二歲，快要死了。 耶穌去的時候，眾人簇擁著他。
LUKE|8|43|有一個女人，患了經血不止的病有十二年，在醫生手裏花盡了一生所有的 ，但沒有人能治好她。
LUKE|8|44|她來到耶穌背後，摸他的衣裳繸子，經血立刻止住了。
LUKE|8|45|耶穌說：「摸我的是誰？」眾人都不承認。 彼得 說：「老師，眾人擁擁擠擠緊靠著你。」
LUKE|8|46|耶穌說：「有人摸了我，因為我覺得有能力從我身上出去。」
LUKE|8|47|那女人知道瞞不住了，就戰戰兢兢地俯伏在耶穌跟前，把摸他的緣故和怎樣立刻痊癒的事，當著眾人都說出來。
LUKE|8|48|耶穌對她說：「女兒，你的信救了你。平安地回去吧！」
LUKE|8|49|耶穌還在說話的時候，有人從會堂主管的家裏來，說：「你的女兒死了，不要勞駕老師了。」
LUKE|8|50|耶穌聽見就對他說：「不要怕，只要信！她必得痊癒。」
LUKE|8|51|耶穌到了他的家，除了 彼得 、 約翰 、 雅各 ，和女兒的父母，不許別人同他進去。
LUKE|8|52|眾人都在為這女孩哀哭捶胸。耶穌說：「不要哭，她不是死了，是睡著了。」
LUKE|8|53|他們知道她已經死了，就嘲笑耶穌。
LUKE|8|54|耶穌拉著她的手，呼叫著：「孩子，起來吧！」
LUKE|8|55|她的靈魂就回來了，她立刻起來。耶穌吩咐給她東西吃。
LUKE|8|56|她的父母非常驚奇；耶穌吩咐他們不要把所發生的事告訴任何人。
LUKE|9|1|耶穌叫齊了十二使徒，給他們能力和權柄制伏一切的鬼，醫治疾病，
LUKE|9|2|又差遣他們宣講上帝的國，醫治病人，
LUKE|9|3|對他們說：「途中甚麼都不要帶；不要帶手杖和行囊，不要帶食物和銀錢，也不要帶兩件內衣 。
LUKE|9|4|你們無論進哪一家，就住在哪裏，也從那裏離開。
LUKE|9|5|凡不接待你們的，你們離開那城的時候，要跺掉你們腳上的塵土，證明他們的不是。」
LUKE|9|6|於是使徒出去，走遍各鄉傳福音，到處治病。
LUKE|9|7|希律 分封王聽見耶穌所做的一切事，就困惑起來，因為有人說：「 約翰 從死人中復活了。」
LUKE|9|8|又有人說：「 以利亞 顯現了。」還有人說：「古時的一個先知又活了。」
LUKE|9|9|希律 說：「 約翰 我已經斬了，但這是甚麼人？關於他，我竟聽到這樣的事！」於是 希律 想要見他。
LUKE|9|10|使徒們回來，把所做的事告訴耶穌，耶穌就私下帶他們離開那裏，往一座叫 伯賽大 的城去。
LUKE|9|11|眾人知道了，就跟著他去；耶穌接待他們，對他們講論上帝國的事，治好那些需要醫治的人。
LUKE|9|12|太陽快要下山，十二使徒進前來對他說：「請叫眾人散去，他們好往四面村莊鄉鎮裏去借宿和找吃的，因為我們這裏地方偏僻。」
LUKE|9|13|耶穌對他們說：「你們給他們吃吧！」他們說：「我們不過有五個餅、兩條魚，若不去為這許多人買食物就不夠。」
LUKE|9|14|那時，男人約有五千。耶穌對門徒說：「叫他們分組坐下，每組大約五十個人。」
LUKE|9|15|門徒就這樣做了，叫眾人都坐下。
LUKE|9|16|耶穌拿著這五個餅和兩條魚，望著天祝福，擘開，遞給門徒，擺在眾人面前。
LUKE|9|17|所有的人都吃，並且吃飽了。他們把剩下的碎屑收拾起來，裝滿了十二個籃子。
LUKE|9|18|耶穌獨自禱告的時候，門徒也同他在那裏。耶穌問他們：「眾人說我是誰？」
LUKE|9|19|他們回答：「是施洗的 約翰 ；有人說是 以利亞 ；還有人說是古時的一個先知又活了。」
LUKE|9|20|耶穌問他們：「你們說我是誰？」 彼得 回答：「是上帝所立的基督。」
LUKE|9|21|耶穌切切吩咐他們，命令他們不可把這事告訴任何人；
LUKE|9|22|又說：「人子必須受許多的苦，被長老、祭司長和文士棄絕，並且被殺，第三天復活。」
LUKE|9|23|耶穌又對眾人說：「若有人要跟從我，就當捨己，天天背起自己的十字架來跟從我。
LUKE|9|24|因為凡要救自己生命的，必喪失生命；凡為我喪失生命的，他必救自己的生命。
LUKE|9|25|人就是賺得全世界，卻喪失了自己，或賠上自己，有甚麼益處呢？
LUKE|9|26|凡把我和我的道當作可恥的，人子在自己的榮耀裏，和天父與聖天使的榮耀裏來臨的時候，也要把那人當作可恥的。
LUKE|9|27|我實在告訴你們，站在這裏的，有人在沒經歷死亡以前，必定看見上帝的國。」
LUKE|9|28|說了這些話以後約有八天，耶穌帶著 彼得 、 約翰 、 雅各 上山去禱告。
LUKE|9|29|正禱告的時候，他的面貌改變了，衣服潔白放光。
LUKE|9|30|忽然有 摩西 和 以利亞 兩個人同耶穌說話；
LUKE|9|31|他們在榮光裏顯現，談論耶穌去世的事，就是他在 耶路撒冷 將要完成的事。
LUKE|9|32|彼得 和他的同伴都打盹，但一清醒，就看見耶穌的榮光和與他一起站著的那兩個人。
LUKE|9|33|二人正要和耶穌分離的時候， 彼得 對耶穌說：「老師，我們在這裏真好！我們來搭三座棚，一座為你，一座為 摩西 ，一座為 以利亞 。」他卻不知道自己在說些甚麼。
LUKE|9|34|說這些話的時候，有一朵雲彩來遮蓋他們；他們一進入雲彩就很懼怕。
LUKE|9|35|有聲音從雲彩裏出來，說：「這是我的兒子，我所揀選的 。你們要聽從他！」
LUKE|9|36|聲音停止後，只見耶穌獨自一人。當那些日子，門徒保持沉默，不把所看見的事告訴任何人。
LUKE|9|37|第二天，他們下了山，有一大群人來迎見耶穌。
LUKE|9|38|其中有一人喊著說：「老師！求你看看我的兒子，因為他是我的獨子。
LUKE|9|39|他被靈拿住就突然喊叫，那靈又使他抽風，口吐白沫，並且重重地傷害他，不輕易放過他。
LUKE|9|40|我求過你的門徒把那靈趕出去，他們卻不能。」
LUKE|9|41|耶穌回答：「唉！這又不信又悖謬的世代啊，我和你們在一起，忍耐你們，要到幾時呢？把你的兒子帶到這裏來！」
LUKE|9|42|他正來的時候，那鬼把他摔倒，使他重重地抽風。耶穌斥責那污靈，把孩子治好了，交給他父親。
LUKE|9|43|眾人都詫異上帝的大能 。 眾人正驚訝於耶穌所做的一切事的時候，耶穌對門徒說：
LUKE|9|44|「你們要把這些話聽進去，因為人子將要被交在人手裏。」
LUKE|9|45|門徒卻不明白這話，其中的意思對他們隱藏著，使他們不能明白，他們也不敢問這話的意思。
LUKE|9|46|門徒互相議論，他們中間誰最大。
LUKE|9|47|耶穌看出他們心中的議論，就領一個小孩子來，叫他站在自己旁邊，
LUKE|9|48|對他們說：「凡為我的名接納這小孩子的，就是接納我；凡接納我的，就是接納那差我來的。你們中間最小的，他就是最大的。」
LUKE|9|49|約翰 回應說：「老師，我們看見一個人奉你的名趕鬼，我們就阻止他，因為他不與我們一同跟從你。」
LUKE|9|50|耶穌對他說：「不要阻止他，因為不抵擋你們的，就是幫助你們的。」
LUKE|9|51|耶穌被接上升的日子將到，他決定面向 耶路撒冷 走去。
LUKE|9|52|他打發使者在他前頭走；他們進了 撒瑪利亞 的一個村莊，要為他作準備。
LUKE|9|53|那裏的人不接待他，因為他面向著 耶路撒冷 去。
LUKE|9|54|他的門徒 雅各 和 約翰 看見了，就說：「主啊！你要我們吩咐火從天上降下來，燒滅他們 嗎？」
LUKE|9|55|耶穌轉身責備兩個門徒。
LUKE|9|56|於是他們就往別的村莊去了。
LUKE|9|57|他們在路上走的時候，有一個人對耶穌說：「你無論往哪裏去，我都要跟從你。」
LUKE|9|58|耶穌對他說：「狐狸有洞，天空的飛鳥有窩，人子卻沒有枕頭的地方。」
LUKE|9|59|他又對另一個人說：「來跟從我！」那人說：「主啊 ，容許我先回去埋葬我的父親。」
LUKE|9|60|耶穌對他說：「讓死人埋葬他們的死人，你只管去傳講上帝的國。」
LUKE|9|61|又有一人說：「主啊，我要跟從你，但容許我先去辭別我家裏的人。」
LUKE|9|62|耶穌對他說：「手扶著犁向後看的人，不配進上帝的國。」
LUKE|10|1|這些事以後，主另外指定七十二個人 ，差遣他們兩個兩個地在他前面，往自己所要到的各城各地去。
LUKE|10|2|他對他們說：「要收的莊稼多，做工的人少。所以，你們要求莊稼的主差遣做工的人出去收他的莊稼。
LUKE|10|3|你們去吧！看！我差你們出去，如同羔羊進入狼群。
LUKE|10|4|不要帶錢囊，不要帶行囊，不要帶鞋子；在路上也不要向人問安。
LUKE|10|5|無論進哪一家，先要說：『願這一家平安。』
LUKE|10|6|那裏若有當得平安的人，你們所求的平安就必臨到那家，不然，將歸還你們。
LUKE|10|7|你們要住在那家，吃喝他們所供給的，因為工人得工錢是應當的；不要從這家搬到那家。
LUKE|10|8|無論進哪一城，人若接待你們，給你們擺上甚麼食物，你們就吃甚麼。
LUKE|10|9|要醫治那城裏的病人，對他們說：『上帝的國臨近你們了。』
LUKE|10|10|無論進哪一城，人若不接待你們，你們就到大街上去，說：
LUKE|10|11|『就是你們城裏的塵土黏在我們的腳上，我們也當著你們擦去。但是，你們該知道上帝的國臨近了。』
LUKE|10|12|我告訴你們，在那日子， 所多瑪 所受的，比那城還容易受呢！」
LUKE|10|13|「 哥拉汛 哪，你有禍了！ 伯賽大 啊，你有禍了！因為在你們中間所行的異能，若行在 推羅 、 西頓 ，他們早已披麻蒙灰，坐在地上悔改了。
LUKE|10|14|在審判的時候， 推羅 和 西頓 所受的，比你們還容易受呢！
LUKE|10|15|迦百農 啊， 你以為要被舉到天上嗎？ 你要被推下陰間！」
LUKE|10|16|耶穌又對門徒說：「聽從你們的就是聽從我；棄絕你們的就是棄絕我；棄絕我的就是棄絕差遣我來的那位。」
LUKE|10|17|那七十二個人歡歡喜喜地回來，說：「主啊，因你的名，就是鬼也服了我們。」
LUKE|10|18|耶穌對他們說：「我看見撒但從天上墜落，像閃電一樣。
LUKE|10|19|我已經給你們權柄可以踐踏蛇和蠍子，又勝過仇敵一切的能力，絕沒有甚麼能害你們。
LUKE|10|20|然而，不要因靈服了你們就歡喜，而要因你們的名記錄在天上歡喜。」
LUKE|10|21|正當那時，耶穌被聖靈感動而歡喜快樂，說：「父啊，天地的主，我感謝你！因為你把這些事向聰明智慧的人隱藏起來，而向嬰孩啟示出來。父啊，是的，因為你的美意本是如此。
LUKE|10|22|一切都是我父交給我的。除了父，沒有人知道子是誰；除了子和子所願意啟示的人，沒有人知道父是誰。」
LUKE|10|23|耶穌轉身私下對門徒說：「看見你們所看見的，那眼睛有福了。
LUKE|10|24|我告訴你們，從前有許多先知和君王要看你們所看的，卻沒有看見，要聽你們所聽的，卻沒有聽見。」
LUKE|10|25|有一個律法師起來試探耶穌，說：「老師！我該做甚麼才可以承受永生？」
LUKE|10|26|耶穌對他說：「律法上寫的是甚麼？你是怎樣念的呢？」
LUKE|10|27|他回答說：「你要盡心、盡性、盡力、盡意愛主—你的上帝，又要愛鄰 如己。」
LUKE|10|28|耶穌對他說：「你回答得正確，你這樣做就會得永生。」
LUKE|10|29|那人要證明自己有理，就對耶穌說：「誰是我的鄰舍呢？」
LUKE|10|30|耶穌回答：「有一個人從 耶路撒冷 下 耶利哥 去，落在強盜手中。他們剝去他的衣裳，把他打個半死，丟下他走了。
LUKE|10|31|偶然有一個祭司從那條路下來，看見他就從另一邊過去了。
LUKE|10|32|又有一個 利未 人來到那裏，看見他，也照樣從另一邊過去了。
LUKE|10|33|可是，有一個 撒瑪利亞 人路過那裏，看見他就動了慈心，
LUKE|10|34|上前用油和酒倒在他的傷處，包裹好了，扶他騎上自己的牲口，帶他到旅店裏去，照應他。
LUKE|10|35|第二天，他拿出兩個銀幣來，交給店主，說：『請你照應他，額外的費用，我回來時會還你。』
LUKE|10|36|你想，這三個人哪一個是落在強盜手中那人的鄰舍呢？」
LUKE|10|37|他說：「是憐憫他的。」耶穌對他說：「你去，照樣做吧！」
LUKE|10|38|他們繼續前行，耶穌進了一個村莊。有一個女人，名叫 馬大 ，接他到自己家裏。
LUKE|10|39|她有一個妹妹，名叫 馬利亞 ，在主的腳前坐著聽他的道。
LUKE|10|40|馬大 伺候的事多，心裏忙亂，進前來，說：「主啊，我的妹妹留下我一個人伺候，你不在意嗎？請吩咐她來幫助我。」
LUKE|10|41|主回答說：「 馬大 ， 馬大 ，你為許多的事操心煩惱，
LUKE|10|42|但是不可少的只有一件 。 馬利亞 已經選擇了那上好的福分，是沒有人能從她奪去的。」
LUKE|11|1|耶穌在一個地方禱告。禱告完了，有個門徒對他說：「主啊，求你教導我們禱告，像 約翰 教導他的門徒一樣。」
LUKE|11|2|耶穌對他們說：「你們禱告的時候，要說： 『父啊， 願人都尊你的名為聖； 願你的國降臨；
LUKE|11|3|我們日用的飲食，天天賜給我們。
LUKE|11|4|赦免我們的罪， 因為我們也赦免凡虧欠我們的人。 不叫我們陷入試探。 』」
LUKE|11|5|耶穌又對他們說：「你們中間誰有一個朋友半夜到他那裏去，對他說：『朋友！請借給我三個餅；
LUKE|11|6|因為我有一個朋友旅途中來到我這裏，我沒有東西招待他。』
LUKE|11|7|那人在裏面回答：『不要打擾我，門已經關了，孩子們也同我在床上了，我不能起來給你。』
LUKE|11|8|我告訴你們，雖不因他是朋友起來給他，也會因他不顧面子地直求，起來照他所需要的給他。
LUKE|11|9|我又告訴你們，祈求，就給你們；尋找，就找到；叩門，就給你們開門。
LUKE|11|10|因為凡祈求的，就得著；尋找的，就找到；叩門的，就給他開門。
LUKE|11|11|你們中間作父親的，誰有兒子 求魚，反拿蛇當魚給他呢？
LUKE|11|12|求雞蛋，反給他蠍子呢？
LUKE|11|13|你們雖然不好，尚且知道拿好東西給兒女，何況 天父，他豈不更要把聖靈賜給求他的人嗎？」
LUKE|11|14|耶穌趕出一個使人成為啞巴的鬼 ，鬼出去了，啞巴就說出話來；眾人都很驚訝。
LUKE|11|15|其中卻有人說：「他是靠著鬼王 別西卜 趕鬼。」
LUKE|11|16|又有人試探耶穌，要他顯個來自天上的神蹟。
LUKE|11|17|他知道他們的意念，就對他們說：「一國自相紛爭，必定荒蕪；一家自相紛爭，就必敗落。
LUKE|11|18|撒但若自相紛爭，他的國怎能立得住呢？因為你們說我是靠著 別西卜 趕鬼。
LUKE|11|19|我若靠著 別西卜 趕鬼，你們的子弟趕鬼又靠著誰呢？這樣，他們要作你們的判官。
LUKE|11|20|我若靠著上帝的能力趕鬼，那麼，上帝的國就已臨到你們了。
LUKE|11|21|壯士全副武裝，看守自己的住宅，他所有的都很安全；
LUKE|11|22|但有一個比他更強的來攻擊他，並且戰勝了他，就奪去他所倚靠的盔甲兵器，又分了他的掠物。
LUKE|11|23|不跟我一起的，就是反對我；不與我一起收聚的，就是在拆散。」
LUKE|11|24|「污靈離了人身，走遍無水之地尋找安歇之處，卻找不到。就說：『我要回到我原來的屋裏去。』
LUKE|11|25|他到了，看見裏面打掃乾淨，修飾好了，
LUKE|11|26|就去另帶了七個比自己更惡的靈來，都進去住在那裏。那人後來的景況比先前更壞了。」
LUKE|11|27|耶穌正說這些話的時候，眾人中間有一個女人高聲對他說：「懷你胎乳養你的有福了！」
LUKE|11|28|耶穌卻說：「更有福的是聽上帝的道而遵守的人！」
LUKE|11|29|當眾人越來越擁擠的時候，耶穌說：「這世代是一個邪惡的世代。他們求看神蹟，除了 約拿 的神蹟以外，再沒有神蹟給他們看了。
LUKE|11|30|約拿 怎樣為 尼尼微 人成了神蹟，人子也要照樣為這世代的人成為神蹟。
LUKE|11|31|在審判的時候，南方的女王要起來定這世代的人的罪，因為她從地極而來，要聽 所羅門 智慧的話。看哪，比 所羅門 更大的在這裏！
LUKE|11|32|在審判的時候， 尼尼微 人要起來定這世代的罪，因為 尼尼微 人聽了 約拿 所傳的就悔改了。看哪，比 約拿 更大的在這裏！」
LUKE|11|33|「沒有人點燈放在地窖裏，或是斗底下 ，總是放在燈臺上，讓進來的人看見亮光。
LUKE|11|34|你的眼睛就是身體的燈。當你的眼睛明亮，全身就光明，當眼睛昏花，全身就黑暗。
LUKE|11|35|所以，你要注意，免得你裏面的光暗了。
LUKE|11|36|若是你全身光明，毫無黑暗，就必全然光明，如同燈的明光照亮你。」
LUKE|11|37|耶穌正說話的時候，有一個法利賽人請他吃飯，耶穌就進去坐席。
LUKE|11|38|這法利賽人看見耶穌飯前不先洗手就很詫異。
LUKE|11|39|主對他說：「如今你們法利賽人洗淨杯盤的外面，你們裏面卻滿了貪婪和邪惡。
LUKE|11|40|無知的人哪！造外面的，不也造了裏面嗎？
LUKE|11|41|只要把杯盤裏面的施捨給人，對你們來說一切就都潔淨了。
LUKE|11|42|「但是你們法利賽人有禍了！因為你們將薄荷、芸香，和各樣蔬菜獻上十分之一，疏忽了公義和愛上帝的事；這原是你們該做的—至於其他也不可忽略。
LUKE|11|43|你們法利賽人有禍了！因為你們喜愛會堂裏的高位，又喜歡人們在街市上向你們問安。
LUKE|11|44|你們有禍了！因為你們如同不顯露的墳墓，走在上面的人並不知道。」
LUKE|11|45|律法師中有一個回答耶穌，說：「老師，你這樣說也把我們侮辱了。」
LUKE|11|46|耶穌說：「你們律法師也有禍了！因為你們把難挑的擔子放在別人身上，自己卻不肯動一個指頭去減輕這些擔子。
LUKE|11|47|你們有禍了！因為你們建造先知的墳墓，那些先知正是你們的祖宗所殺的。
LUKE|11|48|可見你們祖宗所做的事，你們是證人，你們也贊同，因為他們殺了先知，你們建造先知的墳墓。
LUKE|11|49|所以，上帝的智慧也曾說：『我要差遣先知和使徒到他們那裏去，有的他們要殘殺，有的他們要迫害』，
LUKE|11|50|為使創世以來所流眾先知的血的罪都歸在這世代的人身上，
LUKE|11|51|就是從 亞伯 的血起，直到被殺在祭壇和聖所中間的 撒迦利亞 的血為止。是的，我告訴你們，這都要向這世代的人追討。
LUKE|11|52|你們律法師有禍了！因為你們把知識的鑰匙奪了去，自己不進去，要進去的人，你們也阻擋他們。」
LUKE|11|53|耶穌從那裏出來，文士和法利賽人就開始極力地催逼他，盤問他許多事，
LUKE|11|54|伺機要抓他的話柄。
LUKE|12|1|這時，有幾萬人聚集，甚至彼此踐踏。耶穌就先對門徒說：「你們要防備法利賽人的酵，就是假冒為善。
LUKE|12|2|掩蓋的事沒有不顯露出來的，隱藏的事也沒有不被人知道的。
LUKE|12|3|因此，你們在暗中所說的，將要在明處被人聽見；在密室附耳所說的，將要在屋頂上被人宣揚。」
LUKE|12|4|「我的朋友，我對你們說，那最多只能殺人身體而不能再做甚麼的，不要怕他們。
LUKE|12|5|我提醒你們該怕的是誰：該怕那殺了以後又有權柄把人扔在地獄裏的。是的，我告訴你們，正要怕他。
LUKE|12|6|五隻麻雀不是賣二銅錢 嗎？但在上帝面前，一隻也不被忘記；
LUKE|12|7|就是你們的頭髮也都數過了。不要懼怕，你們比許多的麻雀還貴重！」
LUKE|12|8|「我又告訴你們，凡在人面前認我的，人子在上帝的使者面前也必認他；
LUKE|12|9|在人面前不認我的，人子在上帝的使者面前也必不認他。
LUKE|12|10|凡說話干犯人子的，還可得赦免；但是褻瀆聖靈的，總不得赦免。
LUKE|12|11|有人帶你們到會堂、官長和掌權的人面前，不要擔心怎麼答辯，說甚麼話；
LUKE|12|12|因為就在那時候，聖靈要指教你們該說的話。」
LUKE|12|13|人群中有一個人對耶穌說：「老師！請你吩咐我的兄弟和我分家產。」
LUKE|12|14|耶穌對他說：「你這個人！誰立我作你們的判官，或給你們分家產的呢？」
LUKE|12|15|於是他對他們說：「你們要謹慎自守，躲避一切的貪心，因為人的生命不在於家道豐富。」
LUKE|12|16|然後他用比喻對他們說：「有一個財主，田地出產豐富。
LUKE|12|17|他自己心裏想：『我的出產沒有地方儲藏，怎麼辦呢？』
LUKE|12|18|就說：『我要這麼辦：要把我的倉庫拆了，另蓋更大的，在那裏好儲藏我一切的糧食和財物，
LUKE|12|19|然後要對我自己說：你這個人哪，你有許多財物積存，可供多年享用，只管安安逸逸吃喝快樂吧！』
LUKE|12|20|上帝卻對他說：『無知的人哪！今夜就要你的性命，你所預備的要歸誰呢？』
LUKE|12|21|凡為自己積財，在上帝面前卻不富足的，也是這樣。」
LUKE|12|22|耶穌又對門徒說：「所以，我告訴你們，不要為生命憂慮吃甚麼，為身體憂慮穿甚麼。
LUKE|12|23|因為生命勝於飲食，身體勝於衣裳。
LUKE|12|24|你們想一想烏鴉：牠們既不種也不收，既沒有倉又沒有庫，上帝尚且養活牠們。你們比飛鳥要貴重得多呢！
LUKE|12|25|你們哪一個能藉著憂慮使壽數多加一刻呢 ？
LUKE|12|26|這最小的事你們尚且不能做，何必憂慮其餘的事呢？
LUKE|12|27|你們想一想百合花是怎麼長起來的：它也不勞動，也不紡線。然而我告訴你們，就是 所羅門 極榮華的時候，他所穿戴的還不如這些花的一朵呢！
LUKE|12|28|你們這小信的人哪！野地裏的草今天還在，明天就丟在爐裏，上帝還給它這樣的妝飾，何況你們呢？
LUKE|12|29|你們不要求吃甚麼，喝甚麼，也不要掛慮。
LUKE|12|30|這都是世上的外邦人所求的；你們需要這些東西，你們的父都知道。
LUKE|12|31|你們只要求他的國，這些東西就必加給你們了。
LUKE|12|32|你們這小群，不要懼怕，因為你們的父樂意把國賜給你們。
LUKE|12|33|你們要變賣財產賙濟人，為自己預備永不壞的錢囊和用不盡的財寶在天上，就是賊不能近，蟲不能蛀的地方。
LUKE|12|34|因為你們的財寶在哪裏，你們的心也在哪裏。」
LUKE|12|35|「你們要束緊腰帶，燈也要點著，
LUKE|12|36|好像僕人等候自己的主人從婚宴上回來。他來叩門，就立刻給他開門。
LUKE|12|37|主人來了，看見僕人警醒，那些僕人就有福了。我實在告訴你們，主人會叫他們坐席，自己束上腰帶，前來伺候他們。
LUKE|12|38|他或是半夜來，或是天亮之前來，看見僕人這樣，那些僕人就有福了。
LUKE|12|39|你們要知道，一家的主人若知道賊甚麼時候來，就 不容賊挖穿房屋。
LUKE|12|40|你們也要預備，因為在你們想不到的時候，人子就來了。」
LUKE|12|41|彼得 說：「主啊，這比喻是對我們說的呢？還是也對眾人呢？」
LUKE|12|42|主說：「那麼，誰是那忠心又精明的管家，主人要派他管理自己的家僕，按時定量分糧給他們的呢？
LUKE|12|43|主人來到，看見僕人這樣做，那僕人就有福了。
LUKE|12|44|我實在告訴你們，主人要派他管理所有的財產。
LUKE|12|45|如果那僕人心裏說『我的主人會來得遲』，就動手打僮僕和使女，並且吃喝醉酒，
LUKE|12|46|在想不到的日子，不知道的時候，那僕人的主人要來，重重地懲罰他 ，定他和不忠心的人同罪。
LUKE|12|47|僕人知道主人的意思，卻沒預備，又未順他的意思做，那僕人要多受責打；
LUKE|12|48|至於那不知道而做了當受責打的事的，要少受責打。多給誰，就向誰多取；多託誰，就向誰多要。」
LUKE|12|49|「我來是要把火丟在地上，假如已經燒起來，不也是我所希望的嗎？
LUKE|12|50|我有當受的洗還沒有受，在這事完成之前，我是多麼地焦急！
LUKE|12|51|你們以為我來是要使地上太平嗎？不！我告訴你們，是使人紛爭。
LUKE|12|52|從今以後，一家五個人將要紛爭，三個和兩個相爭，兩個和三個相爭：
LUKE|12|53|父親和兒子相爭， 兒子和父親相爭； 母親和女兒相爭， 女兒和母親相爭； 婆婆和媳婦相爭， 媳婦和婆婆相爭。」
LUKE|12|54|耶穌又對眾人說：「你們看見西邊起了雲彩，就說：『要下大雨了』，果然就有；
LUKE|12|55|起了南風，你們就說：『要燥熱了』，也就有了。
LUKE|12|56|假冒為善的人哪，你們知道分辨天地的氣象，怎麼不知道分辨這是甚麼時代呢？」
LUKE|12|57|「你們又為何不自己判斷甚麼是合理的呢？
LUKE|12|58|你同告你的冤家去見官，還在路上，要盡力跟他和解，免得他拉你到法官面前，法官把你交給法警，法警把你下在監裏。
LUKE|12|59|我告訴你，就是最後一小文錢 還沒有還清，你也絕不能從那裏出來。」
LUKE|13|1|正當那時，有些在場的人把 彼拉多 使 加利利 人的血攙雜在他們祭物中的事，告訴耶穌。
LUKE|13|2|耶穌對他們說：「你們以為這些 加利利 人比其他的 加利利 人更有罪，所以受這害嗎？
LUKE|13|3|我告訴你們，不是的！你們若不悔改，都同樣要滅亡！
LUKE|13|4|從前 西羅亞 樓倒塌，壓死了十八個人，你們以為那些人比一切住在 耶路撒冷 的人更有罪嗎？
LUKE|13|5|我告訴你們，不是的！你們若不悔改，都照樣要滅亡！」
LUKE|13|6|於是，耶穌用比喻說：「有一個人在葡萄園裏栽了一棵無花果樹。他前來在樹上找果子，卻找不到，
LUKE|13|7|就對園丁說：『看哪，我這三年來到這棵無花果樹前找果子，竟找不到。把它砍了吧，何必白佔土地呢？』
LUKE|13|8|園丁回答：『主啊，今年且留著，等我在樹周圍掘開土，加上肥料，
LUKE|13|9|以後若結果子便罷，不然再把它砍了。』」
LUKE|13|10|安息日，耶穌在一個會堂裏教導人。
LUKE|13|11|有一個女人被靈附身，病了十八年，腰彎得一點都直不起來。
LUKE|13|12|耶穌看見，就叫她過來，對她說：「婦人，你的病好了！」
LUKE|13|13|於是用雙手按著她，她立刻直起腰來，就歸榮耀給上帝。
LUKE|13|14|會堂的主管因為耶穌在安息日治病，就很生氣，對眾人說：「有六天應當做工，那六天之內可以來求醫，在安息日卻不可。」
LUKE|13|15|主回答他：「假冒為善的人哪，難道你們各人在安息日不解開槽上的牛和驢，牽去喝水嗎？
LUKE|13|16|何況她本是 亞伯拉罕 的後裔，被撒但捆綁了十八年，不該在安息日這天解開她的綁嗎？」
LUKE|13|17|耶穌說這些話，他的敵人都慚愧了；所有的人因他所做一切榮耀的事都很歡喜。
LUKE|13|18|耶穌說：「上帝的國像甚麼？我拿甚麼來比擬呢？
LUKE|13|19|它好比一粒芥菜種，有人拿去種在園子裏，長大成樹，天上的飛鳥在它的枝上築巢。」
LUKE|13|20|他又說：「我拿甚麼來比擬上帝的國呢？
LUKE|13|21|它好比麵酵，有婦人拿來放進三斗麵裏，直到全團都發起來。」
LUKE|13|22|耶穌往 耶路撒冷 去，在所經過的各城各鄉教導人。
LUKE|13|23|有一個人問他：「主啊，得救的人很少吧？」 耶穌對眾人說：
LUKE|13|24|「你們要努力進窄門。我告訴你們，將來有許多人想要進去，卻不能。
LUKE|13|25|等到一家之主起來關了門，你們才站在外面敲門，說：『主啊，給我們開門！』他要回答你們說：『我不認識你們，不知道你們是哪裏來的。』
LUKE|13|26|那時，你們要說：『我們在你面前吃過喝過，你也在我們的街上教導過人。』
LUKE|13|27|他要對你們說：『我 告訴你們，我不知道你們是哪裏來的。你們這一切不義的人，給我走開！』
LUKE|13|28|你們要看見 亞伯拉罕 、 以撒 、 雅各 和眾先知都在上帝的國裏，你們卻被趕到外面，在那裏要哀哭切齒了。
LUKE|13|29|從東從西，從南從北，將有人來，在上帝的國裏坐席。
LUKE|13|30|看吧，在後的，將要在前；在前的，將要在後。」
LUKE|13|31|就在那時，有幾個法利賽人來對耶穌說：「離開這裏到別處去吧，因為 希律 想要殺你。」
LUKE|13|32|耶穌對他們說：「你們去告訴那個狐狸：『你看吧，今天明天我趕鬼治病，第三天我的事就成了。』
LUKE|13|33|雖然這樣，今天明天後天我必須向前走，因為先知是不可能在 耶路撒冷 之外被害的。
LUKE|13|34|耶路撒冷 啊， 耶路撒冷 啊，你常殺害先知，又用石頭打死那奉差遣到你這裏來的人。我多少次想聚集你的兒女，好像母雞把小雞聚集在翅膀底下，可是你們不願意。
LUKE|13|35|看吧，你們的家要被廢棄。我告訴你們，你們絕不會再見到我，直到你們說：『奉主名來的是應當稱頌的！』」
LUKE|14|1|安息日，耶穌到一個法利賽人的領袖家裏去吃飯，他們就窺探他。
LUKE|14|2|這時在他面前有一個患水腫病的人。
LUKE|14|3|耶穌回答律法師和法利賽人，說：「安息日治病合不合法？」
LUKE|14|4|他們卻不說話。耶穌扶著那人，治好了他，叫他走了。
LUKE|14|5|耶穌對他們說：「你們中間誰有兒子 或有牛在安息日掉在井裏，不立刻拉他上來呢？」
LUKE|14|6|他們對這些事不能反駁。
LUKE|14|7|耶穌見所請的客人選擇首位，就用比喻對他們說：
LUKE|14|8|「你被人請去赴婚宴，不要坐在首位上，恐怕主人請了比你尊貴的客人，
LUKE|14|9|請了你和他的那人前來，對你說：『請讓座給這一位吧。』你就羞羞慚慚地退到末位去了。
LUKE|14|10|你被請的時候，去坐在末位上，好讓主人來對你說：『朋友，請上座。』那時，你在同席的人面前就有光彩了。
LUKE|14|11|因為凡自高的，必降為卑；自甘卑微的，必升為高。」
LUKE|14|12|耶穌又對請他的人說：「你準備午飯或晚餐，不要請你的朋友、弟兄、親屬和富足的鄰舍，免得他們回請你，你就得了報答。
LUKE|14|13|你擺設宴席，倒要請那貧窮的、殘疾的、瘸腿的、失明的，
LUKE|14|14|你就有福了！因為他們沒有甚麼可報答你。到義人復活的時候，你要得到報答。」
LUKE|14|15|同席的有一人聽見這些話，就對耶穌說：「在上帝國裏吃飯的有福了！」
LUKE|14|16|耶穌對他說：「有人擺設大宴席，請了許多客人。
LUKE|14|17|到了坐席的時候，他打發僕人去對所請的人說：『請來吧！樣樣都已齊備了。』
LUKE|14|18|眾人異口同聲地推辭。頭一個對他說：『我買了一塊地，必須去看看。請你准我辭了。』
LUKE|14|19|另一個說：『我買了五對牛，要去試一試。請你准我辭了。』
LUKE|14|20|又有一個說：『我才娶了妻子，所以不能去。』
LUKE|14|21|那僕人回來，把這些事都告訴了主人。這家的主人就發怒，對僕人說：『快出去，到城裏大街小巷，領那貧窮的、殘疾的、失明的、瘸腿的來。』
LUKE|14|22|僕人說：『主啊，你所吩咐的已經辦了，還有空位。』
LUKE|14|23|主人對僕人說：『你出去，到大街小巷強拉人進來，坐滿我的屋子。
LUKE|14|24|我告訴你們，先前所請的人沒有一個可以嘗到我的宴席。』」
LUKE|14|25|有一大群人和耶穌同行。他轉過來對他們說：
LUKE|14|26|「無論甚麼人到我這裏來，若不愛我勝過愛 自己的父母、妻子、兒女、兄弟、姊妹，甚至自己的性命，就不能作我的門徒。
LUKE|14|27|凡不背著自己的十字架來跟從我的，也不能作我的門徒。
LUKE|14|28|你們哪一個要蓋一座樓，不先坐下來計算費用，看能不能蓋成？
LUKE|14|29|免得安了地基，不能蓋成，看見的人都笑話他，說：
LUKE|14|30|『這個人開了工，卻不能完工。』
LUKE|14|31|或是一個王出去和別的王打仗，豈不先坐下來酌量，他能不能用一萬兵去抵抗那領二萬兵來攻打他的嗎？
LUKE|14|32|若是不能，他就趁敵人還遠的時候，派使者去談和平的條件。
LUKE|14|33|這樣，你們無論甚麼人，若不撇下一切所有的，就不能作我的門徒。」
LUKE|14|34|「鹽本是好的；鹽若失了味，怎能叫它再鹹呢？
LUKE|14|35|或用在田裏，或堆在糞裏，都不合適，只好丟在外面。有耳可聽的，就應當聽！」
LUKE|15|1|許多稅吏和罪人都挨近耶穌，要聽他講道。
LUKE|15|2|法利賽人和文士私下議論說：「這個人接納罪人，又同他們吃飯。」
LUKE|15|3|耶穌就用比喻對他們說：
LUKE|15|4|「你們中間誰有一百隻羊，失去其中的一隻，不把這九十九隻留在曠野，去找那失去的羊，直到找著呢？
LUKE|15|5|找到了，他就歡歡喜喜地把羊扛在肩上。
LUKE|15|6|他回到家裏，請朋友和鄰舍來，對他們說：『你們和我一同歡喜吧，我失去的羊已經找到了！』
LUKE|15|7|我告訴你們，一個罪人悔改，在天上也要這樣為他歡喜，比為九十九個不用悔改的義人歡喜還大呢！」
LUKE|15|8|「同樣，哪一個婦人有十塊錢 ，若失落一塊，不點上燈，打掃屋子，細細地找，直到找著呢？
LUKE|15|9|找到了，她就請朋友和鄰舍來，對她們說：『你們和我一同歡喜吧，我失落的那塊錢已經找到了！』
LUKE|15|10|我告訴你們，一個罪人悔改，上帝的使者也是這樣為他歡喜。」
LUKE|15|11|耶穌又說：「一個人有兩個兒子。
LUKE|15|12|小兒子對父親說：『父親，請你把我應得的家業分給我。』他父親就把財產分給他們。
LUKE|15|13|過了不多幾天，小兒子把他一切所有的都收拾起來，往遠方去了。在那裏，他任意放蕩，浪費錢財。
LUKE|15|14|他耗盡了一切所有的，又恰逢那地方有大饑荒，就窮困起來。
LUKE|15|15|於是他去投靠當地的一個居民，那人打發他到田裏去放豬。
LUKE|15|16|他恨不得拿豬所吃的豆莢充飢，也沒有人給他甚麼吃的。
LUKE|15|17|他醒悟過來，就說：『我父親有多少雇工，糧食有餘，我倒在這裏餓死嗎？
LUKE|15|18|我要起來，到我父親那裏去，對他說：父親！我得罪了天，又得罪了你，
LUKE|15|19|從今以後，我不配稱為你的兒子，把我當作一個雇工吧。』
LUKE|15|20|於是他起來，往他父親那裏去。相離還遠，他父親看見，就動了慈心，跑去擁抱著他，連連親他。
LUKE|15|21|兒子對他說：『父親！我得罪了天，又得罪了你，從今以後，我不配稱為你的兒子。』
LUKE|15|22|父親卻吩咐僕人：『快把那上好的袍子拿出來給他穿，把戒指戴在他指頭上，把鞋穿在他腳上，
LUKE|15|23|把那肥牛犢牽來宰了，我們來吃喝慶祝；
LUKE|15|24|因為我這個兒子是死而復活，失而復得的。』他們就開始慶祝。
LUKE|15|25|「那時，大兒子正在田裏。他回來，離家不遠時，聽見奏樂跳舞的聲音，
LUKE|15|26|就叫一個僮僕來，問是甚麼事。
LUKE|15|27|僮僕對他說：『你弟弟回來了，你父親因為他無災無病地回來，把肥牛犢宰了。』
LUKE|15|28|大兒子就生氣，不肯進去，他父親出來勸他。
LUKE|15|29|他對父親說：『你看，我服侍你這麼多年，從來沒有違背過你的命令，而你從來沒有給我一隻小山羊，叫我和朋友們一同快樂。
LUKE|15|30|但你這個兒子和娼妓吃光了你的財產，他一回來，你倒為他宰了肥牛犢。』
LUKE|15|31|父親對他說：『兒啊！你常和我同在，我所有的一切都是你的；
LUKE|15|32|可是你這個弟弟是死而復活，失而復得的，所以我們理當歡喜慶祝。』」
LUKE|16|1|耶穌又對門徒說：「某財主有一個管家，有人向主人告管家浪費他的財物。
LUKE|16|2|主人叫他來，對他說：『我聽到了，你做的是甚麼事？把你所經管的交代清楚，你不能再作我的管家了。』
LUKE|16|3|那管家心裏說：『主人辭我，不用我再作管家，我將來做甚麼呢？鋤地嘛，沒有力氣；討飯嘛，怕羞。
LUKE|16|4|我知道怎麼做，好叫人們在我不作管家之後，接我到他們家裏去。』
LUKE|16|5|於是他把欠他主人債的，一個一個地叫了來，問頭一個說：『你欠我主人多少？』
LUKE|16|6|他說：『一百簍 油。』管家對他說：『拿你的賬，快坐下，寫五十。』
LUKE|16|7|他問另一個說：『你欠多少？』他說：『一百石麥子。』管家對他說：『拿你的賬，寫八十。』
LUKE|16|8|主人就誇獎這不義的管家做事精明，因為今世之子應付自己的世代比光明之子更加精明。
LUKE|16|9|我又告訴你們，要藉著那不義的錢財結交朋友，到了錢財無用的時候，他們可以接你們到永遠的住處 去。
LUKE|16|10|人在最小的事上忠心，在大事上也忠心；在最小的事上不義，在大事上也不義。
LUKE|16|11|若是你們在不義的錢財上不忠心，誰還把那真實的錢財託付你們呢？
LUKE|16|12|如果你們在別人的東西上不忠心，誰還把你們自己的東西給你們呢？
LUKE|16|13|一個僕人不能服侍兩個主；他不是恨這個愛那個，就是重這個輕那個。你們不能又服侍上帝，又服侍 瑪門 。」
LUKE|16|14|法利賽人是貪愛錢財的；他們聽見這一切話，就嘲笑耶穌。
LUKE|16|15|耶穌對他們說：「你們是在人面前自稱為義的，你們的心，上帝卻知道；因為人以為尊貴的，是上帝看為可憎惡的。
LUKE|16|16|律法和先知到 約翰 為止，從此上帝國的福音傳開了，人人努力要進去。
LUKE|16|17|天地廢去比律法的一點一畫落空還要容易。
LUKE|16|18|凡休妻另娶的，就是犯姦淫；娶被丈夫休了的婦人的，也是犯姦淫。」
LUKE|16|19|「有一個財主穿著紫色袍和細麻布衣服，天天奢華宴樂。
LUKE|16|20|又有一個討飯的，名叫 拉撒路 ，渾身長瘡，被人放在財主門口，
LUKE|16|21|想得財主桌子上掉下來的碎食充飢，甚至還有狗來舔他的瘡。
LUKE|16|22|後來那討飯的死了，被天使帶去放在 亞伯拉罕 的懷裏。財主也死了，並且埋葬了。
LUKE|16|23|他在陰間受苦，舉目遠遠地望見 亞伯拉罕 ，又望見 拉撒路 在他懷裏，
LUKE|16|24|他就喊著說：『我祖 亞伯拉罕 哪，可憐我吧！請打發 拉撒路 來，用指頭尖蘸點水，涼涼我的舌頭，因為我在這火焰裏，極其痛苦。』
LUKE|16|25|亞伯拉罕 說：『孩子啊，你該回想你生前享過福， 拉撒路 也同樣受過苦，如今他在這裏得安慰，你卻受痛苦。
LUKE|16|26|除此之外，在你們和我們之間，有深淵隔開，以致人要從這邊過到你們那邊是不可能的；要從那邊過到這邊也是不可能的。』
LUKE|16|27|財主說：『我祖啊，既然這樣，求你打發 拉撒路 到我父家去，
LUKE|16|28|因為我還有五個兄弟，他可以警告他們，免得他們也來到這痛苦的地方。』
LUKE|16|29|亞伯拉罕 說：『他們有 摩西 和先知的話可以聽從。』
LUKE|16|30|他說：『不！我祖 亞伯拉罕 哪，假如有一個人從死人中到他們那裏去，他們一定會悔改。』
LUKE|16|31|亞伯拉罕 對他說：『如果他們不聽從 摩西 和先知的話，就是有人從死人中復活，他們也不會信服的。』」
LUKE|17|1|耶穌又對門徒說：「絆倒人的事是免不了的，但那絆倒人的有禍了！
LUKE|17|2|人若把這些小子中的一個絆倒的，還不如把磨石拴在他的頸項上，丟在海裏。
LUKE|17|3|你們要謹慎！若是你的弟兄犯罪，就勸戒他；他若懊悔，就饒恕他。
LUKE|17|4|如果他一天七次得罪你，又七次回頭，說：『我懊悔了』，你總要饒恕他。」
LUKE|17|5|使徒對主說：「請加增我們的信心。」
LUKE|17|6|主說：「你們若有信心像一粒芥菜種，就是對這棵桑樹說：『你要連根拔起，栽在海裏』，它也會聽從你們。」
LUKE|17|7|「你們當中誰有僕人耕地或是放羊，從田裏回來，就對他說『你快來坐下吃飯』呢？
LUKE|17|8|他豈不對僕人說『你給我預備晚飯，束上帶子伺候我，等我吃喝完了，你才可以吃喝』嗎？
LUKE|17|9|僕人照所吩咐的去做，主人還謝謝他嗎？
LUKE|17|10|這樣，你們做完了一切所吩咐的，要說：『我們是無用的僕人，所做的本是我們該做的。』」
LUKE|17|11|耶穌往 耶路撒冷 去，經過 撒瑪利亞 和 加利利 中間的地區。
LUKE|17|12|他進入一個村子，有十個痲瘋病人迎面而來，遠遠地站著，
LUKE|17|13|高聲說：「耶穌，老師啊，可憐我們吧！」
LUKE|17|14|耶穌看見，就對他們說：「你們去，把身體給祭司檢查。」他們正去的時候就潔淨了。
LUKE|17|15|其中有一個見自己已經好了，就回來大聲歸榮耀給上帝，
LUKE|17|16|又俯伏在耶穌腳前感謝他。這人是 撒瑪利亞 人。
LUKE|17|17|耶穌回答說：「潔淨了的不是十個人嗎？那九個在哪裏呢？
LUKE|17|18|除了這外族人，再沒有別人回來歸榮耀給上帝嗎？」
LUKE|17|19|於是他對那人說：「起來，走吧，你的信救了你！」
LUKE|17|20|法利賽人問：「上帝的國幾時來到？」耶穌回答：「上帝的國來到，不是眼睛看得見的。
LUKE|17|21|人也不能說：『看哪，在這裏！』或說：『在那裏！』因為上帝的國就在你們心裏 。」
LUKE|17|22|他又對門徒說：「那些日子將到，你們渴望能看見人子的一個日子，卻看不見。
LUKE|17|23|有人要對你們說：『看哪，在那裏！』或說：『看哪，在這裏！』你們不要出去，也不要追隨他們。
LUKE|17|24|好像閃電從天這邊一閃直照到天那邊，人子在他的日子 也要這樣。
LUKE|17|25|可是他必須先受許多苦，又被這世代所棄絕。
LUKE|17|26|挪亞 的日子怎樣，人子的日子也要怎樣。
LUKE|17|27|那時，人又吃又喝，又娶又嫁，直到 挪亞 進方舟的那日，洪水就來，把他們全都滅了。
LUKE|17|28|同樣，就像在 羅得 的日子，人又吃又喝，又買又賣，又耕種又建造，
LUKE|17|29|到 羅得 離開 所多瑪 的那日，有火與硫磺從天上降下來，把他們全都滅了。
LUKE|17|30|人子顯現的日子也要這樣。
LUKE|17|31|在那日，人在屋頂上，東西在屋裏，不要下來拿；人在田裏，也不要回家。
LUKE|17|32|你們想想 羅得 的妻子吧！
LUKE|17|33|凡想保全性命的，要喪失性命；凡喪失性命的，要保存性命。
LUKE|17|34|我告訴你們，在那一夜，兩個人在一張床上，一個被接去，一個被撇下。
LUKE|17|35|兩個女人一同推磨，一個被接去，一個被撇下。 」
LUKE|17|36|
LUKE|17|37|門徒回答他說：「主啊，在哪裏呢？」耶穌對他們說：「屍首在哪裏，鷹也會聚在哪裏。」
LUKE|18|1|耶穌對門徒講了一個比喻，為了要他們常常禱告，不可灰心。
LUKE|18|2|他說：「某城有一個官，不懼怕上帝，也不尊重人。
LUKE|18|3|那城裏有個寡婦，常到他那裏，說：『我有一個冤家，求你給我伸冤。』
LUKE|18|4|他很久不受理，後來心裏說：『我雖不懼怕上帝，也不尊重人，
LUKE|18|5|只因這寡婦煩擾我，我就給她伸冤吧，免得她常來糾纏我。』」
LUKE|18|6|主說：「你們聽這不義的官所說的話。
LUKE|18|7|上帝的選民晝夜呼籲他，他豈會延遲不給他們伸冤嗎？
LUKE|18|8|我告訴你們，他很快就要給他們伸冤。然而，人子來的時候，能在世上找到這樣的信德嗎？」
LUKE|18|9|耶穌向那些自以為義而藐視別人的人講了這比喻：
LUKE|18|10|「有兩個人上聖殿去禱告，一個是法利賽人，一個是稅吏。
LUKE|18|11|法利賽人獨自站著，自言自語地禱告說：『上帝啊，我感謝你，我不像別人勒索、不義、姦淫，也不像這個稅吏。
LUKE|18|12|我每週禁食兩次，凡我所得的都獻上十分之一。』
LUKE|18|13|那稅吏遠遠地站著，連舉目望天也不敢，只捶著胸，說：『上帝啊，開恩可憐我這個罪人！』
LUKE|18|14|我告訴你們，這人回家去比那人倒算為義了。因為凡自高的，必降為卑；自甘卑微的，必升為高。」
LUKE|18|15|有人甚至連嬰孩也帶來見耶穌，要他摸他們，門徒看見就責備那些人。
LUKE|18|16|耶穌卻叫他們來，說：「讓小孩子到我這裏來，不要阻止他們，因為在上帝國的正是這樣的人。
LUKE|18|17|我實在告訴你們，凡要接受上帝國的，若不像小孩子，絕不能進去。」
LUKE|18|18|有一個官問耶穌說：「善良的老師，我該做甚麼事才能承受永生？」
LUKE|18|19|耶穌對他說：「你為甚麼稱我是善良的？除了上帝一位之外，再沒有善良的。
LUKE|18|20|誡命你是知道的：『不可姦淫；不可殺人；不可偷盜；不可作假見證；當孝敬父母。』」
LUKE|18|21|那人說：「這一切我從小都遵守了。」
LUKE|18|22|耶穌聽見了，就對他說：「你還缺少一件：要變賣你一切所有的，分給窮人，就必有財寶在天上；你還要來跟從我。」
LUKE|18|23|他聽見這些話，就很憂愁，因為他很富有。
LUKE|18|24|耶穌見他變得很憂愁 ，就說：「有錢財的人進上帝的國是何等的難哪！
LUKE|18|25|駱駝穿過針眼比財主進上帝的國還容易呢！」
LUKE|18|26|聽見的人說：「這樣，誰能得救呢？」
LUKE|18|27|耶穌說：「在人所不能的事，在上帝都能。」
LUKE|18|28|彼得 說：「看哪，我們已經撇下自己所有的跟從你了。」
LUKE|18|29|耶穌對他們說：「我實在告訴你們，凡是為上帝的國撇下房屋，或是妻子、兄弟、父母、兒女的，
LUKE|18|30|沒有不在今世得更多倍，而在來世得永生的。」
LUKE|18|31|耶穌把十二使徒帶到一邊，對他們說：「看哪，我們上 耶路撒冷 去，先知所寫的一切事都要成就在人子身上。
LUKE|18|32|他將被交給外邦人；他們要戲弄他，凌辱他，向他吐唾沫，
LUKE|18|33|並要鞭打他，殺害他；第三天他要復活。」
LUKE|18|34|這些事門徒一點也不明白，這話的意思對他們是隱藏的；他們不知道所說的是甚麼。
LUKE|18|35|耶穌將近 耶利哥 的時候，有一個盲人坐在路旁討飯。
LUKE|18|36|他聽見許多人經過，就問是甚麼事。
LUKE|18|37|他們告訴他，是 拿撒勒 人耶穌經過。
LUKE|18|38|他就呼叫說：「 大衛 之子耶穌啊，可憐我吧！」
LUKE|18|39|在前頭走的人就責備他，不許他作聲，他卻越發喊叫：「 大衛 之子啊，可憐我吧！」
LUKE|18|40|耶穌就站住，吩咐把他領過來，他到了跟前，就問他：
LUKE|18|41|「你要我為你做甚麼？」他說：「主啊，我要能看見。」
LUKE|18|42|耶穌對他說：「你看見吧！你的信救了你。」
LUKE|18|43|那盲人立刻看得見了，就跟隨耶穌，一路歸榮耀給上帝。眾人看見這事，也都讚美上帝。
LUKE|19|1|耶穌進了 耶利哥 ，要從那裏經過。
LUKE|19|2|有一個人名叫 撒該 ，作稅吏長，是個財主。
LUKE|19|3|他要看看耶穌是怎樣的人，只因人多，他的身材又矮，所以看不見。
LUKE|19|4|於是他跑到前頭，爬上桑樹，要看耶穌，因為耶穌要從那裏經過。
LUKE|19|5|耶穌到了那裏，抬頭一看，對他說：「 撒該 ，快下來！今天我必須住在你家裏。」
LUKE|19|6|他就急忙下來，歡歡喜喜地接待耶穌。
LUKE|19|7|眾人看見，都私下議論說：「他竟然到罪人家裏去住宿。」
LUKE|19|8|撒該 站著對主說：「主啊，我把所有的一半給窮人；我若勒索了誰，就還他四倍。」
LUKE|19|9|耶穌對他說：「今天救恩到了這家，因為他也是 亞伯拉罕 的子孫。
LUKE|19|10|人子來是要尋找和拯救失喪的人。」
LUKE|19|11|眾人正聽見這些話的時候，耶穌因為將近 耶路撒冷 ，又因他們以為上帝的國快要顯現，就接著講了一個比喻，
LUKE|19|12|說：「有一個貴族往遠方去，為要取得王位，然後回來。
LUKE|19|13|他叫了自己的十個僕人來，交給他們十錠銀子，說：『你們去做生意，直到我回來。』
LUKE|19|14|他本國的百姓卻恨他，打發使者隨後去，說：『我們不願意這個人作我們的王。』
LUKE|19|15|他得了王位回來，就吩咐叫那領了銀子的僕人來，要知道他們做生意賺了多少。
LUKE|19|16|頭一個上來，說：『主啊，你的一錠銀子已經賺了十錠。』
LUKE|19|17|主人對他說：『好，我善良的僕人，你既在最小的事上忠心，你有權柄管十座城。』
LUKE|19|18|第二個來，說：『主啊，你的一錠銀子已經賺了五錠。』
LUKE|19|19|主人也對這個說：『你管五座城。』
LUKE|19|20|又有一個來說：『主啊！看哪，你的一錠銀子在這裏，我把它包在手巾裏存著。
LUKE|19|21|我向來怕你，因為你是嚴厲的人：沒有放的，也要去拿；沒有種的，也要去收。』
LUKE|19|22|主人對他說：『你這惡僕，我要憑你的話定你的罪。你既知道我是嚴厲的人，沒有放的也去拿，沒有種的也去收，
LUKE|19|23|為甚麼不把我的銀子存在銀行，等我來的時候，連本帶利都取回來呢？』
LUKE|19|24|於是他對那些站在旁邊的人說：『把他這一錠奪過來，給那有十錠的。』
LUKE|19|25|他們對他說：『主啊，他已經有十錠了。』
LUKE|19|26|主人說：『我告訴你們，凡有的，還要給他；沒有的，連他所有的也要奪過來。
LUKE|19|27|至於我那些仇敵，不要我作他們王的，把他們拉來，在我面前殺了！』」
LUKE|19|28|耶穌說完了這些話，就走在前面，上 耶路撒冷 去。
LUKE|19|29|快到 伯法其 和 伯大尼 ，在名叫 橄欖山 的地方，他打發兩個門徒，
LUKE|19|30|說：「你們往對面村子裏去，進去的時候會看見一匹驢駒拴在那裏，是從來沒有人騎過的，把牠解開，牽來。
LUKE|19|31|若有人問為甚麼解開牠，你們就這樣說：『主要用牠。』」
LUKE|19|32|被打發的人去了，所遇見的正如耶穌對他們所說的。
LUKE|19|33|他們解開驢駒的時候，主人問他們：「為甚麼解開驢駒？」
LUKE|19|34|他們說：「主要用牠。」
LUKE|19|35|他們把驢駒牽到耶穌那裏，把自己的衣服搭在上面，扶耶穌騎上。
LUKE|19|36|他前進的時候，眾人把衣服鋪在路上。
LUKE|19|37|他將近 耶路撒冷 ，正下 橄欖山 的時候，一大群門徒因所見過的一切異能，都歡呼起來，大聲讚美上帝，
LUKE|19|38|說： 「奉主名來的王 是應當稱頌的！ 在天上有和平； 在至高之處有榮光。」
LUKE|19|39|人群中有幾個法利賽人對耶穌說：「老師，責備你的門徒吧！」
LUKE|19|40|耶穌回答：「我告訴你們，若是這些人閉口不說，石頭也要呼叫起來。」
LUKE|19|41|耶穌快到 耶路撒冷 ，看見那城，就為它哀哭，
LUKE|19|42|說：「但願你在這日子知道有關你平安的事，不過這事現在是隱藏的，你的眼睛看不出來。
LUKE|19|43|因為日子將到，你的仇敵要築起土壘包圍你，四面困住你，
LUKE|19|44|並要消滅你和你裏頭的兒女，連一塊石頭也不留在另一塊石頭上，因為你不知道你蒙眷顧的時候。」
LUKE|19|45|耶穌一進聖殿就趕出在裏面做買賣的人，
LUKE|19|46|對他們說：「經上說： 『我的殿是禱告的殿， 你們倒使它成為賊窩了。』」
LUKE|19|47|耶穌天天在聖殿裏教導人。祭司長、文士和百姓的領袖都想殺他，
LUKE|19|48|但找不出方法來，因為百姓都側耳聽他。
LUKE|20|1|有一天，耶穌在聖殿裏教導百姓，宣講福音的時候，祭司長、文士和長老上前來，
LUKE|20|2|問他說：「你告訴我們，你仗著甚麼權柄做這些事？給你這權柄的是誰呢？」
LUKE|20|3|耶穌回答他們：「我也要問你們一句話，你們告訴我。
LUKE|20|4|約翰 的洗禮是從天上來的，還是從人間來的呢？」
LUKE|20|5|他們彼此商量說：「我們若說『從天上來的』，他會說『這樣，你們為甚麼不信他呢？』
LUKE|20|6|我們若說『從人間來的』，所有的百姓都會用石頭打死我們，因為他們信 約翰 是先知。」
LUKE|20|7|於是他們回答：「我們不知道是從哪裏來的。」
LUKE|20|8|耶穌對他們說：「我也不告訴你們，我仗著甚麼權柄做這些事。」
LUKE|20|9|耶穌用這個比喻對百姓說：「有人開墾了一個葡萄園，租給園戶，就出外遠行，去了許久。
LUKE|20|10|到了時候，他打發一個僕人到園戶那裏去，叫他們把園中當納的果子交給他；園戶竟打了他，叫他空手回去。
LUKE|20|11|園主又打發另一個僕人去，他們也打了他，並且侮辱他，叫他空手回去。
LUKE|20|12|園主又打發第三個僕人去，他們也打傷了他，把他推出去了。
LUKE|20|13|葡萄園主說：『我要怎麼做呢？我要打發我的愛子去，或許他們會尊敬他。』
LUKE|20|14|可是，園戶看見他，彼此說：『這是承受產業的。我們殺了他，產業就歸我們了！』
LUKE|20|15|於是他們把他扔出葡萄園外，殺了。這樣，葡萄園主要怎麼處置他們呢？
LUKE|20|16|他要來除滅那些園戶，將葡萄園轉給別人。」聽見的人說：「絕對不可！」
LUKE|20|17|耶穌看著他們，說：「那麼，經上記著： 『匠人所丟棄的石頭 已作了房角的頭塊石頭。』 這是甚麼意思呢？
LUKE|20|18|凡跌在那石頭上的，一定會跌得粉碎；那石頭掉在誰的身上，就要把誰壓得稀爛。」
LUKE|20|19|文士和祭司長看出這比喻是指著他們說的，當時就想要下手拿他，只是懼怕百姓。
LUKE|20|20|於是他們窺探耶穌，打發奸細裝作好人，要在他的話上抓把柄，好把他交給總督處置。
LUKE|20|21|奸細就問耶穌：「老師，我們知道你所講所教的都很正確，也不看人的面子，而是誠誠實實傳上帝的道。
LUKE|20|22|我們納稅給凱撒合不合法？」
LUKE|20|23|耶穌看出他們的詭詐，就對他們說：
LUKE|20|24|「拿一個銀幣來給我看。這像和這名號是誰的？」他們說：「是凱撒的。」
LUKE|20|25|耶穌對他們說：「這樣，凱撒的歸凱撒，上帝的歸上帝。」
LUKE|20|26|他們無法當著百姓在他的話上抓到把柄，又因他的對答而驚訝，就閉口不言了。
LUKE|20|27|有些撒都該人來見耶穌。他們說沒有復活這回事，於是問耶穌：
LUKE|20|28|「老師， 摩西 為我們寫下這話：『某人的哥哥若死了，有妻無子，他該娶哥哥的妻子，為哥哥生子立後。』
LUKE|20|29|那麼，有兄弟七人，第一個娶了妻，沒有孩子死了。
LUKE|20|30|第二個、
LUKE|20|31|第三個也娶過她；同樣地，七個人都娶過她，沒有留下孩子就死了。
LUKE|20|32|後來，那婦人也死了。
LUKE|20|33|那麼，在復活的時候，那婦人是哪一個的妻子呢？因為他們七個人都娶過她。」
LUKE|20|34|耶穌對他們說：「這世代的人有娶有嫁，
LUKE|20|35|惟有配得那要來的世代和從死人中復活的人不娶也不嫁。
LUKE|20|36|因為他們不能再死，和天使一樣；既然是復活的人，他們就是上帝的兒子。
LUKE|20|37|至於死人復活， 摩西 在《荊棘篇》上就指明了，他稱主是 亞伯拉罕 的上帝， 以撒 的上帝， 雅各 的上帝。
LUKE|20|38|上帝不是死人的上帝，而是活人的上帝，因為對他來說，人都是活的。」
LUKE|20|39|有幾個文士說：「老師，你說得好。」
LUKE|20|40|以後，他們不敢再問他甚麼了。
LUKE|20|41|耶穌對他們說：「人們怎麼說基督是 大衛 的後裔呢？
LUKE|20|42|《詩篇》 上 大衛 自己說： 「主對我主說： 『你坐在我的右邊，
LUKE|20|43|等我使你的仇敵作你的腳凳。』
LUKE|20|44|大衛 既稱他為主，他怎麼又是 大衛 的後裔呢？」
LUKE|20|45|眾百姓聽的時候，耶穌對他的門徒說：
LUKE|20|46|「你們要防備文士。他們好穿長袍走來走去，喜歡人們在街市上向他們問安，又喜愛會堂裏的高位，宴席上的首座。
LUKE|20|47|他們侵吞寡婦的家產，假意作很長的禱告。這些人要受更重的懲罰！」
LUKE|21|1|耶穌抬頭觀看，見財主把捐項投入聖殿銀庫，
LUKE|21|2|又見一個窮寡婦投了兩個小文錢 ，
LUKE|21|3|就說：「我實在告訴你們，這窮寡婦所投的比眾人更多。
LUKE|21|4|因為眾人都是拿有餘的捐獻，但這寡婦，雖然自己不足，卻把一生所有的都投進去了。」
LUKE|21|5|有人談論聖殿是用美石和供物裝飾的，耶穌就說：
LUKE|21|6|「你們所看見的這一切，日子將到，沒有一塊石頭會留在另一塊石頭上而不被拆毀的。」
LUKE|21|7|他們問他：「老師，甚麼時候有這些事呢？這些事將臨到的時候有甚麼預兆呢？」
LUKE|21|8|耶穌說：「你們要謹慎，不要受迷惑，因為將有好些人冒我的名來，說『我是基督』，又說『時候近了』，你們不要跟從他們！
LUKE|21|9|當你們聽見打仗和動亂的事，不要驚惶；因為這些事必須先發生，但終結不會立刻就到。」
LUKE|21|10|於是耶穌對他們說：「民要攻打民，國要攻打國，
LUKE|21|11|將有大地震，多處必有饑荒、瘟疫，又有可怕的異象和大神蹟從天上顯現。
LUKE|21|12|但這一切的事以前，有人要下手拿你們，迫害你們，把你們交給會堂，並且關在監裏，又為我名的緣故拉你們到君王和統治者面前。
LUKE|21|13|但這些事終必成為你們作見證的機會。
LUKE|21|14|所以，你們要立定心意，不要預先考慮怎樣申辯；
LUKE|21|15|因為我必賜你們口才和智慧，是你們一切敵人所敵不住、駁不倒的。
LUKE|21|16|連你們的父母、兄弟、親族、朋友也要把你們交給官府；你們中間也將有被他們害死的。
LUKE|21|17|你們要為我的名被眾人憎恨。
LUKE|21|18|然而，你們連一根頭髮也不會損失。
LUKE|21|19|你們憑著堅忍，就必保全性命。」
LUKE|21|20|「當你們看見 耶路撒冷 被兵圍困，就可知道它成為荒蕪的日子近了。
LUKE|21|21|那時，在 猶太 的，應當逃到山上；在城裏的，應當出來；在鄉下的，不要進城。
LUKE|21|22|因為這是報應的日子，要使經上所寫的都得應驗。
LUKE|21|23|在那些日子，懷孕的和奶孩子的就苦了。因為將有大災難降在這地方，也有憤怒臨到這百姓。
LUKE|21|24|他們要倒在刀下，又被擄到各國去。 耶路撒冷 要被外邦人踐踏，直到外邦人的日子滿了。」
LUKE|21|25|「日月星辰要顯出預兆，地上的邦國也有困苦，因海中波浪的響聲而惶惶不安。
LUKE|21|26|人想到那要臨到世界的事，就都嚇得魂不附體，因為天上的萬象都要震動。
LUKE|21|27|那時，他們要看見人子帶著能力和大榮耀駕雲來臨。
LUKE|21|28|一有這些事，你們就當挺身昂首，因為你們得救贖的日子近了。」
LUKE|21|29|耶穌對他們講了一個比喻說：「你們看無花果樹和各樣的樹，
LUKE|21|30|樹葉一長出來，你們看了自然就知道夏天近了。
LUKE|21|31|同樣，當你們看見這些事發生，就知道上帝的國近了。
LUKE|21|32|我實在告訴你們，這世代還沒有過去，一切都要發生。
LUKE|21|33|天地要廢去，我的話卻絕不廢去。」
LUKE|21|34|「你們要謹慎，免得被貪食、醉酒和今生的憂慮壓住你們的心，那日子就忽然臨到你們，
LUKE|21|35|如同羅網一樣，因為那日子要臨到所有居住在地面上的人。
LUKE|21|36|你們要時時警醒，常常祈求，使你們能逃避這一切要來的事，得以站立在人子面前。」
LUKE|21|37|耶穌每日在聖殿裏教導人，每夜出城到 橄欖山 住宿。
LUKE|21|38|眾百姓清早上聖殿，到耶穌那裏聽他講道。
LUKE|22|1|除酵節，又叫逾越節，近了。
LUKE|22|2|祭司長和文士在想法子怎樣殺害耶穌，因他們懼怕百姓。
LUKE|22|3|這時，撒但入了那稱為 加略 人 猶大 的心。他本是十二使徒裏的一個。
LUKE|22|4|他去跟祭司長和守殿官商量怎樣把耶穌交給他們。
LUKE|22|5|他們很高興，就約定給他銀子。
LUKE|22|6|他應允了，就找機會，要趁眾人不在跟前的時候把耶穌交給他們。
LUKE|22|7|除酵節到了，這一天必須宰逾越節的羔羊。
LUKE|22|8|耶穌打發 彼得 和 約翰 ，說：「你們去為我們預備逾越節的宴席，好讓我們吃。」
LUKE|22|9|他們問他：「你要我們在哪裏預備？」
LUKE|22|10|耶穌對他們說：「你們進了城，會有人拿著一罐水迎面而來，你們就跟著他，到他所進的房子裏去，
LUKE|22|11|對那家的主人說：『老師問：客房在哪裏？我和我的門徒要在那裏吃逾越節的宴席。』
LUKE|22|12|他會帶你們看一間擺設齊全的樓上大廳，你們就在那裏預備。」
LUKE|22|13|他們去了，所看到的正如耶穌所說的。他們就預備了逾越節的宴席。
LUKE|22|14|時候到了，耶穌坐席，使徒們也和他同坐。
LUKE|22|15|耶穌對他們說：「我非常渴望在受害以前和你們吃這逾越節的宴席。
LUKE|22|16|我告訴你們，我不再吃這宴席，直到它實現在上帝的國裏。」
LUKE|22|17|耶穌接過杯來，祝謝了，說：「你們拿這杯，大家分著喝。
LUKE|22|18|我告訴你們，從今以後，我不再喝這葡萄汁，直等上帝的國來到。」
LUKE|22|19|他又拿起餅來，祝謝了，就擘開，遞給他們，說：「這是我的身體，為你們捨的，你們要如此行，為的是記念我。」
LUKE|22|20|飯後他照樣拿起杯來，說：「這杯是用我的血所立的新約，為你們流出來的。
LUKE|22|21|但是，看哪，那出賣我的人的手跟我一同在桌子上。
LUKE|22|22|人子固然要照所預定的離去，但那出賣人子的人有禍了！」
LUKE|22|23|於是他們開始互相追問他們中間哪一個會做這事。
LUKE|22|24|門徒中間也起了爭論：他們中哪一個可算為大。
LUKE|22|25|耶穌對他們說：「外邦人有君王為主治理他們，那掌權管他們的稱為恩主。
LUKE|22|26|但你們不可這樣。你們中間最大的，倒要成為最小的；為領袖的，倒要像服事人的。
LUKE|22|27|是誰為大？是坐席的還是服事人的呢？不是坐席的大嗎？然而，我在你們中間是如同服事人的。
LUKE|22|28|「我在試煉之中，常和我同在的就是你們。
LUKE|22|29|我把國賜給你們，正如我父賜給我一樣，
LUKE|22|30|使你們在我的國裏坐在我的席上吃喝，並且坐在寶座上審判 以色列 十二個支派。」
LUKE|22|31|主又說：「 西門 ， 西門 ！撒但要得著你們，好篩你們像篩麥子一樣；
LUKE|22|32|但我已經為你祈求，使你不至於失了信心。你回頭以後，要堅固你的弟兄。」
LUKE|22|33|彼得 對他說：「主啊，我已準備好要同你坐牢，與你同死。」
LUKE|22|34|耶穌說：「 彼得 ，我告訴你，今日雞還沒有叫，你要三次說不認得我。」
LUKE|22|35|耶穌又對他們說：「我差你們出去的時候，沒有錢囊，沒有行囊，沒有鞋子，你們缺少甚麼沒有？」他們說：「沒有。」
LUKE|22|36|耶穌對他們說：「但如今，有錢囊的要帶著，有行囊的也一樣；沒有刀的要賣衣服買刀。
LUKE|22|37|我告訴你們，經上寫著說：『他被列在罪犯之中。』這話必須應驗在我身上，因為那關於我的事必然成就。」
LUKE|22|38|他們說：「主啊，請看！這裏有兩把刀。」耶穌對他們說：「夠了。」
LUKE|22|39|耶穌出來，照常往 橄欖山 去，門徒也跟隨他。
LUKE|22|40|到了那地方，他就對他們說：「你們要禱告，免得陷入試探。」
LUKE|22|41|於是他離開他們約有一塊石頭扔出去那麼遠，跪下禱告，
LUKE|22|42|說：「父啊！你若願意，求你將這杯撤去；然而，不是照我的意願，而是要成全你的旨意。」 〔
LUKE|22|43|有一位天使從天上顯現，加添他的力量。
LUKE|22|44|耶穌非常痛苦焦慮，禱告更加懇切，汗如大血點滴在地上。 〕
LUKE|22|45|禱告完了，他起來，到門徒那裏，見他們因為憂愁都睡著了，
LUKE|22|46|就對他們說：「你們為甚麼睡覺呢？起來禱告，免得陷入試探！」
LUKE|22|47|耶穌還在說話的時候，來了一群人。十二使徒之一名叫 猶大 的，走在前頭，接近耶穌，要親他。
LUKE|22|48|耶穌對他說：「 猶大 ，你用親吻來出賣人子嗎？」
LUKE|22|49|左右的人見了要發生的事，就說：「主啊，我們拿刀砍好不好？」
LUKE|22|50|其中有一個人把大祭司的僕人砍了一刀，削掉了他的右耳。
LUKE|22|51|耶穌回答說：「算了，住手吧！」就摸那人的耳朵，把他治好了。
LUKE|22|52|耶穌對那些來抓他的祭司長、守殿官和長老說：「你們帶著刀棒出來，如同對付強盜嗎？
LUKE|22|53|我天天同你們在聖殿裏，你們不下手抓我。現在卻是你們的時候，黑暗掌權了。」
LUKE|22|54|他們拿住耶穌，把他帶走，進入大祭司的住宅。 彼得 遠遠地跟著。
LUKE|22|55|他們在院子中間生了火，一同坐著， 彼得 也坐在他們當中。
LUKE|22|56|有一個使女看見 彼得 面向火光坐著，就定睛看他，說：「這個人素來也是同那人一起的。」
LUKE|22|57|彼得 卻不承認，說：「你這個女人，我不認得他！」
LUKE|22|58|過了一會兒，又有一個人看見他，說：「你也是他們一夥的。」 彼得 說：「你這個人，我不是！」
LUKE|22|59|約過了一小時，又有一個人堅持說：「他實在是同那人一起的，因為他也是 加利利 人。」
LUKE|22|60|彼得 說：「你這個人，我不知道你在說甚麼！」正說話之間，雞就叫了。
LUKE|22|61|主轉過身來看 彼得 ， 彼得 就想起主對他所說的話：「今日雞叫以前，你要三次不認我。」
LUKE|22|62|他就出去痛哭。
LUKE|22|63|看守耶穌的人戲弄他，打他，
LUKE|22|64|又蒙著他的眼，問他：「你說預言吧！打你的是誰？」
LUKE|22|65|他們還用許多別的話辱罵他。
LUKE|22|66|天一亮，民間的眾長老、祭司長和文士都聚集，把耶穌帶到他們的議會裏，
LUKE|22|67|說：「如果你是基督，就告訴我們。」耶穌對他們說：「我若告訴你們，你們也不信；
LUKE|22|68|我若問你們，你們也不回答。
LUKE|22|69|從今以後，人子要坐在權能者上帝的右邊。」
LUKE|22|70|他們都說：「那麼，你是上帝的兒子了？」耶穌對他們說：「你們說我是。」
LUKE|22|71|他們說：「我們何必再要見證呢？他親口所說的，我們都親耳聽見了。」
LUKE|23|1|眾人都起來，把耶穌解到 彼拉多 面前。
LUKE|23|2|他們開始控告他說：「我們見這人煽惑我們的國民，禁止我們納稅給凱撒，並說自己是基督，是王。」
LUKE|23|3|彼拉多 問耶穌：「你是 猶太 人的王嗎？」耶穌回答：「是你說的。」
LUKE|23|4|彼拉多 對祭司長們和眾人說：「我查不出這人有甚麼罪來。」
LUKE|23|5|但他們越發竭力地說：「他煽動百姓，在 猶太 全地傳道，從 加利利 起，直到這裏了。」
LUKE|23|6|彼拉多 一聽見，就問：「這人是 加利利 人嗎？」
LUKE|23|7|既知道耶穌屬 希律 所管， 彼拉多 就把他送到 希律 那裏去。那時 希律 正在 耶路撒冷 。
LUKE|23|8|希律 看見耶穌就非常高興；因為聽見過他的事，早就想要見他，並且指望看他行些神蹟，
LUKE|23|9|於是問他許多的話，耶穌卻一言不答。
LUKE|23|10|那些祭司長和文士都站著，竭力控告他。
LUKE|23|11|希律 和他的士兵就藐視耶穌，戲弄他，給他穿上華麗的衣服，把他送回 彼拉多 那裏去。
LUKE|23|12|從前 希律 和 彼拉多 彼此有仇，在那一天竟成了朋友。
LUKE|23|13|彼拉多 傳齊了眾祭司長、官長和百姓，
LUKE|23|14|對他們說：「你們解這人到我這裏，說他是煽惑百姓的。看哪，我也曾在你們面前審問他，並沒有查出這人犯過你們控告他的任何罪；
LUKE|23|15|就是 希律 也是如此，所以把他送回來。可見他沒有做甚麼該死的事。
LUKE|23|16|所以，我要責打他，把他釋放。」
LUKE|23|17|
LUKE|23|18|眾人卻一齊喊著說：「除掉這個人！釋放 巴拉巴 給我們！」
LUKE|23|19|這 巴拉巴 是因在城裏作亂和殺人而下在監裏的。
LUKE|23|20|彼拉多 願意釋放耶穌，就再次向他們講話。
LUKE|23|21|無奈他們喊著說：「把他釘十字架！把他釘十字架！」
LUKE|23|22|彼拉多 第三次對他們說：「為甚麼呢？這人做了甚麼惡事呢？我並沒有查出他有甚麼該死的罪來。所以，我要責打他，把他釋放。」
LUKE|23|23|他們大聲催逼 彼拉多 ，要求他把耶穌釘十字架；他們的聲音終於得勝。
LUKE|23|24|彼拉多 這才照他們的要求定案；
LUKE|23|25|又把他們所要求的那因作亂和殺人而下在監裏的人釋放了，而把耶穌交給他們，隨他們的意思處置。
LUKE|23|26|他們把耶穌帶去的時候，有一個 古利奈 人 西門 從鄉下來，他們就拿住他，把十字架擱在他身上，叫他背著跟在耶穌後面。
LUKE|23|27|有許多百姓跟隨耶穌，其中有好些婦女為他號咷痛哭。
LUKE|23|28|耶穌轉身對她們說：「 耶路撒冷 的女子，不要為我哭，要為你們自己和你們的兒女哭。
LUKE|23|29|因為日子將到，人要說：『不生育的、未曾懷孕的，和未曾哺乳孩子的有福了！』
LUKE|23|30|那時，人要向大山說： 『倒在我們身上！』 向小山說： 『遮蓋我們！』
LUKE|23|31|他們若在樹木青綠的時候做這些事，那麼在枯乾的時候將會怎麼樣呢？」
LUKE|23|32|另外有兩個犯人也被帶來和耶穌一同處死。
LUKE|23|33|到了一個地方，名叫髑髏地，他們就在那裏把耶穌釘在十字架上，又釘了兩個犯人：一個在右邊，一個在左邊。 〔
LUKE|23|34|這時，耶穌說：「父啊！赦免他們，因為他們所做的，他們不知道。」 〕士兵就抽籤分他的衣服。
LUKE|23|35|百姓站在那裏觀看。官長也嘲笑他，說：「他救了別人，他若是基督，是上帝所揀選的，救救他自己吧！」
LUKE|23|36|士兵也戲弄他，上前拿醋送給他喝，
LUKE|23|37|說：「你若是 猶太 人的王，救救你自己吧！」
LUKE|23|38|在耶穌上方有一個牌子寫著：「這是 猶太 人的王。」
LUKE|23|39|同釘的犯人中有一個譏笑他，說：「你不是基督嗎？救救你自己和我們吧！」
LUKE|23|40|另一個就應聲責備他，說：「你是一樣受刑的，還不怕上帝嗎？
LUKE|23|41|我們是應得的，因為我們是自作自受，但這個人沒有做過一件不對的事。」
LUKE|23|42|他對耶穌說：「耶穌啊，你進入你國的時候，求你記念我。」
LUKE|23|43|耶穌對他說：「我實在告訴你，今日你要同我在樂園裏了。」
LUKE|23|44|那時大約是正午，全地都黑暗了，直到下午三點鐘，
LUKE|23|45|太陽變黑了，殿的幔子從當中裂為兩半。
LUKE|23|46|耶穌大聲喊著說：「父啊，我將我的靈交在你手裏！」他說了這話，氣就斷了。
LUKE|23|47|百夫長看見所發生的事，就歸榮耀給上帝，說：「這人真是個義人！」
LUKE|23|48|聚集觀看這事的眾人，見了所發生的事，都捶著胸回去了。
LUKE|23|49|所有與耶穌熟悉的人，和從 加利利 跟著他來的婦女們，都遠遠地站著，看這些事。
LUKE|23|50|有一個人名叫 約瑟 ，是個議員，為人善良正直，
LUKE|23|51|卻沒有附從別人的所謀所為。他是 猶太 的 亞利馬太城 人，素常盼望著上帝的國。
LUKE|23|52|這人去見 彼拉多 ，請求要耶穌的身體。
LUKE|23|53|他把耶穌的身體取下來，用細麻布裹好，安放在鑿巖而成的墳墓裏；那墳墓從來沒有葬過人。
LUKE|23|54|那日是預備日，安息日快到了。
LUKE|23|55|那些從 加利利 和耶穌同來的婦女跟在後面，看見了墳墓和他的身體怎樣安放。
LUKE|23|56|她們就回去，預備了香料香膏。在安息日，她們遵照誡命安息了。
LUKE|24|1|七日的第一日，黎明的時候，那些婦女帶著所預備的香料來到墳墓那裏，
LUKE|24|2|發現石頭已經從墳墓滾開了，
LUKE|24|3|她們就進去，只是不見主耶穌的身體。
LUKE|24|4|正在為這事困惑的時候，忽然有兩個人站在旁邊，衣服放光。
LUKE|24|5|婦女們非常害怕，就俯伏在地上。那兩個人對她們說：「為甚麼在死人中找活人呢？
LUKE|24|6|他不在這裏，已經復活了。要記得他還在 加利利 的時候怎樣告訴你們的，
LUKE|24|7|他說：『人子必須被交在罪人手裏，釘在十字架上，第三天復活。』」
LUKE|24|8|她們就想起耶穌的話來。
LUKE|24|9|於是她們從墳墓那裏回去，把這一切事告訴十一個使徒和其餘的人。
LUKE|24|10|把這些事告訴使徒的有 抹大拉 的 馬利亞 、 約亞拿 ，和 雅各 的母親 馬利亞 ，還有跟她們在一起的婦女。
LUKE|24|11|她們這些話，使徒以為是胡言，就不相信。
LUKE|24|12|彼得 起來，跑到墳墓前，俯身往裏看，只見細麻布，就回去了，因所發生的事而心裏驚訝。
LUKE|24|13|同一天，門徒中有兩個人往一個村子去；這村子名叫 以馬忤斯 ，離 耶路撒冷 約有二十五里 。
LUKE|24|14|他們彼此談論所發生的這一切事。
LUKE|24|15|正交談議論的時候，耶穌親自走近他們，和他們同行，
LUKE|24|16|可是他們的眼睛模糊了，沒認出他。
LUKE|24|17|耶穌對他們說：「你們一邊走一邊談，彼此談論的是甚麼事呢？」他們就站住，臉上帶著愁容。
LUKE|24|18|兩人中有一個名叫 革流巴 的回答：「你是在 耶路撒冷 的旅客中，惟一還不知道這幾天在那裏發生了甚麼事的人嗎？」
LUKE|24|19|耶穌對他們說：「甚麼事呢？」他們對他說：「就是 拿撒勒 人耶穌的事。他是個先知，在上帝和眾百姓面前，說話行事都大有能力。
LUKE|24|20|祭司長們和我們的官長竟把他解去，定了死罪，釘在十字架上。
LUKE|24|21|但我們素來所盼望要救贖 以色列 民的就是他。不但如此，這些事發生到現在已經三天了。
LUKE|24|22|還有，我們中間的幾個婦女使我們驚奇：她們清早去了墳墓，
LUKE|24|23|不見他的身體，就回來告訴我們，說她們看見了天使顯現，說他活了。
LUKE|24|24|又有我們的幾個人往墳墓那裏去，所發現的正如婦女們所說的，只是沒有看見他。」
LUKE|24|25|耶穌對他們說：「無知的人哪，先知所說的一切話，你們的心信得太遲鈍了。
LUKE|24|26|基督不是必須受這些苦難，然後進入他的榮耀嗎？」
LUKE|24|27|於是，他從 摩西 和眾先知起，凡經上所指著自己的話都給他們作了解釋。
LUKE|24|28|他們走近所要去的村子，耶穌好像還要往前走，
LUKE|24|29|他們卻強留他說：「時候晚了，天快黑了，請你同我們住下吧。」耶穌就進去，要同他們住下。
LUKE|24|30|坐下來和他們用餐的時候，耶穌拿起餅來，祝福了，擘開，遞給他們。
LUKE|24|31|他們的眼睛開了，這才認出他來。耶穌卻從他們眼前消失了。
LUKE|24|32|他們彼此說：「在路上他和我們說話，給我們講解聖經的時候，我們的心在我們裏面 豈不是火熱的嗎？」
LUKE|24|33|於是他們立刻起身，回 耶路撒冷 去，看見十一個使徒和與他們正在一起的人聚集在一處，
LUKE|24|34|說：「主果然復活了，已經顯現給 西門 看了。」
LUKE|24|35|於是，兩個人把路上所遇到，和耶穌擘餅的時候怎麼被他們認出來的事，都述說了一遍。
LUKE|24|36|正說這些話的時候，耶穌親自站在他們當中，說：「願你們平安！」
LUKE|24|37|他們卻驚慌害怕，以為所看見的是魂。
LUKE|24|38|耶穌對他們說：「你們為甚麼驚恐不安？為甚麼心裏起疑惑呢？
LUKE|24|39|你們看我的手和我的腳，就知道實在是我了。摸摸我，看，因為魂無骨無肉，你們看，我是有的。」
LUKE|24|40|說了這話，他就把手和腳給他們看。
LUKE|24|41|他們還在又驚又喜、不敢相信的時候，耶穌對他們說：「你們這裏有甚麼吃的沒有？」
LUKE|24|42|他們給了他一片烤魚，
LUKE|24|43|他接過來，在他們面前吃了。
LUKE|24|44|耶穌對他們說：「這就是我從前和你們同在時所告訴你們的話： 摩西 的律法、先知的書，和《 詩篇》 上所記一切指著我的話都必須應驗。」
LUKE|24|45|於是耶穌開他們的心竅，使他們能明白聖經，
LUKE|24|46|又對他們說：「照經上所寫的，基督必受害，第三天從死人中復活，
LUKE|24|47|並且人們要奉他的名傳悔改、使罪得赦的道，從 耶路撒冷 起直傳到萬邦。
LUKE|24|48|你們就是這些事的見證。
LUKE|24|49|我要將我父所應許的降在你們身上，你們要在城裏等候，直到你們領受從上面來的能力。」
LUKE|24|50|耶穌領他們出來，直到 伯大尼 附近，就舉手給他們祝福。
LUKE|24|51|正祝福的時候，他離開他們，被帶到天上去了。
LUKE|24|52|他們就拜他，帶著極大的喜樂回 耶路撒冷 去，
LUKE|24|53|常在聖殿裏稱頌上帝。
JOHN|1|1|太初有道，道與上帝同在，道就是上帝。
JOHN|1|2|這道太初與上帝同在。
JOHN|1|3|萬物都是藉著他造的，沒有一樣不是藉著他造的。凡被造的，
JOHN|1|4|在他裏面有生命 ，這生命就是人的光。
JOHN|1|5|光照在黑暗裏，黑暗卻沒有勝過光 。
JOHN|1|6|有一個人，是從上帝那裏差來的，名叫 約翰 。
JOHN|1|7|這人來是為了作見證，是為那光作見證，要使眾人藉著他而信。
JOHN|1|8|他不是那光，而是要為那光作見證。
JOHN|1|9|那光是真光，來到世上，照亮所有的人 。
JOHN|1|10|他在世界，世界是藉著他造的，世界卻不認識他。
JOHN|1|11|他來到自己的地方，自己的人並不接納他。
JOHN|1|12|凡接納他的，就是信他名的人，他就賜他們權柄作上帝的兒女。
JOHN|1|13|這些人不是從血生的，不是從情慾生的，也不是從人的意願生的，而是從上帝生的。
JOHN|1|14|道成了肉身，住在我們中間，充充滿滿地有恩典有真理，我們也見過他的榮光，正是父獨一兒子 的榮光。
JOHN|1|15|約翰 為他作見證，喊著說：「這就是我曾說：『那在我以後來的先於我，因為在我以前，他已經存在。』」
JOHN|1|16|從他的豐富裏，我們都領受了恩典，而且恩上加恩。
JOHN|1|17|律法是藉著 摩西 頒佈的；恩典和真理卻是由耶穌基督來的。
JOHN|1|18|從來沒有人見過上帝，只有在父懷裏獨一的兒子將他表明出來。
JOHN|1|19|這是 約翰 的見證： 猶太 人從 耶路撒冷 差祭司和 利未 人到 約翰 那裏去問他：「你是誰？」
JOHN|1|20|他就承認，並不隱瞞，承認說：「我不是基督。」
JOHN|1|21|他們又問他：「那麼，你是誰？是 以利亞 嗎？」他說：「我不是。」「是那位先知嗎？」他回答：「不是。」
JOHN|1|22|於是他們對他說：「你到底是誰，好讓我們回覆差我們來的人。你說，你自己是誰？」
JOHN|1|23|他說： 「我就是那在曠野呼喊的聲音： 修直主的道。」 正如 以賽亞 先知所說的。
JOHN|1|24|那些人是法利賽人差來的。
JOHN|1|25|他們就問他：「你既不是基督，不是 以利亞 ，也不是那位先知，那麼，你為甚麼施洗呢？」
JOHN|1|26|約翰 回答：「我是用水施洗，但有一位站在你們中間，是你們不認識的，
JOHN|1|27|就是那在我以後來的，我給他解鞋帶也不配。」
JOHN|1|28|這些事發生在 約旦河 東邊的 伯大尼 ， 約翰 施洗的地方。
JOHN|1|29|第二天， 約翰 看見耶穌來到他那裏，就說：「看哪，上帝的羔羊，除去世人的罪的！
JOHN|1|30|這就是我曾說『那在我以後來的先於我，因為在我以前，他已經存在』的那一位。
JOHN|1|31|我先前不認識他，如今我來用水施洗，為要使他顯明給 以色列 人。」
JOHN|1|32|約翰 又作見證說：「我曾看見聖靈彷彿鴿子從天降下，停留在他的身上。
JOHN|1|33|我先前不認識他，可是那差我來用水施洗的對我說：『你看見聖靈降下來，停留在誰的身上，誰就是用聖靈施洗的。』
JOHN|1|34|我看見了，所以作證：這一位是上帝的兒子。」
JOHN|1|35|又過了一天， 約翰 同兩個門徒站在那裏。
JOHN|1|36|他見耶穌走過，就說：「看哪，上帝的羔羊！」
JOHN|1|37|兩個門徒聽見他的話，就跟從了耶穌。
JOHN|1|38|耶穌轉過身來，看見他們跟著，就對他們說：「你們要甚麼？」他們對他說：「拉比，你在哪裏住？」（「拉比」翻出來就是老師。）
JOHN|1|39|耶穌說：「你們來看。」他們就去看他在哪裏住。這一天他們就跟他同住；那時大約是下午四點鐘。
JOHN|1|40|聽了 約翰 的話而跟從耶穌的那兩個人，其中一個是 西門．彼得 的弟弟 安得烈 。
JOHN|1|41|他先找到自己的哥哥 西門 ，對他說：「我們遇見彌賽亞了。」（「彌賽亞」翻出來就是基督。）
JOHN|1|42|於是 安得烈 領 西門 去見耶穌。耶穌看著他，說：「你是 約翰 的兒子 西門 ，你要稱為 磯法 。」（「磯法」翻出來就是 彼得 。）
JOHN|1|43|又過了一天，耶穌想要往 加利利 去。他找到 腓力 ，就對他說：「來跟從我！」
JOHN|1|44|這 腓力 是 伯賽大 人，是 安得烈 和 彼得 的同鄉。
JOHN|1|45|腓力 找到 拿但業 ，對他說：「 摩西 在律法書上所寫的，和眾先知所記的那一位，我們遇見了，就是 約瑟 的兒子 拿撒勒 人耶穌。」
JOHN|1|46|拿但業 對他說：「 拿撒勒 還能出甚麼好的嗎？」 腓力 說：「你來看。」
JOHN|1|47|耶穌看見 拿但業 向他走來，就論到他說：「看哪，這真是個 以色列 人！他心裏是沒有詭詐的。」
JOHN|1|48|拿但業 對耶穌說：「你從哪裏認識我的？」耶穌回答他說：「 腓力 還沒有呼喚你，你在無花果樹底下，我就看見你了。」
JOHN|1|49|拿但業 回答他說：「拉比！你是上帝的兒子，你是 以色列 的王。」
JOHN|1|50|耶穌回答他說：「因為我說在無花果樹底下看見你，你就信嗎？你將看見比這些更大的事呢！」
JOHN|1|51|他又說：「我實實在在地告訴你們，你們將要看見天開了，上帝的使者在人子身上，上去下來。」
JOHN|2|1|第三日，在 加利利 的 迦拿 有一個婚宴，耶穌的母親在那裏。
JOHN|2|2|耶穌和他的門徒也被請去赴宴。
JOHN|2|3|酒用完了，耶穌的母親對他說：「他們沒有酒了。」
JOHN|2|4|耶穌說：「母親 ，我與你何干呢？我的時候還沒有到。」
JOHN|2|5|他母親對用人說：「他告訴你們甚麼，你們就做吧。」
JOHN|2|6|照 猶太 人潔淨禮的規矩，有六口石缸擺在那裏，每口可以盛兩三桶 水。
JOHN|2|7|耶穌對用人說：「把缸倒滿水。」他們就倒滿了，直到缸口。
JOHN|2|8|耶穌又說：「現在舀出來，送給宴會總管。」他們就送了去。
JOHN|2|9|宴會總管嘗了那水變的酒，並不知道是哪裏來的，只有舀水的用人知道。於是宴會總管叫新郎來，
JOHN|2|10|對他說：「人家都是先擺上好酒，等客人喝夠了才擺上次的，你倒把好酒留到現在！」
JOHN|2|11|這是耶穌所行的第一個神蹟，是在 加利利 的 迦拿 行的，顯出了他的榮耀來，他的門徒就信他了。
JOHN|2|12|這事以後，耶穌與他的母親、兄弟 和門徒 都下 迦百農 去，在那裏住了不多幾天。
JOHN|2|13|猶太 人的逾越節近了，耶穌上 耶路撒冷 去。
JOHN|2|14|他看見聖殿裏有賣牛羊和鴿子的，還有兌換銀錢的人坐著，
JOHN|2|15|耶穌就拿繩子做成鞭子，把所有的，包括牛羊都趕出聖殿，倒出兌換銀錢之人的銀錢，推翻他們的桌子，
JOHN|2|16|又對賣鴿子的說：「把這些東西拿走！不要把我父的殿當作買賣的地方。」
JOHN|2|17|他的門徒就想起經上記著：「我為你的殿心裏焦急，如同火燒。」
JOHN|2|18|因此 猶太 領袖問他：「你能顯甚麼神蹟給我們看，表明你可以做這些事呢？」
JOHN|2|19|耶穌回答他們說：「你們拆毀這殿，我三日內要把它重建。」
JOHN|2|20|猶太 人問：「這殿造了四十六年，你三日內就能重建嗎？」
JOHN|2|21|但耶穌所說的殿是指他的身體。
JOHN|2|22|所以他從死人中復活以後，門徒想起他曾說過這事，就信了聖經和耶穌所說的話。
JOHN|2|23|耶穌在 耶路撒冷 過逾越節的時候，有許多人看見他所行的神蹟，就信了他的名。
JOHN|2|24|耶穌自己卻不信任他們，因為他認識所有的人，
JOHN|2|25|也用不著誰來證明人是怎樣的，因為他自己認識人的內心。
JOHN|3|1|有一個法利賽人，名叫 尼哥德慕 ，是 猶太 人的官。
JOHN|3|2|這人夜裏來見耶穌，對他說：「拉比，我們知道你是由上帝那裏來作老師的；因為你所行的神蹟，若沒有上帝同在，無人能行。」
JOHN|3|3|耶穌回答他說：「我實實在在地告訴你，人若不重生 ，就不能見上帝的國。」
JOHN|3|4|尼哥德慕 對他說：「人已經老了，如何能重生呢？豈能再進母腹生出來嗎？」
JOHN|3|5|耶穌回答：「我實實在在地告訴你，人若不是從水和聖靈生的，就不能進上帝的國。
JOHN|3|6|從肉身生的就是肉身；從靈生的就是靈。
JOHN|3|7|我說『你們必須重生』，你不要驚訝。
JOHN|3|8|風 隨著意思吹，你聽見風的聲音，卻不知道是從哪裏來，往哪裏去；凡從聖靈生的也是如此。」
JOHN|3|9|尼哥德慕 問他：「怎麼能有這些事呢？」
JOHN|3|10|耶穌回答，對他說：「你是 以色列 人的老師，還不明白這些事嗎？
JOHN|3|11|我實實在在地告訴你，我們所說的是我們知道的，我們所見證的是我們見過的，你們卻不領受我們的見證。
JOHN|3|12|我對你們說地上的事，你們尚且不信，若對你們說天上的事，如何能信呢？
JOHN|3|13|除了從天降下 的人子，沒有人升過天。
JOHN|3|14|摩西 在曠野怎樣舉蛇，人子也必須照樣被舉起來，
JOHN|3|15|要使一切信他的人都得永生。
JOHN|3|16|「上帝愛世人，甚至將他獨一的兒子 賜給他們，叫一切信他的人不致滅亡，反得永生。
JOHN|3|17|因為上帝差他的兒子到世上來，不是要定世人的罪 ，而是要使世人因他得救。
JOHN|3|18|信他的人不被定罪；不信的人已經被定罪了，因為他不信上帝獨一兒子的名。
JOHN|3|19|光來到世上，世人因自己的行為是惡的，不愛光，倒愛黑暗，這就定了他們的罪。
JOHN|3|20|凡作惡的人都恨惡光，不來接近光，恐怕他的行為被暴露。
JOHN|3|21|但實行真理的人就來接近光，為要顯明他的行為是靠上帝而行的。」
JOHN|3|22|這些事以後，耶穌和門徒到了 猶太 地區，在那裏他和他們同住，並且施洗。
JOHN|3|23|約翰 也在靠近 撒冷 的 哀嫩 施洗，因為那裏水多，眾人都去受洗。
JOHN|3|24|那時 約翰 還沒有下在監裏。
JOHN|3|25|約翰 的門徒和一個 猶太 人辯論潔淨的禮儀，
JOHN|3|26|就來見 約翰 ，對他說：「拉比，從前同你在 約旦河 的東邊，你所見證的那位，你看，他在施洗，眾人都到他那裏去了。」
JOHN|3|27|約翰 回答說：「若不是從天上賜的，人就不能得到甚麼。
JOHN|3|28|你們自己可以為我作見證，我曾說，我不是基督，只是奉差遣在他前面開路的。
JOHN|3|29|娶新娘的是新郎；新郎的朋友站在一旁聽，一聽見新郎的聲音就歡喜快樂。因此，我這喜樂得以滿足了。
JOHN|3|30|他必興旺；我必衰微。」
JOHN|3|31|「從上頭來的是在萬有之上；出於地的是屬於地，他所說的也是屬於地。從天上來的是在萬有之上。
JOHN|3|32|他把所見所聞的見證出來，只是沒有人領受他的見證。
JOHN|3|33|那領受他見證的，就印證上帝是真實的。
JOHN|3|34|上帝所差來的說上帝的話，因為上帝所賜給他的聖靈是沒有限量的。
JOHN|3|35|父愛子，已把萬有交在他手裏。
JOHN|3|36|信子的人有永生；不信子的人得不到永生，而且上帝的憤怒常在他身上。」
JOHN|4|1|耶穌 知道法利賽人聽見他收門徒和施洗比 約翰 還多， （
JOHN|4|2|其實不是耶穌親自施洗，而是他的門徒施洗，）
JOHN|4|3|他就離開 猶太 ，又回 加利利 去。
JOHN|4|4|他必須經過 撒瑪利亞 ，
JOHN|4|5|於是到了 撒瑪利亞 的一座城，名叫 敘加 ，靠近 雅各 給他兒子 約瑟 的那塊地。
JOHN|4|6|雅各井 就在那裏；耶穌因旅途疲乏，坐在井旁。那時約是正午。
JOHN|4|7|有一個 撒瑪利亞 婦人來打水。耶穌對她說：「請給我水喝。」
JOHN|4|8|因為那時門徒進城買食物去了。
JOHN|4|9|撒瑪利亞 婦人對他說：「你是 猶太 人，怎麼向我一個 撒瑪利亞 女人要水喝呢？」因為 猶太 人和 撒瑪利亞 人沒有來往。
JOHN|4|10|耶穌回答她說：「你若知道上帝的恩賜，和對你說『請給我水喝』的是誰，你早就會求他，他也早就會給了你活水。」
JOHN|4|11|婦人對耶穌說：「先生，你沒有打水的器具，井又深，哪裏去取活水呢？
JOHN|4|12|我們的祖宗 雅各 把這井留給我們，他自己和兒女以及牲畜都喝這井裏的水，難道你比他還大嗎？」
JOHN|4|13|耶穌回答，對她說：「凡喝這水的，還要再渴；
JOHN|4|14|誰喝我所賜的水，就永遠不渴。我所賜的水要在他裏面成為泉源，直湧到永生。」
JOHN|4|15|婦人對他說：「先生，請把這水賜給我，使我不渴，也不用到這裏來打水。」
JOHN|4|16|耶穌對她說：「你去，叫你的丈夫，再到這裏來。」
JOHN|4|17|婦人回答，對耶穌說：「我沒有丈夫。」耶穌說：「你說沒有丈夫是對的。
JOHN|4|18|你已經有過五個丈夫，你現在有的並不是你的丈夫。你這話是真的。」
JOHN|4|19|婦人對他說：「先生，我看你是一位先知。
JOHN|4|20|我們的祖宗在這山上敬拜上帝，你們倒說，應當敬拜的地方是在 耶路撒冷 。」
JOHN|4|21|耶穌對她說：「婦人，你要信我。時候將到，你們敬拜父，既不在這山上，也不在 耶路撒冷 。
JOHN|4|22|你們所敬拜的，你們不知道；我們所敬拜的，我們知道，因為救恩是從 猶太 人出來的。
JOHN|4|23|時候將到，現在就是了，那真正敬拜父的，要用心靈和誠實敬拜他，因為父要這樣的人敬拜他。
JOHN|4|24|上帝是靈，所以敬拜他的必須用心靈和誠實敬拜他。」
JOHN|4|25|婦人對他說：「我知道彌賽亞—就是那稱為基督的—要來；他來了，會把一切的事都告訴我們。」
JOHN|4|26|耶穌對她說：「我就是，正在跟你說話呢！」
JOHN|4|27|正在這時，門徒回來了。他們對耶穌正在和一個婦人說話感到驚訝，可是沒有人說：「你要甚麼？」或說：「你為甚麼和她說話？」
JOHN|4|28|那婦人留下水罐，往城裏去，對眾人說：
JOHN|4|29|「你們來看！有一個人把我素來所做的一切事都說了出來，難道這個人就是基督嗎？」
JOHN|4|30|他們就出城，來到耶穌那裏。
JOHN|4|31|就在這個時候，門徒求耶穌說：「拉比，請吃吧。」
JOHN|4|32|耶穌對他們說：「我有食物吃，是你們不知道的。」
JOHN|4|33|門徒就彼此說：「難道有人拿甚麼給他吃了嗎？」
JOHN|4|34|耶穌對他們說：「我的食物就是要遵行差我來那位的旨意，完成他的工作。
JOHN|4|35|你們不是說『到收割的時候還有四個月』嗎？我告訴你們，舉目向田觀看，莊稼熟了，可以收割了。
JOHN|4|36|收割的人已經得工錢 ，為永生儲存五穀，使撒種的和收割的一同快樂。
JOHN|4|37|『那人撒種，這人收割』，這話可見是真的。
JOHN|4|38|我差你們去收你們所沒有辛勞的；別人辛勞，你們享受他們辛勞的成果。」
JOHN|4|39|那城裏有好些 撒瑪利亞 人信了耶穌，因為那婦人作見證，說：「他把我素來所做的一切事都說了出來。」
JOHN|4|40|於是 撒瑪利亞 人來見耶穌，求他在他們那裏住下，他就在那裏住了兩天。
JOHN|4|41|因為耶穌的話，信的人就更多了。
JOHN|4|42|他們對那婦人說：「現在我們信，不再是因為你的話，而是我們親自聽見了，知道這人真是世界的救主。」
JOHN|4|43|過了那兩天，耶穌離開那地方，往 加利利 去。
JOHN|4|44|因為耶穌自己作過見證說：「先知在自己的家鄉是沒有人尊敬的。」
JOHN|4|45|到了 加利利 ， 加利利 人都歡迎他，因為他們也上 耶路撒冷 去過節，曾經看過他在節期間所做的一切事。
JOHN|4|46|耶穌又到了 加利利 的 迦拿 ，就是他從前變水為酒的地方。有一個大臣，他的兒子在 迦百農 病了。
JOHN|4|47|他聽見耶穌從 猶太 到了 加利利 ，就來見他，求他下去醫治他的兒子，因為他兒子快要死了。
JOHN|4|48|耶穌對他說：「若不看見神蹟奇事，你們總是不信。」
JOHN|4|49|那大臣對他說：「先生，求你趁著我的孩子還沒有死就下去吧。」
JOHN|4|50|耶穌對他說：「回去吧，你的兒子會活！」那人信耶穌所說的話，就回去了。
JOHN|4|51|正下去的時候，他的僕人迎面而來，說他的兒子活了。
JOHN|4|52|他就問甚麼時候見好的。他們對他說：「昨天下午一點鐘熱就退了。」
JOHN|4|53|他就知道這正是耶穌對他說「你的兒子會活」的時候；他自己和全家就都信了。
JOHN|4|54|這是耶穌從 猶太 回到 加利利 後所行的第二個神蹟。
JOHN|5|1|這些事以後，到了 猶太 人的一個節期，耶穌上 耶路撒冷 去。
JOHN|5|2|在 耶路撒冷 ，靠近 羊門 有一個池子， 希伯來 話叫 畢士大 ，旁邊有五個柱廊；
JOHN|5|3|裏面躺著許多病人，有失明的、瘸腿的、癱瘓的 。
JOHN|5|4|
JOHN|5|5|在那裏有一個人，病了三十八年。
JOHN|5|6|耶穌看見他躺著，知道他病了很久，就問他：「你要痊癒嗎？」
JOHN|5|7|病人回答他：「先生，水動的時候，沒有人把我放在池子裏；我正要去的時候，別人比我先下去了。」
JOHN|5|8|耶穌對他說：「起來，拿起你的褥子走吧！」
JOHN|5|9|那人立刻痊癒，就拿起自己的褥子走了。 那天是安息日，
JOHN|5|10|所以 猶太 人對那被治好了的人說：「今天是安息日，你拿褥子是不合法的。」
JOHN|5|11|他卻回答他們：「那使我痊癒的人對我說：『拿起你的褥子走吧！』」
JOHN|5|12|他們問他：「對你說『拿起褥子走』的是甚麼人？」
JOHN|5|13|那治好了的人不知道那人是誰，因為那裏人很多，耶穌已經躲開了。
JOHN|5|14|後來耶穌在聖殿裏找到他，對他說：「你已經痊癒了，不要再犯罪，免得你的遭遇更壞。」
JOHN|5|15|那人就去告訴 猶太 人，使他痊癒的是耶穌。
JOHN|5|16|所以 猶太 人迫害耶穌，因為他在安息日做了這些事。
JOHN|5|17|耶穌就回答他們：「我父做事直到如今，我也做事。」
JOHN|5|18|為了這緣故， 猶太 人越發想要殺他，因為他不但犯了安息日，而且稱上帝為他的父，把自己和上帝看為同等。
JOHN|5|19|於是耶穌回答，對他們說：「我實實在在地告訴你們，子憑著自己不能做甚麼，惟有看見父所做的，他才做；父所做的事，子也照樣做。
JOHN|5|20|父愛子，將自己所做的一切事指示給他看，還要將比這更大的事給他看，使你們驚訝。
JOHN|5|21|父怎樣叫死人復活，賜他們生命，子也照樣隨自己的意願賜人生命。
JOHN|5|22|父不審判任何人，而是把審判的事全交給子，
JOHN|5|23|為要使人都尊敬子，如同尊敬父一樣。不尊敬子的，就是不尊敬差子來的父。
JOHN|5|24|「我實實在在地告訴你們，那聽我話又信差我來那位的，就有永生，不至於被定罪，而是已經出死入生了。
JOHN|5|25|我實實在在地告訴你們，時候將到，現在就是了，死人要聽見上帝兒子的聲音，聽見的人就要活了。
JOHN|5|26|因為父怎樣自己裏面有生命，也照樣賜給他兒子自己裏面有生命，
JOHN|5|27|並且賜給他施行審判的權柄，因為他是人子。
JOHN|5|28|你們不要對這事感到驚訝，因為時候將到，凡在墳墓裏的，都要聽見他的聲音，
JOHN|5|29|並且要出來：行善的，復活得生命；作惡的，復活被定罪。
JOHN|5|30|「我憑著自己不能做甚麼。我怎麼聽見就怎麼審判，而我的審判是公平的，因為我不尋求自己的意願，只尋求差我來那位的旨意。」
JOHN|5|31|「我若為自己作見證，我的見證就不真。
JOHN|5|32|另有一位為我作見證，我也知道他為我作的見證是真的。
JOHN|5|33|你們曾差人到 約翰 那裏，他為真理作過見證。
JOHN|5|34|其實，我所受的見證不是從人來的；然而，我說這些話是為了使你們得救。
JOHN|5|35|約翰 是點亮的明燈，你們情願因他的光歡欣一時。
JOHN|5|36|但我有比 約翰 更大的見證：父交給我去完成的工作，就是我正在做的，為我作證是父差遣了我。
JOHN|5|37|那差我來的父也為我作了見證。你們從來沒有聽見他的聲音，也沒有看見他的形像。
JOHN|5|38|你們並沒有他的道存在心裏，因為你們不信他所差來的那一位。
JOHN|5|39|你們查考聖經，因你們以為其中有永生；而這經正是為我作見證的。
JOHN|5|40|然而，你們不肯到我這裏來得生命。
JOHN|5|41|「我不接受從人來的榮耀，
JOHN|5|42|但我知道，你們沒有愛上帝的心。
JOHN|5|43|我奉我父的名來了，你們並不接納我；若有別人奉自己的名來，你們倒會接納他。
JOHN|5|44|你們互相受榮耀，卻不尋求從獨一上帝來的榮耀，怎能信我呢？
JOHN|5|45|不要以為我會在父面前告你們；有一位告你們的，就是你們所仰望的 摩西 。
JOHN|5|46|如果你們信 摩西 ，也會信我，因為他寫過關於我的事。
JOHN|5|47|你們若不信他的書，怎能信我的話呢？」
JOHN|6|1|這些事以後，耶穌渡過 加利利海 ，就是 提比哩亞海 。
JOHN|6|2|有一大群人因為看見他在病人身上所行的神蹟，就跟隨他。
JOHN|6|3|耶穌上了山，和門徒一同坐在那裏。
JOHN|6|4|那時 猶太 人的逾越節近了。
JOHN|6|5|耶穌舉目看見一大群人來，就對 腓力 說：「我們到哪裏去買餅給這些人吃呢？」
JOHN|6|6|他說這話是要考驗 腓力 ，他自己原知道要怎樣做。
JOHN|6|7|腓力 回答他：「就是兩百個銀幣的餅也不夠給他們每人吃一點點。」
JOHN|6|8|有一個門徒，就是 西門．彼得 的弟弟 安得烈 ，對耶穌說：
JOHN|6|9|「這裏有一個孩子，帶著五個大麥餅和兩條魚，但是分給這麼多人還算甚麼呢？」
JOHN|6|10|耶穌說：「你們叫大家坐下。」那地方的草多，人們就坐下，男人的數目約有五千。
JOHN|6|11|耶穌拿起餅來，祝謝了，就分給坐著的人，也同樣分了魚，都照他們所要的來分。
JOHN|6|12|他們吃飽後，耶穌對門徒說：「把剩下的碎屑收拾起來，免得糟蹋了。」
JOHN|6|13|他們就把那五個大麥餅的碎屑，就是大家吃剩的，收拾起來，裝滿了十二個籃子。
JOHN|6|14|人們看見耶穌所行的神蹟，就說：「這真是那要到世上來的先知！」
JOHN|6|15|耶穌知道他們要來強迫他作王，就獨自又退到山上去了。
JOHN|6|16|到了晚上，他的門徒下到海邊，
JOHN|6|17|上了船，要過海往 迦百農 去。天已經黑了，耶穌還沒有來到他們那裏。
JOHN|6|18|忽然狂風大作，海浪翻騰。
JOHN|6|19|門徒搖櫓，約行了十里多 ，看見耶穌在海面上走，漸漸靠近了船，他們就害怕。
JOHN|6|20|耶穌對他們說：「是我，不要怕！」
JOHN|6|21|門徒就欣然接他上船，船立刻到了他們所要去的地方。
JOHN|6|22|第二天，留在海的對岸的眾人發覺那裏原來只有一條小船，而且耶穌沒有同他的門徒上船，是門徒自己去的。
JOHN|6|23|另外有幾條從 提比哩亞 來的小船，卻停靠在主祝謝後給他們吃餅的地方附近。
JOHN|6|24|這時眾人見耶穌和門徒都不在那裏，就上了船，往 迦百農 去找耶穌。
JOHN|6|25|他們在海的對岸找到他後，對他說：「拉比，你幾時到這裏來的？」
JOHN|6|26|耶穌回答他們說：「我實實在在地告訴你們，你們找我，並不是因見了神蹟，而是因吃餅吃飽了。
JOHN|6|27|不要為那會壞的食物操勞，而要為那存到永生的食物操勞。這食物是人子要賜給你們的，因為父上帝已印證了。」
JOHN|6|28|於是他們問他：「我們該做甚麼才算是做上帝的工作呢？」
JOHN|6|29|耶穌回答，對他們說：「信上帝所差來的，這就是上帝的工作。」
JOHN|6|30|於是他們對他說：「你行甚麼神蹟，好讓我們看見而信你呢？你到底要做甚麼呢？
JOHN|6|31|我們的祖宗在曠野吃過嗎哪，如經上寫著：『他從天上賜下糧食來給他們吃。』」
JOHN|6|32|於是耶穌對他們說：「我實實在在地告訴你們，那從天上來的糧不是 摩西 賜給你們的，那從天上來的真糧是我父賜給你們的。
JOHN|6|33|因為上帝的糧就是那位從天上降下來，並且賜生命給世界的。」
JOHN|6|34|於是他們對他說：「主啊，請常常把這糧賜給我們！」
JOHN|6|35|耶穌對他們說：「我就是生命的糧。到我這裏來的，絕不飢餓；信我的，永不乾渴。
JOHN|6|36|可是，我告訴過你們，你們已經看見我 ，還是不信。
JOHN|6|37|凡父所賜給我的人，必到我這裏來；到我這裏來的，我總不丟棄他。
JOHN|6|38|因為我從天上降下來，不是要按自己的意願行，而是要遵行差我來那位的旨意。
JOHN|6|39|差我來那位的旨意就是：他所賜給我的，要我一個也不失落，並且在末日使他復活。
JOHN|6|40|因為我父的旨意是要使每一個見了子而信的人得永生，並且在末日我要使他復活。」
JOHN|6|41|猶太 人因為耶穌說「我是從天上降下來的糧」，就私下議論他，
JOHN|6|42|說：「這不是 約瑟 的兒子耶穌嗎？我們豈不認得他的父母嗎？現在他怎麼說『我是從天上降下來的』呢？」
JOHN|6|43|耶穌回答，對他們說：「你們不要彼此私下議論。
JOHN|6|44|若不是差我來的父吸引人，就沒有人能到我這裏來；到我這裏來的，在末日我要使他復活。
JOHN|6|45|在先知書上寫著：『他們都要蒙上帝教導。』凡聽了父的教導而學習的，都到我這裏來。
JOHN|6|46|這不是說有人看見過父，惟獨從上帝來的，他才看見過父。
JOHN|6|47|我實實在在地告訴你們，信的人有永生。
JOHN|6|48|我就是生命的糧。
JOHN|6|49|你們的祖宗在曠野吃過嗎哪，還是死了。
JOHN|6|50|這是從天上降下來的糧，使人吃了就不死。
JOHN|6|51|我就是從天上降下來生命的糧；人若吃這糧，必永遠活著。我為世人的生命所賜下的糧就是我的肉。」
JOHN|6|52|因此， 猶太 人彼此爭論說：「這個人怎能把他的肉給我們吃呢？」
JOHN|6|53|耶穌對他們說：「我實實在在地告訴你們，你們若不吃人子的肉，不喝人子的血，在你們裏面就沒有生命。
JOHN|6|54|吃我肉、喝我血的人就有永生，並且在末日我要使他復活。
JOHN|6|55|我的肉是真正可吃的；我的血是真正可喝的。
JOHN|6|56|吃我肉、喝我血的人常在我裏面，我也常在他裏面。
JOHN|6|57|永生的父怎樣差我來，我又怎樣因父活著，照樣，吃我肉的人也要因我活著。
JOHN|6|58|這是從天上降下來的糧，不像你們的祖宗吃過嗎哪還是死了；吃這糧的人將永遠活著。」
JOHN|6|59|這些話是耶穌在 迦百農 會堂裏教導人的時候說的。
JOHN|6|60|他的門徒中有好些人聽見了，就說：「這話很難，誰聽得進呢？」
JOHN|6|61|耶穌心裏知道門徒為這話私下議論，就對他們說：「這話成了你們的絆腳石嗎？
JOHN|6|62|如果你們看見人子升到他原來所在之處，會怎麼樣呢？
JOHN|6|63|聖靈賜人生命，肉體毫無用處。我對你們所說的話就是靈，就是生命。
JOHN|6|64|可是你們中間有些人不信。」耶穌起初就知道哪些人不信他，哪一個要出賣他。
JOHN|6|65|於是耶穌說：「所以，我對你們說過，若不是蒙我父的恩賜，沒有人能到我這裏來。」
JOHN|6|66|從此，他門徒中有很多退卻了，不再和他同行。
JOHN|6|67|耶穌就對那十二使徒說：「你們也要離開嗎？」
JOHN|6|68|西門．彼得 回答他：「主啊，你有永生之道，我們還跟從誰呢？
JOHN|6|69|我們已經信了，又知道你是上帝的聖者。」
JOHN|6|70|耶穌回答他們：「我不是揀選了你們十二個嗎？但你們中間有一個是魔鬼。」
JOHN|6|71|耶穌這話是指著要出賣他的 加略 人 西門 的兒子 猶大 說的；他本是十二使徒裏的一個。
JOHN|7|1|這些事以後，耶穌周遊 加利利 ，不願在 猶太 往來，因為 猶太 人想要殺他。
JOHN|7|2|這時 猶太 人的住棚節近了。
JOHN|7|3|耶穌的兄弟們對他說：「你離開這裏上 猶太 去吧，好讓你的門徒也看見你所做的事。
JOHN|7|4|因為人要揚名，沒有在隱祕的地方行事的，如果你要做這些事，該把自己顯明給世人看。」
JOHN|7|5|原來連他的兄弟們也不信他。
JOHN|7|6|於是耶穌對他們說：「我的時機還沒有到，你們的時機卻隨時都有。
JOHN|7|7|世人不會恨你們，卻是恨我，因為我指證他們的行為是惡的。
JOHN|7|8|你們上去過節吧！我現在不上去過這節 ，因為我的時機還沒有成熟。」
JOHN|7|9|耶穌說了這些話，仍然留在 加利利 。
JOHN|7|10|但他的兄弟們上去過節以後，他也上去，不是公開去，卻似乎 是祕密地去的。
JOHN|7|11|節期間， 猶太 人尋找耶穌，說：「他在哪裏？」
JOHN|7|12|人群中有許多人對他議論紛紛，另有的說：「他是好人。」有的說：「不，他是迷惑群眾的。」
JOHN|7|13|可是沒有人公開談論他，因為他們怕 猶太 人。
JOHN|7|14|節期已過了一半，耶穌上聖殿去教導人。
JOHN|7|15|猶太 人驚訝地說：「這個人沒有學過，怎麼那樣熟悉經典呢？」
JOHN|7|16|於是耶穌回答他們，說：「我的教導不是我自己的，而是差我來那位的。
JOHN|7|17|人若立志要遵行上帝的旨意，就會知道這教導究竟是出於上帝，還是我憑著自己說的。
JOHN|7|18|憑著自己說的人是尋求自己的榮耀；但那尋求差他來那位的榮耀的人，他是真誠的，在他心裏沒有不義。
JOHN|7|19|摩西 不是傳了律法給你們嗎？你們卻沒有一個人守律法。為甚麼想要殺我呢？」
JOHN|7|20|眾人回答：「你是被鬼附了！誰想要殺你呢？」
JOHN|7|21|耶穌回答，對他們說：「我做了一件事，你們都驚訝。
JOHN|7|22|摩西 傳割禮給你們（其實割禮不是從 摩西 開始，而是從列祖開始的），你們就在安息日給人行割禮。
JOHN|7|23|人若在安息日受割禮，是為了不違背 摩西 的律法，我在安息日使一個人痊癒了，你們就向我發怒嗎？
JOHN|7|24|不要憑外表斷定是非，總要按公平斷定是非。」
JOHN|7|25|於是 耶路撒冷 人中有的說：「這個人不是他們想要殺的嗎？
JOHN|7|26|你看，他還公開講道，他們也不對他說甚麼。難道官長真的認為這是基督嗎？
JOHN|7|27|然而，我們知道這個人從哪裏來；可是基督來的時候，沒有人知道他從哪裏來。」
JOHN|7|28|那時，耶穌在聖殿裏教導人，喊著說：「你們認識我，也知道我從哪裏來；我並不是憑著自己來的。但差我來的那位是真實的，你們不認識他。
JOHN|7|29|我卻認識他，因為我從他那裏來，是他差遣了我。」
JOHN|7|30|於是他們想要捉拿耶穌，只是沒有人下手，因為他的時候還沒有到。
JOHN|7|31|但人群中有好些人信他，他們說：「基督來的時候，他所行的神蹟難道會比這人行的更多嗎？」
JOHN|7|32|法利賽人聽見群眾對耶穌這樣議論紛紛，祭司長和法利賽人就打發聖殿警衛去捉拿他。
JOHN|7|33|於是耶穌說：「我跟你們在一起的時候不會太久了，我要回到那差我來的那裏去。
JOHN|7|34|你們要找我，卻找不到；我所在的地方，你們不能去。」
JOHN|7|35|於是 猶太 人彼此問：「這人要往哪裏去，使我們找不到他呢？難道他要往散居在 希臘 的 猶太 人那裏去教導 希臘 人嗎？
JOHN|7|36|他說『你們要找我，卻找不到；我所在的地方，你們不能去』這話是甚麼意思呢？」
JOHN|7|37|節期的最後一天，就是最隆重的一天，耶穌站著，喊著說：「人若渴了，到我這裏來喝！
JOHN|7|38|信我的人，就如經上所說：『從他腹中將流出活水的江河來。』」
JOHN|7|39|耶穌這話是指信他的人要受聖靈說的；那時還沒有賜下聖靈，因為耶穌還沒有得到榮耀。
JOHN|7|40|眾人聽見這些話，有的說：「這真是那先知。」
JOHN|7|41|另有的說：「這是基督。」但也有的說：「難道基督是出自 加利利 嗎？
JOHN|7|42|經上不是說『基督是 大衛 的後裔，出自 大衛 的本鄉 伯利恆 』嗎？」
JOHN|7|43|於是眾人因耶穌而分裂了。
JOHN|7|44|其中有人要捉拿他，只是沒有人下手。
JOHN|7|45|警衛們回到祭司長和法利賽人那裏。他們對警衛說：「你們為甚麼沒有帶他來呢？」
JOHN|7|46|警衛回答：「從來沒有像他這樣說話的！」
JOHN|7|47|於是法利賽人說：「你們也受了迷惑嗎？
JOHN|7|48|難道官長或法利賽人中有信他的嗎？
JOHN|7|49|但這些不明白律法的眾人是被詛咒的！」
JOHN|7|50|其中有 尼哥德慕 ，就是從前去見過耶穌的，對他們說：
JOHN|7|51|「不先聽本人的口供，查明他所做的事，難道我們的律法還定他的罪嗎？」
JOHN|7|52|他們回答他說：「你也是出自 加利利 嗎？你去查考就知道， 加利利 是不出先知的。」 〔
JOHN|7|53|於是各人都回家去了，
JOHN|8|1|耶穌卻到 橄欖山 去。
JOHN|8|2|清早，他又回到聖殿裏。眾百姓都到他那裏去，他就坐下，教導他們。
JOHN|8|3|文士和法利賽人帶著一個犯姦淫時被捉的女人來，叫她站在當中，
JOHN|8|4|然後對耶穌說：「老師，這女人是正在犯姦淫的時候被捉到的。
JOHN|8|5|摩西 在律法書上命令我們把這樣的女人用石頭打死。那麼，你怎麼說呢？」
JOHN|8|6|他們說這話是要試探耶穌，要抓到控告他的把柄。耶穌卻彎下腰，用指頭在地上寫字。
JOHN|8|7|他們還是不住地問他，耶穌就直起腰來，對他們說：「你們中間誰沒有罪，誰就先拿石頭打她！」
JOHN|8|8|於是他又彎著腰，用指頭在地上寫字。
JOHN|8|9|他們聽見這話，從老的開始，一個一個都走開了，只剩下耶穌一人和那仍然站在中間的女人。
JOHN|8|10|耶穌就直起腰來，對她說：「婦人，那些人在哪裏呢？沒有任何人定你的罪嗎？」
JOHN|8|11|她說：「主啊，沒有。」耶穌說：「我也不定你的罪。去吧！從今以後不要再犯罪了。」〕
JOHN|8|12|耶穌又對眾人說：「我就是世界的光。跟從我的，必不在黑暗裏走，卻要得著生命的光。」
JOHN|8|13|法利賽人對他說：「你是為自己作見證，你的見證不真。」
JOHN|8|14|耶穌回答他們，對他們說：「即使我為自己作見證，我的見證還是真的，因為我知道我從哪裏來，到哪裏去。你們卻不知道我從哪裏來，到哪裏去。
JOHN|8|15|你們是以人的標準來判斷人，我不判斷任何人。
JOHN|8|16|即使我判斷人，我的判斷也是真確的，因為不是我獨自在判斷，而是差我來的父與我一同判斷。
JOHN|8|17|你們的律法也記著說：『兩個人的見證才算為真』。
JOHN|8|18|我是為自己作見證，還有差我來的父也為我作見證。」
JOHN|8|19|於是他們問他：「你的父在哪裏？」耶穌回答：「你們不認識我，也不認識我的父；若是認識我，也會認識我的父。」
JOHN|8|20|這些話是耶穌在聖殿的銀庫房裏教導人的時候說的。當時沒有人捉拿他，因為他的時候還沒有到。
JOHN|8|21|於是耶穌又對他們說：「我去了，你們會找我，而你們會死在自己的罪中；我所去的地方，你們不能去。」
JOHN|8|22|猶太 人說：「他說『我所去的地方，你們不能去』，難道他要自殺嗎？」
JOHN|8|23|耶穌對他們說：「你們是從下面來的，我是從上面來的；你們是屬這世界的，我不是屬這世界的。
JOHN|8|24|所以我對你們說，你們會死在自己的罪中，你們若不信我就是那位，就會死在自己的罪中。」
JOHN|8|25|他們就問他：「你到底是誰？」耶穌對他們說：「我從起初就告訴你們了。
JOHN|8|26|我有許多事要講論你們，判斷你們；但差我來的那位是真實的，我從他那裏所聽見的，就告訴世人。」
JOHN|8|27|他們不明白耶穌是對他們講父的事。
JOHN|8|28|所以耶穌說：「你們舉起人子以後就會知道我就是那位了，並且知道我沒有一件事是憑著自己做的。我說這些話是照著父所教導我的。
JOHN|8|29|差我來的那位與我同在；他沒有撇下我獨自一人，因為我一直行他所喜悅的事。」
JOHN|8|30|耶穌說這些話的時候，有許多人信了他。
JOHN|8|31|耶穌對信他的 猶太 人說：「你們若繼續遵守我的道，就真是我的門徒了。
JOHN|8|32|你們將認識真理，真理會使你們自由。」
JOHN|8|33|他們回答他：「我們是 亞伯拉罕 的後裔，從來沒有作過誰的奴隸，你怎麼說『會使你們自由』呢？」
JOHN|8|34|耶穌回答他們：「我實實在在地告訴你們，所有犯罪的人就是罪的奴隸。
JOHN|8|35|奴隸不能永遠住在家裏；兒子才永遠住在家裏。
JOHN|8|36|所以，上帝的兒子若使你們自由，你們就真正自由了。」
JOHN|8|37|「我知道，你們是 亞伯拉罕 的後裔，你們卻想要殺我，因為你們心裏容不下我的道。
JOHN|8|38|我所說的是在我父那裏看見的；你們所做的是在你們的父那裏聽到的。」
JOHN|8|39|他們回答耶穌：「我們的父是 亞伯拉罕 。」耶穌對他們說：「你們若是 亞伯拉罕 的兒女，就會做 亞伯拉罕 所做的事。
JOHN|8|40|我把在上帝那裏所聽見的真理告訴了你們，現在你們卻想要殺我； 亞伯拉罕 沒有做過這樣的事。
JOHN|8|41|你們是做你們父的工作。」他們就對他說：「我們不是從淫亂生的，我們只有一位父，就是上帝。」
JOHN|8|42|耶穌對他們說：「假如上帝是你們的父，你們會愛我，因為我本是出於上帝，也是從上帝而來，我不是憑著自己來，而是他差我來的。
JOHN|8|43|你們為甚麼不明白我的話呢？無非是你們聽不進我的道。
JOHN|8|44|你們是出於你們的父魔鬼，你們寧願隨著你們父的慾念而行。他從起初就是殺人的，不守真理，因他心裏沒有真理。他說謊是出於自己的本性，因他本來是說謊的，也是說謊者之父。
JOHN|8|45|但是，因為我講真理，你們就不信我。
JOHN|8|46|你們中間誰能指證我有罪呢？既然我講真理，你們為甚麼不信我呢？
JOHN|8|47|出於上帝的，必聽上帝的話；你們不聽，因為你們不是出於上帝。」
JOHN|8|48|猶太 人回答他：「我們說你是 撒瑪利亞 人，並且是被鬼附的，這話不是很對嗎？」
JOHN|8|49|耶穌回答：「我沒有被鬼附的；我尊敬我的父，你們卻不尊敬我。
JOHN|8|50|我不尋求自己的榮耀，但有一位為我尋求榮耀，判斷是非。
JOHN|8|51|我實實在在地告訴你們，人若遵守我的道，就永遠不經歷死亡。」
JOHN|8|52|於是 猶太 人對他說：「現在我們知道你是被鬼附了。 亞伯拉罕 死了，眾先知也死了，你還說：『人若遵守我的道，就永遠不經歷死亡。』
JOHN|8|53|難道你比我們的祖宗 亞伯拉罕 還大嗎？他死了，眾先知也死了，你把自己當作甚麼人呢？」
JOHN|8|54|耶穌回答：「我若榮耀自己，我的榮耀就算不了甚麼；榮耀我的是我的父，就是你們所說的你們的上帝。
JOHN|8|55|你們不認識他，我卻認識他。我若說不認識他，我就是說謊的，像你們一樣；但我認識他，也遵守他的道。
JOHN|8|56|你們的祖宗 亞伯拉罕 歡歡喜喜地仰望我的日子，他看見了，就快樂。」
JOHN|8|57|猶太 人就對他說：「你還沒有五十歲，難道見過 亞伯拉罕 嗎？」
JOHN|8|58|耶穌對他們說：「我實實在在地告訴你們，還沒有 亞伯拉罕 我就存在了。」
JOHN|8|59|於是他們拿石頭要打他，耶穌卻躲開，走出了聖殿。
JOHN|9|1|耶穌往前走的時候，看見一個生來就失明的人。
JOHN|9|2|門徒問耶穌：「拉比，這人生來失明，是誰犯了罪？是這人還是他的父母呢？」
JOHN|9|3|耶穌回答：「既不是這人犯了罪，也不是他的父母，而是要在他身上顯出上帝的作為來。
JOHN|9|4|趁著白日，我們 必須做差我 來的那位的工；黑夜來到，就沒有人能做工了。
JOHN|9|5|我在世上的時候，是世上的光。」
JOHN|9|6|耶穌說了這些話，就吐唾沫在地上，用唾沫和了泥抹在盲人的眼睛上，
JOHN|9|7|對他說：「你到 西羅亞 池子裏去洗。」（ 西羅亞 翻出來就是「奉差遣」。）於是他去，洗了，回來就看見了。
JOHN|9|8|他的鄰舍和素常見他討飯的人，就說：「這不是那從前坐著討飯的人嗎？」
JOHN|9|9|有的說：「是他」；又有的說：「不是，卻是像他。」他自己說：「是我。」
JOHN|9|10|於是他們對他說：「你的眼睛是怎麼開的呢？」
JOHN|9|11|那人回答：「有一個名叫耶穌的，他和了泥抹我的眼睛，對我說：『你到 西羅亞 池子去洗。』我去一洗，就看見了。」
JOHN|9|12|他們對他說：「那個人在哪裏？」他說：「我不知道。」
JOHN|9|13|他們把以前失明的那個人帶到法利賽人那裏。
JOHN|9|14|耶穌和泥開他眼睛的那一天是安息日。
JOHN|9|15|法利賽人又問他是怎麼得看見的。他對他們說：「他把泥抹在我的眼睛上，我一洗，就看見了。」
JOHN|9|16|於是法利賽人中有的說：「這個人不是從上帝來的，因為他不守安息日。」另有的說：「一個罪人怎能行這樣的神蹟呢？」他們之間就產生了分裂。
JOHN|9|17|於是他們又對那盲人說：「他開了你的眼睛，你說他是怎樣的人呢？」他說：「他是個先知。」
JOHN|9|18|猶太 人不信他以前是失明，後來能看見的，等到叫了他的父母來，
JOHN|9|19|問他們說：「這是你們的兒子嗎？你們說他生來是失明的，現在怎麼看見了呢？」
JOHN|9|20|他的父母就回答說：「他是我們的兒子，生來就失明，這是我們知道的。
JOHN|9|21|至於他現在怎麼能看見，我們卻不知道；是誰開了他的眼睛，我們也不知道。他已經是成人，你們問他吧，他自己會說。」
JOHN|9|22|他父母說這些話，是怕 猶太 人，因為 猶太 人已經商定，若有宣認耶穌是基督的，要把他趕出會堂。
JOHN|9|23|因此他父母說「他已經是成人，你們問他吧」。
JOHN|9|24|於是法利賽人第二次叫了那以前失明的人來，對他說：「你要將榮耀歸給上帝，我們知道這人是個罪人。」
JOHN|9|25|那人就回答：「他是不是個罪人，我不知道；有一件事我知道，我本來是失明的，現在我看見了。」
JOHN|9|26|他們就問他：「他給你做了甚麼？是怎麼開了你的眼睛？」
JOHN|9|27|他回答他們：「我已經告訴你們了，你們不聽，為甚麼又要聽呢？難道你們也要作他的門徒嗎？」
JOHN|9|28|他們就罵他：「你是他的門徒，而我們是 摩西 的門徒。
JOHN|9|29|上帝對 摩西 說話是我們知道的，可是這個人，我們不知道他從哪裏來。」
JOHN|9|30|那人回答，對他們說：「他開了我的眼睛，你們竟不知道他從哪裏來，這真是奇怪！
JOHN|9|31|我們知道上帝不聽罪人，惟有敬奉上帝、遵行他旨意的，上帝才聽他。
JOHN|9|32|從創世以來，未曾聽見有人開了生來就失明的人的眼睛。
JOHN|9|33|這人若不是從上帝來的，甚麼也不能做。」
JOHN|9|34|他們回答他說：「你完全是生在罪中的，還要來教訓我們嗎？」於是他們把他趕出去了。
JOHN|9|35|耶穌聽說他們把他趕出去，就找到他，說：「你信人子 嗎？」
JOHN|9|36|那人回答說：「主啊，人子是誰？告訴我，好讓我信他。」
JOHN|9|37|耶穌對他說：「你已經看見他，現在和你說話的就是他。」
JOHN|9|38|他說：「主啊，我信！」他就拜耶穌。
JOHN|9|39|耶穌說：「我為審判到這世上來，使不能看見的看見，能看見的反而失明。」
JOHN|9|40|同他在那裏的法利賽人聽見這些話，就對他說：「難道我們也失明了嗎？」
JOHN|9|41|耶穌對他們說：「你們若是失明的，就沒有罪了；但現在你們說『我們能看見』，你們的罪還在。」
JOHN|10|1|「我實實在在地告訴你們，那不從門進羊圈，倒從別處爬進去的，就是賊，就是強盜。
JOHN|10|2|那從門進去的才是羊的牧人。
JOHN|10|3|看門的給他開門，羊也聽他的聲音。他按著名叫自己的羊，把羊領出來。
JOHN|10|4|當他把自己的羊都放出來，就走在前面，羊也跟著他，因為牠們認得他的聲音。
JOHN|10|5|羊絕不跟陌生人，反而會逃走，因為不認得陌生人的聲音。」
JOHN|10|6|耶穌把這比方告訴他們，但他們不明白他所說的是甚麼。
JOHN|10|7|所以，耶穌又對他們說：「我實實在在地告訴你們，我就是羊的門。
JOHN|10|8|凡在我以前 來的都是賊，是強盜；羊沒有聽從他們。
JOHN|10|9|我就是門，凡從我進來的，必得安全 ，並且可進出，找到草吃。
JOHN|10|10|盜賊來，無非要偷竊，殺害，毀壞；我來了，是要羊得生命，並且得的更豐盛。
JOHN|10|11|「我是好牧人，好牧人為羊捨命。
JOHN|10|12|雇工不是牧人，羊不是他自己的，他一看見狼來，就撇下羊群逃跑；狼抓住羊，把牠們趕散。
JOHN|10|13|雇工逃走，因為他是雇工，對羊毫不關心。
JOHN|10|14|我是好牧人；我認識我的羊，我的羊也認識我，
JOHN|10|15|正如父認識我，我也認識父一樣；並且我為羊捨命。
JOHN|10|16|我另外有羊，不屬這圈裏的，我必須領牠們來，牠們也要聽我的聲音，並且要合成一群，歸一個牧人。
JOHN|10|17|為此，我父愛我，因為我把命捨去，好再取回來。
JOHN|10|18|沒有人奪去我的命，是我自己捨的；我有權捨棄，也有權再取回。這是我從我父所受的命令。」
JOHN|10|19|猶太 人為這些話又起了分裂。
JOHN|10|20|其中有好些人說：「他是被鬼附了，而且瘋了，為甚麼聽他的呢？」
JOHN|10|21|另有的說：「這不是被鬼附的人所說的話。鬼豈能開盲人的眼睛呢？」
JOHN|10|22|那時正是冬天，在 耶路撒冷 有獻殿節。
JOHN|10|23|耶穌在聖殿裏的 所羅門 廊下行走。
JOHN|10|24|猶太 人圍著他，對他說：「你讓我們猶豫不定到幾時呢？你若是基督，就明白地告訴我們。」
JOHN|10|25|耶穌回答他們：「我已經告訴你們，你們卻不信。我奉我父的名所行的事可以為我作見證。
JOHN|10|26|但是你們不信，因為你們不是我的羊。
JOHN|10|27|我的羊聽我的聲音，我認識牠們，牠們也跟從我。
JOHN|10|28|並且，我賜給他們永生；他們永不滅亡，誰也不能從我手裏把他們奪去。
JOHN|10|29|我父所賜給我的比萬有都大 ，誰也不能從我父手裏把他們奪去。
JOHN|10|30|我與父原為一。」
JOHN|10|31|猶太 人又拿起石頭來要打他。
JOHN|10|32|耶穌回應他們：「我做了許多從父那裏來的善事給你們看，你們是為哪一件拿石頭打我呢？」
JOHN|10|33|猶太 人回答他：「我們不是為了善事拿石頭打你，而是為了你說褻瀆的話；因為你是個人，卻把自己當作上帝。」
JOHN|10|34|耶穌回答他們：「你們的律法書上不是寫著『我曾說你們是諸神』嗎？
JOHN|10|35|經上的話是不能廢的；如果那些領受上帝的道的人，上帝尚且稱他們為諸神，
JOHN|10|36|那麼父所分別為聖又差到世上來的那位說『我是上帝的兒子』，你們還對他說『你說褻瀆的話』嗎？
JOHN|10|37|我若不做我父的工作，你們就不必信我；
JOHN|10|38|我若做了，你們即使不信我，也當信這些工作，好讓你們知道並且明白父在我裏面，我也在父裏面。」
JOHN|10|39|於是，他們又要捉拿他，他卻從他們手中逃脫了。
JOHN|10|40|耶穌又往 約旦河 的東邊去，到了 約翰 起初施洗的地方，就住在那裏。
JOHN|10|41|有許多人來到他那裏，說：「 約翰 沒有行過一件神蹟，但 約翰 所說有關這人的一切話都是真的。」
JOHN|10|42|在那裏，許多人信了耶穌。
JOHN|11|1|有一個患病的人，名叫 拉撒路 ，住在 伯大尼 ，就是 馬利亞 和她姐姐 馬大 的村莊。
JOHN|11|2|這 馬利亞 就是那用香膏抹主，又用頭髮擦他腳的；患病的 拉撒路 是她的弟弟。
JOHN|11|3|姊妹兩個就打發人去見耶穌，說：「主啊，你所愛的人病了。」
JOHN|11|4|耶穌聽見後卻說：「這病不至於死，而是為了上帝的榮耀，為要使上帝的兒子藉此得榮耀。」
JOHN|11|5|耶穌素來愛 馬大 和她妹妹，以及 拉撒路 。
JOHN|11|6|他聽見 拉撒路 病了，仍在原地住了兩天，
JOHN|11|7|然後對門徒說：「我們再到 猶太 去吧！」
JOHN|11|8|門徒對他說：「拉比， 猶太 人近來要拿石頭打你，你還再到那裏去嗎？」
JOHN|11|9|耶穌回答：「白天不是有十二小時嗎？人若在白天行走，就不致跌倒，因為他看見這世上的光。
JOHN|11|10|人若在黑夜行走，就會跌倒，因為他沒有光。」
JOHN|11|11|耶穌說了這些話，隨後對他們說：「我們的朋友 拉撒路 睡了，我去叫醒他。」
JOHN|11|12|門徒就說：「主啊，他若睡了，就會好的。」
JOHN|11|13|耶穌說這話是指 拉撒路 死了，他們卻以為他是指通常的睡眠。
JOHN|11|14|於是耶穌就明白地告訴他們：「 拉撒路 死了。
JOHN|11|15|為了你們的緣故，我不在那裏反而歡喜，為要使你們信。現在我們到他那裏去吧。」
JOHN|11|16|於是那稱為 低土馬 的 多馬 對其他的門徒說：「我們也去和他同死吧！」
JOHN|11|17|耶穌到了，知道 拉撒路 在墳墓裏已經四天了。
JOHN|11|18|伯大尼 離 耶路撒冷 不遠，約有六里 路。
JOHN|11|19|有好些 猶太 人來看 馬大 和 馬利亞 ，要為她們弟弟的緣故安慰她們。
JOHN|11|20|馬大 聽見耶穌來了，就出去迎接他； 馬利亞 卻仍然坐在家裏。
JOHN|11|21|馬大 對耶穌說：「主啊，你若早在這裏，我弟弟就不會死了。
JOHN|11|22|我也知道，即使現在，你無論向上帝求甚麼，上帝也必賜給你。」
JOHN|11|23|耶穌對她說：「你弟弟會復活的。」
JOHN|11|24|馬大 對他說：「我知道在末日復活的時候，他會復活。」
JOHN|11|25|耶穌對她說：「復活在我，生命也在我 。信我的人雖然死了，也必復活；
JOHN|11|26|凡活著信我的人必永遠不死。你信這話嗎？」
JOHN|11|27|馬大 對他說：「主啊，是的。我信你是基督，是上帝的兒子，就是那要臨到世界的。」
JOHN|11|28|馬大 說了這話就回去，叫她妹妹 馬利亞 ，私下說：「老師來了，他在叫你。」
JOHN|11|29|馬利亞 聽見了，急忙起來，到耶穌那裏去。
JOHN|11|30|那時，耶穌還沒有進村子，仍在 馬大 迎接他的地方。
JOHN|11|31|那些同 馬利亞 在家裏安慰她的 猶太 人，見她急忙起來，出去，就跟著她，以為她要往墳墓那裏去哭。
JOHN|11|32|馬利亞 到了耶穌那裏，看見他，就俯伏在他腳前，對他說：「主啊，你若早在這裏，我弟弟就不會死了。」
JOHN|11|33|耶穌看見她哭，並看見與她同來的 猶太 人也哭，就心裏悲嘆，又甚憂愁，
JOHN|11|34|就說：「你們把他安放在哪裏？」他們對他說：「主啊，請你來看。」
JOHN|11|35|耶穌哭了。
JOHN|11|36|猶太 人就說：「你看，他多麼愛他！」
JOHN|11|37|其中有人說：「他既然開了盲人的眼睛，難道不能叫這人不死嗎？」
JOHN|11|38|耶穌又心裏悲嘆，來到墳墓前。那墳墓是個穴，有一塊石頭擋著。
JOHN|11|39|耶穌說：「把石頭挪開！」那死者的姐姐 馬大 對他說：「主啊，他現在必定臭了，因為他已經死了四天了。」
JOHN|11|40|耶穌對她說：「我不是對你說過，你若信就必看見上帝的榮耀嗎？」
JOHN|11|41|於是他們把石頭挪開。耶穌舉目望天，說：「父啊，我感謝你，因為你已經聽了我。
JOHN|11|42|我知道你常常聽我，但我說這話是為了周圍站著的眾人，要使他們信是你差了我來的。」
JOHN|11|43|說了這些話，他大聲呼叫說：「 拉撒路 ，出來！」
JOHN|11|44|那死了的人就出來了，手腳都裹著布，臉上包著頭巾。耶穌對他們說：「解開他，讓他走！」
JOHN|11|45|於是來看 馬利亞 的 猶太 人中，有很多人見了耶穌所做的事，就信了他。
JOHN|11|46|但其中也有人去見法利賽人，把耶穌所做的事告訴他們。
JOHN|11|47|祭司長和法利賽人召開議會，說：「這人行好些神蹟，我們怎麼辦呢？
JOHN|11|48|若讓他這樣做，人人都要信他； 羅馬 人也要來毀滅我們的聖殿 和我們的民族。」
JOHN|11|49|其中有一個人，名叫 該亞法 ，那年當大祭司，對他們說：「你們甚麼都不知道，
JOHN|11|50|也不想想，一個人替百姓死，免得整個民族滅亡，這對你們是有利的。」
JOHN|11|51|他這話不是出於自己的意思，而是因他那年當大祭司，所以預言耶穌將為這民族而死。
JOHN|11|52|他不但替這民族死，還要把上帝四散的兒女都聚集起來，合成一群。
JOHN|11|53|從那日起，他們就商議要殺耶穌。
JOHN|11|54|所以，耶穌不再公開在 猶太 人中走動，卻離開那裏，往靠近曠野的鄉間去，到了一座城，名叫 以法蓮 ，就在那裏和門徒住下來。
JOHN|11|55|猶太 人的逾越節近了，有許多人從鄉下上 耶路撒冷 去，要在過節前潔淨自己。
JOHN|11|56|於是他們尋找耶穌，站在聖殿裏彼此說：「你們認為怎樣，他不會來過節吧？」
JOHN|11|57|那時，祭司長和法利賽人早已下令，若有人知道耶穌的下落，就要報告，他們好去捉拿他。
JOHN|12|1|逾越節前六天，耶穌來到 伯大尼 ，就是他使 拉撒路 從死人中復活的地方。
JOHN|12|2|有人在那裏為耶穌預備宴席； 馬大 伺候， 拉撒路 也在同耶穌坐席的人中間。
JOHN|12|3|馬利亞 拿著一斤極貴的純哪噠 香膏，抹耶穌的腳，又用自己頭髮去擦，屋裏充滿了膏的香氣。
JOHN|12|4|有一個門徒，就是那將要出賣耶穌的 加略 人 猶大 ，說：
JOHN|12|5|「為甚麼不把這香膏賣三百個銀幣去賙濟窮人呢？」
JOHN|12|6|他說這話，並不是關心窮人，而是因為他是個賊，又管錢囊，常偷取錢囊中所存的。
JOHN|12|7|耶穌說：「由她吧！她這香膏本是為我的安葬之日留著的。
JOHN|12|8|因為常有窮人和你們在一起，但是你們不常有我。」
JOHN|12|9|有一大群 猶太 人知道耶穌在那裏，就來了，不但是為耶穌的緣故，也是要看耶穌使他從死人中復活的 拉撒路 。
JOHN|12|10|於是眾祭司長商議連 拉撒路 也要殺了，
JOHN|12|11|因為有許多 猶太 人為了 拉撒路 的緣故，開始背離他們，信了耶穌。
JOHN|12|12|第二天，有一大群上來過節的人聽見耶穌要來 耶路撒冷 ，
JOHN|12|13|就拿著棕樹枝出去迎接他，喊著： 「和散那 ， 以色列 的王！ 奉主名來的是應當稱頌的！」
JOHN|12|14|耶穌找到了一匹驢駒，就騎上，如經上所記：
JOHN|12|15|「 錫安 的兒女 啊，不要懼怕！ 看哪，你的王來了； 他騎在驢駒上。」
JOHN|12|16|門徒當初不明白這些事，等到耶穌得了榮耀後才想起這些話是指他寫的，並且人們果然對他做了這些事。
JOHN|12|17|當耶穌呼喚 拉撒路 ，使他從死人中復活出墳墓的時候，同耶穌在那裏的眾人就作見證。
JOHN|12|18|眾人因聽見耶穌行了這神蹟，就去迎接他。
JOHN|12|19|法利賽人彼此說：「你們看，你們一事無成，世人都隨著他去了。」
JOHN|12|20|那時，上來過節禮拜的人中，有幾個 希臘 人。
JOHN|12|21|他們來見 加利利 的 伯賽大 人 腓力 ，請求他說：「先生，我們想見耶穌。」
JOHN|12|22|腓力 去告訴 安得烈 ，然後 安得烈 同 腓力 去告訴耶穌。
JOHN|12|23|耶穌回答他們說：「人子得榮耀的時候到了。
JOHN|12|24|我實實在在地告訴你們，一粒麥子不落在地裏死了，仍舊是一粒；若是死了，就結出許多子粒來。
JOHN|12|25|愛惜自己性命的，就喪失性命；那恨惡自己在這世上的性命的，要保全性命到永生。
JOHN|12|26|若有人服事我，就當跟從我；我在哪裏，服事我的人也要在哪裏；若有人服事我，我父必尊重他。」
JOHN|12|27|「我現在心裏憂愁，我說甚麼才好呢？說『父啊，救我脫離這時候』嗎？但我正是為這時候來的。
JOHN|12|28|父啊，願你榮耀你的名！」於是有聲音從天上來，說：「我已經榮耀了我的名，還要再榮耀。」
JOHN|12|29|站在旁邊的眾人聽見，就說：「打雷了。」另有的說：「有天使對他說話。」
JOHN|12|30|耶穌回答說：「這聲音不是為我，而是為你們來的。
JOHN|12|31|現在正是這世界受審判的時候；現在這世界的統治者要被趕出去。
JOHN|12|32|我從地上被舉起來的時候，我要吸引萬人來歸我。」
JOHN|12|33|耶穌這話是指自己將要怎樣死說的。
JOHN|12|34|眾人就回答他：「我們聽見律法書上說，基督是永存的；你怎麼說，人子必須被舉起來呢？這人子是誰呢？」
JOHN|12|35|耶穌對他們說：「光在你們中間為時不多了，應該趁著有光的時候行走，免得黑暗臨到你們；那在黑暗裏行走的，不知道往何處去。
JOHN|12|36|你們趁著有光，要信從這光，使你們成為光明之子。」 耶穌說了這些話，就離開他們隱藏了。
JOHN|12|37|他雖然在他們面前行了許多神蹟，他們還是不信他。
JOHN|12|38|這是要應驗 以賽亞 先知所說的話： 「主啊，我們所傳的有誰信呢？ 主的膀臂向誰顯露呢？」
JOHN|12|39|他們所以不能信，因為 以賽亞 又說：
JOHN|12|40|「主使他們瞎了眼， 使他們硬了心， 免得他們眼睛看見， 他們心裏明白，回轉過來， 我會醫治他們。」
JOHN|12|41|以賽亞 因看見了他的榮耀，就說了關於他的這話。
JOHN|12|42|雖然如此，官長中卻有好些信他的，只因法利賽人的緣故不敢承認，恐怕被趕出會堂。
JOHN|12|43|這是因他們愛人給的尊榮過於愛上帝給的尊榮。
JOHN|12|44|耶穌喊著說：「信我的人不是信我，而是信差我來的那位。
JOHN|12|45|看見我的，就是看見差我來的那位。
JOHN|12|46|我就是來到世上的光，使凡信我的不住在黑暗裏。
JOHN|12|47|若有人聽見我的話而不遵守，我不審判他，因為我來不是要審判世人，而是要拯救世人。
JOHN|12|48|棄絕我、不領受我話的人自有審判他的；我所講的道在末日要審判他。
JOHN|12|49|因為我沒有憑著自己講，而是差我來的父已經給我命令，叫我說甚麼，講甚麼。
JOHN|12|50|我也知道他的命令就是永生。所以，我講的正是照著父所告訴我的，我就這麼講了。」
JOHN|13|1|逾越節以前，耶穌知道自己離世歸父的時候到了。他一向愛世間屬自己的人，就愛他們到底。
JOHN|13|2|晚餐的時候，魔鬼已把出賣耶穌的意思放在 加略 人 西門 的兒子 猶大 心裏。
JOHN|13|3|耶穌知道父已把萬有交在他手裏，且知道自己是從上帝出來的，又要回到上帝那裏去，
JOHN|13|4|就離席站起來，脫了衣服，拿一條手巾束腰，
JOHN|13|5|隨後把水倒在盆裏，開始洗門徒的腳，並用束腰的手巾擦乾。
JOHN|13|6|到了 西門．彼得 跟前， 彼得 對他說：「主啊，你洗我的腳嗎？」
JOHN|13|7|耶穌回答他說：「我所做的，你現在不知道，但以後會明白。」
JOHN|13|8|彼得 對他說：「你絕對不可以洗我的腳！」耶穌回答他：「我若不洗你，你就與我無份了。」
JOHN|13|9|西門．彼得 對他說：「主啊，不僅是我的腳，連手和頭也要洗！」
JOHN|13|10|耶穌對他說：「凡洗過澡的人不需要再洗，只要把腳一洗，全身就乾淨了。你們是乾淨的，然而不都是乾淨的。」
JOHN|13|11|耶穌已知道要出賣他的是誰，因此說「你們不都是乾淨的」。
JOHN|13|12|耶穌洗完了他們的腳，就穿上衣服，又坐下，對他們說：「我為你們所做的，你們明白嗎？
JOHN|13|13|你們稱呼我老師，稱呼我主，你們說的不錯，我本來就是。
JOHN|13|14|我是你們的主，你們的老師，尚且洗你們的腳，你們也應當彼此洗腳。
JOHN|13|15|我給你們作了榜樣，為要你們照著我為你們所做的去做。
JOHN|13|16|我實實在在地告訴你們，僕人不大於主人；奉差的人也不大於差他的人。
JOHN|13|17|你們既知道這些事，若是去實行就有福了。
JOHN|13|18|我不是指著你們眾人說的，我知道我所揀選的是誰；但是要應驗經上的話：『吃我飯的人 用腳踢我。』
JOHN|13|19|事情還沒有發生，我現在先告訴你們，讓你們到事情發生的時候好信我就是那位。
JOHN|13|20|我實實在在地告訴你們，接納我所差遣的就是接納我；接納我的就是接納差遣我的那位。」
JOHN|13|21|耶穌說了這些話，心裏憂愁，於是明確地說：「我實實在在地告訴你們，你們中間有一個人要出賣我。」
JOHN|13|22|門徒彼此相看，猜不出他說的是誰。
JOHN|13|23|門徒中有一個人，是耶穌所愛的，側身挨近耶穌的胸懷。
JOHN|13|24|西門．彼得 就對這個人示意，要問耶穌是指著誰說的。
JOHN|13|25|於是那人緊靠著耶穌的胸膛，問他：「主啊，是誰呢？」
JOHN|13|26|耶穌回答：「我蘸一點餅給誰，就是誰。」耶穌就蘸了一點餅，遞給 加略 人 西門 的兒子 猶大 。
JOHN|13|27|他接 了那餅以後，撒但就進入他的心。於是耶穌對他說：「你要做的，快做吧！」
JOHN|13|28|同席的人沒有一個知道耶穌為甚麼對他說這話。
JOHN|13|29|有人因 猶大 管錢囊，以為耶穌是對他說「你去買我們過節所需要的東西」，或是叫他拿些甚麼給窮人。
JOHN|13|30|猶大 受 了那點餅以後立刻出去。那時候是夜間了。
JOHN|13|31|猶大 出去後，耶穌說：「如今人子得了榮耀，上帝在人子身上也得了榮耀。
JOHN|13|32|如果上帝因人子得了榮耀 ，上帝也要因自己榮耀人子，並且要立刻榮耀他。
JOHN|13|33|孩子們！我與你們同在的時候不多了；你們會找我，但我所去的地方，你們不能去。這話我曾對 猶太 人說過，現在也照樣對你們說。
JOHN|13|34|我賜給你們一條新命令，乃是叫你們彼此相愛；我怎樣愛你們，你們也要怎樣彼此相愛。
JOHN|13|35|你們若彼此相愛，眾人因此就認出你們是我的門徒了。」
JOHN|13|36|西門．彼得 問耶穌：「主啊，你去哪裏？」耶穌回答：「我所去的地方，你現在不能跟我去，以後卻要跟我去。」
JOHN|13|37|彼得 對他說：「主啊，為甚麼我現在不能跟你去？我願意為你捨命。」
JOHN|13|38|耶穌回答：「你願意為我捨命嗎？我實實在在地告訴你，雞叫以前，你要三次不認我。」
JOHN|14|1|「你們心裏不要憂愁；你們信上帝，也當信我。
JOHN|14|2|在我父的家裏有許多住處；若是沒有，我就早已告訴你們了。我去原是為你們預備地去方。
JOHN|14|3|我若去為你們預備了地方，就必再來接你們到我那裏去，我在哪裏，叫你們也在哪裏。
JOHN|14|4|我往哪裏去，你們知道那條路。」
JOHN|14|5|多馬 對他說：「主啊，我們不知道你去哪裏，怎麼能知道那條路呢？」
JOHN|14|6|耶穌對他說：「我就是道路、真理、生命；若不藉著我，沒有人能到父那裏去。
JOHN|14|7|既然你們認識了我，也會認識我的父。從今以後，你們就認識他，並且已經看見他了。」
JOHN|14|8|腓力 對他說：「主啊，將父顯給我們看，我們就知足了。」
JOHN|14|9|耶穌對他說：「 腓力 ，我與你們在一起這麼久了，你還不認識我嗎？看見我的就是看見了父，你怎麼還說『將父顯給我們看』呢？
JOHN|14|10|我在父裏面，父在我裏面，你不信嗎？我對你們所說的話不是憑著自己說的，而是住在我裏面的父在做他的工作。
JOHN|14|11|你們要信我，我在父裏面，父在我裏面；即使不信，也要因我所做的工作信我。
JOHN|14|12|我實實在在地告訴你們，我所做的工作，信我的人也要做，並且要做得比這些更大，因為我到父那裏去。
JOHN|14|13|你們奉我的名無論求甚麼，我必成全，為了使父因兒子得榮耀。
JOHN|14|14|你們若奉我的名向我求甚麼，我必成全。」
JOHN|14|15|「你們若愛我，就會遵守我的命令。
JOHN|14|16|我要求父，父就賜給你們另外一位保惠師 ，使他永遠與你們同在。
JOHN|14|17|他就是真理的靈，是世人不能接受的。因為他們既看不見他，也不認識他；你們卻認識他，因他常與你們同在，也要在你們裏面。
JOHN|14|18|我不會撇下你們為孤兒，我必到你們這裏來。
JOHN|14|19|再過不久，世人不再看見我，你們卻會看見我，因為我活著，你們也要活著。
JOHN|14|20|到那日，你們就會知道我在父裏面，你們在我裏面，我也在你們裏面。
JOHN|14|21|有了我的命令而又遵守的人，就是愛我的；愛我的人，我父要愛他，我也要愛他，並且要親自向他顯現。」
JOHN|14|22|猶大 （不是 加略 人 猶大 ）問耶穌：「主啊，為甚麼親自向我們顯現，而不向世人顯現呢？」
JOHN|14|23|耶穌回答他說：「凡愛我的人就會遵守我的道，我父也會愛他，並且我們要到他那裏去，與他同住。
JOHN|14|24|不愛我的人就不遵守我的道。你們所聽見的道不是我的，而是差我來之父的。
JOHN|14|25|「我還與你們在一起的時候，已對你們說了這些事。
JOHN|14|26|但保惠師，就是父因我的名所要差來的聖靈，他要把一切的事教導你們，並且要使你們想起我對你們所說的一切話。
JOHN|14|27|我留下平安給你們，我把我的平安賜給你們。我所賜給你們的，不像世人所賜的。你們心裏不要憂愁，也不要膽怯。
JOHN|14|28|你們聽見我對你們說過，我去了還要回到你們這裏來。你們若愛我，就會因我到父那裏去而喜樂，因為父比我大。
JOHN|14|29|現在事情還沒有發生，我預先告訴你們，使你們在事情發生的時候會信。
JOHN|14|30|我不再和你們多說了，因為這世界的統治者將到，他在我身上一無所能。
JOHN|14|31|我這麼做是照著父命令我的，為了讓世人知道我愛父。起來，我們走吧！」
JOHN|15|1|「我就是真葡萄樹，我父是栽培的人。
JOHN|15|2|凡屬我不結果子的枝子，他就剪掉；凡結果子的，他就修剪乾淨，使枝子結果子更多。
JOHN|15|3|現在你們因我講給你們的道已經潔淨了。
JOHN|15|4|你們要常在我裏面，我也常在你們裏面。枝子若不常在葡萄樹上，自己就不能結果子；你們若不常在我裏面，也是這樣。
JOHN|15|5|我就是葡萄樹，你們是枝子。常在我裏面的，我也常在他裏面，這人就多結果子，因為離了我，你們就不能做甚麼。
JOHN|15|6|人若不常在我裏面，就像枝子被丟在外面，枯乾了，人撿起來，扔進火裏燒了。
JOHN|15|7|你們若常在我裏面，我的話也常在你們裏面，凡你們想要的，祈求，就給你們成全。
JOHN|15|8|你們多結果子，我父就因此得榮耀，你們也就是 我的門徒了。
JOHN|15|9|我愛你們，正如父愛我一樣；你們要常在我的愛裏。
JOHN|15|10|你們若遵守我的命令，就會常在我的愛裏，正如我遵守了我父的命令，常在他的愛裏。
JOHN|15|11|「我已對你們說了這些事，是要讓我的喜樂存在你們心裏，並讓你們的喜樂得以滿足。
JOHN|15|12|你們要彼此相愛，像我愛你們一樣，這是我的命令。
JOHN|15|13|人為朋友捨命，人的愛心沒有比這個更大的了。
JOHN|15|14|你們若遵行我所命令的，就是我的朋友。
JOHN|15|15|以後我不再稱你們為僕人，因為僕人不知道主人所做的事；但我稱你們為朋友，因為我從我父所聽見的一切都已經讓你們知道了。
JOHN|15|16|不是你們揀選了我，而是我揀選了你們，並且派你們去結果子，讓你們的果子得以長存，好使你們奉我的名，無論向父求甚麼，他會賜給你們。
JOHN|15|17|我這樣命令你們，是要你們彼此相愛。」
JOHN|15|18|「世人若恨你們，你們要知道，他們在恨你們以前已經恨我了。
JOHN|15|19|你們若屬世界，世界會愛屬自己的；只因你們不屬世界，而是我從世界中揀選了你們，所以世界就恨你們。
JOHN|15|20|你們要記得我對你們說過的話：『僕人不大於主人。』他們若迫害了我，也會迫害你們，他們若遵守了我的話，也會遵守你們的話。
JOHN|15|21|但他們要因我的名向你們做這一切的事，因為他們不認識差我來的那位。
JOHN|15|22|我若沒有來教導他們，他們就沒有罪；但如今他們的罪無可推諉了。
JOHN|15|23|恨我的也恨我的父。
JOHN|15|24|我若沒有在他們中間做過別人未曾做的事，他們就沒有罪；但如今連我與我的父，他們也看見了，也恨惡了。
JOHN|15|25|這是要應驗他們律法上所寫的話：『他們無故地恨我。』
JOHN|15|26|「但我要從父那裏差保惠師來，就是從父出來的那真理的靈，他來的時候要為我作見證。
JOHN|15|27|你們也要作見證，因為你們從起初就與我同在。」
JOHN|16|1|「我對你們說了這些事，是要使你們不至於跌倒。
JOHN|16|2|人要把你們趕出會堂，而且時候將到，凡殺你們的還以為是在事奉上帝。
JOHN|16|3|他們這樣做，是因為沒有認識父，也沒有認識我。
JOHN|16|4|我對你們說了這些事，是要在他們做這些事的時候，你們會想起我對你們說過的話。」 「我起先沒有對你們說這些事，因為我一直與你們同在。
JOHN|16|5|現在我要到差我來的父那裏去，你們中間卻沒有人問我『你去哪裏？』
JOHN|16|6|只因我對你們說了這些事，你們就滿心憂愁。
JOHN|16|7|然而，我把真情告訴你們，我去對你們是有益的。我若不去，保惠師就不會到你們這裏來；我若去，就差他到你們這裏來。
JOHN|16|8|他來的時候，要為罪、為義，為審判，指證世人；
JOHN|16|9|為罪，是因他們不信我；
JOHN|16|10|為義，是因我到父那裏去，你們將不再見到我；
JOHN|16|11|為審判，是因這世界的統治者已受了審判。
JOHN|16|12|「我還有好些事要告訴你們，但你們現在擔當不了 。
JOHN|16|13|但真理的靈來的時候，他要引導你們進入一切真理。因為他不是憑著自己說的，而是把他所聽見的都說出來，並且要把將要來的事向你們傳達。
JOHN|16|14|他要榮耀我，因為他要把從我領受的向你們傳達。
JOHN|16|15|凡父所有的都是我的，所以我說，他要把從我領受的向你們傳達。」
JOHN|16|16|「不久，你們將不再見到我；再過不久，你們還要見到我。」
JOHN|16|17|有幾個門徒彼此說：「他對我們說『不久，你們將不再見到我；再過不久，你們還要見到我』；又說『因我到父那裏去』。這是甚麼意思呢？」
JOHN|16|18|於是門徒說：「他說 『不久』到底是甚麼意思呢？我們不明白他說甚麼。」
JOHN|16|19|耶穌看出他們要問他，就對他們說：「我說『不久，你們將不再見到我；再過不久，你們還要見到我』，你們為這話彼此詢問嗎？
JOHN|16|20|我實實在在地告訴你們，你們將要痛哭，哀號，世人反要歡喜。你們將要憂愁，然而你們的憂愁要變成喜樂。
JOHN|16|21|婦人生產的時候會憂愁，因為她的時候到了；但孩子一生出來，就不再記得那痛苦了，因為歡喜有一個人生在世上了。
JOHN|16|22|你們現在也是憂愁，但我要再見到你們，你們的心就會有喜樂了；這喜樂沒有人能奪去。
JOHN|16|23|到那日，你們甚麼也不會問我了。我實實在在地告訴你們，你們奉我的名無論向父求甚麼，他會賜給你們 。
JOHN|16|24|直到現在，你們沒有奉我的名求甚麼，如今你們求就必得著，使你們的喜樂得以滿足。」
JOHN|16|25|「這些事，我是用比方對你們說的；時候將到，我不再用比方對你們說，而是要把父的事明白地告訴你們。
JOHN|16|26|到那日，你們要奉我的名祈求；我並不對你們說，我要為你們向父祈求。
JOHN|16|27|父自己愛你們，因為你們已經愛我，又信我是從上帝 而來的。
JOHN|16|28|我從父而來，到了世界 ，又離開世界，到父那裏去。」
JOHN|16|29|門徒說：「你看，如今你是明說，不用比方了。
JOHN|16|30|現在我們曉得你凡事都知道，也不需要有人問你；從此我們信你是從上帝而來的。」
JOHN|16|31|耶穌回答他們：「現在你們信了嗎？
JOHN|16|32|看哪，時候將到，其實已經到了，你們要分散，各歸自己的地方，留下我獨自一人；然而我不是獨自一人，因為有父與我同在。
JOHN|16|33|我對你們說了這些事，是要使你們在我裏面有平安。在世上你們有苦難，但你們要有勇氣 ，我已經勝過世界。」
JOHN|17|1|耶穌說了這些話，就舉目望天，說：「父啊，時候到了，願你榮耀你的兒子，使兒子也榮耀你；
JOHN|17|2|因為你曾賜給他權柄掌管凡血肉之軀的，使他把永生賜給你所賜給他的人。
JOHN|17|3|認識你—獨一的真神，並且認識你所差來的耶穌基督，這就是永生。
JOHN|17|4|我在地上已經榮耀你，你交給我做的工作，我已完成了。
JOHN|17|5|父啊，現在求你使我在你面前得榮耀，就是在未有世界以前，我同你享有的榮耀。
JOHN|17|6|「你從世上賜給我的人，我已把你的名顯明給他們。他們本是你的，你把他們賜給我，他們也遵守了你的道。
JOHN|17|7|現在他們知道，你所賜給我的一切都是從你那裏來的；
JOHN|17|8|因為你所賜給我的話，我已經賜給他們，他們也領受了，又確實知道，我是從你出來的，並且信你差了我來。
JOHN|17|9|我為他們祈求，不為世人祈求，卻為你所賜給我的人祈求，因他們本是你的。
JOHN|17|10|凡是我的都是你的，你的也是我的，並且我因他們得了榮耀。
JOHN|17|11|我到你那裏去；我不再留在世上，他們卻在世上。聖父啊，求你因你的名，就是你所賜給我的名，保守他們，使他們像我們一樣合而為一。
JOHN|17|12|我與他們同在的時候，我奉你的名，就是你所賜給我的名，保守了他們，我也護衛了他們；其中除了那滅亡之子，沒有一個滅亡的，好使經上的話得以應驗。
JOHN|17|13|現在我到你那裏去，我在世上說這些話，是要他們心裏充滿了我的喜樂。
JOHN|17|14|我已把你的道賜給他們；世界恨他們，因為他們不屬世界，正如我不屬世界一樣。
JOHN|17|15|我不求你把他們從世上接走，只求你保全他們，使他們脫離那惡者。
JOHN|17|16|他們不屬世界，正如我不屬世界一樣。
JOHN|17|17|求你用真理使他們成聖；你的道就是真理。
JOHN|17|18|你怎樣差我到世上，我也照樣差他們到世上。
JOHN|17|19|我為他們的緣故使自己分別為聖，為要使他們也因真理成聖。
JOHN|17|20|「我不但為這些人祈求，也為那些藉著他們的話信我的人祈求，
JOHN|17|21|使他們都合而為一。正如父你在我裏面，我在你裏面，使他們也在我們裏面，好讓世人信是你差我來的。
JOHN|17|22|你所賜給我的榮耀，我已賜給他們，使他們合而為一，像我們合而為一。
JOHN|17|23|我在他們裏面，你在我裏面，使他們完完全全合而為一，讓世人知道是你差我來的，也知道你愛他們，如同愛我一樣。
JOHN|17|24|父啊，我在哪裏，願你所賜給我的人也同我在哪裏，使他們看見你所賜給我的榮耀，因為創世以前，你已經愛我了。
JOHN|17|25|公義的父啊，世人未曾認識你，我卻認識你，這些人也知道是你差我來的。
JOHN|17|26|我已讓他們認識你的名，還要讓他們認識，好讓你愛我的愛在他們裏面，我也在他們裏面。」
JOHN|18|1|耶穌說了這些話，就同門徒出去，過了 汲淪溪 。在那裏有一個園子，他和門徒進去了。
JOHN|18|2|出賣耶穌的 猶大 也知道那地方，因為耶穌和門徒屢次在那裏聚集。
JOHN|18|3|猶大 領了一隊兵，以及祭司長和法利賽人的聖殿警衛，拿著燈籠、火把和兵器來到園裏。
JOHN|18|4|耶穌知道將要臨到自己的一切事，就出來對他們說：「你們找誰？」
JOHN|18|5|他們回答他：「 拿撒勒 人耶穌。」耶穌對他們說：「我就是。」出賣他的 猶大 也同他們站在一起。
JOHN|18|6|耶穌一對他們說「我就是」，他們就退後，倒在地上。
JOHN|18|7|他又問他們：「你們找誰？」他們說：「 拿撒勒 人耶穌。」
JOHN|18|8|耶穌回答：「我已經告訴你們，我就是。你們若找的是我，就讓這些人走吧。」
JOHN|18|9|這要應驗耶穌說過的話：「你所賜給我的人，我一個也不失落。」
JOHN|18|10|西門．彼得 帶著一把刀，就拔出來，把大祭司的僕人砍了一刀，削掉了他的右耳，那僕人名叫 馬勒古 。
JOHN|18|11|於是耶穌對 彼得 說：「收刀入鞘吧！我父給我的杯，我豈可不喝呢？」
JOHN|18|12|那隊兵、千夫長和 猶太 人的警衛拿住耶穌，把他捆綁了，
JOHN|18|13|先帶到 亞那 面前，因為他是那年的大祭司 該亞法 的岳父。
JOHN|18|14|這 該亞法 就是從前向 猶太 人忠告說「一個人替百姓死是有利的」那個人。
JOHN|18|15|西門．彼得 跟著耶穌，另一個門徒也跟著；那門徒是大祭司所認識的，他就同耶穌進了大祭司的院子。
JOHN|18|16|彼得 卻站在門外。大祭司所認識的那個門徒出來，對看門的使女說了一聲，就領 彼得 進去。
JOHN|18|17|那看門的使女對 彼得 說：「你不也是這人的門徒嗎？」他說：「我不是。」
JOHN|18|18|僕人和警衛因為天冷生了炭火，站在那裏取暖； 彼得 也同他們站著取暖。
JOHN|18|19|於是，大祭司盤問耶穌有關他的門徒和他教導的事。
JOHN|18|20|耶穌回答他：「我一向都是公開地對世人講話，我常在會堂和聖殿裏，就是 猶太 人聚集的地方教導人，我私下並沒有講甚麼。
JOHN|18|21|你為甚麼問我呢？去問那些聽過我講話的人，我所說的，他們都知道。」
JOHN|18|22|耶穌說了這些話，旁邊站著的一個警衛打了他一耳光，說：「你這樣回答大祭司嗎？」
JOHN|18|23|耶穌回答他：「假如我說的不對，你指證不對的地方；假如我說的對，你為甚麼打我呢？」
JOHN|18|24|於是 亞那 把耶穌綁著押解到大祭司 該亞法 那裏。
JOHN|18|25|西門．彼得 正站著取暖，有人對他說：「你不也是他的門徒嗎？」 彼得 不承認，說：「我不是。」
JOHN|18|26|大祭司的一個僕人，是被 彼得 削掉耳朵那人的親屬，說：「我不是看見你同他在園子裏嗎？」
JOHN|18|27|彼得 又不承認，立刻雞就叫了。
JOHN|18|28|他們把耶穌從 該亞法 那裏押解到總督府。那時是清早。他們自己卻不進總督府，恐怕染了污穢，不能吃逾越節的宴席。
JOHN|18|29|於是 彼拉多 出來，到他們那裏，說：「你們告這人是為甚麼事呢？」
JOHN|18|30|他們回答他說：「這人若不作惡，我們就不會把他交給你了。」
JOHN|18|31|彼拉多 對他們說：「你們自己帶他去，按著你們的律法問他吧！」 猶太 人說：「我們沒有殺人的權柄。」
JOHN|18|32|這是要應驗耶穌所說，指自己將要怎樣死的話。
JOHN|18|33|於是 彼拉多 又進了總督府，叫耶穌來，對他說：「你是 猶太 人的王嗎？」
JOHN|18|34|耶穌回答：「這話是你說的，還是別人論到我時對你說的呢？」
JOHN|18|35|彼拉多 回答：「難道我是 猶太 人嗎？你的同胞和祭司長把你交給我。你做了甚麼事呢？」
JOHN|18|36|耶穌回答：「我的國不屬於這世界；我的國若屬於這世界，我的部下就會為我戰鬥，使我不至於被交給 猶太 人。只是我的國不屬於這世界。」
JOHN|18|37|於是 彼拉多 對他說：「那麼，你是王了？」耶穌回答：「是你說我是王。我為此而生，也為此來到世界，為了給真理作見證。凡屬真理的人都聽我的話。」
JOHN|18|38|彼拉多 對他說：「真理是甚麼呢？」 說了這話， 彼拉多 又出來到 猶太 人那裏，對他們說：「我查不出他有甚麼罪狀。
JOHN|18|39|但你們有個規矩，在逾越節要我給你們釋放一個人，你們要我給你們釋放這 猶太 人的王嗎？」
JOHN|18|40|他們又再喊著說：「不要這人！要 巴拉巴 ！」這 巴拉巴 是個強盜。
JOHN|19|1|於是， 彼拉多 命令把耶穌帶去鞭打了。
JOHN|19|2|士兵用荊棘編了冠冕，戴在他頭上，給他穿上紫袍，
JOHN|19|3|又走到他面前，說：「萬歲， 猶太 人的王！」他們就打他耳光。
JOHN|19|4|彼拉多 又出來對眾人說：「看，我帶他出來見你們，讓你們知道我查不出他有甚麼罪狀。」
JOHN|19|5|耶穌出來，戴著荊棘冠冕，穿著紫袍。 彼拉多 對他們說：「看哪，這個人！」
JOHN|19|6|祭司長和聖殿警衛看見他，就喊著說：「釘十字架！釘十字架！」 彼拉多 對他們說：「你們自己把他帶去釘十字架吧！我查不出他有甚麼罪狀。」
JOHN|19|7|猶太 人回答他：「我們有律法，按照律法，他是該死的，因為他自以為是上帝的兒子。」
JOHN|19|8|彼拉多 聽見這話，越發害怕，
JOHN|19|9|又進了總督府，對耶穌說：「你是哪裏來的？」耶穌卻不回答。
JOHN|19|10|於是 彼拉多 對他說：「你不對我說話嗎？難道你不知道我有權柄釋放你，也有權柄把你釘十字架嗎？」
JOHN|19|11|耶穌回答他：「若不是從上頭賜給你的，你就毫無權柄辦我，所以，把我交給你的那人罪更重了。」
JOHN|19|12|從此， 彼拉多 想要釋放耶穌，無奈 猶太 人喊著說：「你若釋放這個人，你就不是凱撒的忠臣 。凡自立為王的就是背叛凱撒。」
JOHN|19|13|彼拉多 聽見這些話，就帶耶穌出來，到了一個地方，叫「鋪華石處」， 希伯來 話叫 厄巴大 ，就在那裏坐堂。
JOHN|19|14|那日是逾越節的預備日，約在正午。 彼拉多 對 猶太 人說：「看哪，你們的王！」
JOHN|19|15|他們就喊著：「除掉他！除掉他！把他釘十字架！」 彼拉多 對他們說：「要我把你們的王釘十字架嗎？」祭司長回答：「除了凱撒，我們沒有王。」
JOHN|19|16|於是 彼拉多 把耶穌交給他們去釘十字架。 他們就把耶穌帶了去。
JOHN|19|17|耶穌背著自己的十字架出來，到了一個地方，名叫「髑髏地」， 希伯來 話叫 各各他 。
JOHN|19|18|他們就在那裏把他釘在十字架上，還有兩個人和他一同被釘，一邊一個，耶穌在中間。
JOHN|19|19|彼拉多 又寫了一個牌子，釘在十字架上，寫的是：「 猶太 人的王， 拿撒勒 人耶穌。」
JOHN|19|20|有許多 猶太 人念這牌子，因為耶穌被釘十字架的地方靠近城，而且牌子是用 希伯來 、 羅馬 、 希臘 三種文字寫的。
JOHN|19|21|猶太 人的祭司長就對 彼拉多 說：「不要寫『 猶太 人的王』，要寫『那人說：我是 猶太 人的王』。」
JOHN|19|22|彼拉多 回答：「我寫了就寫了。」
JOHN|19|23|士兵把耶穌釘在十字架上以後，把他的衣服拿來分為四份，每人一份。他們又拿他的內衣，這件內衣沒有縫，是上下一片織成的。
JOHN|19|24|他們就彼此說：「我們不要撕開，我們抽籤，看是誰的。」這要應驗經上的話說： 「他們分了我的外衣， 為我的內衣抽籤。」 士兵果然做了這些事。
JOHN|19|25|站在耶穌十字架旁邊的，有他的母親、姨母、 革羅罷 的妻子 馬利亞 ，和 抹大拉 的 馬利亞 。
JOHN|19|26|耶穌見母親和他所愛的那門徒站在旁邊，就對母親說：「母親 ，看，你的兒子！」
JOHN|19|27|又對那門徒說：「看，你的母親！」從那刻起，那門徒就接她到自己家裏去了。
JOHN|19|28|這事以後，耶穌知道各樣的事已經成了，為使經上的話應驗，就說：「我渴了。」
JOHN|19|29|有一個盛滿了醋的罐子放在那裏，他們就拿海綿蘸滿了醋，綁在牛膝草上，送到他嘴邊。
JOHN|19|30|耶穌嘗了那醋，說：「成了！」就低下頭，斷了氣 。
JOHN|19|31|因為這日是預備日，又因為那安息日是個大日子， 猶太 人就來求 彼拉多 叫人打斷他們的腿，把他們搬走，免得屍首在安息日留在十字架上。
JOHN|19|32|於是士兵來，把第一個人的腿，和與耶穌同釘的另一個人的腿，都打斷了。
JOHN|19|33|當他們來到耶穌那裏，見他已經死了，就沒有打斷他的腿。
JOHN|19|34|然而有一個士兵拿槍扎他的肋旁，立刻有血和水流出來。
JOHN|19|35|看見這事的人作了見證—他的見證是真的，他知道自己所說的是真的—好讓你們也信。
JOHN|19|36|這些事發生，為要應驗經上的話：「他的骨頭一根也不可折斷。」
JOHN|19|37|另有經文也說：「他們要仰望自己所扎的人。」
JOHN|19|38|這些事以後， 亞利馬太 的 約瑟 來求 彼拉多 ，要把耶穌的身體領去。他是耶穌的門徒，只因怕 猶太 人，就暗地裏作門徒。 彼拉多 准許了，他就把耶穌的身體領走。
JOHN|19|39|尼哥德慕 也來了，就是先前夜裏去見耶穌的那位，他帶著約一百斤的沒藥和沉香。
JOHN|19|40|他們照 猶太 人喪葬的規矩，用細麻布加上香料，把耶穌的身體裹好了。
JOHN|19|41|在耶穌釘十字架的地方有一個園子，園子裏有一座新墓穴，是從來沒有葬過人的。
JOHN|19|42|因為那天是 猶太 人的預備日，而那墳墓又在附近，他們就把耶穌安放在那裏。
JOHN|20|1|七日的第一日清早，天還黑的時候， 抹大拉 的 馬利亞 來到墳墓，看見石頭已從墳墓挪開了，
JOHN|20|2|就跑來見 西門．彼得 和耶穌所愛的那個門徒，對他們說：「有人從墳墓裏把主移走了，我們不知道他們把他放在哪裏。」
JOHN|20|3|彼得 和那門徒就出來，往墳墓去。
JOHN|20|4|兩個人同跑，那門徒比 彼得 跑得快，先到了墳墓，
JOHN|20|5|低頭往裏看，看見細麻布還放在那裏，只是沒有進去。
JOHN|20|6|西門．彼得 隨後也到了，進了墳墓，看見細麻布放在那裏，
JOHN|20|7|又看見耶穌的裹頭巾沒有和細麻布放在一起，是另在一處捲著。
JOHN|20|8|然後先到墳墓的那門徒也進去，他看見就信了。
JOHN|20|9|他們還不明白聖經所說耶穌必須從死人中復活的意思。
JOHN|20|10|於是兩個門徒回自己的住處去了。
JOHN|20|11|馬利亞 卻站在墳墓外面哭。她哭的時候，低頭往墳墓裏看，
JOHN|20|12|看見兩個天使穿著白衣，在安放耶穌身體的地方坐著，一個在頭，一個在腳。
JOHN|20|13|天使對她說：「婦人，你為甚麼哭？」她對他們說：「因為有人把我主移走了，我不知道他們把他放在哪裏。」
JOHN|20|14|說了這些話，她轉過身來，看見耶穌站在那裏，卻不知道他是耶穌。
JOHN|20|15|耶穌問她：「婦人，你為甚麼哭？你找誰？」 馬利亞 以為他是看園子的，就對他說：「先生，若是你把他移了去，請告訴我，你把他放在哪裏，我去把他移回來。」
JOHN|20|16|耶穌對她說：「 馬利亞 。」 馬利亞 轉過身來，用 希伯來 話對他說：「拉波尼！」（「拉波尼」就是老師的意思。）
JOHN|20|17|耶穌對她說：「不要拉住我，因為我還沒有升上去見我的父。你到我弟兄那裏去告訴他們，我要升上去見我的父，也是你們的父，見我的上帝，也是你們的上帝。」
JOHN|20|18|抹大拉 的 馬利亞 就向門徒報信：「我已經看見了主。」她又把主對她說的話告訴他們。
JOHN|20|19|那日（就是七日的第一日）晚上，門徒因怕 猶太 人，所在的地方門都關了。耶穌來，站在當中，對他們說：「願你們平安！」
JOHN|20|20|說了這話，他把手和肋旁給他們看。門徒一看見主就喜樂了。
JOHN|20|21|於是耶穌又對他們說：「願你們平安！父怎樣差遣了我，我也照樣差遣你們。」
JOHN|20|22|說了這話，他向他們吹一口氣，說：「領受聖靈吧！
JOHN|20|23|你們赦免誰的罪，誰的罪就得赦免；你們不赦免誰的罪，誰的罪就不得赦免。」
JOHN|20|24|那十二使徒中，有個叫 低土馬 的 多馬 ，耶穌來的時候，他沒有和他們在一起。
JOHN|20|25|其他的門徒就對他說：「我們已經看見主了。」 多馬 卻對他們說：「除非我看見他手上的釘痕，用我的指頭探入那釘痕，用我的手探入他的肋旁，我絕不信。」
JOHN|20|26|過了八日，門徒又在屋裏， 多馬 也和他們在一起。門都關了，耶穌來，站在當中，說：「願你們平安！」
JOHN|20|27|然後他對 多馬 說：「把你的指頭伸到這裏來，看看我的手；把你的手伸過來，探入我的肋旁。不要疑惑，總要信！」
JOHN|20|28|多馬 回答，對他說：「我的主！我的上帝！」
JOHN|20|29|耶穌對他說：「你因為看見了我才信嗎？那沒有看見卻信的有福了。」
JOHN|20|30|耶穌在他門徒面前另外行了許多神蹟，沒有記錄在這書上。
JOHN|20|31|但記載這些事是要使你們信 耶穌是基督，是上帝的兒子，並且使你們信他，好因著他的名得生命。
JOHN|21|1|這些事以後，耶穌在 提比哩亞 海邊又向門徒顯現。他怎樣顯現記在下面。
JOHN|21|2|西門．彼得 、叫 低土馬 的 多馬 、 加利利 的 迦拿 人 拿但業 、 西庇太 的兩個兒子，和另外兩個門徒，都在一起。
JOHN|21|3|西門．彼得 對他們說：「我打魚去。」他們對他說：「我們也和你一起去。」他們就出去，上了船；那一夜並沒有打著甚麼。
JOHN|21|4|天剛亮的時候，耶穌站在岸上，門徒卻不知道他是耶穌。
JOHN|21|5|耶穌就對他們說：「孩子們！你們有吃的沒有？」他們回答他：「沒有。」
JOHN|21|6|耶穌對他們說：「你們把網撒在船的右邊，就會得到。」於是他們撒下網去，竟拉不上來了，因為魚很多。
JOHN|21|7|耶穌所愛的那門徒對 彼得 說：「是主！」那時 西門．彼得 赤著身子，一聽見是主，就束上外衣，跳進海裏。
JOHN|21|8|其餘的門徒因離岸不遠，約有二百肘，就坐著小船把那網魚拉過來。
JOHN|21|9|他們上了岸，看見那裏有炭火，上面有魚和餅。
JOHN|21|10|耶穌對他們說：「把剛才打的魚拿幾條來。」
JOHN|21|11|西門．彼得 就上船，把網拉到岸上，網裏滿了大魚，共一百五十三條；雖然魚這樣多，網卻沒有破。
JOHN|21|12|耶穌對他們說：「你們來吃早飯。」門徒中沒有一個敢問他：「你是誰？」因為他們知道他是主。
JOHN|21|13|耶穌走過來，拿餅給他們，也照樣拿魚給他們。
JOHN|21|14|耶穌從死人中復活後向門徒顯現，這是第三次。
JOHN|21|15|他們吃完了早飯，耶穌對 西門．彼得 說：「 約翰 的兒子 西門 ，你愛我比這些更深嗎？」 彼得 對他說：「主啊，是的，你知道我愛你。」耶穌對他說：「你餵養我的小羊。」
JOHN|21|16|耶穌第二次又對他說：「 約翰 的兒子 西門 ，你愛我嗎？」 彼得 對他說：「主啊，是的，你知道我愛你。」耶穌說：「你牧養我的羊。」
JOHN|21|17|耶穌第三次對他說：「 約翰 的兒子 西門 ，你愛我嗎？」 彼得 因為耶穌第三次對他說「你愛我嗎」，就憂愁，對耶穌說：「主啊，你無所不知，你知道我愛你。」耶穌說：「你餵養我的羊。
JOHN|21|18|我實實在在地告訴你，你年輕的時候，自己束上帶子，隨意往來；但年老的時候，你要伸出手來，別人要把你束上，帶你到不願意去的地方。」
JOHN|21|19|耶穌說這話，是指 彼得 會怎樣死來榮耀上帝。說了這話，耶穌對他說：「你跟從我吧！」
JOHN|21|20|彼得 轉過身來，看見耶穌所愛的那門徒跟著，就是在晚餐時靠著耶穌胸膛說「主啊，出賣你的是誰」的那門徒。
JOHN|21|21|彼得 看見他，就問耶穌：「主啊，這個人怎樣呢？」
JOHN|21|22|耶穌對他說：「假如我要他等到我來的時候還在，跟你有甚麼關係呢？你跟從我吧！」
JOHN|21|23|於是這話在弟兄中間流傳，說那門徒不死。其實，耶穌不是說他不死，而是對 彼得 說：「假如我要他等到我來的時候還在，跟你有甚麼關係呢？ 」
JOHN|21|24|這門徒就是為這些事作見證、並且記載這些事的，我們知道他的見證是真的。
JOHN|21|25|耶穌所行的事還有許多，若是一一都寫出來，我想，就是全世界也容不下所要寫的書。
ACTS|1|1|提阿非羅 啊，我在第一本書中已論到耶穌從開頭所做和所教導的一切事，
ACTS|1|2|直到他藉著聖靈吩咐所揀選的使徒後，被接上升的日子為止。
ACTS|1|3|他受害以後，用許多確據向使徒顯明自己是活著的，在四十天之中向他們顯現，並講說上帝國的事。
ACTS|1|4|耶穌和他們聚集的時候，囑咐他們說：「不要離開 耶路撒冷 ，但要等候父的應許，就是你們聽見我說過的。
ACTS|1|5|約翰 是用水施洗，但過了不多幾天，你們要在聖靈裏受洗。」
ACTS|1|6|他們聚集的時候，問耶穌：「主啊，你就要在這時候復興 以色列 國嗎？」
ACTS|1|7|耶穌對他們說：「父憑著自己的權柄所定的時候和日期，不是你們可以知道的。
ACTS|1|8|但聖靈降臨在你們身上，你們就必得著能力，並要在 耶路撒冷 、 猶太 全地和 撒瑪利亞 ，直到地極，作我的見證。」
ACTS|1|9|說了這些話，他們正看的時候，他被接上升，有一朵雲彩從他們眼前把他接去。
ACTS|1|10|他升上去的時候，他們定睛望天，看哪，有兩個人身穿白衣站在他們旁邊，
ACTS|1|11|說：「 加利利 人哪，你們為甚麼站著望天呢？這離開你們被接升天的耶穌，你們見他怎樣升上天去，他也要怎樣來臨。」
ACTS|1|12|有一座山，名叫 橄欖山 ，離 耶路撒冷 不遠，有安息日可行走的路程 。那時，門徒從那裏回 耶路撒冷 去，
ACTS|1|13|他們一進城，就上了所住的樓房；在那裏有 彼得 、 約翰 、 雅各 、 安得烈 、 腓力 、 多馬 、 巴多羅買 、 馬太 、 亞勒腓 的兒子 雅各 、激進黨的 西門 ，和 雅各 的兒子 猶大 。
ACTS|1|14|這些人和幾個婦人，包括耶穌的母親 馬利亞 ，和耶穌的兄弟，都同心合意地恆切禱告。
ACTS|1|15|那時，有許多人聚會，約有一百二十名， 彼得 在弟兄中間站起來，說：
ACTS|1|16|「諸位弟兄，聖經的話必須應驗。聖經中，聖靈曾藉 大衛 的口預先說到那領人來拿耶穌的 猶大 ；
ACTS|1|17|他本來算是我們中的一個，並且得了這一份使徒的職任。
ACTS|1|18|這人用他不義的代價買了一塊田，以後身子仆倒，肚腹崩裂，腸子都流出來。
ACTS|1|19|住在 耶路撒冷 的人都知道這事，所以按著他們當地的話把那塊田叫 亞革大馬 ，就是「血田」的意思。
ACTS|1|20|因為《詩篇》上寫著： 「願他的住處變為廢墟， 無人在內居住。」 又說： 「願別人得他的職分。」
ACTS|1|21|所以，主耶穌在我們中間出入的整段時間，就是從 約翰 施洗起，直到主離開我們被接上升的日子為止，必須從那常與我們一起的人中，立一位與我們同作耶穌復活的見證。」
ACTS|1|22|
ACTS|1|23|於是他們推舉兩個人，就是那叫 巴撒巴 ，又稱為 猶士都 的 約瑟 ，和 馬提亞 。
ACTS|1|24|眾人禱告說：「主啊，你知道萬人的心，求你從這兩個人中指明你所揀選的是哪一位，
ACTS|1|25|去得這使徒的職任；這職位 猶大 已經丟棄，往自己的地方去了。」
ACTS|1|26|於是眾人為他們搖籤，搖出 馬提亞 來；他就和十一個使徒同列。
ACTS|2|1|五旬節那日到了，他們全都聚集在一起。
ACTS|2|2|忽然，有響聲從天上下來，好像一陣大風吹過，充滿了他們所坐的整座屋子；
ACTS|2|3|又有舌頭如火焰向他們顯現，分開落在他們每個人身上。
ACTS|2|4|他們都被聖靈充滿，就按著聖靈所賜的口才說起別國的話來。
ACTS|2|5|那時，有從天下各國來的虔誠的 猶太 人，住在 耶路撒冷 。
ACTS|2|6|這聲音一響，許多人都來聚集，各人因為聽見門徒用他們各自的鄉談說話，就甚納悶，
ACTS|2|7|都詫異驚奇說：「看哪，這些說話的不都是 加利利 人嗎？
ACTS|2|8|我們每個人怎麼聽見他們說我們生來所用的鄉談呢？
ACTS|2|9|我們 帕提亞 人、 瑪代 人、 以攔 人，和住在 美索不達米亞 、 猶太 、 加帕多家 、 本都 、 亞細亞 、
ACTS|2|10|弗呂家 、 旁非利亞 、 埃及 的人，並靠近 古利奈 的 利比亞 一帶地方的人，僑居的 羅馬 人，
ACTS|2|11|包括 猶太 人和皈依 猶太 教的人， 克里特 人和 阿拉伯 人，都聽見他們用我們的鄉談講論上帝的大作為。」
ACTS|2|12|眾人就都驚奇困惑，彼此說：「這是甚麼意思呢？」
ACTS|2|13|還有人譏誚，說：「他們是灌滿了新酒吧！」
ACTS|2|14|彼得 和十一個使徒站起來，他就高聲向眾人說：「 猶太 人和所有住在 耶路撒冷 的人哪，這件事你們要知道，要側耳聽我的話。
ACTS|2|15|這些人並不像你們所想的喝醉了，因為現在才早晨九點鐘。
ACTS|2|16|這正是藉著先知 約珥 所說的：
ACTS|2|17|『上帝說： 在末後的日子， 我要將我的靈澆灌凡血肉之軀的。 你們的兒女要說預言； 你們的少年要見異象； 你們的老人要做異夢。
ACTS|2|18|在那些日子，我要把我的靈澆灌， 甚至給我的僕人和婢女， 他們要說預言。
ACTS|2|19|在天上，我要顯出奇事， 在地下，我要顯出神蹟， 有血，有火，有煙霧。
ACTS|2|20|太陽要變為黑暗， 月亮要變為血， 這都在主大而光榮的日子未到以前。
ACTS|2|21|那時，凡求告主名的都必得救。』
ACTS|2|22|「 以色列 人哪，你們要聽我這些話： 拿撒勒 人耶穌就是上帝以異能、奇事、神蹟向你們證明出來的人，這些事是上帝藉著他在你們中間施行，正如你們自己知道的。
ACTS|2|23|他既按著上帝確定的旨意和預知被交與人，你們就藉著不法之人的手把他釘在十字架上，殺了。
ACTS|2|24|上帝卻將死的痛苦解除，使他復活了，因為他原不能被死拘禁。
ACTS|2|25|大衛 指著他說： 『我看見 主常在我眼前， 他在我右邊，使我不至於動搖。
ACTS|2|26|所以我心裏歡喜，我的舌頭快樂， 而且我的肉身要安居在指望中。
ACTS|2|27|因你必不將我的靈魂撇在陰間， 也不讓你的聖者見朽壞。
ACTS|2|28|你已將生命的道路指示我， 必使我在你面前充滿快樂。』
ACTS|2|29|「諸位弟兄，先祖 大衛 的事，我可以坦然地對你們說：他死了，也埋葬了，而且他的墳墓直到今日還在我們這裏。
ACTS|2|30|既然 大衛 是先知，他知道上帝曾向他起誓，要從他的後裔中立一位坐在他的寶座上。
ACTS|2|31|他預先看見了，就講論基督的復活，說： 『他不被撇在陰間； 他的肉身也不見朽壞。』
ACTS|2|32|這耶穌，上帝已經使他復活了，我們都是這事的見證人。
ACTS|2|33|他既被高舉在上帝的右邊，又從父受了所應許的聖靈，就把你們所看見所聽見的，澆灌下來。
ACTS|2|34|大衛 並沒有升到天上，但他自己說： 『主對我主說： 你坐在我的右邊，
ACTS|2|35|等我使你的仇敵作你的腳凳。』
ACTS|2|36|故此， 以色列 全家當確實知道，你們釘在十字架上的這位耶穌，上帝已經立他為主，為基督了。」
ACTS|2|37|眾人聽見這話，覺得扎心，就對 彼得 和其餘的使徒說：「諸位弟兄，我們該怎樣做呢？」
ACTS|2|38|彼得 對他們說：「你們各人要悔改，奉耶穌基督的名受洗，使你們的罪得赦免，就會領受所賜的聖靈。
ACTS|2|39|因為這應許是給你們和你們的兒女，並一切在遠方的人，就是給所有主—我們的上帝所召來的人。」
ACTS|2|40|彼得 還用更多別的話作見證，勸勉他們說：「你們當救自己脫離這彎曲的世代。」
ACTS|2|41|於是領受他話的人，都受了洗；那一天，門徒約添了三千人。
ACTS|2|42|他們都專注於使徒的教導和彼此的團契，擘餅和祈禱。
ACTS|2|43|眾人都心存敬畏；使徒們 又行了許多奇事神蹟。
ACTS|2|44|信的人都聚在一處，凡物公用，
ACTS|2|45|又賣了田產和家業，照每一個人所需要的分給他們。
ACTS|2|46|他們天天同心合意恆切地在聖殿裏敬拜，且在家中 擘餅，存著歡喜坦誠的心用飯，
ACTS|2|47|讚美上帝，得全體百姓的喜愛。主將得救的人天天加給他們。
ACTS|3|1|下午三點鐘禱告的時候， 彼得 和 約翰 上聖殿去。
ACTS|3|2|一個從母腹裏就是瘸腿的人正被人抬來，他們天天把他放在聖殿的一個叫 美門 的門口，求進聖殿的人施捨。
ACTS|3|3|他看見 彼得 、 約翰 將要進聖殿，就求他們施捨。
ACTS|3|4|彼得 和 約翰 定睛看他， 彼得 說：「看著我們！」
ACTS|3|5|那人就注目看他們，指望從他們得著甚麼。
ACTS|3|6|彼得 卻說：「金銀我都沒有，但我把我有的給你：奉 拿撒勒 人耶穌基督的名起來 行走！」
ACTS|3|7|於是 彼得 拉著他的右手，扶他起來；他的腳和踝骨立刻健壯了，
ACTS|3|8|就跳起來，站著，又開始行走。他跟他們進了聖殿，邊走邊跳，讚美上帝。
ACTS|3|9|百姓都看見他又行走，又讚美上帝，
ACTS|3|10|認得他是那素常坐在聖殿的 美門 口求人施捨的，就因他所遇到的事滿心驚訝詫異。
ACTS|3|11|那人正在稱為 所羅門 的廊下，拉住 彼得 和 約翰 ，大家都覺得很驚訝，一齊跑到他們那裏。
ACTS|3|12|彼得 看見，就對百姓說：「 以色列 人哪，為甚麼因這事而驚訝呢？為甚麼定睛看我們，以為我們憑自己的能力和虔誠使這人行走呢？
ACTS|3|13|亞伯拉罕 的上帝、 以撒 的上帝、 雅各 的上帝，就是我們列祖的上帝，已經榮耀了他的僕人耶穌，這耶穌就是你們交付官府的那位， 彼拉多 決定要釋放他時，你們卻在 彼拉多 面前棄絕了他。
ACTS|3|14|你們棄絕了那聖潔公義者，反而要求釋放一個兇手給你們。
ACTS|3|15|你們殺了那生命的創始者，上帝卻叫他從死人中復活；我們都是這事的見證人。
ACTS|3|16|因信他的名，他的名使你們所看見所認識的這人健壯了；正是他所賜的信心使這人在你們眾人面前完全好了。
ACTS|3|17|「如今，弟兄們，我知道你們做這事是出於無知，你們的官長也是如此。
ACTS|3|18|但上帝藉著眾先知的口預先宣告過基督將要受害的事，就這樣應驗了。
ACTS|3|19|所以，你們當悔改歸正，使你們的罪得以塗去，
ACTS|3|20|這樣，那安舒的日子就必從主面前來到；主也必差遣所預定給你們的基督耶穌來臨。
ACTS|3|21|他必須留在天上，直到萬物復興的時候，就是上帝自古藉著聖先知的口所說的。
ACTS|3|22|摩西 曾說：『主—你們 的上帝要從你們弟兄中給你們興起一位先知像我，凡他向你們所說的一切，你們都要聽從。
ACTS|3|23|凡不聽從那先知的，必將從民中滅絕。』
ACTS|3|24|從 撒母耳 以來和後繼的眾先知，凡說預言的，也都曾宣告這些日子。
ACTS|3|25|你們是先知的子孫，也是上帝與你們 祖宗所立之約的子孫，就是對 亞伯拉罕 說：『地上萬族都將因你的後裔得福。』
ACTS|3|26|上帝既興起他的僕人，就先差他到你們這裏來，賜福給你們，使各人回轉，離開你們的邪惡。」
ACTS|4|1|彼得 和 約翰 正向百姓說話的時候，祭司們、守殿官和撒都該人來了，
ACTS|4|2|就很煩惱，因為使徒們教導百姓，傳揚在耶穌的事上證明有死人復活，
ACTS|4|3|於是下手拿住他們；因為天已經晚了，就把他們押在拘留所到第二天。
ACTS|4|4|但聽道的人有許多信了，男人的數目約有五千。
ACTS|4|5|第二天，官長、長老和文士在 耶路撒冷 聚集，
ACTS|4|6|又有 亞那 大祭司、 該亞法 、 約翰 、 亞歷山大 ，和大祭司的親族都在那裏。
ACTS|4|7|他們叫使徒站在中間，問他們：「你們憑甚麼能力，奉誰的名做這事呢？」
ACTS|4|8|那時， 彼得 被聖靈充滿，對他們說：「民間的官長和長老啊，
ACTS|4|9|倘若今日我們被查問是因為在殘障的人身上所行的善事，就是這人怎麼得了痊癒，
ACTS|4|10|那麼，你們大家和 以色列 全民都當知道，站在你們面前的這人得痊癒，是因你們所釘在十字架、上帝使他從死人中復活的 拿撒勒 人耶穌基督的名。
ACTS|4|11|這位耶穌是： 『你們匠人所丟棄的石頭， 已成了房角的頭塊石頭。』
ACTS|4|12|除他以外，別無拯救，因為在天下人間，沒有賜下別的名，我們可以靠著得救。」
ACTS|4|13|他們見 彼得 、 約翰 的膽量，又看出他們原是沒有學問的平民，就很驚訝，認出他們曾是跟耶穌一起的；
ACTS|4|14|又看見那治好了的人和他們一同站著，就無話可駁。
ACTS|4|15|於是他們吩咐他們兩人從議會退出，就彼此商議，
ACTS|4|16|說：「我們當怎樣辦這兩個人呢？因為他們誠然行了一件明顯的神蹟，凡住在 耶路撒冷 的人都知道，我們也不能否認。
ACTS|4|17|但為避免這事越發在民間傳揚，我們必須威嚇他們，叫他們不可再奉這名對任何人講論。」
ACTS|4|18|於是他們叫了兩人來，禁止他們，再不可奉耶穌的名講論或教導人。
ACTS|4|19|彼得 和 約翰 回答他們說：「聽從你們，不聽從上帝，在上帝面前合理不合理，你們自己判斷吧！
ACTS|4|20|我們所看見所聽見的，我們不能不說。」
ACTS|4|21|官長為百姓的緣故，想不出任何法子懲罰他們，只好威嚇一番就把他們釋放了；這是因眾人為了所行的奇事都歸榮耀與上帝。
ACTS|4|22|原來經歷這神蹟醫好的人有四十多歲了。
ACTS|4|23|二人既被釋放，就到自己的人那裏去，把祭司長和長老所說的話都告訴他們。
ACTS|4|24|他們聽見了，就同心合意地高聲向上帝說：「主宰啊！你是那創造天、地、海和其中萬物的；
ACTS|4|25|你曾藉著聖靈託你僕人—我們祖宗 大衛 的口說： 『外邦為甚麼擾動？ 萬民為甚麼謀算虛妄的事？
ACTS|4|26|地上的君王都站穩， 臣宰也聚集一處， 要對抗主，對抗主的受膏者 』。
ACTS|4|27|希律 和 本丟．彼拉多 ，同外邦人和 以色列 民，果然在這城裏聚集，要攻打你所膏的聖僕耶穌，
ACTS|4|28|做了你手和你旨意所預定必成就的事。
ACTS|4|29|主啊，現在求你鑒察，他們的威嚇，使你僕人放膽講你的道，
ACTS|4|30|伸出你的手來，讓醫治、神蹟、奇事藉著你聖僕耶穌的名行出來。」
ACTS|4|31|他們禱告完了，聚會的地方震動；他們都被聖靈充滿，放膽傳講上帝的道。
ACTS|4|32|許多信徒都一心一意，沒有一人說他的任何東西是自己的，都是大家公用。
ACTS|4|33|使徒以大能見證主耶穌 復活；眾人也都蒙了大恩。
ACTS|4|34|他們當中沒有一個缺乏的，因為凡有田產房屋的都賣了，把所賣的錢拿來，
ACTS|4|35|放在使徒腳前，照每人所需要的，分給每人。
ACTS|4|36|有一個 利未 人，名叫 約瑟 ，使徒稱他為 巴拿巴 （ 巴拿巴 翻出來就是安慰之子），生在 塞浦路斯 。
ACTS|4|37|他有田地，也賣了，把錢拿來，放在使徒腳前。
ACTS|5|1|有一個人，名叫 亞拿尼亞 ，同他的妻子 撒非喇 ，賣了田產，
ACTS|5|2|把錢私自留下一部分，他的妻子也知道，其餘的部分拿來放在使徒腳前。
ACTS|5|3|彼得 說：「 亞拿尼亞 ！為甚麼撒但充滿了你的心，使你欺騙聖靈，把賣田地的錢私自留下一部分呢？
ACTS|5|4|田地還沒有賣，不是你自己的嗎？既賣了，錢不是你作主嗎？你怎麼心裏會想這樣做呢？你不是欺騙人，是欺騙上帝！」
ACTS|5|5|亞拿尼亞 一聽見這些話，就仆倒，斷了氣；所有聽見的人都非常懼怕。
ACTS|5|6|有些年輕人起來，把他裹好，抬出去埋葬了。
ACTS|5|7|約過了三小時，他的妻子進來，還不知道所發生的事。
ACTS|5|8|彼得 對她說：「你告訴我，你們賣田地的錢就是這些嗎？」她說：「就是這些。」
ACTS|5|9|彼得 對她說：「你們為甚麼同謀來試探主的靈呢？你看，埋葬你丈夫之人的腳已到門口，他們也要把你抬出去。」
ACTS|5|10|她立刻仆倒在 彼得 腳前，斷了氣。那些年輕人進來，見她已經死了，就把她抬出去，埋在她丈夫旁邊。
ACTS|5|11|全教會和所有聽見這些事的人都非常懼怕。
ACTS|5|12|主藉使徒的手在民間行了許多神蹟奇事；他們都同心合意地聚集在 所羅門 的廊下。
ACTS|5|13|其餘的人沒有一個敢接近他們，百姓卻尊重他們。
ACTS|5|14|信主的人越發增添，連男帶女都很多，
ACTS|5|15|甚至有人將病人抬到街上，放在床上或褥子上，好讓 彼得 走過來的時候，或者影子投在一些人身上。
ACTS|5|16|還有許多人帶著病人和被污靈纏磨的，從 耶路撒冷 四圍的城鎮來，他們全都得了醫治。
ACTS|5|17|於是，大祭司採取行動，他和他所有一起的人，就是撒都該派的人，滿心忌恨，
ACTS|5|18|就下手拿住使徒，把他們押在公共拘留所內。
ACTS|5|19|但在夜間主的使者開了監門，領他們出來，說：
ACTS|5|20|「你們去，站在聖殿裏，把這生命的一切話講給百姓聽。」
ACTS|5|21|使徒聽了這話，天將亮的時候就進聖殿裏去教導人。大祭司和他一起的人來了，叫齊議會的人和 以色列 人的眾長老，然後派人到監牢裏去把使徒提出來。
ACTS|5|22|但差役到了，不見他們在監裏，就回來稟報，
ACTS|5|23|說：「我們看見監牢關得很緊，警衛也站在門外，但打開門來，裏面一個人都不見。」
ACTS|5|24|守殿官和祭司長聽了這些話，心裏困惑，不知這事將來如何。
ACTS|5|25|有一個人來稟報說：「你們押在監裏的人，現在站在聖殿裏教導百姓。」
ACTS|5|26|於是守殿官和差役去帶使徒來，並沒有用暴力，因為怕百姓用石頭打他們。
ACTS|5|27|他們把使徒帶來了，就叫他們站在議會前。大祭司問他們，
ACTS|5|28|說：「我們不是嚴嚴地禁止你們，不可奉這名教導人嗎？ 看，你們倒把你們的道理充滿了 耶路撒冷 ，想要叫這人的血歸到我們身上！」
ACTS|5|29|彼得 和眾使徒回答：「我們必須順從上帝，勝於順從人。
ACTS|5|30|你們掛在木頭上殺害的耶穌，我們祖宗的上帝已經使他復活了。
ACTS|5|31|上帝把他高舉在自己的右邊，使他作元帥，作救主，使 以色列 人得以悔改，並且罪得赦免。
ACTS|5|32|我們是這些事的見證人；上帝賜給順從的人的聖靈也為這些事作見證。」
ACTS|5|33|議會的人聽了極其惱怒，想要殺他們。
ACTS|5|34|但有一個法利賽人，名叫 迦瑪列 ，是眾百姓所敬重的律法教師，他在議會中站起來，吩咐人把使徒暫且帶到外面去，
ACTS|5|35|然後對眾人說：「 以色列 人哪，對於這些人，你們應當小心怎樣處理。
ACTS|5|36|從前 杜達 出現，自命不凡，附從他的人數約有四百；他被殺後，附從他的人全都散了，歸於無有。
ACTS|5|37|此後，登記戶籍的時候，又有 加利利 的 猶大 出現，引誘百姓跟從他，他也滅亡，附從他的人也都四散了。
ACTS|5|38|現在，我勸你們不要管這些人，任憑他們吧！他們所謀所為若是出於人，必要敗壞；
ACTS|5|39|若是出於上帝，你們就不能敗壞他們，恐怕你們倒是攻擊上帝了。」 議會的人被他說服了，
ACTS|5|40|就叫使徒來，把他們打了，又吩咐他們不可奉耶穌的名講道，然後把他們釋放了。
ACTS|5|41|他們歡歡喜喜地離開議會，因他們算配為這名受辱。
ACTS|5|42|他們就每日在聖殿裏，在家裏 ，不住地教導人，傳耶穌是基督的福音。
ACTS|6|1|那些日子，門徒增多，有說希臘話的 猶太 人向 希伯來 人發怨言，因為在日常的供給上忽略了他們的寡婦。
ACTS|6|2|十二使徒叫眾門徒來，說：「我們撇下上帝的道去管理飯食，是不合宜的。
ACTS|6|3|所以弟兄們，當從你們中間選出七個有好名聲、滿有聖靈和智慧，我們派他們管理這事。
ACTS|6|4|至於我們，我們要專注於祈禱和傳道的事奉。」
ACTS|6|5|這話使全會眾都喜悅，就揀選了 司提反 —他是一個滿有信心和聖靈的人；他們又揀選了 腓利 、 伯羅哥羅 、 尼迦挪 、 提門 、 巴米拿 ，並皈依 猶太 教的 安提阿 人 尼哥拉 ，
ACTS|6|6|叫他們站在使徒面前，使徒禱告後，就為他們按手。
ACTS|6|7|上帝的道興旺起來；在 耶路撒冷 門徒數目增加得很多，也有許多祭司聽從了這信仰。
ACTS|6|8|司提反 滿有恩惠和能力，在民間行了大奇事和神蹟。
ACTS|6|9|當時有從稱為「自由人」會堂，並 古利奈 、 亞歷山大 會堂來的人，還有些從 基利家 、 亞細亞 來的人，起來和 司提反 辯論。
ACTS|6|10|司提反 是以智慧和聖靈說話，眾人抵擋不住，
ACTS|6|11|就收買人來說：「我們聽見他說褻瀆 摩西 和上帝的話。」
ACTS|6|12|他們又煽動百姓、長老和文士，就突然來捉拿他，把他帶到議會去，
ACTS|6|13|設下假見證，說：「這個人不斷地說話，侮辱神聖的地方和律法。
ACTS|6|14|我們曾聽見他說，這 拿撒勒 人耶穌要毀壞這地方，也要改變 摩西 所交給我們的規矩。」
ACTS|6|15|在議會裏坐著的人都定睛看他，見他的面貌好像天使的面貌。
ACTS|7|1|大祭司說：「果真有這些事嗎？」
ACTS|7|2|司提反 說：「諸位父老弟兄請聽！從前我們的祖宗 亞伯拉罕 在 美索不達米亞 ，還沒有住在 哈蘭 的時候，榮耀的上帝向他顯現，
ACTS|7|3|對他說：『你要離開本地和親族，往我所要指示你的地去。』
ACTS|7|4|他就離開 迦勒底 人的地方，住在 哈蘭 。他父親死了以後，上帝使他從那裏搬到你們現在所住的地方。
ACTS|7|5|在這裏上帝並沒有給他產業，連立足的地方都沒有，但應許要將這地賜給他和他的後裔為業，雖然那時他還沒有兒子。
ACTS|7|6|上帝這樣說：『他的後裔必寄居外邦，那裏的人要使他們作奴隸，苦待他們四百年。』
ACTS|7|7|上帝又說：『但我要懲罰使他們作奴隸的那國。以後他們要出來，在這地方事奉我。』
ACTS|7|8|上帝又賜他割禮的約。於是 亞伯拉罕 生了 以撒 ，在第八日給他行了割禮；後來 以撒 生 雅各 ， 雅各 生十二位先祖。
ACTS|7|9|「先祖嫉妒 約瑟 ，把他賣到 埃及 去，上帝卻與他同在，
ACTS|7|10|救他脫離一切苦難，又使他在 埃及 王法老面前蒙恩，又有智慧。法老派他作 埃及 國的宰相兼管法老的全家。
ACTS|7|11|後來全 埃及 和 迦南 遭遇饑荒和大災難，我們的祖宗絕了糧。
ACTS|7|12|雅各 聽見在 埃及 有糧，就打發我們的祖宗初次往那裏去。
ACTS|7|13|第二次 約瑟 與兄弟們相認，法老才認識他的家族。
ACTS|7|14|約瑟 就打發人，請父親 雅各 和全族七十五個人都來。
ACTS|7|15|於是 雅各 下了 埃及 ，後來他和我們的祖宗都死在那裏；
ACTS|7|16|他們又被遷到 示劍 ，葬於 亞伯拉罕 在 示劍 用銀子從 哈抹 子孫 買來的墳墓裏。
ACTS|7|17|「當上帝應許 亞伯拉罕 的日期將到的時候， 以色列 人在 埃及 人丁興旺，
ACTS|7|18|直到另一位不認識 約瑟 的王興起統治 埃及 。
ACTS|7|19|他用詭計待我們的宗族，苦待我們的祖宗，強迫他們丟棄嬰孩，使嬰孩不能存活。
ACTS|7|20|就在那時， 摩西 生了下來，上帝看為俊美，在父親家裏被撫養了三個月。
ACTS|7|21|他被丟棄的時候，法老的女兒拾了去，當自己的兒子撫養。
ACTS|7|22|摩西 學了 埃及 人一切的學問，說話辦事都有才能。
ACTS|7|23|「他到了四十歲，心中起意去看望他的弟兄 以色列 人。
ACTS|7|24|他見他們中的一個人受冤屈，就庇護他，為那被壓迫的人報仇，打死了那 埃及 人。
ACTS|7|25|他以為他的弟兄們必明白上帝是藉他的手搭救他們，他們卻不明白。
ACTS|7|26|第二天，他遇見有人在打架，就想勸他們和好，說：『二位，你們是弟兄，為甚麼彼此欺負呢？』
ACTS|7|27|那欺負鄰舍的人把他推開，說：『誰立你作我們的領袖和審判官呢？
ACTS|7|28|難道你要殺我像昨天殺那 埃及 人一樣嗎？』
ACTS|7|29|摩西 聽見這話就逃走了，寄居於 米甸 地，在那裏生了兩個兒子。
ACTS|7|30|「過了四十年，在 西奈山 的曠野，有一位天使在荊棘的火焰中向 摩西 顯現。
ACTS|7|31|摩西 見了那異象，覺得很驚訝，正往前觀看的時候，有主的聲音說：
ACTS|7|32|『我是你列祖的上帝，就是 亞伯拉罕 、 以撒 、 雅各 的上帝。』 摩西 戰戰兢兢，不敢觀看。
ACTS|7|33|主對他說：『把你腳上的鞋脫下來，因為你所站的地方是聖地。
ACTS|7|34|我的百姓在 埃及 所受的困苦，我確實看見了；他們悲嘆的聲音，我也聽見了。我下來要救他們。現在，你來，我要差你往 埃及 去。』
ACTS|7|35|「這 摩西 就是有人曾棄絕他說『誰立你作我們的領袖和審判官』的，上帝卻藉那在荊棘中顯現的天使的手差派他作領袖，作解救者。
ACTS|7|36|這人領 以色列 人出來，在 埃及 地，在 紅海 ，在曠野的四十年間行了奇事神蹟。
ACTS|7|37|這人是 摩西 ，就是那曾對 以色列 人說『上帝要從你們弟兄中給你們興起一位先知像我』的。
ACTS|7|38|這人是那曾在曠野的會眾中和 西奈山 上，與那對他說話的天使同在，又與我們祖宗同在的，他領受了活潑的聖言傳給我們。
ACTS|7|39|我們的祖宗不肯聽從，反棄絕他，他們的心轉向 埃及 ，
ACTS|7|40|對 亞倫 說：『你為我們造神明，在我們前面引路，因為領我們出 埃及 地的這個 摩西 ，我們不知道他遭遇了甚麼事。』
ACTS|7|41|那時，他們造了一個牛犢，又拿祭物獻給那像，為自己手所做的工作歡躍。
ACTS|7|42|但是上帝轉臉不顧，任憑他們祭拜天上的日月星辰，正如先知書上所寫的： 『 以色列 家啊，你們四十年間在曠野， 何曾將犧牲和祭物獻給我？
ACTS|7|43|你們抬著 摩洛 的帳幕 和 理番 ──你們神明的星， 就是你們所造為要敬拜的像。 因此，我要把你們遷到 巴比倫 外去。』
ACTS|7|44|「我們的祖宗在曠野，有作證的會幕，是上帝吩咐 摩西 照著他所看見的樣式做的。
ACTS|7|45|這帳幕，我們的祖宗同 約書亞 相繼承受了，當上帝在他們面前趕走外邦人的時候，他們把這帳幕搬進承受為業之地，直存到 大衛 的日子。
ACTS|7|46|大衛 在上帝面前蒙恩，祈求為 雅各 的家 預備居所。
ACTS|7|47|但卻是 所羅門 為上帝造成殿宇。
ACTS|7|48|其實，至高者並不住人手所造的，就如先知所言：
ACTS|7|49|『主說：天是我的寶座， 地是我的腳凳。 你們要為我造怎樣的殿宇？ 哪裏是我安歇的地方呢？
ACTS|7|50|這一切不都是我手所造的嗎？』
ACTS|7|51|「你們這硬著頸項，心與耳未受割禮的人哪，時常抗拒聖靈！你們的祖宗怎樣，你們也怎樣。
ACTS|7|52|先知中有哪一個不是受你們祖宗的迫害呢？他們把預先宣告那義者要來的人殺了。如今你們成了那義者的出賣者和兇手了。
ACTS|7|53|你們領受了天使所傳佈的律法，竟不遵守。」
ACTS|7|54|眾人聽見這些話，心中極其惱怒，向 司提反 咬牙切齒。
ACTS|7|55|但 司提反 滿有聖靈，定睛望天，看見上帝的榮耀，又看見耶穌站在上帝的右邊，
ACTS|7|56|就說：「我看見天開了，人子站在上帝的右邊。」
ACTS|7|57|眾人大聲喊叫，摀著耳朵，齊心衝向他，
ACTS|7|58|把他推到城外，用石頭打他。作見證的人把他們的衣裳放在一個名叫 掃羅 的青年腳前。
ACTS|7|59|他們正用石頭打 司提反 的時候，他呼求說：「主耶穌啊，求你接納我的靈魂！」
ACTS|7|60|然後他跪下來，大聲喊著：「主啊，不要將這罪歸於他們！」說了這話，就長眠了。
ACTS|8|1|掃羅 也贊同處死他。從那一天開始， 耶路撒冷 的教會遭受到大迫害，除了使徒以外，眾門徒都分散在 猶太 和 撒瑪利亞 各處。
ACTS|8|2|有些虔誠的人把 司提反 埋葬了，為他大大哀哭。
ACTS|8|3|掃羅 卻殘害教會，挨家挨戶地進去，拉著男女關在監裏。
ACTS|8|4|那些分散的人往各地去傳福音的道。
ACTS|8|5|腓利 下 撒瑪利亞城 去 ，向當地人宣講基督。
ACTS|8|6|眾人都聚精會神，同心合意地聽 腓利 所說的話，一邊聽他的話，一邊看他所行的神蹟。
ACTS|8|7|因為有許多人被污靈附著，那些污靈大聲呼叫，從他們身上出來；還有許多癱瘓的、瘸腿的都得了醫治。
ACTS|8|8|那城裏，有極大的喜樂。
ACTS|8|9|有一個人名叫 西門 ，向來在那城裏行邪術，自命為大人物，使 撒瑪利亞 的居民驚奇。
ACTS|8|10|所有的人，從小到大都聽從他，說：「這個人就是上帝的能力，那稱為大能者的。」
ACTS|8|11|他們聽從他，因他很久以來用邪術使他們驚奇。
ACTS|8|12|當他們信了 腓利 所傳上帝國的福音和耶穌基督的名，連男帶女都受了洗。
ACTS|8|13|西門 自己也信了；既受了洗，就常與 腓利 在一處，看見他所行的神蹟和大異能，就覺得很驚奇。
ACTS|8|14|在 耶路撒冷 的使徒聽見 撒瑪利亞 人領受了上帝的道，就打發 彼得 和 約翰 到他們那裏去。
ACTS|8|15|兩個人下去，就為他們禱告，要讓他們領受聖靈，
ACTS|8|16|因為聖靈還沒有降在他們任何一個人身上，他們只奉主耶穌的名受了洗。
ACTS|8|17|於是使徒按手在他們頭上，他們就領受了聖靈。
ACTS|8|18|西門 看見使徒一按手，就有聖靈賜下，就拿錢給使徒，
ACTS|8|19|說：「請把這權柄也給我，使我手按著誰，誰就可以領受聖靈。」
ACTS|8|20|彼得 對他說：「你的銀子和你一同滅亡吧！因為你想上帝的恩賜是可以用錢買的。
ACTS|8|21|你在這道上無份無關；因為你在上帝面前心懷不正。
ACTS|8|22|你要為你這樣的惡而悔改，祈求主，或者你心裏的意念可得赦免。
ACTS|8|23|我看出你正在苦膽之中，被不義捆綁著。」
ACTS|8|24|西門 回答說：「請你們為我求主，使你們所說的，沒有一樣臨到我身上。」
ACTS|8|25|使徒既作了見證，並且宣講了主的道，就回 耶路撒冷 去，一路在 撒瑪利亞 好些村莊傳揚福音。
ACTS|8|26|有主的一個使者對 腓利 說：「起來！向南走，往那從 耶路撒冷 下 迦薩 的路上去。」那路是曠野。
ACTS|8|27|腓利 就起身去了。不料，有一個 埃塞俄比亞 人，是個有大權的太監，在 埃塞俄比亞 女王 甘大基 的手下總管銀庫，他上 耶路撒冷 去禮拜。
ACTS|8|28|回程中，他坐在車上，正念著 以賽亞 先知的書，
ACTS|8|29|聖靈對 腓利 說：「你去！靠近那車走。」
ACTS|8|30|腓利 就跑到太監那裏，聽見他正在念 以賽亞 先知的書，就說：「你明白你所念的嗎？」
ACTS|8|31|他說：「沒有人指教我，怎能明白呢？」於是他請 腓利 上車，與他同坐。
ACTS|8|32|他所念的那段經文是這樣： 「他像羊被牽去宰殺， 又像羔羊在剪毛的人手下無聲， 他也是這樣不開口。
ACTS|8|33|他卑微的時候，得不到公義的審判， 誰能述說他的身世？ 因為他的生命從地上被奪去。」
ACTS|8|34|太監回答 腓利 說：「請問，先知說這話是指誰，是指自己，還是指別人呢？」
ACTS|8|35|腓利 就開口，從這段經文開始，對他傳講耶穌的福音。
ACTS|8|36|二人正沿路往前走，到了有水的地方，太監說：「看哪！這裏有水，有甚麼能阻止我受洗呢？」
ACTS|8|37|
ACTS|8|38|於是他吩咐把車停下來， 腓利 和太監二人一同下到水裏， 腓利 就給他施洗。
ACTS|8|39|他們從水裏上來，主的靈把 腓利 提了去，太監再也看不見他了，就歡歡喜喜地上路。
ACTS|8|40|後來有人在 亞鎖都 遇見 腓利 ；他走遍那地方，在各城宣揚福音，一直到 凱撒利亞 。
ACTS|9|1|掃羅 不斷用威嚇兇悍的口氣向主的門徒說話。他去見大祭司，
ACTS|9|2|要求發信給 大馬士革 的各會堂，若是找著信奉這道的人，無論男女，都准他捆綁帶到 耶路撒冷 。
ACTS|9|3|掃羅 在途中，將到 大馬士革 的時候，忽然有一道光從天上下來，四面照射著他，
ACTS|9|4|他就仆倒在地，聽見有聲音對他說：「 掃羅 ！ 掃羅 ！你為甚麼迫害我？」
ACTS|9|5|他說：「主啊！你是誰？」主說：「我就是你所迫害的耶穌。
ACTS|9|6|起來！進城去，你應該做的事，必有人告訴你。」
ACTS|9|7|同行的人站在那裏，說不出話來，因為他們聽見聲音，卻看不見人。
ACTS|9|8|掃羅 從地上起來，睜開眼睛，竟不能看見甚麼。有人拉他的手，領他進了 大馬士革 。
ACTS|9|9|他三天甚麼都看不見，也不吃也不喝。
ACTS|9|10|那時，在 大馬士革 有一個門徒，名叫 亞拿尼亞 。主在異象中對他說：「 亞拿尼亞 ！」他說：「主啊，我在這裏。」
ACTS|9|11|主對他說：「起來！往那叫 直街 的路去，在 猶大 的家裏，去找一個 大數 人，名叫 掃羅 ；他正在禱告，
ACTS|9|12|在異象中 看見了一個人，名叫 亞拿尼亞 ，進來為他按手，讓他能再看得見。」
ACTS|9|13|亞拿尼亞 回答：「主啊，我聽見許多人講到這個人，說他怎樣在 耶路撒冷 多多苦待你的聖徒，
ACTS|9|14|並且他在這裏有從祭司長得來的權柄，要捆綁一切求告你名的人。」
ACTS|9|15|主對他說：「你只管去。他是我所揀選的器皿，要在外邦人、君王和 以色列 人面前宣揚我的名。
ACTS|9|16|我也要指示他，為我的名必須受許多的苦難。」
ACTS|9|17|亞拿尼亞 就去了，進入那家，把手按在 掃羅 身上，說：「 掃羅 弟兄，在你來的路上向你顯現的主，就是耶穌，打發我來，叫你能再看得見，又被聖靈充滿。」
ACTS|9|18|掃羅 的眼睛上立刻好像有鱗一般的東西掉下來，他就能再看得見，於是他起來，受了洗，
ACTS|9|19|吃過飯體力就恢復了。 掃羅 和 大馬士革 的門徒一起住了些日子，
ACTS|9|20|立刻在各會堂裏傳揚耶穌，說他是上帝的兒子。
ACTS|9|21|凡聽見的人都很驚奇，說：「在 耶路撒冷 殘害求告這名的不就是這個人嗎？他不是到這裏來要捆綁他們，帶到祭司長那裏去嗎？」
ACTS|9|22|但 掃羅 越發有能力，駁倒住在 大馬士革 的 猶太 人，證明耶穌是基督。
ACTS|9|23|過了好些日子， 猶太 人商議要殺 掃羅 ，
ACTS|9|24|但他們的計謀被 掃羅 知道了。他們晝夜在城門守候著要殺他。
ACTS|9|25|他的門徒就在夜間用筐子把他從城牆上縋了下去。
ACTS|9|26|掃羅 到了 耶路撒冷 ，想與門徒結交，大家卻都怕他，不信他是門徒。
ACTS|9|27|只有 巴拿巴 接待他，領他去見使徒，把他在路上怎麼看見主，主怎麼向他說話，他在 大馬士革 怎麼奉耶穌的名放膽傳道，都述說出來。
ACTS|9|28|於是 掃羅 在 耶路撒冷 同門徒出入來往，奉主的名放膽傳道，
ACTS|9|29|並和說 希臘 話的 猶太 人講論辯駁，他們卻想法子要殺他。
ACTS|9|30|弟兄們知道了，就帶他下 凱撒利亞 ，送他往 大數 去。
ACTS|9|31|那時， 猶太 、 加利利 、 撒瑪利亞 各處的教會都得平安，建立起來，凡事敬畏主，蒙聖靈的安慰，人數逐漸增多。
ACTS|9|32|彼得 在眾信徒中到處奔波的時候，也到了住在 呂大 的聖徒那裏。
ACTS|9|33|他在那裏遇見一個人，名叫 以尼雅 ，得了癱瘓，在褥子上躺了八年。
ACTS|9|34|彼得 對他說：「 以尼雅 ，耶穌基督醫好你了，起來！整理你的褥子吧。」他立刻就起來了。
ACTS|9|35|凡住 呂大 和 沙崙 的人都看見了他，就歸向主。
ACTS|9|36|在 約帕 有一個女門徒，名叫 大比大 ，翻出來的意思是 多加 ；她廣行善事，多施賙濟。
ACTS|9|37|當時，她患病死了，有人把她清洗後，停在樓上。
ACTS|9|38|呂大 原與 約帕 相近；門徒聽見 彼得 在那裏，就派兩個人去見他，央求他說：「請快到我們那裏去，不要耽延。」
ACTS|9|39|彼得 就起身和他們同去。他到了，就有人領他上樓。眾寡婦都站在 彼得 旁邊哭，拿 多加 與她們同在時所做的內衣外衣給他看。
ACTS|9|40|彼得 叫她們都出去，然後跪下禱告，轉身對著屍體說：「 大比大 ，起來！」她就睜開眼睛，看見 彼得 ，就坐了起來。
ACTS|9|41|彼得 伸手扶她起來，叫那些聖徒和寡婦都進來，把 多加 活活地交給他們。
ACTS|9|42|這事傳遍了 約帕 ，就有許多人信了主。
ACTS|9|43|此後， 彼得 在 約帕 一個皮革匠 西門 的家裏住了好些日子。
ACTS|10|1|在 凱撒利亞 有一個人名叫 哥尼流 ，是 意大利 營的百夫長。
ACTS|10|2|他是個虔誠人，他和全家都敬畏上帝。他多多賙濟百姓，常常向上帝禱告。
ACTS|10|3|有一天，約在下午三點鐘，他在異象中清楚看見上帝的一個使者進來，到他那裏，對他說：「 哥尼流 。」
ACTS|10|4|哥尼流 定睛看他，驚惶地說：「主啊，甚麼事？」天使對他說：「你的禱告和你的賙濟已達到上帝面前，蒙記念了。
ACTS|10|5|現在你要派人往 約帕 去，請一位稱為 彼得 的 西門 來。
ACTS|10|6|他住在一個皮革匠 西門 的家裏，房子就在海邊。」
ACTS|10|7|向他說話的天使離開後， 哥尼流 叫了兩個僕人和常伺候他的一個虔誠的兵來，
ACTS|10|8|把一切的事都講給他們聽，然後就派他們往 約帕 去。
ACTS|10|9|第二天，他們走路將近那城，約在正午， 彼得 上房頂去禱告。
ACTS|10|10|他覺得餓了，想要吃。那家的人正預備飯的時候， 彼得 魂遊象外，
ACTS|10|11|看見天開了，有一塊好像大布的東西降下，四角 吊著縋在地上，
ACTS|10|12|裏面有地上各樣四腳的走獸、爬蟲和天上的飛鳥。
ACTS|10|13|又有聲音對他說：「 彼得 ，起來！宰了吃。」
ACTS|10|14|彼得 卻說：「主啊，絕對不可！凡污俗和不潔淨的東西，我從來沒有吃過。」
ACTS|10|15|第二次有聲音再對他說：「上帝所潔淨的，你不可當作污俗的。」
ACTS|10|16|這樣一連三次，那東西隨即收回天上去了。
ACTS|10|17|正當 彼得 心裏困惑，不知所看見的異象是甚麼意思時， 哥尼流 所差來的人已經找到了 西門 的家，站在門外，
ACTS|10|18|喊著問有沒有一位稱為 彼得 的 西門 住在這裏。
ACTS|10|19|彼得 還在思考那異象的時候，聖靈對他說：「有三個人來找你。
ACTS|10|20|起來，下去，跟他們同去，不要疑惑，因為是我差他們來的。」
ACTS|10|21|於是 彼得 下去見那些人，說：「我就是你們要找的人，你們是為了甚麼緣故在這裏？」
ACTS|10|22|他們說：「百夫長 哥尼流 是個義人，敬畏上帝，為 猶太 全民族所稱讚。他蒙一位聖天使指示，叫他請你到他家裏去，要聽你講話。」
ACTS|10|23|彼得 就請他們進去住宿。 次日，他起身和他們同去，還有 約帕 的幾個弟兄跟他一起去。
ACTS|10|24|又次日，他 進入 凱撒利亞 ， 哥尼流 已經請了他的親朋好友在等候他們。
ACTS|10|25|彼得 一進去， 哥尼流 就迎接他，俯伏在他腳前拜他。
ACTS|10|26|但是 彼得 拉他起來，說：「你起來，我自己也不過是人。」
ACTS|10|27|彼得 和他一邊說話一邊進去，見有好些人聚集，
ACTS|10|28|就對他們說：「你們知道， 猶太 人和別國的人結交來往本是不合規矩的，但上帝已經指示我，無論甚麼人都不可看作污俗或不潔淨的。
ACTS|10|29|所以，我一被邀請，沒有推辭就來了。現在請問，你們為甚麼叫我來呢？」
ACTS|10|30|哥尼流 說：「四天前，這個時候，我在家中守著下午三點鐘的禱告，忽然有一個人穿著明亮的衣裳站在我面前，
ACTS|10|31|說：『 哥尼流 ，你的禱告已蒙垂聽，你的賙濟在上帝面前已蒙記念了。
ACTS|10|32|你要派人往 約帕 去，請那稱為 彼得 的 西門 來，他住在海邊一個皮革匠 西門 的家裏。』
ACTS|10|33|所以我立刻派人去請你。你來了真好。現在我們都在上帝面前，要聽主 吩咐你的一切話。」
ACTS|10|34|彼得 開口說：「我真的看出上帝是不偏待人的。
ACTS|10|35|不但如此，在各國中那敬畏他而行義的人都為他所悅納。
ACTS|10|36|上帝藉著耶穌基督—他是萬有的主—傳和平的福音，把這道傳給 以色列 人。
ACTS|10|37|這話在 約翰 傳揚洗禮以後，從 加利利 起，傳遍了 猶太 。上帝怎樣以聖靈和能力膏了 拿撒勒 人耶穌，這都是你們知道的。他到處奔波，行善事，醫好凡被魔鬼壓制的人，因為上帝與他同在。
ACTS|10|38|
ACTS|10|39|他在 猶太 人之地和 耶路撒冷 所行的一切事，有我們作見證人。他們竟把他掛在木頭上殺了。
ACTS|10|40|第三天，上帝使他復活，使他顯現出來；
ACTS|10|41|不是顯現給所有的人看，而是顯現給上帝預先所揀選為他作見證的人看，就是我們這些在他從死人中復活以後和他同吃同喝的人。
ACTS|10|42|他吩咐我們傳道給眾人，證明他是上帝所立定，要作審判活人、死人的審判者。
ACTS|10|43|眾先知也為這人作見證：凡信他的人，必藉著他的名得蒙赦罪。」
ACTS|10|44|彼得 還在說這些話的時候，聖靈降在一切聽道的人身上。
ACTS|10|45|那些奉割禮的信徒和 彼得 同來，見聖靈的恩賜也澆在外邦人身上，就都驚奇；
ACTS|10|46|因聽見他們說方言 ，稱讚上帝為大。於是 彼得 回答：
ACTS|10|47|「這些人既受了聖靈，跟我們一樣，誰能阻止用水給他們施洗呢？」
ACTS|10|48|他就吩咐奉耶穌基督的名給他們施洗。於是他們請 彼得 住了幾天。
ACTS|11|1|使徒和在 猶太 的眾弟兄聽到外邦人也領受了上帝的道。
ACTS|11|2|等到 彼得 上了 耶路撒冷 ，那些奉割禮的信徒和他爭辯，
ACTS|11|3|說：「你竟進入未受割禮之人當中，和他們一同吃飯！」
ACTS|11|4|彼得 就開始把這事逐一向他們解釋，說：
ACTS|11|5|「我在 約帕城 裏禱告的時候，魂遊象外，看見異象，有一塊好像大布的東西降下，四角吊著從天縋下，直來到我跟前。
ACTS|11|6|我定睛觀看，見內中有地上四腳的牲畜、野獸、爬蟲和天上的飛鳥。
ACTS|11|7|我還聽見有聲音對我說：『 彼得 ，起來！宰了吃。』
ACTS|11|8|我說：『主啊，絕對不可！凡污俗或不潔淨的東西從來沒有進過我的口。』
ACTS|11|9|第二次，有聲音從天上回答：『上帝所潔淨的，你不可當作污俗的。』
ACTS|11|10|這樣一連三次，然後一切就都收回天上去了。
ACTS|11|11|正當那時，有三個從 凱撒利亞 差來見我的人，站在我們 所住的屋子門前。
ACTS|11|12|聖靈吩咐我和他們同去，不要疑惑，還有這六位弟兄也跟我一起去，我們進了那人的家。
ACTS|11|13|那人就告訴我們，他如何看見一位天使站在他家裏，說：『你派人往 約帕 去，請那稱為 彼得 的 西門 來，
ACTS|11|14|他有話要告訴你，因這些話你和你的全家都可以得救。』
ACTS|11|15|我一開始講話，聖靈就降在他們身上，正像當初降在我們身上一樣。
ACTS|11|16|我就想起主的話如何說：『 約翰 用水施洗，但你們要在聖靈裏受洗。』
ACTS|11|17|既然上帝給他們恩賜，像在我們信主耶穌基督的時候給了我們一樣，我是誰，能攔阻上帝嗎？」
ACTS|11|18|眾人聽見這些話，就不說話了，只歸榮耀給上帝，說：「這樣看來，上帝也賜恩給外邦人，使他們悔改得生命了。」
ACTS|11|19|那些因 司提反 的事遭患難而四處分散的門徒，直走到 腓尼基 、 塞浦路斯 和 安提阿 。他們不向別人講道，只向 猶太 人講。
ACTS|11|20|但內中有 塞浦路斯 和 古利奈 人，他們到了 安提阿 也向 希臘 人傳講主耶穌的福音 。
ACTS|11|21|主的手與他們同在，信而歸主的人數很多。
ACTS|11|22|這風聲傳到 耶路撒冷 教會的人耳中，他們就打發 巴拿巴 到 安提阿 去。
ACTS|11|23|他到了那裏，看見上帝所賜的恩就歡喜，勸勉眾人要立定心志，恆久靠主。
ACTS|11|24|這 巴拿巴 原是個好人，滿有聖靈和信心，於是有許多人歸服了主。
ACTS|11|25|他又往 大數 去找 掃羅 ，
ACTS|11|26|找著了，就帶他到 安提阿 去。他們足有一年和教會一同聚集，教導了許多人。門徒稱為「基督徒」是從 安提阿 開始的。
ACTS|11|27|當那些日子，有幾位先知從 耶路撒冷 下到 安提阿 。
ACTS|11|28|內中有一位，名叫 亞迦布 ，站起來，藉著聖靈指示普天下將有大饑荒；這事在 克勞第 年間果然實現了。
ACTS|11|29|於是門徒決定，照各人的力量捐錢，送去供給住在 猶太 的弟兄。
ACTS|11|30|他們就這樣做了，託 巴拿巴 和 掃羅 的手送到眾長老那裏。
ACTS|12|1|約在那時候， 希律 王下手苦待教會中的一些人，
ACTS|12|2|用刀殺了 約翰 的哥哥 雅各 。
ACTS|12|3|他見 猶太 人喜歡這事，也去拿住 彼得 。那時候正是除酵節期間。
ACTS|12|4|希律 捉了 彼得 ，押在監裏，交給四班士兵看守，每班四個人，企圖要在逾越節後把他提出來，當著百姓辦他。
ACTS|12|5|於是 彼得 被囚在監裏，教會卻為他切切禱告上帝。
ACTS|12|6|希律 將要提他出來的前一夜， 彼得 被兩條鐵鏈鎖著，睡在兩個士兵當中；門前還有警衛看守。
ACTS|12|7|忽然，有主的一個使者顯現，牢房裏有光照耀；天使拍 彼得 的肋旁，叫醒了他，說：「快起來！」鐵鏈就從他手上脫落下來。
ACTS|12|8|天使對他說：「束上腰帶，穿上鞋子。」他就照著做了。天使又對他說：「披上外衣，跟我來。」
ACTS|12|9|彼得 就出來跟著他走，不知道天使所做是真的，以為見了異象。
ACTS|12|10|他們經過了第一層和第二層監牢，就來到往城內的鐵門，那門就自動給他們開了。他們出來，走過一條街，忽然天使離開他去了。
ACTS|12|11|彼得 清醒過來，說：「現在我真知道主差遣他的使者，救我脫離 希律 的手，和 猶太 人所期待的一切。」
ACTS|12|12|他明白了，就到那稱為 馬可 的 約翰 的母親 馬利亞 家去，在那裏已有好些人聚集禱告。
ACTS|12|13|彼得 敲外門時，有一個使女，名叫 羅大 ，出來應門，
ACTS|12|14|認出是 彼得 的聲音，歡喜得顧不了開門，就跑進去報信，說 彼得 站在門外。
ACTS|12|15|他們對她說：「你瘋了！」使女堅持真有其事。他們說：「那是他的天使。」
ACTS|12|16|彼得 不停地敲門；他們開了門，一見是他，就很驚奇。
ACTS|12|17|彼得 做個手勢，要他們不作聲，就告訴他們主怎樣領他出監；又說：「你們要把這些事告訴 雅各 和眾弟兄。」然後，他離開往別處去了。
ACTS|12|18|到了天亮，士兵中起了不少騷動，不知道 彼得 到哪裏去了。
ACTS|12|19|希律 找他，找不著，就審問警衛，下令帶走他們處死。後來 希律 離開 猶太 ，下 凱撒利亞 去，住在那裏。
ACTS|12|20|希律 向 推羅 和 西頓 的人發怒。他們那一帶地方是從王的土地供應糧食的，因此就託了王的內侍大臣 伯拉斯都 的情，一心來求和。
ACTS|12|21|希律 在所定的日子，穿上朝服，坐在位上，對他們演講。
ACTS|12|22|民眾一直喊著：「這是神明的聲音，不是人的聲音。」
ACTS|12|23|希律 不歸榮耀給上帝，所以主的使者立刻擊打他，他被蟲咬，就斷了氣。
ACTS|12|24|上帝的道日見興旺，越發廣傳。
ACTS|12|25|巴拿巴 和 掃羅 完成了供給的事，就回到 耶路撒冷 ，帶著稱為 馬可 的 約翰 同去。
ACTS|13|1|在 安提阿 的教會中，有幾位先知和教師，就是 巴拿巴 和稱為 尼結 的 西面 、 古利奈 人 路求 ，與 希律 分封王一起長大的 馬念 ，和 掃羅 。
ACTS|13|2|他們在事奉主和禁食的時候，聖靈說：「要為我分派 巴拿巴 和 掃羅 去做我召他們做的工作。」
ACTS|13|3|於是他們禁食禱告後，給 巴拿巴 和 掃羅 按手，然後派遣他們走了。
ACTS|13|4|他們既蒙聖靈差遣，就下到 西流基 ，從那裏坐船往 塞浦路斯 去，
ACTS|13|5|到了 撒拉米 ，就在 猶太 人各會堂裏宣講上帝的道，也有 約翰 作他們的幫手。
ACTS|13|6|他們走遍全島，直到 帕弗 ，在那裏遇見一個術士— 猶太 人的假先知，名叫 巴耶穌 。
ACTS|13|7|這人常和 士求．保羅 省長在一起。 士求．保羅 是個通達人，他請 巴拿巴 和 掃羅 來，要聽上帝的道。
ACTS|13|8|只是術士 以呂馬 (他的名字翻出來就是行法術的意思)敵對使徒，設法使省長遠離這信仰。
ACTS|13|9|掃羅 ，又名 保羅 ，被聖靈充滿，定睛看他，
ACTS|13|10|說：「你這充滿各樣詭詐奸惡，魔鬼的兒子，一切正義的仇敵，你還不停止扭曲主的正道嗎？
ACTS|13|11|現在你看，主的手臨到你身上，你會瞎眼，暫時看不見日光。」立刻迷濛和黑暗籠罩著他，他到處摸索，求人拉著手領他。
ACTS|13|12|省長看見所發生的事就信了，因對主的教導感到驚奇。
ACTS|13|13|保羅 和他的同伴從 帕弗 開船，來到 旁非利亞 的 別加 ， 約翰 卻離開他們，回 耶路撒冷 去了。
ACTS|13|14|他們從 別加 往前行，來到 彼西底 的 安提阿 。在安息日，他們進了會堂就坐下。
ACTS|13|15|在讀完了律法和先知的書，會堂主管們叫人過去，對他們說：「二位弟兄，你們若有甚麼勸勉眾人的話，請說。」
ACTS|13|16|保羅 就站起來，做個手勢，說：「諸位 以色列 人和一切敬畏上帝的人，請聽。
ACTS|13|17|這 以色列 民的上帝揀選了我們的祖宗，當百姓寄居 埃及 的時候抬舉他們，用大能的手領他們從那地出來。
ACTS|13|18|他在曠野容忍 他們，約有四十年。
ACTS|13|19|他消滅了 迦南 地七族的人後，把那地分給他們為業，
ACTS|13|20|約有四百五十年。此後 ，他給他們設立士師，直到 撒母耳 先知的時候。
ACTS|13|21|從那時起，他們要求立一個王，上帝就將 便雅憫 支派中 基士 的兒子 掃羅 給他們作王，共四十年。
ACTS|13|22|他廢了 掃羅 之後，就興起 大衛 作他們的王，又為他作見證說：『我尋得 耶西 的兒子 大衛 ，他是合我心意的人，他要遵行我一切的旨意。』
ACTS|13|23|從這人的後裔中，上帝已經照著所應許的為 以色列 人興起一位救主，就是耶穌。
ACTS|13|24|在他沒有出來以前， 約翰 已向 以色列 全民宣講悔改的洗禮。
ACTS|13|25|約翰 快走完他的人生路程時，說：『你們以為我是誰？我不是 ；但是有一位在我以後來的，我就是解他腳上的鞋帶也不配。』
ACTS|13|26|「諸位弟兄— 亞伯拉罕 的子孫和你們中間敬畏上帝的人哪，這救世的道是傳給我們的。
ACTS|13|27|耶路撒冷 的居民和他們的官長，因為不認識這基督，也不明白每安息日所讀的先知的書，把他定了死罪，正應驗了先知的預言。
ACTS|13|28|雖然他們查不出他有該死的罪狀，還是要求 彼拉多 把他殺了。
ACTS|13|29|他們既實現了經上指著他所記的一切話，就從木頭上把他取下來，放在墳墓裏。
ACTS|13|30|上帝卻使他從死人中復活。
ACTS|13|31|有許多日子，他向那些從 加利利 同他上 耶路撒冷 的人顯現，這些人如今在民間成為他的見證人。
ACTS|13|32|我們報好信息給你們，就是那應許祖宗的話，
ACTS|13|33|上帝已經向我們這些作他們兒女的 應驗，使耶穌復活了。正如《詩篇》第二篇上記著： 『你是我的兒子， 我今日生了你。』
ACTS|13|34|論到上帝使他從死人中復活，不再歸於朽壞，他曾這樣說： 『我必將所應許 大衛 那聖潔、 可靠的恩典賜給你們。』
ACTS|13|35|所以他也在另一篇說： 『你必不讓你的聖者見朽壞。』
ACTS|13|36|大衛 在世的時候，遵行了上帝的旨意就長眠了 ，歸到他祖宗那裏，已見朽壞；
ACTS|13|37|惟獨上帝使他復活的那一位，他並未見朽壞。
ACTS|13|38|所以弟兄們，你們當知道：赦罪的道是由這人傳給你們的，
ACTS|13|39|你們靠 摩西 的律法在不得稱義的一切事上，每一個信靠這位耶穌的都得稱義了。
ACTS|13|40|所以，你們要小心，免得先知書上所說的臨到你們：
ACTS|13|41|『要觀看，你們這些藐視的人， 要驚訝，要滅亡， 因為在你們的日子，我行一件事， 雖有人告訴你們，你們總是不信。』」
ACTS|13|42|他們走出會堂的時候，眾人請他們在下一個安息日再講這些話給他們聽。
ACTS|13|43|散會以後，有許多 猶太 人和敬虔的皈依 猶太 教的人跟從了 保羅 和 巴拿巴 。二人對他們講話，勸他們務要恆久倚靠上帝的恩典。
ACTS|13|44|到下一個安息日，全城的人幾乎都聚集起來，要聽主的道 。
ACTS|13|45|但 猶太 人看見這麼多的人，就滿心嫉妒，辯駁 保羅 所說的話，並且毀謗他。
ACTS|13|46|於是 保羅 和 巴拿巴 放膽說：「上帝的道本應先傳給你們；只因你們棄絕這道，斷定自己不配得永生，我們就轉向外邦人。
ACTS|13|47|因為主曾這樣吩咐我們： 『我已經立你作萬邦之光， 使你施行我的救恩，直到地極。』」
ACTS|13|48|外邦人聽見這話很歡喜，讚美主的道，凡被指定得永生的人都信了。
ACTS|13|49|於是主的道傳遍了那一帶地方。
ACTS|13|50|但 猶太 人挑唆虔敬尊貴的婦女和城內有名望的人，迫害 保羅 和 巴拿巴 ，把他們趕出境外。
ACTS|13|51|二人對著眾人跺掉腳上的塵土，然後往 以哥念 去了。
ACTS|13|52|門徒滿心喜樂，又被聖靈充滿。
ACTS|14|1|同樣的事也發生在 以哥念 。 保羅 和 巴拿巴 進了 猶太 人的會堂，在那裏講道，所以有很多 猶太 人和 希臘 人都信了。
ACTS|14|2|但那不順從的 猶太 人煽動外邦人，使他們心裏仇恨弟兄。
ACTS|14|3|二人在那裏住了好些日子，倚靠主放膽講道，主藉他們的手施行神蹟奇事，證明他恩惠的道。
ACTS|14|4|城裏的眾人卻分裂了：有依附 猶太 人的，有依附使徒的。
ACTS|14|5|那時，外邦人、 猶太 人和他們的官長，一齊擁上來，要凌辱使徒，用石頭打他們。
ACTS|14|6|使徒知道了，就逃到 呂高尼 的 路司得 和 特庇 兩個城，以及周圍地方去，
ACTS|14|7|在那裏繼續傳福音。
ACTS|14|8|路司得城 裏有一個兩腳無力的人，他從母腹裏就是瘸腿的，老是坐著，從來沒有走過。
ACTS|14|9|他聽 保羅 講道； 保羅 定睛看他，見他有信心，可得痊癒，
ACTS|14|10|就大聲說：「起來！兩腳站直。」那人就跳起來，開始行走。
ACTS|14|11|眾人看見 保羅 所做的事，就用 呂高尼 話大聲說：「有神明藉著人形降臨在我們中間了。」
ACTS|14|12|於是他們稱 巴拿巴 為 宙斯 ，稱 保羅 為 希耳米 ，因為他總是帶頭說話。
ACTS|14|13|城外有 宙斯 廟的祭司牽著牛，拿著花環，來到門前，要同眾人一起獻祭。
ACTS|14|14|巴拿巴 和 保羅 二位使徒聽見，就撕開衣裳，跳進眾人中間，喊著：
ACTS|14|15|「諸位，為甚麼做這些事呢？我們也是人，性情和你們一樣。我們傳福音給你們，是要你們離棄這些虛妄的事，歸向那創造天、地、海和其中萬物的永生的上帝。
ACTS|14|16|他在從前的世代，任憑萬國各行其道；
ACTS|14|17|然而他未嘗不為自己留下證據來，就如常行善事，從天降雨，賞賜豐年，使你們飲食飽足，滿心喜樂。」
ACTS|14|18|二人說了這些話，總算攔住眾人不獻祭給他們。
ACTS|14|19|但有些 猶太 人，從 安提阿 和 以哥念 來，挑唆眾人，並且用石頭打 保羅 ，以為他死了，就把他拖到城外。
ACTS|14|20|當門徒圍著他的時候，他站了起來，走進城去。第二天， 保羅 同 巴拿巴 往 特庇 去。
ACTS|14|21|保羅 和 巴拿巴 對那城裏的人傳了福音，使好些人成為門徒後，又回 路司得 、 以哥念 、 安提阿 去，
ACTS|14|22|堅固門徒的心，勸他們持守他們的信仰，說：「我們進入上帝的國，必須經歷許多艱難。」
ACTS|14|23|二人在各教會中選立了長老，禁食禱告後，把他們交託給他們所信的主。
ACTS|14|24|二人經過 彼西底 來到 旁非利亞 ，
ACTS|14|25|在 別加 講了道，就下 亞大利 去，
ACTS|14|26|從那裏坐船回 安提阿 去。當初，眾人就在這地方，把他們交託在上帝的恩典中，要完成現在所做的工。
ACTS|14|27|他們一到那裏，就聚集了會眾，述說上帝藉他們所行的一切事，並且上帝怎樣為外邦人開了信道的門。
ACTS|14|28|二人在那裏同門徒住了一段日子。
ACTS|15|1|有幾個人從 猶太 下來，教導弟兄們說：「你們若不按照 摩西 的規矩受割禮，不能得救。」
ACTS|15|2|保羅 和 巴拿巴 跟他們發生了激烈的爭執和辯論；大家就決定指派 保羅 、 巴拿巴 和本會的幾個人，為所辯論的事上 耶路撒冷 去見使徒和長老。
ACTS|15|3|於是教會為他們送行。他們經過 腓尼基 、 撒瑪利亞 ，沿途敘說外邦人歸主的事，使眾弟兄都非常歡喜。
ACTS|15|4|他們到了 耶路撒冷 ，教會、使徒和長老都接待他們，他們就述說上帝同他們所做的一切事。
ACTS|15|5|惟有幾個法利賽派的信徒起來，說：「必須給外邦人行割禮，吩咐他們遵守 摩西 的律法。」
ACTS|15|6|使徒和長老聚集商議這事。
ACTS|15|7|辯論了許久後， 彼得 站起來，對他們說：「諸位弟兄，你們知道上帝早已在你們中間揀選了我，讓外邦人從我口中得聽福音之道，而且相信。
ACTS|15|8|知道人心的上帝也為他們作了見證，賜聖靈給他們，正如給我們一樣；
ACTS|15|9|又藉著信潔淨了他們的心，他們和我們之間並沒有甚麼分別。
ACTS|15|10|現在你們為甚麼試探上帝，要把我們祖宗和我們所不能負的軛放在門徒的頸項上呢？
ACTS|15|11|相反地，我們相信，我們得救是因主耶穌的恩典，和他們一樣。」
ACTS|15|12|眾人都默默無聲，聽 巴拿巴 和 保羅 述說上帝藉著他們在外邦人中所行的神蹟和奇事。
ACTS|15|13|他們講完了， 雅各 回答說：「諸位弟兄，請聽我說。
ACTS|15|14|剛才 西門 述說上帝當初怎樣眷顧外邦人，從他們中間選取人民歸於自己的名下；
ACTS|15|15|眾先知的話也與這意思相符合。
ACTS|15|16|正如經上所寫的： 『此後，我要回來， 重新修造 大衛 倒塌了的帳幕， 從廢墟中重新修造， 把它建立起來，
ACTS|15|17|使剩餘的人， 就是凡稱我名的外邦人， 都尋求主。 這話是自古以來顯明這些事的主說的。』
ACTS|15|18|
ACTS|15|19|所以，我的意見是不可難為那歸向上帝的外邦人；
ACTS|15|20|但是要寫信吩咐他們禁戒偶像所玷污的東西、血和勒死的牲畜 ，禁戒淫亂。
ACTS|15|21|因為歷代以來， 摩西 的書在各城都有人宣講，每逢安息日，也在會堂裏誦讀。」
ACTS|15|22|那時，使徒、長老和全教會認為應從他們中間揀選人，差他們和 保羅 、 巴拿巴 一同到 安提阿 去，所揀選的就是稱為 巴撒巴 的 猶大 和 西拉 。這二人在弟兄中是領袖。
ACTS|15|23|他們帶去的信說：「使徒和作長老的弟兄們向 安提阿 、 敘利亞 、 基利家 外邦眾弟兄問安。
ACTS|15|24|我們聽說，有幾個人從我們這裏出去 ，用一些話騷擾你們，使你們的心困惑， 其實我們並沒有吩咐他們。
ACTS|15|25|我們認為，既然我們同心定意，就揀選幾個人，派他們同我們所親愛的 巴拿巴 和 保羅 到你們那裏去。
ACTS|15|26|這二人曾為我主耶穌基督的名不顧自己的性命。
ACTS|15|27|所以我們派 猶大 和 西拉 去，他們也會親口述說這些事。
ACTS|15|28|因為聖靈和我們決定除了這幾件重要的事，不將別的重擔放在你們身上，
ACTS|15|29|就是禁戒偶像所玷污的東西、血和勒死的牲畜，禁戒淫亂。這幾件你們若能自己禁戒就好了。祝你們安康！」
ACTS|15|30|他們既奉了差遣就下 安提阿 去，聚集會眾，把書信交給他們。
ACTS|15|31|眾人念了，因為信上鼓勵的話而感到欣慰。
ACTS|15|32|猶大 和 西拉 自己也是先知，就用許多話勸勉弟兄，堅固他們。
ACTS|15|33|二人住了些日子，弟兄們打發他們平平安安地回到差遣他們的人那裏去。
ACTS|15|34|
ACTS|15|35|但 保羅 和 巴拿巴 仍留在 安提阿 ，和許多別的人一同教導，並傳揚主的道。
ACTS|15|36|過了些日子， 保羅 對 巴拿巴 說：「讓我們回到從前宣揚主道的各城，看看弟兄們的情況如何。」
ACTS|15|37|巴拿巴 有意要帶稱為 馬可 的 約翰 同去；
ACTS|15|38|但 保羅 認為不宜帶他去，因為 馬可 從前在 旁非利亞 離開他們，不和他們一起工作。
ACTS|15|39|於是二人起了爭執，甚至彼此分手。 巴拿巴 帶著 馬可 ，坐船往 塞浦路斯 去；
ACTS|15|40|保羅 則揀選了 西拉 ，也出發了，蒙弟兄們把他交於主的恩典中。
ACTS|15|41|他就走遍了 敘利亞 、 基利家 ，堅固眾教會。
ACTS|16|1|後來， 保羅 來到 特庇 ，又到 路司得 。在那裏有一個門徒，名叫 提摩太 ，是信主的 猶太 婦人的兒子，他父親卻是 希臘 人。
ACTS|16|2|路司得 和 以哥念 的弟兄都稱讚他。
ACTS|16|3|保羅 要帶他同去，只因那些地方的 猶太 人都知道他父親是 希臘 人，就給他行了割禮。
ACTS|16|4|他們經過各城，把 耶路撒冷 使徒和長老所決定的規條交給門徒遵守。
ACTS|16|5|於是眾教會信心越發堅固，人數天天增加。
ACTS|16|6|因為聖靈禁止他們在 亞細亞 講道，他們就經過 弗呂家 、 加拉太 一帶地方。
ACTS|16|7|到了 每西亞 的邊界，他們想要往 庇推尼 去，耶穌的靈卻不許。
ACTS|16|8|他們就越過 每西亞 ，下 特羅亞 去。
ACTS|16|9|夜間，有異象向 保羅 顯現。有一個 馬其頓 人站著求他說：「請你過來，到 馬其頓 來幫助我們！」
ACTS|16|10|保羅 既看見這異象，我們就立即設法往 馬其頓 去，認為上帝呼召我們傳福音給那裏的人。
ACTS|16|11|我們從 特羅亞 開船，直行駛到 撒摩特喇 ，第二天到了 尼亞坡里 ；
ACTS|16|12|從那裏來到 腓立比 ，就是 馬其頓 這一帶的一個重要城市 ，也是 羅馬 的駐防城。我們在這城裏住了幾天。
ACTS|16|13|在安息日，我們出城門，到了河邊，知道那裏有一個禱告的地方 ，我們就坐下來對那些聚會的婦女講道。
ACTS|16|14|有一個賣紫色布的婦人，名叫 呂底亞 ，是 推雅推喇城 的人，素來敬拜上帝。她在聽著，主就開導她的心，使她留心聽 保羅 所講的話。
ACTS|16|15|她和她一家都領了洗，就求我們說：「你們若以為我是真心信主的 ，請到我家裏來住。」於是她堅決請我們留下。
ACTS|16|16|後來，我們往那禱告的地方去時，有一個被占卜的靈附身的使女迎面走來，她使用法術使她的主人們發了大財。
ACTS|16|17|她跟隨 保羅 和我們，喊著說：「這些人是至高上帝的僕人，對你們傳講救人的道路。」
ACTS|16|18|她一連好幾天這樣喊叫， 保羅 就心中厭煩，轉身對那靈說：「我奉耶穌基督的名吩咐你從她身上出來！」那靈立刻出來了。
ACTS|16|19|使女的主人們見發財的指望沒有了，就揪住 保羅 和 西拉 ，拉他們到市上去見官；
ACTS|16|20|又帶他們到行政官長們面前，說：「這些騷擾我們城的，他們是 猶太 人，
ACTS|16|21|竟傳佈我們 羅馬 人所不可接受、不可遵守的規矩。」
ACTS|16|22|群眾就一齊起來攻擊他們。官長們吩咐撕開他們的衣裳，用棍子打；
ACTS|16|23|打了許多棍，就把他們下在監裏，囑咐獄警嚴緊看守。
ACTS|16|24|獄警領了這樣的命令，就把他們下在內監，兩腳拴在木架上。
ACTS|16|25|約在半夜， 保羅 和 西拉 正在禱告，唱詩讚美上帝，眾囚犯也側耳聽著的時候，
ACTS|16|26|忽然，地大震動，甚至監牢的地基都搖動了，監門立刻全開，眾囚犯的鎖鏈也都解開了。
ACTS|16|27|獄警一醒，看見監門全開，以為囚犯已經逃走，就拔刀要自殺。
ACTS|16|28|保羅 大聲呼叫：「不要傷害自己！我們都在這裏。」
ACTS|16|29|獄警叫人拿燈來，就衝進去，戰戰兢兢地俯伏在 保羅 和 西拉 面前。
ACTS|16|30|然後獄警領他們出來，說：「二位先生，我必須做甚麼才可以得救？」
ACTS|16|31|他們說：「當信主耶穌，你和你一家都必得救 。」
ACTS|16|32|他們就把主的道講給他和他全家的人聽。
ACTS|16|33|當夜，就在那時候，獄警把他們帶去，洗他們的傷；他和他所有的家人立刻都受了洗。
ACTS|16|34|於是獄警領他們上自己的家裏去，給他們擺上飯。他和全家的人，因為信了上帝，都滿心喜樂。
ACTS|16|35|到了天亮，官長們打發差役來，說：「釋放那兩個人吧。」
ACTS|16|36|獄警就把這些話告訴 保羅 ：「官長們打發人來，要釋放你們，現在可以出監，平平安安去吧。」
ACTS|16|37|保羅 卻說：「我們是 羅馬 人，並沒有定罪，他們竟在公眾面前打了我們，又把我們下在監裏；現在要私下趕我們出去嗎？這不行！叫他們自己來領我們出去吧！」
ACTS|16|38|差役把這些話回稟官長們；官長們聽見他們是 羅馬 人，就害怕了，
ACTS|16|39|於是來勸他們，領他們出來，請他們離開那城。
ACTS|16|40|二人出了監牢，往 呂底亞 家裏去，見了弟兄們，勸慰他們一番，就離開了。
ACTS|17|1|保羅 和 西拉 經過 暗妃坡里 、 亞波羅尼亞 ，來到 帖撒羅尼迦 ，在那裏有 猶太 人的會堂。
ACTS|17|2|保羅 照他素常的規矩進去，一連三個安息日，根據聖經與他們辯論，
ACTS|17|3|講解和說明基督必須受害，從死人中復活；又說：「我所傳給你們的這位耶穌就是基督。」
ACTS|17|4|他們中間有些人聽了勸，就跟從 保羅 和 西拉 ，還有許多虔敬的 希臘 人，尊貴的婦女也不少。
ACTS|17|5|但不信的 猶太 人心裏嫉妒，聚集了些市井流氓，搭夥成群，煽動全城的人闖進 耶孫 的家，要把 保羅 和 西拉 帶到民眾那裏。
ACTS|17|6|那些人找不著他們，就把 耶孫 和幾個弟兄拉到地方官那裏，喊叫著：「這些攪亂天下的人也到這裏來了，
ACTS|17|7|耶孫 竟收留他們。這些人都違背凱撒的命令，說另有一個王耶穌。」
ACTS|17|8|眾人和地方官聽見這些話，就惶恐了，
ACTS|17|9|於是收了 耶孫 和其餘的人的保證金後，釋放了他們。
ACTS|17|10|當夜，弟兄們立刻送 保羅 和 西拉 往 庇哩亞 去；二人到了，就進入 猶太 人的會堂。
ACTS|17|11|這地方的 猶太 人比 帖撒羅尼迦 的人開明，熱心領受這道，天天查考聖經，要知道這道是否真實。
ACTS|17|12|所以，他們中間有許多信了，又有 希臘 的尊貴婦人，男人也不少。
ACTS|17|13|但 帖撒羅尼迦 的 猶太 人知道 保羅 又在 庇哩亞 傳上帝的道，就往那裏去，煽動挑撥群眾。
ACTS|17|14|於是，弟兄們立刻送 保羅 到海邊去， 西拉 和 提摩太 卻仍留在 庇哩亞 。
ACTS|17|15|護送 保羅 的人帶他到了 雅典 ，他們領了 保羅 的命令，叫 西拉 和 提摩太 趕快到他那裏來，然後回去了。
ACTS|17|16|保羅 在 雅典 等候他們的時候，看見滿城都是偶像，就心裏非常難過。
ACTS|17|17|於是他在會堂裏與 猶太 人和虔敬的人，以及每日在市場上所遇見的人辯論。
ACTS|17|18|還有 伊壁鳩魯 和 斯多亞 兩派的哲學家也與他爭辯。有的說：「這胡言亂語的要說甚麼？」有的說：「他似乎是宣傳外邦鬼神的。」這是因 保羅 傳講耶穌與復活的福音。
ACTS|17|19|他們就把他帶到 亞略巴古 ，說：「你所講的這新學說，我們也可以知道嗎？
ACTS|17|20|因為你有些奇怪的事傳到我們耳中，我們想知道這些事是甚麼意思。」
ACTS|17|21|原來所有的 雅典 人和居住在那裏的外國人都無暇管別的事，只是談談或聽聽新聞。
ACTS|17|22|保羅 站在 亞略巴古 當中，說：「諸位 雅典 人！我看你們凡事很敬畏鬼神。
ACTS|17|23|我到處走走的時候，仔細觀察你們所敬拜的，發現一座壇，上面寫著『獻給未識之神明』。你們所不認識而敬拜的，我現在向你們宣告：
ACTS|17|24|他是創造宇宙和其中萬物的上帝；他既是天地的主，就不住在人手所造的殿宇裏，
ACTS|17|25|也不用人手去服侍，好像缺少甚麼似的；自己倒將生命、氣息、萬物賜給萬人。
ACTS|17|26|他從一人 造出萬族，居住在全地面上，並且預先定準他們的年限和所住的疆界，
ACTS|17|27|為要使他們尋求上帝，或者可以揣摩而找到他，其實他離我們各人不遠。
ACTS|17|28|我們生活、行動、存在都在於他。就如你們的詩人也有人說：『我們也是他所生的。』
ACTS|17|29|既然我們是上帝所生的，就不應該以為上帝的神性像人用手藝和心思所雕刻的金、銀、石像一般。
ACTS|17|30|世人蒙昧無知的時候，上帝並不追究，如今卻吩咐各處的人都要悔改。
ACTS|17|31|因為他已經定了日子，要藉著他所設立的人按公義審判天下，並且使他從死人中復活，給萬人作可信的憑據。」
ACTS|17|32|眾人聽見死人復活的話，就有人譏誚他；又有人說：「我們會再聽你講這事。」
ACTS|17|33|於是 保羅 從他們當中出去了。
ACTS|17|34|但有幾個人依附他，信了主，其中有 亞略巴古 的議員 丟尼修 ，和一個名叫 大馬哩 的婦人，還有幾個與他們一起的人。
ACTS|18|1|這些事以後， 保羅 離開 雅典 ，來到 哥林多 。
ACTS|18|2|他遇見一個生在 本都 的 猶太 人，名叫 亞居拉 。不久前，他帶著妻子 百基拉 從 意大利 來，因為 克勞第 命令所有的 猶太 人都離開 羅馬 。 保羅 去投靠他們。
ACTS|18|3|他們本是製造帳棚為業。 保羅 因與他們同業，就和他們同住，一同做工。
ACTS|18|4|每逢安息日， 保羅 在會堂裏辯論，勸導 猶太 人和 希臘 人。
ACTS|18|5|西拉 和 提摩太 從 馬其頓 來的時候， 保羅 正專心傳道，向 猶太 人證明耶穌是基督。
ACTS|18|6|當他們抗拒他、毀謗他的時候，他就抖掉衣裳的灰塵，對他們說：「你們的罪歸到你們自己的頭上，與我無干。從今以後，我要往外邦人那裏去。」
ACTS|18|7|於是他離開那裏，到了一個人的家裏，他名叫 提多．猶士都 ，是敬拜上帝的人，他的家靠近會堂。
ACTS|18|8|會堂的主管 基利司布 和全家都信了主，還有許多 哥林多 人聽了就信，而且受了洗。
ACTS|18|9|夜間，主在異象中對 保羅 說：「不要怕，只管講，不要沉默，
ACTS|18|10|有我與你同在，沒有人會下手害你，因為在這城裏有許多屬我的人。」
ACTS|18|11|保羅 在那裏住了一年六個月，將上帝的道教導他們。
ACTS|18|12|到 迦流 作 亞該亞 省長的時候， 猶太 人齊心起來攻擊 保羅 ，拉他到法庭，
ACTS|18|13|說：「這個人教唆人不按著律法敬拜上帝。」
ACTS|18|14|保羅 剛要開口， 迦流 對 猶太 人說：「你們這些 猶太 人哪！如果是為冤枉或奸惡的事，我理當耐性聽你們。
ACTS|18|15|既然你們所爭論的是關乎用字、名目和你們的律法，你們自己去辦吧！這樣的事我不願意審問。」
ACTS|18|16|於是，他把他們逐出法庭。
ACTS|18|17|眾人就揪住會堂的主管 所提尼 ，在法庭前打他。這些事 迦流 都不管。
ACTS|18|18|保羅 又住了好些日子，就辭別了弟兄，坐船到 敘利亞 去。 百基拉 、 亞居拉 和他同去。他因為許過願，就在 堅革哩 剃了頭髮。
ACTS|18|19|到了 以弗所 ， 保羅 就把他們留在那裏，自己進了會堂，和 猶太 人辯論。
ACTS|18|20|眾人請他多住些日子，他沒有答應，
ACTS|18|21|就辭別他們，說：「上帝若許可，我還要回到你們這裏來。」於是他上船離開 以弗所 。
ACTS|18|22|他在 凱撒利亞 下了船，上 耶路撒冷 去問候教會，隨後下 安提阿 去。
ACTS|18|23|他在那裏住了些日子，又離開了那裏，逐一經過 加拉太 和 弗呂家 各地方，堅固眾門徒。
ACTS|18|24|有一個生在 亞歷山大 的 猶太 人，名叫 亞波羅 ，來到 以弗所 ，他很有口才，很會講解聖經。
ACTS|18|25|這人已經在主的道路上受了訓練，心裏火熱，精確地講論和教導耶穌的事；可是他只知道 約翰 的洗禮。
ACTS|18|26|他開始在會堂裏放膽講道； 百基拉 、 亞居拉 聽見，就接他來，將上帝的道路 給他更精確地講解。
ACTS|18|27|他想要往 亞該亞 去，弟兄們就勉勵他，並寫信請門徒們接待他，他到了那裏，多多幫助那些蒙恩信主的人，
ACTS|18|28|因為他在公眾面前極力駁倒 猶太 人，引聖經證明耶穌是基督。
ACTS|19|1|亞波羅 在 哥林多 的時候， 保羅 經過了內陸地區，來到 以弗所 ，在那裏他遇見幾個門徒，
ACTS|19|2|問他們：「你們信的時候領受了聖靈沒有？」他們說：「沒有，我們連甚麼是聖靈都沒有聽過。」
ACTS|19|3|保羅 說：「這樣，你們受的是甚麼洗呢？」他們說：「是受了 約翰 的洗。」
ACTS|19|4|保羅 說：「 約翰 所施的是悔改的洗禮，他告訴百姓當信那在他以後要來的那位，就是耶穌。」
ACTS|19|5|他們聽見這話以後，就奉主耶穌的名受洗。
ACTS|19|6|保羅 給他們按手，聖靈就降在他們身上，他們開始說方言 和說預言。
ACTS|19|7|他們約有十二個人。
ACTS|19|8|保羅 進會堂，一連三個月放膽講道，辯論上帝國的事，勸導眾人。
ACTS|19|9|後來，有些人心裏剛硬不信，在眾人面前毀謗這道； 保羅 就離開他們，也叫門徒與他們分開，就在 推喇奴 的講堂天天辯論。
ACTS|19|10|這樣有兩年之久，使一切住在 亞細亞 的，無論是 猶太 人是 希臘 人，都聽見主的道。
ACTS|19|11|上帝藉 保羅 的手行了些奇異的神蹟，
ACTS|19|12|甚至有人從 保羅 身上拿走手巾或圍裙放在病人身上，病就消除了，邪靈也出去了。
ACTS|19|13|那時，有幾個巡迴各處念咒趕鬼的 猶太 人，擅自利用主耶穌的名，向那些被邪靈所附的人說：「我奉 保羅 所傳的耶穌命令你們出來！」
ACTS|19|14|做這事的是 猶太 祭司長 士基瓦 的七個兒子。
ACTS|19|15|但邪靈回答他們：「耶穌我知道， 保羅 我也認識，你們卻是誰呢？」
ACTS|19|16|被邪靈所附的人就撲到他們身上，制伏他們，勝過他們，使他們赤著身子，受了傷，從那房子裏逃出去了。
ACTS|19|17|凡住在 以弗所 的，無論是 猶太 人是 希臘 人，都知道這件事，也都懼怕；主耶穌的名從此就更被尊為大了。
ACTS|19|18|許多已經信的人來承認並公開自己所行的事。
ACTS|19|19|又有許多平素行邪術的人把他們的書都拿來，堆積在眾人面前焚燒。他們計算書價，得知共值五萬塊銀錢。
ACTS|19|20|這樣，主的道大大興旺，而且普遍傳開了。
ACTS|19|21|這些事過後， 保羅 心裏決定要經過 馬其頓 、 亞該亞 ，就往 耶路撒冷 去。他說：「我到了那裏以後，也必須到 羅馬 去看看。」
ACTS|19|22|於是他差遣兩個助手 提摩太 和 以拉都 往 馬其頓 去，自己暫時留在 亞細亞 。
ACTS|19|23|那時，因這道路而起的騷動不小。
ACTS|19|24|有一個銀匠，名叫 底米丟 ，是製造 亞底米 神銀龕的，他使從事這手藝的人生意發達。
ACTS|19|25|他聚集他們和同行的工人，說：「諸位，你們知道我們是倚靠這生意發財的。
ACTS|19|26|你們看到，也聽見這 保羅 不但在 以弗所 ，也幾乎在 亞細亞 全地，引誘迷惑了許多人，說：『人手所做的不是神明。』
ACTS|19|27|這樣，不僅我們這行業陷入被藐視的危險，就是大女神 亞底米 的廟也要被人輕看，連 亞細亞 全地和普天下所敬拜的女神的威望也受損害了。」
ACTS|19|28|眾人聽見，就怒氣沖沖，喊著說：「大哉， 以弗所 人的 亞底米 ！」
ACTS|19|29|於是滿城都騷動起來。眾人抓住與 保羅 同行的 馬其頓 人 該猶 和 亞里達古 ，齊心衝進劇場。
ACTS|19|30|保羅 想要進到民眾那裏，門徒卻不許他去。
ACTS|19|31|連 亞細亞 的幾位官員，是 保羅 的朋友，也打發人來勸他不要冒險到劇場裏去。
ACTS|19|32|聚集的人亂成一團，有的喊這個，有的喊那個，大半不知道為了甚麼聚集。
ACTS|19|33|猶太 人把 亞歷山大 推出去，人群中有人慫恿他，他就做手勢，要向民眾申訴。
ACTS|19|34|但他們一認出他是 猶太 人，大家就異口同聲喊著：「大哉， 以弗所 人的 亞底米 ！」約喊了兩小時。
ACTS|19|35|城裏的書記官安撫了群眾後，說：「 以弗所 人哪，誰不知道 以弗所 人的城是看守大 亞底米 的廟和從 宙斯 那裏落下來的像的守護者呢？
ACTS|19|36|既然這些事是駁不倒的，你們就要安靜下來，不可妄動。
ACTS|19|37|你們把這些人帶來，他們並沒有偷竊廟中之物，也沒有褻瀆我們的女神。
ACTS|19|38|如果 底米丟 和他同行的手藝人有控告的事，自有公堂，也有省長，他們可以彼此控告。
ACTS|19|39|你們若有別的事請求，可以在合法的集會裏解決。
ACTS|19|40|今日的擾亂本是無緣無故的，有被控告的危險。這次的騷動，我們也說不出理由來。」
ACTS|19|41|他說完這些話，就叫眾人散會。
ACTS|20|1|騷亂平定以後， 保羅 請門徒來，勸勉了他們，就辭別他們，往 馬其頓 去。
ACTS|20|2|他走遍那一帶地方，用許多話勸勉門徒，然後來到 希臘 ，
ACTS|20|3|在那裏住了三個月。他快要坐船往 敘利亞 去的時候， 猶太 人設計害他，他就決定從 馬其頓 回去。
ACTS|20|4|同他到 亞細亞 去的，有 庇哩亞 人 畢羅斯 的兒子 所巴特 ， 帖撒羅尼迦 人 亞里達古 和 西公都 ，還有 特庇 人 該猶 和 提摩太 ，又有 亞細亞 人 推基古 和 特羅非摩 。
ACTS|20|5|這些人先走，在 特羅亞 等候我們。
ACTS|20|6|過了除酵節的日子，我們從 腓立比 開船，五天以後到了 特羅亞 ，和他們相會，在那裏住了七天。
ACTS|20|7|七日的第一日，我們聚會擘餅的時候， 保羅 因次日要起行，就為他們講道，直講到半夜。
ACTS|20|8|我們聚會的那座樓上有好些燈火。
ACTS|20|9|有一個少年，名叫 猶推古 ，坐在窗口上，沉沉入睡。 保羅 講了多時，少年睡熟了，從三層樓上掉下去，扶起來時已經死了。
ACTS|20|10|保羅 下去，伏在他身上，抱著他，說：「你們不要慌亂，他還有氣呢！」
ACTS|20|11|保羅 又上樓去，擘餅，吃了，再講了許久，直到天亮才離開。
ACTS|20|12|他們把那活過來的孩子帶走，大家得到很大的安慰。
ACTS|20|13|我們先上船，起航往 亞朔 去，想要在那裏接 保羅 ；因為他是這樣安排的，他自己本來打算要走陸路。
ACTS|20|14|他既在 亞朔 與我們相會，我們就接他上船，來到 米推利尼 。
ACTS|20|15|我們從那裏開船，第二天到了 基阿 的對岸；再下一天，在 撒摩 靠岸，又過了一天，到了 米利都 。
ACTS|20|16|因為 保羅 早已決定要越過 以弗所 ，免得在 亞細亞 耽延，他急忙前行，假如可能的話，在五旬節前能趕到 耶路撒冷 。
ACTS|20|17|保羅 從 米利都 打發人往 以弗所 去，請教會的長老來。
ACTS|20|18|他們來了， 保羅 對他們說：「你們自己知道，自從我到 亞細亞 的第一天，我怎樣跟你們相處，
ACTS|20|19|怎樣凡事謙卑，以眼淚服侍主，又因 猶太 人的謀害經歷試煉。
ACTS|20|20|你們也知道，凡對你們有益的，我沒有一樣隱瞞不說的，或在公眾面前，或在每一個人的家裏，我都教導你們，
ACTS|20|21|不論 猶太 人和 希臘 人，我都已證明他們當在上帝面前悔改，信靠我們的主耶穌。
ACTS|20|22|現在我被聖靈催迫 要往 耶路撒冷 去，雖然不知道在那裏會遭遇甚麼事，
ACTS|20|23|但知道聖靈在各城裏向我指證，說有捆鎖與患難等著我。
ACTS|20|24|我卻不以性命為念，只要走完我的路程，完成我從主耶穌所領受的職分，為上帝恩典的福音作見證。
ACTS|20|25|「我素常在你們中間到處傳講上帝的國；現在我知道，你們眾人以後不會再見到我的面了。
ACTS|20|26|所以我今日向你們作證，你們中間無論何人死亡，罪不在我。
ACTS|20|27|因為上帝一切的旨意，我並沒有退縮不傳給你們的。
ACTS|20|28|聖靈立你們作全群的監督，你們就當為自己謹慎，也為全群謹慎，牧養上帝 的教會，就是他用自己血所買來的 。
ACTS|20|29|我知道，在我離開以後必有兇暴的豺狼進入你們中間，不顧惜羊群。
ACTS|20|30|就是你們中間也必有人起來，說悖謬的話，要引誘門徒跟從他們。
ACTS|20|31|所以你們要警醒，記念我三年之久，晝夜不斷地流淚勸戒你們各人。
ACTS|20|32|現在我把你們交託給上帝和他恩惠的道；這道能建立你們，使你們和一切成聖的人同得基業。
ACTS|20|33|我未曾貪圖一個人的金、銀或衣服。
ACTS|20|34|你們自己知道，我靠兩隻手工作來供給我和同工的需用。
ACTS|20|35|我凡事給你們作榜樣，叫你們知道應當這樣勞苦，扶助軟弱的人，又當記念主耶穌的話，說：『施比受更為有福。』」
ACTS|20|36|保羅 說完了這些話，就和大家跪下來禱告。
ACTS|20|37|眾人痛哭，抱著 保羅 的頸項跟他親吻。
ACTS|20|38|叫他們最傷心的，就是他說「以後不會再見到我的面」那句話。於是他們送他上船去了。
ACTS|21|1|我們離別了眾人，就開船直航到 哥士 ，第二天到了 羅底 ，又從那裏到 帕大喇 。
ACTS|21|2|我們遇見一隻船要往 腓尼基 去，就上船起航。
ACTS|21|3|我們望見 塞浦路斯 ，就從南邊行過，往 敘利亞 去，在 推羅 上岸，因為船要在那裏卸貨。
ACTS|21|4|我們在那裏找到了一些門徒，就住了七天。他們藉著聖靈的感動，告訴 保羅 不要上 耶路撒冷 去。
ACTS|21|5|幾天之後，我們又出發前行。他們眾人同妻子兒女都送我們到城外，我們都跪在灘上禱告，彼此辭別。
ACTS|21|6|我們上了船，他們就回家去了。
ACTS|21|7|我們從 推羅 行完航程，來到了 多利買 ，問候那裏的弟兄，和他們同住了一天。
ACTS|21|8|第二天，我們離開那裏，來到 凱撒利亞 ，就進了傳福音的 腓利 家裏，和他同住；他是那七個執事裏的一個。
ACTS|21|9|他有四個女兒，都是未出嫁的，都會說預言。
ACTS|21|10|我們在那裏多住了好幾天，有一個先知，名叫 亞迦布 ，從 猶太 下來。
ACTS|21|11|他到了我們這裏，就拿 保羅 的腰帶，捆上自己的手腳，說：「聖靈這樣說：『 猶太 人在 耶路撒冷 要如此捆綁這腰帶的主人，把他交在外邦人手裏。』」
ACTS|21|12|我們聽見這些話，就跟當地的人苦勸 保羅 不要上 耶路撒冷 去。
ACTS|21|13|於是 保羅 回答：「你們為甚麼這樣痛哭，使我心碎呢？我為主耶穌的名，不但被人捆綁，就是死在 耶路撒冷 也是願意的。」
ACTS|21|14|既然 保羅 不聽勸，我們就住了口，只說：「願主的旨意成就。」
ACTS|21|15|過了這幾天，我們收拾行李上 耶路撒冷 去。
ACTS|21|16|有 凱撒利亞 的幾個門徒和我們同去，帶我們到一個早期的門徒 塞浦路斯 人 拿孫 的家裏，請我們與他同住。
ACTS|21|17|我們到了 耶路撒冷 ，弟兄們歡歡喜喜地接待我們。
ACTS|21|18|第二天， 保羅 同我們去見 雅各 ；所有的長老也都在場。
ACTS|21|19|保羅 向他們問安，然後將上帝用他在外邦人中所做的事奉，一一述說了。
ACTS|21|20|他們聽見了，就歸榮耀給上帝，對 保羅 說：「弟兄，你看 猶太 人中有數以萬計的信徒，而他們都是熱心於律法的人。
ACTS|21|21|他們曾聽見人說，你教導所有在外邦的 猶太 人離棄 摩西 ，對他們說，不要給孩子行割禮，也不要遵守規矩。
ACTS|21|22|眾人必聽見你來了，這可怎麼辦呢？
ACTS|21|23|你就照著我們的話做吧！我們這裏有四個人，都有願在身。
ACTS|21|24|你帶他們去，與他們一同行潔淨的禮，替他們繳納規費，讓他們得以剃頭。這樣，眾人就會知道，先前所聽見關於你的事都是假的；而且也知道，你自己為人循規蹈矩，遵行律法。
ACTS|21|25|至於信主的外邦人， 我們已經根據我們的決議寫信，叫他們要禁戒偶像所玷污的東西、血和勒死的牲畜，禁戒淫亂。」
ACTS|21|26|於是 保羅 帶著那四個人，第二天與他們一同行了潔淨禮，進了聖殿，報告潔淨期滿的日子，等候祭司為他們各人獻上祭物。
ACTS|21|27|那七日將完，從 亞細亞 來的 猶太 人看見 保羅 在聖殿裏，就煽動所有的群眾，下手拿住他，
ACTS|21|28|喊著：「 以色列 人哪，來幫忙！這就是在各處教導眾人糟蹋我們百姓、律法和這地方的人。不但如此，他還帶了 希臘 人進聖殿，污穢了這聖地。」
ACTS|21|29|這話是因他們曾看見 以弗所 人 特羅非摩 跟 保羅 一起在城裏，以為 保羅 帶他進了聖殿。
ACTS|21|30|於是全城都騷動，百姓一齊跑來，拿住 保羅 ，拉他出聖殿，殿門立刻都關了。
ACTS|21|31|他們正想要殺他，有人報信給營裏的千夫長，說 耶路撒冷 全城都亂了。
ACTS|21|32|千夫長立刻帶著士兵和幾個百夫長，跑下去到他們那裏。他們見了千夫長和士兵，就停下來不打 保羅 。
ACTS|21|33|於是千夫長上前拿住他，吩咐用兩條鐵鏈捆鎖，又問他是甚麼人，做了甚麼事。
ACTS|21|34|群眾中有的喊這個，有的喊那個；因為這樣亂嚷，千夫長無法知道實情，就下令將 保羅 帶進營樓去。
ACTS|21|35|保羅 一走上臺階，群眾擠得兇猛，士兵只得將 保羅 抬起來。
ACTS|21|36|一群人跟在後面，喊著：「除掉他！」
ACTS|21|37|保羅 快要被帶進營樓時，對千夫長說：「我可以對你說句話嗎？」千夫長說：「你懂得 希臘 話嗎？
ACTS|21|38|那你就不是從前作亂、帶領四千兇徒往曠野去的那 埃及 人了。」
ACTS|21|39|保羅 說：「我本是 猶太 人，生在 基利家 的 大數 ，並不是無名小城的公民。求你准我對百姓說話。」
ACTS|21|40|千夫長准了。 保羅 就站在臺階上，向百姓做了個手勢，要他們靜下來， 保羅 就用 希伯來 話對他們說：
ACTS|22|1|「諸位父老弟兄，請聽我現在對你們的申辯。」
ACTS|22|2|他們聽 保羅 說的是 希伯來 話，就更加安靜了。
ACTS|22|3|保羅 說：「我原是 猶太 人，生在 基利家 的 大數 ，但在這城裏長大，在 迦瑪列 門下按著我們祖宗嚴緊的律法受教，熱心事奉上帝，就如你們大家今日一樣。
ACTS|22|4|我也曾迫害信奉這道路的人，置他們於死地，無論男女都捆綁，關在監裏。
ACTS|22|5|這是大祭司和議會的眾長老都可以給我作證的。我又從他們那裏領了致弟兄們的書信，往 大馬士革 去，要把在那裏的信徒綁起來，帶到 耶路撒冷 受刑。」
ACTS|22|6|「當我走近 大馬士革 的時候，約在中午，忽然有一道大光從天上下來，照射在我周圍。
ACTS|22|7|我就仆倒在地，聽見有聲音對我說：『 掃羅 ！ 掃羅 ！你為甚麼迫害我？』
ACTS|22|8|我回答：『主啊！你是誰？』他對我說：『我就是你所迫害的 拿撒勒 人耶穌。』
ACTS|22|9|跟我一起的人看見了那光，卻沒有聽見那位對我說話的聲音。
ACTS|22|10|我說：『主啊，我該做甚麼？』主說：『起來，進 大馬士革 去，在那裏有人會把指派你做的一切事告訴你。』
ACTS|22|11|我因那光的閃耀不能看見，跟我一起的人就拉著我的手進了 大馬士革 。
ACTS|22|12|「那裏有一個人，名叫 亞拿尼亞 ，按著律法是虔誠人，為所有住在那裏的 猶太 人所稱讚。
ACTS|22|13|他來見我，站在旁邊，對我說：『 掃羅 弟兄，你看見吧！』就在那時，我恢復視覺，看見了他。
ACTS|22|14|他又說：『我們祖宗的上帝揀選了你，讓你明白他的旨意，又看見那義者，聽見他口中所出的聲音。
ACTS|22|15|因為你要將所看見的、所聽見的，對著萬人作他的見證人。
ACTS|22|16|現在你為甚麼耽延呢？起來，受洗，求告他的名，洗去你的罪。』」
ACTS|22|17|「後來，我回到 耶路撒冷 ，在聖殿裏禱告的時候，魂遊象外，
ACTS|22|18|看見主對我說：『你趕緊離開 耶路撒冷 ，越快越好，因為這裏的人不接受你為我作的見證。』
ACTS|22|19|我就說：『主啊，他們都知道，我從前在各會堂裏把信你的人監禁，又鞭打他們。
ACTS|22|20|當你的見證人 司提反 被害流血的時候，我也站在一旁贊同；又為打死他的人看守衣裳。』
ACTS|22|21|主對我說：『你去吧！我要差你到遠方外邦人那裏去。』」
ACTS|22|22|眾人聽他說到這句話，就高聲說：「這樣的人，從地上除掉他吧！他是該死的。」
ACTS|22|23|大家一邊喧嚷一邊摔衣裳，向空中撒灰塵。
ACTS|22|24|千夫長下令把 保羅 帶進營樓，叫人用鞭子拷問他，要知道他們向他這樣喧嚷是甚麼緣故。
ACTS|22|25|他們剛用皮條把他捆上的時候， 保羅 對站在旁邊的百夫長說：「一個 羅馬 人，又未被定罪，你們就鞭打他是合法的嗎？」
ACTS|22|26|百夫長聽見這話，就去見千夫長，報告說：「你要怎麼辦呢？這個人是 羅馬 人。」
ACTS|22|27|千夫長就來問 保羅 ：「你告訴我，你是 羅馬 人嗎？」 保羅 說：「是。」
ACTS|22|28|千夫長回答：「我用了許多銀子才得到 羅馬 公民的身份。」 保羅 說：「我生來就是。」
ACTS|22|29|於是那些要拷問 保羅 的人立刻離開他走了。千夫長一知道他是 羅馬 人，又因為曾捆綁了他，也害怕起來。
ACTS|22|30|第二天，千夫長為要知道 猶太 人控告 保羅 的實情，就解開他，下令祭司長們和全議會的人都聚集，然後將 保羅 帶下來，叫他站在他們面前。
ACTS|23|1|保羅 定睛看著議會的人，說：「諸位弟兄，我在上帝面前，行事為人都是憑著清白的良心，直到今日。」
ACTS|23|2|亞拿尼亞 大祭司就吩咐旁邊站著的人打他的嘴。
ACTS|23|3|這時， 保羅 對他說：「你這粉飾的牆，上帝要打你！你坐堂是要按律法審問我，你竟違背律法，命令人打我嗎？」
ACTS|23|4|站在旁邊的人說：「你竟敢辱罵上帝的大祭司嗎？」
ACTS|23|5|保羅 說：「弟兄們，我不知道他是大祭司；因為經上記著：『不可毀謗你百姓的官長。』」
ACTS|23|6|保羅 看出他們一部分是撒都該人，一部分是法利賽人，就在議會中喊著：「諸位弟兄，我是法利賽人，也是法利賽人的子孫。我現在受審問是為有關死人復活的盼望。」
ACTS|23|7|說了這話，法利賽人和撒都該人爭論起來，會眾分為兩派。
ACTS|23|8|因為撒都該人一方面說沒有復活，另一方面沒有天使和鬼魂；法利賽人卻承認兩方面都有。
ACTS|23|9|於是大大地爭吵起來；有幾個法利賽派的文士站起來爭辯說：「我們看不出這人有甚麼錯處；說不定有鬼魂或者天使對他說過話呢！」
ACTS|23|10|那時爭辯越來越大，千夫長恐怕 保羅 被他們扯碎了，就命令士兵下去，把他從眾人當中搶出來，帶進營樓去。
ACTS|23|11|當夜，主站在 保羅 旁邊，說：「放心吧！你怎樣在 耶路撒冷 為我作見證，也必怎樣在 羅馬 為我作見證。」
ACTS|23|12|到了天亮， 猶太 人同謀起誓，說「若不先殺 保羅 就不吃不喝」。
ACTS|23|13|參與這陰謀的有四十多人。
ACTS|23|14|他們來見祭司長和長老，說：「我們已經發了重誓，若不先殺 保羅 就甚麼也不吃。
ACTS|23|15|現在你們和議會要通知千夫長，叫他把 保羅 帶到你們這裏來，假裝要詳細調查他的事；我們已經預備好，在他來到這裏以前就殺掉他。」
ACTS|23|16|保羅 的外甥聽見他們設下埋伏，就來到營樓裏告訴 保羅 。
ACTS|23|17|保羅 請一個百夫長來，說：「你領這青年去見千夫長，他有事告訴他。」
ACTS|23|18|於是百夫長把他領去見千夫長，說：「被囚的 保羅 請我到他那裏，求我領這青年來見你；他有事告訴你。」
ACTS|23|19|千夫長就拉著他的手，走到一旁，私下問他：「你有甚麼事告訴我呢？」
ACTS|23|20|他說：「 猶太 人已經約定，要求你明天把 保羅 帶到議會去，假裝要詳細查問他的事。
ACTS|23|21|你切不要隨從他們，因為他們有四十多人埋伏，已經起誓，若不先殺掉 保羅 就不吃不喝。現在都預備好了，只等你的允准。」
ACTS|23|22|於是千夫長打發那青年走，囑咐他：「不要告訴人，你已將這些事報告我了。」
ACTS|23|23|於是，千夫長叫了兩個百夫長來，說：「預備步兵二百、騎兵七十、長槍手二百，今夜九點往 凱撒利亞 去；
ACTS|23|24|也要預備牲口讓 保羅 騎上，護送到 腓力斯 總督那裏去。」
ACTS|23|25|千夫長又寫了公文，大略說：
ACTS|23|26|「 克勞第．呂西亞 向 腓力斯 總督大人請安。
ACTS|23|27|這個人被 猶太 人拿住，快被殺害時，我得知他是 羅馬 人，就帶士兵下去，把他救了出來。
ACTS|23|28|因為我要知道他們告他的罪狀，就帶他下到他們的議會去。
ACTS|23|29|我查知他被告發是因他們律法上的爭論，並沒有甚麼該死或該監禁的罪名。
ACTS|23|30|後來有人把要害他的計謀告訴我，我立刻把他解到你那裏去，又命令告他的人在你面前告他。 」
ACTS|23|31|於是士兵照所命令他們的，連夜把 保羅 帶到 安提帕底 。
ACTS|23|32|第二天，由騎兵護送 保羅 ，他們就回營樓去。
ACTS|23|33|騎兵來到 凱撒利亞 ，把公文呈給總督，就叫 保羅 站在他面前。
ACTS|23|34|總督讀了公文，問 保羅 是哪一省的人；一知道他是 基利家 人，
ACTS|23|35|就說：「等告你的人來到，我才詳細聽你。」於是他命令把 保羅 拘留在 希律 的衙門裏。
ACTS|24|1|過了五天， 亞拿尼亞 大祭司、幾個長老和一個叫 帖土羅 的律師下來，向總督控告 保羅 。
ACTS|24|2|保羅 一被傳來， 帖土羅 就開始控告他，說：「 腓力斯 大人，我們因你得以享受國泰民安，並且這一國的弊病，因著你的遠見得以改革。
ACTS|24|3|我們隨時隨地都滿心感激不盡。
ACTS|24|4|為了不敢耽擱你太久，我只求你寬容一下，聽我們說幾句話。
ACTS|24|5|我們看這個人如同瘟疫一般，是鼓動普天下所有的 猶太 人作亂的人，又是 拿撒勒 教派裏的一個頭目。
ACTS|24|6|他甚至連聖殿也要污穢，我們就把他捉拿了。
ACTS|24|7|
ACTS|24|8|你自己審問他，就可以知道我們所控告他的一切事了。」
ACTS|24|9|眾 猶太 人也隨著控告他，說：「這些事情確是這樣。」
ACTS|24|10|總督示意叫 保羅 說話， 保羅 就回答：「我知道你在本國作法官多年，所以我樂意為自己申辯。
ACTS|24|11|你查問就可以知道，從我上 耶路撒冷 去禮拜到今日不過十二天。
ACTS|24|12|他們並沒有看見我在聖殿裏跟人辯論，或在會堂裏、在城裏煽動群眾。
ACTS|24|13|也不能對你證實他們現在所控告我的事。
ACTS|24|14|但有一件事我向你承認，就是我正按著他們所稱為異端的道事奉我祖宗的上帝，又信合乎律法和先知書上所記載的一切。
ACTS|24|15|我對上帝存著這些人自己也接受的盼望，就是義人和不義的人都要復活。
ACTS|24|16|因此，我勉勵自己，對上帝對人，時常存著無虧的良心。
ACTS|24|17|過了幾年，我帶著賙濟本國的捐項和供物上去。
ACTS|24|18|正獻的時候，他們看見我在聖殿裏已經潔淨了，並沒有聚眾，也沒有吵嚷，
ACTS|24|19|惟有幾個從 亞細亞 來的 猶太 人—他們若有控告我的事，應當到你面前來告我。
ACTS|24|20|不然，讓這些人自己說，他們看出我站在議會前的時間，有甚麼不對的地方。
ACTS|24|21|縱然有，也不過是為了一句話，就是我站在他們中間喊說：『我今日在你們面前受審，是為了死人復活。』」
ACTS|24|22|腓力斯 本是詳細認識這道，就拖延他們，說：「且等 呂西亞 千夫長下來，我再審判你們的案。」
ACTS|24|23|於是他下令百夫長看守 保羅 ，要從寬待他，不可攔阻他的親友來供給他。
ACTS|24|24|過了幾天， 腓力斯 和他夫人 猶太 女子 土西拉 一同來到，就叫 保羅 來，聽他講論信基督耶穌的事。
ACTS|24|25|保羅 講論公義、節制和將來的審判， 腓力斯 害怕起來，就回答：「你暫且去吧！等我有機會時再來叫你。」
ACTS|24|26|腓力斯 又指望 保羅 送他銀錢，所以屢次叫他來，和他談論。
ACTS|24|27|過了兩年， 波求．非斯都 接了 腓力斯 的任； 腓力斯 要討 猶太 人的喜歡，就把 保羅 留在監裏。
ACTS|25|1|非斯都 到省裏上任，過了三天，就從 凱撒利亞 上 耶路撒冷 去。
ACTS|25|2|祭司長和 猶太 人的領袖向他控告 保羅 ；又央求他，
ACTS|25|3|向他求情要對付 保羅 ，把他提到 耶路撒冷 來，他們要在路上埋伏殺害他。
ACTS|25|4|非斯都 就回答：「 保羅 押在 凱撒利亞 ，我自己快要往那裏去。」
ACTS|25|5|他又說：「所以，你們中間有權的人與我一同下去，那人若有甚麼不是，就讓他們控告他。」
ACTS|25|6|非斯都 在他們那裏住了不超過八天或十天，就下 凱撒利亞 去；第二天開庭，下令把 保羅 提上來。
ACTS|25|7|保羅 來了，那些從 耶路撒冷 下來的 猶太 人周圍站著，提出許多嚴重而不能證實的事控告他。
ACTS|25|8|保羅 申辯說：「無論 猶太 人的律法，或是聖殿，或是凱撒，我都沒有干犯。」
ACTS|25|9|但 非斯都 要討 猶太 人的喜歡，就回答 保羅 說：「你願意上 耶路撒冷 去，在那裏為這些事受我的審判嗎？」
ACTS|25|10|保羅 說：「我現在站在凱撒的審判臺前，這就是我應當受審的地方。我並沒有對 猶太 人做過甚麼不對的事，這也是你明明知道的。
ACTS|25|11|我若做了不對的事，犯了甚麼該死的罪，就是死我也不辭。他們所控告我的事若都不實，就沒有人能把我交給他們。我要向凱撒上訴。」
ACTS|25|12|非斯都 和議會商量了，就回答：「既然你要向凱撒上訴，你就到凱撒那裏去吧。」
ACTS|25|13|過了些日子， 亞基帕 王和 百妮基 來到 凱撒利亞 ，拜訪 非斯都 。
ACTS|25|14|他們在那裏住了好些日子， 非斯都 將 保羅 的案件向王陳述，說：「這裏有一個人，是 腓力斯 留在監裏的。
ACTS|25|15|我在 耶路撒冷 的時候，祭司長和 猶太 的長老把他的事稟報了，要求定他的罪。
ACTS|25|16|我回覆他們，無論甚麼人，被告還沒有和原告當面對質，沒有機會為所控告的事申辯，就先定他罪的，這不是 羅馬 人的規矩。
ACTS|25|17|及至他們都來到這裏，我沒有耽誤，第二天就開庭，下令把那人提上來。
ACTS|25|18|控告他的人站起來告他，所控告的並沒有任何我所預料的那等惡 事。
ACTS|25|19|不過，有幾樣辯論是有關他們自己敬鬼神的事，以及一個名叫耶穌的人，他已經死了， 保羅 卻說他是活著的。
ACTS|25|20|我對這些事不知該怎樣處理，所以問他是否願意上 耶路撒冷 去，在那裏為這些事接受審判。
ACTS|25|21|但 保羅 要求我留下他，要聽皇上判斷，我就下令把他留下，等我解他到凱撒那裏去。」
ACTS|25|22|亞基帕 對 非斯都 說：「我也願意親自聽聽這個人。」 非斯都 說：「明天你就可以聽他。」
ACTS|25|23|第二天， 亞基帕 和 百妮基 大張旗鼓而來，與眾千夫長和城裏的顯要進了大廳。 非斯都 一聲令下，就有人將 保羅 帶進來。
ACTS|25|24|非斯都 說：「 亞基帕 王和在這裏的諸位，你們看這個人，他就是所有在 耶路撒冷 和這裏的 猶太 人曾向我懇求呼叫，說不可容他再活著的。
ACTS|25|25|但我查明他並沒有犯甚麼該死的罪，並且他自己也已向皇帝上訴了，所以我決定把他解去。
ACTS|25|26|論到這個人，我沒有確實的事可以奏明主上。因此，我帶他到你們面前，尤其到你 亞基帕 王面前，為要在查問之後有所呈奏。
ACTS|25|27|因為據我看，解送囚犯而不指明他的罪狀是不合理的。」
ACTS|26|1|亞基帕 對 保羅 說：「准你為自己申訴。」於是 保羅 伸手辯護說：
ACTS|26|2|「 亞基帕 王啊， 猶太 人所控告我的一切事，今日得以在你面前辯護，實為萬幸。
ACTS|26|3|更慶幸的是你熟悉 猶太 人的規矩和他們的爭論；所以，求你耐心聽我。
ACTS|26|4|「我自幼為人如何，從起初在本國的同胞中，以及在 耶路撒冷 ，所有的 猶太 人都知道。
ACTS|26|5|他們若肯作見證，就知道我從起初是按著我們教中最嚴緊的教門作了法利賽人。
ACTS|26|6|現在我站在這裏受審，是為了對上帝向我們祖宗的應許存著盼望。
ACTS|26|7|這應許，我們十二個支派，晝夜切切地事奉上帝，都指望得著。王啊，我正是因這指望被 猶太 人控告。
ACTS|26|8|上帝使死人復活，你們為甚麼判斷為不可信呢？
ACTS|26|9|「從前我自己認為必須竭力反對 拿撒勒 人耶穌的名，
ACTS|26|10|我在 耶路撒冷 也曾這樣做過；我不但從祭司長得了權柄，把許多聖徒收在監裏，而且他們被殺，我也表示 贊成。
ACTS|26|11|在各會堂，我屢次用刑強迫他們說褻瀆的話，我非常厭惡他們，甚至追逼他們，直到外邦的城鎮。」
ACTS|26|12|「那時，我帶著祭司長的權柄和命令往 大馬士革 去。
ACTS|26|13|王啊！我在路上，中午的時候，看見從天上有一道光，比太陽還亮，四面照射著我和跟我同行的人。
ACTS|26|14|我們都仆倒在地，我就聽見有聲音用 希伯來 話對我說：『 掃羅 ！ 掃羅 ！你為甚麼迫害我？你用腳踢刺棒是自找苦吃的！』
ACTS|26|15|我說：『主啊，你是誰？』主說：『我就是你所迫害的耶穌。
ACTS|26|16|起來，站著，我向你顯現的目的是要派你作僕役，為你所看見我 的事，和我將要指示你的事作見證人。
ACTS|26|17|我也要救你脫離百姓和外邦人的手。我差你到他們那裏去，
ACTS|26|18|要開他們的眼睛，使他們從黑暗中轉向光明，從撒但權下歸向上帝；使他們因信我而得蒙赦罪，和一切成聖的人同得基業。』」
ACTS|26|19|「因此， 亞基帕 王啊！我沒有違背那從天上來的異象；
ACTS|26|20|我先在 大馬士革 ，後在 耶路撒冷 和 猶太 全地，以及外邦，勸勉他們應當悔改歸向上帝，行事與悔改的心相稱。
ACTS|26|21|為這緣故， 猶太 人在聖殿裏拿住我，想要殺我。
ACTS|26|22|然而，我蒙上帝的幫助，直到今日還站立得穩，向尊貴的和卑微的作見證。我所講的，並不外乎眾先知和 摩西 所說將來必成的事，
ACTS|26|23|就是基督必須受害，並且首先從死人中復活，把亮光傳給 猶太 人和外邦人。」
ACTS|26|24|保羅 這樣申訴時， 非斯都 大聲說：「 保羅 ，你瘋了！你的學問太大，反使你瘋了！」
ACTS|26|25|保羅 說：「 非斯都 大人，我不是瘋了，我說的乃是真實和清醒的話。
ACTS|26|26|王也知道這些事，所以對王大膽直言，我深信這些事沒有一件能向王隱瞞的，因為都不是在背地裏做的。
ACTS|26|27|亞基帕 王啊，你信先知嗎？我知道你是信的。」
ACTS|26|28|亞基帕 對 保羅 說：「你想稍微勸一勸就能說服我作基督徒了嗎？」
ACTS|26|29|保羅 說：「無論少勸還是多勸，我向上帝所求的，不但你一個人，就是今天所有聽我說話的人都要像我一樣，只是不要有這些鎖鏈。」
ACTS|26|30|於是，王和總督以及 百妮基 跟同坐的人都站起來，
ACTS|26|31|退到裏面，彼此談論說：「這個人並沒有犯甚麼該死該監禁的罪。」
ACTS|26|32|亞基帕 對 非斯都 說：「這人若沒有向凱撒上訴，早就被釋放了。」
ACTS|27|1|既然 非斯都 決定要我們坐船往 意大利 去，就將 保羅 和別的囚犯交給御營裏的一個名叫 猶流 的百夫長。
ACTS|27|2|有一隻 亞大米田 的船要開往 亞細亞 沿海一帶地方去，我們上了那船，就起航了；有 馬其頓 的 帖撒羅尼迦 人 亞里達古 和我們同去。
ACTS|27|3|第二天，我們到了 西頓 。 猶流 寬待 保羅 ，准他往朋友那裏去，受他們的照應。
ACTS|27|4|我們又從那裏開船，因為遇到逆風，就貼著 塞浦路斯 的背風岸航行，
ACTS|27|5|渡過了 基利家 、 旁非利亞 一帶的海面，就到了 呂家 的 每拉 。
ACTS|27|6|在那裏，百夫長找到一隻 亞歷山大 的船要往 意大利 去，就叫我們上了那船。
ACTS|27|7|一連多日，船行得很慢，我們好不容易才來到 革尼土 的對面；又因被風攔阻，我們就貼著 克里特 島背風岸，從 撒摩尼 對面航行。
ACTS|27|8|我們沿岸前進，十分艱難，來到一個名叫 佳澳 的地方，離那裏不遠有 拉西亞城 。
ACTS|27|9|航行的日子久了，已經過了禁食的節期，行船又危險， 保羅 就建議，
ACTS|27|10|對眾人說：「諸位，我看這次航行，不但貨物和船要受損傷，大遭破壞，連我們的性命也難保。」
ACTS|27|11|但百夫長信從船長和船主，不信 保羅 所說的。
ACTS|27|12|且因在這港口不適宜過冬，船上大多數的人都主張開船離開這地方，或者能到 非尼基 去過冬。 非尼基 是 克里特 的一個港口，一面朝西南，一面朝西北。
ACTS|27|13|當南風微微吹起時，他們以為對目的地已有了把握，就起錨，貼近 克里特 開去。
ACTS|27|14|過了不久，有一股叫「友拉革羅」的東北巨風從島上撲來，
ACTS|27|15|船被風抓住，無法頂風航行，我們只好任它漂流。
ACTS|27|16|我們貼著一個叫 高大 的小島的背風岸急航，好不容易才保住了救生艇。
ACTS|27|17|既然把救生艇拉上來，他們就用纜索捆綁船底，又恐怕在 賽耳底 淺灘上擱淺，就落了篷，任船漂流。
ACTS|27|18|我們被風浪逼得很急，第二天眾人就把貨物拋在海裏。
ACTS|27|19|第三天，他們又親手把船上的器具拋棄了。
ACTS|27|20|許多天都沒有看到太陽和星辰，又有狂風大浪催逼，我們獲救的指望都放棄了。
ACTS|27|21|眾人已有好幾天沒有吃東西， 保羅 就出來站在他們中間，說：「諸位，你們本該聽我的話不離開 克里特 島，就不致遭到這樣的損失和破壞。
ACTS|27|22|現在我勸你們放心，除了損失這條船，你們中間沒有一人會喪失性命。
ACTS|27|23|因為昨夜，我所屬所事奉的上帝的使者站在我旁邊，
ACTS|27|24|說：『 保羅 ，不要害怕，你必定站在凱撒面前；並且上帝已把安全賜給與你同船的人了。』
ACTS|27|25|所以，諸位可以放心，我信上帝怎樣對我說，事情也要怎樣成就；
ACTS|27|26|只是我們必須在一個島上擱淺。」
ACTS|27|27|到了第十四天夜間，船在 亞得里亞海 漂來漂去。約在半夜，水手以為漸近旱地，
ACTS|27|28|就去探測深淺，探得有十二丈 ；稍往前行，又探深淺，探得有九丈。
ACTS|27|29|恐怕我們撞到礁石，他們就從船尾拋下四個錨，盼望天亮。
ACTS|27|30|水手想棄船逃走，把救生艇縋下海裏，假裝要從船頭拋錨的樣子。
ACTS|27|31|保羅 對百夫長和士兵說：「這些人若不留在船上，你們就不能獲救。」
ACTS|27|32|於是士兵砍斷救生艇的繩子，由它漂去。
ACTS|27|33|天快亮的時候， 保羅 勸眾人都用餐，說：「你們一直捱餓等候，不吃甚麼，已經十四天了。
ACTS|27|34|所以我勸你們吃點東西，這是關乎你們獲救的，因為你們各人連一根頭髮也不至於掉落。」
ACTS|27|35|保羅 說了這話，就拿起餅來，在眾人面前祝謝了上帝，然後擘開來吃。
ACTS|27|36|於是他們都放心，就吃了。
ACTS|27|37|我們在船上的共有二百七十六個人。
ACTS|27|38|他們吃飽了，為要使船輕一點，就把船上的麥子拋到海裏。
ACTS|27|39|天亮的時候，他們不認得那地方，只見一個有岸可登的海灣，就想法子看能不能把船靠岸。
ACTS|27|40|於是他們砍斷纜索，把錨丟到海裏，同時也鬆開舵繩，拉起頭篷，順風向著岸行去。
ACTS|27|41|但碰到兩水夾流的地方，就擱了淺，船頭膠住不動，船尾被浪的猛力衝壞了 。
ACTS|27|42|士兵的意思要把囚犯都殺了，免得有游水脫逃的。
ACTS|27|43|但百夫長要救 保羅 ，不准他們任意而行，就吩咐會游水的，跳下水去，先上岸；
ACTS|27|44|其餘的人則用板子或船的碎片上岸。這樣，眾人都獲救，上了岸。
ACTS|28|1|我們既已獲救，才知道那島名叫 馬耳他 。
ACTS|28|2|當地人非常友善地接待我們；因為正在下雨，天氣又冷，他們就生了火歡迎我們眾人。
ACTS|28|3|那時， 保羅 拾起一捆柴，放在火中，有一條毒蛇，因為熱的緣故鑽了出來，纏住他的手。
ACTS|28|4|當地的人看見那毒蛇懸在他手上，就彼此說：「這人必是個兇手，雖然他從海裏獲救，天理仍不容他活著。」
ACTS|28|5|保羅 竟把那毒蛇甩在火裏，並沒有受傷。
ACTS|28|6|當地的人想他快要腫起來，或是忽然倒下死了，但等了好久，見他沒有甚麼異樣，就轉念說他是個神明。
ACTS|28|7|離那地方不遠有一些田產，是島長 部百流 的。他接納我們，盡情款待了我們三日。
ACTS|28|8|當時， 部百流 的父親臥病不起，患了熱病和痢疾。 保羅 進去見他，為他禱告按手，治好了他。
ACTS|28|9|從此，島上其餘的病人也都來，得了醫治。
ACTS|28|10|他們又多方面尊敬我們，到了開船的時候，又把我們所需用的東西送到船上。
ACTS|28|11|過了三個月，我們上了 亞歷山大 的船起航。這船以「 宙斯 雙子」為記，是在那海島過冬的。
ACTS|28|12|我們到了 敘拉古 ，停泊了三日；
ACTS|28|13|又從那裏起錨開船， 來到 利基翁 。過了一天，起了南風，第二天就來到 部丟利 。
ACTS|28|14|我們在那裏遇見一些弟兄，他們請我們同住了七天。就這樣，我們來到 羅馬 。
ACTS|28|15|那裏的弟兄們一聽見我們的消息，就到 亞比烏 市和 三館 來迎接我們。 保羅 見了他們，就感謝上帝，越發壯膽。
ACTS|28|16|我們進了 羅馬城 ， 保羅 蒙准和那個看守他的兵另住在一處。
ACTS|28|17|過了三天， 保羅 請當地 猶太 人的領袖來。他們來了， 保羅 對他們說：「諸位弟兄，雖然我沒有做甚麼事干犯本國的百姓和我們祖宗的規矩，卻在 耶路撒冷 被囚禁，交在 羅馬 人的手裏。
ACTS|28|18|他們審問了我，有意要釋放我，因為在我身上並沒有該死的罪狀。
ACTS|28|19|但 猶太 人反對，我不得已只好上訴於凱撒，並不是有甚麼事要控告我本國的百姓。
ACTS|28|20|為這緣故，我請你們來見我當面談話，我原是為 以色列 人所指望的那位才被這鐵鏈捆綁的。」
ACTS|28|21|他們對他說：「我們並沒有接到從 猶太 寄來有關於你的信，也沒有弟兄到這裏來向我們報告，或說你有甚麼不好的地方。
ACTS|28|22|但我們願意聽聽你的意見，因為我們知道這教門是到處遭人反對的。」
ACTS|28|23|他們和 保羅 約定了日子，就有許多人到他的住處來。 保羅 從早到晚向他們講解這事，為上帝的國作證，並引 摩西 的律法和先知的書勸導他們信從耶穌。
ACTS|28|24|他所說的話，有的信，有的不信。
ACTS|28|25|他們間彼此不合，就分散了；未散以先， 保羅 說了一句話：「聖靈藉 以賽亞 先知向你們祖宗所說的話是對的。
ACTS|28|26|他說： 『你去對這百姓說： 你們聽了又聽，卻不明白； 看了又看，卻看不清。
ACTS|28|27|因為這百姓的心麻木， 耳朵塞著， 眼睛閉著， 免得眼睛看見， 耳朵聽見， 心裏明白，回轉過來， 我會醫治他們。』
ACTS|28|28|所以，你們當知道，上帝這救恩已經傳給外邦人；他們會聽的。」
ACTS|28|29|
ACTS|28|30|保羅 在自己所租的房子裏住了足足兩年。凡來見他的人，他都接待，
ACTS|28|31|放膽傳講上帝的國，並教導主耶穌基督的事，沒有人禁止。
ROM|1|1|基督耶穌的僕人 保羅 ，蒙召為使徒，奉派傳上帝的福音。
ROM|1|2|這福音是上帝從前藉眾先知，在聖經上所應許的。
ROM|1|3|論到他兒子－我主耶穌基督，按肉體說，是從 大衛 後裔生的；按神聖的靈說，因從死人中復活，用大能顯明他是上帝的兒子。
ROM|1|4|
ROM|1|5|我們從他蒙恩受了使徒的職分，為他的名在萬國中使人因信而順服，
ROM|1|6|其中也有你們這蒙召屬耶穌基督的人。
ROM|1|7|我寫信給你們在 羅馬 、為上帝所愛、蒙召作聖徒的眾人。願恩惠、平安 從我們的父上帝和主耶穌基督歸給你們！
ROM|1|8|首先，我靠著耶穌基督，為你們眾人感謝我的上帝，因你們的信德傳遍了天下。
ROM|1|9|我在他兒子的福音上，用心靈所事奉的上帝可以見證，我怎樣不住地提到你們，
ROM|1|10|在我的禱告中常常懇求，或許照上帝的旨意，最終我能毫無阻礙地往你們那裏去。
ROM|1|11|因為我迫切地想見你們，要把一些屬靈的恩賜分給你們，使你們得以堅固，
ROM|1|12|也可以說，我在你們中間，因你我彼此的信心而同得安慰。
ROM|1|13|弟兄們，我不願意你們不知道，我屢次計劃往你們那裏去，要在你們中間得些果子，如同在其餘的外邦人中一樣，只是到如今仍有攔阻。
ROM|1|14|無論是 希臘 人、未開化的人、聰明人、愚拙人，我都欠他們的債，
ROM|1|15|所以願意盡我的力量把福音也傳給你們在 羅馬 的人。
ROM|1|16|我不以福音為恥；這福音本是上帝的大能，要救一切相信的，先是 猶太 人，後是 希臘 人。
ROM|1|17|因為上帝的義正在這福音上顯明出來；這義是本於信，以至於信。如經上所記：「義人必因信得生。」
ROM|1|18|原來，上帝的憤怒從天上顯明在一切不虔不義的人身上，就是那些行不義壓制真理的人。
ROM|1|19|上帝的事情，人所能知道的，原顯明在人心裏，因為上帝已經向他們顯明。
ROM|1|20|自從造天地以來，上帝的永能和神性是明明可知的，雖然眼不能見，但藉著所造之物就可以了解看見，叫人無可推諉。
ROM|1|21|因為，他們雖然知道上帝，卻不把他當作上帝榮耀他，也不感謝他。他們的思想變為虛妄，無知的心昏暗了。
ROM|1|22|他們自以為聰明，反成了愚昧，
ROM|1|23|將不能朽壞之上帝的榮耀變為偶像，仿照必朽壞的人、飛禽、走獸、爬蟲的形像。
ROM|1|24|所以，上帝任憑他們隨著心裏的情慾行污穢的事，以致彼此羞辱自己的身體。
ROM|1|25|他們將上帝的真實變為虛謊，去敬拜事奉受造之物，不敬奉那造物的主—主是可稱頌的，直到永遠。阿們！
ROM|1|26|因此，上帝任憑他們放縱可羞恥的情慾。他們的女人把自然的關係變成違反自然的；
ROM|1|27|男人也是如此，放棄了和女人自然的關係，慾火攻心，男的和男的彼此貪戀，行可恥的事，就在自己身上受這逆性行為當得的報應。
ROM|1|28|他們既然故意不認識上帝，上帝就任憑他們存扭曲的心，做那些不該做的事，
ROM|1|29|裝滿了各樣不義 、邪惡、貪婪、惡毒，滿心是嫉妒、兇殺、紛爭、詭詐、毒恨，又是毀謗的、
ROM|1|30|說人壞話的、怨恨上帝的 、侮辱人的、狂傲的、自誇的、製造是非的、忤逆父母的、
ROM|1|31|頑梗不化的、言而無信的、無情無義的、不憐憫人的。
ROM|1|32|他們雖知道上帝判定做這樣事的人是該死的，然而他們不但自己去做，還贊同別人去做。
ROM|2|1|所以，你這評斷人的人哪，無論你是誰，都無可推諉。你在甚麼事上評斷人，就在甚麼事上定自己的罪。因你這評斷人的，自己所做的卻和別人一樣。
ROM|2|2|我們知道這樣做的人，上帝必公平地審判他。
ROM|2|3|你這個人哪，你評斷做這樣事的人，自己所做的卻和別人一樣，你以為能逃脫上帝的審判嗎？
ROM|2|4|還是你藐視他豐富的恩慈、寬容、忍耐，不知道他的恩慈是領你悔改嗎？
ROM|2|5|你竟放任你剛硬不悔改的心，為自己累積憤怒！在憤怒的日子，上帝公義的審判要顯示出來。
ROM|2|6|他要照各人的行為報應各人。
ROM|2|7|凡恆心行善，尋求榮耀、尊貴和不能朽壞的，就有永生報償他們；
ROM|2|8|但是那些自私自利、不順從真理、反順從不義的人，就有惱恨、憤怒報應他們。
ROM|2|9|他要把患難、困苦加給一切作惡的人，先是 猶太 人，後是 希臘 人；
ROM|2|10|卻把榮耀、尊貴、平安加給一切行善的人，先是 猶太 人，後是 希臘 人。
ROM|2|11|因為上帝不偏待人。
ROM|2|12|凡在律法之外犯了罪的，將在律法之外滅亡；凡在律法之內犯了罪的，將按律法受審判。
ROM|2|13|原來在上帝面前，不是聽律法的為義，而是行律法的稱義。
ROM|2|14|沒有律法的外邦人若順著本性行律法上的事，他們雖然沒有律法，自己就是自己的律法。
ROM|2|15|他們顯明律法的功用刻在他們心裏，他們的良心一同作證—他們的內心掙扎，有時自責，有時為自己辯護。
ROM|2|16|在那日，上帝要藉著基督耶穌 ，按照我所傳的福音，審判人隱藏的事。
ROM|2|17|但是你，你既自稱為 猶太 人，倚靠律法，以上帝誇口，
ROM|2|18|知道上帝的旨意，從律法受了教導而能分辨是非；
ROM|2|19|你既深信自己是給盲人領路的，是在黑暗中人的光，
ROM|2|20|是無知的人的師傅，是小孩子的老師，體現了律法中的知識和真理；
ROM|2|21|那麼，你這教導別人的，還不教導自己嗎？你這宣講不可偷竊的，自己還偷竊嗎？
ROM|2|22|你這說不可姦淫的，自己還姦淫嗎？你這厭惡偶像的，自己還搶劫廟中之物嗎？
ROM|2|23|你這以律法誇口的，自己倒違犯律法，羞辱上帝！
ROM|2|24|上帝的名在外邦人中因你們受了褻瀆，正如經上所記的。
ROM|2|25|你若遵行律法，割禮固然於你有益；若違犯律法，你的割禮就算不得割禮。
ROM|2|26|所以，那未受割禮的，若遵守律法的要求，他雖然未受割禮，豈不算是受了割禮嗎？
ROM|2|27|而且那本來未受割禮的，若能全守律法，豈不是要審判你這有儀文和割禮，竟違犯律法的人嗎？
ROM|2|28|因為外表是 猶太 人的不是真 猶太 人；外表肉身的割禮也不是真割禮。
ROM|2|29|惟有內心作 猶太 人的才是真 猶太 人，真割禮也是心裏的，在乎聖靈 ，不在乎儀文。這樣的人所受的稱讚不是從人來的，而是從上帝來的。
ROM|3|1|這樣說來， 猶太 人有甚麼比別人強呢？割禮有甚麼益處呢？
ROM|3|2|很多，各方面都有。首先，上帝的聖言交託他們。
ROM|3|3|即使有不信的，這又何妨呢？難道他們的不信就廢掉上帝的信實嗎？
ROM|3|4|絕對不會！不如說，上帝是真實的，而人都是虛謊的。如經上所記： 「以致你責備的時候顯為公義； 你被指控的時候一定勝訴。」
ROM|3|5|我姑且照著人的看法來說，我們的不義若顯出上帝的義來，我們要怎麼說呢？上帝降怒是他不義嗎？
ROM|3|6|絕對不是！若是這樣，上帝怎能審判世界呢？
ROM|3|7|若上帝的真實因我的虛謊越發顯出他的榮耀，為甚麼我還像罪人一樣受審判呢？
ROM|3|8|為甚麼不說，我們可以作惡以成善呢？有人毀謗我們，說我們講過這話；這等人被定罪是應該的。
ROM|3|9|那又怎麼樣呢？我們比他們強嗎？絕不是！因我們已經指證： 猶太 人和 希臘 人都在罪惡之下。
ROM|3|10|就如經上所記： 「沒有義人，連一個也沒有。
ROM|3|11|沒有明白的， 沒有尋求上帝的。
ROM|3|12|人人偏離正路，一同走向敗壞。 沒有行善的，連一個也沒有 。
ROM|3|13|他們的喉嚨是敞開的墳墓； 他們的舌頭玩弄詭詐。 他們的嘴唇裏有毒蛇的毒液，
ROM|3|14|滿口是咒罵苦毒。
ROM|3|15|他們的腳為殺人流血飛跑；
ROM|3|16|他們的路留下毀壞和災難。
ROM|3|17|和平的路，他們不認識；
ROM|3|18|他們眼中不怕上帝。」
ROM|3|19|我們知道律法所說的話都是對律法之下的人說的，好塞住各人的口，使普世的人都伏在上帝的審判之下。
ROM|3|20|所以，凡血肉之軀沒有一個能因律法的行為而在上帝面前稱義，因為律法本是要人認識罪。
ROM|3|21|但如今，上帝的義在律法之外已經顯明出來，有律法和先知為證：
ROM|3|22|就是上帝的義，因信耶穌基督 加給一切信的人。這並沒有分別，
ROM|3|23|因為世人都犯了罪，虧缺了上帝的榮耀，
ROM|3|24|如今卻蒙上帝的恩典，藉著在基督耶穌裏的救贖，就白白地得稱為義。
ROM|3|25|上帝設立耶穌作贖罪祭，是憑耶穌的血，藉著信，要顯明上帝的義；因為他用忍耐的心寬容人先前所犯的罪，好使今時顯明他的義，讓人知道他自己為義，也稱信耶穌的人為義 。
ROM|3|26|
ROM|3|27|既是這樣，哪裏可誇口呢？沒有可誇的。是藉甚麼法呢？功德嗎？不是！是藉信主之法。
ROM|3|28|所以我們認定，人稱義是因著信，不在於律法的行為。
ROM|3|29|難道上帝只是 猶太 人的嗎？不也是外邦人的嗎？是的，他也是外邦人的上帝。
ROM|3|30|既然上帝是一位，他就要本於信稱那受割禮的為義，也要藉著信稱那未受割禮的為義。
ROM|3|31|這樣，我們藉著信廢了律法嗎？絕對不是！更是鞏固律法。
ROM|4|1|這樣，那按肉體作我們祖宗的 亞伯拉罕 ，我們要怎麼說呢？
ROM|4|2|倘若 亞伯拉罕 是因行為稱義，他就有可誇的，但是在上帝面前他一無可誇。
ROM|4|3|經上說甚麼呢？「 亞伯拉罕 信了上帝，這就算他為義。」
ROM|4|4|做工的得工資不算是恩典，而是應得的；
ROM|4|5|但那不做工的，只信那位稱不敬虔之人為義的，他的信就算為義。
ROM|4|6|正如 大衛 稱那在行為之外蒙上帝算為義的人是有福的：
ROM|4|7|「過犯得赦免，罪惡蒙遮蓋的人有福了！
ROM|4|8|主不算為有罪的，這樣的人有福了！」
ROM|4|9|如此看來，這福只加給那受割禮的人嗎？不也加給那未受割禮的人嗎？我們說，因著信，就算 亞伯拉罕 為義。
ROM|4|10|那麼，這是怎麼算的呢？是在他受割禮的時候呢？還是在他未受割禮的時候呢？不是在受割禮的時候，而是在未受割禮的時候。
ROM|4|11|並且，他受了割禮的記號，作他未受割禮的時候因信稱義的印證，為使他作一切未受割禮而信之人的父，使他們也算為義，
ROM|4|12|也使他作受割禮之人的父，就是那些不但受割禮，而且跟隨我們的祖宗 亞伯拉罕 未受割禮而信的足跡的人。
ROM|4|13|因為上帝給 亞伯拉罕 和他後裔承受世界的應許不是藉著律法，而是藉著信而得的義。
ROM|4|14|若是屬於律法的人才是後嗣，信就落空了，應許也就失效了。
ROM|4|15|因為律法是惹動憤怒的，哪裏沒有律法，哪裏就沒有過犯。
ROM|4|16|所以，人作後嗣是出於信，因此就屬乎恩，以致應許保證歸給所有的後裔，不但歸給那屬於律法的，也歸給那效法 亞伯拉罕 之信的人。 亞伯拉罕 所信的是那叫死人復活、使無變為有的上帝，在這位上帝面前 亞伯拉罕 成為我們眾人的父，如經上所記：「我已經立你作多國之父。」
ROM|4|17|
ROM|4|18|他在沒有盼望的時候，仍存著盼望來相信，就得以作多國之父，正如先前所說：「你的後裔將要如此。」
ROM|4|19|他將近百歲的時候，雖然想到 自己的身體如同已死， 撒拉 也不可能生育，他的信心還是不軟弱，
ROM|4|20|仍仰望上帝的應許，總沒有因不信而起疑惑，反倒因信而剛強，將榮耀歸給上帝，
ROM|4|21|且滿心相信上帝所應許的必能成就。
ROM|4|22|所以這也 就算他為義。
ROM|4|23|「算他為義」這句話不是單為他寫的，
ROM|4|24|也是為我們將來得算為義的人寫的，就是為我們這些信上帝使我們的主耶穌從死人中復活的人寫的。
ROM|4|25|耶穌被出賣，是為我們的過犯；他復活，是為使我們稱義。
ROM|5|1|所以，我們既因信稱義，就藉著我們的主耶穌基督得以與上帝和好。
ROM|5|2|我們又藉著他，因信 得以進入現在所站立的這恩典中，並且歡歡喜喜盼望上帝的榮耀。
ROM|5|3|不但如此，就是在患難中也是歡歡喜喜的，因為知道患難生忍耐，
ROM|5|4|忍耐生老練，老練生盼望，
ROM|5|5|盼望不至於落空，因為上帝的愛，已藉著所賜給我們的聖靈，澆灌在我們心裏。
ROM|5|6|我們還軟弱的時候，基督就在特定的時刻為不敬虔之人死。
ROM|5|7|為義人死，是少有的；為仁人死，也者有敢做的。
ROM|5|8|惟有基督在我們還作罪人的時候為我們死，上帝的愛就在此向我們顯明了。
ROM|5|9|現在我們既靠著他的血稱義，就更要藉著他得救，免受上帝的憤怒。
ROM|5|10|因為我們作仇敵的時候，尚且藉著上帝兒子的死得以與上帝和好，既已和好，就更要因他的生得救了。
ROM|5|11|不但如此，我們既藉著我們的主耶穌基督得以與上帝和好，也就藉著他以上帝為樂。
ROM|5|12|為此，正如罪是從一人進入世界，死又從罪而來，於是死就臨到所有的人，因為人人都犯了罪。
ROM|5|13|沒有律法之前，罪已經在世上，但沒有律法，罪也不算罪。
ROM|5|14|然而，從 亞當 到 摩西 ，死就掌了權，連那些不與 亞當 犯一樣罪過的，也在死的權下。 亞當 是那以後要來之人的預像。
ROM|5|15|但是過犯不如恩賜，若因一人的過犯，眾人都死了，那麼，上帝的恩典，與那因耶穌基督一人而來的恩典中的賞賜，豈不加倍地臨到眾人嗎？
ROM|5|16|因一人犯罪而來的後果，也不如賞賜，原來審判是由一人而定罪，恩賜乃是由許多過犯而稱義。
ROM|5|17|若因一人的過犯，死就因這一人掌權，那些受洪恩又蒙所賜之義的，豈不更要因耶穌基督一人在他們生命中掌權嗎？
ROM|5|18|這樣看來，因一次的過犯，所有的人都被定罪；照樣，因一次的義行，所有的人也就被稱義而得生命了。
ROM|5|19|因一人的悖逆，眾人成為罪人；照樣，因一人的順從，眾人也成為義了。
ROM|5|20|而且加添了律法，使得過犯增加，只是罪在哪裏增加，恩典就在哪裏越發豐盛了。
ROM|5|21|所以，正如罪藉著死掌權；照樣，恩典也藉著義掌權，使人因我們的主耶穌基督得永生。
ROM|6|1|這樣，我們要怎麼說呢？我們可以仍在罪中使恩典增多嗎？
ROM|6|2|絕對不可！我們向罪死了的人，豈可仍在罪中活著呢？
ROM|6|3|難道你們不知道，我們這受洗歸入基督耶穌的人，就是受洗歸入他的死嗎？
ROM|6|4|所以，我們藉著洗禮歸入死，和他一同埋葬，是要我們行事為人都有新生的樣子，像基督藉著父的榮耀從死人中復活一樣。
ROM|6|5|我們若與他合一，經歷與他一樣的死，也將經歷與他一樣的復活。
ROM|6|6|我們知道，我們的舊人和他同釘十字架，使罪身滅絕，叫我們不再作罪的奴隸，
ROM|6|7|因為已死的人是脫離了罪。
ROM|6|8|我們若與基督同死，我們信也必與他同活，
ROM|6|9|因為知道基督既從死人中復活，就不再死，死也不再作他的主了。
ROM|6|10|他死了，是對罪死，只這一次；他活，是對上帝活著。
ROM|6|11|這樣，你們也要看自己對罪是死的，在基督耶穌裏對上帝卻是活的。
ROM|6|12|所以，不要讓罪在你們必死的身上掌權，使你們順從身體的私慾。
ROM|6|13|也不要把你們的肢體獻給罪作不義的工具，倒要像從死人中活著的人，把自己獻給上帝，並把你們的肢體獻給上帝作義的工具。
ROM|6|14|罪必不能作你們的主，因你們不在律法之下，而是在恩典之下。
ROM|6|15|那又怎麼樣呢？我們在恩典之下，不在律法之下，就可以犯罪嗎？絕對不可！
ROM|6|16|難道你們不知道，你們獻自己作奴僕，順從誰就作誰的奴僕嗎？或作罪的奴隸，以至於死；或作順服的奴僕，以至於成義。
ROM|6|17|感謝上帝！因為你們從前雖然作罪的奴隸，現在卻從心裏順服了所傳給你們教導的典範。
ROM|6|18|你們既從罪裏得了釋放，就作了義的奴僕。
ROM|6|19|我因你們肉體的軟弱，就以人的觀點來說。你們從前怎樣把肢體獻給不潔不法作奴隸，以至於不法；現在也要照樣將肢體獻給義作奴僕，以至於成聖。
ROM|6|20|因為你們作罪的奴隸時，不被義所約束。
ROM|6|21|那麼，你們現在所看為羞恥的事，當時有甚麼果子呢？那些事的結局就是死。
ROM|6|22|但如今，你們既從罪裏得了釋放，作了上帝的奴僕，就結出果子，以至於成聖，那結局就是永生。
ROM|6|23|因為罪的工價乃是死；惟有上帝的恩賜，在我們的主基督耶穌裏，乃是永生。
ROM|7|1|弟兄們，我對你們這些明白律法的人說，你們豈不知道律法約束人是在他活著的時候嗎？
ROM|7|2|就如女人有了丈夫，丈夫還活著，她就被律法約束；丈夫若死了，她就從丈夫的律法中解脫了。
ROM|7|3|所以丈夫還活著，她若跟了別的男人，就叫淫婦；丈夫若死了，她就脫離了律法，雖然跟了別的男人，也不是淫婦。
ROM|7|4|我的弟兄們，這樣說來，你們藉著基督的身體對律法也是死了，使你們歸於另一位，就是歸於那從死人中復活的，為要使我們結果子給上帝。
ROM|7|5|因為我們屬肉體的時候，那因律法而生犯罪的慾望在我們肢體中發動，以致結出死亡的果子。
ROM|7|6|但如今，我們既然在捆綁我們的律法上死了，就從律法中解脫，使我們服侍主，要按著聖靈 的新樣，不按著儀文的舊樣。
ROM|7|7|這樣，我們要怎麼說呢？律法是罪嗎？絕對不是！但是，若不是藉著律法，我就不知何為罪；若不是律法說「不可貪心」，我就不知何為貪心。
ROM|7|8|然而，罪趁著機會，藉著誡命，使各樣的貪心在我裏頭發動，因為沒有律法，罪是死的。
ROM|7|9|以前沒有律法的時候，我是活的；但是誡命來到，罪活起來，
ROM|7|10|我就死了。那本該叫人活的誡命反而叫我死。
ROM|7|11|因為罪趁著機會，藉著誡命誘惑我，並且藉著誡命殺了我。
ROM|7|12|這樣看來，律法是聖的，誡命也是聖的、義的、善的。
ROM|7|13|那麼，那善的是叫我死嗎？絕對不是！叫我死的是罪。罪藉著那善的叫我死，為要顯出這真是罪，以致罪藉著誡命更顯出是惡極了。
ROM|7|14|我們原知道律法是屬靈的，我卻是屬肉體的，是已經賣給罪了。
ROM|7|15|因為我所做的，我自己不明白。我所願意的，我並不做；我所恨惡的，我反而去做。
ROM|7|16|如果我所做的是我所不願意的，我得承認律法是善的。
ROM|7|17|事實上，這不是我做的，而是住在我裏面的罪做的。
ROM|7|18|我也知道，住在我裏面的，就是我肉體之中，沒有善。因為立志為善由得我，只是行出來由不得我。
ROM|7|19|我所願意的善，我不去做；我所不願意的惡，我反而去做。
ROM|7|20|如果我去做我不願意做的，就不是我做的，而是住在我裏面的罪做的。
ROM|7|21|我覺得有個律，就是我願意行善的時候，就有惡纏著我。
ROM|7|22|因為，按著我裏面的人，我喜歡上帝的律，
ROM|7|23|但我看出肢體中另有個律和我內心的律交戰，把我擄去，使我附從那肢體中罪的律。
ROM|7|24|我真苦啊！誰能救我脫離這必死的身體呢？
ROM|7|25|感謝上帝，靠著我們的主耶穌基督就能！這樣看來，一方面，我內心順服上帝的律，另一方面，肉體卻順服罪的律了。
ROM|8|1|如今，那些在基督耶穌裏的人就不被定罪了。
ROM|8|2|因為賜生命的聖靈的律，在基督耶穌裏從罪和死的律中把你釋放出來。
ROM|8|3|律法既因肉體軟弱而無能為力，上帝就差遣自己的兒子成為罪身的樣子，為了對付罪 ，在肉體中定了罪，
ROM|8|4|為要使律法要求的義，實現在我們這不隨從肉體、只隨從聖靈去行的人身上。
ROM|8|5|因為，隨從肉體的人體貼肉體的事；隨從聖靈的人體貼聖靈的事。
ROM|8|6|體貼肉體就是死；體貼聖靈就是生命和平安 。
ROM|8|7|因為體貼肉體就是與上帝為敵，對上帝的律法不順服，事實上也無法順服。
ROM|8|8|屬肉體的人無法使上帝喜悅。
ROM|8|9|如果上帝的靈住在你們裏面，你們就不屬肉體，而是屬聖靈了。人若沒有基督的靈，就不是屬基督的。
ROM|8|10|基督若在你們裏面，身體就因罪而死，靈卻因義而活。
ROM|8|11|然而，使耶穌從死人中復活的上帝的靈若住在你們裏面，那使基督從死人中復活的，也必藉著住在你們裏面的聖靈使你們必死的身體又活過來。
ROM|8|12|弟兄們，這樣看來，我們不是欠肉體的債去順從肉體而活。
ROM|8|13|你們若順從肉體活著，必定會死；若靠著聖靈把身體的惡行處死，就必存活。
ROM|8|14|因為凡被上帝的靈引導的都是上帝的兒子。
ROM|8|15|你們所領受的不是奴僕的靈，仍舊害怕；所領受的是兒子名分的靈，因此我們呼叫：「阿爸，父！」
ROM|8|16|聖靈自己與我們的靈一同見證我們是上帝的兒女。
ROM|8|17|若是兒女，就是後嗣，是上帝的後嗣，和基督同作後嗣。如果我們和他一同受苦，是要我們和他一同得榮耀。
ROM|8|18|我認為，現在的苦楚，若比起將來要顯示給我們的榮耀，是不足介意的。
ROM|8|19|受造之物切望等候上帝的眾子顯出來。
ROM|8|20|因為受造之物屈服在虛空之下，不是自己願意，而是因那使它屈服的叫他如此。但受造之物仍然指望從敗壞的轄制下得釋放，得享上帝兒女榮耀的自由。
ROM|8|21|
ROM|8|22|我們知道，一切受造之物一同呻吟，一同忍受陣痛，直到如今。
ROM|8|23|不但如此，就是我們這有聖靈作初熟果子的，也是自己內心呻吟，等候得著兒子的名分，就是我們的身體得救贖。
ROM|8|24|我們得救是在於盼望；可是看得見的盼望就不是盼望。誰還去盼望他所看得見的呢？
ROM|8|25|但我們若盼望那看不見的，我們就耐心等候。
ROM|8|26|同樣，我們的軟弱有聖靈幫助。我們本不知道當怎樣禱告，但是聖靈親自用無可言喻的嘆息替我們祈求。
ROM|8|27|那鑒察人心的知道聖靈所體貼的，因為聖靈照著上帝的旨意替聖徒祈求。
ROM|8|28|我們知道，萬事 都互相效力，叫愛上帝的人得益處，就是按他旨意被召的人。
ROM|8|29|因為他所預知的人，他也預定他們效法他兒子的榜樣，使他兒子在許多弟兄中作長子 。
ROM|8|30|他所預定的人，他又召他們來；所召來的人，他又稱他們為義；所稱為義的人，他又叫他們得榮耀。
ROM|8|31|既是這樣，我們對這些事還要怎麼說呢？上帝若幫助我們，誰能抵擋我們呢？
ROM|8|32|上帝既不顧惜自己的兒子，為我們眾人捨了他，豈不也把萬物和他一同白白地賜給我們嗎？
ROM|8|33|誰能控告上帝所揀選的人呢？有上帝稱他們為義了。
ROM|8|34|誰能定他們的罪呢？有基督耶穌 已經死了，而且復活了，現今在上帝的右邊，也替我們祈求。
ROM|8|35|誰能使我們與基督的愛隔絕呢？難道是患難嗎？是困苦嗎？是迫害嗎？是飢餓嗎？是赤身露體嗎？是危險嗎？是刀劍嗎？
ROM|8|36|如經上所記： 「我們為你的緣故終日被殺； 人看我們如將宰的羊。」
ROM|8|37|然而，靠著愛我們的主，在這一切的事上，我們已經得勝有餘了。
ROM|8|38|因為我深信，無論是死，是活，是天使，是掌權的，是有權能的 ，是現在的事，是將來的事，
ROM|8|39|是高處的，是深處的，是別的受造之物，都不能使我們與上帝的愛隔絕，這愛是在我們的主基督耶穌裏的。
ROM|9|1|我在基督裏說真話，不說謊話；我的良心被聖靈感動為我作證。
ROM|9|2|我非常憂愁，心裏時常傷痛。
ROM|9|3|為我弟兄，我骨肉之親，就是自己被詛咒，與基督分離，我也願意。
ROM|9|4|他們是 以色列 人，那兒子的名分、榮耀、諸約、律法的頒佈、敬拜的禮儀、應許都是給他們的。
ROM|9|5|列祖是他們的，基督按肉體說也是從他們出來的。願在萬有之上的上帝被稱頌，直到永遠 。阿們！
ROM|9|6|這不是說上帝的話落了空。因為從 以色列 生的不都是 以色列 人，
ROM|9|7|也不因為是 亞伯拉罕 的後裔就都是他的兒女；惟獨「從 以撒 生的才要稱為你的後裔。」
ROM|9|8|這就是說，肉身所生的兒女不是上帝的兒女，惟獨那應許的兒女才算是後裔。
ROM|9|9|因為所應許的話是這樣：「到明年這時候我要來， 撒拉 必會生一個兒子。」
ROM|9|10|不但如此， 利百加 也是這樣。她從一個人，就是從我們的祖宗 以撒 懷了孕。
ROM|9|11|雙胞胎還沒有生下來，善惡還沒有行出來，為要貫徹上帝揀選人的旨意，
ROM|9|12|不是憑著人的行為，而是憑著那呼召人的，上帝就對 利百加 說：「將來，大的要服侍小的。」
ROM|9|13|正如經上所記：「 雅各 是我所愛的； 以掃 是我所惡的。」
ROM|9|14|這樣，我們要怎麼說呢？難道上帝有甚麼不義嗎？絕對沒有！
ROM|9|15|因他對 摩西 說： 「我要憐憫誰就憐憫誰， 要恩待誰就恩待誰。」
ROM|9|16|由此看來，這不靠人的意願，也不靠人的努力，只靠上帝的憐憫。
ROM|9|17|因為經上有話對法老說：「我將你興起來，特要在你身上彰顯我的權能，為要使我的名傳遍全地。」
ROM|9|18|由此看來，上帝要憐憫誰就憐憫誰，要使誰剛硬就使誰剛硬。
ROM|9|19|這樣，你會對我說：「那麼，他為甚麼還指責人呢？有誰能抗拒他的旨意呢？」
ROM|9|20|你這個人哪，你是誰，竟敢向上帝頂嘴呢？受造之物豈會對造他的說：「你為甚麼把我造成這樣呢？」
ROM|9|21|難道陶匠沒有權從一團泥裏拿一塊做成貴重的器皿，又拿一塊做成卑賤的器皿嗎？
ROM|9|22|倘若上帝要顯明他的憤怒，彰顯他的權能，難道不可多多忍耐寬容那應受憤怒、預備遭毀滅的器皿嗎？
ROM|9|23|這是為了要把他豐盛的榮耀彰顯在那蒙憐憫、早預備得榮耀的器皿上。
ROM|9|24|這器皿也就是我們這些蒙上帝所召的，不但是從 猶太 人中，也是從外邦人中召來的。
ROM|9|25|正如上帝在《何西阿書》上說： 「那本來不是我子民的， 我要稱為『我的子民』； 本來不是蒙愛的， 我要稱為『蒙愛的』。
ROM|9|26|從前在甚麼地方對他們說： 你們不是我的子民， 將來就在那裏稱他們為『永生上帝的兒子』。」
ROM|9|27|關於 以色列 人， 以賽亞 喊著：「雖然 以色列 人多如海沙，得救的將是剩下的餘數，
ROM|9|28|因為主要在地上施行他的話，徹底而又迅速。」
ROM|9|29|又如 以賽亞 先前說過： 「若不是萬軍之主給我們存留餘種， 我們早已變成 所多瑪 ，像 蛾摩拉 一樣了。」
ROM|9|30|這樣，我們要怎麼說呢？那不追求義的外邦人卻獲得了義，就是因信而獲得的義。
ROM|9|31|但 以色列 人追求律法的義，反而達不到律法的義。
ROM|9|32|這是甚麼緣故呢？是因為他們不憑著信心，而是憑著行為，他們正跌在那絆腳石上。
ROM|9|33|就如經上所記： 「我在 錫安 放一塊絆腳的石頭，使人跌倒的磐石； 信靠他的人必不蒙羞。」
ROM|10|1|弟兄們，我心裏所渴望的和向上帝所求的，是要 以色列 人得救。
ROM|10|2|我為他們作證，他們對上帝有熱心，但不是按著真知識。
ROM|10|3|因為不明白上帝的義，想要立自己的義，他們就不服上帝的義了。
ROM|10|4|律法的總結就是基督，使所有信他的人都得著義。
ROM|10|5|論到出於律法的義， 摩西 寫著：「行這些事的人，就必因此得生。」
ROM|10|6|但出於信的義卻如此說：「你不要心裏說：誰要升到天上去呢？（就是說，把基督領下來。）
ROM|10|7|或說：誰要下到陰間去呢？（就是說，把基督從死人中領上來。）」
ROM|10|8|他到底怎麼說呢？ 「這話語就離你近， 就在你口中，在你心裏，」 （就是說，我們傳揚所信的話語。）
ROM|10|9|你若口裏宣認耶穌為主，心裏信上帝叫他從死人中復活，就必得救。
ROM|10|10|因為，人心裏信就可以稱義，口裏宣認就可以得救。
ROM|10|11|經上說：「凡信靠他的人必不蒙羞。」
ROM|10|12|猶太 人和 希臘 人並沒有分別，因為人人都有同一位主，他也厚待求告他的每一個人。
ROM|10|13|因為「凡求告主名的就必得救」。
ROM|10|14|然而，人未曾信他，怎能求告他呢？未曾聽見他，怎能信他呢？沒有傳道的，怎能聽見呢？
ROM|10|15|若沒有奉差遣，怎能傳道呢？如經上所記：「報福音、傳喜信的人，他們的腳蹤何等佳美！」
ROM|10|16|但不是每一個人都聽從福音，因為 以賽亞 說：「主啊，我們所傳的有誰信呢？」
ROM|10|17|可見，信道是從聽道來的，聽道是從基督的話來的。
ROM|10|18|但我要問，人沒有聽見嗎？當然聽見了。 「他們的聲音傳遍全地； 他們的言語傳到地極。」
ROM|10|19|我再問， 以色列 人不知道嗎？先有 摩西 說： 「我要以不成國的激起你們嫉妒； 我要以愚頑的國惹起你們發怒。」
ROM|10|20|又有 以賽亞 放膽說： 「沒有尋找我的，我要讓他們尋見； 沒有求問我的，我要向他們顯現。」
ROM|10|21|關於 以色列 人，他說：「我整天向那悖逆頂嘴的百姓招手。」
ROM|11|1|那麼，我要問，上帝棄絕了他的百姓嗎？絕對沒有！因為我也是 以色列 人， 亞伯拉罕 的後裔，屬 便雅憫 支派的。
ROM|11|2|上帝並沒有棄絕他預先所知道的百姓。你們豈不知道經上論到 以利亞 是怎麼說的呢？他在上帝面前怎樣控告 以色列 人說：
ROM|11|3|「主啊，他們殺了你的先知，拆了你的祭壇，只剩下我一個人，他們還要我的命。」
ROM|11|4|但上帝的指示是怎麼對他說的呢？他說：「我為自己留下七千人，是未曾向 巴力 屈膝的。」
ROM|11|5|現在這時刻也是這樣，照著出於恩典的揀選，還有所留的餘數。
ROM|11|6|既是靠恩典，就不憑行為，不然，恩典就不再是恩典了。
ROM|11|7|那又怎麼說呢？ 以色列 人所尋求的，他們沒有得著。但是蒙揀選的人得著了，其餘的人卻成了頑梗不化的。
ROM|11|8|如經上所記： 「上帝給他們昏沉的靈， 眼睛看不見， 耳朵聽不到， 直到今日。」
ROM|11|9|大衛 也說： 「願他們的宴席變為羅網，變為陷阱， 變為絆腳石，作他們的報應。
ROM|11|10|願他們的眼睛昏花，看不見； 願你時常彎下他們的腰。」
ROM|11|11|那麼，我再問，他們失足是要他們跌倒嗎？絕對不是！因他們的過犯，救恩反而臨到外邦人，要激起他們嫉妒的心。
ROM|11|12|如果他們的過犯成為世界的富足，他們的缺乏成為外邦人的富足，更何況他們全數得救呢？
ROM|11|13|我對你們外邦人說，正因為我是外邦人的使徒，我敬重我的職分，
ROM|11|14|希望可以激起我骨肉之親的嫉妒，好救他們一些人。
ROM|11|15|如果他們被丟棄，世界因而得以與上帝和好；他們被收納，豈不就是從死人中復生嗎？
ROM|11|16|所獻的新麵若聖潔，整個麵團都聖潔了；樹根若聖潔，樹枝也聖潔了。
ROM|11|17|若有幾根枝子被折下來，你這野橄欖枝接上去，同享橄欖根的肥汁，
ROM|11|18|你就不可向舊枝子誇口；若是誇口，該知道不是你托著根，而是根托著你。
ROM|11|19|你會說，那些枝子被折下來是為了使我接上去。
ROM|11|20|不錯。他們因為不信，所以被折下來；你因為信，所以立得住。你不可自高，反要戰戰兢兢。
ROM|11|21|上帝既然不顧惜原來的枝子，豈會顧惜你？
ROM|11|22|可見，上帝又恩慈又嚴厲：對那跌倒的人是嚴厲的；對你是恩慈的，只要你長久在他的恩慈裏，不然，你也要被砍下來。
ROM|11|23|而且，他們若不是長久不信，仍要被接上，因為上帝能夠重新把他們接上去。
ROM|11|24|你是從那天生的野橄欖上砍下來的，尚且違反自然地接在好橄欖上，何況這些原來的枝子豈不更要接在原樹上嗎？
ROM|11|25|弟兄們，我不願意你們不知道這奧祕，恐怕你們自以為聰明。這奧祕就是有一部分 以色列 人是硬心的，等到外邦人的數目添滿了，
ROM|11|26|以色列 全家都要得救。如經上所記： 「必有一位救主從 錫安 出來， 要消除 雅各 家一切不虔不敬。」
ROM|11|27|「這就是我與他們所立的約， 那時我要除去他們的罪。」
ROM|11|28|就福音來說，他們為你們的緣故是仇敵；就揀選來說，他們因列祖的緣故是蒙愛的。
ROM|11|29|因為上帝的恩賜和選召是不會撤回的。
ROM|11|30|你們從前不順服上帝，如今因他們的不順服，你們倒蒙了憐憫。
ROM|11|31|同樣，他們現在也是不順服，叫他們因著施給你們的憐憫，現在 也就蒙憐憫。
ROM|11|32|因為上帝把眾人都圈在不順服中，為的是要憐憫眾人。
ROM|11|33|深哉，上帝的豐富、智慧和知識！ 他的判斷何其難測！ 他的蹤跡何其難尋！
ROM|11|34|誰知道主的心？ 誰作過他的謀士？
ROM|11|35|誰先給了他， 使他後來償還呢？
ROM|11|36|因為萬有都是本於他， 倚靠他，歸於他。 願榮耀歸給他，直到永遠。阿們！
ROM|12|1|所以，弟兄們，我以上帝的慈悲勸你們，將身體獻上當作活祭，是聖潔的，是上帝所喜悅的，你們如此事奉乃是理所當然的 。
ROM|12|2|不要效法這個世界，只要心意更新而變化，叫你們察驗何為上帝的善良、純全、可喜悅的旨意。
ROM|12|3|我憑著所賜我的恩對你們每一位說：不要把自己看得太高，要照著上帝所分給各人的信心來衡量，看得合乎中道。
ROM|12|4|正如我們一個身子上有好些肢體，肢體也不都有一樣的用處。
ROM|12|5|這樣，我們許多人在基督裏是一個身體，互相聯絡作肢體。
ROM|12|6|按著所得的恩典，我們各有不同的恩賜：或說預言，要按著信心的程度說預言；
ROM|12|7|或服事的，要專一服事；或教導的，要專一教導；
ROM|12|8|或勸勉的，要專一勸勉；施捨的，要誠實；治理的，要殷勤；憐憫人的，要樂意。
ROM|12|9|愛，不可虛假；惡，要厭惡；善，要親近。
ROM|12|10|愛弟兄，要相親相愛；恭敬人，要彼此推讓；
ROM|12|11|殷勤，不可懶惰。要靈裏火熱；常常服侍主。
ROM|12|12|在盼望中要喜樂；在患難中要忍耐；禱告要恆切。
ROM|12|13|聖徒有缺乏，要供給；異鄉客，要殷勤款待。
ROM|12|14|要祝福迫害你們 的，要祝福，不可詛咒。
ROM|12|15|要與喜樂的人同樂；要與哀哭的人同哭。
ROM|12|16|要彼此同心，不要心高氣傲，倒要俯就卑微的人。不要自以為聰明。
ROM|12|17|不要以惡報惡，眾人以為美的事要留心去做。
ROM|12|18|若是可行，總要盡力與眾人和睦。
ROM|12|19|各位親愛的，不要自己伸冤，寧可給主的憤怒留地步，因為經上記著：「主說：『伸冤在我，我必報應。』」
ROM|12|20|不但如此，「你的仇敵若餓了，就給他吃；若渴了，就給他喝。因為你這樣做，就是把炭火堆在他的頭上。」
ROM|12|21|不要被惡所勝，反要以善勝惡。
ROM|13|1|在上有權柄的，人人要順服，因為沒有權柄不是來自上帝的。掌權的都是上帝所立的。
ROM|13|2|所以，抗拒掌權的就是抗拒上帝所立的；抗拒的人必自招審判。
ROM|13|3|作官的原不是要使行善的懼怕，而是要使作惡的懼怕。你願意不懼怕掌權的嗎？只要行善，你就可得他的稱讚；
ROM|13|4|因為他是上帝的用人，是與你有益的。你若作惡，就該懼怕，因為他不是徒然佩劍；他是上帝的用人，為上帝的憤怒，報應作惡的。
ROM|13|5|所以，你們必須順服，不但是因上帝的憤怒，也是因著良心。
ROM|13|6|你們納糧也為這個緣故，因他們是上帝的僕役，專管這事。
ROM|13|7|凡人所當得的，就給他。當得糧的，給他納糧；當得稅的，給他上稅；當懼怕的，懼怕他；當恭敬的，恭敬他。
ROM|13|8|你們除了彼此相愛，對任何人都不可虧欠甚麼，因為那愛人的就成全了律法。
ROM|13|9|那不可姦淫，不可殺人，不可偷盜，不可貪婪，或別的誡命，都包括在「愛鄰 如己」這一句話之內了。
ROM|13|10|愛是不對鄰人作惡，所以愛就成全了律法。
ROM|13|11|還有，你們要知道，現在正是該從睡夢中醒來的時候了；因為我們得救，現在比初信的時候更近了。
ROM|13|12|黑夜已深，白晝將近。所以我們該除去暗昧的行為，帶上光明的兵器。
ROM|13|13|行事為人要端正，好像在白晝行走。不可荒宴醉酒；不可好色淫蕩；不可紛爭嫉妒。
ROM|13|14|總要披戴主耶穌基督，不要只顧滿足肉體，去放縱私慾。
ROM|14|1|信心軟弱的，你們要接納，不同的意見，不要爭論。
ROM|14|2|有人信甚麼都可吃；但那軟弱的，只吃蔬菜。
ROM|14|3|吃的人不可輕看不吃的人；不吃的人也不可評斷吃的人，因為上帝已經接納他了。
ROM|14|4|你是誰，竟評斷別人的僕人呢？他或站立或跌倒，自有他的主人在，而且他也必會站立，因為主能使他站穩。
ROM|14|5|有人看這日比那日強；有人看日日都是一樣。只是各人要在自己的心意上堅定。
ROM|14|6|守日子的人是為主守的。吃的人是為主吃的，因他感謝上帝；不吃的人是為主不吃的，他也感謝上帝。
ROM|14|7|我們沒有一個人為自己而活，也沒有一個人為自己而死。
ROM|14|8|我們若活，是為主而活；我們若死，是為主而死。所以，我們或死或活總是主的人。
ROM|14|9|為此，基督死了，又活了，為要作死人和活人的主。
ROM|14|10|可是你，你為甚麼評斷弟兄呢？你又為甚麼輕看弟兄呢？因我們都要站在上帝的審判臺前。
ROM|14|11|經上寫著： 「主說，我指著我的永生起誓： 萬膝必向我跪拜； 萬口必稱頌上帝。」
ROM|14|12|這樣看來，我們各人一定要把自己的事在上帝面前 交代。
ROM|14|13|所以，我們不可再彼此評斷，寧可決意不給弟兄放置障礙或絆腳石。
ROM|14|14|我憑著主耶穌確知深信，凡物本來沒有不潔淨的，除非人以為不潔淨的，在他就不潔淨了。
ROM|14|15|你若因食物使弟兄憂愁，就不是按著愛心行事。基督已經為他死，你不可因你的食物使他敗壞。
ROM|14|16|所以，不可讓你們的善被人毀謗。
ROM|14|17|因為上帝的國不在乎飲食，而在乎公義、和平及聖靈中的喜樂 。
ROM|14|18|凡這樣服侍基督的，就為上帝所喜悅，又為人所讚許。
ROM|14|19|所以，我們務要追求 和平與彼此造就的事。
ROM|14|20|不可因食物毀壞上帝的工作。一切都是潔淨的，但有人因食物使人跌倒，這在他就是惡了。
ROM|14|21|無論是吃肉是喝酒，是甚麼別的事，使弟兄跌倒，一概不做，才是善的。
ROM|14|22|你有信心，就要在上帝面前持守。人能在自己以為可行的事上不自責就有福了。
ROM|14|23|若有人疑惑而吃的，就被定罪，因為他吃不是出於信心。凡不出於信心的都是罪。
ROM|15|1|我們堅強的人應該分擔不堅強的人的軟弱，不求自己的喜悅。
ROM|15|2|我們各人務必要讓鄰人喜悅，使他得益處，得造就。
ROM|15|3|因為基督也不求自己的喜悅，如經上所記：「辱罵你的人的辱罵都落在我身上。」
ROM|15|4|從前所寫的聖經都是為教導我們寫的，要使我們藉著忍耐和因聖經所生的安慰，得著盼望。
ROM|15|5|但願賜忍耐和安慰的上帝使你們彼此同心，效法基督耶穌，
ROM|15|6|為使你們同心同聲榮耀我們主耶穌基督的父上帝！
ROM|15|7|所以，你們要彼此接納，如同基督接納你們一樣，歸榮耀給上帝。
ROM|15|8|我說，基督是為上帝真理作了受割禮的人的執事，要證實所應許列祖的話，
ROM|15|9|並使外邦人，因他的憐憫，榮耀上帝。如經上所記： 「因此，我要在外邦中稱頌你， 歌頌你的名。」
ROM|15|10|又說： 「外邦人哪，你們要與主的子民一同歡樂。」
ROM|15|11|又說： 「列邦啊，你們要讚美主！ 萬民哪，你們都要頌讚他！」
ROM|15|12|又有 以賽亞 說： 「將來有 耶西 的根， 就是那興起來要治理列邦的； 外邦人要仰望他。」
ROM|15|13|願賜盼望的上帝，因你們的信把各樣的喜樂、平安 充滿你們的心，使你們藉著聖靈的能力大有盼望！
ROM|15|14|我的弟兄們，我本人也深信你們自己充滿良善，有各種豐富的知識，也能彼此勸戒。
ROM|15|15|但我更大膽寫信給你們，是要在一些事上提醒你們，我因上帝所賜我的恩，
ROM|15|16|使我為外邦人作基督耶穌的僕役，作上帝福音的祭司，使所獻上的外邦人因著聖靈成為聖潔，可蒙悅納。
ROM|15|17|所以，有關上帝面前的事奉，我在基督耶穌裏是有可誇的。
ROM|15|18|除了基督藉我做的那些事，我甚麼都不敢提，只提他藉我的言語作為，用神蹟奇事的能力，並上帝的靈 的能力，使外邦人順服；甚至我從 耶路撒冷 ，直轉到 以利哩古 ，到處傳了基督的福音。
ROM|15|19|
ROM|15|20|這樣，我立了志向，不在基督的名已經傳揚過的地方傳福音，免得建造在別人的根基上；
ROM|15|21|卻如經上所記： 「未曾傳給他們的，他們必看見； 未曾聽見過的事，他們要明白。」
ROM|15|22|因此我多次被攔阻，不能到你們那裏去。
ROM|15|23|但如今，在這一帶再沒有可傳的地方，而且這許多年來，我迫切想去你們那裏，
ROM|15|24|盼望到 西班牙 去的時候經過，得見你們，先與你們彼此交往，心裏稍得滿足，然後蒙你們為我送行。
ROM|15|25|但如今我要到 耶路撒冷 去，供應聖徒的需要。
ROM|15|26|因為 馬其頓 和 亞該亞 人樂意湊出一些捐款給 耶路撒冷 聖徒中的窮人。
ROM|15|27|這固然是他們樂意的，其實也算是所欠的債；因為外邦人既然分享了他們靈性上的好處，就當把肉體上的需用供給他們。
ROM|15|28|等我辦完了這事，把這筆捐款 交付給他們，我就要路過你們那裏，到 西班牙 去。
ROM|15|29|我也知道去你們那裏的時候，我將帶著基督豐盛的恩典去。
ROM|15|30|弟兄們，我藉著我們的主耶穌基督，又藉著聖靈的愛，勸你們與我一同竭力為我祈求上帝，
ROM|15|31|使我脫離在 猶太 不順從的人，也讓我在 耶路撒冷 的事奉可蒙聖徒悅納，
ROM|15|32|並使我照著上帝的旨意歡歡喜喜地到你們那裏，與你們同得安息。
ROM|15|33|願賜平安的上帝與你們眾人同在。阿們！
ROM|16|1|我對你們推薦我們的姊妹 非比 ，她是 堅革哩 教會中的執事。
ROM|16|2|請你們在主裏用合乎聖徒的方式來接待她。她在任何事上需要你們幫助，你們就幫助她；因她素來幫助許多人，也幫助了我。
ROM|16|3|請向 百基拉 和 亞居拉 問安。他們在基督耶穌裏作我的同工，
ROM|16|4|也為我的性命把自己的生死置之度外；不但我感謝他們，就是外邦的眾教會也感謝他們。
ROM|16|5|又向在他們家中的教會問安。向我所親愛的 以拜尼土 問安，他是 亞細亞 歸於基督的初結果子。
ROM|16|6|又向 馬利亞 問安，她為你們非常辛勞。
ROM|16|7|又向與我一同坐監的親戚 安多尼古 和 猶尼亞 問安，他們在使徒中是有名望的，也是比我先在基督裏的。
ROM|16|8|又向我在主裏面所親愛的 暗伯利 問安。
ROM|16|9|又向我們在基督裏的同工 耳巴奴 和我所親愛的 士大古 問安。
ROM|16|10|又向在基督裏經過考驗的 亞比利 問安。向 亞利多布 家裏的人問安。
ROM|16|11|又向我親戚 希羅天 問安。向 拿其數 家在主裏的人問安。
ROM|16|12|又向為主辛勞的 土非拿 和 土富撒 問安。向所親愛、為主非常辛勞的 彼息 問安。
ROM|16|13|又向在主裏蒙揀選的 魯孚 和他母親問安，他的母親就是我的母親。
ROM|16|14|又向 亞遜其土 、 弗勒干 、 黑米 、 八羅巴 、 黑馬 ，和跟他們在一起的弟兄們問安。
ROM|16|15|又向 非羅羅古 和 猶利亞 ， 尼利亞 和他姊妹， 阿林巴 和跟他們在一起的眾聖徒問安。
ROM|16|16|你們要以聖潔的吻彼此問安。基督的眾教會都向你們問安！
ROM|16|17|弟兄們，那些離間你們、使你們跌倒、違背所學之道的人，我勸你們要留意躲避他們。
ROM|16|18|因為這樣的人不服侍我們的主基督，只服侍自己的肚腹，用花言巧語誘惑老實人的心。
ROM|16|19|你們的順服已經傳於眾人，所以我為你們歡喜；但我願你們在善上聰明，在惡上愚拙。
ROM|16|20|那賜平安 的上帝快要把撒但踐踏在你們腳下。願我們主耶穌基督的恩與你們同在！
ROM|16|21|我的同工 提摩太 ，和我的親戚 路求 、 耶孫 、 所西巴德 ，向你們問安。
ROM|16|22|我這代筆寫信的 德提 ，在主裏向你們問安。
ROM|16|23|那接待我，也接待全教會的 該猶 ，向你們問安。城裏的財務官 以拉都 和弟兄 括土 向你們問安。
ROM|16|24|
ROM|16|25|惟有上帝能照我所傳的福音和所講的耶穌基督，並照歷代以來隱藏的奧祕的啟示，堅固你們。
ROM|16|26|這奧祕如今顯示出來，而且按著永生上帝的命令，藉眾先知的書指示萬民，使他們因信而順服。
ROM|16|27|願榮耀，藉著耶穌基督，歸給獨一全智的上帝，直到永遠。阿們！
1COR|1|1|奉上帝旨意，蒙召作基督耶穌使徒的 保羅 ，同弟兄 所提尼 ，
1COR|1|2|寫信給在 哥林多 上帝的教會—就是在基督耶穌裏成聖、蒙召作聖徒的—以及所有在各處求告我主耶穌基督之名的人。基督是他們的主，也是我們的主。
1COR|1|3|願恩惠、平安 從我們的父上帝並主耶穌基督歸給你們！
1COR|1|4|我常為你們感謝我的上帝，因上帝在基督耶穌裏所賜給你們的恩惠。
1COR|1|5|因為你們在他裏面凡事富足，具有各種口才、各樣知識，
1COR|1|6|正如我為基督作的見證在你們心裏得以堅固，
1COR|1|7|以致你們在恩賜上一無欠缺，切切等候我們主耶穌基督的顯現。
1COR|1|8|他也必堅固你們到底，使你們在我們主耶穌基督 的日子無可指責。
1COR|1|9|上帝是信實的，他呼召你們好與他兒子—我們的主耶穌基督—共享團契。
1COR|1|10|弟兄們，我藉我們主耶穌基督的名勸你們說話要一致。你們中間不可分裂，只要一心一意彼此團結。
1COR|1|11|我的弟兄們， 革來 氏家裏的人曾對我提起你們，說你們中間有紛爭。
1COR|1|12|我的意思是，你們各人說：「我是屬 保羅 的」；「我是屬 亞波羅 的」；「我是屬 磯法 的」；「我是屬基督的。」
1COR|1|13|基督是分裂的嗎？ 保羅 為你們釘了十字架嗎？你們是奉 保羅 的名受了洗嗎？
1COR|1|14|我感謝上帝 ，除了 基利司布 和 該猶 以外，我沒有給你們中的任何一個人施洗，
1COR|1|15|免得有人說你們是奉我的名受洗的。
1COR|1|16|我曾為 司提法那 家施過洗；此外我已記不清有沒有給別人施過洗。
1COR|1|17|因為基督差遣我不是為施洗，而是為傳福音；並不是用智慧的言論，免得基督的十字架落了空。
1COR|1|18|因為十字架的道理，在那滅亡的人是愚拙，在我們得救的人卻是上帝的大能。
1COR|1|19|就如經上所記： 「我要摧毀智慧人的智慧， 廢棄聰明人的聰明。」
1COR|1|20|智慧人在哪裏？文士在哪裏？這世上的辯士在哪裏？上帝豈不是已使這世上的智慧變成愚拙了嗎？
1COR|1|21|既然世人憑自己的智慧不認識上帝，上帝就本著自己的智慧樂意藉著人所傳愚拙的話拯救那些信的人。
1COR|1|22|猶太 人要的是神蹟， 希臘 人求的是智慧，
1COR|1|23|我們卻是傳被釘十字架的基督，這對 猶太 人是絆腳石，對外邦人是愚拙；
1COR|1|24|但對那蒙召的，無論是 猶太 人、 希臘 人，基督總是上帝的大能，上帝的智慧。
1COR|1|25|因為，上帝的愚拙總比人智慧；上帝的軟弱總比人強壯。
1COR|1|26|弟兄們哪，想一想你們的蒙召，按著人的觀點，有智慧的不多，有能力的不多，有尊貴地位的也不多。
1COR|1|27|但是，上帝揀選了世上愚拙的，為了使有智慧的羞愧；又揀選了世上軟弱的，為了使強壯的羞愧。
1COR|1|28|上帝也揀選了世上卑賤的，被人厭惡的，以及那一無所有的，為要廢掉那樣樣都有的，
1COR|1|29|使凡血肉之軀的，在上帝面前，一個也不能自誇。
1COR|1|30|但你們得以在基督耶穌裏是本乎上帝，他使基督成為我們的智慧，成為公義、聖潔、救贖。
1COR|1|31|如經上所記：「要誇耀的，該誇耀主。」
1COR|2|1|弟兄們，從前我到你們那裏去，並沒有用高言大智對你們宣講上帝的奧祕。
1COR|2|2|因為我曾定了主意，在你們中間不知道別的，只知道耶穌基督並他釘十字架。
1COR|2|3|我在你們那裏時，又軟弱，又懼怕，又戰戰兢兢。
1COR|2|4|我說的話、講的道不是用委婉智慧的言語 ，而是以聖靈的大能來證明，
1COR|2|5|為要使你們的信不靠著人的智慧，而是靠著上帝的大能。
1COR|2|6|然而，在成熟的人中，我們也講智慧，但不是今世的智慧，也不是今世有權有位、將要滅亡的人的智慧。
1COR|2|7|我們講的是從前隱藏的、上帝奧祕的智慧，就是上帝在萬世以前預定使我們得榮耀的智慧；
1COR|2|8|這智慧，今世有權有位的人沒有一個知道，若知道，他們就不會把榮耀的主釘在十字架上了。
1COR|2|9|如經上所記： 「上帝為愛他的人所預備的 是眼睛未曾看見，耳朵未曾聽見， 人心也未曾想到的。」
1COR|2|10|只有上帝藉著聖靈把這事向我們顯明了；因為聖靈參透萬事，就是上帝深奧的事也參透了。
1COR|2|11|除了在人裏頭的靈，誰知道人的事？照樣，除了上帝的靈，也沒有人知道上帝的事。
1COR|2|12|我們所領受的並不是世上的靈，而是從上帝來的靈，為使我們知道上帝把恩賜賞給我們的事。
1COR|2|13|我們也講說這些事，不是用人的智慧所教的言語，而是用聖靈所教的言語，用屬靈的話解釋屬靈的事 。
1COR|2|14|然而，屬血氣的人不接受上帝的靈的事，他反倒以這為愚拙，並且他不能了解，因為這些事惟有屬靈的人才能領悟。
1COR|2|15|屬靈的人能看透萬事，卻沒有一人能看透他。
1COR|2|16|「誰曾知道主的心？ 誰會教導他？」 至於我們，我們有基督的心。
1COR|3|1|弟兄們，我從前對你們說話，還不能把你們當作屬靈的，只能把你們當作屬肉體的，你們在基督裏僅是嬰孩。
1COR|3|2|我用奶餵你們，沒有用飯餵你們，因為那時你們不能吃。就是如今還是不能，
1COR|3|3|因為你們仍是屬肉體的。你們中間有嫉妒、紛爭，這豈不是屬乎肉體，照著世人的樣子生活嗎？
1COR|3|4|有人說：「我是屬 保羅 的」；有人說：「我是屬 亞波羅 的」；這樣你們豈不是和世人一樣嗎？
1COR|3|5|亞波羅 算甚麼？ 保羅 算甚麼？我們都是上帝的執事，藉著我們，你們信了；這不過是照著主給各人的恩賜去做罷了。
1COR|3|6|我栽種了， 亞波羅 澆灌了，惟有上帝使它生長。
1COR|3|7|可見，栽種的算不了甚麼，澆灌的也算不了甚麼；惟有上帝能使它生長。
1COR|3|8|栽種的和澆灌的都是一樣，但將來各人要照自己的勞苦得到自己的報酬。
1COR|3|9|因為我們是上帝的同工，而你們是上帝的田地、上帝的房屋。
1COR|3|10|我照上帝所給我的恩典，好像一個聰明的工頭，立好了根基，別人在上面建造；只是各人要謹慎怎樣在上面建造。
1COR|3|11|因為，那已經立好的根基就是耶穌基督，此外沒有人能立別的根基。
1COR|3|12|若有人用金銀、寶石，草木、禾秸，在這根基上建造，
1COR|3|13|各人的工程必將顯露，因為那日子要將它顯明，有火把它暴露出來，這火要試煉各人的工程怎樣。
1COR|3|14|人在那根基上所建造的工程若能保得住，他將要得賞賜。
1COR|3|15|人的工程若被燒了，他將損失，雖然他自己將得救，卻要像從火裏經過一樣。
1COR|3|16|難道不知你們是上帝的殿，上帝的靈住在你們裏面嗎？
1COR|3|17|若有人毀壞上帝的殿，上帝一定要毀滅那人；因為上帝的殿是神聖的，這殿就是你們。
1COR|3|18|誰都不可自欺。你們中間若有人自以為在今世有智慧，倒不如變為愚拙，好成為有智慧的。
1COR|3|19|因為這世界的智慧在上帝看來是愚拙的。如經上記著： 「主使有智慧的人中了自己的詭計；」
1COR|3|20|又說： 「主知道智慧人的意念， 因為它們是虛妄的。」
1COR|3|21|所以，無論誰都不可誇耀人；因為萬有都是你們的，
1COR|3|22|或 保羅 ，或 亞波羅 ，或 磯法 ，或世界，或生，或死，或現今的事，或將來的事，全是你們的，
1COR|3|23|而你們是屬基督的，基督是屬上帝的。
1COR|4|1|人應該把我們看為基督的執事，為上帝的奧祕的管家。
1COR|4|2|所求於管家的，是要他忠心。
1COR|4|3|我被你們評斷，或被別人評斷，我都以為是極小的事；連我自己也不評斷自己。
1COR|4|4|雖然我不覺得自己有錯，卻也不能因此判為無罪；審斷我的是主。
1COR|4|5|所以，時候未到，在主來以前甚麼都不要評斷，他要照出暗中的隱情，揭發人的動機。那時，各人要從上帝那裏得著稱讚。
1COR|4|6|弟兄們，為你們的緣故，我拿這些事應用到我自己和 亞波羅 身上，讓你們從我們學到「不可過於聖經所記」這話的意思，免得你們自高自大，看重這個，看輕那個。
1COR|4|7|使你與人不同的是誰呢？你所有的有哪一個不是領受的呢？若是領受的，為何自誇，彷彿不是領受的呢？
1COR|4|8|你們已經飽足了，已經富足了，用不著我們，自己就作王了。我願意你們果真作王，讓我們也可以與你們一同作王！
1COR|4|9|我想，上帝把我們作使徒的明顯地列在末後，好像定死罪的囚犯，因為我們成了一臺戲，給世界、天使和眾人觀看。
1COR|4|10|我們為基督的緣故成為愚拙的；你們在基督裏倒是聰明的。我們軟弱，你們倒強壯；你們有榮耀，我們倒被藐視。
1COR|4|11|直到如今，我們還是又飢又渴，又赤身露體，又挨打，又到處漂泊，
1COR|4|12|並且勞碌，親手做工；被人咒罵，我們就祝福；被人迫害，我們就忍受；
1COR|4|13|被人毀謗，我們就勸導。直到如今，人還把我們看作世上的污穢，萬物中的渣滓。
1COR|4|14|我寫這些話，不是要使你們羞愧，而是要警戒你們，好像我所愛的兒女一樣。
1COR|4|15|雖然你們在基督裏有無數的導師，卻沒有許多父親，因我是在基督耶穌裏用福音生了你們。
1COR|4|16|所以，我求你們要效法我。
1COR|4|17|因此，我已差 提摩太 到你們那裏去。他在主裏面是我親愛和忠心的兒子；他要提醒你們，我在基督耶穌 裏怎樣行事為人，在各處各教會中怎樣教導人。
1COR|4|18|有些人以為我不到你們那裏去而自高自大。
1COR|4|19|但是，主若准許，我會很快到你們那裏去；我所要知道的，不是那些自高自大者的言語，而是他們的權能。
1COR|4|20|因為上帝的國不在乎言語，而在乎權能。
1COR|4|21|你們願意怎麼樣呢？要我帶著棍子到你們那裏去呢，還是帶著慈愛溫柔的心呢？
1COR|5|1|我確實聽說在你們中間有淫亂的事；這種淫亂連外邦人中也沒有，就是有人和他的繼母同居。
1COR|5|2|你們還自高自大！你們不是該覺得痛心，把做這事的人從你們中間趕出去嗎？
1COR|5|3|我人雖然不在你們那裏，心卻在你們那裏，好像親自與你們同在。我奉我們主耶穌 的名，已經判斷了做這事的人。你們聚會的時候，我的心和你們同在。你們藉著我們主耶穌的權能，
1COR|5|4|
1COR|5|5|要把這樣的人交給撒但，使他的肉體敗壞，好讓他的靈魂在主的日子可以得救。
1COR|5|6|你們這樣自誇是不好的。你們不知道一點麵酵能使全團發起來嗎？
1COR|5|7|既然你們是無酵的麵，要把舊酵除淨，好使你們成為新團；因為我們逾越節的羔羊—基督已經被殺獻為祭牲了。
1COR|5|8|所以，我們來守這節，不可用舊酵，就是不可用惡毒、邪惡的酵，只用純潔真實的無酵餅。
1COR|5|9|我先前寫信告訴過你們，不可與淫亂的人交往。
1COR|5|10|此話不是泛指這世上所有行淫亂的，或貪婪的，勒索的，或拜偶像的；若是這樣，你們非離開這世界不可。
1COR|5|11|但現在，我寫信告訴你們，若有稱為弟兄的人卻仍犯淫亂，或貪婪，或拜偶像，或辱罵，或醉酒，或勒索，這樣的人不可跟他交往，就是跟他吃飯都不可以。
1COR|5|12|因為審判教外的人與我何干？教內的人豈不是你們要審判嗎？
1COR|5|13|至於外人有上帝審判他們。如經上說：「要從你們中間把那邪惡的人趕出去。」
1COR|6|1|你們中間有彼此爭吵的事，怎敢告到不義的人面前，而不告到聖徒面前呢？
1COR|6|2|你們豈不知聖徒要審判世界嗎？若世界要受你們的審判，難道你們不配審判這最小的事嗎？
1COR|6|3|你們豈不知我們要審判天使嗎？何況今生的事呢！
1COR|6|4|既是這樣，你們若有今生當審判的事，會讓教會所輕看的人來審判嗎？
1COR|6|5|我說這話是要使你們慚愧。難道你們中間沒有一個有智慧的人能審斷弟兄中的事嗎？
1COR|6|6|你們竟然有弟兄去告弟兄，而且告到不信主的人面前。
1COR|6|7|你們彼此告狀，這已經是你們的大錯了。為甚麼不情願受冤屈呢？為甚麼不情願吃虧呢？
1COR|6|8|你們反倒去冤枉人，虧負人，況且所冤枉所虧負的就是弟兄。
1COR|6|9|你們豈不知不義的人不能承受上帝的國嗎？不要自欺！無論是淫亂的、拜偶像的、姦淫的、作娼妓 的，親男色的、
1COR|6|10|偷竊的、貪婪的、醉酒的、辱罵的、勒索的，都不能承受上帝的國。
1COR|6|11|從前你們中間也有人是這樣；但現在你們奉主耶穌基督 的名，並藉著我們上帝的靈，已經洗淨，已經成聖，已經稱義了。
1COR|6|12|「凡事我都可行」，但不是凡事都有益處。「凡事我都可行」，但無論哪一件，我都不受它的轄制。
1COR|6|13|「食物是為肚腹，肚腹是為食物」；但上帝要使這兩樣都毀壞。身體不是為淫亂，而是為主；主也是為身體。
1COR|6|14|上帝已經使主復活，也要用他自己的能力使我們復活。
1COR|6|15|你們豈不知道你們的身體是基督的肢體嗎？我可以把基督的肢體作為娼妓的肢體嗎？絕對不可！
1COR|6|16|你們豈不知道與娼妓苟合的，就是與她成為一體嗎？因為主說：「二人要成為一體。」
1COR|6|17|但與主聯合的，就是與主成為一靈。
1COR|6|18|你們要遠避淫行。人所犯的，無論甚麼罪，都在身體以外；惟有行淫的，是得罪自己的身體。
1COR|6|19|你們豈不知道你們的身體是聖靈的殿嗎？這聖靈是從上帝而來，住在你們裏面的。而且你們不是屬自己的人，
1COR|6|20|因為你們是重價買來的。所以，要在你們的身體上榮耀上帝。
1COR|7|1|關於你們信上所提的事，男人不親近女人倒好。
1COR|7|2|但為了避免淫亂的事，男人當各有自己的妻子，女人也當各有自己的丈夫。
1COR|7|3|丈夫對妻子要盡本分；妻子對丈夫也要如此。
1COR|7|4|妻子對自己的身體沒有主張的權柄，權柄在丈夫；丈夫對自己的身體也沒有主張的權柄，權柄在妻子。
1COR|7|5|夫妻不可忽略對方的需求，除非為了要專心禱告，在兩相情願下暫時分房；以後仍要同房，免得撒但趁著你們情不自禁而引誘你們。
1COR|7|6|我說這話是出於容忍，不是命令。
1COR|7|7|我願眾人像我一樣；但是各人都有來自上帝的恩賜，一個是這樣，一個是那樣。
1COR|7|8|我對沒有嫁娶的和寡婦說，他們若能維持獨身像我一樣就好。
1COR|7|9|但他們若不能自制，就應該嫁娶，與其慾火攻心，倒不如結婚為妙。
1COR|7|10|至於那已經嫁娶的，我吩咐他們—其實不是我，而是主吩咐的：妻子不可離開丈夫，
1COR|7|11|若是離開了，不可再嫁，不然要跟丈夫復和；丈夫也不可離棄妻子。
1COR|7|12|我對其餘的人說—是我，不是主說—倘若某弟兄有不信的妻子，妻子也情願和他一起生活，他就不可離棄妻子。
1COR|7|13|妻子有不信的丈夫，丈夫也情願和她一起生活，她就不可離棄丈夫。
1COR|7|14|因為不信的丈夫會因著妻子成了聖潔；不信的妻子也會因著丈夫 成了聖潔。不然，你們的兒女就不潔淨了，但現在他們是聖潔的。
1COR|7|15|倘若那不信的人要離開，就由他離開吧！無論是弟兄是姊妹，遇著這樣的事都不必拘束。上帝召你們原是要你們和睦。
1COR|7|16|你這作妻子的怎麼知道不能救你的丈夫呢？你這作丈夫的怎麼知道不能救你的妻子呢？
1COR|7|17|無論如何，要照主所分給各人的恩賜和上帝所召各人的情況生活。我在各教會裏都是這樣規定的。
1COR|7|18|有人受割禮後才蒙召，他就不必除去割禮的記號。有人未受割禮前蒙召，他就不必受割禮。
1COR|7|19|受割禮算不了甚麼，不受割禮也算不了甚麼，只要謹守上帝的誡命就是了。
1COR|7|20|各人蒙召的時候是甚麼身份，要守住這身份。
1COR|7|21|你是作奴隸時蒙召的嗎？不要介意；若能獲得自由，就爭取自由更好。
1COR|7|22|因為，蒙主呼召的奴僕是主所釋放的人；蒙主呼召的自由之人是基督的奴僕。
1COR|7|23|你們是重價買來的；不要作人的奴僕。
1COR|7|24|弟兄們，你們各人蒙召的時候是甚麼身份，要在上帝面前守住這身份。
1COR|7|25|關於未婚女子，我沒有主的命令，但我既蒙主憐憫、作為一個可信靠的人，把自己的意見告訴你們。
1COR|7|26|因現今的艱難，據我看來，人不如安於現狀。
1COR|7|27|你已經有了妻子，就不要求擺脫；你還沒有妻子，就不要想娶妻。
1COR|7|28|你若娶妻，並不是犯罪；未婚女子若出嫁，也不是犯罪。然而，這等人會遭受肉身上的苦難，我寧願你們免受這苦難。
1COR|7|29|弟兄們，我是說：時候不多了。從此以後，那有妻子的，要像沒有一樣；
1COR|7|30|哀哭的，不像在哀哭；快樂的，不像在快樂；購買的，像一無所得；
1COR|7|31|享受這世界的，不像在享受這世界；因為這世界的局面將要過去了。
1COR|7|32|我願你們一無掛慮。沒有結婚的是為主的事掛慮，想怎樣令主喜悅；
1COR|7|33|結了婚的是為世上的事掛慮，想怎樣讓妻子喜悅，
1COR|7|34|於是，他就分心了。沒有結婚的和未婚的女子是為主的事掛慮，為要身體和心靈都聖潔；已經出嫁的是為世上的事掛慮，想怎樣讓丈夫喜悅。
1COR|7|35|我說這話是為你們的益處，不是要限制你們，而是要你們做合宜的事，得以不分心地對主忠誠。
1COR|7|36|若有人認為自己待他的女兒 不合宜，女兒也過了適婚年齡 ，他可以隨意處理，不算有罪，讓兩人結婚就是了。
1COR|7|37|倘若有人心裏堅定，沒有不得已的事，並且由得自己作主，心裏又決定了不讓女兒結婚 ，這樣做也好。
1COR|7|38|這樣看來，讓自己的女兒結婚 固然是好，不讓她結婚更好。
1COR|7|39|丈夫活著的時候，妻子是受約束的；丈夫若長眠了，妻子就自由了，可以隨意再嫁，只是要嫁給主裏面的人。
1COR|7|40|然而，按我的意見，她若能守節就更有福氣。我想我自己也有上帝的靈的感動。
1COR|8|1|關於祭過偶像的食物，我們曉得「我們都有知識」，但知識使人自高自大，惟有愛心能造就人。
1COR|8|2|若有人自以為知道甚麼，他其實仍不知道他所應當知道的。
1COR|8|3|若有人愛上帝，他就是上帝所認識的人了。
1COR|8|4|關於吃祭過偶像的食物，我們知道「偶像在世上算不得甚麼」；也知道「上帝只有一位，沒有別的」。
1COR|8|5|雖然在天上或地上有許多所謂的神明，就如他們中間有許多的神明，許多的主，
1COR|8|6|但是我們只有一位上帝，就是父，萬物都出於他，我們也歸於他；並只有一位主，就是耶穌基督，萬物都是藉著他而有，我們也是藉著他而有。
1COR|8|7|可是，不是人人都有這知識。有人到現在因拜慣了偶像，仍以為所吃的是祭過偶像的食物；既然他們的良心軟弱，也就污穢了。
1COR|8|8|其實，食物不能使我們更接近上帝，因為我們不吃也無損，吃也無益。
1COR|8|9|可是，你們要謹慎，免得你們這自由竟成了軟弱人的絆腳石。
1COR|8|10|若有人見你這有知識的在偶像的廟裏坐席，而這人的良心是軟弱的，他豈不放膽去吃那祭過偶像的食物嗎？
1COR|8|11|因此，基督為他死的那軟弱弟兄，也就因你的知識沉淪了。
1COR|8|12|你們這樣得罪弟兄，傷了他們軟弱的良心，就是得罪基督。
1COR|8|13|所以，食物若使我的弟兄跌倒，我就永遠不吃肉，免得使我的弟兄跌倒了。
1COR|9|1|我不是自由的嗎？我不是使徒嗎？我不是見過我們的主耶穌嗎？你們不是我在主裏面工作的成果嗎？
1COR|9|2|假若對別人來說，我不是使徒，對你們來說，我總是使徒；因為你們在主裏正是我作使徒的印證。
1COR|9|3|對那些質問我的人，這就是我的答辯。
1COR|9|4|難道我們沒有權利靠著傳福音吃喝嗎？
1COR|9|5|難道我們沒有權利帶著信主的妻子一起出入，如同其餘的使徒，和主的兄弟們，和 磯法 一樣嗎？
1COR|9|6|只有我和 巴拿巴 沒有權利不做工嗎？
1COR|9|7|有誰當兵而自備糧餉呢？有誰栽葡萄園而不吃園裏的果子呢？有誰牧養牛羊而不喝牛羊的奶呢？
1COR|9|8|我說這些話豈是照一般人的看法？律法不也是這樣說嗎？
1COR|9|9|就如 摩西 的律法記著：「牛在踹穀的時候，不可籠住牠的嘴。」難道上帝所掛念的是牛嗎？
1COR|9|10|他不全是為我們說的嗎？的確是為我們說的！因為耕種的要存著指望去耕種；收割的也要存著分享穀物的指望去收割。
1COR|9|11|我們既然把屬靈的種子撒在你們中間，若從你們收取養生之物，這還算大事嗎？
1COR|9|12|假如別人在你們身上享有這權利，何況我們呢？ 然而，我們並沒有用過這權利，倒是凡事忍受，免得基督的福音受到阻礙。
1COR|9|13|你們豈不知在聖殿供職的人吃聖殿中的食物嗎？在祭壇伺候的人分享壇上的供物嗎？
1COR|9|14|主也是這樣命令，要傳福音的人靠著福音養生。
1COR|9|15|但這權利我全然沒有用過。我寫這些話，並非要你們這樣待我，因為我寧可死也不讓人使我所誇的落了空。
1COR|9|16|我傳福音原沒有可誇耀的，因為我是不得已的，若不傳福音，我就有禍了。
1COR|9|17|我若甘心做這事，就有賞賜；若不甘心，責任卻已經託付給我了。
1COR|9|18|這樣，我的賞賜是甚麼呢？就是我傳福音的時候，使人不花錢得福音，免得我用盡了傳福音的權利。
1COR|9|19|我雖然是自由的，不受人管轄，但我甘心作了眾人的僕人，為贏得更多的人。
1COR|9|20|對 猶太 人，我就作 猶太 人，為要贏得 猶太 人；對律法以下的人，我雖不在律法以下，還是作律法以下的人，為要贏得律法以下的人。
1COR|9|21|對沒有律法的人，我就作沒有律法的人，為要贏得沒有律法的人；其實我在上帝面前，不是沒有律法，而是在基督的律法之下。
1COR|9|22|對軟弱的人，我就作軟弱的人，為要贏得軟弱的人。對甚麼樣的人，我就作甚麼樣的人。無論如何我總要救一些人。
1COR|9|23|凡我所做的，都是為福音的緣故，為要與人共享這福音的好處。
1COR|9|24|你們不知道在運動場上賽跑的，大家都跑，但得獎賞的只有一人？你們也要這樣跑，好使你們得著獎賞。
1COR|9|25|凡參加競賽的，在各方面都要有節制，他們不過是要得會朽壞的冠冕；我們卻是要得不會朽壞的冠冕。
1COR|9|26|所以，我奔跑，不像無目標的；我鬥拳，不像打空氣的。
1COR|9|27|我克制己身，使它完全順服，免得我傳福音給別人，自己反而被淘汰了。
1COR|10|1|弟兄們，我不願意你們不知道，我們的祖宗從前都在雲下，都從海中經過，
1COR|10|2|都在雲裏、海裏受洗 歸了 摩西 ，
1COR|10|3|並且都吃了一樣的靈糧，
1COR|10|4|也都喝了一樣的靈水，所喝的是出於跟隨著他們的靈磐石；那磐石就是基督。
1COR|10|5|但他們中間多半是上帝不喜歡的人，所以倒斃在曠野裏了。
1COR|10|6|這些事都是我們的鑒戒，使我們不要貪戀惡事，像他們貪戀過的一樣。
1COR|10|7|也不要拜偶像，像他們中有些人曾經拜過。如經上所記：「百姓坐下吃喝，起來玩樂。」
1COR|10|8|我們也不可犯姦淫，像他們中有些人曾經犯過，一天就倒斃了二萬三千人。
1COR|10|9|也不可試探主 ，像他們中有些人曾試探主就被蛇咬死。
1COR|10|10|你們也不可發怨言，像他們中有些人曾經發過，就被毀滅者所滅。
1COR|10|11|這些事發生在他們身上，要作為鑒戒，而且寫下來正是要警戒我們這末世的人。
1COR|10|12|所以，自以為站得穩的人必須謹慎，免得跌倒。
1COR|10|13|你們所受的考驗無非是人所承受得了的。上帝是信實的，他不會讓你們遭受無法承受的考驗，在受考驗的時候，總會給你們開一條出路，讓你們能忍受得了。
1COR|10|14|所以，我親愛的，你們要遠避拜偶像的事。
1COR|10|15|我好像對精明人說的；你們要辨別我的話。
1COR|10|16|我們所祝謝的杯，豈不是同領基督的血嗎？我們所擘開的餅，豈不是同領基督的身體嗎？
1COR|10|17|因為餅只是一個，我們雖然人多，仍是一體，我們同享一個餅。
1COR|10|18|你們看那按肉體是 以色列 人的，那些吃祭物的人豈不是與祭壇有份嗎？
1COR|10|19|那麼，我怎麼說呢？是說祭偶像之物算得了甚麼嗎？或說偶像算得了甚麼嗎？
1COR|10|20|不，我是說，他們 所獻的祭是祭鬼，不是祭上帝；我不願意你們與鬼來往。
1COR|10|21|你們不能喝主的杯，又喝鬼的杯；不能吃主的筵席，又吃鬼的筵席。
1COR|10|22|我們要惹主的嫉恨嗎？我們比他更強嗎？
1COR|10|23|「凡事都可行」，但不都有益處。「凡事都可行」，但不都造就人。
1COR|10|24|無論甚麼人，不要求自己的益處，而要求別人的益處。
1COR|10|25|凡市場上所賣的，你們只管吃，不要為良心的緣故問甚麼，
1COR|10|26|「因為地和其中所充滿的都屬於主」。
1COR|10|27|倘若有一個不信的人請你們吃飯，而你們也願意去，凡擺在你們面前的，只管吃，不要為良心的緣故問甚麼。
1COR|10|28|若有人對你們說：「這是獻過祭的物」，那麼為了那告訴你們的人，並為了良心的緣故就不吃。
1COR|10|29|我說的良心不是你自己的，而是他的。我的自由為甚麼被別人的良心評斷呢？
1COR|10|30|我若謝恩而吃，為甚麼因我謝恩的物被人毀謗呢？
1COR|10|31|所以，你們或吃或喝，無論做甚麼，都要為榮耀上帝而做。
1COR|10|32|你們不要使 猶太 人、 希臘 人，或上帝教會中的人跌倒；
1COR|10|33|但要像我一樣，凡事都使眾人喜歡，不求自己的益處，只求眾人的益處，使他們得救。
1COR|11|1|你們該效法我，像我效法基督一樣。
1COR|11|2|我稱讚你們，因為你們凡事記得我，又堅守我所傳授給你們的。
1COR|11|3|但是我要你們知道：基督是男人的頭；男人是女人的頭 ；上帝是基督的頭。
1COR|11|4|凡男人禱告或講道 ，若蒙著頭，就是羞辱自己的頭。
1COR|11|5|凡女人禱告或講道，若不蒙著頭，就是羞辱自己的頭，因為這就如同剃了頭髮一樣。
1COR|11|6|女人若不蒙著頭，就該剪了頭髮；女人若以剪髮剃髮為羞愧，就該蒙著頭。
1COR|11|7|男人本不該蒙著頭，因為他是上帝的形像和榮耀；但女人是男人的榮耀。
1COR|11|8|起初，男人不是由女人而出，女人卻是由男人而出。
1COR|11|9|而且男人不是為女人造的，女人卻是為男人造的。
1COR|11|10|因此，女人為天使的緣故應當在頭上有服權柄的記號。
1COR|11|11|然而，照主的安排，女人不可沒有男人，男人也不可沒有女人。
1COR|11|12|因為女人原是由男人而出，男人是藉著女人而生；但萬有都是出於上帝。
1COR|11|13|你們自己要判斷，女人禱告上帝，不蒙著頭合宜嗎？
1COR|11|14|你們的本性不也教導你們，男人若留長頭髮是他的羞辱嗎？
1COR|11|15|但女人留長頭髮是她的榮耀，因為這頭髮是給她蓋頭的 。
1COR|11|16|若有人想要辯駁，我們卻沒有這樣的規矩，上帝的眾教會也沒有。
1COR|11|17|我現在吩咐你們這話不是在稱讚你們，因為你們聚會是有損無益的。
1COR|11|18|首先，我聽說你們教會聚會的時候有分裂的事，我也有些相信這話。
1COR|11|19|在你們中間必然有分門結黨的事，好使那些經得起考驗的人顯明出來。
1COR|11|20|你們聚會的時候，不是在吃主的晚餐，
1COR|11|21|因為吃的時候，各人先吃自己的飯，甚至有人飢餓，有人酒醉。
1COR|11|22|難道你們沒有家可以吃喝嗎？還是你們藐視上帝的教會，使那沒有的羞愧呢？我該對你們說甚麼呢？我要稱讚你們嗎？在這事上我絕不稱讚你們！
1COR|11|23|我當日傳給你們的是從主所領受的。主耶穌被出賣的那一夜，拿起餅來，
1COR|11|24|祝謝了，就擘開，說：「這是我的身體，為你們捨 的；你們要如此行，為的是記念我。」
1COR|11|25|飯後，他也照樣拿起杯來，說：「這杯是用我的血所立的新約；你們每逢喝的時候，要如此行，來記念我。」
1COR|11|26|你們每逢吃這餅，喝這杯，是宣告主的死，直到他來。
1COR|11|27|所以，任何不按規矩吃了主的餅，喝了主的杯，就是干犯主的身體和主的血了。
1COR|11|28|人應該省察自己，然後吃這餅，喝這杯。
1COR|11|29|因為人吃喝，若不分辨是主的身體，他的吃喝就是定自己的罪了。
1COR|11|30|因此，在你們中間有好些軟弱的與患病的，長眠了的也不少。
1COR|11|31|我們若是先省察自己，就不至於受審判。
1COR|11|32|我們受審判的時候，就是被主管教，這樣就免得和世人一同被定罪。
1COR|11|33|所以，我的弟兄們，你們聚會吃晚餐的時候，要彼此等待。
1COR|11|34|若有人餓了，要在家裏先吃，免得你們聚會，反被定罪。其餘的事等我來的時候再安排。
1COR|12|1|弟兄們，關於屬靈的恩賜 ，我不願意你們不明白。
1COR|12|2|你們知道，你們作外邦人的時候，隨事被引誘，受了迷惑去拜不會出聲的偶像。
1COR|12|3|所以，我要你們知道，被上帝的靈感動的，沒有人會說「耶穌該受詛咒」；若不是被聖靈感動的，也沒有人能說「耶穌是主」。
1COR|12|4|恩賜有許多種，卻是同一位聖靈所賜。
1COR|12|5|事奉有許多種，卻是事奉同一位主。
1COR|12|6|工作有許多種，卻是同一位上帝在萬人中運行萬事。
1COR|12|7|聖靈彰顯在各人身上，是要使人得益處。
1COR|12|8|有人藉著聖靈領受智慧的言語；有人也靠著同一位聖靈領受知識的言語；
1COR|12|9|又有人由同一位聖靈領受信心；還有人由同一位聖靈領受醫病的恩賜；
1COR|12|10|又有人能行異能，又有人能作先知，又有人能辨別諸靈，又有人能說方言 ，又有人能翻方言。
1COR|12|11|這一切都是由惟一的、同一位聖靈所運行，隨著自己的旨意分給各人的。
1COR|12|12|就如身體是一個，卻有許多肢體，身體的肢體雖多，仍是一個身體；基督也是這樣。
1COR|12|13|我們無論是 猶太 人是 希臘 人，是為奴的是自主的，都從一位聖靈受洗成了一個身體，並且共享這位聖靈。
1COR|12|14|身體原不只是一個肢體，而是許多肢體。
1COR|12|15|假如腳說：「我不是手，所以不屬於身體」，它不能因此就不屬於身體。
1COR|12|16|假如耳朵說：「我不是眼睛，所以不屬於身體」，它也不能因此就不屬於身體。
1COR|12|17|假如全身是眼睛，聽覺在哪裏呢？假如全身是耳朵，嗅覺在哪裏呢？
1COR|12|18|但現在上帝隨自己的意思把肢體一一安置在身體上了。
1COR|12|19|假如全都是一個肢體，身體在哪裏呢？
1COR|12|20|但現在肢體雖多，身體還是一個。
1COR|12|21|眼睛不能對手說：「我用不著你。」頭也不能對腳說：「我用不著你。」
1COR|12|22|不但如此，身上的肢體，人以為軟弱的，更是不可缺少的；
1COR|12|23|身上的肢體，我們認為不體面的，越發給它加上體面；我們不雅觀的，越發裝飾得雅觀。
1COR|12|24|我們雅觀的肢體自然用不著裝飾；但上帝配搭這身子，把加倍的體面給那有缺欠的肢體，
1COR|12|25|免得身體不協調，總要肢體彼此照顧。
1COR|12|26|假如一個肢體受苦，所有的肢體就一同受苦；假如一個肢體得光榮，所有的肢體就一同快樂。
1COR|12|27|你們是基督的身體，並且各自都是肢體。
1COR|12|28|上帝在教會所設立的：第一是使徒；第二是先知；第三是教師；其次是行異能的；再次是醫病的恩賜，幫助人的，治理事的，說方言的。
1COR|12|29|難道個個都是使徒嗎？難道個個都是先知嗎？難道個個都是教師嗎？難道個個都是行異能的嗎？
1COR|12|30|難道個個都是有醫病的恩賜嗎？難道個個都是說方言的嗎？難道個個都是翻方言的嗎？
1COR|12|31|你們要追求那更大的恩賜。 我現今把最妙的道指示你們。
1COR|13|1|我若能說人間的方言，甚至天使的語言，卻沒有愛，我就成為鳴的鑼、響的鈸一般。
1COR|13|2|我若有先知講道的能力，也明白各樣的奧祕，各樣的知識，而且有齊備的信心，使我能夠移山，卻沒有愛，我就算不了甚麼。
1COR|13|3|我若將所有的財產救濟窮人，又犧牲自己的身體讓人誇讚 ，卻沒有愛，仍然對我無益。
1COR|13|4|愛是恆久忍耐；又有恩慈；愛是不嫉妒；愛是不自誇，不張狂，
1COR|13|5|不做害羞的事，不求自己的益處，不輕易發怒，不計算人的惡，
1COR|13|6|不喜歡不義，只喜歡真理；
1COR|13|7|凡事包容，凡事相信，凡事盼望，凡事忍耐。
1COR|13|8|愛是永不止息。先知講道之能終必歸於無有；說方言 之能終必停止；知識也終必歸於無有。
1COR|13|9|我們現在所知道的有限，先知所講的也有限，
1COR|13|10|等那完全的來到，這有限的必消逝。
1COR|13|11|我作孩子的時候，說話像孩子，心思像孩子，意念像孩子；既長大成人，就把孩子的事丟棄了。
1COR|13|12|我們現在是對著鏡子觀看，模糊不清 ；到那時，就要面對面了。我如今所認識的有限，到那時就全認識，如同主認識我一樣。
1COR|13|13|如今常存的有信，有望，有愛這三樣，其中最大的是愛。
1COR|14|1|你們要追求愛，也要切慕屬靈的恩賜，尤其是作先知講道 。
1COR|14|2|那說方言 的，不是對人說，而是對上帝說，因為沒有人聽得懂；他是藉著聖靈說各樣的奧祕。
1COR|14|3|但作先知講道的，是對人說，要造就、安慰、勸勉人。
1COR|14|4|說方言的，是造就自己；作先知講道的，是造就教會。
1COR|14|5|我希望你們都說方言，更希望你們作先知講道；因為說方言的，若不解釋出來，使教會得造就，那作先知講道的就比他強了。
1COR|14|6|弟兄們，我到你們那裏去，若只說方言，不用啟示，或知識，或預言，或教導，給你們講解，我對你們有甚麼益處呢？
1COR|14|7|就連那有聲而沒有生命的東西，如簫，如琴，發出來的音若沒有分別，怎能知道所吹所彈的是甚麼呢？
1COR|14|8|號角吹出來的音若不清楚，誰會預備打仗呢？
1COR|14|9|你們也是如此；若用舌頭說聽不懂的信息，怎能知道所說的是甚麼呢？你們就是向空氣說話了。
1COR|14|10|世上有許多種語言，卻沒有一樣是無意思的。
1COR|14|11|我若不明白那語言的意思，說話的人必以我為未開化的人，我也以他為未開化的人。
1COR|14|12|你們也是如此，既然你們切慕屬靈的恩賜，就當追求多得造就教會的恩賜。
1COR|14|13|所以，那說方言的，就當祈求有翻方言的恩賜。
1COR|14|14|我若用方言禱告，是我的靈在禱告；但我的理智沒有效果。
1COR|14|15|我應該怎麼做呢？我要用靈禱告，也要用理智禱告；我要用靈歌唱，也要用理智歌唱。
1COR|14|16|不然，你用靈祝謝，那在座不通方言的人，既然不明白你的話，怎能在你感謝的時候說「阿們」呢？
1COR|14|17|你的感謝固然是好，不過不能造就別人。
1COR|14|18|我感謝上帝，我說方言比你們眾人還多；
1COR|14|19|但在教會中，我寧可用理智說五句教導人的話，強過說萬句方言。
1COR|14|20|弟兄們，在心志上不要作小孩子。但是，在惡事上要作嬰孩，而在心志上總要作大人。
1COR|14|21|律法上記著：「主說： 我要用外邦人的舌頭 和外邦人的嘴唇 向這百姓說話； 雖然如此，他們還是不聽從我。」
1COR|14|22|這樣看來，說方言不是為信的人作標記，而是為不信的人；作先知講道不是為不信的人作標記，而是為信的人。
1COR|14|23|所以，全教會聚在一處的時候，若都說方言，偶然有不通方言的或是不信的人進來，豈不會說你們瘋了嗎？
1COR|14|24|若個個都作先知講道，偶然有不信的或是不懂方言的人進來，就被眾人勸戒，被眾人審問，
1COR|14|25|他心裏的隱情被顯露出來，就必將臉伏地，敬拜上帝，宣告說：「上帝真的是在你們中間了。」
1COR|14|26|弟兄們，那麼，你們該怎麼做呢？你們聚會的時候，各人或有詩歌，或有教導，或有啟示，或有方言，或有翻出來，凡事都應當造就人。
1COR|14|27|若有說方言的，只可有兩個人，至多三個人，且要輪流著說，也要有一個人翻出來。
1COR|14|28|若沒有人翻，就當在會中閉口，只對自己和上帝說就是了。
1COR|14|29|至於作先知講道的，只可有兩個人或是三個人，其餘的人當慎思明辨。
1COR|14|30|假如旁邊坐著的得了啟示，那先說話的就當閉口不言。
1COR|14|31|因為你們都可以一個一個地作先知講道，使眾人都可以學習，使眾人都得勸勉。
1COR|14|32|先知的靈是順服先知的，
1COR|14|33|因為上帝不是叫人混亂，而是叫人和諧的上帝。 在聖徒的眾教會中，
1COR|14|34|婦女應該閉口不言；因為，不准她們說話，總要順服，正如律法所說的。
1COR|14|35|她們若要學甚麼，應該在家裏問自己的丈夫，因為婦女在會中說話是可恥的。
1COR|14|36|難道上帝的話是從你們出來的嗎？難道是單臨到你們的嗎？
1COR|14|37|若有人自以為是先知，或是屬靈的，就應該知道，我所寫給你們的是主的命令。
1COR|14|38|若有不理會的，你們也不必理會他。
1COR|14|39|所以，我的弟兄們，你們要切慕作先知講道的恩賜，不要禁止說方言。
1COR|14|40|凡事都要規規矩矩地按著次序行。
1COR|15|1|弟兄們，我要你們認清我先前傳給你們的福音；這福音你們領受了，又靠著它站立得住，
1COR|15|2|你們若能夠持守我傳給你們的信息，就必因這福音得救，否則你們是徒然相信。
1COR|15|3|我當日所領受又傳給你們的，最重要的就是：照聖經所說，基督為我們的罪死了，
1COR|15|4|而且埋葬了；又照聖經所說，第三天復活了，
1COR|15|5|還顯給 磯法 看，又顯給十二使徒看，
1COR|15|6|後來一次顯給五百多弟兄看，其中一大半到現在還在，卻也有已經睡了的。
1COR|15|7|以後他顯給 雅各 看，再顯給眾使徒看，
1COR|15|8|最後也顯給我看；我如同未到產期而生的人一般。
1COR|15|9|我原是使徒中最小的，不配稱為使徒，因為我曾迫害過上帝的教會。
1COR|15|10|然而，由於上帝的恩典，我才成了今日的我，並且他所賜給我的恩典不是徒然的。我比眾使徒格外勞苦；其實不是我，而是上帝的恩典與我同在。
1COR|15|11|無論是我或是其他使徒，我們都如此傳，你們也都如此信了。
1COR|15|12|既然我們傳基督是從死人中復活了，怎麼在你們中間有人說沒有死人復活的事呢？
1COR|15|13|若沒有死人復活的事，基督就沒有復活了。
1COR|15|14|基督若沒有復活，我們所傳的就是枉然，你們所信的也是枉然。
1COR|15|15|這樣，我們甚至被當作是為上帝妄作見證的，因為我們見證上帝是使基督復活了。如果死人真的沒有復活，上帝就沒有使基督復活了。
1COR|15|16|因為死人若不復活，基督也就沒有復活了。
1COR|15|17|基督若沒有復活，你們的信就是徒然，你們仍活在罪裏。
1COR|15|18|就是在基督裏睡了的人也滅亡了。
1COR|15|19|我們若靠基督只在今生有指望，就比所有的人更可憐了。
1COR|15|20|其實，基督已經從死人中復活，成為睡了之人初熟的果子。
1COR|15|21|既然死是因一人而來，死人復活也因一人而來。
1COR|15|22|在 亞當 裏眾人都死了；同樣，在基督裏眾人也都要復活。
1COR|15|23|但各人是按著自己的次序復活：初熟的果子是基督；然後在他來的時候，是那些屬於基督的。
1COR|15|24|再後，終結到了，那時基督既將一切執政的、掌權的、有權能的都毀滅了，就把國交給父上帝。
1COR|15|25|因為基督必須掌權，等上帝把一切仇敵都放在他的腳下。
1COR|15|26|他要毀滅的最後仇敵就是死亡。
1COR|15|27|因為經上說：「上帝使萬物都服在他的腳下。」既然說萬物都服了他，那使萬物屈服的，很明顯地是不在其內了。
1COR|15|28|既然萬物服了他，那時，子也要自己順服那叫萬物服他的，好使上帝在萬物之中，在萬物之上。
1COR|15|29|不然，那些為死人受洗的，能做甚麼呢？如果死人不會復活，為甚麼替他們受洗呢？
1COR|15|30|我們為甚麼要時刻冒險呢？
1COR|15|31|弟兄們 ，我在我們的主基督耶穌裏，指著你們—我所誇的極力地說，我天天冒死。
1COR|15|32|從人的觀點看來，我當日在 以弗所 同野獸搏鬥，對我有甚麼益處呢？如果死人沒有復活， 「讓我們吃吃喝喝吧！ 因為明天要死了。」
1COR|15|33|不要被欺騙了； 「濫交朋友敗壞品德。」
1COR|15|34|你們要醒悟為善，不再犯罪；因為有人不認識上帝。我說這話是要使你們羞愧。
1COR|15|35|但是有人會問：「死人怎樣復活呢？他們帶著甚麼身體來呢？」
1COR|15|36|無知的人哪，你所種的若不死就不能生。
1COR|15|37|並且你所種的不是那將來要有的形體，無論是麥子或別樣穀物，都不過是子粒。
1COR|15|38|但上帝隨自己的意思給它一個形體，並叫各樣子粒各有自己的形體。
1COR|15|39|不是所有的肉體都是同樣的：人是一個樣子，獸又是一個樣子，鳥又是一個樣子，魚又是一個樣子。
1COR|15|40|有天上的形體，也有地上的形體；但天上形體的榮光是一個樣子，地上形體的榮光又是一個樣子。
1COR|15|41|日有日的光輝，月有月的光輝，星有星的光輝；這星和那星的光輝也有區別。
1COR|15|42|死人復活也是這樣。所種的是會朽壞的，復活的是不朽壞的；
1COR|15|43|所種的是羞辱的，復活的是榮耀的；所種的是軟弱的，復活的是強壯的；
1COR|15|44|所種的是血肉的身體，復活的是靈性的身體。既有血肉的身體，也就有靈性的身體。
1COR|15|45|經上也是這樣記著說：「首先的人 亞當 成了有生命的人」；末後的 亞當 成了賜生命的靈。
1COR|15|46|但是，不是屬靈的在先，而是屬血肉的在先，然後才是屬靈的。
1COR|15|47|第一個人是出於地，是屬於塵土；第二個人是出於天。
1COR|15|48|那屬塵土的怎樣，凡屬塵土的也都怎樣；屬天的怎樣，凡屬天的也都怎樣。
1COR|15|49|就如我們既有屬塵土的形像，將來也必有屬天的形像。
1COR|15|50|弟兄們，我要告訴你們的是：血肉之軀不能承受上帝的國，必朽壞的也不能承受不朽壞的。
1COR|15|51|我如今把一件奧祕的事告訴你們：我們不是都要睡覺，而是都要改變，
1COR|15|52|就在一剎那，眨眼之間，號筒末次吹響的時候。因號筒要吹響，死人要復活成為不朽壞的，我們也要改變。
1COR|15|53|這會朽壞的必須變成 不朽壞的；這會死的總要變成不會死的。
1COR|15|54|當這會朽壞的變成不朽壞的，這會死的變成不會死的，那時經上所記「死亡已被勝利吞滅了」的話就應驗了。
1COR|15|55|「死亡啊！你得勝的權勢在哪裏？ 死亡啊！你的毒刺在哪裏？」
1COR|15|56|死亡的毒刺就是罪，罪的權勢就是律法。
1COR|15|57|感謝上帝，他使我們藉著我們的主耶穌基督得勝。
1COR|15|58|所以，我親愛的弟兄們，你們務要堅固，不可動搖，常常竭力多做主工，因為你們知道，你們在主裏的勞苦不是徒然的。
1COR|16|1|關於為聖徒捐款的事，我從前怎樣吩咐 加拉太 的眾教會，你們也該怎樣做。
1COR|16|2|每逢七日的第一日，每人要照自己的收入抽出若干，保留起來，免得我來的時候現湊。
1COR|16|3|等到我來了，你們寫信舉薦誰，我就差遣他們，把你們的款項送到 耶路撒冷 去。
1COR|16|4|如果我也該去，他們可以和我同去。
1COR|16|5|我想穿越 馬其頓 ；我經過了 馬其頓 後，就到你們那裏去，
1COR|16|6|可能會和你們同住一些時候，甚至和你們一起過冬。這樣無論我往哪裏去，你們可以給我送行。
1COR|16|7|我現在不願意在路過的時候見你們；主若允許，我就指望和你們同住一些時候。
1COR|16|8|不過我要仍舊住在 以弗所 ，直到五旬節，
1COR|16|9|因為有又寬大又有效的門為我開了，雖然反對的人也多。
1COR|16|10|若是 提摩太 來到，你們要留心照顧他，使他在你們那裏無所懼怕，因為他做主的工作像我一樣。
1COR|16|11|所以，無論誰都不可藐視他。只要送他平安前行，讓他到我這裏來，因為我等著他和弟兄們同來。
1COR|16|12|至於 亞波羅 弟兄，我再三勸他同弟兄們到你們那裏去；但現在他絕不願意去，等有機會他就會去。
1COR|16|13|你們要警醒，在信仰上要站穩，要勇敢，要剛強。
1COR|16|14|你們所做的一切都要憑愛心而做。
1COR|16|15|弟兄們，你們知道 司提法那 一家，是 亞該亞 初結的果子；他們專以服事聖徒為念。
1COR|16|16|我勸你們順服這樣的人，和一切與他同工同勞的人。
1COR|16|17|司提法那 、 福徒拿都 和 亞該古 到這裏來，我很高興，因為他們補上了你們不在我身邊的遺憾。
1COR|16|18|他們使我和你們心裏都快慰；這樣的人，你們務要敬重。
1COR|16|19|亞細亞 的眾教會向你們問安。 亞居拉 、 百基拉 ，和在他們家裏的教會，在主裏熱切地向你們問安。
1COR|16|20|眾弟兄都向你們問安。要用聖潔的吻彼此問安。
1COR|16|21|我— 保羅 親筆問安。
1COR|16|22|若有人不愛主，這人該受詛咒。主啊，願你來！
1COR|16|23|願主耶穌基督的恩常與你們眾人同在。
1COR|16|24|我在基督耶穌裏的愛與你們同在！
2COR|1|1|奉上帝旨意作基督耶穌使徒的 保羅 和弟兄 提摩太 ，寫信給在 哥林多 上帝的教會和全 亞該亞 的眾聖徒。
2COR|1|2|願恩惠、平安 從我們的父上帝和主耶穌基督歸給你們！
2COR|1|3|願頌讚歸於上帝—我們主耶穌基督的父；他是發慈悲的父，賜各樣安慰的上帝。
2COR|1|4|我們在一切患難中，他安慰我們，使我們能用上帝所賜的安慰去安慰那些遭各樣患難的人。
2COR|1|5|正如我們跟基督同受許多苦楚，我們也靠基督得許多安慰。
2COR|1|6|如果我們受患難，那是為使你們得安慰，得拯救；如果我們得安慰，那也是為使你們得安慰，這安慰能使你們忍受我們所受同樣的苦楚。
2COR|1|7|我們為你們所存的盼望是確定的，因為知道你們分擔了我們的痛苦，也要分享我們的安慰。
2COR|1|8|弟兄們，我們不要你們不知道，我們從前在 亞細亞 遭遇苦難，因受到無法忍受的壓力，甚至連活命的指望都沒有了。
2COR|1|9|自己心裏也斷定是必死無疑，這是要使我們不依靠自己，只依靠使死人復活的上帝。
2COR|1|10|他曾救我們脫離那極大的死亡，他要繼續救我們，而且我們指望他將來還要救我們。
2COR|1|11|你們也要一同用祈禱來幫助我們，好使許多人為我們感恩，因著他們許多的禱告，我們獲得了恩賜。
2COR|1|12|我們所誇的是：我們在世為人，特別是跟你們的關係，是憑著上帝所賜的坦率和真誠，不是靠人的聰明，而是靠上帝的恩惠；這是我們的良心可以作證的。
2COR|1|13|我們現在寫給你們的話，無非是你們所能誦讀、所能明白的，我也盼望你們真能徹底明白。
2COR|1|14|你們已經有幾分認識我們，在我們主耶穌 的日子，你們會以我們為榮，正像我們也以你們為榮。
2COR|1|15|既然我這樣深信，早就有意先到你們那裏去，讓你們得加倍的益處。
2COR|1|16|我要路過你們那裏往 馬其頓 去，再從 馬其頓 回到你們那裏，讓你們給我送行往 猶太 去。
2COR|1|17|我有此意，難道是反覆不定嗎？難道我的意願是從私慾起的，以致我忽是忽非嗎？
2COR|1|18|我指著信實的上帝說，我們向你們所傳的道並非又是又非的。
2COR|1|19|因為，我、 西拉 和 提摩太 在你們中間傳上帝的兒子耶穌基督，從沒有「又是又非」的；在他只有一個「是」。
2COR|1|20|上帝的應許，不論有多少，在基督都是「是」的。所以，我們藉著他說「阿們」，使上帝因我們得榮耀。
2COR|1|21|那在基督裏堅固我們和你們，並且膏抹我們的，就是上帝。
2COR|1|22|他在我們身上蓋了印，並賜聖靈在我們心裏作憑據。
2COR|1|23|我指著我的性命求告上帝作證，我沒有再往 哥林多 去是為了要寬容你們。
2COR|1|24|我們並不是要控制你們的信心，而是要作你們的同工，讓你們得快樂，因為你們在信仰上已經站得穩了。
2COR|2|1|我自己定了主意，下次不再帶著悲傷到你們那裏去。
2COR|2|2|我若使你們悲傷，除了因我而使他悲傷的那人以外，誰能使我喜樂呢？
2COR|2|3|我曾把這事寫給你們，免得我到的時候，那該令我喜樂的人反倒令我悲傷。我也深信，你們眾人都以我的喜樂為自己的喜樂。
2COR|2|4|我先前憂心忡忡、眼淚汪汪地給你們寫了信，並非要使你們悲傷，而是要你們知道我格外疼愛你們。
2COR|2|5|如果有人使人悲傷，他不但使我悲傷，也是使你們眾人有些悲傷。我說有些，恐怕說得太重了。
2COR|2|6|這樣的人受了大多數人的責備也就夠了，
2COR|2|7|倒不如赦免他，安慰他，免得他過分悲傷，甚至受不了啦！
2COR|2|8|所以，我勸你們，要向他肯定你們的愛心。
2COR|2|9|為此，我先前也寫信給你們，正是要考驗你們，看你們是否在一切事上都順從我。
2COR|2|10|你們赦免誰，我也赦免誰。我若有所赦免，是在基督面前為你們的緣故赦免的，
2COR|2|11|免得撒但趁著機會勝過我們，因我們並非不知道他的詭計。
2COR|2|12|我從前為基督的福音到了 特羅亞 ，主給我開了門。
2COR|2|13|那時，因為沒有遇見我的弟兄 提多 ，我心裏不安，就辭別那裏的人，往 馬其頓 去了。
2COR|2|14|感謝上帝！他常率領我們在基督裏得勝，並藉著我們在各處顯揚那因認識基督而有的香氣。
2COR|2|15|因為無論在得救的人或在滅亡的人當中，我們都是基督馨香之氣，是獻給上帝的。
2COR|2|16|對滅亡的人，這是死而又死的氣味；對得救的人，這是生而又生的氣味。這些事誰能當得起呢？
2COR|2|17|我們不像許多人，把上帝的道當商品販賣，而是由於真誠，而是受命於上帝，在上帝面前憑著基督講道。
2COR|3|1|難道我們又開始推薦自己嗎？難道我們像某些人那樣要用人的推薦信介紹給你們，或用你們的推薦信給人嗎？
2COR|3|2|你們就是我們的推薦信，寫在我們心裏，被眾人所知道、所誦讀的，
2COR|3|3|而你們顯明自己是基督的書信，藉著我們寫成的。不是用墨寫的，而是用永生上帝的靈寫的；不是寫在石版上，而是寫在心版上的。
2COR|3|4|我們藉著基督才對上帝有這樣的信心。
2COR|3|5|並不是我們憑自己配做甚麼事，我們之所以配做是出於上帝；
2COR|3|6|他使我們能配作新約的執事，不是文字上的約，而是聖靈的約；因為文字使人死，聖靈能使人活。
2COR|3|7|那用字刻在石頭上屬死的事奉尚且有榮光，以致 以色列 人因 摩西 臉上那逐漸褪色的榮光不能定睛看他的臉，
2COR|3|8|那屬聖靈的事奉不是更有榮光嗎？
2COR|3|9|若是那使人定罪的事奉有榮光，那使人稱義的事奉的榮光就越發大了。
2COR|3|10|那從前有榮光的，因這更大的榮光，就算不得有榮光了；
2COR|3|11|若是那逐漸褪色的有榮光，這長存的就更有榮光了。
2COR|3|12|既然我們有這樣的盼望，就大有膽量，
2COR|3|13|不像 摩西 將面紗蒙在臉上，使 以色列 人不能定睛看到那逐漸褪色的榮光的結局。
2COR|3|14|但他們的心地剛硬，直到今日誦讀舊約的時候，這同樣的面紗還沒有揭去；因為這面紗在基督裏才被廢去。
2COR|3|15|然而直到今日，每逢誦讀 摩西 書的時候，面紗還在他們心上。
2COR|3|16|但他們的心何時歸向主，面紗就何時除去。
2COR|3|17|主就是那靈；主的靈在哪裏，哪裏就有自由。
2COR|3|18|既然我們眾人以揭去面紗的臉得以看見 主的榮光，好像從鏡子裏返照，就變成了與主有同樣的形像，榮上加榮，如同從主的靈 變成的。
2COR|4|1|所以，既然我們蒙憐憫受了這事奉的責任，就不喪膽，
2COR|4|2|反而把那些暗昧可恥的事棄絕了，不行詭詐，不曲解上帝的道，只將真理顯揚出來，好在上帝面前把自己推薦給各人的良心。
2COR|4|3|即使我們的福音被遮蔽，那只是對滅亡的人遮蔽。
2COR|4|4|這些不信的人被這世界的神明弄瞎了心眼，使他們看不見基督榮耀的福音。基督本是上帝的像。
2COR|4|5|我們不是傳自己，而是傳耶穌基督為主，並且自己因耶穌作你們的僕人。
2COR|4|6|那吩咐光從黑暗裏照出來的上帝已經照在我們心裏，使我們知道上帝榮耀的光顯在耶穌基督的臉上。
2COR|4|7|我們有這寶貝放在瓦器裏，為要顯明這莫大的能力是出於上帝，不是出於我們。
2COR|4|8|我們處處受困，卻不被捆住；內心困擾，卻沒有絕望；
2COR|4|9|遭受迫害，卻不被撇棄；擊倒在地，卻不致滅亡。
2COR|4|10|我們身上常帶著耶穌的死，使耶穌的生也在我們身上顯明。
2COR|4|11|因為我們這活著的人常為耶穌被置於死地，使耶穌的生命在我們這必死的人身上顯明出來。
2COR|4|12|這樣看來，死是在我們身上運作，生卻在你們身上運作。
2COR|4|13|但我們既然有從同一位靈而來的信心，正如經上記著：「我信，故我說話」，我們也信，所以也說話；
2COR|4|14|因為知道，那使主耶穌復活的也必使我們與耶穌一同復活，並且使我們與你們一起站在他面前。
2COR|4|15|凡事都是為了你們，好使恩惠既藉著更多的人而加增，感恩也格外顯多，好歸榮耀給上帝。
2COR|4|16|所以，我們不喪膽。雖然我們外在的人日漸朽壞，內在的人卻日日更新。
2COR|4|17|我們這短暫而輕微的苦楚要為我們成就極重、無比、永遠的榮耀。
2COR|4|18|因為我們不是顧念看得見的，而是顧念看不見的；原來看得見的是暫時的，看不見的才是永遠的。
2COR|5|1|因為我們知道，我們這地上的帳篷若拆毀了，我們將有上帝所造的居所，不是人手所造的，而是在天上永存的。
2COR|5|2|我們在這帳篷裏嘆息，渴望得到那從天上來的居所，好像穿上衣服；
2COR|5|3|倘若脫下也 不至於赤身了。
2COR|5|4|其實，我們在這帳篷裏的人勞苦嘆息，並不是願意脫下地上的帳篷，而是願意穿上天上的居所，好使這必死的被生命吞滅了。
2COR|5|5|那為我們安排這事的是上帝，他賜給我們聖靈作憑據 。
2COR|5|6|所以，我們總是勇敢的，並且知道，只要我們住在這身體內就是離開了主。
2COR|5|7|因為我們行事為人是憑著信心，不是憑著眼見。
2COR|5|8|我們勇敢，更情願離開身體，與主同住。
2COR|5|9|所以，無論是住在身內或住在身外，我們都立了志向要得主的喜悅。
2COR|5|10|因為我們眾人必須站在基督審判臺前受審，為使各人按著本身所行的，或善或惡受報。
2COR|5|11|既然我們知道主是可畏的，就勸導人；但是上帝是認識我們的，我盼望你們的良心也認識我們。
2COR|5|12|我們不是向你們再推薦自己，而是要讓你們有誇耀我們的機會，使你們好面對那憑外貌、不憑內心誇耀的人。
2COR|5|13|如果我們癲狂，是為上帝；如果我們清醒，是為你們。
2COR|5|14|原來基督的愛激勵我們；因我們這樣斷定，一人既替眾人死了，眾人就都死了。
2COR|5|15|並且他替眾人死，是叫那些活著的人不再為自己活，乃為替他們死而復活的主活。
2COR|5|16|所以，從今以後，我們不再按照人的看法來認識人，縱使我們曾經按照人的看法認識基督，如今卻不再這樣認識他了。
2COR|5|17|所以，若有人在基督裏，他就是新造的人：舊事已過，都變成新的了。
2COR|5|18|一切都是出於上帝；他藉著基督使我們與他和好，又將勸人與他和好的使命賜給我們。
2COR|5|19|這就是：上帝在基督裏使世人與自己和好，不將他們的過犯歸到他們身上，並且將這和好的信息託付了我們。
2COR|5|20|所以，我們作基督的特使，就好像上帝藉我們勸你們一般。我們替基督求你們，與上帝和好吧！
2COR|5|21|上帝使那無罪 的，替我們成為罪，好使我們在他裏面成為上帝的義。
2COR|6|1|我們與上帝同工的也勸你們，不可白受他的恩典；
2COR|6|2|因為他說： 「在悅納的時候，我應允了你； 在拯救的日子，我幫助了你。」 看哪，現在正是悅納的時候！看哪，現在正是拯救的日子！
2COR|6|3|我們不在任何事上妨礙任何人，免得這使命被人毀謗；
2COR|6|4|反倒在各樣的事上表明自己是上帝的用人：就如在持久的忍耐、患難、困苦、災難、
2COR|6|5|鞭打、監禁、動亂、勞碌、失眠、飢餓、
2COR|6|6|廉潔、知識、堅忍、恩慈、聖靈的感化、無偽的愛心、
2COR|6|7|真實的言語、上帝的大能、藉著仁義的兵器在左在右、
2COR|6|8|榮譽或羞辱、惡名或美名。我們似乎是誘惑人的，卻是誠實的；
2COR|6|9|似乎不為人所知，卻是人所共知；似乎是死了，卻是活著；似乎受懲罰，卻沒有被處死；
2COR|6|10|似乎憂愁，卻常有喜樂；似乎貧窮，卻使許多人富足；似乎一無所有，卻樣樣都有。
2COR|6|11|哥林多 人哪，我們對你們，口是誠實的，心是寬宏的。
2COR|6|12|你們的狹窄不是由於我們，而是由於你們自己的心腸狹窄。
2COR|6|13|你們也要照樣用寬宏的心報答我；我這話正像對自己的孩子說的。
2COR|6|14|你們不要和不信的人同負一軛。義和不義有甚麼相關？光明和黑暗有甚麼相連？
2COR|6|15|基督和 彼列 有甚麼相和？信主的和不信主的有甚麼相干？
2COR|6|16|上帝的殿和偶像有甚麼相同？因為我們是永生上帝的殿，就如上帝曾說： 「我要在他們中間居住來往； 我要作他們的上帝， 他們要作我的子民。」
2COR|6|17|所以主說： 「你們務要從他們中間出來， 跟他們分別； 不要沾不潔淨的東西， 我就收納你們。
2COR|6|18|我要作你們的父， 你們要作我的兒女。 這是全能的主說的。」
2COR|7|1|所以，親愛的，既然我們有這樣的應許，就當潔淨自己，除去身體和靈魂一切的污穢，藉著敬畏上帝，得以成聖。
2COR|7|2|寬宏大量地接納我們吧！我們未曾虧負誰，未曾敗壞誰，未曾佔誰的便宜。
2COR|7|3|我說這話，不是要定你們的罪，我已經說過，你們常在我們心裏，我們情願與你們同生共死。
2COR|7|4|我對你們很是放心，多多誇耀你們；我滿有安慰，在我們一切患難中格外喜樂。
2COR|7|5|我們從前到了 馬其頓 的時候，身體沒有絲毫安寧，反而到處遭患難，外有紛爭，內有懼怕。
2COR|7|6|但那安慰灰心之人的上帝藉著 提多 來安慰了我們；
2COR|7|7|不但藉著他來，也藉著他從你們所得的安慰安慰了我們，因為他把你們的思念，你們的哀慟，你們對我的熱忱，都告訴了我，使我更加歡喜。
2COR|7|8|即使我先前那封信使你們憂愁，後來我曾懊悔，如今卻不懊悔；因為我知道，那封信使你們憂愁，不過是暫時的。
2COR|7|9|如今我歡喜，不是因你們曾憂愁，而是因憂愁導致你們的悔改。你們依著上帝的意思憂愁，凡事就不至於因我們受虧損了。
2COR|7|10|因為依著上帝的意思而憂愁，就生出沒有懊悔的悔改來，以致得救；但世俗的憂愁叫人死。
2COR|7|11|你看，你們依著上帝的意思而憂愁，這在你們當中產生了何等的殷勤、甚至辯白、甚至憤慨、甚至恐懼、甚至渴望、甚至熱忱、甚至責罰。在這一切事上，你們都表明自己是無可指責的。
2COR|7|12|所以，雖然我從前寫信給你們，卻不是為那虧負人的，也不是為那受人虧負的，而是要在上帝面前把你們顧念我們的熱忱表現出來。
2COR|7|13|因此，我們得了安慰。 在我們所得的安慰之外，又因你們眾人使 提多 心裏暢快喜樂，我們就更加歡喜了。
2COR|7|14|我若對 提多 誇獎過你們甚麼，也不覺得慚愧，因為我對 提多 誇獎你們的話是真的，正如我對你們所說的話也向來都是真的。
2COR|7|15|提多 一想起你們眾人的順服，怎樣恐懼戰兢地接待他，他愛你們的心就越發熱切了。
2COR|7|16|我如今歡喜，因為我在一切事上對你們有信心。
2COR|8|1|弟兄們，我們要把上帝賜給 馬其頓 眾教會的恩惠告訴你們：
2COR|8|2|他們在患難中受大考驗的時候，仍然滿有喜樂，在極度貧窮中還格外顯出他們樂捐的慷慨。
2COR|8|3|我可以證明，他們是按著能力，而且超過了能力來捐助，主動
2COR|8|4|再三懇求我們，准他們在這供給聖徒的善事上有份；
2COR|8|5|並且他們所做的，不但照我們所期望的，更照上帝的旨意先把自己獻給主，又給了我們。
2COR|8|6|因此，我們勸 提多 ，既然在你們中間開始這慈善的事，就當把它辦成。
2COR|8|7|既然你們在信心、口才、知識、萬分的熱忱，以及我們對你們 的愛心上，都勝人一等，那麼，當在這慈善的事上也要勝人一等。
2COR|8|8|我說這話，並不是命令你們，而是藉著別人的熱忱來考驗你們愛心的真誠。
2COR|8|9|你們知道我們主耶穌基督的恩典：他本是富足，卻為你們成了貧窮，好使你們因他的貧窮而成為富足。
2COR|8|10|我在這事上把我的意見告訴你們，是對你們有益，因為你們開始辦這事，而且起此心意已經有一年了。
2COR|8|11|如今就當辦成這事，既然有願做的心，也當照你們所有的去辦成。
2COR|8|12|因為人只要有願做的心，必照他所有的蒙悅納，並不是照他所沒有的。
2COR|8|13|我不是要別人輕鬆，你們受累，而是要均勻：
2COR|8|14|就是要你們現在的富餘補他們的不足，使他們的富餘將來也可以補你們的不足，這就均勻了。
2COR|8|15|如經上所記： 多收的沒有餘， 少收的也沒有缺。
2COR|8|16|感謝上帝，把我對你們的熱忱同樣放在 提多 心裏。
2COR|8|17|他固然聽了我的勸告，但自己更加熱心，自願往你們那裏去。
2COR|8|18|我們還差遣一位弟兄和他同去，這人在傳福音的事上得了眾教會的稱讚；
2COR|8|19|不但這樣，他也被眾教會選派跟我們同行，把所交託我們的這捐款送到了，為的是榮耀主，也表明我們的好意。
2COR|8|20|我們這樣做，免得有人因我們收的捐款多而挑剔我們。
2COR|8|21|我們留心做好事，不但在主面前，就是在人面前也是這樣。
2COR|8|22|我們又差遣一位弟兄同去。這人的熱忱，我們在許多事上屢次考驗過，現在他因為深深信任你們，就更加熱心了。
2COR|8|23|至於 提多 ，他是我的夥伴，為服事你們作我的同工。至於那兩位弟兄，他們是眾教會的使者，是基督的榮耀。
2COR|8|24|所以，你們務要在眾教會面前向他們顯明你們的愛心和我所誇獎你們的憑據。
2COR|9|1|關於供給聖徒的事，我本來不必寫信給你們；
2COR|9|2|因為我知道你們的好意，常對 馬其頓 人誇獎你們，說 亞該亞 人預備好已經有一年了。你們的熱心感動了許多人。
2COR|9|3|但我差遣那幾位弟兄去，要使你們照我的話預備妥當，免得我們在這事上誇獎你們的話落了空。
2COR|9|4|萬一有 馬其頓 人與我同去，見你們沒有預備好，就使我們所確信的反成了羞愧；你們的羞愧更不用說了。
2COR|9|5|因此，我想必須鼓勵那幾位弟兄先到你們那裏去，把從前所應許的捐款預備妥當，好顯出你們所捐的是出於樂意，不是出於勉強。
2COR|9|6|還有一點：「少種的少收；多種的多收。」
2COR|9|7|各人要隨心所願，不要為難，不要勉強，因為上帝愛樂捐的人。
2COR|9|8|上帝能將各樣的恩惠多多加給你們，使你們凡事常常充足，能多做各樣善事。
2COR|9|9|如經上所記： 「他施捨，賙濟貧窮； 他的義行存到永遠。」
2COR|9|10|那賜種子給撒種的，賜糧食給人吃的，必多多加給你們種地的種子，又增添你們仁義的果子。
2COR|9|11|你們必凡事富足，能多多施捨，使人藉著我們而生感謝上帝的心。
2COR|9|12|因為辦這供給的事，不但補聖徒的缺乏，而且使許多人對上帝充滿更多的感謝。
2COR|9|13|他們從這供給的事上得了憑據，知道你們宣認基督，順服他的福音，慷慨捐助給他們和眾人，把榮耀歸給上帝。
2COR|9|14|他們也因上帝極大的恩賜顯在你們身上而切切想念你們，為你們祈禱。
2COR|9|15|感謝上帝，因他有說不盡的恩賜！
2COR|10|1|我－ 保羅 與你們見面的時候是溫和的，不在你們那裏的時候向你們是勇敢的，如今親自藉著基督的溫柔和慈祥勸你們。
2COR|10|2|有人認為我們是憑著血氣行事，我認為必須敢於對付這等人；我但求在那裏的時候，不必這樣勇敢。
2COR|10|3|我們雖然在血氣中行事，卻不憑著血氣爭戰。
2COR|10|4|因為我們爭戰的兵器本不是屬血氣的，而是憑著上帝的能力，能夠攻破堅固的營壘。我們攻破各樣的計謀，
2COR|10|5|和各樣攔阻人認識上帝的高壘，又奪回人心來順服基督。
2COR|10|6|我已經預備好了，等你們完全順服的時候來懲罰所有不順服的人。
2COR|10|7|你們只看事情的外表。倘若有人自信是屬基督的，他要再想想，他屬基督，我們也屬基督。
2COR|10|8|主賜給我們權柄，是要造就你們，並不是要拆毀你們；我就是為這權柄稍微誇口也不覺得慚愧。
2COR|10|9|我說這話，免得你們以為我寫信是要恐嚇你們。
2COR|10|10|因為有人說：「他信上的語氣既嚴厲又強硬，他本人卻軟弱無能，言語粗俗。」
2COR|10|11|這等人當明白，我們不在那裏時信上怎麼說，見面時也必怎麼做。
2COR|10|12|因為我們不敢將自己和某些自我推薦的人並列相比；他們用自己度量自己，用自己比較自己，是不明智的。
2COR|10|13|我們不願意過分誇口，但是我們只在上帝劃定的界限內誇口。這界限甚至擴展到你們那裏。
2COR|10|14|我們擴展到你們那裏時並沒有越過了自己的界限，其實我們是首先到你們那裏傳基督福音的。
2COR|10|15|我們不靠別人所勞碌的過分誇口；我們只希望你們信心增長的時候，所劃定給我們的範圍也能夠因著你們更加擴展，
2COR|10|16|使福音得以傳到你們以外的地方，而不在別人的範圍之內，以別人所成就的事誇口。
2COR|10|17|但「要誇耀的，該誇耀主」。
2COR|10|18|因為蒙悅納的，不是自我稱許的，而是主所稱許的。
2COR|11|1|但願你們容忍我小小的愚蠢；請你們務必容忍我。
2COR|11|2|我以上帝嫉妒的愛來愛你們，因為我曾把你們許配給一個丈夫，要把你們如同貞潔的童女獻給基督。
2COR|11|3|我只怕你們的心偏邪了，失去那向基督所獻誠懇貞潔 的心，就像蛇用詭詐誘惑了 夏娃 一樣。
2COR|11|4|假如有人來，傳另一個耶穌，不是我們所傳過的；或者你們另受一個靈，不是你們所受過的聖靈；或者接納另一個福音，不是你們所接納過的；你們居然容忍了！
2COR|11|5|但我想，我一點也不在那些超級使徒以下。
2COR|11|6|雖然我不擅長說話，我的知識卻不如此。這點我們已經在每一方面各樣事上向你們表明了。
2COR|11|7|我貶低自己，為了使你們高升，因為我白白地傳上帝的福音給你們，難道這算是我犯了錯嗎？
2COR|11|8|我剝奪了別的教會，向他們取了報酬來效勞你們。
2COR|11|9|我在你們那裏有缺乏的時候，並沒有連累你們一個人，因為我所缺乏的，那些從 馬其頓 來的弟兄都補足了。我向來凡事謹慎，將來也必謹慎，總不要連累你們。
2COR|11|10|既有基督的真誠在我裏面，在 亞該亞 一帶地方就沒有人能阻止我這樣自誇。
2COR|11|11|為甚麼呢？是因我不愛你們嗎？上帝知道，我愛你們！
2COR|11|12|我現在所做的，將來還要做，為要斷絕那些尋機會之人的機會，不讓他們在所誇耀的事上被人認為與我們一樣。
2COR|11|13|那樣的人是假使徒，行事詭詐，裝作基督的使徒。
2COR|11|14|這也不足為奇，因為連撒但也裝作光明的天使。
2COR|11|15|所以，他的差役若裝作公義的差役也沒有甚麼大不了。他們的結局必然跟他們的行為相符。
2COR|11|16|我再說，誰都不可把我看作愚蠢的；即使你們把我當作愚蠢人，那麼，也讓我稍微誇誇口吧。
2COR|11|17|我說的話不是奉主的權柄說的，而是像愚蠢人具有自信地放膽誇口。
2COR|11|18|既然有好些人憑著血氣在誇口，我也要誇口了。
2COR|11|19|你們是聰明人，竟能甘心容忍愚蠢人！
2COR|11|20|假若有人奴役你們，或侵吞你們，或壓榨你們，或侮辱你們，或打你們的臉，你們居然都能容忍。
2COR|11|21|說來慚愧，在這方面好像我們是太軟弱了。 然而，我說句蠢話，人在甚麼事上敢誇口，我也敢誇口。
2COR|11|22|他們是 希伯來 人嗎？我也是。他們是 以色列 人嗎？我也是。他們是 亞伯拉罕 的後裔嗎？我也是。
2COR|11|23|他們是基督的用人嗎？我說句狂話，我更是。我比他們忍受更多勞苦，坐過更多次監牢，受過無數次的鞭打，常常冒死。
2COR|11|24|我被 猶太 人鞭打五次，每次四十減去一下；
2COR|11|25|被棍打了三次，被石頭打了一次，遭海難三次，一晝一夜在深海裏掙扎。
2COR|11|26|我又屢次行遠路，遭江河的危險，盜賊的危險，同族人的危險，外族人的危險，城裏的危險，曠野的危險，海中的危險，假弟兄的危險。
2COR|11|27|我勞碌困苦，常常失眠，又飢又渴，忍飢耐寒，赤身露體。
2COR|11|28|除了這些外表的事以外，我還有為眾教會操心的事天天壓在我身上。
2COR|11|29|有誰軟弱，我不軟弱呢？有誰跌倒，我不焦急呢？
2COR|11|30|我若必須誇口，就誇我軟弱的事好了。
2COR|11|31|那永遠可稱頌之主耶穌的父上帝知道我不說謊。
2COR|11|32|在 大馬士革 的 亞哩達 王手下的提督把守 大馬士革城 ，要捉拿我，
2COR|11|33|我被人用筐子從城牆上的窗口縋下，逃脫了他的手。
2COR|12|1|雖然自誇無益，我還是不得不誇。我現在要提到主的異象和啟示。
2COR|12|2|我認識一個在基督裏的人，他在十四年前被提到第三層天上去；或在身內，我不知道，或在身外，我也不知道，只有上帝知道。
2COR|12|3|我認識的這樣的一個人—或在身內，或在身外，我都不知道，只有上帝知道—
2COR|12|4|他被提到樂園裏，聽見隱祕的言語，是人不可說的。
2COR|12|5|為這人，我要誇口；但是為我自己，除了我的軟弱以外，我並不誇口。
2COR|12|6|就是我願意誇口也不算狂，因為我會說實話；只是我絕口不談，恐怕有人把我看得太高了，過於他在我身上所看見所聽見的；
2COR|12|7|又恐怕我因所得的啟示太高深，就過於高抬自己，所以 有一根刺加在我身上，就是撒但的差役來折磨我，免得我過於高抬自己。
2COR|12|8|為了這事，我曾三次求主使這根刺離開我。
2COR|12|9|他對我說：「我的恩典是夠你用的，因為我的能力是在人的軟弱上顯得完全。」所以，我更喜歡誇耀自己的軟弱，好使基督的能力覆庇我。
2COR|12|10|為基督的緣故，我以軟弱、凌辱、艱難、迫害、困苦為可喜樂的事；因為我甚麼時候軟弱，甚麼時候就剛強了。
2COR|12|11|我成了愚蠢人，是被你們逼出來的，因為我本該被你們讚許才是。雖然我算不了甚麼，卻沒有一件事在那些超級使徒以下。
2COR|12|12|我在你們中間，用百般的忍耐，藉著神蹟、奇事、異能顯出使徒的憑據來。
2COR|12|13|除了我不曾連累你們這一件事，你們還有甚麼事不及別的教會呢？這不公平之處，請你們饒恕我吧。
2COR|12|14|如今，我準備第三次到你們那裏去。我仍不會連累你們，因為我所求的是你們，不是你們的財物。兒女不該為父母積財，父母該為兒女積財。
2COR|12|15|我也甘心樂意為你們的靈魂費財費力。難道我越愛你們，就越少得你們的愛嗎？
2COR|12|16|罷了，我自己並沒有連累你們，你們卻有人說，我施詭詐，用心計牢籠你們。
2COR|12|17|我所差遣到你們那裏去的人，我何曾藉著他們中的任何人佔過你們的便宜呢？
2COR|12|18|我勸 提多 到你們那裏去，又差遣那位弟兄與他同去， 提多 佔過你們的便宜嗎？我們的行事為人不是同一心靈 嗎？不是同一步伐嗎？
2COR|12|19|你們一直認為我們是在你們面前為自己辯護嗎？其實，我們本是在基督裏當著上帝面前說話。親愛的，一切的事都是為了造就你們。
2COR|12|20|我怕我再來的時候，見你們不合我所期望的，而你們見我也不合你們所期望的。我怕有紛爭、嫉妒、憤怒、自私、毀謗、讒言、狂傲、動亂的事。
2COR|12|21|我怕我再來的時候，我的上帝使我在你們面前蒙羞，並且又因許多人從前犯罪，行污穢、淫亂、放蕩的事，不肯悔改而悲傷。
2COR|13|1|這是我第三次要到你們那裏去。「任何指控都要憑兩個或三個證人的口述才能成立」。
2COR|13|2|對那些犯了罪的人和其餘所有的人，正如我第二次見你們的時候曾說過，現在不在你們那裏再次說：「我若再來，必不寬容。」
2COR|13|3|因為你們想求證基督是否藉著我說話。基督對你們並不是軟弱的，而是在你們裏面大有能力的。
2COR|13|4|他因軟弱被釘在十字架上，卻因上帝的大能仍然活著。我們在他裏面也成為軟弱的，但對你們，我們將因上帝的大能而與他一同活著。
2COR|13|5|你們總要省察自己是否在信仰中生活；你們要考驗自己。除非你們經不起考驗，你們自己豈不應該知道有耶穌基督在你們裏面嗎？
2COR|13|6|我希望你們知道，我們並不是經不起考驗的人。
2COR|13|7|我們祈求上帝使你們不做任何惡事；這不是要顯明我們是經得起考驗的，而是要你們行事端正，即使我們似乎經不起考驗也沒有關係。
2COR|13|8|我們不能做任何對抗真理的事，只能維護真理。
2COR|13|9|當我們軟弱而你們剛強時，我們也歡喜。我們所祈求的是：你們能成為完全人。
2COR|13|10|所以，我不在你們那裏的時候，把這些話寫給你們，好使我見你們的時候不用照主所給我的權柄嚴厲地待你們；這權柄原是為造就人，而不是為摧毀人。
2COR|13|11|末了，弟兄們，願你們喜樂。要追求完全；要接受鼓勵；要同心合意；要彼此和睦。如此，慈愛和平的上帝必與你們同在。
2COR|13|12|你們要用聖潔的吻彼此問安。眾聖徒都向你們問安。
2COR|13|13|願主耶穌基督的恩惠、上帝的慈愛、聖靈的感動常與你們眾人同在！
GAL|1|1|我使徒 保羅 和所有跟我一起的弟兄，寫信給 加拉太 的眾教會。我作使徒不是由於人，也不是藉著人，而是藉著耶穌基督與使他從死人中復活的父上帝。
GAL|1|2|
GAL|1|3|願恩惠、平安 從我們的父上帝和主耶穌基督歸給你們！
GAL|1|4|基督照我們父上帝的旨意，為我們的罪捨己，要救我們脫離現今這罪惡的世代。
GAL|1|5|願榮耀歸給上帝，直到永永遠遠。阿們！
GAL|1|6|我很驚訝你們這麼快就離開那位藉著基督之 恩呼召你們的上帝，而去隨從別的福音；
GAL|1|7|其實並沒有另一個福音，不過有些人騷擾你們，要把基督的福音更改了。
GAL|1|8|但無論是我們或是天上來的使者，若傳福音給你們 ，與我們所傳給你們的不同，他該受詛咒！
GAL|1|9|我們已經說了，現在我再說，若有人傳福音給你們，與你們以往所領受的不同，他該受詛咒！
GAL|1|10|我現在是要得人的心，還是要得上帝的心呢？難道我在討人的喜歡嗎？我若仍舊想討人的喜歡，我就不是基督的僕人了。
GAL|1|11|弟兄們，我要你們知道，我所傳的福音不是按照人的意思；
GAL|1|12|因為我不是從人領受的，也不是人教導我的，而是藉著耶穌基督的啟示而來。
GAL|1|13|你們聽說過從前我在 猶太 教中的行徑，我怎樣竭力壓迫殘害上帝的教會。
GAL|1|14|在 猶太 教中，我比本國許多同輩的人更激進，為我祖宗的傳統更熱心。
GAL|1|15|然而，那位把我從母腹裏分別出來、又施恩呼召我的上帝 ，既然樂意
GAL|1|16|把他兒子啟示在我心裏，讓我在外邦人中傳揚他，我就沒有跟有血有肉的人商量，
GAL|1|17|也沒有上 耶路撒冷 去見那些比我先作使徒的，惟獨到 阿拉伯 去，後來又回到 大馬士革 。
GAL|1|18|過了三年，我才上 耶路撒冷 去見 磯法 ，和他同住了十五天。
GAL|1|19|至於別的使徒，除了主的兄弟 雅各 ，我都沒有見過。
GAL|1|20|我現在寫給你們的是在上帝面前說的，不說謊話。
GAL|1|21|以後我到了 敘利亞 和 基利家 一帶；
GAL|1|22|那時，在基督裏的 猶太 各教會都沒有見過我的面。
GAL|1|23|不過他們聽說「那從前壓迫我們的，現在竟傳揚他原先所殘害的信仰」。
GAL|1|24|他們就為我的緣故歸榮耀給上帝。
GAL|2|1|過了十四年，我再上 耶路撒冷 去， 巴拿巴 同行，也帶了 提多 一起去。
GAL|2|2|我是奉了啟示上去的；我把在外邦人中所傳的福音對弟兄們說明，我是私下對那些有名望的人說的，免得我現在或是從前都徒然奔跑了。
GAL|2|3|但跟我同去的 提多 ，雖是 希臘 人，也沒有勉強他受割禮；
GAL|2|4|因為有偷著混進來的假弟兄，暗中窺探我們在基督耶穌裏擁有的自由，要使我們作奴隸，
GAL|2|5|可是，為要使福音的真理仍存在你們中間，我們一點也沒有讓步順服他們。
GAL|2|6|至於那些有名望的，不論他們是何等人，都與我無關；上帝不以外貌取人。那些有名望的，並沒有加增我甚麼。
GAL|2|7|相反地，他們看見了主託付我傳福音給未受割禮的人，正如主託付 彼得 傳福音給受割禮的人；
GAL|2|8|那感動 彼得 、叫他為受割禮的人作使徒的，也感動我，叫我為外邦人作使徒。
GAL|2|9|那些被認為是教會柱石的 雅各 、 磯法 、 約翰 知道上帝所賜給我的恩典，就跟我和 巴拿巴 握右手以示合作，同意我們往外邦人那裏去，他們往受割禮的人那裏去。
GAL|2|10|他們只要求我們記念窮人，這也是我一向熱心在做的。
GAL|2|11|後來， 磯法 到了 安提阿 ，因為他有可責之處，我就當面反對他。
GAL|2|12|從 雅各 那裏來的人未到以前，他和外邦人一同吃飯，及至他們來到，他因怕奉割禮的人就退出，跟外邦人疏遠了。
GAL|2|13|其餘的 猶太 人也都隨著他裝假，甚至連 巴拿巴 也隨夥裝假。
GAL|2|14|但我一看見他們做得不對，與福音的真理不合，就在眾人面前對 磯法 說：「你既是 猶太 人，卻按照外邦人的樣子，不按照 猶太 人的樣子生活，怎麼能勉強外邦人按照 猶太 人的樣子生活呢？」
GAL|2|15|我們生來就是 猶太 人，不是外邦罪人；
GAL|2|16|可是我們知道，人稱義不是因律法的行為，而是因信耶穌基督 ，我們也信了基督耶穌，為要使我們因信基督稱義，不因律法的行為稱義，因為，凡血肉之軀沒有一個能因律法的行為稱義。
GAL|2|17|我們若求在基督裏稱義，自己卻還被視為罪人，那麼，基督是罪的用人嗎？絕對不是！
GAL|2|18|如果我重新建造我所拆毀的，這就證明自己是違犯律法的人。
GAL|2|19|我因律法而向律法死了，使我可以向上帝活著。我已經與基督同釘十字架，
GAL|2|20|現在活著的不再是我，乃是基督在我裏面活著；並且我如今在肉身活著，是因信上帝的兒子而活；他是愛我，為我捨己。
GAL|2|21|我不廢掉上帝的恩；如果義是藉著律法而獲得，那麼基督就白白死了。
GAL|3|1|無知的 加拉太 人哪，耶穌基督釘十字架，已經活現在你們眼前，誰又迷惑了你們呢？
GAL|3|2|這是我惟一要問你們的：你們領受了聖靈，是因律法的行為或是因聽信福音呢？
GAL|3|3|你們既然以聖靈開始，如今竟要以肉身終結嗎？你們是這樣的無知嗎？
GAL|3|4|你們受這麼多的苦都是徒然的嗎？如果真是徒然的，
GAL|3|5|那麼，上帝賜給你們聖靈，又在你們中間行異能，是因律法的行為或是因聽信福音呢？
GAL|3|6|正如 亞伯拉罕 「信了上帝，這就算他為義」。
GAL|3|7|所以，你們知道：有信心的人才是 亞伯拉罕 的子孫。
GAL|3|8|聖經既然預先看見上帝要使外邦人因信稱義，預先傳福音給 亞伯拉罕 ，說：「萬國都必因你得福。」
GAL|3|9|可見，那有信心的人和有信心的 亞伯拉罕 一同得福。
GAL|3|10|凡出於律法的行為都是受詛咒的，因為經上記著：「凡不持守律法書上所記的一切而去行的，都是受詛咒的。」
GAL|3|11|沒有一個人靠著律法在上帝面前稱義，這是明顯的，因為經上說：「義人必因信得生。」
GAL|3|12|律法並不出於信，而是說：「行這些事的就必因此得生。」
GAL|3|13|既然基督為我們成了詛咒，就把我們從律法的詛咒中贖出來。因為經上記著：「凡掛在木頭上的都是受詛咒的。」
GAL|3|14|這是要使 亞伯拉罕 的福，因著基督耶穌臨到外邦人，使我們能因信得著所應許的聖靈。
GAL|3|15|弟兄們，我照著人的觀點說，人的遺囑一經確定，沒有人能廢棄或加增。
GAL|3|16|那些應許原是向 亞伯拉罕 和他後裔說的，並不是說「和眾後裔」，指許多人，而是說「和你那個後裔」，指一個人，就是基督。
GAL|3|17|我是這麼說，上帝預先所立的約不能被四百三十年以後的律法廢掉，使應許失效。
GAL|3|18|因為承受產業若是出於律法，就不再是出於應許；但上帝是憑著應許把產業賜給 亞伯拉罕 。
GAL|3|19|這樣說來，為甚麼要有律法呢？律法是為過犯的緣故而加上去的，等候那蒙應許的子孫來到才結束，是藉著天使經中保之手而設立的。
GAL|3|20|但中保本不是為單方設立的；上帝卻是一位。
GAL|3|21|這樣，律法是與上帝的 應許對立嗎？絕對不是！如果律法的頒佈能使人得生命，義就誠然出於律法了。
GAL|3|22|但聖經把萬物都圈在罪裏，為要使因信耶穌基督 而來的應許歸給信的人。
GAL|3|23|但這「信」還未來以前，我們被看守在律法之下，像被圈住，直到那將來的「信」顯明出來。
GAL|3|24|這樣，律法是我們的啟蒙教師，直到基督來了 ，好使我們因信稱義。
GAL|3|25|但這「信」既然來到，我們從此就不在啟蒙教師的手下了。
GAL|3|26|其實，你們藉著信，在基督耶穌裏都成為上帝的兒女。
GAL|3|27|你們凡受洗歸入基督的都披戴基督了：
GAL|3|28|不再分 猶太 人或 希臘 人，不再分為奴的自主的，不再分男的女的，因為你們在基督耶穌裏都成為一了。
GAL|3|29|既然你們屬於基督，你們就是 亞伯拉罕 的子孫，是照著應許承受產業的了。
GAL|4|1|我說，雖然那承受產業的是整個產業的主人，但在未成年的時候卻與奴隸毫無分別，
GAL|4|2|仍是在監護人和管家的手下，直等他父親預定的時候來到。
GAL|4|3|我們也是一樣，在未成年的時候，被世上粗淺的學說 所奴役，也是如此。
GAL|4|4|等到時候成熟，上帝就差遣他的兒子，為女子所生，且生在律法之下，
GAL|4|5|為要把律法之下的人贖出來，使我們獲得兒子的名分。
GAL|4|6|因為你們是兒子，上帝就差他兒子的靈進入我們 的心，呼叫：「阿爸，父！」
GAL|4|7|可見，你不再是奴隸，而是兒子了，既然是兒子，就靠著上帝也成為後嗣了。
GAL|4|8|但從前不認識上帝的時候，你們是給那些本來不是上帝的神明作奴隸；
GAL|4|9|現在你們既然認識上帝，更可說是被上帝所認識的，怎麼還要轉回那懦弱無用的粗淺學說 ，情願再給它們作奴隸呢？
GAL|4|10|你們竟又謹守日子、月份、節期、年份，
GAL|4|11|我為你們擔心，惟恐我在你們身上是枉費工夫了。
GAL|4|12|弟兄們，我勸你們，要像我一樣，因為我也像你們一樣。你們一點沒有虧負我。
GAL|4|13|你們知道，我因為身體有疾病才有第一次傳福音給你們的機會。
GAL|4|14|雖然你們為我身體的緣故受試煉，卻沒有輕看我，也沒有厭棄我，反倒接待我如同上帝的使者，如同基督耶穌。
GAL|4|15|你們當日的好意哪裏去了呢？那時若辦得到，你們就是把自己的眼睛挖出來給我，也都情願。這是我可以給你們作證的。
GAL|4|16|如今我把真理告訴你們，倒成了你們的仇敵嗎？
GAL|4|17|那些熱心待你們的人，不懷好意，是要隔絕你們，好使你們熱心待他們。
GAL|4|18|在善事上，時刻熱心待別人原是好的，卻不只是我與你們同在的時候才這樣。
GAL|4|19|我的孩子們哪，我為你們再受生產之苦，直等到基督成形在你們心裏 。
GAL|4|20|我期望現今就在你們那裏，可以改變我的口氣，因為我為你們心裏難過。
GAL|4|21|你們這願意在律法之下的人，請告訴我，你們沒有聽見律法嗎？
GAL|4|22|因為律法上記著， 亞伯拉罕 有兩個兒子，一個是使女生的，一個是自由的婦人生的。
GAL|4|23|那使女所生的是按著肉體生的；那自由的婦人所生的是憑著應許生的。
GAL|4|24|這是比方：那兩個婦人就是兩個約；一個婦人是出於 西奈山 ，生子為奴，就是 夏甲 。
GAL|4|25|這 夏甲 是指著 阿拉伯 的 西奈山 ，與現在的 耶路撒冷 同類，因為 耶路撒冷 和她的兒女都是為奴的。
GAL|4|26|但另一婦人就是在上的 耶路撒冷 ，是自由的，她是我們的母親。
GAL|4|27|因為經上記著： 不懷孕、不生養的，你要歡樂； 未曾經過產難的，你要高聲歡呼； 因為沒有丈夫的，比有丈夫的有更多的兒女。
GAL|4|28|弟兄們，你們是憑著應許作兒女的，如同 以撒 一樣。
GAL|4|29|當時，那按著肉體生的迫害了那按著聖靈生的，現在也是這樣。
GAL|4|30|然而經上是怎麼說的呢？是說：「把使女和她兒子趕出去！因為使女的兒子絕不能與自由婦人的兒子一同承受產業。」
GAL|4|31|弟兄們，這樣看來，我們不是使女的兒女，而是自由婦人的兒女了。
GAL|5|1|基督釋放了我們，為使我們得自由。所以要站穩了，不要再被奴隸的軛挾制。
GAL|5|2|我— 保羅 告訴你們，你們若受割禮，基督就對你們無益了。
GAL|5|3|我再指著凡受割禮的人確實地說，他有義務遵行全部的律法。
GAL|5|4|你們這要靠律法稱義的是與基督隔絕，從恩典中墜落了。
GAL|5|5|至於我們，我們是靠著聖靈，憑著信心，等候所盼望的義。
GAL|5|6|因為在基督耶穌裏，受割禮不受割禮都沒有功效，惟獨使人發出仁愛的信心才有功效。
GAL|5|7|你們向來跑得好，誰攔阻了你們，使你們不順從真理呢？
GAL|5|8|這樣的勸導不是出於那召你們的。
GAL|5|9|一點麵酵能使全團都發起來。
GAL|5|10|我在主裏深信你們必不懷別樣的心；但騷擾你們的，無論是誰，必須承受懲罰。
GAL|5|11|弟兄們，我若仍舊傳割禮，為甚麼還受迫害呢？若是這樣，十字架絆倒人的地方就沒有了。
GAL|5|12|恨不得那騷擾你們的人把自己閹割了。
GAL|5|13|弟兄們，你們蒙召是要得自由；只是不可把這自由當作放縱情慾的機會，總要用愛心互相服侍。
GAL|5|14|因為全部律法都包括在「愛鄰 如己」這一句話之內了。
GAL|5|15|你們要謹慎，你們若相咬相吞，恐怕要彼此消滅了。
GAL|5|16|我說，你們要順著聖靈而行，絕不可滿足肉體的情慾。
GAL|5|17|因為肉體的情慾和聖靈相爭，聖靈和肉體相爭，這兩個彼此敵對，使你們不能做所願意做的。
GAL|5|18|但你們若被聖靈引導，就不在律法之下。
GAL|5|19|情慾的事都是顯而易見的；就如淫亂、污穢、放蕩、
GAL|5|20|拜偶像、行邪術、仇恨、紛爭、忌恨、憤怒、自私、分派、結黨、
GAL|5|21|嫉妒 、醉酒、荒宴等類。我從前告訴過你們，現在又告訴你們，做這樣事的人必不能承受上帝的國。
GAL|5|22|聖靈的果子就是仁愛、喜樂、和平、忍耐、恩慈、良善、信實、
GAL|5|23|溫柔、節制。這樣的事沒有律法禁止。
GAL|5|24|凡屬基督耶穌 的人，是已經把肉體與肉體的邪情私慾同釘在十字架上了。
GAL|5|25|我們若靠著聖靈而活，也要靠著聖靈行事。
GAL|5|26|不要貪圖虛名，彼此惹氣，互相嫉妒。
GAL|6|1|弟兄們，若有人偶然被過犯所勝，你們屬靈的人就要用溫柔的心把他挽回過來；自己也要留意，免得也被引誘。
GAL|6|2|你們各人的重擔要互相擔當，這樣就會成全 基督的律法。
GAL|6|3|人若沒有甚麼了不起，還自以為了不起的，就是自欺。
GAL|6|4|各人要省察自己的行為；這樣，他所誇口的只在自己，而不在別人。
GAL|6|5|因為人人必須擔當自己的擔子。
GAL|6|6|在真道上受教的，要把一切美好的東西與施教的人分享。
GAL|6|7|不要自欺；上帝是輕慢不得的，因為人種的是甚麼，收的也是甚麼。
GAL|6|8|順著肉體撒種的，必從肉體收敗壞；順著聖靈撒種的，必從聖靈收永生。
GAL|6|9|我們行善不可喪志，因為若不灰心，到了適當的時候就有收成。
GAL|6|10|所以，一有機會就要向眾人行善，向信徒一家的人更要這樣。
GAL|6|11|你們看我親手寫給你們的字是何等的大！
GAL|6|12|那些想要炫耀外表的人才勉強你們受割禮，無非是怕自己為基督的十字架受迫害。
GAL|6|13|他們那些受割禮的，連自己也不守律法；他們要你們受割禮，不過是要拿你們的肉體誇口。
GAL|6|14|但我絕不以別的誇口，只誇我們主耶穌基督的十字架；因這十字架 ，就我而論，世界已經釘在十字架上；就世界而論，我已經釘在十字架上。
GAL|6|15|受割禮或不受割禮都無關緊要，要緊的就是作新造的人。
GAL|6|16|凡照這準則行的人，願平安 憐憫，加給他們，和上帝的 以色列 民。
GAL|6|17|從今以後，不要有人再攪擾我，因為我身上帶著耶穌的印記。
GAL|6|18|弟兄們，願我們主耶穌基督的恩與你們的靈同在。阿們！
EPH|1|1|奉上帝旨意作基督耶穌使徒的 保羅 ，寫信給在 以弗所 的 眾聖徒，就是在基督耶穌裏忠心的人。
EPH|1|2|願恩惠、平安 從我們的父上帝和主耶穌基督歸給你們！
EPH|1|3|願頌讚歸給我們主耶穌基督的父上帝。他在基督裏曾把天上各樣屬靈的福氣賜給我們。
EPH|1|4|因為他從創世以前，在基督裏揀選了我們，使我們在他面前成為聖潔，沒有瑕疵，滿有愛心。
EPH|1|5|他按著自己旨意所喜悅的 ，預定我們藉著耶穌基督得兒子的名分，
EPH|1|6|使他榮耀的恩典得到稱讚；這恩典是他在愛子裏白白賜給我們的。
EPH|1|7|我們藉著這愛子的血得蒙救贖，過犯得以赦免，這是照他豐富的恩典，
EPH|1|8|充充足足地賞給我們的。他以諸般的智慧聰明，
EPH|1|9|照自己在基督裏所立定的美意，使我們知道他旨意的奧祕，
EPH|1|10|要照著所安排的，在時機成熟的時候，使天上、地上、一切所有的，都在基督裏面同歸於一。
EPH|1|11|我們也在他裏面得了基業；這原是那位隨己意行萬事的上帝照著自己的旨意所預定的，
EPH|1|12|為要使我們，這些首先把希望寄託在基督裏的人，頌讚他的榮耀。
EPH|1|13|在基督裏你們聽見真理的道，就是那使你們得救的福音，你們也信了他，就受了所應許的聖靈為印記。
EPH|1|14|這聖靈是我們得基業的憑據，直等到上帝的子民得救贖，使他的榮耀得到稱讚。
EPH|1|15|因此，我既然聽見你們對主耶穌有信心，對眾聖徒有愛心，
EPH|1|16|就不住地為你們感謝上帝，禱告的時候常常提到你們，
EPH|1|17|求我們主耶穌基督的上帝，榮耀的父，把那賜人智慧和啟示的靈賜給你們，使你們真正認識他，
EPH|1|18|照亮你們心中的眼睛，使你們知道他呼召你們來得的指望是甚麼，他在聖徒中所得榮耀的基業是何等豐盛，
EPH|1|19|並知道他向我們這些信的人所顯的能力是何等浩大，這是照他的大能大力運行的。
EPH|1|20|這大能曾運行在基督身上，使他從死人中復活，又使他在天上坐在自己的右邊，
EPH|1|21|遠超越一切執政的、掌權的、有權能的、統治的和一切有名號的；不但是今世的，連來世的也都超越了。
EPH|1|22|上帝使萬有服在他的腳下，又使他為了教會作萬有之首；
EPH|1|23|教會是他的身體，是那充滿萬有者所充滿的。
EPH|2|1|從前，你們因著自己的過犯罪惡而死了。
EPH|2|2|那時，你們在過犯罪惡中生活，隨從今世的風俗，順服空中掌權者的領袖，就是現今在悖逆的人心中運行的邪靈。
EPH|2|3|我們從前也都生活在他們當中，放縱肉體的私慾，隨著肉體和心中的意念去做，和別人一樣，生來就是該受懲罰的人。
EPH|2|4|然而，上帝有豐富的憐憫，因著他愛我們的大愛，
EPH|2|5|竟在我們因過犯而死了的時候，使我們與基督一同活過來—可見你們得救是本乎恩—
EPH|2|6|他又使我們在基督耶穌裏與他一同復活，一同坐在天上，
EPH|2|7|為要把他極豐富的恩典，就是他在基督耶穌裏向我們所施的恩慈，顯明給後來的世代。
EPH|2|8|你們得救是本乎恩，也因著信；這並不是出於自己，而是上帝所賜的；
EPH|2|9|也不是出於行為，免得有人自誇。
EPH|2|10|我們是他所造之物，在基督耶穌裏創造的，為要使我們行善，就是上帝早已預備好要我們做的。
EPH|2|11|所以，你們要記得：從前你們按肉體是外邦人，是「沒受割禮的」；這名字是那些憑人手在肉身上「受割禮的人」所取的。
EPH|2|12|要記得那時候，你們與基督無關，與 以色列 選民團體隔絕，在所應許的約上是局外人，而且在世上沒有指望，沒有上帝。
EPH|2|13|從前你們是遠離上帝的人，如今卻在基督耶穌裏，靠著他的血，已經得以親近了。
EPH|2|14|因為他自己是我們的和平 ，使雙方合而為一，拆毀了中間隔絕的牆，而且以自己的身體終止了冤仇，
EPH|2|15|廢掉那記在律法上的規條，為要使兩方藉著自己造成一個新人，促成了和平；
EPH|2|16|既在十字架上消滅了冤仇，就藉這十字架使雙方歸為一體，與上帝和好，
EPH|2|17|並且來傳和平的福音給你們遠處的人，也傳和平給那些近處的人，
EPH|2|18|因為我們雙方藉著他，在同一位聖靈裏得以進到父面前。
EPH|2|19|這樣，你們不再是外人或客旅，是與聖徒同國，是上帝家裏的人了，
EPH|2|20|被建造在使徒和先知的根基上，而基督耶穌自己為房角石，
EPH|2|21|靠著他整座房子連接得緊湊，漸漸成為在主裏的聖殿。
EPH|2|22|你們也靠他同被建造，成為上帝藉著聖靈居住的所在。
EPH|3|1|因此，我— 保羅 為你們外邦人作了基督耶穌 囚徒的，替你們祈禱 。
EPH|3|2|想你們必曾聽見上帝賜恩給我，把關切你們的職分託付我，
EPH|3|3|用啟示讓我知道福音的奧祕，正如我以前略略寫過的。
EPH|3|4|你們讀了，就會知道我深深了解基督的奧祕；
EPH|3|5|這奧祕在以前的世代沒有讓人知道，像如今藉著聖靈向他的聖使徒和先知啟示一樣，
EPH|3|6|就是外邦人在基督耶穌裏，藉著福音，得以同為後嗣，同為一體，同為蒙應許的人。
EPH|3|7|我作了這福音的僕役，是照著上帝的恩賜，是照他運行的大能賜給我的。
EPH|3|8|雖然我比眾聖徒中最小的還小，他還賜我這恩典，讓我把基督那測不透的豐富傳給外邦人，
EPH|3|9|又使眾人都明白 甚麼是歷代以來隱藏在創造萬物之上帝裏的奧祕，
EPH|3|10|為要在現今藉著教會使天上執政的、掌權的知道上帝百般的智慧。
EPH|3|11|這是照著上帝在我們主基督耶穌裏所完成的永恆的計劃。
EPH|3|12|我們因信耶穌 ，就在他裏面放膽無懼，滿有自信地進到上帝面前。
EPH|3|13|所以我求你們，不要因我為你們所受的患難喪膽；這原是你們的光榮。
EPH|3|14|因此，我在父面前屈膝—
EPH|3|15|天上地上的各家都是從他得名的－
EPH|3|16|為要他按著他豐盛的榮耀，藉著他的靈，使你們內心的力量剛強起來；
EPH|3|17|又要他使基督因著你們的信住在你們心裏，使你們既在愛中生根立基，
EPH|3|18|能夠和眾聖徒一同明白基督的愛是何等的長、闊、高、深，並知道這愛是超過人的知識所能測度的，為要使你們充滿上帝一切的豐盛。
EPH|3|19|
EPH|3|20|上帝能照著運行在我們心裏的大能充充足足地成就一切，超過我們所求所想的。
EPH|3|21|願他在教會中，並在基督耶穌裏，得著榮耀，直到世世代代，永永遠遠。阿們！
EPH|4|1|我為主作囚徒的勸你們，既然蒙召，行事為人就要與你們所蒙的呼召相稱。
EPH|4|2|凡事要謙虛、溫柔、忍耐，用愛心互相寬容，
EPH|4|3|以和平彼此聯繫，竭力保持聖靈所賜的合一。
EPH|4|4|身體只有一個，聖靈只有一位，正如你們蒙召，是為同有一個指望而蒙召，
EPH|4|5|一主，一信，一洗，
EPH|4|6|一上帝－就是萬人之父，超越萬有之上，貫通萬有，在萬有之中。
EPH|4|7|我們每個人蒙恩都是照基督所量給每個人的恩賜。
EPH|4|8|所以有話說： 「他升上高天的時候，擄掠了俘虜， 將各樣的恩賜賞給人。」
EPH|4|9|既說「他升上」，豈不是指他曾降到地底下嗎？
EPH|4|10|那降下的，就是高升遠超越諸天之上的，為要充滿萬有。
EPH|4|11|他所賜的有使徒，有先知，有傳福音的，有牧者和教師，
EPH|4|12|為要裝備聖徒，做事奉的工作，建立基督的身體，
EPH|4|13|直等到我們眾人在信仰上同歸於一，認識上帝的兒子，得以長大成人，達到基督完全長成的身量。
EPH|4|14|這樣，我們不再作小孩子，中了人的詭計和欺騙的法術，被一切邪說之風搖動，飄來飄去。
EPH|4|15|我們反而要用愛心說誠實話，各方面向著基督長進，連於元首基督，
EPH|4|16|靠著他全身都連接得緊湊，百節各按各職，照著各體的功用彼此相助，使身體漸漸增長，在愛中建立自己。
EPH|4|17|所以我這樣說，且在主裏鄭重地說，你們行事為人，不要再像外邦人存虛妄的心而活。
EPH|4|18|他們心地昏昧，因自己無知，心裏剛硬而與上帝所賜的生命隔絕了。
EPH|4|19|既然他們已經麻木，就放縱情慾，貪婪地行種種污穢的事。
EPH|4|20|但你們從基督學的不是這樣。
EPH|4|21|如果你們聽過他的道，領了他的教，因為真理就在耶穌裏，
EPH|4|22|你們要脫去從前的行為，脫去舊我；這舊我是因私慾的迷惑而漸漸敗壞的。
EPH|4|23|你們要把自己的心志更新，
EPH|4|24|並且穿上新我；這新我是照著上帝的形像造的，有從真理來的公義和聖潔。
EPH|4|25|所以，你們要棄絕謊言，每個人要與鄰舍說誠實話，因為我們是互為肢體。
EPH|4|26|即使生氣也不要犯罪；不可含怒到日落，
EPH|4|27|不可給魔鬼留地步。
EPH|4|28|偷竊的，不要再偷；總要勤勞，親手 做正當的事，這樣才可以把自己有的，分給有缺乏的人。
EPH|4|29|一句壞話也不可出口，只要隨著需要說造就人的好話，讓聽見的人得益處。
EPH|4|30|不要使上帝的聖靈擔憂，你們原是受了他的印記，等候得救贖的日子來到。
EPH|4|31|一切苦毒、憤怒、惱恨、嚷鬧、毀謗，和一切的惡毒都要從你們中間除掉。
EPH|4|32|要仁慈相待，存憐憫的心，彼此饒恕，正如上帝在基督裏饒恕了你們一樣。
EPH|5|1|所以，作為蒙慈愛的兒女，你們該效法上帝。
EPH|5|2|要憑愛心行事，正如基督愛我們，為我們捨了自己，當作馨香的供物和祭物獻給上帝。
EPH|5|3|至於淫亂和一切污穢，或是貪婪，在你們中間連提都不可，這才合乎聖徒的體統。
EPH|5|4|淫詞、妄語和粗俗的俏皮話都不合宜；總要說感謝的話。
EPH|5|5|要確實知道，無論是淫亂的，是污穢的，是貪心的（貪心的就是拜偶像的），在基督和上帝的國裏都得不到基業。
EPH|5|6|不要被人虛浮的話欺騙了，因這些事，上帝的憤怒必臨到那些悖逆的人。
EPH|5|7|所以，不要與他們同夥。
EPH|5|8|從前你們是暗昧的，但如今在主裏面是光明的，行事為人要像光明的子女—
EPH|5|9|光明所結的果子就是一切的良善、公義、誠實。
EPH|5|10|總要察驗甚麼是主所喜悅的事。
EPH|5|11|那暗昧無益的事，不可參與，倒要把這種事揭發出來。
EPH|5|12|因為，他們暗中所做的，就是連提起來都是可恥的。
EPH|5|13|凡被光所照明的都顯露出來，
EPH|5|14|因為使一切顯露出來的就是光。所以有話說： 「你這睡著的人醒過來吧！ 要從死人中復活， 基督要光照你了。」
EPH|5|15|你們要謹慎行事，不要像無知的人，要像智慧的人。
EPH|5|16|要把握時機 ，因為現今的世代邪惡。
EPH|5|17|不要作糊塗人，要明白主的旨意如何。
EPH|5|18|不要醉酒，酒能使人放蕩；要被聖靈充滿。
EPH|5|19|要用詩篇、讚美詩、靈歌彼此對說，口唱心和地讚美主。
EPH|5|20|凡事要奉我們主耶穌基督的名常常感謝父上帝。
EPH|5|21|要存敬畏基督的心彼此順服。
EPH|5|22|作妻子的，你們要順服自己的丈夫，如同順服主。
EPH|5|23|因為丈夫是妻子的頭，如同基督是教會的頭；他又是這身體的救主。
EPH|5|24|教會怎樣順服基督，妻子也要怎樣凡事順服丈夫。
EPH|5|25|作丈夫的，你們要愛自己的妻子，正如基督愛教會，為教會捨己，
EPH|5|26|以水藉著道把教會洗淨，使她成為聖潔，
EPH|5|27|好獻給自己，作榮耀的教會，毫無玷污、皺紋等類的缺陷，而是聖潔沒有瑕疵的。
EPH|5|28|丈夫也應當照樣愛妻子，如同愛自己的身體；愛妻子就是愛自己了。
EPH|5|29|從來沒有人恨惡自己的身體，總是保養愛惜，正像基督待教會一樣，
EPH|5|30|因我們是他身體的肢體。
EPH|5|31|「為這個緣故，人要離開父母，與妻子結合，二人成為一體。」
EPH|5|32|這是極大的奧祕，而我是指基督和教會說的。
EPH|5|33|然而，你們每個人都要愛妻子，如同愛自己一樣；妻子也要敬重她的丈夫。
EPH|6|1|作兒女的，你們要在主裏 聽從父母，這是理所當然的。
EPH|6|2|當孝敬父母，使你得福，在世長壽。這是第一條帶應許的誡命。
EPH|6|3|
EPH|6|4|作父親的，你們不要激怒兒女，但要照著主的教導和勸戒養育他們。
EPH|6|5|作僕人的，你們要懼怕戰兢，用誠實的心聽從你們肉身的主人，好像聽從基督一般；
EPH|6|6|不要只在人的眼前這樣做，像僅是討人的喜歡，而是作基督的僕人，從心裏遵行上帝的旨意，
EPH|6|7|甘心服侍，好像服侍主，不像服侍人，
EPH|6|8|因為知道每個人所做的善事，不論是為奴的或是自主的，都必按所做的從主得到賞賜。
EPH|6|9|作主人的，你們待僕人也是一樣，不要威嚇他們，因為知道他們和你們在天上同有一位主，他並不偏待人。
EPH|6|10|最後，你們要靠著主，依賴他的大能大力作剛強的人。
EPH|6|11|要穿戴上帝所賜的全副軍裝，好抵擋魔鬼的詭計。
EPH|6|12|因為我們的爭戰並不是對抗有血有肉的人，而是對抗那些執政的、掌權的、管轄這幽暗世界的，以及天空靈界的惡魔。
EPH|6|13|所以，要拿起上帝所賜的全副軍裝，好在邪惡的日子能抵擋仇敵，並且完成了一切後還能站立得住。
EPH|6|14|所以，要站穩了，用真理當作帶子束腰，用公義當作護心鏡遮胸，
EPH|6|15|又用和平的福音當作預備走路的鞋穿在腳上。
EPH|6|16|此外，要拿信德當作盾牌，用來撲滅那惡者一切燒著的箭。
EPH|6|17|要戴上救恩的頭盔，拿著聖靈的寶劍—就是上帝的道。
EPH|6|18|要靠著聖靈，隨時多方禱告祈求，並要為此警醒不倦，為眾聖徒祈求。
EPH|6|19|也要為我祈求，讓我有口才，能放膽開口講明福音的奧祕，
EPH|6|20|我為這福音的奧祕作了帶鐵鏈的使者，讓我能照著當盡的本分放膽宣講。
EPH|6|21|今有親愛、忠心服事主的弟兄 推基古 ，為了你們也明白我的事情和我的景況，他會讓你們知道一切的事。
EPH|6|22|我特意打發他到你們那裏去，好讓你們知道我們的情況，又讓他安慰你們的心。
EPH|6|23|願平安 、慈愛、信心從父上帝和主耶穌基督歸給弟兄們。
EPH|6|24|願所有恆心愛我們主耶穌基督的人都蒙恩惠。
PHIL|1|1|基督耶穌的僕人 保羅 和 提摩太 寫信給住 腓立比 、在基督耶穌裏的眾聖徒，以及諸位監督和執事。
PHIL|1|2|願恩惠、平安 從我們的父上帝和主耶穌基督歸給你們！
PHIL|1|3|我每逢想念你們，就感謝我的上帝，
PHIL|1|4|每逢為你們眾人祈求的時候，總是歡歡喜喜地祈求，
PHIL|1|5|因為從第一天直到如今，你們都同心合意興旺福音。
PHIL|1|6|我深信，那在你們心裏動了美好工作的，到了耶穌基督的日子必完成這工作。
PHIL|1|7|我為你們眾人有這樣的想法原是應當的，因為你們常在我心裏；無論我是在捆鎖中，在辯明並證實福音的時候，你們都與我一同蒙恩。
PHIL|1|8|我以基督耶穌的心腸切切想念你們眾人，這是上帝可以為我作證的。
PHIL|1|9|我所禱告的就是：要你們的愛心，在知識和各樣見識上，不斷增長，
PHIL|1|10|使你們能分辨是非，在基督的日子作真誠無可指責的人，
PHIL|1|11|更靠著耶穌基督結滿仁義的果子，歸榮耀稱讚給上帝。
PHIL|1|12|弟兄們，我要你們知道，我所遭遇的事反而使福音更興旺，
PHIL|1|13|以致御營全軍和其餘的人都知道我是為基督的緣故受捆鎖的；
PHIL|1|14|而且那在主裏的弟兄，多半都因我受的捆鎖而篤信不疑，越發放膽無所懼怕地傳道。
PHIL|1|15|有些人傳基督是出於嫉妒紛爭；有些人是出於好意。
PHIL|1|16|後者是出於愛心，知道我奉差遣是為福音辯護的。
PHIL|1|17|前者傳基督是出於自私，動機不純，企圖要加增我捆鎖的苦楚。
PHIL|1|18|這又何妨呢？或是假意或是真心，無論如何，只要基督被傳開了，為此我就歡喜。 我還要歡喜，
PHIL|1|19|因為我知道，這事藉著你們的祈禱和耶穌基督的靈的幫助，終必使我得到釋放。
PHIL|1|20|這就是我所切慕、所盼望的：沒有一事能使我羞愧；反倒凡事坦然無懼，無論是生是死，總要讓基督在我身上照常顯大。
PHIL|1|21|因為我活著就是基督，死了就有益處。
PHIL|1|22|但是，我在肉身活著，若能有工作的成果，我就不知道該挑選甚麼。
PHIL|1|23|我處在兩難之間：我情願離世與基督同在，因為這是好得無比的；
PHIL|1|24|然而，我為你們肉身活著更加要緊。
PHIL|1|25|既然我這樣深信，就知道仍要留在世間，且與你們眾人一起存留，使你們在所信的道上又長進又喜樂，
PHIL|1|26|為了我再到你們那裏時，你們在基督耶穌裏的誇耀越發加增。
PHIL|1|27|最重要的是：你們行事為人要與基督的福音相稱，這樣，無論我來見你們，或不在你們那裏，都可以聽到你們的景況，知道你們同有一個心志，站立得穩，為福音的信仰齊心努力，
PHIL|1|28|絲毫不怕敵人的威脅；以此證明他們會沉淪，你們會得救，這是出於上帝。
PHIL|1|29|因為你們蒙恩，不但得以信服基督，而且要為他受苦。
PHIL|1|30|你們的爭戰，就與你們曾在我身上見過、現在所聽到的是一樣的。
PHIL|2|1|所以，在基督裏若有任何勸勉，若有任何愛心的安慰，若有任何聖靈的團契，若有任何慈悲憐憫，
PHIL|2|2|你們就要意志相同，愛心相同，有一致的心思，一致的想法，使我的喜樂得以滿足。
PHIL|2|3|凡事不可自私自利，不可貪圖虛榮；只要心存謙卑，各人看別人比自己強。
PHIL|2|4|各人不要單顧自己的事，也要顧別人的事。
PHIL|2|5|你們當以基督耶穌的心為心：
PHIL|2|6|他本有上帝的形像， 卻不堅持自己與上帝同等 ；
PHIL|2|7|反倒虛己， 取了奴僕的形像， 成為人的樣式； 既有人的樣子，
PHIL|2|8|就謙卑自己， 存心順服，以至於死， 且死在十字架上。
PHIL|2|9|所以上帝把他升為至高， 又賜給他超乎萬名之上的名，
PHIL|2|10|使一切在天上的、地上的和地底下的， 因耶穌的名， 眾膝都要跪下，
PHIL|2|11|眾口都要宣認： 耶穌基督是主， 歸榮耀給父上帝。
PHIL|2|12|我親愛的，這樣看來，你們向來是順服的，不但我在你們那裏，就是我現在不在你們那裏的時候更是順服的，就當恐懼戰兢完成你們自己得救的事；
PHIL|2|13|因為是上帝在你們心裏運行，使你們又立志又實行，為要成就他的美意。
PHIL|2|14|你們無論做甚麼事，都不要發怨言起爭論，
PHIL|2|15|好使你們無可指責，誠實無偽，在這彎曲悖謬的世代作上帝無瑕疵的兒女。你們在這世代中要像明光照耀，
PHIL|2|16|將生命的道顯明出來，使我在基督的日子得以誇耀我沒有白跑，也沒有徒勞。
PHIL|2|17|我以你們的信心為供獻的祭物，我若被澆獻在其上也是喜樂，並且與你們眾人一同喜樂。
PHIL|2|18|你們也要照樣喜樂，並且與我一同喜樂。
PHIL|2|19|我靠主耶穌希望很快能差 提摩太 去見你們，好讓我知道你們的事而心裏得著安慰。
PHIL|2|20|因為我沒有別人與我同心，真正關懷你們的事。
PHIL|2|21|其他的人都求自己的事，並不求耶穌基督的事。
PHIL|2|22|但你們知道 提摩太 是經得起考驗的，他與我為了福音一同服侍，待我像兒子待父親一樣。
PHIL|2|23|所以，我一看出我的事怎樣了結，我希望立刻差他去，
PHIL|2|24|但我靠著主自信我不久也會去。
PHIL|2|25|然而，我想必須差 以巴弗提 到你們那裏去。他是我的弟兄、同工和戰友，是你們差遣來供應我需要的。
PHIL|2|26|他很想念 你們眾人，並且極其難過，因為你們聽見他病了。
PHIL|2|27|他真的生病了，幾乎要死。然而上帝憐憫他，不但憐憫他，也憐憫我，免得我憂上加憂。
PHIL|2|28|所以，我更要盡快送他回去，好讓你們再見到他而喜樂，我也可以減少憂愁。
PHIL|2|29|故此，你們要在主裏歡歡喜喜地接待他，而且要尊重這樣的人，
PHIL|2|30|因他為做基督的工作不顧性命，幾乎至死，為要補足你們供應我不夠的地方。
PHIL|3|1|末了，我的弟兄們，你們要靠主喜樂。我把這些話再寫給你們，對我並不困難，對你們卻是妥當的。
PHIL|3|2|應當防備犬類，防備作惡的，防備妄自行割的。
PHIL|3|3|因為真受割禮的，就是我們這藉著上帝的靈敬拜、以基督耶穌為誇耀、不依靠肉體的。
PHIL|3|4|其實，我也可以靠肉體；若是別人以為他可以依靠肉體，我更可以。
PHIL|3|5|我出生後第八天受割禮；我是 以色列 族、 便雅憫 支派的人，是 希伯來 人所生的 希伯來 人。就律法說，我是法利賽人；
PHIL|3|6|就熱心說，我是迫害教會的；就律法上的義說，我是無可指責的。
PHIL|3|7|只是我先前以為對我是有益的，我現在因基督的緣故而當作是有損的。
PHIL|3|8|不但如此，我已把萬事當作是有損的，因我以認識我主基督耶穌為至寶。我為他已經丟棄萬事，看作糞土，為要贏得基督，
PHIL|3|9|並且得以在他裏面，不是有自己因律法而得的義，而是有信基督的義 ，就是基於信，從上帝而來的義，
PHIL|3|10|使我認識基督，知道他復活的大能，並且知道和他一同受苦，效法他的死，
PHIL|3|11|或許我也得以從死人中復活。
PHIL|3|12|這不是說我已經得著了，已經完全了；而是竭力追求，或許可以得著基督耶穌 所要我得著的 。
PHIL|3|13|弟兄們，我不是以為自己已經得著了；我只有一件事，就是忘記背後，努力面前的，
PHIL|3|14|向著標竿直跑，要得上帝在基督耶穌裏從上面召我來得的獎賞。
PHIL|3|15|所以，我們中間凡是成熟的人，總要存這樣的心；若在甚麼事上存別樣的心，上帝也會把這些事指示你們。
PHIL|3|16|然而，我們達到甚麼地步，就當照這個地步行。
PHIL|3|17|弟兄們，你們要一同效法我，也當留意看那些效法我們榜樣的人。
PHIL|3|18|因為，我屢次告訴你們，現在又流淚告訴你們：許多人行事是基督十字架的仇敵。
PHIL|3|19|他們的結局就是滅亡。他們的神明是自己的肚腹；他們以自己的羞辱為光榮，專以地上的事為念。
PHIL|3|20|我們卻是天上的國民，並且等候救主，就是主耶穌基督從天上降臨。
PHIL|3|21|他要按著那能使萬有歸服自己的大能，把我們這卑賤的身體改變形狀，和他自己榮耀的身體相似。
PHIL|4|1|我所親愛、所想念的弟兄們，你們就是我的喜樂，我的冠冕。我親愛的，你們應當靠主站立得穩。
PHIL|4|2|我勸 友阿蝶 和 循都基 要在主裏同心。
PHIL|4|3|我也求你這真實同負一軛的，要幫助這兩個女人，因為她們在福音上曾與我、 革利免 和我其餘的同工一同勞苦，他們的名字都在生命冊上。
PHIL|4|4|你們要靠主常常喜樂。我再說，你們要喜樂。
PHIL|4|5|要讓眾人知道你們謙讓的心。主已經近了。
PHIL|4|6|應當一無掛慮，只要凡事藉著禱告、祈求和感謝，將你們所要的告訴上帝。
PHIL|4|7|上帝所賜那超越人所能了解的平安 ，必在基督耶穌裏，保守你們的心懷意念。
PHIL|4|8|末了，弟兄們，凡是真實的、凡是可敬的、凡是公義的、凡是清潔的、凡是可愛的、凡是有美名的，若有甚麼德行，若有甚麼稱讚，你們都要留意。
PHIL|4|9|你們從我所學習的，所領受的，所聽見的，所看見的事，你們都要繼續去做，賜平安的上帝就必與你們同在。
PHIL|4|10|我靠主大大喜樂，因為你們關懷我的心如今又表現了出來；其實你們一直都關懷我，只是沒有機會罷了。
PHIL|4|11|我並不是因缺乏而說這話，因為我已經學會無論在甚麼景況都可以知足。
PHIL|4|12|我知道怎樣處卑賤，也知道怎樣處豐富；或飽足或飢餓，或有餘或缺乏，任何事情，任何景況，我都得了祕訣。
PHIL|4|13|我靠著那加給我力量的，凡事都能做。
PHIL|4|14|然而，你們能和我分擔憂患是一件好事。
PHIL|4|15|腓立比 人哪，你們也知道我開始傳福音、離開 馬其頓 的時候，在收支的事上，除了你們以外，並沒有別的教會和我分擔。
PHIL|4|16|就是我在 帖撒羅尼迦 ，你們也一再差人來供給我的需用。
PHIL|4|17|我並不求甚麼饋贈，只求你們的果子不斷增多，歸在你們的賬上。
PHIL|4|18|但我已經如數收到，並且有餘；我已經充足，因我從 以巴弗提 受了你們的饋贈，當作極美的香氣，為上帝所接納、所喜悅的祭物。
PHIL|4|19|我的上帝必照他榮耀的豐富，在基督耶穌裏，使你們一切所需用的都充足。
PHIL|4|20|願榮耀歸給我們的父上帝，直到永永遠遠。阿們！
PHIL|4|21|請問候在基督耶穌裏的各位聖徒。跟我一起的眾弟兄都問候你們。
PHIL|4|22|眾聖徒都問候你們，特別在凱撒家裏的人問候你們。
PHIL|4|23|願主耶穌基督的恩與你們的靈同在！
COL|1|1|奉上帝旨意，作基督耶穌使徒的 保羅 ，和我們的弟兄 提摩太 ，
COL|1|2|寫信給 歌羅西 的聖徒，在基督裏忠心的弟兄。願恩惠、平安 從我們的父上帝歸給你們！
COL|1|3|我們為你們禱告的時候，常常感謝我們主耶穌基督的父上帝 ，
COL|1|4|因為聽見你們對基督耶穌的信心，並對眾聖徒有的愛心。
COL|1|5|這都是因著那給你們存在天上的盼望，它就是你們從前所聽見真理的道，就是福音；
COL|1|6|這福音傳到你們那裏，也傳到普天下，並且繼續增長，不斷結果，正如自從你們聽見福音，真正知道上帝恩惠的日子起，在你們中間也是這樣。
COL|1|7|這福音是你們從我們所親愛、一同作僕人的 以巴弗 學到的。他為我們 作了基督的忠心僕役，
COL|1|8|也把聖靈賜給你們的愛告訴我們。
COL|1|9|因此，我們自從聽見的日子就不住地為你們禱告和祈求，願你們滿有一切屬靈的智慧和悟性，真正知道上帝的旨意，
COL|1|10|好使你們行事為人對得起主，凡事蒙他喜悅，在一切善事上結果子，對上帝的認識更有長進。
COL|1|11|願你們從他榮耀的權能中，得以在一切事上力上加力，好使你們凡事歡歡喜喜地忍耐寬容，
COL|1|12|又感謝父，使你們配與眾聖徒在光明中分享基業。
COL|1|13|他救了我們脫離黑暗的權勢，遷移到他愛子的國度裏。
COL|1|14|藉著他的愛子，我們得蒙救贖，罪得赦免。
COL|1|15|愛子是那看不見的上帝之像， 是首生的 ，在一切被造的以先。
COL|1|16|因為萬有都是在他裏面 造的， 無論是天上的、地上的， 能看見的、不能看見的， 或是有權位的、統治的， 或是執政的、掌權的， 一概都是藉著他為著他造的。
COL|1|17|他在萬有之先； 萬有也靠他而存在。
COL|1|18|他是身體（教會）的頭； 他是元始， 是從死人中復活的首生者， 好讓他在萬有中居首位。
COL|1|19|因為上帝喜歡使一切的豐盛在他裏面居住，
COL|1|20|藉著他 ，上帝使萬有與自己和好， 無論是地上的、天上的， 都藉著他在十字架上所流的血促成了和平。
COL|1|21|從前你們與上帝隔絕，心思上與他為敵，行為邪惡；
COL|1|22|但如今，他藉著他兒子肉身的死，已經使你們與他自己和好了 ，把你們獻在他的面前，成為聖潔，沒有瑕疵，無可指責。
COL|1|23|只要你們持守信仰，根基穩固，堅定不移，不致動搖，離開了你們從前所聽見的福音的盼望；這福音也是傳給天下一切被造之物的，我— 保羅 作了這福音的僕役。
COL|1|24|現在我為你們受苦，倒很快樂；並且為基督的身體，就是為教會，我要在自己的肉身上補滿基督未盡的苦難。
COL|1|25|我照上帝為你們所賜我的職分作了教會的僕役，要把上帝的道傳得完滿；
COL|1|26|這道就是歷世歷代所隱藏的奧祕，但如今向他的聖徒顯明了。
COL|1|27|上帝要讓他們知道，這奧祕在外邦人中有何等豐盛的榮耀；就是基督在你們心裏 成了得榮耀的盼望。
COL|1|28|我們傳揚他，是用諸般的智慧，勸戒各人，教導各人，要把各人在基督裏完完全全地獻上 。
COL|1|29|我也為此勞苦，照著他在我裏面運用的大能盡心竭力。
COL|2|1|我要你們知道，我為你們和 老底嘉 人，和所有沒有與我見過面的人，是何等地勤奮；
COL|2|2|為要使他們的心得安慰，因愛心互相聯絡，以致有從確實了解所產生的豐盛，好深知上帝的奧祕，就是基督；
COL|2|3|在他裏面蘊藏著一切智慧和知識。
COL|2|4|我說這話，免得有人用花言巧語迷惑你們。
COL|2|5|雖然我身體不在你們那裏，心卻與你們同在，很高興見你們循規蹈矩，對基督的信心也堅固。
COL|2|6|既然你們接受了主基督耶穌，就要靠著他而生活，
COL|2|7|照著你們所領受的教導，在他裏面生根建造，信心堅固，充滿著感謝的心。
COL|2|8|你們要謹慎，免得有人用他的哲學和虛空的廢話，不照著基督，而是照人間的傳統和世上粗淺的學說 ，把你們擄去。
COL|2|9|因為上帝本性一切的豐盛都有形有體地居住在基督裏面；
COL|2|10|你們在他裏面也已經成為豐盛。他是所有執政掌權者的元首。
COL|2|11|你們也在他裏面受了不是人手所行的割禮，而是使你們脫去肉體情慾的基督的割禮。
COL|2|12|你們既受洗與他一同埋葬，也就在此禮上，因信那使他從死人中復活的上帝的作為跟他一同復活。
COL|2|13|你們從前在過犯和未受割禮的肉體中死了，上帝卻赦免了你們一切的過犯，使你們與基督一同活過來，
COL|2|14|塗去了在律例上所寫、敵對我們、束縛我們的字據，把它撤去，釘在十字架上。
COL|2|15|基督既將一切執政者、掌權者的權勢解除了，就在凱旋的行列中，將他們公開示眾，仗著十字架誇勝。
COL|2|16|所以，不要讓任何人在飲食上，或節期、初一、安息日等事上評斷你們。
COL|2|17|這些原是未來的事的影子，真體卻是屬基督的。
COL|2|18|不要讓人藉著故作謙虛和敬拜天使奪去你們的獎賞。這等人拘泥在所見過的幻象 ，隨著自己的慾望無故地自高自大，
COL|2|19|不緊隨元首；其實，由於他全身藉著關節筋絡才得到滋養，互相聯絡，靠上帝所賜的成長而成長。
COL|2|20|既然你們與基督同死而脫離了世上粗淺的學說，為甚麼仍像生活在世俗中一樣，去服從那「不可拿、不可嘗、不可摸」等類的規條呢？
COL|2|21|
COL|2|22|這些都是根據人的命令和教導，論到這一切都是一經使用就都敗壞了。
COL|2|23|這些規條使人徒有智慧之名，用私意崇拜，自表謙卑，苦待己身，其實在克制肉體的情慾上毫無功效。
COL|3|1|所以，既然你們已經與基督一同復活，就當求上面的事；那裏有基督，坐在上帝的右邊。
COL|3|2|你們要思考上面的事，不要思考地上的事。
COL|3|3|因為你們已經死了，你們的生命與基督一同藏在上帝裏面。
COL|3|4|基督是你們的生命，他顯現的時候，你們也要與他一同在榮耀裏顯現。
COL|3|5|所以，要治死你們在地上的肢體；就如淫亂、污穢、邪情、惡慾和貪婪—貪婪就是拜偶像。
COL|3|6|因這些事，上帝的憤怒必臨到那些悖逆的人 。
COL|3|7|當你們在這些事中活著的時候，你們的行為也曾是這樣的。
COL|3|8|但現在你們要棄絕這一切的事，就是惱恨、憤怒、惡毒、毀謗和口中污穢的言語。
COL|3|9|不要彼此說謊，因為你們已經脫去舊人和舊人的行為，
COL|3|10|穿上了新人，這新人照著造他的主的形像在知識上不斷地更新。
COL|3|11|在這事上並不分 希臘 人和 猶太 人，受割禮的和未受割禮的，未開化的人、 西古提 人、為奴的、自主的；惟獨基督是一切，又在一切之內。
COL|3|12|所以，你們既是上帝的選民，聖潔、蒙愛的人，要穿上憐憫、恩慈、謙虛、溫柔和忍耐。
COL|3|13|倘若這人與那人有嫌隙，總要彼此容忍，彼此饒恕；主 怎樣饒恕了你們，你們也要怎樣饒恕人。
COL|3|14|除此以外，還要穿上愛心，因為愛是貫通全德的。
COL|3|15|你們要讓基督所賜的和平在你們心裏作主，也為此蒙召，歸為一體。你們還要存感謝的心。
COL|3|16|當用各樣的智慧，把基督的道豐豐富富的存在心裏，用詩篇、讚美詩、靈歌，彼此教導，互相勸戒，以感恩的心歌頌上帝。
COL|3|17|你們無論做甚麼，或說話或行事，都要奉主耶穌的名，藉著他感謝父上帝。
COL|3|18|你們作妻子的，要順服自己的丈夫，這在主裏面是合宜的。
COL|3|19|你們作丈夫的，要愛你們的妻子，不可虐待她們。
COL|3|20|你們作兒女的，要凡事聽從父母，因為這是主所喜悅的。
COL|3|21|你們作父親的，不要惹兒女生氣，恐怕他們會灰心。
COL|3|22|你們作僕人的，要凡事聽從你們肉身的主人，不要只在眼前服事，像是討人喜歡的，總要心存誠實，因為你們敬畏主。
COL|3|23|你們無論做甚麼，都要從心裏做，像是為主做的，不是為人做的；
COL|3|24|因為你們知道，從主那裏必得著基業作為賞賜。你們要服侍的是主基督。
COL|3|25|行不義的人必受不義的報應；主並不偏待人。
COL|4|1|你們作主人的，待僕人要公正，因為知道，你們也有一位主在天上。
COL|4|2|你們要恆切禱告，在禱告中警醒感恩。
COL|4|3|同時，也要為我們禱告，求上帝給我們開傳道的門，能宣講基督的奧祕，
COL|4|4|使我能按著所該說的話將這奧祕顯明出來，我為此而被捆鎖。
COL|4|5|你們要把握時機，用智慧與外人來往。
COL|4|6|你們的言談要時常帶著溫和，好像用鹽調味，讓你們知道該怎樣應對每一個人。
COL|4|7|推基古 是我親愛的弟兄，忠心的僕役，和我一同作主的僕人；他要把我一切的事都告訴你們。
COL|4|8|我特意打發他到你們那裏去，好讓你們知道我們的情況，又讓他安慰你們的心。
COL|4|9|我又打發一位親愛忠心的弟兄 阿尼西謀 同去；他也是你們那裏的人。他們會把這裏一切的事都告訴你們。
COL|4|10|與我一同坐牢的 亞里達古 問候你們。 巴拿巴 的表弟 馬可 也問候你們。關於他，你們已經得到指示；他若到你們那裏，你們要接待他。
COL|4|11|稱為 猶士都 的 耶數 也問候你們。奉割禮的人中，只有這三個人是為上帝的國與我作同工的，也是使我心裏得安慰的。
COL|4|12|有一位你們那裏的人，作基督耶穌 僕人的 以巴弗 問候你們。他禱告的時候常為你們竭力祈求，願你們能站穩而成熟，充分確信上帝一切的旨意。
COL|4|13|他為你們、 老底嘉 和 希拉坡里 的弟兄多多勞苦，這是我可以為他作見證的。
COL|4|14|親愛的醫生 路加 和 底馬 問候你們。
COL|4|15|請問候 老底嘉 的弟兄以及 寧法 ，和她家裏 的教會。
COL|4|16|你們宣讀了這書信，也要交給 老底嘉 的教會宣讀；你們也要宣讀從 老底嘉 轉來的書信。
COL|4|17|你們要對 亞基布 說：「務要完成你從主所領受的職分。」
COL|4|18|我— 保羅 親筆問候你們。要記念我在捆鎖中。願恩惠與你們同在！
1THESS|1|1|保羅 、 西拉 、 提摩太 寫信給 帖撒羅尼迦 在父上帝和主耶穌基督裏的教會。願恩惠、平安 歸給你們！
1THESS|1|2|我們為你們眾人常常感謝上帝，禱告的時候提到你們，
1THESS|1|3|在我們的父上帝面前，不住地記念你們因信心所做的工作，因愛心所受的勞苦，因盼望我們主耶穌基督所存的堅忍。
1THESS|1|4|上帝所愛的弟兄啊，我知道你們是蒙揀選的；
1THESS|1|5|因為我們的福音傳到你們那裏，不僅在言語，也在能力，也在聖靈和充足的確信。你們知道，我們在你們那裏，為你們的緣故是怎樣為人。
1THESS|1|6|你們成為效法我們，更效法主的人，因聖靈所激發的喜樂，在大患難中領受了真道，
1THESS|1|7|從此你們作了 馬其頓 和 亞該亞 所有信主的人的榜樣。
1THESS|1|8|因為主的道已經從你們那裏傳播出去，你們向上帝的信心不只在 馬其頓 和 亞該亞 ，就是在各處也都傳開了，所以不用我們說甚麼話。
1THESS|1|9|因為他們自己已經傳講我們是怎樣進到你們那裏，你們是怎樣離棄偶像，歸向上帝來服侍那又真又活的上帝，
1THESS|1|10|等候他兒子從天降臨，就是上帝使他從死人中復活的那位救我們脫離將來憤怒的耶穌。
1THESS|2|1|弟兄們，你們自己知道我們來到你們那裏並不是徒然的。
1THESS|2|2|我們從前在 腓立比 蒙難受辱，這是你們知道的，可是我們還是靠著上帝給我們的勇氣，在強烈反對中把上帝的福音傳給你們。
1THESS|2|3|我們的勸勉不是出於錯誤，也不是出於污穢，也不是用詭詐。
1THESS|2|4|但上帝既然認定我們經得起考驗，把福音託付我們，我們就照著傳講，不是要討人喜歡，而是要討那考驗我們的心的上帝喜歡。
1THESS|2|5|因為我們從來沒有用過諂媚的話，這是你們知道的，也沒有藏著貪心，這是上帝可以作證的。
1THESS|2|6|我們作為基督的使徒，雖然可以受人尊重，卻沒有向你們或向別人求榮耀，反而在你們當中心存溫柔，如同母親哺乳自己的孩子。
1THESS|2|7|
1THESS|2|8|既然我們這樣愛你們，不但樂意將上帝的福音給你們，連自己的性命也樂意給你們，因為你們是我們所疼愛的。
1THESS|2|9|弟兄們，你們記念我們的辛苦勞碌，晝夜做工，傳上帝的福音給你們，免得你們任何人受累。
1THESS|2|10|我們對你們信主的人是何等聖潔、正直、無可指責，這有你們作證，也有上帝作證。
1THESS|2|11|正如你們知道，我們待你們好像父親待自己的兒女一樣。
1THESS|2|12|我們勸勉你們，安慰你們，囑咐你們，使你們行事對得起那召你們進他自己的國、得他榮耀的上帝。
1THESS|2|13|為此，我們也不斷地感謝上帝，因為你們聽見我們所傳上帝的道的時候，你們領受了，不以為這是人的道，而以為這確實是上帝的道，而且在你們信主的人當中運行著。
1THESS|2|14|弟兄們，你們與 猶太 地區上帝的各教會，就是在基督耶穌裏的各教會，有同樣的遭遇，因為你們也受了同胞的迫害，像他們受了 猶太 人的迫害一樣。
1THESS|2|15|這些 猶太 人不但殺了主耶穌和先知們，又把我們趕出去。他們令上帝不悅，且與眾人為敵，
1THESS|2|16|阻撓我們傳道給外邦人，使他們得救，以致常常惡貫滿盈，但上帝的憤怒終於臨到他們身上。
1THESS|2|17|弟兄們，我們被迫暫時與你們分離，身體離開，心卻沒有；我們極力想法子，渴望見你們的面。
1THESS|2|18|所以我們很想到你們那裏去。我－ 保羅 有一兩次要去，只是撒但阻擋了我們。
1THESS|2|19|當我們的主耶穌再來，我們站在他面前的時候，我們的盼望、喜樂和所誇的冠冕是甚麼呢？不正是你們嗎？
1THESS|2|20|你們就是我們的榮耀和喜樂！
1THESS|3|1|既然我們不能再忍，就決定獨自留在 雅典 ，
1THESS|3|2|於是差派我們在基督福音上作上帝同工的弟兄 提摩太 前去，在你們所信的道上堅固你們，勸勉你們，
1THESS|3|3|免得有人被這些患難動搖。因為你們自己知道，我們受患難原是命定的。
1THESS|3|4|我們在你們那裏的時候，曾預先告訴你們，我們必受患難；你們知道，這果然發生了。
1THESS|3|5|為此，既然我不能再忍，就差派人去，要知道你們的信心如何，恐怕那誘惑人的果真誘惑了你們，以致我們的勞苦歸於徒然。
1THESS|3|6|但是， 提摩太 剛從你們那裏回來，將你們信心和愛心的好消息報給我們，又說你們常常記念我們，切切想見我們，如同我們想見你們一樣。
1THESS|3|7|所以，弟兄們，我們在一切困苦患難中，因著你們的信心得到鼓勵。
1THESS|3|8|如今你們若靠主站立得穩，我們就得生了。
1THESS|3|9|我們在上帝面前，因著你們滿有喜樂。為這一切喜樂，我們能用怎樣的感謝為你們報答上帝呢？
1THESS|3|10|我們晝夜切切祈求要見你們的面，來補足你們信心的不足。
1THESS|3|11|願我們的父上帝自己和我們的主耶穌，為我們開路到你們那裏去。
1THESS|3|12|又願主使你們彼此相愛的心，和愛眾人的心，都能增長，充足，如同我們愛你們一樣，
1THESS|3|13|好堅固你們的心，使你們在我們的主耶穌同他眾聖徒來臨的時候，在我們父上帝面前，成為聖潔，無可指責。阿們！
1THESS|4|1|末了，弟兄們，我們靠著主耶穌求你們，勸你們，既然你們領受了我們的教導，知道該怎樣行事為人，討上帝的喜悅，其實你們也正這樣行，我勸你們要更加努力。
1THESS|4|2|你們原知道，我們憑主耶穌傳給你們甚麼命令。
1THESS|4|3|上帝的旨意就是要你們成為聖潔，遠避淫行；
1THESS|4|4|要你們各人知道怎樣用聖潔、尊貴控制自己的身體 ，
1THESS|4|5|不放縱私慾的邪情，像不認識上帝的外邦人。
1THESS|4|6|不准有人在這事上越軌，佔他弟兄的便宜；因為這一類的事，主必報應，正如我預先對你們說過，又切切警告過你們的。
1THESS|4|7|上帝召我們本不是要我們沾染污穢，而是要我們聖潔。
1THESS|4|8|所以，那棄絕這教導的不是棄絕人，而是棄絕那把自己的聖靈賜給你們的上帝。
1THESS|4|9|有關弟兄間的手足之情，不用人寫信給你們，因為你們自己蒙了上帝的教導要彼此相愛。
1THESS|4|10|你們向全 馬其頓 的眾弟兄固然是這樣行，但我勸弟兄們要更加努力。
1THESS|4|11|要立志過安靜的生活，管自己的事，親手 做工，正如我們從前吩咐你們的，
1THESS|4|12|好使你們的行為能得外人的尊敬，同時也不依賴任何人。
1THESS|4|13|弟兄們，至於已睡了的人，我們不願意你們不知道，恐怕你們憂傷，像那些沒有指望的人一樣。
1THESS|4|14|既然我們信耶穌死了，復活了，那些已經在耶穌裏睡了的人，上帝也必將他們與耶穌一同帶來。
1THESS|4|15|我們照主的話告訴你們一件事：我們這活著還存留到主來臨的人，絕不會在那已經睡了的人之先。
1THESS|4|16|因為，召集令一發，天使長的呼聲一叫，上帝的號角一吹，主必親自從天降臨；那在基督裏死了的人必先復活，
1THESS|4|17|然後我們這些活著還存留的人必和他們一同被提到雲裏，在空中與主相會。這樣，我們就要和主永遠同在。
1THESS|4|18|所以，你們當用這些話彼此勸勉。
1THESS|5|1|弟兄們，關於那時候和日期，不用人寫信給你們，
1THESS|5|2|因為你們自己明明知道，主的日子來到會像賊在夜間突然來到一樣。
1THESS|5|3|人正說平安穩定的時候，災禍忽然臨到他們，如同陣痛臨到懷胎的婦人一樣，他們絕逃脫不了。
1THESS|5|4|弟兄們，你們並不在黑暗裏，那日子不會像賊一樣臨到你們。
1THESS|5|5|你們都是光明之子，都是白晝之子；我們不屬黑夜，也不屬幽暗。
1THESS|5|6|所以，我們不要沉睡，像別人一樣，總要警醒謹慎。
1THESS|5|7|因為睡了的人是在夜間睡，醉了的人是在夜間醉。
1THESS|5|8|但既然我們屬於白晝，就應當謹慎，把信和愛當作護心鏡遮胸，把得救的盼望當作頭盔戴上。
1THESS|5|9|因為上帝不是預定我們受懲罰，而是預定我們藉著我們的主耶穌基督得救。
1THESS|5|10|他替我們死，讓我們無論醒著、睡著，都與他同活。
1THESS|5|11|所以，你們該彼此勸勉，互相造就，正如你們素常做的。
1THESS|5|12|弟兄們，我們勸你們要敬重那些在你們中間勞苦的，就是在主裏面督導你們、勸戒你們的人。
1THESS|5|13|又因他們所做的工作，要以愛心格外尊重他們。你們也要彼此和睦。
1THESS|5|14|弟兄們，我們勸你們，要警戒不守規矩的人，勉勵灰心的人，扶助軟弱的人，對眾人要有耐心。
1THESS|5|15|你們要謹慎，無論是誰都不要以惡報惡，彼此間和對眾人都要追求做好事。
1THESS|5|16|要常常喜樂，
1THESS|5|17|不住地禱告，
1THESS|5|18|凡事謝恩，因為這是上帝在基督耶穌裏向你們所定的旨意。
1THESS|5|19|不要熄滅聖靈；
1THESS|5|20|不要藐視先知的講論。
1THESS|5|21|但凡事要察驗：美善的事要持守，
1THESS|5|22|各樣惡事要禁戒。
1THESS|5|23|願賜平安 的上帝親自使你們完全成聖！願你們的靈、魂、體得蒙保守，在我們的主耶穌基督來臨的時候，完全無可指責。
1THESS|5|24|那召你們的本是信實的，他必成就這事。
1THESS|5|25|弟兄們，請也為 我們禱告。
1THESS|5|26|用聖潔的吻向眾弟兄問安。
1THESS|5|27|我指著主囑咐你們，要把這信宣讀給眾弟兄聽。
1THESS|5|28|願我們的主耶穌基督的恩惠與你們同在！
2THESS|1|1|保羅 、 西拉 和 提摩太 寫信給 帖撒羅尼迦 、在我們的父上帝與主耶穌基督裏的教會。
2THESS|1|2|願恩惠、平安 從我們的 父上帝和主耶穌基督歸給你們！
2THESS|1|3|弟兄們，我們該常常為你們感謝上帝，這本是合宜的；因為你們的信心格外增長，你們眾人彼此相愛的心也都增加。
2THESS|1|4|所以，我們在上帝的各教會裏為你們誇耀，因為你們在所受的一切壓迫患難中仍牢守著耐心和信心。
2THESS|1|5|這正是上帝公義判斷的明證，使你們配得上他的國，你們就是為這國受苦。
2THESS|1|6|既然上帝是公義的，他必以患難報復那加患難給你們的人，
2THESS|1|7|也必使你們這受患難的人與我們同得平安。那時，主耶穌同他有權能的天使從天上在火焰中顯現，要報應那些不認識上帝和不聽從我們的主耶穌福音的人。
2THESS|1|8|
2THESS|1|9|他們要受懲罰，永遠沉淪，與主的面和他權能的榮光隔絕。
2THESS|1|10|這正是主再來，要在他聖徒的身上得榮耀，就是要使一切信的人感到驚訝的那日子，因為你們信了我們對你們作的見證。
2THESS|1|11|為此，我們常為你們禱告，願我們的上帝看你們與他的呼召相配，又用大能成就你們一切良善的美意和因信心所做的工作，
2THESS|1|12|使我們主耶穌的名，照著我們的上帝和主耶穌基督的恩，在你們身上得榮耀，你們也在他身上得榮耀。
2THESS|2|1|弟兄們，關於我們主耶穌基督的來臨和我們到他那裏聚集，我勸你們：
2THESS|2|2|無論藉著靈，藉著言語，藉著冒我的名寫的書信，說主的日子已經到了，不要輕易動心，也不要驚慌。
2THESS|2|3|不要讓任何人用甚麼法子欺騙你們，因為那日子以前必有叛教的事，並有那不法的人，那沉淪之子出現。
2THESS|2|4|那抵擋者高抬自己超過一切稱為神明的，和一切受人敬拜的，甚至坐在上帝的殿裏，自稱為上帝。
2THESS|2|5|我還在你們那裏的時候曾把這些事告訴你們，你們不記得嗎？
2THESS|2|6|現在你們也知道那攔阻他的是甚麼，為要使他到了時機才出現。
2THESS|2|7|因為那不法的隱祕已經運作，只是現在有一個阻擋的，要等到那阻擋的被除去才會發作，
2THESS|2|8|那時這不法的人必出現，主耶穌 要用口中的氣滅絕他，以自己來臨的光輝摧毀他。
2THESS|2|9|這不法的人來，是靠撒但的運作，行各樣的異能、神蹟和一切虛假的奇事，
2THESS|2|10|並且在那沉淪的人身上行各樣不義的詭詐，因為他們不領受愛真理的心，好讓他們得救。
2THESS|2|11|故此，上帝就給他們一個引發錯誤的心，叫他們信從虛謊，
2THESS|2|12|使一切不信真理、倒喜愛不義的人都被定罪。
2THESS|2|13|主所愛的弟兄們哪，我們本該常為你們感謝上帝，因為他揀選你們為初熟的果子 ，使你們因信真道，又蒙聖靈感化成聖，得到拯救。
2THESS|2|14|為此，上帝藉著我們所傳的福音呼召你們，好得著我們主耶穌基督的榮光。
2THESS|2|15|所以，弟兄們，你們要站立得穩，凡所領受的教導，無論是我們口傳的，是信上寫的，都要堅守。
2THESS|2|16|願我們主耶穌基督自己，和那愛我們、開恩將永遠的安慰及美好的盼望賜給我們的父上帝，
2THESS|2|17|安慰你們的心，並且在一切善行善言上堅固你們！
2THESS|3|1|末了，弟兄們，請你們為我們禱告，好讓主的道快快傳開，得著榮耀，正如在你們中間一樣，
2THESS|3|2|也讓我們能脫離無理和邪惡人的手，因為不是人人都有信仰。
2THESS|3|3|但主是信實的，他要堅固你們，保護你們脫離那邪惡者。
2THESS|3|4|我們靠主對你們有信心，你們現在遵行，以後也必遵行我們所吩咐的。
2THESS|3|5|願主引導你們的心去愛上帝，並學基督的忍耐！
2THESS|3|6|弟兄們，我們奉主耶穌基督的名吩咐你們，凡有弟兄懶散，不遵守我們所傳授的教導，要遠離他。
2THESS|3|7|你們自己知道該怎樣效法我們。因為我們在你們當中從未懶散過，
2THESS|3|8|也從未白吃人的飯，倒是辛苦勞碌，晝夜做工，免得使你們中間有人受累。
2THESS|3|9|這並不是因我們沒有權柄，而是要給你們作榜樣，好讓你們效法我們。
2THESS|3|10|我們在你們那裏的時候曾吩咐你們，說若有人不肯做工，就不可吃飯。
2THESS|3|11|因為我們聽說，在你們中間有人懶散，甚麼工都不做，反倒專管閒事。
2THESS|3|12|我們靠主耶穌基督吩咐並勸戒這樣的人，要安分做工，自食其力。
2THESS|3|13|弟兄們，你們行善不可喪志。
2THESS|3|14|若有人不聽從我們這信上的話，要把他記下，不和他交往，使他自覺羞愧；
2THESS|3|15|但不要把他當仇人，要勸他如勸弟兄。
2THESS|3|16|願賜平安 的主隨時隨事親自賜給你們平安！願主與你們眾人同在！
2THESS|3|17|我— 保羅 親筆向你們問安。凡我的信都以此為記，我的筆跡就是這樣。
2THESS|3|18|願我們主耶穌基督的恩惠與你們眾人同在！
1TIM|1|1|奉我們的救主上帝，和我們的盼望基督耶穌的命令，作基督耶穌使徒的 保羅 ，
1TIM|1|2|寫信給那因信主作我真兒子的 提摩太 。願恩惠、憐憫、平安 從父上帝和我們主基督耶穌歸給你！
1TIM|1|3|我往 馬其頓 去的時候，曾勸你留在 以弗所 ，好囑咐某些人不可傳別的教義，
1TIM|1|4|也不要聽從無稽的傳說和冗長的家譜；這樣的事只會引起爭論，無助於上帝的計劃，這計劃是憑著信才能了解的。
1TIM|1|5|但命令的目的就是愛；這愛是出於清潔的心、無愧的良心和無偽的信心。
1TIM|1|6|有人偏離了這些而轉向空談，
1TIM|1|7|想要作律法教師，卻不明白自己所講的是甚麼，也不知道所主張的是甚麼。
1TIM|1|8|我們知道，只要人善用律法，律法是好的；
1TIM|1|9|因為知道律法不是為義人訂立的，而是為不法和叛逆的，不虔誠和犯罪的，不聖潔和戀世俗的，弒父母和殺人的，
1TIM|1|10|犯淫亂和親男色的，拐賣人口和說謊話的，並起假誓的，或是為任何違背健全教義的事訂立的。
1TIM|1|11|這是按照可稱頌、榮耀之上帝交託我的福音說的。
1TIM|1|12|我感謝那賜給我力量的我們的主基督耶穌，因為他認為我可信任，派我服事他。
1TIM|1|13|我從前是褻瀆、迫害、侮慢上帝的人；然而我還蒙了憐憫，因為我是在不信、不明白的時候做的。
1TIM|1|14|而且我們的主的恩典格外豐盛，使我在基督耶穌裏有信心和愛心。
1TIM|1|15|這話可信，值得完全接受：「基督耶穌到世上來是要拯救罪人」，而在罪人中我是個罪魁。
1TIM|1|16|然而，我蒙了憐憫，好讓基督耶穌在我這罪魁身上顯明他完全的忍耐，給後來信他得永生的人作榜樣。
1TIM|1|17|願尊貴、榮耀歸給永世的君王，那不朽壞、看不見、獨一的上帝，直到永永遠遠。阿們！
1TIM|1|18|我兒 提摩太 啊，我照從前指著你的預言把這命令交託你，使你能藉著這些預言打那美好的仗，
1TIM|1|19|常存信心和無愧的良心。有些人丟棄良心，在信仰上觸了礁；
1TIM|1|20|其中有 許米乃 和 亞歷山大 ，我已經把他們交給撒但，讓他們學會不再褻瀆。
1TIM|2|1|所以，我勸你，首先要為人人祈求、禱告、代求、感謝；
1TIM|2|2|為君王和一切在位的，也要如此，使我們能夠敬虔端正地過平穩寧靜的生活。
1TIM|2|3|這是好的，在我們的救主上帝面前可蒙悅納。
1TIM|2|4|他願意人人得救，並得以認識真理。
1TIM|2|5|因為只有一位上帝， 在上帝和人之間也只有一位中保， 是成為人的基督耶穌。
1TIM|2|6|他獻上自己作人人的贖價； 在適當的時候這事已經證實了。
1TIM|2|7|我為此奉派作傳道，作使徒，在信仰和真理上作外邦人的教師。我說的是真話，不是說謊。
1TIM|2|8|我希望男人舉起聖潔的手隨處禱告，不發怒，不爭論。
1TIM|2|9|我也希望女人以端正、克制和合乎體統的服裝打扮自己，不以編髮、金飾、珍珠和名貴衣裳來打扮。
1TIM|2|10|要有善行，這才與自稱為敬畏上帝的女人相稱。
1TIM|2|11|女人要事事順服地安靜學習。
1TIM|2|12|我不許女人教導，也不許她管轄男人，只要安靜。
1TIM|2|13|因為 亞當 先被造，然後才是 夏娃 ；
1TIM|2|14|亞當 並沒有受騙，而是女人受騙，陷在過犯裏。
1TIM|2|15|然而，女人若持守信心、愛心，又聖潔克制，就必藉著生產而得救。
1TIM|3|1|「若有人想望監督的職分，他是在羨慕一件好事」，這話是可信的。
1TIM|3|2|監督必須無可指責，只作一個婦人的丈夫，有節制、克己、端正，樂意接待外人，善於教導，
1TIM|3|3|不酗酒，不打人；要溫和，不好鬥，不貪財。
1TIM|3|4|要好好管理自己的家，使兒女順服，凡事莊重。
1TIM|3|5|人若不知道管理自己的家，怎能照管上帝的教會呢？
1TIM|3|6|剛信主的，不可作監督，恐怕他自高自大，落在魔鬼所受的懲罰裏。
1TIM|3|7|監督也必須在教外有好名聲，免得被人毀謗，落在魔鬼的羅網裏。
1TIM|3|8|同樣，執事也必須莊重，不一口兩舌，不好酒，不貪不義之財；
1TIM|3|9|要存清白的良心固守信仰的奧祕。
1TIM|3|10|這些人也要先受考驗，若沒有可責之處，才讓他們作執事。
1TIM|3|11|同樣，女執事 也必須莊重，不說閒話，有節制，凡事忠心。
1TIM|3|12|執事只作一個婦人的丈夫，要好好管兒女和自己的家。
1TIM|3|13|因為善於作執事的，為自己得到美好的地位，並且無懼地堅信在基督耶穌裏的信仰。
1TIM|3|14|我希望盡快到你那裏去，所以先把這些事寫給你；
1TIM|3|15|倘若我延誤了，你也可以知道在上帝的家中該怎樣做。這家就是永生上帝的教會，真理的柱石和根基。
1TIM|3|16|敬虔的奧祕是公認為偉大的： 上帝在肉身顯現， 被聖靈稱義， 被天使看見， 被傳於外邦， 被世人信服， 被接在榮耀裏。
1TIM|4|1|聖靈明說，在末後的時期必有人離棄信仰，去聽信那誘惑人的邪靈和鬼魔的教訓。
1TIM|4|2|這是出於撒謊者的假冒；這些人的良心如同被熱鐵烙了一般。
1TIM|4|3|他們禁止嫁娶，又禁戒食物—就是上帝所造、讓那信而明白真理的人存感謝的心領受的。
1TIM|4|4|上帝所造之物樣樣都是好的，若存感謝的心領受，沒有一樣是不可吃的，
1TIM|4|5|都因上帝的話和人的祈禱而成為聖潔了。
1TIM|4|6|你若把這些事提醒弟兄們，就是基督耶穌的好執事，在信仰的話語和你向來所服從的正確教義上得到了栽培。
1TIM|4|7|要棄絕那世俗的言語和老婦的無稽傳說。要在敬虔上操練自己：
1TIM|4|8|因操練身體有些益處；但敬虔在各方面都有益，它有現今和未來的生命的應許。
1TIM|4|9|這話可信，值得完全接受。
1TIM|4|10|我們勞苦，努力 正是為此，因為我們的指望在乎永生的上帝。他是人人的救主，更是信徒的救主。
1TIM|4|11|你要囑咐和教導這些事。
1TIM|4|12|不可叫人小看你年輕，總要在言語、行為、愛心、信心、清潔上，都作信徒的榜樣。
1TIM|4|13|要以宣讀聖經，勸勉，教導為念，直等到我來。
1TIM|4|14|不要忽略你所得的恩賜，就是從前藉著預言、在眾長老按手的時候賜給你的。
1TIM|4|15|這些事你要殷勤去做，並要在這些事上專心，讓眾人看出你的長進來。
1TIM|4|16|要謹慎自己和自己的教導，要在這些事上恆心，因為這樣做，既能救自己，又能救聽你的人。
1TIM|5|1|不可嚴責老年人，要勸他如同父親。要待年輕人如同弟兄，
1TIM|5|2|年老婦女如同母親。要清清潔潔地待年輕婦女如同姊妹。
1TIM|5|3|要尊敬真正守寡的婦人。
1TIM|5|4|寡婦若有兒女，或有孫兒女，要讓兒孫先在自己家中學習行孝，報答親恩，因為這在上帝面前是可蒙悅納的。
1TIM|5|5|獨居無靠的真寡婦只仰賴上帝，晝夜不住地祈求禱告。
1TIM|5|6|但好宴樂的寡婦活著也算是死了。
1TIM|5|7|這些事，你要囑咐她們，讓她們無可指責。
1TIM|5|8|若有人不照顧親屬，尤其是自己家裏的人，就是背棄信仰，還不如不信的人。
1TIM|5|9|寡婦登記，年齡必須在六十歲以上，只作一個丈夫的妻子，
1TIM|5|10|又有行善的名聲，就如養育兒女，收留外人，洗聖徒的腳，救濟遭難的人，竭力行各樣善事。
1TIM|5|11|至於年輕的寡婦，你要拒絕登記，因為她們情慾衝動、背棄基督的時候，就想嫁人，
1TIM|5|12|她們因廢棄了當初所許的願而被定罪。
1TIM|5|13|同時，她們又學了懶惰，習慣於挨家閒逛；不但懶惰，而且說長道短，好管閒事，說些不該說的話。
1TIM|5|14|所以，我希望年輕的寡婦嫁人，生養兒女，治理家務，不讓敵人有辱罵的把柄，
1TIM|5|15|因為已經有一些人轉去隨從撒但了。
1TIM|5|16|信主的婦女若有親戚是寡婦，要救濟她們，不可拖累教會，好使教會能救濟真正無助的寡婦。
1TIM|5|17|善於督導教會的長老，尤其是勤勞講道教導人的，應該得到加倍的敬奉。
1TIM|5|18|因為經上說：「牛在踹穀的時候，不可籠住牠的嘴」；又說：「工人得工資是應當的。」
1TIM|5|19|有控告長老的案件，非有兩三個證人就不要受理。
1TIM|5|20|繼續犯罪的人，要在眾人面前責備他，使其餘的人也有所懼怕。
1TIM|5|21|我在上帝、基督耶穌和蒙揀選的天使面前囑咐你要遵守這些話，不可存成見，做事也不可偏心。
1TIM|5|22|不可急於給人行按手禮；也不可在別人的罪上有份，要保守自己純潔。
1TIM|5|23|為了你的胃，又常患病，不要只喝水，要稍微喝點酒。
1TIM|5|24|有些人的罪是明顯的，已先受審判了；有些人的罪是隨後跟著來。
1TIM|5|25|同樣，善行也有明顯的，就是那不明顯的也不能隱藏。
1TIM|6|1|凡負軛作奴隸的，要認為自己的主人配受各樣的尊敬，免得上帝的名和教導被人褻瀆。
1TIM|6|2|奴隸若有信主的主人，不可因他是主內弟兄就輕看他們，更要越發服侍他們，因為得到服侍的益處的正是信徒，是蒙愛的人。 你要教導人和勸勉這些事。
1TIM|6|3|若有人傳別的教義，不符合我們主耶穌基督純正的話語與合乎敬虔的教導，
1TIM|6|4|他是自高自大，一無所知，專好爭辯，擅於舌戰，因而生出嫉妒、紛爭、毀謗、惡意猜疑，
1TIM|6|5|和心術不正與喪失真理的人不停地爭吵，以敬虔為得利的門路。
1TIM|6|6|其實，敬虔加上知足就是大利。
1TIM|6|7|因為我們沒有帶甚麼到世上來， 也不能帶甚麼去；
1TIM|6|8|只要有衣有食， 我們就該知足。
1TIM|6|9|但那些想要發財的人就陷在誘惑、羅網和許多無知有害的慾望中，使人沉淪，以致敗壞和滅亡。
1TIM|6|10|貪財是萬惡之根。有人因貪戀錢財而背離信仰，用許多愁苦把自己刺透了。
1TIM|6|11|但你這屬上帝的人哪，要逃避這些事；要追求公義、敬虔、信心、愛心、忍耐、溫柔。
1TIM|6|12|你要為信仰打那美好的仗；要持定永生，你為此被召，也已經在許多見證人面前作了那美好的見證。
1TIM|6|13|我在那賜生命給萬物的上帝面前，並在向 本丟．彼拉多 作過那美好見證的基督耶穌面前囑咐你 ：
1TIM|6|14|要守這命令，毫不玷污，無可指責，直到我們的主耶穌基督顯現。
1TIM|6|15|到了適當的時候都要顯明出來： 他是那可稱頌、獨一的權能者， 萬王之王， 萬主之主，
1TIM|6|16|就是那獨一不死、 住在人不能靠近的光裏， 是人未曾看見，也是不能看見的。 願尊貴和永遠的權能都歸給他。阿們！
1TIM|6|17|至於那些今世富足的人，你要囑咐他們不要自高，也不要倚賴靠不住的錢財；要倚靠那厚賜萬物給我們享受的上帝。
1TIM|6|18|又要囑咐他們行善，在好事上富足，甘心施捨，樂意分享，
1TIM|6|19|為自己積存財富，而為將來打美好的根基，好使他們能把握那真正的生命。
1TIM|6|20|提摩太 啊，要持守所給你的託付。要躲避世俗的空談和那假冒知識的矛盾言論。
1TIM|6|21|有人自稱有這知識而偏離了信仰。 願恩惠與你們同在！
2TIM|1|1|奉上帝旨意，按照基督耶穌裏所應許的生命，作基督耶穌使徒的 保羅 ，
2TIM|1|2|寫信給我親愛的兒子 提摩太 。願恩惠、憐憫、平安 從父上帝和我們的主基督耶穌歸給你！
2TIM|1|3|我感謝上帝，就是我接續祖先用純潔的良心所事奉的上帝，在祈禱中晝夜不停地想念你。
2TIM|1|4|我一想起你的眼淚，就急切想見你，好讓我滿心快樂。
2TIM|1|5|我記得你無偽的信心，這信心先存在你外祖母 羅以 和你母親 友妮基 的心裏，我深信也存在你的心裏。
2TIM|1|6|為這緣故，我提醒你要把上帝藉著我按手所給你的恩賜再如火挑旺起來。
2TIM|1|7|因為上帝賜給我們的不是膽怯的心，而是剛強、仁愛、自制的心。
2TIM|1|8|所以，不要以給我們的主作見證為恥，也不要以我這為主被囚的為恥；總要靠著上帝的大能，與我為福音同受苦難。
2TIM|1|9|上帝救了我們， 以聖召召我們， 不是按我們的行為， 而是按他的旨意和恩典； 這恩典是萬古之先 在基督耶穌裏賜給我們的，
2TIM|1|10|但如今 藉著我們的救主基督耶穌的顯現已經表明出來； 他把死廢去， 藉著福音，將不朽的生命彰顯出來。
2TIM|1|11|我為這福音奉派作傳道，作使徒，作教師。
2TIM|1|12|為這緣故，我也受這些苦難。然而，我不以為恥，因為我知道我所信的是誰，也深信他能保全他所交託我的 ，直到那日。
2TIM|1|13|你從我聽到那健全的言論，要用在基督耶穌裏的信心和愛心常常守著，作為規範。
2TIM|1|14|你要靠著那住在我們裏面的聖靈，牢牢守住所交託給你那美好的事。
2TIM|1|15|你知道，所有在 亞細亞 的人都離棄了我，其中有 腓吉路 和 黑摩其尼 。
2TIM|1|16|願主憐憫 阿尼色弗 一家的人，因為他屢次令我欣慰。他不以我的鐵鏈為恥，
2TIM|1|17|反而一到 羅馬 就急切尋找我，並且找到了。
2TIM|1|18|願主使他在那日能蒙主的憐憫。他在 以弗所 怎樣多服事我，你是清楚知道的。
2TIM|2|1|我兒啊，你要在基督耶穌的恩典上剛強起來。
2TIM|2|2|你在許多見證人面前聽見我所教導的，也要交託給那忠心而又能教導別人的人。
2TIM|2|3|你要和我同受苦難，作基督耶穌的精兵。
2TIM|2|4|凡當兵的，不讓世務纏身，好使那招他當兵的人喜悅。
2TIM|2|5|運動員在比賽的時候，不按規則就不能得冠冕。
2TIM|2|6|勤勞的農夫理當先得糧食。
2TIM|2|7|我所說的話，你要考慮，因為主必在凡事上給你聰明。
2TIM|2|8|要記得耶穌基督，他是 大衛 的後裔，從死人中復活；這就是我所傳的福音。
2TIM|2|9|我為這福音受苦難，甚至像犯人一樣被捆綁，然而上帝的話沒有被捆綁。
2TIM|2|10|所以，我為了選民事事忍耐，為使他們也能得到那在基督耶穌裏的救恩和永遠的榮耀。
2TIM|2|11|這話是可信的： 我們若與基督同死，也必與他同活；
2TIM|2|12|我們若忍耐到底，也必和他一同作王。 我們若不認他，他也必不認我們；
2TIM|2|13|我們縱然失信，他仍是可信的， 因為他不能否認自己。
2TIM|2|14|你要向眾人提醒這些事，在上帝 面前囑咐他們不可在言詞上爭辯；這是沒有益處的，只能傷害聽的人。
2TIM|2|15|你當竭力在上帝面前作一個經得起考驗、無愧的工人，按著正意講解真理的話。
2TIM|2|16|要遠避世俗的空談，因為這等空談會使人進到更不敬虔的地步。
2TIM|2|17|他們的話如同毒瘡越爛越大；其中有 許米乃 和 腓理徒 ，
2TIM|2|18|他們偏離了真理，說復活的事已過去，敗壞了好些人的信心。
2TIM|2|19|然而，上帝堅固的根基屹立不移；上面有這印記說：「主認得他自己的人」，又說：「凡稱呼主名的人總要離開不義。」
2TIM|2|20|大戶人家不但有金器銀器，也有木器瓦器；有作為貴重之用的，有作為卑賤之用的。
2TIM|2|21|人若自潔，脫離卑賤的事，必成為貴重的器皿，成為聖潔，合乎主用，預備行各樣的善事。
2TIM|2|22|你要逃避年輕人的私慾，同那以純潔的心求告主的人追求公義、信實、仁愛、和平。
2TIM|2|23|但要棄絕那愚拙無知的辯論，因為你知道這等事只會引起爭辯。
2TIM|2|24|主的僕人不可爭辯，只要溫和待人，善於教導，恆心忍耐，
2TIM|2|25|用溫柔勸導反對的人。也許上帝會給他們悔改的心能明白真理，
2TIM|2|26|讓他們這些已被魔鬼擄去順從他詭計的人能醒悟過來，脫離他的羅網。
2TIM|3|1|你該知道，末世必有艱難的日子來到。
2TIM|3|2|那時人會專愛自己，貪愛錢財，自誇，狂傲，毀謗，違背父母，忘恩負義，心不聖潔，
2TIM|3|3|沒有親情，抗拒和解，好說讒言，不能節制，性情兇暴，不愛良善，
2TIM|3|4|賣主賣友，任意妄為，自高自大，愛好宴樂，不愛上帝，
2TIM|3|5|有敬虔的外貌，卻背棄了敬虔的實質，這等人你要避開。
2TIM|3|6|他們當中有人潛入別人家裏，操縱無知的婦女；這些婦女被罪惡壓制，被各樣的私慾引誘，
2TIM|3|7|雖然常常學習，終久無法達到明白真理的地步。
2TIM|3|8|從前 雅尼 和 佯庇 怎樣反對 摩西 ，這等人也怎樣抵擋真理；他們的心地敗壞，信仰經不起考驗。
2TIM|3|9|然而，他們沒有進步，因為他們的愚昧必在眾人面前顯露出來，像那兩人一樣。
2TIM|3|10|但你已經追隨了我的教導、行為、志向、信心、寬容、愛心、忍耐，
2TIM|3|11|以及我在 安提阿 、 以哥念 、 路司得 所遭遇的迫害和苦難。我忍受了何等的迫害！但從這一切苦難中，主都把我救了出來。
2TIM|3|12|其實，凡立志在基督耶穌裏敬虔度日的，也都將受迫害。
2TIM|3|13|只是作惡的和騙人的將變本加厲，迷惑人也被人迷惑。
2TIM|3|14|至於你，你要持守所學習的和所確信的，因為你知道是跟誰學的，
2TIM|3|15|並且知道你從小明白聖經，這聖經能使你因在基督耶穌裏的信 有得救的智慧。
2TIM|3|16|聖經都是上帝所默示的 ，於教訓、督責、使人歸正、教導人學義都是有益的，
2TIM|3|17|叫屬上帝的人得以完全，預備行各樣的善事。
2TIM|4|1|我在上帝面前，並在將來審判活人死人的基督耶穌面前，憑著他的顯現和他的國度鄭重地勸戒你：
2TIM|4|2|務要傳道；無論得時不得時總要專心，並以百般的忍耐和各樣的教導責備人，警戒人，勸勉人。
2TIM|4|3|因為時候將到，那時人會厭煩健全的教導，耳朵發癢，就隨心所欲地增添好些教師，
2TIM|4|4|並且掩耳不聽真理，偏向無稽的傳說。
2TIM|4|5|至於你，凡事要謹慎，忍受苦難，做傳福音的工作，盡你的職分。
2TIM|4|6|至於我，我已經被澆獻，離世的時候到了。
2TIM|4|7|那美好的仗我已經打過了，當跑的路我已經跑盡了，該信的道我已經守住了。
2TIM|4|8|從此以後，有公義的冠冕為我存留，就是按著公義審判的主到了那日要賜給我的；不但賜給我，也賜給凡愛慕他顯現的人。
2TIM|4|9|你要趕緊到我這裏來。
2TIM|4|10|因為 底馬 貪愛現今的世界，已經離棄我，往 帖撒羅尼迦 去了； 革勒士 往 加拉太 去； 提多 往 撻馬太 去；
2TIM|4|11|只有 路加 在我這裏。你來的時候把 馬可 帶來，因為他在服事 上於我有益。
2TIM|4|12|我已經打發 推基古 往 以弗所 去。
2TIM|4|13|我在 特羅亞 留給 加布 的那件外衣，你來的時候要帶來，那些書也帶來，特別是那幾卷羊皮的書。
2TIM|4|14|銅匠 亞歷山大 多方害我；主必照他所行的報應他。
2TIM|4|15|你也要防備他，因為他極力抗拒我們的話。
2TIM|4|16|我初次上訴時，沒有人前來幫助，竟都離棄了我，但願這罪不歸在他們身上。
2TIM|4|17|惟有主站在我身邊，加給我力量，使我能把福音完整地傳開，讓所有的外邦人都聽見；我也從獅子口裏被救出來。
2TIM|4|18|主必救我脫離一切的兇惡，也必救我進他的天國。願榮耀歸給他，直到永永遠遠。阿們！
2TIM|4|19|請向 百基拉 、 亞居拉 和 阿尼色弗 一家的人問安。
2TIM|4|20|以拉都 在 哥林多 住下了。 特羅非摩 病了，我把他留在 米利都 。
2TIM|4|21|你要趕緊在冬天以前到我這裏來。 友布羅 、 布田 、 利奴 、 革老底亞 和眾弟兄都向你問安。
2TIM|4|22|願主與你的靈同在！願恩惠與你們同在！
TITUS|1|1|上帝的僕人、耶穌基督的使徒 保羅 ，為了使上帝的選民信從與認識合乎敬虔的真理—
TITUS|1|2|這真理是在盼望那無謊言的上帝在萬古之先所應許的永生，
TITUS|1|3|到了適當的時機，藉著傳揚福音，把他的道顯明了；這傳揚的責任是按著我們的救主上帝的命令交託給我的—
TITUS|1|4|我寫信給在共同的信仰上作我真兒子的 提多 。願恩惠、平安 從父上帝和我們的救主基督耶穌歸給你！
TITUS|1|5|我從前把你留在 克里特 ，是要你將那沒有辦完的事都辦妥，又照我所吩咐你的，在各城設立長老。
TITUS|1|6|若有無可指責的人，只作一個婦人的丈夫，兒女也是信主的，沒有人告他們放蕩，不受約束，就可以設立。
TITUS|1|7|監督既然是上帝的管家，必須無可指責、不自負、不暴躁、不酗酒、不好鬥、不貪財；
TITUS|1|8|卻要樂意接待外人、好善、克己、正直、聖潔、節制，
TITUS|1|9|堅守合乎教義的可靠之道，就能將健全的教導勸勉人，又能駁倒爭辯的人。
TITUS|1|10|因為也有許多人不受約束，說空話欺哄人，尤其是那些奉割禮的人。
TITUS|1|11|這些人的口必須堵住，因為他們貪不義之財，將不該教導的事教導人，敗壞人的全家。
TITUS|1|12|克里特 人中有一個本地的先知說：「 克里特 人常說謊話，是惡獸，貪吃懶做。」
TITUS|1|13|這個見證是真的。為這緣故，你要嚴厲地責備他們，使他們在信仰上健全。
TITUS|1|14|不要聽 猶太 人無稽的傳說和背棄真理之人的命令。
TITUS|1|15|在潔淨的人，凡物都潔淨；在污穢不信的人，甚麼都不潔淨，連心地和天良也都污穢了。
TITUS|1|16|他們宣稱認識上帝，卻在行為上否認他；他們是可憎惡的，是悖逆的，不配做任何好事。
TITUS|2|1|至於你，你所講的總要合乎那健全的教導。
TITUS|2|2|勸老年人要有節制、端正、克己，在信心、愛心、耐心上都要健全。
TITUS|2|3|又要勸年長的婦女在操守上恭正，不說讒言，不作酒的奴隸，用善道教導人，
TITUS|2|4|好指教年輕的婦女愛丈夫，愛兒女，
TITUS|2|5|克己，貞潔，理家，善良，順服自己的丈夫，免得上帝的道被毀謗。
TITUS|2|6|同樣，要勸年輕人凡事克己。
TITUS|2|7|你要顯出自己是好行為的榜樣，在教導上要正直、莊重，
TITUS|2|8|言語健全，無可指責，使那反對的人，因說不出我們有甚麼不好而自覺羞愧。
TITUS|2|9|要勸僕人順服自己的主人，凡事討他的喜悅，不可頂撞他，
TITUS|2|10|不可私竊財物；要凡事顯出完美的忠誠，好事事都能榮耀我們救主上帝的教導。
TITUS|2|11|因為，上帝救眾人的恩典已經顯明出來，
TITUS|2|12|訓練我們除去不敬虔的心和世俗的情慾，在今世過克己、正直、敬虔的生活，
TITUS|2|13|等候福樂的盼望，並等候至大的上帝和我們的救主 耶穌基督的榮耀顯現。
TITUS|2|14|他為我們的緣故捨己，為了要贖我們脫離一切罪惡，又潔淨我們作他自己的子民，熱心為善。
TITUS|2|15|這些事你要講明，要充分運用你的職權勸勉人，責備人。不要讓任何人輕看你。
TITUS|3|1|你要提醒眾人，叫他們順服執政的、掌權的，要服從，預備行各樣善事。
TITUS|3|2|不要毀謗，不要爭吵，要和氣，對眾人總要顯出溫柔。
TITUS|3|3|我們從前也是無知、悖逆、受迷惑，作各樣私慾和宴樂的奴隸，在惡毒、嫉妒中度日，是可恨的，而且彼此相恨。
TITUS|3|4|但到了我們救主上帝的恩慈和慈愛顯明的時候，
TITUS|3|5|他救了我們，並不是因我們自己所行的義，而是照他的憐憫，藉著重生的洗和聖靈的更新。
TITUS|3|6|聖靈就是上帝藉著我們的救主耶穌基督厚厚地澆灌在我們身上的，
TITUS|3|7|好讓我們因他的恩得稱為義，可以憑著永生的盼望成為後嗣 。
TITUS|3|8|這話是可信的。 我願你堅持這些事，使那些已信上帝的人留心行善 。這都是美好且對人有益的。
TITUS|3|9|要遠避愚拙的辯論、家譜、紛爭和因律法而起的爭辯，因為這都是虛妄無益的。
TITUS|3|10|分門結黨的人，警戒過一兩次後就要拒絕跟他來往；
TITUS|3|11|因為你知道這樣的人已經背道，常常犯罪，自己定自己的罪了。
TITUS|3|12|我打發 亞提馬 或 推基古 到你那裏去的時候，你要趕緊往 尼哥坡里 來見我，因為我已經決定在那裏過冬。
TITUS|3|13|你要趕緊給 西納 律師和 亞波羅 送行，讓他們沒有缺乏。
TITUS|3|14|我們的人也該學習行善，幫助有迫切需要的人，這樣才不會不結果子。
TITUS|3|15|跟我同在一起的人都向你問安。請代向在信仰上愛我們的人問安。願恩惠與你們眾人同在！
PHLM|1|1|為基督耶穌被囚的 保羅 ，同弟兄 提摩太 ，寫信給我們所親愛的同工 腓利門 、
PHLM|1|2|亞腓亞 姊妹，和我們的戰友 亞基布 ，以及在你家裏的教會。
PHLM|1|3|願恩惠、平安 從我們的父上帝和主耶穌基督歸給你們！
PHLM|1|4|我在禱告中記念你的時候，常為你感謝我的上帝，
PHLM|1|5|因聽說你對眾聖徒的愛心，和你對主耶穌的信心。
PHLM|1|6|願你與人分享信心的時候，能產生功效，讓人知道我們 所行的各樣善事都是為基督做的。
PHLM|1|7|弟兄啊，由於你的愛心，我得到極大的快樂和安慰，因為眾聖徒的心從你得到舒暢。
PHLM|1|8|雖然我靠著基督能放膽吩咐你做該做的事，
PHLM|1|9|可是像我這上了年紀的 保羅 ，現在又是為基督耶穌被囚的，寧可憑著愛心求你，
PHLM|1|10|就是為我在捆鎖中所生的兒子 阿尼西謀 求你。
PHLM|1|11|從前他與你沒有益處，但如今與你我都有益處。
PHLM|1|12|我現在打發他回到你那裏去，他是我心肝。
PHLM|1|13|我本來有意將他留下，在我為福音所受的捆鎖中替你伺候我。
PHLM|1|14|但不知道你的意見，我不願意這樣做，好使你的善行不是出於勉強，而是出於自願。
PHLM|1|15|他暫時離開你，也許是要讓你永遠得著他，
PHLM|1|16|不再是奴隸，而是高過奴隸，是親愛的弟兄；對我確實如此，何況對你呢！無論在肉身或在主裏更是如此。
PHLM|1|17|所以，你若以我為同伴，就接納他，如同接納我一樣。
PHLM|1|18|他若虧負你，或欠你甚麼，都算在我的賬上吧，
PHLM|1|19|我必償還。這是我— 保羅 親筆寫的。我並不用對你說，甚至你自己也虧欠我呢！
PHLM|1|20|弟兄啊，希望你使我在主裏因你得益處，讓我的心在基督裏得到舒暢。
PHLM|1|21|我寫信給你，深信你必順服，知道你所要做的，必過於我所說的。
PHLM|1|22|此外，還請給我預備住處，因為我盼望藉著你們的禱告，必蒙恩回到你們那裏去。
PHLM|1|23|為基督耶穌與我一同坐監的 以巴弗 問候你。
PHLM|1|24|我的同工 馬可 、 亞里達古 、 底馬 、 路加 也都問候你。
PHLM|1|25|願 主耶穌基督的恩與你們的靈同在。
HEB|1|1|古時候，上帝藉著眾先知多次多方向列祖說話，
HEB|1|2|末世，藉著他兒子向我們說話，又立他為承受萬有的，也藉著他創造宇宙。
HEB|1|3|他是上帝榮耀的光輝，是上帝本體的真像，常用他大能的命令托住萬有。他洗淨了人的罪，就坐在高天至大者的右邊。
HEB|1|4|他所承受的名比天使的名更尊貴，所以他遠比天使崇高。
HEB|1|5|上帝曾對哪一個天使說過： 「你是我的兒子； 我今日生了你」？ 又說過： 「我要作他的父； 他要作我的子」呢？
HEB|1|6|再者，上帝引領他長子 進入世界的時候，說： 「上帝的使者都要拜他。」
HEB|1|7|關於使者，他說： 「上帝以風為使者， 以火焰為僕役。」
HEB|1|8|關於子，他卻說： 「上帝啊，你的寶座是永永遠遠的； 你國度的權杖是正直的權杖。
HEB|1|9|你喜愛公義，恨惡罪惡； 所以上帝，就是你的上帝，用喜樂油膏你， 勝過膏你的同伴。」
HEB|1|10|他又說： 「主啊，你起初立了地的根基， 天也是你手所造的。
HEB|1|11|天地都會消滅，你卻長存； 天地都會像衣服漸漸舊了；
HEB|1|12|你要將天地捲起來，像捲一件外衣， 天地像衣服都會改變。 你卻永不改變； 你的年數沒有窮盡。」
HEB|1|13|上帝曾對哪一個天使說： 「你坐在我的右邊， 等我使你的仇敵作你的腳凳」？
HEB|1|14|眾天使不都是事奉的靈，奉差遣為那將要承受救恩的人服務的嗎？
HEB|2|1|所以，我們必須越發注意所聽見的道，免得我們隨流失去。
HEB|2|2|既然那藉著天使所傳的話是確定的，凡違背不聽從的，都受了該受的報應；
HEB|2|3|我們若忽略這麼大的救恩，怎能逃避呢？這拯救起先是主親自講的，後來是聽見的人給我們證實了。
HEB|2|4|上帝又按自己的旨意，更用神蹟奇事、百般的異能，和聖靈所給的恩賜，與他們一同作見證。
HEB|2|5|我們所說將來的世界，上帝沒有交給天使管轄。
HEB|2|6|但有人在某處證明說： 「人算甚麼，你竟顧念他； 世人算甚麼，你竟眷顧他。
HEB|2|7|你使他暫時比天使微小 ， 賜他榮耀尊貴為冠冕， 你派他管理你手所造的，
HEB|2|8|使萬物都服在他的腳下。」 既然使萬物都服他 ，就沒有剩下一樣不服他的了。只是如今我們還不見萬物都服他；
HEB|2|9|惟獨見那成為暫時比天使微小的耶穌，因為受了死的痛苦，得了尊貴榮耀為冠冕，好使他因著上帝的恩，為人人經歷了死亡。
HEB|2|10|原來那為萬物所屬、為萬物所本的，為要領許多兒子進入榮耀，使救他們的元帥因受苦難而得以完全，本是合宜的。
HEB|2|11|因那使人成聖的，和那些得以成聖的，都是出於一。為這緣故，他稱他們為弟兄也不以為恥，
HEB|2|12|說： 「我要將你的名傳給我的弟兄， 在會眾中我要頌揚你。」
HEB|2|13|他又說： 「我要依賴他。」 他又說： 「看哪！我與上帝所給我的兒女都在這裏。」
HEB|2|14|既然兒女同有血肉之軀，他也照樣親自成了血肉之軀，為能藉著死敗壞那掌管死權的，就是魔鬼，
HEB|2|15|並要釋放那些一生因怕死而作奴隸的人。
HEB|2|16|誠然，他並沒有幫助天使，而是幫助了 亞伯拉罕 的後裔。
HEB|2|17|所以，他凡事應當與他的弟兄相同，為要在上帝的事上成為慈悲忠信的大祭司，為百姓的罪獻上贖罪祭。
HEB|2|18|既然他自己被試探而受苦，他能幫助被試探的人。
HEB|3|1|同蒙天召的聖潔弟兄啊，要思想我們所宣認為使者、為大祭司的耶穌；
HEB|3|2|他向指派他的盡忠，如同 摩西 向上帝的全 家盡忠一樣。
HEB|3|3|他比 摩西 配得更多的榮耀，好像建造房屋的人比房屋更尊榮；
HEB|3|4|因為房屋都必有人建造，但建造萬物的是上帝。
HEB|3|5|摩西 作為僕人，向上帝的全家盡忠，為將來要談論的事作證；
HEB|3|6|但是基督作為兒子，治理上帝的家。我們若堅持因盼望而有的膽量和誇耀，我們就是他的家了。
HEB|3|7|所以，正如聖靈所說： 「今日，你們若聽他的話，
HEB|3|8|就不可硬著心，像在背叛之時， 就如在曠野受試探之日。
HEB|3|9|在那裏，你們的祖宗試探我， 並且觀看我的作為，
HEB|3|10|有四十年之久。 所以，我厭煩那世代， 說：他們的心常常迷糊， 竟不知道我的道路！
HEB|3|11|我在怒中起誓： 他們斷不可進入我的安息！」
HEB|3|12|弟兄們，你們要謹慎，免得你們中間有人存著邪惡不信的心，離棄了永生的上帝。
HEB|3|13|總要趁著還有今日，天天彼此相勸，免得你們中間有人被罪迷惑，心腸剛硬了。
HEB|3|14|只要我們將起初確實的信心堅持到底，就在基督裏有份了。
HEB|3|15|經上說： 「今日，你們若聽他的話， 就不可硬著心，像在背叛之時。」
HEB|3|16|聽見他而又背叛他的是誰呢？豈不是跟著 摩西 從 埃及 出來的眾人嗎？
HEB|3|17|上帝向誰發怒四十年之久呢？豈不是那些犯罪而陳屍在曠野的人嗎？
HEB|3|18|他向誰起誓，不容他們進入他的安息呢？豈不是向那些不信從的人嗎？
HEB|3|19|這樣看來，他們不能進入安息是因為不信的緣故了。
HEB|4|1|所以，既然進入他安息的應許依舊存在，我們就該存畏懼的心，免得我們 中間有人似乎沒有得到安息。
HEB|4|2|因為的確有福音傳給我們像傳給他們一樣；只是所聽見的道對他們無益，因為他們沒有以信心與所聽見的道配合。
HEB|4|3|但我們已經信的人進入安息，正如上帝所說： 「我在怒中起誓： 他們斷不可進入我的安息！」 其實造物之工，從創世以來已經完成了。
HEB|4|4|論到第七日，有一處說：「到第七日，上帝就歇了他一切工作。」
HEB|4|5|又有一處說：「他們斷不可進入我的安息！」
HEB|4|6|既有這安息保留著讓一些人進入，那些先前聽見福音的人，因不信從而不得進去，
HEB|4|7|所以上帝多年後藉著 大衛 的書，又定了一天—「今日」，如以上所引的說： 「今日，你們若聽他的話， 就不可硬著心。」
HEB|4|8|若是 約書亞 已使他們享了安息，後來上帝就不會再提別的日子了。
HEB|4|9|這樣看來，另有一安息日的安息為上帝的子民保留著。
HEB|4|10|因為那些進入安息的，也是歇了自己的工作，正如上帝歇了他的工作一樣。
HEB|4|11|所以，我們務必竭力進入那安息，免得有人學了不順從而跌倒了。
HEB|4|12|上帝的道是活潑的，是有功效的，比一切兩刃的劍更鋒利，甚至魂與靈、骨節與骨髓，都能刺入、剖開，連心中的思念和主意都能辨明。
HEB|4|13|被造的，沒有一樣在他面前不是顯露的；萬物在他眼前都是赤露敞開的，我們必須向他交賬。
HEB|4|14|既然我們有一位偉大、進入高天的大祭司，就是耶穌—上帝的兒子，我們應當持定所宣認的道。
HEB|4|15|因為我們的大祭司並非不能體恤我們的軟弱；他也在各方面受過試探，與我們一樣，只是他沒有犯罪。
HEB|4|16|所以，我們只管坦然無懼地來到施恩的寶座前，為要得憐憫，蒙恩惠，作及時的幫助。
HEB|5|1|凡從人間挑選的大祭司都是奉派替人辦理屬上帝的事，要為罪獻上禮物和祭物 。
HEB|5|2|他能體諒無知和迷失的人，因為他自己也是被軟弱所困，
HEB|5|3|因此他理當為百姓和自己的罪獻祭。
HEB|5|4|沒有人可擅自取得大祭司的尊榮，惟有蒙上帝所選召的才可以，像 亞倫 一樣。
HEB|5|5|同樣，基督也沒有自取作大祭司的榮耀，而是在乎向他說話的那一位，他說： 「你是我的兒子， 我今日生了你。」
HEB|5|6|就如又有一處說： 「你是照著 麥基洗德 的體系 永遠為祭司。」
HEB|5|7|基督在他肉身的日子，曾大聲哀哭，流淚禱告，懇求那能救他免死的上帝，就因他的虔誠蒙了應允。
HEB|5|8|他雖然為兒子，還是因所受的苦難學了順從。
HEB|5|9|既然他得以完全，就為凡順從他的人成了永遠得救的根源，
HEB|5|10|並蒙上帝照著 麥基洗德 的體系宣稱他為大祭司。
HEB|5|11|論到這事，我們有好些話要說，可是很難解釋，因為你們聽不進去。
HEB|5|12|按時間說，你們早該作教師了，誰知還需要有人再將上帝聖言基礎的要道教導你們；你們成了那需要吃奶、不能吃乾糧的人。
HEB|5|13|凡只能吃奶的，就不熟練仁義的道理，因為他是嬰孩。
HEB|5|14|惟獨長大成人的才能吃乾糧，他們的心竅因練習而靈活，能分辨善惡了。
HEB|6|1|所以，我們應當離開基督道理的基礎，竭力進到成熟的地步；不必再立根基，就如懊悔致死的行為、信靠上帝、
HEB|6|2|各樣洗禮、按手禮、死人復活，以及永遠的審判等的教導。
HEB|6|3|上帝若准許，我們就這樣做。
HEB|6|4|論到那些已經蒙了光照、嘗過天恩的滋味、又於聖靈有份、並嘗過上帝的話的美味，和來世權能的人，若再離棄真道，就不可能使他們重新懊悔了；因為他們親自把上帝的兒子重釘十字架，公然羞辱他。
HEB|6|5|
HEB|6|6|
HEB|6|7|就如一塊田地吸收過屢次下的雨水，生長蔬菜，合乎耕種的人用，就從上帝得福。
HEB|6|8|這塊田地若長荊棘和蒺藜，必被廢棄，近於詛咒，結局就是焚燒。
HEB|6|9|親愛的，雖然這樣說，我們仍深信你們有更好的情況，更接近救恩。
HEB|6|10|因為上帝並非不公義，竟忘記你們的工作和你們為他的名所顯的愛心，就是你們過去和現在伺候聖徒的愛心。
HEB|6|11|我們盼望你們各人都顯出同樣的熱忱，一直到底，好達成所確信的指望。
HEB|6|12|這樣你們才不會懶惰，卻成為效法那些藉著信和忍耐承受應許的人。
HEB|6|13|當初上帝應許 亞伯拉罕 的時候，因為沒有比自己更大的可以指著起誓，就指著自己起誓，
HEB|6|14|說：「我必多多賜福給你；我必使你大大增多。」
HEB|6|15|這樣， 亞伯拉罕 因恆心等待而得了所應許的。
HEB|6|16|人都是指著比自己大的起誓，並且以起誓作保證，了結各樣的爭論。
HEB|6|17|照樣，上帝願意為那承受應許的人更有力地顯明他的旨意不可更改，他以起誓作保證。
HEB|6|18|藉這兩件不可更改的事—在這些事上，上帝絕不會說謊—我們這些逃往避難所的人能得到強有力的鼓勵，去抓住那擺在我們前頭的指望。
HEB|6|19|我們有這指望，如同靈魂的錨，又堅固又牢靠，進入幔子後面的至聖所。
HEB|6|20|為我們作先鋒的耶穌，既照著 麥基洗德 的體系成了永遠的大祭司，已經進入了。
HEB|7|1|這 麥基洗德 就是 撒冷 王，是至高上帝的祭司。他在 亞伯拉罕 打敗諸王回來的時候迎接他，並給他祝福。
HEB|7|2|亞伯拉罕 也將自己所得來的一切，取十分之一給他。他頭一個名字翻譯出來是「公義的王」，他又名「 撒冷 王」，是和平王的意思。
HEB|7|3|他無父、無母、無族譜、無生之始、無命之終，是與上帝的兒子相似，他永遠作祭司。
HEB|7|4|你們想一想，這個人多麼偉大啊！連先祖 亞伯拉罕 都拿戰利品的十分之一給他。
HEB|7|5|那得祭司職分的 利未 子孫，奉命照例向百姓取十分之一，這百姓是自己的弟兄，雖是從 亞伯拉罕 親身生的，還是照例取十分之一。
HEB|7|6|惟獨 麥基洗德 那不與他們同族譜的，從 亞伯拉罕 收取了十分之一，並且給蒙應許的 亞伯拉罕 祝福。
HEB|7|7|向來位分大的給位分小的祝福，這是無可爭議的。
HEB|7|8|在這事上，一方面，收取十分之一的都是必死的人；另一方面，收取十分之一的卻是那位被證實是活著的。
HEB|7|9|我們可以說，那接受十分之一的 利未 也是藉著 亞伯拉罕 納了十分之一，
HEB|7|10|因為 麥基洗德 迎接 亞伯拉罕 的時候， 利未 還在他先祖的身體裏面。
HEB|7|11|那麼，如果百姓藉著 利未 人的祭司職任能達到完全—因為百姓是在這職分下領受律法的—為甚麼還需要按照 麥基洗德 的體系另外興起一位祭司，而不按照 亞倫 的體系呢？
HEB|7|12|既然祭司的職分已更改，律法也需要更改。
HEB|7|13|因為這些話所指的人本屬別的支派，那支派裏從來沒有一人在祭壇前事奉的。
HEB|7|14|很明顯地，我們的主是從 猶大 出來的；但關於這支派， 摩西 並沒有提到祭司。
HEB|7|15|倘若有另一位像 麥基洗德 的祭司興起來，我的話就更顯而易見了。
HEB|7|16|他成為祭司，並不是照屬肉身的條例，而是照無窮 生命的大能。
HEB|7|17|因為有給他作見證的說： 「你是照著 麥基洗德 的體系 永遠為祭司。」
HEB|7|18|一方面，先前的誡命因軟弱無能而廢掉了，
HEB|7|19|（律法本來就不能成就甚麼）；另一方面，一個更好的指望被引進來，靠這指望，我們就可以親近上帝。
HEB|7|20|再者，耶穌成為祭司，並不是沒有上帝的誓言；其他的祭司被指派時並沒有這種誓言，
HEB|7|21|只有耶穌是起誓立的，因為那位立他的對他說： 「主起了誓， 絕不改變。 你是永遠為祭司。」
HEB|7|22|既是起誓立的，耶穌也作了更美之約的中保。
HEB|7|23|一方面，那些成為祭司的數目本來多，是因為受死亡限制不能長久留住。
HEB|7|24|另一方面，這位既是永遠留住的，他具有不可更換的祭司職任。
HEB|7|25|所以，凡靠著他進到上帝面前的人，他都能拯救到底，因為他長遠活著為他們祈求。
HEB|7|26|這樣一位聖潔、無邪惡、無玷污、遠離罪人、高過諸天的大祭司，對我們是最合適的；
HEB|7|27|他不像那些大祭司，每日必須先為自己的罪，後為百姓的罪獻祭，因為他只一次將自己獻上就把這事成全了。
HEB|7|28|律法所立的大祭司本是有弱點的人，但在律法以後，上帝以起誓的話立了兒子為大祭司，成為完全，直到永遠。
HEB|8|1|我們所講的事，其中第一要緊的就是：我們有這樣一位大祭司，他已經坐在天上至大者寶座的右邊，
HEB|8|2|在聖所，就是在真帳幕裏作僕役；這帳幕是主所支搭的，不是人所支搭的。
HEB|8|3|凡大祭司都是為獻禮物和祭物設立的，所以這位大祭司也必須有所獻上。
HEB|8|4|他若在地上，就不用作祭司，因為已經有照律法獻禮物的祭司了。
HEB|8|5|他們所供奉的本是天上之事的樣式和影像，正如 摩西 將要造帳幕的時候，上帝警戒他，說：「要謹慎，一切都要照著在山上指示你的樣式去做。」
HEB|8|6|如今耶穌已經得了更優越的事奉，正如他作更美之約的中保；這約原是憑更美之應許立的。
HEB|8|7|第一個約若沒有瑕疵，就無須尋求第二個約了。
HEB|8|8|所以上帝指責他們說： 「主說，看哪，日子將到， 我要與 以色列 家 和 猶大 家另立新的約；
HEB|8|9|不像我拉著他們祖宗的手 領他們出 埃及 地的時候， 與他們所立的約； 因為他們不恆心守我的約， 所以我也不理他們；這是主說的。
HEB|8|10|主又說： 那些日子以後， 我與 以色列 家所立的約是這樣： 我要將我的律法放在他們的心思裏， 寫在他們的心上； 我要作他們的上帝， 他們要作我的子民。
HEB|8|11|他們各人不用教導自己的鄉親和自己的弟兄，說：你要認識主； 因為從最小的到最大的， 他們都要認識我。
HEB|8|12|我要寬恕他們的不義， 絕不再記得他們的罪惡。」
HEB|8|13|既然上帝提到「新的約」，那麼第一個約就成為舊的了；而那漸舊漸衰的必然很快消逝了。
HEB|9|1|原來連第一個約都有敬拜的禮儀和屬世界的聖幕。
HEB|9|2|因為那預備好了的帳幕，第一層叫聖所，裏面有燈臺、供桌和供餅。
HEB|9|3|第二層幔子後又有一層帳幕，叫至聖所，
HEB|9|4|有金香壇和四周包金的約櫃，櫃裏有盛嗎哪的金罐、 亞倫 那根發過芽的杖和兩塊約版；
HEB|9|5|櫃上面有榮耀的基路伯罩著施恩座。有關這一切我現在不能一一細說。
HEB|9|6|這些物件既如此預備齊了，眾祭司就不斷地進第一層帳幕行拜上帝的禮。
HEB|9|7|至於第二層帳幕，惟有大祭司一年一次獨自進去，沒有一次不帶著血，為自己獻上，也為百姓無意所犯的過錯獻上。
HEB|9|8|聖靈藉此指明，第一層帳幕仍存在的時候，進入至聖所的路還沒有顯示。
HEB|9|9|那第一層帳幕是現今時代的一個預表，表示所獻的禮物和祭物都不能使敬拜的人在良心上得以完全。
HEB|9|10|這些事只不過是有關飲食和各種潔淨的規矩，是屬肉體的條例，它的功效是直到新次序的時期來到為止。
HEB|9|11|但現在基督已經來到，作了已實現的美事的大祭司，經過那更大更全備的帳幕，不是人手所造，也不是屬於這世界的；
HEB|9|12|他不用山羊和牛犢的血，而是用自己的血，只一次進入至聖所就獲得了永遠的贖罪。
HEB|9|13|若山羊和公牛的血，以及母牛犢的灰，灑在不潔的人身上，尚且使人成聖，身體潔淨，
HEB|9|14|何況基督的血，他藉著永遠的靈把自己無瑕疵地獻給上帝，更能洗淨我們 的良心，除去致死的行為，好事奉那位永生的上帝。
HEB|9|15|為此，基督作了新約的中保；因為他的死，贖了人在第一個約之時所犯的罪過，使蒙召的人能得著所應許永遠的產業。
HEB|9|16|凡有遺囑，必須證實立遺囑的人已經死了。
HEB|9|17|因為人死了，遺囑才有效力；立遺囑的人尚在，遺囑就不能生效。
HEB|9|18|所以，第一個約也是用血立的。
HEB|9|19|因為 摩西 當日照著律法將各樣誡命傳給眾百姓，就拿朱紅色絨和牛膝草，把牛犢、山羊 的血和水灑在書上，又灑在眾百姓身上，
HEB|9|20|說：「這血就是上帝與你們立約的憑據。」
HEB|9|21|他又照樣把血灑在帳幕和敬拜用的各樣器皿上。
HEB|9|22|按著律法，幾乎每樣東西都是用血潔淨的；沒有流血，就沒有赦罪。
HEB|9|23|這樣，照著天上樣式做的物件必須用這些禮儀去潔淨，但那天上的一切，自然當用更美的祭物去潔淨。
HEB|9|24|因為基督並沒有進了人手所造的聖所—這不過是真聖所的影像—而是進到天上，如今為我們出現在上帝面前。
HEB|9|25|他也無須多次將自己獻上，像大祭司每年帶著牛羊的血進入至聖所。
HEB|9|26|如果這樣，他從創世以來就必須多次受苦了。但如今，他在今世的末期顯現，僅一次把自己獻為祭，好除掉罪。
HEB|9|27|按著命定，人人都有一死，死後且有審判。
HEB|9|28|同樣，基督既然一次獻上，擔當了許多人的罪，將來要第二次顯現，與罪無關，而是為了拯救熱切等候他的人。
HEB|10|1|既然律法只不過是未來美好事物的影子，不是本體的真像，就不能藉著每年常獻一樣的祭物，使那些進前來的人完全。
HEB|10|2|若不然，獻祭的事豈不早已停止了嗎？因為敬拜的人僅只一次潔淨，良心就不再覺得有罪了。
HEB|10|3|但是這些祭物使人每年都想起罪來，
HEB|10|4|因為公牛和山羊的血不能除罪。
HEB|10|5|所以，基督到世上來的時候，就說： 「祭物和禮物不是你所要的， 但你曾給我預備了身體。
HEB|10|6|燔祭和贖罪祭 是你不喜歡的。
HEB|10|7|那時我說： 看哪！我來了，我的事在經卷上已經記載了； 上帝啊！我來為要照你的旨意行。」
HEB|10|8|以上說：「祭物和禮物，以及燔祭和贖罪祭，不是你所要的，也不是你喜歡的。」這都是按著律法獻的。
HEB|10|9|他接著說：「看哪！我來了，為要照你的旨意行。」可見他除去在先的，為要立定在後的。
HEB|10|10|我們憑著這旨意，藉著耶穌基督，僅只一次獻上他的身體就得以成聖。
HEB|10|11|所有的祭司天天站著事奉上帝，屢次獻上一樣的祭物，這祭物永不能除罪。
HEB|10|12|但基督獻了一次永遠有效的贖罪祭，就坐在上帝的右邊，
HEB|10|13|從此等候他的仇敵成為他的腳凳。
HEB|10|14|因為他僅只一次獻祭，就使那些得以成聖的人永遠完全。
HEB|10|15|聖靈也對我們作證，因為他說過：
HEB|10|16|「主說：那些日子以後， 我與他們所立的約是這樣的： 我要將我的律法放在他們的心上， 又要寫在他們的心思裏。」
HEB|10|17|並說： 「他們的罪惡和他們的過犯， 我絕不再記得。」
HEB|10|18|這些罪過既已蒙赦免，就不用再為罪獻祭了。
HEB|10|19|所以，弟兄們，既然我們靠著耶穌的血得以坦然進入至聖所，
HEB|10|20|是藉著他給我們開了一條又新又活的路，從幔子經過，這幔子就是他的身體。
HEB|10|21|既然我們有一位偉大祭司治理上帝的家，
HEB|10|22|那麼，我們該用誠心和充足的信心，同已蒙潔淨、無虧的良心，和清水洗淨了的身體來親近上帝。
HEB|10|23|我們要堅守所宣認的指望，毫不動搖，因為應許我們的那位是信實的。
HEB|10|24|我們要彼此相顧，激發愛心，勉勵行善；
HEB|10|25|不可停止聚會，好像那些停止慣了的人，倒要彼此勸勉，既然知道那日子臨近，就更當如此。
HEB|10|26|如果我們領受真理的知識以後仍故意犯罪，就不再有贖罪的祭物，
HEB|10|27|惟有戰戰兢兢等候審判和那將吞滅眾敵人的烈火了。
HEB|10|28|任何人干犯 摩西 的律法，憑兩個或三個證人，尚且必須處死，不得寬赦，
HEB|10|29|更何況踐踏上帝兒子的人，他們將那使他成聖之約的血當作不潔淨，又褻慢施恩的聖靈的人，你們想，他不該受更嚴厲的懲罰嗎？
HEB|10|30|因為我們知道誰說： 「伸冤在我， 我必報應。」 又說： 「主要審判他的百姓。」
HEB|10|31|落在永生上帝的手裏真是可怕呀！
HEB|10|32|你們要追念往日；你們蒙了光照以後，忍受了許多痛苦的掙扎：
HEB|10|33|一面在眾人面前公然被毀謗，遭患難；一面陪伴那些受這樣苦難的人。
HEB|10|34|你們同情那些遭監禁的人，也欣然忍受你們的家業被人搶去，因為你們知道自己有更美好更長存的家業。
HEB|10|35|所以，不可丟棄你們無懼的心，存這樣的心必得大賞賜。
HEB|10|36|你們必須忍耐，使你們行完了上帝的旨意，可以獲得所應許的。
HEB|10|37|因為 「還有一點點時候， 那要來的就來，必不遲延。
HEB|10|38|只是我的義人必因信得生； 他若退縮，我心就不喜歡他。」
HEB|10|39|我們卻不是退縮以致沉淪的那等人，而是有信心以致得生命的人。
HEB|11|1|信就是對所盼望之事有把握，對未見之事有確據。
HEB|11|2|古人因著這信獲得了讚許。
HEB|11|3|因著信，我們知道這宇宙是藉上帝的話造成的。這樣，看得見的是從看不見的造出來的。
HEB|11|4|因著信， 亞伯 獻祭給上帝比 該隱 所獻的更美，因此獲得了讚許為義人，上帝親自悅納了他的禮物。他雖然死了，卻因這信仍舊在說話。
HEB|11|5|因著信， 以諾 被接去，得以不見死，人也找不著他，因為上帝已經把他接去了；只是他被接去以前，已討得上帝的喜悅而蒙讚許。
HEB|11|6|沒有信，就不能討上帝的喜悅，因為到上帝面前來的人必須信有上帝，並且信他會賞賜尋求他的人。
HEB|11|7|因著信， 挪亞 既蒙上帝指示他未見的事，動了敬畏的心，造了方舟，使他全家得救。藉此他定了那世代的罪，自己也承受了那從信而來的義。
HEB|11|8|因著信， 亞伯拉罕 蒙召的時候就遵命出去，往將來要承受為基業的地方去；他出去的時候還不知往哪裏去。
HEB|11|9|因著信，他就在所應許之地作客，好像在異鄉，居住在帳棚裏，與蒙同一個應許的 以撒 和 雅各 一樣。
HEB|11|10|因為他等候著那座有根基的城，就是上帝所設計和建造的。
HEB|11|11|因著信， 撒拉 自己已過了生育的年齡還能懷孕，因為她認為應許她的那位是可信的 ；
HEB|11|12|所以，從一個彷彿已死的人竟生出子孫，如同天上的星那樣眾多，海邊的沙那樣無數。
HEB|11|13|這些人都是存著信心死的，並沒有得著所應許的，卻從遠處觀望，且歡喜迎接。他們承認自己在地上是客旅，是寄居的。
HEB|11|14|說這樣話的人是表明自己要尋找一個家鄉。
HEB|11|15|他們若想念所離開的家鄉，還有回去的機會。
HEB|11|16|其實他們所羨慕的是一個更美的，就是在天上的家鄉。所以，上帝並不因他們稱他為上帝 而覺得羞恥，因為他已經為他們預備了一座城。
HEB|11|17|因著信， 亞伯拉罕 被考驗的時候把 以撒 獻上，這就是那領受了應許的人甘心把自己獨生的兒子獻上。
HEB|11|18|論到這兒子，上帝曾說：「從 以撒 生的才要稱為你的後裔。」
HEB|11|19|他認為上帝甚至能使人從死人中復活，意味著他得回了他的兒子。
HEB|11|20|因著信， 以撒 指著將來的事給 雅各 、 以掃 祝福。
HEB|11|21|因著信， 雅各 臨死的時候給 約瑟 的兩個兒子個別祝福，扶著枴杖敬拜上帝。
HEB|11|22|因著信， 約瑟 臨終的時候提到 以色列 人將來要出 埃及 ，並為自己的骸骨留下遺言。
HEB|11|23|因著信， 摩西 生下來，他的父母見他是個俊美的孩子，把他藏了三個月，並不怕王的命令。
HEB|11|24|因著信， 摩西 長大了不肯稱為法老女兒之子。
HEB|11|25|他寧可和上帝的百姓一同受苦，也不願在罪中享受片刻的歡樂。
HEB|11|26|他把為彌賽亞受凌辱看得比 埃及 的財物更寶貴，因為他想望所要得的賞賜。
HEB|11|27|因著信，他離開 埃及 ，不怕王的憤怒，因為他恆心忍耐，如同看見那不能看見的上帝。
HEB|11|28|因著信，他設立逾越節，在門上灑血，免得那毀滅者加害 以色列 人的長子。
HEB|11|29|因著信，他們過 紅海 如行乾地； 埃及 人試著要過去就被淹沒了。
HEB|11|30|因著信， 以色列 人圍繞 耶利哥城 七日，城牆就倒塌了。
HEB|11|31|因著信，妓女 喇合 曾友善地接待探子，就沒有跟那些不順從的人一同滅亡。
HEB|11|32|我還要說甚麼呢？若要一一細說 基甸 、 巴拉 、 參孫 、 耶弗他 、 大衛 、 撒母耳 和眾先知的事，時間就不夠了。
HEB|11|33|他們藉著信，制伏了敵國，行了公義，得了應許，堵住了獅子的口，
HEB|11|34|滅了烈火的威力，在鋒利的刀劍下逃生，從軟弱變為剛強，爭戰中顯出勇猛，打退外邦的全軍。
HEB|11|35|有些婦人得回從死人中復活的親人。又有人忍受嚴刑，拒絕被釋放，為要得著更美好的復活。
HEB|11|36|又有人忍受戲弄、鞭打、捆鎖、監禁、各等的磨煉；
HEB|11|37|他們被石頭打死，被鋸鋸死， 被刀殺，披著綿羊山羊的皮各處奔跑，受貧窮、患難、虐待。
HEB|11|38|這世界配不上他們，他們在曠野、山嶺、山洞、地穴，飄流無定。
HEB|11|39|這些人都是因信獲得了讚許，卻仍未得著所應許的，
HEB|11|40|因為上帝給我們預備了更美好的事，若沒有我們，他們就不能達到完全。
HEB|12|1|所以，既然我們有這許多見證人如同雲彩圍繞著我們，就該卸下各樣重擔和緊緊纏累的罪，以堅忍的心奔那擺在我們前頭的路程，
HEB|12|2|仰望我們信心的創始成終者耶穌，他因那擺在前面的喜樂，輕看羞辱，忍受了十字架的苦難，如今已坐在上帝寶座的右邊。
HEB|12|3|你們要仔細想想這位忍受了罪人如此頂撞的耶穌，你們就不致心灰意懶了。
HEB|12|4|你們與罪惡爭鬥，還沒有抵抗到流血的地步。
HEB|12|5|你們又忘了上帝勸你們如同勸兒女的那些話，說： 「我兒啊，不可輕看主的管教， 被他責備的時候不可灰心；
HEB|12|6|因為主所愛的，他必管教， 又鞭打他所接納的每一個孩子。」
HEB|12|7|為了受管教，你們要忍受。上帝待你們如同待兒女。哪有兒女不被父親管教的呢？
HEB|12|8|管教原是眾兒女共同所領受的；你們若不受管教，就是私生子，不是兒女了。
HEB|12|9|再者，我們曾有肉身之父管教我們，我們尚且敬重他，何況靈性之父，我們豈不更當順服他而得生命嗎？
HEB|12|10|肉身之父都是短時間隨己意管教我們，惟有靈性之父管教我們是要我們得益處，使我們在他的聖潔上有份。
HEB|12|11|凡管教的事，當時不覺得快樂，反覺得痛苦；後來卻為那經過鍛鍊的人結出平安的果子，就是義的果子。
HEB|12|12|所以，你們要把下垂的手舉起來，發酸的腿挺直；
HEB|12|13|要為自己的腳把道路修直了，使瘸了的腿不再脫臼，反而得到痊癒。
HEB|12|14|你們要追求與眾人和睦，並要追求聖潔；人非聖潔不能見主。
HEB|12|15|要謹慎，免得有人失去了上帝的恩典；免得有毒根生出來擾亂你們，因而使許多人沾染污穢，
HEB|12|16|免得有人淫亂，或不敬虔如 以掃 ，他因一點點食物把自己長子的名分賣了。
HEB|12|17|後來你們知道，他想要承受父親的祝福，竟被拒絕，雖然流著淚苦求，卻得不著門路使他父親回心轉意。
HEB|12|18|你們不是來到那可觸摸的山，那裏有火焰、密雲、黑暗、暴風、
HEB|12|19|角聲，和說話的聲音；當時那些聽見這聲音的，都求不要再向他們說話，
HEB|12|20|因為他們擔當不起所命令他們的話，說：「靠近這山的，即使是走獸，也要用石頭打死。」
HEB|12|21|所見的景象極其可怕，以致 摩西 說：「我恐懼戰兢。」
HEB|12|22|但是你們是來到 錫安山 ，永生上帝的城，就是天上的 耶路撒冷 ，那裏有千千萬萬的天使，
HEB|12|23|有名字記錄在天上眾長子的盛會，有審判眾人的上帝和成為完全的義人的靈魂，
HEB|12|24|並新約的中保耶穌，以及所灑的血；這血所說的信息比 亞伯 的血所說的更美。
HEB|12|25|你們總要謹慎，不可拒絕那向你們說話的，因為那些拒絕了在地上警戒他們的，尚且不能逃罪，何況我們違背那從天上警戒我們的呢？
HEB|12|26|當時他的聲音震動了地，但如今他應許說：「再一次我不單要震動地，還要震動天。」
HEB|12|27|這「再一次」的話是指明被震動的要像受造之物一樣被挪去，使那不被震動的能常存。
HEB|12|28|所以，既然我們得了不能被震動的國度，就要感恩，照著上帝所喜悅的，用虔誠、敬畏的心事奉上帝，
HEB|12|29|因為我們的上帝是吞滅的火。
HEB|13|1|你們務要常存弟兄相愛的心。
HEB|13|2|不可忘記用愛心接待旅客，因為曾經有人這樣做，在無意中接待了天使。
HEB|13|3|要記念受監禁的人，好像與他們同受監禁；要記念受虐待的人，好像你們也親身受虐待一樣。
HEB|13|4|婚姻，人人都當尊重，共眠的床也不可污穢，因為淫亂和通姦的人，上帝必審判。
HEB|13|5|不可貪愛錢財，要以自己所有的為滿足，因為上帝曾說：「我絕不撇下你，也絕不丟棄你。」
HEB|13|6|所以，我們可以勇敢地說： 「主是我的幫助， 我必不懼怕。 人能把我怎麼樣呢？」
HEB|13|7|從前引導你們、傳上帝的道給你們的人，你們要記念他們，效法他們的信心，回顧他們為人的結局。
HEB|13|8|耶穌基督昨日、今日，一直到永遠，是一樣的。
HEB|13|9|你們不要被種種怪異的教訓勾引了去，因為人的心靠恩典得堅固才是好的，並不是靠飲食。那在飲食上用心的，從來沒有得到益處。
HEB|13|10|我們有一祭壇，上面的祭物是那些在會幕中供職的人無權可吃的。
HEB|13|11|因為牲畜的血被大祭司帶入至聖所作贖罪祭，牲畜的體卻在營外燒掉。
HEB|13|12|所以，耶穌也在城門外受苦，為要用自己的血使百姓成聖。
HEB|13|13|這樣，我們也當走出營外，到他那裏去，忍受他所受的凌辱。
HEB|13|14|在這裏，我們本沒有永存的城，而是在尋求那將要來的城。
HEB|13|15|我們應當藉著耶穌，常常以頌讚為祭獻給上帝，這是那宣認他名的人嘴唇所結的果子。
HEB|13|16|只是不可忘記行善和分享，因為這樣的祭物是上帝所喜悅的。
HEB|13|17|你們要服從那些引導你們的，並且要順服，因為他們為你們的靈魂時刻警醒，像在上帝面前交賬的人，讓他們在交賬的時候有喜樂，而不是嘆息，嘆息就對你們無益了。
HEB|13|18|請你們為我們禱告；因為我們自覺良心無虧，願意凡事按正道而行。
HEB|13|19|我更求你們為我禱告，使我快些回到你們那裏去。
HEB|13|20|但願賜平安 的上帝，就是那憑永約之血，把群羊的大牧人—我們主耶穌從死人中領出來的上帝，
HEB|13|21|在各樣善事上裝備你們，使你們遵行他的旨意；又藉著耶穌基督在我們 裏面行他所喜悅的事。願榮耀歸給他，直到永永遠遠 。阿們！
HEB|13|22|弟兄們，我簡略地寫信給你們，希望你們聽我勸勉的話。
HEB|13|23|你們該知道，我們的弟兄 提摩太 已經重獲自由了；他若很快就來，我必同他去見你們。
HEB|13|24|請你們向帶領你們的諸位和眾聖徒問安。從 意大利 來的人也向你們問安。
HEB|13|25|願恩惠與你們眾人同在。
JAS|1|1|上帝和主耶穌基督的僕人 雅各 問候散居在各處的十二個支派的人。
JAS|1|2|我的弟兄們，你們遭受各種試煉時，都要認為是大喜樂，
JAS|1|3|因為知道你們的信心經過考驗，就生忍耐。
JAS|1|4|但要讓忍耐發揮完全的功用，使你們能又完全又完整，一無所缺。
JAS|1|5|你們中間若有缺少智慧的，該求那厚賜與眾人又不斥責人的上帝，上帝必賜給他。
JAS|1|6|只要憑著信心求，一點也不疑惑；因為那疑惑的人，就像海中的波浪被風吹動翻騰。
JAS|1|7|這樣的人不要想從主那裏得到甚麼。
JAS|1|8|三心二意的人，在他一切所行的路上都搖擺不定。
JAS|1|9|卑微的弟兄要因高升而誇耀，
JAS|1|10|富足的卻要因被降卑而誇耀，因為富足的人要消逝，如同草上的花一樣。
JAS|1|11|太陽出來，熱風颳起，草就枯乾，花也凋謝，它美麗的樣子就消失了；那富足的人在他一生的奔波中也要這樣衰殘。
JAS|1|12|忍受試煉的人有福了，因為他經過考驗以後必得生命的冠冕，這是主應許給愛他之人的。
JAS|1|13|人被誘惑，不可說：「我是被上帝誘惑」；因為上帝是不被惡誘惑的，他也不誘惑人。
JAS|1|14|但每一個人被誘惑是因自己的私慾牽引而被誘惑的。
JAS|1|15|私慾既懷了胎，就生出罪來；罪既長成，就生出死來。
JAS|1|16|我親愛的弟兄們，不要被欺騙了。
JAS|1|17|各樣美善的恩澤和各樣完美的賞賜都是從上頭來的，從眾光之父那裏降下來的；在他並沒有改變，也沒有轉動的影兒。
JAS|1|18|他按自己的旨意，用真理的道生了我們，使我們在他所造的萬物中成為初熟的果子。
JAS|1|19|我親愛的弟兄們，你們要明白：你們每一個人要快快地聽，慢慢地說，慢慢地動怒，
JAS|1|20|因為人的怒氣並不能實現上帝的義。
JAS|1|21|所以，你們要除去一切的污穢和累積的惡毒，要存溫柔的心領受所栽種的道，就是能救你們靈魂的道。
JAS|1|22|但是，你們要作行道的人，不要只作聽道的人，自己欺騙自己。
JAS|1|23|因為只聽道而不行道的，就像人對著鏡子觀看自己本來的面目，
JAS|1|24|注視後，就離開，立刻忘了自己的相貌如何。
JAS|1|25|惟有查看那完美、使人自由的律法，並且時常遵守的，他不是聽了就忘，而是切實行出來，這樣的人在所行的事上必然蒙福。
JAS|1|26|若有人自以為虔誠，卻不勒住自己的舌頭，反欺騙自己的心，這人的虔誠是徒然的。
JAS|1|27|在上帝—我們的父面前，清潔沒有玷污的虔誠就是看顧在患難中的孤兒寡婦，並且保守自己不沾染世俗。
JAS|2|1|我的弟兄們，你們信奉我們榮耀的主耶穌基督，就不可按著外貌待人。
JAS|2|2|若有一個人戴著金戒指，穿著華麗的衣服，進入你們的會堂，又有一個窮人穿著骯髒的衣服也進去，
JAS|2|3|而你們只看重那穿華麗衣服的人，說：「請坐在這裏」，又對那窮人說：「你站在那裏」，或「坐在我腳凳旁」；
JAS|2|4|這豈不是你們偏心待人，用惡意評斷人嗎？
JAS|2|5|我親愛的弟兄們，請聽，上帝豈不是揀選了世上的貧窮人，使他們在信心上富足，並承受他所應許給那些愛他之人的國嗎？
JAS|2|6|你們卻羞辱貧窮的人。欺壓你們，拉你們到公堂去的，不就是這些富有的人嗎？
JAS|2|7|毀謗為你們求告時所奉的尊名的，不就是他們嗎？
JAS|2|8|經上記著：「要愛鄰 如己」，你們若切實守這至尊的律法，你們就做得很好。
JAS|2|9|但你們若按外貌待人就是犯罪，是被律法定為犯法的。
JAS|2|10|因為凡遵守全部律法的，只違背了一條就是違犯了所有的律法。
JAS|2|11|原來那說「不可姦淫」的，也說「不可殺人」。你就是不姦淫，卻殺人，也是成為違犯律法的。
JAS|2|12|既然你們要按使人自由的律法受審判，就要照這律法說話行事。
JAS|2|13|因為對那不憐憫人的，他們要受沒有憐憫的審判；憐憫勝過審判。
JAS|2|14|我的弟兄們，若有人說自己有信心，卻沒有行為，有甚麼益處呢？這信心能救他嗎？
JAS|2|15|若是弟兄或是姊妹沒有衣服穿，又缺少日用的飲食；
JAS|2|16|你們中間有人對他們說：「平平安安地去吧！願你們穿得暖，吃得飽」，卻不給他們身體所需要的，這有甚麼益處呢？
JAS|2|17|信心也是這樣，若沒有行為是死的。
JAS|2|18|但是有人會說：「你有信心，我有行為。」把你沒有行為的信心給我看，我就藉著我的行為把我的信心給你看。
JAS|2|19|你信上帝只有一位，你信得很好；連鬼魔也信，且怕得發抖。
JAS|2|20|你這虛浮的人哪，你願意知道沒有行為的信心是沒有用的嗎？
JAS|2|21|我們的祖宗 亞伯拉罕 把他兒子 以撒 獻在壇上，豈不是因行為得稱義嗎？
JAS|2|22|可見信心是與他的行為相輔並行，而且信心是因著行為才得以成全的。
JAS|2|23|這正應驗了經上所說：「 亞伯拉罕 信了上帝，這就算他為義」；他又得稱為上帝的朋友。
JAS|2|24|這樣看來，人稱義是因著行為，不是單因著信。
JAS|2|25|同樣，妓女 喇合 接待使者，又放他們從另一條路出去，不也是因行為稱義嗎？
JAS|2|26|所以，就如身體沒有靈魂是死的，信心沒有行為也是死的。
JAS|3|1|我的弟兄們，不要許多人做教師，因為你們知道，我們做教師的要接受更嚴厲的審判。
JAS|3|2|原來我們在許多事上都有過失；若有人在言語上沒有過失，他就是完全的人，也能勒住自己的全身。
JAS|3|3|我們若把嚼環放在馬嘴裏使牠們馴服，就能控制牠們的全身。
JAS|3|4|再看船隻，雖然甚大，又被強風猛吹，只用小小的舵就隨著掌舵的意思轉動。
JAS|3|5|同樣，舌頭是小肢體，卻能說大話。 看哪，最小的火能點燃最大的樹林。
JAS|3|6|舌頭就是火。在我們百體中，舌頭是個不義的世界，能玷污全身，也能燒燬生命的輪子，而且是被地獄的火點燃的。
JAS|3|7|各類的走獸、飛禽、爬蟲、水族，本來都可以制伏，也已經被人制伏了；
JAS|3|8|惟獨舌頭沒有人能制伏，是永不靜止的邪惡，充滿了害死人的毒氣。
JAS|3|9|我們用舌頭頌讚我們的主—我們的天父，又用舌頭詛咒照著上帝形像被造的人。
JAS|3|10|頌讚和詛咒從同一個口出來。我的弟兄們，這是不應該的。
JAS|3|11|泉源能從一個出口發出甜苦兩樣的水嗎？
JAS|3|12|我的弟兄們，無花果樹能生橄欖嗎？葡萄樹能結無花果嗎？鹹水也不能流出甜水來。
JAS|3|13|你們中間誰是有智慧有見識的呢？他就當在智慧的溫柔上顯出他的善行來。
JAS|3|14|你們心裏若懷著惡毒的嫉妒和自私，就不可自誇，不可說謊話抵擋真理。
JAS|3|15|這樣的智慧不是從上頭下來的，而是屬地上的，屬情慾的，屬鬼魔的。
JAS|3|16|在何處有嫉妒、自私，在何處就有動亂和各樣的壞事。
JAS|3|17|惟獨從上頭來的智慧，先是清潔，後是和平、溫良、柔順，滿有憐憫和美善的果子，沒有偏私，沒有虛偽。
JAS|3|18|正義的果實是為促進和平的人用和平栽種出來的。
JAS|4|1|你們中間的衝突是哪裏來的？爭執是哪裏來的？不是從你們肢體中交戰著的私慾來的嗎？
JAS|4|2|你們貪戀，得不著就殺人；你們嫉妒，不能得手就起爭執和衝突；你們得不著，是因為你們不求。
JAS|4|3|你們求也得不著，是因為你們妄求，為了要浪費在你們的宴樂中。
JAS|4|4|你們這些淫亂的人哪，豈不知道與世俗為友就是與上帝為敵嗎？所以，凡想要與世俗為友的，就是與上帝為敵了。
JAS|4|5|經上說：「上帝愛安置在我們裏面的靈，愛到嫉妒的地步。」 你們以為這話是徒然的嗎？
JAS|4|6|但是他賜更多的恩典，正如經上說： 「上帝抵擋驕傲的人， 但賜恩給謙卑的人。」
JAS|4|7|所以，要順服上帝。要抵擋魔鬼，魔鬼就必逃避你們；
JAS|4|8|要親近上帝，上帝就必親近你們。有罪的人哪，要潔淨你們的手！心懷二意的人哪，要清潔你們的心！
JAS|4|9|你們要愁苦，悲哀，哭泣；要將歡笑變為悲哀，歡樂變為愁悶。
JAS|4|10|要在主面前謙卑，他就使你們高升。
JAS|4|11|弟兄們，不可彼此詆毀。詆毀弟兄或評斷弟兄的人，就是詆毀律法，評斷律法；你若評斷律法，就不是遵行律法，而是評斷者了。
JAS|4|12|立法者和審判者只有一位；他就是那能拯救人也能毀滅人的。你是誰，竟敢評斷你的鄰舍！
JAS|4|13|注意！有人說：「今天或明天我們要往某城去，在那裏住一年，做買賣賺錢。」
JAS|4|14|其實明天如何，你們還不知道。你們的生命是甚麼呢？你們 原來是一片雲霧，出現片刻就不見了。
JAS|4|15|你們倒應當說：「主若願意，我們就能活著，也可以做這事或那事。」
JAS|4|16|現今你們竟然狂傲自誇；凡這樣的自誇都是邪惡的。
JAS|4|17|所以，人若知道該行善而不去行，這就是他的罪了。
JAS|5|1|注意！你們這些富足人哪，要為將要臨到你們身上的災難哭泣、號咷。
JAS|5|2|你們的財物腐爛了，你們的衣服被蟲子蛀了。
JAS|5|3|你們的金銀都生銹了；這銹要證明你們的不是，又要像火一樣吞吃你們的肉。你們在這末世只知道積蓄錢財。
JAS|5|4|工人給你們收割莊稼，你們剋扣他們的工錢；這工錢在喊冤，而且收割工人的冤聲已經進入萬軍之主的耳朵了。
JAS|5|5|你們在地上享奢華宴樂，把自己養肥了，等候宰殺的日子。
JAS|5|6|你們定了義人的罪，把他殺害，他沒有抵抗你們。
JAS|5|7|所以弟兄們，你們要忍耐，直到主來。看哪，農夫等候著地裏寶貴的出產，耐心地等到它得了秋霖春雨。
JAS|5|8|你們也要忍耐，堅固你們的心，因為主來的日子近了。
JAS|5|9|弟兄們，你們不要彼此埋怨，免得受審判。看哪，審判的主站在門口了。
JAS|5|10|弟兄們，你們要把那先前奉主名說話的眾先知作能受苦、能忍耐的榜樣。
JAS|5|11|看哪，那些忍耐的人，我們稱他們是有福的。你們聽見過 約伯 的忍耐，也看見主給他的結局，知道主是充滿憐憫和慈悲的。
JAS|5|12|我的弟兄們，最要緊的是不可起誓；不可指著天起誓，也不可指著地起誓，任何誓都不可起。你們說話，是，就說是；不是，就說不是，免得你們落在審判之下。
JAS|5|13|你們中間若有人受苦，他該禱告；有人喜樂，他該歌頌。
JAS|5|14|你們中間若有人病了，他該請教會的長老們來為他禱告，奉主的名為他抹油。
JAS|5|15|出於信心的祈禱必能救那病人，主必叫他起來；他若犯了罪，也必蒙赦免。
JAS|5|16|所以，你們要彼此認罪，互相代求，使你們得醫治。義人祈禱所發的力量是大有功效的。
JAS|5|17|以利亞 與我們是同樣性情的人，他懇切地祈求不要下雨，地上就三年六個月沒有下雨。
JAS|5|18|他又禱告，天就降下雨來，地就有了出產。
JAS|5|19|我的弟兄們，你們中間若有人迷失了真理而有人使他回轉，
JAS|5|20|這人該知道，使一個罪人從迷途中回轉，會從死亡中把他的靈魂救回來，而且遮蓋許多的罪。
1PET|1|1|耶穌基督的使徒 彼得 寫信給那些被揀選，分散在 本都 、 加拉太 、 加帕多家 、 亞細亞 、 庇推尼 寄居的人，
1PET|1|2|就是照父上帝的預知，藉著聖靈得以成聖，以致順服耶穌基督，又蒙他血所灑的人。願恩惠、平安 多多地賜給你們！
1PET|1|3|願頌讚歸於我們主耶穌基督的父上帝！他曾照自己的大憐憫，藉著耶穌基督從死人中復活，重生了我們，使我們有活的盼望，
1PET|1|4|好得到不朽壞、不玷污、不衰殘、為你們存留在天上的基業，
1PET|1|5|就是為你們這些藉著信、蒙上帝大能保守的人，能獲得他所預備、到末世要顯現的救恩。
1PET|1|6|雖然你們必須在百般試煉中暫時憂愁，你們要為此喜樂 ，
1PET|1|7|使你們的信心既被考驗，就比那被火試煉仍然能壞的金子更顯寶貴，可以在耶穌基督顯現的時候得著稱讚、榮耀、尊貴。
1PET|1|8|雖然你們沒有見過他，卻是愛他；如今雖看不見，你們卻因信他而有說不出來、滿有榮光的喜樂，
1PET|1|9|因為你們 得到信心的效果，就是靈魂的得救。
1PET|1|10|論到這救恩，那預先說你們要得恩典的眾先知已經詳細地搜索查考過，
1PET|1|11|查考在他們心裏的基督的靈預先證明基督受苦難，後來得榮耀，是指甚麼時候，甚麼樣的情況。
1PET|1|12|他們得了啟示，知道他們所服事的不是自己，而是你們。那藉著從天上差來的聖靈傳福音給你們的人，現在將這些事傳給你們；這些事連天使也都切望察看呢！
1PET|1|13|所以，要準備 好你們的心，謹慎自守，專心盼望耶穌基督顯現的時候帶給你們的恩惠。
1PET|1|14|作為順服的兒女，就不要效法從前蒙昧無知的時候那放縱私慾的樣子。
1PET|1|15|但那召你們的既是聖潔，你們在一切所行的事上也要聖潔；
1PET|1|16|因為經上記著：「你們要成為聖，因為我是神聖的。」
1PET|1|17|既然你們稱那不偏待人、按各人行為審判人的主為父 ，就當存敬畏的心，度你們在世寄居的日子。
1PET|1|18|你們知道，你們得以從你們祖先傳下來虛妄的行為中救贖出來，不是靠著會朽壞的金銀等物，
1PET|1|19|而是憑著基督的寶血，如同無瑕疵、無玷污的羔羊的血。
1PET|1|20|基督是上帝在創世以前所預知，而在這末世才為你們顯現的。
1PET|1|21|你們也因著他而信那使他從死人中復活、又給他榮耀的上帝，好讓你們的信心和盼望都在於上帝。
1PET|1|22|既然你們因順從真理而潔淨了自己的心靈，能真誠愛弟兄，就該以清潔的心 彼此切實相愛。
1PET|1|23|你們蒙了重生，不是由於會朽壞的種子，而是由於不會朽壞的種子，是藉著上帝永活常存的道。
1PET|1|24|因為 「凡血肉之軀的盡都如草， 他的一切榮美像草上的花； 草必枯乾，花必凋謝，
1PET|1|25|惟有主的道永遠常存。」 這話就是傳給你們的福音。
1PET|2|1|所以，你們要除去一切的惡毒，一切詭詐、假善、嫉妒，和一切毀謗的話。
1PET|2|2|要愛慕那純淨的靈奶，像初生的嬰孩愛慕奶一樣，好使你們藉著它成長，以致得救，
1PET|2|3|因為你們已經嘗過主恩的滋味。
1PET|2|4|要親近主，他是活石，雖然被人所丟棄，卻是上帝所揀選、所珍貴的。
1PET|2|5|你們作為活石，要被建造成屬靈的殿，成為聖潔的祭司，藉著耶穌基督獻上蒙上帝悅納的屬靈祭物。
1PET|2|6|因為經上說： 「看哪，我把一塊石頭放在 錫安 — 一塊蒙揀選、珍貴的房角石； 信靠他的人必不蒙羞。」
1PET|2|7|所以，這石頭在你們信的人是珍貴的；在那不信的人卻有話說： 「匠人所丟棄的石頭 已作了房角的頭塊石頭。」
1PET|2|8|又說： 「作了絆腳的石頭， 使人跌倒的磐石。」 他們絆跌，因為不順從這道，這也是預定的。
1PET|2|9|不過，你們是被揀選的一族，是君尊的祭司，是神聖的國度，是屬上帝的子民，要使你們宣揚那召你們出黑暗入奇妙光明者的美德。
1PET|2|10|「你們從前不是子民， 現在卻成了上帝的子民； 從前未曾蒙憐憫， 現在卻蒙了憐憫。」
1PET|2|11|親愛的，你們是客旅，是寄居的，我勸你們要禁戒肉體的情慾；這情慾是與靈魂爭戰的。
1PET|2|12|你們在外邦人中要品行端正，好讓那些人，雖然毀謗你們是作惡的，會因看見你們的好行為而在鑒察 的日子歸榮耀給上帝。
1PET|2|13|你們為主的緣故要順服人的一切制度，或是在上的君王，
1PET|2|14|或是君王所派懲惡賞善的官員。
1PET|2|15|因為上帝的旨意原是要你們以行善來堵住糊塗無知人的口。
1PET|2|16|雖然你們是自由的，卻不可藉著自由遮蓋惡毒，總要作上帝的僕人。
1PET|2|17|務要尊重眾人；要敬愛教中的弟兄姊妹；要敬畏上帝；要尊敬君王。
1PET|2|18|你們作奴僕的，凡事要存敬畏的心順服主人；不但順服善良溫和的，就是乖僻的也要順服。
1PET|2|19|倘若你們為使良心對得起上帝，忍受冤屈的痛苦，這是可讚許的。
1PET|2|20|你們若因犯罪受責打而忍耐，有甚麼可稱讚的呢？但你們若因行善受苦而忍耐，這在上帝看來是可讚許的。
1PET|2|21|你們蒙召就是為此，因為基督也為你們受過苦，給你們留下榜樣，為要使你們跟隨他的腳蹤。
1PET|2|22|「他並沒有犯罪， 口裏也沒有詭詐。」
1PET|2|23|他被辱罵不還口，受害也不說威嚇的話，只將自己交託給公義的審判者。
1PET|2|24|他被掛在木頭上，親身擔當了我們的罪，使我們既然在罪上死，就得以在義上活。因他受的鞭傷，你們得了醫治。
1PET|2|25|你們從前好像迷路的羊，如今卻歸回你們靈魂的牧人和監督了。
1PET|3|1|同樣，你們作妻子的，要順服自己的丈夫，這樣，即使有不信從道理的丈夫，也會因妻子的品行，並非言語，而感化過來，
1PET|3|2|因為看見了你們敬虔純潔的品行。
1PET|3|3|你們不要藉外表來妝飾自己，如編頭髮，戴金飾，穿美麗的衣裳等，
1PET|3|4|而要有蘊藏在人內心不衰退的美，以溫柔嫻靜的心妝飾自己；這在上帝面前是極寶貴的。
1PET|3|5|因為古時仰賴上帝的聖潔婦人正是以此為妝飾，順服自己的丈夫。
1PET|3|6|就如 撒拉 聽從 亞伯拉罕 ，稱他為主。你們只要行善，不怕任何恐嚇，就成為 撒拉 的女兒了。
1PET|3|7|同樣，你們作丈夫的，要按情理 跟妻子共同生活，體貼女性是比較軟弱的器皿；要尊重她，因為她也與你一同承受生命之恩。這樣，你們的禱告就不會受阻礙。
1PET|3|8|總而言之，你們都要同心，彼此體恤，相愛如弟兄，存憐憫和謙卑的心。
1PET|3|9|不要以惡報惡，以辱罵還辱罵，倒要祝福，因為你們正是為此蒙召的，好使你們承受福氣。
1PET|3|10|因為經上說： 「凡要愛惜生命、 享受好日子的人， 要禁止舌頭不出惡言， 嘴唇不說詭詐的話。
1PET|3|11|也要棄惡行善， 尋求和睦，一心追求。
1PET|3|12|因為主的眼看顧義人， 他的耳聽他們的祈禱； 但主向行惡的人變臉。」
1PET|3|13|你們若熱心行善，有誰會害你們呢？
1PET|3|14|即使你們為義受苦，也是有福的。不要怕人的威嚇，也不要驚慌；
1PET|3|15|只要心裏奉主基督為聖，尊他為主。有人問你們心中盼望的理由，要隨時準備答覆；
1PET|3|16|不過，要以溫柔、敬畏的心回答。要存無虧的良心，使你們在何事上被毀謗，就在何事上使那些凌辱你們在基督裏有好品行的人自覺羞愧。
1PET|3|17|上帝的旨意若是要你們因行善受苦，這總比因行惡受苦好。
1PET|3|18|因為基督也曾一次為罪受苦 ， 就是義的代替不義的， 為要引領你們 到上帝面前。 在肉體裏，他被治死； 但在靈裏，他復活了。
1PET|3|19|他藉這靈也曾去向那些在監獄裏的靈傳道，
1PET|3|20|就是那些從前在 挪亞 預備方舟、上帝容忍等待的時候不信從的人。當時進入方舟，藉著水得救的不多，只有八個人。
1PET|3|21|這水所預表的洗禮，現在藉著耶穌基督的復活拯救你們，不是除掉肉體的污穢，而是向上帝懇求有無虧的良心。
1PET|3|22|耶穌已經到天上去，在上帝的右邊，眾天使、有權柄的、有權能的都服從了他。
1PET|4|1|既然基督在肉身受苦，你們也該將這樣的心志作為兵器，因為在肉身受過苦的已經與罪斷絕了，
1PET|4|2|使你們從今以後不再隨從人的情慾，只順從上帝的旨意，在世度餘下的光陰。
1PET|4|3|因為你們從前隨從外邦人的心意，生活在淫蕩、情慾、醉酒、荒宴、狂飲和可憎的偶像崇拜中，時候已經夠了。
1PET|4|4|在這些事上，他們見你們不與他們同奔放蕩無度的路就以為怪，毀謗你們。
1PET|4|5|他們必須在那位將要審判活人死人的主面前交賬。
1PET|4|6|為此，死人也曾有福音傳給他們，要使他們的肉體按著人受審判，他們的靈卻靠上帝活著。
1PET|4|7|萬物的結局近了。所以你們要謹慎自守，要警醒禱告。
1PET|4|8|最要緊的是彼此切實相愛，因為愛能遮掩許多的罪。
1PET|4|9|你們要互相款待，不發怨言。
1PET|4|10|人人要照自己所得的恩賜彼此服事，作上帝各種恩賜的好管家。
1PET|4|11|若有人講道，他要按著上帝的聖言講；若有人服事，他要按著上帝所賜的力量服事，好讓上帝在凡事上因耶穌基督得榮耀。願榮耀和權能都歸給他，直到永永遠遠。阿們！
1PET|4|12|親愛的，有火一般的考驗臨到你們，不要奇怪，似乎是遭遇非常的事；
1PET|4|13|倒要歡喜，因為你們是與基督一同受苦，使你們在他榮耀顯現的時候也可以歡喜快樂。
1PET|4|14|你們若為基督的名受辱罵是有福的，因為榮耀的靈，就是上帝的靈，在你們身上。
1PET|4|15|你們中間，不可有人因為殺人、偷竊、作惡、好管閒事而受苦。
1PET|4|16|若有人因是基督徒而受苦，不要引以為恥，倒要因這名而歸榮耀給上帝。
1PET|4|17|因為時候到了，審判要從上帝的家開始；若是先從我們開始，那麼，不信從上帝福音的人將有何等的結局呢？
1PET|4|18|「若是義人還僅僅得救， 不虔敬和犯罪的人將有何地可站呢？」
1PET|4|19|所以，照上帝旨意受苦的人要一心為善，將自己的靈魂交給那信實的造物主。
1PET|5|1|所以，我這同作長老，作基督受苦的證人和分享將來所要顯現的榮耀的人，勉勵在你們中間的長老們：
1PET|5|2|務要牧養在你們當中上帝的群羊，按著上帝的旨意照顧他們 ，不是出於勉強，而是出於甘心；也不是因為貪財，而是出於樂意。
1PET|5|3|不要轄制所託付你們的群羊，而是要作他們的榜樣。
1PET|5|4|到了大牧人顯現的時候，你們必得到那永不衰殘、榮耀的冠冕。
1PET|5|5|同樣，你們年輕的，要順服年長的。你們大家都要以謙卑當衣服穿上，彼此順服，因為 「上帝抵擋驕傲的人， 但賜恩給謙卑的人。」
1PET|5|6|所以，你們要謙卑服在上帝大能的手下，這樣，到了適當的時候，他必使你們升高。
1PET|5|7|你們要將一切的憂慮卸給上帝，因為他顧念你們。
1PET|5|8|務要謹慎，要警醒。因為你們的仇敵魔鬼，如同咆哮的獅子，走來走去，尋找可吞吃的人。
1PET|5|9|你們要用堅固的信心抵擋他，因為知道你們在世上的眾弟兄也正在經歷這樣的苦難。
1PET|5|10|那賜一切恩典的上帝曾在基督 裏召了你們，得享他永遠的榮耀，在你們暫受苦難之後，必要親自成全你們，堅固你們，賜力量給你們，建立你們 。
1PET|5|11|願權能歸給他，直到永永遠遠。阿們！
1PET|5|12|我簡單地寫了這信，託我所看為忠心的弟兄 西拉 交給你們，勸勉你們，又證明這恩是上帝真實的恩典；你們務要在這恩上站立得住。
1PET|5|13|在 巴比倫 與你們同蒙揀選的教會向你們問安。我兒子 馬可 也向你們問安。
1PET|5|14|你們要用愛心彼此親吻問安。願平安 歸給你們所有在基督裏的人！
2PET|1|1|耶穌基督的僕人和使徒 西門．彼得 寫信給那因我們的上帝和 救主耶穌基督的義，與我們同得一樣寶貴信心的人。
2PET|1|2|願恩惠、平安 ，因你們認識上帝和我們的主耶穌，多多加給你們！
2PET|1|3|上帝的神能已把一切關乎生命和虔敬的事賜給我們，因我們認識那用自己榮耀和美德召我們的上帝。
2PET|1|4|因此，他已把又寶貴又極大的應許賜給我們，使我們既脫離世上從情慾來的敗壞，就得分享上帝的本性。
2PET|1|5|正因這緣故，你們要分外地努力。有了信心，又要加上德行；有了德行，又要加上知識；
2PET|1|6|有了知識，又要加上節制；有了節制，又要加上忍耐；有了忍耐，又要加上虔敬；
2PET|1|7|有了虔敬，又要加上愛弟兄的心；有了愛弟兄的心，又要加上愛眾人的心。
2PET|1|8|你們有了這幾樣，再繼續增長，就必使你們在認識我們的主耶穌基督上，不至於懶散和不結果子了。
2PET|1|9|沒有這幾樣的人就是瞎眼，是短視，忘了他過去的罪已經得了潔淨。
2PET|1|10|所以，弟兄們，要更加努力，使你們的蒙召和被選堅定不移。你們實行這幾樣，就永不失腳。
2PET|1|11|這樣，必叫你們豐豐富富地得以進入我們主－救主耶穌基督永遠的國度。
2PET|1|12|雖然你們已經知道這些事，並且在你們已有的真道上得到堅固，我還是要常常提醒你們這些事。
2PET|1|13|我認為趁我還在這帳棚的時候，應該激發你們的記憶，
2PET|1|14|因為知道我脫離這帳棚的時候快到了，正如我們的主耶穌基督所指示我的。
2PET|1|15|我也要盡心竭力，使你們在我去世以後時常記念這些事。
2PET|1|16|我們從前把我們主耶穌基督的大能和他來臨的事告訴你們，並不是隨從一些捏造出來的無稽傳說，我們是曾經親眼見過他的威榮的人。
2PET|1|17|他從父上帝得尊貴榮耀的時候，從至高無上的榮耀有聲音出來，對他說：「這是我的愛子，我所喜悅的。」
2PET|1|18|我們同他在聖山的時候，親自聽見這聲音從天上出來。
2PET|1|19|我們有先知更確實的信息，你們要好好地留意這信息，如同留意照耀在暗處的明燈，直等到天亮，晨星在你們心裏升起的時候。
2PET|1|20|第一要緊的，你們要知道，經上所有的預言是不可隨私意解釋的，
2PET|1|21|因為預言從來沒有出於人意的，而是人被聖靈感動說出上帝的話來。
2PET|2|1|從前在民間有假先知起來；同樣，將來在你們中間也會有假教師，偷偷地引進使人滅亡的異端。他們甚至不認買他們的主人，自取迅速滅亡。
2PET|2|2|許多人會隨從他們淫蕩的行為，以致真理之道因他們的緣故被毀謗。
2PET|2|3|他們因貪婪，要用捏造的言語在你們身上取得利益。他們的懲罰，自古以來並不遲延；他們的滅亡也必迅速來到。
2PET|2|4|既然上帝沒有寬容犯了罪的天使，反而把他們丟在地獄裏，囚禁在幽暗中等候審判；
2PET|2|5|既然上帝也沒有寬容上古的世界，曾叫洪水臨到那不敬虔的世界，只保護了報公義信息的 挪亞 一家八口；
2PET|2|6|既然上帝判決了 所多瑪 和 蛾摩拉 ，將二城傾覆 ，焚燒成灰，作為後世不敬虔人的鑒戒，
2PET|2|7|只搭救了那常為惡人的淫蕩憂傷的義人 羅得 —
2PET|2|8|因為那義人住在他們當中，他正義的心因天天看見和聽見他們不法的事而傷痛；
2PET|2|9|那麼，主知道搭救敬虔的人脫離試煉，把不義的人留在懲罰之下等候審判的日子，
2PET|2|10|尤其那些隨從肉體、放縱污穢的情慾、藐視主的權威的人更是如此。 他們膽大任性，無懼地毀謗眾尊榮者；
2PET|2|11|就是天使，雖然力量權能更大，在對他們宣告從主來的審判的時候還不用毀謗的話 。
2PET|2|12|但這些人好像沒有理性的牲畜，生來就是要被捉拿宰殺的。他們毀謗自己所不知道的事，正在敗壞人的時候，自己也遭遇敗壞，
2PET|2|13|為所行的不義受不義的工錢。他們喜愛白晝狂歡，他們已被玷污，又有瑕疵，正與你們一同歡宴，以自己的詭詐為樂。
2PET|2|14|他們滿眼是淫色，是止不住的罪，引誘心不堅定的人，心中習慣了貪婪，正是被詛咒的種類。
2PET|2|15|他們離棄了正路，走入歧途，隨從 比珥 的兒子 巴蘭 的路； 巴蘭 就是那貪愛不義的工錢的人，
2PET|2|16|他卻為自己的過犯受了責備，而那不能說話的驢以人的聲音阻止了先知的狂妄。
2PET|2|17|這些人是無水的泉源，是狂風催逼的霧氣，有漆黑的幽暗為他們存留。
2PET|2|18|他們說虛妄誇大的話，用肉體的情慾和淫蕩的事引誘那些剛脫離錯謬生活的人。
2PET|2|19|他們應許人自由，自己卻作了腐敗的奴隸，因為人被誰制伏就是誰的奴隸。
2PET|2|20|倘若他們因認識我們的主和救主耶穌基督而得以脫離世上的污穢，後來又被污穢纏住，被制伏，他們末後的景況就比先前更不好了。
2PET|2|21|他們知道義路，竟背棄了傳授給他們那神聖的誡命，倒不如不知道為妙。
2PET|2|22|俗語說得好，這話正印證在他們身上了： 「狗轉過來吃自己所吐的；」 又說： 「豬洗淨了，又回到爛泥裏打滾。」
2PET|3|1|親愛的，我現在寫給你們的是第二封信。在這兩封信裏，我都提醒你們，激發你們真誠的心，
2PET|3|2|要你們記得聖先知預先所說的話和主—救主的命令，就是使徒所傳給你們的。
2PET|3|3|第一要緊的，你們要知道，在末世必有好譏誚的人隨從自己的私慾出來譏誚，
2PET|3|4|說：「他要來臨的應許在哪裏呢？因為從列祖長眠以來，萬物與起初創造的時候仍是一樣啊！」
2PET|3|5|他們故意忘記這事，就是從太古憑上帝的話有了天，並由水而出和藉著水而成的地；
2PET|3|6|藉著水，當時的世界被水淹沒而消滅了。
2PET|3|7|但現在的天地還是憑著上帝的話存留，直留到不敬虔之人受審判遭沉淪的日子，用火焚燒。
2PET|3|8|親愛的，有一件事你們不可忘記，就是：主看一日如千年，千年如一日。
2PET|3|9|主沒有遲延他的應許，就如有人以為他是遲延，其實他是寬容你們，不願一人沉淪，而是人人都來悔改。
2PET|3|10|但主的日子要像賊一樣來到；那日，天必在轟然一聲中消失，天體都要被烈火熔化，地和地上的萬物都要燒盡 。
2PET|3|11|既然這一切都要如此消失，你們 處世為人必須聖潔敬虔，
2PET|3|12|等候並催促上帝的日子來到。因為在那日，天要被火燒而消滅，天體都要被烈火熔化。
2PET|3|13|但照他的應許，我們等候新天新地，其中有正義常住。
2PET|3|14|所以，親愛的，既然你們等候這些事，就要竭力使自己沒有玷污，無可指責，在主前和睦；
2PET|3|15|並且要以我們主的容忍作為你們得救的機會，就如我們所親愛的弟兄 保羅 ，照著所賜給他的智慧寫信給你們。
2PET|3|16|他一切的信上都談到這事。信中有些難明白的，那無學問、不堅定的人加以曲解，如曲解別的經書一樣，自取滅亡。
2PET|3|17|所以，親愛的，既然你們預先知道這事，就當防備，免得被惡人的錯謬誘惑，從自己穩定的立場上墜落。
2PET|3|18|你們倒要在我們的主和救主耶穌基督的恩典和知識上有長進。願榮耀歸給他，從今直到永遠之日。阿們！
1JOHN|1|1|論到從起初原有的生命之道，就是我們所聽見、所看見、親眼看過、親手摸過的－
1JOHN|1|2|這生命已經顯現出來，我們看見了，現在又作見證，把原與父同在，並且向我們顯現過的那永遠的生命傳揚給你們－
1JOHN|1|3|我們把所看見、所聽見的傳揚給你們，為要使你們也與我們有團契，而我們的團契是與父和他兒子耶穌基督所共有的。
1JOHN|1|4|我們把這些事寫給你們，使我們 的喜樂得以滿足。
1JOHN|1|5|上帝就是光，在他毫無黑暗；這是我們從主所聽見，又報給你們的信息。
1JOHN|1|6|我們若說，我們與上帝有團契，卻仍在黑暗裏行走，就是說謊話，不實行真理了。
1JOHN|1|7|我們若在光明中行走，如同上帝在光明中，就彼此有團契，他兒子耶穌的血就洗淨我們一切的罪。
1JOHN|1|8|我們若說自己沒有罪，就是欺騙自己，真理就不在我們裏面了。
1JOHN|1|9|我們若認自己的罪，上帝是信實的，是公義的，必要赦免我們的罪，洗淨我們一切的不義。
1JOHN|1|10|我們若說自己沒有犯過罪，就是把上帝當作說謊的，他的道就不在我們裏面了。
1JOHN|2|1|我的孩子們哪，我把這些話寫給你們，是要你們不犯罪。若有人犯罪，在父那裏我們有一位中保，就是那義者耶穌基督。
1JOHN|2|2|他為我們的罪作了贖罪祭，不單是為我們的罪，也是為普天下人的罪。
1JOHN|2|3|我們若遵守上帝的命令，就知道我們確實認識他。
1JOHN|2|4|人若說「我認識他」，卻不遵守他的命令，就是說謊話的，真理就不在他裏面了。
1JOHN|2|5|凡遵守他的道的，愛上帝的心確實地在他裏面達到完全了。由此我們知道我們是在他裏面。
1JOHN|2|6|凡說自己住在他裏面的，就該照著他所行的去行。
1JOHN|2|7|親愛的，我寫給你們的不是一條新命令，而是你們從起初所受的舊命令；這舊命令就是你們所聽過的道。
1JOHN|2|8|然而，我寫給你們的是一條新命令，在基督裏是真實的，在你們也是真實的，因為黑暗漸漸消逝，真光已經在照耀。
1JOHN|2|9|人若說自己在光明中，卻恨他的弟兄，他到如今還是在黑暗裏。
1JOHN|2|10|那愛弟兄的，就是住在光明中，他不會使人失足犯罪 。
1JOHN|2|11|惟獨那恨弟兄的，是在黑暗裏，也在黑暗裏行走，不知道往哪裏去，因為黑暗使他的眼睛瞎了。
1JOHN|2|12|孩子們哪，我寫信給你們， 因為你們的罪藉著基督的名得了赦免。
1JOHN|2|13|父老們啊，我寫信給你們， 因為你們認識從起初就有的那一位。 青年們哪，我寫信給你們， 因為你們勝過了那惡者。
1JOHN|2|14|孩子們哪，我曾寫信給你們， 因為你們認識父。 父老們啊，我曾寫信給你們， 因為你們認識從起初就有的那一位。 青年們哪，我曾寫信給你們， 因為你們剛強， 上帝的道常存在你們心裏， 你們也勝過了那惡者。
1JOHN|2|15|不要愛世界和世界上的東西，若有人愛世界，愛父的心就不在他裏面了。
1JOHN|2|16|因為凡世界上的東西，好比肉體的情慾、眼目的情慾和今生的驕傲，都不是從父來的，而是從世界來的。
1JOHN|2|17|這世界和世上的情慾都要消逝，惟獨那遵行上帝旨意的人永遠常存。
1JOHN|2|18|孩子們哪，如今是末世的時光了。你們曾聽過那敵基督者要來，現在有好些敵基督者已經出來了；由此我們就知道，如今是末世的時光了。
1JOHN|2|19|他們從我們中間出去，卻不是屬我們的，若是屬我們的，就必仍舊與我們同在。他們出去，這就顯明他們都不是屬我們的。
1JOHN|2|20|你們從那聖者受了恩膏，並且你們大家都知道 。
1JOHN|2|21|我寫信給你們，不是因你們不認識真理，而是因你們認識，並且知道一切虛謊都不是從真理出來的。
1JOHN|2|22|誰是說謊話的呢？不就是那不認耶穌為基督的嗎？那不認父與子的，這個人就是敵基督的。
1JOHN|2|23|凡不認子的，就沒有父；宣認子的，連父也有了。
1JOHN|2|24|論到你們，務要將那從起初所聽見的常存在心裏；若將從起初所聽見的存在心裏，你們就會住在子裏面，也會住在父裏面。
1JOHN|2|25|基督所應許我們的就是永生。
1JOHN|2|26|我將這些話寫給你們，是論到那些迷惑你們的人說的。
1JOHN|2|27|至於你們，你們從基督所受的恩膏常存在你們心裏，並不用人教導你們，自有他的恩膏在凡事上教導你們。這恩膏是真的，不是假的，你們要按這恩膏的教導住在他裏面。
1JOHN|2|28|孩子們哪，你們要住在基督裏面。這樣，他若顯現，我們就可以坦然無懼；當他來臨的時候，在他面前不至於慚愧。
1JOHN|2|29|你們若知道他是公義的，就知道凡行公義的人都是他所生的。
1JOHN|3|1|你們看父賜給我們的是何等的慈愛，讓我們得以稱為上帝的兒女；我們也真是他的兒女。世人不認識我們 的理由，是因他們未曾認識父。
1JOHN|3|2|親愛的，我們現在是上帝的兒女，將來如何還未顯明。我們所知道的是：基督顯現的時候，我們會像他，因為我們將見到他的本相。
1JOHN|3|3|凡對他有這指望的，就潔淨自己，像他是潔淨的一樣。
1JOHN|3|4|凡犯罪的，就是做違背律法的事；違背律法就是罪。
1JOHN|3|5|你們知道，基督曾顯現是要除掉罪 ；在他並沒有罪。
1JOHN|3|6|凡住在他裏面的，不犯罪；凡犯罪的，未曾看見他，也未曾認識他。
1JOHN|3|7|孩子們哪，不要讓人迷惑了你們；行義的才是義人，正如基督是義的。
1JOHN|3|8|犯罪的是出於魔鬼，因為魔鬼從起初就犯罪。上帝的兒子顯現出來，是為了要毀滅魔鬼的作為。
1JOHN|3|9|凡從上帝生的，不犯罪，因上帝的道 存在他裏面，他也不能犯罪，因為他是由上帝所生的。
1JOHN|3|10|這就顯明誰是上帝的兒女，誰是魔鬼的兒女了。凡不行義的，不是出於上帝，不愛他弟兄的，也是如此。
1JOHN|3|11|我們要彼此相愛。這就是你們從起初所聽到的信息。
1JOHN|3|12|不要像 該隱 ；他是屬那邪惡者，殺了自己的弟弟。為甚麼殺了他呢？因為自己的行為是邪惡的，而弟弟的行為是正直的。
1JOHN|3|13|弟兄們，世人若恨你們，不要驚訝。
1JOHN|3|14|我們知道，我們已經出死入生了，因為我們愛弟兄。沒有愛心的，仍住在死中。
1JOHN|3|15|凡恨自己弟兄的，就是殺人的；你們知道，凡殺人的，沒有永生住在他裏面。
1JOHN|3|16|基督為我們捨命，我們從此就知道何為愛；我們也當為弟兄捨命。
1JOHN|3|17|凡有世上財物的，看見弟兄缺乏，卻關閉了惻隱的心，上帝的愛怎能住在他裏面呢？
1JOHN|3|18|孩子們哪，我們相愛，不要只在言語或舌頭上，總要以行為和真誠表現出來。
1JOHN|3|19|從這一點，我們會知道，我們是出於真理的，並且我們在上帝面前可以安心，
1JOHN|3|20|即使我們的心責備自己，上帝比我們的心大，他知道一切。
1JOHN|3|21|親愛的，我們的心若不責備我們，在上帝面前就可以坦然無懼了。
1JOHN|3|22|我們一切所求的，就從他得著，因為我們遵守他的命令，行他所喜悅的事。
1JOHN|3|23|上帝的命令就是：我們要信他兒子耶穌基督的名，並且照他所賜給我們的命令彼此相愛。
1JOHN|3|24|遵守上帝命令的，住在上帝裏面，而上帝也住在他裏面。從這一點，我們知道上帝住在我們裏面，這是由於他所賜給我們的聖靈。
1JOHN|4|1|親愛的，一切的靈不可都信，總要察驗那些靈是否出於上帝，因為有許多假先知已經來到世上。
1JOHN|4|2|凡宣認耶穌基督是成了肉身而來的靈就是出於上帝的，由此你們可以認出上帝的靈來；
1JOHN|4|3|凡不宣認耶穌的靈，不是出於上帝。這是那敵基督者的靈；你們從前聽見他要來，現在他已經在世上了。
1JOHN|4|4|孩子們哪，你們是屬上帝的，並且勝過了假先知，因為那在你們裏面的比那在世界上的更大。
1JOHN|4|5|他們是屬世界的，所以講論世界的事，而世人也聽從他們。
1JOHN|4|6|我們是屬上帝的，認識上帝的就聽從我們；不屬上帝的就不聽從我們。從此我們可以認出真理的靈和錯謬的靈來。
1JOHN|4|7|親愛的，我們要彼此相愛，因為愛是從上帝來的。凡有愛的都是由上帝而生，並且認識上帝。
1JOHN|4|8|沒有愛的就不認識上帝，因為上帝就是愛。
1JOHN|4|9|上帝差他獨一的兒子到世上來，使我們藉著他得生命；由此，上帝對我們的愛就顯明了。
1JOHN|4|10|不是我們愛上帝，而是上帝愛我們，差他的兒子為我們的罪作了贖罪祭；這就是愛。
1JOHN|4|11|親愛的，既然上帝這樣愛我們，我們也要彼此相愛。
1JOHN|4|12|從來沒有人見過上帝，我們若彼此相愛，上帝就住在我們裏面，他的愛在我們裏面得以完滿了。
1JOHN|4|13|因為上帝將他的靈賜給我們，由此我們知道我們是住在他裏面，而他也住在我們裏面。
1JOHN|4|14|父差子作世人的救主，這是我們所看見並且作見證的。
1JOHN|4|15|凡宣認耶穌為上帝兒子的，上帝就住在他裏面，而他也住在上帝裏面。
1JOHN|4|16|我們知道並且深信上帝是愛我們的。 上帝就是愛，住在愛裏面的就是住在上帝裏面；上帝也住在他裏面。
1JOHN|4|17|由此，愛在我們裏面得以完滿：我們可以在審判的日子坦然無懼，因為基督如何，我們在這世上也如何。
1JOHN|4|18|在愛裏沒有懼怕；完滿的愛把懼怕驅逐出去，因為懼怕裏含著懲罰，懼怕的人在愛裏尚未得到完滿。
1JOHN|4|19|我們愛，因為上帝先愛我們。
1JOHN|4|20|人若說「我愛上帝」，卻恨他的弟兄，就是說謊了；不愛他看得見的弟兄，就不能愛看不見的上帝 。
1JOHN|4|21|愛上帝的，也要愛弟兄；這是我們從上帝所受的命令。
1JOHN|5|1|凡信耶穌是基督的，都是從上帝生的；凡愛生他之上帝的，也必愛從上帝生的 。
1JOHN|5|2|我們愛上帝，又實行 他的命令，由此就知道我們愛上帝的兒女了。
1JOHN|5|3|我們遵守上帝的命令，這就是愛他了，而且他的命令並不是難守的。
1JOHN|5|4|因為凡從上帝生的就勝過世界；使我們勝過世界的就是我們的信心。
1JOHN|5|5|勝過世界的是誰呢？不就是那信耶穌是上帝兒子的嗎？
1JOHN|5|6|這藉著水和血而來的，就是耶穌基督，不是單用水，而是用水又用血，並且有聖靈作見證，因為聖靈就是真理。
1JOHN|5|7|作見證的有三：
1JOHN|5|8|就是聖靈、水與血，這三樣也都是一致的。
1JOHN|5|9|既然我們領受人的見證，上帝的見證更該領受 了，因為上帝的見證是為他兒子作的。
1JOHN|5|10|信上帝兒子的，就有這見證在他心裏；不信上帝的，就是把上帝當作說謊的，因為不信上帝為他兒子作的見證。
1JOHN|5|11|這見證就是：上帝賜給我們永生，而這永生是在他兒子裏面的。
1JOHN|5|12|那有上帝兒子的，就有生命；沒有上帝兒子的，就沒有生命。
1JOHN|5|13|我把這些話寫給你們信奉上帝兒子之名的人，要讓你們知道自己有永生。
1JOHN|5|14|我們若照著上帝的旨意祈求，他就垂聽我們；這就是我們對他所存坦然無懼的心。
1JOHN|5|15|既然我們知道他聽我們一切所求的，就知道我們所求於他的，無不得著。
1JOHN|5|16|人若看見弟兄犯了不至於死的罪，就要為他祈求，上帝必將生命賜給他—有些人犯的罪是不至於死的；有的是至於死的罪，我不是說要為這罪祈求。
1JOHN|5|17|一切不義的事都是罪，但也有不至於死的罪。
1JOHN|5|18|我們知道，凡從上帝生的，必不犯罪；從上帝生的那一位，必保守他，那邪惡者無法加害於他。
1JOHN|5|19|我們知道，我們是屬上帝的，而全世界都伏在那邪惡者的權勢之下。
1JOHN|5|20|我們知道，上帝的兒子已經來到，並且將悟性賜給我們，使我們認識那位真實者，我們也在那位真實者裏面，就是在他兒子耶穌基督裏面。這是真神，也是永生。
1JOHN|5|21|孩子們哪，你們要遠避偶像。
2JOHN|1|1|我作長老的寫信給蒙揀選的夫人 和她的兒女，就是我真心所愛的；不但我愛，也是一切認識真理的人所愛的，
2JOHN|1|2|這是因為真理住在我們裏面，也必與我們同在直到永遠。
2JOHN|1|3|願恩惠、憐憫、平安 從父上帝和他兒子耶穌基督，在真理和愛中必與我們同在。
2JOHN|1|4|我非常歡喜見你的兒女，有照我們從父所受之命令遵行真理的。
2JOHN|1|5|夫人哪，我現在請求你，我們大家要彼此相愛。我寫給你的，並不是一條新命令，而是我們從起初就有的。
2JOHN|1|6|這就是愛，就是照他的命令行事；這就是命令，你們要照這命令行，正如你們從起初所聽見的。
2JOHN|1|7|有許多迷惑人的已經來到世上，他們不宣認耶穌基督是成了肉身來的；這樣的人是迷惑人的，是敵基督的。
2JOHN|1|8|你們要小心，不要失去你們 所完成的工作，而要得到充足的賞賜。
2JOHN|1|9|凡越過基督的教導而不持守的，就沒有上帝；凡持守這教導的，就有父又有子。
2JOHN|1|10|若有人到你們那裏而不傳這教導，不要接他到家裏，也不要向他問安；
2JOHN|1|11|因為向他問安的，就在他的惡行上有份。
2JOHN|1|12|我還有許多事要寫給你們，卻不願意用紙用墨，但盼望到你們那裏，與你們面對面談論，使我們的喜樂得以滿足。
2JOHN|1|13|你那蒙揀選的姊妹的兒女向你問安。
3JOHN|1|1|我作長老的寫信給親愛的 該猶 ，就是我真心所愛的。
3JOHN|1|2|親愛的，我願你事事安寧，身體健康，正如你的心神安寧一樣。
3JOHN|1|3|我非常歡喜，有弟兄到這裏來，證實你對真理的忠誠，就是你按著真理而行。
3JOHN|1|4|我聽見我的兒女按真理而行，我的歡喜沒有比這個更大的。
3JOHN|1|5|親愛的，你對弟兄，特別是對作客旅的弟兄所做的都是忠誠的。
3JOHN|1|6|他們在教會面前證實了你的愛；你若以對得起上帝的方式，為他們送行就好了；
3JOHN|1|7|因為他們是為基督的名 出外，並沒有從未信的人接受甚麼。
3JOHN|1|8|所以，我們應當接待這樣的人，好讓我們與他們在真理上成為同工。
3JOHN|1|9|我曾寫過一些東西給教會，但他們中間那好作領袖的 丟特腓 不接納我們。
3JOHN|1|10|為此，我若去，要提起他所做的事，就是他用惡言攻擊我們，還不滿足，他自己不接納弟兄，有人願意接納，他還阻止，並且把接納弟兄的人趕出教會。
3JOHN|1|11|親愛的，不要效法惡，只要效法善。行善的人屬乎上帝；行惡的人未曾見過上帝。
3JOHN|1|12|低米丟 行善，有眾人給他作見證，又有真理給他作見證，就是我們也給他作見證，你知道我們的見證是真的。
3JOHN|1|13|我還有許多事要寫給你，卻不願意用筆墨來寫給你，
3JOHN|1|14|但盼望很快見到你，我們好面對面談論。
3JOHN|1|15|願你平安！朋友們都向你問安。請你替我按著名字一一向朋友們問安。
JUDE|1|1|耶穌基督的僕人、 雅各 的兄弟 猶大 ，寫信給那些被召、在父上帝裏蒙愛、為耶穌基督保守的人。
JUDE|1|2|願憐憫、平安 、慈愛多多加給你們！
JUDE|1|3|親愛的，我一直很迫切地想要寫信給你們，論到我們同享的救恩，但我覺得有必要現在就寫信勸你們，要為從前一次交付給聖徒的真道竭力奮鬥。
JUDE|1|4|因為有些人偷偷地進來，就是早就被判定受懲罰的不虔誠的人，他們把我們上帝的恩典變為放縱情慾的機會，並且不認獨一的主宰—我們的主耶穌基督。
JUDE|1|5|這一切的事，你們雖然知道，我卻仍要提醒你們：從前主 只一次就 救了他的百姓出 埃及 地，後來卻把那些不信的滅絕了。
JUDE|1|6|至於那些不守本位、離開自己住處的天使，主用鎖鏈把他們永遠拘留在黑暗裏，等候大日子的審判。
JUDE|1|7|同樣， 所多瑪 、 蛾摩拉 和周圍城鎮的人也跟著他們一樣犯淫亂，隨從逆性的情慾，以致遭受永不熄滅之火的懲罰，作為眾人的鑒戒。
JUDE|1|8|照樣，這些做夢的人也污穢身體，輕慢掌權者，毀謗眾尊榮者。
JUDE|1|9|天使長 米迦勒 為 摩西 的屍首與魔鬼爭辯的時候，尚且不敢用毀謗的話譴責他，只說：「主責備你吧！」
JUDE|1|10|但這些人毀謗他們所不知道的。他們與那些沒有理性的牲畜一樣，只做本性所知道的事，敗壞了自己。
JUDE|1|11|他們有禍了！因為他們走 該隱 的道路，又為財利往 巴蘭 的錯謬裏直奔，並在 可拉 的背叛中滅亡了。
JUDE|1|12|這樣的人是你們愛筵上的污點 ；他們無所懼怕地同你們宴樂，彷彿牧人只顧餵飽自己。他們是無雨的浮雲，被風飄蕩；是秋天沒有果子的樹，死而又死，連根被拔出來；
JUDE|1|13|是海裏的狂浪，湧出自己可恥的沫子來；是流蕩的星，有漆黑的幽暗永遠為他們保留著。
JUDE|1|14|亞當 的七世孫 以諾 曾預言這些人說：「看哪，主帶著他的千萬聖者來臨，
JUDE|1|15|要審判眾人，證實一切不敬虔的人所妄行一切不敬虔的事，又證實不敬虔的罪人所說頂撞他的剛愎的話。」
JUDE|1|16|這些人喜出怨言，責怪他人，隨從自己的情慾而行，口說誇大的話，為自己的利益諂媚人。
JUDE|1|17|親愛的，至於你們，要記得我們主耶穌基督的使徒從前所說的話。
JUDE|1|18|他們曾對你們說過，末世必有好嘲弄的人隨從自己不敬虔的私慾而行。
JUDE|1|19|這就是那些好結黨分派、屬乎血氣、沒有聖靈的人。
JUDE|1|20|親愛的，至於你們，要在至聖的真道上造就自己，藉著聖靈禱告，
JUDE|1|21|保守自己常在上帝的愛中，仰望我們主耶穌基督的憐憫，進入永生。
JUDE|1|22|有些人心中猶疑 ，你們要憐憫 他們；
JUDE|1|23|有些人你們要從火中搶出來，搭救他們 ；有些人你們要存懼怕的心憐憫他們，連那被情慾污染的衣服也要厭惡。
JUDE|1|24|願那能保守你們不失腳，使你們無瑕無疵、歡歡喜喜站在他榮耀之前的、
JUDE|1|25|我們的救主獨一的上帝，藉著我們的主耶穌基督，得享榮耀、威嚴、能力、權柄，從萬古以前，到現今，直到永永遠遠。阿們！
REV|1|1|耶穌基督的啟示，就是上帝賜給他，要他將必須快要發生的事指示他的眾僕人。他差遣使者指明給他的僕人 約翰 ，
REV|1|2|約翰 就將上帝的道和耶穌基督的見證，凡自己所看見的，都見證出來。
REV|1|3|誦讀這書上預言的，和那些聽見又遵守其中所記載的，都是有福的，因為時候近了。
REV|1|4|約翰 寫信給 亞細亞 的七個教會。願那位今在、昔在、以後永在的上帝，與他寶座前的七靈，和那忠信的見證者、從死人中復活的首生者 、世上君王的元首耶穌基督，賜恩惠和平安 給你們。 他愛我們，用自己的血使我們從罪中得釋放 ，
REV|1|5|
REV|1|6|又使我們成為國度，作他父上帝的祭司。願榮耀、權能歸給他，直到永永遠遠 。阿們！
REV|1|7|「看哪，他駕雲降臨； 眾目都要看見他， 連刺他的人也要看見他； 地上的萬族要因他哀哭。」 這是真實的。阿們！
REV|1|8|主上帝說：「我是阿拉法，我是俄梅戛 ，是今在、昔在、以後永在的全能者。」
REV|1|9|我— 約翰 就是你們的弟兄，在耶穌裏和你們一同在患難、國度、忍耐裏有份的，為上帝的道，並為給耶穌作的見證，曾在那名叫 拔摩 的海島上。
REV|1|10|有一主日我被聖靈感動，聽見在我後面有大聲音如吹號，
REV|1|11|說：「把你所看見的寫在書上，寄給 以弗所 、 士每拿 、 別迦摩 、 推雅推喇 、 撒狄 、 非拉鐵非 、 老底嘉 那七個教會。」
REV|1|12|我轉過身來要看看是誰的聲音在跟我說話。我一轉過來，看見了七個金燈臺；
REV|1|13|在燈臺中間有一位好像人子的，身穿垂到腳的長袍，胸間束著金帶。
REV|1|14|他的頭與髮皆白，如白羊毛，如雪；他的眼睛好像火焰，
REV|1|15|雙腳好像在爐中鍛鍊得發亮的銅，聲音好像眾水的聲音。
REV|1|16|他右手拿著七顆星，從他口中吐出一把兩刃的利劍，面貌好像烈日放光。
REV|1|17|我看見了他，就仆倒在他腳前，像死人一樣。他用右手按著我說：「不要怕。我是首先的，是末後的，
REV|1|18|又是永活的。我曾死過，看哪，我是活著的，直到永永遠遠；並且我拿著死亡和陰間的鑰匙。
REV|1|19|所以，你要把所看見的事、現在的事和以後將發生的事，都寫下來。
REV|1|20|至於你所看見、在我右手中的七顆星和那七個金燈臺的奧祕就是：七顆星是七個教會的使者，七個燈臺是七個教會。」
REV|2|1|「你要寫信給 以弗所 教會的使者，說：『那右手拿著七顆星，在七個金燈臺中間行走的這樣說：
REV|2|2|我知道你的行為、勞碌、忍耐，也知道你不容忍惡人。你也曾察驗那自稱為使徒卻不是使徒的，看出他們是假的。
REV|2|3|你能忍耐，曾為我的名勞苦而不困倦。
REV|2|4|然而，有一件事我要責備你，就是你把起初的愛心拋棄了。
REV|2|5|所以你要回想你是從哪裏墜落的，並且要悔改，做起初所做的工作。你若不悔改，我要到你那裏去，把你的燈臺從原處挪去。
REV|2|6|然而你還有一件可取的事，就是你恨惡 尼哥拉 派的行為，這種行為也是我所恨惡的。
REV|2|7|凡有耳朵的都應當聽聖靈向眾教會所說的話。得勝的，我必將上帝樂園中生命樹的果子賜給他吃。』」
REV|2|8|「你要寫信給 士每拿 教會的使者，說：『那首先的、末後的，死過又活了的這樣說：
REV|2|9|我知道你的患難和貧窮—其實你卻是富足的，也知道那自稱是 猶太 人的所說毀謗的話，其實他們不是 猶太 人，而是撒但會堂的人。
REV|2|10|你將要受的苦，你不用怕。看哪！魔鬼要把你們中間幾個人下在監裏，使你們受考驗，你們要遭受苦難十日。你務要至死忠心，我就賜給你那生命的冠冕。
REV|2|11|凡有耳朵的都應當聽聖靈向眾教會所說的話。得勝的必不受第二次死的害。』」
REV|2|12|「你要寫信給 別迦摩 教會的使者，說：『那有兩刃利劍的這樣說：
REV|2|13|我知道你的居所，就是有撒但座位之處；當我忠心的見證人 安提帕 在你們中間，在撒但所住的地方被殺之時，你還堅守我的名，沒有否認對我的信仰。
REV|2|14|然而，有幾件事我要責備你，就是在你那裏有人服從了 巴蘭 的教訓；這 巴蘭 曾教唆 巴勒 將絆腳石放在 以色列 人面前，使他們吃祭過偶像之物，並且犯淫亂。
REV|2|15|同樣，你那裏也有人服從了 尼哥拉 派的教訓。
REV|2|16|所以，你當悔改；若不悔改，我很快就到你那裏來，用我口中的劍攻擊他們。
REV|2|17|凡有耳朵的都應當聽聖靈向眾教會所說的話。得勝的，我必將那隱藏的嗎哪賜給他，並賜他一塊白石，石上寫著新的名字，除了那領受的以外，沒有人認識。』」
REV|2|18|「你要寫信給 推雅推喇 教會的使者，說：『上帝的兒子，那位眼睛如火焰、雙腳像發亮的銅的這樣說：
REV|2|19|我知道你的行為：愛心、信心、勤勞、忍耐；又知道你末後所行的善事比起初所行的更多。
REV|2|20|然而，有一件事我要責備你，就是你容忍那自稱是先知的婦人 耶洗別 教唆我的僕人，引誘他們犯淫亂，吃祭過偶像之物。
REV|2|21|我曾給她悔改的機會，她卻不肯悔改她的淫行。
REV|2|22|看吧，我要使她病倒在床上。那些與她犯姦淫的人若不悔改他們的行為，我也要使他們同受大患難。
REV|2|23|我又要殺死她的兒女，眾教會就知道，我是那察看人肺腑心腸的，我要照你們的行為報應各人。
REV|2|24|至於你們其餘的 推雅推喇 人，就是一切不隨從這教訓，不明白他們所謂撒但深奧之理的人，我告訴你們，我不會再把別的擔子放在你們身上。
REV|2|25|你們只要持守那已經有的，直到我來。
REV|2|26|那得勝又遵守我命令到底的， 我要賜給他權柄制伏列國；
REV|2|27|他必用鐵杖管轄他們， 如同打碎陶器，
REV|2|28|像我也從我父領受了權柄一樣。我又要把晨星賜給他。
REV|2|29|凡有耳朵的都應當聽聖靈向眾教會所說的話。』」
REV|3|1|「你要寫信給 撒狄 教會的使者，說：『那有上帝的七靈和七顆星的這樣說：我知道你的行為，就是名義上你是活的，實際上你是死的。
REV|3|2|你要警醒，堅固那些剩下、快要死的，因為我發現你的行為，在我上帝面前沒有一樣是完全的。
REV|3|3|所以，要記得你所領受和聽見的；要遵守，並要悔改。你若不警醒，我必如賊一樣來到；我幾時來到你那裏，你絕不會知道。
REV|3|4|然而，在 撒狄 你還有幾位是未曾污穢自己衣服的，他們會穿白衣與我同行，因為他們是配穿的。
REV|3|5|得勝的必這樣穿白衣，我也不從生命冊上塗去他的名；我要在我父面前，和我父的眾使者面前，宣認他的名。
REV|3|6|凡有耳朵的都應當聽聖靈向眾教會所說的話。』」
REV|3|7|「你要寫信給 非拉鐵非 教會的使者，說： 『那神聖、真實的， 拿著 大衛 的鑰匙， 開了就沒有人能關， 關了就沒有人能開的這樣說：
REV|3|8|我知道你的行為。看哪，我在你面前給你一個敞開的門，是沒有人能關的。我知道你有一點力量，也遵守我的道，沒有否認我的名。
REV|3|9|那屬撒但會堂的，自稱是 猶太 人，其實不是 猶太 人，而是說謊話的，我要使他們來到你腳前下拜，使他們知道我已經愛你了。
REV|3|10|因為你遵守了我堅忍的道，我也必在普天下人受試煉的時候保守你免受試煉。
REV|3|11|我必快來，你要持守你所有的，免得人奪去你的冠冕。
REV|3|12|得勝的，我要使他在我上帝的殿中作柱子，他必不再從那裏出去。我又要把我上帝的名和我上帝城的名—從天上我上帝那裏降下來的新 耶路撒冷 ，和我的新名，都寫在他上面。
REV|3|13|凡有耳朵的都應當聽聖靈向眾教會所說的話。』」
REV|3|14|「你要寫信給 老底嘉 教會的使者，說：『那位阿們、誠信真實的見證者、上帝創造的根源這樣說：
REV|3|15|我知道你的行為，你也不冷也不熱；我巴不得你或冷或熱。
REV|3|16|既然你如溫水，也不冷也不熱，我要從我口中把你吐出去。
REV|3|17|你說：我是富足的，已經發了財，一樣都不缺，卻不知道你是困苦、可憐、貧窮、瞎眼、赤身的。
REV|3|18|我勸你向我買從火中鍛鍊出來的金子，使你富足；又買白衣穿上，使你赤身的羞恥不露出來；又買眼藥抹你的眼睛，使你能看見。
REV|3|19|凡我所疼愛的，我就責備管教。所以，你要發熱心，也要悔改。
REV|3|20|看哪，我站在門外叩門，若有聽見我聲音而開門的，我要進到他那裏去，我與他，他與我一起吃飯。
REV|3|21|得勝的，我要賜他在我寶座上與我同坐，就如我得了勝，在我父的寶座上與他同坐一般。
REV|3|22|凡有耳朵的都應當聽聖靈向眾教會所說的話。』」
REV|4|1|這些事以後，我觀看，看見天上有一道門開著。我頭一次聽見的那好像吹號的聲音對我說：「你上這裏來，我要把此後必須發生的事指示你。」
REV|4|2|我立刻被聖靈感動，見有一個寶座安置在天上，有一位坐在寶座上。
REV|4|3|那坐著的，看來好像碧玉和紅寶石；又有彩虹圍著寶座，光彩好像綠寶石。
REV|4|4|寶座的周圍又有二十四個座位，上面坐著二十四位長老，身穿白衣，頭上戴著金冠冕。
REV|4|5|有閃電、聲音、雷轟從寶座中發出。在寶座前點著七支火炬，就是上帝的七靈。
REV|4|6|寶座前有一個如同水晶的玻璃海。 寶座的周圍，四邊有四個活物，遍體前後都長滿了眼睛。
REV|4|7|第一個活物像獅子，第二個像牛犢，第三個的臉像人臉，第四個像飛鷹。
REV|4|8|四個活物各有六個翅膀，遍體內外都長滿了眼睛。他們晝夜不住地說： 「聖哉！聖哉！聖哉！ 主—全能的上帝； 昔在、今在、以後永在！」
REV|4|9|每逢四活物將榮耀、尊貴、感謝歸給那坐在寶座上、活到永永遠遠者的時候，
REV|4|10|二十四位長老就俯伏敬拜坐在寶座上活到永永遠遠的那一位，又把他們的冠冕放在寶座前，說：
REV|4|11|「我們的主，我們的上帝， 你配得榮耀、尊貴、權柄， 因為你創造了萬物， 萬物因你的旨意被創造而存在。」
REV|5|1|我看見坐在寶座那位的右手中有書卷，正反面都寫著字，用七個印密封著。
REV|5|2|我又看見一位大力的天使大聲宣告說：「有誰配展開那書卷，揭開那七個印呢？」
REV|5|3|在天上、地上、地底下，沒有人能展開、能閱覽那書卷。
REV|5|4|因為沒有人配展開、閱覽那書卷，我就大哭。
REV|5|5|長老中有一位對我說：「不要哭。看哪， 猶大 支派中的獅子， 大衛 的根，他已得勝，能展開那書卷，揭開那七個印。」
REV|5|6|我又看見寶座和四個活物，以及長老之中有羔羊站著，像是被殺的，有七個角七隻眼睛，就是上帝的七 靈，奉差遣往普天下去的。
REV|5|7|這羔羊前來，從坐在寶座上那位的右手中拿了書卷。
REV|5|8|他一拿了書卷，四活物和二十四位長老就俯伏在羔羊面前，各拿著琴和盛滿了香的金爐；這香就是眾聖徒的祈禱。
REV|5|9|他們唱新歌，說： 「你配拿書卷， 配揭開它的七印； 因為你曾被殺，用自己的血 從各支派、各語言、各民族、各邦國中買了人來，使他們歸於上帝，
REV|5|10|又使他們成為國民和祭司，歸於我們的上帝； 他們將在地上執掌王權。」
REV|5|11|我又觀看，我聽見寶座和活物及長老的周圍有許多天使的聲音；他們的數目有千千萬萬，
REV|5|12|大聲說： 「被殺的羔羊配得 權能、豐富、智慧、力量、 尊貴、榮耀、頌讚。
REV|5|13|我又聽見在天上、地上、地底下、滄海裏和天地間一切所有被造之物，都說： 「願頌讚、尊貴、榮耀、權勢， 都歸給坐在寶座上的那位和羔羊， 直到永永遠遠！」
REV|5|14|四活物就說：「阿們！」眾長老也俯伏敬拜。
REV|6|1|我看見羔羊揭開七個印中第一個印的時候，聽見四活物中的一個活物，聲音如雷，說：「你來！」
REV|6|2|我就觀看，看見一匹白馬，騎在馬上的拿著弓，並有冠冕賜給他。他出來征服，勝而又勝。
REV|6|3|羔羊揭開第二個印的時候，我聽見第二個活物說：「你來！」
REV|6|4|就另有一匹馬出來，是紅色的；有權柄賜給了那騎馬的，要從地上奪去太平，使人彼此相殺；他又接受了一把大刀。
REV|6|5|羔羊揭開第三個印的時候，我聽見第三個活物說：「你來！」我就觀看，看見一匹黑馬；騎在馬上的，手裏拿著天平。
REV|6|6|我聽見在四個活物中似乎有聲音說：「一個銀幣買一升麥子，一個銀幣買三升大麥；油和酒不可糟蹋。」
REV|6|7|羔羊揭開第四個印的時候，我聽見第四個活物說：「你來！」
REV|6|8|我就觀看，看見一匹灰色馬；騎在馬上的，名字叫作「死」，陰間也隨著他；有權柄賜給他們，可以用刀劍、饑荒、瘟疫、野獸，殺害地上四分之一的人。
REV|6|9|羔羊揭開第五個印的時候，我看見在祭壇底下有曾為上帝的道，並為作見證而被殺的人的靈魂，
REV|6|10|大聲喊著說：「神聖真實的主宰啊，你不審判住在地上的人，為我們所流的血伸冤，要到幾時呢？」
REV|6|11|於是有白袍賜給他們各人；又有話吩咐他們還要歇息片刻，等到與他們同作僕人的，和他們的弟兄，像他們一樣被殺的人的數目湊足的時候。
REV|6|12|羔羊揭開第六個印的時候，我看見地大震動，太陽變黑像粗麻布，整個月亮變紅像血，
REV|6|13|天上的星辰墜落在地上，如同無花果樹被大風搖動，落下未熟的果子一樣。
REV|6|14|天就裂開，好像書卷被捲起來；山嶺海島都被移動離開原位。
REV|6|15|地上的君王、臣宰、將軍、富戶、壯士，和一切為奴的、自主的，都藏在山洞和巖石穴裏，
REV|6|16|向山和巖石說：「倒在我們身上吧！把我們藏起來，躲避坐寶座者的臉面和羔羊的憤怒；
REV|6|17|因為他們遭憤怒的大日子到了，誰能站得住呢？」
REV|7|1|此後，我看見四位天使站在地的四角，執掌地上四方的風，使風不吹在地上、海上和各種樹上。
REV|7|2|我又看見另有一位天使從日出之地上來，拿著永生上帝的印。他向那得到權柄能傷害地和海的四位天使大聲喊著，
REV|7|3|說：「你們不可傷害地、海和樹林，等我們在我們上帝眾僕人的額上蓋了印。」
REV|7|4|我聽見 以色列 人各支派中受印的數目有十四萬四千；
REV|7|5|猶大 支派中受印的有一萬二千； 呂便 支派中有一萬二千； 迦得 支派中有一萬二千；
REV|7|6|亞設 支派中有一萬二千； 拿弗他利 支派中有一萬二千； 瑪拿西 支派中有一萬二千；
REV|7|7|西緬 支派中有一萬二千； 利未 支派中有一萬二千； 以薩迦 支派中有一萬二千；
REV|7|8|西布倫 支派中有一萬二千； 約瑟 支派中有一萬二千； 便雅憫 支派中受印的有一萬二千。
REV|7|9|此後，我觀看，看見有許多人，沒有人能計算，是從各邦國、各支派、各民族、各語言來的，站在寶座和羔羊面前，身穿白衣，手拿棕樹枝，
REV|7|10|大聲喊著說： 「願救恩歸於坐在寶座上我們的上帝， 也歸於羔羊！」
REV|7|11|眾天使都站在寶座和眾長老，以及四個活物的周圍，俯伏在寶座前，敬拜上帝，
REV|7|12|說： 「阿們！頌讚、榮耀、智慧、 感謝、尊貴、權能、 力量都歸於我們的上帝， 直到永永遠遠。阿們！」
REV|7|13|長老中有一位回應我說：「這些穿白衣的是誰？是從哪裏來的？」
REV|7|14|我對他說：「我主啊，你是知道的。」他向我說：「這些人是從大患難中出來的，他們曾用羔羊的血把衣裳洗得潔白。
REV|7|15|所以，他們在上帝寶座前， 晝夜在他殿中事奉他； 那坐在寶座上的要用帳幕覆庇他們。
REV|7|16|他們不再飢，不再渴； 太陽必不傷害他們， 任何炎熱也不傷害他們，
REV|7|17|因為寶座中的羔羊必牧養他們， 領他們到生命水的泉源； 上帝必擦去他們一切的眼淚。」
REV|8|1|羔羊揭開第七個印的時候，天上寂靜約有半小時。
REV|8|2|我看見那站在上帝面前的七位天使，有七枝號賜給他們。
REV|8|3|另有一位天使拿著金香爐來，站在祭壇旁邊；有許多香賜給他，要和眾聖徒的祈禱一同獻在寶座前的金壇上。
REV|8|4|那香的煙和眾聖徒的祈禱從天使的手中一同升到上帝面前。
REV|8|5|天使拿著香爐，盛滿了壇上的火，倒在地上；就有雷轟、響聲、閃電、地震。
REV|8|6|拿著七枝號筒的七位天使預備好要吹號。
REV|8|7|第一位天使吹號，就有冰雹和火攙著血扔在地上；地的三分之一和樹的三分之一被燒掉了，一切的青草也被燒掉了。
REV|8|8|第二位天使吹號，就有像火燒著的大山扔在海中；海的三分之一變成血，
REV|8|9|海中有生命的被造之物死了三分之一，船隻也毀壞了三分之一。
REV|8|10|第三位天使吹號，就有燒著的大星好像火把從天上墜下來，落在江河的三分之一和眾水的泉源上。
REV|8|11|這星名叫「苦艾」；眾水的三分之一變為苦艾，許多人因水變苦而死了。
REV|8|12|第四位天使吹號，太陽的三分之一、月亮的三分之一、星辰的三分之一都被擊打，以致日月星的三分之一變黑了，白晝的三分之一沒有光，黑夜也是這樣。
REV|8|13|我觀看，聽見一隻在空中飛的鷹大聲說：「禍哉！禍哉！禍哉！地上的居民哪，其餘的三位天使快要吹號了！」
REV|9|1|第五位天使吹號，我就看見一顆星從天上墜落到地上；有無底坑的鑰匙賜給它。
REV|9|2|它開了無底坑，就有煙從坑裏往上冒，好像大火爐的煙；太陽和天空都因這煙昏暗了。
REV|9|3|有蝗蟲從煙中出來，飛到地上，有權柄賜給牠們，好像地上的蠍子有權柄一樣。
REV|9|4|牠們奉命不可傷害地上的草、各樣綠色植物和各種樹木，惟獨可傷害額上沒有上帝印記的人；
REV|9|5|但是不許蝗蟲害死他們，只可使他們受痛苦五個月；這痛苦就像人被蠍子螫了的痛苦一樣。
REV|9|6|在那些日子，人求死，卻死不了；想死，死卻避開他們。
REV|9|7|蝗蟲的形狀好像預備上陣的戰馬一樣，頭上戴的好像金冠冕，臉面好像男人的臉面，
REV|9|8|頭髮像女人的頭髮，牙齒像獅子的牙齒；
REV|9|9|牠們胸前有甲，好像鐵甲；又有翅膀的響聲，好像許多車馬奔跑上陣的聲音。
REV|9|10|牠們有尾巴像蠍子，長著毒刺，尾巴上的毒刺有能力傷害人五個月。
REV|9|11|牠們有無底坑的使者作牠們的王，按著 希伯來 話名叫 亞巴頓 ， 希臘 話名話叫 亞玻倫 。
REV|9|12|第一樣災禍過去了；看哪，還有兩樣災禍要來。
REV|9|13|第六位天使吹號，我聽見有聲音從上帝面前金壇的四 角發出來，
REV|9|14|吩咐那吹號的第六位天使，說：「把那捆綁在 幼發拉底 大河的四個使者釋放了。」
REV|9|15|那四個使者就被釋放；他們原是預備好，在特定的年、月、日、時，要殺人類的三分之一。
REV|9|16|騎兵有二億；他們的數目我聽見了。
REV|9|17|我在異象中看見那些馬和騎馬的：騎馬的穿著火紅、紫瑪瑙及硫磺色的胸甲；馬的頭好像獅子的頭，有火、有煙、有硫磺從馬的口中噴出來。
REV|9|18|從馬的口中所噴出來的火、煙和硫磺這三樣災害殺了人類的三分之一。
REV|9|19|馬的能力在於牠們的口和尾巴；牠們的尾巴像蛇，有頭，用頭來傷害人。
REV|9|20|其餘未曾被這些災難所殺的人仍舊不為自己手所做的悔改，還是去拜鬼魔和那些不能看、不能聽、不能走，用金、銀、銅、木、石所造的偶像。
REV|9|21|他們也不為自己所犯的那些兇殺、邪術、淫亂、偷竊的事悔改。
REV|10|1|我又看見另一位大力的天使從天降下，披著雲彩，頭上有彩虹，臉面像太陽，兩腳像火柱。
REV|10|2|他手裏拿著展開的小書卷。他右腳踏海，左腳踏地，
REV|10|3|大聲呼喊，好像獅子吼叫。呼喊完了，就有七個雷發出聲音。
REV|10|4|七個雷發聲後，我正要寫出來，就聽見從天上有聲音說：「七個雷所說的，你要封上，不可寫出來。」
REV|10|5|我所看見的那踏海踏地的天使向天舉起右手，
REV|10|6|指著創造天和天上之物、地和地上之物、海和海中之物、直活到永永遠遠的那位起誓，說：「不再有時日了 。」
REV|10|7|但在第七位天使要吹號的日子，上帝的奧祕就要成全了，正如上帝向他僕人眾先知所宣告的。
REV|10|8|我先前從天上所聽見的那聲音又吩咐我說：「你去，把那踏海踏地之天使手中展開的小書卷拿過來。」
REV|10|9|我就走到天使那裏，對他說，請他把小書卷給我。他對我說：「你拿去，把它吃光。它會使你肚子發苦，然而在你口中會甘甜如蜜。」
REV|10|10|於是我從天使手中把小書卷接過來，把它吃光了，在我口中果然甘甜如蜜，吃了以後，我肚子覺得發苦。
REV|10|11|天使們對我說：「你必須指著許多民族、邦國、語言、君王再說預言。」
REV|11|1|有一根蘆葦，像丈量的杖，賜給我；且有話說：「起來！將上帝的殿和祭壇，以及在殿中禮拜的人，都量一量。
REV|11|2|只是殿外的院子不用量，因為這是要給外邦人的；他們將踐踏聖城四十二個月。
REV|11|3|「我要賜權柄給我那兩個見證人，穿著粗麻衣說預言一千二百六十天。」
REV|11|4|他們就是那站在世界之主面前的兩棵橄欖樹和兩個燈臺。
REV|11|5|若有人想要害他們，就有火從他們口中噴出來，燒滅仇敵；凡想要害他們的都必須這樣被殺。
REV|11|6|這二人有權柄關閉天空，使他們說預言的日子不下雨；又有權柄使水變為血，並且能隨時隨意用各樣的災害擊打大地世界。
REV|11|7|他們作完見證的時候，那從無底坑裏上來的獸要跟他們交戰，並且得勝，把他們殺了。
REV|11|8|他們的屍首將倒在大城的街道上；這城按著靈意叫 所多瑪 ，又叫 埃及 ，就是他們的主釘十字架的地方。
REV|11|9|從各民族、支派、語言、邦國中有人觀看他們的屍首三天半，又不許人把屍首安放在墳墓裏。
REV|11|10|住在地上的人會因他們而歡喜快樂，互相饋送禮物，因為這兩位先知曾使住在地上的人受痛苦。
REV|11|11|過了這三天半，有生命的氣息從上帝那裏進入他們裏面，他們就站起來；看見他們的人都大大懼怕。
REV|11|12|兩位先知聽見有大聲音從天上對他們說：「上這裏來。」他們就駕著雲上了天，他們的仇敵也看見了。
REV|11|13|正在那時候，地大震動，城倒塌了十分之一；因地震而死的有七千人，其餘的都恐懼，歸榮耀給天上的上帝。
REV|11|14|第二樣災禍過去了；看哪，第三樣災禍快到了。
REV|11|15|第七位天使吹號，天上就有大聲音說： 「世上的國已成了我們的主和他所立的基督的國了。 他要作王直到永永遠遠！」
REV|11|16|在上帝面前，坐在自己座位上的二十四位長老都俯伏在地上敬拜上帝，
REV|11|17|說： 「今在昔在的主—全能的上帝啊， 我們感謝你！ 因你執掌大權作王了。
REV|11|18|外邦發怒， 你的憤怒臨到了。 審判死人的時候也到了； 你的僕人眾先知、眾聖徒及敬畏你名的人， 連大帶小得賞賜的時候到了； 你毀滅那些毀滅大地者的時候也到了。」
REV|11|19|於是，上帝天上的聖所開了，在他聖所中，他的約櫃出現了；隨後有閃電、響聲、雷轟、地震、大冰雹。
REV|12|1|天上出現了一個大兆頭：有一個婦人身披太陽，腳踏月亮，頭戴十二顆星的冠冕；
REV|12|2|她懷了孕，在生產的陣痛中疼痛地喊叫。
REV|12|3|天上又出現了另一個兆頭：有一條大紅龍 ，有七個頭十個角；七個頭上戴著七個冠冕。
REV|12|4|牠的尾巴拖拉著天上星辰的三分之一，把它們摔在地上。然後龍站在那將要生產的婦人面前，等她生產後要吞吃她的孩子。
REV|12|5|婦人生了一個男孩子，就是將來要用鐵杖管轄 萬國的；她的孩子被提到上帝和他寶座那裏去。
REV|12|6|婦人就逃到曠野，在那裏有上帝給她預備的地方，使她在那裏被供養一千二百六十天。
REV|12|7|天上發生了爭戰。 米迦勒 同他的使者與龍作戰，龍同牠的使者也起來應戰，
REV|12|8|牠們都打敗了，天上再也沒有牠們的地方。
REV|12|9|大龍就是那古蛇，名叫魔鬼，又叫撒但，是迷惑普天下的；牠被摔在地上，牠的使者也一同被摔下去。
REV|12|10|我聽見在天上有大聲音說： 「我上帝的救恩、能力、國度， 和他所立的基督的權柄現在都來到了。 因為那個在我們上帝面前、 晝夜控告我們弟兄的， 已經被摔下去了。
REV|12|11|弟兄勝過那條龍是因羔羊的血， 和因自己所見證的道。 雖然至於死，他們也不惜自己的性命。
REV|12|12|所以，諸天和住在其中的， 你們都快樂吧！ 只是地和海有禍了！ 因為魔鬼知道自己的時候不多， 就氣憤憤地下到你們那裏去了。」
REV|12|13|龍見自己被摔在地上，就迫害那生男孩子的婦人。
REV|12|14|於是有大鷹的兩個翅膀賜給婦人，讓她能飛到曠野，到自己的地方，躲避那蛇。她在那裏受供養一載二載半載。
REV|12|15|蛇在婦人背後，從口中噴出水來，像河一樣，要將婦人沖走。
REV|12|16|地卻幫助了婦人，開口吞了從龍口噴出來的水。
REV|12|17|於是龍向婦人發怒，去與她其餘的兒女作戰，就是與那些遵守上帝命令 、為耶穌作見證的 。
REV|12|18|那時龍站在海邊沙灘上。
REV|13|1|我又看見一隻獸從海裏上來，有十個角七個頭；在十個角上戴著十個冠冕，七個頭上有褻瀆的名號。
REV|13|2|我所看見的獸，形狀像豹，腳像熊的腳，口像獅子的口。那條龍將自己的能力、座位和大權柄都給了牠。
REV|13|3|我看見獸的七個頭中，有一個似乎受了致命傷，那傷卻醫好了。全地的人都很驚訝，跟從了那隻獸。
REV|13|4|他們都拜那條龍，因為牠把自己的權柄給了獸；又拜那隻獸，說：「誰能比這隻獸，誰能與牠交戰呢？」
REV|13|5|龍又賜給那隻獸說誇大褻瀆話的口，又賜給牠權柄可以任意行事四十二個月。
REV|13|6|那獸就開口向上帝說褻瀆的話，褻瀆上帝的名和他的帳幕，就是那些住在天上的。
REV|13|7|牠又被准許與聖徒作戰，並且得勝，也賜給牠權柄，可以制伏各支派、各民族、各語言、各邦國。
REV|13|8|凡住在地上、名字從創世以來沒有記在被殺羔羊的生命冊上的人都要拜牠。
REV|13|9|凡有耳朵的都聽吧！
REV|13|10|該被擄掠的，必被擄掠； 該被刀殺的，必被刀殺。 在此，聖徒要有耐心和信心。
REV|13|11|我又看見另一隻獸從地裏上來。牠有兩個角如同羔羊，說話好像龍。
REV|13|12|牠在第一隻獸面前施行第一隻獸所有的權柄，並且使地和住在地上的人拜那致命傷被醫好了的第一隻獸。
REV|13|13|這隻獸又行大奇事，甚至在人面前使火從天降在地上。
REV|13|14|牠得了權柄在第一隻獸面前能行奇事，迷惑住在地上的人，告訴他們要為那受過刀傷還活著的獸造個像。
REV|13|15|又有權柄賜給牠，讓那隻獸的像有生氣，並且能說話，又使所有不拜獸像的人都被殺害。
REV|13|16|牠又使眾人，無論大小、貧富，自主的、為奴的，都在右手上，或是在額上，打一個印記；
REV|13|17|這樣，除了那有印記，有獸的名或有獸名數字的，都不得買或賣。
REV|13|18|在此，要有智慧：讓有悟性的人解開獸的數目吧，因為這是一個人的數字，那數字是六百六十六。
REV|14|1|我又觀看，看見羔羊站在 錫安山 ，和他在一起的有十四萬四千人，都有他的名和他父親的名寫在額上。
REV|14|2|我聽見從天上有聲音，像眾水的聲音和大雷的聲音，我所聽見的聲音好像琴師所彈的琴聲。
REV|14|3|他們在寶座前，和在四活物及眾長老前唱新歌，除了從地上買來的那十四萬四千人以外，沒有人能學這歌。
REV|14|4|這些人未曾沾染婦女，他們原是童身。羔羊無論往哪裏去，他們都跟隨他。他們是從人間買來的，作為初熟的果子歸給上帝和羔羊。
REV|14|5|在他們口中找不出謊言，他們是沒有瑕疵的。
REV|14|6|我又看見另一位天使在空中飛翔，有永遠的福音要傳給住在地上的人，就是各邦國、各支派、各語言、各民族。
REV|14|7|他大聲說：「要敬畏上帝，把榮耀歸給他，因為他施行審判的時候已經到了。要敬拜那創造天、地、海和水源的主。」
REV|14|8|另有第二位天使接著說：「傾覆了！那曾叫列國喝淫亂、烈怒之酒的大 巴比倫 傾覆了！」
REV|14|9|另有第三位天使接著他們，大聲說：「若有人拜那隻獸和獸像，在額上或在手上受了印記，
REV|14|10|他也必喝上帝烈怒的酒；這酒是斟在上帝憤怒的杯中的純酒。他要在聖天使和羔羊面前，在火與硫磺之中受痛苦。
REV|14|11|使他們受痛苦的煙往上冒，直到永永遠遠。那些拜獸和獸像，受了牠名字的印記的人，晝夜不得安寧。」
REV|14|12|在此，遵守上帝命令 和堅信耶穌真道的聖徒要有耐心。
REV|14|13|我聽見從天上有聲音說：「你要寫下：從今以後，在主裏死去的人有福了。」聖靈說：「是的，他們要從自己的勞苦中得安息，因為工作的成果永隨著他們。」
REV|14|14|我又觀看，看見有一片白雲，雲上坐著一位好像是人子的，頭上戴著金冠冕，手裏拿著鋒利的鐮刀。
REV|14|15|另有一位天使從聖所出來，向那坐在雲上的大聲喊著：「伸出你的鐮刀來收割吧，因為收割的時候已經到了，地上的莊稼已經熟透了。」
REV|14|16|於是那坐在雲上的把鐮刀向地上揮去，地上的莊稼就收割了。
REV|14|17|另有一位天使從天上的聖所出來，他也拿著鋒利的鐮刀。
REV|14|18|另有一位天使從祭壇出來，是有權柄管火的，向那拿著鋒利鐮刀的大聲喊著說：「伸出鋒利的鐮刀來，收取地上葡萄樹的果子，因為葡萄熟透了。」
REV|14|19|那天使就把鐮刀向地上揮去，收取了地上的葡萄，扔進上帝憤怒的大醡酒池裏。
REV|14|20|那醡酒池在城外被踹踏，有血從醡酒池裏流出來，漲到馬的嚼環那麼高，約有一千六百斯他迪 那麼遠。
REV|15|1|我看見在天上有另一兆頭，大而且奇，就是七位天使掌管末了的七種災難，因為上帝的烈怒在這七種災難中發盡了。
REV|15|2|我看見彷彿有攙雜火的玻璃海；又看見那些勝了那獸和獸像，以及牠名字的數字的人，都站在玻璃海上，拿著上帝的豎琴。
REV|15|3|他們唱上帝僕人 摩西 的歌和羔羊的歌，說： 「主—全能的上帝啊， 你的作為又偉大又奇妙！ 萬國之王啊， 你的道路又公義又真實！
REV|15|4|主啊，誰敢不敬畏你， 不把榮耀歸於你的名？ 因為只有你是神聖的。 萬民都要來， 在你面前敬拜， 因你公義的作為已經彰顯了。」
REV|15|5|此後，我看見在天上那存放法櫃的聖所開了。
REV|15|6|那掌管七種災難的七位天使從聖所出來，穿著潔白明亮的細麻衣 ，胸間束著金帶。
REV|15|7|四個活物中，有一個把盛滿了活到永永遠遠之上帝烈怒的七個金碗給了那七位天使。
REV|15|8|聖所中充滿了上帝的榮耀和權能而來的煙。沒有人能進入聖所，直等到那七位天使降完了七種災難。
REV|16|1|我聽見有大聲音從聖所裏出來，向那七位天使說：「你們去，把盛著上帝烈怒的七碗傾倒在地上。」
REV|16|2|第一位天使去，把碗傾倒在地上，就有又臭又毒的瘡生在那些有獸的印記和拜獸像的人身上。
REV|16|3|第二位天使把碗傾倒在海裏，海就變成像死人的血一樣，海裏所有的活物都死了。
REV|16|4|第三位天使把碗傾倒在河流和水源裏，水就變成血了。
REV|16|5|我聽見掌管眾水的天使說： 「昔在、今在的聖者啊， 你做的判斷公義；
REV|16|6|因他們曾流過聖徒與先知的血， 現在你給他們血喝， 這是他們該受的。」
REV|16|7|我又聽見祭壇中有聲音說： 「是的，主—全能的上帝啊， 你的判斷又真實又公義！」
REV|16|8|第四位天使把碗傾倒在太陽上，使太陽可用火烤人。
REV|16|9|人被炎熱所烤，就褻瀆那有權掌管這些災難的上帝的名，他們沒有悔改，也沒有把榮耀歸給上帝。
REV|16|10|第五位天使把碗傾倒在獸的座位上，獸的國就變成黑暗。人因疼痛而咬自己的舌頭；
REV|16|11|又因所受的疼痛和生的瘡，就褻瀆天上的上帝，也沒有為他們的行為悔改。
REV|16|12|第六位天使把碗傾倒在大 幼發拉底河 上，河水就乾了，為要給從日出之地所來的眾王預備道路。
REV|16|13|我又看見三個污穢的靈，好像青蛙，從龍的口、獸的口和假先知的口中出來。
REV|16|14|他們本是鬼魔的靈，施行奇事，到普天下眾王那裏去，召集他們在全能者上帝的大日子作戰。
REV|16|15|看哪，我來像賊一樣。那警醒、穿著衣服的人有福了；他不至於赤身而行，給人看見他的羞恥。
REV|16|16|於是，那三個鬼魔把眾王聚集在 希伯來 話叫作 哈米吉多頓 的地方。
REV|16|17|第七位天使把碗傾倒在空中，就有大聲音從聖所的寶座上出來，說：「成了！」
REV|16|18|又有閃電、響聲、雷轟、大地震，自從地上有人以來沒有這樣大、這樣厲害的地震。
REV|16|19|那大城裂為三段，列國的城也都倒塌了。上帝記起了大 巴比倫城 ，把那盛自己烈怒的酒杯遞給她。
REV|16|20|各海島都逃避了，眾山也不見了。
REV|16|21|又有大冰雹從天掉落在人身上，每一個約重一他連得，以致人因冰雹的災難而褻瀆上帝，因為那災難太大了。
REV|17|1|拿著七個碗的七位天使中，有一位前來對我說：「來，我要讓你看那坐在眾水之上的大淫婦所要受的懲罰；
REV|17|2|地上的君王都曾與她行淫，住在地上的人也喝醉了她淫亂的酒。」
REV|17|3|我在聖靈感動下，被天使帶到曠野去，我看見一個女人騎在朱紅色的獸上；那隻獸有七個頭十個角，遍體有褻瀆的名號。
REV|17|4|那女人穿著紫色和朱紅色的衣服，用金子、寶石、珍珠作妝飾，手拿著金杯，杯中盛滿了可憎之物和她淫亂的污穢。
REV|17|5|在她額上寫著奧祕的名字，說：「大 巴比倫 ，世上的淫婦和一切可憎之物的母。」
REV|17|6|我又看見那女人喝醉了聖徒的血和為耶穌作見證的人的血。 我看見她，非常詫異。
REV|17|7|天使對我說：「你為甚麼詫異呢？我要把這女人和馱著她那七頭十角的獸的奧祕告訴你。
REV|17|8|你曾看見的獸，以前有，現在沒有，將來要從無底坑裏上來，又歸於沉淪。凡住在地上、名字從創世以來沒有記在生命冊上的人看見那隻獸都要詫異，因為牠以前有，現在沒有，以後再有。
REV|17|9|在此要有智慧的心思：那七個頭就是女人所坐的七座山；他們又是七個王，
REV|17|10|五個已經倒了，一個還在，一個還沒有來到；他來的時候必須只暫時停留。
REV|17|11|那以前有、現在沒有的獸就是第八個，他也和那七個同列，正歸於沉淪。
REV|17|12|你曾看見的那十個角就是十個王；他們還沒有得到國度，但他們要和那隻獸同得權柄作王一個時辰。
REV|17|13|他們同心把自己的能力權柄交給那隻獸。
REV|17|14|他們將與羔羊作戰，羔羊必勝過他們，因為羔羊是萬主之主、萬王之王，而同羔羊在一起的是蒙召、被選、忠心的人。」
REV|17|15|天使又對我說：「你所看見那淫婦坐的眾水，就是許多民族、人民、邦國、語言。
REV|17|16|你所看見的那十個角與獸必恨這淫婦，他們要使她孤獨赤身，又要吃她的肉，用火將她燒盡。
REV|17|17|因為上帝使諸王同心執行他的旨意，把他們自己的國交給那隻獸，直等到上帝的話都應驗了。
REV|17|18|你所看見的那女人就是管轄地上眾王的大城。」
REV|18|1|此後，我看見另一位有大權柄的天使從天降下，地由於他的榮耀而發光。
REV|18|2|他以強而有力的聲音喊著說： 「傾覆了！大 巴比倫 傾覆了！ 她成了鬼魔的住處， 各樣污穢之靈的巢穴， 各樣污穢之鳥的窩， 各樣污穢可憎之獸的出沒處 。
REV|18|3|因為列國都喝了她淫亂大怒的酒 ； 地上的君王和她行淫； 地上的商人因她極度奢華而發了財。」
REV|18|4|我又聽見另一個聲音從天上說： 「我的民哪，從那城出來吧！ 免得和她在罪上有份， 受她所受的災殃；
REV|18|5|因她的罪惡滔天， 上帝已經記得她的不義。
REV|18|6|她怎樣待人，也要怎樣待她， 按她所行的加倍地報應她； 用她調酒的杯加倍調給她喝。
REV|18|7|她怎樣榮耀自己，怎樣奢華， 也要使她照樣痛苦悲哀。 因她心裏說： 『我坐了皇后的位， 並不是寡婦， 絕不至於悲哀。』
REV|18|8|所以在一天之內，她的災殃要一齊來到， 就是死亡、悲哀、饑荒。 她將被火燒盡， 因為審判她的主上帝大有能力。」
REV|18|9|地上的君王，與她行淫、一同奢華的，看見燒她的煙，就必為她哭泣哀號；
REV|18|10|因怕她的痛苦，就遠遠地站著，說： 「禍哉，禍哉，這大城！ 堅固的 巴比倫城 啊！ 一時之間，你的審判要來到了。」
REV|18|11|地上的商人也都為她哭泣悲哀，因為沒有人再買他們的貨物了；
REV|18|12|這貨物就是金、銀、寶石、珍珠、細麻布、絲綢、紫色和朱紅色衣料、各樣香木、各樣象牙的器皿、各樣極寶貴的木頭和銅、鐵、大理石的器皿，
REV|18|13|和肉桂、豆蔻、香料、香膏、乳香、酒、油、細麵、麥子、牛、羊、馬、馬車，以及奴隸、人口。
REV|18|14|「你所貪愛的果子離開了你； 你一切的珍饈美味和華美的物件 都從你那裏毀滅， 絕對見不到了。」
REV|18|15|販賣這些貨物、藉著她發財的商人，因怕她的痛苦，就遠遠地站著哭泣悲哀，
REV|18|16|說： 「禍哉，禍哉，這大城！ 她穿著細麻、 紫色、朱紅色的衣服， 用金子、寶石、珍珠為妝飾。
REV|18|17|一時之間，這麼多的財富就歸於無有了。」 所有的船長和到處航海的，水手以及所有靠海為業的，都遠遠地站著，
REV|18|18|看見燒她的煙，就喊著說：「有哪一個城能跟這大城比呢？」
REV|18|19|於是他們把灰塵撒在頭上，哭泣悲哀地喊著說： 「禍哉，禍哉，這大城！ 凡有船在海中的， 都因她的珍寶成了富足。 她在一時之間就成為荒蕪。
REV|18|20|天哪，眾聖徒、眾使徒、眾先知啊！ 你們都要因她歡喜， 因為上帝已經在她身上為你們伸了冤。」
REV|18|21|有一位大力的天使舉起一塊石頭，好像大磨石，扔在海裏，說： 「 巴比倫 大城 也必這樣猛力地被扔下去， 絕對見不到了。
REV|18|22|彈琴、歌唱、 吹笛、吹號的聲音， 在你中間絕對聽不見了； 各行手藝的技工 在你中間絕對見不到了； 推磨的聲音 在你中間絕對聽不見了；
REV|18|23|燈臺的光 在你中間絕對不再照耀了； 新郎和新娘的聲音 在你中間絕對聽不見了。 你的商人原來是地上的顯要； 萬國也被你的邪術迷惑了。
REV|18|24|先知、聖徒和地上一切被殺的人的血都在這城裏找到了。」
REV|19|1|此後，我聽見好像有一大群人在天上大聲說： 「哈利路亞 ！ 救恩、榮耀、權能都屬於我們的上帝。
REV|19|2|他的判斷又真實又公義； 因他判斷了那大淫婦， 她用淫行敗壞了世界。 上帝為他的僕人伸冤， 向淫婦討流僕人血的罪。」
REV|19|3|他們又一次說： 「哈利路亞！ 燒淫婦的煙往上冒，直到永永遠遠。」
REV|19|4|那二十四位長老和四活物就俯伏敬拜坐在寶座上的上帝，說： 「阿們。哈利路亞！」
REV|19|5|接著，有聲音從寶座出來說： 「上帝的眾僕人哪， 凡敬畏他的， 無論大小， 都要讚美我們的上帝！」
REV|19|6|我聽見好像一大群人的聲音，像眾水的聲音，像大雷的聲音，說： 「哈利路亞！ 因為主─我們的上帝 、 全能者，作王了。
REV|19|7|我們要歡喜快樂， 將榮耀歸給他； 因為羔羊的婚期到了， 他的新娘也自己預備好了，
REV|19|8|她蒙恩得穿明亮潔白的細麻衣： 這細麻衣就是聖徒們的義行。」
REV|19|9|天使對我說：「你要寫下來：凡被請赴羔羊婚宴的人有福了！」他又對我說：「這些都是上帝真實的話。」
REV|19|10|我就俯伏在他腳前要拜他。他對我說：「千萬不可！我和你，以及那些為耶穌作見證的弟兄同是僕人。你要敬拜上帝。」因為那些為耶穌作見證的人有預言的靈。
REV|19|11|後來我看見天開了。有一匹白馬，騎在馬上的稱為 「誠信」、「真實」，他審判和爭戰都憑著公義。
REV|19|12|他的眼睛如 火焰，頭上戴著許多冠冕；他身上寫著一個名字，除了他自己沒有人知道。
REV|19|13|他穿著浸過血的衣服；他的名稱為「上帝之道」。
REV|19|14|眾天軍都騎著白馬，穿著又白又潔淨的細麻衣跟隨他。
REV|19|15|有利劍從他口中出來，用來擊打列國。他要用鐵杖管轄 他們，並且要踹全能上帝烈怒的醡酒池。
REV|19|16|在他衣服和大腿上寫著「萬王之王，萬主之主」的名號。
REV|19|17|我又看見一位天使站在太陽中，向天空一切的飛鳥大聲喊著說：「你們聚集來赴上帝的大宴席，
REV|19|18|為要吃君王的肉、將軍的肉、壯士的肉、馬和騎士的肉、一切自主的和為奴的，以及尊貴的和卑賤的肉。」
REV|19|19|我又看見那獸和地上的君王，和他們的軍隊都聚集，要與白馬騎士和他的軍隊作戰。
REV|19|20|那獸被擒拿了；那在獸面前曾行奇事、迷惑了接受獸的印記和拜獸像的人的假先知，也與獸同被擒拿。他們兩個就活生生地被扔進燒著硫磺的火湖裏，
REV|19|21|其餘的人被白馬騎士口中吐出來的劍殺了；所有的飛鳥都吃飽了他們的肉。
REV|20|1|我又看見一位天使從天降下，手裏拿著無底坑的鑰匙和一條大鐵鏈。
REV|20|2|他抓住那龍，那古蛇，就是魔鬼、撒但，把牠捆綁了一千年，
REV|20|3|扔在無底坑裏，把無底坑關閉，用印封上，使牠不再迷惑列國，等到那一千年滿了。這些事以後，牠必須暫時被釋放。
REV|20|4|我又看見一些寶座，坐在上面的有審判的權柄賜給他們。我又看見那些因為給耶穌作見證，並為上帝之道被斬首的人的靈魂，和沒有拜過那獸與獸像、也沒有在額上和手上打過牠印記的人的靈魂。他們都復活了，與基督一同作王一千年。
REV|20|5|這是頭一次的復活。其餘的死人還沒有復活，直等那一千年滿了。
REV|20|6|在頭一次復活有份的有福了，聖潔了！第二次的死在他們身上沒有權柄，但他們要作上帝和基督的祭司，也要與基督一同作王一千年。
REV|20|7|那一千年滿了，撒但會從監牢裏被釋放，
REV|20|8|出來要迷惑地上四方的列國，就是 歌革 和 瑪各 ，使他們聚集爭戰。他們的人數多如海沙。
REV|20|9|他們上來佈滿了全地，圍住聖徒的營與蒙愛的城，就有火從天降下，燒滅了他們。
REV|20|10|那迷惑他們的魔鬼被扔進硫磺的火湖裏，就是那獸和假先知所在的地方，他們會晝夜受折磨，直到永永遠遠。
REV|20|11|我又看見一個白色的大寶座和那坐在上面的；天和地都從他面前逃避，再也找不到它們的位置了。
REV|20|12|我又看見死了的人，無論大小，都站在寶座前。案卷都展開了，並另有一卷展開，就是生命冊。死了的人都憑著這些案卷所記載的，照他們所行的受審判。
REV|20|13|於是海交出其中的死人，死亡和陰間也交出其中的死人；他們都照各人所行的受審判。
REV|20|14|死亡和陰間也被扔進火湖裏，這火湖就是第二次的死。
REV|20|15|凡名字沒有記在生命冊上的人，就被扔進火湖裏。
REV|21|1|我又看見一個新天新地，因為先前的天和先前的地已經過去了，海也不再有了。
REV|21|2|我又看見聖城，新 耶路撒冷 由上帝那裏，從天而降，預備好了，就如新娘打扮整齊，等候丈夫。
REV|21|3|我聽見有大聲音從寶座出來，說： 「看哪，上帝的帳幕在人間！ 他要和他們同住， 他們要作他的子民。 上帝要親自與他們同在。
REV|21|4|上帝要擦去他們一切的眼淚； 不再有死亡， 也不再有悲哀、哭號、痛苦， 因為先前的事都過去了。」
REV|21|5|那位坐在寶座上的說：「看哪，我把一切都更新了！」他又說：「你要寫下來，因為這些話是可信靠的，是真實的。」
REV|21|6|他又對我說：「成了！我是阿拉法，我是俄梅戛；我是開始，我是終結。我要把生命的泉水白白賜給那口渴的人喝。
REV|21|7|得勝的要承受這些為業；我要作他的上帝，他要作我的兒子。
REV|21|8|至於膽怯的、不信的、可憎的、殺人的、淫亂的、行邪術的、拜偶像的和一切說謊話的人，他們將在燒著硫磺的火湖裏有份；這是第二次的死。」
REV|21|9|拿著七個金碗、盛滿末後七種災禍的七位天使中，有一位來對我說：「你來，我要給你看新娘，就是羔羊的妻子。」
REV|21|10|我在聖靈感動下，天使帶我到一座高大的山，給我看由上帝那裏、從天而降的聖城 耶路撒冷 ，
REV|21|11|這城有上帝的榮耀，它光輝如同極貴的寶石，好像碧玉，明如水晶。
REV|21|12|它有高大的牆，有十二個門，門上有十二位天使，門上又寫著 以色列 人十二個支派的名字 。
REV|21|13|東邊有三個門，北邊有三個門，南邊有三個門，西邊有三個門。
REV|21|14|城牆有十二個根基，根基上有羔羊十二使徒的名字。
REV|21|15|那對我說話的天使拿著金的蘆葦當尺，要量那城、城門和城牆。
REV|21|16|城是四方的，長寬一樣。天使用蘆葦量那城，共有一萬二千斯他迪，長、寬、高都是一樣。
REV|21|17|他又量了城牆，按著人的尺寸，就是天使的尺寸，共有一百四十四肘。
REV|21|18|牆是碧玉造的；城是純金的，如同明淨的玻璃。
REV|21|19|城牆的根基是用各樣寶石修飾的：第一個根基是碧玉，第二是藍寶石，第三是綠瑪瑙，第四是綠寶石，
REV|21|20|第五是紅瑪瑙，第六是紅寶石，第七是黃璧璽，第八是水蒼玉，第九是紅璧璽，第十是翡翠，第十一是紫瑪瑙，第十二是紫晶。
REV|21|21|十二個門是十二顆珍珠；每一個門是一顆珍珠造的。城內的街道是純金的，好像透明的玻璃。
REV|21|22|我沒有看見城內有殿，因主—全能者上帝和羔羊就是城的殿。
REV|21|23|那城內不用日月光照，因為有上帝的榮耀光照，又有羔羊為城的燈。
REV|21|24|列國要藉著城的光行走；地上的君王要把自己的榮耀帶給那城。
REV|21|25|城門白晝總不關閉，在那裏沒有黑夜。
REV|21|26|人要將列國的榮耀尊貴帶給那城。
REV|21|27|凡不潔淨的，和那行可憎與虛謊之事的人，都不得進那城，只有名字寫在羔羊生命冊上的才得進去。
REV|22|1|天使又讓我看一道生命水的河，明亮如水晶，從上帝和羔羊的寶座流出來，
REV|22|2|經過城內街道的中央；在河的兩邊有生命樹，結十二樣 的果子，每月都結果子；樹上的葉子可作醫治萬民之用。
REV|22|3|以後不再有任何詛咒。在城裏將有上帝和羔羊的寶座。他的僕人都要事奉他，
REV|22|4|也要見他的面。他的名字將寫在他們的額上。
REV|22|5|不再有黑夜；他們也不需要燈光或日光，因為主上帝要光照他們。他們要作王，直到永永遠遠。
REV|22|6|天使又對我說：「這些話是可信靠的，是真實的。主，就是賜靈感給眾先知的上帝，差遣他的使者，要將必須快要發生的事指示他的眾僕人。」
REV|22|7|「看哪，我必快來！凡遵守這書上預言的有福了。」
REV|22|8|這些事是我－ 約翰 所聽見所看見的。當我聽見看見時，就俯伏在指示我的天使腳前要拜他。
REV|22|9|他對我說：「千萬不可！我與你和你的弟兄眾先知，以及那些守這書上的話的人，同是作僕人。你要敬拜上帝。」
REV|22|10|他又對我說：「不可封了這書上的預言，因為時候近了。
REV|22|11|不義的，讓他仍舊不義；污穢的，讓他仍舊污穢；為義的，讓他仍舊為義；聖潔的，讓他仍舊聖潔。」
REV|22|12|「看哪，我必快來！賞罰在我，要照每個人所行的報應他。
REV|22|13|我是阿拉法，我是俄梅戛；我是首先的，我是末後的；我是開始，我是終結。」
REV|22|14|那些洗淨自己衣服的有福了！他們可得權柄到生命樹那裏，也能從門進城。
REV|22|15|城外有犬類、行邪術的、淫亂的、殺人的、拜偶像的，以及所有喜愛和行虛謊的人。
REV|22|16|「我－耶穌差遣我的使者，為了眾教會向你們證明這些事。我是 大衛 的根，是他的後裔；我是明亮的晨星。」
REV|22|17|聖靈和新娘都說：「來！」聽見的人也要說：「來！」口渴的人也要來，願意的人都可以白白取生命的水喝。
REV|22|18|我警告一切聽見這書上預言的人：若有人在這預言上加添甚麼，上帝必將記在這書上的災禍加在他身上。
REV|22|19|這書上的預言，若有人刪去甚麼，上帝必從這書上所記的生命樹和聖城刪去他的份。
REV|22|20|證明這些事的說：「是的，我必快來！」阿們！主耶穌啊，我願你來！
REV|22|21|願主耶穌的恩惠與眾聖徒同在。阿們！
