REV|1|1|耶穌基督的啟示，就是上帝賜給他，要他將必須快要發生的事指示他的眾僕人。他差遣使者指明給他的僕人 約翰 ，
REV|1|2|約翰 就將上帝的道和耶穌基督的見證，凡自己所看見的，都見證出來。
REV|1|3|誦讀這書上預言的，和那些聽見又遵守其中所記載的，都是有福的，因為時候近了。
REV|1|4|約翰 寫信給 亞細亞 的七個教會。願那位今在、昔在、以後永在的上帝，與他寶座前的七靈，和那忠信的見證者、從死人中復活的首生者 、世上君王的元首耶穌基督，賜恩惠和平安 給你們。 他愛我們，用自己的血使我們從罪中得釋放 ，
REV|1|5|
REV|1|6|又使我們成為國度，作他父上帝的祭司。願榮耀、權能歸給他，直到永永遠遠 。阿們！
REV|1|7|「看哪，他駕雲降臨； 眾目都要看見他， 連刺他的人也要看見他； 地上的萬族要因他哀哭。」 這是真實的。阿們！
REV|1|8|主上帝說：「我是阿拉法，我是俄梅戛 ，是今在、昔在、以後永在的全能者。」
REV|1|9|我— 約翰 就是你們的弟兄，在耶穌裏和你們一同在患難、國度、忍耐裏有份的，為上帝的道，並為給耶穌作的見證，曾在那名叫 拔摩 的海島上。
REV|1|10|有一主日我被聖靈感動，聽見在我後面有大聲音如吹號，
REV|1|11|說：「把你所看見的寫在書上，寄給 以弗所 、 士每拿 、 別迦摩 、 推雅推喇 、 撒狄 、 非拉鐵非 、 老底嘉 那七個教會。」
REV|1|12|我轉過身來要看看是誰的聲音在跟我說話。我一轉過來，看見了七個金燈臺；
REV|1|13|在燈臺中間有一位好像人子的，身穿垂到腳的長袍，胸間束著金帶。
REV|1|14|他的頭與髮皆白，如白羊毛，如雪；他的眼睛好像火焰，
REV|1|15|雙腳好像在爐中鍛鍊得發亮的銅，聲音好像眾水的聲音。
REV|1|16|他右手拿著七顆星，從他口中吐出一把兩刃的利劍，面貌好像烈日放光。
REV|1|17|我看見了他，就仆倒在他腳前，像死人一樣。他用右手按著我說：「不要怕。我是首先的，是末後的，
REV|1|18|又是永活的。我曾死過，看哪，我是活著的，直到永永遠遠；並且我拿著死亡和陰間的鑰匙。
REV|1|19|所以，你要把所看見的事、現在的事和以後將發生的事，都寫下來。
REV|1|20|至於你所看見、在我右手中的七顆星和那七個金燈臺的奧祕就是：七顆星是七個教會的使者，七個燈臺是七個教會。」
REV|2|1|「你要寫信給 以弗所 教會的使者，說：『那右手拿著七顆星，在七個金燈臺中間行走的這樣說：
REV|2|2|我知道你的行為、勞碌、忍耐，也知道你不容忍惡人。你也曾察驗那自稱為使徒卻不是使徒的，看出他們是假的。
REV|2|3|你能忍耐，曾為我的名勞苦而不困倦。
REV|2|4|然而，有一件事我要責備你，就是你把起初的愛心拋棄了。
REV|2|5|所以你要回想你是從哪裏墜落的，並且要悔改，做起初所做的工作。你若不悔改，我要到你那裏去，把你的燈臺從原處挪去。
REV|2|6|然而你還有一件可取的事，就是你恨惡 尼哥拉 派的行為，這種行為也是我所恨惡的。
REV|2|7|凡有耳朵的都應當聽聖靈向眾教會所說的話。得勝的，我必將上帝樂園中生命樹的果子賜給他吃。』」
REV|2|8|「你要寫信給 士每拿 教會的使者，說：『那首先的、末後的，死過又活了的這樣說：
REV|2|9|我知道你的患難和貧窮—其實你卻是富足的，也知道那自稱是 猶太 人的所說毀謗的話，其實他們不是 猶太 人，而是撒但會堂的人。
REV|2|10|你將要受的苦，你不用怕。看哪！魔鬼要把你們中間幾個人下在監裏，使你們受考驗，你們要遭受苦難十日。你務要至死忠心，我就賜給你那生命的冠冕。
REV|2|11|凡有耳朵的都應當聽聖靈向眾教會所說的話。得勝的必不受第二次死的害。』」
REV|2|12|「你要寫信給 別迦摩 教會的使者，說：『那有兩刃利劍的這樣說：
REV|2|13|我知道你的居所，就是有撒但座位之處；當我忠心的見證人 安提帕 在你們中間，在撒但所住的地方被殺之時，你還堅守我的名，沒有否認對我的信仰。
REV|2|14|然而，有幾件事我要責備你，就是在你那裏有人服從了 巴蘭 的教訓；這 巴蘭 曾教唆 巴勒 將絆腳石放在 以色列 人面前，使他們吃祭過偶像之物，並且犯淫亂。
REV|2|15|同樣，你那裏也有人服從了 尼哥拉 派的教訓。
REV|2|16|所以，你當悔改；若不悔改，我很快就到你那裏來，用我口中的劍攻擊他們。
REV|2|17|凡有耳朵的都應當聽聖靈向眾教會所說的話。得勝的，我必將那隱藏的嗎哪賜給他，並賜他一塊白石，石上寫著新的名字，除了那領受的以外，沒有人認識。』」
REV|2|18|「你要寫信給 推雅推喇 教會的使者，說：『上帝的兒子，那位眼睛如火焰、雙腳像發亮的銅的這樣說：
REV|2|19|我知道你的行為：愛心、信心、勤勞、忍耐；又知道你末後所行的善事比起初所行的更多。
REV|2|20|然而，有一件事我要責備你，就是你容忍那自稱是先知的婦人 耶洗別 教唆我的僕人，引誘他們犯淫亂，吃祭過偶像之物。
REV|2|21|我曾給她悔改的機會，她卻不肯悔改她的淫行。
REV|2|22|看吧，我要使她病倒在床上。那些與她犯姦淫的人若不悔改他們的行為，我也要使他們同受大患難。
REV|2|23|我又要殺死她的兒女，眾教會就知道，我是那察看人肺腑心腸的，我要照你們的行為報應各人。
REV|2|24|至於你們其餘的 推雅推喇 人，就是一切不隨從這教訓，不明白他們所謂撒但深奧之理的人，我告訴你們，我不會再把別的擔子放在你們身上。
REV|2|25|你們只要持守那已經有的，直到我來。
REV|2|26|那得勝又遵守我命令到底的， 我要賜給他權柄制伏列國；
REV|2|27|他必用鐵杖管轄他們， 如同打碎陶器，
REV|2|28|像我也從我父領受了權柄一樣。我又要把晨星賜給他。
REV|2|29|凡有耳朵的都應當聽聖靈向眾教會所說的話。』」
REV|3|1|「你要寫信給 撒狄 教會的使者，說：『那有上帝的七靈和七顆星的這樣說：我知道你的行為，就是名義上你是活的，實際上你是死的。
REV|3|2|你要警醒，堅固那些剩下、快要死的，因為我發現你的行為，在我上帝面前沒有一樣是完全的。
REV|3|3|所以，要記得你所領受和聽見的；要遵守，並要悔改。你若不警醒，我必如賊一樣來到；我幾時來到你那裏，你絕不會知道。
REV|3|4|然而，在 撒狄 你還有幾位是未曾污穢自己衣服的，他們會穿白衣與我同行，因為他們是配穿的。
REV|3|5|得勝的必這樣穿白衣，我也不從生命冊上塗去他的名；我要在我父面前，和我父的眾使者面前，宣認他的名。
REV|3|6|凡有耳朵的都應當聽聖靈向眾教會所說的話。』」
REV|3|7|「你要寫信給 非拉鐵非 教會的使者，說： 『那神聖、真實的， 拿著 大衛 的鑰匙， 開了就沒有人能關， 關了就沒有人能開的這樣說：
REV|3|8|我知道你的行為。看哪，我在你面前給你一個敞開的門，是沒有人能關的。我知道你有一點力量，也遵守我的道，沒有否認我的名。
REV|3|9|那屬撒但會堂的，自稱是 猶太 人，其實不是 猶太 人，而是說謊話的，我要使他們來到你腳前下拜，使他們知道我已經愛你了。
REV|3|10|因為你遵守了我堅忍的道，我也必在普天下人受試煉的時候保守你免受試煉。
REV|3|11|我必快來，你要持守你所有的，免得人奪去你的冠冕。
REV|3|12|得勝的，我要使他在我上帝的殿中作柱子，他必不再從那裏出去。我又要把我上帝的名和我上帝城的名—從天上我上帝那裏降下來的新 耶路撒冷 ，和我的新名，都寫在他上面。
REV|3|13|凡有耳朵的都應當聽聖靈向眾教會所說的話。』」
REV|3|14|「你要寫信給 老底嘉 教會的使者，說：『那位阿們、誠信真實的見證者、上帝創造的根源這樣說：
REV|3|15|我知道你的行為，你也不冷也不熱；我巴不得你或冷或熱。
REV|3|16|既然你如溫水，也不冷也不熱，我要從我口中把你吐出去。
REV|3|17|你說：我是富足的，已經發了財，一樣都不缺，卻不知道你是困苦、可憐、貧窮、瞎眼、赤身的。
REV|3|18|我勸你向我買從火中鍛鍊出來的金子，使你富足；又買白衣穿上，使你赤身的羞恥不露出來；又買眼藥抹你的眼睛，使你能看見。
REV|3|19|凡我所疼愛的，我就責備管教。所以，你要發熱心，也要悔改。
REV|3|20|看哪，我站在門外叩門，若有聽見我聲音而開門的，我要進到他那裏去，我與他，他與我一起吃飯。
REV|3|21|得勝的，我要賜他在我寶座上與我同坐，就如我得了勝，在我父的寶座上與他同坐一般。
REV|3|22|凡有耳朵的都應當聽聖靈向眾教會所說的話。』」
REV|4|1|這些事以後，我觀看，看見天上有一道門開著。我頭一次聽見的那好像吹號的聲音對我說：「你上這裏來，我要把此後必須發生的事指示你。」
REV|4|2|我立刻被聖靈感動，見有一個寶座安置在天上，有一位坐在寶座上。
REV|4|3|那坐著的，看來好像碧玉和紅寶石；又有彩虹圍著寶座，光彩好像綠寶石。
REV|4|4|寶座的周圍又有二十四個座位，上面坐著二十四位長老，身穿白衣，頭上戴著金冠冕。
REV|4|5|有閃電、聲音、雷轟從寶座中發出。在寶座前點著七支火炬，就是上帝的七靈。
REV|4|6|寶座前有一個如同水晶的玻璃海。 寶座的周圍，四邊有四個活物，遍體前後都長滿了眼睛。
REV|4|7|第一個活物像獅子，第二個像牛犢，第三個的臉像人臉，第四個像飛鷹。
REV|4|8|四個活物各有六個翅膀，遍體內外都長滿了眼睛。他們晝夜不住地說： 「聖哉！聖哉！聖哉！ 主—全能的上帝； 昔在、今在、以後永在！」
REV|4|9|每逢四活物將榮耀、尊貴、感謝歸給那坐在寶座上、活到永永遠遠者的時候，
REV|4|10|二十四位長老就俯伏敬拜坐在寶座上活到永永遠遠的那一位，又把他們的冠冕放在寶座前，說：
REV|4|11|「我們的主，我們的上帝， 你配得榮耀、尊貴、權柄， 因為你創造了萬物， 萬物因你的旨意被創造而存在。」
REV|5|1|我看見坐在寶座那位的右手中有書卷，正反面都寫著字，用七個印密封著。
REV|5|2|我又看見一位大力的天使大聲宣告說：「有誰配展開那書卷，揭開那七個印呢？」
REV|5|3|在天上、地上、地底下，沒有人能展開、能閱覽那書卷。
REV|5|4|因為沒有人配展開、閱覽那書卷，我就大哭。
REV|5|5|長老中有一位對我說：「不要哭。看哪， 猶大 支派中的獅子， 大衛 的根，他已得勝，能展開那書卷，揭開那七個印。」
REV|5|6|我又看見寶座和四個活物，以及長老之中有羔羊站著，像是被殺的，有七個角七隻眼睛，就是上帝的七 靈，奉差遣往普天下去的。
REV|5|7|這羔羊前來，從坐在寶座上那位的右手中拿了書卷。
REV|5|8|他一拿了書卷，四活物和二十四位長老就俯伏在羔羊面前，各拿著琴和盛滿了香的金爐；這香就是眾聖徒的祈禱。
REV|5|9|他們唱新歌，說： 「你配拿書卷， 配揭開它的七印； 因為你曾被殺，用自己的血 從各支派、各語言、各民族、各邦國中買了人來，使他們歸於上帝，
REV|5|10|又使他們成為國民和祭司，歸於我們的上帝； 他們將在地上執掌王權。」
REV|5|11|我又觀看，我聽見寶座和活物及長老的周圍有許多天使的聲音；他們的數目有千千萬萬，
REV|5|12|大聲說： 「被殺的羔羊配得 權能、豐富、智慧、力量、 尊貴、榮耀、頌讚。
REV|5|13|我又聽見在天上、地上、地底下、滄海裏和天地間一切所有被造之物，都說： 「願頌讚、尊貴、榮耀、權勢， 都歸給坐在寶座上的那位和羔羊， 直到永永遠遠！」
REV|5|14|四活物就說：「阿們！」眾長老也俯伏敬拜。
REV|6|1|我看見羔羊揭開七個印中第一個印的時候，聽見四活物中的一個活物，聲音如雷，說：「你來！」
REV|6|2|我就觀看，看見一匹白馬，騎在馬上的拿著弓，並有冠冕賜給他。他出來征服，勝而又勝。
REV|6|3|羔羊揭開第二個印的時候，我聽見第二個活物說：「你來！」
REV|6|4|就另有一匹馬出來，是紅色的；有權柄賜給了那騎馬的，要從地上奪去太平，使人彼此相殺；他又接受了一把大刀。
REV|6|5|羔羊揭開第三個印的時候，我聽見第三個活物說：「你來！」我就觀看，看見一匹黑馬；騎在馬上的，手裏拿著天平。
REV|6|6|我聽見在四個活物中似乎有聲音說：「一個銀幣買一升麥子，一個銀幣買三升大麥；油和酒不可糟蹋。」
REV|6|7|羔羊揭開第四個印的時候，我聽見第四個活物說：「你來！」
REV|6|8|我就觀看，看見一匹灰色馬；騎在馬上的，名字叫作「死」，陰間也隨著他；有權柄賜給他們，可以用刀劍、饑荒、瘟疫、野獸，殺害地上四分之一的人。
REV|6|9|羔羊揭開第五個印的時候，我看見在祭壇底下有曾為上帝的道，並為作見證而被殺的人的靈魂，
REV|6|10|大聲喊著說：「神聖真實的主宰啊，你不審判住在地上的人，為我們所流的血伸冤，要到幾時呢？」
REV|6|11|於是有白袍賜給他們各人；又有話吩咐他們還要歇息片刻，等到與他們同作僕人的，和他們的弟兄，像他們一樣被殺的人的數目湊足的時候。
REV|6|12|羔羊揭開第六個印的時候，我看見地大震動，太陽變黑像粗麻布，整個月亮變紅像血，
REV|6|13|天上的星辰墜落在地上，如同無花果樹被大風搖動，落下未熟的果子一樣。
REV|6|14|天就裂開，好像書卷被捲起來；山嶺海島都被移動離開原位。
REV|6|15|地上的君王、臣宰、將軍、富戶、壯士，和一切為奴的、自主的，都藏在山洞和巖石穴裏，
REV|6|16|向山和巖石說：「倒在我們身上吧！把我們藏起來，躲避坐寶座者的臉面和羔羊的憤怒；
REV|6|17|因為他們遭憤怒的大日子到了，誰能站得住呢？」
REV|7|1|此後，我看見四位天使站在地的四角，執掌地上四方的風，使風不吹在地上、海上和各種樹上。
REV|7|2|我又看見另有一位天使從日出之地上來，拿著永生上帝的印。他向那得到權柄能傷害地和海的四位天使大聲喊著，
REV|7|3|說：「你們不可傷害地、海和樹林，等我們在我們上帝眾僕人的額上蓋了印。」
REV|7|4|我聽見 以色列 人各支派中受印的數目有十四萬四千；
REV|7|5|猶大 支派中受印的有一萬二千； 呂便 支派中有一萬二千； 迦得 支派中有一萬二千；
REV|7|6|亞設 支派中有一萬二千； 拿弗他利 支派中有一萬二千； 瑪拿西 支派中有一萬二千；
REV|7|7|西緬 支派中有一萬二千； 利未 支派中有一萬二千； 以薩迦 支派中有一萬二千；
REV|7|8|西布倫 支派中有一萬二千； 約瑟 支派中有一萬二千； 便雅憫 支派中受印的有一萬二千。
REV|7|9|此後，我觀看，看見有許多人，沒有人能計算，是從各邦國、各支派、各民族、各語言來的，站在寶座和羔羊面前，身穿白衣，手拿棕樹枝，
REV|7|10|大聲喊著說： 「願救恩歸於坐在寶座上我們的上帝， 也歸於羔羊！」
REV|7|11|眾天使都站在寶座和眾長老，以及四個活物的周圍，俯伏在寶座前，敬拜上帝，
REV|7|12|說： 「阿們！頌讚、榮耀、智慧、 感謝、尊貴、權能、 力量都歸於我們的上帝， 直到永永遠遠。阿們！」
REV|7|13|長老中有一位回應我說：「這些穿白衣的是誰？是從哪裏來的？」
REV|7|14|我對他說：「我主啊，你是知道的。」他向我說：「這些人是從大患難中出來的，他們曾用羔羊的血把衣裳洗得潔白。
REV|7|15|所以，他們在上帝寶座前， 晝夜在他殿中事奉他； 那坐在寶座上的要用帳幕覆庇他們。
REV|7|16|他們不再飢，不再渴； 太陽必不傷害他們， 任何炎熱也不傷害他們，
REV|7|17|因為寶座中的羔羊必牧養他們， 領他們到生命水的泉源； 上帝必擦去他們一切的眼淚。」
REV|8|1|羔羊揭開第七個印的時候，天上寂靜約有半小時。
REV|8|2|我看見那站在上帝面前的七位天使，有七枝號賜給他們。
REV|8|3|另有一位天使拿著金香爐來，站在祭壇旁邊；有許多香賜給他，要和眾聖徒的祈禱一同獻在寶座前的金壇上。
REV|8|4|那香的煙和眾聖徒的祈禱從天使的手中一同升到上帝面前。
REV|8|5|天使拿著香爐，盛滿了壇上的火，倒在地上；就有雷轟、響聲、閃電、地震。
REV|8|6|拿著七枝號筒的七位天使預備好要吹號。
REV|8|7|第一位天使吹號，就有冰雹和火攙著血扔在地上；地的三分之一和樹的三分之一被燒掉了，一切的青草也被燒掉了。
REV|8|8|第二位天使吹號，就有像火燒著的大山扔在海中；海的三分之一變成血，
REV|8|9|海中有生命的被造之物死了三分之一，船隻也毀壞了三分之一。
REV|8|10|第三位天使吹號，就有燒著的大星好像火把從天上墜下來，落在江河的三分之一和眾水的泉源上。
REV|8|11|這星名叫「苦艾」；眾水的三分之一變為苦艾，許多人因水變苦而死了。
REV|8|12|第四位天使吹號，太陽的三分之一、月亮的三分之一、星辰的三分之一都被擊打，以致日月星的三分之一變黑了，白晝的三分之一沒有光，黑夜也是這樣。
REV|8|13|我觀看，聽見一隻在空中飛的鷹大聲說：「禍哉！禍哉！禍哉！地上的居民哪，其餘的三位天使快要吹號了！」
REV|9|1|第五位天使吹號，我就看見一顆星從天上墜落到地上；有無底坑的鑰匙賜給它。
REV|9|2|它開了無底坑，就有煙從坑裏往上冒，好像大火爐的煙；太陽和天空都因這煙昏暗了。
REV|9|3|有蝗蟲從煙中出來，飛到地上，有權柄賜給牠們，好像地上的蠍子有權柄一樣。
REV|9|4|牠們奉命不可傷害地上的草、各樣綠色植物和各種樹木，惟獨可傷害額上沒有上帝印記的人；
REV|9|5|但是不許蝗蟲害死他們，只可使他們受痛苦五個月；這痛苦就像人被蠍子螫了的痛苦一樣。
REV|9|6|在那些日子，人求死，卻死不了；想死，死卻避開他們。
REV|9|7|蝗蟲的形狀好像預備上陣的戰馬一樣，頭上戴的好像金冠冕，臉面好像男人的臉面，
REV|9|8|頭髮像女人的頭髮，牙齒像獅子的牙齒；
REV|9|9|牠們胸前有甲，好像鐵甲；又有翅膀的響聲，好像許多車馬奔跑上陣的聲音。
REV|9|10|牠們有尾巴像蠍子，長著毒刺，尾巴上的毒刺有能力傷害人五個月。
REV|9|11|牠們有無底坑的使者作牠們的王，按著 希伯來 話名叫 亞巴頓 ， 希臘 話名話叫 亞玻倫 。
REV|9|12|第一樣災禍過去了；看哪，還有兩樣災禍要來。
REV|9|13|第六位天使吹號，我聽見有聲音從上帝面前金壇的四 角發出來，
REV|9|14|吩咐那吹號的第六位天使，說：「把那捆綁在 幼發拉底 大河的四個使者釋放了。」
REV|9|15|那四個使者就被釋放；他們原是預備好，在特定的年、月、日、時，要殺人類的三分之一。
REV|9|16|騎兵有二億；他們的數目我聽見了。
REV|9|17|我在異象中看見那些馬和騎馬的：騎馬的穿著火紅、紫瑪瑙及硫磺色的胸甲；馬的頭好像獅子的頭，有火、有煙、有硫磺從馬的口中噴出來。
REV|9|18|從馬的口中所噴出來的火、煙和硫磺這三樣災害殺了人類的三分之一。
REV|9|19|馬的能力在於牠們的口和尾巴；牠們的尾巴像蛇，有頭，用頭來傷害人。
REV|9|20|其餘未曾被這些災難所殺的人仍舊不為自己手所做的悔改，還是去拜鬼魔和那些不能看、不能聽、不能走，用金、銀、銅、木、石所造的偶像。
REV|9|21|他們也不為自己所犯的那些兇殺、邪術、淫亂、偷竊的事悔改。
REV|10|1|我又看見另一位大力的天使從天降下，披著雲彩，頭上有彩虹，臉面像太陽，兩腳像火柱。
REV|10|2|他手裏拿著展開的小書卷。他右腳踏海，左腳踏地，
REV|10|3|大聲呼喊，好像獅子吼叫。呼喊完了，就有七個雷發出聲音。
REV|10|4|七個雷發聲後，我正要寫出來，就聽見從天上有聲音說：「七個雷所說的，你要封上，不可寫出來。」
REV|10|5|我所看見的那踏海踏地的天使向天舉起右手，
REV|10|6|指著創造天和天上之物、地和地上之物、海和海中之物、直活到永永遠遠的那位起誓，說：「不再有時日了 。」
REV|10|7|但在第七位天使要吹號的日子，上帝的奧祕就要成全了，正如上帝向他僕人眾先知所宣告的。
REV|10|8|我先前從天上所聽見的那聲音又吩咐我說：「你去，把那踏海踏地之天使手中展開的小書卷拿過來。」
REV|10|9|我就走到天使那裏，對他說，請他把小書卷給我。他對我說：「你拿去，把它吃光。它會使你肚子發苦，然而在你口中會甘甜如蜜。」
REV|10|10|於是我從天使手中把小書卷接過來，把它吃光了，在我口中果然甘甜如蜜，吃了以後，我肚子覺得發苦。
REV|10|11|天使們對我說：「你必須指著許多民族、邦國、語言、君王再說預言。」
REV|11|1|有一根蘆葦，像丈量的杖，賜給我；且有話說：「起來！將上帝的殿和祭壇，以及在殿中禮拜的人，都量一量。
REV|11|2|只是殿外的院子不用量，因為這是要給外邦人的；他們將踐踏聖城四十二個月。
REV|11|3|「我要賜權柄給我那兩個見證人，穿著粗麻衣說預言一千二百六十天。」
REV|11|4|他們就是那站在世界之主面前的兩棵橄欖樹和兩個燈臺。
REV|11|5|若有人想要害他們，就有火從他們口中噴出來，燒滅仇敵；凡想要害他們的都必須這樣被殺。
REV|11|6|這二人有權柄關閉天空，使他們說預言的日子不下雨；又有權柄使水變為血，並且能隨時隨意用各樣的災害擊打大地世界。
REV|11|7|他們作完見證的時候，那從無底坑裏上來的獸要跟他們交戰，並且得勝，把他們殺了。
REV|11|8|他們的屍首將倒在大城的街道上；這城按著靈意叫 所多瑪 ，又叫 埃及 ，就是他們的主釘十字架的地方。
REV|11|9|從各民族、支派、語言、邦國中有人觀看他們的屍首三天半，又不許人把屍首安放在墳墓裏。
REV|11|10|住在地上的人會因他們而歡喜快樂，互相饋送禮物，因為這兩位先知曾使住在地上的人受痛苦。
REV|11|11|過了這三天半，有生命的氣息從上帝那裏進入他們裏面，他們就站起來；看見他們的人都大大懼怕。
REV|11|12|兩位先知聽見有大聲音從天上對他們說：「上這裏來。」他們就駕著雲上了天，他們的仇敵也看見了。
REV|11|13|正在那時候，地大震動，城倒塌了十分之一；因地震而死的有七千人，其餘的都恐懼，歸榮耀給天上的上帝。
REV|11|14|第二樣災禍過去了；看哪，第三樣災禍快到了。
REV|11|15|第七位天使吹號，天上就有大聲音說： 「世上的國已成了我們的主和他所立的基督的國了。 他要作王直到永永遠遠！」
REV|11|16|在上帝面前，坐在自己座位上的二十四位長老都俯伏在地上敬拜上帝，
REV|11|17|說： 「今在昔在的主—全能的上帝啊， 我們感謝你！ 因你執掌大權作王了。
REV|11|18|外邦發怒， 你的憤怒臨到了。 審判死人的時候也到了； 你的僕人眾先知、眾聖徒及敬畏你名的人， 連大帶小得賞賜的時候到了； 你毀滅那些毀滅大地者的時候也到了。」
REV|11|19|於是，上帝天上的聖所開了，在他聖所中，他的約櫃出現了；隨後有閃電、響聲、雷轟、地震、大冰雹。
REV|12|1|天上出現了一個大兆頭：有一個婦人身披太陽，腳踏月亮，頭戴十二顆星的冠冕；
REV|12|2|她懷了孕，在生產的陣痛中疼痛地喊叫。
REV|12|3|天上又出現了另一個兆頭：有一條大紅龍 ，有七個頭十個角；七個頭上戴著七個冠冕。
REV|12|4|牠的尾巴拖拉著天上星辰的三分之一，把它們摔在地上。然後龍站在那將要生產的婦人面前，等她生產後要吞吃她的孩子。
REV|12|5|婦人生了一個男孩子，就是將來要用鐵杖管轄 萬國的；她的孩子被提到上帝和他寶座那裏去。
REV|12|6|婦人就逃到曠野，在那裏有上帝給她預備的地方，使她在那裏被供養一千二百六十天。
REV|12|7|天上發生了爭戰。 米迦勒 同他的使者與龍作戰，龍同牠的使者也起來應戰，
REV|12|8|牠們都打敗了，天上再也沒有牠們的地方。
REV|12|9|大龍就是那古蛇，名叫魔鬼，又叫撒但，是迷惑普天下的；牠被摔在地上，牠的使者也一同被摔下去。
REV|12|10|我聽見在天上有大聲音說： 「我上帝的救恩、能力、國度， 和他所立的基督的權柄現在都來到了。 因為那個在我們上帝面前、 晝夜控告我們弟兄的， 已經被摔下去了。
REV|12|11|弟兄勝過那條龍是因羔羊的血， 和因自己所見證的道。 雖然至於死，他們也不惜自己的性命。
REV|12|12|所以，諸天和住在其中的， 你們都快樂吧！ 只是地和海有禍了！ 因為魔鬼知道自己的時候不多， 就氣憤憤地下到你們那裏去了。」
REV|12|13|龍見自己被摔在地上，就迫害那生男孩子的婦人。
REV|12|14|於是有大鷹的兩個翅膀賜給婦人，讓她能飛到曠野，到自己的地方，躲避那蛇。她在那裏受供養一載二載半載。
REV|12|15|蛇在婦人背後，從口中噴出水來，像河一樣，要將婦人沖走。
REV|12|16|地卻幫助了婦人，開口吞了從龍口噴出來的水。
REV|12|17|於是龍向婦人發怒，去與她其餘的兒女作戰，就是與那些遵守上帝命令 、為耶穌作見證的 。
REV|12|18|那時龍站在海邊沙灘上。
REV|13|1|我又看見一隻獸從海裏上來，有十個角七個頭；在十個角上戴著十個冠冕，七個頭上有褻瀆的名號。
REV|13|2|我所看見的獸，形狀像豹，腳像熊的腳，口像獅子的口。那條龍將自己的能力、座位和大權柄都給了牠。
REV|13|3|我看見獸的七個頭中，有一個似乎受了致命傷，那傷卻醫好了。全地的人都很驚訝，跟從了那隻獸。
REV|13|4|他們都拜那條龍，因為牠把自己的權柄給了獸；又拜那隻獸，說：「誰能比這隻獸，誰能與牠交戰呢？」
REV|13|5|龍又賜給那隻獸說誇大褻瀆話的口，又賜給牠權柄可以任意行事四十二個月。
REV|13|6|那獸就開口向上帝說褻瀆的話，褻瀆上帝的名和他的帳幕，就是那些住在天上的。
REV|13|7|牠又被准許與聖徒作戰，並且得勝，也賜給牠權柄，可以制伏各支派、各民族、各語言、各邦國。
REV|13|8|凡住在地上、名字從創世以來沒有記在被殺羔羊的生命冊上的人都要拜牠。
REV|13|9|凡有耳朵的都聽吧！
REV|13|10|該被擄掠的，必被擄掠； 該被刀殺的，必被刀殺。 在此，聖徒要有耐心和信心。
REV|13|11|我又看見另一隻獸從地裏上來。牠有兩個角如同羔羊，說話好像龍。
REV|13|12|牠在第一隻獸面前施行第一隻獸所有的權柄，並且使地和住在地上的人拜那致命傷被醫好了的第一隻獸。
REV|13|13|這隻獸又行大奇事，甚至在人面前使火從天降在地上。
REV|13|14|牠得了權柄在第一隻獸面前能行奇事，迷惑住在地上的人，告訴他們要為那受過刀傷還活著的獸造個像。
REV|13|15|又有權柄賜給牠，讓那隻獸的像有生氣，並且能說話，又使所有不拜獸像的人都被殺害。
REV|13|16|牠又使眾人，無論大小、貧富，自主的、為奴的，都在右手上，或是在額上，打一個印記；
REV|13|17|這樣，除了那有印記，有獸的名或有獸名數字的，都不得買或賣。
REV|13|18|在此，要有智慧：讓有悟性的人解開獸的數目吧，因為這是一個人的數字，那數字是六百六十六。
REV|14|1|我又觀看，看見羔羊站在 錫安山 ，和他在一起的有十四萬四千人，都有他的名和他父親的名寫在額上。
REV|14|2|我聽見從天上有聲音，像眾水的聲音和大雷的聲音，我所聽見的聲音好像琴師所彈的琴聲。
REV|14|3|他們在寶座前，和在四活物及眾長老前唱新歌，除了從地上買來的那十四萬四千人以外，沒有人能學這歌。
REV|14|4|這些人未曾沾染婦女，他們原是童身。羔羊無論往哪裏去，他們都跟隨他。他們是從人間買來的，作為初熟的果子歸給上帝和羔羊。
REV|14|5|在他們口中找不出謊言，他們是沒有瑕疵的。
REV|14|6|我又看見另一位天使在空中飛翔，有永遠的福音要傳給住在地上的人，就是各邦國、各支派、各語言、各民族。
REV|14|7|他大聲說：「要敬畏上帝，把榮耀歸給他，因為他施行審判的時候已經到了。要敬拜那創造天、地、海和水源的主。」
REV|14|8|另有第二位天使接著說：「傾覆了！那曾叫列國喝淫亂、烈怒之酒的大 巴比倫 傾覆了！」
REV|14|9|另有第三位天使接著他們，大聲說：「若有人拜那隻獸和獸像，在額上或在手上受了印記，
REV|14|10|他也必喝上帝烈怒的酒；這酒是斟在上帝憤怒的杯中的純酒。他要在聖天使和羔羊面前，在火與硫磺之中受痛苦。
REV|14|11|使他們受痛苦的煙往上冒，直到永永遠遠。那些拜獸和獸像，受了牠名字的印記的人，晝夜不得安寧。」
REV|14|12|在此，遵守上帝命令 和堅信耶穌真道的聖徒要有耐心。
REV|14|13|我聽見從天上有聲音說：「你要寫下：從今以後，在主裏死去的人有福了。」聖靈說：「是的，他們要從自己的勞苦中得安息，因為工作的成果永隨著他們。」
REV|14|14|我又觀看，看見有一片白雲，雲上坐著一位好像是人子的，頭上戴著金冠冕，手裏拿著鋒利的鐮刀。
REV|14|15|另有一位天使從聖所出來，向那坐在雲上的大聲喊著：「伸出你的鐮刀來收割吧，因為收割的時候已經到了，地上的莊稼已經熟透了。」
REV|14|16|於是那坐在雲上的把鐮刀向地上揮去，地上的莊稼就收割了。
REV|14|17|另有一位天使從天上的聖所出來，他也拿著鋒利的鐮刀。
REV|14|18|另有一位天使從祭壇出來，是有權柄管火的，向那拿著鋒利鐮刀的大聲喊著說：「伸出鋒利的鐮刀來，收取地上葡萄樹的果子，因為葡萄熟透了。」
REV|14|19|那天使就把鐮刀向地上揮去，收取了地上的葡萄，扔進上帝憤怒的大醡酒池裏。
REV|14|20|那醡酒池在城外被踹踏，有血從醡酒池裏流出來，漲到馬的嚼環那麼高，約有一千六百斯他迪 那麼遠。
REV|15|1|我看見在天上有另一兆頭，大而且奇，就是七位天使掌管末了的七種災難，因為上帝的烈怒在這七種災難中發盡了。
REV|15|2|我看見彷彿有攙雜火的玻璃海；又看見那些勝了那獸和獸像，以及牠名字的數字的人，都站在玻璃海上，拿著上帝的豎琴。
REV|15|3|他們唱上帝僕人 摩西 的歌和羔羊的歌，說： 「主—全能的上帝啊， 你的作為又偉大又奇妙！ 萬國之王啊， 你的道路又公義又真實！
REV|15|4|主啊，誰敢不敬畏你， 不把榮耀歸於你的名？ 因為只有你是神聖的。 萬民都要來， 在你面前敬拜， 因你公義的作為已經彰顯了。」
REV|15|5|此後，我看見在天上那存放法櫃的聖所開了。
REV|15|6|那掌管七種災難的七位天使從聖所出來，穿著潔白明亮的細麻衣 ，胸間束著金帶。
REV|15|7|四個活物中，有一個把盛滿了活到永永遠遠之上帝烈怒的七個金碗給了那七位天使。
REV|15|8|聖所中充滿了上帝的榮耀和權能而來的煙。沒有人能進入聖所，直等到那七位天使降完了七種災難。
REV|16|1|我聽見有大聲音從聖所裏出來，向那七位天使說：「你們去，把盛著上帝烈怒的七碗傾倒在地上。」
REV|16|2|第一位天使去，把碗傾倒在地上，就有又臭又毒的瘡生在那些有獸的印記和拜獸像的人身上。
REV|16|3|第二位天使把碗傾倒在海裏，海就變成像死人的血一樣，海裏所有的活物都死了。
REV|16|4|第三位天使把碗傾倒在河流和水源裏，水就變成血了。
REV|16|5|我聽見掌管眾水的天使說： 「昔在、今在的聖者啊， 你做的判斷公義；
REV|16|6|因他們曾流過聖徒與先知的血， 現在你給他們血喝， 這是他們該受的。」
REV|16|7|我又聽見祭壇中有聲音說： 「是的，主—全能的上帝啊， 你的判斷又真實又公義！」
REV|16|8|第四位天使把碗傾倒在太陽上，使太陽可用火烤人。
REV|16|9|人被炎熱所烤，就褻瀆那有權掌管這些災難的上帝的名，他們沒有悔改，也沒有把榮耀歸給上帝。
REV|16|10|第五位天使把碗傾倒在獸的座位上，獸的國就變成黑暗。人因疼痛而咬自己的舌頭；
REV|16|11|又因所受的疼痛和生的瘡，就褻瀆天上的上帝，也沒有為他們的行為悔改。
REV|16|12|第六位天使把碗傾倒在大 幼發拉底河 上，河水就乾了，為要給從日出之地所來的眾王預備道路。
REV|16|13|我又看見三個污穢的靈，好像青蛙，從龍的口、獸的口和假先知的口中出來。
REV|16|14|他們本是鬼魔的靈，施行奇事，到普天下眾王那裏去，召集他們在全能者上帝的大日子作戰。
REV|16|15|看哪，我來像賊一樣。那警醒、穿著衣服的人有福了；他不至於赤身而行，給人看見他的羞恥。
REV|16|16|於是，那三個鬼魔把眾王聚集在 希伯來 話叫作 哈米吉多頓 的地方。
REV|16|17|第七位天使把碗傾倒在空中，就有大聲音從聖所的寶座上出來，說：「成了！」
REV|16|18|又有閃電、響聲、雷轟、大地震，自從地上有人以來沒有這樣大、這樣厲害的地震。
REV|16|19|那大城裂為三段，列國的城也都倒塌了。上帝記起了大 巴比倫城 ，把那盛自己烈怒的酒杯遞給她。
REV|16|20|各海島都逃避了，眾山也不見了。
REV|16|21|又有大冰雹從天掉落在人身上，每一個約重一他連得，以致人因冰雹的災難而褻瀆上帝，因為那災難太大了。
REV|17|1|拿著七個碗的七位天使中，有一位前來對我說：「來，我要讓你看那坐在眾水之上的大淫婦所要受的懲罰；
REV|17|2|地上的君王都曾與她行淫，住在地上的人也喝醉了她淫亂的酒。」
REV|17|3|我在聖靈感動下，被天使帶到曠野去，我看見一個女人騎在朱紅色的獸上；那隻獸有七個頭十個角，遍體有褻瀆的名號。
REV|17|4|那女人穿著紫色和朱紅色的衣服，用金子、寶石、珍珠作妝飾，手拿著金杯，杯中盛滿了可憎之物和她淫亂的污穢。
REV|17|5|在她額上寫著奧祕的名字，說：「大 巴比倫 ，世上的淫婦和一切可憎之物的母。」
REV|17|6|我又看見那女人喝醉了聖徒的血和為耶穌作見證的人的血。 我看見她，非常詫異。
REV|17|7|天使對我說：「你為甚麼詫異呢？我要把這女人和馱著她那七頭十角的獸的奧祕告訴你。
REV|17|8|你曾看見的獸，以前有，現在沒有，將來要從無底坑裏上來，又歸於沉淪。凡住在地上、名字從創世以來沒有記在生命冊上的人看見那隻獸都要詫異，因為牠以前有，現在沒有，以後再有。
REV|17|9|在此要有智慧的心思：那七個頭就是女人所坐的七座山；他們又是七個王，
REV|17|10|五個已經倒了，一個還在，一個還沒有來到；他來的時候必須只暫時停留。
REV|17|11|那以前有、現在沒有的獸就是第八個，他也和那七個同列，正歸於沉淪。
REV|17|12|你曾看見的那十個角就是十個王；他們還沒有得到國度，但他們要和那隻獸同得權柄作王一個時辰。
REV|17|13|他們同心把自己的能力權柄交給那隻獸。
REV|17|14|他們將與羔羊作戰，羔羊必勝過他們，因為羔羊是萬主之主、萬王之王，而同羔羊在一起的是蒙召、被選、忠心的人。」
REV|17|15|天使又對我說：「你所看見那淫婦坐的眾水，就是許多民族、人民、邦國、語言。
REV|17|16|你所看見的那十個角與獸必恨這淫婦，他們要使她孤獨赤身，又要吃她的肉，用火將她燒盡。
REV|17|17|因為上帝使諸王同心執行他的旨意，把他們自己的國交給那隻獸，直等到上帝的話都應驗了。
REV|17|18|你所看見的那女人就是管轄地上眾王的大城。」
REV|18|1|此後，我看見另一位有大權柄的天使從天降下，地由於他的榮耀而發光。
REV|18|2|他以強而有力的聲音喊著說： 「傾覆了！大 巴比倫 傾覆了！ 她成了鬼魔的住處， 各樣污穢之靈的巢穴， 各樣污穢之鳥的窩， 各樣污穢可憎之獸的出沒處 。
REV|18|3|因為列國都喝了她淫亂大怒的酒 ； 地上的君王和她行淫； 地上的商人因她極度奢華而發了財。」
REV|18|4|我又聽見另一個聲音從天上說： 「我的民哪，從那城出來吧！ 免得和她在罪上有份， 受她所受的災殃；
REV|18|5|因她的罪惡滔天， 上帝已經記得她的不義。
REV|18|6|她怎樣待人，也要怎樣待她， 按她所行的加倍地報應她； 用她調酒的杯加倍調給她喝。
REV|18|7|她怎樣榮耀自己，怎樣奢華， 也要使她照樣痛苦悲哀。 因她心裏說： 『我坐了皇后的位， 並不是寡婦， 絕不至於悲哀。』
REV|18|8|所以在一天之內，她的災殃要一齊來到， 就是死亡、悲哀、饑荒。 她將被火燒盡， 因為審判她的主上帝大有能力。」
REV|18|9|地上的君王，與她行淫、一同奢華的，看見燒她的煙，就必為她哭泣哀號；
REV|18|10|因怕她的痛苦，就遠遠地站著，說： 「禍哉，禍哉，這大城！ 堅固的 巴比倫城 啊！ 一時之間，你的審判要來到了。」
REV|18|11|地上的商人也都為她哭泣悲哀，因為沒有人再買他們的貨物了；
REV|18|12|這貨物就是金、銀、寶石、珍珠、細麻布、絲綢、紫色和朱紅色衣料、各樣香木、各樣象牙的器皿、各樣極寶貴的木頭和銅、鐵、大理石的器皿，
REV|18|13|和肉桂、豆蔻、香料、香膏、乳香、酒、油、細麵、麥子、牛、羊、馬、馬車，以及奴隸、人口。
REV|18|14|「你所貪愛的果子離開了你； 你一切的珍饈美味和華美的物件 都從你那裏毀滅， 絕對見不到了。」
REV|18|15|販賣這些貨物、藉著她發財的商人，因怕她的痛苦，就遠遠地站著哭泣悲哀，
REV|18|16|說： 「禍哉，禍哉，這大城！ 她穿著細麻、 紫色、朱紅色的衣服， 用金子、寶石、珍珠為妝飾。
REV|18|17|一時之間，這麼多的財富就歸於無有了。」 所有的船長和到處航海的，水手以及所有靠海為業的，都遠遠地站著，
REV|18|18|看見燒她的煙，就喊著說：「有哪一個城能跟這大城比呢？」
REV|18|19|於是他們把灰塵撒在頭上，哭泣悲哀地喊著說： 「禍哉，禍哉，這大城！ 凡有船在海中的， 都因她的珍寶成了富足。 她在一時之間就成為荒蕪。
REV|18|20|天哪，眾聖徒、眾使徒、眾先知啊！ 你們都要因她歡喜， 因為上帝已經在她身上為你們伸了冤。」
REV|18|21|有一位大力的天使舉起一塊石頭，好像大磨石，扔在海裏，說： 「 巴比倫 大城 也必這樣猛力地被扔下去， 絕對見不到了。
REV|18|22|彈琴、歌唱、 吹笛、吹號的聲音， 在你中間絕對聽不見了； 各行手藝的技工 在你中間絕對見不到了； 推磨的聲音 在你中間絕對聽不見了；
REV|18|23|燈臺的光 在你中間絕對不再照耀了； 新郎和新娘的聲音 在你中間絕對聽不見了。 你的商人原來是地上的顯要； 萬國也被你的邪術迷惑了。
REV|18|24|先知、聖徒和地上一切被殺的人的血都在這城裏找到了。」
REV|19|1|此後，我聽見好像有一大群人在天上大聲說： 「哈利路亞 ！ 救恩、榮耀、權能都屬於我們的上帝。
REV|19|2|他的判斷又真實又公義； 因他判斷了那大淫婦， 她用淫行敗壞了世界。 上帝為他的僕人伸冤， 向淫婦討流僕人血的罪。」
REV|19|3|他們又一次說： 「哈利路亞！ 燒淫婦的煙往上冒，直到永永遠遠。」
REV|19|4|那二十四位長老和四活物就俯伏敬拜坐在寶座上的上帝，說： 「阿們。哈利路亞！」
REV|19|5|接著，有聲音從寶座出來說： 「上帝的眾僕人哪， 凡敬畏他的， 無論大小， 都要讚美我們的上帝！」
REV|19|6|我聽見好像一大群人的聲音，像眾水的聲音，像大雷的聲音，說： 「哈利路亞！ 因為主─我們的上帝 、 全能者，作王了。
REV|19|7|我們要歡喜快樂， 將榮耀歸給他； 因為羔羊的婚期到了， 他的新娘也自己預備好了，
REV|19|8|她蒙恩得穿明亮潔白的細麻衣： 這細麻衣就是聖徒們的義行。」
REV|19|9|天使對我說：「你要寫下來：凡被請赴羔羊婚宴的人有福了！」他又對我說：「這些都是上帝真實的話。」
REV|19|10|我就俯伏在他腳前要拜他。他對我說：「千萬不可！我和你，以及那些為耶穌作見證的弟兄同是僕人。你要敬拜上帝。」因為那些為耶穌作見證的人有預言的靈。
REV|19|11|後來我看見天開了。有一匹白馬，騎在馬上的稱為 「誠信」、「真實」，他審判和爭戰都憑著公義。
REV|19|12|他的眼睛如 火焰，頭上戴著許多冠冕；他身上寫著一個名字，除了他自己沒有人知道。
REV|19|13|他穿著浸過血的衣服；他的名稱為「上帝之道」。
REV|19|14|眾天軍都騎著白馬，穿著又白又潔淨的細麻衣跟隨他。
REV|19|15|有利劍從他口中出來，用來擊打列國。他要用鐵杖管轄 他們，並且要踹全能上帝烈怒的醡酒池。
REV|19|16|在他衣服和大腿上寫著「萬王之王，萬主之主」的名號。
REV|19|17|我又看見一位天使站在太陽中，向天空一切的飛鳥大聲喊著說：「你們聚集來赴上帝的大宴席，
REV|19|18|為要吃君王的肉、將軍的肉、壯士的肉、馬和騎士的肉、一切自主的和為奴的，以及尊貴的和卑賤的肉。」
REV|19|19|我又看見那獸和地上的君王，和他們的軍隊都聚集，要與白馬騎士和他的軍隊作戰。
REV|19|20|那獸被擒拿了；那在獸面前曾行奇事、迷惑了接受獸的印記和拜獸像的人的假先知，也與獸同被擒拿。他們兩個就活生生地被扔進燒著硫磺的火湖裏，
REV|19|21|其餘的人被白馬騎士口中吐出來的劍殺了；所有的飛鳥都吃飽了他們的肉。
REV|20|1|我又看見一位天使從天降下，手裏拿著無底坑的鑰匙和一條大鐵鏈。
REV|20|2|他抓住那龍，那古蛇，就是魔鬼、撒但，把牠捆綁了一千年，
REV|20|3|扔在無底坑裏，把無底坑關閉，用印封上，使牠不再迷惑列國，等到那一千年滿了。這些事以後，牠必須暫時被釋放。
REV|20|4|我又看見一些寶座，坐在上面的有審判的權柄賜給他們。我又看見那些因為給耶穌作見證，並為上帝之道被斬首的人的靈魂，和沒有拜過那獸與獸像、也沒有在額上和手上打過牠印記的人的靈魂。他們都復活了，與基督一同作王一千年。
REV|20|5|這是頭一次的復活。其餘的死人還沒有復活，直等那一千年滿了。
REV|20|6|在頭一次復活有份的有福了，聖潔了！第二次的死在他們身上沒有權柄，但他們要作上帝和基督的祭司，也要與基督一同作王一千年。
REV|20|7|那一千年滿了，撒但會從監牢裏被釋放，
REV|20|8|出來要迷惑地上四方的列國，就是 歌革 和 瑪各 ，使他們聚集爭戰。他們的人數多如海沙。
REV|20|9|他們上來佈滿了全地，圍住聖徒的營與蒙愛的城，就有火從天降下，燒滅了他們。
REV|20|10|那迷惑他們的魔鬼被扔進硫磺的火湖裏，就是那獸和假先知所在的地方，他們會晝夜受折磨，直到永永遠遠。
REV|20|11|我又看見一個白色的大寶座和那坐在上面的；天和地都從他面前逃避，再也找不到它們的位置了。
REV|20|12|我又看見死了的人，無論大小，都站在寶座前。案卷都展開了，並另有一卷展開，就是生命冊。死了的人都憑著這些案卷所記載的，照他們所行的受審判。
REV|20|13|於是海交出其中的死人，死亡和陰間也交出其中的死人；他們都照各人所行的受審判。
REV|20|14|死亡和陰間也被扔進火湖裏，這火湖就是第二次的死。
REV|20|15|凡名字沒有記在生命冊上的人，就被扔進火湖裏。
REV|21|1|我又看見一個新天新地，因為先前的天和先前的地已經過去了，海也不再有了。
REV|21|2|我又看見聖城，新 耶路撒冷 由上帝那裏，從天而降，預備好了，就如新娘打扮整齊，等候丈夫。
REV|21|3|我聽見有大聲音從寶座出來，說： 「看哪，上帝的帳幕在人間！ 他要和他們同住， 他們要作他的子民。 上帝要親自與他們同在。
REV|21|4|上帝要擦去他們一切的眼淚； 不再有死亡， 也不再有悲哀、哭號、痛苦， 因為先前的事都過去了。」
REV|21|5|那位坐在寶座上的說：「看哪，我把一切都更新了！」他又說：「你要寫下來，因為這些話是可信靠的，是真實的。」
REV|21|6|他又對我說：「成了！我是阿拉法，我是俄梅戛；我是開始，我是終結。我要把生命的泉水白白賜給那口渴的人喝。
REV|21|7|得勝的要承受這些為業；我要作他的上帝，他要作我的兒子。
REV|21|8|至於膽怯的、不信的、可憎的、殺人的、淫亂的、行邪術的、拜偶像的和一切說謊話的人，他們將在燒著硫磺的火湖裏有份；這是第二次的死。」
REV|21|9|拿著七個金碗、盛滿末後七種災禍的七位天使中，有一位來對我說：「你來，我要給你看新娘，就是羔羊的妻子。」
REV|21|10|我在聖靈感動下，天使帶我到一座高大的山，給我看由上帝那裏、從天而降的聖城 耶路撒冷 ，
REV|21|11|這城有上帝的榮耀，它光輝如同極貴的寶石，好像碧玉，明如水晶。
REV|21|12|它有高大的牆，有十二個門，門上有十二位天使，門上又寫著 以色列 人十二個支派的名字 。
REV|21|13|東邊有三個門，北邊有三個門，南邊有三個門，西邊有三個門。
REV|21|14|城牆有十二個根基，根基上有羔羊十二使徒的名字。
REV|21|15|那對我說話的天使拿著金的蘆葦當尺，要量那城、城門和城牆。
REV|21|16|城是四方的，長寬一樣。天使用蘆葦量那城，共有一萬二千斯他迪，長、寬、高都是一樣。
REV|21|17|他又量了城牆，按著人的尺寸，就是天使的尺寸，共有一百四十四肘。
REV|21|18|牆是碧玉造的；城是純金的，如同明淨的玻璃。
REV|21|19|城牆的根基是用各樣寶石修飾的：第一個根基是碧玉，第二是藍寶石，第三是綠瑪瑙，第四是綠寶石，
REV|21|20|第五是紅瑪瑙，第六是紅寶石，第七是黃璧璽，第八是水蒼玉，第九是紅璧璽，第十是翡翠，第十一是紫瑪瑙，第十二是紫晶。
REV|21|21|十二個門是十二顆珍珠；每一個門是一顆珍珠造的。城內的街道是純金的，好像透明的玻璃。
REV|21|22|我沒有看見城內有殿，因主—全能者上帝和羔羊就是城的殿。
REV|21|23|那城內不用日月光照，因為有上帝的榮耀光照，又有羔羊為城的燈。
REV|21|24|列國要藉著城的光行走；地上的君王要把自己的榮耀帶給那城。
REV|21|25|城門白晝總不關閉，在那裏沒有黑夜。
REV|21|26|人要將列國的榮耀尊貴帶給那城。
REV|21|27|凡不潔淨的，和那行可憎與虛謊之事的人，都不得進那城，只有名字寫在羔羊生命冊上的才得進去。
REV|22|1|天使又讓我看一道生命水的河，明亮如水晶，從上帝和羔羊的寶座流出來，
REV|22|2|經過城內街道的中央；在河的兩邊有生命樹，結十二樣 的果子，每月都結果子；樹上的葉子可作醫治萬民之用。
REV|22|3|以後不再有任何詛咒。在城裏將有上帝和羔羊的寶座。他的僕人都要事奉他，
REV|22|4|也要見他的面。他的名字將寫在他們的額上。
REV|22|5|不再有黑夜；他們也不需要燈光或日光，因為主上帝要光照他們。他們要作王，直到永永遠遠。
REV|22|6|天使又對我說：「這些話是可信靠的，是真實的。主，就是賜靈感給眾先知的上帝，差遣他的使者，要將必須快要發生的事指示他的眾僕人。」
REV|22|7|「看哪，我必快來！凡遵守這書上預言的有福了。」
REV|22|8|這些事是我－ 約翰 所聽見所看見的。當我聽見看見時，就俯伏在指示我的天使腳前要拜他。
REV|22|9|他對我說：「千萬不可！我與你和你的弟兄眾先知，以及那些守這書上的話的人，同是作僕人。你要敬拜上帝。」
REV|22|10|他又對我說：「不可封了這書上的預言，因為時候近了。
REV|22|11|不義的，讓他仍舊不義；污穢的，讓他仍舊污穢；為義的，讓他仍舊為義；聖潔的，讓他仍舊聖潔。」
REV|22|12|「看哪，我必快來！賞罰在我，要照每個人所行的報應他。
REV|22|13|我是阿拉法，我是俄梅戛；我是首先的，我是末後的；我是開始，我是終結。」
REV|22|14|那些洗淨自己衣服的有福了！他們可得權柄到生命樹那裏，也能從門進城。
REV|22|15|城外有犬類、行邪術的、淫亂的、殺人的、拜偶像的，以及所有喜愛和行虛謊的人。
REV|22|16|「我－耶穌差遣我的使者，為了眾教會向你們證明這些事。我是 大衛 的根，是他的後裔；我是明亮的晨星。」
REV|22|17|聖靈和新娘都說：「來！」聽見的人也要說：「來！」口渴的人也要來，願意的人都可以白白取生命的水喝。
REV|22|18|我警告一切聽見這書上預言的人：若有人在這預言上加添甚麼，上帝必將記在這書上的災禍加在他身上。
REV|22|19|這書上的預言，若有人刪去甚麼，上帝必從這書上所記的生命樹和聖城刪去他的份。
REV|22|20|證明這些事的說：「是的，我必快來！」阿們！主耶穌啊，我願你來！
REV|22|21|願主耶穌的恩惠與眾聖徒同在。阿們！
