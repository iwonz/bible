2THESS|1|1|保羅 、 西拉 和 提摩太 寫信給 帖撒羅尼迦 、在我們的父上帝與主耶穌基督裏的教會。
2THESS|1|2|願恩惠、平安 從我們的 父上帝和主耶穌基督歸給你們！
2THESS|1|3|弟兄們，我們該常常為你們感謝上帝，這本是合宜的；因為你們的信心格外增長，你們眾人彼此相愛的心也都增加。
2THESS|1|4|所以，我們在上帝的各教會裏為你們誇耀，因為你們在所受的一切壓迫患難中仍牢守著耐心和信心。
2THESS|1|5|這正是上帝公義判斷的明證，使你們配得上他的國，你們就是為這國受苦。
2THESS|1|6|既然上帝是公義的，他必以患難報復那加患難給你們的人，
2THESS|1|7|也必使你們這受患難的人與我們同得平安。那時，主耶穌同他有權能的天使從天上在火焰中顯現，要報應那些不認識上帝和不聽從我們的主耶穌福音的人。
2THESS|1|8|
2THESS|1|9|他們要受懲罰，永遠沉淪，與主的面和他權能的榮光隔絕。
2THESS|1|10|這正是主再來，要在他聖徒的身上得榮耀，就是要使一切信的人感到驚訝的那日子，因為你們信了我們對你們作的見證。
2THESS|1|11|為此，我們常為你們禱告，願我們的上帝看你們與他的呼召相配，又用大能成就你們一切良善的美意和因信心所做的工作，
2THESS|1|12|使我們主耶穌的名，照著我們的上帝和主耶穌基督的恩，在你們身上得榮耀，你們也在他身上得榮耀。
2THESS|2|1|弟兄們，關於我們主耶穌基督的來臨和我們到他那裏聚集，我勸你們：
2THESS|2|2|無論藉著靈，藉著言語，藉著冒我的名寫的書信，說主的日子已經到了，不要輕易動心，也不要驚慌。
2THESS|2|3|不要讓任何人用甚麼法子欺騙你們，因為那日子以前必有叛教的事，並有那不法的人，那沉淪之子出現。
2THESS|2|4|那抵擋者高抬自己超過一切稱為神明的，和一切受人敬拜的，甚至坐在上帝的殿裏，自稱為上帝。
2THESS|2|5|我還在你們那裏的時候曾把這些事告訴你們，你們不記得嗎？
2THESS|2|6|現在你們也知道那攔阻他的是甚麼，為要使他到了時機才出現。
2THESS|2|7|因為那不法的隱祕已經運作，只是現在有一個阻擋的，要等到那阻擋的被除去才會發作，
2THESS|2|8|那時這不法的人必出現，主耶穌 要用口中的氣滅絕他，以自己來臨的光輝摧毀他。
2THESS|2|9|這不法的人來，是靠撒但的運作，行各樣的異能、神蹟和一切虛假的奇事，
2THESS|2|10|並且在那沉淪的人身上行各樣不義的詭詐，因為他們不領受愛真理的心，好讓他們得救。
2THESS|2|11|故此，上帝就給他們一個引發錯誤的心，叫他們信從虛謊，
2THESS|2|12|使一切不信真理、倒喜愛不義的人都被定罪。
2THESS|2|13|主所愛的弟兄們哪，我們本該常為你們感謝上帝，因為他揀選你們為初熟的果子 ，使你們因信真道，又蒙聖靈感化成聖，得到拯救。
2THESS|2|14|為此，上帝藉著我們所傳的福音呼召你們，好得著我們主耶穌基督的榮光。
2THESS|2|15|所以，弟兄們，你們要站立得穩，凡所領受的教導，無論是我們口傳的，是信上寫的，都要堅守。
2THESS|2|16|願我們主耶穌基督自己，和那愛我們、開恩將永遠的安慰及美好的盼望賜給我們的父上帝，
2THESS|2|17|安慰你們的心，並且在一切善行善言上堅固你們！
2THESS|3|1|末了，弟兄們，請你們為我們禱告，好讓主的道快快傳開，得著榮耀，正如在你們中間一樣，
2THESS|3|2|也讓我們能脫離無理和邪惡人的手，因為不是人人都有信仰。
2THESS|3|3|但主是信實的，他要堅固你們，保護你們脫離那邪惡者。
2THESS|3|4|我們靠主對你們有信心，你們現在遵行，以後也必遵行我們所吩咐的。
2THESS|3|5|願主引導你們的心去愛上帝，並學基督的忍耐！
2THESS|3|6|弟兄們，我們奉主耶穌基督的名吩咐你們，凡有弟兄懶散，不遵守我們所傳授的教導，要遠離他。
2THESS|3|7|你們自己知道該怎樣效法我們。因為我們在你們當中從未懶散過，
2THESS|3|8|也從未白吃人的飯，倒是辛苦勞碌，晝夜做工，免得使你們中間有人受累。
2THESS|3|9|這並不是因我們沒有權柄，而是要給你們作榜樣，好讓你們效法我們。
2THESS|3|10|我們在你們那裏的時候曾吩咐你們，說若有人不肯做工，就不可吃飯。
2THESS|3|11|因為我們聽說，在你們中間有人懶散，甚麼工都不做，反倒專管閒事。
2THESS|3|12|我們靠主耶穌基督吩咐並勸戒這樣的人，要安分做工，自食其力。
2THESS|3|13|弟兄們，你們行善不可喪志。
2THESS|3|14|若有人不聽從我們這信上的話，要把他記下，不和他交往，使他自覺羞愧；
2THESS|3|15|但不要把他當仇人，要勸他如勸弟兄。
2THESS|3|16|願賜平安 的主隨時隨事親自賜給你們平安！願主與你們眾人同在！
2THESS|3|17|我— 保羅 親筆向你們問安。凡我的信都以此為記，我的筆跡就是這樣。
2THESS|3|18|願我們主耶穌基督的恩惠與你們眾人同在！
