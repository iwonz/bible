PS|1|1|不从恶人的计谋， 不站罪人的道路， 不坐傲慢人的座位， 惟喜爱耶和华的律法， 昼夜思想 他的律法； 这人便为有福！
PS|1|2|
PS|1|3|他要像一棵树栽在溪水旁， 按时候结果子， 叶子也不枯干。 凡他所做的尽都顺利。
PS|1|4|恶人并不是这样， 却像糠秕被风吹散。
PS|1|5|因此，当审判的时候恶人必站立不住， 罪人在义人的会众中也是如此。
PS|1|6|因为耶和华知道义人的道路， 恶人的道路却必灭亡。
PS|2|1|列国为什么争闹？ 万民为什么图谋虚妄？
PS|2|2|世上的君王都站稳， 臣宰一同算计， 要对抗耶和华， 对抗他的受膏者：
PS|2|3|“我们要挣脱他们的捆绑， 脱去他们的绳索。”
PS|2|4|那坐在天上的必讥笑， 主必嗤笑他们。
PS|2|5|那时，他要在怒中责备他们， 在烈怒中惊吓他们：
PS|2|6|“我已经在 锡安 －我的圣山 膏立了我的君王。”
PS|2|7|我要传耶和华的圣旨， 他对我说：“你是我的儿子， 我今日生了你。
PS|2|8|你求我，我就将列国赐你为基业， 将地极赐你为田产。
PS|2|9|你必用铁杖打破他们， 把他们如同陶匠的瓦器摔碎。”
PS|2|10|现在，君王啊，应当谨慎！ 世上的审判官哪，要听劝戒！
PS|2|11|当存敬畏的心事奉耶和华， 又当战兢而快乐。
PS|2|12|当亲吻儿子，免得他发怒， 你们就在半途中灭亡， 因为他的怒气快要发作。 凡投靠他的，都是有福的。
PS|3|1|耶和华啊，我的敌人何其增多！ 许多人起来攻击我。
PS|3|2|许多人议论我： “他得不到上帝的帮助。”（细拉）
PS|3|3|但你－耶和华是我四围的盾牌， 是我的荣耀，又是令我抬起头来的。
PS|3|4|我用我的声音求告耶和华， 他就从他的圣山上应允我。（细拉）
PS|3|5|我躺下，我睡觉，我醒来， 耶和华都保佑我。
PS|3|6|虽有成万的百姓周围攻击我， 我也不惧怕。
PS|3|7|耶和华啊，求你兴起！ 我的上帝啊，求你救我！ 因为你打断我所有仇敌的腮骨， 敲碎了恶人的牙齿。
PS|3|8|救恩属于耶和华； 愿你赐福给你的百姓。（细拉）
PS|4|1|显我为义的上帝啊， 我呼求的时候，求你应允我！ 我在困境中，你曾使我宽畅； 求你怜悯我，听我的祷告！
PS|4|2|你们这些人哪，你们把我的尊荣变为羞辱，要到几时呢？ 你们喜爱虚妄，寻找虚假，要到几时呢？ （细拉）
PS|4|3|你们要知道，耶和华已将虔诚人分别出来归他自己； 我求告耶和华，他必垂听。
PS|4|4|应当畏惧，不可犯罪； 在床上的时候，要心里思想，并要安静。（细拉）
PS|4|5|当献上公义的祭， 又当倚靠耶和华。
PS|4|6|有许多人说：“谁能指示我们什么好处？ 耶和华啊，求你用你脸上的光照耀我们。”
PS|4|7|你使我心里喜乐， 胜过那丰收五谷新酒的人。
PS|4|8|我必平安地躺下睡觉， 因为独有你－耶和华使我安然居住。
PS|5|1|耶和华啊，求你侧耳听我的言语， 顾念我的心思！
PS|5|2|我的王，我的上帝啊，求你留心听我呼求的声音！ 因为我向你祈祷。
PS|5|3|耶和华啊，早晨你必听我的声音； 早晨我要向你陈明我的心思，并要警醒。
PS|5|4|因为你不是喜爱邪恶的上帝， 恶人不能与你同住。
PS|5|5|狂傲的人不能站在你眼前； 凡作恶的，都是你所恨恶的。
PS|5|6|说谎言的，你必灭绝； 好流人血、玩弄诡诈的，都为耶和华所憎恶。
PS|5|7|至于我，我必凭你丰盛的慈爱进入你的居所， 我要存敬畏你的心向你的圣殿下拜。
PS|5|8|耶和华啊，求你因我仇敌的缘故，凭你的公义引领我， 使你的道路在我面前正直。
PS|5|9|因为他们口中没有诚实， 心里充满邪恶， 他们的喉咙是敞开的坟墓； 他们用舌头谄媚人。
PS|5|10|上帝啊，求你定他们的罪！ 愿他们因自己的计谋跌倒； 求你因他们过犯众多赶逐他们， 因为他们背叛了你。
PS|5|11|凡投靠你的，愿他们喜乐，时常欢呼， 因为你庇护他们； 又愿那爱你名的人都靠你欢欣。
PS|5|12|耶和华啊，因为你必赐福给义人， 你必用恩惠如同盾牌四面护卫他。
PS|6|1|耶和华啊，求你不要在怒中责备我， 不要在烈怒中惩罚我！
PS|6|2|耶和华啊，求你怜悯我，因为我软弱。 耶和华啊，求你医治我，因为我的骨头战抖。
PS|6|3|我的心也大大惊惶。 耶和华啊，你要等到几时呢？
PS|6|4|耶和华啊，求你转回搭救我， 因你的慈爱拯救我。
PS|6|5|因为死了的人不会记念你， 在阴间有谁称谢你？
PS|6|6|我因呻吟而困乏； 我每夜流泪，使床铺漂起， 把褥子湿透。
PS|6|7|我的眼睛因忧愁而昏花， 因敌人的缘故，我的眼目模糊不清。
PS|6|8|你们所有作恶的人，离开我吧！ 因为耶和华听了我哀哭的声音。
PS|6|9|耶和华听了我的恳求， 耶和华必接纳我的祷告。
PS|6|10|我所有的仇敌都必羞愧，大大惊惶； 转眼之间，他们要羞愧撤退。
PS|7|1|耶和华－我的上帝啊，我投靠你！ 求你救我脱离所有追赶我的人，搭救我出来！
PS|7|2|免得他们像狮子撕裂我， 甚至撕碎，无人搭救。
PS|7|3|耶和华－我的上帝啊，我若行了这事， 若有罪孽在我手里，
PS|7|4|我若以恶回报我的朋友， 连那无故与我为敌的，我也救了他 ，
PS|7|5|就任凭仇敌追赶我，直到追上， 把我的性命踏在地上， 使我的荣耀归于灰尘。（细拉）
PS|7|6|耶和华啊，求你在怒中起来， 挺身而立，抵挡我敌人的烈怒！ 求你为我兴起！你已经发令施行审判。
PS|7|7|愿万民聚集环绕你！ 愿你居高位统治他们！
PS|7|8|耶和华向万民施行审判； 耶和华啊，求你按我的公义 和我心中的纯正判断我。
PS|7|9|愿恶人的恶断绝！ 愿你坚立义人！ 因为公义的上帝察验人的心肠肺腑。
PS|7|10|上帝是我的盾牌， 他拯救心里正直的人。
PS|7|11|上帝是公义的审判者， 又是天天向恶人发怒的上帝。
PS|7|12|若有人不回头，他的刀必磨快， 弓必上弦，预备妥当。
PS|7|13|他也预备了致死的兵器， 他所射的是火箭。
PS|7|14|看哪，恶人怀邪恶， 养毒害，生虚假。
PS|7|15|他掘了坑，挖得太深， 竟掉在自己所挖的陷阱里。
PS|7|16|他的毒害必回到自己头上， 他的残暴必落到自己的脑袋上。
PS|7|17|我要照着耶和华的公义称谢他， 要歌颂耶和华至高者的名。
PS|8|1|耶和华－我们的主啊， 你的名在全地何其美！ 你将你的荣耀彰显于天 。
PS|8|2|你因敌人的缘故， 从孩童和吃奶的口中建立了能力， 使仇敌和报仇的闭口无言。
PS|8|3|我观看你手指所造的天， 并你所陈设的月亮星宿。
PS|8|4|人算什么，你竟顾念他！ 世人算什么，你竟眷顾他！
PS|8|5|你使他比上帝 微小一点， 赐他荣耀尊贵为冠冕。
PS|8|6|你派他管理你手所造的， 使万物，就是一切的牛羊、 田野的牲畜、空中的鸟、海里的鱼， 凡游在水里的，都服在他的脚下。
PS|8|7|
PS|8|8|
PS|8|9|耶和华－我们的主啊， 你的名在全地何其美！
PS|9|1|我要一心称谢耶和华， 传扬你一切奇妙的作为。
PS|9|2|我要因你欢喜快乐； 至高者啊，我要歌颂你的名！
PS|9|3|我的仇敌回转撤退的时候， 他们在你面前跌倒灭亡。
PS|9|4|因你已经为我伸冤，为我辩护； 你坐在宝座上，按公义审判。
PS|9|5|你曾斥责列国，灭绝恶人； 你曾涂去他们的名，直到永永远远。
PS|9|6|仇敌到了尽头； 他们遭毁坏，直到永远。 你拆毁他们的城镇， 连他们的名字 也都消灭！
PS|9|7|惟耶和华坐在王位上，直到永远； 他已经为审判摆设宝座。
PS|9|8|他要按公义审判世界， 按正直判断万民。
PS|9|9|耶和华要作受欺压者的庇护所， 在患难时的庇护所。
PS|9|10|耶和华啊，认识你名的人要倚靠你， 因你没有离弃寻求你的人。
PS|9|11|应当歌颂居于 锡安 的耶和华， 将他所做的传扬在万民中。
PS|9|12|那位追讨流人血的， 他记念受屈的人， 不忘记困苦人的哀求。
PS|9|13|耶和华啊，求你怜悯我！ 你是从死门把我提升起来的， 求你看那恨我的人所加给我的苦难，
PS|9|14|好让我述说你一切的美德。 我要在 锡安 的城门因你的救恩欢乐。
PS|9|15|外邦人陷在自己所掘的坑中， 他们的脚被自己暗设的网罗缠住了。
PS|9|16|耶和华已将自己显明，他已施行审判； 恶人被自己手所做的缠住了 。（细拉）
PS|9|17|恶人，就是忘记上帝的外邦人， 都必归到阴间。
PS|9|18|贫穷人必不永久被忘， 困苦人的指望必不永远落空。
PS|9|19|耶和华啊，求你兴起，不容世人得胜！ 愿外邦人在你面前受审判！
PS|9|20|耶和华啊，求你使他们恐惧， 愿外邦人知道自己不过是人。（细拉）
PS|10|1|耶和华啊，你为什么站在远处？ 在患难的时候为什么隐藏？
PS|10|2|恶人骄横地追逼困苦人； 愿他们陷在自己所设的计谋里。
PS|10|3|因为恶人以自己的心愿自夸， 贪财的背弃耶和华，并且轻慢他 。
PS|10|4|恶人面带骄傲，不寻找耶和华； 他的思想中全无上帝。
PS|10|5|他的路时常亨通， 你的审判不在他眼里。 至于他所有的敌人，他都向他们发怒气。
PS|10|6|他心里说：“我必不动摇， 世世代代不遭灾难。”
PS|10|7|他满口咒骂、诡诈、欺压， 舌底尽是毒害、奸恶。
PS|10|8|他在村庄埋伏等候， 在隐密处杀害无辜的人， 他的眼睛窥探无倚无靠的人。
PS|10|9|他埋伏在暗地，如狮子蹲在洞中。 他埋伏，要俘掳困苦人； 他拉网，就把困苦人掳去。
PS|10|10|他屈身蹲伏， 无倚无靠的人就倒在他的暴力之下。
PS|10|11|他心里说：“上帝竟忘记了， 上帝转脸永不观看。”
PS|10|12|耶和华啊，求你兴起！ 上帝啊，求你举手！ 不要忘记困苦人！
PS|10|13|恶人为何轻慢上帝， 心里说“你必不追究”？
PS|10|14|你已经察看， 顾念人的忧患和愁苦， 放在你的手中。 无倚无靠的人把自己交托给你， 你向来是帮助孤儿的。
PS|10|15|求你打断恶人的膀臂， 至于坏人，求你追究他的恶，直到净尽。
PS|10|16|耶和华永永远远为王， 外邦人从他的地已经灭绝了。
PS|10|17|耶和华啊，困苦人的心愿你早已听见； 你必坚固他们的心，也必侧耳听他们的祈求，
PS|10|18|为要给孤儿和受欺压的人伸冤， 使世上的人不再威吓他们。
PS|11|1|我投靠耶和华； 你们怎么对我说：“你当像鸟逃到你们的山去；
PS|11|2|看哪，恶人弯弓，把箭搭在弦上， 要在暗中射那心里正直的人。
PS|11|3|根基若毁坏， 义人还能做什么呢？”
PS|11|4|耶和华在他的圣殿里， 耶和华在天上的宝座上； 他的眼睛察看， 他的眼目 察验世人。
PS|11|5|耶和华考验义人； 惟有恶人和喜爱暴力的人，他心里恨恶。
PS|11|6|他要向恶人密布罗网， 烈火、硫磺、热风作他们杯中的份。
PS|11|7|因为耶和华是公义的，他喜爱义行， 正直人必得见他的面。
PS|12|1|耶和华啊，求你帮助，因虔诚人断绝了， 世人中间忠信的人消失了。
PS|12|2|人人向邻舍说谎； 他们说话嘴唇油滑，心口不一。
PS|12|3|愿耶和华剪除一切油滑的嘴唇， 夸大的舌头。
PS|12|4|他们说：“我们必能以舌头取胜， 我们的嘴唇是自己的， 谁能作我们的主呢？”
PS|12|5|耶和华说：“因为困苦人的冤屈 和贫穷人的叹息， 我现在要起来， 把他安置在他所切慕的稳妥之地。”
PS|12|6|耶和华的言语是纯净的言语， 如同银子在泥做的炉中炼过七次。
PS|12|7|耶和华啊，你必保护他们， 你必保佑他们永远脱离这世代的人。
PS|12|8|卑鄙的人在世人中高升时， 就有恶人四处横行。
PS|13|1|耶和华啊，你忘记我要到几时呢？要到永远吗？ 你转脸不顾我要到几时呢？
PS|13|2|我心里筹算，终日愁苦，要到几时呢？ 我的仇敌升高压制我，要到几时呢？
PS|13|3|耶和华－我的上帝啊，求你看顾我，应允我！ 求你使我眼目明亮，免得我沉睡至死；
PS|13|4|免得我的仇敌说“我胜了他”； 免得我的敌人在我动摇的时候喜乐。
PS|13|5|但我倚靠你的慈爱， 我的心因你的救恩快乐。
PS|13|6|我要向耶和华歌唱， 因他厚厚地恩待我。
PS|14|1|愚顽人心里说：“没有上帝。” 他们都败坏，行了可憎恶的事， 没有一个人行善。
PS|14|2|耶和华从天上垂看世人， 要看有明白的没有， 有寻求上帝的没有。
PS|14|3|他们都偏离正路，一同变为污秽， 没有行善的， 连一个也没有。
PS|14|4|作恶的都没有知识吗？ 他们吞吃我的百姓如同吃饭一样， 并不求告耶和华。
PS|14|5|他们在那里大大害怕， 因为上帝在义人的族类中。
PS|14|6|你们叫困苦人的筹算变为羞辱， 然而耶和华是他的避难所。
PS|14|7|但愿 以色列 的救恩出自 锡安 。 当耶和华救回他被掳子民的时候， 雅各 要快乐， 以色列 要欢喜。
PS|15|1|耶和华啊，谁能寄居你的帐幕？ 谁能居住你的圣山？
PS|15|2|就是行为正直、做事公义、 心里说实话的人。
PS|15|3|他不以舌头谗害人， 不恶待朋友， 也不随伙毁谤邻舍。
PS|15|4|他眼中藐视匪类， 却尊重那敬畏耶和华的人。 他发了誓，虽然自己吃亏也不更改。
PS|15|5|他不放债取利， 不受贿赂以害无辜。 做这些事的人必永不动摇。
PS|16|1|上帝啊，求你保佑我， 因为我投靠你。
PS|16|2|我 曾对耶和华说：“你是我的主， 我的福气惟独从你而来。”
PS|16|3|论到世上的圣民，他们是尊贵的人， 是我最喜悦的。
PS|16|4|追逐 别神的， 他们的愁苦必增加； 他们所浇奠的血我不献上， 我嘴唇也不提别神的名号。
PS|16|5|耶和华是我的产业，是我杯中的福分； 我所得的，你为我持守。
PS|16|6|用绳量给我的地界，坐落在佳美之处； 我的产业实在美好。
PS|16|7|我要称颂那指引我的耶和华， 在夜间我的心肠也指教我。
PS|16|8|我让耶和华常在我面前， 因他在我右边，我就不致动摇。
PS|16|9|因此，我的心欢喜，我的灵 快乐； 我的肉身也要安然居住。
PS|16|10|因为你必不将我的灵魂 撇在阴间， 也不让你的圣者见地府 。
PS|16|11|你必将生命的道路指示我。 在你面前有满足的喜乐， 在你右手中有永远的福乐。
PS|17|1|耶和华啊，求你垂听公义的呼声， 留心听我的呼求！ 求你侧耳听我这没有诡诈的嘴唇的祈祷！
PS|17|2|愿判我公正的话从你面前发出， 愿你的眼睛察看正直。
PS|17|3|你已经考验我的心， 你在夜间鉴察我。 你熬炼我，却找不到错失， 我立志叫我口中没有过失。
PS|17|4|论到人的行为，我谨守你嘴唇的言语， 不走残暴人的道路。
PS|17|5|我的脚紧紧跟随你的脚踪， 我的两脚未曾滑跌。
PS|17|6|上帝啊，我求告你，因为你必应允我； 求你向我侧耳，听我的言语。
PS|17|7|求你显出你奇妙的慈爱， 你用右手拯救投靠你的人，脱离那起来攻击他们的人。
PS|17|8|求你保护我，如同保护眼中的瞳人， 把我隐藏在你翅膀的荫下，
PS|17|9|使我脱离欺压我的恶人， 脱离那围困我要害我命的仇敌。
PS|17|10|他们的心被油脂包裹， 用口说骄傲的话。
PS|17|11|他们追逼我 ，现在他们围困了我们， 瞪着眼，要把我们推倒在地。
PS|17|12|他像狮子要贪吃猎物， 又像少壮狮子蹲伏在暗处。
PS|17|13|耶和华啊，求你兴起，前去迎敌，把他打倒！ 求你用你的刀救我的命脱离恶人。
PS|17|14|耶和华啊，求你用手救我脱离世人， 脱离那只在今生有福分的世人！ 你以财宝充满他们的肚腹， 他们因有儿女就满足， 将其余的财物留给他们的孩子。
PS|17|15|至于我，我必因公正得见你的面； 我醒了的时候，你的形像使我满足。
PS|18|1|耶和华我的力量啊，我爱你！
PS|18|2|耶和华是我的岩石、我的山寨、我的救主、 我的上帝、我的磐石、我所投靠的。 他是我的盾牌， 是拯救我的角，是我的碉堡。
PS|18|3|我要求告当赞美的耶和华， 我必从仇敌手中被救出来。
PS|18|4|死亡的绳索勒住我， 毁灭的急流惊吓我，
PS|18|5|阴间的绳索缠绕我， 死亡的圈套临到我。
PS|18|6|我在急难中求告耶和华， 向我的上帝呼求。 他从殿中听了我的声音， 我在他面前的呼求必进入他耳中。
PS|18|7|那时，因他发怒地就震动战抖， 山的根基也震动挪移。
PS|18|8|他的鼻孔冒烟上腾， 他的口发火焚烧，连煤炭也烧着了。
PS|18|9|他使天垂下，亲自降临， 黑云在他脚下。
PS|18|10|他乘坐基路伯飞行， 藉着风的翅膀快飞，
PS|18|11|以黑暗为藏身之处， 以水的黑暗、天空的密云作四围的行宫。
PS|18|12|因他发出光辉， 冰雹和火炭穿透密云。
PS|18|13|耶和华在天上打雷， 至高者发出声音，就有冰雹和火炭 。
PS|18|14|他射出箭来，使仇敌四散； 发出连串的闪电，击溃他们。
PS|18|15|耶和华啊，你的斥责一发， 你鼻孔的气一出， 海底就显现， 大地的根基也暴露。
PS|18|16|他从高天伸手抓住我， 把我从大水中拉上来。
PS|18|17|他救我脱离强敌和那些恨我的人， 因为他们比我强盛。
PS|18|18|我遭遇灾难的日子，他们来攻击我； 但耶和华是我的倚靠。
PS|18|19|他领我到宽阔之处， 他救拔我，因他喜爱我。
PS|18|20|耶和华必按我的公义报答我， 按我手中的清洁赏赐我。
PS|18|21|因为我遵守耶和华的道， 未曾作恶离开我的上帝。
PS|18|22|他的一切典章常在我面前， 他的律例我也未曾丢弃。
PS|18|23|我在他面前作了完全人， 我也保护自己远离罪孽。
PS|18|24|所以耶和华按我的公义， 在他眼前按我手中的清洁赏赐我。
PS|18|25|慈爱的人，你以慈爱待他； 完全的人，你以完善待他。
PS|18|26|清洁的人，你以清洁待他； 歪曲的人，你以弯曲待他。
PS|18|27|困苦的百姓，你必拯救； 高傲的眼目，你使他降卑。
PS|18|28|你必点亮我的灯； 耶和华－我的上帝必照明我的黑暗。
PS|18|29|我藉着你冲入敌军， 藉着我的上帝跳过城墙。
PS|18|30|至于上帝，他的道是完全的； 耶和华的话是纯净的。 凡投靠他的，他就作他们的盾牌。
PS|18|31|除了耶和华，谁是上帝呢？ 除了我们的上帝，谁是磐石呢？
PS|18|32|惟有那以力量束我的腰、 使我行为完全的，他是上帝。
PS|18|33|他使我的脚快如母鹿， 使我站稳在高处。
PS|18|34|他教导我的手能争战， 我的膀臂能开铜造的弓。
PS|18|35|你赐救恩给我作盾牌， 你的右手扶持我， 你的庇护 使我为大。
PS|18|36|你使我脚步宽阔， 我的脚踝未曾滑跌。
PS|18|37|我要追赶我的仇敌，且要追上他们； 若不将他们灭绝，我总不归回。
PS|18|38|我要打伤他们，使他们站不起来； 他们必倒在我的脚下。
PS|18|39|你曾以力量束我的腰，使我能争战； 也曾使那起来攻击我的，都服在我以下。
PS|18|40|你又使我的仇敌在我面前转身逃跑， 使我剪除那恨我的人。
PS|18|41|他们呼求，却无人拯救； 就是呼求耶和华，他也不应允。
PS|18|42|我捣碎他们，如同风前的灰尘； 倾倒 他们，如同街上的泥土。
PS|18|43|你救我脱离百姓的纷争， 立我作列国的元首； 我素不认识的百姓必事奉我。
PS|18|44|他们一听见我的名声就必顺从我， 外邦人要投降我。
PS|18|45|外邦人要丧胆， 战战兢兢地出营寨。
PS|18|46|耶和华永远活着。 愿我的磐石被称颂， 愿救我的上帝受尊崇。
PS|18|47|这位上帝为我伸冤， 使万民服在我以下。
PS|18|48|他拯救我脱离仇敌， 又把我举起，高过那些起来攻击我的人， 救我脱离残暴的人。
PS|18|49|耶和华啊，因此我要在外邦中称谢你， 歌颂你的名。
PS|18|50|耶和华赐极大的救恩给他所立的王， 施慈爱给他的受膏者， 就是给 大卫 和他的后裔，直到永远。
PS|19|1|诸天述说上帝的荣耀， 穹苍传扬他手的作为。
PS|19|2|这日到那日发出言语， 这夜到那夜传出知识。
PS|19|3|无言无语， 也无声音可听。
PS|19|4|它们的声浪 传遍天下， 它们的言语传到地极。 上帝在其中为太阳安设帐幕，
PS|19|5|太阳如同新郎步出洞房， 又如勇士欢然奔路。
PS|19|6|它从天这边出来，绕到天那边， 没有一物可隐藏得不到它的热气。
PS|19|7|耶和华的律法全备，使人苏醒； 耶和华的法度确定，使愚蒙人有智慧。
PS|19|8|耶和华的训词正直，使人心快活； 耶和华的命令清洁，使人眼目明亮。
PS|19|9|耶和华的典章真实，全然公义， 敬畏耶和华是纯洁的，存到永远，
PS|19|10|比金子可羡慕，比极多的纯金可羡慕； 比蜜甘甜，比蜂房下滴的蜜甘甜。
PS|19|11|因此你的仆人受警戒， 遵守这些有极大的赏赐。
PS|19|12|谁能察觉自己的错失呢？ 求你赦免我隐藏的过犯。
PS|19|13|求你拦阻仆人不犯任意妄为的罪， 不容这罪辖制我， 我就完全，免犯大罪。
PS|19|14|耶和华－我的磐石，我的救赎主啊， 愿我口中的言语，心里的意念在你面前蒙悦纳。
PS|20|1|愿耶和华在你患难的日子应允你， 愿 雅各 的上帝的名保护你。
PS|20|2|愿他从圣所救助你， 从 锡安 坚固你，
PS|20|3|记念你的一切祭物， 悦纳你的燔祭，（细拉）
PS|20|4|将你心所愿的赐给你， 成就你的一切筹算。
PS|20|5|我们要因你的救恩夸胜， 要奉我们上帝的名竖立旌旗。 愿耶和华成就你一切所求的！
PS|20|6|现在我知道耶和华必救护他的受膏者， 从他神圣的天上应允他， 用右手的能力救护他。
PS|20|7|有人靠车，有人靠马， 但我们要提耶和华－我们上帝的名。
PS|20|8|他们都屈身仆倒， 我们却起来，坚立不移。
PS|20|9|耶和华啊，求你拯救； 我们呼求的时候，愿王应允我们！
PS|21|1|耶和华啊，王必因你的能力欢喜； 因你的救恩，他的快乐何其大！
PS|21|2|他心里所愿的，你已经赐给他； 他嘴唇所求的，你未尝不应允。（细拉）
PS|21|3|你以美善的福气迎接他， 把纯金的冠冕戴在他头上。
PS|21|4|他向你祈求长寿，你就赐给他， 就是日子长久，直到永远。
PS|21|5|他因你的救恩大有荣耀， 你将尊荣威严加在他身上。
PS|21|6|你使他有洪福，直到永远， 又使他在你面前欢喜快乐。
PS|21|7|王倚靠耶和华， 因至高者的慈爱，王必不动摇。
PS|21|8|你的手要搜出所有的仇敌， 你的右手要搜出那些恨你的人。
PS|21|9|你的脸出现的时候，要使他们如在炎热的火炉中。 耶和华要在他的震怒中吞灭他们， 那火要把他们烧尽。
PS|21|10|你必从世上灭绝他们的幼苗， 从人间灭绝他们的后裔。
PS|21|11|因为他们有意加害于你； 他们想出计谋，却不能做成。
PS|21|12|你必使他们转身逃跑， 向着他们的脸搭箭在弦。
PS|21|13|耶和华啊，愿你因自己的能力显为至高！ 这样，我们就唱诗，歌颂你的大能。
PS|22|1|我的上帝，我的上帝，为什么离弃我？ 为什么远离不救我，不听我的呻吟？
PS|22|2|我的上帝啊，我白日呼求，你不应允； 夜间呼求，也不得安宁。
PS|22|3|但你是神圣的， 用 以色列 的赞美为宝座。
PS|22|4|我们的祖宗倚靠你； 他们倚靠你，你解救他们。
PS|22|5|他们哀求你，就蒙解救； 他们倚靠你，就不羞愧。
PS|22|6|但我是虫，不是人， 被众人羞辱，被百姓藐视。
PS|22|7|凡看见我的都嗤笑我； 他们撇嘴摇头：
PS|22|8|“他把自己交托给耶和华，让耶和华救他吧！ 耶和华既喜爱他，可以搭救他吧！”
PS|22|9|但你是叫我出母腹的， 我在母怀里，你就使我有倚靠的心。
PS|22|10|我自出母胎就交在你手里， 自我出母腹，你就是我的上帝。
PS|22|11|求你不要远离我！ 因为灾难临头，无人帮助。
PS|22|12|许多公牛环绕我， 巴珊 大力的公牛四面围困我。
PS|22|13|它们向我张口， 好像猎食吼叫的狮子。
PS|22|14|我如水被倒出， 我的骨头都脱了节， 我的心如蜡，在我里面熔化。
PS|22|15|我的精力枯干，如同瓦片， 我的舌头紧贴上颚。 你将我安置在死灰中。
PS|22|16|犬类围着我，恶党环绕我； 他们扎了我的手、我的脚。
PS|22|17|我数遍我的骨头； 他们瞪着眼看我。
PS|22|18|他们分我的外衣， 为我的内衣抽签。
PS|22|19|耶和华啊，求你不要远离我！ 我的救主啊，求你快来帮助我！
PS|22|20|求你救我的性命脱离刀剑， 使我仅有的 脱离犬类，
PS|22|21|求你救我脱离狮子的口； 你已经应允我，使我脱离野牛的角。
PS|22|22|我要将你的名传给我的弟兄， 在会众中我要赞美你。
PS|22|23|敬畏耶和华的人哪，要赞美他！ 雅各 的后裔啊，要荣耀他！ 以色列 的后裔啊，要惧怕他！
PS|22|24|因为他没有藐视、憎恶受苦的人， 也没有转脸不顾他们； 那受苦之人呼求的时候，他就垂听。
PS|22|25|我在大会中赞美你的话是从你而来， 我要在敬畏耶和华的人面前还我的愿。
PS|22|26|愿困苦的人吃得饱足， 愿寻求耶和华的人赞美他。 愿你们的心永远活着！
PS|22|27|地的四极都要想念耶和华，并且归顺他， 列国的万族都要在你面前敬拜。
PS|22|28|因为国度属于耶和华， 他是管理列国的。
PS|22|29|地上富足的人都必吃喝而敬拜， 凡下到尘土中不能存活自己性命的人， 都要在他面前下拜 ；
PS|22|30|必有后裔事奉他， 主所做的事必传给后代。
PS|22|31|他们必来传他的公义给尚未出生的子民， 这是他的作为。
PS|23|1|耶和华是我的牧者， 我必不致缺乏。
PS|23|2|他使我躺卧在青草地上， 领我在可安歇的水边。
PS|23|3|他使我的灵魂苏醒 ， 为自己的名引导我走义路。
PS|23|4|我虽然行过死荫的幽谷， 也不怕遭害， 因为你与我同在； 你的杖、你的竿，都安慰我。
PS|23|5|在我敌人面前，你为我摆设筵席； 你用油膏了我的头，使我的福杯满溢。
PS|23|6|我一生一世必有恩惠慈爱随着我； 我且要住在 耶和华的殿中，直到永远。
PS|24|1|地和其中所充满的， 世界和住在其中的，都属耶和华。
PS|24|2|他把地建立在海上， 安定在江河之上。
PS|24|3|谁能登耶和华的山？ 谁能站在他的圣所？
PS|24|4|就是手洁心清，意念不向虚妄， 起誓不怀诡诈的人。
PS|24|5|他必蒙耶和华赐福， 又蒙救他的上帝使他成义。
PS|24|6|这是寻求耶和华的族类， 是寻求你面的 雅各 。（细拉）
PS|24|7|众城门哪，要抬起头来！ 永久的门户啊，你们要被举起！ 荣耀的王将要进来！
PS|24|8|这荣耀的王是谁呢？ 就是有力有能的耶和华， 在战场上大有能力的耶和华！
PS|24|9|众城门哪，要抬起头来！ 永久的门户啊，你们要高举！ 荣耀的王将要进来！
PS|24|10|这荣耀的王是谁呢？ 万军之耶和华是荣耀的王！（细拉）
PS|25|1|耶和华啊，我的心仰望你。
PS|25|2|我的上帝啊，我素来倚靠你； 求你不要叫我羞愧， 不要叫我的仇敌向我夸胜。
PS|25|3|凡等候你的必不羞愧， 惟有那无故行奸诈的必要羞愧。
PS|25|4|耶和华啊，求你将你的道指示我， 将你的路指教我！
PS|25|5|求你指教我，引导我进入你的真理， 因为你是救我的上帝。 我整日等候你。
PS|25|6|耶和华啊，求你记念你的怜悯和慈爱， 因为这是亘古以来所常有的。
PS|25|7|求你不要记得我幼年的罪愆和我的过犯； 耶和华啊，求你因你的良善，按你的慈爱记念我。
PS|25|8|耶和华是良善正直的， 因此，他必教导罪人走正路。
PS|25|9|他要按公平引领谦卑人， 将他的道指教他们。
PS|25|10|凡遵守他的约和他法度的人， 耶和华都以慈爱信实待他。
PS|25|11|耶和华啊，求你因你名的缘故赦免我的罪， 因我的罪重大。
PS|25|12|谁敬畏耶和华， 耶和华必教导他当选择的道路。
PS|25|13|他要安然居住， 他的后裔必承受土地。
PS|25|14|耶和华与敬畏他的人亲密， 他要将自己的约指示他们。
PS|25|15|我的眼目时常仰望耶和华， 因他必将我的脚从网里拉出来。
PS|25|16|求你转向我，怜悯我， 因我孤独困苦。
PS|25|17|我心里愁苦甚多， 求你救我脱离我的祸患。
PS|25|18|求你看顾我的困苦、我的艰难， 赦免我一切的罪。
PS|25|19|求你察看我的仇敌， 因为他们人数众多，并且痛恨我。
PS|25|20|求你保护我的性命，搭救我， 使我不致羞愧，因为我投靠你。
PS|25|21|愿纯全、正直保护我， 因为我等候你。
PS|25|22|上帝啊，求你救赎 以色列 脱离他一切的愁苦。
PS|26|1|耶和华啊，求你为我伸冤， 因我向来行事纯正； 我倚靠耶和华，必不动摇。
PS|26|2|耶和华啊，求你察看我，考验我， 熬炼我的肺腑心肠。
PS|26|3|因为你的慈爱常在我眼前， 我也按你的真理而行。
PS|26|4|我未曾与虚妄的人同坐， 也不与伪善的人来往。
PS|26|5|我痛恨恶人的集会， 必不与恶人同坐。
PS|26|6|耶和华啊，我要洗手表明无辜， 才环绕你的祭坛；
PS|26|7|我好发出称谢的声音， 述说你一切奇妙的作为。
PS|26|8|耶和华啊，我喜爱你所住的殿 和你显荣耀的居所。
PS|26|9|不要把我的性命和罪人一同除掉， 不要把我的生命和好流人血的一同除掉。
PS|26|10|他们的手中有奸恶， 他们的右手满有贿赂。
PS|26|11|至于我，却要行事纯正； 求你救赎我，怜悯我！
PS|26|12|我的脚站在平坦的地方， 在聚会中我要称颂耶和华！
PS|27|1|耶和华是我的亮光，是我的拯救， 我还怕谁呢？ 耶和华是我生命的保障， 我还惧谁呢？
PS|27|2|那作恶的就是我的仇敌， 前来吃我肉的时候就绊跌仆倒。
PS|27|3|虽有军队安营攻击我，我的心也不害怕； 虽然兴起战争攻击我，我仍旧安稳。
PS|27|4|有一件事，我曾求耶和华，我仍要寻求， 就是一生一世住在耶和华的殿中， 瞻仰他的荣美，在他的殿宇里求问。
PS|27|5|因为我遭遇患难，他必将我隐藏在他的帐棚里， 把我藏在他帐幕的隐密处， 将我高举在磐石上。
PS|27|6|现在我得以昂首，高过四面的仇敌。 我要在他的帐幕里欢然献祭， 我要唱诗歌颂耶和华。
PS|27|7|耶和华啊，我呼求的时候，求你垂听我的声音； 求你怜悯我，应允我。
PS|27|8|你说：“你们当寻求我的面。” 那时我的心向你说： “耶和华啊，你的面我正要寻求。”
PS|27|9|求你不要转脸不顾我， 不要发怒赶逐你的仆人， 你向来是帮助我的。 救我的上帝啊，不要离开我， 也不要撇弃我。
PS|27|10|即使我的父母撇弃我， 耶和华终必收留我。
PS|27|11|耶和华啊，求你将你的道指教我， 因我仇敌的缘故引导我走平坦的路。
PS|27|12|求你不要把我交给敌人，遂其所愿； 因为妄作见证的和口吐凶言的都起来攻击我。
PS|27|13|我深信在活人之地 必得见耶和华的恩惠。
PS|27|14|要等候耶和华， 当壮胆，坚固你的心， 要等候耶和华！
PS|28|1|耶和华啊，我要求告你！ 我的磐石啊，求你不要向我缄默！ 倘若你向我闭口， 我就如下入地府的人一样。
PS|28|2|我呼求你，向你至圣所举手的时候， 求你垂听我恳求的声音！
PS|28|3|不要把我和坏人并作恶的一同除掉； 他们跟邻舍说平安，心里却是奸恶。
PS|28|4|求你按着他们所做的， 按他们的恶行对待他们； 求你照着他们手所做的对待他们， 将他们应得的报应加给他们。
PS|28|5|他们既然不尊重耶和华的作为， 也不尊重他手所做的， 耶和华就必毁坏他们，不建立他们。
PS|28|6|耶和华是应当称颂的， 因为他听了我恳求的声音。
PS|28|7|耶和华是我的力量，是我的盾牌， 我心里倚靠他就得帮助。 我心中欢乐， 我要用诗歌称谢他。
PS|28|8|耶和华是他百姓的力量， 又是他受膏者得救的保障。
PS|28|9|求你拯救你的百姓，赐福给你的产业； 求你牧养他们，扶持他们，直到永远。
PS|29|1|上帝的子民 哪，你们要将荣耀、能力归给耶和华， 都归给耶和华！
PS|29|2|要将耶和华的名的荣耀归给他， 要敬拜神圣荣耀的耶和华 。
PS|29|3|耶和华的声音在众水上， 荣耀的上帝打雷； 耶和华打雷在大水之上。
PS|29|4|耶和华的声音大有能力， 耶和华的声音满有威严。
PS|29|5|耶和华的声音震碎香柏树， 耶和华震碎 黎巴嫩 的香柏树。
PS|29|6|他使 黎巴嫩 跳跃如牛犊， 使 西连 跳跃如野牛犊。
PS|29|7|耶和华的声音使火焰分岔。
PS|29|8|耶和华的声音震动旷野， 耶和华震动 加低斯 的旷野。
PS|29|9|耶和华的声音惊动母鹿落胎， 树林也脱落净光。 凡在他殿中的，都述说他的荣耀。
PS|29|10|耶和华坐在洪水之上为王； 耶和华坐着为王，直到永远。
PS|29|11|耶和华必赐力量给他的百姓， 耶和华必赐平安的福给他的百姓。
PS|30|1|耶和华啊，我要尊崇你， 因为你救了我，不让仇敌向我夸耀。
PS|30|2|耶和华－我的上帝啊， 我呼求你，你医治了我。
PS|30|3|耶和华啊，你救我的性命脱离阴间， 使我存活，不至于下入地府。
PS|30|4|耶和华的圣民哪，你们要歌颂他， 要颂扬他神圣的名字 。
PS|30|5|因为，他的怒气不过是转眼之间； 他的恩典乃是一生之久。 一宿虽然有哭泣， 早晨便必欢呼。
PS|30|6|至于我，我凡事顺利，就说： “我永不动摇。”
PS|30|7|耶和华啊，你曾施恩，使我稳固如山； 你转脸不顾，我就惊惶。
PS|30|8|耶和华啊，我曾求告你； 我向耶和华恳求：
PS|30|9|“我被害流血，下到地府，有何益处呢？ 尘土岂能称谢你、传扬你的信实吗？
PS|30|10|耶和华啊，求你应允我，怜悯我！ 耶和华啊，求你帮助我！”
PS|30|11|你将我的哀哭变为跳舞， 脱去我的麻衣，为我披上喜乐，
PS|30|12|使我的灵 歌颂你，不致缄默。 耶和华－我的上帝啊，我要称谢你，直到永远！
PS|31|1|耶和华啊，我投靠你， 求你使我永不羞愧， 凭你的公义搭救我！
PS|31|2|求你侧耳听我， 快快救我！ 求你作我坚固的磐石， 拯救我的保障！
PS|31|3|你真是我的岩石、我的山寨， 求你为你名的缘故引导我，指教我。
PS|31|4|求你救我脱离人为我暗设的网罗， 因为你是我的保障。
PS|31|5|我将我的灵交在你手里； 耶和华─信实的上帝啊，你救赎了我。
PS|31|6|我 恨恶那信奉虚无神明 的人； 我却倚靠耶和华。
PS|31|7|我要因你的慈爱欢喜快乐， 因为你见过我的困苦， 知道我心中的艰难。
PS|31|8|你未曾把我交在仇敌手里， 你使我的脚站在宽阔的地方。
PS|31|9|耶和华啊，求你怜悯我， 因为我在急难之中； 我的眼睛因忧愁而昏花， 我的身心也已耗尽。
PS|31|10|我的生命为愁苦所消耗， 我的年岁为叹息所荒废； 我的力量因我的罪孽 衰败， 我的骨头也枯干。
PS|31|11|我因所有的敌人成了羞辱， 在我邻舍跟前更加羞辱； 那认识我的都惧怕我， 在街上看见我的都躲避我。
PS|31|12|我被遗忘，如同死人，无人记念； 我好像破碎的器皿。
PS|31|13|我听见许多人的毁谤， 四围尽是惊吓； 他们一同商议攻击我， 图谋害我的性命。
PS|31|14|耶和华啊，我仍要倚靠你； 我说：“你是我的上帝。”
PS|31|15|我终生的事在你手中， 求你救我脱离仇敌的手和那些迫害我的人。
PS|31|16|求你使你的脸向仆人发光， 凭你的慈爱拯救我。
PS|31|17|耶和华啊，求你叫我不致羞愧， 因为我曾呼求你； 求你使恶人羞愧， 使他们在阴间缄默无声。
PS|31|18|那撒谎的人逞骄傲轻慢， 出狂妄的话攻击义人， 愿他的嘴哑而无言。
PS|31|19|在世人眼前， 你为敬畏你的人所积存的， 为投靠你的人所施行的， 是何等大的恩惠啊！
PS|31|20|你必将他们藏在你面前的隐密处， 免得遭人暗算； 你要隐藏他们在棚子里， 免受口舌的争闹。
PS|31|21|耶和华是应当称颂的， 因为我在围城里，他向我施展奇妙的慈爱。
PS|31|22|至于我，我曾惊惶地说： “我从你眼前被隔绝。” 然而，我呼求你的时候， 你仍听我恳求的声音。
PS|31|23|耶和华的圣民哪，你们都要爱他！ 耶和华保护诚实可靠的人， 却加倍报应行事骄傲的人。
PS|31|24|凡仰望耶和华的人， 你们都要壮胆，坚固你们的心！
PS|32|1|过犯得赦免， 罪恶蒙遮盖的人有福了！
PS|32|2|耶和华不算为有罪， 内心没有诡诈的人有福了！
PS|32|3|我闭口不认罪的时候， 因终日呻吟而骨头枯干。
PS|32|4|黑夜白日，你的手压在我身上沉重； 我的精力耗尽 ，如同夏天的干旱。（细拉）
PS|32|5|我向你陈明我的罪， 不隐瞒我的恶。 我说：“我要向耶和华承认我的过犯”； 你就赦免我的罪恶。（细拉）
PS|32|6|为此，凡虔诚人都当趁你可寻找 的时候向你祷告； 大水泛滥的时候，必不临到他。
PS|32|7|你是我藏身之处， 你必保佑我脱离苦难， 以得救的欢呼 四面环绕我。（细拉）
PS|32|8|我要教导你，指示你当行的路， 我要定睛在你身上劝戒你。
PS|32|9|你不可像那无知的骡马， 须用嚼环缰绳勒住， 不然，它就不会靠近你。
PS|32|10|恶人必多受苦楚； 惟独倚靠耶和华的，必有慈爱四面环绕他。
PS|32|11|义人哪，你们应当靠耶和华欢喜快乐， 心里正直的人哪，你们都当欢呼。
PS|33|1|义人哪，你们当因耶和华欢呼， 正直人理当赞美耶和华。
PS|33|2|你们要弹琴称谢耶和华， 用十弦瑟歌颂他。
PS|33|3|应当向他唱新歌， 弹得巧妙，声音洪亮。
PS|33|4|因为耶和华的言语正直， 他的作为尽都信实。
PS|33|5|他喜爱公义和公平， 遍地满了耶和华的慈爱。
PS|33|6|诸天藉耶和华的话而造， 万象藉他口中的气而成。
PS|33|7|他聚集海水如垒， 收藏深洋在仓库。
PS|33|8|愿全地都敬畏耶和华！ 愿世上的居民都惧怕他！
PS|33|9|因为他说有，就有， 命立，就立。
PS|33|10|耶和华使列国的筹算归于无有， 使万民的计谋全无功效。
PS|33|11|耶和华的筹算永远立定， 他心中的计划万代长存。
PS|33|12|以耶和华为上帝的，那国有福了！ 耶和华拣选为自己产业的，那民有福了！
PS|33|13|耶和华从天上观看， 看见所有的人，
PS|33|14|从他的居所察看地上每一个居民，
PS|33|15|他塑造他们的心， 洞察他们一切的作为。
PS|33|16|君王不能因兵多得胜， 勇士不能因力大得救。
PS|33|17|靠马得救是枉然的， 马也不能因力大救人。
PS|33|18|看哪，耶和华的眼目看顾敬畏他的人 和仰望他慈爱的人，
PS|33|19|要救他们的性命脱离死亡， 使他们在饥荒中存活。
PS|33|20|我们的心向来等候耶和华； 他是我们的帮助，是我们的盾牌。
PS|33|21|我们的心必靠他欢喜， 因为我们向来倚靠他的圣名。
PS|33|22|耶和华啊，求你照着我们所仰望你的， 向我们施行慈爱！
PS|34|1|我要时时称颂耶和华， 赞美他的话常在我口中。
PS|34|2|我的心必因耶和华夸耀， 谦卑的人听见就喜乐。
PS|34|3|你们要和我一同尊耶和华为大， 让我们一同高举他的名。
PS|34|4|我曾寻求耶和华，他就应允我， 救我脱离一切的恐惧。
PS|34|5|仰望他的人，就有光荣； 他们 的脸必不蒙羞。
PS|34|6|这困苦人呼求，耶和华就垂听， 救他脱离一切的患难。
PS|34|7|耶和华的使者在敬畏他的人四围安营， 要搭救他们。
PS|34|8|你们要尝尝主恩的滋味，便知道他是美善； 投靠他的人有福了！
PS|34|9|耶和华的圣民哪，你们当敬畏他， 因敬畏他的一无所缺。
PS|34|10|少壮狮子尚且缺食忍饿， 但寻求耶和华的什么好处都不缺。
PS|34|11|孩子们哪，来听我！ 我要将敬畏耶和华的道教导你们。
PS|34|12|有谁喜爱生命， 爱慕长寿，得享美福？
PS|34|13|你要禁止舌头不出恶言， 嘴唇不说诡诈的话。
PS|34|14|要弃恶行善， 寻求和睦，一心追求。
PS|34|15|耶和华的眼目看顾义人， 他的耳朵听他们的呼求。
PS|34|16|耶和华向行恶的人变脸， 要从地上除灭他们的名字 。
PS|34|17|义人呼求，耶和华听见了， 就拯救他们脱离一切患难。
PS|34|18|耶和华靠近伤心的人， 拯救心灵痛悔的人。
PS|34|19|义人多有苦难， 但耶和华救他脱离这一切，
PS|34|20|又保护他全身的骨头， 连一根也不折断。
PS|34|21|恶必害死恶人， 恨恶义人的，必被定罪。
PS|34|22|耶和华救赎他仆人的性命， 凡投靠他的，必不致定罪。
PS|35|1|耶和华啊，与我相争的，求你与他们相争！ 与我争战的，求你与他们争战！
PS|35|2|求你拿着大小盾牌， 起来帮助我；
PS|35|3|举起枪来，抵挡那追赶我的。 求你对我说：“我是拯救你的。”
PS|35|4|愿那寻索我命的，蒙羞受辱！ 愿那谋害我的，退后羞愧！
PS|35|5|愿他们像风前的糠秕， 有耶和华的使者赶逐他们。
PS|35|6|愿他们的道路又暗又滑， 有耶和华的使者追赶他们。
PS|35|7|因他们无故为我暗设网罗， 无故挖坑，要害我的命。
PS|35|8|愿灾祸忽然临到他身上！ 愿他暗设的网罗缠住自己！ 愿他落在其中遭灾祸！
PS|35|9|我的心必靠耶和华快乐， 靠他的救恩欢喜。
PS|35|10|我全身的骨头要说： “耶和华啊，谁能像你 救护困苦人脱离那比他强壮的， 救护困苦贫穷人脱离那抢夺他的？”
PS|35|11|凶恶的见证人起来， 盘问我所不知道的事。
PS|35|12|他们向我以恶报善， 使我丧失儿子。
PS|35|13|至于我，他们有病的时候， 我穿麻衣，禁食，刻苦己心； 我所求的都归到自己身上。
PS|35|14|我如此行，好像他是我的朋友，我的兄弟； 我屈身悲哀，如同哀悼自己的母亲。
PS|35|15|我在患难中，他们却欢喜，大家聚集， 我所不认识的卑贱人 聚集攻击我， 他们不住地撕裂我。
PS|35|16|他们试探我，不断嘲笑我 ， 向我咬牙切齿。
PS|35|17|主啊，你看着不理要到几时呢？ 求你救我的性命脱离他们的残害， 救我仅有的 脱离少壮狮子！
PS|35|18|我在大会中要称谢你， 在许多百姓中要赞美你。
PS|35|19|求你不容那无理与我为仇的向我夸耀！ 不容那无故恨我的向我瞪眼！
PS|35|20|因为他们不说平安， 倒想出诡诈的言语扰害地上安静的人。
PS|35|21|他们大大张口攻击我，说： “啊哈，啊哈，我们已经亲眼看见了！”
PS|35|22|耶和华啊，你已经看见了，求你不要沉默！ 主啊，求你不要远离我！
PS|35|23|我的上帝─我的主啊，求你醒来，求你奋起， 还我公正，伸明我冤！
PS|35|24|耶和华－我的上帝啊，求你按你的公义判断我， 不容他们向我夸耀！
PS|35|25|不容他们心里说：“啊哈，遂我们的心愿了！” 不容他们说：“我们已经把他吞了！”
PS|35|26|愿那喜欢我遭难的一同抱愧蒙羞！ 愿那向我妄自尊大的披戴惭愧，蒙受羞辱！
PS|35|27|愿那喜悦我被判为义 的欢呼快乐； 愿他们常说：“当尊耶和华为大！ 耶和华喜悦他的仆人平安。”
PS|35|28|我的舌头要论说你的公义， 要常常赞美你。
PS|36|1|过犯在恶人的心底向他说话 ， 他的眼中不怕上帝。
PS|36|2|他自夸自媚， 以致罪孽无法察觉，不被恨恶。
PS|36|3|他口中的言语尽是罪孽诡诈， 他不再有智慧，也不再行善。
PS|36|4|他在床上图谋罪孽， 定意行不善的道，不憎恶恶事。
PS|36|5|耶和华啊，你的慈爱上及诸天， 你的信实达到穹苍，
PS|36|6|你的公义好像高山， 你的判断如同深渊； 耶和华啊，人民、牲畜，你都救护。
PS|36|7|上帝啊，你的慈爱何其宝贵！ 世人投靠在你翅膀的荫下。
PS|36|8|他们必因你殿里的丰盛得以饱足， 你也必叫他们喝你那喜乐的泉水。
PS|36|9|因为在你那里有生命的泉源， 在你的光中，我们必得见光。
PS|36|10|愿你常施慈爱给认识你的人， 常以公义待心里正直的人。
PS|36|11|不容骄傲人的脚践踏我， 不容凶恶人的手赶逐我。
PS|36|12|在那里，作恶的人已经仆倒； 他们被推倒，不能再起来。
PS|37|1|不要为作恶的心怀不平， 也不要嫉妒那行不义的人。
PS|37|2|因为他们如草快被割下， 又如绿色的嫩草快要枯干。
PS|37|3|你当倚靠耶和华而行善， 安居地上，以他的信实为粮；
PS|37|4|又当以耶和华为乐， 他就将你心里所求的赐给你。
PS|37|5|当将你的道路交托耶和华， 并倚靠他，他就必成全。
PS|37|6|他要使你的公义如光发出， 使你的公平明如正午。
PS|37|7|你当安心倚靠耶和华，耐性等候他， 不要因那道路通达的和那恶谋成就的心怀不平。
PS|37|8|当止住怒气，离弃愤怒； 不要心怀不平，以致作恶。
PS|37|9|因为作恶的必被剪除； 惟有等候耶和华的必承受土地。
PS|37|10|还有片时，恶人要归于无有； 你就是细察他的住处，也不存在。
PS|37|11|但谦卑的人必承受土地， 以丰盛的平安为乐。
PS|37|12|恶人设谋要害义人， 向他咬牙。
PS|37|13|但主必笑他， 因见他受罚的日子将要来到。
PS|37|14|恶人刀已出鞘，弓已上弦， 要砍倒困苦贫穷的人， 要杀害行为正直的人。
PS|37|15|他们的刀必刺入自己的心， 他们的弓必折断。
PS|37|16|一个义人所有的虽少， 强过许多恶人的富余。
PS|37|17|因为恶人的膀臂必折断； 但耶和华扶持义人。
PS|37|18|耶和华知道完全人的日子， 他们的产业要存到永远。
PS|37|19|他们在患难的时候必不致羞愧， 在饥荒的日子必得饱足。
PS|37|20|恶人却要灭亡。 耶和华的仇敌要像草地的华美 ； 他们要毁灭，在烟中消失 。
PS|37|21|恶人借贷却不偿还； 义人恩待人，并且施舍。
PS|37|22|蒙耶和华赐福的必承受土地； 他所诅咒的必被剪除。
PS|37|23|义人的脚步为耶和华所稳定； 他的道路，耶和华也喜爱。
PS|37|24|他虽失脚也不致全身仆倒， 因为耶和华搀扶他的手。
PS|37|25|我从前年幼，现在年老， 却未见过义人被弃， 也未见过他的后裔求乞。
PS|37|26|他常常恩待人，借贷给人， 他的后裔也必蒙福。
PS|37|27|你当离恶行善， 就可永远安居。
PS|37|28|因为耶和华喜爱公平， 不撇弃他的圣民， 他们永蒙保佑； 但恶人的后裔必被剪除。
PS|37|29|义人必承受土地， 永居其上。
PS|37|30|义人的口发出智慧， 他的舌头讲说公平。
PS|37|31|上帝的律法在他心里， 他的步伐总不摇动。
PS|37|32|恶人窥探义人， 想要杀他。
PS|37|33|耶和华必不把他交在恶人手中， 当审判的时候，也不定他的罪。
PS|37|34|你当等候耶和华，遵守他的道， 他就抬举你，使你承受土地； 你必看到恶人被剪除。
PS|37|35|我见过恶人大有势力， 高耸如本地青翠的树木。
PS|37|36|有人 从那里经过，看哪，他已不存在， 我寻找他，却寻不着了。
PS|37|37|你要细察那完全人，观看那正直人， 因为和平的人有好结局。
PS|37|38|至于罪人，必一同灭绝， 恶人的结局必被剪除。
PS|37|39|义人得救是出于耶和华， 在患难时耶和华作他们的避难所。
PS|37|40|耶和华帮助他们，解救他们； 他解救他们脱离恶人，把他们救出来， 因为他们投靠他。
PS|38|1|耶和华啊，求你不要在怒中责备我， 不要在烈怒中惩罚我！
PS|38|2|因为你的箭射入我身， 你的手压住我。
PS|38|3|因你的恼怒，我的肉无一完全； 因我的罪过，我的骨头也不安宁。
PS|38|4|我的罪孽高过我的头， 如同重担叫我担当不起。
PS|38|5|因我的愚昧， 我的伤发臭流脓。
PS|38|6|我疼痛，大大蜷曲， 整日哀痛。
PS|38|7|我满腰灼热， 我的肉无一完全。
PS|38|8|我被压碎，身心虚弱； 因心里痛苦，我就呻吟。
PS|38|9|主啊，我的心愿都在你面前， 我的叹息不向你隐瞒。
PS|38|10|我心颤栗，体力衰微， 眼中无光。
PS|38|11|我遭遇灾病，良朋密友都袖手旁观， 我的亲戚本家也远远站立。
PS|38|12|那寻索我命的设下罗网， 那想要害我的口出恶言， 整日思想诡计。
PS|38|13|但我如聋子听不见， 像哑巴不能开口。
PS|38|14|我如听不见的人， 无法用口答辩。
PS|38|15|耶和华啊，我仰望你！ 主－我的上帝啊，你必应允我！
PS|38|16|我曾说：“恐怕他们向我夸耀， 我失脚的时候，他们向我夸口。”
PS|38|17|我就要跌倒， 我的痛苦常在我面前。
PS|38|18|我要承认我的罪孽， 要因我的罪忧愁。
PS|38|19|但我的仇敌又活泼又强壮， 无理恨我的增多了。
PS|38|20|以恶报善的与我作对， 但我追求良善。
PS|38|21|耶和华啊，求你不要撇弃我！ 我的上帝啊，求你不要远离我！
PS|38|22|拯救我的主啊， 求你快快帮助我！
PS|39|1|我曾说：“我要谨慎我的言行， 免得我的舌头犯罪； 恶人在我面前的时候， 我要用嚼环勒住我的口。”
PS|39|2|我默然无声，连好话也不出口， 我的愁苦就更加深。
PS|39|3|我的心在我里面发热； 我默想的时候，火就烧起， 我用舌头说话：
PS|39|4|“耶和华啊，求你让我晓得我的结局， 我的寿数几何， 使我知道我的生命何等短暂！
PS|39|5|看哪，你使我的年日窄如手掌， 我一生的年数，在你面前如同无有； 各人最稳妥的时候，真是全然虚幻。（细拉）
PS|39|6|世人行动实系幻影， 他们忙乱，真是枉然， 积蓄财宝，不知将来有谁收取。
PS|39|7|“主啊，如今我等什么呢？ 我的指望在乎你！
PS|39|8|求你救我脱离一切的过犯， 不要使我受愚顽人的羞辱。
PS|39|9|我保持沉默，闭口不言， 因为这一切都是你所做的。
PS|39|10|求你从我身上免去你的责罚； 因你手的责打，我就消灭。
PS|39|11|因人的罪恶你惩罚管教他的时候， 如蛀虫一般，吃掉他所喜爱的。 世人真是虚幻！（细拉）
PS|39|12|“耶和华啊，求你听我的祷告， 侧耳听我的呼求！ 我流泪，求你不要静默无声！ 因为在你面前我是客旅， 是寄居的，像我列祖一般。
PS|39|13|求你宽容我， 使我在去而不返之先可以喜乐。”
PS|40|1|我曾耐性等候耶和华， 他垂听我的呼求。
PS|40|2|他从泥坑里， 从淤泥中，把我拉上来， 使我的脚立在磐石上， 使我脚步稳健。
PS|40|3|他使我口唱新歌， 就是赞美我们上帝的话。 许多人必看见而惧怕， 并要倚靠耶和华。
PS|40|4|那倚靠耶和华、 不理会狂傲和偏向虚假的， 这人有福了！
PS|40|5|耶和华－我的上帝啊，你所行的奇事 和你为我们设想的计划，多到无法尽述； 若要述说陈明，不可胜数。
PS|40|6|祭物和礼物，你不喜爱， 你已经开通我的耳朵； 燔祭和赎罪祭非你所要。
PS|40|7|那时我说：“看哪，我来了！ 我的事在经卷上已经记载了。
PS|40|8|我的上帝啊，我乐意照你的旨意行， 你的律法在我心里。”
PS|40|9|我在大会中传讲公义的佳音， 看哪，必不制止我的嘴唇； 耶和华啊，这一切你都知道。
PS|40|10|我未曾把你的公义藏在心里， 我已陈明你的信实和你的救恩； 在大会中我未曾隐瞒你的慈爱和信实。
PS|40|11|耶和华啊，求你不要向我止住你的怜悯！ 愿你的慈爱和信实常常保佑我！
PS|40|12|因有无数的祸患围困我， 我的罪孽追上了我，使我不能看见， 这罪孽比我的头发还多， 我的胆量丧失了。
PS|40|13|耶和华啊，求你开恩搭救我！ 耶和华啊，求你速速帮助我！
PS|40|14|愿那些寻找我、要灭我命的，一同抱愧蒙羞！ 愿那些喜悦我遭害的，退后受辱！
PS|40|15|愿那些对我说“啊哈、啊哈”的， 因羞愧而败亡！
PS|40|16|愿一切寻求你的，因你欢喜快乐！ 愿那些喜爱你救恩的，常说：“当尊耶和华为大！”
PS|40|17|我本是困苦贫穷的，主却顾念我。 你是帮助我的，搭救我的； 我的上帝啊，求你不要耽延！
PS|41|1|眷顾贫寒人的有福了 ！ 在患难的日子，耶和华必搭救他。
PS|41|2|耶和华必保全他，使他存活， 他要在地上享福。 求你不要把他交给仇敌，遂其所愿。
PS|41|3|他病重在榻，耶和华必扶持他； 他在病中，你必使他离开病床。
PS|41|4|我曾说：“耶和华啊，求你怜悯我， 医治我，因为我得罪了你。”
PS|41|5|我的仇敌用恶言议论我： “他几时才会死，他的名几时才会消灭呢？”
PS|41|6|当他来看我的时候，说的是假话； 他心存奸恶，走到外边才说出来。
PS|41|7|所有恨我的，都一同交头接耳议论我， 他们设计要害我。
PS|41|8|他们说：“他有怪病缠身， 他已躺下，必不能再起来。”
PS|41|9|连我知己的朋友， 我所信赖、吃我饭的人也用脚踢我。
PS|41|10|耶和华啊，求你怜悯我， 使我起来，好报复他们！
PS|41|11|我因此就知道你喜爱我， 我的仇敌不得向我夸胜。
PS|41|12|你因我纯正就扶持我， 使我永远站立在你面前。
PS|41|13|耶和华－ 以色列 的上帝是应当称颂的， 从亘古直到永远。阿们！阿们！ 可拉后裔的诗。交给圣咏团长。
PS|42|1|上帝啊，我的心切慕你， 如鹿切慕溪水。
PS|42|2|我的心渴想上帝，就是永生上帝， 我几时得朝见上帝呢？
PS|42|3|我昼夜以眼泪当食物， 人不住地对我说：“你的上帝在哪里呢？”
PS|42|4|我从前与众人同往， 领他们到上帝的殿里， 大家用欢呼称颂的声音守节； 我追想这些事， 我的心极其悲伤。
PS|42|5|我的心哪，你为何忧闷？ 为何在我里面烦躁？ 应当仰望上帝， 因我还要称谢他，我当面的拯救，
PS|42|6|我的上帝。我的心在我里面忧闷， 所以我从 约旦 地， 从 黑门岭 ，从 米萨山 记念你。
PS|42|7|你的瀑布发声，深渊就与深渊响应， 你的波浪洪涛漫过我身。
PS|42|8|白昼，耶和华必施慈爱； 黑夜，我要歌颂祈祷赐我生命的上帝。
PS|42|9|我要对上帝－我的磐石说： “你为何忘记我呢？ 我为何因仇敌的欺压时常哀痛呢？”
PS|42|10|我的敌人辱骂我， 好像敲碎我的骨头， 他们不住地对我说： “你的上帝在哪里呢？”
PS|42|11|我的心哪，你为何忧闷？ 为何在我里面烦躁？ 应当仰望上帝， 因我还要称谢他，我当面的拯救，我的上帝。
PS|43|1|上帝啊，求你为我伸冤， 向不虔诚的国为我辩护； 求你救我脱离诡诈不义的人。
PS|43|2|你是作我保障 的上帝，为何丢弃我呢？ 我为何因仇敌的欺压时常哀痛呢？
PS|43|3|求你发出你的亮光和信实，好引导我， 带我到你的圣山，到你的居所！
PS|43|4|我就走到上帝的祭坛， 到赐我喜乐的上帝那里。 上帝，我的上帝啊， 我要弹琴称谢你！
PS|43|5|我的心哪，你为何忧闷？ 为何在我里面烦躁？ 应当仰望上帝， 我还要称谢他，我当面的拯救，我的上帝。
PS|44|1|上帝啊，你在古时， 我们列祖的日子所做的事， 我们亲耳听见了， 我们的列祖曾为我们述说。
PS|44|2|你曾用手赶出外邦人， 却栽培了我们的列祖； 你苦待万民， 却叫我们的列祖发达。
PS|44|3|因为他们不是靠自己的刀剑承受土地， 也不是靠自己的膀臂得胜， 而是靠你的右手、你的膀臂， 和你脸上的亮光， 因为你喜爱他们。
PS|44|4|上帝啊，你是我的君王， 求你发命令使 雅各 得胜。
PS|44|5|靠你，我们要推倒我们的敌人； 靠你的名，我们要践踏那兴起攻击我们的人。
PS|44|6|因为我必不倚靠我的弓， 我的刀也不能使我得胜。
PS|44|7|惟有你拯救我们脱离敌人， 使恨我们的人羞愧。
PS|44|8|我们要常常因上帝夸耀， 要永远颂扬你的名。（细拉）
PS|44|9|但如今你丢弃了我们，使我们受辱， 不和我们的军队同去。
PS|44|10|你使我们在敌人前转身撤退， 使那恨我们的人任意抢夺。
PS|44|11|你使我们如羊当作食物， 把我们分散在列国中。
PS|44|12|你卖了你的子民也不获利， 所得的并未加添你的资财。
PS|44|13|你使我们受邻国的羞辱， 被四围的人嗤笑讥讽。
PS|44|14|你使我们在列国中成了笑柄， 在万民中使人摇头。
PS|44|15|因辱骂者和毁谤者的声音， 因仇敌和报仇者的缘故， 我的凌辱常常在我面前， 我脸上的羞愧将我遮蔽，
PS|44|16|
PS|44|17|这些事都临到我们身上， 我们却没有忘记你， 也没有违背你的约；
PS|44|18|我们的心并未退缩， 我们的脚也没有偏离你的路。
PS|44|19|你在野狗出没之处压伤我们， 以死荫笼罩我们。
PS|44|20|倘若我们忘记上帝的名， 或向外邦神明举手，
PS|44|21|上帝岂不鉴察这事吗？ 因为他晓得人心里的隐秘。
PS|44|22|我们为你的缘故终日被杀， 人看我们如将宰的羊。
PS|44|23|主啊，求你睡醒，为何尽睡呢？ 求你醒来，不要永远丢弃我们！
PS|44|24|你为何转脸， 不顾我们所遭的苦难和所受的欺压呢？
PS|44|25|我们俯伏在尘土上， 我们的肚腹紧贴地面。
PS|44|26|求你兴起帮助我们！ 因你的慈爱救赎我们！
PS|45|1|我心里涌出美辞， 我为王朗诵我的诗章， 我的舌头是敏捷文士的手笔。
PS|45|2|你比世人更美， 你嘴里满有恩惠； 所以上帝赐福给你，直到永远。
PS|45|3|勇士啊，愿你腰间佩刀， 大展荣耀和威严，
PS|45|4|为真理、谦卑、公义威严地驾车前进，无不得胜； 愿你的右手显明可畏的事。
PS|45|5|你的箭锋快，射中王的仇敌的心， 万民仆倒在你之下。
PS|45|6|上帝啊，你的宝座是永永远远的， 你国度的权杖是正直的权杖。
PS|45|7|你喜爱公义，恨恶罪恶， 所以上帝，就是你的上帝，用喜乐油膏你， 胜过膏你的同伴。
PS|45|8|你的衣服散发没药、沉香、肉桂的香气， 象牙宫中丝弦乐器的声音使你欢喜。
PS|45|9|你的妃嫔之中有列王的女儿， 王后佩戴 俄斐 金饰站立在你右边。
PS|45|10|女子啊，要倾听，要思想，要侧耳而听！ 不要记念你本族和你父家，
PS|45|11|王就羡慕你的美貌； 因为他是你的主，你当向他下拜。
PS|45|12|推罗 必来送礼， 百姓中富足的人也必向你求恩。
PS|45|13|君王的女儿在宫里极其荣华， 她的衣服是金线绣的；
PS|45|14|她穿锦绣的衣服，引到王面前， 陪伴她的童女随从她，也被带到你面前。
PS|45|15|她们要欢喜快乐， 被引导进入王宫。
PS|45|16|你的子孙要接续你列祖， 你要立他们在各地作王。
PS|45|17|我必使万代记念你的名， 万民要永永远远称谢你。
PS|46|1|上帝是我们的避难所，是我们的力量， 是我们在患难中随时的帮助。
PS|46|2|所以，地虽改变， 山虽摇动到海心，
PS|46|3|其中的水虽澎湃翻腾， 山虽因海涨而战抖， 我们也不害怕。（细拉）
PS|46|4|有一道河，这河的分汊使上帝的城欢喜， 这城就是至高者居住的圣所。
PS|46|5|上帝在其中，城必不动摇； 到天一亮，上帝必帮助这城。
PS|46|6|万邦喧嚷，国度动摇； 上帝出声，地就熔化。
PS|46|7|万军之耶和华与我们同在， 雅各 的上帝是我们的避难所！（细拉）
PS|46|8|你们来看耶和华的作为， 看他使地怎样荒凉。
PS|46|9|他止息战争，直到地极； 他折弓、断枪，把战车焚烧在火中。
PS|46|10|你们要休息，要知道我是上帝！ 我必在列国中受尊崇，在全地也受尊崇。
PS|46|11|万军之耶和华与我们同在， 雅各 的上帝是我们的避难所！
PS|47|1|万民哪，你们都要鼓掌！ 用欢呼的声音向上帝呼喊！
PS|47|2|因为耶和华至高者是可畏的， 他是治理全地的大君王。
PS|47|3|他使万民服在我们以下， 又使万族服在我们脚下。
PS|47|4|他为我们选择产业， 就是他所爱之 雅各 的荣耀。（细拉）
PS|47|5|上帝上升，有喊声相送； 耶和华上升，有角声相送。
PS|47|6|你们要向上帝歌颂，歌颂！ 向我们的王歌颂，歌颂！
PS|47|7|因为上帝是全地的王， 你们要用圣诗歌颂！
PS|47|8|上帝作王治理列国， 上帝坐在他的圣宝座上。
PS|47|9|万民的君王聚集， 要作 亚伯拉罕 的上帝的子民， 因为地上的盾牌是属上帝的， 他为至高！
PS|48|1|耶和华本为大！ 在我们上帝的城中， 在他的圣山上， 当受大赞美。
PS|48|2|锡安山 －大君王的城， 在北面居高华美， 为全地所喜悦。
PS|48|3|上帝在城的宫殿中， 自显为避难所。
PS|48|4|看哪，诸王会合， 一同经过。
PS|48|5|他们见了这城就惊奇丧胆， 急忙逃跑。
PS|48|6|战兢在那里抓住他们， 他们好像临产的妇人一样阵痛。
PS|48|7|上帝啊，你用东风击破 他施 的船只。
PS|48|8|我们在万军之耶和华的城里， 就是我们上帝的城里， 所看见的正如我们所听见的。 上帝必坚立这城，直到永远。（细拉）
PS|48|9|上帝啊，我们在你的殿中 想念你的慈爱。
PS|48|10|上帝啊，你受的赞美正与你的名相称，直到地极！ 你的右手满了公义。
PS|48|11|因你的判断， 锡安山 应当欢喜， 犹大 的城镇 应当快乐。
PS|48|12|你们当周游 锡安 ， 四围环绕，数点城楼，
PS|48|13|细看它的城郭， 察看它的宫殿， 为要传扬给后代。
PS|48|14|因为这上帝永永远远为我们的上帝， 他必作我们引路的，直到死时 。
PS|49|1|万民哪，你们都当听这话！ 世上所有的居民， 无论贵贱贫富， 都当侧耳而听！
PS|49|2|
PS|49|3|我口要说智慧的言语， 我心思想通达的道理。
PS|49|4|我要侧耳听比喻， 用琴解谜语。
PS|49|5|在患难的日子，追逼我的人的奸恶 环绕我， 我何必惧怕？
PS|49|6|他们那些倚靠财货， 自夸钱财多的人，
PS|49|7|没有一个能赎自己的弟兄 ， 能将赎价给上帝，
PS|49|8|让他长远活着，不见地府 ； 因为赎生命的价值极贵， 只可永远罢休。
PS|49|9|
PS|49|10|他要见智慧人死， 愚昧人和畜牲一般的人一同灭亡， 把他们的财货留给别人。
PS|49|11|他们虽以自己的名叫自己的地， 坟墓却作他们永远的家， 作他们世世代代的居所。
PS|49|12|人居尊贵中不能长久， 如同死亡的畜类一样。
PS|49|13|他们所行之道本为自己的愚昧， 后来的人却还佩服他们的话语。（细拉）
PS|49|14|他们如同羊群注定要下阴间， 死亡必作他们的牧者； 到了早晨，正直人必管辖他们。 他们的形像必被阴间所灭，无处可容身。
PS|49|15|然而上帝必救赎我的命脱离阴间的掌控， 因他必收纳我。（细拉）
PS|49|16|见人发财、家室日益显赫的时候， 你不要惧怕；
PS|49|17|因为他死的时候什么也不能带去， 他的荣耀不能随他下去。
PS|49|18|他活着的时候，虽然自夸为有福 ─你若自己行得好，人必夸奖你─
PS|49|19|他仍必与历代的祖宗一样同归死亡， 永不见光。
PS|49|20|人在尊贵中而不醒悟， 就如死亡的畜类一样。
PS|50|1|大能者上帝－耶和华已经发言呼召天下， 从日出之地到日落之处。
PS|50|2|从全然美丽的 锡安 中， 上帝已经发光了。
PS|50|3|我们的上帝要来，绝不闭口； 有烈火在他面前吞灭， 有暴风在他四围刮起。
PS|50|4|他呼召上天下地， 为要审判他的子民：
PS|50|5|“召集我的圣民， 就是那些用祭物与我立约的人，到我这里来。”
PS|50|6|诸天必表明他的公义， 因为上帝是施行审判的。（细拉）
PS|50|7|“听啊，我的子民，我要说话！ 以色列 啊，我要审问你； 我是上帝，是你的上帝！
PS|50|8|我并不因你的祭物责备你； 你的燔祭常在我面前。
PS|50|9|我不从你家中取公牛， 也不从你圈内取公山羊；
PS|50|10|因为，林中的百兽是我的， 千山的牲畜也是我的。
PS|50|11|山中 的飞鸟，我都知道， 田野的走兽也都属我。
PS|50|12|“我若是饥饿，不用告诉你， 因为世界和其中所充满的都是我的。
PS|50|13|我岂吃公牛的肉呢？ 我岂喝公山羊的血呢？
PS|50|14|你们要以感谢为祭献给上帝， 又要向至高者还你的愿，
PS|50|15|并要在患难之日求告我， 我必搭救你，你也要荣耀我。”
PS|50|16|但上帝对恶人说：“你怎敢传讲我的律例， 口中提到我的约呢？
PS|50|17|其实你恨恶管教， 将我的言语抛在脑后。
PS|50|18|你见了盗贼就乐意与他同伙， 又和行奸淫的人同流合污。
PS|50|19|“你的口出恶言， 你的舌编造诡诈。
PS|50|20|你坐着，毁谤你的兄弟， 谗害你亲母的儿子。
PS|50|21|你做了这些事，我闭口不言， 你想我正如你一样； 其实我要责备你，将这些事摆在你眼前。
PS|50|22|“你们忘记上帝的，要思想这事， 免得我把你们撕碎，无人搭救。
PS|50|23|凡以感谢献祭的就是荣耀我； 那按正路而行的，我必使他得着上帝的救恩。”
PS|51|1|上帝啊，求你按你的慈爱恩待我！ 按你丰盛的怜悯涂去我的过犯！
PS|51|2|求你将我的罪孽洗涤净尽， 洁除我的罪！
PS|51|3|因为我知道我的过犯； 我的罪常在我面前。
PS|51|4|我向你犯罪，惟独得罪了你， 在你眼前行了这恶， 以致你责备的时候显为公义， 判断的时候显为清白。
PS|51|5|看哪，我是在罪孽里生的， 在我母亲怀胎的时候就有了罪。
PS|51|6|你所喜爱的是内心的诚实； 求你在我隐密处使我得智慧。
PS|51|7|求你用牛膝草洁净我，我就干净； 求你洗涤我，我就比雪更白。
PS|51|8|求你使我得听欢喜快乐的声音， 使你所压伤的骨头可以踊跃。
PS|51|9|求你转脸不看我的罪， 涂去我一切的罪孽。
PS|51|10|上帝啊，求你为我造清洁的心， 使我里面重新有正直 的灵。
PS|51|11|不要丢弃我，使我离开你的面； 不要从我收回你的圣灵。
PS|51|12|求你使我重得救恩之乐， 以乐意的灵来扶持我，
PS|51|13|我就把你的道指教有过犯的人， 罪人必归顺你。
PS|51|14|上帝啊，你是拯救我的上帝； 求你救我脱离流人血的罪！ 我的舌头就高唱你的公义。
PS|51|15|主啊，求你使我嘴唇张开， 我的口就传扬赞美你的话！
PS|51|16|你本不喜爱祭物，若喜爱，我就献上； 燔祭你也不喜悦。
PS|51|17|上帝所要的祭就是忧伤的灵； 上帝啊，忧伤痛悔的心，你必不轻看。
PS|51|18|求你随你的美意善待 锡安 ， 建造 耶路撒冷 的城墙。
PS|51|19|那时，你必喜爱公义的祭 和燔祭，全牲的燔祭； 那时，人必将公牛献在你坛上。
PS|52|1|勇士啊，你为何作恶自夸？ 上帝的慈爱是常存的。
PS|52|2|你这行诡诈的人哪， 你的舌头像快利的剃刀，图谋毁灭。
PS|52|3|你爱恶胜似爱善， 又爱说谎，胜于爱说公义。（细拉）
PS|52|4|诡诈的舌头啊， 你爱说一切毁灭的话！
PS|52|5|上帝也要毁灭你，直到永远。 他要抓住你，从帐棚中拉你出来， 从活人之地将你拔除。（细拉）
PS|52|6|义人要看见而惧怕， 并要笑他。
PS|52|7|看哪，这就是那不以上帝为保障的人， 他只倚靠丰富的财物，在邪恶上坚立自己。
PS|52|8|至于我，就像上帝殿中的青橄榄树， 我永永远远倚靠上帝的慈爱。
PS|52|9|我要称谢你，直到永远， 因为你做了这事。 我也要在你圣民面前仰望你的名， 这名本为美好。
PS|53|1|愚顽人心里说：“没有上帝。” 他们都败坏，行了可憎恶的罪孽， 没有一个人行善。
PS|53|2|上帝从天上垂看世人， 要看有明白的没有， 有寻求上帝的没有。
PS|53|3|他们全都退后，一同变为污秽， 没有行善的， 连一个也没有。
PS|53|4|作恶的都没有知识吗？ 他们吞吃我的百姓如同吃饭一样， 并不求告上帝。
PS|53|5|他们在无可惧怕之处就大大害怕， 因为上帝使那安营攻击你之人的骨头散开了。 你使他们蒙羞，因为上帝弃绝了他们。
PS|53|6|但愿 以色列 的救恩出自 锡安 。 当上帝救回他被掳子民的时候， 雅各 要快乐， 以色列 要欢喜。
PS|54|1|上帝啊，求你因你的名拯救我， 凭你的大能为我伸冤。
PS|54|2|上帝啊，求你听我的祷告， 侧耳听我口中的言语。
PS|54|3|因为陌生人兴起攻击我， 强横的人寻索我的性命； 他们眼中没有上帝。（细拉）
PS|54|4|看哪，上帝是帮助我的， 主是扶持我性命的，
PS|54|5|他要报应我仇敌所作的恶； 求你凭你的信实灭绝他们。
PS|54|6|我要把甘心祭献给你； 耶和华啊，我要颂扬你的名，这名本为美好。
PS|54|7|他从一切的急难中把我救出来， 我的眼睛也看见了我的仇敌遭报。
PS|55|1|上帝啊，求你侧耳听我的祷告， 不要隐藏不听我的恳求！
PS|55|2|求你留心听我，应允我。 我哀叹不安，发出呻吟，
PS|55|3|都因仇敌的声音，恶人的欺压； 他们将罪孽加在我身上，发怒气加害我。
PS|55|4|我的心在我里面阵痛， 死亡的恐怖落在我身。
PS|55|5|恐惧战兢临到了我， 惊恐笼罩我。
PS|55|6|我说：“但愿我有翅膀像鸽子， 我就飞去，得享安息。
PS|55|7|看哪，我要远走高飞， 宿在旷野。（细拉）
PS|55|8|我要速速逃到避难之所， 脱离狂风暴雨。”
PS|55|9|主啊，求你吞灭他们，变乱他们的言语！ 因为我在城中见了凶暴争吵的事。
PS|55|10|他们昼夜在城墙上绕行， 城内也有罪孽和奸恶。
PS|55|11|邪恶在其中， 欺压和诡诈不离街市。
PS|55|12|原来，不是仇敌辱骂我， 若是仇敌，还可忍受； 也不是恨我的人向我狂妄自大， 若是恨我的人，我必躲避他。
PS|55|13|不料是你；你原与我同等， 是我的朋友，是我的知己！
PS|55|14|我们素常彼此交谈，以为甘甜； 我们结伴在上帝的殿中同行。
PS|55|15|愿死亡忽然临到他们！ 愿他们活生生地下入阴间！ 因为他们的住处都是邪恶， 他们的内心充满奸恶。
PS|55|16|至于我，我要求告上帝， 耶和华必拯救我。
PS|55|17|晚上、早晨、中午我要哀声悲叹， 他就垂听我的声音。
PS|55|18|他救赎我的命脱离攻击我的人， 使我得享平安， 因为与我相争的人很多。
PS|55|19|那不愿改变、不敬畏上帝的人， 从太古常存的上帝必听见而使他受苦。（细拉）
PS|55|20|他背了约， 伸手攻击与他和好的人。
PS|55|21|他的口如奶油光滑， 他的心却怀着敌意； 他的话比油柔和， 其实是拔出的刀。
PS|55|22|你要把你的重担卸给耶和华， 他必扶持你， 他永不叫义人动摇。
PS|55|23|上帝啊，你必使恶人坠入灭亡的坑； 那好流人血、行诡诈的人必活不过半生， 但我要倚靠你。
PS|56|1|上帝啊，求你怜悯我，因为有人践踏我， 终日攻击欺压我。
PS|56|2|我的仇敌终日践踏我， 逞骄傲攻击我的人很多。
PS|56|3|我惧怕的时候要倚靠你。
PS|56|4|我倚靠上帝，我要赞美他的话语； 我倚靠上帝，必不惧怕。 血肉之躯能把我怎么样呢？
PS|56|5|他们终日扭曲我的话， 千方百计加害于我。
PS|56|6|他们聚集，埋伏，窥探我的脚踪， 等候要害我的命。
PS|56|7|他们岂能脱罪呢 ？ 上帝啊，求你在怒中使万民败落！
PS|56|8|我几次流离，你都数算； 求你把我的眼泪装在你的皮袋里。 这一切不都记在你的册子上吗？
PS|56|9|我呼求的日子，仇敌都要转身撤退。 上帝帮助我，这是我所知道的。
PS|56|10|我倚靠上帝，我要赞美他的话语； 我倚靠耶和华，我要赞美他的话语。
PS|56|11|我倚靠上帝，必不惧怕。 人能把我怎么样呢？
PS|56|12|上帝啊，我要向你还所许的愿， 我要以感谢祭回报你；
PS|56|13|因为你救我的命脱离死亡。 你保护我的脚不跌倒， 使我在生命的光中行在上帝面前。
PS|57|1|上帝啊，求你怜悯我，怜悯我， 因为我的心投靠你。 我要投靠在你翅膀荫下， 直等到灾害过去。
PS|57|2|我要求告至高的上帝， 就是为我成全万事的上帝。
PS|57|3|那践踏我的人辱骂我的时候， 上帝必从天上施恩救我，(细拉) 他必向我施行慈爱和信实。
PS|57|4|至于我的性命， 我好像躺卧在吞噬人的狮子当中； 他们的牙齿是枪、箭， 他们的舌头是快刀。
PS|57|5|上帝啊，愿你崇高过于诸天！ 愿你的荣耀高过全地！
PS|57|6|他们为我的脚设下网罗，压迫我； 他们在我面前掘了坑，自己反掉在其中。（细拉）
PS|57|7|上帝啊，我心坚定，我心坚定； 我要唱诗，我要歌颂！
PS|57|8|我的灵 啊，你当醒起！ 琴瑟啊，当醒起！ 我自己要极早醒起！
PS|57|9|主啊，我要在万民中称谢你， 在万族中歌颂你！
PS|57|10|因为你的慈爱高及诸天， 你的信实达到穹苍。
PS|57|11|上帝啊，愿你崇高过于诸天！ 愿你的荣耀高过全地！
PS|58|1|你们缄默不语，真合公义吗？ 你们审判世人，岂按正直吗？
PS|58|2|不然！你们心中作恶， 量出你们在地上手中的残暴。
PS|58|3|恶人一出母胎就与上帝疏远， 一离母腹就走错路，说谎话。
PS|58|4|他们的毒气好像蛇的毒气， 他们好像聋的毒蛇塞住耳朵，
PS|58|5|听不见弄蛇者的声音， 也听不见魔术师的咒语。
PS|58|6|上帝啊，求你敲碎他们口中的牙！ 耶和华啊，求你敲掉少壮狮子的大牙！
PS|58|7|愿他们消灭，如急流的水一般； 他们瞄准射箭的时候，箭头仿佛折断。
PS|58|8|愿他们像蜗牛腐烂消失， 又像妇人流掉的胎儿，未见天日。
PS|58|9|你们用荆棘烧火，锅还未热， 上帝就用旋风把未烧着的和已烧着的一齐刮去。
PS|58|10|义人见仇敌遭报就欢喜， 他要在恶人的血中洗脚。
PS|58|11|因此，人必说：“义人诚然有善报， 在地上果然有施行审判的上帝！”
PS|59|1|我的上帝啊，求你救我脱离仇敌， 把我安置在高处，脱离那些起来攻击我的人。
PS|59|2|求你救我脱离作恶的人， 救我脱离好流人血的人！
PS|59|3|因为他们埋伏要害我命， 强悍的人聚集攻击我， 耶和华啊，不是为我的过犯， 也不是为我的罪愆。
PS|59|4|我虽然无过，他们急忙摆阵攻击我。 求你兴起，来帮助我，来鉴察！
PS|59|5|万军之耶和华上帝－ 以色列 的上帝啊， 求你醒起，惩治万国！ 不要怜悯行诡诈的恶人！（细拉）
PS|59|6|他们晚上转回， 叫号如狗，围城绕行。
PS|59|7|看哪，他们口中喷吐恶言， 嘴里有刀： “有谁听见呢？”
PS|59|8|但你－耶和华必讥笑他们， 你要嗤笑万国。
PS|59|9|我 的力量啊，我要等候你， 因为上帝是我的庇护所。
PS|59|10|我的上帝要以慈爱 迎接我， 上帝要叫我看见我的仇敌遭报。
PS|59|11|主，我们的盾牌啊， 不要杀他们，免得我的子民遗忘； 求你用你的能力使他们四散， 使他们降为卑。
PS|59|12|愿他们因口中的罪和嘴唇的言语， 被自己的骄傲抓住， 他们所说的尽是咒骂和谎话。
PS|59|13|求你发怒，使他们消灭， 求你使他们消灭，归于无有， 使他们知道上帝在 雅各 中间掌权， 直到地极。（细拉）
PS|59|14|他们晚上转回， 叫号如狗，围城绕行。
PS|59|15|他们到处走动觅食， 若不饱足就咆哮不已。
PS|59|16|但我要歌颂你的能力， 早晨要高唱你的慈爱； 因为你是我的庇护所， 在急难的日子作过我的避难所。
PS|59|17|我的力量啊，我要歌颂你； 因为上帝是我的庇护所， 是赐恩给我的上帝。
PS|60|1|上帝啊，你丢弃了我们，破坏了我们； 你曾发怒，求你使我们复兴！
PS|60|2|你使地震动，崩裂； 求你将裂口补好，因为地在摇动。
PS|60|3|你让你的子民遇见艰难， 使我们喝那令人东倒西歪的酒。
PS|60|4|你把旌旗赐给敬畏你的人， 可以躲避弓箭 。（细拉）
PS|60|5|求你应允我们 ，用右手施行拯救， 好让你所亲爱的人得救。
PS|60|6|上帝在他的圣所 说： “我要欢乐； 要划分 示剑 ， 丈量 疏割谷 。
PS|60|7|基列 是我的， 玛拿西 是我的。 以法莲 是护卫我头的， 犹大 是我的权杖。
PS|60|8|摩押 是我的沐浴盆， 我要向 以东 扔鞋。 非利士 啊，你还能因我欢呼吗？”
PS|60|9|谁能领我进坚固城？ 谁能引我到 以东 地？
PS|60|10|上帝啊，你真的丢弃了我们吗？ 上帝啊，你不和我们的军队同去吗？
PS|60|11|求你帮助我们攻击敌人， 因为人的帮助是枉然的。
PS|60|12|我们倚靠上帝才得施展大能， 因为践踏我们敌人的就是他。
PS|61|1|上帝啊，求你听我的呼求， 留心听我的祷告！
PS|61|2|我心里发昏的时候， 要从地极求告你。 求你领我到那比我更高的磐石，
PS|61|3|因为你是我的避难所， 是我的坚固台，使我脱离仇敌。
PS|61|4|我要永远住在你的帐幕里！ 我要投靠在你翅膀下的隐密处！（细拉）
PS|61|5|上帝啊，你听了我所许的愿； 你将产业赐给敬畏你名的人。
PS|61|6|求你加添王的寿数， 使他的年岁存到世世代代。
PS|61|7|愿他在上帝面前永远坐在王位上， 求你预备慈爱和信实保佑他！
PS|61|8|这样，我要歌颂你的名，直到永远， 天天还我所许的愿。
PS|62|1|我的心默默无声，专等候上帝， 我的救恩从他而来。
PS|62|2|惟独他是我的磐石，我的拯救； 他是我的庇护所，我必不大大动摇。
PS|62|3|你们大家攻击一人，使他被杀， 如歪斜的墙、将倒的壁，要到几时呢？
PS|62|4|他们彼此商议，要把他从高位上拉下来； 他们喜爱谎话，口虽祝福，心却诅咒。（细拉）
PS|62|5|我的心哪，你当默默无声，专等候上帝， 因为我的盼望是从他而来。
PS|62|6|惟独他是我的磐石，我的拯救； 他是我的庇护所，我必不动摇。
PS|62|7|我的拯救、我的荣耀都在于上帝； 我力量的磐石、我的避难所都在于上帝。
PS|62|8|百姓啊，要时时倚靠他， 在他面前倾心吐意； 上帝是我们的避难所。（细拉）
PS|62|9|人真是虚空， 人真是虚假； 放在天平里就必浮起， 他们一共比空气还轻。
PS|62|10|不要仗势欺人， 也不要因抢夺而骄傲； 若财宝加增，不要放在心上。
PS|62|11|上帝说了一次、两次，我都听见了， 就是能力属乎上帝。
PS|62|12|主啊，慈爱也是属乎你， 因为你照着各人所做的报应他。
PS|63|1|上帝啊，你是我的上帝， 我要切切寻求你； 在干旱疲乏无水之地， 我的心灵渴想你，我的肉身切慕你。
PS|63|2|我在圣所中曾如此瞻仰你， 为要见你的能力和你的荣耀。
PS|63|3|因你的慈爱比生命更好， 我的嘴唇要颂赞你。
PS|63|4|我还活着的时候要这样称颂你， 我要奉你的名举手。
PS|63|5|我在床上记念你， 在夜更的时候思念你； 我的心像吃饱了骨髓肥油， 我也要以欢乐的嘴唇赞美你。
PS|63|6|
PS|63|7|因为你曾帮助了我， 我要在你翅膀的荫下欢呼。
PS|63|8|我的心紧紧跟随你； 你的右手扶持了我。
PS|63|9|但那些寻索要灭我命的人 必往地底下去；
PS|63|10|他们必被刀剑所杀， 成为野狗的食物。
PS|63|11|但是王必因上帝欢喜， 凡指着他发誓的都要夸耀， 因为说谎之人的口必被塞住。
PS|64|1|上帝啊，我哀叹的时候，求你听我的声音！ 求你保护我的性命，不受仇敌的惊吓！
PS|64|2|求你把我隐藏， 使我脱离作恶之人的暗谋， 脱离作孽之人的扰乱。
PS|64|3|他们磨舌如刀， 发出苦毒的言语，好像瞄准了的箭，
PS|64|4|要在暗地里射完全人； 他们忽然射他，并不惧怕。
PS|64|5|他们彼此勉励，设下恶计； 他们商量，暗设圈套， 说：“谁能看见呢？”
PS|64|6|他们图谋奸恶： “我们完成了精密的策划。” 各人的意念心思是深沉的。
PS|64|7|但上帝要用箭射他们， 他们忽然受了伤。
PS|64|8|他们必然绊跌，被自己的舌头所害； 凡看见他们的都必摇头。
PS|64|9|众人都要害怕， 要传扬上帝的工作， 并且明白他的作为。
PS|64|10|义人必因耶和华欢喜，并要投靠他； 凡心里正直的人都必夸耀。
PS|65|1|上帝啊，在 锡安 ，人都等候赞美你， 也要向你还所许的愿。
PS|65|2|听祷告的主啊， 凡有血肉之躯的都要来就你。
PS|65|3|罪孽胜了我； 至于我们的过犯，你都要赦免。
PS|65|4|你所拣选、使他亲近你、住在你院中的， 这人有福了！ 我们要因你居所、你圣殿的美福知足。
PS|65|5|拯救我们的上帝啊，你必以威严秉公义应允我们； 地极和海角远方的人都倚靠你。
PS|65|6|你既以大能束腰， 就用力量安定诸山，
PS|65|7|使诸海的响声和其中波浪的响声， 并万民的喧哗，都平静了。
PS|65|8|住在地极的人因你的神迹惧怕， 你使日出日落之地都欢呼。
PS|65|9|你眷顾地， 降雨使地大大肥沃。 上帝的河满了水； 你这样浇灌了地， 好为人预备五谷。
PS|65|10|你浇透地的犁沟，润泽犁脊， 降甘霖，使地松软； 其中生长的，蒙你赐福。
PS|65|11|你以恩惠为年岁的冠冕， 你的路径都滴下油脂，
PS|65|12|滴在旷野的草场上。 小山以欢乐束腰，
PS|65|13|草场以羊群为衣， 谷中也长满了五谷； 这一切都欢呼歌唱。
PS|66|1|全地都当向上帝欢呼！
PS|66|2|当歌颂他名的荣耀， 使赞美他的话大有荣耀！
PS|66|3|当对上帝说：“你的作为何等可畏！ 因你的大能，仇敌要向你投降。
PS|66|4|全地要敬拜你，歌颂你， 要歌颂你的名。”（细拉）
PS|66|5|你们来看上帝所做的， 他向世人所做之事是可畏的。
PS|66|6|他将海变成干地，使百姓步行过河； 我们在那里要因他欢喜。
PS|66|7|他用权能治理，直到永远。 他的眼睛鉴察万民； 悖逆的人不可自高。（细拉）
PS|66|8|万民哪，你们当称颂我们的上帝， 使人得听赞美他的声音。
PS|66|9|他使我们的性命存活， 不叫我们的脚摇动。
PS|66|10|上帝啊，你曾考验我们， 你熬炼我们，如炼银子一样。
PS|66|11|你使我们进入罗网， 把重担放在我们身上。
PS|66|12|你使人坐车轧我们的头； 我们经过水火， 你却使我们到丰富之地。
PS|66|13|我要带着燔祭进你的殿， 向你还我的愿，
PS|66|14|就是在急难时我嘴唇所发的、 口中所许的。
PS|66|15|我要将肥牛的燔祭 和公羊的香祭献给你， 又要把公牛和公山羊献上。（细拉）
PS|66|16|敬畏上帝的人哪，你们都来听！ 我要述说他为我所做的事。
PS|66|17|我曾用口求告他， 我的舌头也称他为高。
PS|66|18|我若心里注重罪孽， 主必不听。
PS|66|19|但上帝实在听见了， 他留心听了我祷告的声音。
PS|66|20|上帝是应当称颂的！ 他没有推却我的祷告， 也没有使他的慈爱离开我。
PS|67|1|愿上帝怜悯我们，赐福给我们， 使他的脸向我们发光，（细拉）
PS|67|2|好让全地得知你的道路， 万国得知你的救恩。
PS|67|3|上帝啊，愿万民称谢你！ 愿万民都称谢你！
PS|67|4|愿万族都快乐欢呼； 因为你必按公正审判万民， 引导地上的万族。（细拉）
PS|67|5|上帝啊，愿万民称谢你！ 愿万民都称谢你！
PS|67|6|地已经出了土产， 上帝，我们的上帝，要赐福给我们。
PS|67|7|上帝要赐福给我们， 地的四极都要敬畏他！
PS|68|1|愿上帝兴起，使他的仇敌四散， 使那恨他的人从他面前逃跑。
PS|68|2|你驱逐他们 ，如烟被吹散； 恶人见上帝的面就消灭，如蜡被火熔化。
PS|68|3|惟有义人必然欢喜， 在上帝面前快乐， 他们要在喜乐中欢欣。
PS|68|4|你们当向上帝唱诗，歌颂他的名； 为那驾车经过旷野的修平道路 。 他的名是耶和华， 你们要在他面前欢乐！
PS|68|5|上帝在他的圣所作孤儿的父， 作寡妇的伸冤者。
PS|68|6|上帝使孤独的有家， 使被囚的出来享福； 惟有悖逆的要住在干旱之地。
PS|68|7|上帝啊，当你走在百姓前头， 在旷野行进，（细拉）
PS|68|8|地见上帝的面就震动，天也降雨； 西奈山 见 以色列 上帝的面也震动。
PS|68|9|上帝啊，你降下大雨； 你的产业 以色列 疲乏的时候，你使他坚固。
PS|68|10|你的会众住在境内； 上帝啊，你在恩惠中为困苦人预备所需的。
PS|68|11|主发命令， 传好信息的妇女成了大群：
PS|68|12|“统领大军的君王逃跑了，逃跑了！” 在家等候的妇女也分得了掠物。
PS|68|13|你们躺卧在羊圈， 好像鸽子的翅膀镀银，翎毛镀金一般。
PS|68|14|全能者在境内赶散列王的时候， 势如飘雪在 撒们 。
PS|68|15|巴珊山 是极其宏伟 的山， 巴珊山 是多峰多岭的山。
PS|68|16|你们多峰多岭的山哪， 为何以妒忌的眼光看上帝所愿居住的山？ 耶和华必住这山，直到永远！
PS|68|17|上帝的车辇累万盈千； 主在其中，好像在 西奈 圣山一样。
PS|68|18|你已经升上高天，掳掠了俘虏； 你在人间，就是在悖逆的人中，受了供献， 使耶和华上帝可以与他们同住。
PS|68|19|天天背负我们重担的主， 就是拯救我们的上帝， 是应当称颂的！（细拉）
PS|68|20|上帝是为我们施行拯救的上帝； 人能脱离死亡是在乎主─耶和华。
PS|68|21|但上帝要打破他仇敌的头， 就是那常犯罪之人的头颅。
PS|68|22|主说：“我要使百姓从 巴珊 归来， 使他们从深海转回，
PS|68|23|好叫你打碎仇敌，使你的脚踹在血中， 使你狗的舌头也有份。”
PS|68|24|上帝啊，你是我的上帝，我的王； 人已经看见你行走，进入圣所。
PS|68|25|歌唱的行在前，作乐的随在后， 都在击鼓的童女中间：
PS|68|26|“从 以色列 源头而来的啊， 你们当在各会中称颂上帝─耶和华！”
PS|68|27|在那里，有统管他们的小 便雅悯 ， 有 犹大 的领袖和他们的一群人， 有 西布伦 的领袖， 有 拿弗他利 的领袖。
PS|68|28|你的上帝已赐给你力量 ； 上帝啊，求你坚固你为我们所成全的事！
PS|68|29|因你 耶路撒冷 的殿， 列王必带贡物献给你。
PS|68|30|求你斥责芦苇中的野兽和公牛群， 并万民中的牛犊。 直到他们带着银块来朝贡 ； 上帝已经赶散好战的万民 。
PS|68|31|埃及 的使臣要出来， 古实 人要急忙向上帝伸出手来。
PS|68|32|地上的国度啊， 你们要向上帝歌唱， 要歌颂主，（细拉）
PS|68|33|就是那驾行在亘古的诸天之上的主！ 听啊，他发出声音，是极大的声音。
PS|68|34|你们要将能力归给上帝； 他的威荣在 以色列 之上， 他的能力显在天上。
PS|68|35|上帝啊，你从圣所显为可畏， 以色列 的上帝是那将力量权能赐给他百姓的。 上帝是应当称颂的！
PS|69|1|上帝啊，求你救我！ 因为众水就要淹没我。
PS|69|2|我深陷在淤泥中，没有立脚之地； 我到了深水之中，波涛漫过我身。
PS|69|3|我因呼求困乏，喉咙发干； 我因等候上帝，眼睛失明。
PS|69|4|无故恨我的，比我的头发还多； 无理与我为仇、要把我剪除的，甚为强盛。 我没有抢夺，他们竟然要我偿还！
PS|69|5|上帝啊，我的愚昧，你原知道， 我的罪愆不能向你隐瞒。
PS|69|6|万军之主耶和华啊， 求你不要让那等候你的因我蒙羞！ 以色列 的上帝啊， 求你不要让那寻求你的因我受辱！
PS|69|7|因我为你的缘故受了辱骂， 满面羞愧。
PS|69|8|我的兄弟把我当陌生人， 我母亲的儿子把我当外邦人。
PS|69|9|因我为你的殿心里焦急，如同火烧， 并且辱骂你的人的辱骂都落在我身上。
PS|69|10|我哭泣，以禁食刻苦我心； 这倒成了我的羞辱。
PS|69|11|我拿麻布当衣裳， 却成了他们的笑柄。
PS|69|12|坐在城门口的谈论我， 酒徒也以我为歌曲。
PS|69|13|至于我，耶和华啊，在悦纳的时候我向你祈祷。 上帝啊，求你按你丰盛的慈爱， 凭你拯救的信实应允我！
PS|69|14|求你搭救我脱离淤泥， 不叫我陷在其中； 求你使我脱离那些恨我的人， 使我脱离深水。
PS|69|15|求你不容波涛漫过我， 不容深渊吞灭我， 不容深坑在我以上合口。
PS|69|16|耶和华啊，求你应允我！ 因为你的慈爱本为美好； 求你按你丰盛的怜悯转回眷顾我！
PS|69|17|不要转脸不顾你的仆人； 我在急难之中，求你速速应允我！
PS|69|18|求你亲近我，救赎我！ 求你因我仇敌的缘故将我赎回！
PS|69|19|你知道我所受的辱骂、欺凌、羞辱； 我的敌人都在你面前。
PS|69|20|辱骂刺伤我的心， 使我忧愁。 我指望有人体恤，却没有一个； 指望有人安慰，却找不着一个。
PS|69|21|他们拿苦胆给我当食物； 我渴了，他们拿醋给我喝。
PS|69|22|愿他们的筵席在他们面前变为罗网， 在他们平安的时候 变为圈套。
PS|69|23|愿他们的眼睛昏花，看不见； 求你使他们的腰常常战抖。
PS|69|24|求你将你的恼恨倒在他们身上， 使你的烈怒追上他们。
PS|69|25|愿他们的住处变为废墟， 他们的帐棚无人居住。
PS|69|26|因为你所击打的，他们就迫害； 你所击伤的，他们述说 他的愁苦。
PS|69|27|求你使他们罪上加罪， 不容他们在你面前称义。
PS|69|28|愿他们从生命册上被涂去， 不得名列在义人之中。
PS|69|29|但我困苦忧伤； 上帝啊，愿你的救恩将我安置在高处。
PS|69|30|我要以诗歌赞美上帝的名， 以感谢尊他为大！
PS|69|31|这就让耶和华喜悦，胜似献牛， 献有角有蹄的公牛。
PS|69|32|谦卑的人看见了就喜乐； 寻求上帝的人，愿你们的心苏醒。
PS|69|33|因为耶和华听了穷乏的人， 不藐视被囚的人。
PS|69|34|愿天和地、 海洋和其中一切的动物都赞美他！
PS|69|35|因为上帝要拯救 锡安 ，建造 犹大 的城镇； 他的子民要在那里居住，得地为业。
PS|69|36|他仆人的后裔要承受这地， 爱他名的人要住在其中。
PS|70|1|上帝啊，求你快快搭救我！ 耶和华啊，求你速速帮助我！
PS|70|2|愿那些寻索我命的，抱愧蒙羞； 愿那些喜悦我遭害的，退后受辱。
PS|70|3|愿那些对我说“啊哈、啊哈”的， 因羞愧退后。
PS|70|4|愿所有寻求你的，因你欢喜快乐； 愿那些喜爱你救恩的，常说：“当尊上帝为大！”
PS|70|5|但我是困苦贫穷的； 上帝啊，求你速速到我这里来！ 你是帮助我的，搭救我的； 耶和华啊，求你不要耽延！
PS|71|1|耶和华啊，我投靠你， 求你叫我永不羞愧！
PS|71|2|求你凭你的公义搭救我，救拔我； 侧耳听我，拯救我！
PS|71|3|求你作我常来栖身 的磐石， 你已经吩咐要救我， 因为你是我的岩石、我的山寨。
PS|71|4|我的上帝啊，求你救我脱离恶人的手， 脱离不义和残暴之人的手。
PS|71|5|主耶和华啊，你是我所盼望的； 自我年幼，你是我所倚靠的。
PS|71|6|我自出母胎被你扶持， 使我出母腹的是你。 我要常常赞美你！
PS|71|7|许多人看我为异类， 但你是我坚固的避难所。
PS|71|8|我要满口述说赞美你的话 终日荣耀你。
PS|71|9|我年老的时候，求你不要丢弃我！ 我体力衰弱时，求你不要离弃我！
PS|71|10|我的仇敌议论我， 那些窥探要害我命的一同商议，
PS|71|11|说：“上帝已经离弃他； 你们去追赶他，捉拿他吧！ 因为没有人搭救。”
PS|71|12|上帝啊，求你不要远离我！ 我的上帝啊，求你速速帮助我！
PS|71|13|愿那与我为敌的，羞愧灭亡； 愿那谋害我的，受辱蒙羞。
PS|71|14|我却要常常仰望， 并要越发赞美你。
PS|71|15|我的口要终日述说你的公义和你的救恩， 因我无从计算其数。
PS|71|16|我要述说主耶和华的大能， 我单要提说你的公义。
PS|71|17|上帝啊，自我年幼，你就教导我； 直到如今，我传扬你奇妙的作为。
PS|71|18|上帝啊，我年老发白的时候， 求你不要离弃我！ 等我宣扬你的能力给下一代， 宣扬你的大能给后世的人。
PS|71|19|上帝啊，你的公义极高； 行过大事的上帝啊，谁能像你？
PS|71|20|你是叫我多经历重大急难的， 必使我再活过来， 从地的深处救我上来。
PS|71|21|你必使我越发昌大， 又转来安慰我。
PS|71|22|我的上帝啊，我要鼓瑟称谢你， 称谢你的信实！ 以色列 的圣者啊，我要弹琴歌颂你！
PS|71|23|我歌颂你的时候，我的嘴唇要欢呼； 我的性命，就是你所救赎的，也要欢呼。
PS|71|24|我的舌头也必终日讲论你的公义， 因为那些谋害我的人已经蒙羞受辱了。
PS|72|1|上帝啊，求你将你的公平赐给王， 将你的公义赐给王的儿子。
PS|72|2|使他按公义审判你的子民， 按公平审判你的困苦人。
PS|72|3|大山小山都要因公义 使百姓得享平安。
PS|72|4|他必为百姓中困苦的人伸冤， 拯救贫穷之辈， 压碎那欺压人的人。
PS|72|5|太阳还存，月亮犹在， 人要敬畏你 ，直到万代！
PS|72|6|他必降临，像雨降在已割的草地上， 如甘霖滋润田地。
PS|72|7|在他的日子，公义 要兴旺， 大有平安，除非月亮不在。
PS|72|8|他要执掌权柄，从这海直到那海， 从 大河 直到地极。
PS|72|9|住在旷野的必在他面前下拜， 他的仇敌必要舔土。
PS|72|10|他施 和海岛的王要进贡， 示巴 和 西巴 的王要献礼物。
PS|72|11|众王都要叩拜他， 万国都要事奉他。
PS|72|12|贫穷人呼求，他要搭救， 无人帮助的困苦人，他也搭救。
PS|72|13|他要怜悯贫寒和贫穷的人， 拯救贫穷人的性命。
PS|72|14|他要救赎他们脱离欺压和残暴， 他们的血在他眼中看为宝贵。
PS|72|15|愿他永远活着， 示巴 的金子要献给他； 愿人常常为他祷告，终日祝福他。
PS|72|16|在地的山顶上，愿五谷茂盛， 所结的谷实响动，如 黎巴嫩 的树林； 愿城里的人兴旺，如地上的草。
PS|72|17|愿他的名存到永远， 他的名如太阳之长久 ； 愿人因他蒙福， 万国称他为有福。
PS|72|18|惟独耶和华－ 以色列 的上帝能行奇事， 他是应当称颂的！
PS|72|19|他荣耀的名也当称颂，直到永远。 愿他的荣耀充满全地！ 阿们！阿们！
PS|72|20|耶西 的儿子－ 大卫 的祈祷完毕。 亚萨的诗。
PS|73|1|上帝实在恩待 以色列 那些清心的人！
PS|73|2|至于我，我的脚几乎失闪， 我的步伐险些走偏；
PS|73|3|因为我嫉妒狂傲的人， 我看见恶人享平安。
PS|73|4|他们的力气强壮， 他们死的时候也没有疼痛。
PS|73|5|他们不像别人受苦， 也不像别人遭灾。
PS|73|6|所以，骄傲如链子戴在他们项上， 残暴像衣裳覆盖在他们身上。
PS|73|7|他们的眼睛 因体胖而凸出， 他们的内心放任不羁 。
PS|73|8|他们讥笑人，凭恶意说欺压人的话。 他们说话自高；
PS|73|9|他们的口亵渎上天， 他们的舌毁谤全地。
PS|73|10|所以他的百姓归到这里， 享受满杯的水 。
PS|73|11|他们说：“上帝怎能晓得？ 至高者哪会知道呢？”
PS|73|12|看哪，这就是恶人， 他们常享安逸，财宝增多。
PS|73|13|我实在徒然洁净了我的心， 徒然洗手表明我的无辜，
PS|73|14|因为我终日遭灾难， 每日早晨受惩治。
PS|73|15|我若说“我要这样讲”， 就是愧对这世代的众儿女了。
PS|73|16|我思索要明白这事， 眼看实系为难，
PS|73|17|直到我进了上帝的圣所， 思想他们的结局。
PS|73|18|你实在把他们安放在滑地， 使他们跌倒灭亡；
PS|73|19|他们转眼之间成了何等荒凉！ 他们被惊恐灭尽了。
PS|73|20|人睡醒了，怎样看梦， 主啊，你醒了也必照样轻看他们的影像。
PS|73|21|因此，我心里苦恼， 肺腑被刺。
PS|73|22|我这样愚昧无知， 在你面前如同畜牲。
PS|73|23|然而，我常与你同在； 你搀扶我的右手。
PS|73|24|你要以你的训言引导我， 以后你必接我到荣耀里。
PS|73|25|除你以外，在天上我有谁呢？ 除你以外，在地上我也没有所爱慕的。
PS|73|26|我的肉体和我的心肠衰残； 但上帝是我心里的力量， 又是我的福分，直到永远。
PS|73|27|看哪，远离你的，必要死亡； 凡离弃你行淫的，你都灭绝了。
PS|73|28|但我亲近上帝是于我有益； 我以主耶和华为我的避难所， 好叫我述说你一切的作为。
PS|74|1|上帝啊，你为何永远丢弃我们呢？ 为何向你草场的羊发怒，如烟冒出呢？
PS|74|2|求你记念你古时得来的会众， 就是你所赎、作你产业支派的， 并记念你向来居住的 锡安山 。
PS|74|3|求你举步去看那日久荒凉之地， 看仇敌在圣所中所做的一切恶事。
PS|74|4|你的敌人在你会中吼叫， 他们竖起自己的标帜为记号，
PS|74|5|好像人扬起斧子 对着林中的树，
PS|74|6|现在将圣所中的雕刻 ， 全都用斧子锤子打坏。
PS|74|7|他们用火焚烧你的圣所， 亵渎你名的居所于地。
PS|74|8|他们心里说“我们要尽行毁灭”； 就在遍地烧毁敬拜上帝聚会的所在。
PS|74|9|我们看不见自己的标帜，不再有先知， 我们当中也无人知道这灾祸要到几时。
PS|74|10|上帝啊，敌人辱骂要到几时呢？ 仇敌藐视你的名要到永远吗？
PS|74|11|你为什么缩回你的右手？ 求你从怀中伸出手来，毁灭他们。
PS|74|12|上帝自古以来是我的王， 在这地上施行拯救。
PS|74|13|你曾用能力将海分开， 你打破水里大鱼的头。
PS|74|14|你曾压碎 力威亚探 的头， 把它给旷野的禽兽作食物。
PS|74|15|你曾分裂泉源和溪流； 使长流的江河枯干。
PS|74|16|白昼属你，黑夜也属你； 亮光和太阳是你预备的。
PS|74|17|地的一切疆界是你立的， 夏天和冬天是你定的。
PS|74|18|耶和华啊，仇敌辱骂，愚顽之辈藐视你的名； 求你记念这事。
PS|74|19|不要将属你的斑鸠 交给野兽， 不要永远忘记你困苦人的性命。
PS|74|20|求你顾念所立的约， 因为地上黑暗之处遍满了凶暴。
PS|74|21|不要让受欺压的人蒙羞回去； 要使困苦贫穷的人赞美你的名。
PS|74|22|上帝啊，求你起来为自己辩护！ 求你记念愚顽人怎样终日辱骂你。
PS|74|23|不要忘记你敌人的喧闹， 就是那时常上升、起来对抗你之人的喧哗。
PS|75|1|上帝啊，我们称谢你，我们称谢你！ 你的名临近，人 都述说你奇妙的作为。
PS|75|2|我选定了日期， 必按正直施行审判。
PS|75|3|地和其上的居民都熔化了； 我亲自坚立地的柱子。（细拉）
PS|75|4|我对狂傲的人说：“不要狂傲！” 对凶恶的人说：“不要举角！”
PS|75|5|不要把你们的角高举， 不要挺着颈项 说话。
PS|75|6|因为高举非从东，非从西， 也非从南而来。
PS|75|7|惟有上帝断定， 他使这人降卑，使那人升高。
PS|75|8|耶和华的手里有杯， 杯内满了调和起沫的酒； 他倒出来， 地上的恶人都必喝，直到喝尽它的渣滓。
PS|75|9|但我要宣扬，直到永远！ 我要歌颂 雅各 的上帝！
PS|75|10|恶人一切的角，我要砍断； 惟有义人的角必被高举。
PS|76|1|在 犹大 ，上帝为人所认识； 在 以色列 ，他的名为大。
PS|76|2|在 撒冷 有他的住处， 在 锡安 有他的居所。
PS|76|3|他在那里折断弓上的火箭、 盾牌、刀剑和战争的兵器。（细拉）
PS|76|4|你是光荣的， 比猎物 之山更威严。
PS|76|5|心中勇敢的人都被掠夺； 他们睡了长觉，没有一个英雄能措手。
PS|76|6|雅各 的上帝啊，你的斥责一发， 战车和战马都沉睡了。
PS|76|7|你，惟独你是可畏的！ 你的怒气一发，谁能在你面前站得住呢？
PS|76|8|你从天上使人听判断。 上帝起来施行审判， 要救地上所有困苦的人； 那时地就惧怕而静默。（细拉）
PS|76|9|
PS|76|10|人的愤怒终必称谢你， 你要以人的余怒束腰。
PS|76|11|你们当向耶和华－你们的上帝许愿，还愿； 在他四围的人都当拿贡物献给那可畏的主。
PS|76|12|他要挫折王子的骄气， 向地上的君王显为可畏。
PS|77|1|我要向上帝发声呼求； 我向上帝发声，他必侧耳听我。
PS|77|2|我在患难之日寻求主， 在夜间不住地举手祷告 ， 我的心不肯受安慰。
PS|77|3|我想念上帝，就烦躁不安； 我沉思默想，心灵发昏。（细拉）
PS|77|4|你使我不能闭眼； 我心烦乱，甚至不能说话。
PS|77|5|我追想古时之日， 上古之年。
PS|77|6|夜间我想起我的歌曲 ， 我的心默想，我的灵仔细省察：
PS|77|7|“难道主要永远丢弃我， 不再施恩吗？
PS|77|8|难道他的慈爱永远穷尽， 他的应许世世废弃吗？
PS|77|9|难道上帝忘记施恩， 因发怒就止住他的怜悯吗？”（细拉）
PS|77|10|我说，至高者右手的能力已改变， 这是我的悲哀。
PS|77|11|我要记念耶和华所做的， 要记念你古时的奇事；
PS|77|12|我要思想你所做的， 默念你的作为。
PS|77|13|上帝啊，你的道是神圣的； 有何神明大如上帝呢？
PS|77|14|你是行奇事的上帝， 你曾在万民中彰显能力。
PS|77|15|你曾用膀臂赎了你的子民， 就是 雅各 和 约瑟 的子孙。（细拉）
PS|77|16|上帝啊，众水见你， 众水一见你就都惊惶， 深渊也都战抖。
PS|77|17|密云倒出水来， 天空发出响声， 你的箭也飞行四方。
PS|77|18|你的雷声在旋风之中， 闪电照亮世界， 大地战抖震动。
PS|77|19|你的道在海中， 你的路在大水之中， 你的脚踪无人知道。
PS|77|20|你曾藉 摩西 和 亚伦 的手引导你的百姓， 好像领羊群一般。
PS|78|1|我的子民哪，要侧耳听我的训诲， 竖起耳朵听我口中的言语。
PS|78|2|我要开口说比喻， 我要解开古时的谜语，
PS|78|3|是我们所听见、所知道， 我们的祖宗告诉我们的。
PS|78|4|我们不要向子孙隐瞒这些事， 而要将耶和华的美德和他的能力， 并他所行的奇事，述说给后代听。
PS|78|5|他在 雅各 中立法度， 在 以色列 中设律法； 他吩咐我们的祖宗要传给子孙，
PS|78|6|使将要生的后代子孙可以晓得。 他们也要起来告诉他们的子孙，
PS|78|7|好让他们仰望上帝， 不忘记上帝的作为， 惟遵守他的命令；
PS|78|8|不要像他们的祖宗， 是顽梗悖逆、心不坚定， 向上帝心不忠实之辈。
PS|78|9|以法莲 人带着兵器，拿着弓， 临阵之日转身退后。
PS|78|10|他们不遵守上帝的约， 不肯照他的律法行；
PS|78|11|又忘记他的作为 和他所彰显的奇事。
PS|78|12|他在 埃及 地，在 琐安 田， 在他们祖宗眼前施行奇事。
PS|78|13|他把海分开，使他们过去， 又叫水立起如垒。
PS|78|14|他白日用云彩， 终夜用火光引导他们。
PS|78|15|他在旷野使磐石裂开， 多多地给他们水喝，如从深渊而出。
PS|78|16|他使水从磐石涌出， 叫水如江河下流。
PS|78|17|他们却仍旧得罪他， 在干旱之地悖逆至高者。
PS|78|18|他们心中试探上帝， 随自己所欲的求食物，
PS|78|19|并且妄论上帝说： “上帝岂能在旷野摆设筵席吗？
PS|78|20|他虽曾击打磐石，使水涌出，如江河泛滥； 他还能赐粮食吗？ 还能为他的百姓预备吃的肉吗？”
PS|78|21|所以，耶和华听见就发怒， 有烈火向 雅各 点燃， 有怒气向 以色列 上腾；
PS|78|22|因为他们不信服上帝， 不倚赖他的拯救。
PS|78|23|然而他却吩咐天空， 又敞开天上的门，
PS|78|24|降吗哪像雨，给他们吃， 将天上的粮食赐给他们。
PS|78|25|各人就吃大能者的食物； 他赐下粮食，使他们饱足。
PS|78|26|他令东风吹在天空， 用能力引来南风。
PS|78|27|他降肉像雨，多如尘土， 降飞鸟，多如海沙，
PS|78|28|落在他自己的营中， 在他帐幕的四周围。
PS|78|29|他们吃了，而且饱足； 这样就随了他们所欲的。
PS|78|30|但在他们满足食欲以前， 食物还在他们口中的时候，
PS|78|31|上帝的怒气就向他们上腾， 杀了他们当中肥壮的人， 打倒 以色列 的青年。
PS|78|32|虽是这样，他们仍旧犯罪， 不信他奇妙的作为。
PS|78|33|因此，他使他们的日子全归虚空， 叫他们的年岁尽属惊恐。
PS|78|34|他杀他们的时候，他们才求问他， 回心转意，切切寻求上帝。
PS|78|35|他们追念上帝是他们的磐石， 至高的上帝是他们的救赎主。
PS|78|36|他们却用口谄媚他， 用舌向他说谎。
PS|78|37|他们的心向他不坚定， 不忠于他的约。
PS|78|38|但他有怜悯， 赦免他们的罪孽， 没有灭绝他们， 而且屡次撤销他的怒气， 不发尽他的愤怒。
PS|78|39|他想念他们不过是血肉之躯， 是一阵去而不返的风。
PS|78|40|他们在旷野悖逆他， 在荒地令他担忧，何其多呢！
PS|78|41|他们再三试探上帝， 惹动 以色列 的圣者。
PS|78|42|他们不追念他手的能力， 和他救赎他们脱离敌人的日子；
PS|78|43|他怎样在 埃及 显神迹， 在 琐安 田显奇事，
PS|78|44|把江河并河汊的水都变为血， 使他们不能喝。
PS|78|45|他使苍蝇成群落在他们当中，吃尽他们， 又叫青蛙灭了他们，
PS|78|46|将他们的果实交给蚂蚱， 把他们劳碌得来的交给蝗虫。
PS|78|47|他降冰雹打坏他们的葡萄树， 下寒霜打坏他们的桑树，
PS|78|48|将他们的牲畜交给冰雹， 把他们的群畜交给闪电。
PS|78|49|他使猛烈的怒气和愤怒、恼恨、苦难， 成了一群降灾的使者，临到他们。
PS|78|50|他为自己的怒气修平了路， 将他们的性命交给瘟疫， 使他们死亡，
PS|78|51|在 埃及 击杀所有的长子， 在 含 的帐棚中击杀他们壮年时头生的。
PS|78|52|他却领出自己的子民如羊， 在旷野引导他们如羊群。
PS|78|53|他领他们稳稳妥妥地，使他们不致害怕； 海却淹没他们的仇敌。
PS|78|54|他带他们到自己圣地的边界， 到他右手所得的这山地。
PS|78|55|他在他们面前赶出外邦人， 用绳子抽签量地给他们为业， 让 以色列 支派的人住在自己的帐棚里。
PS|78|56|他们仍旧试探，悖逆至高的上帝， 不遵守他的法度，
PS|78|57|反倒退后，行诡诈，像他们的祖宗一样， 他们翻转，如同松弛的弓，
PS|78|58|以丘坛惹他发怒， 以雕刻的偶像使他忌恨。
PS|78|59|上帝听见就发怒， 全然弃绝了 以色列 ，
PS|78|60|甚至离弃 示罗 的帐幕， 就是他在人间所搭的帐棚；
PS|78|61|又将他有能力的约柜 交给人掳去， 将他的荣耀交在敌人手中；
PS|78|62|并将他的百姓交给刀剑， 向他的产业发怒。
PS|78|63|壮丁被火烧灭， 童女也无婚礼颂歌。
PS|78|64|祭司倒在刀下， 寡妇却不哀哭。
PS|78|65|那时，主像睡觉的人醒来， 如勇士饮酒呼喊。
PS|78|66|他击退敌人， 叫他们永蒙羞辱。
PS|78|67|他撇弃 约瑟 的帐棚， 不拣选 以法莲 支派，
PS|78|68|却拣选 犹大 支派， 拣选他所喜爱的 锡安山 ；
PS|78|69|建造他的圣所如同高峰， 又像他所建立的永存之地。
PS|78|70|他拣选他的仆人 大卫 ， 从羊圈中将他召来，
PS|78|71|叫他不再牧放那些母羊， 为要牧养自己的百姓 雅各 和自己的产业 以色列 。
PS|78|72|于是，他以纯正的心牧养他们， 用巧妙的手引导他们。
PS|79|1|上帝啊，外邦人侵犯你的产业， 玷污你的圣殿，使 耶路撒冷 变成废墟，
PS|79|2|将你仆人的尸首交给天空的飞鸟为食， 把你圣民的肉交给地上的走兽，
PS|79|3|耶路撒冷 的周围流出他们的血如水， 无人埋葬。
PS|79|4|我们成为邻国羞辱的对象， 被四围的人嗤笑讥刺。
PS|79|5|耶和华啊，你发怒要到几时呢？ 要到永远吗？ 你的忌恨要如火焚烧吗？
PS|79|6|求你将你的愤怒倾倒在那不认识你的万邦 和那不求告你名的国度。
PS|79|7|因为他们吞了 雅各 ， 将他的住处变为废墟。
PS|79|8|求你不要记得我们先前世代的罪孽； 愿你的怜悯速速临到我们， 因为我们落到极卑微的地步。
PS|79|9|拯救我们的上帝啊，求你因你名的荣耀帮助我们！ 为你名的缘故搭救我们，赦免我们的罪。
PS|79|10|为何让列国说“他们的上帝在哪里”呢？ 求你让列国知道， 你在我们眼前伸你仆人流血的冤。
PS|79|11|愿被囚之人的叹息达到你面前， 求你以强大的膀臂存留那些将死的人。
PS|79|12|主啊，求你将我们邻邦所加给你的羞辱 七倍归到他们身上。
PS|79|13|这样，你的子民，你草场的羊， 要称谢你，直到永远； 要述说赞美你的话，直到万代。
PS|80|1|领 约瑟 如领羊群的 以色列 牧者啊，求你侧耳而听！ 在基路伯之上坐宝座的啊，求你发出光来！
PS|80|2|在 以法莲 、 便雅悯 、 玛拿西 面前 求你施展你的大能，拯救我们。
PS|80|3|上帝啊，求你使我们回转 ， 使你的脸发光，我们就会得救！
PS|80|4|耶和华─万军之上帝啊， 你因你百姓的祷告发怒，要到几时呢？
PS|80|5|你以眼泪当食物给他们吃， 量出满碗的眼泪给他们喝。
PS|80|6|你使邻邦因我们纷争， 我们的仇敌彼此戏笑。
PS|80|7|万军之上帝啊，求你使我们回转， 使你的脸发光，我们就会得救！
PS|80|8|你从 埃及 拔出一棵葡萄树， 赶出外邦人，把这树栽上。
PS|80|9|你在它面前清除杂物， 它就深深扎根，蔓延满地。
PS|80|10|它的影子遮蔽群山， 枝子好像高大的香柏树。
PS|80|11|它长出枝子，直到大海， 伸展嫩枝，延到 大河 。
PS|80|12|你为何拆毁这树的篱笆， 任凭路人摘取？
PS|80|13|林中的野猪践踏它， 田里的走兽吞吃它。
PS|80|14|万军之上帝啊，求你转回， 从天上垂看观察，眷顾这葡萄树；
PS|80|15|保护你右手所栽的根， 你为自己所坚固的幼苗。
PS|80|16|这树已经被火焚烧，被刀砍伐， 因你脸上的怒容就灭亡了。
PS|80|17|愿你的手扶持你右边的人， 你为自己所坚固的人子。
PS|80|18|这样，我们就不背离你； 求你救活我们，让我们得以求告你的名。
PS|80|19|耶和华─万军之上帝啊，求你使我们回转， 使你的脸发光，我们就会得救！
PS|81|1|你们当向上帝－我们的力量大声歌唱， 向 雅各 的上帝欢呼！
PS|81|2|高唱诗歌，击打手鼓， 弹奏悦耳的琴瑟。
PS|81|3|当在新月和满月－ 我们过节的日期吹角，
PS|81|4|因这是为 以色列 所定的律例， 是 雅各 上帝的典章。
PS|81|5|他攻击 埃及 地的时候， 曾立此为 约瑟 的法度。 我听见我所不明白的语言：
PS|81|6|“我使你 的肩头得脱重担， 使你的手放下筐子。
PS|81|7|你在急难中呼求，我就搭救你， 在雷的隐密处应允你， 在 米利巴 水那里考验你。（细拉）
PS|81|8|听啊，我的子民，我要劝戒你； 以色列 啊，我真愿你肯听从我。
PS|81|9|在你当中，不可有外族的神明； 外邦的神明，你也不可下拜。
PS|81|10|我是耶和华－你的上帝， 曾将你从 埃及 地领上来； 你要大大张口，我就使你满足。
PS|81|11|“无奈，我的子民不听我的声音， 以色列 不肯听从我。
PS|81|12|我就任凭他们心里顽梗， 随自己的计谋而行。
PS|81|13|我的子民若肯听从我， 以色列 肯行我的道，
PS|81|14|我就速速制伏他们的仇敌， 反手攻击他们的敌人。
PS|81|15|恨耶和华的人必来投降， 愿他们的厄运直到永远。
PS|81|16|他必拿上好的麦子给 以色列 吃， 又拿磐石出的蜂蜜使你饱足。 ”
PS|82|1|上帝站立在神圣的会中， 在诸神中施行审判。
PS|82|2|你们审判不秉公义， 抬举恶人的脸面，要到几时呢？（细拉）
PS|82|3|当为贫寒的人和孤儿伸冤， 为困苦和穷乏的人施行公义。
PS|82|4|当保护贫寒和贫穷的人， 救他们脱离恶人的手。
PS|82|5|他们愚昧，他们无知， 在黑暗中走来走去； 地的根基都摇动了。
PS|82|6|我曾说：“你们是诸神， 都是至高者的儿子。
PS|82|7|然而，你们要死去，与世人一样， 要仆倒，像任何一位王子一般。”
PS|82|8|上帝啊，求你起来审判全地， 因为你必得万国为业。
PS|83|1|上帝啊，求你不要静默！ 上帝啊，求你不要闭口，不要不作声！
PS|83|2|因为你的仇敌喧嚷， 恨你的抬起头来。
PS|83|3|他们同谋奸诈要害你的百姓， 彼此商议要害你所保护的人。
PS|83|4|他们说：“来吧，我们将他们除灭， 使他们不再成国！ 使 以色列 的名不再被人记念！”
PS|83|5|他们同心商议， 彼此结盟，要抵挡你；
PS|83|6|他们就是住帐棚的 以东 和 以实玛利 人， 摩押 和 夏甲 人，
PS|83|7|迦巴勒 、 亚扪 、 亚玛力 、 非利士 和 推罗 的居民。
PS|83|8|亚述 也与他们联合， 作 罗得 子孙的帮手。（细拉）
PS|83|9|求你待他们，如待 米甸 ， 如在 基顺河 待 西西拉 和 耶宾 一样。
PS|83|10|他们在 隐．多珥 灭亡， 成了地上的粪土。
PS|83|11|求你使他们的贵族像 俄立 和 西伊伯 ， 使他们的王子都像 西巴 和 撒慕拿 。
PS|83|12|因为他们说：“我们要得上帝的住处， 作自己的产业。”
PS|83|13|我的上帝啊，求你使他们像旋风中的尘土， 如风前的碎秸。
PS|83|14|火怎样焚烧树林， 火焰怎样烧着山岭，
PS|83|15|求你也照样用狂风追赶他们， 用暴雨恐吓他们。
PS|83|16|耶和华啊，求你使他们满面羞耻， 好叫他们寻求你的名！
PS|83|17|愿他们永远羞愧惊惶！ 愿他们惭愧灭亡！
PS|83|18|愿他们认识你的名是耶和华， 惟独你是掌管全地的至高者！
PS|84|1|万军之耶和华啊， 你的居所何等可爱！
PS|84|2|我羡慕渴想耶和华的院宇， 我的内心，我的肉体向永生上帝欢呼。
PS|84|3|万军之耶和华－我的王，我的上帝啊， 在你祭坛那里，麻雀为自己找到了家， 燕子为自己找着菢雏之窝。
PS|84|4|如此住在你殿中的有福了！ 他们不断地赞美你。（细拉）
PS|84|5|靠你有力量、心中向往 锡安 大道的， 这人有福了！
PS|84|6|他们经过“流泪谷” ，叫这谷变为泉源之地； 且有秋雨之福盖满了全谷。
PS|84|7|他们行走，力上加力， 各人到 锡安 朝见上帝。
PS|84|8|万军之耶和华上帝啊，求你听我的祷告！ 雅各 的上帝啊，求你侧耳而听！（细拉）
PS|84|9|上帝啊，我们的盾牌，求你观看， 求你垂顾你受膏者的面！
PS|84|10|在你的院宇一日， 胜似千日； 宁可在我上帝的殿中看门， 不愿住在恶人的帐棚里。
PS|84|11|因为耶和华上帝是太阳，是盾牌， 耶和华要赐下恩惠和荣耀。 他未尝留下福气不给那些行动正直的人。
PS|84|12|万军之耶和华啊， 倚靠你的人有福了！
PS|85|1|耶和华啊，你已经向你的地施恩， 救回被掳的 雅各 。
PS|85|2|你赦免了你百姓的罪孽， 遮盖了他们一切的过犯。（细拉）
PS|85|3|你收回所发的愤怒， 撤销你猛烈的怒气。
PS|85|4|拯救我们的上帝啊，求你使我们回转， 使你向我们所发的愤怒止息。
PS|85|5|你要向我们发怒到永远吗？ 要将你的怒气延留到万代吗？
PS|85|6|你不再将我们救活， 使你的百姓因你欢喜吗？
PS|85|7|耶和华啊，求你使我们得见你的慈爱， 又将你的救恩赐给我们。
PS|85|8|我要听上帝－耶和华所说的话， 因为他必应许赐平安给他的百姓，就是他的圣民； 他们却不可再转向愚昧 。
PS|85|9|他的救恩诚然与敬畏他的人相近， 使荣耀住在我们的地上。
PS|85|10|慈爱和诚实彼此相遇， 公义与和平彼此相亲。
PS|85|11|诚实从地而生， 公义从天而现。
PS|85|12|耶和华必赐福气给我们； 我们的地也要出土产。
PS|85|13|公义要行在他面前， 使他的脚踪有可走之路。
PS|86|1|耶和华啊，求你侧耳应允我， 因我是困苦贫穷的。
PS|86|2|求你保住我的性命，因我是虔诚的人。 我的上帝啊，求你拯救我这倚靠你的仆人！
PS|86|3|主啊，求你怜悯我， 因我终日求告你。
PS|86|4|主啊，求你使你的仆人心里欢喜， 因为我的心仰望你。
PS|86|5|主啊，你本为良善，乐于饶恕人， 以丰盛的慈爱对待凡求告你的人。
PS|86|6|耶和华啊，求你侧耳听我的祷告， 留心听我恳求的声音。
PS|86|7|我在患难之日要求告你， 因为你必应允我。
PS|86|8|主啊，诸神之中没有可与你相比的， 你的作为也无以为比。
PS|86|9|主啊，你所造的万民都要来敬拜你， 他们要荣耀你的名。
PS|86|10|因你本为大，且行奇妙的事， 惟独你是上帝。
PS|86|11|耶和华啊，求你将你的道指教我， 我要照你的真理而行； 求你使我专心敬畏你的名！
PS|86|12|主－我的上帝啊，我要一心称谢你； 我要荣耀你的名，直到永远。
PS|86|13|因为你的慈爱在我身上浩大， 你救了我的性命免入阴间的深处。
PS|86|14|上帝啊，骄傲的人起来攻击我， 又有一群强横的人寻索我的命； 他们没有将你放在眼里。
PS|86|15|主啊，你是有怜悯，有恩惠的上帝， 不轻易发怒，并有丰盛的慈爱和信实。
PS|86|16|求你转向我，怜悯我， 将你的力量赐给仆人，拯救你使女的儿子。
PS|86|17|求你向我显出恩待我的凭据， 使恨我的人看见就羞愧， 因为你－耶和华帮助我，安慰了我。
PS|87|1|耶和华所立的根基在圣山上。
PS|87|2|耶和华爱 锡安 的门， 胜于爱 雅各 一切的住处。
PS|87|3|上帝的城啊， 有荣耀的事是指着你说的。（细拉）
PS|87|4|我要提起 拉哈伯 和 巴比伦 人， 是在认识我之中的； 看哪， 非利士 、 推罗 和 古实 人， 个个生在那里。
PS|87|5|论到 锡安 ，必有话说： “这一个、那一个都生在其中”； 而且至高者必亲自坚立这城。
PS|87|6|当耶和华记录万民的时候， 他要写出人的出生地。（细拉）
PS|87|7|歌唱的、跳舞的，都要说： “我的泉源都在你里面。”
PS|88|1|耶和华－拯救我的上帝啊， 我昼夜在你面前呼求；
PS|88|2|愿我的祷告达到你面前， 求你侧耳听我的恳求！
PS|88|3|因为我心里满了患难， 我的性命临近阴间；
PS|88|4|我与下到地府的人同列， 如同无人帮助的人一样。
PS|88|5|我被丢在死人中， 好像被杀的人躺在坟墓里， 不再被你记得， 与你的手隔绝了。
PS|88|6|你把我放在极深的地府里， 在黑暗地，在深处。
PS|88|7|你的愤怒重压我身， 你用一切的波浪困住我。（细拉）
PS|88|8|你把我所认识的人隔在远处， 使我为他们所憎恶； 我被拘禁，不能出来。
PS|88|9|我的眼睛因困苦而昏花； 耶和华啊，我天天求告你，向你举手。
PS|88|10|你岂要行奇事给死人看吗？ 阴魂还能起来称谢你吗？（细拉）
PS|88|11|你的慈爱岂能在坟墓里被人述说吗？ 你的信实岂能在冥府 被人传扬吗？
PS|88|12|你的奇事岂能在幽暗里为人所知吗？ 你的公义岂能在遗忘之地为人所识吗？
PS|88|13|耶和华啊，至于我，我要呼求你； 每早晨，我的祷告要达到你面前。
PS|88|14|耶和华啊，你为何丢弃我？ 为何转脸不顾我？
PS|88|15|我自幼受苦，几乎死亡； 你使我惊恐，烦乱不安。
PS|88|16|你的烈怒漫过我身， 你用惊吓把我除灭。
PS|88|17|这些如水终日环绕我， 一起围困我。
PS|88|18|你把我的良朋密友隔在远处， 使我所认识的人都在黑暗里 。
PS|89|1|我要歌唱耶和华的慈爱，直到永远， 我要用口将你的信实传到万代。
PS|89|2|因我曾说：“你的慈爱必建立到永远， 你的信实必坚立在天上。”
PS|89|3|“我与我所拣选的人立了约， 向我的仆人 大卫 起了誓：
PS|89|4|‘我要坚立你的后裔，直到永远， 要建立你的宝座，直到万代。’”（细拉）
PS|89|5|耶和华啊，诸天要称谢你的奇事； 在圣者的会中，要称谢你的信实。
PS|89|6|因在天空谁能比耶和华呢？ 诸神之中，谁能像耶和华呢？
PS|89|7|在圣者的会中，他是大有威严的上帝， 比在他四围所有的更可畏惧。
PS|89|8|耶和华－万军之上帝啊， 哪一个大能者像耶和华？ 你的信实在你四围。
PS|89|9|你管辖海的狂傲； 波浪翻腾，你使它平静了。
PS|89|10|你打碎了 拉哈伯 ，使它如遭刺杀的人； 你用大能的膀臂打散了你的仇敌。
PS|89|11|天属你，地也属你； 世界和其中所充满的都为你所建立。
PS|89|12|南北为你所创造； 他泊 和 黑门 都因你的名欢呼。
PS|89|13|你有大能的膀臂， 你的手有力，你的右手也高举。
PS|89|14|公义和公平是你宝座的根基， 慈爱和信实行在你前面。
PS|89|15|知道向你欢呼的，那民有福了！ 耶和华啊，他们要行走在你脸的光中。
PS|89|16|他们因你的名终日欢乐， 因你的公义得以高举。
PS|89|17|你是他们力量的荣耀。 我们的角必被高举，因为你喜爱我们。
PS|89|18|我们的盾牌是耶和华， 我们的王是 以色列 的圣者。
PS|89|19|当时，你在异象中吩咐你的圣民，说： “我已把救助之力加在壮士身上， 高举了那从百姓中所拣选的人。
PS|89|20|我寻得我的仆人 大卫 ， 用我的圣膏膏他。
PS|89|21|我的手必使他坚立， 我的膀臂也必坚固他。
PS|89|22|仇敌必不勒索他， 凶恶之子也不苦害他。
PS|89|23|我要在他面前打碎他的敌人， 击杀那些恨他的人。
PS|89|24|我的信实和我的慈爱要与他同在； 因我的名，他的角必被高举。
PS|89|25|我要使他的手伸到海上， 右手伸到河上。
PS|89|26|他要称呼我说：‘你是我的父， 是我的上帝，是拯救我的磐石。’
PS|89|27|我也要立他为长子， 为世上最高的君王。
PS|89|28|我要为他存留我的慈爱，直到永远， 我与他所立的约必坚定不移。
PS|89|29|我也要使他的后裔存到永远， 使他的宝座如天之久。
PS|89|30|“倘若他的子孙离弃我的律法， 不照我的典章行，
PS|89|31|背弃我的律例， 不遵守我的诫命，
PS|89|32|我就要用杖责罚他们的过犯， 用鞭责罚他们的罪孽。
PS|89|33|只是我不将我的慈爱全然收回， 也不叫我的信实废除。
PS|89|34|我必不毁损我的约， 也不改变我口中所出的话。
PS|89|35|我仅此一次指着自己的神圣起誓， 我绝不向 大卫 说谎！
PS|89|36|他的后裔要存到永远， 他的宝座在我面前如太阳，
PS|89|37|又如月亮永远坚立； 天上的见证是确实的。”（细拉）
PS|89|38|但你恼怒你的受膏者， 拒绝他，离弃了他。
PS|89|39|你厌恶与你仆人所立的约， 将他的冠冕践踏于地。
PS|89|40|你拆毁了他一切的围墙， 使他的堡垒变为废墟。
PS|89|41|过路的人都抢夺他， 他成了邻邦羞辱的对象。
PS|89|42|你高举了他敌人的右手， 使他所有的仇敌欢喜。
PS|89|43|你叫他的刀剑卷刃， 使他在战争中站立不住。
PS|89|44|你使他的光辉止息， 将他的宝座推倒于地。
PS|89|45|你减少他年轻的日子， 又使他蒙羞。（细拉）
PS|89|46|耶和华啊，这要到几时呢？ 你要隐藏自己到永远吗？ 你的愤怒如火焚烧要到几时呢？
PS|89|47|求你想念我的生命是何等短暂。 你创造世人，要使他们归于何等的虚空呢？
PS|89|48|谁能常活不见死亡、 救自己脱离阴间的掌控呢？（细拉）
PS|89|49|主啊，你从前凭你的信实 向 大卫 起誓要施行的慈爱在哪里呢？
PS|89|50|主啊，求你记念仆人们所受的羞辱， 记念我怎样将万族所加的羞辱都放在我的胸怀。
PS|89|51|耶和华啊，这是你仇敌所加的羞辱， 羞辱了你受膏者的脚踪。
PS|89|52|耶和华是应当称颂的，直到永远。 阿们！阿们！ 神人摩西的祈祷。
PS|90|1|主啊，你世世代代作我们的居所。
PS|90|2|诸山未曾生出， 地与世界你未曾造成， 从亘古到永远，你是上帝。
PS|90|3|你使人归于尘土，说： “世人哪，你们要归回。”
PS|90|4|在你看来，千年如已过的昨日， 又如夜间的一更。
PS|90|5|你叫他们如水冲去， 他们如睡一觉。 早晨，他们如生长的草；
PS|90|6|早晨发芽生长， 晚上割下枯干。
PS|90|7|我们因你的怒气而消灭， 因你的愤怒而惊惶。
PS|90|8|你将我们的罪孽摆在你面前， 将我们的隐恶摆在你面光之中。
PS|90|9|我们经过的日子，都在你震怒之下， 我们度尽的年岁，好像一声叹息。
PS|90|10|我们一生的年日是七十岁， 若是强壮可到八十岁； 但其中所矜夸的不过是劳苦愁烦， 转眼即逝，我们便如飞而去。
PS|90|11|谁晓得你怒气的权势？ 谁因着敬畏你而晓得你的愤怒呢？
PS|90|12|求你指教我们怎样数算自己的日子， 好叫我们得着智慧的心。
PS|90|13|耶和华啊，我们要等到几时呢？ 求你转回，怜悯你的仆人们。
PS|90|14|求你使我们早早饱得你的慈爱， 好叫我们一生一世欢呼喜乐。
PS|90|15|求你照着你使我们受苦的日子， 和我们遭难的年岁，使我们喜乐。
PS|90|16|愿你的作为向你仆人们显现， 愿你的荣耀向他们子孙显明。
PS|90|17|愿主－我们上帝的恩宠归于我们身上。 愿你坚立我们手所做的工， 我们手所做的工，愿你坚立。
PS|91|1|住在至高者隐密处的， 必住在全能者的荫下。
PS|91|2|我要向耶和华说： “我的避难所、我的山寨、 我的上帝，你是我所倚靠的。”
PS|91|3|他必救你脱离捕鸟者的罗网 和毁灭人的瘟疫。
PS|91|4|他必用自己的翎毛遮蔽你； 你要投靠在他翅膀底下， 他的信实是大小的盾牌。
PS|91|5|你必不怕黑夜的惊骇， 或是白日飞的箭，
PS|91|6|也不怕黑夜流行的瘟疫， 或是午间灭人的灾害。
PS|91|7|虽有千人仆倒在你旁边， 万人仆倒在你右边， 这灾却不得临近你。
PS|91|8|你惟亲眼观看， 见恶人遭报。
PS|91|9|因为耶和华是我的避难所， 你以至高者为居所，
PS|91|10|祸患必不临到你， 灾害也不挨近你的帐棚。
PS|91|11|因他要为你命令他的使者， 在你所行的一切道路上保护你。
PS|91|12|他们要用手托住你， 免得你的脚碰在石头上。
PS|91|13|你要踹踏狮子和毒蛇， 践踏少壮狮子和大蛇。
PS|91|14|“因为他专心爱我，我要搭救他； 因为他认识我的名，我要把他安置在高处。
PS|91|15|他若求告我，我就应允他； 他在急难中，我与他同在； 我要搭救他，使他尊贵。
PS|91|16|我要使他享足长寿， 将我的救恩显明给他。”
PS|92|1|这是多么好啊！ 称谢耶和华， 歌颂你至高者的名，
PS|92|2|早晨传扬你的慈爱， 每夜传扬你的信实。
PS|92|3|用十弦的乐器和瑟， 用琴优雅的声音；
PS|92|4|因你－耶和华藉着你的作为使我高兴， 我要因你手的工作欢呼。
PS|92|5|耶和华啊，你的工作何其大！ 你的心思极其深！
PS|92|6|畜牲一般的人不晓得， 愚昧人也不明白。
PS|92|7|恶人虽茂盛如草， 作恶的人虽全都兴旺， 他们却要灭亡， 直到永远。
PS|92|8|耶和华啊，惟有你是至高， 直到永远。
PS|92|9|耶和华啊，看哪，你的仇敌， 看哪，你的仇敌都要灭亡； 作恶的全都要离散。
PS|92|10|你却高举了我的角，如野牛的角； 我是被新油膏抹的。
PS|92|11|我的眼睛看见我的仇敌遭报， 我的耳朵听见那些起来攻击我的恶人受罚。
PS|92|12|义人要兴旺如棕树， 生长如 黎巴嫩 的香柏树。
PS|92|13|他们栽于耶和华的殿中， 发旺在我们上帝的院里。
PS|92|14|他们发白的时候仍结果子， 而且鲜美多汁，
PS|92|15|好显明耶和华是正直的； 他是我的磐石，在他毫无不义。
PS|93|1|耶和华作王！ 他以威严为衣穿上； 耶和华以能力为衣，以能力束腰， 世界就坚定，不得动摇。
PS|93|2|你的宝座从太初立定， 你从亘古就有。
PS|93|3|耶和华啊，大水扬起， 大水发声，大水澎湃。
PS|93|4|耶和华在高处大有威力， 胜过诸水的响声，洋海的大浪。
PS|93|5|耶和华啊，你的法度最为确定； 你的殿宜称为圣，直到永远。
PS|94|1|耶和华啊，你是伸冤的上帝； 伸冤的上帝啊，求你发出光来！
PS|94|2|审判世界的主啊，求你挺身而立， 使骄傲的人受应得的报应！
PS|94|3|耶和华啊，恶人夸胜要到几时呢？ 要到几时呢？
PS|94|4|他们咆哮，说狂妄的话， 作恶的人全都夸耀自己。
PS|94|5|耶和华啊，他们强压你的百姓， 苦害你的产业。
PS|94|6|他们杀死寡妇和寄居的人， 又杀害孤儿。
PS|94|7|他们说：“耶和华必不看见， 雅各 的上帝必不留意。”
PS|94|8|百姓中像畜牲一般的人当思想， 你们愚昧人要到几时才有智慧呢？
PS|94|9|造耳朵的，难道自己听不见吗？ 造眼睛的，难道自己看不见吗？
PS|94|10|管教列国的，就是叫人得知识的， 难道自己不惩治人吗？
PS|94|11|耶和华知道人的意念是虚妄的。
PS|94|12|耶和华啊，你所管教、 用律法教导的人有福了！
PS|94|13|你使他在遭难的日子仍得平安， 直到为恶人挖好了坑。
PS|94|14|因为耶和华必不丢弃他的百姓， 也不离弃他的产业。
PS|94|15|审判要回复公义， 心里正直的，都必跟随它。
PS|94|16|谁肯为我起来攻击邪恶的？ 谁肯为我站起抵挡作恶的？
PS|94|17|若不是耶和华帮助我， 我早就住在寂静 之中了。
PS|94|18|我若说：“我失了脚！” 耶和华啊，你的慈爱必扶持我。
PS|94|19|我心里多忧多疑， 你的安慰使我欢乐。
PS|94|20|那藉着律例玩弄奸恶、 以权位肆行残害的，岂能与你交往呢？
PS|94|21|他们大家聚集攻击义人， 将无辜的人定了死罪。
PS|94|22|但耶和华向来作我的碉堡， 我的上帝作了我投靠的磐石。
PS|94|23|他叫他们的罪孽归到自己身上， 要因他们的邪恶剪除他们； 耶和华－我们的上帝要把他们剪除。
PS|95|1|来啊，我们要向耶和华歌唱， 向拯救我们的磐石欢呼！
PS|95|2|我们要以感谢来到他面前， 用诗歌向他欢呼！
PS|95|3|因耶和华是伟大的上帝， 是超越万神的大君王。
PS|95|4|地的深处在他手中； 山的高峰也属他。
PS|95|5|海洋属他，是他造的； 旱地也是他手造成的。
PS|95|6|来啊，我们要俯伏敬拜， 在造我们的耶和华面前跪拜。
PS|95|7|因为他是我们的上帝； 我们是他草场的百姓，是他手中的羊。 惟愿你们今天听他的话！
PS|95|8|你们不可硬着心，像在 米利巴 ， 就是在旷野 玛撒 的日子。
PS|95|9|那时，你们的祖宗试我，探我， 并且观看我的作为。
PS|95|10|四十年之久，我厌烦那世代，说： “这是心里迷糊的百姓， 竟不知道我的道路！”
PS|95|11|所以，我在怒中起誓： “他们断不可进入我的安息！”
PS|96|1|你们要向耶和华唱新歌！ 全地都要向耶和华歌唱！
PS|96|2|要向耶和华歌唱，称颂他的名！ 天天传扬他的救恩！
PS|96|3|在列国中述说他的荣耀！ 在万民中述说他的奇事！
PS|96|4|因耶和华本为大，当受极大的赞美； 他在万神之上，当受敬畏。
PS|96|5|因万民的神明都属虚无； 惟独耶和华创造诸天。
PS|96|6|有尊荣和威严在他面前， 有能力与华美在他圣所。
PS|96|7|民中的万族啊，要将荣耀、能力归给耶和华， 都归给耶和华！
PS|96|8|要将耶和华的名所当得的荣耀归给他， 拿供物来进入他的院宇。
PS|96|9|当敬拜神圣荣耀的耶和华 ， 全地都要在他面前战抖！
PS|96|10|要在列国中说：“耶和华作王了！ 世界坚定，不得动摇； 他要按公正审判万民。”
PS|96|11|愿天欢喜，愿地快乐！ 愿海和其中所充满的澎湃！
PS|96|12|愿田和其中所有的都欢乐！ 那时，林中的树木都要在耶和华面前欢呼。
PS|96|13|因为他来了，他来要审判全地。 他要按公义审判世界， 按信实审判万民。
PS|97|1|耶和华作王！愿地快乐！ 愿众海岛欢喜！
PS|97|2|密云和幽暗在他四围， 公义和公平是他宝座的根基。
PS|97|3|烈火在他前头行， 烧灭他四围的敌人。
PS|97|4|他的闪电光照世界， 大地看见就震动。
PS|97|5|诸山见耶和华的面， 就是全地之主的面，就如蜡熔化。
PS|97|6|诸天表明他的公义， 万民看见他的荣耀。
PS|97|7|愿所有事奉雕刻偶像、 靠虚无神明自夸的，都蒙羞愧。 万神哪，你们都当拜他。
PS|97|8|耶和华啊，因你的判断， 锡安 听见就欢喜； 犹大 的城镇 也都快乐。
PS|97|9|因为你－耶和华至高，超乎全地； 受尊崇，远超万神之上。
PS|97|10|你们爱耶和华的，都当恨恶罪恶； 他保护圣民的性命， 搭救他们脱离恶人的手。
PS|97|11|散播亮光是为义人 ， 喜乐归于心里正直的人。
PS|97|12|义人哪，你们当靠耶和华欢喜， 当颂扬他神圣的名字 。
PS|98|1|你们要向耶和华唱新歌！ 因为他行过奇妙的事， 他的右手和圣臂施行救恩。
PS|98|2|耶和华显明了他的救恩， 在列国眼前显出公义；
PS|98|3|记念他对 以色列 家的慈爱和信实。 地的四极都看见我们上帝的救恩。
PS|98|4|全地都要向耶和华欢呼， 要扬声，欢唱，歌颂！
PS|98|5|用琴歌颂耶和华， 用琴和诗歌的声音歌颂他！
PS|98|6|用号筒和角声， 在大君王耶和华面前欢呼！
PS|98|7|愿海和其中所充满的澎湃， 愿世界和住在其间的发声。
PS|98|8|愿大水拍掌， 愿诸山在耶和华面前一同欢呼；
PS|98|9|因为他来要审判全地。 他要按公义审判世界， 按公正审判万民。
PS|99|1|耶和华作王，万民当战抖！ 他坐在基路伯的宝座上，地当动摇。
PS|99|2|耶和华在 锡安 为大， 他超越万民之上。
PS|99|3|愿他们颂扬他大而可畏的名， 他本为圣！
PS|99|4|喜爱公平、大能的王啊，你坚立公正， 在 雅各 中施行公平和公义。
PS|99|5|当尊崇耶和华－我们的上帝， 在他脚凳前下拜。 他本为圣！
PS|99|6|在他的祭司中有 摩西 和 亚伦 ， 在求告他名的人中有 撒母耳 。 他们求告耶和华，他就应允他们。
PS|99|7|他在云柱中向他们说话， 他们遵守他的法度和他所赐给他们的律例。
PS|99|8|耶和华－我们的上帝啊，你应允了他们； 你是赦免他们的上帝， 却按他们所做的报应他们。
PS|99|9|当尊崇耶和华－我们的上帝， 在他的圣山下拜， 因为耶和华－我们的上帝本为圣！
PS|100|1|普天下当向耶和华欢呼！
PS|100|2|当乐意事奉耶和华， 当欢唱来到他面前！
PS|100|3|当认识耶和华是上帝！ 我们是他造的，也是属他的； 我们是他的民，是他草场的羊。
PS|100|4|当称谢进入他的门， 当赞美进入他的院。 当感谢他，称颂他的名！
PS|100|5|因为耶和华本为善； 他的慈爱存到永远， 他的信实直到万代。
PS|101|1|我要歌唱慈爱和公平， 耶和华啊，我要向你歌颂！
PS|101|2|我要用智慧行完全的道。 你几时到我这里来呢？ 我要以纯正的心行在我家中。
PS|101|3|邪僻的事，我都不摆在我眼前； 悖逆的人所做的事，我甚恨恶， 不容沾在我身上。
PS|101|4|歪曲的心思，我必远离； 邪恶的事情，我不知道。
PS|101|5|暗中谗害他邻居的，我必将他灭绝； 眼目高傲、心里骄纵的，我必不容忍。
PS|101|6|我眼要看顾地上诚实可靠的人，使他们与我同住； 行正直路的，他要侍候我。
PS|101|7|行诡诈的，必不得住在我家里； 说谎言的，必不得立在我眼前。
PS|101|8|我每日早晨要灭绝地上所有的恶人， 把作恶的从耶和华的城里全都剪除。
PS|102|1|耶和华啊，求你听我的祷告， 愿我的呼求达到你面前！
PS|102|2|我急难的日子，求你不要转脸不顾我！ 我呼求的日子，求你向我侧耳，快快应允我！
PS|102|3|因为我的年日在烟中消失 ， 我的骨头如火把烧着。
PS|102|4|我的心如草被踩碎而枯干， 甚至我忘记吃饭。
PS|102|5|因我叹息的声音， 我的肉紧贴骨头。
PS|102|6|我如同旷野的鹈鹕， 好像荒地的猫头鹰。
PS|102|7|我清醒难以入眠， 如同房顶上孤单的麻雀。
PS|102|8|我的仇敌整日辱骂我， 向我叫号的人指着我赌咒。
PS|102|9|我吃灰烬如同吃饭， 我喝的有眼泪搀杂。
PS|102|10|这都因你的恼恨和愤怒， 你把我举起，又把我摔下。
PS|102|11|我的年日如夕阳， 我也如草枯干。
PS|102|12|惟你－耶和华必永远坐在宝座上， 你的名 存到万代。
PS|102|13|你必起来怜悯 锡安 ； 因现在是可怜它的时候， 因所定的日期已经到了。
PS|102|14|你的仆人们喜爱 锡安 的石头， 怜悯它的尘土。
PS|102|15|列国要敬畏耶和华的名， 地上众王都要敬畏你的荣耀。
PS|102|16|因为耶和华建造了 锡安 ， 在他的荣耀里显现。
PS|102|17|他垂听穷乏人的祷告， 不藐视他们的祈求。
PS|102|18|这必为后代的人记下， 将来受造的百姓要赞美耶和华。
PS|102|19|因为他从至高的圣所垂看； 耶和华从天向地观看，
PS|102|20|要垂听被囚之人的叹息， 要释放将死的人，
PS|102|21|使人在 锡安 传扬耶和华的名， 在 耶路撒冷 传扬赞美他的话，
PS|102|22|就是在万民和列国 聚集事奉耶和华的时候。
PS|102|23|他使我的力量半途衰弱， 使我的年日短少。
PS|102|24|我说：“我的上帝啊， 不要使我中年去世。 你的年数世世无穷！”
PS|102|25|你起初立了地的根基， 天也是你手所造的。
PS|102|26|天地都会消灭，你却长存； 天地都会像外衣渐渐旧了。 你要将天地如内衣更换， 天地就都改变了。
PS|102|27|惟有你永不改变， 你的年数没有穷尽。
PS|102|28|你仆人的子孙要安然居住， 他们的后裔要坚立在你面前。
PS|103|1|我的心哪，你要称颂耶和华！ 凡在我里面的，都要称颂他的圣名！
PS|103|2|我的心哪，你要称颂耶和华！ 不可忘记他一切的恩惠！
PS|103|3|他赦免你一切的罪孽， 医治你一切的疾病。
PS|103|4|他救赎你的命脱离地府， 以仁爱和怜悯为你的冠冕。
PS|103|5|他用美物使你的生命 得以满足， 以致你如鹰返老还童。
PS|103|6|耶和华施行公义， 为所有受欺压的人伸冤。
PS|103|7|他使 摩西 知道他的法则， 使 以色列 人晓得他的作为。
PS|103|8|耶和华有怜悯，有恩惠， 不轻易发怒，且有丰盛的慈爱。
PS|103|9|他不长久责备， 也不永远怀怒。
PS|103|10|他没有按我们的罪待我们， 也没有照我们的罪孽报应我们。
PS|103|11|天离地何等的高， 他的慈爱向敬畏他的人也是何等的大！
PS|103|12|东离西有多远， 他叫我们的过犯离我们也有多远！
PS|103|13|父亲怎样怜悯他的儿女， 耶和华也怎样怜悯敬畏他的人！
PS|103|14|因为他知道我们的本体， 思念我们不过是尘土。
PS|103|15|至于世人，他的年日如草一样。 他兴旺如野地的花，
PS|103|16|经风一吹，就归无有， 它的原处也不再认识它。
PS|103|17|但耶和华的慈爱归于敬畏他的人， 从亘古到永远； 他的公义也归于子子孙孙，
PS|103|18|就是那些遵守他的约、 记念他的训词而遵行的人。
PS|103|19|耶和华在天上立定宝座， 他的国统管万有。
PS|103|20|听从他命令、成全他旨意、 有大能的天使啊，你们都要称颂耶和华！
PS|103|21|你们行他所喜悦的， 作他诸军，作他仆役的啊，都要称颂耶和华！
PS|103|22|你们一切被他造的， 在他所治理的各处， 都要称颂耶和华！ 我的心哪，你要称颂耶和华！
PS|104|1|我的心哪，你要称颂耶和华！ 耶和华－我的上帝啊，你为至大！ 你以尊荣威严为衣，
PS|104|2|披上亮光，如披外袍， 铺张穹苍，如铺幔子，
PS|104|3|在水中立楼阁的栋梁， 用云彩为车辇， 藉着风的翅膀而行，
PS|104|4|以风为使者， 以火焰为仆役，
PS|104|5|将地立在根基上， 使地永不动摇。
PS|104|6|你用深水遮盖地面，犹如衣裳； 诸水高过山岭。
PS|104|7|你的斥责一发，水就奔逃； 你的雷声一发，水就奔流。
PS|104|8|诸山上升，诸谷下沉， 归你为它所立定之地。
PS|104|9|你定了界限，使水不能超越， 不再转回淹没大地。
PS|104|10|耶和华使泉源涌在山谷， 流在山间，
PS|104|11|使野地的走兽有水喝， 野驴得解其渴。
PS|104|12|天上的飞鸟在水旁住宿， 在枝干间啼叫。
PS|104|13|他从楼阁中浇灌山岭； 因他作为的功效，地就丰足。
PS|104|14|他使草生长，给牲畜吃， 使菜蔬生长，供给人用 ， 使人从地里得食物，
PS|104|15|得酒能悦人心， 得油能润人面， 得粮能养人心。
PS|104|16|佳美的树木， 就是耶和华所栽种的 黎巴嫩 的香柏树， 都满了汁浆。
PS|104|17|雀鸟在其上搭窝， 鹳以松树 为家。
PS|104|18|高山为野山羊的居所， 岩石为石的藏身处。
PS|104|19|你安置月亮以定季节， 太阳自知沉落。
PS|104|20|你造黑暗为夜， 林中的百兽就都爬出来。
PS|104|21|少壮狮子吼叫觅食， 向上帝寻求食物。
PS|104|22|太阳一出，兽就躲避， 躺卧在洞里。
PS|104|23|人出去做工， 劳碌直到晚上。
PS|104|24|耶和华啊，你所造的何其多！ 都是你用智慧造成的， 全地遍满了你所造之物。
PS|104|25|那里有海，又大又广， 其中有无数的动物， 大小活物都有。
PS|104|26|那里有船行走， 有你所造的 力威亚探 悠游在其中。
PS|104|27|这些都仰望你按时给它们食物。
PS|104|28|你给它们，它们就拾起来； 你张手，它们就饱得美食。
PS|104|29|你转脸，它们就惊惶； 你收回它们的气，它们就死亡，归于尘土。
PS|104|30|你差遣你的灵，它们就受造； 你使地面更换为新。
PS|104|31|愿耶和华的荣耀存到永远！ 愿耶和华喜爱自己所造的！
PS|104|32|他看地，地便震动； 他摸山，山就冒烟。
PS|104|33|我一生要向耶和华唱诗！ 我还活的时候，要向我的上帝歌颂！
PS|104|34|愿他悦纳我的默念！ 我要因耶和华欢喜！
PS|104|35|愿罪人从世上消灭！ 愿恶人归于无有！ 我的心哪，你要称颂耶和华！ 哈利路亚 ！
PS|105|1|你们要称谢耶和华，求告他的名， 在万民中传扬他的作为！
PS|105|2|要向他唱诗，向他歌颂， 述说他一切奇妙的作为！
PS|105|3|要夸耀他的圣名！ 愿寻求耶和华的人心中欢喜！
PS|105|4|要寻求耶和华与他的能力， 时常寻求他的面。
PS|105|5|他仆人 亚伯拉罕 的后裔， 他所拣选 雅各 的子孙哪， 要记念他奇妙的作为和他的奇事， 并他口中的判语。
PS|105|6|
PS|105|7|他是耶和华－我们的上帝， 全地都有他的判断。
PS|105|8|他记念他的约，直到永远； 记念他吩咐的话，直到千代，
PS|105|9|就是与 亚伯拉罕 所立的约， 向 以撒 所起的誓。
PS|105|10|他将这约向 雅各 定为律例， 向 以色列 定为永远的约，
PS|105|11|说：“我必将 迦南 地赐给你， 作你们应得的产业。”
PS|105|12|当时，他们人丁有限， 数目稀少，在那地寄居。
PS|105|13|他们从这邦游到那邦， 从这国去到另一民族。
PS|105|14|他不容人欺负他们， 为他们的缘故责备君王：
PS|105|15|“不可伤害我的受膏者， 也不可恶待我的先知。”
PS|105|16|他命饥荒降在那地， 断绝日用的粮食 ，
PS|105|17|在他们以先差遣一个人前往， 约瑟 被卖为奴。
PS|105|18|人用脚镣伤他的脚， 他被铁的项链捆锁。
PS|105|19|耶和华的话试炼他， 直等所说的应验了。
PS|105|20|王差人将他解开， 治理万民的把他释放，
PS|105|21|立他为王家之主， 掌管他一切所有的，
PS|105|22|使他随意捆绑他的臣宰， 将智慧教导他的长老。
PS|105|23|以色列 也到了 埃及 ， 雅各 在 含 地寄居。
PS|105|24|耶和华使他的百姓生养众多， 使他们比敌人强盛，
PS|105|25|他使敌人的心转去恨他的百姓， 用诡计待他的仆人。
PS|105|26|他差遣他的仆人 摩西 和他所拣选的 亚伦 ，
PS|105|27|在敌人中间显他的神迹， 在 含 地显他的奇事。
PS|105|28|他差遣黑暗，就有黑暗； 他们没有违背他的话。
PS|105|29|他使 埃及 的水变为血， 令他们的鱼死了。
PS|105|30|在他们的地上，青蛙多多滋生， 王宫的内室也是如此。
PS|105|31|他一吩咐，苍蝇就成群飞来， 并有蚊子进入他们四境。
PS|105|32|他给他们降下冰雹为雨， 在他们的地上降下火焰。
PS|105|33|他击打他们的葡萄树和无花果树， 毁坏他们境内的树木。
PS|105|34|他一吩咐，就有蝗虫蝻子上来， 不计其数，
PS|105|35|吃光他们地上各样的菜蔬， 吞尽他们田地的出产。
PS|105|36|他又击杀他们国内 所有的长子， 就是他们强壮时头生的。
PS|105|37|他却带领自己的百姓带着金子银子出来， 他支派中没有一个走不动的。
PS|105|38|他们出来的时候， 埃及 人就欢喜； 因为 埃及 人惧怕他们。
PS|105|39|他铺张云彩当遮蔽， 夜间使火光照。
PS|105|40|他们祈求，他就使鹌鹑飞来， 并用天上的粮食使他们饱足。
PS|105|41|他敲开磐石，水就涌出； 在干旱之处，水流成河。
PS|105|42|这都因他记念他的圣言 和他的仆人 亚伯拉罕 。
PS|105|43|他带领自己的百姓欢乐而出， 带领自己的选民欢呼前往。
PS|105|44|他把列国的地赐给他们， 他们就承受万民劳碌得来的，
PS|105|45|好让他们遵他的律例， 守他的律法。 哈利路亚！
PS|106|1|哈利路亚！ 你们要称谢耶和华，因他本为善， 他的慈爱永远长存！
PS|106|2|谁能传扬耶和华的大能？ 谁能表明他一切的美德？
PS|106|3|凡遵守公平、常行公义的， 这人有福了！
PS|106|4|耶和华啊，你恩待你百姓的时候，求你记念我； 你拯救他们的时候，求你眷顾我，
PS|106|5|好使我经历你选民的福分， 享受你国民的喜乐， 与你的产业一同夸耀。
PS|106|6|我们与我们的祖宗一同犯罪， 偏邪行恶。
PS|106|7|我们的祖宗在 埃及 不明白你的奇事， 不记念你丰盛的慈爱， 反倒在 红海 行了悖逆。
PS|106|8|然而，他因自己的名拯救他们， 为要彰显他的大能。
PS|106|9|他斥责 红海 ，海就干了， 带领他们走过深海，如走旷野。
PS|106|10|他拯救他们脱离恨他们之人的手， 从仇敌手中救赎他们。
PS|106|11|水淹没他们的敌人， 没有一个存留。
PS|106|12|那时，他们才信他的话， 歌唱赞美他。
PS|106|13|很快地，他们就忘了他的作为， 不仰望他的指引，
PS|106|14|反倒在旷野起了贪婪之心， 在荒地试探上帝。
PS|106|15|他将他们所求的赐给他们， 却使他们心灵软弱。
PS|106|16|他们在营中嫉妒 摩西 和耶和华的圣者 亚伦 。
PS|106|17|地就裂开，吞下 大坍 ， 掩盖 亚比兰 一伙的人。
PS|106|18|有火在他们党中点燃， 有火焰烧毁了恶人。
PS|106|19|他们在 何烈山 造了牛犊， 叩拜铸成的像，
PS|106|20|将他们荣耀的主 换为吃草之牛的像，
PS|106|21|忘了上帝－他们的救主， 就是曾在 埃及 行大事，
PS|106|22|在 含 地行奇事， 在 红海 行可畏之事的那位。
PS|106|23|因此，他说要灭绝他们； 若非他所拣选的 摩西 在他面前站在破裂之处， 使他的愤怒转消， 恐怕他就灭绝他们了。
PS|106|24|他们又藐视那美地， 不信他的话，
PS|106|25|在自己帐棚内发怨言， 不听耶和华的声音。
PS|106|26|所以他向他们起誓， 必叫他们倒在旷野，
PS|106|27|叫他们的后裔倒在列国之中， 分散在各地。
PS|106|28|他们又与 巴力．毗珥 连合， 吃了祭死人的物。
PS|106|29|他们这样行，惹耶和华发怒， 就有瘟疫流行在他们中间。
PS|106|30|那时， 非尼哈 起而干预， 瘟疫这才止息。
PS|106|31|那就算他为义， 世世代代，直到永远。
PS|106|32|他们在 米利巴 水又惹耶和华发怒， 甚至 摩西 也因他们的缘故受亏损，
PS|106|33|是因他们触怒了他的灵， 摩西就用嘴说了急躁的话。
PS|106|34|他们不照耶和华所吩咐的 灭绝外邦人，
PS|106|35|反倒与列国相交， 学习他们的行为，
PS|106|36|事奉他们的偶像， 这就成了自己的圈套。
PS|106|37|他们把自己的儿女祭祀鬼魔，
PS|106|38|流无辜人的血， 就是自己儿女的血， 用他们祭祀 迦南 的偶像， 那地就被血玷污了。
PS|106|39|这样，他们被自己所做的玷污了， 在行为上犯了淫乱。
PS|106|40|耶和华的怒气向他的百姓发作， 他憎恶自己的产业，
PS|106|41|将他们交在外邦人手里， 恨他们的人就辖制他们。
PS|106|42|他们的仇敌欺压他们， 他们伏在敌人手下。
PS|106|43|他屡次搭救他们， 他们却图谋悖逆， 就因自己的罪孽降为卑下。
PS|106|44|然而，他听见他们哀告的时候， 就眷顾他们的急难，
PS|106|45|为了他们，他记念自己的约， 照他丰盛的慈爱改变心意，
PS|106|46|使他们在凡掳掠他们的人面前蒙怜悯。
PS|106|47|耶和华－我们的上帝啊，求你拯救我们， 从列国中召集我们， 我们好颂扬你的圣名， 以赞美你为夸胜。
PS|106|48|耶和华－ 以色列 的上帝是应当称颂的， 从亘古直到永远。 愿全体百姓都说：“阿们！” 哈利路亚！
PS|107|1|你们要称谢耶和华，因他本为善， 他的慈爱永远长存！
PS|107|2|愿耶和华救赎的百姓说这话， 就是他从敌人手中所救赎，
PS|107|3|从各地，从东从西， 从北从海那边召集来的。
PS|107|4|他们在旷野、在荒地飘流， 找不到可居住的城，
PS|107|5|又饥又渴， 心里发昏。
PS|107|6|于是他们在急难中哀求耶和华， 他就搭救他们脱离祸患，
PS|107|7|又领他们行走直路， 前往可居住的城。
PS|107|8|但愿人因耶和华的慈爱 和他向人所做的奇事都称谢他；
PS|107|9|因他使心里渴慕的人得以满足， 使饥饿的人得饱美食。
PS|107|10|那些坐在黑暗中、死荫里的人， 被困苦和铁链捆锁，
PS|107|11|是因他们违背上帝的言语， 藐视至高者的旨意。
PS|107|12|所以，他用劳苦制伏他们的心； 他们仆倒，无人扶助。
PS|107|13|于是他们在急难中哀求耶和华， 他就拯救他们脱离祸患。
PS|107|14|他从黑暗中、从死荫里领他们出来， 扯断他们的捆绑。
PS|107|15|但愿人因耶和华的慈爱 和他向人所做的奇事都称谢他；
PS|107|16|因为他打破了铜门， 砍断了铁闩。
PS|107|17|愚妄人因自己叛逆的行径 和自己的罪孽受苦楚。
PS|107|18|他们心里厌恶各样的食物， 就临近死亡之门。
PS|107|19|于是他们在急难中哀求耶和华， 他就拯救他们脱离祸患。
PS|107|20|他发出自己的话语医治他们， 救他们脱离阴府。
PS|107|21|但愿人因耶和华的慈爱 和他向人所做的奇事都称谢他。
PS|107|22|愿他们以感谢为祭献给他， 欢呼述说他的作为！
PS|107|23|那些搭船出海， 在大水中做生意的，
PS|107|24|他们看见耶和华的作为， 并他在深海中的奇事。
PS|107|25|他一出令，狂风卷起， 波浪翻腾。
PS|107|26|他们上到天空，下到海底， 他们的心因患难而消沉。
PS|107|27|他们摇摇晃晃，东倒西歪，好像醉酒的人， 他们的智慧无法可施。
PS|107|28|于是他们在急难中哀求耶和华， 他就领他们脱离祸患。
PS|107|29|他使狂风止息， 波浪平静，
PS|107|30|既平静了，他们就欢喜， 他就领他们到想要去的海港。
PS|107|31|但愿人因耶和华的慈爱 和他向人所做的奇事都称谢他。
PS|107|32|愿他们在百姓的会中尊崇他， 在长老的座位上赞美他！
PS|107|33|他使江河变为旷野， 叫水泉变为干涸之地，
PS|107|34|使肥沃之地变为荒芜的盐地， 都因当地居民的邪恶。
PS|107|35|他使旷野变为水潭， 叫旱地变为水泉，
PS|107|36|使饥饿的人住在那里， 建造可居住的城，
PS|107|37|又种田地，栽葡萄园， 得享所出产的果实。
PS|107|38|他赐福给他们，使他们生养众多， 也不叫他们的牲畜减少。
PS|107|39|但他们因欺压、患难、愁苦， 人口减少而且卑微。
PS|107|40|他使贵族蒙羞受辱， 使他们迷失在荒凉无路之地；
PS|107|41|却将穷乏人安置在高处，脱离苦难， 使他的家属多如羊群。
PS|107|42|正直的人看见就欢喜， 罪孽之辈却要哑口无言。
PS|107|43|凡有智慧的必在这些事上留心， 他必思想耶和华的慈爱。
PS|108|1|上帝啊，我心坚定； 我口 要唱诗歌颂！
PS|108|2|琴瑟啊，当醒起！ 我要唤起曙光！
PS|108|3|耶和华啊，我要在万民中称谢你， 在万族中歌颂你！
PS|108|4|因为你的慈爱大过诸天， 你的信实达到穹苍。
PS|108|5|上帝啊，愿你崇高过于诸天！ 愿你的荣耀高过全地！
PS|108|6|求你应允我，用右手施行拯救， 好让你所亲爱的人得救。
PS|108|7|上帝在他的圣所 说： “我要欢乐； 要划分 示剑 ， 丈量 疏割谷 。
PS|108|8|基列 是我的， 玛拿西 是我的， 以法莲 是护卫我头的， 犹大 是我的权杖。
PS|108|9|摩押 是我的沐浴盆， 我要向 以东 扔鞋， 我必因胜 非利士 而欢呼。”
PS|108|10|谁能领我进坚固城？ 谁能引我到 以东 地？
PS|108|11|上帝啊，你真的丢弃了我们吗？ 上帝啊，你不和我们的军队同去吗？
PS|108|12|求你帮助我们攻击敌人， 因为人的帮助是枉然的。
PS|108|13|我们倚靠上帝才得施展大能， 因为践踏我们敌人的就是他。
PS|109|1|我所赞美的上帝啊， 求你不要闭口不言。
PS|109|2|因为恶人的嘴和诡诈人的口张开攻击我， 他们用撒谎的舌头对我说话。
PS|109|3|他们围绕我，说怨恨的话， 又无故地攻打我。
PS|109|4|他们与我作对回报我的爱， 但我专心祈祷。
PS|109|5|他们向我以恶报善， 以恨报爱。
PS|109|6|求你派恶人辖制他， 派对头站在他右边！
PS|109|7|他受审判的时候， 愿他背负罪名而出！ 愿他的祈祷反成为罪！
PS|109|8|愿他的年岁短少！ 愿别人得他的职分！
PS|109|9|愿他的儿女成为孤儿， 他的妻子成为寡妇！
PS|109|10|愿他的儿女飘流讨饭， 从荒凉之处出来求乞 ！
PS|109|11|愿债主牢笼他一切所有的！ 愿陌生人抢走他劳碌得来的！
PS|109|12|愿无人向他布施恩惠， 无人恩待他的孤儿！
PS|109|13|愿他的后人断绝， 名字被涂去，不传于下代！
PS|109|14|愿耶和华记得他祖宗的罪孽， 不涂去他母亲的罪过！
PS|109|15|愿这些罪常在耶和华面前！ 愿他们的名字 从地上除灭！
PS|109|16|因为他从未想过要施恩， 却迫害困苦贫穷的和伤心的人， 把他们处死。
PS|109|17|他爱咒骂，咒骂就临到他； 他不喜爱祝福，祝福就远离他！
PS|109|18|他拿咒骂当衣服穿上； 这咒骂就如水进到他里面， 如油进入他骨头。
PS|109|19|愿这咒骂当他遮身的衣服， 作他经常束腰的带子！
PS|109|20|这就是那些与我作对、用恶言议论我的人 从耶和华所受的报应。
PS|109|21|但是你，主－耶和华啊， 求你因你的名采取行动； 因你的慈爱美好，求你搭救我！
PS|109|22|因为我困苦贫穷， 内心受伤。
PS|109|23|我如日影偏斜而去， 如蝗虫被抖出来。
PS|109|24|我因禁食，膝盖软弱； 我身体消瘦，不再丰润。
PS|109|25|我受他们的羞辱， 他们看见我就摇头。
PS|109|26|耶和华－我的上帝啊，求你帮助我， 照你的慈爱拯救我，
PS|109|27|好让他们知道这是你的手， 是你－耶和华所做的事。
PS|109|28|任凭他们咒骂，你却要赐福； 他们几时起来就必蒙羞， 你的仆人却要欢喜。
PS|109|29|愿与我作对的人披戴羞辱！ 愿他们以自己的羞愧作外袍遮身！
PS|109|30|我要用口极力称谢耶和华， 我要在众人中间赞美他；
PS|109|31|因为他必站在贫穷人的右边， 救他脱离定他死罪的人。
PS|110|1|耶和华对我主说： “你坐在我的右边， 等我使你仇敌作你的脚凳。”
PS|110|2|耶和华必使你从 锡安 伸出你能力的权杖； 你务要在仇敌中掌权。
PS|110|3|你在圣山上 掌权的日子， 你的子民必甘心跟随 ； 从晨曦初现， 你就有清晨 的甘露。
PS|110|4|耶和华起了誓，绝不改变： “你是照着 麦基洗德 的体系永远为祭司。”
PS|110|5|在你右边的主， 当他发怒的日子，必打伤列王。
PS|110|6|他要审判列国， 尸首就布满各处； 他要痛击遍地的领袖。
PS|110|7|他要喝路旁的河水， 因此必抬起头来。
PS|111|1|哈利路亚！ 我要在正直人的大会和会众中 一心称谢耶和华。
PS|111|2|耶和华的作为本为大， 被所有喜爱的人所探寻。
PS|111|3|他所做的是尊荣和威严， 他的公义存到永远。
PS|111|4|他行了奇事，使人记念； 耶和华有恩惠，有怜悯。
PS|111|5|他赐粮食给敬畏他的人， 他必永远记念他的约。
PS|111|6|他向百姓显出大能的作为， 将列国赐给他们为业。
PS|111|7|他手所做的信实公平， 他的训词全然可靠，
PS|111|8|是永永远远坚定的， 是按信实正直设立的。
PS|111|9|他向百姓施行救赎， 颁布他的约，直到永远； 他的名圣而可畏。
PS|111|10|敬畏耶和华是智慧的开端， 凡遵行他命令的有美好的见识。 耶和华是永远当赞美的！
PS|112|1|哈利路亚！ 敬畏耶和华，甚喜爱他命令的， 这人有福了！
PS|112|2|他的后裔在世必强盛， 正直人的后代必蒙福。
PS|112|3|他的家中有金银财宝， 他的义行存到永远。
PS|112|4|正直人在黑暗中有光向他照耀， 他有恩惠，有怜悯，有公义。
PS|112|5|施恩与人、借贷与人、秉公处事的人 必享美福，
PS|112|6|他永不动摇。 义人被记念，直到永远。
PS|112|7|他不惧怕凶恶的信息， 他的心坚定，倚靠耶和华。
PS|112|8|他的心确定，总不惧怕， 直到他看见敌人遭报。
PS|112|9|他施舍，赒济贫穷， 他的义行存到永远， 他的角必被高举，大有荣耀。
PS|112|10|恶人看见就愤怒，必咬牙而消亡， 恶人的心愿要归于幻灭。
PS|113|1|哈利路亚！ 耶和华的仆人哪，你们要赞美， 赞美耶和华的名！
PS|113|2|耶和华的名是应当称颂的， 从今时直到永远！
PS|113|3|从日出之地到日落之处， 耶和华的名是应当赞美的！
PS|113|4|耶和华超乎万国之上， 他的荣耀高过诸天。
PS|113|5|谁像耶和华－我们的上帝呢？ 他坐在至高之处，
PS|113|6|自己谦卑， 观看天上地下的事。
PS|113|7|他从灰尘里抬举贫寒的人， 从粪堆中提拔贫穷的人，
PS|113|8|使他们与贵族同坐， 与本国的贵族同坐。
PS|113|9|他使不孕的妇女安居家中， 成为快乐的母亲，儿女成群。 哈利路亚！
PS|114|1|以色列 出 埃及 ， 雅各 家离开说陌生语言之民时，
PS|114|2|犹大 作主的圣所， 以色列 为他所治理的国。
PS|114|3|沧海看见就奔逃， 约旦河 也倒流。
PS|114|4|大山踊跃如公羊， 小山跳舞如羔羊。
PS|114|5|沧海啊，你为何奔逃？ 约旦 哪，你为何倒流？
PS|114|6|大山哪，你为何踊跃如公羊？ 小山哪，你为何跳舞如羔羊？
PS|114|7|大地啊，在主的面前， 在 雅各 的上帝的面前，震动吧！
PS|114|8|他叫磐石变为水池， 使坚石变为泉源。
PS|115|1|耶和华啊，荣耀不要归与我们， 不要归与我们； 要因你的慈爱和信实归在你的名下！
PS|115|2|为何让列国说 “他们的上帝在哪里”呢？
PS|115|3|但是，我们的上帝在天上， 万事都随自己的旨意而行。
PS|115|4|他们的偶像是金的，是银的， 是人手所造的，
PS|115|5|有口却不能言， 有眼却不能看，
PS|115|6|有耳却不能听， 有鼻却不能闻，
PS|115|7|有手却不能摸， 有脚却不能走， 有喉却不能说话。
PS|115|8|造它们的要像它们一样， 凡靠它们的也必如此。
PS|115|9|以色列 啊，要倚靠耶和华！ 他是人的帮助和盾牌。
PS|115|10|亚伦 家啊，要倚靠耶和华！ 他是人的帮助和盾牌。
PS|115|11|敬畏耶和华的人哪，要倚靠耶和华！ 他是人的帮助和盾牌。
PS|115|12|耶和华向来眷念我们， 他还要赐福， 赐福给 以色列 家， 赐福给 亚伦 家。
PS|115|13|凡敬畏耶和华的，无论大小， 主必赐福给他。
PS|115|14|愿耶和华使你们 和你们的子孙日见增加。
PS|115|15|你们蒙了耶和华的福， 他是创造天地的主宰。
PS|115|16|天，是耶和华的天； 地，他却给了世人。
PS|115|17|死人不能赞美耶和华， 下到寂静 中的也都不能。
PS|115|18|但我们要称颂耶和华， 从今时直到永远。 哈利路亚！
PS|116|1|我爱耶和华， 因为他听了我的声音和我的恳求。
PS|116|2|他既向我侧耳， 我一生要求告他。
PS|116|3|死亡的绳索勒住我， 阴间的痛苦抓住我， 我遭遇患难愁苦。
PS|116|4|那时，我求告耶和华的名： “耶和华啊，求你救我！”
PS|116|5|耶和华有恩惠，有公义， 我们的上帝有怜悯。
PS|116|6|耶和华保护愚蒙的人； 我落到卑微的地步，他救了我。
PS|116|7|我的心哪！你要复归安宁， 因为耶和华用厚恩待你。
PS|116|8|主啊，你救我的命脱离死亡， 使我的眼不再流泪， 使我的脚不致跌倒。
PS|116|9|我行在耶和华面前， 走在活人之地。
PS|116|10|我信，尽管我说： “我受了极大的困苦。”
PS|116|11|我曾惊惶地说： “人都是说谎的！”
PS|116|12|耶和华向我赏赐一切厚恩， 我拿什么来报答他呢？
PS|116|13|我要举起救恩的杯， 称扬耶和华的名。
PS|116|14|我要在他的全体百姓面前 向耶和华还我所许的愿。
PS|116|15|在耶和华眼中， 圣民之死极为宝贵。
PS|116|16|耶和华啊，哦，我是你的仆人； 我是你的仆人，是你使女的儿子。 你已经解开我的捆索。
PS|116|17|我要以感谢为祭献给你， 又要求告耶和华的名。
PS|116|18|我要在 耶路撒冷 当中， 在耶和华殿的院内， 在他的全体百姓面前， 向耶和华还我所许的愿。 哈利路亚！
PS|116|19|
PS|117|1|万国啊，你们要赞美耶和华！ 万族啊，你们都要颂赞他！
PS|117|2|因为他向我们大施慈爱， 耶和华的信实存到永远。 哈利路亚！
PS|118|1|你们要称谢耶和华，因他本为善； 他的慈爱永远长存！
PS|118|2|愿 以色列 说： “他的慈爱永远长存！”
PS|118|3|愿 亚伦 家说： “他的慈爱永远长存！”
PS|118|4|愿敬畏耶和华的人说： “他的慈爱永远长存！”
PS|118|5|我在急难中求告耶和华， 耶和华就应允我，把我安置在宽阔之地。
PS|118|6|耶和华在我这边 ，我必不惧怕， 人能把我怎么样呢？
PS|118|7|在那帮助我的人中，有耶和华帮助我， 所以我要看见那些恨我的人遭报。
PS|118|8|投靠耶和华， 强似倚赖人；
PS|118|9|投靠耶和华， 强似倚赖权贵。
PS|118|10|列邦围绕我， 我靠耶和华的名必剿灭他们。
PS|118|11|他们围绕我，围困我， 我靠耶和华的名必剿灭他们。
PS|118|12|他们如同蜜蜂一般地围绕我， 他们熄灭，好像烧荆棘的火； 我靠耶和华的名，必剿灭他们。
PS|118|13|你用力推我，要叫我跌倒， 但耶和华帮助了我。
PS|118|14|耶和华是我的力量，是我的诗歌， 他也成了我的拯救。
PS|118|15|在义人的帐棚里，有欢呼拯救的声音， 耶和华的右手施展大能。
PS|118|16|耶和华的右手高举， 耶和华的右手施展大能。
PS|118|17|我不至于死，仍要存活， 并要传扬耶和华的作为。
PS|118|18|耶和华虽严严地惩治我， 却未曾将我交于死亡。
PS|118|19|给我敞开义门， 我要进去称谢耶和华！
PS|118|20|这是耶和华的门， 义人要进去！
PS|118|21|我要称谢你，因为你已经应允我， 又成了我的拯救！
PS|118|22|匠人所丢弃的石头 已成了房角的头块石头。
PS|118|23|这是耶和华所做的， 在我们眼中看为奇妙。
PS|118|24|这是耶和华所定的日子， 我们在其中要高兴欢喜！
PS|118|25|耶和华啊，求你拯救 ！ 耶和华啊，求你使我们顺利！
PS|118|26|奉耶和华的名来的是应当称颂的！ 我们从耶和华的殿中为你们祝福！
PS|118|27|耶和华是上帝， 他光照了我们。 你们要用绳索把祭牲拴住， 直牵到坛角。
PS|118|28|你是我的上帝，我要称谢你！ 我的上帝啊，我要尊崇你 ！
PS|118|29|你们要称谢耶和华，因他本为善； 他的慈爱永远长存！
PS|119|1|行为正直、遵行耶和华律法的， 这人有福了！
PS|119|2|遵守他的法度、一心寻求他的， 这人有福了！
PS|119|3|他们不做不义的事， 但遵行他的道。
PS|119|4|耶和华啊，你曾将你的训词吩咐我们， 为要我们切实遵守。
PS|119|5|但愿我行事坚定， 得以遵守你的律例。
PS|119|6|我看重你的一切命令， 就不致羞愧。
PS|119|7|我学习你公义的典章， 要以正直的心称谢你。
PS|119|8|我必遵守你的律例， 求你不要把我全然弃绝！
PS|119|9|青年要如何保持纯洁呢？ 是要遵行你的话！
PS|119|10|我曾一心寻求你， 求你不要使我偏离你的命令。
PS|119|11|我将你的话藏在心里， 免得我得罪你。
PS|119|12|耶和华啊，你是应当称颂的！ 求你将你的律例教导我！
PS|119|13|我用嘴唇传扬 你口中一切的典章。
PS|119|14|我喜爱你的法度， 如同喜爱一切的财物。
PS|119|15|我要默想你的训词， 看重你的道路。
PS|119|16|我要以你的律例为乐， 我不忘记你的话。
PS|119|17|求你用厚恩待你的仆人，使我存活， 我就遵守你的话。
PS|119|18|求你开我的眼睛， 使我看出你律法中的奇妙。
PS|119|19|我在地上是寄居的人， 求你不要向我隐藏你的命令！
PS|119|20|我时常切慕你的典章， 耗尽心力。
PS|119|21|受诅咒、偏离你命令的骄傲人， 你已经责备他们。
PS|119|22|求你除掉我所受的羞辱和藐视， 因我遵守你的法度。
PS|119|23|虽有掌权者坐着妄论我， 你仆人却思想你的律例。
PS|119|24|你的法度也是我的喜乐， 我的导师 。
PS|119|25|我的性命几乎归于尘土， 求你照你的话将我救活！
PS|119|26|我述说我所做的，你应允了我； 求你将你的律例教导我！
PS|119|27|求你使我明白你的训词， 我要默想你的奇事。
PS|119|28|我因愁苦身心耗尽， 求你照你的话使我坚立！
PS|119|29|求你使我离开奸诈的道路， 开恩将你的律法赐给我！
PS|119|30|我选择了忠信的道路， 将你的典章摆在我面前。
PS|119|31|我持守你的法度； 耶和华啊，求你不要叫我羞愧！
PS|119|32|你使我心胸开阔的时候， 我就往你命令的道路直奔。
PS|119|33|耶和华啊，求你将你的律例指教我， 我必遵守到底！
PS|119|34|求你赐我悟性，我就遵守你的律法， 且要一心遵守。
PS|119|35|求你叫我遵行你的命令， 因为这是我所喜爱的。
PS|119|36|求你使我的心趋向你的法度， 不趋向不义之财。
PS|119|37|求你叫我转眼不看虚假， 使我活在你的道路 中。
PS|119|38|求你向敬畏你的仆人 坚守你的话！
PS|119|39|求你使我所惧怕的羞辱远离我， 因你的典章本为美。
PS|119|40|看哪，我切慕你的训词， 求你因你的公义赐我生命 ！
PS|119|41|耶和华啊，求你使你的慈爱临到我， 照你的话使你的救恩临到我，
PS|119|42|我就有话回答那羞辱我的， 因我倚靠你的话。
PS|119|43|求你叫真理的话总不离开我的口， 因我仰望你的典章。
PS|119|44|我要常守你的律法， 直到永永远远。
PS|119|45|我要自由而行 ， 因我寻求了你的训词。
PS|119|46|我要在列王面前宣讲你的法度， 也不致羞愧。
PS|119|47|我以你的命令为乐， 这命令是我所喜爱的。
PS|119|48|我向我所爱的，就是你的命令高举双手 ， 我也要默想你的律例。
PS|119|49|求你记念你向仆人所说的话， 这话使我有盼望。
PS|119|50|你的话将我救活了； 这是我在患难中的安慰。
PS|119|51|骄傲的人极度地侮慢我， 我却未曾偏离你的律法。
PS|119|52|耶和华啊，我记念你从古以来的典章， 就得了安慰。
PS|119|53|我因恶人离弃你的律法， 怒火中烧。
PS|119|54|我在世寄居， 以你的律例为诗歌。
PS|119|55|耶和华啊，我夜间记念你的名， 我也要遵守你的律法。
PS|119|56|这临到我， 是因我谨守你的训词。
PS|119|57|耶和华是我的福分； 我曾说，我要遵守你的话。
PS|119|58|我一心恳求你的面， 求你照你的话怜悯我！
PS|119|59|我思想自己所行的道路， 我的脚步就转向你的法度。
PS|119|60|我速速遵守你的命令， 并不迟延。
PS|119|61|恶人的绳索缠绕我， 我却没有忘记你的律法。
PS|119|62|我因你公义的典章， 夜半起来称谢你。
PS|119|63|凡敬畏你、守你训词的人， 我都与他作伴。
PS|119|64|耶和华啊，遍地满了你的慈爱； 求你将你的律例教导我！
PS|119|65|耶和华啊，你照你的话， 善待你的仆人。
PS|119|66|求你教我明辨和知识， 因我信靠你的命令。
PS|119|67|我未受苦以先曾经迷失， 现在却遵守你的话。
PS|119|68|你本为善，所行的也善； 求你将你的律例教导我！
PS|119|69|骄傲的人编造谎言攻击我， 我却要一心遵守你的训词。
PS|119|70|他们的心蒙昧如蒙油脂， 我却喜爱你的律法。
PS|119|71|我受苦是与我有益， 为要使我学习你的律例。
PS|119|72|你口中的律法与我有益， 胜于千万金银。
PS|119|73|你的手造了我，塑造我； 求你赐我悟性学习你的命令！
PS|119|74|敬畏你的人看见我就欢喜， 因我仰望你的话。
PS|119|75|耶和华啊，我知道你的典章是公义的； 你使我受苦是以信实待我。
PS|119|76|求你照着你向仆人所说的话， 以慈爱安慰我。
PS|119|77|求你的怜悯临到我，使我存活， 因你的律法是我的喜乐。
PS|119|78|愿骄傲的人蒙羞，因为他们无理倾覆我； 但我要默想你的训词。
PS|119|79|愿敬畏你的人和知道你法度的人 都归向我。
PS|119|80|愿我的心在你的律例上完全， 使我不致蒙羞。
PS|119|81|我渴想你的救恩身心耗尽， 我仰望你的话。
PS|119|82|我因渴望你的话眼睛失明，说： “你何时安慰我呢？”
PS|119|83|我虽像烟薰的皮囊， 却不忘记你的律例。
PS|119|84|你仆人的年日有多少呢？ 你几时向迫害我的人施行审判呢？
PS|119|85|不顺从你律法的骄傲人 为我掘了坑。
PS|119|86|你的命令尽都信实； 他们无理迫害我，求你帮助我！
PS|119|87|他们几乎把我从世上除灭； 但我没有离弃你的训词。
PS|119|88|求你照你的慈爱将我救活， 我就遵守你口中的法度。
PS|119|89|耶和华啊，你的话安定在天， 直到永远。
PS|119|90|你的信实存到万代； 你坚立了地，地就长存。
PS|119|91|天地照你的典章存到今日； 万物都是你的仆役。
PS|119|92|我若不以你的律法为乐， 早就在苦难中灭绝了！
PS|119|93|我永不忘记你的训词， 因你用这训词将我救活。
PS|119|94|我是属你的，求你救我， 因我寻求了你的训词。
PS|119|95|恶人等着要灭绝我， 我却要揣摩你的法度。
PS|119|96|我看万事尽都有限， 惟有你的命令极其宽广。
PS|119|97|我何等爱慕你的律法， 终日不住地思想。
PS|119|98|你的命令常存在我心里， 使我比仇敌有智慧。
PS|119|99|我比我的教师更通达， 因我思想你的法度。
PS|119|100|我比年老的更明白， 因我谨守你的训词。
PS|119|101|我阻止我的脚走一切邪路， 为要遵守你的话。
PS|119|102|我没有偏离你的典章， 因为你教导了我。
PS|119|103|你的言语在我上膛何等甘美， 在我口中比蜜更甜！
PS|119|104|我藉着你的训词得以明白， 因此，我恨恶一切虚假的行径。
PS|119|105|你的话是我脚前的灯， 是我路上的光。
PS|119|106|你公义的典章，我曾起誓遵守， 我必按着誓言而行。
PS|119|107|我极其痛苦； 耶和华啊，求你照你的话将我救活！
PS|119|108|耶和华啊，求你悦纳我口中的赞美为甘心祭， 又将你的典章教导我！
PS|119|109|我的性命常在我手掌中 ， 我却不忘记你的律法。
PS|119|110|恶人为我设下罗网， 我却没有偏离你的训词。
PS|119|111|我以你的法度为永远的产业， 因这是我心中所喜爱的。
PS|119|112|我的心倾向你的律例， 谨守到底，直到永远。
PS|119|113|心怀二意的人为我所恨； 但你的律法为我所爱。
PS|119|114|你是我藏身之处，是我的盾牌； 我仰望你的话。
PS|119|115|作恶的人哪，你们离开我吧！ 我要遵守我上帝的命令。
PS|119|116|求你照你的话扶持我，使我存活， 不要叫我因失望而蒙羞。
PS|119|117|求你扶持我，使我得救， 时常看重你的律例。
PS|119|118|凡偏离你律例的人，你都轻看他们， 因为他们的诡诈必归虚空。
PS|119|119|你除掉地上所有的恶人，好像除掉渣滓 ； 因此我喜爱你的法度。
PS|119|120|我因惧怕你，肉体战栗； 我害怕你的典章。
PS|119|121|我行公平和公义， 求你不要撇下我，交给欺压我的人！
PS|119|122|求你保证你的仆人得福， 不容骄傲的人欺压我！
PS|119|123|我因盼望你的救恩 和你公义的言语眼睛失明。
PS|119|124|求你照你的慈爱待仆人， 将你的律例教导我。
PS|119|125|我是你的仆人，求你赐我悟性， 得以认识你的法度。
PS|119|126|这是耶和华采取行动的时候， 因人废弃了你的律法。
PS|119|127|所以，我喜爱你的命令胜于金子， 更胜于纯金。
PS|119|128|你的一切训词，在万事上我都以为正直； 我恨恶一切虚假的行径。
PS|119|129|你的法度奇妙， 所以我一心谨守。
PS|119|130|你的话一开启就发出亮光， 使愚蒙人通达。
PS|119|131|我大大张口，呼吸急促， 因我切慕你的命令。
PS|119|132|求你转向我，怜悯我， 就像你待那些喜爱你名的人。
PS|119|133|求你用你的言语使我脚步稳健， 不容罪孽辖制我。
PS|119|134|求你救我脱离人的欺压， 我要遵守你的训词。
PS|119|135|求你使你的脸向仆人发光， 又将你的律例教导我。
PS|119|136|我的眼睛流泪成河， 因为他们不守你的律法。
PS|119|137|耶和华啊，你是公义的； 你的典章正直！
PS|119|138|你所颁布的法度是公义的， 极其可靠。
PS|119|139|我的狂热把我烧灭， 因我敌人忘记你的话。
PS|119|140|你的言语极其精炼， 令你仆人喜爱。
PS|119|141|我渺小，被人藐视， 却不忘记你的训词。
PS|119|142|你的公义永远公义， 你的律法是确实的。
PS|119|143|我遭遇患难愁苦， 你的命令是我的喜乐。
PS|119|144|你的法度永远公义； 求你赐我悟性，使我存活。
PS|119|145|耶和华啊，我一心呼求你，求你应允我！ 我必谨守你的律例。
PS|119|146|我向你呼求，求你救我！ 我要遵守你的法度。
PS|119|147|天尚未亮我呼喊求救， 我仰望你的话。
PS|119|148|我终夜双眼睁开， 为要思想你的言语。
PS|119|149|求你按你的慈爱听我的声音， 耶和华啊，求你照你的典章将我救活！
PS|119|150|追逐奸恶的人 迫近了， 他们远离你的律法。
PS|119|151|耶和华啊，你就在我身边， 你一切的命令是确实的！
PS|119|152|我从你的法度早已知道， 这法度是你永远立定的。
PS|119|153|求你看顾我的苦难，搭救我， 因我不忘记你的律法。
PS|119|154|求你为我的冤屈辩护，救赎我， 照你的言语将我救活。
PS|119|155|救恩远离恶人， 因为他们不寻求你的律例。
PS|119|156|耶和华啊，你的怜悯本为大； 求你照你的典章将我救活。
PS|119|157|迫害我的、抵挡我的甚多， 我却没有偏离你的法度。
PS|119|158|我看见奸恶的人就憎恶， 因为他们不遵守你的言语。
PS|119|159|你看我何等喜爱你的训词！ 耶和华啊，求你按你的慈爱将我救活！
PS|119|160|你话语的精髓是真实的， 你一切公义的典章永远长存。
PS|119|161|掌权者无故迫害我， 然而我的心畏惧你的话。
PS|119|162|我喜爱你的言语， 好像人得到许多战利品。
PS|119|163|我恨恶，憎恶虚假； 惟喜爱你的律法。
PS|119|164|我因你公义的典章 一天七次赞美你。
PS|119|165|喜爱你律法的人大有平安， 任何事都不能使他们跌倒。
PS|119|166|耶和华啊，我仰望你的救恩， 遵行你的命令。
PS|119|167|我心谨守你的法度， 这法度我极其喜爱。
PS|119|168|我遵守你的训词和法度， 因我所行的道路都在你的面前。
PS|119|169|耶和华啊，愿我的呼求达到你面前， 求你照你的话赐我悟性。
PS|119|170|愿我的恳求达到你面前， 求你照你的言语搭救我。
PS|119|171|愿我的嘴唇发出赞美， 因为你将律例教导我。
PS|119|172|愿我的舌头歌唱你的言语， 因你一切的命令尽都公义。
PS|119|173|求你用你的手帮助我， 因我选择你的训词。
PS|119|174|耶和华啊，我切慕你的救恩！ 你的律法是我的喜乐。
PS|119|175|愿我的性命存活，得以赞美你！ 愿你的典章帮助我！
PS|119|176|我走迷了路如同失丧的羊，求你寻找你的仆人， 因我不忘记你的命令。
PS|120|1|我在急难中求告耶和华， 他就应允我。
PS|120|2|耶和华啊，求你救我脱离 说谎的嘴唇和诡诈的舌头！
PS|120|3|诡诈的舌头啊，他会给你什么呢？ 会加给你什么呢？
PS|120|4|就是勇士的利箭、 罗腾木 的炭火。
PS|120|5|祸哉！我寄居在 米设 ， 住在 基达 帐棚之中。
PS|120|6|我与那恨恶和平的人 许久同住。
PS|120|7|我愿和平， 当我发言，他们却要战争。
PS|121|1|我要向山举目， 我的帮助从何而来？
PS|121|2|我的帮助 从造天地的耶和华而来。
PS|121|3|他不叫你的脚摇动， 保护你的必不打盹！
PS|121|4|保护 以色列 的 必不打盹，也不睡觉。
PS|121|5|保护你的是耶和华， 耶和华在你右边荫庇你。
PS|121|6|白日，太阳必不伤你； 夜间，月亮也不害你。
PS|121|7|耶和华要保护你，免受一切的灾害， 他要保护你的性命。
PS|121|8|你出你入，耶和华要保护你， 从今时直到永远。
PS|122|1|我喜乐， 因人对我说：“我们到耶和华的殿去。”
PS|122|2|耶路撒冷 啊， 我们的脚站在你门内。
PS|122|3|耶路撒冷 被建造， 如同连结整齐的一座城。
PS|122|4|众支派就是耶和华的支派，上那里去， 按 以色列 的法度颂扬耶和华的名。
PS|122|5|他们在那里设立审判的宝座， 就是 大卫 家的宝座。
PS|122|6|你们要为 耶路撒冷 求平安： “愿爱你的人兴旺！
PS|122|7|愿你城中有平安！ 愿你宫内得平静！”
PS|122|8|为我弟兄和同伴的缘故，我要说： “愿你平安！”
PS|122|9|为耶和华－我们上帝殿的缘故， 我要为你求福！
PS|123|1|坐在天上的主啊， 我向你举目。
PS|123|2|看哪，仆人的眼睛怎样仰望主人的手， 婢女的眼睛怎样仰望女主人的手， 我们的眼睛也照样仰望耶和华－我们的上帝， 直到他怜悯我们。
PS|123|3|耶和华啊，求你怜悯我们，怜悯我们！ 因为我们受尽了藐视。
PS|123|4|我们受尽了安逸人的讥诮 和骄傲人的藐视。
PS|124|1|说吧， 以色列 ： “若不是耶和华帮助我们，
PS|124|2|若不是耶和华帮助我们， 当人起来攻击我们，
PS|124|3|那时，人向我们发怒， 就把我们活活吞了；
PS|124|4|那时，波涛必漫过我们， 河水必淹没我们；
PS|124|5|那时，狂傲的水 必淹没我们。”
PS|124|6|耶和华是应当称颂的！ 他没有把我们交给他们，作牙齿的猎物。
PS|124|7|我们好像雀鸟，从捕鸟人的罗网里逃脱， 罗网破裂，我们就逃脱了。
PS|124|8|我们得帮助， 是因造天地之耶和华的名。
PS|125|1|倚靠耶和华的人好像 锡安山 ， 安稳坐镇，永不动摇。
PS|125|2|众山怎样围绕 耶路撒冷 ， 耶和华也照样围绕他的百姓，从今时直到永远。
PS|125|3|恶人的杖必不在义人的土地上停留， 免得义人伸手作恶。
PS|125|4|耶和华啊，求你善待 行善和心里正直的人。
PS|125|5|至于那偏行弯曲道路的人， 耶和华必将他们和作恶的人一同驱逐出去。 愿平安归于 以色列 ！
PS|126|1|当耶和华使 锡安 被掳的人归回的时候， 我们好像做梦的人。
PS|126|2|那时，我们满口喜笑、 满舌欢呼； 那时，列国中就有人说： “耶和华为他们行了大事！”
PS|126|3|耶和华果然为我们行了大事， 我们就欢喜。
PS|126|4|耶和华啊，求你使我们这些被掳的人归回， 好像 尼革夫 的河水复流。
PS|126|5|流泪撒种的， 必欢呼收割！
PS|126|6|那带种流泪出去的， 必欢呼地带禾捆回来！
PS|127|1|若不是耶和华建造房屋， 建造的人就枉然劳力； 若不是耶和华看守城池， 看守的人就枉然警醒。
PS|127|2|你们清晨早起，夜晚安歇， 吃劳碌得来的饭，本是枉然； 惟有耶和华所亲爱的， 必叫他安然睡觉。
PS|127|3|看哪，儿女是耶和华所赐的产业， 所怀的胎是他所给的赏赐。
PS|127|4|人在年轻时生的儿女 好像勇士手中的箭。
PS|127|5|箭袋充满的人有福了！ 他们在城门口和仇敌争论时必不蒙羞。
PS|128|1|凡敬畏耶和华、 遵行他道的人有福了！
PS|128|2|你要吃劳碌得来的； 你要享福，凡事顺利。
PS|128|3|你妻子在你内室，好像多结果子的葡萄树； 你儿女围绕你的桌子，如同橄榄树苗。
PS|128|4|看哪，敬畏耶和华的人 必要这样蒙福！
PS|128|5|愿耶和华从 锡安 赐福给你！ 愿你一生一世看见 耶路撒冷 兴旺！
PS|128|6|愿你看见 你的子子孙孙！ 愿平安归于 以色列 ！
PS|129|1|说吧， 以色列 ： “从我幼年以来，人屡次苦害我；
PS|129|2|从我幼年以来，人屡次苦害我， 却没有胜过我。
PS|129|3|扶犁的人在我背上扶犁而耕， 耕的犁沟很长。”
PS|129|4|耶和华是公义的， 他砍断了恶人的绳索。
PS|129|5|愿恨恶 锡安 的 都蒙羞退后！
PS|129|6|愿他们像房顶上的草， 一发芽就枯干，
PS|129|7|收割的不够用手抓一把， 捆禾的也不够抱满怀。
PS|129|8|过路的也不说：“愿耶和华所赐的福归与你们！ 我们奉耶和华的名给你们祝福！”
PS|130|1|耶和华啊， 我从深处求告你！
PS|130|2|主啊，求你听我的声音！ 求你侧耳听我恳求的声音！
PS|130|3|耶和华啊，你若究察罪孽， 主啊，谁能站得住呢？
PS|130|4|但在你有赦免之恩， 要叫人敬畏你。
PS|130|5|我等候耶和华，我的心等候； 我也仰望他的话。
PS|130|6|我的心等候主，胜于守夜的等候天亮， 胜于守夜的等候天亮。
PS|130|7|以色列 啊，你当仰望耶和华， 因耶和华有慈爱，有丰盛的救恩。
PS|130|8|他必救赎 以色列 脱离一切的罪孽。
PS|131|1|耶和华啊，我的心不狂妄， 我的眼不高傲； 重大和测不透的事， 我也不敢行。
PS|131|2|我使我心安稳平静，好像母亲怀中断奶的孩子； 我的心在我里面如同断过奶的孩子。
PS|131|3|以色列 啊，你当仰望耶和华， 从今时直到永远！
PS|132|1|耶和华啊，求你记念 大卫 ， 记念他所受的一切苦难！
PS|132|2|他怎样向耶和华起誓， 向 雅各 的大能者许愿：
PS|132|3|“我必不进我的帐幕， 也不上我的床铺；
PS|132|4|我不容我的眼睛睡觉， 也不容我的眼皮打盹；
PS|132|5|直等到我为耶和华寻得所在， 为 雅各 的大能者寻得居所。”
PS|132|6|我们听说约柜在 以法他 ， 我们在 雅珥 的田野寻见它。
PS|132|7|“我们要进他的居所， 在他脚凳前下拜。”
PS|132|8|耶和华啊，求你兴起， 与你有能力的约柜同入安歇之所！
PS|132|9|愿你的祭司披上公义！ 愿你的圣民欢呼！
PS|132|10|求你因你仆人 大卫 的缘故， 不要厌弃你的受膏者！
PS|132|11|耶和华凭信实向 大卫 起了誓，绝不改变： “我要立你身所生的 坐在你的宝座上。
PS|132|12|你的众子若谨守我的约和我所教导他们的法度， 他们的子孙必永远坐在你的宝座上。”
PS|132|13|因为耶和华拣选了 锡安 ， 愿意当作自己的居所：
PS|132|14|“这是我永远安歇之所； 我要住在这地方，因为我愿意在这里。
PS|132|15|我要赐福使粮食丰足， 使其中的贫穷人饱享食物。
PS|132|16|我要使祭司披上救恩， 圣民就要大声欢呼！
PS|132|17|在那里我要使 大卫 的角茁壮， 为我的受膏者预备明灯。
PS|132|18|我要使他的仇敌披上羞耻； 但他的冠冕要在他头上发光。”
PS|133|1|看哪，弟兄和睦同住 是何等的善，何等的美！
PS|133|2|这好比那贵重的油浇在 亚伦 的头上， 流到胡须，又流到他的衣襟；
PS|133|3|又好比 黑门 的甘露降在 锡安山 ； 因为在那里有耶和华所命定的福，就是永远的生命。
PS|134|1|来，称颂耶和华！ 夜间侍立在耶和华殿中，耶和华的仆人，
PS|134|2|当向圣所举手， 称颂耶和华！
PS|134|3|愿造天地的耶和华 从 锡安 赐福给你们！
PS|135|1|哈利路亚！ 你们要赞美耶和华的名！ 侍立在耶和华殿中，耶和华的仆人， 侍立在我们上帝殿院中的，要赞美他！
PS|135|2|
PS|135|3|你们要赞美耶和华， 因耶和华本为善； 要歌颂他的名， 因为这是美好的。
PS|135|4|耶和华拣选 雅各 归自己， 拣选 以色列 作他宝贵的产业。
PS|135|5|我知道耶和华本为大， 也知道我们的主超乎万神之上。
PS|135|6|在天，在地，在海洋，在各深渊， 耶和华都随自己的旨意而行。
PS|135|7|他使云雾从地极上腾， 造电随雨而闪， 从仓库中吹出风来。
PS|135|8|他将 埃及 头生的， 连人带牲畜都击杀了。
PS|135|9|埃及 啊，他施行神迹奇事， 在你们中间，在法老和他所有臣仆身上。
PS|135|10|他击打许多国家， 杀戮大能的君王，
PS|135|11|就是 亚摩利 王 西宏 、 巴珊 王 噩 ， 和 迦南 一切的国度，
PS|135|12|他赏赐他们的地为业， 作为自己百姓 以色列 的产业。
PS|135|13|耶和华啊，你的名字存到永远！ 耶和华啊，你的称号 存到万代！
PS|135|14|耶和华要为自己的百姓伸冤， 为自己的仆人发怜悯。
PS|135|15|外邦的偶像是金的，是银的， 是人手所造的，
PS|135|16|有口却不能言， 有眼却不能看，
PS|135|17|有耳却不能听， 口中也没有气息。
PS|135|18|造它们的要像它们一样， 凡靠它们的也必如此。
PS|135|19|以色列 家啊，要称颂耶和华！ 亚伦 家啊，要称颂耶和华！
PS|135|20|利未 家啊，要称颂耶和华！ 你们敬畏耶和华的，要称颂耶和华！
PS|135|21|住在 耶路撒冷 的、 锡安 的耶和华， 是应当称颂的。 哈利路亚！
PS|136|1|你们要称谢耶和华，因他本为善； 他的慈爱永远长存。
PS|136|2|你们要称谢万神之神， 因他的慈爱永远长存。
PS|136|3|你们要称谢万主之主， 因他的慈爱永远长存。
PS|136|4|称谢那惟一能行大 奇事的， 因他的慈爱永远长存。
PS|136|5|称谢那用智慧造天的， 因他的慈爱永远长存。
PS|136|6|称谢那铺地在水以上的， 因他的慈爱永远长存。
PS|136|7|称谢那造成大光的， 因他的慈爱永远长存。
PS|136|8|他造太阳管白昼， 因他的慈爱永远长存。
PS|136|9|他造月亮星宿管黑夜， 因他的慈爱永远长存。
PS|136|10|称谢那击杀 埃及 凡是头生的， 因他的慈爱永远长存。
PS|136|11|他以大能的手和伸出来的膀臂， 因他的慈爱永远长存。 领 以色列 人从 埃及 人中出来， 因他的慈爱永远长存。
PS|136|12|
PS|136|13|称谢那分裂 红海 的， 因他的慈爱永远长存。
PS|136|14|他领 以色列 从其中经过， 因他的慈爱永远长存；
PS|136|15|却把法老和他的军队推落 红海 里， 因他的慈爱永远长存。
PS|136|16|称谢那引导自己子民行走旷野的， 因他的慈爱永远长存。
PS|136|17|称谢那击杀大君王的， 因他的慈爱永远长存。
PS|136|18|他杀戮威武的君王， 因他的慈爱永远长存；
PS|136|19|杀戮 亚摩利 王 西宏 ， 因他的慈爱永远长存；
PS|136|20|杀戮 巴珊 王 噩 ， 因他的慈爱永远长存。
PS|136|21|他赏赐他们的地为业， 因他的慈爱永远长存；
PS|136|22|作为他仆人 以色列 的产业， 因他的慈爱永远长存。
PS|136|23|我们身处卑微，他顾念我们， 因他的慈爱永远长存。
PS|136|24|他搭救我们脱离敌人， 因他的慈爱永远长存。
PS|136|25|凡有血有肉的，他赐粮食， 因他的慈爱永远长存。
PS|136|26|你们要称谢天上的上帝， 因他的慈爱永远长存。
PS|137|1|我们在 巴比伦 河边， 坐在那里，追想 锡安 ，就哭了。
PS|137|2|在一排柳树中， 我们挂上我们的竖琴。
PS|137|3|掳掠我们的在那里 要我们唱歌； 抢夺我们的要我们为他们作乐： “给我们唱一首 锡安 的歌吧！”
PS|137|4|我们怎能在外邦之土 唱耶和华的歌呢？
PS|137|5|耶路撒冷 啊，我若忘记你， 宁愿我的右手枯萎；
PS|137|6|我若不记得你，不看你过于我最喜乐的， 宁愿我的舌头贴于上膛！
PS|137|7|耶路撒冷 攻破的日子， 以东 人说：“拆毁！拆毁！ 直拆到根基！” 耶和华啊，求你记得！
PS|137|8|将要被灭的 巴比伦 哪， 用你待我们的恶行报复你的，那人有福了。
PS|137|9|抓起你的婴孩摔在磐石上的， 那人有福了。
PS|138|1|我要一心称谢你 ， 在诸神面前歌颂你。
PS|138|2|我要向你的圣殿下拜， 我要因你的慈爱和信实颂扬你的名； 因你使你的名和你的言语显为大， 超乎一切 。
PS|138|3|我呼求的日子，你应允我， 使我壮胆，心里有能力。
PS|138|4|耶和华啊，地上的君王都要称谢你， 因他们听见了你口中的言语。
PS|138|5|他们要歌颂耶和华的作为， 因耶和华大有荣耀。
PS|138|6|耶和华虽崇高，却看顾卑微的人； 骄傲的人，他从远处即能认出。
PS|138|7|我虽困在患难中，你必将我救活； 我的仇敌发怒，你必伸手抵挡他们， 你的右手也必拯救我。
PS|138|8|耶和华必成全他在我身上的旨意； 耶和华啊，你的慈爱永远长存！ 求你不要离弃你手所造的。
PS|139|1|耶和华啊，你已经鉴察我， 认识我。
PS|139|2|我坐下，我起来，你都晓得； 你从远处知道我的意念。
PS|139|3|我行路，我躺卧，你都细察； 你也深知我一切所行的。
PS|139|4|耶和华啊，我舌头上的话， 你没有一句不知道的。
PS|139|5|你前后环绕我， 按手在我身上。
PS|139|6|这样的知识奇妙，是我不能测的； 至高，是我不能及的。
PS|139|7|我往哪里去，躲避你的灵？ 我往哪里逃，躲避你的面？
PS|139|8|我若升到天上，你在那里； 我若躺在阴间，你也在那里。
PS|139|9|我若展开清晨的翅膀， 飞到海极居住，
PS|139|10|就是在那里，你的手必引导我， 你的右手也必扶持我。
PS|139|11|我若说“黑暗必定压碎我， 我周围的亮光必成为黑夜”，
PS|139|12|黑暗对你不再是黑暗， 黑夜却如白昼发亮。 黑暗和光明， 在你看来都是一样。
PS|139|13|我的肺腑是你所造的， 我在母腹中，你已编织 我。
PS|139|14|我要称谢你，因我受造奇妙可畏， 你的作为奇妙，这是我心深知道的。
PS|139|15|我在暗中受造，在地的深处被塑造； 那时，我的形体并不向你隐藏。
PS|139|16|我未成形的体质， 你的眼早已看见了； 你所定的日子，我尚未度一日， 都在你的册子写上了。
PS|139|17|上帝啊，你的意念向我何等宝贵！ 其数何等众多！
PS|139|18|我若数点，比海沙更多； 我睡醒的时候，仍和你同在。
PS|139|19|上帝啊，惟愿你杀戮恶人； 你们好流人血的，离开我去吧！
PS|139|20|他们说恶言顶撞你， 你的仇敌妄称你的名 。
PS|139|21|耶和华啊，恨恶你的，我岂不恨恶他们吗？ 攻击你的，我岂不憎恶他们吗？
PS|139|22|我恨恶他们到极点， 以他们为我的仇敌。
PS|139|23|上帝啊，求你鉴察我，知道我的心思， 试炼我，知道我的意念；
PS|139|24|看在我里面有什么恶行没有， 引导我走永生的道路。
PS|140|1|耶和华啊，求你救我脱离邪恶的人， 保护我脱离残暴的人！
PS|140|2|他们心中图谋奸恶， 日日不停挑起战争。
PS|140|3|他们的舌头锐利如蛇， 嘴唇里有毒蛇的毒液。（细拉）
PS|140|4|耶和华啊，求你庇护我脱离恶人的手， 保护我脱离残暴的人，他们想要推倒我。
PS|140|5|骄傲的人为我暗设罗网和绳索； 他们在路旁张开网，为我设下圈套。（细拉）
PS|140|6|我曾对耶和华说：“你是我的上帝。” 耶和华啊，求你侧耳听我恳求的声音！
PS|140|7|主－耶和华、我救恩的力量啊， 在战争的日子，你遮蔽了我的头。
PS|140|8|耶和华啊，求你不要遂恶人的心愿； 不要成就他们的计谋，免得他们自高。（细拉）
PS|140|9|至于那些昂首围困我的人， 愿他们嘴唇的奸恶陷害 自己！
PS|140|10|愿他们被丢在火中，火炭落在他们身上； 愿他们被抛在深坑里，不能再起来！
PS|140|11|愿说恶言的人在地上站立不住； 愿祸患猎取残暴的人，把他打倒。
PS|140|12|我知道耶和华必为困苦人伸冤， 为贫穷人辩护。
PS|140|13|义人必颂扬你的名， 正直人要在你面前居住。
PS|141|1|耶和华啊，我曾求告你， 求你快快临到我这里！ 我求告你的时候， 求你侧耳听我的声音！
PS|141|2|愿我的祷告如香呈到你面前！ 愿我的手举起 ，如献晚祭！
PS|141|3|耶和华啊，求你看守我的口， 把守我的嘴唇！
PS|141|4|不要使我的心偏向邪恶的事， 以致我和作恶的人一同行恶； 也不叫我吃他们的美食。
PS|141|5|任凭义人击打我，这算为仁慈； 任凭他责备我，这算为头上的膏油； 我的头不躲闪。 人正行恶的时候，我仍要祈祷。
PS|141|6|他们的审判官被扔在岩下， 他们就要听我的话，因为这话甘甜。
PS|141|7|我们的 骨头散落在阴间的口， 就像人耕田刨地 一样。
PS|141|8|主－耶和华啊，我的眼目仰望你； 我投靠你，求你不要使我的性命陷入危险！
PS|141|9|求你保护我脱离恶人为我设的罗网 和作恶之人的圈套！
PS|141|10|愿恶人落在自己的网中， 我却得以逃脱。
PS|142|1|我出声哀告耶和华， 出声恳求耶和华。
PS|142|2|我在他面前倾诉我的苦情， 在他面前陈说我的患难。
PS|142|3|我的灵在我里面发昏的时候， 你知道我的道路。 在我所行的路上， 人为我暗设罗网。
PS|142|4|求你留意向我右边观看， 无人认识我； 我无避难之处， 也无人眷顾我。
PS|142|5|耶和华啊，我曾向你哀求。 我说：“你是我的避难所， 在活人之地，你是我的福分。”
PS|142|6|求你留心听我的呼求， 因我落到极卑微之地； 求你救我脱离迫害我的人， 因为他们比我强盛。
PS|142|7|求你从被囚之地领我出来， 我好颂扬你的名。 义人必环绕我， 因为你用厚恩待我。
PS|143|1|耶和华啊，求你听我的祷告， 侧耳听我的恳求，凭你的信实和公义应允我。
PS|143|2|求你不要审问仆人， 因为在你面前，凡活着的人没有一个是义的。
PS|143|3|因为仇敌迫害我， 将我打倒在地， 使我住在幽暗之处， 像死了许久的人一样。
PS|143|4|我的灵在我里面发昏， 我的心在我里面颤栗。
PS|143|5|我追想古时之日，思想你的一切作为， 默念你手的工作。
PS|143|6|我向你举手， 我的心渴想你，如干旱之地盼雨一样。（细拉）
PS|143|7|耶和华啊，求你速速应允我！ 我的心神耗尽！ 求你不要转脸不顾我， 免得我像那些下入地府的人一样。
PS|143|8|求你使我清晨得听你慈爱的声音， 因我倚靠你； 求你使我知道当走的路， 因我的心仰望你。
PS|143|9|耶和华啊，求你救我脱离我的仇敌！ 我往你那里藏身。
PS|143|10|求你指教我遵行你的旨意， 因你是我的上帝； 愿你至善的灵 引我到平坦之地。
PS|143|11|耶和华啊，求你为你名的缘故将我救活， 凭你的公义，将我从患难中领出来，
PS|143|12|凭你的慈爱剪除我的仇敌， 灭绝所有苦待我的人，因我是你的仆人。
PS|144|1|耶和华─我的磐石是应当称颂的！ 他教导我的手争战， 教导我的指头打仗。
PS|144|2|他是我慈爱的主、我的山寨、 我的碉堡、我的救主、 我的盾牌，是我所投靠的。 他使我的百姓 服在我以下。
PS|144|3|耶和华啊，人算什么，你竟认识他！ 世人算什么，你竟顾念他！
PS|144|4|人不过像一口气， 他的年日如影消逝。
PS|144|5|耶和华啊，求你使天下垂，亲自降临； 求你摸山，使山冒烟。
PS|144|6|求你发出闪电，使仇敌四散， 射出你的箭，使他们混乱。
PS|144|7|求你从高处伸手救拔我， 救我脱离大水，脱离外邦人的手。
PS|144|8|他们的口说谎话， 他们的右手起假誓。
PS|144|9|上帝啊，我要向你唱新歌， 用十弦瑟向你歌颂。
PS|144|10|你是那拯救君王的， 你是那救仆人 大卫 脱离害命之刀的。
PS|144|11|求你救拔我， 救我脱离外邦人的手。 他们的口说谎话， 他们的右手起假誓。
PS|144|12|我们的儿子从幼年好像树苗长大， 我们的女儿如同房角石，按照建宫殿的样式凿成。
PS|144|13|我们的仓盈满，能供应各种粮食； 我们的羊在田野孳生千万。
PS|144|14|我们的牲口驮满货物， 没有人闯进来抢夺， 也没有人出去争战； 我们的街市上也没有哭号的声音。
PS|144|15|这样情况的百姓有福了！ 以耶和华为他们上帝的百姓有福了！
PS|145|1|我的上帝、我的王啊、我要尊崇你！ 我要永永远远称颂你的名！
PS|145|2|我要天天称颂你， 也要永永远远赞美你的名！
PS|145|3|耶和华本为大，该受大赞美， 其大无法测度。
PS|145|4|这一代要对那一代颂赞你的作为， 他们要传扬你的大能。
PS|145|5|他们要述说你威严荣耀的尊荣， 我要默念你奇妙的作为 。
PS|145|6|人要传讲你可畏的能力， 我也要传扬你的伟大。
PS|145|7|他们要将你可记念的大恩传开， 并要高唱你的公义。
PS|145|8|耶和华有恩惠，有怜悯， 不轻易发怒，大有慈爱。
PS|145|9|耶和华善待万有， 他的怜悯覆庇他一切所造的。
PS|145|10|耶和华啊，你一切所造的都要称谢你， 你的圣民也要称颂你。
PS|145|11|他们要传讲你国度的荣耀， 谈论你的大能，
PS|145|12|好让世人知道你大能的作为 和你国度威严的荣耀。
PS|145|13|你的国是永远的国！ 你执掌的权柄存到万代！ 耶和华一切的话信实可靠， 他一切的作为都有慈爱 。
PS|145|14|耶和华扶起所有跌倒的， 扶起所有被压下的。
PS|145|15|万有的眼目都仰望你， 你按时给他们食物。
PS|145|16|你张手， 使一切有生命的都随愿饱足。
PS|145|17|耶和华一切所行的，无不公义， 一切所做的，都有慈爱。
PS|145|18|耶和华临近凡求告他的， 临近所有诚心求告他的人。
PS|145|19|敬畏他的，他必成就他们的心愿， 也必听他们的呼求，拯救他们。
PS|145|20|耶和华保护凡爱他的人， 却要灭绝所有的恶人。
PS|145|21|我的口要述说赞美耶和华的话； 惟愿有血肉之躯的都永永远远称颂他的圣名。
PS|146|1|哈利路亚！ 我的心哪，你要赞美耶和华！
PS|146|2|我一生要赞美耶和华！ 我还活着的时候要歌颂我的上帝！
PS|146|3|你们不要倚靠君王，不要倚靠世人， 他一点也不能帮助。
PS|146|4|他的气一断，就归回尘土， 他所打算的，当日就消灭了。
PS|146|5|以 雅各 的上帝为帮助、 仰望耶和华－他上帝的，这人有福了！
PS|146|6|耶和华造天、地、海和其中的万物， 他守信实，直到永远。
PS|146|7|他为受欺压的伸冤， 赐食物给饥饿的人。 耶和华释放被囚的，
PS|146|8|耶和华开了盲人的眼睛， 耶和华扶起被压下的人， 耶和华喜爱义人。
PS|146|9|耶和华保护寄居的，扶持孤儿和寡妇， 却使恶人的道路弯曲。
PS|146|10|耶和华要作王，直到永远！ 锡安 哪，你的上帝要作王，直到万代！ 哈利路亚！
PS|147|1|哈利路亚！ 歌颂我们的上帝是美善的， 因为他是美好的，赞美他是合宜的。
PS|147|2|耶和华建造 耶路撒冷 ， 聚集 以色列 中被赶散的人。
PS|147|3|他医好伤心的人， 包扎他们的伤处。
PS|147|4|他数点星宿的数目， 一一称它们的名。
PS|147|5|我们的主本为大，大有能力， 他的智慧无法测度。
PS|147|6|耶和华扶持谦卑的人， 将恶人倾覆于地。
PS|147|7|你们要以感谢向耶和华歌唱， 用琴向我们的上帝歌颂。
PS|147|8|他用密云遮天，为地预备雨水， 使草生长在山上。
PS|147|9|他赐食物给走兽 和啼叫的小乌鸦。
PS|147|10|他不喜悦马的力大， 不喜爱人的腿快。
PS|147|11|耶和华喜爱敬畏他 和盼望他慈爱的人。
PS|147|12|耶路撒冷 啊，要颂赞耶和华！ 锡安 哪，要赞美你的上帝！
PS|147|13|因为他坚固了你的门闩， 赐福给你中间的儿女。
PS|147|14|他使你境内平安， 用上好的麦子使你满足。
PS|147|15|他向大地发出命令， 他的话速速颁行。
PS|147|16|他降雪如羊毛， 撒霜如灰烬。
PS|147|17|他掷下冰雹如碎渣， 他发出寒冷，谁能当得起呢？
PS|147|18|他一出令，这些就都融化， 他使风刮起，水便流动。
PS|147|19|他将他的道指示 雅各 ， 将他的律例典章指示 以色列 。
PS|147|20|他未曾这样对待别国， 至于他的典章，他们向来都不知道 。 哈利路亚！
PS|148|1|哈利路亚！ 你们要从天上赞美耶和华， 在高处赞美他！
PS|148|2|他的众使者啊，要赞美他！ 他的诸军啊，都要赞美他！
PS|148|3|太阳月亮啊，要赞美他！ 放光的星宿啊，都要赞美他！
PS|148|4|天上的天和天上的水啊， 你们都要赞美他！
PS|148|5|愿这些都赞美耶和华的名！ 因他一吩咐就都造成。
PS|148|6|他将这些设定，直到永永远远； 他订了律例，不能废去。
PS|148|7|你们哪，都当赞美耶和华： 地上一切所有的，大鱼和深洋，
PS|148|8|火和冰雹，雪和雾气， 成就他命令的狂风，
PS|148|9|大山和小山， 结果子的树木和一切香柏树，
PS|148|10|野兽和一切牲畜， 昆虫和飞鸟，
PS|148|11|世上的君王和万民， 领袖和世上所有的审判官，
PS|148|12|少年和少女， 老人和孩童，
PS|148|13|愿这些都赞美耶和华的名！ 因为独有他的名被尊崇，他的荣耀在天地之上。
PS|148|14|他高举自己百姓的角， 使他的圣民 以色列 人，就是与他相近的百姓得荣耀 。 哈利路亚！
PS|149|1|哈利路亚！ 你们要向耶和华唱新歌， 在圣民的会中赞美他！
PS|149|2|愿 以色列 因造他的主欢喜！ 愿 锡安 的民因他们的王快乐！
PS|149|3|愿他们跳舞赞美他的名， 击鼓弹琴歌颂他！
PS|149|4|因为耶和华喜爱自己的百姓， 他要用救恩当作谦卑人的妆饰。
PS|149|5|愿圣民因所得的荣耀欢乐！ 愿他们在床上也欢呼！
PS|149|6|愿他们口中称颂上帝为至高， 手里有两刃的剑，
PS|149|7|为要报复列国， 惩罚万民。
PS|149|8|要用链子捆他们的君王， 用铁镣锁他们的贵族，
PS|149|9|要在他们身上施行所记录的审判。 他的圣民都享荣耀。 哈利路亚！
PS|150|1|哈利路亚！ 你们要在上帝的圣所赞美他！ 在他显能力的穹苍赞美他！
PS|150|2|要因他大能的作为赞美他， 因他极其伟大赞美他！
PS|150|3|要用角声赞美他， 鼓瑟弹琴赞美他！
PS|150|4|击鼓跳舞赞美他！ 用丝弦的乐器和箫的声音赞美他！
PS|150|5|用大响的钹赞美他！ 用高声的钹赞美他！
PS|150|6|凡有生命的都要赞美耶和华！ 哈利路亚！
