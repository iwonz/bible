GAL|1|1|我使徒 保罗 和所有跟我一起的弟兄，写信给 加拉太 的众教会。我作使徒不是由于人，也不是藉着人，而是藉着耶稣基督与使他从死人中复活的父上帝。
GAL|1|2|
GAL|1|3|愿恩惠、平安 从我们的父上帝和主耶稣基督归给你们！
GAL|1|4|基督照我们父上帝的旨意，为我们的罪舍己，要救我们脱离现今这罪恶的世代。
GAL|1|5|愿荣耀归给上帝，直到永永远远。阿们！
GAL|1|6|我很惊讶你们这么快就离开那位藉着基督之 恩呼召你们的上帝，而去随从别的福音；
GAL|1|7|其实并没有另一个福音，不过有些人骚扰你们，要把基督的福音更改了。
GAL|1|8|但无论是我们或是天上来的使者，若传福音给你们 ，与我们所传给你们的不同，他该受诅咒！
GAL|1|9|我们已经说了，现在我再说，若有人传福音给你们，与你们以往所领受的不同，他该受诅咒！
GAL|1|10|我现在是要得人的心，还是要得上帝的心呢？难道我在讨人的喜欢吗？我若仍旧想讨人的喜欢，我就不是基督的仆人了。
GAL|1|11|弟兄们，我要你们知道，我所传的福音不是按照人的意思；
GAL|1|12|因为我不是从人领受的，也不是人教导我的，而是藉着耶稣基督的启示而来。
GAL|1|13|你们听说过从前我在 犹太 教中的行径，我怎样竭力压迫残害上帝的教会。
GAL|1|14|在 犹太 教中，我比本国许多同辈的人更激进，为我祖宗的传统更热心。
GAL|1|15|然而，那位把我从母腹里分别出来、又施恩呼召我的上帝 ，既然乐意
GAL|1|16|把他儿子启示在我心里，让我在外邦人中传扬他，我就没有跟有血有肉的人商量，
GAL|1|17|也没有上 耶路撒冷 去见那些比我先作使徒的，惟独到 阿拉伯 去，后来又回到 大马士革 。
GAL|1|18|过了三年，我才上 耶路撒冷 去见 矶法 ，和他同住了十五天。
GAL|1|19|至于别的使徒，除了主的兄弟 雅各 ，我都没有见过。
GAL|1|20|我现在写给你们的是在上帝面前说的，不说谎话。
GAL|1|21|以后我到了 叙利亚 和 基利家 一带；
GAL|1|22|那时，在基督里的 犹太 各教会都没有见过我的面。
GAL|1|23|不过他们听说“那从前压迫我们的，现在竟传扬他原先所残害的信仰”。
GAL|1|24|他们就为我的缘故归荣耀给上帝。
GAL|2|1|过了十四年，我再上 耶路撒冷 去， 巴拿巴 同行，也带了 提多 一起去。
GAL|2|2|我是奉了启示上去的；我把在外邦人中所传的福音对弟兄们说明，我是私下对那些有名望的人说的，免得我现在或是从前都徒然奔跑了。
GAL|2|3|但跟我同去的 提多 ，虽是 希腊 人，也没有勉强他受割礼；
GAL|2|4|因为有偷着混进来的假弟兄，暗中窥探我们在基督耶稣里拥有的自由，要使我们作奴隶，
GAL|2|5|可是，为要使福音的真理仍存在你们中间，我们一点也没有让步顺服他们。
GAL|2|6|至于那些有名望的，不论他们是何等人，都与我无关；上帝不以外貌取人。那些有名望的，并没有加增我什么。
GAL|2|7|相反地，他们看见了主托付我传福音给未受割礼的人，正如主托付 彼得 传福音给受割礼的人；
GAL|2|8|那感动 彼得 、叫他为受割礼的人作使徒的，也感动我，叫我为外邦人作使徒。
GAL|2|9|那些被认为是教会柱石的 雅各 、 矶法 、 约翰 知道上帝所赐给我的恩典，就跟我和 巴拿巴 握右手以示合作，同意我们往外邦人那里去，他们往受割礼的人那里去。
GAL|2|10|他们只要求我们记念穷人，这也是我一向热心在做的。
GAL|2|11|后来， 矶法 到了 安提阿 ，因为他有可责之处，我就当面反对他。
GAL|2|12|从 雅各 那里来的人未到以前，他和外邦人一同吃饭，及至他们来到，他因怕奉割礼的人就退出，跟外邦人疏远了。
GAL|2|13|其余的 犹太 人也都随着他装假，甚至连 巴拿巴 也随伙装假。
GAL|2|14|但我一看见他们做得不对，与福音的真理不合，就在众人面前对 矶法 说：“你既是 犹太 人，却按照外邦人的样子，不按照 犹太 人的样子生活，怎么能勉强外邦人按照 犹太 人的样子生活呢？”
GAL|2|15|我们生来就是 犹太 人，不是外邦罪人；
GAL|2|16|可是我们知道，人称义不是因律法的行为，而是因信耶稣基督 ，我们也信了基督耶稣，为要使我们因信基督称义，不因律法的行为称义，因为，凡血肉之躯没有一个能因律法的行为称义。
GAL|2|17|我们若求在基督里称义，自己却还被视为罪人，那么，基督是罪的用人吗？绝对不是！
GAL|2|18|如果我重新建造我所拆毁的，这就证明自己是违犯律法的人。
GAL|2|19|我因律法而向律法死了，使我可以向上帝活着。我已经与基督同钉十字架，
GAL|2|20|现在活着的不再是我，乃是基督在我里面活着；并且我如今在肉身活着，是因信上帝的儿子而活；他是爱我，为我舍己。
GAL|2|21|我不废掉上帝的恩；如果义是藉着律法而获得，那么基督就白白死了。
GAL|3|1|无知的 加拉太 人哪，耶稣基督钉十字架，已经活现在你们眼前，谁又迷惑了你们呢？
GAL|3|2|这是我惟一要问你们的：你们领受了圣灵，是因律法的行为或是因听信福音呢？
GAL|3|3|你们既然以圣灵开始，如今竟要以肉身终结吗？你们是这样的无知吗？
GAL|3|4|你们受这么多的苦都是徒然的吗？如果真是徒然的，
GAL|3|5|那么，上帝赐给你们圣灵，又在你们中间行异能，是因律法的行为或是因听信福音呢？
GAL|3|6|正如 亚伯拉罕 “信了上帝，这就算他为义”。
GAL|3|7|所以，你们知道：有信心的人才是 亚伯拉罕 的子孙。
GAL|3|8|圣经既然预先看见上帝要使外邦人因信称义，预先传福音给 亚伯拉罕 ，说：“万国都必因你得福。”
GAL|3|9|可见，那有信心的人和有信心的 亚伯拉罕 一同得福。
GAL|3|10|凡出于律法的行为都是受诅咒的，因为经上记着：“凡不持守律法书上所记的一切而去行的，都是受诅咒的。”
GAL|3|11|没有一个人靠着律法在上帝面前称义，这是明显的，因为经上说：“义人必因信得生。”
GAL|3|12|律法并不出于信，而是说：“行这些事的就必因此得生。”
GAL|3|13|既然基督为我们成了诅咒，就把我们从律法的诅咒中赎出来。因为经上记着：“凡挂在木头上的都是受诅咒的。”
GAL|3|14|这是要使 亚伯拉罕 的福，因着基督耶稣临到外邦人，使我们能因信得着所应许的圣灵。
GAL|3|15|弟兄们，我照着人的观点说，人的遗嘱一经确定，没有人能废弃或加增。
GAL|3|16|那些应许原是向 亚伯拉罕 和他后裔说的，并不是说“和众后裔”，指许多人，而是说“和你那个后裔”，指一个人，就是基督。
GAL|3|17|我是这么说，上帝预先所立的约不能被四百三十年以后的律法废掉，使应许失效。
GAL|3|18|因为承受产业若是出于律法，就不再是出于应许；但上帝是凭着应许把产业赐给 亚伯拉罕 。
GAL|3|19|这样说来，为什么要有律法呢？律法是为过犯的缘故而加上去的，等候那蒙应许的子孙来到才结束，是藉着天使经中保之手而设立的。
GAL|3|20|但中保本不是为单方设立的；上帝却是一位。
GAL|3|21|这样，律法是与上帝的 应许对立吗？绝对不是！如果律法的颁布能使人得生命，义就诚然出于律法了。
GAL|3|22|但圣经把万物都圈在罪里，为要使因信耶稣基督 而来的应许归给信的人。
GAL|3|23|但这“信”还未来以前，我们被看守在律法之下，像被圈住，直到那将来的“信”显明出来。
GAL|3|24|这样，律法是我们的启蒙教师，直到基督来了 ，好使我们因信称义。
GAL|3|25|但这“信”既然来到，我们从此就不在启蒙教师的手下了。
GAL|3|26|其实，你们藉着信，在基督耶稣里都成为上帝的儿女。
GAL|3|27|你们凡受洗归入基督的都披戴基督了：
GAL|3|28|不再分 犹太 人或 希腊 人，不再分为奴的自主的，不再分男的女的，因为你们在基督耶稣里都成为一了。
GAL|3|29|既然你们属于基督，你们就是 亚伯拉罕 的子孙，是照着应许承受产业的了。
GAL|4|1|我说，虽然那承受产业的是整个产业的主人，但在未成年的时候却与奴隶毫无分别，
GAL|4|2|仍是在监护人和管家的手下，直等他父亲预定的时候来到。
GAL|4|3|我们也是一样，在未成年的时候，被世上粗浅的学说 所奴役，也是如此。
GAL|4|4|等到时候成熟，上帝就差遣他的儿子，为女子所生，且生在律法之下，
GAL|4|5|为要把律法之下的人赎出来，使我们获得儿子的名分。
GAL|4|6|因为你们是儿子，上帝就差他儿子的灵进入我们 的心，呼叫：“阿爸，父！”
GAL|4|7|可见，你不再是奴隶，而是儿子了，既然是儿子，就靠着上帝也成为后嗣了。
GAL|4|8|但从前不认识上帝的时候，你们是给那些本来不是上帝的神明作奴隶；
GAL|4|9|现在你们既然认识上帝，更可说是被上帝所认识的，怎么还要转回那懦弱无用的粗浅学说 ，情愿再给它们作奴隶呢？
GAL|4|10|你们竟又谨守日子、月份、节期、年份，
GAL|4|11|我为你们担心，惟恐我在你们身上是枉费工夫了。
GAL|4|12|弟兄们，我劝你们，要像我一样，因为我也像你们一样。你们一点没有亏负我。
GAL|4|13|你们知道，我因为身体有疾病才有第一次传福音给你们的机会。
GAL|4|14|虽然你们为我身体的缘故受试炼，却没有轻看我，也没有厌弃我，反倒接待我如同上帝的使者，如同基督耶稣。
GAL|4|15|你们当日的好意哪里去了呢？那时若办得到，你们就是把自己的眼睛挖出来给我，也都情愿。这是我可以给你们作证的。
GAL|4|16|如今我把真理告诉你们，倒成了你们的仇敌吗？
GAL|4|17|那些热心待你们的人，不怀好意，是要隔绝你们，好使你们热心待他们。
GAL|4|18|在善事上，时刻热心待别人原是好的，却不只是我与你们同在的时候才这样。
GAL|4|19|我的孩子们哪，我为你们再受生产之苦，直等到基督成形在你们心里 。
GAL|4|20|我期望现今就在你们那里，可以改变我的口气，因为我为你们心里难过。
GAL|4|21|你们这愿意在律法之下的人，请告诉我，你们没有听见律法吗？
GAL|4|22|因为律法上记着， 亚伯拉罕 有两个儿子，一个是使女生的，一个是自由的妇人生的。
GAL|4|23|那使女所生的是按着肉体生的；那自由的妇人所生的是凭着应许生的。
GAL|4|24|这是比方：那两个妇人就是两个约；一个妇人是出于 西奈山 ，生子为奴，就是 夏甲 。
GAL|4|25|这 夏甲 是指着 阿拉伯 的 西奈山 ，与现在的 耶路撒冷 同类，因为 耶路撒冷 和她的儿女都是为奴的。
GAL|4|26|但另一妇人就是在上的 耶路撒冷 ，是自由的，她是我们的母亲。
GAL|4|27|因为经上记着： 不怀孕、不生养的，你要欢乐； 未曾经过产难的，你要高声欢呼； 因为没有丈夫的，比有丈夫的有更多的儿女。
GAL|4|28|弟兄们，你们是凭着应许作儿女的，如同 以撒 一样。
GAL|4|29|当时，那按着肉体生的迫害了那按着圣灵生的，现在也是这样。
GAL|4|30|然而经上是怎么说的呢？是说：“把使女和她儿子赶出去！因为使女的儿子绝不能与自由妇人的儿子一同承受产业。”
GAL|4|31|弟兄们，这样看来，我们不是使女的儿女，而是自由妇人的儿女了。
GAL|5|1|基督释放了我们，为使我们得自由。所以要站稳了，不要再被奴隶的轭挟制。
GAL|5|2|我— 保罗 告诉你们，你们若受割礼，基督就对你们无益了。
GAL|5|3|我再指着凡受割礼的人确实地说，他有义务遵行全部的律法。
GAL|5|4|你们这要靠律法称义的是与基督隔绝，从恩典中坠落了。
GAL|5|5|至于我们，我们是靠着圣灵，凭着信心，等候所盼望的义。
GAL|5|6|因为在基督耶稣里，受割礼不受割礼都没有功效，惟独使人发出仁爱的信心才有功效。
GAL|5|7|你们向来跑得好，谁拦阻了你们，使你们不顺从真理呢？
GAL|5|8|这样的劝导不是出于那召你们的。
GAL|5|9|一点面酵能使全团都发起来。
GAL|5|10|我在主里深信你们必不怀别样的心；但骚扰你们的，无论是谁，必须承受惩罚。
GAL|5|11|弟兄们，我若仍旧传割礼，为什么还受迫害呢？若是这样，十字架绊倒人的地方就没有了。
GAL|5|12|恨不得那骚扰你们的人把自己阉割了。
GAL|5|13|弟兄们，你们蒙召是要得自由；只是不可把这自由当作放纵情欲的机会，总要用爱心互相服侍。
GAL|5|14|因为全部律法都包括在“爱邻 如己”这一句话之内了。
GAL|5|15|你们要谨慎，你们若相咬相吞，恐怕要彼此消灭了。
GAL|5|16|我说，你们要顺着圣灵而行，绝不可满足肉体的情欲。
GAL|5|17|因为肉体的情欲和圣灵相争，圣灵和肉体相争，这两个彼此敌对，使你们不能做所愿意做的。
GAL|5|18|但你们若被圣灵引导，就不在律法之下。
GAL|5|19|情欲的事都是显而易见的；就如淫乱、污秽、放荡、
GAL|5|20|拜偶像、行邪术、仇恨、纷争、忌恨、愤怒、自私、分派、结党、
GAL|5|21|嫉妒 、醉酒、荒宴等类。我从前告诉过你们，现在又告诉你们，做这样事的人必不能承受上帝的国。
GAL|5|22|圣灵的果子就是仁爱、喜乐、和平、忍耐、恩慈、良善、信实、
GAL|5|23|温柔、节制。这样的事没有律法禁止。
GAL|5|24|凡属基督耶稣 的人，是已经把肉体与肉体的邪情私欲同钉在十字架上了。
GAL|5|25|我们若靠着圣灵而活，也要靠着圣灵行事。
GAL|5|26|不要贪图虚名，彼此惹气，互相嫉妒。
GAL|6|1|弟兄们，若有人偶然被过犯所胜，你们属灵的人就要用温柔的心把他挽回过来；自己也要留意，免得也被引诱。
GAL|6|2|你们各人的重担要互相担当，这样就会成全 基督的律法。
GAL|6|3|人若没有什么了不起，还自以为了不起的，就是自欺。
GAL|6|4|各人要省察自己的行为；这样，他所夸口的只在自己，而不在别人。
GAL|6|5|因为人人必须担当自己的担子。
GAL|6|6|在真道上受教的，要把一切美好的东西与施教的人分享。
GAL|6|7|不要自欺；上帝是轻慢不得的，因为人种的是什么，收的也是什么。
GAL|6|8|顺着肉体撒种的，必从肉体收败坏；顺着圣灵撒种的，必从圣灵收永生。
GAL|6|9|我们行善不可丧志，因为若不灰心，到了适当的时候就有收成。
GAL|6|10|所以，一有机会就要向众人行善，向信徒一家的人更要这样。
GAL|6|11|你们看我亲手写给你们的字是何等的大！
GAL|6|12|那些想要炫耀外表的人才勉强你们受割礼，无非是怕自己为基督的十字架受迫害。
GAL|6|13|他们那些受割礼的，连自己也不守律法；他们要你们受割礼，不过是要拿你们的肉体夸口。
GAL|6|14|但我绝不以别的夸口，只夸我们主耶稣基督的十字架；因这十字架 ，就我而论，世界已经钉在十字架上；就世界而论，我已经钉在十字架上。
GAL|6|15|受割礼或不受割礼都无关紧要，要紧的就是作新造的人。
GAL|6|16|凡照这准则行的人，愿平安 怜悯，加给他们，和上帝的 以色列 民。
GAL|6|17|从今以后，不要有人再搅扰我，因为我身上带着耶稣的印记。
GAL|6|18|弟兄们，愿我们主耶稣基督的恩与你们的灵同在。阿们！
