LAM|1|1|How deserted lies the city, once so full of people! How like a widow is she, who once was great among the nations! She who was queen among the provinces has now become a slave.
LAM|1|2|Bitterly she weeps at night, tears are upon her cheeks. Among all her lovers there is none to comfort her. All her friends have betrayed her; they have become her enemies.
LAM|1|3|After affliction and harsh labor, Judah has gone into exile. She dwells among the nations; she finds no resting place. All who pursue her have overtaken her in the midst of her distress.
LAM|1|4|The roads to Zion mourn, for no one comes to her appointed feasts. All her gateways are desolate, her priests groan, her maidens grieve, and she is in bitter anguish.
LAM|1|5|Her foes have become her masters; her enemies are at ease. The LORD has brought her grief because of her many sins. Her children have gone into exile, captive before the foe.
LAM|1|6|All the splendor has departed from the Daughter of Zion. Her princes are like deer that find no pasture; in weakness they have fled before the pursuer.
LAM|1|7|In the days of her affliction and wandering Jerusalem remembers all the treasures that were hers in days of old. When her people fell into enemy hands, there was no one to help her. Her enemies looked at her and laughed at her destruction.
LAM|1|8|Jerusalem has sinned greatly and so has become unclean. All who honored her despise her, for they have seen her nakedness; she herself groans and turns away.
LAM|1|9|Her filthiness clung to her skirts; she did not consider her future. Her fall was astounding; there was none to comfort her. "Look, O LORD, on my affliction, for the enemy has triumphed."
LAM|1|10|The enemy laid hands on all her treasures; she saw pagan nations enter her sanctuary- those you had forbidden to enter your assembly.
LAM|1|11|All her people groan as they search for bread; they barter their treasures for food to keep themselves alive. "Look, O LORD, and consider, for I am despised."
LAM|1|12|"Is it nothing to you, all you who pass by? Look around and see. Is any suffering like my suffering that was inflicted on me, that the LORD brought on me in the day of his fierce anger?
LAM|1|13|"From on high he sent fire, sent it down into my bones. He spread a net for my feet and turned me back. He made me desolate, faint all the day long.
LAM|1|14|"My sins have been bound into a yoke; by his hands they were woven together. They have come upon my neck and the Lord has sapped my strength. He has handed me over to those I cannot withstand.
LAM|1|15|"The Lord has rejected all the warriors in my midst; he has summoned an army against me to crush my young men. In his winepress the Lord has trampled the Virgin Daughter of Judah.
LAM|1|16|"This is why I weep and my eyes overflow with tears. No one is near to comfort me, no one to restore my spirit. My children are destitute because the enemy has prevailed."
LAM|1|17|Zion stretches out her hands, but there is no one to comfort her. The LORD has decreed for Jacob that his neighbors become his foes; Jerusalem has become an unclean thing among them.
LAM|1|18|"The LORD is righteous, yet I rebelled against his command. Listen, all you peoples; look upon my suffering. My young men and maidens have gone into exile.
LAM|1|19|"I called to my allies but they betrayed me. My priests and my elders perished in the city while they searched for food to keep themselves alive.
LAM|1|20|"See, O LORD, how distressed I am! I am in torment within, and in my heart I am disturbed, for I have been most rebellious. Outside, the sword bereaves; inside, there is only death.
LAM|1|21|"People have heard my groaning, but there is no one to comfort me. All my enemies have heard of my distress; they rejoice at what you have done. May you bring the day you have announced so they may become like me.
LAM|1|22|"Let all their wickedness come before you; deal with them as you have dealt with me because of all my sins. My groans are many and my heart is faint."
LAM|2|1|How the Lord has covered the Daughter of Zion with the cloud of his anger! He has hurled down the splendor of Israel from heaven to earth; he has not remembered his footstool in the day of his anger.
LAM|2|2|Without pity the Lord has swallowed up all the dwellings of Jacob; in his wrath he has torn down the strongholds of the Daughter of Judah. He has brought her kingdom and its princes down to the ground in dishonor.
LAM|2|3|In fierce anger he has cut off every horn of Israel. He has withdrawn his right hand at the approach of the enemy. He has burned in Jacob like a flaming fire that consumes everything around it.
LAM|2|4|Like an enemy he has strung his bow; his right hand is ready. Like a foe he has slain all who were pleasing to the eye; he has poured out his wrath like fire on the tent of the Daughter of Zion.
LAM|2|5|The Lord is like an enemy; he has swallowed up Israel. He has swallowed up all her palaces and destroyed her strongholds. He has multiplied mourning and lamentation for the Daughter of Judah.
LAM|2|6|He has laid waste his dwelling like a garden; he has destroyed his place of meeting. The LORD has made Zion forget her appointed feasts and her Sabbaths; in his fierce anger he has spurned both king and priest.
LAM|2|7|The Lord has rejected his altar and abandoned his sanctuary. He has handed over to the enemy the walls of her palaces; they have raised a shout in the house of the LORD as on the day of an appointed feast.
LAM|2|8|The LORD determined to tear down the wall around the Daughter of Zion. He stretched out a measuring line and did not withhold his hand from destroying. He made ramparts and walls lament; together they wasted away.
LAM|2|9|Her gates have sunk into the ground; their bars he has broken and destroyed. Her king and her princes are exiled among the nations, the law is no more, and her prophets no longer find visions from the LORD.
LAM|2|10|The elders of the Daughter of Zion sit on the ground in silence; they have sprinkled dust on their heads and put on sackcloth. The young women of Jerusalem have bowed their heads to the ground.
LAM|2|11|My eyes fail from weeping, I am in torment within, my heart is poured out on the ground because my people are destroyed, because children and infants faint in the streets of the city.
LAM|2|12|They say to their mothers, "Where is bread and wine?" as they faint like wounded men in the streets of the city, as their lives ebb away in their mothers' arms.
LAM|2|13|What can I say for you? With what can I compare you, O Daughter of Jerusalem? To what can I liken you, that I may comfort you, O Virgin Daughter of Zion? Your wound is as deep as the sea. Who can heal you?
LAM|2|14|The visions of your prophets were false and worthless; they did not expose your sin to ward off your captivity. The oracles they gave you were false and misleading.
LAM|2|15|All who pass your way clap their hands at you; they scoff and shake their heads at the Daughter of Jerusalem: "Is this the city that was called the perfection of beauty, the joy of the whole earth?"
LAM|2|16|All your enemies open their mouths wide against you; they scoff and gnash their teeth and say, "We have swallowed her up. This is the day we have waited for; we have lived to see it."
LAM|2|17|The LORD has done what he planned; he has fulfilled his word, which he decreed long ago. He has overthrown you without pity, he has let the enemy gloat over you, he has exalted the horn of your foes.
LAM|2|18|The hearts of the people cry out to the Lord. O wall of the Daughter of Zion, let your tears flow like a river day and night; give yourself no relief, your eyes no rest.
LAM|2|19|Arise, cry out in the night, as the watches of the night begin; pour out your heart like water in the presence of the Lord. Lift up your hands to him for the lives of your children, who faint from hunger at the head of every street.
LAM|2|20|"Look, O LORD, and consider: Whom have you ever treated like this? Should women eat their offspring, the children they have cared for? Should priest and prophet be killed in the sanctuary of the Lord?
LAM|2|21|"Young and old lie together in the dust of the streets; my young men and maidens have fallen by the sword. You have slain them in the day of your anger; you have slaughtered them without pity.
LAM|2|22|"As you summon to a feast day, so you summoned against me terrors on every side. In the day of the LORD's anger no one escaped or survived; those I cared for and reared, my enemy has destroyed."
LAM|3|1|I am the man who has seen affliction by the rod of his wrath.
LAM|3|2|He has driven me away and made me walk in darkness rather than light;
LAM|3|3|indeed, he has turned his hand against me again and again, all day long.
LAM|3|4|He has made my skin and my flesh grow old and has broken my bones.
LAM|3|5|He has besieged me and surrounded me with bitterness and hardship.
LAM|3|6|He has made me dwell in darkness like those long dead.
LAM|3|7|He has walled me in so I cannot escape; he has weighed me down with chains.
LAM|3|8|Even when I call out or cry for help, he shuts out my prayer.
LAM|3|9|He has barred my way with blocks of stone; he has made my paths crooked.
LAM|3|10|Like a bear lying in wait, like a lion in hiding,
LAM|3|11|he dragged me from the path and mangled me and left me without help.
LAM|3|12|He drew his bow and made me the target for his arrows.
LAM|3|13|He pierced my heart with arrows from his quiver.
LAM|3|14|I became the laughingstock of all my people; they mock me in song all day long.
LAM|3|15|He has filled me with bitter herbs and sated me with gall.
LAM|3|16|He has broken my teeth with gravel; he has trampled me in the dust.
LAM|3|17|I have been deprived of peace; I have forgotten what prosperity is.
LAM|3|18|So I say, "My splendor is gone and all that I had hoped from the LORD."
LAM|3|19|I remember my affliction and my wandering, the bitterness and the gall.
LAM|3|20|I well remember them, and my soul is downcast within me.
LAM|3|21|Yet this I call to mind and therefore I have hope:
LAM|3|22|Because of the LORD's great love we are not consumed, for his compassions never fail.
LAM|3|23|They are new every morning; great is your faithfulness.
LAM|3|24|I say to myself, "The LORD is my portion; therefore I will wait for him."
LAM|3|25|The LORD is good to those whose hope is in him, to the one who seeks him;
LAM|3|26|it is good to wait quietly for the salvation of the LORD.
LAM|3|27|It is good for a man to bear the yoke while he is young.
LAM|3|28|Let him sit alone in silence, for the LORD has laid it on him.
LAM|3|29|Let him bury his face in the dust- there may yet be hope.
LAM|3|30|Let him offer his cheek to one who would strike him, and let him be filled with disgrace.
LAM|3|31|For men are not cast off by the Lord forever.
LAM|3|32|Though he brings grief, he will show compassion, so great is his unfailing love.
LAM|3|33|For he does not willingly bring affliction or grief to the children of men.
LAM|3|34|To crush underfoot all prisoners in the land,
LAM|3|35|to deny a man his rights before the Most High,
LAM|3|36|to deprive a man of justice- would not the Lord see such things?
LAM|3|37|Who can speak and have it happen if the Lord has not decreed it?
LAM|3|38|Is it not from the mouth of the Most High that both calamities and good things come?
LAM|3|39|Why should any living man complain when punished for his sins?
LAM|3|40|Let us examine our ways and test them, and let us return to the LORD.
LAM|3|41|Let us lift up our hearts and our hands to God in heaven, and say:
LAM|3|42|"We have sinned and rebelled and you have not forgiven.
LAM|3|43|"You have covered yourself with anger and pursued us; you have slain without pity.
LAM|3|44|You have covered yourself with a cloud so that no prayer can get through.
LAM|3|45|You have made us scum and refuse among the nations.
LAM|3|46|"All our enemies have opened their mouths wide against us.
LAM|3|47|We have suffered terror and pitfalls, ruin and destruction."
LAM|3|48|Streams of tears flow from my eyes because my people are destroyed.
LAM|3|49|My eyes will flow unceasingly, without relief,
LAM|3|50|until the LORD looks down from heaven and sees.
LAM|3|51|What I see brings grief to my soul because of all the women of my city.
LAM|3|52|Those who were my enemies without cause hunted me like a bird.
LAM|3|53|They tried to end my life in a pit and threw stones at me;
LAM|3|54|the waters closed over my head, and I thought I was about to be cut off.
LAM|3|55|I called on your name, O LORD, from the depths of the pit.
LAM|3|56|You heard my plea: "Do not close your ears to my cry for relief."
LAM|3|57|You came near when I called you, and you said, "Do not fear."
LAM|3|58|O Lord, you took up my case; you redeemed my life.
LAM|3|59|You have seen, O LORD, the wrong done to me. Uphold my cause!
LAM|3|60|You have seen the depth of their vengeance, all their plots against me.
LAM|3|61|O LORD, you have heard their insults, all their plots against me-
LAM|3|62|what my enemies whisper and mutter against me all day long.
LAM|3|63|Look at them! Sitting or standing, they mock me in their songs.
LAM|3|64|Pay them back what they deserve, O LORD, for what their hands have done.
LAM|3|65|Put a veil over their hearts, and may your curse be on them!
LAM|3|66|Pursue them in anger and destroy them from under the heavens of the LORD.
LAM|4|1|How the gold has lost its luster, the fine gold become dull! The sacred gems are scattered at the head of every street.
LAM|4|2|How the precious sons of Zion, once worth their weight in gold, are now considered as pots of clay, the work of a potter's hands!
LAM|4|3|Even jackals offer their breasts to nurse their young, but my people have become heartless like ostriches in the desert.
LAM|4|4|Because of thirst the infant's tongue sticks to the roof of its mouth; the children beg for bread, but no one gives it to them.
LAM|4|5|Those who once ate delicacies are destitute in the streets. Those nurtured in purple now lie on ash heaps.
LAM|4|6|The punishment of my people is greater than that of Sodom, which was overthrown in a moment without a hand turned to help her.
LAM|4|7|Their princes were brighter than snow and whiter than milk, their bodies more ruddy than rubies, their appearance like sapphires.
LAM|4|8|But now they are blacker than soot; they are not recognized in the streets. Their skin has shriveled on their bones; it has become as dry as a stick.
LAM|4|9|Those killed by the sword are better off than those who die of famine; racked with hunger, they waste away for lack of food from the field.
LAM|4|10|With their own hands compassionate women have cooked their own children, who became their food when my people were destroyed.
LAM|4|11|The LORD has given full vent to his wrath; he has poured out his fierce anger. He kindled a fire in Zion that consumed her foundations.
LAM|4|12|The kings of the earth did not believe, nor did any of the world's people, that enemies and foes could enter the gates of Jerusalem.
LAM|4|13|But it happened because of the sins of her prophets and the iniquities of her priests, who shed within her the blood of the righteous.
LAM|4|14|Now they grope through the streets like men who are blind. They are so defiled with blood that no one dares to touch their garments.
LAM|4|15|"Go away! You are unclean!" men cry to them. "Away! Away! Don't touch us!" When they flee and wander about, people among the nations say, "They can stay here no longer."
LAM|4|16|The LORD himself has scattered them; he no longer watches over them. The priests are shown no honor, the elders no favor.
LAM|4|17|Moreover, our eyes failed, looking in vain for help; from our towers we watched for a nation that could not save us.
LAM|4|18|Men stalked us at every step, so we could not walk in our streets. Our end was near, our days were numbered, for our end had come.
LAM|4|19|Our pursuers were swifter than eagles in the sky; they chased us over the mountains and lay in wait for us in the desert.
LAM|4|20|The LORD's anointed, our very life breath, was caught in their traps. We thought that under his shadow we would live among the nations.
LAM|4|21|Rejoice and be glad, O Daughter of Edom, you who live in the land of Uz. But to you also the cup will be passed; you will be drunk and stripped naked.
LAM|4|22|O Daughter of Zion, your punishment will end; he will not prolong your exile. But, O Daughter of Edom, he will punish your sin and expose your wickedness.
LAM|5|1|Remember, O LORD, what has happened to us; look, and see our disgrace.
LAM|5|2|Our inheritance has been turned over to aliens, our homes to foreigners.
LAM|5|3|We have become orphans and fatherless, our mothers like widows.
LAM|5|4|We must buy the water we drink; our wood can be had only at a price.
LAM|5|5|Those who pursue us are at our heels; we are weary and find no rest.
LAM|5|6|We submitted to Egypt and Assyria to get enough bread.
LAM|5|7|Our fathers sinned and are no more, and we bear their punishment.
LAM|5|8|Slaves rule over us, and there is none to free us from their hands.
LAM|5|9|We get our bread at the risk of our lives because of the sword in the desert.
LAM|5|10|Our skin is hot as an oven, feverish from hunger.
LAM|5|11|Women have been ravished in Zion, and virgins in the towns of Judah.
LAM|5|12|Princes have been hung up by their hands; elders are shown no respect.
LAM|5|13|Young men toil at the millstones; boys stagger under loads of wood.
LAM|5|14|The elders are gone from the city gate; the young men have stopped their music.
LAM|5|15|Joy is gone from our hearts; our dancing has turned to mourning.
LAM|5|16|The crown has fallen from our head. Woe to us, for we have sinned!
LAM|5|17|Because of this our hearts are faint, because of these things our eyes grow dim
LAM|5|18|for Mount Zion, which lies desolate, with jackals prowling over it.
LAM|5|19|You, O LORD, reign forever; your throne endures from generation to generation.
LAM|5|20|Why do you always forget us? Why do you forsake us so long?
LAM|5|21|Restore us to yourself, O LORD, that we may return; renew our days as of old
LAM|5|22|unless you have utterly rejected us and are angry with us beyond measure.
