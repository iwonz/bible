ZEPH|1|1|The word of the LORD which came unto Zephaniah the son of Cushi, the son of Gedaliah, the son of Amariah, the son of Hizkiah, in the days of Josiah the son of Amon, king of Judah.
ZEPH|1|2|I will utterly consume all things from off the land, saith the LORD.
ZEPH|1|3|I will consume man and beast; I will consume the fowls of the heaven, and the fishes of the sea, and the stumblingblocks with the wicked: and I will cut off man from off the land, saith the LORD.
ZEPH|1|4|I will also stretch out mine hand upon Judah, and upon all the inhabitants of Jerusalem; and I will cut off the remnant of Baal from this place, and the name of the Chemarims with the priests;
ZEPH|1|5|And them that worship the host of heaven upon the housetops; and them that worship and that swear by the LORD, and that swear by Malcham;
ZEPH|1|6|And them that are turned back from the LORD; and those that have not sought the LORD, nor enquired for him.
ZEPH|1|7|Hold thy peace at the presence of the Lord GOD: for the day of the LORD is at hand: for the LORD hath prepared a sacrifice, he hath bid his guests.
ZEPH|1|8|And it shall come to pass in the day of the LORD's sacrifice, that I will punish the princes, and the king's children, and all such as are clothed with strange apparel.
ZEPH|1|9|In the same day also will I punish all those that leap on the threshold, which fill their masters' houses with violence and deceit.
ZEPH|1|10|And it shall come to pass in that day, saith the LORD, that there shall be the noise of a cry from the fish gate, and an howling from the second, and a great crashing from the hills.
ZEPH|1|11|Howl, ye inhabitants of Maktesh, for all the merchant people are cut down; all they that bear silver are cut off.
ZEPH|1|12|And it shall come to pass at that time, that I will search Jerusalem with candles, and punish the men that are settled on their lees: that say in their heart, The LORD will not do good, neither will he do evil.
ZEPH|1|13|Therefore their goods shall become a booty, and their houses a desolation: they shall also build houses, but not inhabit them; and they shall plant vineyards, but not drink the wine thereof.
ZEPH|1|14|The great day of the LORD is near, it is near, and hasteth greatly, even the voice of the day of the LORD: the mighty man shall cry there bitterly.
ZEPH|1|15|That day is a day of wrath, a day of trouble and distress, a day of wasteness and desolation, a day of darkness and gloominess, a day of clouds and thick darkness,
ZEPH|1|16|A day of the trumpet and alarm against the fenced cities, and against the high towers.
ZEPH|1|17|And I will bring distress upon men, that they shall walk like blind men, because they have sinned against the LORD: and their blood shall be poured out as dust, and their flesh as the dung.
ZEPH|1|18|Neither their silver nor their gold shall be able to deliver them in the day of the LORD's wrath; but the whole land shall be devoured by the fire of his jealousy: for he shall make even a speedy riddance of all them that dwell in the land.
ZEPH|2|1|Gather yourselves together, yea, gather together, O nation not desired;
ZEPH|2|2|Before the decree bring forth, before the day pass as the chaff, before the fierce anger of the LORD come upon you, before the day of the LORD's anger come upon you.
ZEPH|2|3|Seek ye the LORD, all ye meek of the earth, which have wrought his judgment; seek righteousness, seek meekness: it may be ye shall be hid in the day of the LORD's anger.
ZEPH|2|4|For Gaza shall be forsaken, and Ashkelon a desolation: they shall drive out Ashdod at the noon day, and Ekron shall be rooted up.
ZEPH|2|5|Woe unto the inhabitants of the sea coast, the nation of the Cherethites! the word of the LORD is against you; O Canaan, the land of the Philistines, I will even destroy thee, that there shall be no inhabitant.
ZEPH|2|6|And the sea coast shall be dwellings and cottages for shepherds, and folds for flocks.
ZEPH|2|7|And the coast shall be for the remnant of the house of Judah; they shall feed thereupon: in the houses of Ashkelon shall they lie down in the evening: for the LORD their God shall visit them, and turn away their captivity.
ZEPH|2|8|I have heard the reproach of Moab, and the revilings of the children of Ammon, whereby they have reproached my people, and magnified themselves against their border.
ZEPH|2|9|Therefore as I live, saith the LORD of hosts, the God of Israel, Surely Moab shall be as Sodom, and the children of Ammon as Gomorrah, even the breeding of nettles, and saltpits, and a perpetual desolation: the residue of my people shall spoil them, and the remnant of my people shall possess them.
ZEPH|2|10|This shall they have for their pride, because they have reproached and magnified themselves against the people of the LORD of hosts.
ZEPH|2|11|The LORD will be terrible unto them: for he will famish all the gods of the earth; and men shall worship him, every one from his place, even all the isles of the heathen.
ZEPH|2|12|Ye Ethiopians also, ye shall be slain by my sword.
ZEPH|2|13|And he will stretch out his hand against the north, and destroy Assyria; and will make Nineveh a desolation, and dry like a wilderness.
ZEPH|2|14|And flocks shall lie down in the midst of her, all the beasts of the nations: both the cormorant and the bittern shall lodge in the upper lintels of it; their voice shall sing in the windows; desolation shall be in the thresholds; for he shall uncover the cedar work.
ZEPH|2|15|This is the rejoicing city that dwelt carelessly, that said in her heart, I am, and there is none beside me: how is she become a desolation, a place for beasts to lie down in! every one that passeth by her shall hiss, and wag his hand.
ZEPH|3|1|Woe to her that is filthy and polluted, to the oppressing city!
ZEPH|3|2|She obeyed not the voice; she received not correction; she trusted not in the LORD; she drew not near to her God.
ZEPH|3|3|Her princes within her are roaring lions; her judges are evening wolves; they gnaw not the bones till the morrow.
ZEPH|3|4|Her prophets are light and treacherous persons: her priests have polluted the sanctuary, they have done violence to the law.
ZEPH|3|5|The just LORD is in the midst thereof; he will not do iniquity: every morning doth he bring his judgment to light, he faileth not; but the unjust knoweth no shame.
ZEPH|3|6|I have cut off the nations: their towers are desolate; I made their streets waste, that none passeth by: their cities are destroyed, so that there is no man, that there is none inhabitant.
ZEPH|3|7|I said, Surely thou wilt fear me, thou wilt receive instruction; so their dwelling should not be cut off, howsoever I punished them: but they rose early, and corrupted all their doings.
ZEPH|3|8|Therefore wait ye upon me, saith the LORD, until the day that I rise up to the prey: for my determination is to gather the nations, that I may assemble the kingdoms, to pour upon them mine indignation, even all my fierce anger: for all the earth shall be devoured with the fire of my jealousy.
ZEPH|3|9|For then will I turn to the people a pure language, that they may all call upon the name of the LORD, to serve him with one consent.
ZEPH|3|10|From beyond the rivers of Ethiopia my suppliants, even the daughter of my dispersed, shall bring mine offering.
ZEPH|3|11|In that day shalt thou not be ashamed for all thy doings, wherein thou hast transgressed against me: for then I will take away out of the midst of thee them that rejoice in thy pride, and thou shalt no more be haughty because of my holy mountain.
ZEPH|3|12|I will also leave in the midst of thee an afflicted and poor people, and they shall trust in the name of the LORD.
ZEPH|3|13|The remnant of Israel shall not do iniquity, nor speak lies; neither shall a deceitful tongue be found in their mouth: for they shall feed and lie down, and none shall make them afraid.
ZEPH|3|14|Sing, O daughter of Zion; shout, O Israel; be glad and rejoice with all the heart, O daughter of Jerusalem.
ZEPH|3|15|The LORD hath taken away thy judgments, he hath cast out thine enemy: the king of Israel, even the LORD, is in the midst of thee: thou shalt not see evil any more.
ZEPH|3|16|In that day it shall be said to Jerusalem, Fear thou not: and to Zion, Let not thine hands be slack.
ZEPH|3|17|The LORD thy God in the midst of thee is mighty; he will save, he will rejoice over thee with joy; he will rest in his love, he will joy over thee with singing.
ZEPH|3|18|I will gather them that are sorrowful for the solemn assembly, who are of thee, to whom the reproach of it was a burden.
ZEPH|3|19|Behold, at that time I will undo all that afflict thee: and I will save her that halteth, and gather her that was driven out; and I will get them praise and fame in every land where they have been put to shame.
ZEPH|3|20|At that time will I bring you again, even in the time that I gather you: for I will make you a name and a praise among all people of the earth, when I turn back your captivity before your eyes, saith the LORD.
