2COR|1|1|奉上帝旨意作基督耶穌使徒的 保羅 和弟兄 提摩太 ，寫信給在 哥林多 上帝的教會和全 亞該亞 的眾聖徒。
2COR|1|2|願恩惠、平安 從我們的父上帝和主耶穌基督歸給你們！
2COR|1|3|願頌讚歸於上帝—我們主耶穌基督的父；他是發慈悲的父，賜各樣安慰的上帝。
2COR|1|4|我們在一切患難中，他安慰我們，使我們能用上帝所賜的安慰去安慰那些遭各樣患難的人。
2COR|1|5|正如我們跟基督同受許多苦楚，我們也靠基督得許多安慰。
2COR|1|6|如果我們受患難，那是為使你們得安慰，得拯救；如果我們得安慰，那也是為使你們得安慰，這安慰能使你們忍受我們所受同樣的苦楚。
2COR|1|7|我們為你們所存的盼望是確定的，因為知道你們分擔了我們的痛苦，也要分享我們的安慰。
2COR|1|8|弟兄們，我們不要你們不知道，我們從前在 亞細亞 遭遇苦難，因受到無法忍受的壓力，甚至連活命的指望都沒有了。
2COR|1|9|自己心裏也斷定是必死無疑，這是要使我們不依靠自己，只依靠使死人復活的上帝。
2COR|1|10|他曾救我們脫離那極大的死亡，他要繼續救我們，而且我們指望他將來還要救我們。
2COR|1|11|你們也要一同用祈禱來幫助我們，好使許多人為我們感恩，因著他們許多的禱告，我們獲得了恩賜。
2COR|1|12|我們所誇的是：我們在世為人，特別是跟你們的關係，是憑著上帝所賜的坦率和真誠，不是靠人的聰明，而是靠上帝的恩惠；這是我們的良心可以作證的。
2COR|1|13|我們現在寫給你們的話，無非是你們所能誦讀、所能明白的，我也盼望你們真能徹底明白。
2COR|1|14|你們已經有幾分認識我們，在我們主耶穌 的日子，你們會以我們為榮，正像我們也以你們為榮。
2COR|1|15|既然我這樣深信，早就有意先到你們那裏去，讓你們得加倍的益處。
2COR|1|16|我要路過你們那裏往 馬其頓 去，再從 馬其頓 回到你們那裏，讓你們給我送行往 猶太 去。
2COR|1|17|我有此意，難道是反覆不定嗎？難道我的意願是從私慾起的，以致我忽是忽非嗎？
2COR|1|18|我指著信實的上帝說，我們向你們所傳的道並非又是又非的。
2COR|1|19|因為，我、 西拉 和 提摩太 在你們中間傳上帝的兒子耶穌基督，從沒有「又是又非」的；在他只有一個「是」。
2COR|1|20|上帝的應許，不論有多少，在基督都是「是」的。所以，我們藉著他說「阿們」，使上帝因我們得榮耀。
2COR|1|21|那在基督裏堅固我們和你們，並且膏抹我們的，就是上帝。
2COR|1|22|他在我們身上蓋了印，並賜聖靈在我們心裏作憑據。
2COR|1|23|我指著我的性命求告上帝作證，我沒有再往 哥林多 去是為了要寬容你們。
2COR|1|24|我們並不是要控制你們的信心，而是要作你們的同工，讓你們得快樂，因為你們在信仰上已經站得穩了。
2COR|2|1|我自己定了主意，下次不再帶著悲傷到你們那裏去。
2COR|2|2|我若使你們悲傷，除了因我而使他悲傷的那人以外，誰能使我喜樂呢？
2COR|2|3|我曾把這事寫給你們，免得我到的時候，那該令我喜樂的人反倒令我悲傷。我也深信，你們眾人都以我的喜樂為自己的喜樂。
2COR|2|4|我先前憂心忡忡、眼淚汪汪地給你們寫了信，並非要使你們悲傷，而是要你們知道我格外疼愛你們。
2COR|2|5|如果有人使人悲傷，他不但使我悲傷，也是使你們眾人有些悲傷。我說有些，恐怕說得太重了。
2COR|2|6|這樣的人受了大多數人的責備也就夠了，
2COR|2|7|倒不如赦免他，安慰他，免得他過分悲傷，甚至受不了啦！
2COR|2|8|所以，我勸你們，要向他肯定你們的愛心。
2COR|2|9|為此，我先前也寫信給你們，正是要考驗你們，看你們是否在一切事上都順從我。
2COR|2|10|你們赦免誰，我也赦免誰。我若有所赦免，是在基督面前為你們的緣故赦免的，
2COR|2|11|免得撒但趁著機會勝過我們，因我們並非不知道他的詭計。
2COR|2|12|我從前為基督的福音到了 特羅亞 ，主給我開了門。
2COR|2|13|那時，因為沒有遇見我的弟兄 提多 ，我心裏不安，就辭別那裏的人，往 馬其頓 去了。
2COR|2|14|感謝上帝！他常率領我們在基督裏得勝，並藉著我們在各處顯揚那因認識基督而有的香氣。
2COR|2|15|因為無論在得救的人或在滅亡的人當中，我們都是基督馨香之氣，是獻給上帝的。
2COR|2|16|對滅亡的人，這是死而又死的氣味；對得救的人，這是生而又生的氣味。這些事誰能當得起呢？
2COR|2|17|我們不像許多人，把上帝的道當商品販賣，而是由於真誠，而是受命於上帝，在上帝面前憑著基督講道。
2COR|3|1|難道我們又開始推薦自己嗎？難道我們像某些人那樣要用人的推薦信介紹給你們，或用你們的推薦信給人嗎？
2COR|3|2|你們就是我們的推薦信，寫在我們心裏，被眾人所知道、所誦讀的，
2COR|3|3|而你們顯明自己是基督的書信，藉著我們寫成的。不是用墨寫的，而是用永生上帝的靈寫的；不是寫在石版上，而是寫在心版上的。
2COR|3|4|我們藉著基督才對上帝有這樣的信心。
2COR|3|5|並不是我們憑自己配做甚麼事，我們之所以配做是出於上帝；
2COR|3|6|他使我們能配作新約的執事，不是文字上的約，而是聖靈的約；因為文字使人死，聖靈能使人活。
2COR|3|7|那用字刻在石頭上屬死的事奉尚且有榮光，以致 以色列 人因 摩西 臉上那逐漸褪色的榮光不能定睛看他的臉，
2COR|3|8|那屬聖靈的事奉不是更有榮光嗎？
2COR|3|9|若是那使人定罪的事奉有榮光，那使人稱義的事奉的榮光就越發大了。
2COR|3|10|那從前有榮光的，因這更大的榮光，就算不得有榮光了；
2COR|3|11|若是那逐漸褪色的有榮光，這長存的就更有榮光了。
2COR|3|12|既然我們有這樣的盼望，就大有膽量，
2COR|3|13|不像 摩西 將面紗蒙在臉上，使 以色列 人不能定睛看到那逐漸褪色的榮光的結局。
2COR|3|14|但他們的心地剛硬，直到今日誦讀舊約的時候，這同樣的面紗還沒有揭去；因為這面紗在基督裏才被廢去。
2COR|3|15|然而直到今日，每逢誦讀 摩西 書的時候，面紗還在他們心上。
2COR|3|16|但他們的心何時歸向主，面紗就何時除去。
2COR|3|17|主就是那靈；主的靈在哪裏，哪裏就有自由。
2COR|3|18|既然我們眾人以揭去面紗的臉得以看見 主的榮光，好像從鏡子裏返照，就變成了與主有同樣的形像，榮上加榮，如同從主的靈 變成的。
2COR|4|1|所以，既然我們蒙憐憫受了這事奉的責任，就不喪膽，
2COR|4|2|反而把那些暗昧可恥的事棄絕了，不行詭詐，不曲解上帝的道，只將真理顯揚出來，好在上帝面前把自己推薦給各人的良心。
2COR|4|3|即使我們的福音被遮蔽，那只是對滅亡的人遮蔽。
2COR|4|4|這些不信的人被這世界的神明弄瞎了心眼，使他們看不見基督榮耀的福音。基督本是上帝的像。
2COR|4|5|我們不是傳自己，而是傳耶穌基督為主，並且自己因耶穌作你們的僕人。
2COR|4|6|那吩咐光從黑暗裏照出來的上帝已經照在我們心裏，使我們知道上帝榮耀的光顯在耶穌基督的臉上。
2COR|4|7|我們有這寶貝放在瓦器裏，為要顯明這莫大的能力是出於上帝，不是出於我們。
2COR|4|8|我們處處受困，卻不被捆住；內心困擾，卻沒有絕望；
2COR|4|9|遭受迫害，卻不被撇棄；擊倒在地，卻不致滅亡。
2COR|4|10|我們身上常帶著耶穌的死，使耶穌的生也在我們身上顯明。
2COR|4|11|因為我們這活著的人常為耶穌被置於死地，使耶穌的生命在我們這必死的人身上顯明出來。
2COR|4|12|這樣看來，死是在我們身上運作，生卻在你們身上運作。
2COR|4|13|但我們既然有從同一位靈而來的信心，正如經上記著：「我信，故我說話」，我們也信，所以也說話；
2COR|4|14|因為知道，那使主耶穌復活的也必使我們與耶穌一同復活，並且使我們與你們一起站在他面前。
2COR|4|15|凡事都是為了你們，好使恩惠既藉著更多的人而加增，感恩也格外顯多，好歸榮耀給上帝。
2COR|4|16|所以，我們不喪膽。雖然我們外在的人日漸朽壞，內在的人卻日日更新。
2COR|4|17|我們這短暫而輕微的苦楚要為我們成就極重、無比、永遠的榮耀。
2COR|4|18|因為我們不是顧念看得見的，而是顧念看不見的；原來看得見的是暫時的，看不見的才是永遠的。
2COR|5|1|因為我們知道，我們這地上的帳篷若拆毀了，我們將有上帝所造的居所，不是人手所造的，而是在天上永存的。
2COR|5|2|我們在這帳篷裏嘆息，渴望得到那從天上來的居所，好像穿上衣服；
2COR|5|3|倘若脫下也 不至於赤身了。
2COR|5|4|其實，我們在這帳篷裏的人勞苦嘆息，並不是願意脫下地上的帳篷，而是願意穿上天上的居所，好使這必死的被生命吞滅了。
2COR|5|5|那為我們安排這事的是上帝，他賜給我們聖靈作憑據 。
2COR|5|6|所以，我們總是勇敢的，並且知道，只要我們住在這身體內就是離開了主。
2COR|5|7|因為我們行事為人是憑著信心，不是憑著眼見。
2COR|5|8|我們勇敢，更情願離開身體，與主同住。
2COR|5|9|所以，無論是住在身內或住在身外，我們都立了志向要得主的喜悅。
2COR|5|10|因為我們眾人必須站在基督審判臺前受審，為使各人按著本身所行的，或善或惡受報。
2COR|5|11|既然我們知道主是可畏的，就勸導人；但是上帝是認識我們的，我盼望你們的良心也認識我們。
2COR|5|12|我們不是向你們再推薦自己，而是要讓你們有誇耀我們的機會，使你們好面對那憑外貌、不憑內心誇耀的人。
2COR|5|13|如果我們癲狂，是為上帝；如果我們清醒，是為你們。
2COR|5|14|原來基督的愛激勵我們；因我們這樣斷定，一人既替眾人死了，眾人就都死了。
2COR|5|15|並且他替眾人死，是叫那些活著的人不再為自己活，乃為替他們死而復活的主活。
2COR|5|16|所以，從今以後，我們不再按照人的看法來認識人，縱使我們曾經按照人的看法認識基督，如今卻不再這樣認識他了。
2COR|5|17|所以，若有人在基督裏，他就是新造的人：舊事已過，都變成新的了。
2COR|5|18|一切都是出於上帝；他藉著基督使我們與他和好，又將勸人與他和好的使命賜給我們。
2COR|5|19|這就是：上帝在基督裏使世人與自己和好，不將他們的過犯歸到他們身上，並且將這和好的信息託付了我們。
2COR|5|20|所以，我們作基督的特使，就好像上帝藉我們勸你們一般。我們替基督求你們，與上帝和好吧！
2COR|5|21|上帝使那無罪 的，替我們成為罪，好使我們在他裏面成為上帝的義。
2COR|6|1|我們與上帝同工的也勸你們，不可白受他的恩典；
2COR|6|2|因為他說： 「在悅納的時候，我應允了你； 在拯救的日子，我幫助了你。」 看哪，現在正是悅納的時候！看哪，現在正是拯救的日子！
2COR|6|3|我們不在任何事上妨礙任何人，免得這使命被人毀謗；
2COR|6|4|反倒在各樣的事上表明自己是上帝的用人：就如在持久的忍耐、患難、困苦、災難、
2COR|6|5|鞭打、監禁、動亂、勞碌、失眠、飢餓、
2COR|6|6|廉潔、知識、堅忍、恩慈、聖靈的感化、無偽的愛心、
2COR|6|7|真實的言語、上帝的大能、藉著仁義的兵器在左在右、
2COR|6|8|榮譽或羞辱、惡名或美名。我們似乎是誘惑人的，卻是誠實的；
2COR|6|9|似乎不為人所知，卻是人所共知；似乎是死了，卻是活著；似乎受懲罰，卻沒有被處死；
2COR|6|10|似乎憂愁，卻常有喜樂；似乎貧窮，卻使許多人富足；似乎一無所有，卻樣樣都有。
2COR|6|11|哥林多 人哪，我們對你們，口是誠實的，心是寬宏的。
2COR|6|12|你們的狹窄不是由於我們，而是由於你們自己的心腸狹窄。
2COR|6|13|你們也要照樣用寬宏的心報答我；我這話正像對自己的孩子說的。
2COR|6|14|你們不要和不信的人同負一軛。義和不義有甚麼相關？光明和黑暗有甚麼相連？
2COR|6|15|基督和 彼列 有甚麼相和？信主的和不信主的有甚麼相干？
2COR|6|16|上帝的殿和偶像有甚麼相同？因為我們是永生上帝的殿，就如上帝曾說： 「我要在他們中間居住來往； 我要作他們的上帝， 他們要作我的子民。」
2COR|6|17|所以主說： 「你們務要從他們中間出來， 跟他們分別； 不要沾不潔淨的東西， 我就收納你們。
2COR|6|18|我要作你們的父， 你們要作我的兒女。 這是全能的主說的。」
2COR|7|1|所以，親愛的，既然我們有這樣的應許，就當潔淨自己，除去身體和靈魂一切的污穢，藉著敬畏上帝，得以成聖。
2COR|7|2|寬宏大量地接納我們吧！我們未曾虧負誰，未曾敗壞誰，未曾佔誰的便宜。
2COR|7|3|我說這話，不是要定你們的罪，我已經說過，你們常在我們心裏，我們情願與你們同生共死。
2COR|7|4|我對你們很是放心，多多誇耀你們；我滿有安慰，在我們一切患難中格外喜樂。
2COR|7|5|我們從前到了 馬其頓 的時候，身體沒有絲毫安寧，反而到處遭患難，外有紛爭，內有懼怕。
2COR|7|6|但那安慰灰心之人的上帝藉著 提多 來安慰了我們；
2COR|7|7|不但藉著他來，也藉著他從你們所得的安慰安慰了我們，因為他把你們的思念，你們的哀慟，你們對我的熱忱，都告訴了我，使我更加歡喜。
2COR|7|8|即使我先前那封信使你們憂愁，後來我曾懊悔，如今卻不懊悔；因為我知道，那封信使你們憂愁，不過是暫時的。
2COR|7|9|如今我歡喜，不是因你們曾憂愁，而是因憂愁導致你們的悔改。你們依著上帝的意思憂愁，凡事就不至於因我們受虧損了。
2COR|7|10|因為依著上帝的意思而憂愁，就生出沒有懊悔的悔改來，以致得救；但世俗的憂愁叫人死。
2COR|7|11|你看，你們依著上帝的意思而憂愁，這在你們當中產生了何等的殷勤、甚至辯白、甚至憤慨、甚至恐懼、甚至渴望、甚至熱忱、甚至責罰。在這一切事上，你們都表明自己是無可指責的。
2COR|7|12|所以，雖然我從前寫信給你們，卻不是為那虧負人的，也不是為那受人虧負的，而是要在上帝面前把你們顧念我們的熱忱表現出來。
2COR|7|13|因此，我們得了安慰。 在我們所得的安慰之外，又因你們眾人使 提多 心裏暢快喜樂，我們就更加歡喜了。
2COR|7|14|我若對 提多 誇獎過你們甚麼，也不覺得慚愧，因為我對 提多 誇獎你們的話是真的，正如我對你們所說的話也向來都是真的。
2COR|7|15|提多 一想起你們眾人的順服，怎樣恐懼戰兢地接待他，他愛你們的心就越發熱切了。
2COR|7|16|我如今歡喜，因為我在一切事上對你們有信心。
2COR|8|1|弟兄們，我們要把上帝賜給 馬其頓 眾教會的恩惠告訴你們：
2COR|8|2|他們在患難中受大考驗的時候，仍然滿有喜樂，在極度貧窮中還格外顯出他們樂捐的慷慨。
2COR|8|3|我可以證明，他們是按著能力，而且超過了能力來捐助，主動
2COR|8|4|再三懇求我們，准他們在這供給聖徒的善事上有份；
2COR|8|5|並且他們所做的，不但照我們所期望的，更照上帝的旨意先把自己獻給主，又給了我們。
2COR|8|6|因此，我們勸 提多 ，既然在你們中間開始這慈善的事，就當把它辦成。
2COR|8|7|既然你們在信心、口才、知識、萬分的熱忱，以及我們對你們 的愛心上，都勝人一等，那麼，當在這慈善的事上也要勝人一等。
2COR|8|8|我說這話，並不是命令你們，而是藉著別人的熱忱來考驗你們愛心的真誠。
2COR|8|9|你們知道我們主耶穌基督的恩典：他本是富足，卻為你們成了貧窮，好使你們因他的貧窮而成為富足。
2COR|8|10|我在這事上把我的意見告訴你們，是對你們有益，因為你們開始辦這事，而且起此心意已經有一年了。
2COR|8|11|如今就當辦成這事，既然有願做的心，也當照你們所有的去辦成。
2COR|8|12|因為人只要有願做的心，必照他所有的蒙悅納，並不是照他所沒有的。
2COR|8|13|我不是要別人輕鬆，你們受累，而是要均勻：
2COR|8|14|就是要你們現在的富餘補他們的不足，使他們的富餘將來也可以補你們的不足，這就均勻了。
2COR|8|15|如經上所記： 多收的沒有餘， 少收的也沒有缺。
2COR|8|16|感謝上帝，把我對你們的熱忱同樣放在 提多 心裏。
2COR|8|17|他固然聽了我的勸告，但自己更加熱心，自願往你們那裏去。
2COR|8|18|我們還差遣一位弟兄和他同去，這人在傳福音的事上得了眾教會的稱讚；
2COR|8|19|不但這樣，他也被眾教會選派跟我們同行，把所交託我們的這捐款送到了，為的是榮耀主，也表明我們的好意。
2COR|8|20|我們這樣做，免得有人因我們收的捐款多而挑剔我們。
2COR|8|21|我們留心做好事，不但在主面前，就是在人面前也是這樣。
2COR|8|22|我們又差遣一位弟兄同去。這人的熱忱，我們在許多事上屢次考驗過，現在他因為深深信任你們，就更加熱心了。
2COR|8|23|至於 提多 ，他是我的夥伴，為服事你們作我的同工。至於那兩位弟兄，他們是眾教會的使者，是基督的榮耀。
2COR|8|24|所以，你們務要在眾教會面前向他們顯明你們的愛心和我所誇獎你們的憑據。
2COR|9|1|關於供給聖徒的事，我本來不必寫信給你們；
2COR|9|2|因為我知道你們的好意，常對 馬其頓 人誇獎你們，說 亞該亞 人預備好已經有一年了。你們的熱心感動了許多人。
2COR|9|3|但我差遣那幾位弟兄去，要使你們照我的話預備妥當，免得我們在這事上誇獎你們的話落了空。
2COR|9|4|萬一有 馬其頓 人與我同去，見你們沒有預備好，就使我們所確信的反成了羞愧；你們的羞愧更不用說了。
2COR|9|5|因此，我想必須鼓勵那幾位弟兄先到你們那裏去，把從前所應許的捐款預備妥當，好顯出你們所捐的是出於樂意，不是出於勉強。
2COR|9|6|還有一點：「少種的少收；多種的多收。」
2COR|9|7|各人要隨心所願，不要為難，不要勉強，因為上帝愛樂捐的人。
2COR|9|8|上帝能將各樣的恩惠多多加給你們，使你們凡事常常充足，能多做各樣善事。
2COR|9|9|如經上所記： 「他施捨，賙濟貧窮； 他的義行存到永遠。」
2COR|9|10|那賜種子給撒種的，賜糧食給人吃的，必多多加給你們種地的種子，又增添你們仁義的果子。
2COR|9|11|你們必凡事富足，能多多施捨，使人藉著我們而生感謝上帝的心。
2COR|9|12|因為辦這供給的事，不但補聖徒的缺乏，而且使許多人對上帝充滿更多的感謝。
2COR|9|13|他們從這供給的事上得了憑據，知道你們宣認基督，順服他的福音，慷慨捐助給他們和眾人，把榮耀歸給上帝。
2COR|9|14|他們也因上帝極大的恩賜顯在你們身上而切切想念你們，為你們祈禱。
2COR|9|15|感謝上帝，因他有說不盡的恩賜！
2COR|10|1|我－ 保羅 與你們見面的時候是溫和的，不在你們那裏的時候向你們是勇敢的，如今親自藉著基督的溫柔和慈祥勸你們。
2COR|10|2|有人認為我們是憑著血氣行事，我認為必須敢於對付這等人；我但求在那裏的時候，不必這樣勇敢。
2COR|10|3|我們雖然在血氣中行事，卻不憑著血氣爭戰。
2COR|10|4|因為我們爭戰的兵器本不是屬血氣的，而是憑著上帝的能力，能夠攻破堅固的營壘。我們攻破各樣的計謀，
2COR|10|5|和各樣攔阻人認識上帝的高壘，又奪回人心來順服基督。
2COR|10|6|我已經預備好了，等你們完全順服的時候來懲罰所有不順服的人。
2COR|10|7|你們只看事情的外表。倘若有人自信是屬基督的，他要再想想，他屬基督，我們也屬基督。
2COR|10|8|主賜給我們權柄，是要造就你們，並不是要拆毀你們；我就是為這權柄稍微誇口也不覺得慚愧。
2COR|10|9|我說這話，免得你們以為我寫信是要恐嚇你們。
2COR|10|10|因為有人說：「他信上的語氣既嚴厲又強硬，他本人卻軟弱無能，言語粗俗。」
2COR|10|11|這等人當明白，我們不在那裏時信上怎麼說，見面時也必怎麼做。
2COR|10|12|因為我們不敢將自己和某些自我推薦的人並列相比；他們用自己度量自己，用自己比較自己，是不明智的。
2COR|10|13|我們不願意過分誇口，但是我們只在上帝劃定的界限內誇口。這界限甚至擴展到你們那裏。
2COR|10|14|我們擴展到你們那裏時並沒有越過了自己的界限，其實我們是首先到你們那裏傳基督福音的。
2COR|10|15|我們不靠別人所勞碌的過分誇口；我們只希望你們信心增長的時候，所劃定給我們的範圍也能夠因著你們更加擴展，
2COR|10|16|使福音得以傳到你們以外的地方，而不在別人的範圍之內，以別人所成就的事誇口。
2COR|10|17|但「要誇耀的，該誇耀主」。
2COR|10|18|因為蒙悅納的，不是自我稱許的，而是主所稱許的。
2COR|11|1|但願你們容忍我小小的愚蠢；請你們務必容忍我。
2COR|11|2|我以上帝嫉妒的愛來愛你們，因為我曾把你們許配給一個丈夫，要把你們如同貞潔的童女獻給基督。
2COR|11|3|我只怕你們的心偏邪了，失去那向基督所獻誠懇貞潔 的心，就像蛇用詭詐誘惑了 夏娃 一樣。
2COR|11|4|假如有人來，傳另一個耶穌，不是我們所傳過的；或者你們另受一個靈，不是你們所受過的聖靈；或者接納另一個福音，不是你們所接納過的；你們居然容忍了！
2COR|11|5|但我想，我一點也不在那些超級使徒以下。
2COR|11|6|雖然我不擅長說話，我的知識卻不如此。這點我們已經在每一方面各樣事上向你們表明了。
2COR|11|7|我貶低自己，為了使你們高升，因為我白白地傳上帝的福音給你們，難道這算是我犯了錯嗎？
2COR|11|8|我剝奪了別的教會，向他們取了報酬來效勞你們。
2COR|11|9|我在你們那裏有缺乏的時候，並沒有連累你們一個人，因為我所缺乏的，那些從 馬其頓 來的弟兄都補足了。我向來凡事謹慎，將來也必謹慎，總不要連累你們。
2COR|11|10|既有基督的真誠在我裏面，在 亞該亞 一帶地方就沒有人能阻止我這樣自誇。
2COR|11|11|為甚麼呢？是因我不愛你們嗎？上帝知道，我愛你們！
2COR|11|12|我現在所做的，將來還要做，為要斷絕那些尋機會之人的機會，不讓他們在所誇耀的事上被人認為與我們一樣。
2COR|11|13|那樣的人是假使徒，行事詭詐，裝作基督的使徒。
2COR|11|14|這也不足為奇，因為連撒但也裝作光明的天使。
2COR|11|15|所以，他的差役若裝作公義的差役也沒有甚麼大不了。他們的結局必然跟他們的行為相符。
2COR|11|16|我再說，誰都不可把我看作愚蠢的；即使你們把我當作愚蠢人，那麼，也讓我稍微誇誇口吧。
2COR|11|17|我說的話不是奉主的權柄說的，而是像愚蠢人具有自信地放膽誇口。
2COR|11|18|既然有好些人憑著血氣在誇口，我也要誇口了。
2COR|11|19|你們是聰明人，竟能甘心容忍愚蠢人！
2COR|11|20|假若有人奴役你們，或侵吞你們，或壓榨你們，或侮辱你們，或打你們的臉，你們居然都能容忍。
2COR|11|21|說來慚愧，在這方面好像我們是太軟弱了。 然而，我說句蠢話，人在甚麼事上敢誇口，我也敢誇口。
2COR|11|22|他們是 希伯來 人嗎？我也是。他們是 以色列 人嗎？我也是。他們是 亞伯拉罕 的後裔嗎？我也是。
2COR|11|23|他們是基督的用人嗎？我說句狂話，我更是。我比他們忍受更多勞苦，坐過更多次監牢，受過無數次的鞭打，常常冒死。
2COR|11|24|我被 猶太 人鞭打五次，每次四十減去一下；
2COR|11|25|被棍打了三次，被石頭打了一次，遭海難三次，一晝一夜在深海裏掙扎。
2COR|11|26|我又屢次行遠路，遭江河的危險，盜賊的危險，同族人的危險，外族人的危險，城裏的危險，曠野的危險，海中的危險，假弟兄的危險。
2COR|11|27|我勞碌困苦，常常失眠，又飢又渴，忍飢耐寒，赤身露體。
2COR|11|28|除了這些外表的事以外，我還有為眾教會操心的事天天壓在我身上。
2COR|11|29|有誰軟弱，我不軟弱呢？有誰跌倒，我不焦急呢？
2COR|11|30|我若必須誇口，就誇我軟弱的事好了。
2COR|11|31|那永遠可稱頌之主耶穌的父上帝知道我不說謊。
2COR|11|32|在 大馬士革 的 亞哩達 王手下的提督把守 大馬士革城 ，要捉拿我，
2COR|11|33|我被人用筐子從城牆上的窗口縋下，逃脫了他的手。
2COR|12|1|雖然自誇無益，我還是不得不誇。我現在要提到主的異象和啟示。
2COR|12|2|我認識一個在基督裏的人，他在十四年前被提到第三層天上去；或在身內，我不知道，或在身外，我也不知道，只有上帝知道。
2COR|12|3|我認識的這樣的一個人—或在身內，或在身外，我都不知道，只有上帝知道—
2COR|12|4|他被提到樂園裏，聽見隱祕的言語，是人不可說的。
2COR|12|5|為這人，我要誇口；但是為我自己，除了我的軟弱以外，我並不誇口。
2COR|12|6|就是我願意誇口也不算狂，因為我會說實話；只是我絕口不談，恐怕有人把我看得太高了，過於他在我身上所看見所聽見的；
2COR|12|7|又恐怕我因所得的啟示太高深，就過於高抬自己，所以 有一根刺加在我身上，就是撒但的差役來折磨我，免得我過於高抬自己。
2COR|12|8|為了這事，我曾三次求主使這根刺離開我。
2COR|12|9|他對我說：「我的恩典是夠你用的，因為我的能力是在人的軟弱上顯得完全。」所以，我更喜歡誇耀自己的軟弱，好使基督的能力覆庇我。
2COR|12|10|為基督的緣故，我以軟弱、凌辱、艱難、迫害、困苦為可喜樂的事；因為我甚麼時候軟弱，甚麼時候就剛強了。
2COR|12|11|我成了愚蠢人，是被你們逼出來的，因為我本該被你們讚許才是。雖然我算不了甚麼，卻沒有一件事在那些超級使徒以下。
2COR|12|12|我在你們中間，用百般的忍耐，藉著神蹟、奇事、異能顯出使徒的憑據來。
2COR|12|13|除了我不曾連累你們這一件事，你們還有甚麼事不及別的教會呢？這不公平之處，請你們饒恕我吧。
2COR|12|14|如今，我準備第三次到你們那裏去。我仍不會連累你們，因為我所求的是你們，不是你們的財物。兒女不該為父母積財，父母該為兒女積財。
2COR|12|15|我也甘心樂意為你們的靈魂費財費力。難道我越愛你們，就越少得你們的愛嗎？
2COR|12|16|罷了，我自己並沒有連累你們，你們卻有人說，我施詭詐，用心計牢籠你們。
2COR|12|17|我所差遣到你們那裏去的人，我何曾藉著他們中的任何人佔過你們的便宜呢？
2COR|12|18|我勸 提多 到你們那裏去，又差遣那位弟兄與他同去， 提多 佔過你們的便宜嗎？我們的行事為人不是同一心靈 嗎？不是同一步伐嗎？
2COR|12|19|你們一直認為我們是在你們面前為自己辯護嗎？其實，我們本是在基督裏當著上帝面前說話。親愛的，一切的事都是為了造就你們。
2COR|12|20|我怕我再來的時候，見你們不合我所期望的，而你們見我也不合你們所期望的。我怕有紛爭、嫉妒、憤怒、自私、毀謗、讒言、狂傲、動亂的事。
2COR|12|21|我怕我再來的時候，我的上帝使我在你們面前蒙羞，並且又因許多人從前犯罪，行污穢、淫亂、放蕩的事，不肯悔改而悲傷。
2COR|13|1|這是我第三次要到你們那裏去。「任何指控都要憑兩個或三個證人的口述才能成立」。
2COR|13|2|對那些犯了罪的人和其餘所有的人，正如我第二次見你們的時候曾說過，現在不在你們那裏再次說：「我若再來，必不寬容。」
2COR|13|3|因為你們想求證基督是否藉著我說話。基督對你們並不是軟弱的，而是在你們裏面大有能力的。
2COR|13|4|他因軟弱被釘在十字架上，卻因上帝的大能仍然活著。我們在他裏面也成為軟弱的，但對你們，我們將因上帝的大能而與他一同活著。
2COR|13|5|你們總要省察自己是否在信仰中生活；你們要考驗自己。除非你們經不起考驗，你們自己豈不應該知道有耶穌基督在你們裏面嗎？
2COR|13|6|我希望你們知道，我們並不是經不起考驗的人。
2COR|13|7|我們祈求上帝使你們不做任何惡事；這不是要顯明我們是經得起考驗的，而是要你們行事端正，即使我們似乎經不起考驗也沒有關係。
2COR|13|8|我們不能做任何對抗真理的事，只能維護真理。
2COR|13|9|當我們軟弱而你們剛強時，我們也歡喜。我們所祈求的是：你們能成為完全人。
2COR|13|10|所以，我不在你們那裏的時候，把這些話寫給你們，好使我見你們的時候不用照主所給我的權柄嚴厲地待你們；這權柄原是為造就人，而不是為摧毀人。
2COR|13|11|末了，弟兄們，願你們喜樂。要追求完全；要接受鼓勵；要同心合意；要彼此和睦。如此，慈愛和平的上帝必與你們同在。
2COR|13|12|你們要用聖潔的吻彼此問安。眾聖徒都向你們問安。
2COR|13|13|願主耶穌基督的恩惠、上帝的慈愛、聖靈的感動常與你們眾人同在！
