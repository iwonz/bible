1TIM|1|1|Павел, Апостол Иисуса Христа по повелению Бога, Спасителя нашего, и Господа Иисуса Христа, надежды нашей,
1TIM|1|2|Тимофею, истинному сыну в вере: благодать, милость, мир от Бога, Отца нашего, и Христа Иисуса, Господа нашего.
1TIM|1|3|Отходя в Македонию, я просил тебя пребыть в Ефесе и увещевать некоторых, чтобы они не учили иному
1TIM|1|4|и не занимались баснями и родословиями бесконечными, которые производят больше споры, нежели Божие назидание в вере.
1TIM|1|5|Цель же увещания есть любовь от чистого сердца и доброй совести и нелицемерной веры,
1TIM|1|6|от чего отступив, некоторые уклонились в пустословие,
1TIM|1|7|желая быть законоучителями, но не разумея ни того, о чем говорят, ни того, что утверждают.
1TIM|1|8|А мы знаем, что закон добр, если кто законно употребляет его,
1TIM|1|9|зная, что закон положен не для праведника, но для беззаконных и непокоривых, нечестивых и грешников, развратных и оскверненных, для оскорбителей отца и матери, для человекоубийц,
1TIM|1|10|для блудников, мужеложников, человекохищников, (клеветников, скотоложников,) лжецов, клятвопреступников, и для всего, что противно здравому учению,
1TIM|1|11|по славному благовестию блаженного Бога, которое мне вверено.
1TIM|1|12|Благодарю давшего мне силу, Христа Иисуса, Господа нашего, что Он признал меня верным, определив на служение,
1TIM|1|13|меня, который прежде был хулитель и гонитель и обидчик, но помилован потому, что [так] поступал по неведению, в неверии;
1TIM|1|14|благодать же Господа нашего (Иисуса Христа) открылась [во мне] обильно с верою и любовью во Христе Иисусе.
1TIM|1|15|Верно и всякого принятия достойно слово, что Христос Иисус пришел в мир спасти грешников, из которых я первый.
1TIM|1|16|Но для того я и помилован, чтобы Иисус Христос во мне первом показал все долготерпение, в пример тем, которые будут веровать в Него к жизни вечной.
1TIM|1|17|Царю же веков нетленному, невидимому, единому премудрому Богу честь и слава во веки веков. Аминь.
1TIM|1|18|Преподаю тебе, сын [мой] Тимофей, сообразно с бывшими о тебе пророчествами, такое завещание, чтобы ты воинствовал согласно с ними, как добрый воин,
1TIM|1|19|имея веру и добрую совесть, которую некоторые отвергнув, потерпели кораблекрушение в вере;
1TIM|1|20|таковы Именей и Александр, которых я предал сатане, чтобы они научились не богохульствовать.
1TIM|2|1|Итак прежде всего прошу совершать молитвы, прошения, моления, благодарения за всех человеков,
1TIM|2|2|за царей и за всех начальствующих, дабы проводить нам жизнь тихую и безмятежную во всяком благочестии и чистоте,
1TIM|2|3|ибо это хорошо и угодно Спасителю нашему Богу,
1TIM|2|4|Который хочет, чтобы все люди спаслись и достигли познания истины.
1TIM|2|5|Ибо един Бог, един и посредник между Богом и человеками, человек Христос Иисус,
1TIM|2|6|предавший Себя для искупления всех. [Таково было] в свое время свидетельство,
1TIM|2|7|для которого я поставлен проповедником и Апостолом, – истину говорю во Христе, не лгу, – учителем язычников в вере и истине.
1TIM|2|8|Итак желаю, чтобы на всяком месте произносили молитвы мужи, воздевая чистые руки без гнева и сомнения;
1TIM|2|9|чтобы также и жены, в приличном одеянии, со стыдливостью и целомудрием, украшали себя не плетением [волос], не золотом, не жемчугом, не многоценною одеждою,
1TIM|2|10|но добрыми делами, как прилично женам, посвящающим себя благочестию.
1TIM|2|11|Жена да учится в безмолвии, со всякою покорностью;
1TIM|2|12|а учить жене не позволяю, ни властвовать над мужем, но быть в безмолвии.
1TIM|2|13|Ибо прежде создан Адам, а потом Ева;
1TIM|2|14|и не Адам прельщен; но жена, прельстившись, впала в преступление;
1TIM|2|15|впрочем спасется через чадородие, если пребудет в вере и любви и в святости с целомудрием.
1TIM|3|1|Верно слово: если кто епископства желает, доброго дела желает.
1TIM|3|2|Но епископ должен быть непорочен, одной жены муж, трезв, целомудрен, благочинен, честен, страннолюбив, учителен,
1TIM|3|3|не пьяница, не бийца, не сварлив, не корыстолюбив, но тих, миролюбив, не сребролюбив,
1TIM|3|4|хорошо управляющий домом своим, детей содержащий в послушании со всякою честностью;
1TIM|3|5|ибо, кто не умеет управлять собственным домом, тот будет ли пещись о Церкви Божией?
1TIM|3|6|Не [должен быть] из новообращенных, чтобы не возгордился и не подпал осуждению с диаволом.
1TIM|3|7|Надлежит ему также иметь доброе свидетельство от внешних, чтобы не впасть в нарекание и сеть диавольскую.
1TIM|3|8|Диаконы также [должны быть] честны, не двоязычны, не пристрастны к вину, не корыстолюбивы,
1TIM|3|9|хранящие таинство веры в чистой совести.
1TIM|3|10|И таких надобно прежде испытывать, потом, если беспорочны, [допускать] до служения.
1TIM|3|11|Равно и жены [их должны быть] честны, не клеветницы, трезвы, верны во всем.
1TIM|3|12|Диакон должен быть муж одной жены, хорошо управляющий детьми и домом своим.
1TIM|3|13|Ибо хорошо служившие приготовляют себе высшую степень и великое дерзновение в вере во Христа Иисуса.
1TIM|3|14|Сие пишу тебе, надеясь вскоре придти к тебе,
1TIM|3|15|чтобы, если замедлю, ты знал, как должно поступать в доме Божием, который есть Церковь Бога живаго, столп и утверждение истины.
1TIM|3|16|И беспрекословно – великая благочестия тайна: Бог явился во плоти, оправдал Себя в Духе, показал Себя Ангелам, проповедан в народах, принят верою в мире, вознесся во славе.
1TIM|4|1|Дух же ясно говорит, что в последние времена отступят некоторые от веры, внимая духам обольстителям и учениям бесовским,
1TIM|4|2|через лицемерие лжесловесников, сожженных в совести своей,
1TIM|4|3|запрещающих вступать в брак [и] употреблять в пищу то, что Бог сотворил, дабы верные и познавшие истину вкушали с благодарением.
1TIM|4|4|Ибо всякое творение Божие хорошо, и ничто не предосудительно, если принимается с благодарением,
1TIM|4|5|потому что освящается словом Божиим и молитвою.
1TIM|4|6|Внушая сие братиям, будешь добрый служитель Иисуса Христа, питаемый словами веры и добрым учением, которому ты последовал.
1TIM|4|7|Негодных же и бабьих басен отвращайся, а упражняй себя в благочестии,
1TIM|4|8|ибо телесное упражнение мало полезно, а благочестие на все полезно, имея обетование жизни настоящей и будущей.
1TIM|4|9|Слово сие верно и всякого принятия достойно.
1TIM|4|10|Ибо мы для того и трудимся и поношения терпим, что уповаем на Бога живаго, Который есть Спаситель всех человеков, а наипаче верных.
1TIM|4|11|Проповедуй сие и учи.
1TIM|4|12|Никто да не пренебрегает юностью твоею; но будь образцом для верных в слове, в житии, в любви, в духе, в вере, в чистоте.
1TIM|4|13|Доколе не приду, занимайся чтением, наставлением, учением.
1TIM|4|14|Не неради о пребывающем в тебе даровании, которое дано тебе по пророчеству с возложением рук священства.
1TIM|4|15|О сем заботься, в сем пребывай, дабы успех твой для всех был очевиден.
1TIM|4|16|Вникай в себя и в учение; занимайся сим постоянно: ибо, так поступая, и себя спасешь и слушающих тебя.
1TIM|5|1|Старца не укоряй, но увещевай, как отца; младших, как братьев;
1TIM|5|2|стариц, как матерей; молодых, как сестер, со всякою чистотою.
1TIM|5|3|Вдовиц почитай, истинных вдовиц.
1TIM|5|4|Если же какая вдовица имеет детей или внучат, то они прежде пусть учатся почитать свою семью и воздавать должное родителям, ибо сие угодно Богу.
1TIM|5|5|Истинная вдовица и одинокая надеется на Бога и пребывает в молениях и молитвах день и ночь;
1TIM|5|6|а сластолюбивая заживо умерла.
1TIM|5|7|И сие внушай им, чтобы были беспорочны.
1TIM|5|8|Если же кто о своих и особенно о домашних не печется, тот отрекся от веры и хуже неверного.
1TIM|5|9|Вдовица должна быть избираема не менее, как шестидесятилетняя, бывшая женою одного мужа,
1TIM|5|10|известная по добрым делам, если она воспитала детей, принимала странников, умывала ноги святым, помогала бедствующим и была усердна ко всякому доброму делу.
1TIM|5|11|Молодых же вдовиц не принимай, ибо они, впадая в роскошь в противность Христу, желают вступать в брак.
1TIM|5|12|Они подлежат осуждению, потому что отвергли прежнюю веру;
1TIM|5|13|притом же они, будучи праздны, приучаются ходить по домам и [бывают] не только праздны, но и болтливы, любопытны, и говорят, чего не должно.
1TIM|5|14|Итак я желаю, чтобы молодые вдовы вступали в брак, рождали детей, управляли домом и не подавали противнику никакого повода к злоречию;
1TIM|5|15|ибо некоторые уже совратились вслед сатаны.
1TIM|5|16|Если какой верный или верная имеет вдов, то должны их довольствовать и не обременять Церкви, чтобы она могла довольствовать истинных вдовиц.
1TIM|5|17|Достойно начальствующим пресвитерам должно оказывать сугубую честь, особенно тем, которые трудятся в слове и учении.
1TIM|5|18|Ибо Писание говорит: не заграждай рта у вола молотящего; и: трудящийся достоин награды своей.
1TIM|5|19|Обвинение на пресвитера не иначе принимай, как при двух или трех свидетелях.
1TIM|5|20|Согрешающих обличай перед всеми, чтобы и прочие страх имели.
1TIM|5|21|Пред Богом и Господом Иисусом Христом и избранными Ангелами заклинаю тебя сохранить сие без предубеждения, ничего не делая по пристрастию.
1TIM|5|22|Рук ни на кого не возлагай поспешно, и не делайся участником в чужих грехах. Храни себя чистым.
1TIM|5|23|Впредь пей не [одну] воду, но употребляй немного вина, ради желудка твоего и частых твоих недугов.
1TIM|5|24|Грехи некоторых людей явны и прямо ведут к осуждению, а некоторых [открываются] впоследствии.
1TIM|5|25|Равным образом и добрые дела явны; а если и не таковы, скрыться не могут.
1TIM|6|1|Рабы, под игом находящиеся, должны почитать господ своих достойными всякой чести, дабы не было хулы на имя Божие и учение.
1TIM|6|2|Те, которые имеют господами верных, не должны обращаться с ними небрежно, потому что они братья; но тем более должны служить им, что они верные и возлюбленные и благодетельствуют [им]. Учи сему и увещевай.
1TIM|6|3|Кто учит иному и не следует здравым словам Господа нашего Иисуса Христа и учению о благочестии,
1TIM|6|4|тот горд, ничего не знает, но заражен [страстью] к состязаниям и словопрениям, от которых происходят зависть, распри, злоречия, лукавые подозрения.
1TIM|6|5|Пустые споры между людьми поврежденного ума, чуждыми истины, которые думают, будто благочестие служит для прибытка. Удаляйся от таких.
1TIM|6|6|Великое приобретение – быть благочестивым и довольным.
1TIM|6|7|Ибо мы ничего не принесли в мир; явно, что ничего не можем и вынести [из него].
1TIM|6|8|Имея пропитание и одежду, будем довольны тем.
1TIM|6|9|А желающие обогащаться впадают в искушение и в сеть и во многие безрассудные и вредные похоти, которые погружают людей в бедствие и пагубу;
1TIM|6|10|ибо корень всех зол есть сребролюбие, которому предавшись, некоторые уклонились от веры и сами себя подвергли многим скорбям.
1TIM|6|11|Ты же, человек Божий, убегай сего, а преуспевай в правде, благочестии, вере, любви, терпении, кротости.
1TIM|6|12|Подвизайся добрым подвигом веры, держись вечной жизни, к которой ты и призван, и исповедал доброе исповедание перед многими свидетелями.
1TIM|6|13|Пред Богом, все животворящим, и пред Христом Иисусом, Который засвидетельствовал пред Понтием Пилатом доброе исповедание, завещеваю тебе
1TIM|6|14|соблюсти заповедь чисто и неукоризненно, даже до явления Господа нашего Иисуса Христа,
1TIM|6|15|которое в свое время откроет блаженный и единый сильный Царь царствующих и Господь господствующих,
1TIM|6|16|единый имеющий бессмертие, Который обитает в неприступном свете, Которого никто из человеков не видел и видеть не может. Ему честь и держава вечная! Аминь.
1TIM|6|17|Богатых в настоящем веке увещевай, чтобы они не высоко думали [о] [себе] и уповали не на богатство неверное, но на Бога живаго, дающего нам все обильно для наслаждения;
1TIM|6|18|чтобы они благодетельствовали, богатели добрыми делами, были щедры и общительны,
1TIM|6|19|собирая себе сокровище, доброе основание для будущего, чтобы достигнуть вечной жизни.
1TIM|6|20|О, Тимофей! храни преданное тебе, отвращаясь негодного пустословия и прекословий лжеименного знания,
1TIM|6|21|которому предавшись, некоторые уклонились от веры. Благодать с тобою. Аминь.
