2JOHN|1|1|我作長老的寫信給蒙揀選的夫人 和她的兒女，就是我真心所愛的；不但我愛，也是一切認識真理的人所愛的，
2JOHN|1|2|這是因為真理住在我們裏面，也必與我們同在直到永遠。
2JOHN|1|3|願恩惠、憐憫、平安 從父上帝和他兒子耶穌基督，在真理和愛中必與我們同在。
2JOHN|1|4|我非常歡喜見你的兒女，有照我們從父所受之命令遵行真理的。
2JOHN|1|5|夫人哪，我現在請求你，我們大家要彼此相愛。我寫給你的，並不是一條新命令，而是我們從起初就有的。
2JOHN|1|6|這就是愛，就是照他的命令行事；這就是命令，你們要照這命令行，正如你們從起初所聽見的。
2JOHN|1|7|有許多迷惑人的已經來到世上，他們不宣認耶穌基督是成了肉身來的；這樣的人是迷惑人的，是敵基督的。
2JOHN|1|8|你們要小心，不要失去你們 所完成的工作，而要得到充足的賞賜。
2JOHN|1|9|凡越過基督的教導而不持守的，就沒有上帝；凡持守這教導的，就有父又有子。
2JOHN|1|10|若有人到你們那裏而不傳這教導，不要接他到家裏，也不要向他問安；
2JOHN|1|11|因為向他問安的，就在他的惡行上有份。
2JOHN|1|12|我還有許多事要寫給你們，卻不願意用紙用墨，但盼望到你們那裏，與你們面對面談論，使我們的喜樂得以滿足。
2JOHN|1|13|你那蒙揀選的姊妹的兒女向你問安。
