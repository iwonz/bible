3JOHN|1|1|The elder unto the wellbeloved Gaius, whom I love in the truth.
3JOHN|1|2|Beloved, I wish above all things that thou mayest prosper and be in health, even as thy soul prospereth.
3JOHN|1|3|For I rejoiced greatly, when the brethren came and testified of the truth that is in thee, even as thou walkest in the truth.
3JOHN|1|4|I have no greater joy than to hear that my children walk in truth.
3JOHN|1|5|Beloved, thou doest faithfully whatsoever thou doest to the brethren, and to strangers;
3JOHN|1|6|Which have borne witness of thy charity before the church: whom if thou bring forward on their journey after a godly sort, thou shalt do well:
3JOHN|1|7|Because that for his name's sake they went forth, taking nothing of the Gentiles.
3JOHN|1|8|We therefore ought to receive such, that we might be fellowhelpers to the truth.
3JOHN|1|9|I wrote unto the church: but Diotrephes, who loveth to have the preeminence among them, receiveth us not.
3JOHN|1|10|Wherefore, if I come, I will remember his deeds which he doeth, prating against us with malicious words: and not content therewith, neither doth he himself receive the brethren, and forbiddeth them that would, and casteth them out of the church.
3JOHN|1|11|Beloved, follow not that which is evil, but that which is good. He that doeth good is of God: but he that doeth evil hath not seen God.
3JOHN|1|12|Demetrius hath good report of all men, and of the truth itself: yea, and we also bear record; and ye know that our record is true.
3JOHN|1|13|I had many things to write, but I will not with ink and pen write unto thee:
3JOHN|1|14|But I trust I shall shortly see thee, and we shall speak face to face. Peace be to thee. Our friends salute thee. Greet the friends by name.
