ACTS|1|1|提阿非罗 啊，我在第一本书中已论到耶稣从开头所做和所教导的一切事，
ACTS|1|2|直到他藉着圣灵吩咐所拣选的使徒后，被接上升的日子为止。
ACTS|1|3|他受害以后，用许多确据向使徒显明自己是活着的，在四十天之中向他们显现，并讲说上帝国的事。
ACTS|1|4|耶稣和他们聚集的时候，嘱咐他们说：“不要离开 耶路撒冷 ，但要等候父的应许，就是你们听见我说过的。
ACTS|1|5|约翰 是用水施洗，但过了不多几天，你们要在圣灵里受洗。”
ACTS|1|6|他们聚集的时候，问耶稣：“主啊，你就要在这时候复兴 以色列 国吗？”
ACTS|1|7|耶稣对他们说：“父凭着自己的权柄所定的时候和日期，不是你们可以知道的。
ACTS|1|8|但圣灵降临在你们身上，你们就必得着能力，并要在 耶路撒冷 、 犹太 全地和 撒玛利亚 ，直到地极，作我的见证。”
ACTS|1|9|说了这些话，他们正看的时候，他被接上升，有一朵云彩从他们眼前把他接去。
ACTS|1|10|他升上去的时候，他们定睛望天，看哪，有两个人身穿白衣站在他们旁边，
ACTS|1|11|说：“ 加利利 人哪，你们为什么站着望天呢？这离开你们被接升天的耶稣，你们见他怎样升上天去，他也要怎样来临。”
ACTS|1|12|有一座山，名叫 橄榄山 ，离 耶路撒冷 不远，有安息日可行走的路程 。那时，门徒从那里回 耶路撒冷 去，
ACTS|1|13|他们一进城，就上了所住的楼房；在那里有 彼得 、 约翰 、 雅各 、 安得烈 、 腓力 、 多马 、 巴多罗买 、 马太 、 亚勒腓 的儿子 雅各 、激进党的 西门 ，和 雅各 的儿子 犹大 。
ACTS|1|14|这些人和几个妇人，包括耶稣的母亲 马利亚 ，和耶稣的兄弟，都同心合意地恒切祷告。
ACTS|1|15|那时，有许多人聚会，约有一百二十名， 彼得 在弟兄中间站起来，说：
ACTS|1|16|“诸位弟兄，圣经的话必须应验。圣经中，圣灵曾藉 大卫 的口预先说到那领人来拿耶稣的 犹大 ；
ACTS|1|17|他本来算是我们中的一个，并且得了这一份使徒的职任。
ACTS|1|18|这人用他不义的代价买了一块田，以后身子仆倒，肚腹崩裂，肠子都流出来。
ACTS|1|19|住在 耶路撒冷 的人都知道这事，所以按着他们当地的话把那块田叫 亚革大马 ，就是“血田”的意思。
ACTS|1|20|因为《诗篇》上写着： “愿他的住处变为废墟， 无人在内居住。” 又说： “愿别人得他的职分。”
ACTS|1|21|所以，主耶稣在我们中间出入的整段时间，就是从 约翰 施洗起，直到主离开我们被接上升的日子为止，必须从那常与我们一起的人中，立一位与我们同作耶稣复活的见证。”
ACTS|1|22|
ACTS|1|23|于是他们推举两个人，就是那叫 巴撒巴 ，又称为 犹士都 的 约瑟 ，和 马提亚 。
ACTS|1|24|众人祷告说：“主啊，你知道万人的心，求你从这两个人中指明你所拣选的是哪一位，
ACTS|1|25|去得这使徒的职任；这职位 犹大 已经丢弃，往自己的地方去了。”
ACTS|1|26|于是众人为他们摇签，摇出 马提亚 来；他就和十一个使徒同列。
ACTS|2|1|五旬节那日到了，他们全都聚集在一起。
ACTS|2|2|忽然，有响声从天上下来，好像一阵大风吹过，充满了他们所坐的整座屋子；
ACTS|2|3|又有舌头如火焰向他们显现，分开落在他们每个人身上。
ACTS|2|4|他们都被圣灵充满，就按着圣灵所赐的口才说起别国的话来。
ACTS|2|5|那时，有从天下各国来的虔诚的 犹太 人，住在 耶路撒冷 。
ACTS|2|6|这声音一响，许多人都来聚集，各人因为听见门徒用他们各自的乡谈说话，就甚纳闷，
ACTS|2|7|都诧异惊奇说：“看哪，这些说话的不都是 加利利 人吗？
ACTS|2|8|我们每个人怎么听见他们说我们生来所用的乡谈呢？
ACTS|2|9|我们 帕提亚 人、 玛代 人、 以拦 人，和住在 美索不达米亚 、 犹太 、 加帕多家 、 本都 、 亚细亚 、
ACTS|2|10|弗吕家 、 旁非利亚 、 埃及 的人，并靠近 古利奈 的 利比亚 一带地方的人，侨居的 罗马 人，
ACTS|2|11|包括 犹太 人和皈依 犹太 教的人， 克里特 人和 阿拉伯 人，都听见他们用我们的乡谈讲论上帝的大作为。”
ACTS|2|12|众人就都惊奇困惑，彼此说：“这是什么意思呢？”
ACTS|2|13|还有人讥诮，说：“他们是灌满了新酒吧！”
ACTS|2|14|彼得 和十一个使徒站起来，他就高声向众人说：“ 犹太 人和所有住在 耶路撒冷 的人哪，这件事你们要知道，要侧耳听我的话。
ACTS|2|15|这些人并不像你们所想的喝醉了，因为现在才早晨九点钟。
ACTS|2|16|这正是藉着先知 约珥 所说的：
ACTS|2|17|‘上帝说： 在末后的日子， 我要将我的灵浇灌凡血肉之躯的。 你们的儿女要说预言； 你们的少年要见异象； 你们的老人要做异梦。
ACTS|2|18|在那些日子，我要把我的灵浇灌， 甚至给我的仆人和婢女， 他们要说预言。
ACTS|2|19|在天上，我要显出奇事， 在地下，我要显出神迹， 有血，有火，有烟雾。
ACTS|2|20|太阳要变为黑暗， 月亮要变为血， 这都在主大而光荣的日子未到以前。
ACTS|2|21|那时，凡求告主名的都必得救。’
ACTS|2|22|“ 以色列 人哪，你们要听我这些话： 拿撒勒 人耶稣就是上帝以异能、奇事、神迹向你们证明出来的人，这些事是上帝藉着他在你们中间施行，正如你们自己知道的。
ACTS|2|23|他既按着上帝确定的旨意和预知被交与人，你们就藉着不法之人的手把他钉在十字架上，杀了。
ACTS|2|24|上帝却将死的痛苦解除，使他复活了，因为他原不能被死拘禁。
ACTS|2|25|大卫 指着他说： ‘我看见 主常在我眼前， 他在我右边，使我不至于动摇。
ACTS|2|26|所以我心里欢喜，我的舌头快乐， 而且我的肉身要安居在指望中。
ACTS|2|27|因你必不将我的灵魂撇在阴间， 也不让你的圣者见朽坏。
ACTS|2|28|你已将生命的道路指示我， 必使我在你面前充满快乐。’
ACTS|2|29|“诸位弟兄，先祖 大卫 的事，我可以坦然地对你们说：他死了，也埋葬了，而且他的坟墓直到今日还在我们这里。
ACTS|2|30|既然 大卫 是先知，他知道上帝曾向他起誓，要从他的后裔中立一位坐在他的宝座上。
ACTS|2|31|他预先看见了，就讲论基督的复活，说： ‘他不被撇在阴间； 他的肉身也不见朽坏。’
ACTS|2|32|这耶稣，上帝已经使他复活了，我们都是这事的见证人。
ACTS|2|33|他既被高举在上帝的右边，又从父受了所应许的圣灵，就把你们所看见所听见的，浇灌下来。
ACTS|2|34|大卫 并没有升到天上，但他自己说： ‘主对我主说： 你坐在我的右边，
ACTS|2|35|等我使你的仇敌作你的脚凳。’
ACTS|2|36|故此， 以色列 全家当确实知道，你们钉在十字架上的这位耶稣，上帝已经立他为主，为基督了。”
ACTS|2|37|众人听见这话，觉得扎心，就对 彼得 和其余的使徒说：“诸位弟兄，我们该怎样做呢？”
ACTS|2|38|彼得 对他们说：“你们各人要悔改，奉耶稣基督的名受洗，使你们的罪得赦免，就会领受所赐的圣灵。
ACTS|2|39|因为这应许是给你们和你们的儿女，并一切在远方的人，就是给所有主—我们的上帝所召来的人。”
ACTS|2|40|彼得 还用更多别的话作见证，劝勉他们说：“你们当救自己脱离这弯曲的世代。”
ACTS|2|41|于是领受他话的人，都受了洗；那一天，门徒约添了三千人。
ACTS|2|42|他们都专注于使徒的教导和彼此的团契，擘饼和祈祷。
ACTS|2|43|众人都心存敬畏；使徒们 又行了许多奇事神迹。
ACTS|2|44|信的人都聚在一处，凡物公用，
ACTS|2|45|又卖了田产和家业，照每一个人所需要的分给他们。
ACTS|2|46|他们天天同心合意恒切地在圣殿里敬拜，且在家中 擘饼，存着欢喜坦诚的心用饭，
ACTS|2|47|赞美上帝，得全体百姓的喜爱。主将得救的人天天加给他们。
ACTS|3|1|下午三点钟祷告的时候， 彼得 和 约翰 上圣殿去。
ACTS|3|2|一个从母腹里就是瘸腿的人正被人抬来，他们天天把他放在圣殿的一个叫 美门 的门口，求进圣殿的人施舍。
ACTS|3|3|他看见 彼得 、 约翰 将要进圣殿，就求他们施舍。
ACTS|3|4|彼得 和 约翰 定睛看他， 彼得 说：“看着我们！”
ACTS|3|5|那人就注目看他们，指望从他们得着什么。
ACTS|3|6|彼得 却说：“金银我都没有，但我把我有的给你：奉 拿撒勒 人耶稣基督的名起来 行走！”
ACTS|3|7|于是 彼得 拉着他的右手，扶他起来；他的脚和踝骨立刻健壮了，
ACTS|3|8|就跳起来，站着，又开始行走。他跟他们进了圣殿，边走边跳，赞美上帝。
ACTS|3|9|百姓都看见他又行走，又赞美上帝，
ACTS|3|10|认得他是那素常坐在圣殿的 美门 口求人施舍的，就因他所遇到的事满心惊讶诧异。
ACTS|3|11|那人正在称为 所罗门 的廊下，拉住 彼得 和 约翰 ，大家都觉得很惊讶，一齐跑到他们那里。
ACTS|3|12|彼得 看见，就对百姓说：“ 以色列 人哪，为什么因这事而惊讶呢？为什么定睛看我们，以为我们凭自己的能力和虔诚使这人行走呢？
ACTS|3|13|亚伯拉罕 的上帝、 以撒 的上帝、 雅各 的上帝，就是我们列祖的上帝，已经荣耀了他的仆人耶稣，这耶稣就是你们交付官府的那位， 彼拉多 决定要释放他时，你们却在 彼拉多 面前弃绝了他。
ACTS|3|14|你们弃绝了那圣洁公义者，反而要求释放一个凶手给你们。
ACTS|3|15|你们杀了那生命的创始者，上帝却叫他从死人中复活；我们都是这事的见证人。
ACTS|3|16|因信他的名，他的名使你们所看见所认识的这人健壮了；正是他所赐的信心使这人在你们众人面前完全好了。
ACTS|3|17|“如今，弟兄们，我知道你们做这事是出于无知，你们的官长也是如此。
ACTS|3|18|但上帝藉着众先知的口预先宣告过基督将要受害的事，就这样应验了。
ACTS|3|19|所以，你们当悔改归正，使你们的罪得以涂去，
ACTS|3|20|这样，那安舒的日子就必从主面前来到；主也必差遣所预定给你们的基督耶稣来临。
ACTS|3|21|他必须留在天上，直到万物复兴的时候，就是上帝自古藉着圣先知的口所说的。
ACTS|3|22|摩西 曾说：‘主—你们 的上帝要从你们弟兄中给你们兴起一位先知像我，凡他向你们所说的一切，你们都要听从。
ACTS|3|23|凡不听从那先知的，必将从民中灭绝。’
ACTS|3|24|从 撒母耳 以来和后继的众先知，凡说预言的，也都曾宣告这些日子。
ACTS|3|25|你们是先知的子孙，也是上帝与你们 祖宗所立之约的子孙，就是对 亚伯拉罕 说：‘地上万族都将因你的后裔得福。’
ACTS|3|26|上帝既兴起他的仆人，就先差他到你们这里来，赐福给你们，使各人回转，离开你们的邪恶。”
ACTS|4|1|彼得 和 约翰 正向百姓说话的时候，祭司们、守殿官和撒都该人来了，
ACTS|4|2|就很烦恼，因为使徒们教导百姓，传扬在耶稣的事上证明有死人复活，
ACTS|4|3|于是下手拿住他们；因为天已经晚了，就把他们押在拘留所到第二天。
ACTS|4|4|但听道的人有许多信了，男人的数目约有五千。
ACTS|4|5|第二天，官长、长老和文士在 耶路撒冷 聚集，
ACTS|4|6|又有 亚那 大祭司、 该亚法 、 约翰 、 亚历山大 ，和大祭司的亲族都在那里。
ACTS|4|7|他们叫使徒站在中间，问他们：“你们凭什么能力，奉谁的名做这事呢？”
ACTS|4|8|那时， 彼得 被圣灵充满，对他们说：“民间的官长和长老啊，
ACTS|4|9|倘若今日我们被查问是因为在残障的人身上所行的善事，就是这人怎么得了痊愈，
ACTS|4|10|那么，你们大家和 以色列 全民都当知道，站在你们面前的这人得痊愈，是因你们所钉在十字架、上帝使他从死人中复活的 拿撒勒 人耶稣基督的名。
ACTS|4|11|这位耶稣是： ‘你们匠人所丢弃的石头， 已成了房角的头块石头。’
ACTS|4|12|除他以外，别无拯救，因为在天下人间，没有赐下别的名，我们可以靠着得救。”
ACTS|4|13|他们见 彼得 、 约翰 的胆量，又看出他们原是没有学问的平民，就很惊讶，认出他们曾是跟耶稣一起的；
ACTS|4|14|又看见那治好了的人和他们一同站着，就无话可驳。
ACTS|4|15|于是他们吩咐他们两人从议会退出，就彼此商议，
ACTS|4|16|说：“我们当怎样办这两个人呢？因为他们诚然行了一件明显的神迹，凡住在 耶路撒冷 的人都知道，我们也不能否认。
ACTS|4|17|但为避免这事越发在民间传扬，我们必须威吓他们，叫他们不可再奉这名对任何人讲论。”
ACTS|4|18|于是他们叫了两人来，禁止他们，再不可奉耶稣的名讲论或教导人。
ACTS|4|19|彼得 和 约翰 回答他们说：“听从你们，不听从上帝，在上帝面前合理不合理，你们自己判断吧！
ACTS|4|20|我们所看见所听见的，我们不能不说。”
ACTS|4|21|官长为百姓的缘故，想不出任何法子惩罚他们，只好威吓一番就把他们释放了；这是因众人为了所行的奇事都归荣耀与上帝。
ACTS|4|22|原来经历这神迹医好的人有四十多岁了。
ACTS|4|23|二人既被释放，就到自己的人那里去，把祭司长和长老所说的话都告诉他们。
ACTS|4|24|他们听见了，就同心合意地高声向上帝说：“主宰啊！你是那创造天、地、海和其中万物的；
ACTS|4|25|你曾藉着圣灵托你仆人—我们祖宗 大卫 的口说： ‘外邦为什么扰动？ 万民为什么谋算虚妄的事？
ACTS|4|26|地上的君王都站稳， 臣宰也聚集一处， 要对抗主，对抗主的受膏者 ’。
ACTS|4|27|希律 和 本丢．彼拉多 ，同外邦人和 以色列 民，果然在这城里聚集，要攻打你所膏的圣仆耶稣，
ACTS|4|28|做了你手和你旨意所预定必成就的事。
ACTS|4|29|主啊，现在求你鉴察，他们的威吓，使你仆人放胆讲你的道，
ACTS|4|30|伸出你的手来，让医治、神迹、奇事藉着你圣仆耶稣的名行出来。”
ACTS|4|31|他们祷告完了，聚会的地方震动；他们都被圣灵充满，放胆传讲上帝的道。
ACTS|4|32|许多信徒都一心一意，没有一人说他的任何东西是自己的，都是大家公用。
ACTS|4|33|使徒以大能见证主耶稣 复活；众人也都蒙了大恩。
ACTS|4|34|他们当中没有一个缺乏的，因为凡有田产房屋的都卖了，把所卖的钱拿来，
ACTS|4|35|放在使徒脚前，照每人所需要的，分给每人。
ACTS|4|36|有一个 利未 人，名叫 约瑟 ，使徒称他为 巴拿巴 （ 巴拿巴 翻出来就是安慰之子），生在 塞浦路斯 。
ACTS|4|37|他有田地，也卖了，把钱拿来，放在使徒脚前。
ACTS|5|1|有一个人，名叫 亚拿尼亚 ，同他的妻子 撒非喇 ，卖了田产，
ACTS|5|2|把钱私自留下一部分，他的妻子也知道，其余的部分拿来放在使徒脚前。
ACTS|5|3|彼得 说：“ 亚拿尼亚 ！为什么撒但充满了你的心，使你欺骗圣灵，把卖田地的钱私自留下一部分呢？
ACTS|5|4|田地还没有卖，不是你自己的吗？既卖了，钱不是你作主吗？你怎么心里会想这样做呢？你不是欺骗人，是欺骗上帝！”
ACTS|5|5|亚拿尼亚 一听见这些话，就仆倒，断了气；所有听见的人都非常惧怕。
ACTS|5|6|有些年轻人起来，把他裹好，抬出去埋葬了。
ACTS|5|7|约过了三小时，他的妻子进来，还不知道所发生的事。
ACTS|5|8|彼得 对她说：“你告诉我，你们卖田地的钱就是这些吗？”她说：“就是这些。”
ACTS|5|9|彼得 对她说：“你们为什么同谋来试探主的灵呢？你看，埋葬你丈夫之人的脚已到门口，他们也要把你抬出去。”
ACTS|5|10|她立刻仆倒在 彼得 脚前，断了气。那些年轻人进来，见她已经死了，就把她抬出去，埋在她丈夫旁边。
ACTS|5|11|全教会和所有听见这些事的人都非常惧怕。
ACTS|5|12|主藉使徒的手在民间行了许多神迹奇事；他们都同心合意地聚集在 所罗门 的廊下。
ACTS|5|13|其余的人没有一个敢接近他们，百姓却尊重他们。
ACTS|5|14|信主的人越发增添，连男带女都很多，
ACTS|5|15|甚至有人将病人抬到街上，放在床上或褥子上，好让 彼得 走过来的时候，或者影子投在一些人身上。
ACTS|5|16|还有许多人带着病人和被污灵缠磨的，从 耶路撒冷 四围的城镇来，他们全都得了医治。
ACTS|5|17|于是，大祭司采取行动，他和他所有一起的人，就是撒都该派的人，满心忌恨，
ACTS|5|18|就下手拿住使徒，把他们押在公共拘留所内。
ACTS|5|19|但在夜间主的使者开了监门，领他们出来，说：
ACTS|5|20|“你们去，站在圣殿里，把这生命的一切话讲给百姓听。”
ACTS|5|21|使徒听了这话，天将亮的时候就进圣殿里去教导人。大祭司和他一起的人来了，叫齐议会的人和 以色列 人的众长老，然后派人到监牢里去把使徒提出来。
ACTS|5|22|但差役到了，不见他们在监里，就回来禀报，
ACTS|5|23|说：“我们看见监牢关得很紧，警卫也站在门外，但打开门来，里面一个人都不见。”
ACTS|5|24|守殿官和祭司长听了这些话，心里困惑，不知这事将来如何。
ACTS|5|25|有一个人来禀报说：“你们押在监里的人，现在站在圣殿里教导百姓。”
ACTS|5|26|于是守殿官和差役去带使徒来，并没有用暴力，因为怕百姓用石头打他们。
ACTS|5|27|他们把使徒带来了，就叫他们站在议会前。大祭司问他们，
ACTS|5|28|说：“我们不是严严地禁止你们，不可奉这名教导人吗？ 看，你们倒把你们的道理充满了 耶路撒冷 ，想要叫这人的血归到我们身上！”
ACTS|5|29|彼得 和众使徒回答：“我们必须顺从上帝，胜于顺从人。
ACTS|5|30|你们挂在木头上杀害的耶稣，我们祖宗的上帝已经使他复活了。
ACTS|5|31|上帝把他高举在自己的右边，使他作元帅，作救主，使 以色列 人得以悔改，并且罪得赦免。
ACTS|5|32|我们是这些事的见证人；上帝赐给顺从的人的圣灵也为这些事作见证。”
ACTS|5|33|议会的人听了极其恼怒，想要杀他们。
ACTS|5|34|但有一个法利赛人，名叫 迦玛列 ，是众百姓所敬重的律法教师，他在议会中站起来，吩咐人把使徒暂且带到外面去，
ACTS|5|35|然后对众人说：“ 以色列 人哪，对于这些人，你们应当小心怎样处理。
ACTS|5|36|从前 杜达 出现，自命不凡，附从他的人数约有四百；他被杀后，附从他的人全都散了，归于无有。
ACTS|5|37|此后，登记户籍的时候，又有 加利利 的 犹大 出现，引诱百姓跟从他，他也灭亡，附从他的人也都四散了。
ACTS|5|38|现在，我劝你们不要管这些人，任凭他们吧！他们所谋所为若是出于人，必要败坏；
ACTS|5|39|若是出于上帝，你们就不能败坏他们，恐怕你们倒是攻击上帝了。” 议会的人被他说服了，
ACTS|5|40|就叫使徒来，把他们打了，又吩咐他们不可奉耶稣的名讲道，然后把他们释放了。
ACTS|5|41|他们欢欢喜喜地离开议会，因他们算配为这名受辱。
ACTS|5|42|他们就每日在圣殿里，在家里 ，不住地教导人，传耶稣是基督的福音。
ACTS|6|1|那些日子，门徒增多，有说希腊话的 犹太 人向 希伯来 人发怨言，因为在日常的供给上忽略了他们的寡妇。
ACTS|6|2|十二使徒叫众门徒来，说：“我们撇下上帝的道去管理饭食，是不合宜的。
ACTS|6|3|所以弟兄们，当从你们中间选出七个有好名声、满有圣灵和智慧，我们派他们管理这事。
ACTS|6|4|至于我们，我们要专注于祈祷和传道的事奉。”
ACTS|6|5|这话使全会众都喜悦，就拣选了 司提反 —他是一个满有信心和圣灵的人；他们又拣选了 腓利 、 伯罗哥罗 、 尼迦挪 、 提门 、 巴米拿 ，并皈依 犹太 教的 安提阿 人 尼哥拉 ，
ACTS|6|6|叫他们站在使徒面前，使徒祷告后，就为他们按手。
ACTS|6|7|上帝的道兴旺起来；在 耶路撒冷 门徒数目增加得很多，也有许多祭司听从了这信仰。
ACTS|6|8|司提反 满有恩惠和能力，在民间行了大奇事和神迹。
ACTS|6|9|当时有从称为“自由人”会堂，并 古利奈 、 亚历山大 会堂来的人，还有些从 基利家 、 亚细亚 来的人，起来和 司提反 辩论。
ACTS|6|10|司提反 是以智慧和圣灵说话，众人抵挡不住，
ACTS|6|11|就收买人来说：“我们听见他说亵渎 摩西 和上帝的话。”
ACTS|6|12|他们又煽动百姓、长老和文士，就突然来捉拿他，把他带到议会去，
ACTS|6|13|设下假见证，说：“这个人不断地说话，侮辱神圣的地方和律法。
ACTS|6|14|我们曾听见他说，这 拿撒勒 人耶稣要毁坏这地方，也要改变 摩西 所交给我们的规矩。”
ACTS|6|15|在议会里坐着的人都定睛看他，见他的面貌好像天使的面貌。
ACTS|7|1|大祭司说：“果真有这些事吗？”
ACTS|7|2|司提反 说：“诸位父老弟兄请听！从前我们的祖宗 亚伯拉罕 在 美索不达米亚 ，还没有住在 哈兰 的时候，荣耀的上帝向他显现，
ACTS|7|3|对他说：‘你要离开本地和亲族，往我所要指示你的地去。’
ACTS|7|4|他就离开 迦勒底 人的地方，住在 哈兰 。他父亲死了以后，上帝使他从那里搬到你们现在所住的地方。
ACTS|7|5|在这里上帝并没有给他产业，连立足的地方都没有，但应许要将这地赐给他和他的后裔为业，虽然那时他还没有儿子。
ACTS|7|6|上帝这样说：‘他的后裔必寄居外邦，那里的人要使他们作奴隶，苦待他们四百年。’
ACTS|7|7|上帝又说：‘但我要惩罚使他们作奴隶的那国。以后他们要出来，在这地方事奉我。’
ACTS|7|8|上帝又赐他割礼的约。于是 亚伯拉罕 生了 以撒 ，在第八日给他行了割礼；后来 以撒 生 雅各 ， 雅各 生十二位先祖。
ACTS|7|9|“先祖嫉妒 约瑟 ，把他卖到 埃及 去，上帝却与他同在，
ACTS|7|10|救他脱离一切苦难，又使他在 埃及 王法老面前蒙恩，又有智慧。法老派他作 埃及 国的宰相兼管法老的全家。
ACTS|7|11|后来全 埃及 和 迦南 遭遇饥荒和大灾难，我们的祖宗绝了粮。
ACTS|7|12|雅各 听见在 埃及 有粮，就打发我们的祖宗初次往那里去。
ACTS|7|13|第二次 约瑟 与兄弟们相认，法老才认识他的家族。
ACTS|7|14|约瑟 就打发人，请父亲 雅各 和全族七十五个人都来。
ACTS|7|15|于是 雅各 下了 埃及 ，后来他和我们的祖宗都死在那里；
ACTS|7|16|他们又被迁到 示剑 ，葬于 亚伯拉罕 在 示剑 用银子从 哈抹 子孙 买来的坟墓里。
ACTS|7|17|“当上帝应许 亚伯拉罕 的日期将到的时候， 以色列 人在 埃及 人丁兴旺，
ACTS|7|18|直到另一位不认识 约瑟 的王兴起统治 埃及 。
ACTS|7|19|他用诡计待我们的宗族，苦待我们的祖宗，强迫他们丢弃婴孩，使婴孩不能存活。
ACTS|7|20|就在那时， 摩西 生了下来，上帝看为俊美，在父亲家里被抚养了三个月。
ACTS|7|21|他被丢弃的时候，法老的女儿拾了去，当自己的儿子抚养。
ACTS|7|22|摩西 学了 埃及 人一切的学问，说话办事都有才能。
ACTS|7|23|“他到了四十岁，心中起意去看望他的弟兄 以色列 人。
ACTS|7|24|他见他们中的一个人受冤屈，就庇护他，为那被压迫的人报仇，打死了那 埃及 人。
ACTS|7|25|他以为他的弟兄们必明白上帝是藉他的手搭救他们，他们却不明白。
ACTS|7|26|第二天，他遇见有人在打架，就想劝他们和好，说：‘二位，你们是弟兄，为什么彼此欺负呢？’
ACTS|7|27|那欺负邻舍的人把他推开，说：‘谁立你作我们的领袖和审判官呢？
ACTS|7|28|难道你要杀我像昨天杀那 埃及 人一样吗？’
ACTS|7|29|摩西 听见这话就逃走了，寄居于 米甸 地，在那里生了两个儿子。
ACTS|7|30|“过了四十年，在 西奈山 的旷野，有一位天使在荆棘的火焰中向 摩西 显现。
ACTS|7|31|摩西 见了那异象，觉得很惊讶，正往前观看的时候，有主的声音说：
ACTS|7|32|‘我是你列祖的上帝，就是 亚伯拉罕 、 以撒 、 雅各 的上帝。’ 摩西 战战兢兢，不敢观看。
ACTS|7|33|主对他说：‘把你脚上的鞋脱下来，因为你所站的地方是圣地。
ACTS|7|34|我的百姓在 埃及 所受的困苦，我确实看见了；他们悲叹的声音，我也听见了。我下来要救他们。现在，你来，我要差你往 埃及 去。’
ACTS|7|35|“这 摩西 就是有人曾弃绝他说‘谁立你作我们的领袖和审判官’的，上帝却藉那在荆棘中显现的天使的手差派他作领袖，作解救者。
ACTS|7|36|这人领 以色列 人出来，在 埃及 地，在 红海 ，在旷野的四十年间行了奇事神迹。
ACTS|7|37|这人是 摩西 ，就是那曾对 以色列 人说‘上帝要从你们弟兄中给你们兴起一位先知像我’的。
ACTS|7|38|这人是那曾在旷野的会众中和 西奈山 上，与那对他说话的天使同在，又与我们祖宗同在的，他领受了活泼的圣言传给我们。
ACTS|7|39|我们的祖宗不肯听从，反弃绝他，他们的心转向 埃及 ，
ACTS|7|40|对 亚伦 说：‘你为我们造神明，在我们前面引路，因为领我们出 埃及 地的这个 摩西 ，我们不知道他遭遇了什么事。’
ACTS|7|41|那时，他们造了一个牛犊，又拿祭物献给那像，为自己手所做的工作欢跃。
ACTS|7|42|但是上帝转脸不顾，任凭他们祭拜天上的日月星辰，正如先知书上所写的： ‘ 以色列 家啊，你们四十年间在旷野， 何曾将牺牲和祭物献给我？
ACTS|7|43|你们抬着 摩洛 的帐幕 和 理番 ──你们神明的星， 就是你们所造为要敬拜的像。 因此，我要把你们迁到 巴比伦 外去。’
ACTS|7|44|“我们的祖宗在旷野，有作证的会幕，是上帝吩咐 摩西 照着他所看见的样式做的。
ACTS|7|45|这帐幕，我们的祖宗同 约书亚 相继承受了，当上帝在他们面前赶走外邦人的时候，他们把这帐幕搬进承受为业之地，直存到 大卫 的日子。
ACTS|7|46|大卫 在上帝面前蒙恩，祈求为 雅各 的家 预备居所。
ACTS|7|47|但却是 所罗门 为上帝造成殿宇。
ACTS|7|48|其实，至高者并不住人手所造的，就如先知所言：
ACTS|7|49|‘主说：天是我的宝座， 地是我的脚凳。 你们要为我造怎样的殿宇？ 哪里是我安歇的地方呢？
ACTS|7|50|这一切不都是我手所造的吗？’
ACTS|7|51|“你们这硬着颈项，心与耳未受割礼的人哪，时常抗拒圣灵！你们的祖宗怎样，你们也怎样。
ACTS|7|52|先知中有哪一个不是受你们祖宗的迫害呢？他们把预先宣告那义者要来的人杀了。如今你们成了那义者的出卖者和凶手了。
ACTS|7|53|你们领受了天使所传布的律法，竟不遵守。”
ACTS|7|54|众人听见这些话，心中极其恼怒，向 司提反 咬牙切齿。
ACTS|7|55|但 司提反 满有圣灵，定睛望天，看见上帝的荣耀，又看见耶稣站在上帝的右边，
ACTS|7|56|就说：“我看见天开了，人子站在上帝的右边。”
ACTS|7|57|众人大声喊叫，捂着耳朵，齐心冲向他，
ACTS|7|58|把他推到城外，用石头打他。作见证的人把他们的衣裳放在一个名叫 扫罗 的青年脚前。
ACTS|7|59|他们正用石头打 司提反 的时候，他呼求说：“主耶稣啊，求你接纳我的灵魂！”
ACTS|7|60|然后他跪下来，大声喊着：“主啊，不要将这罪归于他们！”说了这话，就长眠了。
ACTS|8|1|扫罗 也赞同处死他。从那一天开始， 耶路撒冷 的教会遭受到大迫害，除了使徒以外，众门徒都分散在 犹太 和 撒玛利亚 各处。
ACTS|8|2|有些虔诚的人把 司提反 埋葬了，为他大大哀哭。
ACTS|8|3|扫罗 却残害教会，挨家挨户地进去，拉着男女关在监里。
ACTS|8|4|那些分散的人往各地去传福音的道。
ACTS|8|5|腓利 下 撒玛利亚城 去 ，向当地人宣讲基督。
ACTS|8|6|众人都聚精会神，同心合意地听 腓利 所说的话，一边听他的话，一边看他所行的神迹。
ACTS|8|7|因为有许多人被污灵附着，那些污灵大声呼叫，从他们身上出来；还有许多瘫痪的、瘸腿的都得了医治。
ACTS|8|8|那城里，有极大的喜乐。
ACTS|8|9|有一个人名叫 西门 ，向来在那城里行邪术，自命为大人物，使 撒玛利亚 的居民惊奇。
ACTS|8|10|所有的人，从小到大都听从他，说：“这个人就是上帝的能力，那称为大能者的。”
ACTS|8|11|他们听从他，因他很久以来用邪术使他们惊奇。
ACTS|8|12|当他们信了 腓利 所传上帝国的福音和耶稣基督的名，连男带女都受了洗。
ACTS|8|13|西门 自己也信了；既受了洗，就常与 腓利 在一处，看见他所行的神迹和大异能，就觉得很惊奇。
ACTS|8|14|在 耶路撒冷 的使徒听见 撒玛利亚 人领受了上帝的道，就打发 彼得 和 约翰 到他们那里去。
ACTS|8|15|两个人下去，就为他们祷告，要让他们领受圣灵，
ACTS|8|16|因为圣灵还没有降在他们任何一个人身上，他们只奉主耶稣的名受了洗。
ACTS|8|17|于是使徒按手在他们头上，他们就领受了圣灵。
ACTS|8|18|西门 看见使徒一按手，就有圣灵赐下，就拿钱给使徒，
ACTS|8|19|说：“请把这权柄也给我，使我手按着谁，谁就可以领受圣灵。”
ACTS|8|20|彼得 对他说：“你的银子和你一同灭亡吧！因为你想上帝的恩赐是可以用钱买的。
ACTS|8|21|你在这道上无份无关；因为你在上帝面前心怀不正。
ACTS|8|22|你要为你这样的恶而悔改，祈求主，或者你心里的意念可得赦免。
ACTS|8|23|我看出你正在苦胆之中，被不义捆绑着。”
ACTS|8|24|西门 回答说：“请你们为我求主，使你们所说的，没有一样临到我身上。”
ACTS|8|25|使徒既作了见证，并且宣讲了主的道，就回 耶路撒冷 去，一路在 撒玛利亚 好些村庄传扬福音。
ACTS|8|26|有主的一个使者对 腓利 说：“起来！向南走，往那从 耶路撒冷 下 迦萨 的路上去。”那路是旷野。
ACTS|8|27|腓利 就起身去了。不料，有一个 埃塞俄比亚 人，是个有大权的太监，在 埃塞俄比亚 女王 甘大基 的手下总管银库，他上 耶路撒冷 去礼拜。
ACTS|8|28|回程中，他坐在车上，正念着 以赛亚 先知的书，
ACTS|8|29|圣灵对 腓利 说：“你去！靠近那车走。”
ACTS|8|30|腓利 就跑到太监那里，听见他正在念 以赛亚 先知的书，就说：“你明白你所念的吗？”
ACTS|8|31|他说：“没有人指教我，怎能明白呢？”于是他请 腓利 上车，与他同坐。
ACTS|8|32|他所念的那段经文是这样： “他像羊被牵去宰杀， 又像羔羊在剪毛的人手下无声， 他也是这样不开口。
ACTS|8|33|他卑微的时候，得不到公义的审判， 谁能述说他的身世？ 因为他的生命从地上被夺去。”
ACTS|8|34|太监回答 腓利 说：“请问，先知说这话是指谁，是指自己，还是指别人呢？”
ACTS|8|35|腓利 就开口，从这段经文开始，对他传讲耶稣的福音。
ACTS|8|36|二人正沿路往前走，到了有水的地方，太监说：“看哪！这里有水，有什么能阻止我受洗呢？”
ACTS|8|37|
ACTS|8|38|于是他吩咐把车停下来， 腓利 和太监二人一同下到水里， 腓利 就给他施洗。
ACTS|8|39|他们从水里上来，主的灵把 腓利 提了去，太监再也看不见他了，就欢欢喜喜地上路。
ACTS|8|40|后来有人在 亚锁都 遇见 腓利 ；他走遍那地方，在各城宣扬福音，一直到 凯撒利亚 。
ACTS|9|1|扫罗 不断用威吓凶悍的口气向主的门徒说话。他去见大祭司，
ACTS|9|2|要求发信给 大马士革 的各会堂，若是找着信奉这道的人，无论男女，都准他捆绑带到 耶路撒冷 。
ACTS|9|3|扫罗 在途中，将到 大马士革 的时候，忽然有一道光从天上下来，四面照射着他，
ACTS|9|4|他就仆倒在地，听见有声音对他说：“ 扫罗 ！ 扫罗 ！你为什么迫害我？”
ACTS|9|5|他说：“主啊！你是谁？”主说：“我就是你所迫害的耶稣。
ACTS|9|6|起来！进城去，你应该做的事，必有人告诉你。”
ACTS|9|7|同行的人站在那里，说不出话来，因为他们听见声音，却看不见人。
ACTS|9|8|扫罗 从地上起来，睁开眼睛，竟不能看见什么。有人拉他的手，领他进了 大马士革 。
ACTS|9|9|他三天什么都看不见，也不吃也不喝。
ACTS|9|10|那时，在 大马士革 有一个门徒，名叫 亚拿尼亚 。主在异象中对他说：“ 亚拿尼亚 ！”他说：“主啊，我在这里。”
ACTS|9|11|主对他说：“起来！往那叫 直街 的路去，在 犹大 的家里，去找一个 大数 人，名叫 扫罗 ；他正在祷告，
ACTS|9|12|在异象中 看见了一个人，名叫 亚拿尼亚 ，进来为他按手，让他能再看得见。”
ACTS|9|13|亚拿尼亚 回答：“主啊，我听见许多人讲到这个人，说他怎样在 耶路撒冷 多多苦待你的圣徒，
ACTS|9|14|并且他在这里有从祭司长得来的权柄，要捆绑一切求告你名的人。”
ACTS|9|15|主对他说：“你只管去。他是我所拣选的器皿，要在外邦人、君王和 以色列 人面前宣扬我的名。
ACTS|9|16|我也要指示他，为我的名必须受许多的苦难。”
ACTS|9|17|亚拿尼亚 就去了，进入那家，把手按在 扫罗 身上，说：“ 扫罗 弟兄，在你来的路上向你显现的主，就是耶稣，打发我来，叫你能再看得见，又被圣灵充满。”
ACTS|9|18|扫罗 的眼睛上立刻好像有鳞一般的东西掉下来，他就能再看得见，于是他起来，受了洗，
ACTS|9|19|吃过饭体力就恢复了。 扫罗 和 大马士革 的门徒一起住了些日子，
ACTS|9|20|立刻在各会堂里传扬耶稣，说他是上帝的儿子。
ACTS|9|21|凡听见的人都很惊奇，说：“在 耶路撒冷 残害求告这名的不就是这个人吗？他不是到这里来要捆绑他们，带到祭司长那里去吗？”
ACTS|9|22|但 扫罗 越发有能力，驳倒住在 大马士革 的 犹太 人，证明耶稣是基督。
ACTS|9|23|过了好些日子， 犹太 人商议要杀 扫罗 ，
ACTS|9|24|但他们的计谋被 扫罗 知道了。他们昼夜在城门守候着要杀他。
ACTS|9|25|他的门徒就在夜间用筐子把他从城墙上缒了下去。
ACTS|9|26|扫罗 到了 耶路撒冷 ，想与门徒结交，大家却都怕他，不信他是门徒。
ACTS|9|27|只有 巴拿巴 接待他，领他去见使徒，把他在路上怎么看见主，主怎么向他说话，他在 大马士革 怎么奉耶稣的名放胆传道，都述说出来。
ACTS|9|28|于是 扫罗 在 耶路撒冷 同门徒出入来往，奉主的名放胆传道，
ACTS|9|29|并和说 希腊 话的 犹太 人讲论辩驳，他们却想法子要杀他。
ACTS|9|30|弟兄们知道了，就带他下 凯撒利亚 ，送他往 大数 去。
ACTS|9|31|那时， 犹太 、 加利利 、 撒玛利亚 各处的教会都得平安，建立起来，凡事敬畏主，蒙圣灵的安慰，人数逐渐增多。
ACTS|9|32|彼得 在众信徒中到处奔波的时候，也到了住在 吕大 的圣徒那里。
ACTS|9|33|他在那里遇见一个人，名叫 以尼雅 ，得了瘫痪，在褥子上躺了八年。
ACTS|9|34|彼得 对他说：“ 以尼雅 ，耶稣基督医好你了，起来！整理你的褥子吧。”他立刻就起来了。
ACTS|9|35|凡住 吕大 和 沙仑 的人都看见了他，就归向主。
ACTS|9|36|在 约帕 有一个女门徒，名叫 大比大 ，翻出来的意思是 多加 ；她广行善事，多施周济。
ACTS|9|37|当时，她患病死了，有人把她清洗后，停在楼上。
ACTS|9|38|吕大 原与 约帕 相近；门徒听见 彼得 在那里，就派两个人去见他，央求他说：“请快到我们那里去，不要耽延。”
ACTS|9|39|彼得 就起身和他们同去。他到了，就有人领他上楼。众寡妇都站在 彼得 旁边哭，拿 多加 与她们同在时所做的内衣外衣给他看。
ACTS|9|40|彼得 叫她们都出去，然后跪下祷告，转身对着尸体说：“ 大比大 ，起来！”她就睁开眼睛，看见 彼得 ，就坐了起来。
ACTS|9|41|彼得 伸手扶她起来，叫那些圣徒和寡妇都进来，把 多加 活活地交给他们。
ACTS|9|42|这事传遍了 约帕 ，就有许多人信了主。
ACTS|9|43|此后， 彼得 在 约帕 一个皮革匠 西门 的家里住了好些日子。
ACTS|10|1|在 凯撒利亚 有一个人名叫 哥尼流 ，是 意大利 营的百夫长。
ACTS|10|2|他是个虔诚人，他和全家都敬畏上帝。他多多周济百姓，常常向上帝祷告。
ACTS|10|3|有一天，约在下午三点钟，他在异象中清楚看见上帝的一个使者进来，到他那里，对他说：“ 哥尼流 。”
ACTS|10|4|哥尼流 定睛看他，惊惶地说：“主啊，什么事？”天使对他说：“你的祷告和你的周济已达到上帝面前，蒙记念了。
ACTS|10|5|现在你要派人往 约帕 去，请一位称为 彼得 的 西门 来。
ACTS|10|6|他住在一个皮革匠 西门 的家里，房子就在海边。”
ACTS|10|7|向他说话的天使离开后， 哥尼流 叫了两个仆人和常伺候他的一个虔诚的兵来，
ACTS|10|8|把一切的事都讲给他们听，然后就派他们往 约帕 去。
ACTS|10|9|第二天，他们走路将近那城，约在正午， 彼得 上房顶去祷告。
ACTS|10|10|他觉得饿了，想要吃。那家的人正预备饭的时候， 彼得 魂游象外，
ACTS|10|11|看见天开了，有一块好像大布的东西降下，四角 吊着缒在地上，
ACTS|10|12|里面有地上各样四脚的走兽、爬虫和天上的飞鸟。
ACTS|10|13|又有声音对他说：“ 彼得 ，起来！宰了吃。”
ACTS|10|14|彼得 却说：“主啊，绝对不可！凡污俗和不洁净的东西，我从来没有吃过。”
ACTS|10|15|第二次有声音再对他说：“上帝所洁净的，你不可当作污俗的。”
ACTS|10|16|这样一连三次，那东西随即收回天上去了。
ACTS|10|17|正当 彼得 心里困惑，不知所看见的异象是什么意思时， 哥尼流 所差来的人已经找到了 西门 的家，站在门外，
ACTS|10|18|喊着问有没有一位称为 彼得 的 西门 住在这里。
ACTS|10|19|彼得 还在思考那异象的时候，圣灵对他说：“有三个人来找你。
ACTS|10|20|起来，下去，跟他们同去，不要疑惑，因为是我差他们来的。”
ACTS|10|21|于是 彼得 下去见那些人，说：“我就是你们要找的人，你们是为了什么缘故在这里？”
ACTS|10|22|他们说：“百夫长 哥尼流 是个义人，敬畏上帝，为 犹太 全民族所称赞。他蒙一位圣天使指示，叫他请你到他家里去，要听你讲话。”
ACTS|10|23|彼得 就请他们进去住宿。 次日，他起身和他们同去，还有 约帕 的几个弟兄跟他一起去。
ACTS|10|24|又次日，他 进入 凯撒利亚 ， 哥尼流 已经请了他的亲朋好友在等候他们。
ACTS|10|25|彼得 一进去， 哥尼流 就迎接他，俯伏在他脚前拜他。
ACTS|10|26|但是 彼得 拉他起来，说：“你起来，我自己也不过是人。”
ACTS|10|27|彼得 和他一边说话一边进去，见有好些人聚集，
ACTS|10|28|就对他们说：“你们知道， 犹太 人和别国的人结交来往本是不合规矩的，但上帝已经指示我，无论什么人都不可看作污俗或不洁净的。
ACTS|10|29|所以，我一被邀请，没有推辞就来了。现在请问，你们为什么叫我来呢？”
ACTS|10|30|哥尼流 说：“四天前，这个时候，我在家中守着下午三点钟的祷告，忽然有一个人穿着明亮的衣裳站在我面前，
ACTS|10|31|说：‘ 哥尼流 ，你的祷告已蒙垂听，你的周济在上帝面前已蒙记念了。
ACTS|10|32|你要派人往 约帕 去，请那称为 彼得 的 西门 来，他住在海边一个皮革匠 西门 的家里。’
ACTS|10|33|所以我立刻派人去请你。你来了真好。现在我们都在上帝面前，要听主 吩咐你的一切话。”
ACTS|10|34|彼得 开口说：“我真的看出上帝是不偏待人的。
ACTS|10|35|不但如此，在各国中那敬畏他而行义的人都为他所悦纳。
ACTS|10|36|上帝藉着耶稣基督—他是万有的主—传和平的福音，把这道传给 以色列 人。
ACTS|10|37|这话在 约翰 传扬洗礼以后，从 加利利 起，传遍了 犹太 。上帝怎样以圣灵和能力膏了 拿撒勒 人耶稣，这都是你们知道的。他到处奔波，行善事，医好凡被魔鬼压制的人，因为上帝与他同在。
ACTS|10|38|
ACTS|10|39|他在 犹太 人之地和 耶路撒冷 所行的一切事，有我们作见证人。他们竟把他挂在木头上杀了。
ACTS|10|40|第三天，上帝使他复活，使他显现出来；
ACTS|10|41|不是显现给所有的人看，而是显现给上帝预先所拣选为他作见证的人看，就是我们这些在他从死人中复活以后和他同吃同喝的人。
ACTS|10|42|他吩咐我们传道给众人，证明他是上帝所立定，要作审判活人、死人的审判者。
ACTS|10|43|众先知也为这人作见证：凡信他的人，必藉着他的名得蒙赦罪。”
ACTS|10|44|彼得 还在说这些话的时候，圣灵降在一切听道的人身上。
ACTS|10|45|那些奉割礼的信徒和 彼得 同来，见圣灵的恩赐也浇在外邦人身上，就都惊奇；
ACTS|10|46|因听见他们说方言 ，称赞上帝为大。于是 彼得 回答：
ACTS|10|47|“这些人既受了圣灵，跟我们一样，谁能阻止用水给他们施洗呢？”
ACTS|10|48|他就吩咐奉耶稣基督的名给他们施洗。于是他们请 彼得 住了几天。
ACTS|11|1|使徒和在 犹太 的众弟兄听到外邦人也领受了上帝的道。
ACTS|11|2|等到 彼得 上了 耶路撒冷 ，那些奉割礼的信徒和他争辩，
ACTS|11|3|说：“你竟进入未受割礼之人当中，和他们一同吃饭！”
ACTS|11|4|彼得 就开始把这事逐一向他们解释，说：
ACTS|11|5|“我在 约帕城 里祷告的时候，魂游象外，看见异象，有一块好像大布的东西降下，四角吊着从天缒下，直来到我跟前。
ACTS|11|6|我定睛观看，见内中有地上四脚的牲畜、野兽、爬虫和天上的飞鸟。
ACTS|11|7|我还听见有声音对我说：‘ 彼得 ，起来！宰了吃。’
ACTS|11|8|我说：‘主啊，绝对不可！凡污俗或不洁净的东西从来没有进过我的口。’
ACTS|11|9|第二次，有声音从天上回答：‘上帝所洁净的，你不可当作污俗的。’
ACTS|11|10|这样一连三次，然后一切就都收回天上去了。
ACTS|11|11|正当那时，有三个从 凯撒利亚 差来见我的人，站在我们 所住的屋子门前。
ACTS|11|12|圣灵吩咐我和他们同去，不要疑惑，还有这六位弟兄也跟我一起去，我们进了那人的家。
ACTS|11|13|那人就告诉我们，他如何看见一位天使站在他家里，说：‘你派人往 约帕 去，请那称为 彼得 的 西门 来，
ACTS|11|14|他有话要告诉你，因这些话你和你的全家都可以得救。’
ACTS|11|15|我一开始讲话，圣灵就降在他们身上，正像当初降在我们身上一样。
ACTS|11|16|我就想起主的话如何说：‘ 约翰 用水施洗，但你们要在圣灵里受洗。’
ACTS|11|17|既然上帝给他们恩赐，像在我们信主耶稣基督的时候给了我们一样，我是谁，能拦阻上帝吗？”
ACTS|11|18|众人听见这些话，就不说话了，只归荣耀给上帝，说：“这样看来，上帝也赐恩给外邦人，使他们悔改得生命了。”
ACTS|11|19|那些因 司提反 的事遭患难而四处分散的门徒，直走到 腓尼基 、 塞浦路斯 和 安提阿 。他们不向别人讲道，只向 犹太 人讲。
ACTS|11|20|但内中有 塞浦路斯 和 古利奈 人，他们到了 安提阿 也向 希腊 人传讲主耶稣的福音 。
ACTS|11|21|主的手与他们同在，信而归主的人数很多。
ACTS|11|22|这风声传到 耶路撒冷 教会的人耳中，他们就打发 巴拿巴 到 安提阿 去。
ACTS|11|23|他到了那里，看见上帝所赐的恩就欢喜，劝勉众人要立定心志，恒久靠主。
ACTS|11|24|这 巴拿巴 原是个好人，满有圣灵和信心，于是有许多人归服了主。
ACTS|11|25|他又往 大数 去找 扫罗 ，
ACTS|11|26|找着了，就带他到 安提阿 去。他们足有一年和教会一同聚集，教导了许多人。门徒称为“基督徒”是从 安提阿 开始的。
ACTS|11|27|当那些日子，有几位先知从 耶路撒冷 下到 安提阿 。
ACTS|11|28|内中有一位，名叫 亚迦布 ，站起来，藉着圣灵指示普天下将有大饥荒；这事在 克劳第 年间果然实现了。
ACTS|11|29|于是门徒决定，照各人的力量捐钱，送去供给住在 犹太 的弟兄。
ACTS|11|30|他们就这样做了，托 巴拿巴 和 扫罗 的手送到众长老那里。
ACTS|12|1|约在那时候， 希律 王下手苦待教会中的一些人，
ACTS|12|2|用刀杀了 约翰 的哥哥 雅各 。
ACTS|12|3|他见 犹太 人喜欢这事，也去拿住 彼得 。那时候正是除酵节期间。
ACTS|12|4|希律 捉了 彼得 ，押在监里，交给四班士兵看守，每班四个人，企图要在逾越节后把他提出来，当着百姓办他。
ACTS|12|5|于是 彼得 被囚在监里，教会却为他切切祷告上帝。
ACTS|12|6|希律 将要提他出来的前一夜， 彼得 被两条铁链锁着，睡在两个士兵当中；门前还有警卫看守。
ACTS|12|7|忽然，有主的一个使者显现，牢房里有光照耀；天使拍 彼得 的肋旁，叫醒了他，说：“快起来！”铁链就从他手上脱落下来。
ACTS|12|8|天使对他说：“束上腰带，穿上鞋子。”他就照着做了。天使又对他说：“披上外衣，跟我来。”
ACTS|12|9|彼得 就出来跟着他走，不知道天使所做是真的，以为见了异象。
ACTS|12|10|他们经过了第一层和第二层监牢，就来到往城内的铁门，那门就自动给他们开了。他们出来，走过一条街，忽然天使离开他去了。
ACTS|12|11|彼得 清醒过来，说：“现在我真知道主差遣他的使者，救我脱离 希律 的手，和 犹太 人所期待的一切。”
ACTS|12|12|他明白了，就到那称为 马可 的 约翰 的母亲 马利亚 家去，在那里已有好些人聚集祷告。
ACTS|12|13|彼得 敲外门时，有一个使女，名叫 罗大 ，出来应门，
ACTS|12|14|认出是 彼得 的声音，欢喜得顾不了开门，就跑进去报信，说 彼得 站在门外。
ACTS|12|15|他们对她说：“你疯了！”使女坚持真有其事。他们说：“那是他的天使。”
ACTS|12|16|彼得 不停地敲门；他们开了门，一见是他，就很惊奇。
ACTS|12|17|彼得 做个手势，要他们不作声，就告诉他们主怎样领他出监；又说：“你们要把这些事告诉 雅各 和众弟兄。”然后，他离开往别处去了。
ACTS|12|18|到了天亮，士兵中起了不少骚动，不知道 彼得 到哪里去了。
ACTS|12|19|希律 找他，找不着，就审问警卫，下令带走他们处死。后来 希律 离开 犹太 ，下 凯撒利亚 去，住在那里。
ACTS|12|20|希律 向 推罗 和 西顿 的人发怒。他们那一带地方是从王的土地供应粮食的，因此就托了王的内侍大臣 伯拉斯都 的情，一心来求和。
ACTS|12|21|希律 在所定的日子，穿上朝服，坐在位上，对他们演讲。
ACTS|12|22|民众一直喊着：“这是神明的声音，不是人的声音。”
ACTS|12|23|希律 不归荣耀给上帝，所以主的使者立刻击打他，他被虫咬，就断了气。
ACTS|12|24|上帝的道日见兴旺，越发广传。
ACTS|12|25|巴拿巴 和 扫罗 完成了供给的事，就回到 耶路撒冷 ，带著称为 马可 的 约翰 同去。
ACTS|13|1|在 安提阿 的教会中，有几位先知和教师，就是 巴拿巴 和称为 尼结 的 西面 、 古利奈 人 路求 ，与 希律 分封王一起长大的 马念 ，和 扫罗 。
ACTS|13|2|他们在事奉主和禁食的时候，圣灵说：“要为我分派 巴拿巴 和 扫罗 去做我召他们做的工作。”
ACTS|13|3|于是他们禁食祷告后，给 巴拿巴 和 扫罗 按手，然后派遣他们走了。
ACTS|13|4|他们既蒙圣灵差遣，就下到 西流基 ，从那里坐船往 塞浦路斯 去，
ACTS|13|5|到了 撒拉米 ，就在 犹太 人各会堂里宣讲上帝的道，也有 约翰 作他们的帮手。
ACTS|13|6|他们走遍全岛，直到 帕弗 ，在那里遇见一个术士— 犹太 人的假先知，名叫 巴耶稣 。
ACTS|13|7|这人常和 士求．保罗 省长在一起。 士求．保罗 是个通达人，他请 巴拿巴 和 扫罗 来，要听上帝的道。
ACTS|13|8|只是术士 以吕马 (他的名字翻出来就是行法术的意思)敌对使徒，设法使省长远离这信仰。
ACTS|13|9|扫罗 ，又名 保罗 ，被圣灵充满，定睛看他，
ACTS|13|10|说：“你这充满各样诡诈奸恶，魔鬼的儿子，一切正义的仇敌，你还不停止扭曲主的正道吗？
ACTS|13|11|现在你看，主的手临到你身上，你会瞎眼，暂时看不见日光。”立刻迷濛和黑暗笼罩着他，他到处摸索，求人拉着手领他。
ACTS|13|12|省长看见所发生的事就信了，因对主的教导感到惊奇。
ACTS|13|13|保罗 和他的同伴从 帕弗 开船，来到 旁非利亚 的 别加 ， 约翰 却离开他们，回 耶路撒冷 去了。
ACTS|13|14|他们从 别加 往前行，来到 彼西底 的 安提阿 。在安息日，他们进了会堂就坐下。
ACTS|13|15|在读完了律法和先知的书，会堂主管们叫人过去，对他们说：“二位弟兄，你们若有什么劝勉众人的话，请说。”
ACTS|13|16|保罗 就站起来，做个手势，说：“诸位 以色列 人和一切敬畏上帝的人，请听。
ACTS|13|17|这 以色列 民的上帝拣选了我们的祖宗，当百姓寄居 埃及 的时候抬举他们，用大能的手领他们从那地出来。
ACTS|13|18|他在旷野容忍 他们，约有四十年。
ACTS|13|19|他消灭了 迦南 地七族的人后，把那地分给他们为业，
ACTS|13|20|约有四百五十年。此后 ，他给他们设立士师，直到 撒母耳 先知的时候。
ACTS|13|21|从那时起，他们要求立一个王，上帝就将 便雅悯 支派中 基士 的儿子 扫罗 给他们作王，共四十年。
ACTS|13|22|他废了 扫罗 之后，就兴起 大卫 作他们的王，又为他作见证说：‘我寻得 耶西 的儿子 大卫 ，他是合我心意的人，他要遵行我一切的旨意。’
ACTS|13|23|从这人的后裔中，上帝已经照着所应许的为 以色列 人兴起一位救主，就是耶稣。
ACTS|13|24|在他没有出来以前， 约翰 已向 以色列 全民宣讲悔改的洗礼。
ACTS|13|25|约翰 快走完他的人生路程时，说：‘你们以为我是谁？我不是 ；但是有一位在我以后来的，我就是解他脚上的鞋带也不配。’
ACTS|13|26|“诸位弟兄— 亚伯拉罕 的子孙和你们中间敬畏上帝的人哪，这救世的道是传给我们的。
ACTS|13|27|耶路撒冷 的居民和他们的官长，因为不认识这基督，也不明白每安息日所读的先知的书，把他定了死罪，正应验了先知的预言。
ACTS|13|28|虽然他们查不出他有该死的罪状，还是要求 彼拉多 把他杀了。
ACTS|13|29|他们既实现了经上指着他所记的一切话，就从木头上把他取下来，放在坟墓里。
ACTS|13|30|上帝却使他从死人中复活。
ACTS|13|31|有许多日子，他向那些从 加利利 同他上 耶路撒冷 的人显现，这些人如今在民间成为他的见证人。
ACTS|13|32|我们报好信息给你们，就是那应许祖宗的话，
ACTS|13|33|上帝已经向我们这些作他们儿女的 应验，使耶稣复活了。正如《诗篇》第二篇上记着： ‘你是我的儿子， 我今日生了你。’
ACTS|13|34|论到上帝使他从死人中复活，不再归于朽坏，他曾这样说： ‘我必将所应许 大卫 那圣洁、 可靠的恩典赐给你们。’
ACTS|13|35|所以他也在另一篇说： ‘你必不让你的圣者见朽坏。’
ACTS|13|36|大卫 在世的时候，遵行了上帝的旨意就长眠了 ，归到他祖宗那里，已见朽坏；
ACTS|13|37|惟独上帝使他复活的那一位，他并未见朽坏。
ACTS|13|38|所以弟兄们，你们当知道：赦罪的道是由这人传给你们的，
ACTS|13|39|你们靠 摩西 的律法在不得称义的一切事上，每一个信靠这位耶稣的都得称义了。
ACTS|13|40|所以，你们要小心，免得先知书上所说的临到你们：
ACTS|13|41|‘要观看，你们这些藐视的人， 要惊讶，要灭亡， 因为在你们的日子，我行一件事， 虽有人告诉你们，你们总是不信。’”
ACTS|13|42|他们走出会堂的时候，众人请他们在下一个安息日再讲这些话给他们听。
ACTS|13|43|散会以后，有许多 犹太 人和敬虔的皈依 犹太 教的人跟从了 保罗 和 巴拿巴 。二人对他们讲话，劝他们务要恒久倚靠上帝的恩典。
ACTS|13|44|到下一个安息日，全城的人几乎都聚集起来，要听主的道 。
ACTS|13|45|但 犹太 人看见这么多的人，就满心嫉妒，辩驳 保罗 所说的话，并且毁谤他。
ACTS|13|46|于是 保罗 和 巴拿巴 放胆说：“上帝的道本应先传给你们；只因你们弃绝这道，断定自己不配得永生，我们就转向外邦人。
ACTS|13|47|因为主曾这样吩咐我们： ‘我已经立你作万邦之光， 使你施行我的救恩，直到地极。’”
ACTS|13|48|外邦人听见这话很欢喜，赞美主的道，凡被指定得永生的人都信了。
ACTS|13|49|于是主的道传遍了那一带地方。
ACTS|13|50|但 犹太 人挑唆虔敬尊贵的妇女和城内有名望的人，迫害 保罗 和 巴拿巴 ，把他们赶出境外。
ACTS|13|51|二人对着众人跺掉脚上的尘土，然后往 以哥念 去了。
ACTS|13|52|门徒满心喜乐，又被圣灵充满。
ACTS|14|1|同样的事也发生在 以哥念 。 保罗 和 巴拿巴 进了 犹太 人的会堂，在那里讲道，所以有很多 犹太 人和 希腊 人都信了。
ACTS|14|2|但那不顺从的 犹太 人煽动外邦人，使他们心里仇恨弟兄。
ACTS|14|3|二人在那里住了好些日子，倚靠主放胆讲道，主藉他们的手施行神迹奇事，证明他恩惠的道。
ACTS|14|4|城里的众人却分裂了：有依附 犹太 人的，有依附使徒的。
ACTS|14|5|那时，外邦人、 犹太 人和他们的官长，一齐拥上来，要凌辱使徒，用石头打他们。
ACTS|14|6|使徒知道了，就逃到 吕高尼 的 路司得 和 特庇 两个城，以及周围地方去，
ACTS|14|7|在那里继续传福音。
ACTS|14|8|路司得城 里有一个两脚无力的人，他从母腹里就是瘸腿的，老是坐着，从来没有走过。
ACTS|14|9|他听 保罗 讲道； 保罗 定睛看他，见他有信心，可得痊愈，
ACTS|14|10|就大声说：“起来！两脚站直。”那人就跳起来，开始行走。
ACTS|14|11|众人看见 保罗 所做的事，就用 吕高尼 话大声说：“有神明藉着人形降临在我们中间了。”
ACTS|14|12|于是他们称 巴拿巴 为 宙斯 ，称 保罗 为 希耳米 ，因为他总是带头说话。
ACTS|14|13|城外有 宙斯 庙的祭司牵着牛，拿着花环，来到门前，要同众人一起献祭。
ACTS|14|14|巴拿巴 和 保罗 二位使徒听见，就撕开衣裳，跳进众人中间，喊着：
ACTS|14|15|“诸位，为什么做这些事呢？我们也是人，性情和你们一样。我们传福音给你们，是要你们离弃这些虚妄的事，归向那创造天、地、海和其中万物的永生的上帝。
ACTS|14|16|他在从前的世代，任凭万国各行其道；
ACTS|14|17|然而他未尝不为自己留下证据来，就如常行善事，从天降雨，赏赐丰年，使你们饮食饱足，满心喜乐。”
ACTS|14|18|二人说了这些话，总算拦住众人不献祭给他们。
ACTS|14|19|但有些 犹太 人，从 安提阿 和 以哥念 来，挑唆众人，并且用石头打 保罗 ，以为他死了，就把他拖到城外。
ACTS|14|20|当门徒围着他的时候，他站了起来，走进城去。第二天， 保罗 同 巴拿巴 往 特庇 去。
ACTS|14|21|保罗 和 巴拿巴 对那城里的人传了福音，使好些人成为门徒后，又回 路司得 、 以哥念 、 安提阿 去，
ACTS|14|22|坚固门徒的心，劝他们持守他们的信仰，说：“我们进入上帝的国，必须经历许多艰难。”
ACTS|14|23|二人在各教会中选立了长老，禁食祷告后，把他们交托给他们所信的主。
ACTS|14|24|二人经过 彼西底 来到 旁非利亚 ，
ACTS|14|25|在 别加 讲了道，就下 亚大利 去，
ACTS|14|26|从那里坐船回 安提阿 去。当初，众人就在这地方，把他们交托在上帝的恩典中，要完成现在所做的工。
ACTS|14|27|他们一到那里，就聚集了会众，述说上帝藉他们所行的一切事，并且上帝怎样为外邦人开了信道的门。
ACTS|14|28|二人在那里同门徒住了一段日子。
ACTS|15|1|有几个人从 犹太 下来，教导弟兄们说：“你们若不按照 摩西 的规矩受割礼，不能得救。”
ACTS|15|2|保罗 和 巴拿巴 跟他们发生了激烈的争执和辩论；大家就决定指派 保罗 、 巴拿巴 和本会的几个人，为所辩论的事上 耶路撒冷 去见使徒和长老。
ACTS|15|3|于是教会为他们送行。他们经过 腓尼基 、 撒玛利亚 ，沿途叙说外邦人归主的事，使众弟兄都非常欢喜。
ACTS|15|4|他们到了 耶路撒冷 ，教会、使徒和长老都接待他们，他们就述说上帝同他们所做的一切事。
ACTS|15|5|惟有几个法利赛派的信徒起来，说：“必须给外邦人行割礼，吩咐他们遵守 摩西 的律法。”
ACTS|15|6|使徒和长老聚集商议这事。
ACTS|15|7|辩论了许久后， 彼得 站起来，对他们说：“诸位弟兄，你们知道上帝早已在你们中间拣选了我，让外邦人从我口中得听福音之道，而且相信。
ACTS|15|8|知道人心的上帝也为他们作了见证，赐圣灵给他们，正如给我们一样；
ACTS|15|9|又藉着信洁净了他们的心，他们和我们之间并没有什么分别。
ACTS|15|10|现在你们为什么试探上帝，要把我们祖宗和我们所不能负的轭放在门徒的颈项上呢？
ACTS|15|11|相反地，我们相信，我们得救是因主耶稣的恩典，和他们一样。”
ACTS|15|12|众人都默默无声，听 巴拿巴 和 保罗 述说上帝藉着他们在外邦人中所行的神迹和奇事。
ACTS|15|13|他们讲完了， 雅各 回答说：“诸位弟兄，请听我说。
ACTS|15|14|刚才 西门 述说上帝当初怎样眷顾外邦人，从他们中间选取人民归于自己的名下；
ACTS|15|15|众先知的话也与这意思相符合。
ACTS|15|16|正如经上所写的： ‘此后，我要回来， 重新修造 大卫 倒塌了的帐幕， 从废墟中重新修造， 把它建立起来，
ACTS|15|17|使剩余的人， 就是凡称我名的外邦人， 都寻求主。 这话是自古以来显明这些事的主说的。’
ACTS|15|18|
ACTS|15|19|所以，我的意见是不可难为那归向上帝的外邦人；
ACTS|15|20|但是要写信吩咐他们禁戒偶像所玷污的东西、血和勒死的牲畜 ，禁戒淫乱。
ACTS|15|21|因为历代以来， 摩西 的书在各城都有人宣讲，每逢安息日，也在会堂里诵读。”
ACTS|15|22|那时，使徒、长老和全教会认为应从他们中间拣选人，差他们和 保罗 、 巴拿巴 一同到 安提阿 去，所拣选的就是称为 巴撒巴 的 犹大 和 西拉 。这二人在弟兄中是领袖。
ACTS|15|23|他们带去的信说：“使徒和作长老的弟兄们向 安提阿 、 叙利亚 、 基利家 外邦众弟兄问安。
ACTS|15|24|我们听说，有几个人从我们这里出去 ，用一些话骚扰你们，使你们的心困惑， 其实我们并没有吩咐他们。
ACTS|15|25|我们认为，既然我们同心定意，就拣选几个人，派他们同我们所亲爱的 巴拿巴 和 保罗 到你们那里去。
ACTS|15|26|这二人曾为我主耶稣基督的名不顾自己的性命。
ACTS|15|27|所以我们派 犹大 和 西拉 去，他们也会亲口述说这些事。
ACTS|15|28|因为圣灵和我们决定除了这几件重要的事，不将别的重担放在你们身上，
ACTS|15|29|就是禁戒偶像所玷污的东西、血和勒死的牲畜，禁戒淫乱。这几件你们若能自己禁戒就好了。祝你们安康！”
ACTS|15|30|他们既奉了差遣就下 安提阿 去，聚集会众，把书信交给他们。
ACTS|15|31|众人念了，因为信上鼓励的话而感到欣慰。
ACTS|15|32|犹大 和 西拉 自己也是先知，就用许多话劝勉弟兄，坚固他们。
ACTS|15|33|二人住了些日子，弟兄们打发他们平平安安地回到差遣他们的人那里去。
ACTS|15|34|
ACTS|15|35|但 保罗 和 巴拿巴 仍留在 安提阿 ，和许多别的人一同教导，并传扬主的道。
ACTS|15|36|过了些日子， 保罗 对 巴拿巴 说：“让我们回到从前宣扬主道的各城，看看弟兄们的情况如何。”
ACTS|15|37|巴拿巴 有意要带称为 马可 的 约翰 同去；
ACTS|15|38|但 保罗 认为不宜带他去，因为 马可 从前在 旁非利亚 离开他们，不和他们一起工作。
ACTS|15|39|于是二人起了争执，甚至彼此分手。 巴拿巴 带着 马可 ，坐船往 塞浦路斯 去；
ACTS|15|40|保罗 则拣选了 西拉 ，也出发了，蒙弟兄们把他交于主的恩典中。
ACTS|15|41|他就走遍了 叙利亚 、 基利家 ，坚固众教会。
ACTS|16|1|后来， 保罗 来到 特庇 ，又到 路司得 。在那里有一个门徒，名叫 提摩太 ，是信主的 犹太 妇人的儿子，他父亲却是 希腊 人。
ACTS|16|2|路司得 和 以哥念 的弟兄都称赞他。
ACTS|16|3|保罗 要带他同去，只因那些地方的 犹太 人都知道他父亲是 希腊 人，就给他行了割礼。
ACTS|16|4|他们经过各城，把 耶路撒冷 使徒和长老所决定的规条交给门徒遵守。
ACTS|16|5|于是众教会信心越发坚固，人数天天增加。
ACTS|16|6|因为圣灵禁止他们在 亚细亚 讲道，他们就经过 弗吕家 、 加拉太 一带地方。
ACTS|16|7|到了 每西亚 的边界，他们想要往 庇推尼 去，耶稣的灵却不许。
ACTS|16|8|他们就越过 每西亚 ，下 特罗亚 去。
ACTS|16|9|夜间，有异象向 保罗 显现。有一个 马其顿 人站着求他说：“请你过来，到 马其顿 来帮助我们！”
ACTS|16|10|保罗 既看见这异象，我们就立即设法往 马其顿 去，认为上帝呼召我们传福音给那里的人。
ACTS|16|11|我们从 特罗亚 开船，直行驶到 撒摩特喇 ，第二天到了 尼亚坡里 ；
ACTS|16|12|从那里来到 腓立比 ，就是 马其顿 这一带的一个重要城市 ，也是 罗马 的驻防城。我们在这城里住了几天。
ACTS|16|13|在安息日，我们出城门，到了河边，知道那里有一个祷告的地方 ，我们就坐下来对那些聚会的妇女讲道。
ACTS|16|14|有一个卖紫色布的妇人，名叫 吕底亚 ，是 推雅推喇城 的人，素来敬拜上帝。她在听着，主就开导她的心，使她留心听 保罗 所讲的话。
ACTS|16|15|她和她一家都领了洗，就求我们说：“你们若以为我是真心信主的 ，请到我家里来住。”于是她坚决请我们留下。
ACTS|16|16|后来，我们往那祷告的地方去时，有一个被占卜的灵附身的使女迎面走来，她使用法术使她的主人们发了大财。
ACTS|16|17|她跟随 保罗 和我们，喊着说：“这些人是至高上帝的仆人，对你们传讲救人的道路。”
ACTS|16|18|她一连好几天这样喊叫， 保罗 就心中厌烦，转身对那灵说：“我奉耶稣基督的名吩咐你从她身上出来！”那灵立刻出来了。
ACTS|16|19|使女的主人们见发财的指望没有了，就揪住 保罗 和 西拉 ，拉他们到市上去见官；
ACTS|16|20|又带他们到行政官长们面前，说：“这些骚扰我们城的，他们是 犹太 人，
ACTS|16|21|竟传布我们 罗马 人所不可接受、不可遵守的规矩。”
ACTS|16|22|群众就一齐起来攻击他们。官长们吩咐撕开他们的衣裳，用棍子打；
ACTS|16|23|打了许多棍，就把他们下在监里，嘱咐狱警严紧看守。
ACTS|16|24|狱警领了这样的命令，就把他们下在内监，两脚拴在木架上。
ACTS|16|25|约在半夜， 保罗 和 西拉 正在祷告，唱诗赞美上帝，众囚犯也侧耳听着的时候，
ACTS|16|26|忽然，地大震动，甚至监牢的地基都摇动了，监门立刻全开，众囚犯的锁链也都解开了。
ACTS|16|27|狱警一醒，看见监门全开，以为囚犯已经逃走，就拔刀要自杀。
ACTS|16|28|保罗 大声呼叫：“不要伤害自己！我们都在这里。”
ACTS|16|29|狱警叫人拿灯来，就冲进去，战战兢兢地俯伏在 保罗 和 西拉 面前。
ACTS|16|30|然后狱警领他们出来，说：“二位先生，我必须做什么才可以得救？”
ACTS|16|31|他们说：“当信主耶稣，你和你一家都必得救 。”
ACTS|16|32|他们就把主的道讲给他和他全家的人听。
ACTS|16|33|当夜，就在那时候，狱警把他们带去，洗他们的伤；他和他所有的家人立刻都受了洗。
ACTS|16|34|于是狱警领他们上自己的家里去，给他们摆上饭。他和全家的人，因为信了上帝，都满心喜乐。
ACTS|16|35|到了天亮，官长们打发差役来，说：“释放那两个人吧。”
ACTS|16|36|狱警就把这些话告诉 保罗 ：“官长们打发人来，要释放你们，现在可以出监，平平安安去吧。”
ACTS|16|37|保罗 却说：“我们是 罗马 人，并没有定罪，他们竟在公众面前打了我们，又把我们下在监里；现在要私下赶我们出去吗？这不行！叫他们自己来领我们出去吧！”
ACTS|16|38|差役把这些话回禀官长们；官长们听见他们是 罗马 人，就害怕了，
ACTS|16|39|于是来劝他们，领他们出来，请他们离开那城。
ACTS|16|40|二人出了监牢，往 吕底亚 家里去，见了弟兄们，劝慰他们一番，就离开了。
ACTS|17|1|保罗 和 西拉 经过 暗妃坡里 、 亚波罗尼亚 ，来到 帖撒罗尼迦 ，在那里有 犹太 人的会堂。
ACTS|17|2|保罗 照他素常的规矩进去，一连三个安息日，根据圣经与他们辩论，
ACTS|17|3|讲解和说明基督必须受害，从死人中复活；又说：“我所传给你们的这位耶稣就是基督。”
ACTS|17|4|他们中间有些人听了劝，就跟从 保罗 和 西拉 ，还有许多虔敬的 希腊 人，尊贵的妇女也不少。
ACTS|17|5|但不信的 犹太 人心里嫉妒，聚集了些市井流氓，搭伙成群，煽动全城的人闯进 耶孙 的家，要把 保罗 和 西拉 带到民众那里。
ACTS|17|6|那些人找不着他们，就把 耶孙 和几个弟兄拉到地方官那里，喊叫着：“这些搅乱天下的人也到这里来了，
ACTS|17|7|耶孙 竟收留他们。这些人都违背凯撒的命令，说另有一个王耶稣。”
ACTS|17|8|众人和地方官听见这些话，就惶恐了，
ACTS|17|9|于是收了 耶孙 和其余的人的保证金后，释放了他们。
ACTS|17|10|当夜，弟兄们立刻送 保罗 和 西拉 往 庇哩亚 去；二人到了，就进入 犹太 人的会堂。
ACTS|17|11|这地方的 犹太 人比 帖撒罗尼迦 的人开明，热心领受这道，天天查考圣经，要知道这道是否真实。
ACTS|17|12|所以，他们中间有许多信了，又有 希腊 的尊贵妇人，男人也不少。
ACTS|17|13|但 帖撒罗尼迦 的 犹太 人知道 保罗 又在 庇哩亚 传上帝的道，就往那里去，煽动挑拨群众。
ACTS|17|14|于是，弟兄们立刻送 保罗 到海边去， 西拉 和 提摩太 却仍留在 庇哩亚 。
ACTS|17|15|护送 保罗 的人带他到了 雅典 ，他们领了 保罗 的命令，叫 西拉 和 提摩太 赶快到他那里来，然后回去了。
ACTS|17|16|保罗 在 雅典 等候他们的时候，看见满城都是偶像，就心里非常难过。
ACTS|17|17|于是他在会堂里与 犹太 人和虔敬的人，以及每日在市场上所遇见的人辩论。
ACTS|17|18|还有 伊壁鸠鲁 和 斯多亚 两派的哲学家也与他争辩。有的说：“这胡言乱语的要说什么？”有的说：“他似乎是宣传外邦鬼神的。”这是因 保罗 传讲耶稣与复活的福音。
ACTS|17|19|他们就把他带到 亚略巴古 ，说：“你所讲的这新学说，我们也可以知道吗？
ACTS|17|20|因为你有些奇怪的事传到我们耳中，我们想知道这些事是什么意思。”
ACTS|17|21|原来所有的 雅典 人和居住在那里的外国人都无暇管别的事，只是谈谈或听听新闻。
ACTS|17|22|保罗 站在 亚略巴古 当中，说：“诸位 雅典 人！我看你们凡事很敬畏鬼神。
ACTS|17|23|我到处走走的时候，仔细观察你们所敬拜的，发现一座坛，上面写着‘献给未识之神明’。你们所不认识而敬拜的，我现在向你们宣告：
ACTS|17|24|他是创造宇宙和其中万物的上帝；他既是天地的主，就不住在人手所造的殿宇里，
ACTS|17|25|也不用人手去服侍，好像缺少什么似的；自己倒将生命、气息、万物赐给万人。
ACTS|17|26|他从一人 造出万族，居住在全地面上，并且预先定准他们的年限和所住的疆界，
ACTS|17|27|为要使他们寻求上帝，或者可以揣摩而找到他，其实他离我们各人不远。
ACTS|17|28|我们生活、行动、存在都在于他。就如你们的诗人也有人说：‘我们也是他所生的。’
ACTS|17|29|既然我们是上帝所生的，就不应该以为上帝的神性像人用手艺和心思所雕刻的金、银、石像一般。
ACTS|17|30|世人蒙昧无知的时候，上帝并不追究，如今却吩咐各处的人都要悔改。
ACTS|17|31|因为他已经定了日子，要藉着他所设立的人按公义审判天下，并且使他从死人中复活，给万人作可信的凭据。”
ACTS|17|32|众人听见死人复活的话，就有人讥诮他；又有人说：“我们会再听你讲这事。”
ACTS|17|33|于是 保罗 从他们当中出去了。
ACTS|17|34|但有几个人依附他，信了主，其中有 亚略巴古 的议员 丢尼修 ，和一个名叫 大马哩 的妇人，还有几个与他们一起的人。
ACTS|18|1|这些事以后， 保罗 离开 雅典 ，来到 哥林多 。
ACTS|18|2|他遇见一个生在 本都 的 犹太 人，名叫 亚居拉 。不久前，他带着妻子 百基拉 从 意大利 来，因为 克劳第 命令所有的 犹太 人都离开 罗马 。 保罗 去投靠他们。
ACTS|18|3|他们本是制造帐棚为业。 保罗 因与他们同业，就和他们同住，一同做工。
ACTS|18|4|每逢安息日， 保罗 在会堂里辩论，劝导 犹太 人和 希腊 人。
ACTS|18|5|西拉 和 提摩太 从 马其顿 来的时候， 保罗 正专心传道，向 犹太 人证明耶稣是基督。
ACTS|18|6|当他们抗拒他、毁谤他的时候，他就抖掉衣裳的灰尘，对他们说：“你们的罪归到你们自己的头上，与我无干。从今以后，我要往外邦人那里去。”
ACTS|18|7|于是他离开那里，到了一个人的家里，他名叫 提多．犹士都 ，是敬拜上帝的人，他的家靠近会堂。
ACTS|18|8|会堂的主管 基利司布 和全家都信了主，还有许多 哥林多 人听了就信，而且受了洗。
ACTS|18|9|夜间，主在异象中对 保罗 说：“不要怕，只管讲，不要沉默，
ACTS|18|10|有我与你同在，没有人会下手害你，因为在这城里有许多属我的人。”
ACTS|18|11|保罗 在那里住了一年六个月，将上帝的道教导他们。
ACTS|18|12|到 迦流 作 亚该亚 省长的时候， 犹太 人齐心起来攻击 保罗 ，拉他到法庭，
ACTS|18|13|说：“这个人教唆人不按着律法敬拜上帝。”
ACTS|18|14|保罗 刚要开口， 迦流 对 犹太 人说：“你们这些 犹太 人哪！如果是为冤枉或奸恶的事，我理当耐性听你们。
ACTS|18|15|既然你们所争论的是关乎用字、名目和你们的律法，你们自己去办吧！这样的事我不愿意审问。”
ACTS|18|16|于是，他把他们逐出法庭。
ACTS|18|17|众人就揪住会堂的主管 所提尼 ，在法庭前打他。这些事 迦流 都不管。
ACTS|18|18|保罗 又住了好些日子，就辞别了弟兄，坐船到 叙利亚 去。 百基拉 、 亚居拉 和他同去。他因为许过愿，就在 坚革哩 剃了头发。
ACTS|18|19|到了 以弗所 ， 保罗 就把他们留在那里，自己进了会堂，和 犹太 人辩论。
ACTS|18|20|众人请他多住些日子，他没有答应，
ACTS|18|21|就辞别他们，说：“上帝若许可，我还要回到你们这里来。”于是他上船离开 以弗所 。
ACTS|18|22|他在 凯撒利亚 下了船，上 耶路撒冷 去问候教会，随后下 安提阿 去。
ACTS|18|23|他在那里住了些日子，又离开了那里，逐一经过 加拉太 和 弗吕家 各地方，坚固众门徒。
ACTS|18|24|有一个生在 亚历山大 的 犹太 人，名叫 亚波罗 ，来到 以弗所 ，他很有口才，很会讲解圣经。
ACTS|18|25|这人已经在主的道路上受了训练，心里火热，精确地讲论和教导耶稣的事；可是他只知道 约翰 的洗礼。
ACTS|18|26|他开始在会堂里放胆讲道； 百基拉 、 亚居拉 听见，就接他来，将上帝的道路 给他更精确地讲解。
ACTS|18|27|他想要往 亚该亚 去，弟兄们就勉励他，并写信请门徒们接待他，他到了那里，多多帮助那些蒙恩信主的人，
ACTS|18|28|因为他在公众面前极力驳倒 犹太 人，引圣经证明耶稣是基督。
ACTS|19|1|亚波罗 在 哥林多 的时候， 保罗 经过了内陆地区，来到 以弗所 ，在那里他遇见几个门徒，
ACTS|19|2|问他们：“你们信的时候领受了圣灵没有？”他们说：“没有，我们连什么是圣灵都没有听过。”
ACTS|19|3|保罗 说：“这样，你们受的是什么洗呢？”他们说：“是受了 约翰 的洗。”
ACTS|19|4|保罗 说：“ 约翰 所施的是悔改的洗礼，他告诉百姓当信那在他以后要来的那位，就是耶稣。”
ACTS|19|5|他们听见这话以后，就奉主耶稣的名受洗。
ACTS|19|6|保罗 给他们按手，圣灵就降在他们身上，他们开始说方言 和说预言。
ACTS|19|7|他们约有十二个人。
ACTS|19|8|保罗 进会堂，一连三个月放胆讲道，辩论上帝国的事，劝导众人。
ACTS|19|9|后来，有些人心里刚硬不信，在众人面前毁谤这道； 保罗 就离开他们，也叫门徒与他们分开，就在 推喇奴 的讲堂天天辩论。
ACTS|19|10|这样有两年之久，使一切住在 亚细亚 的，无论是 犹太 人是 希腊 人，都听见主的道。
ACTS|19|11|上帝藉 保罗 的手行了些奇异的神迹，
ACTS|19|12|甚至有人从 保罗 身上拿走手巾或围裙放在病人身上，病就消除了，邪灵也出去了。
ACTS|19|13|那时，有几个巡回各处念咒赶鬼的 犹太 人，擅自利用主耶稣的名，向那些被邪灵所附的人说：“我奉 保罗 所传的耶稣命令你们出来！”
ACTS|19|14|做这事的是 犹太 祭司长 士基瓦 的七个儿子。
ACTS|19|15|但邪灵回答他们：“耶稣我知道， 保罗 我也认识，你们却是谁呢？”
ACTS|19|16|被邪灵所附的人就扑到他们身上，制伏他们，胜过他们，使他们赤着身子，受了伤，从那房子里逃出去了。
ACTS|19|17|凡住在 以弗所 的，无论是 犹太 人是 希腊 人，都知道这件事，也都惧怕；主耶稣的名从此就更被尊为大了。
ACTS|19|18|许多已经信的人来承认并公开自己所行的事。
ACTS|19|19|又有许多平素行邪术的人把他们的书都拿来，堆积在众人面前焚烧。他们计算书价，得知共值五万块银钱。
ACTS|19|20|这样，主的道大大兴旺，而且普遍传开了。
ACTS|19|21|这些事过后， 保罗 心里决定要经过 马其顿 、 亚该亚 ，就往 耶路撒冷 去。他说：“我到了那里以后，也必须到 罗马 去看看。”
ACTS|19|22|于是他差遣两个助手 提摩太 和 以拉都 往 马其顿 去，自己暂时留在 亚细亚 。
ACTS|19|23|那时，因这道路而起的骚动不小。
ACTS|19|24|有一个银匠，名叫 底米丢 ，是制造 亚底米 神银龛的，他使从事这手艺的人生意发达。
ACTS|19|25|他聚集他们和同行的工人，说：“诸位，你们知道我们是倚靠这生意发财的。
ACTS|19|26|你们看到，也听见这 保罗 不但在 以弗所 ，也几乎在 亚细亚 全地，引诱迷惑了许多人，说：‘人手所做的不是神明。’
ACTS|19|27|这样，不仅我们这行业陷入被藐视的危险，就是大女神 亚底米 的庙也要被人轻看，连 亚细亚 全地和普天下所敬拜的女神的威望也受损害了。”
ACTS|19|28|众人听见，就怒气冲冲，喊着说：“大哉， 以弗所 人的 亚底米 ！”
ACTS|19|29|于是满城都骚动起来。众人抓住与 保罗 同行的 马其顿 人 该犹 和 亚里达古 ，齐心冲进剧场。
ACTS|19|30|保罗 想要进到民众那里，门徒却不许他去。
ACTS|19|31|连 亚细亚 的几位官员，是 保罗 的朋友，也打发人来劝他不要冒险到剧场里去。
ACTS|19|32|聚集的人乱成一团，有的喊这个，有的喊那个，大半不知道为了什么聚集。
ACTS|19|33|犹太 人把 亚历山大 推出去，人群中有人怂恿他，他就做手势，要向民众申诉。
ACTS|19|34|但他们一认出他是 犹太 人，大家就异口同声喊着：“大哉， 以弗所 人的 亚底米 ！”约喊了两小时。
ACTS|19|35|城里的书记官安抚了群众后，说：“ 以弗所 人哪，谁不知道 以弗所 人的城是看守大 亚底米 的庙和从 宙斯 那里落下来的像的守护者呢？
ACTS|19|36|既然这些事是驳不倒的，你们就要安静下来，不可妄动。
ACTS|19|37|你们把这些人带来，他们并没有偷窃庙中之物，也没有亵渎我们的女神。
ACTS|19|38|如果 底米丢 和他同行的手艺人有控告的事，自有公堂，也有省长，他们可以彼此控告。
ACTS|19|39|你们若有别的事请求，可以在合法的集会里解决。
ACTS|19|40|今日的扰乱本是无缘无故的，有被控告的危险。这次的骚动，我们也说不出理由来。”
ACTS|19|41|他说完这些话，就叫众人散会。
ACTS|20|1|骚乱平定以后， 保罗 请门徒来，劝勉了他们，就辞别他们，往 马其顿 去。
ACTS|20|2|他走遍那一带地方，用许多话劝勉门徒，然后来到 希腊 ，
ACTS|20|3|在那里住了三个月。他快要坐船往 叙利亚 去的时候， 犹太 人设计害他，他就决定从 马其顿 回去。
ACTS|20|4|同他到 亚细亚 去的，有 庇哩亚 人 毕罗斯 的儿子 所巴特 ， 帖撒罗尼迦 人 亚里达古 和 西公都 ，还有 特庇 人 该犹 和 提摩太 ，又有 亚细亚 人 推基古 和 特罗非摩 。
ACTS|20|5|这些人先走，在 特罗亚 等候我们。
ACTS|20|6|过了除酵节的日子，我们从 腓立比 开船，五天以后到了 特罗亚 ，和他们相会，在那里住了七天。
ACTS|20|7|七日的第一日，我们聚会擘饼的时候， 保罗 因次日要起行，就为他们讲道，直讲到半夜。
ACTS|20|8|我们聚会的那座楼上有好些灯火。
ACTS|20|9|有一个少年，名叫 犹推古 ，坐在窗口上，沉沉入睡。 保罗 讲了多时，少年睡熟了，从三层楼上掉下去，扶起来时已经死了。
ACTS|20|10|保罗 下去，伏在他身上，抱着他，说：“你们不要慌乱，他还有气呢！”
ACTS|20|11|保罗 又上楼去，擘饼，吃了，再讲了许久，直到天亮才离开。
ACTS|20|12|他们把那活过来的孩子带走，大家得到很大的安慰。
ACTS|20|13|我们先上船，起航往 亚朔 去，想要在那里接 保罗 ；因为他是这样安排的，他自己本来打算要走陆路。
ACTS|20|14|他既在 亚朔 与我们相会，我们就接他上船，来到 米推利尼 。
ACTS|20|15|我们从那里开船，第二天到了 基阿 的对岸；再下一天，在 撒摩 靠岸，又过了一天，到了 米利都 。
ACTS|20|16|因为 保罗 早已决定要越过 以弗所 ，免得在 亚细亚 耽延，他急忙前行，假如可能的话，在五旬节前能赶到 耶路撒冷 。
ACTS|20|17|保罗 从 米利都 打发人往 以弗所 去，请教会的长老来。
ACTS|20|18|他们来了， 保罗 对他们说：“你们自己知道，自从我到 亚细亚 的第一天，我怎样跟你们相处，
ACTS|20|19|怎样凡事谦卑，以眼泪服侍主，又因 犹太 人的谋害经历试炼。
ACTS|20|20|你们也知道，凡对你们有益的，我没有一样隐瞒不说的，或在公众面前，或在每一个人的家里，我都教导你们，
ACTS|20|21|不论 犹太 人和 希腊 人，我都已证明他们当在上帝面前悔改，信靠我们的主耶稣。
ACTS|20|22|现在我被圣灵催迫 要往 耶路撒冷 去，虽然不知道在那里会遭遇什么事，
ACTS|20|23|但知道圣灵在各城里向我指证，说有捆锁与患难等着我。
ACTS|20|24|我却不以性命为念，只要走完我的路程，完成我从主耶稣所领受的职分，为上帝恩典的福音作见证。
ACTS|20|25|“我素常在你们中间到处传讲上帝的国；现在我知道，你们众人以后不会再见到我的面了。
ACTS|20|26|所以我今日向你们作证，你们中间无论何人死亡，罪不在我。
ACTS|20|27|因为上帝一切的旨意，我并没有退缩不传给你们的。
ACTS|20|28|圣灵立你们作全群的监督，你们就当为自己谨慎，也为全群谨慎，牧养上帝 的教会，就是他用自己血所买来的 。
ACTS|20|29|我知道，在我离开以后必有凶暴的豺狼进入你们中间，不顾惜羊群。
ACTS|20|30|就是你们中间也必有人起来，说悖谬的话，要引诱门徒跟从他们。
ACTS|20|31|所以你们要警醒，记念我三年之久，昼夜不断地流泪劝戒你们各人。
ACTS|20|32|现在我把你们交托给上帝和他恩惠的道；这道能建立你们，使你们和一切成圣的人同得基业。
ACTS|20|33|我未曾贪图一个人的金、银或衣服。
ACTS|20|34|你们自己知道，我靠两只手工作来供给我和同工的需用。
ACTS|20|35|我凡事给你们作榜样，叫你们知道应当这样劳苦，扶助软弱的人，又当记念主耶稣的话，说：‘施比受更为有福。’”
ACTS|20|36|保罗 说完了这些话，就和大家跪下来祷告。
ACTS|20|37|众人痛哭，抱着 保罗 的颈项跟他亲吻。
ACTS|20|38|叫他们最伤心的，就是他说“以后不会再见到我的面”那句话。于是他们送他上船去了。
ACTS|21|1|我们离别了众人，就开船直航到 哥士 ，第二天到了 罗底 ，又从那里到 帕大喇 。
ACTS|21|2|我们遇见一只船要往 腓尼基 去，就上船起航。
ACTS|21|3|我们望见 塞浦路斯 ，就从南边行过，往 叙利亚 去，在 推罗 上岸，因为船要在那里卸货。
ACTS|21|4|我们在那里找到了一些门徒，就住了七天。他们藉着圣灵的感动，告诉 保罗 不要上 耶路撒冷 去。
ACTS|21|5|几天之后，我们又出发前行。他们众人同妻子儿女都送我们到城外，我们都跪在滩上祷告，彼此辞别。
ACTS|21|6|我们上了船，他们就回家去了。
ACTS|21|7|我们从 推罗 行完航程，来到了 多利买 ，问候那里的弟兄，和他们同住了一天。
ACTS|21|8|第二天，我们离开那里，来到 凯撒利亚 ，就进了传福音的 腓利 家里，和他同住；他是那七个执事里的一个。
ACTS|21|9|他有四个女儿，都是未出嫁的，都会说预言。
ACTS|21|10|我们在那里多住了好几天，有一个先知，名叫 亚迦布 ，从 犹太 下来。
ACTS|21|11|他到了我们这里，就拿 保罗 的腰带，捆上自己的手脚，说：“圣灵这样说：‘ 犹太 人在 耶路撒冷 要如此捆绑这腰带的主人，把他交在外邦人手里。’”
ACTS|21|12|我们听见这些话，就跟当地的人苦劝 保罗 不要上 耶路撒冷 去。
ACTS|21|13|于是 保罗 回答：“你们为什么这样痛哭，使我心碎呢？我为主耶稣的名，不但被人捆绑，就是死在 耶路撒冷 也是愿意的。”
ACTS|21|14|既然 保罗 不听劝，我们就住了口，只说：“愿主的旨意成就。”
ACTS|21|15|过了这几天，我们收拾行李上 耶路撒冷 去。
ACTS|21|16|有 凯撒利亚 的几个门徒和我们同去，带我们到一个早期的门徒 塞浦路斯 人 拿孙 的家里，请我们与他同住。
ACTS|21|17|我们到了 耶路撒冷 ，弟兄们欢欢喜喜地接待我们。
ACTS|21|18|第二天， 保罗 同我们去见 雅各 ；所有的长老也都在场。
ACTS|21|19|保罗 向他们问安，然后将上帝用他在外邦人中所做的事奉，一一述说了。
ACTS|21|20|他们听见了，就归荣耀给上帝，对 保罗 说：“弟兄，你看 犹太 人中有数以万计的信徒，而他们都是热心于律法的人。
ACTS|21|21|他们曾听见人说，你教导所有在外邦的 犹太 人离弃 摩西 ，对他们说，不要给孩子行割礼，也不要遵守规矩。
ACTS|21|22|众人必听见你来了，这可怎么办呢？
ACTS|21|23|你就照着我们的话做吧！我们这里有四个人，都有愿在身。
ACTS|21|24|你带他们去，与他们一同行洁净的礼，替他们缴纳规费，让他们得以剃头。这样，众人就会知道，先前所听见关于你的事都是假的；而且也知道，你自己为人循规蹈矩，遵行律法。
ACTS|21|25|至于信主的外邦人， 我们已经根据我们的决议写信，叫他们要禁戒偶像所玷污的东西、血和勒死的牲畜，禁戒淫乱。”
ACTS|21|26|于是 保罗 带着那四个人，第二天与他们一同行了洁净礼，进了圣殿，报告洁净期满的日子，等候祭司为他们各人献上祭物。
ACTS|21|27|那七日将完，从 亚细亚 来的 犹太 人看见 保罗 在圣殿里，就煽动所有的群众，下手拿住他，
ACTS|21|28|喊着：“ 以色列 人哪，来帮忙！这就是在各处教导众人糟蹋我们百姓、律法和这地方的人。不但如此，他还带了 希腊 人进圣殿，污秽了这圣地。”
ACTS|21|29|这话是因他们曾看见 以弗所 人 特罗非摩 跟 保罗 一起在城里，以为 保罗 带他进了圣殿。
ACTS|21|30|于是全城都骚动，百姓一齐跑来，拿住 保罗 ，拉他出圣殿，殿门立刻都关了。
ACTS|21|31|他们正想要杀他，有人报信给营里的千夫长，说 耶路撒冷 全城都乱了。
ACTS|21|32|千夫长立刻带着士兵和几个百夫长，跑下去到他们那里。他们见了千夫长和士兵，就停下来不打 保罗 。
ACTS|21|33|于是千夫长上前拿住他，吩咐用两条铁链捆锁，又问他是什么人，做了什么事。
ACTS|21|34|群众中有的喊这个，有的喊那个；因为这样乱嚷，千夫长无法知道实情，就下令将 保罗 带进营楼去。
ACTS|21|35|保罗 一走上台阶，群众挤得凶猛，士兵只得将 保罗 抬起来。
ACTS|21|36|一群人跟在后面，喊着：“除掉他！”
ACTS|21|37|保罗 快要被带进营楼时，对千夫长说：“我可以对你说句话吗？”千夫长说：“你懂得 希腊 话吗？
ACTS|21|38|那你就不是从前作乱、带领四千凶徒往旷野去的那 埃及 人了。”
ACTS|21|39|保罗 说：“我本是 犹太 人，生在 基利家 的 大数 ，并不是无名小城的公民。求你准我对百姓说话。”
ACTS|21|40|千夫长准了。 保罗 就站在台阶上，向百姓做了个手势，要他们静下来， 保罗 就用 希伯来 话对他们说：
ACTS|22|1|“诸位父老弟兄，请听我现在对你们的申辩。”
ACTS|22|2|他们听 保罗 说的是 希伯来 话，就更加安静了。
ACTS|22|3|保罗 说：“我原是 犹太 人，生在 基利家 的 大数 ，但在这城里长大，在 迦玛列 门下按着我们祖宗严紧的律法受教，热心事奉上帝，就如你们大家今日一样。
ACTS|22|4|我也曾迫害信奉这道路的人，置他们于死地，无论男女都捆绑，关在监里。
ACTS|22|5|这是大祭司和议会的众长老都可以给我作证的。我又从他们那里领了致弟兄们的书信，往 大马士革 去，要把在那里的信徒绑起来，带到 耶路撒冷 受刑。”
ACTS|22|6|“当我走近 大马士革 的时候，约在中午，忽然有一道大光从天上下来，照射在我周围。
ACTS|22|7|我就仆倒在地，听见有声音对我说：‘ 扫罗 ！ 扫罗 ！你为什么迫害我？’
ACTS|22|8|我回答：‘主啊！你是谁？’他对我说：‘我就是你所迫害的 拿撒勒 人耶稣。’
ACTS|22|9|跟我一起的人看见了那光，却没有听见那位对我说话的声音。
ACTS|22|10|我说：‘主啊，我该做什么？’主说：‘起来，进 大马士革 去，在那里有人会把指派你做的一切事告诉你。’
ACTS|22|11|我因那光的闪耀不能看见，跟我一起的人就拉着我的手进了 大马士革 。
ACTS|22|12|“那里有一个人，名叫 亚拿尼亚 ，按着律法是虔诚人，为所有住在那里的 犹太 人所称赞。
ACTS|22|13|他来见我，站在旁边，对我说：‘ 扫罗 弟兄，你看见吧！’就在那时，我恢复视觉，看见了他。
ACTS|22|14|他又说：‘我们祖宗的上帝拣选了你，让你明白他的旨意，又看见那义者，听见他口中所出的声音。
ACTS|22|15|因为你要将所看见的、所听见的，对着万人作他的见证人。
ACTS|22|16|现在你为什么耽延呢？起来，受洗，求告他的名，洗去你的罪。’”
ACTS|22|17|“后来，我回到 耶路撒冷 ，在圣殿里祷告的时候，魂游象外，
ACTS|22|18|看见主对我说：‘你赶紧离开 耶路撒冷 ，越快越好，因为这里的人不接受你为我作的见证。’
ACTS|22|19|我就说：‘主啊，他们都知道，我从前在各会堂里把信你的人监禁，又鞭打他们。
ACTS|22|20|当你的见证人 司提反 被害流血的时候，我也站在一旁赞同；又为打死他的人看守衣裳。’
ACTS|22|21|主对我说：‘你去吧！我要差你到远方外邦人那里去。’”
ACTS|22|22|众人听他说到这句话，就高声说：“这样的人，从地上除掉他吧！他是该死的。”
ACTS|22|23|大家一边喧嚷一边摔衣裳，向空中撒灰尘。
ACTS|22|24|千夫长下令把 保罗 带进营楼，叫人用鞭子拷问他，要知道他们向他这样喧嚷是什么缘故。
ACTS|22|25|他们刚用皮条把他捆上的时候， 保罗 对站在旁边的百夫长说：“一个 罗马 人，又未被定罪，你们就鞭打他是合法的吗？”
ACTS|22|26|百夫长听见这话，就去见千夫长，报告说：“你要怎么办呢？这个人是 罗马 人。”
ACTS|22|27|千夫长就来问 保罗 ：“你告诉我，你是 罗马 人吗？” 保罗 说：“是。”
ACTS|22|28|千夫长回答：“我用了许多银子才得到 罗马 公民的身份。” 保罗 说：“我生来就是。”
ACTS|22|29|于是那些要拷问 保罗 的人立刻离开他走了。千夫长一知道他是 罗马 人，又因为曾捆绑了他，也害怕起来。
ACTS|22|30|第二天，千夫长为要知道 犹太 人控告 保罗 的实情，就解开他，下令祭司长们和全议会的人都聚集，然后将 保罗 带下来，叫他站在他们面前。
ACTS|23|1|保罗 定睛看着议会的人，说：“诸位弟兄，我在上帝面前，行事为人都是凭着清白的良心，直到今日。”
ACTS|23|2|亚拿尼亚 大祭司就吩咐旁边站着的人打他的嘴。
ACTS|23|3|这时， 保罗 对他说：“你这粉饰的墙，上帝要打你！你坐堂是要按律法审问我，你竟违背律法，命令人打我吗？”
ACTS|23|4|站在旁边的人说：“你竟敢辱骂上帝的大祭司吗？”
ACTS|23|5|保罗 说：“弟兄们，我不知道他是大祭司；因为经上记着：‘不可毁谤你百姓的官长。’”
ACTS|23|6|保罗 看出他们一部分是撒都该人，一部分是法利赛人，就在议会中喊着：“诸位弟兄，我是法利赛人，也是法利赛人的子孙。我现在受审问是为有关死人复活的盼望。”
ACTS|23|7|说了这话，法利赛人和撒都该人争论起来，会众分为两派。
ACTS|23|8|因为撒都该人一方面说没有复活，另一方面没有天使和鬼魂；法利赛人却承认两方面都有。
ACTS|23|9|于是大大地争吵起来；有几个法利赛派的文士站起来争辩说：“我们看不出这人有什么错处；说不定有鬼魂或者天使对他说过话呢！”
ACTS|23|10|那时争辩越来越大，千夫长恐怕 保罗 被他们扯碎了，就命令士兵下去，把他从众人当中抢出来，带进营楼去。
ACTS|23|11|当夜，主站在 保罗 旁边，说：“放心吧！你怎样在 耶路撒冷 为我作见证，也必怎样在 罗马 为我作见证。”
ACTS|23|12|到了天亮， 犹太 人同谋起誓，说“若不先杀 保罗 就不吃不喝”。
ACTS|23|13|参与这阴谋的有四十多人。
ACTS|23|14|他们来见祭司长和长老，说：“我们已经发了重誓，若不先杀 保罗 就什么也不吃。
ACTS|23|15|现在你们和议会要通知千夫长，叫他把 保罗 带到你们这里来，假装要详细调查他的事；我们已经预备好，在他来到这里以前就杀掉他。”
ACTS|23|16|保罗 的外甥听见他们设下埋伏，就来到营楼里告诉 保罗 。
ACTS|23|17|保罗 请一个百夫长来，说：“你领这青年去见千夫长，他有事告诉他。”
ACTS|23|18|于是百夫长把他领去见千夫长，说：“被囚的 保罗 请我到他那里，求我领这青年来见你；他有事告诉你。”
ACTS|23|19|千夫长就拉着他的手，走到一旁，私下问他：“你有什么事告诉我呢？”
ACTS|23|20|他说：“ 犹太 人已经约定，要求你明天把 保罗 带到议会去，假装要详细查问他的事。
ACTS|23|21|你切不要随从他们，因为他们有四十多人埋伏，已经起誓，若不先杀掉 保罗 就不吃不喝。现在都预备好了，只等你的允准。”
ACTS|23|22|于是千夫长打发那青年走，嘱咐他：“不要告诉人，你已将这些事报告我了。”
ACTS|23|23|于是，千夫长叫了两个百夫长来，说：“预备步兵二百、骑兵七十、长枪手二百，今夜九点往 凯撒利亚 去；
ACTS|23|24|也要预备牲口让 保罗 骑上，护送到 腓力斯 总督那里去。”
ACTS|23|25|千夫长又写了公文，大略说：
ACTS|23|26|“ 克劳第．吕西亚 向 腓力斯 总督大人请安。
ACTS|23|27|这个人被 犹太 人拿住，快被杀害时，我得知他是 罗马 人，就带士兵下去，把他救了出来。
ACTS|23|28|因为我要知道他们告他的罪状，就带他下到他们的议会去。
ACTS|23|29|我查知他被告发是因他们律法上的争论，并没有什么该死或该监禁的罪名。
ACTS|23|30|后来有人把要害他的计谋告诉我，我立刻把他解到你那里去，又命令告他的人在你面前告他。 ”
ACTS|23|31|于是士兵照所命令他们的，连夜把 保罗 带到 安提帕底 。
ACTS|23|32|第二天，由骑兵护送 保罗 ，他们就回营楼去。
ACTS|23|33|骑兵来到 凯撒利亚 ，把公文呈给总督，就叫 保罗 站在他面前。
ACTS|23|34|总督读了公文，问 保罗 是哪一省的人；一知道他是 基利家 人，
ACTS|23|35|就说：“等告你的人来到，我才详细听你。”于是他命令把 保罗 拘留在 希律 的衙门里。
ACTS|24|1|过了五天， 亚拿尼亚 大祭司、几个长老和一个叫 帖土罗 的律师下来，向总督控告 保罗 。
ACTS|24|2|保罗 一被传来， 帖土罗 就开始控告他，说：“ 腓力斯 大人，我们因你得以享受国泰民安，并且这一国的弊病，因着你的远见得以改革。
ACTS|24|3|我们随时随地都满心感激不尽。
ACTS|24|4|为了不敢耽搁你太久，我只求你宽容一下，听我们说几句话。
ACTS|24|5|我们看这个人如同瘟疫一般，是鼓动普天下所有的 犹太 人作乱的人，又是 拿撒勒 教派里的一个头目。
ACTS|24|6|他甚至连圣殿也要污秽，我们就把他捉拿了。
ACTS|24|7|
ACTS|24|8|你自己审问他，就可以知道我们所控告他的一切事了。”
ACTS|24|9|众 犹太 人也随着控告他，说：“这些事情确是这样。”
ACTS|24|10|总督示意叫 保罗 说话， 保罗 就回答：“我知道你在本国作法官多年，所以我乐意为自己申辩。
ACTS|24|11|你查问就可以知道，从我上 耶路撒冷 去礼拜到今日不过十二天。
ACTS|24|12|他们并没有看见我在圣殿里跟人辩论，或在会堂里、在城里煽动群众。
ACTS|24|13|也不能对你证实他们现在所控告我的事。
ACTS|24|14|但有一件事我向你承认，就是我正按着他们所称为异端的道事奉我祖宗的上帝，又信合乎律法和先知书上所记载的一切。
ACTS|24|15|我对上帝存着这些人自己也接受的盼望，就是义人和不义的人都要复活。
ACTS|24|16|因此，我勉励自己，对上帝对人，时常存着无亏的良心。
ACTS|24|17|过了几年，我带着周济本国的捐项和供物上去。
ACTS|24|18|正献的时候，他们看见我在圣殿里已经洁净了，并没有聚众，也没有吵嚷，
ACTS|24|19|惟有几个从 亚细亚 来的 犹太 人—他们若有控告我的事，应当到你面前来告我。
ACTS|24|20|不然，让这些人自己说，他们看出我站在议会前的时间，有什么不对的地方。
ACTS|24|21|纵然有，也不过是为了一句话，就是我站在他们中间喊说：‘我今日在你们面前受审，是为了死人复活。’”
ACTS|24|22|腓力斯 本是详细认识这道，就拖延他们，说：“且等 吕西亚 千夫长下来，我再审判你们的案。”
ACTS|24|23|于是他下令百夫长看守 保罗 ，要从宽待他，不可拦阻他的亲友来供给他。
ACTS|24|24|过了几天， 腓力斯 和他夫人 犹太 女子 土西拉 一同来到，就叫 保罗 来，听他讲论信基督耶稣的事。
ACTS|24|25|保罗 讲论公义、节制和将来的审判， 腓力斯 害怕起来，就回答：“你暂且去吧！等我有机会时再来叫你。”
ACTS|24|26|腓力斯 又指望 保罗 送他银钱，所以屡次叫他来，和他谈论。
ACTS|24|27|过了两年， 波求．非斯都 接了 腓力斯 的任； 腓力斯 要讨 犹太 人的喜欢，就把 保罗 留在监里。
ACTS|25|1|非斯都 到省里上任，过了三天，就从 凯撒利亚 上 耶路撒冷 去。
ACTS|25|2|祭司长和 犹太 人的领袖向他控告 保罗 ；又央求他，
ACTS|25|3|向他求情要对付 保罗 ，把他提到 耶路撒冷 来，他们要在路上埋伏杀害他。
ACTS|25|4|非斯都 就回答：“ 保罗 押在 凯撒利亚 ，我自己快要往那里去。”
ACTS|25|5|他又说：“所以，你们中间有权的人与我一同下去，那人若有什么不是，就让他们控告他。”
ACTS|25|6|非斯都 在他们那里住了不超过八天或十天，就下 凯撒利亚 去；第二天开庭，下令把 保罗 提上来。
ACTS|25|7|保罗 来了，那些从 耶路撒冷 下来的 犹太 人周围站着，提出许多严重而不能证实的事控告他。
ACTS|25|8|保罗 申辩说：“无论 犹太 人的律法，或是圣殿，或是凯撒，我都没有干犯。”
ACTS|25|9|但 非斯都 要讨 犹太 人的喜欢，就回答 保罗 说：“你愿意上 耶路撒冷 去，在那里为这些事受我的审判吗？”
ACTS|25|10|保罗 说：“我现在站在凯撒的审判台前，这就是我应当受审的地方。我并没有对 犹太 人做过什么不对的事，这也是你明明知道的。
ACTS|25|11|我若做了不对的事，犯了什么该死的罪，就是死我也不辞。他们所控告我的事若都不实，就没有人能把我交给他们。我要向凯撒上诉。”
ACTS|25|12|非斯都 和议会商量了，就回答：“既然你要向凯撒上诉，你就到凯撒那里去吧。”
ACTS|25|13|过了些日子， 亚基帕 王和 百妮基 来到 凯撒利亚 ，拜访 非斯都 。
ACTS|25|14|他们在那里住了好些日子， 非斯都 将 保罗 的案件向王陈述，说：“这里有一个人，是 腓力斯 留在监里的。
ACTS|25|15|我在 耶路撒冷 的时候，祭司长和 犹太 的长老把他的事禀报了，要求定他的罪。
ACTS|25|16|我回覆他们，无论什么人，被告还没有和原告当面对质，没有机会为所控告的事申辩，就先定他罪的，这不是 罗马 人的规矩。
ACTS|25|17|及至他们都来到这里，我没有耽误，第二天就开庭，下令把那人提上来。
ACTS|25|18|控告他的人站起来告他，所控告的并没有任何我所预料的那等恶 事。
ACTS|25|19|不过，有几样辩论是有关他们自己敬鬼神的事，以及一个名叫耶稣的人，他已经死了， 保罗 却说他是活着的。
ACTS|25|20|我对这些事不知该怎样处理，所以问他是否愿意上 耶路撒冷 去，在那里为这些事接受审判。
ACTS|25|21|但 保罗 要求我留下他，要听皇上判断，我就下令把他留下，等我解他到凯撒那里去。”
ACTS|25|22|亚基帕 对 非斯都 说：“我也愿意亲自听听这个人。” 非斯都 说：“明天你就可以听他。”
ACTS|25|23|第二天， 亚基帕 和 百妮基 大张旗鼓而来，与众千夫长和城里的显要进了大厅。 非斯都 一声令下，就有人将 保罗 带进来。
ACTS|25|24|非斯都 说：“ 亚基帕 王和在这里的诸位，你们看这个人，他就是所有在 耶路撒冷 和这里的 犹太 人曾向我恳求呼叫，说不可容他再活着的。
ACTS|25|25|但我查明他并没有犯什么该死的罪，并且他自己也已向皇帝上诉了，所以我决定把他解去。
ACTS|25|26|论到这个人，我没有确实的事可以奏明主上。因此，我带他到你们面前，尤其到你 亚基帕 王面前，为要在查问之后有所呈奏。
ACTS|25|27|因为据我看，解送囚犯而不指明他的罪状是不合理的。”
ACTS|26|1|亚基帕 对 保罗 说：“准你为自己申诉。”于是 保罗 伸手辩护说：
ACTS|26|2|“ 亚基帕 王啊， 犹太 人所控告我的一切事，今日得以在你面前辩护，实为万幸。
ACTS|26|3|更庆幸的是你熟悉 犹太 人的规矩和他们的争论；所以，求你耐心听我。
ACTS|26|4|“我自幼为人如何，从起初在本国的同胞中，以及在 耶路撒冷 ，所有的 犹太 人都知道。
ACTS|26|5|他们若肯作见证，就知道我从起初是按着我们教中最严紧的教门作了法利赛人。
ACTS|26|6|现在我站在这里受审，是为了对上帝向我们祖宗的应许存着盼望。
ACTS|26|7|这应许，我们十二个支派，昼夜切切地事奉上帝，都指望得着。王啊，我正是因这指望被 犹太 人控告。
ACTS|26|8|上帝使死人复活，你们为什么判断为不可信呢？
ACTS|26|9|“从前我自己认为必须竭力反对 拿撒勒 人耶稣的名，
ACTS|26|10|我在 耶路撒冷 也曾这样做过；我不但从祭司长得了权柄，把许多圣徒收在监里，而且他们被杀，我也表示 赞成。
ACTS|26|11|在各会堂，我屡次用刑强迫他们说亵渎的话，我非常厌恶他们，甚至追逼他们，直到外邦的城镇。”
ACTS|26|12|“那时，我带着祭司长的权柄和命令往 大马士革 去。
ACTS|26|13|王啊！我在路上，中午的时候，看见从天上有一道光，比太阳还亮，四面照射着我和跟我同行的人。
ACTS|26|14|我们都仆倒在地，我就听见有声音用 希伯来 话对我说：‘ 扫罗 ！ 扫罗 ！你为什么迫害我？你用脚踢刺棒是自找苦吃的！’
ACTS|26|15|我说：‘主啊，你是谁？’主说：‘我就是你所迫害的耶稣。
ACTS|26|16|起来，站着，我向你显现的目的是要派你作仆役，为你所看见我 的事，和我将要指示你的事作见证人。
ACTS|26|17|我也要救你脱离百姓和外邦人的手。我差你到他们那里去，
ACTS|26|18|要开他们的眼睛，使他们从黑暗中转向光明，从撒但权下归向上帝；使他们因信我而得蒙赦罪，和一切成圣的人同得基业。’”
ACTS|26|19|“因此， 亚基帕 王啊！我没有违背那从天上来的异象；
ACTS|26|20|我先在 大马士革 ，后在 耶路撒冷 和 犹太 全地，以及外邦，劝勉他们应当悔改归向上帝，行事与悔改的心相称。
ACTS|26|21|为这缘故， 犹太 人在圣殿里拿住我，想要杀我。
ACTS|26|22|然而，我蒙上帝的帮助，直到今日还站立得稳，向尊贵的和卑微的作见证。我所讲的，并不外乎众先知和 摩西 所说将来必成的事，
ACTS|26|23|就是基督必须受害，并且首先从死人中复活，把亮光传给 犹太 人和外邦人。”
ACTS|26|24|保罗 这样申诉时， 非斯都 大声说：“ 保罗 ，你疯了！你的学问太大，反使你疯了！”
ACTS|26|25|保罗 说：“ 非斯都 大人，我不是疯了，我说的乃是真实和清醒的话。
ACTS|26|26|王也知道这些事，所以对王大胆直言，我深信这些事没有一件能向王隐瞒的，因为都不是在背地里做的。
ACTS|26|27|亚基帕 王啊，你信先知吗？我知道你是信的。”
ACTS|26|28|亚基帕 对 保罗 说：“你想稍微劝一劝就能说服我作基督徒了吗？”
ACTS|26|29|保罗 说：“无论少劝还是多劝，我向上帝所求的，不但你一个人，就是今天所有听我说话的人都要像我一样，只是不要有这些锁链。”
ACTS|26|30|于是，王和总督以及 百妮基 跟同坐的人都站起来，
ACTS|26|31|退到里面，彼此谈论说：“这个人并没有犯什么该死该监禁的罪。”
ACTS|26|32|亚基帕 对 非斯都 说：“这人若没有向凯撒上诉，早就被释放了。”
ACTS|27|1|既然 非斯都 决定要我们坐船往 意大利 去，就将 保罗 和别的囚犯交给御营里的一个名叫 犹流 的百夫长。
ACTS|27|2|有一只 亚大米田 的船要开往 亚细亚 沿海一带地方去，我们上了那船，就起航了；有 马其顿 的 帖撒罗尼迦 人 亚里达古 和我们同去。
ACTS|27|3|第二天，我们到了 西顿 。 犹流 宽待 保罗 ，准他往朋友那里去，受他们的照应。
ACTS|27|4|我们又从那里开船，因为遇到逆风，就贴着 塞浦路斯 的背风岸航行，
ACTS|27|5|渡过了 基利家 、 旁非利亚 一带的海面，就到了 吕家 的 每拉 。
ACTS|27|6|在那里，百夫长找到一只 亚历山大 的船要往 意大利 去，就叫我们上了那船。
ACTS|27|7|一连多日，船行得很慢，我们好不容易才来到 革尼土 的对面；又因被风拦阻，我们就贴着 克里特岛 背风岸，从 撒摩尼 对面航行。
ACTS|27|8|我们沿岸前进，十分艰难，来到一个名叫 佳澳 的地方，离那里不远有 拉西亚城 。
ACTS|27|9|航行的日子久了，已经过了禁食的节期，行船又危险， 保罗 就建议，
ACTS|27|10|对众人说：“诸位，我看这次航行，不但货物和船要受损伤，大遭破坏，连我们的性命也难保。”
ACTS|27|11|但百夫长信从船长和船主，不信 保罗 所说的。
ACTS|27|12|且因在这港口不适宜过冬，船上大多数的人都主张开船离开这地方，或者能到 非尼基 去过冬。 非尼基 是 克里特 的一个港口，一面朝西南，一面朝西北。
ACTS|27|13|当南风微微吹起时，他们以为对目的地已有了把握，就起锚，贴近 克里特 开去。
ACTS|27|14|过了不久，有一股叫“友拉革罗”的东北巨风从岛上扑来，
ACTS|27|15|船被风抓住，无法顶风航行，我们只好任它漂流。
ACTS|27|16|我们贴着一个叫 高大 的小岛的背风岸急航，好不容易才保住了救生艇。
ACTS|27|17|既然把救生艇拉上来，他们就用缆索捆绑船底，又恐怕在 赛耳底 浅滩上搁浅，就落了篷，任船漂流。
ACTS|27|18|我们被风浪逼得很急，第二天众人就把货物抛在海里。
ACTS|27|19|第三天，他们又亲手把船上的器具抛弃了。
ACTS|27|20|许多天都没有看到太阳和星辰，又有狂风大浪催逼，我们获救的指望都放弃了。
ACTS|27|21|众人已有好几天没有吃东西， 保罗 就出来站在他们中间，说：“诸位，你们本该听我的话不离开 克里特 岛，就不致遭到这样的损失和破坏。
ACTS|27|22|现在我劝你们放心，除了损失这条船，你们中间没有一人会丧失性命。
ACTS|27|23|因为昨夜，我所属所事奉的上帝的使者站在我旁边，
ACTS|27|24|说：‘ 保罗 ，不要害怕，你必定站在凯撒面前；并且上帝已把安全赐给与你同船的人了。’
ACTS|27|25|所以，诸位可以放心，我信上帝怎样对我说，事情也要怎样成就；
ACTS|27|26|只是我们必须在一个岛上搁浅。”
ACTS|27|27|到了第十四天夜间，船在 亚得里亚海 漂来漂去。约在半夜，水手以为渐近旱地，
ACTS|27|28|就去探测深浅，探得有十二丈 ；稍往前行，又探深浅，探得有九丈。
ACTS|27|29|恐怕我们撞到礁石，他们就从船尾抛下四个锚，盼望天亮。
ACTS|27|30|水手想弃船逃走，把救生艇缒下海里，假装要从船头抛锚的样子。
ACTS|27|31|保罗 对百夫长和士兵说：“这些人若不留在船上，你们就不能获救。”
ACTS|27|32|于是士兵砍断救生艇的绳子，由它漂去。
ACTS|27|33|天快亮的时候， 保罗 劝众人都用餐，说：“你们一直捱饿等候，不吃什么，已经十四天了。
ACTS|27|34|所以我劝你们吃点东西，这是关乎你们获救的，因为你们各人连一根头发也不至于掉落。”
ACTS|27|35|保罗 说了这话，就拿起饼来，在众人面前祝谢了上帝，然后擘开来吃。
ACTS|27|36|于是他们都放心，就吃了。
ACTS|27|37|我们在船上的共有二百七十六个人。
ACTS|27|38|他们吃饱了，为要使船轻一点，就把船上的麦子抛到海里。
ACTS|27|39|天亮的时候，他们不认得那地方，只见一个有岸可登的海湾，就想法子看能不能把船靠岸。
ACTS|27|40|于是他们砍断缆索，把锚丢到海里，同时也松开舵绳，拉起头篷，顺风向着岸行去。
ACTS|27|41|但碰到两水夹流的地方，就搁了浅，船头胶住不动，船尾被浪的猛力冲坏了 。
ACTS|27|42|士兵的意思要把囚犯都杀了，免得有游水脱逃的。
ACTS|27|43|但百夫长要救 保罗 ，不准他们任意而行，就吩咐会游水的，跳下水去，先上岸；
ACTS|27|44|其余的人则用板子或船的碎片上岸。这样，众人都获救，上了岸。
ACTS|28|1|我们既已获救，才知道那岛名叫 马耳他 。
ACTS|28|2|当地人非常友善地接待我们；因为正在下雨，天气又冷，他们就生了火欢迎我们众人。
ACTS|28|3|那时， 保罗 拾起一捆柴，放在火中，有一条毒蛇，因为热的缘故钻了出来，缠住他的手。
ACTS|28|4|当地的人看见那毒蛇悬在他手上，就彼此说：“这人必是个凶手，虽然他从海里获救，天理仍不容他活着。”
ACTS|28|5|保罗 竟把那毒蛇甩在火里，并没有受伤。
ACTS|28|6|当地的人想他快要肿起来，或是忽然倒下死了，但等了好久，见他没有什么异样，就转念说他是个神明。
ACTS|28|7|离那地方不远有一些田产，是岛长 部百流 的。他接纳我们，尽情款待了我们三日。
ACTS|28|8|当时， 部百流 的父亲卧病不起，患了热病和痢疾。 保罗 进去见他，为他祷告按手，治好了他。
ACTS|28|9|从此，岛上其余的病人也都来，得了医治。
ACTS|28|10|他们又多方面尊敬我们，到了开船的时候，又把我们所需用的东西送到船上。
ACTS|28|11|过了三个月，我们上了 亚历山大 的船起航。这船以“ 宙斯 双子”为记，是在那海岛过冬的。
ACTS|28|12|我们到了 叙拉古 ，停泊了三日；
ACTS|28|13|又从那里起锚开船， 来到 利基翁 。过了一天，起了南风，第二天就来到 部丢利 。
ACTS|28|14|我们在那里遇见一些弟兄，他们请我们同住了七天。就这样，我们来到 罗马 。
ACTS|28|15|那里的弟兄们一听见我们的消息，就到 亚比乌 市和 三馆 来迎接我们。 保罗 见了他们，就感谢上帝，越发壮胆。
ACTS|28|16|我们进了 罗马城 ， 保罗 蒙准和那个看守他的兵另住在一处。
ACTS|28|17|过了三天， 保罗 请当地 犹太 人的领袖来。他们来了， 保罗 对他们说：“诸位弟兄，虽然我没有做什么事干犯本国的百姓和我们祖宗的规矩，却在 耶路撒冷 被囚禁，交在 罗马 人的手里。
ACTS|28|18|他们审问了我，有意要释放我，因为在我身上并没有该死的罪状。
ACTS|28|19|但 犹太 人反对，我不得已只好上诉于凯撒，并不是有什么事要控告我本国的百姓。
ACTS|28|20|为这缘故，我请你们来见我当面谈话，我原是为 以色列 人所指望的那位才被这铁链捆绑的。”
ACTS|28|21|他们对他说：“我们并没有接到从 犹太 寄来有关于你的信，也没有弟兄到这里来向我们报告，或说你有什么不好的地方。
ACTS|28|22|但我们愿意听听你的意见，因为我们知道这教门是到处遭人反对的。”
ACTS|28|23|他们和 保罗 约定了日子，就有许多人到他的住处来。 保罗 从早到晚向他们讲解这事，为上帝的国作证，并引 摩西 的律法和先知的书劝导他们信从耶稣。
ACTS|28|24|他所说的话，有的信，有的不信。
ACTS|28|25|他们间彼此不合，就分散了；未散以先， 保罗 说了一句话：“圣灵藉 以赛亚 先知向你们祖宗所说的话是对的。
ACTS|28|26|他说： ‘你去对这百姓说： 你们听了又听，却不明白； 看了又看，却看不清。
ACTS|28|27|因为这百姓的心麻木， 耳朵塞着， 眼睛闭着， 免得眼睛看见， 耳朵听见， 心里明白，回转过来， 我会医治他们。’
ACTS|28|28|所以，你们当知道，上帝这救恩已经传给外邦人；他们会听的。”
ACTS|28|29|
ACTS|28|30|保罗 在自己所租的房子里住了足足两年。凡来见他的人，他都接待，
ACTS|28|31|放胆传讲上帝的国，并教导主耶稣基督的事，没有人禁止。
