2COR|1|1|Павел, волею Божиею Апостол Иисуса Христа, и Тимофей брат, церкви Божией, находящейся в Коринфе, со всеми святыми по всей Ахаии:
2COR|1|2|благодать вам и мир от Бога Отца нашего и Господа Иисуса Христа.
2COR|1|3|Благословен Бог и Отец Господа нашего Иисуса Христа, Отец милосердия и Бог всякого утешения,
2COR|1|4|утешающий нас во всякой скорби нашей, чтобы и мы могли утешать находящихся во всякой скорби тем утешением, которым Бог утешает нас самих!
2COR|1|5|Ибо по мере, как умножаются в нас страдания Христовы, умножается Христом и утешение наше.
2COR|1|6|Скорбим ли мы, [скорбим] для вашего утешения и спасения, которое совершается перенесением тех же страданий, какие и мы терпим.
2COR|1|7|И надежда наша о вас тверда. Утешаемся ли, [утешаемся] для вашего утешения и спасения, зная, что вы участвуете как в страданиях наших, так и в утешении.
2COR|1|8|Ибо мы не хотим оставить вас, братия, в неведении о скорби нашей, бывшей с нами в Асии, потому что мы отягчены были чрезмерно и сверх силы, так что не надеялись остаться в живых.
2COR|1|9|Но сами в себе имели приговор к смерти, для того, чтобы надеяться не на самих себя, но на Бога, воскрешающего мертвых,
2COR|1|10|Который и избавил нас от столь [близкой] смерти, и избавляет, и на Которого надеемся, что и еще избавит,
2COR|1|11|при содействии и вашей молитвы за нас, дабы за дарованное нам, по ходатайству многих, многие возблагодарили за нас.
2COR|1|12|Ибо похвала наша сия есть свидетельство совести нашей, что мы в простоте и богоугодной искренности, не по плотской мудрости, но по благодати Божией, жили в мире, особенно же у вас.
2COR|1|13|И мы пишем вам не иное, как то, что вы читаете или разумеете, и что, как надеюсь, до конца уразумеете,
2COR|1|14|так как вы отчасти и уразумели уже, что мы будем вашею похвалою, равно и вы нашею, в день Господа нашего Иисуса Христа.
2COR|1|15|И в этой уверенности я намеревался придти к вам ранее, чтобы вы вторично получили благодать,
2COR|1|16|и через вас пройти в Македонию, из Македонии же опять придти к вам; а вы проводили бы меня в Иудею.
2COR|1|17|Имея такое намерение, легкомысленно ли я поступил? Или, что я предпринимаю, по плоти предпринимаю, так что у меня то "да, да", то "нет, нет"?
2COR|1|18|Верен Бог, что слово наше к вам не было то "да", то "нет".
2COR|1|19|Ибо Сын Божий, Иисус Христос, проповеданный у вас нами, мною и Силуаном и Тимофеем, не был "да" и "нет"; но в Нем было "да", –
2COR|1|20|ибо все обетования Божии в Нем "да" и в Нем "аминь", – в славу Божию, через нас.
2COR|1|21|Утверждающий же нас с вами во Христе и помазавший нас [есть] Бог,
2COR|1|22|Который и запечатлел нас и дал залог Духа в сердца наши.
2COR|1|23|Бога призываю во свидетели на душу мою, что, щадя вас, я доселе не приходил в Коринф,
2COR|1|24|не потому, будто мы берем власть над верою вашею; но мы споспешествуем радости вашей: ибо верою вы тверды.
2COR|2|1|Итак я рассудил сам в себе не приходить к вам опять с огорчением.
2COR|2|2|Ибо если я огорчаю вас, то кто обрадует меня, как не тот, кто огорчен мною?
2COR|2|3|Это самое и писал я вам, дабы, придя, не иметь огорчения от тех, о которых мне надлежало радоваться: ибо я во всех вас уверен, что моя радость есть [радость] и для всех вас.
2COR|2|4|От великой скорби и стесненного сердца я писал вам со многими слезами, не для того, чтобы огорчить вас, но чтобы вы познали любовь, какую я в избытке имею к вам.
2COR|2|5|Если же кто огорчил, то не меня огорчил, но частью, – чтобы не сказать много, – и всех вас.
2COR|2|6|Для такого довольно сего наказания от многих,
2COR|2|7|так что вам лучше уже простить его и утешить, дабы он не был поглощен чрезмерною печалью.
2COR|2|8|И потому прошу вас оказать ему любовь.
2COR|2|9|Ибо я для того и писал, чтобы узнать на опыте, во всем ли вы послушны.
2COR|2|10|А кого вы в чем прощаете, того и я; ибо и я, если в чем простил кого, простил для вас от лица Христова,
2COR|2|11|чтобы не сделал нам ущерба сатана, ибо нам не безызвестны его умыслы.
2COR|2|12|Придя в Троаду для благовествования о Христе, хотя мне и отверста была дверь Господом,
2COR|2|13|я не имел покоя духу моему, потому что не нашел [там] брата моего Тита; но, простившись с ними, я пошел в Македонию.
2COR|2|14|Но благодарение Богу, Который всегда дает нам торжествовать во Христе и благоухание познания о Себе распространяет нами во всяком месте.
2COR|2|15|Ибо мы Христово благоухание Богу в спасаемых и в погибающих:
2COR|2|16|для одних запах смертоносный на смерть, а для других запах живительный на жизнь. И кто способен к сему?
2COR|2|17|Ибо мы не повреждаем слова Божия, как многие, но проповедуем искренно, как от Бога, пред Богом, во Христе.
2COR|3|1|Неужели нам снова знакомиться с вами? Неужели нужны для нас, как для некоторых, одобрительные письма к вам или от вас?
2COR|3|2|Вы – наше письмо, написанное в сердцах наших, узнаваемое и читаемое всеми человеками;
2COR|3|3|вы показываете собою, что вы – письмо Христово, через служение наше написанное не чернилами, но Духом Бога живаго, не на скрижалях каменных, но на плотяных скрижалях сердца.
2COR|3|4|Такую уверенность мы имеем в Боге через Христа,
2COR|3|5|не потому, чтобы мы сами способны были помыслить что от себя, как бы от себя, но способность наша от Бога.
2COR|3|6|Он дал нам способность быть служителями Нового Завета, не буквы, но духа, потому что буква убивает, а дух животворит.
2COR|3|7|Если же служение смертоносным буквам, начертанное на камнях, было так славно, что сыны Израилевы не могли смотреть на лице Моисеево по причине славы лица его преходящей, –
2COR|3|8|то не гораздо ли более должно быть славно служение духа?
2COR|3|9|Ибо если служение осуждения славно, то тем паче изобилует славою служение оправдания.
2COR|3|10|То прославленное даже не оказывается славным с сей стороны, по причине преимущественной славы [последующего].
2COR|3|11|Ибо, если преходящее славно, тем более славно пребывающее.
2COR|3|12|Имея такую надежду, мы действуем с великим дерзновением,
2COR|3|13|а не так, как Моисей, [который] полагал покрывало на лице свое, чтобы сыны Израилевы не взирали на конец преходящего.
2COR|3|14|Но умы их ослеплены: ибо то же самое покрывало доныне остается неснятым при чтении Ветхого Завета, потому что оно снимается Христом.
2COR|3|15|Доныне, когда они читают Моисея, покрывало лежит на сердце их;
2COR|3|16|но когда обращаются к Господу, тогда это покрывало снимается.
2COR|3|17|Господь есть Дух; а где Дух Господень, там свобода.
2COR|3|18|Мы же все открытым лицем, как в зеркале, взирая на славу Господню, преображаемся в тот же образ от славы в славу, как от Господня Духа.
2COR|4|1|Посему, имея по милости [Божией] такое служение, мы не унываем;
2COR|4|2|но, отвергнув скрытные постыдные [дела], не прибегая к хитрости и не искажая слова Божия, а открывая истину, представляем себя совести всякого человека пред Богом.
2COR|4|3|Если же и закрыто благовествование наше, то закрыто для погибающих,
2COR|4|4|для неверующих, у которых бог века сего ослепил умы, чтобы для них не воссиял свет благовествования о славе Христа, Который есть образ Бога невидимого.
2COR|4|5|Ибо мы не себя проповедуем, но Христа Иисуса, Господа; а мы – рабы ваши для Иисуса,
2COR|4|6|потому что Бог, повелевший из тьмы воссиять свету, озарил наши сердца, дабы просветить [нас] познанием славы Божией в лице Иисуса Христа.
2COR|4|7|Но сокровище сие мы носим в глиняных сосудах, чтобы преизбыточная сила была [приписываема] Богу, а не нам.
2COR|4|8|Мы отовсюду притесняемы, но не стеснены; мы в отчаянных обстоятельствах, но не отчаиваемся;
2COR|4|9|мы гонимы, но не оставлены; низлагаемы, но не погибаем.
2COR|4|10|Всегда носим в теле мертвость Господа Иисуса, чтобы и жизнь Иисусова открылась в теле нашем.
2COR|4|11|Ибо мы живые непрестанно предаемся на смерть ради Иисуса, чтобы и жизнь Иисусова открылась в смертной плоти нашей,
2COR|4|12|так что смерть действует в нас, а жизнь в вас.
2COR|4|13|Но, имея тот же дух веры, как написано: я веровал и потому говорил, и мы веруем, потому и говорим,
2COR|4|14|зная, что Воскресивший Господа Иисуса воскресит через Иисуса и нас и поставит перед [Собою] с вами.
2COR|4|15|Ибо все для вас, дабы обилие благодати тем большую во многих произвело благодарность во славу Божию.
2COR|4|16|Посему мы не унываем; но если внешний наш человек и тлеет, то внутренний со дня на день обновляется.
2COR|4|17|Ибо кратковременное легкое страдание наше производит в безмерном преизбытке вечную славу,
2COR|4|18|когда мы смотрим не на видимое, но на невидимое: ибо видимое временно, а невидимое вечно.
2COR|5|1|Ибо знаем, что, когда земной наш дом, эта хижина, разрушится, мы имеем от Бога жилище на небесах, дом нерукотворенный, вечный.
2COR|5|2|От того мы и воздыхаем, желая облечься в небесное наше жилище;
2COR|5|3|только бы нам и одетым не оказаться нагими.
2COR|5|4|Ибо мы, находясь в этой хижине, воздыхаем под бременем, потому что не хотим совлечься, но облечься, чтобы смертное поглощено было жизнью.
2COR|5|5|На сие самое и создал нас Бог и дал нам залог Духа.
2COR|5|6|Итак мы всегда благодушествуем; и как знаем, что, водворяясь в теле, мы устранены от Господа, –
2COR|5|7|ибо мы ходим верою, а не видением, –
2COR|5|8|то мы благодушествуем и желаем лучше выйти из тела и водвориться у Господа.
2COR|5|9|И потому ревностно стараемся, водворяясь ли, выходя ли, быть Ему угодными;
2COR|5|10|ибо всем нам должно явиться пред судилище Христово, чтобы каждому получить [соответственно тому], что он делал, живя в теле, доброе или худое.
2COR|5|11|Итак, зная страх Господень, мы вразумляем людей, Богу же мы открыты; надеюсь, что открыты и вашим совестям.
2COR|5|12|Не снова представляем себя вам, но даем вам повод хвалиться нами, дабы имели вы [что сказать] тем, которые хвалятся лицем, а не сердцем.
2COR|5|13|Если мы выходим из себя, то для Бога; если же скромны, то для вас.
2COR|5|14|Ибо любовь Христова объемлет нас, рассуждающих так: если один умер за всех, то все умерли.
2COR|5|15|А Христос за всех умер, чтобы живущие уже не для себя жили, но для умершего за них и воскресшего.
2COR|5|16|Потому отныне мы никого не знаем по плоти; если же и знали Христа по плоти, то ныне уже не знаем.
2COR|5|17|Итак, кто во Христе, [тот] новая тварь; древнее прошло, теперь все новое.
2COR|5|18|Все же от Бога, Иисусом Христом примирившего нас с Собою и давшего нам служение примирения,
2COR|5|19|потому что Бог во Христе примирил с Собою мир, не вменяя [людям] преступлений их, и дал нам слово примирения.
2COR|5|20|Итак мы – посланники от имени Христова, и как бы Сам Бог увещевает через нас; от имени Христова просим: примиритесь с Богом.
2COR|5|21|Ибо не знавшего греха Он сделал для нас [жертвою за] грех, чтобы мы в Нем сделались праведными пред Богом.
2COR|6|1|Мы же, как споспешники, умоляем вас, чтобы благодать Божия не тщетно была принята вами.
2COR|6|2|Ибо сказано: во время благоприятное Я услышал тебя и в день спасения помог тебе. Вот, теперь время благоприятное, вот, теперь день спасения.
2COR|6|3|Мы никому ни в чем не полагаем претыкания, чтобы не было порицаемо служение,
2COR|6|4|но во всем являем себя, как служители Божии, в великом терпении, в бедствиях, в нуждах, в тесных обстоятельствах,
2COR|6|5|под ударами, в темницах, в изгнаниях, в трудах, в бдениях, в постах,
2COR|6|6|в чистоте, в благоразумии, в великодушии, в благости, в Духе Святом, в нелицемерной любви,
2COR|6|7|в слове истины, в силе Божией, с оружием правды в правой и левой руке,
2COR|6|8|в чести и бесчестии, при порицаниях и похвалах: нас почитают обманщиками, но мы верны;
2COR|6|9|мы неизвестны, но нас узнают; нас почитают умершими, но вот, мы живы; нас наказывают, но мы не умираем;
2COR|6|10|нас огорчают, а мы всегда радуемся; мы нищи, но многих обогащаем; мы ничего не имеем, но всем обладаем.
2COR|6|11|Уста наши отверсты к вам, Коринфяне, сердце наше расширено.
2COR|6|12|Вам не тесно в нас; но в сердцах ваших тесно.
2COR|6|13|В равное возмездие, – говорю, как детям, – распространитесь и вы.
2COR|6|14|Не преклоняйтесь под чужое ярмо с неверными, ибо какое общение праведности с беззаконием? Что общего у света с тьмою?
2COR|6|15|Какое согласие между Христом и Велиаром? Или какое соучастие верного с неверным?
2COR|6|16|Какая совместность храма Божия с идолами? Ибо вы храм Бога живаго, как сказал Бог: вселюсь в них и буду ходить [в них]; и буду их Богом, и они будут Моим народом.
2COR|6|17|И потому выйдите из среды их и отделитесь, говорит Господь, и не прикасайтесь к нечистому; и Я прииму вас.
2COR|6|18|И буду вам Отцем, и вы будете Моими сынами и дщерями, говорит Господь Вседержитель.
2COR|7|1|Итак, возлюбленные, имея такие обетования, очистим себя от всякой скверны плоти и духа, совершая святыню в страхе Божием.
2COR|7|2|Вместите нас. Мы никого не обидели, никому не повредили, ни от кого не искали корысти.
2COR|7|3|Не в осуждение говорю; ибо я прежде сказал, что вы в сердцах наших, так чтобы вместе и умереть и жить.
2COR|7|4|Я много надеюсь на вас, много хвалюсь вами; я исполнен утешением, преизобилую радостью, при всей скорби нашей.
2COR|7|5|Ибо, когда пришли мы в Македонию, плоть наша не имела никакого покоя, но мы были стеснены отовсюду: отвне – нападения, внутри – страхи.
2COR|7|6|Но Бог, утешающий смиренных, утешил нас прибытием Тита,
2COR|7|7|и не только прибытием его, но и утешением, которым он утешался о вас, пересказывая нам о вашем усердии, о вашем плаче, о вашей ревности по мне, так что я еще более обрадовался.
2COR|7|8|Посему, если я опечалил вас посланием, не жалею, хотя и пожалел было; ибо вижу, что послание то опечалило вас, впрочем на время.
2COR|7|9|Теперь я радуюсь не потому, что вы опечалились, но что вы опечалились к покаянию; ибо опечалились ради Бога, так что нисколько не понесли от нас вреда.
2COR|7|10|Ибо печаль ради Бога производит неизменное покаяние ко спасению, а печаль мирская производит смерть.
2COR|7|11|Ибо то самое, что вы опечалились ради Бога, смотрите, какое произвело в вас усердие, какие извинения, какое негодование [на виновного], какой страх, какое желание, какую ревность, какое взыскание! По всему вы показали себя чистыми в этом деле.
2COR|7|12|Итак, если я писал к вам, то не ради оскорбителя и не ради оскорбленного, но чтобы вам открылось попечение наше о вас пред Богом.
2COR|7|13|Посему мы утешились утешением вашим; а еще более обрадованы мы радостью Тита, что вы все успокоили дух его.
2COR|7|14|Итак я не остался в стыде, если чем–либо о вас похвалился перед ним, но как вам мы говорили все истину, так и перед Титом похвала наша оказалась истинною;
2COR|7|15|и сердце его весьма расположено к вам, при воспоминании о послушании всех вас, как вы приняли его со страхом и трепетом.
2COR|7|16|Итак радуюсь, что во всем могу положиться на вас.
2COR|8|1|Уведомляем вас, братия, о благодати Божией, данной церквам Македонским,
2COR|8|2|ибо они среди великого испытания скорбями преизобилуют радостью; и глубокая нищета их преизбыточествует в богатстве их радушия.
2COR|8|3|Ибо они доброхотны по силам и сверх сил – я свидетель:
2COR|8|4|они весьма убедительно просили нас принять дар и участие [их] в служении святым;
2COR|8|5|и не только то, чего мы надеялись, но они отдали самих себя, во–первых, Господу, [потом] и нам по воле Божией;
2COR|8|6|поэтому мы просили Тита, чтобы он, как начал, так и окончил у вас и это доброе дело.
2COR|8|7|А как вы изобилуете всем: верою и словом, и познанием, и всяким усердием, и любовью вашею к нам, – так изобилуйте и сею добродетелью.
2COR|8|8|Говорю это не в виде повеления, но усердием других испытываю искренность и вашей любви.
2COR|8|9|Ибо вы знаете благодать Господа нашего Иисуса Христа, что Он, будучи богат, обнищал ради вас, дабы вы обогатились Его нищетою.
2COR|8|10|Я даю на это совет: ибо это полезно вам, которые не только начали делать сие, но и желали того еще с прошедшего года.
2COR|8|11|Совершите же теперь самое дело, дабы, чего усердно желали, то и исполнено было по достатку.
2COR|8|12|Ибо если есть усердие, то оно принимается смотря по тому, кто что имеет, а не по тому, чего не имеет.
2COR|8|13|Не [требуется], чтобы другим [было] облегчение, а вам тяжесть, но чтобы была равномерность.
2COR|8|14|Ныне ваш избыток в [восполнение] их недостатка; а после их избыток в [восполнение] вашего недостатка, чтобы была равномерность,
2COR|8|15|как написано: кто собрал много, не имел лишнего; и кто мало, не имел недостатка.
2COR|8|16|Благодарение Богу, вложившему в сердце Титово такое усердие к вам.
2COR|8|17|Ибо, хотя и я просил его, впрочем он, будучи очень усерден, пошел к вам добровольно.
2COR|8|18|С ним послали мы также брата, во всех церквах похваляемого за благовествование,
2COR|8|19|и притом избранного от церквей сопутствовать нам для сего благотворения, которому мы служим во славу Самого Господа и [в] [соответствие] вашему усердию,
2COR|8|20|остерегаясь, чтобы нам не подвергнуться от кого нареканию при таком обилии приношений, вверяемых нашему служению;
2COR|8|21|ибо мы стараемся о добром не только пред Господом, но и пред людьми.
2COR|8|22|Мы послали с ними и брата нашего, которого усердие много раз испытали во многом и который ныне еще усерднее по великой уверенности в вас.
2COR|8|23|Что касается до Тита, это – мой товарищ и сотрудник у вас; а что до братьев наших, это – посланники церквей, слава Христова.
2COR|8|24|Итак перед лицем церквей дайте им доказательство любви вашей и того, что мы [справедливо] хвалимся вами.
2COR|9|1|Для меня впрочем излишне писать вам о вспоможении святым,
2COR|9|2|ибо я знаю усердие ваше и хвалюсь вами перед Македонянами, что Ахаия приготовлена еще с прошедшего года; и ревность ваша поощрила многих.
2COR|9|3|Братьев же послал я для того, чтобы похвала моя о вас не оказалась тщетною в сем случае, но чтобы вы, как я говорил, были приготовлены,
2COR|9|4|[и] чтобы, когда придут со мною Македоняне и найдут вас неготовыми, не остались в стыде мы, – не говорю "вы", – похвалившись с такою уверенностью.
2COR|9|5|Посему я почел за нужное упросить братьев, чтобы они наперед пошли к вам и предварительно озаботились, дабы возвещенное уже благословение ваше было готово, как благословение, а не как побор.
2COR|9|6|При сем скажу: кто сеет скупо, тот скупо и пожнет; а кто сеет щедро, тот щедро и пожнет.
2COR|9|7|Каждый [уделяй] по расположению сердца, не с огорчением и не с принуждением; ибо доброхотно дающего любит Бог.
2COR|9|8|Бог же силен обогатить вас всякою благодатью, чтобы вы, всегда и во всем имея всякое довольство, были богаты на всякое доброе дело,
2COR|9|9|как написано: расточил, раздал нищим; правда его пребывает в век.
2COR|9|10|Дающий же семя сеющему и хлеб в пищу подаст обилие посеянному вами и умножит плоды правды вашей,
2COR|9|11|так чтобы вы всем богаты были на всякую щедрость, которая через нас производит благодарение Богу.
2COR|9|12|Ибо дело служения сего не только восполняет скудость святых, но и производит во многих обильные благодарения Богу;
2COR|9|13|ибо, видя опыт сего служения, они прославляют Бога за покорность исповедуемому вами Евангелию Христову и за искреннее общение с ними и со всеми,
2COR|9|14|молясь за вас, по расположению к вам, за преизбыточествующую в вас благодать Божию.
2COR|9|15|Благодарение Богу за неизреченный дар Его!
2COR|10|1|Я же, Павел, который лично между вами скромен, а заочно против вас отважен, убеждаю вас кротостью и снисхождением Христовым.
2COR|10|2|Прошу, чтобы мне по пришествии моем не прибегать к той твердой смелости, которую думаю употребить против некоторых, помышляющих о нас, что мы поступаем по плоти.
2COR|10|3|Ибо мы, ходя во плоти, не по плоти воинствуем.
2COR|10|4|Оружия воинствования нашего не плотские, но сильные Богом на разрушение твердынь: [ими] ниспровергаем замыслы
2COR|10|5|и всякое превозношение, восстающее против познания Божия, и пленяем всякое помышление в послушание Христу,
2COR|10|6|и готовы наказать всякое непослушание, когда ваше послушание исполнится.
2COR|10|7|На личность ли смотрите? Кто уверен в себе, что он Христов, тот сам по себе суди, что, как он Христов, так и мы Христовы.
2COR|10|8|Ибо если бы я и более стал хвалиться нашею властью, которую Господь дал нам к созиданию, а не к расстройству вашему, то не остался бы в стыде.
2COR|10|9|Впрочем, да не покажется, что я устрашаю вас [только] посланиями.
2COR|10|10|Так как [некто] говорит: в посланиях он строг и силен, а в личном присутствии слаб, и речь [его] незначительна, –
2COR|10|11|такой пусть знает, что, каковы мы на словах в посланиях заочно, таковы и на деле лично.
2COR|10|12|Ибо мы не смеем сопоставлять или сравнивать себя с теми, которые сами себя выставляют: они измеряют себя самими собою и сравнивают себя с собою неразумно.
2COR|10|13|А мы не без меры хвалиться будем, но по мере удела, какой назначил нам Бог в такую меру, чтобы достигнуть и до вас.
2COR|10|14|Ибо мы не напрягаем себя, как не достигшие до вас, потому что достигли и до вас благовествованием Христовым.
2COR|10|15|Мы не без меры хвалимся, не чужими трудами, но надеемся, с возрастанием веры вашей, с избытком увеличить в вас удел наш,
2COR|10|16|так чтобы и далее вас проповедывать Евангелие, а не хвалиться готовым в чужом уделе.
2COR|10|17|Хвалящийся хвались о Господе.
2COR|10|18|Ибо не тот достоин, кто сам себя хвалит, но кого хвалит Господь.
2COR|11|1|О, если бы вы несколько были снисходительны к моему неразумию! Но вы и снисходите ко мне.
2COR|11|2|Ибо я ревную о вас ревностью Божиею; потому что я обручил вас единому мужу, чтобы представить Христу чистою девою.
2COR|11|3|Но боюсь, чтобы, как змий хитростью своею прельстил Еву, так и ваши умы не повредились, [уклонившись] от простоты во Христе.
2COR|11|4|Ибо если бы кто, придя, начал проповедывать другого Иисуса, которого мы не проповедывали, или если бы вы получили иного Духа, которого не получили, или иное благовестие, которого не принимали, – то вы были бы очень снисходительны [к тому].
2COR|11|5|Но я думаю, что у меня ни в чем нет недостатка против высших Апостолов:
2COR|11|6|хотя я и невежда в слове, но не в познании. Впрочем мы во всем совершенно известны вам.
2COR|11|7|Согрешил ли я тем, что унижал себя, чтобы возвысить вас, потому что безмездно проповедывал вам Евангелие Божие?
2COR|11|8|Другим церквам я причинял издержки, получая [от них] содержание для служения вам; и, будучи у вас, хотя терпел недостаток, никому не докучал,
2COR|11|9|ибо недостаток мой восполнили братия, пришедшие из Македонии; да и во всем я старался и постараюсь не быть вам в тягость.
2COR|11|10|По истине Христовой во мне [скажу], что похвала сия не отнимется у меня в странах Ахаии.
2COR|11|11|Почему же [так поступаю]? Потому ли, что не люблю вас? Богу известно! Но как поступаю, так и буду поступать,
2COR|11|12|чтобы не дать повода ищущим повода, дабы они, чем хвалятся, в том оказались [такими же], как и мы.
2COR|11|13|Ибо таковые лжеапостолы, лукавые делатели, принимают вид Апостолов Христовых.
2COR|11|14|И неудивительно: потому что сам сатана принимает вид Ангела света,
2COR|11|15|а потому не великое дело, если и служители его принимают вид служителей правды; но конец их будет по делам их.
2COR|11|16|Еще скажу: не почти кто–нибудь меня неразумным; а если не так, то примите меня, хотя как неразумного, чтобы и мне сколько–нибудь похвалиться.
2COR|11|17|Что скажу, то скажу не в Господе, но как бы в неразумии при такой отважности на похвалу.
2COR|11|18|Как многие хвалятся по плоти, то и я буду хвалиться.
2COR|11|19|Ибо вы, люди разумные, охотно терпите неразумных:
2COR|11|20|вы терпите, когда кто вас порабощает, когда кто объедает, когда кто обирает, когда кто превозносится, когда кто бьет вас в лицо.
2COR|11|21|К стыду говорю, что [на это] у нас недоставало сил. А если кто смеет [хвалиться] чем–либо, то (скажу по неразумию) смею и я.
2COR|11|22|Они Евреи? и я. Израильтяне? и я. Семя Авраамово? и я.
2COR|11|23|Христовы служители? (в безумии говорю:) я больше. Я гораздо более [был] в трудах, безмерно в ранах, более в темницах и многократно при смерти.
2COR|11|24|От Иудеев пять раз дано мне было по сорока [ударов] без одного;
2COR|11|25|три раза меня били палками, однажды камнями побивали, три раза я терпел кораблекрушение, ночь и день пробыл во глубине [морской];
2COR|11|26|много раз [был] в путешествиях, в опасностях на реках, в опасностях от разбойников, в опасностях от единоплеменников, в опасностях от язычников, в опасностях в городе, в опасностях в пустыне, в опасностях на море, в опасностях между лжебратиями,
2COR|11|27|в труде и в изнурении, часто в бдении, в голоде и жажде, часто в посте, на стуже и в наготе.
2COR|11|28|Кроме посторонних [приключений], у меня ежедневно стечение [людей], забота о всех церквах.
2COR|11|29|Кто изнемогает, с кем бы и я не изнемогал? Кто соблазняется, за кого бы я не воспламенялся?
2COR|11|30|Если должно мне хвалиться, то буду хвалиться немощью моею.
2COR|11|31|Бог и Отец Господа нашего Иисуса Христа, благословенный во веки, знает, что я не лгу.
2COR|11|32|В Дамаске областной правитель царя Ареты стерег город Дамаск, чтобы схватить меня;
2COR|11|33|и я в корзине был спущен из окна по стене и избежал его рук.
2COR|12|1|Не полезно хвалиться мне, ибо я приду к видениям и откровениям Господним.
2COR|12|2|Знаю человека во Христе, который назад тому четырнадцать лет (в теле ли – не знаю, вне ли тела – не знаю: Бог знает) восхищен был до третьего неба.
2COR|12|3|И знаю о таком человеке ([только] не знаю – в теле, или вне тела: Бог знает),
2COR|12|4|что он был восхищен в рай и слышал неизреченные слова, которых человеку нельзя пересказать.
2COR|12|5|Таким [человеком] могу хвалиться; собою же не похвалюсь, разве только немощами моими.
2COR|12|6|Впрочем, если захочу хвалиться, не буду неразумен, потому что скажу истину; но я удерживаюсь, чтобы кто не подумал о мне более, нежели сколько во мне видит или слышит от меня.
2COR|12|7|И чтобы я не превозносился чрезвычайностью откровений, дано мне жало в плоть, ангел сатаны, удручать меня, чтобы я не превозносился.
2COR|12|8|Трижды молил я Господа о том, чтобы удалил его от меня.
2COR|12|9|Но [Господь] сказал мне: "довольно для тебя благодати Моей, ибо сила Моя совершается в немощи". И потому я гораздо охотнее буду хвалиться своими немощами, чтобы обитала во мне сила Христова.
2COR|12|10|Посему я благодушествую в немощах, в обидах, в нуждах, в гонениях, в притеснениях за Христа, ибо, когда я немощен, тогда силен.
2COR|12|11|Я дошел до неразумия, хвалясь; вы меня [к сему] принудили. Вам бы надлежало хвалить меня, ибо у меня ни в чем нет недостатка против высших Апостолов, хотя я и ничто.
2COR|12|12|Признаки Апостола оказались перед вами всяким терпением, знамениями, чудесами и силами.
2COR|12|13|Ибо чего у вас недостает перед прочими церквами, разве только того, что сам я не был вам в тягость? Простите мне такую вину.
2COR|12|14|Вот, в третий раз я готов идти к вам, и не буду отягощать вас, ибо я ищу не вашего, а вас. Не дети должны собирать имение для родителей, но родители для детей.
2COR|12|15|Я охотно буду издерживать [свое] и истощать себя за души ваши, несмотря на то, что, чрезвычайно любя вас, я менее любим вами.
2COR|12|16|Положим, [что] сам я не обременял вас, но, будучи хитр, лукавством брал с вас.
2COR|12|17|Но пользовался ли я [чем] от вас через кого–нибудь из тех, кого посылал к вам?
2COR|12|18|Я упросил Тита и послал с ним одного из братьев: Тит воспользовался ли чем от вас? Не в одном ли духе мы действовали? Не одним ли путем ходили?
2COR|12|19|Не думаете ли еще, что мы [только] оправдываемся перед вами? Мы говорим пред Богом, во Христе, и все это, возлюбленные, к вашему назиданию.
2COR|12|20|Ибо я опасаюсь, чтобы мне, по пришествии моем, не найти вас такими, какими не желаю, также чтобы и вам не найти меня таким, каким не желаете: чтобы [не найти у вас] раздоров, зависти, гнева, ссор, клевет, ябед, гордости, беспорядков,
2COR|12|21|чтобы опять, когда приду, не уничижил меня у вас Бог мой и [чтобы] не оплакивать мне многих, которые согрешили прежде и не покаялись в нечистоте, блудодеянии и непотребстве, какое делали.
2COR|13|1|В третий уже раз иду к вам. При устах двух или трех свидетелей будет твердо всякое слово.
2COR|13|2|Я предварял и предваряю, как бы находясь [у вас] во второй раз, и теперь, отсутствуя, пишу прежде согрешившим и всем прочим, что, когда опять приду, не пощажу.
2COR|13|3|Вы ищете доказательства на то, Христос ли говорит во мне: Он не бессилен для вас, но силен в вас.
2COR|13|4|Ибо, хотя Он и распят в немощи, но жив силою Божиею; и мы также, [хотя] немощны в Нем, но будем живы с Ним силою Божиею в вас.
2COR|13|5|Испытывайте самих себя, в вере ли вы; самих себя исследывайте. Или вы не знаете самих себя, что Иисус Христос в вас? Разве только вы не то, чем должны быть.
2COR|13|6|О нас же, надеюсь, узнаете, что мы то, чем быть должны.
2COR|13|7|Молим Бога, чтобы вы не делали никакого зла, не для того, чтобы нам показаться, чем должны быть; но чтобы вы делали добро, хотя бы мы казались и не тем, чем должны быть.
2COR|13|8|Ибо мы не сильны против истины, но сильны за истину.
2COR|13|9|Мы радуемся, когда мы немощны, а вы сильны; о сем–то и молимся, о вашем совершенстве.
2COR|13|10|Для того я и пишу сие в отсутствии, чтобы в присутствии не употребить строгости по власти, данной мне Господом к созиданию, а не к разорению.
2COR|13|11|Впрочем, братия, радуйтесь, усовершайтесь, утешайтесь, будьте единомысленны, мирны, – и Бог любви и мира будет с вами.
2COR|13|12|Приветствуйте друг друга лобзанием святым. Приветствуют вас все святые.
2COR|13|13|Благодать Господа нашего Иисуса Христа, и любовь Бога Отца, и общение Святаго Духа со всеми вами. Аминь.
