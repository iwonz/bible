JONAH|1|1|The word of the LORD came to Jonah son of Amittai:
JONAH|1|2|"Go to the great city of Nineveh and preach against it, because its wickedness has come up before me."
JONAH|1|3|But Jonah ran away from the LORD and headed for Tarshish. He went down to Joppa, where he found a ship bound for that port. After paying the fare, he went aboard and sailed for Tarshish to flee from the LORD.
JONAH|1|4|Then the LORD sent a great wind on the sea, and such a violent storm arose that the ship threatened to break up.
JONAH|1|5|All the sailors were afraid and each cried out to his own god. And they threw the cargo into the sea to lighten the ship. But Jonah had gone below deck, where he lay down and fell into a deep sleep.
JONAH|1|6|The captain went to him and said, "How can you sleep? Get up and call on your god! Maybe he will take notice of us, and we will not perish."
JONAH|1|7|Then the sailors said to each other, "Come, let us cast lots to find out who is responsible for this calamity." They cast lots and the lot fell on Jonah.
JONAH|1|8|So they asked him, "Tell us, who is responsible for making all this trouble for us? What do you do? Where do you come from? What is your country? From what people are you?"
JONAH|1|9|He answered, "I am a Hebrew and I worship the LORD, the God of heaven, who made the sea and the land."
JONAH|1|10|This terrified them and they asked, "What have you done?" (They knew he was running away from the LORD, because he had already told them so.)
JONAH|1|11|The sea was getting rougher and rougher. So they asked him, "What should we do to you to make the sea calm down for us?"
JONAH|1|12|"Pick me up and throw me into the sea," he replied, "and it will become calm. I know that it is my fault that this great storm has come upon you."
JONAH|1|13|Instead, the men did their best to row back to land. But they could not, for the sea grew even wilder than before.
JONAH|1|14|Then they cried to the LORD, "O LORD, please do not let us die for taking this man's life. Do not hold us accountable for killing an innocent man, for you, O LORD, have done as you pleased."
JONAH|1|15|Then they took Jonah and threw him overboard, and the raging sea grew calm.
JONAH|1|16|At this the men greatly feared the LORD, and they offered a sacrifice to the LORD and made vows to him.
JONAH|1|17|But the LORD provided a great fish to swallow Jonah, and Jonah was inside the fish three days and three nights.
JONAH|2|1|From inside the fish Jonah prayed to the LORD his God.
JONAH|2|2|He said: "In my distress I called to the LORD, and he answered me. From the depths of the grave I called for help, and you listened to my cry.
JONAH|2|3|You hurled me into the deep, into the very heart of the seas, and the currents swirled about me; all your waves and breakers swept over me.
JONAH|2|4|I said, 'I have been banished from your sight; yet I will look again toward your holy temple.'
JONAH|2|5|The engulfing waters threatened me, the deep surrounded me; seaweed was wrapped around my head.
JONAH|2|6|To the roots of the mountains I sank down; the earth beneath barred me in forever. But you brought my life up from the pit, O LORD my God.
JONAH|2|7|"When my life was ebbing away, I remembered you, LORD, and my prayer rose to you, to your holy temple.
JONAH|2|8|"Those who cling to worthless idols forfeit the grace that could be theirs.
JONAH|2|9|But I, with a song of thanksgiving, will sacrifice to you. What I have vowed I will make good. Salvation comes from the LORD."
JONAH|2|10|And the LORD commanded the fish, and it vomited Jonah onto dry land.
JONAH|3|1|Then the word of the LORD came to Jonah a second time:
JONAH|3|2|"Go to the great city of Nineveh and proclaim to it the message I give you."
JONAH|3|3|Jonah obeyed the word of the LORD and went to Nineveh. Now Nineveh was a very important city-a visit required three days.
JONAH|3|4|On the first day, Jonah started into the city. He proclaimed: "Forty more days and Nineveh will be overturned."
JONAH|3|5|The Ninevites believed God. They declared a fast, and all of them, from the greatest to the least, put on sackcloth.
JONAH|3|6|When the news reached the king of Nineveh, he rose from his throne, took off his royal robes, covered himself with sackcloth and sat down in the dust.
JONAH|3|7|Then he issued a proclamation in Nineveh: "By the decree of the king and his nobles: Do not let any man or beast, herd or flock, taste anything; do not let them eat or drink.
JONAH|3|8|But let man and beast be covered with sackcloth. Let everyone call urgently on God. Let them give up their evil ways and their violence.
JONAH|3|9|Who knows? God may yet relent and with compassion turn from his fierce anger so that we will not perish."
JONAH|3|10|When God saw what they did and how they turned from their evil ways, he had compassion and did not bring upon them the destruction he had threatened.
JONAH|4|1|But Jonah was greatly displeased and became angry.
JONAH|4|2|He prayed to the LORD, "O LORD, is this not what I said when I was still at home? That is why I was so quick to flee to Tarshish. I knew that you are a gracious and compassionate God, slow to anger and abounding in love, a God who relents from sending calamity.
JONAH|4|3|Now, O LORD, take away my life, for it is better for me to die than to live."
JONAH|4|4|But the LORD replied, "Have you any right to be angry?"
JONAH|4|5|Jonah went out and sat down at a place east of the city. There he made himself a shelter, sat in its shade and waited to see what would happen to the city.
JONAH|4|6|Then the LORD God provided a vine and made it grow up over Jonah to give shade for his head to ease his discomfort, and Jonah was very happy about the vine.
JONAH|4|7|But at dawn the next day God provided a worm, which chewed the vine so that it withered.
JONAH|4|8|When the sun rose, God provided a scorching east wind, and the sun blazed on Jonah's head so that he grew faint. He wanted to die, and said, "It would be better for me to die than to live."
JONAH|4|9|But God said to Jonah, "Do you have a right to be angry about the vine?I do," he said. "I am angry enough to die."
JONAH|4|10|But the LORD said, "You have been concerned about this vine, though you did not tend it or make it grow. It sprang up overnight and died overnight.
JONAH|4|11|But Nineveh has more than a hundred and twenty thousand people who cannot tell their right hand from their left, and many cattle as well. Should I not be concerned about that great city?"
