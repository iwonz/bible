ECCL|1|1|verba Ecclesiastes filii David regis Hierusalem
ECCL|1|2|vanitas vanitatum dixit Ecclesiastes vanitas vanitatum omnia vanitas
ECCL|1|3|quid habet amplius homo de universo labore suo quod laborat sub sole
ECCL|1|4|generatio praeterit et generatio advenit terra vero in aeternum stat
ECCL|1|5|oritur sol et occidit et ad locum suum revertitur ibique renascens
ECCL|1|6|gyrat per meridiem et flectitur ad aquilonem lustrans universa circuitu pergit spiritus et in circulos suos regreditur
ECCL|1|7|omnia flumina intrant mare et mare non redundat ad locum unde exeunt flumina revertuntur ut iterum fluant
ECCL|1|8|cunctae res difficiles non potest eas homo explicare sermone non saturatur oculus visu nec auris impletur auditu
ECCL|1|9|quid est quod fuit ipsum quod futurum est quid est quod factum est ipsum quod fiendum est
ECCL|1|10|nihil sub sole novum nec valet quisquam dicere ecce hoc recens est iam enim praecessit in saeculis quae fuerunt ante nos
ECCL|1|11|non est priorum memoria sed nec eorum quidem quae postea futura sunt erit recordatio apud eos qui futuri sunt in novissimo
ECCL|1|12|ego Ecclesiastes fui rex Israhel in Hierusalem
ECCL|1|13|et proposui in animo meo quaerere et investigare sapienter de omnibus quae fiunt sub sole hanc occupationem pessimam dedit Deus filiis hominum ut occuparentur in ea
ECCL|1|14|vidi quae fiunt cuncta sub sole et ecce universa vanitas et adflictio spiritus
ECCL|1|15|perversi difficile corriguntur et stultorum infinitus est numerus
ECCL|1|16|locutus sum in corde meo dicens ecce magnus effectus sum et praecessi sapientia omnes qui fuerunt ante me in Hierusalem et mens mea contemplata est multa sapienter et didicit
ECCL|1|17|dedique cor meum ut scirem prudentiam atque doctrinam erroresque et stultitiam et agnovi quod in his quoque esset labor et adflictio spiritus
ECCL|1|18|eo quod in multa sapientia multa sit indignatio et qui addit scientiam addat et laborem
ECCL|2|1|dixi ego in corde meo vadam et affluam deliciis et fruar bonis et vidi quod hoc quoque esset vanitas
ECCL|2|2|risum reputavi errorem et gaudio dixi quid frustra deciperis
ECCL|2|3|cogitavi in corde meo abstrahere a vino carnem meam ut animum meum transferrem ad sapientiam devitaremque stultitiam donec viderem quid esset utile filiis hominum quod facto opus est sub sole numero dierum vitae suae
ECCL|2|4|magnificavi opera mea aedificavi mihi domos plantavi vineas
ECCL|2|5|feci hortos et pomeria et consevi ea cuncti generis arboribus
ECCL|2|6|extruxi mihi piscinas aquarum ut inrigarem silvam lignorum germinantium
ECCL|2|7|possedi servos et ancillas multamque familiam habui armenta quoque et magnos ovium greges ultra omnes qui fuerunt ante me in Hierusalem
ECCL|2|8|coacervavi mihi argentum et aurum et substantias regum ac provinciarum feci mihi cantores et cantrices et delicias filiorum hominum scyphos et urceos in ministerio ad vina fundenda
ECCL|2|9|et supergressus sum opibus omnes qui fuerunt ante me in Hierusalem sapientia quoque perseveravit mecum
ECCL|2|10|et omnia quae desideraverunt oculi mei non negavi eis nec prohibui cor quin omni voluptate frueretur et oblectaret se in his quae paraveram et hanc ratus sum partem meam si uterer labore meo
ECCL|2|11|cumque me convertissem ad universa opera quae fecerant manus meae et ad labores in quibus frustra sudaveram vidi in omnibus vanitatem et adflictionem animi et nihil permanere sub sole
ECCL|2|12|transivi ad contemplandam sapientiam erroresque et stultitiam quid est inquam homo ut sequi possit regem factorem suum
ECCL|2|13|et vidi quia tantum praecederet sapientia stultitiam quantum differt lux tenebris
ECCL|2|14|sapientis oculi in capite eius stultus in tenebris ambulat et didici quod unus utriusque esset interitus
ECCL|2|15|et dixi in corde meo si unus et stulti et meus occasus erit quid mihi prodest quod maiorem sapientiae dedi operam locutusque cum mente mea animadverti quod hoc quoque esset vanitas
ECCL|2|16|non enim erit memoria sapientis similiter ut stulti in perpetuum et futura tempora oblivione cuncta pariter obruent moritur doctus similiter et indoctus
ECCL|2|17|et idcirco taeduit me vitae meae videntem mala esse universa sub sole et cuncta vanitatem atque adflictionem spiritus
ECCL|2|18|rursum detestatus sum omnem industriam meam quae sub sole studiosissime laboravi habiturus heredem post me
ECCL|2|19|quem ignoro utrum sapiens an stultus futurus sit et dominabitur in laboribus meis quibus desudavi et sollicitus fui et est quicquam tam vanum
ECCL|2|20|unde cessavi renuntiavitque cor meum ultra laborare sub sole
ECCL|2|21|nam cum alius laboret in sapientia et doctrina et sollicitudine homini otioso quaesita dimittit et hoc ergo vanitas et magnum malum
ECCL|2|22|quid enim proderit homini de universo labore suo et adflictione spiritus qua sub sole cruciatus est
ECCL|2|23|cuncti dies eius doloribus et aerumnis pleni sunt nec per noctem mente requiescit et haec non vanitas est
ECCL|2|24|nonne melius est comedere et bibere et ostendere animae suae bona de laboribus suis et hoc de manu Dei est
ECCL|2|25|quis ita vorabit et deliciis affluet ut ego
ECCL|2|26|homini bono in conspectu suo dedit Deus sapientiam et scientiam et laetitiam peccatori autem dedit adflictionem et curam superfluam ut addat et congreget et tradat ei qui placuit Deo sed et hoc vanitas et cassa sollicitudo mentis
ECCL|3|1|omnia tempus habent et suis spatiis transeunt universa sub caelo
ECCL|3|2|tempus nascendi et tempus moriendi tempus plantandi et tempus evellendi quod plantatum est
ECCL|3|3|tempus occidendi et tempus sanandi tempus destruendi et tempus aedificandi
ECCL|3|4|tempus flendi et tempus ridendi tempus plangendi et tempus saltandi
ECCL|3|5|tempus spargendi lapides et tempus colligendi tempus amplexandi et tempus longe fieri a conplexibus
ECCL|3|6|tempus adquirendi et tempus perdendi tempus custodiendi et tempus abiciendi
ECCL|3|7|tempus scindendi et tempus consuendi tempus tacendi et tempus loquendi
ECCL|3|8|tempus dilectionis et tempus odii tempus belli et tempus pacis
ECCL|3|9|quid habet amplius homo de labore suo
ECCL|3|10|vidi adflictionem quam dedit Deus filiis hominum ut distendantur in ea
ECCL|3|11|cuncta fecit bona in tempore suo et mundum tradidit disputationi eorum ut non inveniat homo opus quod operatus est Deus ab initio usque ad finem
ECCL|3|12|et cognovi quod non esset melius nisi laetari et facere bene in vita sua
ECCL|3|13|omnis enim homo qui comedit et bibit et videt bonum de labore suo hoc donum Dei est
ECCL|3|14|didici quod omnia opera quae fecit Deus perseverent in perpetuum non possumus eis quicquam addere nec auferre quae fecit Deus ut timeatur
ECCL|3|15|quod factum est ipsum permanet quae futura sunt iam fuerunt et Deus instaurat quod abiit
ECCL|3|16|vidi sub sole in loco iudicii impietatem et in loco iustitiae iniquitatem
ECCL|3|17|et dixi in corde meo iustum et impium iudicabit Deus et tempus omni rei tunc erit
ECCL|3|18|dixi in corde meo de filiis hominum ut probaret eos Deus et ostenderet similes esse bestiis
ECCL|3|19|idcirco unus interitus est hominis et iumentorum et aequa utriusque condicio sicut moritur homo sic et illa moriuntur similiter spirant omnia et nihil habet homo iumento amplius cuncta subiacent vanitati
ECCL|3|20|et omnia pergunt ad unum locum de terra facta sunt et in terram pariter revertentur
ECCL|3|21|quis novit si spiritus filiorum Adam ascendat sursum et si spiritus iumentorum descendat deorsum
ECCL|3|22|et deprehendi nihil esse melius quam laetari hominem in opere suo et hanc esse partem illius quis enim eum adducet ut post se futura cognoscat
ECCL|4|1|verti me ad alia et vidi calumnias quae sub sole geruntur et lacrimas innocentum et consolatorem neminem nec posse resistere eorum violentiae cunctorum auxilio destitutos
ECCL|4|2|et laudavi magis mortuos quam viventes
ECCL|4|3|et feliciorem utroque iudicavi qui necdum natus est nec vidit mala quae sub sole fiunt
ECCL|4|4|rursum contemplatus omnes labores hominum et industrias animadverti patere invidiae proximi et in hoc ergo vanitas et cura superflua est
ECCL|4|5|stultus conplicat manus suas et comedit carnes suas dicens
ECCL|4|6|melior est pugillus cum requie quam plena utraque manus cum labore et adflictione animi
ECCL|4|7|considerans repperi et aliam vanitatem sub sole
ECCL|4|8|unus est et secundum non habet non filium non fratrem et tamen laborare non cessat nec satiantur oculi eius divitiis nec recogitat dicens cui laboro et fraudo animam meam bonis in hoc quoque vanitas est et adflictio pessima
ECCL|4|9|melius ergo est duos simul esse quam unum habent enim emolumentum societatis suae
ECCL|4|10|si unus ceciderit ab altero fulcietur vae soli quia cum ruerit non habet sublevantem
ECCL|4|11|et si dormierint duo fovebuntur mutuo unus quomodo calefiet
ECCL|4|12|et si quispiam praevaluerit contra unum duo resistent ei funiculus triplex difficile rumpitur
ECCL|4|13|melior est puer pauper et sapiens rege sene et stulto qui nescit providere in posterum
ECCL|4|14|quod et de carcere catenisque interdum quis egrediatur ad regnum et alius natus in regno inopia consumatur
ECCL|4|15|vidi cunctos viventes qui ambulant sub sole cum adulescente secundo qui consurgit pro eo
ECCL|4|16|infinitus numerus est populi omnium qui fuerunt ante eum et qui postea futuri sunt non laetabuntur in eo sed et hoc vanitas et adflictio spiritus
ECCL|4|17|custodi pedem tuum ingrediens domum Dei multo enim melior est oboedientia quam stultorum victimae qui nesciunt quid faciant mali
ECCL|5|1|ne temere quid loquaris neque cor tuum sit velox ad proferendum sermonem coram Deo Deus enim in caelo et tu super terram idcirco sint pauci sermones tui
ECCL|5|2|multas curas sequuntur somnia et in multis sermonibus invenitur stultitia
ECCL|5|3|si quid vovisti Deo ne moreris reddere displicet enim ei infidelis et stulta promissio sed quodcumque voveris redde
ECCL|5|4|multoque melius est non vovere quam post votum promissa non conplere
ECCL|5|5|ne dederis os tuum ut peccare faciat carnem tuam neque dicas coram angelo non est providentia ne forte iratus Deus super sermone tuo dissipet cuncta opera manuum tuarum
ECCL|5|6|ubi multa sunt somnia plurimae vanitates et sermones innumeri tu vero Deum time
ECCL|5|7|si videris calumnias egenorum et violenta iudicia et subverti iustitiam in provincia non mireris super hoc negotio quia excelso alius excelsior est et super hos quoque eminentiores sunt alii
ECCL|5|8|et insuper universae terrae rex imperat servienti
ECCL|5|9|avarus non implebitur pecunia et qui amat divitias fructus non capiet ex eis et hoc ergo vanitas
ECCL|5|10|ubi multae sunt opes multi et qui comedant eas et quid prodest possessori nisi quod cernit divitias oculis suis
ECCL|5|11|dulcis est somnus operanti sive parum sive multum comedat saturitas autem divitis non sinit dormire eum
ECCL|5|12|est et alia infirmitas pessima quam vidi sub sole divitiae conservatae in malum domini sui
ECCL|5|13|pereunt enim in adflictione pessima generavit filium qui in summa egestate erit
ECCL|5|14|sicut egressus est nudus de utero matris suae sic revertetur et nihil auferet secum de labore suo
ECCL|5|15|miserabilis prorsus infirmitas quomodo venit sic revertetur quid ergo prodest ei quod laboravit in ventum
ECCL|5|16|cunctis diebus vitae suae comedit in tenebris et in curis multis et in aerumna atque tristitia
ECCL|5|17|hoc itaque mihi visum est bonum ut comedat quis et bibat et fruatur laetitia ex labore suo quod laboravit ipse sub sole numerum dierum vitae suae quos dedit ei Deus et haec est pars illius
ECCL|5|18|et omni homini cui dedit Deus divitias atque substantiam potestatemque ei tribuit ut comedat ex eis et fruatur parte sua et laetetur de labore suo hoc est donum Dei
ECCL|5|19|non enim satis recordabitur dierum vitae suae eo quod Deus occupet deliciis cor eius
ECCL|6|1|est et aliud malum quod vidi sub sole et quidem frequens apud homines
ECCL|6|2|vir cui dedit Deus divitias et substantiam et honorem et nihil deest animae eius ex omnibus quae desiderat nec tribuit ei potestatem Deus ut comedat ex eo sed homo extraneus vorabit illud hoc vanitas et magna miseria est
ECCL|6|3|si genuerit quispiam centum et vixerit multos annos et plures dies aetatis habuerit et anima illius non utatur bonis substantiae suae sepulturaque careat de hoc ego pronuntio quod melior illo sit abortivus
ECCL|6|4|frustra enim venit et pergit ad tenebras et oblivione delebitur nomen eius
ECCL|6|5|non vidit solem neque cognovit distantiam boni et mali
ECCL|6|6|etiam si duobus milibus annis vixerit et non fuerit perfruitus bonis nonne ad unum locum properant omnia
ECCL|6|7|omnis labor hominis in ore eius sed anima illius non impletur
ECCL|6|8|quid habet amplius sapiens ab stulto et quid pauper nisi ut pergat illuc ubi est vita
ECCL|6|9|melius est videre quod cupias quam desiderare quod nescias sed et hoc vanitas est et praesumptio spiritus
ECCL|6|10|qui futurus est iam vocatum est nomen eius et scitur quod homo sit et non possit contra fortiorem se in iudicio contendere
ECCL|6|11|verba sunt plurima multa in disputando habentia vanitatem
ECCL|7|1|quid necesse est homini maiora se quaerere cum ignoret quid conducat sibi in vita sua numero dierum peregrinationis suae et tempore quo velut umbra praeterit aut quis ei poterit indicare quid post eum futurum sub sole sit
ECCL|7|2|melius est nomen bonum quam unguenta pretiosa et dies mortis die nativitatis
ECCL|7|3|melius est ire ad domum luctus quam ad domum convivii in illa enim finis cunctorum admonetur hominum et vivens cogitat quid futurum sit
ECCL|7|4|melior est ira risu quia per tristitiam vultus corrigitur animus delinquentis
ECCL|7|5|cor sapientium ubi tristitia est et cor stultorum ubi laetitia
ECCL|7|6|melius est a sapiente corripi quam stultorum adulatione decipi
ECCL|7|7|quia sicut sonitus spinarum ardentium sub olla sic risus stulti sed et hoc vanitas
ECCL|7|8|calumnia conturbat sapientem et perdet robur cordis illius
ECCL|7|9|melior est finis orationis quam principium melior est patiens arrogante
ECCL|7|10|ne velox sis ad irascendum quia ira in sinu stulti requiescit
ECCL|7|11|ne dicas quid putas causae est quod priora tempora meliora fuere quam nunc sunt stulta est enim huiuscemodi interrogatio
ECCL|7|12|utilior est sapientia cum divitiis et magis prodest videntibus solem
ECCL|7|13|sicut enim protegit sapientia sic protegit pecunia hoc autem plus habet eruditio et sapientia quod vitam tribuunt possessori suo
ECCL|7|14|considera opera Dei quod nemo possit corrigere quem ille despexerit
ECCL|7|15|in die bona fruere bonis et malam diem praecave sicut enim hanc sic et illam fecit Deus ut non inveniat homo contra eum iustas querimonias
ECCL|7|16|haec quoque vidi in diebus vanitatis meae iustus perit in iustitia sua et impius multo vivit tempore in malitia sua
ECCL|7|17|noli esse iustus multum neque plus sapias quam necesse est ne obstupescas
ECCL|7|18|ne impie agas multum et noli esse stultus ne moriaris in tempore non tuo
ECCL|7|19|bonum est te sustentare iustum sed et ab illo ne subtrahas manum tuam quia qui Deum timet nihil neglegit
ECCL|7|20|sapientia confortabit sapientem super decem principes civitatis
ECCL|7|21|non est enim homo iustus in terra qui faciat bonum et non peccet
ECCL|7|22|sed et cunctis sermonibus qui dicuntur ne accommodes cor tuum ne forte audias servum tuum maledicentem tibi
ECCL|7|23|scit enim tua conscientia quia et tu crebro maledixisti aliis
ECCL|7|24|cuncta temptavi in sapientia dixi sapiens efficiar et ipsa longius recessit a me
ECCL|7|25|multo magis quam erat et alta profunditas quis inveniet eam
ECCL|7|26|lustravi universa animo meo ut scirem et considerarem et quaererem sapientiam et rationem et ut cognoscerem impietatem stulti et errorem inprudentium
ECCL|7|27|et inveni amariorem morte mulierem quae laqueus venatorum est et sagena cor eius vincula sunt manus illius qui placet Deo effugiet eam qui autem peccator est capietur ab illa
ECCL|7|28|ecce hoc inveni dicit Ecclesiastes unum et alterum ut invenirem rationem
ECCL|7|29|quam adhuc quaerit anima mea et non inveni virum de mille unum repperi mulierem ex omnibus non inveni
ECCL|7|30|solummodo hoc inveni quod fecerit Deus hominem rectum et ipse se infinitis miscuerit quaestionibus quis talis ut sapiens est et quis cognovit solutionem verbi
ECCL|8|1|sapientia hominis lucet in vultu eius et potentissimus faciem illius commutavit
ECCL|8|2|ego os regis observo et praecepta iuramenti Dei
ECCL|8|3|ne festines recedere a facie eius neque permaneas in opere malo quia omne quod voluerit faciet
ECCL|8|4|et sermo illius potestate plenus est nec dicere ei quisquam potest quare ita facis
ECCL|8|5|qui custodit praeceptum non experietur quicquam mali tempus et responsionem cor sapientis intellegit
ECCL|8|6|omni negotio tempus est et oportunitas et multa hominis adflictio
ECCL|8|7|quia ignorat praeterita et ventura nullo scire potest nuntio
ECCL|8|8|non est in hominis dicione prohibere spiritum nec habet potestatem in die mortis nec sinitur quiescere ingruente bello neque salvabit impietas impium
ECCL|8|9|omnia haec consideravi et dedi cor meum in cunctis operibus quae fiunt sub sole interdum dominatur homo homini in malum suum
ECCL|8|10|vidi impios sepultos qui etiam cum adviverent in loco sancto erant et laudabantur in civitate quasi iustorum operum sed et hoc vanitas est
ECCL|8|11|etenim quia non profertur cito contra malos sententia absque ullo timore filii hominum perpetrant mala
ECCL|8|12|attamen ex eo quod peccator centies facit malum et per patientiam sustentatur ego cognovi quod erit bonum timentibus Deum qui verentur faciem eius
ECCL|8|13|non sit bonum impio nec prolongentur dies eius sed quasi umbra transeant qui non timent faciem Dei
ECCL|8|14|est et alia vanitas quae fit super terram sunt iusti quibus multa proveniunt quasi opera egerint impiorum et sunt impii qui ita securi sunt quasi iustorum facta habeant sed et hoc vanissimum iudico
ECCL|8|15|laudavi igitur laetitiam quod non esset homini bonum sub sole nisi quod comederet et biberet atque gauderet et hoc solum secum auferret de labore suo in diebus vitae quos dedit ei Deus sub sole
ECCL|8|16|et adposui cor meum ut scirem sapientiam et intellegerem distentionem quae versatur in terra est homo qui diebus ac noctibus somnum oculis non capit
ECCL|8|17|et intellexi quod omnium operum Dei nullam possit homo invenire rationem eorum quae fiunt sub sole et quanto plus laboraverit ad quaerendum tanto minus inveniat etiam si dixerit sapiens se nosse non poterit repperire
ECCL|9|1|omnia haec tractavi in corde meo ut curiose intellegerem sunt iusti atque sapientes et opera eorum in manu Dei et tamen nescit homo utrum amore an odio dignus sit
ECCL|9|2|sed omnia in futuro servantur incerta eo quod universa aeque eveniant iusto et impio bono et malo mundo et inmundo immolanti victimas et sacrificia contemnenti sicut bonus sic et peccator ut periurus ita et ille qui verum deierat
ECCL|9|3|hoc est pessimum inter omnia quae sub sole fiunt quia eadem cunctis eveniunt unde et corda filiorum hominum implentur malitia et contemptu in vita sua et post haec ad inferos deducentur
ECCL|9|4|nemo est qui semper vivat et qui huius rei habeat fiduciam melior est canis vivens leone mortuo
ECCL|9|5|viventes enim sciunt se esse morituros mortui vero nihil noverunt amplius nec habent ultra mercedem quia oblivioni tradita est memoria eorum
ECCL|9|6|amor quoque et odium et invidia simul perierunt nec habent partem in hoc saeculo et in opere quod sub sole geritur
ECCL|9|7|vade ergo et comede in laetitia panem tuum et bibe cum gaudio vinum tuum quia Deo placent opera tua
ECCL|9|8|omni tempore sint vestimenta tua candida et oleum de capite tuo non deficiat
ECCL|9|9|perfruere vita cum uxore quam diligis cunctis diebus vitae instabilitatis tuae qui dati sunt tibi sub sole omni tempore vanitatis tuae haec est enim pars in vita et in labore tuo quod laboras sub sole
ECCL|9|10|quodcumque potest manus tua facere instanter operare quia nec opus nec ratio nec scientia nec sapientia erunt apud inferos quo tu properas
ECCL|9|11|verti me alio vidique sub sole nec velocium esse cursum nec fortium bellum nec sapientium panem nec doctorum divitias nec artificum gratiam sed tempus casumque in omnibus
ECCL|9|12|nescit homo finem suum sed sicut pisces capiuntur hamo et sicut aves conprehenduntur laqueo sic capiuntur homines tempore malo cum eis extemplo supervenerit
ECCL|9|13|hanc quoque vidi sub sole sapientiam et probavi maximam
ECCL|9|14|civitas parva et pauci in ea viri venit contra eam rex magnus et vallavit eam extruxitque munitiones per gyrum et perfecta est obsidio
ECCL|9|15|inventusque in ea vir pauper et sapiens liberavit urbem per sapientiam suam et nullus deinceps recordatus est hominis illius pauperis
ECCL|9|16|et dicebam ego meliorem esse sapientiam fortitudine quomodo ergo sapientia pauperis contempta est et verba eius non sunt audita
ECCL|9|17|verba sapientium audiuntur in silentio plus quam clamor principis inter stultos
ECCL|9|18|melior est sapientia quam arma bellica et qui in uno peccaverit multa bona perdet
ECCL|10|1|muscae morientes perdunt suavitatem unguenti pretiosior est sapientia et gloria parva ad tempus stultitia
ECCL|10|2|cor sapientis in dextera eius et cor stulti in sinistra illius
ECCL|10|3|sed et in via stultus ambulans cum ipse insipiens sit omnes stultos aestimat
ECCL|10|4|si spiritus potestatem habentis ascenderit super te locum tuum ne dimiseris quia curatio cessare faciet peccata maxima
ECCL|10|5|est malum quod vidi sub sole quasi per errorem egrediens a facie principis
ECCL|10|6|positum stultum in dignitate sublimi et divites sedere deorsum
ECCL|10|7|vidi servos in equis et principes ambulantes quasi servos super terram
ECCL|10|8|qui fodit foveam incidet in eam et qui dissipat sepem mordebit eum coluber
ECCL|10|9|qui transfert lapides adfligetur in eis et qui scindit ligna vulnerabitur ab eis
ECCL|10|10|si retunsum fuerit ferrum et hoc non ut prius sed hebetatum erit multo labore exacuatur et post industriam sequitur sapientia
ECCL|10|11|si mordeat serpens in silentio nihil eo minus habet qui occulte detrahit
ECCL|10|12|verba oris sapientis gratia et labia insipientis praecipitabunt eum
ECCL|10|13|initium verborum eius stultitia et novissimum oris illius error pessimus
ECCL|10|14|stultus verba multiplicat ignorat homo quid ante se fuerit et quod post futurum est quis illi poterit indicare
ECCL|10|15|labor stultorum adfliget eos qui nesciunt in urbem pergere
ECCL|10|16|vae tibi terra cuius rex est puer et cuius principes mane comedunt
ECCL|10|17|beata terra cuius rex nobilis est et cuius principes vescuntur in tempore suo ad reficiendum et non ad luxuriam
ECCL|10|18|in pigritiis humiliabitur contignatio et in infirmitate manuum perstillabit domus
ECCL|10|19|in risu faciunt panem ac vinum ut epulentur viventes et pecuniae oboedient omnia
ECCL|10|20|in cogitatione tua regi ne detrahas et in secreto cubiculi tui ne maledixeris diviti quia avis caeli portabit vocem tuam et qui habet pinnas adnuntiabit sententiam
ECCL|11|1|mitte panem tuum super transeuntes aquas quia post multa tempora invenies illum
ECCL|11|2|da partem septem necnon et octo quia ignoras quid futurum sit mali super terram
ECCL|11|3|si repletae fuerint nubes imbrem super terram effundent si ceciderit lignum ad austrum aut ad aquilonem in quocumque loco ceciderit ibi erit
ECCL|11|4|qui observat ventum non seminat et qui considerat nubes numquam metet
ECCL|11|5|quomodo ignoras quae sit via spiritus et qua ratione conpingantur ossa in ventre praegnatis sic nescis opera Dei qui fabricator est omnium
ECCL|11|6|mane semina sementem tuam et vespere ne cesset manus tua quia nescis quid magis oriatur hoc an illud et si utrumque simul melius erit
ECCL|11|7|dulce lumen et delectabile est oculis videre solem
ECCL|11|8|si annis multis vixerit homo et in omnibus his laetatus fuerit meminisse debet tenebrosi temporis et dierum multorum qui cum venerint vanitatis arguentur praeterita
ECCL|11|9|laetare ergo iuvenis in adulescentia tua et in bono sit cor tuum in diebus iuventutis tuae et ambula in viis cordis tui et in intuitu oculorum tuorum et scito quod pro omnibus his adducet te Deus in iudicium
ECCL|11|10|aufer iram a corde tuo et amove malitiam a carne tua adulescentia enim et voluptas vana sunt
ECCL|12|1|memento creatoris tui in diebus iuventutis tuae antequam veniat tempus adflictionis et adpropinquent anni de quibus dicas non mihi placent
ECCL|12|2|antequam tenebrescat sol et lumen et luna et stellae et revertantur nubes post pluviam
ECCL|12|3|quando commovebuntur custodes domus et nutabuntur viri fortissimi et otiosae erunt molentes inminuto numero et tenebrescent videntes per foramina
ECCL|12|4|et claudent ostia in platea in humilitate vocis molentis et consurgent ad vocem volucris et obsurdescent omnes filiae carminis
ECCL|12|5|excelsa quoque timebunt et formidabunt in via florebit amigdalum inpinguabitur lucusta et dissipabitur capparis quoniam ibit homo in domum aeternitatis suae et circumibunt in platea plangentes
ECCL|12|6|antequam rumpatur funis argenteus et recurrat vitta aurea et conteratur hydria super fontem et confringatur rota super cisternam
ECCL|12|7|et revertatur pulvis in terram suam unde erat et spiritus redeat ad Deum qui dedit illum
ECCL|12|8|vanitas vanitatum dixit Ecclesiastes omnia vanitas
ECCL|12|9|cumque esset sapientissimus Ecclesiastes docuit populum et enarravit quae fecerit et investigans conposuit parabolas multas
ECCL|12|10|quaesivit verba utilia et conscripsit sermones rectissimos ac veritate plenos
ECCL|12|11|verba sapientium sicut stimuli et quasi clavi in altum defixi quae per magistrorum concilium data sunt a pastore uno
ECCL|12|12|his amplius fili mi ne requiras faciendi plures libros nullus est finis frequensque meditatio carnis adflictio est
ECCL|12|13|finem loquendi omnes pariter audiamus Deum time et mandata eius observa hoc est enim omnis homo
ECCL|12|14|et cuncta quae fiunt adducet Deus in iudicium pro omni errato sive bonum sive malum sit
