OBAD|1|1|俄巴底亞 所見的異象。 我們從耶和華那裏得到消息， 有使者被差往列國去： 「起來吧， 我們要起來與 以東 爭戰！」 主耶和華論 以東 如此說：
OBAD|1|2|看哪，我要使你在列國中為最小， 被人大大藐視。
OBAD|1|3|你狂傲的心欺騙了你， 你住在巖穴， 居所在高處， 心裏說： 「誰能把我拉下來到地上呢？」
OBAD|1|4|你雖如鷹高飛， 在星宿之間搭窩， 我必從那裏拉你下來。 這是耶和華說的。
OBAD|1|5|盜賊若來到你那裏， 小偷夜間來到， 豈不是只偷他們所需要的嗎？ 摘葡萄的若來到你那裏， 豈不留下幾串嗎？ 你竟全然滅絕！
OBAD|1|6|以掃 遭到搜查， 他隱藏的寶物竟被尋出！
OBAD|1|7|與你結盟的都驅趕你，直到邊界， 與你和好的欺騙你，勝過你， 吃你飯的人設下圈套陷害你─ 他卻毫無聰明 。
OBAD|1|8|到那日， 我豈不從 以東 除滅智慧人？ 從 以掃山 除滅聰明人？ 這是耶和華說的。
OBAD|1|9|提幔 哪， 你的勇士必驚惶， 以致 以掃山 的人都被殺戮剪除。
OBAD|1|10|因你向兄弟 雅各 施暴， 你必蒙羞， 永被剪除。
OBAD|1|11|當陌生人擄掠 雅各 的財物， 當外邦人進入他的城門， 為 耶路撒冷 抽籤分取財物的日子， 你竟站在一旁，像與他們同夥。
OBAD|1|12|你兄弟遭難的日子， 你不該瞪著眼看； 猶大 人被滅的日子， 你不該幸災樂禍； 他們遭難的日子， 你不該說狂傲的話。
OBAD|1|13|我子民遭災的日子， 你不該進他們的城門； 他們遭災的日子， 你不該瞪著眼看他們受苦； 他們遭災的日子， 你不該伸手搶他們的財物。
OBAD|1|14|他們遭難的日子， 你不該站在岔路口 剪除他們逃脫的人， 你不該交出他們的倖存者。
OBAD|1|15|耶和華的日子臨近萬國； 你所做的，人也必向你照樣做， 你的報應必歸到自己頭上。
OBAD|1|16|你們在我聖山怎樣喝了苦杯， 萬國必照樣不停地喝， 且喝且吞， 他們就必歸於無有。
OBAD|1|17|但在 錫安山 必有逃脫的人， 那山必成為聖； 雅各 家必得原有的產業 。
OBAD|1|18|雅各 家必成為大火， 約瑟 家成為火焰； 以掃 家必如碎秸， 遭燃燒，被吞滅， 以掃 家必無倖存者。 這是耶和華說的。
OBAD|1|19|他們必得 尼革夫 和 以掃山 ， 得 謝非拉 ， 非利士 人之地， 他們必得 以法蓮 地和 撒瑪利亞 地， 得 便雅憫 和 基列 ；
OBAD|1|20|被擄的 以色列 大軍 必得 迦南 人的地，直到 撒勒法 ， 在 西法拉 被擄的 耶路撒冷 人 必得 尼革夫 的城鎮。
OBAD|1|21|必有一些解救者 上到 錫安山 ，審判 以掃山 ， 國度就歸耶和華了。
