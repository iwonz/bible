DEUT|1|1|Сии суть слова, которые говорил Моисей всем Израильтянам за Иорданом в пустыне на равнине против Суфа, между Фараном и Тофелом, и Лаваном, и Асирофом, и Дизагавом,
DEUT|1|2|в расстоянии одиннадцати дней пути от Хорива, по дороге от горы Сеир к Кадес–Варни.
DEUT|1|3|Сорокового года, одиннадцатого месяца, в первый [день] месяца говорил Моисей сынам Израилевым все, что заповедал ему Господь о них.
DEUT|1|4|По убиении им Сигона, царя Аморрейского, который жил в Есевоне, и Ога, царя Васанского, который жил в Аштерофе в Едреи,
DEUT|1|5|за Иорданом, в земле Моавитской, начал Моисей изъяснять закон сей и сказал:
DEUT|1|6|Господь, Бог наш, говорил нам в Хориве и сказал: "полно вам жить на горе сей!
DEUT|1|7|обратитесь, отправьтесь в путь и пойдите на гору Аморреев и ко всем соседям их, на равнину, на гору, на низкие места и на южный край и к берегам моря, в землю Ханаанскую и к Ливану, даже до реки великой, реки Евфрата;
DEUT|1|8|вот, Я даю вам землю сию, пойдите, возьмите в наследие землю, которую Господь с клятвою обещал дать отцам вашим, Аврааму, Исааку и Иакову, им и потомству их".
DEUT|1|9|И я сказал вам в то время: не могу один водить вас;
DEUT|1|10|Господь, Бог ваш, размножил вас, и вот, вы ныне многочисленны, как звезды небесные;
DEUT|1|11|Господь, Бог отцов ваших, да умножит вас в тысячу крат против того, сколько вас [теперь], и да благословит вас, как Он говорил вам:
DEUT|1|12|как же мне одному носить тягости ваши, бремена ваши и распри ваши?
DEUT|1|13|изберите себе по коленам вашим мужей мудрых, разумных и испытанных, и я поставлю их начальниками вашими.
DEUT|1|14|Вы отвечали мне и сказали: хорошее дело велишь ты сделать.
DEUT|1|15|И взял я главных из колен ваших, мужей мудрых, и испытанных, и сделал их начальниками над вами, тысяченачальниками, стоначальниками, пятидесятиначальниками, десятиначальниками и надзирателями по коленам вашим.
DEUT|1|16|И дал я повеление судьям вашим в то время, говоря: выслушивайте братьев ваших и судите справедливо, как брата с братом, так и пришельца его;
DEUT|1|17|не различайте лиц на суде, как малого, так и великого выслушивайте: не бойтесь лица человеческого, ибо суд – дело Божие; а дело, которое для вас трудно, доводите до меня, и я выслушаю его.
DEUT|1|18|И дал я вам в то время повеления обо всем, что надлежит вам делать.
DEUT|1|19|И отправились мы от Хорива, и шли по всей этой великой и страшной пустыне, которую вы видели, по пути к горе Аморрейской, как повелел Господь, Бог наш, и пришли в Кадес–Варни.
DEUT|1|20|И сказал я вам: вы пришли к горе Аморрейской, которую Господь, Бог наш, дает нам;
DEUT|1|21|вот, Господь, Бог твой, отдает тебе землю сию, иди, возьми ее во владение, как говорил тебе Господь, Бог отцов твоих, не бойся и не ужасайся.
DEUT|1|22|Но вы все подошли ко мне и сказали: пошлем пред собою людей, чтоб они исследовали нам землю и принесли нам известие о дороге, по которой идти нам, и о городах, в которые идти нам.
DEUT|1|23|Слово это мне понравилось, и я взял из вас двенадцать человек, по одному человеку от [каждого] колена.
DEUT|1|24|Они пошли, взошли на гору и дошли до долины Есхол, и обозрели ее;
DEUT|1|25|и взяли в руки свои плодов земли и доставили нам, и принесли нам известие и сказали: хороша земля, которую Господь, Бог наш, дает нам.
DEUT|1|26|Но вы не захотели идти и воспротивились повелению Господа, Бога вашего,
DEUT|1|27|и роптали в шатрах ваших и говорили: Господь, по ненависти к нам, вывел нас из земли Египетской, чтоб отдать нас в руки Аморреев [и] истребить нас;
DEUT|1|28|куда мы пойдем? братья наши расслабили сердце наше, говоря: народ тот более, и выше нас, города [там] большие и с укреплениями до небес, да и сынов Енаковых видели мы там.
DEUT|1|29|И я сказал вам: не страшитесь и не бойтесь их;
DEUT|1|30|Господь, Бог ваш, идет перед вами; Он будет сражаться за вас, как Он сделал с вами в Египте, пред глазами вашими,
DEUT|1|31|и в пустыне сей, где, как ты видел, Господь, Бог твой, носил тебя, как человек носит сына своего, на всем пути, которым вы проходили до пришествия вашего на сие место.
DEUT|1|32|Но и при этом вы не верили Господу, Богу вашему,
DEUT|1|33|Который шел перед вами путем – искать вам места, где остановиться вам, ночью в огне, чтобы указывать вам дорогу, по которой идти, а днем в облаке.
DEUT|1|34|И Господь услышал слова ваши, и разгневался, и поклялся, говоря:
DEUT|1|35|никто из людей сих, из сего злого рода, не увидит доброй земли, которую Я клялся дать отцам вашим;
DEUT|1|36|только Халев, сын Иефонниин, увидит ее; ему дам Я землю, по которой он проходил, и сынам его, за то, что он повиновался Господу.
DEUT|1|37|И на меня прогневался Господь за вас, говоря: и ты не войдешь туда;
DEUT|1|38|Иисус, сын Навин, который при тебе, он войдет туда; его утверди, ибо он введет Израиля во владение ею;
DEUT|1|39|дети ваши, о которых вы говорили, что они достанутся в добычу [врагам], и сыновья ваши, которые не знают ныне ни добра ни зла, они войдут туда, им дам ее, и они овладеют ею;
DEUT|1|40|а вы обратитесь и отправьтесь в пустыню по дороге к Чермному морю.
DEUT|1|41|И вы отвечали тогда и сказали мне: согрешили мы пред Господом, пойдем и сразимся, как повелел нам Господь, Бог наш. И препоясались вы, каждый ратным оружием своим, и безрассудно решились взойти на гору.
DEUT|1|42|Но Господь сказал мне: скажи им: не всходите и не сражайтесь, потому что нет Меня среди вас, чтобы не поразили вас враги ваши.
DEUT|1|43|И я говорил вам, но вы не послушали и воспротивились повелению Господню и по упорству своему взошли на гору.
DEUT|1|44|И выступил против вас Аморрей, живший на горе той, и преследовали вас так, как делают пчелы, и поражали вас на Сеире до самой Хормы.
DEUT|1|45|И возвратились вы и плакали пред Господом: но Господь не услышал вопля вашего и не внял вам.
DEUT|1|46|И пробыли вы в Кадесе много времени, сколько времени вы [там] были.
DEUT|2|1|И обратились мы и отправились в пустыню к Чермному морю, как говорил мне Господь, и много времени ходили вокруг горы Сеира.
DEUT|2|2|И сказал мне Господь, говоря:
DEUT|2|3|полно вам ходить вокруг этой горы, обратитесь к северу;
DEUT|2|4|и народу дай повеление и скажи: вы будете проходить пределы братьев ваших, сынов Исавовых, живущих на Сеире, и они убоятся вас; но остерегайтесь
DEUT|2|5|начинать с ними войну, ибо Я не дам вам земли их ни на стопу ноги, потому что гору Сеир Я дал во владение Исаву;
DEUT|2|6|пищу покупайте у них за серебро и ешьте; и воду покупайте у них за серебро и пейте;
DEUT|2|7|ибо Господь, Бог твой, благословил тебя во всяком деле рук твоих, покровительствовал [тебе] во время путешествия твоего по великой пустыне сей; вот, сорок лет Господь, Бог твой, с тобою; ты ни в чем не терпел недостатка.
DEUT|2|8|И шли мы мимо братьев наших, сынов Исавовых, живущих на Сеире, путем равнины, от Елафа и Ецион–Гавера, и поворотили, и шли к пустыне Моава.
DEUT|2|9|И сказал мне Господь: не вступай во вражду с Моавом и не начинай с ними войны; ибо Я не дам тебе ничего от земли его во владение, потому что Ар отдал Я во владение сынам Лотовым;
DEUT|2|10|прежде жили там Эмимы, народ великий, многочисленный и высокий, как [сыны] Енаковы,
DEUT|2|11|и они считались между Рефаимами, как [сыны] Енаковы; Моавитяне же называют их Эмимами;
DEUT|2|12|а на Сеире жили прежде Хорреи; но сыны Исавовы прогнали их и истребили их от лица своего и поселились вместо их – так, как поступил Израиль с землею наследия своего, которую дал им Господь;
DEUT|2|13|итак встаньте и пройдите долину Заред. И прошли мы долину Заред.
DEUT|2|14|С тех пор, как мы пошли в Кадес–Варни и как прошли долину Заред, [минуло] тридцать восемь лет, и у нас перевелся из среды стана весь род ходящих на войну, как клялся им Господь;
DEUT|2|15|да и рука Господня была на них, чтоб истреблять их из среды стана, пока не вымерли.
DEUT|2|16|Когда же перевелись все ходящие на войну и вымерли из среды народа,
DEUT|2|17|тогда сказал мне Господь, говоря:
DEUT|2|18|ты проходишь ныне мимо пределов Моава, мимо Ара,
DEUT|2|19|и приблизился к Аммонитянам; не вступай с ними во вражду, и не начинай с ними войны, ибо Я не дам тебе ничего от земли сынов Аммоновых во владение, потому что Я отдал ее во владение сынам Лотовым;
DEUT|2|20|и она считалась землею Рефаимов; прежде жили на ней Рефаимы; Аммонитяне же называют их Замзумимами;
DEUT|2|21|народ великий, многочисленный и высокий, как [сыны] Енаковы, и истребил их Господь пред лицем их, и изгнали они их и поселились на месте их,
DEUT|2|22|как Он сделал для сынов Исавовых, живущих на Сеире, истребив пред лицем их Хорреев, и они изгнали их, и поселились на месте их, и [живут] до сего дня;
DEUT|2|23|и Аввеев, живших в селениях до самой Газы, Кафторимы, исшедшие из Кафтора, истребили и поселились на месте их.
DEUT|2|24|Встаньте, отправьтесь и перейдите поток Арнон; вот, Я предаю в руку твою Сигона, царя Есевонского, Аморреянина, и землю его; начинай овладевать ею, и веди с ним войну;
DEUT|2|25|с сего дня Я начну распространять страх и ужас пред тобою на народы под всем небом; те, которые услышат о тебе, вострепещут и ужаснутся тебя.
DEUT|2|26|И послал я послов из пустыни Кедемоф к Сигону, царю Есевонскому, с словами мирными, чтобы сказать:
DEUT|2|27|позволь пройти мне землею твоею; я пойду дорогою, не сойду ни направо, ни налево;
DEUT|2|28|пищу продавай мне за серебро, и я буду есть, и воду для питья давай мне за серебро, и я буду пить, только ногами моими пройду –
DEUT|2|29|так, как сделали мне сыны Исава, живущие на Сеире, и Моавитяне, живущие в Аре, доколе не перейду чрез Иордан в землю, которую Господь, Бог наш, дает нам.
DEUT|2|30|Но Сигон, царь Есевонский, не согласился позволить пройти нам через свою [землю], потому что Господь, Бог твой, ожесточил дух его и сердце его сделал упорным, чтобы предать его в руку твою, как [это видно] ныне.
DEUT|2|31|И сказал мне Господь: вот, Я начинаю предавать тебе Сигона и землю его; начинай овладевать землею его.
DEUT|2|32|И Сигон со всем народом своим выступил против нас на сражение к Яаце;
DEUT|2|33|и предал его Господь, Бог наш, [в руки наши], и мы поразили его и сынов его и весь народ его,
DEUT|2|34|и взяли в то время все города его, и предали заклятию все города, мужчин и женщин и детей, не оставили никого в живых;
DEUT|2|35|только взяли мы себе в добычу скот их и захваченное во взятых нами городах.
DEUT|2|36|От Ароера, который на берегу потока Арнона, и от города, который на долине, до Галаада не было города, который был бы неприступен для нас: все предал Господь, Бог наш, [в руки наши].
DEUT|2|37|Только к земле Аммонитян ты не подходил, ни к [местам лежащим] близ потока Иавока, ни к городам на горе, ни ко всему, к чему не повелел [нам] Господь, Бог наш.
DEUT|3|1|И обратились мы оттуда, и шли к Васану, и выступил против нас на войну Ог, царь Васанский, со всем народом своим, при Едреи.
DEUT|3|2|И сказал мне Господь: не бойся его, ибо Я отдам в руку твою его, и весь народ его, и всю землю его, и ты поступишь с ним так, как поступил с Сигоном, царем Аморрейским, который жил в Есевоне.
DEUT|3|3|И предал Господь, Бог наш, в руки наши и Ога, царя Васанского, и весь народ его; и мы поразили его, так что никого не осталось у него в живых;
DEUT|3|4|и взяли мы в то время все города его; не было города, которого мы не взяли бы у них: шестьдесят городов, всю область Аргов, царство Ога Васанского;
DEUT|3|5|все эти города укреплены были высокими стенами, воротами и запорами, кроме городов неукрепленных, весьма многих;
DEUT|3|6|и предали мы их заклятию, как поступили с Сигоном, царем Есевонским, предав заклятию всякий город с мужчинами, женщинами и детьми;
DEUT|3|7|но весь скот и захваченное в городах взяли себе в добычу.
DEUT|3|8|И взяли мы в то время из руки двух царей Аморрейских землю сию, которая по эту сторону Иордана, от потока Арнона до горы Ермона, –
DEUT|3|9|Сидоняне Ермон называют Сирионом, а Аморреи называют его Сениром, –
DEUT|3|10|все города на равнине, весь Галаад и весь Васан до Салхи и Едреи, города царства Ога Васанского;
DEUT|3|11|ибо только Ог, царь Васанский, оставался из Рефаимов. Вот, одр его, одр железный, и теперь в Равве, у сынов Аммоновых: длина его девять локтей, а ширина его четыре локтя, локтей мужеских.
DEUT|3|12|Землю сию взяли мы в то время начиная от Ароера, который у потока Арнона; и половину горы Галаада с городами ее отдал я [колену] Рувимову и Гадову;
DEUT|3|13|а остаток Галаада и весь Васан, царство Ога, отдал я половине колена Манассиина, всю область Аргов со всем Васаном.
DEUT|3|14|Иаир, сын Манассиин, взял всю область Аргов, до пределов Гесурских и Маахских, и назвал Васан, по имени своему, селениями Иаировыми, что и доныне;
DEUT|3|15|Махиру дал я Галаад;
DEUT|3|16|а [колену] Рувимову и Гадову дал от Галаада до потока Арнона, [землю] между потоком и пределом, до потока Иавока, предела сынов Аммоновых,
DEUT|3|17|также равнину и Иордан, [который есть] и предел, от Киннерефа до моря равнины, моря Соленого, при подошве [горы] Фасги к востоку.
DEUT|3|18|И дал я вам в то время повеление, говоря: Господь, Бог ваш, дал вам землю сию во владение; все способные к войне, вооружившись, идите впереди братьев ваших, сынов Израилевых;
DEUT|3|19|только жены ваши и дети ваши и скот ваш пусть останутся в городах ваших, которые я дал вам,
DEUT|3|20|доколе Господь не даст покоя братьям вашим, как вам, и доколе и они не получат во владение землю, которую Господь, Бог ваш, дает им за Иорданом; тогда возвратитесь каждый в свое владение, которое я дал вам.
DEUT|3|21|И Иисусу заповедал я в то время, говоря: глаза твои видели все, что сделал Господь, Бог ваш, с двумя царями сими; то же сделает Господь со всеми царствами, которые ты будешь проходить;
DEUT|3|22|не бойтесь их, ибо Господь, Бог ваш, Сам сражается за вас.
DEUT|3|23|И молился я Господу в то время, говоря:
DEUT|3|24|Владыко Господи, Ты начал показывать рабу Твоему величие Твое и крепкую руку Твою; ибо какой бог есть на небе, или на земле, который мог бы делать такие дела, как Твои, и с могуществом таким, как Твое?
DEUT|3|25|дай мне перейти и увидеть ту добрую землю, которая за Иорданом, и ту прекрасную гору и Ливан.
DEUT|3|26|Но Господь гневался на меня за вас и не послушал меня, и сказал мне Господь: полно тебе, впредь не говори Мне более об этом;
DEUT|3|27|взойди на вершину Фасги и взгляни глазами твоими к морю и к северу, и к югу и к востоку, и посмотри глазами твоими, потому что ты не перейдешь за Иордан сей;
DEUT|3|28|и дай наставление Иисусу, и укрепи его, и утверди его; ибо он будет предшествовать народу сему и он разделит им на уделы землю, на которую ты посмотришь.
DEUT|3|29|И остановились мы на долине, напротив Беф–Фегора.
DEUT|4|1|Итак, Израиль, слушай постановления и законы, которые я научаю вас исполнять, дабы вы были живы, и пошли и наследовали ту землю, которую Господь, Бог отцов ваших, дает вам.
DEUT|4|2|не прибавляйте к тому, что я заповедую вам, и не убавляйте от того; соблюдайте заповеди Господа, Бога вашего, которые я вам заповедую.
DEUT|4|3|Глаза ваши видели [все], что сделал Господь с Ваал–Фегором: всякого человека, последовавшего Ваал–Фегору, истребил Господь, Бог твой, из среды тебя;
DEUT|4|4|а вы, прилепившиеся к Господу, Богу вашему, живы все доныне.
DEUT|4|5|Вот, я научил вас постановлениям и законам, как повелел мне Господь, Бог мой, дабы вы так поступали в той земле, в которую вы вступаете, чтоб овладеть ею;
DEUT|4|6|итак храните и исполняйте их, ибо в этом мудрость ваша и разум ваш пред глазами народов, которые, услышав о всех сих постановлениях, скажут: только этот великий народ есть народ мудрый и разумный.
DEUT|4|7|Ибо есть ли какой великий народ, к которому боги [его] были бы столь близки, как близок к нам Господь, Бог наш, когда ни призовем Его?
DEUT|4|8|и есть ли какой великий народ, у которого были бы такие справедливые постановления и законы, как весь закон сей, который я предлагаю вам сегодня?
DEUT|4|9|Только берегись и тщательно храни душу твою, чтобы тебе не забыть тех дел, которые видели глаза твои, и чтобы они не выходили из сердца твоего во все дни жизни твоей; и поведай о них сынам твоим и сынам сынов твоих, –
DEUT|4|10|о том дне, когда ты стоял пред Господом, Богом твоим, при Хориве, и когда сказал Господь мне: собери ко Мне народ, и Я возвещу им слова Мои, из которых они научатся бояться Меня во все дни жизни своей на земле и научат сыновей своих.
DEUT|4|11|Вы приблизились и стали под горою, а гора горела огнем до самых небес, [и была] тьма, облако и мрак.
DEUT|4|12|И говорил Господь к вам из среды огня; глас слов [Его] вы слышали, но образа не видели, а только глас;
DEUT|4|13|и объявил Он вам завет Свой, который повелел вам исполнять, десятословие, и написал его на двух каменных скрижалях;
DEUT|4|14|и повелел мне Господь в то время научить вас постановлениям и законам, дабы вы исполняли их в той земле, в которую вы входите, чтоб овладеть ею.
DEUT|4|15|Твердо держите в душах ваших, что вы не видели никакого образа в тот день, когда говорил к вам Господь на Хориве из среды огня,
DEUT|4|16|дабы вы не развратились и не сделали себе изваяний, изображений какого–либо кумира, представляющих мужчину или женщину,
DEUT|4|17|изображения какого–либо скота, который на земле, изображения какой–либо птицы крылатой, которая летает под небесами,
DEUT|4|18|изображения какого–либо [гада], ползающего по земле, изображения какой–либо рыбы, которая в водах ниже земли;
DEUT|4|19|и дабы ты, взглянув на небо и увидев солнце, луну и звезды [и] все воинство небесное, не прельстился и не поклонился им и не служил им, так как Господь, Бог твой, уделил их всем народам под всем небом.
DEUT|4|20|А вас взял Господь и вывел вас из печи железной, из Египта, дабы вы были народом Его удела, как это ныне [видно].
DEUT|4|21|И Господь прогневался на меня за вас, и клялся, что я не перейду за Иордан и не войду в ту добрую землю, которую Господь, Бог твой, дает тебе в удел;
DEUT|4|22|я умру в сей земле, не перейдя за Иордан, а вы перейдете и овладеете тою доброю землею.
DEUT|4|23|Берегитесь, чтобы не забыть вам завета Господа, Бога вашего, который Он поставил с вами, и чтобы не делать себе кумиров, изображающих что–либо, как повелел тебе Господь, Бог твой;
DEUT|4|24|ибо Господь, Бог твой, есть огнь поядающий, Бог ревнитель.
DEUT|4|25|Если же родятся у тебя сыны и сыны у сынов [твоих], и, долго жив на земле, вы развратитесь и сделаете изваяние, изображающее что–либо, и сделаете зло сие пред очами Господа, Бога вашего, и раздражите Его,
DEUT|4|26|то свидетельствуюсь вам сегодня небом и землею, что скоро потеряете землю, для наследования которой вы переходите за Иордан; не пробудете много времени на ней, но погибнете;
DEUT|4|27|и рассеет вас Господь по [всем] народам, и останетесь в малом числе между народами, к которым отведет вас Господь;
DEUT|4|28|и будете там служить богам, сделанным руками человеческими из дерева и камня, которые не видят и не слышат, и не едят и не обоняют.
DEUT|4|29|Но когда ты взыщешь там Господа, Бога твоего, то найдешь [Его], если будешь искать Его всем сердцем твоим и всею душею твоею.
DEUT|4|30|Когда ты будешь в скорби, и когда все это постигнет тебя в последствие времени, то обратишься к Господу, Богу твоему, и послушаешь гласа Его.
DEUT|4|31|Господь, Бог твой, есть Бог милосердый; Он не оставит тебя и не погубит тебя, и не забудет завета с отцами твоими, который Он клятвою утвердил им.
DEUT|4|32|Ибо спроси у времен прежних, бывших прежде тебя, с того дня, в который сотворил Бог человека на земле, и от края неба до края неба: бывало ли что–нибудь такое, как сие великое дело, или слыхано ли подобное сему?
DEUT|4|33|слышал ли [какой] народ глас Бога, говорящего из среды огня, и остался жив, как слышал ты?
DEUT|4|34|или покушался ли [какой] бог пойти, взять себе народ из среды [другого] народа казнями, знамениями и чудесами, и войною, и рукою крепкою, и мышцею высокою, и великими ужасами, как сделал для вас Господь, Бог ваш, в Египте пред глазами твоими?
DEUT|4|35|Тебе дано видеть [это], чтобы ты знал, что [только] Господь есть Бог, [и] нет еще кроме Его;
DEUT|4|36|с неба дал Он слышать тебе глас Свой, дабы научить тебя, и на земле показал тебе великий огнь Свой, и ты слышал слова Его из среды огня;
DEUT|4|37|и так как Он возлюбил отцов твоих и избрал [вас], потомство их после них, то и вывел тебя Сам великою силою Своею из Египта,
DEUT|4|38|чтобы прогнать от лица твоего народы, которые больше и сильнее тебя, [и] ввести тебя [и] дать тебе землю их в удел, как это ныне [видно].
DEUT|4|39|Итак знай ныне и положи на сердце твое, что Господь есть Бог на небе вверху и на земле внизу, [и] нет еще [кроме Его];
DEUT|4|40|и храни постановления Его и заповеди Его, которые я заповедую тебе ныне, чтобы хорошо было тебе и сынам твоим после тебя, и чтобы ты много времени пробыл на той земле, которую Господь, Бог твой, дает тебе навсегда.
DEUT|4|41|Тогда отделил Моисей три города по эту сторону Иордана на восток солнца,
DEUT|4|42|чтоб убегал туда убийца, который убьет ближнего своего без намерения, не быв врагом ему ни вчера, ни третьего дня, [и] чтоб, убежав в один из этих городов, остался жив:
DEUT|4|43|Бецер в пустыне, на равнине в [колене] Рувимовом, и Рамоф в Галааде в [колене] Гадовом, и Голан в Васане в [колене] Манассиином.
DEUT|4|44|Вот закон, который предложил Моисей сынам Израилевым;
DEUT|4|45|вот повеления, постановления и уставы, которые изрек Моисей сынам Израилевым, по исшествии их из Египта,
DEUT|4|46|за Иорданом, на долине против Беф–Фегора, в земле Сигона, царя Аморрейского, жившего в Есевоне, которого поразил Моисей с сынами Израилевыми, по исшествии их из Египта.
DEUT|4|47|И овладели они землею его и землею Ога, царя Васанского, двух царей Аморрейских, которая за Иорданом к востоку солнца,
DEUT|4|48|[начиная] от Ароера, который [лежит] на берегу потока Арнона, до горы Сиона, она же Ермон,
DEUT|4|49|и всею равниною по эту сторону Иордана к востоку, до самого моря равнины при подошве Фасги.
DEUT|5|1|И созвал Моисей весь Израиль и сказал им: слушай, Израиль, постановления и законы, которые я изреку сегодня в уши ваши, и выучите их и старайтесь исполнять их.
DEUT|5|2|Господь, Бог наш, поставил с нами завет на Хориве;
DEUT|5|3|не с отцами нашими поставил Господь завет сей, но с нами, [которые] здесь сегодня все живы.
DEUT|5|4|Лицем к лицу говорил Господь с вами на горе из среды огня;
DEUT|5|5|я же стоял между Господом и между вами в то время, дабы пересказывать вам слово Господа, ибо вы боялись огня и не восходили на гору. Он [тогда] сказал:
DEUT|5|6|Я Господь, Бог твой, Который вывел тебя из земли Египетской, из дома рабства;
DEUT|5|7|да не будет у тебя других богов перед лицем Моим.
DEUT|5|8|Не делай себе кумира и никакого изображения того, что на небе вверху и что на земле внизу, и что в водах ниже земли,
DEUT|5|9|не поклоняйся им и не служи им; ибо Я Господь, Бог твой, Бог ревнитель, за вину отцов наказывающий детей до третьего и четвертого рода, ненавидящих Меня,
DEUT|5|10|и творящий милость до тысячи [родов] любящим Меня и соблюдающим заповеди Мои.
DEUT|5|11|Не произноси имени Господа, Бога твоего, напрасно; ибо не оставит Господь без наказания того, кто употребляет имя Его напрасно.
DEUT|5|12|Наблюдай день субботний, чтобы свято хранить его, как заповедал тебе Господь, Бог твой;
DEUT|5|13|шесть дней работай и делай всякие дела твои,
DEUT|5|14|а день седьмой – суббота Господу, Богу твоему. Не делай [в оный] никакого дела, ни ты, ни сын твой, ни дочь твоя, ни раб твой, ни раба твоя, ни вол твой, ни осел твой, ни всякий скот твой, ни пришелец твой, который у тебя, чтобы отдохнул раб твой, и раба твоя, как и ты;
DEUT|5|15|и помни, что [ты] был рабом в земле Египетской, но Господь, Бог твой, вывел тебя оттуда рукою крепкою и мышцею высокою, потому и повелел тебе Господь, Бог твой, соблюдать день субботний.
DEUT|5|16|Почитай отца твоего и матерь твою, как повелел тебе Господь, Бог твой, чтобы продлились дни твои, и чтобы хорошо тебе было на той земле, которую Господь, Бог твой, дает тебе.
DEUT|5|17|Не убивай.
DEUT|5|18|Не прелюбодействуй.
DEUT|5|19|Не кради.
DEUT|5|20|Не произноси ложного свидетельства на ближнего твоего.
DEUT|5|21|Не желай жены ближнего твоего и не желай дома ближнего твоего, ни поля его, ни раба его, ни рабы его, ни вола его, ни осла его, ни всего, что есть у ближнего твоего.
DEUT|5|22|Слова сии изрек Господь ко всему собранию вашему на горе из среды огня, облака и мрака громогласно, и более не говорил, и написал их на двух каменных скрижалях, и дал их мне.
DEUT|5|23|И когда вы услышали глас из среды мрака, и гора горела огнем, то вы подошли ко мне, все начальники колен ваших и старейшины ваши,
DEUT|5|24|и сказали: вот, показал нам Господь, Бог наш, славу Свою и величие Свое, и глас Его слышали мы из среды огня; сегодня видели мы, что Бог говорит с человеком, и сей остается жив;
DEUT|5|25|но теперь для чего нам умирать? ибо великий огонь сей пожрет нас; если мы еще услышим глас Господа, Бога нашего, то умрем,
DEUT|5|26|ибо есть ли какая плоть, которая слышала бы глас Бога живаго, говорящего из среды огня, как мы, и осталась жива?
DEUT|5|27|приступи ты и слушай все, что скажет [тебе] Господь, Бог наш, и ты пересказывай нам все, что будет говорить тебе Господь, Бог наш, и мы будем слушать и исполнять.
DEUT|5|28|И Господь услышал слова ваши, как вы разговаривали со мною, и сказал мне Господь: слышал Я слова народа сего, которые они говорили тебе; все, что ни говорили они, хорошо;
DEUT|5|29|о, если бы сердце их было у них таково, чтобы бояться Меня и соблюдать все заповеди Мои во все дни, дабы хорошо было им и сынам их вовек!
DEUT|5|30|пойди, скажи им: "возвратитесь в шатры свои";
DEUT|5|31|а ты здесь останься со Мною, и Я изреку тебе все заповеди и постановления и законы, которым ты должен научить их, чтобы они [так] поступали на той земле, которую Я даю им во владение.
DEUT|5|32|Смотрите, поступайте так, как повелел вам Господь, Бог ваш; не уклоняйтесь ни направо, ни налево;
DEUT|5|33|ходите по тому пути, по которому повелел вам Господь, Бог ваш, дабы вы были живы, и хорошо было вам, и прожили много времени на той земле, которую получите во владение.
DEUT|6|1|Вот заповеди, постановления и законы, которым повелел Господь, Бог ваш, научить вас, чтобы вы поступали [так] в той земле, в которую вы идете, чтоб овладеть ею;
DEUT|6|2|дабы ты боялся Господа, Бога твоего, и все постановления Его и заповеди Его, которые заповедую тебе, соблюдал ты и сыны твои и сыны сынов твоих во все дни жизни твоей, дабы продлились дни твои.
DEUT|6|3|Итак слушай, Израиль, и старайся исполнить это, чтобы тебе хорошо было, и чтобы вы весьма размножились, как Господь, Бог отцов твоих, говорил тебе, [что Он даст тебе] землю, где течет молоко и мед.
DEUT|6|4|Слушай, Израиль: Господь, Бог наш, Господь един есть;
DEUT|6|5|и люби Господа, Бога твоего, всем сердцем твоим, и всею душею твоею и всеми силами твоими.
DEUT|6|6|И да будут слова сии, которые Я заповедую тебе сегодня, в сердце твоем.
DEUT|6|7|и внушай их детям твоим и говори о них, сидя в доме твоем и идя дорогою, и ложась и вставая;
DEUT|6|8|и навяжи их в знак на руку твою, и да будут они повязкою над глазами твоими,
DEUT|6|9|и напиши их на косяках дома твоего и на воротах твоих.
DEUT|6|10|Когда же введет тебя Господь, Бог твой, в ту землю, которую Он клялся отцам твоим, Аврааму, Исааку и Иакову, дать тебе с большими и хорошими городами, которых ты не строил,
DEUT|6|11|и с домами, наполненными всяким добром, которых ты не наполнял, и с колодезями, высеченными [из камня], которых ты не высекал, с виноградниками и маслинами, которых ты не садил, и будешь есть и насыщаться,
DEUT|6|12|тогда берегись, чтобы не забыл ты Господа, Который вывел тебя из земли Египетской, из дома рабства.
DEUT|6|13|Господа, Бога твоего, бойся, и Ему [одному] служи, и Его именем клянись.
DEUT|6|14|Не последуйте иным богам, богам тех народов, которые будут вокруг вас;
DEUT|6|15|ибо Господь, Бог твой, Который среди тебя, есть Бог ревнитель; чтобы не воспламенился гнев Господа, Бога твоего, на тебя, и не истребил Он тебя с лица земли.
DEUT|6|16|Не искушайте Господа, Бога вашего, как вы искушали Его в Массе.
DEUT|6|17|Твердо храните заповеди Господа, Бога вашего, и уставы Его и постановления, которые Он заповедал тебе;
DEUT|6|18|и делай справедливое и доброе пред очами Господа, дабы хорошо тебе было, и дабы ты вошел и овладел доброю землею, которую Господь с клятвою обещал отцам твоим,
DEUT|6|19|и чтобы Он прогнал всех врагов твоих от лица твоего, как говорил Господь.
DEUT|6|20|Если спросит у тебя сын твой в последующее время, говоря: "что [значат] сии уставы, постановления и законы, которые заповедал вам Господь, Бог ваш?"
DEUT|6|21|то скажи сыну твоему: "рабами были мы у фараона в Египте, но Господь вывел нас из Египта рукою крепкою;
DEUT|6|22|и явил Господь знамения и чудеса великие и казни над Египтом, над фараоном и над всем домом его пред глазами нашими;
DEUT|6|23|а нас вывел оттуда чтобы ввести нас и дать нам землю, которую клялся отцам нашим [дать нам];
DEUT|6|24|и заповедал нам Господь исполнять все постановления сии, чтобы мы боялись Господа, Бога нашего, дабы хорошо было нам во все дни, дабы сохранить нашу жизнь, как и теперь;
DEUT|6|25|и в сем будет наша праведность, если мы будем стараться исполнять все сии заповеди пред лицем Господа, Бога нашего, как Он заповедал нам".
DEUT|7|1|Когда введет тебя Господь, Бог твой, в землю, в которую ты идешь, чтоб овладеть ею, и изгонит от лица твоего многочисленные народы, Хеттеев, Гергесеев, Аморреев, Хананеев, Ферезеев, Евеев и Иевусеев, семь народов, которые многочисленнее и сильнее тебя,
DEUT|7|2|и предаст их тебе Господь, Бог твой, и поразишь их, тогда предай их заклятию, не вступай с ними в союз и не щади их;
DEUT|7|3|и не вступай с ними в родство: дочери твоей не отдавай за сына его, и дочери его не бери за сына твоего;
DEUT|7|4|ибо они отвратят сынов твоих от Меня, чтобы служить иным богам, и [тогда] воспламенится на вас гнев Господа, и Он скоро истребит тебя.
DEUT|7|5|Но поступите с ними так: жертвенники их разрушьте, столбы их сокрушите, и рощи их вырубите, и истуканов их сожгите огнем;
DEUT|7|6|ибо ты народ святый у Господа, Бога твоего: тебя избрал Господь, Бог твой, чтобы ты был собственным Его народом из всех народов, которые на земле.
DEUT|7|7|Не потому, чтобы вы были многочисленнее всех народов, принял вас Господь и избрал вас, – ибо вы малочисленнее всех народов, –
DEUT|7|8|но потому, что любит вас Господь, и для того, чтобы сохранить клятву, которою Он клялся отцам вашим, вывел вас Господь рукою крепкою и освободил тебя из дома рабства, из руки фараона, царя Египетского.
DEUT|7|9|Итак знай, что Господь, Бог твой, есть Бог, Бог верный, Который хранит завет [Свой] и милость к любящим Его и сохраняющим заповеди Его до тысячи родов,
DEUT|7|10|и воздает ненавидящим Его в лице их, погубляя их; Он не замедлит, ненавидящему Его самому лично воздаст.
DEUT|7|11|Итак, соблюдай заповеди и постановления и законы, которые сегодня заповедую тебе исполнять.
DEUT|7|12|И если вы будете слушать законы сии и хранить и исполнять их, то Господь, Бог твой, будет хранить завет и милость к тебе, как Он клялся отцам твоим,
DEUT|7|13|и возлюбит тебя, и благословит тебя, и размножит тебя, и благословит плод чрева твоего и плод земли твоей, и хлеб твой, и вино твое, и елей твой, рождаемое от крупного скота твоего и от стада овец твоих, на той земле, которую Он клялся отцам твоим дать тебе;
DEUT|7|14|благословен ты будешь больше всех народов; не будет ни бесплодного, ни бесплодной, ни у тебя, ни в скоте твоем;
DEUT|7|15|и отдалит от тебя Господь всякую немощь, и никаких лютых болезней Египетских, которые ты знаешь, не наведет на тебя, но наведет их на всех, ненавидящих тебя;
DEUT|7|16|и истребишь все народы, которые Господь, Бог твой, дает тебе: да не пощадит их глаз твой; и не служи богам их, ибо это сеть для тебя.
DEUT|7|17|Если скажешь в сердце твоем: "народы сии многочисленнее меня; как я могу изгнать их?"
DEUT|7|18|Не бойся их, вспомни то, что сделал Господь, Бог твой, с фараоном и всем Египтом,
DEUT|7|19|те великие испытания, которые видели глаза твои, знамения, чудеса, и руку крепкую и мышцу высокую, с какими вывел тебя Господь, Бог твой; то же сделает Господь, Бог твой, со всеми народами, которых ты боишься;
DEUT|7|20|и шершней нашлет Господь, Бог твой, на них, доколе не погибнут оставшиеся и скрывшиеся от лица твоего;
DEUT|7|21|не страшись их, ибо Господь, Бог твой, среди тебя, Бог великий и страшный.
DEUT|7|22|И будет Господь, Бог твой, изгонять пред тобою народы сии мало–помалу; не можешь ты истребить их скоро, чтобы не умножились против тебя полевые звери;
DEUT|7|23|но предаст их тебе Господь, Бог твой, и приведет их в великое смятение, так что они погибнут;
DEUT|7|24|и предаст царей их в руки твои, и ты истребишь имя их из поднебесной: не устоит никто против тебя, доколе не искоренишь их.
DEUT|7|25|Кумиры богов их сожгите огнем; не пожелай взять себе серебра или золота, которое на них, дабы это не было для тебя сетью, ибо это мерзость для Господа, Бога твоего;
DEUT|7|26|и не вноси мерзости в дом твой, дабы не подпасть заклятию, как она; отвращайся сего и гнушайся сего, ибо это заклятое.
DEUT|8|1|Все заповеди, которые я заповедую вам сегодня, старайтесь исполнять, дабы вы были живы и размножились, и пошли и завладели землею, которую с клятвою обещал Господь отцам вашим.
DEUT|8|2|И помни весь путь, которым вел тебя Господь, Бог твой, по пустыне, вот уже сорок лет, чтобы смирить тебя, чтобы испытать тебя и узнать, что в сердце твоем, будешь ли хранить заповеди Его, или нет;
DEUT|8|3|Он смирял тебя, томил тебя голодом и питал тебя манною, которой не знал ты и не знали отцы твои, дабы показать тебе, что не одним хлебом живет человек, но всяким [словом], исходящим из уст Господа, живет человек;
DEUT|8|4|одежда твоя не ветшала на тебе, и нога твоя не пухла, вот уже сорок лет.
DEUT|8|5|И знай в сердце твоем, что Господь, Бог твой, учит тебя, как человек учит сына своего.
DEUT|8|6|Итак храни заповеди Господа, Бога твоего, ходя путями Его и боясь Его.
DEUT|8|7|Ибо Господь, Бог твой, ведет тебя в землю добрую, в землю, [где] потоки вод, источники и озера выходят из долин и гор,
DEUT|8|8|в землю, [где] пшеница, ячмень, виноградные лозы, смоковницы и гранатовые деревья, в землю, [где] масличные деревья и мед,
DEUT|8|9|в землю, в которой без скудости будешь есть хлеб твой и ни в чем не будешь иметь недостатка, в землю, в которой камни – железо, и из гор которой будешь высекать медь.
DEUT|8|10|И когда будешь есть и насыщаться, тогда благословляй Господа, Бога твоего, за добрую землю, которую Он дал тебе.
DEUT|8|11|Берегись, чтобы ты не забыл Господа, Бога твоего, не соблюдая заповедей Его, и законов Его, и постановлений Его, которые сегодня заповедую тебе.
DEUT|8|12|Когда будешь есть и насыщаться, и построишь хорошие домы и будешь жить [в них],
DEUT|8|13|и когда будет у тебя много крупного и мелкого скота, и будет много серебра и золота, и всего у тебя будет много, –
DEUT|8|14|то смотри, чтобы не надмилось сердце твое и не забыл ты Господа, Бога твоего, Который вывел тебя из земли Египетской, из дома рабства;
DEUT|8|15|Который провел тебя по пустыне великой и страшной, [где] змеи, василиски, скорпионы и места сухие, на которых нет воды; Который источил для тебя [источник] воды из скалы гранитной,
DEUT|8|16|питал тебя в пустыне манною, которой не знали отцы твои, дабы смирить тебя и испытать тебя, чтобы впоследствии сделать тебе добро,
DEUT|8|17|и чтобы ты не сказал в сердце твоем: "моя сила и крепость руки моей приобрели мне богатство сие",
DEUT|8|18|но чтобы помнил Господа, Бога твоего, ибо Он дает тебе силу приобретать богатство, дабы исполнить, как ныне, завет Свой, который Он клятвою утвердил отцам твоим.
DEUT|8|19|Если же ты забудешь Господа, Бога твоего, и пойдешь вслед богов других, и будешь служить им и поклоняться им, то свидетельствуюсь вам сегодня, что вы погибнете;
DEUT|8|20|как народы, которые Господь истребляет от лица вашего, так погибнете [и вы] за то, что не послушаете гласа Господа, Бога вашего.
DEUT|9|1|Слушай, Израиль: ты теперь идешь за Иордан, чтобы пойти овладеть народами, которые больше и сильнее тебя, городами большими, с укреплениями до небес,
DEUT|9|2|народом многочисленным и великорослым, сынами Енаковыми, о которых ты знаешь и слышал: "кто устоит против сынов Енаковых?"
DEUT|9|3|Знай же ныне, что Господь, Бог твой, идет пред тобою, [как] огнь поядающий; Он будет истреблять их и низлагать их пред тобою, и ты изгонишь их, и погубишь их скоро, как говорил тебе Господь.
DEUT|9|4|Когда будет изгонять их Господь, Бог твой, от лица твоего, не говори в сердце твоем, что за праведность мою привел меня Господь овладеть сею землею, и что за нечестие народов сих Господь изгоняет их от лица твоего;
DEUT|9|5|не за праведность твою и не за правоту сердца твоего идешь ты наследовать землю их, но за нечестие народов сих Господь, Бог твой, изгоняет их от лица твоего, и дабы исполнить слово, которым клялся Господь отцам твоим Аврааму, Исааку и Иакову;
DEUT|9|6|посему знай, что не за праведность твою Господь, Бог твой, дает тебе овладеть сею доброю землею, ибо ты народ жестоковыйный.
DEUT|9|7|Помни, не забудь, сколько ты раздражал Господа, Бога твоего, в пустыне: с самого того дня, как вышел ты из земли Египетской, и до самого прихода вашего на место сие вы противились Господу.
DEUT|9|8|И при Хориве вы раздражали Господа, и прогневался на вас Господь, так что [хотел] истребить вас,
DEUT|9|9|когда я взошел на гору, чтобы принять скрижали каменные, скрижали завета, который поставил Господь с вами, и пробыл на горе сорок дней и сорок ночей, хлеба не ел и воды не пил,
DEUT|9|10|и дал мне Господь две скрижали каменные, написанные перстом Божиим, а на них все слова, которые изрек вам Господь на горе из среды огня в день собрания.
DEUT|9|11|По окончании же сорока дней и сорока ночей дал мне Господь две скрижали каменные, скрижали завета,
DEUT|9|12|и сказал мне Господь: встань, пойди скорее отсюда, ибо развратился народ твой, который ты вывел из Египта; скоро уклонились они от пути, который Я заповедал им; они сделали себе литый истукан.
DEUT|9|13|И сказал мне Господь: вижу Я народ сей, вот он народ жестоковыйный;
DEUT|9|14|не удерживай Меня, и Я истреблю их, и изглажу имя их из поднебесной, а от тебя произведу народ, [который будет] сильнее и многочисленнее их.
DEUT|9|15|Я обратился и пошел с горы, гора же горела огнем; две скрижали завета [были] в обеих руках моих;
DEUT|9|16|и видел я, что вы согрешили против Господа, Бога вашего, сделали себе литого тельца, скоро уклонились от пути, которого [держаться] заповедал вам Господь;
DEUT|9|17|и взял я обе скрижали, и бросил их из обеих рук своих, и разбил их пред глазами вашими.
DEUT|9|18|И повергшись пред Господом, молился я, как прежде, сорок дней и сорок ночей, хлеба не ел и воды не пил, за все грехи ваши, которыми вы согрешили, сделав зло в очах Господа и раздражив Его;
DEUT|9|19|ибо я страшился гнева и ярости, которыми Господь прогневался на вас [и хотел] погубить вас. И послушал меня Господь и на сей раз.
DEUT|9|20|И на Аарона весьма прогневался Господь [и хотел] погубить его; но я молился и за Аарона в то время.
DEUT|9|21|Грех же ваш, который вы сделали, – тельца я взял, сожег его в огне, разбил его и всего истер до того, что он стал мелок, как прах, и я бросил прах сей в поток, текущий с горы.
DEUT|9|22|И в Тавере, в Массе и в Киброт–Гаттааве вы раздражили Господа.
DEUT|9|23|И когда посылал вас Господь из Кадес–Варни, говоря: пойдите, овладейте землею, которую Я даю вам, – то вы воспротивились повелению Господа Бога вашего, и не поверили Ему, и не послушали гласа Его.
DEUT|9|24|Вы были непокорны Господу с того самого дня, как я стал знать вас.
DEUT|9|25|И повергшись пред Господом, умолял я сорок дней и сорок ночей, в которые я молился, ибо Господь хотел погубить вас;
DEUT|9|26|и молился я Господу и сказал: Владыка Господи, не погубляй народа Твоего и удела Твоего, который Ты избавил величием [крепости] Твоей, который вывел Ты из Египта рукою сильною.
DEUT|9|27|вспомни рабов Твоих, Авраама, Исаака и Иакова; не смотри на ожесточение народа сего и на нечестие его и на грехи его,
DEUT|9|28|дабы [живущие] в той земле, откуда Ты вывел нас, не сказали: "Господь не мог ввести их в землю, которую обещал им, и, ненавидя их, вывел Он их, чтоб умертвить их в пустыне".
DEUT|9|29|А они Твой народ и Твой удел, который Ты вывел [из земли Египетской] силою Твоею великою и мышцею Твоею высокою.
DEUT|10|1|В то время сказал мне Господь: вытеши себе две скрижали каменные, подобные первым, и взойди ко Мне на гору, и сделай себе деревянный ковчег;
DEUT|10|2|и Я напишу на скрижалях те слова, которые были на прежних скрижалях, которые ты разбил; и положи их в ковчег.
DEUT|10|3|И сделал я ковчег из дерева ситтим, и вытесал две каменные скрижали, как прежние, и пошел на гору; и две сии скрижали [были] в руках моих.
DEUT|10|4|И написал Он на скрижалях, как написано было прежде, те десять слов, которые изрек вам Господь на горе из среды огня в день собрания, и отдал их Господь мне.
DEUT|10|5|И обратился я, и сошел с горы, и положил скрижали в ковчег, который я сделал, чтоб они там были, как повелел мне Господь.
DEUT|10|6|И сыны Израилевы отправились из Беероф–Бене–Яакана в Мозер; там умер Аарон и погребен там, и стал священником вместо него сын его Елеазар.
DEUT|10|7|Оттуда отправились в Гудгод, из Гудгода в Иотвафу, в землю, где потоки вод.
DEUT|10|8|В то время отделил Господь колено Левиино, чтобы носить ковчег завета Господня, предстоять пред Господом, служить Ему и благословлять именем Его, [как это продолжается] до сего дня;
DEUT|10|9|потому нет левиту части и удела с братьями его: Сам Господь есть удел его, как говорил ему Господь, Бог твой.
DEUT|10|10|И пробыл я на горе, как и в прежнее время, сорок дней и сорок ночей; и послушал меня Господь и на сей раз, [и] не восхотел Господь погубить тебя;
DEUT|10|11|и сказал мне Господь: встань, пойди в путь пред народом [сим]; пусть они пойдут и овладеют землею, которую Я клялся отцам их дать им.
DEUT|10|12|Итак, Израиль, чего требует от тебя Господь, Бог твой? Того только, чтобы ты боялся Господа, Бога твоего, ходил всеми путями Его, и любил Его, и служил Господу, Богу твоему, от всего сердца твоего и от всей души твоей,
DEUT|10|13|чтобы соблюдал заповеди Господа и постановления Его, которые сегодня заповедую тебе, дабы тебе было хорошо.
DEUT|10|14|Вот у Господа, Бога твоего, небо и небеса небес, земля и все, что на ней;
DEUT|10|15|но только отцов твоих принял Господь и возлюбил их, и избрал вас, семя их после них, из всех народов, как ныне [видишь].
DEUT|10|16|Итак обрежьте крайнюю плоть сердца вашего и не будьте впредь жестоковыйны;
DEUT|10|17|ибо Господь, Бог ваш, есть Бог богов и Владыка владык, Бог великий, сильный и страшный, Который не смотрит на лица и не берет даров,
DEUT|10|18|Который дает суд сироте и вдове, и любит пришельца, и дает ему хлеб и одежду.
DEUT|10|19|Любите и вы пришельца, ибо [сами] были пришельцами в земле Египетской.
DEUT|10|20|Господа, Бога твоего, бойся [и] Ему [одному] служи, и к Нему прилепись и Его именем клянись:
DEUT|10|21|Он хвала твоя и Он Бог твой, Который сделал с тобою те великие и страшные [дела], какие видели глаза твои;
DEUT|10|22|в семидесяти душах пришли отцы твои в Египет, а ныне Господь Бог твой, сделал тебя многочисленным, как звезды небесные.
DEUT|11|1|Итак люби Господа, Бога твоего, и соблюдай, что повелено Им соблюдать, и постановления Его и законы Его и заповеди Его во все дни.
DEUT|11|2|И вспомните ныне, – ибо [я говорю] не с сынами вашими, которые не знают и не видели наказания Господа Бога вашего, – Его величие Его крепкую руку и высокую мышцу его,
DEUT|11|3|знамения Его и дела Его, которые Он сделал среди Египта с фараоном, царем Египетским, и со всею землею его,
DEUT|11|4|и что Он сделал с войском Египетским, с конями его и колесницами его, которых Он потопил в водах Чермного моря, когда они гнались за вами, – и погубил их Господь даже до сего дня;
DEUT|11|5|и что Он делал для вас в пустыне, доколе вы не дошли до места сего,
DEUT|11|6|и что Он сделал с Дафаном и Авироном, сынами Елиава, сына Рувимова, когда земля разверзла уста свои и среди всего Израиля поглотила их и семейства их, и шатры их, и все имущество их, которое было у них;
DEUT|11|7|ибо глаза ваши видели все великие дела Господа, которые Он сделал.
DEUT|11|8|Итак соблюдайте все заповеди [Его], которые я заповедую вам сегодня, дабы вы укрепились и пошли и овладели землею, в которую вы переходите, чтоб овладеть ею;
DEUT|11|9|и дабы вы жили много времени на той земле, которую клялся Господь отцам вашим дать им и семени их, на земле, в которой течет молоко и мед.
DEUT|11|10|Ибо земля, в которую ты идешь, чтоб овладеть ею, не такова, как земля Египетская, из которой вышли вы, где ты, посеяв семя твое, поливал [ее] при помощи ног твоих, как масличный сад;
DEUT|11|11|но земля, в которую вы переходите, чтоб овладеть ею, есть земля с горами и долинами, и от дождя небесного напояется водою, –
DEUT|11|12|земля, о которой Господь, Бог твой, печется: очи Господа, Бога твоего, непрестанно на ней, от начала года и до конца года.
DEUT|11|13|Если вы будете слушать заповеди Мои, которые заповедую вам сегодня, любить Господа, Бога вашего, и служить Ему от всего сердца вашего и от всей души вашей,
DEUT|11|14|то дам земле вашей дождь в свое время, ранний и поздний; и ты соберешь хлеб твой и вино твое и елей твой;
DEUT|11|15|и дам траву на поле твоем для скота твоего, и будешь есть и насыщаться.
DEUT|11|16|Берегитесь, чтобы не обольстилось сердце ваше, и вы не уклонились и не стали служить иным богам и не поклонились им;
DEUT|11|17|и тогда воспламенится гнев Господа на вас, и заключит Он небо, и не будет дождя, и земля не принесет произведений своих, и вы скоро погибнете с доброй земли, которую Господь дает вам.
DEUT|11|18|Итак положите сии слова Мои в сердце ваше и в душу вашу, и навяжите их в знак на руку свою, и да будут они повязкою над глазами вашими;
DEUT|11|19|и учите им сыновей своих, говоря о них, когда ты сидишь в доме твоем, и когда идешь дорогою, и когда ложишься, и когда встаешь;
DEUT|11|20|и напиши их на косяках дома твоего и на воротах твоих,
DEUT|11|21|дабы столько же много было дней ваших и дней детей ваших на той земле, которую Господь клялся дать отцам вашим, сколько дней небо будет над землею.
DEUT|11|22|Ибо если вы будете соблюдать все заповеди сии, которые заповедую вам исполнять, будете любить Господа, Бога вашего, ходить всеми путями Его и прилепляться к Нему,
DEUT|11|23|то изгонит Господь все народы сии от лица вашего, и вы овладеете народами, которые больше и сильнее вас;
DEUT|11|24|всякое место, на которое ступит нога ваша, будет ваше; от пустыни и Ливана, от реки, реки Евфрата, даже до моря западного будут пределы ваши;
DEUT|11|25|никто не устоит против вас: Господь, Бог ваш, наведет страх и трепет пред вами на всякую землю, на которую вы ступите, как Он говорил вам.
DEUT|11|26|Вот, я предлагаю вам сегодня благословение и проклятие:
DEUT|11|27|благословение, если послушаете заповедей Господа, Бога вашего, которые я заповедую вам сегодня,
DEUT|11|28|а проклятие, если не послушаете заповедей Господа, Бога вашего, и уклонитесь от пути, который заповедую вам сегодня, и пойдете вслед богов иных, которых вы не знаете.
DEUT|11|29|Когда введет тебя Господь, Бог твой, в ту землю, в которую ты идешь, чтоб овладеть ею, тогда произнеси благословение на горе Гаризим, а проклятие на горе Гевал:
DEUT|11|30|вот они за Иорданом, по дороге к захождению солнца, в земле Хананеев, живущих на равнине, против Галгала, близ дубравы Море.
DEUT|11|31|Ибо вы переходите Иордан, чтобы пойти овладеть землею, которую Господь, Бог ваш, дает вам, и овладеете ею и будете жить на ней.
DEUT|11|32|Итак старайтесь соблюдать все постановления и законы [Его], которые предлагаю я вам сегодня.
DEUT|12|1|Вот постановления и законы, которые вы должны стараться исполнять в земле, которую Господь, Бог отцов твоих, дает тебе во владение, во все дни, которые вы будете жить на той земле.
DEUT|12|2|Истребите все места, где народы, которыми вы овладеете, служили богам своим, на высоких горах и на холмах, и под всяким ветвистым деревом;
DEUT|12|3|и разрушьте жертвенники их, и сокрушите столбы их, и сожгите огнем рощи их, и разбейте истуканы богов их, и истребите имя их от места того.
DEUT|12|4|Не то должны вы делать для Господа, Бога вашего;
DEUT|12|5|но к месту, какое изберет Господь, Бог ваш, из всех колен ваших, чтобы пребывать имени Его там, обращайтесь и туда приходите,
DEUT|12|6|и туда приносите всесожжения ваши, и жертвы ваши, и десятины ваши, и возношение рук ваших, и обеты ваши, и добровольные приношения ваши, и первенцев крупного скота вашего и мелкого скота вашего;
DEUT|12|7|и ешьте там пред Господом, Богом вашим, и веселитесь вы и семейства ваши о всем, что делалось руками вашими, чем благословил тебя Господь, Бог твой.
DEUT|12|8|Там вы не должны делать всего, как мы теперь здесь делаем, каждый, что ему кажется правильным;
DEUT|12|9|ибо вы ныне еще не вступили в место покоя и в удел, который Господь, Бог твой, дает тебе.
DEUT|12|10|Но когда перейдете Иордан и поселитесь на земле, которую Господь, Бог ваш, дает вам в удел, и когда Он успокоит вас от всех врагов ваших, окружающих [вас], и будете жить безопасно,
DEUT|12|11|тогда, какое место изберет Господь, Бог ваш, чтобы пребывать имени Его там, туда приносите все, что я заповедую вам: всесожжения ваши и жертвы ваши, десятины ваши и возношение рук ваших, и все, избранное по обетам вашим, что вы обещали Господу;
DEUT|12|12|и веселитесь пред Господом, Богом вашим, вы и сыны ваши, и дочери ваши, и рабы ваши, и рабыни ваши, и левит, который посреди жилищ ваших, ибо нет ему части и удела с вами.
DEUT|12|13|Берегись приносить всесожжения твои на всяком месте, которое ты увидишь;
DEUT|12|14|но на том только месте, которое изберет Господь, в одном из колен твоих, приноси всесожжения твои и делай все, что заповедую тебе.
DEUT|12|15|Впрочем, когда только пожелает душа твоя, можешь заколать и есть, по благословению Господа, Бога твоего, мясо, которое Он дал тебе, во всех жилищах твоих: нечистый и чистый могут есть сие, как серну и как оленя;
DEUT|12|16|только крови не ешьте: на землю выливайте ее, как воду.
DEUT|12|17|Нельзя тебе есть в жилищах твоих десятины хлеба твоего, и вина твоего, и елея твоего, и первенцев крупного скота твоего и мелкого скота твоего, и всех обетов твоих, которые ты обещал, и добровольных приношений твоих, и возношения рук твоих;
DEUT|12|18|но ешь сие пред Господом, Богом твоим, на том месте, которое изберет Господь, Бог твой, – ты и сын твой, и дочь твоя, и раб твой, и раба твоя, и левит, [и пришелец], который в жилищах твоих, и веселись пред Господом, Богом твоим, о всем, что делалось руками твоими.
DEUT|12|19|Смотри, не оставляй левита во все дни, [которые будешь жить] на земле твоей.
DEUT|12|20|Когда распространит Господь, Бог твой, пределы твои, как Он говорил тебе, и ты скажешь: "поем я мяса", потому что душа твоя пожелает есть мяса, – тогда, по желанию души твоей, ешь мясо.
DEUT|12|21|Если далеко будет от тебя то место, которое изберет Господь, Бог твой, чтобы пребывать имени Его там, то заколай из крупного и мелкого скота твоего, который дал тебе Господь, как я повелел тебе, и ешь в жилищах твоих, по желанию души твоей;
DEUT|12|22|но ешь их так, как едят серну и оленя; нечистый как и чистый могут есть сие;
DEUT|12|23|только строго наблюдай, чтобы не есть крови, потому что кровь есть душа: не ешь души вместе с мясом;
DEUT|12|24|не ешь ее: выливай ее на землю, как воду;
DEUT|12|25|не ешь ее, дабы хорошо было тебе и детям твоим после тебя, если будешь делать справедливое пред очами Господа.
DEUT|12|26|Только святыни твои, какие будут у тебя, и обеты твои приноси, и приходи на то место, которое изберет Господь.
DEUT|12|27|и совершай всесожжения твои, мясо и кровь, на жертвеннике Господа, Бога твоего; но кровь [других] жертв твоих должна быть проливаема у жертвенника Господа, Бога твоего, а мясо ешь.
DEUT|12|28|Слушай и исполняй все слова сии, которые заповедую тебе, дабы хорошо было тебе и детям твоим после тебя во век, если будешь делать доброе и угодное пред очами Господа, Бога твоего.
DEUT|12|29|Когда Господь, Бог твой, истребит от лица твоего народы, к которым ты идешь, чтобы взять их во владение, и ты, взяв их, поселишься в земле их;
DEUT|12|30|тогда берегись, чтобы ты не попал в сеть, последуя им, по истреблении их от лица твоего, и не искал богов их, говоря: "как служили народы сии богам своим, так буду и я делать";
DEUT|12|31|не делай так Господу, Богу твоему, ибо все, чего гнушается Господь, что ненавидит Он, они делают богам своим: они и сыновей своих и дочерей своих сожигают на огне богам своим.
DEUT|13|1|Все, что я заповедую вам, старайтесь исполнить; не прибавляй к тому и не убавляй от того.
DEUT|13|2|Если восстанет среди тебя пророк, или сновидец, и представит тебе знамение или чудо,
DEUT|13|3|и сбудется то знамение или чудо, о котором он говорил тебе, и скажет притом: "пойдем вслед богов иных, которых ты не знаешь, и будем служить им", –
DEUT|13|4|то не слушай слов пророка сего, или сновидца сего; ибо [чрез] [сие] искушает вас Господь, Бог ваш, чтобы узнать, любите ли вы Господа, Бога вашего, от всего сердца вашего и от всей души вашей;
DEUT|13|5|Господу, Богу вашему, последуйте и Его бойтесь, заповеди Его соблюдайте и гласа Его слушайте, и Ему служите, и к Нему прилепляйтесь;
DEUT|13|6|а пророка того или сновидца того должно предать смерти за то, что он уговаривал вас отступить от Господа, Бога вашего, выведшего вас из земли Египетской и избавившего тебя из дома рабства, желая совратить тебя с пути, по которому заповедал тебе идти Господь, Бог твой; и [так] истреби зло из среды себя.
DEUT|13|7|Если будет уговаривать тебя тайно брат твой, сын матери твоей, или сын твой, или дочь твоя, или жена на лоне твоем, или друг твой, который для тебя, как душа твоя, говоря: "пойдем и будем служить богам иным, которых не знал ты и отцы твои",
DEUT|13|8|богам тех народов, которые вокруг тебя, близких к тебе или отдаленных от тебя, от одного края земли до другого, –
DEUT|13|9|то не соглашайся с ним и не слушай его; и да не пощадит его глаз твой, не жалей его и не прикрывай его,
DEUT|13|10|но убей его; твоя рука прежде [всех] должна быть на нем, чтоб убить его, а потом руки всего народа;
DEUT|13|11|побей его камнями до смерти, ибо он покушался отвратить тебя от Господа, Бога твоего, Который вывел тебя из земли Египетской, из дома рабства;
DEUT|13|12|весь Израиль услышит сие и убоится, и не станут впредь делать среди тебя такого зла.
DEUT|13|13|Если услышишь о каком–либо из городов твоих, которые Господь, Бог твой, дает тебе для жительства,
DEUT|13|14|что появились в нем нечестивые люди из среды тебя и соблазнили жителей города их, говоря: "пойдем и будем служить богам иным, которых вы не знали", –
DEUT|13|15|то ты разыщи, исследуй и хорошо расспроси; и если это точная правда, что случилась мерзость сия среди тебя,
DEUT|13|16|порази жителей того города острием меча, предай заклятию его и все, что в нем, и скот его [порази] острием меча;
DEUT|13|17|всю же добычу его собери на средину площади его и сожги огнем город и всю добычу его во всесожжение Господу, Богу твоему, и да будет он вечно в развалинах, не должно никогда вновь созидать его;
DEUT|13|18|ничто из заклятого да не прилипнет к руке твоей, дабы укротил Господь ярость гнева Своего, и дал тебе милость и помиловал тебя, и размножил тебя, как клялся отцам твоим,
DEUT|13|19|если будешь слушать гласа Господа, Бога твоего, соблюдая все заповеди Его, которые ныне заповедую тебе, делая угодное пред очами Господа, Бога твоего.
DEUT|14|1|Вы сыны Господа Бога вашего; не делайте нарезов [на теле] [вашем] и не выстригайте волос над глазами вашими по умершем;
DEUT|14|2|ибо ты народ святой у Господа Бога твоего, и тебя избрал Господь, чтобы ты был собственным Его народом из всех народов, которые на земле.
DEUT|14|3|Не ешь никакой мерзости.
DEUT|14|4|Вот скот, который вам можно есть: волы, овцы, козы,
DEUT|14|5|олень и серна, и буйвол, и лань, и зубр, и орикс, и камелопард.
DEUT|14|6|Всякий скот, у которого раздвоены копыта и на обоих копытах глубокий разрез, и который скот жует жвачку, тот ешьте;
DEUT|14|7|только сих не ешьте из жующих жвачку и имеющих раздвоенные копыта с глубоким разрезом: верблюда, зайца и тушканчика, потому что, хотя они жуют жвачку, но копыта у них не раздвоены: нечисты они для вас;
DEUT|14|8|и свиньи, потому что копыта у нее раздвоены, но не жует жвачки: нечиста она для вас; не ешьте мяса их, и к трупам их не прикасайтесь.
DEUT|14|9|Из всех [животных], которые в воде, ешьте всех, у которых есть перья и чешуя;
DEUT|14|10|а всех тех, у которых нет перьев и чешуи, не ешьте: нечисто это для вас.
DEUT|14|11|Всякую птицу чистую ешьте;
DEUT|14|12|но сих не должно вам есть из них: орла, грифа и морского орла,
DEUT|14|13|и коршуна, и сокола, и кречета с породою их,
DEUT|14|14|и всякого ворона с породою его,
DEUT|14|15|и страуса, и совы, и чайки, и ястреба с породою его,
DEUT|14|16|и филина, и ибиса, и лебедя,
DEUT|14|17|и пеликана, и сипа, и рыболова,
DEUT|14|18|и цапли, и зуя с породою его, и удода, и нетопыря.
DEUT|14|19|Все крылатые пресмыкающиеся нечисты для вас, не ешьте [их].
DEUT|14|20|Всякую птицу чистую ешьте.
DEUT|14|21|Не ешьте никакой мертвечины; иноземцу, который [случится] в жилищах твоих, отдай ее, он пусть ест ее, или продай ему, ибо ты народ святой у Господа Бога твоего. Не вари козленка в молоке матери его.
DEUT|14|22|Отделяй десятину от всего произведения семян твоих, которое приходит с поля [твоего] каждогодно,
DEUT|14|23|и ешь пред Господом, Богом твоим, на том месте, которое изберет Он, чтобы пребывать имени Его там; десятину хлеба твоего, вина твоего и елея твоего, и первенцев крупного скота твоего и мелкого скота твоего, дабы ты научился бояться Господа, Бога твоего, во все дни.
DEUT|14|24|Если же длинна будет для тебя дорога, так что ты не можешь нести сего, потому что далеко от тебя то место, которое изберет Господь, Бог твой, чтоб положить там имя Свое, и Господь, Бог твой, благословил тебя,
DEUT|14|25|то променяй это на серебро и возьми серебро в руку твою и приходи на место, которое изберет Господь, Бог твой;
DEUT|14|26|и покупай на серебро сие всего, чего пожелает душа твоя, волов, овец, вина, сикера и всего, чего потребует от тебя душа твоя; и ешь там пред Господом, Богом твоим, и веселись ты и семейство твое.
DEUT|14|27|И левита, который в жилищах твоих, не оставь, ибо нет ему части и удела с тобою.
DEUT|14|28|По прошествии же трех лет отделяй все десятины произведений твоих в тот год и клади [сие] в жилищах твоих;
DEUT|14|29|и пусть придет левит, ибо ему нет части и удела с тобою, и пришелец, и сирота, и вдова, которые [находятся] в жилищах твоих, и пусть едят и насыщаются, дабы благословил тебя Господь, Бог твой, во всяком деле рук твоих, которое ты будешь делать.
DEUT|15|1|В седьмой год делай прощение.
DEUT|15|2|Прощение же состоит в том, чтобы всякий заимодавец, который дал взаймы ближнему своему, простил [долг] и не взыскивал с ближнего своего или с брата своего, ибо провозглашено прощение ради Господа.
DEUT|15|3|с иноземца взыскивай, а что будет твое у брата твоего, прости.
DEUT|15|4|Разве только не будет у тебя нищего: ибо благословит тебя Господь на той земле, которую Господь, Бог твой, дает тебе в удел, чтобы ты взял ее в наследство,
DEUT|15|5|если только будешь слушать гласа Господа, Бога твоего, и стараться исполнять все заповеди сии, которые я сегодня заповедую тебе;
DEUT|15|6|ибо Господь, Бог твой, благословит тебя, как Он говорил тебе, и ты будешь давать взаймы многим народам, а сам не будешь брать взаймы; и господствовать будешь над многими народами, а они над тобою не будут господствовать.
DEUT|15|7|Если же будет у тебя нищий кто–либо из братьев твоих, в одном из жилищ твоих, на земле твоей, которую Господь, Бог твой, дает тебе, то не ожесточи сердца твоего и не сожми руки твоей пред нищим братом твоим,
DEUT|15|8|но открой ему руку твою и дай ему взаймы, смотря по его нужде, в чем он нуждается;
DEUT|15|9|берегись, чтобы не вошла в сердце твое беззаконная мысль: "приближается седьмой год, год прощения", и чтоб [от того] глаз твой не сделался немилостив к нищему брату твоему, и ты не отказал ему; ибо он возопиет на тебя к Господу, и будет на тебе грех;
DEUT|15|10|дай ему [взаймы] и когда будешь давать ему, не должно скорбеть сердце твое, ибо за то благословит тебя Господь, Бог твой, во всех делах твоих и во всем, что будет делаться твоими руками;
DEUT|15|11|ибо нищие всегда будут среди земли [твоей]; потому я и повелеваю тебе: отверзай руку твою брату твоему, бедному твоему и нищему твоему на земле твоей.
DEUT|15|12|Если продастся тебе брат твой, Еврей, или Евреянка, то шесть лет должен он быть рабом тебе, а в седьмой год отпусти его от себя на свободу;
DEUT|15|13|когда же будешь отпускать его от себя на свободу, не отпусти его с пустыми [руками],
DEUT|15|14|но снабди его от стад твоих, от гумна твоего и от точила твоего: дай ему, чем благословил тебя Господь, Бог твой:
DEUT|15|15|помни, что [и] ты был рабом в земле Египетской и избавил тебя Господь, Бог твой, потому я сегодня и заповедую тебе сие.
DEUT|15|16|Если же он скажет тебе: "не пойду я от тебя, потому что я люблю тебя и дом твой", потому что хорошо ему у тебя,
DEUT|15|17|то возьми шило и проколи ухо его к двери; и будет он рабом твоим на век. Так поступай и с рабою твоею.
DEUT|15|18|Не считай этого для себя тяжким, что ты должен отпустить его от себя на свободу, ибо он в шесть лет заработал тебе вдвое против платы наемника; и благословит тебя Господь, Бог твой, во всем, что ни будешь делать.
DEUT|15|19|Все первородное мужеского пола, что родится от крупного скота твоего и от мелкого скота твоего, посвящай Господу, Богу твоему: не работай на первородном воле твоем и не стриги первородного из мелкого скота твоего;
DEUT|15|20|пред Господом, Богом твоим, каждогодно съедай это ты и семейство твое, на месте, которое изберет Господь.
DEUT|15|21|если же будет на нем порок, хромота или слепота [или] другой какой–нибудь порок, то не приноси его в жертву Господу, Богу твоему,
DEUT|15|22|но в жилищах твоих ешь его; нечистый, как и чистый, [могут есть], как серну и как оленя;
DEUT|15|23|только крови его не ешь: на землю выливай ее, как воду.
DEUT|16|1|Наблюдай месяц Авив, и совершай Пасху Господу, Богу твоему, потому что в месяце Авиве вывел тебя Господь, Бог твой, из Египта ночью.
DEUT|16|2|И заколай Пасху Господу, Богу твоему, из мелкого и крупного скота на месте, которое изберет Господь, чтобы пребывало там имя Его.
DEUT|16|3|Не ешь с нею квасного; семь дней ешь с нею опресноки, хлебы бедствия, ибо ты с поспешностью вышел из земли Египетской, дабы ты помнил день исшествия своего из земли Египетской во все дни жизни твоей;
DEUT|16|4|не должно находиться у тебя ничто квасное во всем уделе твоем в продолжение семи дней, и из мяса, которое ты принес в жертву вечером в первый день, ничто не должно оставаться до утра.
DEUT|16|5|Не можешь ты заколать Пасху в котором–нибудь из жилищ твоих, которые Господь, Бог твой, даст тебе;
DEUT|16|6|но только на том месте, которое изберет Господь, Бог твой, чтобы пребывало там имя Его, заколай Пасху вечером при захождении солнца, в то самое время, в которое ты вышел из Египта;
DEUT|16|7|и испеки и съешь на том месте, которое изберет Господь, Бог твой, а на другой день можешь возвратиться и войти в шатры твои.
DEUT|16|8|Шесть дней ешь пресные хлебы, а в седьмой день отдание праздника Господу, Богу твоему; не занимайся работою.
DEUT|16|9|Семь седмиц отсчитай себе; начинай считать семь седмиц с того времени, как появится серп на жатве;
DEUT|16|10|тогда совершай праздник седмиц Господу, Богу твоему, по усердию руки твоей, сколько ты дашь, смотря по тому, чем благословит тебя Господь, Бог твой;
DEUT|16|11|и веселись пред Господом, Богом твоим, ты, и сын твой, и дочь твоя, и раб твой, и раба твоя, и левит, который в жилищах твоих, и пришелец, и сирота, и вдова, которые среди тебя, на месте, которое изберет Господь, Бог твой, чтобы пребывало там имя Его;
DEUT|16|12|помни, что ты был рабом в Египте, и соблюдай и исполняй постановления сии.
DEUT|16|13|Праздник кущей совершай у себя семь дней, когда уберешь с гумна твоего и из точила твоего;
DEUT|16|14|и веселись в праздник твой ты и сын твой, и дочь твоя, и раб твой, и раба твоя, и левит, и пришелец, и сирота, и вдова, которые в жилищах твоих;
DEUT|16|15|семь дней празднуй Господу, Богу твоему, на месте, которое изберет Господь, Бог твой; ибо благословит тебя Господь, Бог твой, во всех произведениях твоих и во всяком деле рук твоих, и ты будешь только веселиться.
DEUT|16|16|Три раза в году весь мужеский пол должен являться пред лице Господа, Бога твоего, на место, которое изберет Он: в праздник опресноков, в праздник седмиц и в праздник кущей; и [никто] не должен являться пред лице Господа с пустыми [руками],
DEUT|16|17|но каждый с даром в руке своей, смотря по благословению Господа, Бога твоего, какое Он дал тебе.
DEUT|16|18|Во всех жилищах твоих, которые Господь, Бог твой, даст тебе, поставь себе судей и надзирателей по коленам твоим, чтоб они судили народ судом праведным;
DEUT|16|19|не извращай закона, не смотри на лица и не бери даров, ибо дары ослепляют глаза мудрых и превращают дело правых;
DEUT|16|20|правды, правды ищи, дабы ты был жив и овладел землею, которую Господь, Бог твой, дает тебе.
DEUT|16|21|Не сади себе рощи из каких–либо дерев при жертвеннике Господа, Бога твоего, который ты сделаешь себе,
DEUT|16|22|и не ставь себе столба, что ненавидит Господь Бог твой.
DEUT|17|1|Не приноси в жертву Господу, Богу твоему, вола, или овцы, на которой будет порок, [или] что–нибудь худое, ибо это мерзость для Господа, Бога твоего.
DEUT|17|2|Если найдется среди тебя в каком–либо из жилищ твоих, которые Господь, Бог твой, дает тебе, мужчина или женщина, кто сделает зло пред очами Господа, Бога твоего, преступив завет Его,
DEUT|17|3|и пойдет и станет служить иным богам, и поклонится им, или солнцу, или луне, или всему воинству небесному, чего я не повелел,
DEUT|17|4|и тебе возвещено будет, и ты услышишь, то ты хорошо разыщи; и если это точная правда, если сделана мерзость сия в Израиле,
DEUT|17|5|то выведи мужчину того, или женщину ту, которые сделали зло сие, к воротам твоим и побей их камнями до смерти.
DEUT|17|6|По словам двух свидетелей, или трех свидетелей, должен умереть осуждаемый на смерть: не должно предавать смерти по словам одного свидетеля;
DEUT|17|7|рука свидетелей должна быть на нем прежде [всех], чтоб убить его, потом рука всего народа; и [так] истреби зло из среды себя.
DEUT|17|8|Если по какому делу затруднительным будет для тебя рассудить между кровью и кровью, между судом и судом, между побоями и побоями, [и] [будут] несогласные мнения в воротах твоих, то встань и пойди на место, которое изберет Господь, Бог твой,
DEUT|17|9|и приди к священникам левитам и к судье, который будет в те дни, и спроси их, и они скажут тебе, как рассудить;
DEUT|17|10|и поступи по слову, какое они скажут тебе, на том месте, которое изберет Господь, и постарайся исполнить все, чему они научат тебя;
DEUT|17|11|по закону, которому научат они тебя, и по определению, какое они скажут тебе, поступи, и не уклоняйся ни направо, ни налево от того, что они скажут тебе.
DEUT|17|12|А кто поступит так дерзко, что не послушает священника, стоящего там на служении пред Господом, Богом твоим, или судьи, тот должен умереть, – и [так] истреби зло от Израиля;
DEUT|17|13|и весь народ услышит и убоится, и не будут впредь поступать дерзко.
DEUT|17|14|Когда ты придешь в землю, которую Господь, Бог твой, дает тебе, и овладеешь ею, и поселишься на ней, и скажешь: "поставлю я над собою царя, подобно прочим народам, которые вокруг меня",
DEUT|17|15|то поставь над собою царя, которого изберет Господь, Бог твой; из среды братьев твоих поставь над собою царя; не можешь поставить над собою [царем] иноземца, который не брат тебе.
DEUT|17|16|Только чтоб он не умножал себе коней и не возвращал народа в Египет для умножения себе коней, ибо Господь сказал вам: "не возвращайтесь более путем сим";
DEUT|17|17|и чтобы не умножал себе жен, дабы не развратилось сердце его, и чтобы серебра и золота не умножал себе чрезмерно.
DEUT|17|18|Но когда он сядет на престоле царства своего, должен списать для себя список закона сего с книги, [находящейся] у священников левитов,
DEUT|17|19|и пусть он будет у него, и пусть он читает его во все дни жизни своей, дабы научался бояться Господа, Бога своего, и старался исполнять все слова закона сего и постановления сии;
DEUT|17|20|чтобы не надмевалось сердце его пред братьями его, и чтобы не уклонялся он от закона ни направо, ни налево, дабы долгие дни пребыл на царстве своем он и сыновья его посреди Израиля.
DEUT|18|1|Священникам левитам, всему колену Левиину, не будет части и удела с Израилем: они должны питаться жертвами Господа и Его частью;
DEUT|18|2|удела же не будет ему между братьями его: Сам Господь удел его, как говорил Он ему.
DEUT|18|3|Вот что должно быть положено священникам от народа, от приносящих в жертву волов или овец: должно отдавать священнику плечо, челюсти и желудок;
DEUT|18|4|также начатки от хлеба твоего, вина твоего и елея твоего, и начатки от шерсти овец твоих отдавай ему,
DEUT|18|5|ибо его избрал Господь Бог твой из всех колен твоих, чтобы он предстоял [пред Господом, Богом твоим], служил во имя Господа, сам и сыны его во все дни.
DEUT|18|6|И если левит придет из одного из жилищ твоих, из всей [земли сынов] Израилевых, где он жил, и придет по желанию души своей на место, которое изберет Господь,
DEUT|18|7|и будет служить во имя Господа Бога своего, как и все братья его левиты, предстоящие там пред Господом, –
DEUT|18|8|то пусть они пользуются одинаковою частью, сверх полученного от продажи отцовского [имущества].
DEUT|18|9|Когда ты войдешь в землю, которую дает тебе Господь Бог твой, тогда не научись делать мерзости, какие делали народы сии:
DEUT|18|10|не должен находиться у тебя проводящий сына своего или дочь свою чрез огонь, прорицатель, гадатель, ворожея, чародей,
DEUT|18|11|обаятель, вызывающий духов, волшебник и вопрошающий мертвых;
DEUT|18|12|ибо мерзок пред Господом всякий, делающий это, и за сии–то мерзости Господь Бог твой изгоняет их от лица твоего;
DEUT|18|13|будь непорочен пред Господом Богом твоим;
DEUT|18|14|ибо народы сии, которых ты изгоняешь, слушают гадателей и прорицателей, а тебе не то дал Господь Бог твой.
DEUT|18|15|Пророка из среды тебя, из братьев твоих, как меня, воздвигнет тебе Господь Бог твой, – Его слушайте, –
DEUT|18|16|так как ты просил у Господа Бога твоего при Хориве в день собрания, говоря: да не услышу впредь гласа Господа Бога моего и огня сего великого да не увижу более, дабы мне не умереть.
DEUT|18|17|И сказал мне Господь: хорошо то, что они говорили.
DEUT|18|18|Я воздвигну им Пророка из среды братьев их, такого как ты, и вложу слова Мои в уста Его, и Он будет говорить им все, что Я повелю Ему;
DEUT|18|19|а кто не послушает слов Моих, которые [Пророк тот] будет говорить Моим именем, с того Я взыщу;
DEUT|18|20|но пророка, который дерзнет говорить Моим именем то, чего Я не повелел ему говорить, и который будет говорить именем богов иных, такого пророка предайте смерти.
DEUT|18|21|И если скажешь в сердце твоем: "как мы узнаем слово, которое не Господь говорил?"
DEUT|18|22|Если пророк скажет именем Господа, но слово то не сбудется и не исполнится, то не Господь говорил сие слово, но говорил сие пророк по дерзости своей, – не бойся его.
DEUT|19|1|Когда Господь Бог твой истребит народы, которых землю дает тебе Господь Бог твой и ты вступишь в наследие после них, и поселишься в городах их и домах их,
DEUT|19|2|тогда отдели себе три города среди земли твоей, которую Господь Бог твой дает тебе во владение;
DEUT|19|3|устрой себе дорогу и раздели на три части всю землю твою, которую Господь Бог твой дает тебе в удел; они будут служить убежищем всякому убийце.
DEUT|19|4|И вот какой убийца может убегать туда и остаться жив: кто убьет ближнего своего без намерения, не быв врагом ему вчера и третьего дня;
DEUT|19|5|кто пойдет с ближним своим в лес рубить дрова, и размахнется рука его с топором, чтобы срубить дерево, и соскочит железо с топорища и попадет в ближнего, и он умрет, – такой пусть убежит в один из городов тех, чтоб остаться живым,
DEUT|19|6|дабы мститель за кровь в горячности сердца своего не погнался за убийцею и не настиг его, если далек будет путь, и не убил его, между тем как он не [подлежит] осуждению на смерть, ибо не был врагом ему вчера и третьего дня;
DEUT|19|7|посему я и дал тебе повеление, говоря: отдели себе три города.
DEUT|19|8|Когда же Господь Бог твой распространит пределы твои, как Он клялся отцам твоим, и даст тебе всю землю, которую Он обещал дать отцам твоим,
DEUT|19|9|если ты будешь стараться исполнять все сии заповеди, которые я заповедую тебе сегодня, любить Господа Бога твоего и ходить путями Его во все дни, – тогда к сим трем городам прибавь еще три города,
DEUT|19|10|дабы не проливалась кровь невинного среди земли твоей, которую Господь Бог твой дает тебе в удел, и чтобы не было на тебе [вины] крови.
DEUT|19|11|Но если кто будет врагом ближнему своему и будет подстерегать его, и восстанет на него и убьет его до смерти, и убежит в один из городов тех,
DEUT|19|12|то старейшины города его должны послать, чтобы взять его оттуда и предать его в руки мстителя за кровь, чтоб он умер;
DEUT|19|13|да не пощадит его глаз твой; смой с Израиля кровь невинного, и будет тебе хорошо.
DEUT|19|14|Не нарушай межи ближнего твоего, которую положили предки в уделе твоем, доставшемся тебе в земле, которую Господь Бог твой дает тебе во владение.
DEUT|19|15|Недостаточно одного свидетеля против кого–либо в какой – нибудь вине и в каком–нибудь преступлении и в каком–нибудь грехе, которым он согрешит: при словах двух свидетелей, или при словах трех свидетелей состоится дело.
DEUT|19|16|Если выступит против кого свидетель несправедливый, обвиняя его в преступлении,
DEUT|19|17|то пусть предстанут оба сии человека, у которых тяжба, пред Господа, пред священников и пред судей, которые будут в те дни;
DEUT|19|18|судьи должны хорошо исследовать, и если свидетель тот свидетель ложный, ложно донес на брата своего,
DEUT|19|19|то сделайте ему то, что он умышлял сделать брату своему; и [так] истреби зло из среды себя;
DEUT|19|20|и прочие услышат, и убоятся, и не станут впредь делать такое зло среди тебя;
DEUT|19|21|да не пощадит [его] глаз твой: душу за душу, глаз за глаз, зуб за зуб, руку за руку, ногу за ногу.
DEUT|20|1|Когда ты выйдешь на войну против врага твоего и увидишь коней и колесницы [и] народа более, нежели у тебя, то не бойся их, ибо с тобою Господь Бог твой, Который вывел тебя из земли Египетской.
DEUT|20|2|Когда же приступаете к сражению, тогда пусть подойдет священник, и говорит народу,
DEUT|20|3|и скажет ему: слушай, Израиль! вы сегодня вступаете в сражение с врагами вашими, да не ослабеет сердце ваше, не бойтесь, не смущайтесь и не ужасайтесь их,
DEUT|20|4|ибо Господь Бог ваш идет с вами, чтобы сразиться за вас с врагами вашими [и] спасти вас.
DEUT|20|5|Надзиратели же пусть объявят народу, говоря: кто построил новый дом и не обновил его, тот пусть идет и возвратится в дом свой, дабы не умер на сражении, и другой не обновил его;
DEUT|20|6|и кто насадил виноградник и не пользовался им, тот пусть идет и возвратится в дом свой, дабы не умер на сражении, и другой не воспользовался им;
DEUT|20|7|и кто обручился с женою и не взял ее, тот пусть идет и возвратится в дом свой, дабы не умер на сражении, и другой не взял ее.
DEUT|20|8|И еще объявят надзиратели народу, и скажут: кто боязлив и малодушен, тот пусть идет и возвратится в дом свой, дабы он не сделал робкими сердца братьев его, как его сердце.
DEUT|20|9|Когда надзиратели скажут все это народу, тогда должно поставить военных начальников в вожди народу.
DEUT|20|10|Когда подойдешь к городу, чтобы завоевать его, предложи ему мир;
DEUT|20|11|если он согласится на мир с тобою и отворит тебе [ворота], то весь народ, который найдется в нем, будет платить тебе дань и служить тебе;
DEUT|20|12|если же он не согласится на мир с тобою и будет вести с тобою войну, то осади его,
DEUT|20|13|и [когда] Господь Бог твой предаст его в руки твои, порази в нем весь мужеский пол острием меча;
DEUT|20|14|только жен и детей и скот и все, что в городе, всю добычу его возьми себе и пользуйся добычею врагов твоих, которых предал тебе Господь Бог твой;
DEUT|20|15|так поступай со всеми городами, которые от тебя весьма далеко, которые не из [числа] городов народов сих.
DEUT|20|16|А в городах сих народов, которых Господь Бог твой дает тебе во владение, не оставляй в живых ни одной души,
DEUT|20|17|но предай их заклятию: Хеттеев и Аморреев, и Хананеев, и Ферезеев, и Евеев, и Иевусеев, как повелел тебе Господь Бог твой,
DEUT|20|18|дабы они не научили вас делать такие же мерзости, какие они делали для богов своих, и дабы вы не грешили пред Господом Богом вашим.
DEUT|20|19|Если долгое время будешь держать в осаде [какой–нибудь] город, чтобы завоевать его и взять его, то не порти дерев его, от которых можно питаться, и не опустошай окрестностей, ибо дерево на поле не человек, чтобы могло уйти от тебя в укрепление;
DEUT|20|20|только те дерева, о которых ты знаешь, что они ничего не приносят в пищу, можешь портить и рубить, и строить укрепление против города, который ведет с тобою войну, доколе не покоришь его.
DEUT|21|1|Если в земле, которую Господь Бог твой, дает тебе во владение, найден будет убитый, лежащий на поле, и неизвестно, кто убил его,
DEUT|21|2|то пусть выйдут старейшины твои и судьи твои и измерят [расстояние] до городов, которые вокруг убитого;
DEUT|21|3|и старейшины города того, который будет ближайшим к убитому, пусть возьмут телицу, на которой не работали, [и] которая не носила ярма,
DEUT|21|4|и пусть старейшины того города отведут сию телицу в дикую долину, которая не разработана и не засеяна, и заколют там телицу в долине;
DEUT|21|5|и придут священники, сыны Левиины;
DEUT|21|6|и все старейшины города того, ближайшие к убитому, пусть омоют руки свои над [головою] телицы, зарезанной в долине,
DEUT|21|7|и объявят и скажут: руки наши не пролили крови сей, и глаза наши не видели;
DEUT|21|8|очисти народ Твой, Израиля, который Ты, Господи, освободил, и не вмени народу Твоему, Израилю, невинной крови. И они очистятся от крови.
DEUT|21|9|[Так] должен ты смывать у себя кровь невинного, если хочешь делать [доброе и] справедливое пред очами Господа.
DEUT|21|10|Когда выйдешь на войну против врагов твоих, и Господь Бог твой предаст их в руки твои, и возьмешь их в плен,
DEUT|21|11|и увидишь между пленными женщину, красивую видом, и полюбишь ее, и захочешь взять ее себе в жену,
DEUT|21|12|то приведи ее в дом свой, и пусть она острижет голову свою и обрежет ногти свои,
DEUT|21|13|и снимет с себя пленническую одежду свою, и живет в доме твоем, и оплакивает отца своего и матерь свою в продолжение месяца; и после того ты можешь войти к ней и сделаться ее мужем, и она будет твоею женою;
DEUT|21|14|если же она [после] не понравится тебе, то отпусти ее, [куда] она захочет, но не продавай ее за серебро и не обращай ее в рабство, потому что ты смирил ее.
DEUT|21|15|Если у кого будут две жены – одна любимая, а другая нелюбимая, и как любимая, [так] и нелюбимая родят ему сыновей, и первенцем будет сын нелюбимой, –
DEUT|21|16|то, при разделе сыновьям своим имения своего, он не может сыну жены любимой дать первенство пред первородным сыном нелюбимой;
DEUT|21|17|но первенцем должен признать сына нелюбимой [и] дать ему двойную часть из всего, что у него найдется, ибо он есть начаток силы его, ему [принадлежит] право первородства.
DEUT|21|18|Если у кого будет сын буйный и непокорный, неповинующийся голосу отца своего и голосу матери своей, и они наказывали его, но он не слушает их, –
DEUT|21|19|то отец его и мать его пусть возьмут его и приведут его к старейшинам города своего и к воротам своего местопребывания
DEUT|21|20|и скажут старейшинам города своего: "сей сын наш буен и непокорен, не слушает слов наших, мот и пьяница";
DEUT|21|21|тогда все жители города его пусть побьют его камнями до смерти; и [так] истреби зло из среды себя, и все Израильтяне услышат и убоятся.
DEUT|21|22|Если в ком найдется преступление, достойное смерти, и он будет умерщвлен, и ты повесишь его на дереве,
DEUT|21|23|то тело его не должно ночевать на дереве, но погреби его в тот же день, ибо проклят пред Богом [всякий] повешенный [на дереве], и не оскверняй земли твоей, которую Господь Бог твой дает тебе в удел.
DEUT|22|1|Когда увидишь вола брата твоего или овцу его заблудившихся, не оставляй их, но возврати их брату твоему;
DEUT|22|2|если же не близко будет к тебе брат твой, или ты не знаешь его, то прибери их в дом свой, и пусть они будут у тебя, доколе брат твой не будет искать их, и тогда возврати ему их;
DEUT|22|3|так поступай и с ослом его, так поступай с одеждой его, так поступай со всякою потерянною [вещью] брата твоего, которая будет им потеряна и которую ты найдешь; нельзя тебе уклоняться [от сего].
DEUT|22|4|Когда увидишь осла брата твоего или вола его упадших на пути, не оставляй их, но подними их с ним вместе.
DEUT|22|5|На женщине не должно быть мужской одежды, и мужчина не должен одеваться в женское платье, ибо мерзок пред Господом Богом твоим всякий делающий сие.
DEUT|22|6|Если попадется тебе на дороге птичье гнездо на каком–либо дереве или на земле, с птенцами или яйцами, и мать сидит на птенцах или на яйцах, то не бери матери вместе с детьми:
DEUT|22|7|мать пусти, а детей возьми себе, чтобы тебе было хорошо, и чтобы продлились дни твои.
DEUT|22|8|Если будешь строить новый дом, то сделай перила около кровли твоей, чтобы не навести тебе крови на дом твой, когда кто – нибудь упадет с него.
DEUT|22|9|Не засевай виноградника своего двумя родами семян, чтобы не сделать тебе заклятым сбора семян, которые ты посеешь вместе с плодами виноградника [своего].
DEUT|22|10|Не паши на воле и осле вместе.
DEUT|22|11|Не надевай одежды, сделанной из разных веществ, из шерсти и льна вместе.
DEUT|22|12|Сделай себе кисточки на четырех углах покрывала твоего, которым ты покрываешься.
DEUT|22|13|Если кто возьмет жену, и войдет к ней, и возненавидит ее,
DEUT|22|14|и будет возводить на нее порочные дела, и пустит о ней худую молву, и скажет: "я взял сию жену, и вошел к ней, и не нашел у нее девства",
DEUT|22|15|то отец отроковицы и мать ее пусть возьмут и вынесут [признаки] девства отроковицы к старейшинам города, к воротам;
DEUT|22|16|и отец отроковицы скажет старейшинам: дочь мою я отдал в жену сему человеку, и [ныне] он возненавидел ее,
DEUT|22|17|и вот, он взводит [на нее] порочные дела, говоря: "я не нашел у дочери твоей девства"; но вот признаки девства дочери моей. И расстелют одежду пред старейшинами города.
DEUT|22|18|Тогда старейшины того города пусть возьмут мужа и накажут его,
DEUT|22|19|и наложат на него сто [сиклей] серебра пени и отдадут отцу отроковицы за то, что он пустил худую молву о девице Израильской; она же пусть останется его женою, и он не может развестись с нею во всю жизнь свою.
DEUT|22|20|Если же сказанное будет истинно, и не найдется девства у отроковицы,
DEUT|22|21|то отроковицу пусть приведут к дверям дома отца ее, и жители города ее побьют ее камнями до смерти, ибо она сделала срамное дело среди Израиля, блудодействовав в доме отца своего; и [так] истреби зло из среды себя.
DEUT|22|22|Если найден будет кто лежащий с женою замужнею, то должно предать смерти обоих: и мужчину, лежавшего с женщиною, и женщину; и [так] истреби зло от Израиля.
DEUT|22|23|Если будет молодая девица обручена мужу, и кто–нибудь встретится с нею в городе и ляжет с нею,
DEUT|22|24|то обоих их приведите к воротам того города, и побейте их камнями до смерти: отроковицу за то, что она не кричала в городе, а мужчину за то, что он опорочил жену ближнего своего; и [так] истреби зло из среды себя.
DEUT|22|25|Если же кто в поле встретится с отроковицею обрученною и, схватив ее, ляжет с нею, то должно предать смерти только мужчину, лежавшего с нею,
DEUT|22|26|а отроковице ничего не делай; на отроковице нет преступления смертного: ибо это то же, как если бы кто восстал на ближнего своего и убил его;
DEUT|22|27|ибо он встретился с нею в поле, и [хотя] отроковица обрученная кричала, но некому было спасти ее.
DEUT|22|28|Если кто–нибудь встретится с девицею необрученною, и схватит ее и ляжет с нею, и застанут их,
DEUT|22|29|то лежавший с нею должен дать отцу отроковицы пятьдесят [сиклей] серебра, а она пусть будет его женою, потому что он опорочил ее; во всю жизнь свою он не может развестись с нею.
DEUT|23|1|Никто не должен брать жены отца своего и открывать край [одежды] отца своего.
DEUT|23|2|У кого раздавлены ятра или отрезан детородный член, тот не может войти в общество Господне.
DEUT|23|3|Сын блудницы не может войти в общество Господне, и десятое поколение его не может войти в общество Господне.
DEUT|23|4|Аммонитянин и Моавитянин не может войти в общество Господне, и десятое поколение их не может войти в общество Господне во веки,
DEUT|23|5|потому что они не встретили вас с хлебом и водою на пути, когда вы шли из Египта, и потому что они наняли против тебя Валаама, сына Веорова, из Пефора Месопотамского, чтобы проклясть тебя;
DEUT|23|6|но Господь, Бог твой, не восхотел слушать Валаама и обратил Господь Бог твой проклятие его в благословение тебе, ибо Господь Бог твой любит тебя.
DEUT|23|7|Не желай им мира и благополучия во все дни твои, во веки.
DEUT|23|8|Не гнушайся Идумеянином, ибо он брат твой; не гнушайся Египтянином, ибо ты был пришельцем в земле его;
DEUT|23|9|дети, которые у них родятся, в третьем поколении могут войти в общество Господне.
DEUT|23|10|Когда пойдешь в поход против врагов твоих, берегись всего худого.
DEUT|23|11|Если у тебя будет кто нечист от случившегося [ему] ночью, то он должен выйти вон из стана и не входить в стан,
DEUT|23|12|а при наступлении вечера должен омыть [тело свое] водою, и по захождении солнца может войти в стан.
DEUT|23|13|Место должно быть у тебя вне стана, куда бы тебе выходить;
DEUT|23|14|кроме оружия твоего должна быть у тебя лопатка; и когда будешь садиться вне [стана], выкопай ею [яму] и опять зарой [ею] испражнение твое;
DEUT|23|15|ибо Господь Бог твой ходит среди стана твоего, чтобы избавлять тебя и предавать врагов твоих [в руки твои], а [посему] стан твой должен быть свят, чтобы Он не увидел у тебя чего срамного и не отступил от тебя.
DEUT|23|16|Не выдавай раба господину его, когда он прибежит к тебе от господина своего;
DEUT|23|17|пусть он у тебя живет, среди вас на месте, которое он изберет в каком–нибудь из жилищ твоих, где ему понравится; не притесняй его.
DEUT|23|18|Не должно быть блудницы из дочерей Израилевых и не должно быть блудника из сынов Израилевых.
DEUT|23|19|Не вноси платы блудницы и цены пса в дом Господа Бога твоего ни по какому обету, ибо то и другое есть мерзость пред Господом Богом твоим.
DEUT|23|20|Не отдавай в рост брату твоему ни серебра, ни хлеба, ни чего–либо другого, что [можно] отдавать в рост;
DEUT|23|21|иноземцу отдавай в рост, а брату твоему не отдавай в рост, чтобы Господь Бог твой благословил тебя во всем, что делается руками твоими, на земле, в которую ты идешь, чтобы овладеть ею.
DEUT|23|22|Если дашь обет Господу Богу твоему, немедленно исполни его, ибо Господь Бог твой взыщет его с тебя, и на тебе будет грех;
DEUT|23|23|если же ты не дал обета, то не будет на тебе греха.
DEUT|23|24|Что вышло из уст твоих, соблюдай и исполняй так, как обещал ты Господу Богу твоему добровольное приношение, о котором сказал ты устами своими.
DEUT|23|25|Когда войдешь в виноградник ближнего твоего, можешь есть ягоды досыта, сколько [хочет] душа твоя, а в сосуд твой не клади.
DEUT|23|26|Когда придешь на жатву ближнего твоего, срывай колосья руками твоими, но серпа не заноси на жатву ближнего твоего.
DEUT|24|1|Если кто возьмет жену и сделается ее мужем, и она не найдет благоволения в глазах его, потому что он находит в ней что–нибудь противное, и напишет ей разводное письмо, и даст ей в руки, и отпустит ее из дома своего,
DEUT|24|2|и она выйдет из дома его, пойдет, и выйдет за другого мужа,
DEUT|24|3|но и сей последний муж возненавидит ее и напишет ей разводное письмо, и даст ей в руки, и отпустит ее из дома своего, или умрет сей последний муж ее, взявший ее себе в жену, –
DEUT|24|4|то не может первый ее муж, отпустивший ее, опять взять ее себе в жену, после того как она осквернена, ибо сие есть мерзость пред Господом, и не порочь земли, которую Господь Бог твой дает тебе в удел.
DEUT|24|5|Если кто взял жену недавно, то пусть не идет на войну, и ничего не должно возлагать на него; пусть он остается свободен в доме своем в продолжение одного года и увеселяет жену свою, которую взял.
DEUT|24|6|Никто не должен брать в залог верхнего и нижнего жернова, ибо таковой берет в залог душу.
DEUT|24|7|Если найдут кого, что он украл кого–нибудь из братьев своих, из сынов Израилевых, и поработил его, и продал его, то такого вора должно предать смерти; и [так] истреби зло из среды себя.
DEUT|24|8|Смотри, в язве проказы тщательно соблюдай и исполняй весь [закон], которому научат вас священники левиты; тщательно исполняйте, что я повелел им;
DEUT|24|9|помни, что Господь Бог твой сделал Мариами на пути, когда вы шли из Египта.
DEUT|24|10|Если ты ближнему твоему дашь что–нибудь взаймы, то не ходи к нему в дом, чтобы взять у него залог,
DEUT|24|11|постой на улице, а тот, которому ты дал взаймы, вынесет тебе залог свой на улицу;
DEUT|24|12|если же он будет человек бедный, то ты не ложись спать, имея залог его:
DEUT|24|13|возврати ему залог при захождении солнца, чтоб он лег спать в одежде своей и благословил тебя, – и тебе поставится [сие] в праведность пред Господом Богом твоим.
DEUT|24|14|Не обижай наемника, бедного и нищего, из братьев твоих или из пришельцев твоих, которые в земле твоей, в жилищах твоих;
DEUT|24|15|в тот же день отдай плату его, чтобы солнце не зашло прежде того, ибо он беден, и ждет ее душа его; чтоб он не возопил на тебя к Господу, и не было на тебе греха.
DEUT|24|16|Отцы не должны быть наказываемы смертью за детей, и дети не должны быть наказываемы смертью за отцов; каждый должен быть наказываем смертью за свое преступление.
DEUT|24|17|Не суди превратно пришельца, сироту; и у вдовы не бери одежды в залог;
DEUT|24|18|помни, что и ты был рабом в Египте, и Господь освободил тебя оттуда: посему я и повелеваю тебе делать сие.
DEUT|24|19|Когда будешь жать на поле твоем, и забудешь сноп на поле, то не возвращайся взять его; пусть он остается пришельцу, сироте и вдове, чтобы Господь Бог твой благословил тебя во всех делах рук твоих.
DEUT|24|20|Когда будешь обивать маслину твою, то не пересматривай за собою ветвей: пусть остается пришельцу, сироте и вдове.
DEUT|24|21|Когда будешь снимать плоды в винограднике твоем, не собирай остатков за собою: пусть остается пришельцу, сироте и вдове;
DEUT|24|22|и помни, что ты был рабом в земле Египетской: посему я и повелеваю тебе делать сие.
DEUT|25|1|Если будет тяжба между людьми, то пусть приведут их в суд и рассудят их, правого пусть оправдают, а виновного осудят;
DEUT|25|2|и если виновный достоин будет побоев, то судья пусть прикажет положить его и бить при себе, смотря по вине его, по счету;
DEUT|25|3|сорок ударов можно дать ему, а не более, чтобы от многих ударов брат твой не был обезображен пред глазами твоими.
DEUT|25|4|Не заграждай рта волу, когда он молотит.
DEUT|25|5|Если братья живут вместе и один из них умрет, не имея у себя сына, то жена умершего не должна выходить на сторону за человека чужого, но деверь ее должен войти к ней и взять ее себе в жену, и жить с нею, –
DEUT|25|6|и первенец, которого она родит, останется с именем брата его умершего, чтоб имя его не изгладилось в Израиле.
DEUT|25|7|Если же он не захочет взять невестку свою, то невестка его пойдет к воротам, к старейшинам, и скажет: "деверь мой отказывается восставить имя брата своего в Израиле, не хочет жениться на мне";
DEUT|25|8|тогда старейшины города его должны призвать его и уговаривать его, и если он станет и скажет: "не хочу взять ее",
DEUT|25|9|[тогда] невестка его пусть пойдет к нему в глазах старейшин, и снимет сапог его с ноги его, и плюнет в лице его, и скажет: "так поступают с человеком, который не созидает дома брату своему".
DEUT|25|10|и нарекут ему имя в Израиле: дом разутого.
DEUT|25|11|Когда дерутся между собою мужчины, и жена одного подойдет, чтобы отнять мужа своего из рук бьющего его, и протянув руку свою, схватит его за срамный уд,
DEUT|25|12|то отсеки руку ее: да не пощадит [ее] глаз твой.
DEUT|25|13|В кисе твоей не должны быть двоякие гири, большие и меньшие;
DEUT|25|14|в доме твоем не должна быть двоякая ефа, большая и меньшая;
DEUT|25|15|гиря у тебя должна быть точная и правильная, и ефа у тебя должна быть точная и правильная, чтобы продлились дни твои на земле, которую Господь Бог твой дает тебе.
DEUT|25|16|ибо мерзок пред Господом Богом твоим всякий делающий неправду.
DEUT|25|17|Помни, как поступил с тобою Амалик на пути, когда вы шли из Египта:
DEUT|25|18|как он встретил тебя на пути, и побил сзади тебя всех ослабевших, когда ты устал и утомился, и не побоялся он Бога;
DEUT|25|19|итак, когда Господь Бог твой успокоит тебя от всех врагов твоих со всех сторон, на земле, которую Господь Бог твой дает тебе в удел, чтоб овладеть ею, изгладь память Амалика из поднебесной; не забудь.
DEUT|26|1|Когда ты придешь в землю, которую Господь Бог твой дает тебе в удел, и овладеешь ею, и поселишься в ней;
DEUT|26|2|то возьми начатков всех плодов земли, которые ты получишь от земли твоей, которую Господь Бог твой дает тебе, и положи в корзину, и пойди на то место, которое Господь Бог твой изберет, чтобы пребывало там имя Его;
DEUT|26|3|и приди к священнику, который будет в те дни, и скажи ему: сегодня исповедую пред Господом Богом твоим, что я вошел в ту землю, которую Господь клялся отцам нашим дать нам.
DEUT|26|4|Священник возьмет корзину из руки твоей и поставит ее пред жертвенником Господа Бога твоего.
DEUT|26|5|Ты же отвечай и скажи пред Господом Богом твоим: отец мой был странствующий Арамеянин, и пошел в Египет и поселился там с немногими людьми, и произошел там от него народ великий, сильный и многочисленный;
DEUT|26|6|но Египтяне худо поступали с нами, и притесняли нас, и налагали на нас тяжкие работы;
DEUT|26|7|и возопили мы к Господу Богу отцов наших, и услышал Господь вопль наш и увидел бедствие наше, труды наши и угнетение наше;
DEUT|26|8|и вывел нас Господь из Египта рукою сильною и мышцею простертою, великим ужасом, знамениями и чудесами,
DEUT|26|9|и привел нас на место сие, и дал нам землю сию, землю, в которой течет молоко и мед;
DEUT|26|10|итак вот, я принес начатки плодов от земли, которую Ты, Господи, дал мне. И поставь это пред Господом Богом твоим, и поклонись пред Господом Богом твоим,
DEUT|26|11|и веселись о всех благах, которые Господь Бог твой дал тебе и дому твоему, ты и левит и пришелец, который будет у тебя.
DEUT|26|12|Когда ты отделишь все десятины произведений [земли] твоей в третий год, год десятин, и отдашь левиту, пришельцу, сироте и вдове, чтоб они ели в жилищах твоих и насыщались,
DEUT|26|13|тогда скажи пред Господом Богом твоим: я отобрал от дома [моего] святыню и отдал ее левиту, пришельцу, сироте и вдове, по всем повелениям Твоим, которые Ты заповедал мне: я не преступил заповедей Твоих и не забыл;
DEUT|26|14|я не ел от нее в печали моей, и не отделял ее в нечистоте, и не давал из нее для мертвого; я повиновался гласу Господа Бога моего, исполнил все, что Ты заповедал мне;
DEUT|26|15|призри от святого жилища Твоего, с небес, и благослови народ Твой, Израиля, и землю, которую Ты дал нам – так как Ты клялся отцам нашим [дать нам] землю, в которой течет молоко и мед.
DEUT|26|16|В день сей Господь Бог твой завещевает тебе исполнять постановления сии и законы: соблюдай и исполняй их от всего сердца твоего и от всей души твоей.
DEUT|26|17|Господу сказал ты ныне, что Он будет твоим Богом, и что ты будешь ходить путями Его и хранить постановления Его и заповеди Его и законы Его, и слушать гласа Его;
DEUT|26|18|и Господь обещал тебе ныне, что ты будешь собственным Его народом, как Он говорил тебе, если ты будешь хранить все заповеди Его,
DEUT|26|19|и что Он поставит тебя выше всех народов, которых Он сотворил, в чести, славе и великолепии, что ты будешь святым народом у Господа Бога твоего, как Он говорил.
DEUT|27|1|И заповедал Моисей и старейшины [сынов] Израилевых народу, говоря: исполняйте все заповеди, которые заповедую вам ныне.
DEUT|27|2|И когда перейдете за Иордан, в землю, которую Господь Бог твой дает тебе, тогда поставь себе большие камни и обмажь их известью;
DEUT|27|3|и напиши на [камнях] сих все слова закона сего, когда перейдешь [Иордан], чтобы вступить в землю, которую Господь Бог твой дает тебе, в землю, где течет молоко и мед, как говорил тебе Господь Бог отцов твоих.
DEUT|27|4|Когда перейдете Иордан, поставьте камни те, как я повелеваю вам сегодня, на горе Гевал, и обмажьте их известью;
DEUT|27|5|и устрой там жертвенник Господу Богу твоему, жертвенник из камней, не поднимая на них железа;
DEUT|27|6|из камней цельных устрой жертвенник Господа Бога твоего, и возноси на нем всесожжения Господу Богу твоему,
DEUT|27|7|и приноси жертвы мирные, и ешь там, и веселись пред Господом Богом твоим;
DEUT|27|8|и напиши на камнях все слова закона сего очень явственно.
DEUT|27|9|И сказал Моисей и священники левиты всему Израилю, говоря: внимай и слушай, Израиль: в день сей ты сделался народом Господа Бога твоего;
DEUT|27|10|итак слушай гласа Господа Бога твоего и исполняй заповеди Его и постановления Его, которые заповедую тебе сегодня.
DEUT|27|11|И заповедал Моисей народу в день тот, говоря:
DEUT|27|12|сии должны стать на горе Гаризим, чтобы благословлять народ, когда перейдете Иордан: Симеон, Левий, Иуда, Иссахар, Иосиф и Вениамин;
DEUT|27|13|а сии должны стать на горе Гевал, чтобы [произносить] проклятие: Рувим, Гад, Асир, Завулон, Дан и Неффалим.
DEUT|27|14|Левиты возгласят и скажут всем Израильтянам громким голосом:
DEUT|27|15|проклят, кто сделает изваянный или литый кумир, мерзость пред Господом, произведение рук художника, и поставит его в тайном месте! Весь народ возгласит и скажет: аминь.
DEUT|27|16|Проклят злословящий отца своего или матерь свою! И весь народ скажет: аминь.
DEUT|27|17|Проклят нарушающий межи ближнего своего! И весь народ скажет: аминь.
DEUT|27|18|Проклят, кто слепого сбивает с пути! И весь народ скажет: аминь.
DEUT|27|19|Проклят, кто превратно судит пришельца, сироту и вдову! И весь народ скажет: аминь.
DEUT|27|20|Проклят, кто ляжет с женою отца своего, ибо он открыл край [одежды] отца своего! И весь народ скажет: аминь.
DEUT|27|21|Проклят, кто ляжет с каким–либо скотом! И весь народ скажет: аминь.
DEUT|27|22|Проклят, кто ляжет с сестрою своею, с дочерью отца своего, или дочерью матери своей! И весь народ скажет: аминь.
DEUT|27|23|Проклят, кто ляжет с тещею своею! И весь народ скажет: аминь.
DEUT|27|24|Проклят, кто тайно убивает ближнего своего! И весь народ скажет: аминь.
DEUT|27|25|Проклят, кто берет подкуп, чтоб убить душу [и пролить] кровь невинную! И весь народ скажет: аминь.
DEUT|27|26|Проклят, кто не исполнит слов закона сего и не будет поступать по ним! И весь народ скажет: аминь.
DEUT|28|1|Если ты, когда перейдете [за Иордан], будешь слушать гласа Господа Бога твоего, тщательно исполнять все заповеди Его, которые заповедую тебе сегодня, то Господь Бог твой поставит тебя выше всех народов земли;
DEUT|28|2|и придут на тебя все благословения сии и исполнятся на тебе, если будешь слушать гласа Господа, Бога твоего.
DEUT|28|3|Благословен ты в городе и благословен на поле.
DEUT|28|4|Благословен плод чрева твоего, и плод земли твоей, и плод скота твоего, и плод твоих волов, и плод овец твоих.
DEUT|28|5|Благословенны житницы твои и кладовые твои.
DEUT|28|6|Благословен ты при входе твоем и благословен ты при выходе твоем.
DEUT|28|7|Поразит пред тобою Господь врагов твоих, восстающих на тебя; одним путем они выступят против тебя, а семью путями побегут от тебя.
DEUT|28|8|Пошлет Господь тебе благословение в житницах твоих и во всяком деле рук твоих; и благословит тебя на земле, которую Господь Бог твой дает тебе.
DEUT|28|9|Поставит тебя Господь народом святым Своим, как Он клялся тебе, если ты будешь соблюдать заповеди Господа Бога твоего и будешь ходить путями Его;
DEUT|28|10|и увидят все народы земли, что имя Господа нарицается на тебе, и убоятся тебя.
DEUT|28|11|И даст тебе Господь изобилие во всех благах, в плоде чрева твоего, и в плоде скота твоего, и в плоде полей твоих на земле, которую Господь клялся отцам твоим дать тебе.
DEUT|28|12|Откроет тебе Господь добрую сокровищницу Свою, небо, чтоб оно давало дождь земле твоей во время свое, и чтобы благословлять все дела рук твоих: и будешь давать взаймы многим народам, а сам не будешь брать взаймы.
DEUT|28|13|Сделает тебя Господь главою, а не хвостом, и будешь только на высоте, а не будешь внизу, если будешь повиноваться заповедям Господа Бога твоего, которые заповедую тебе сегодня хранить и исполнять,
DEUT|28|14|и не отступишь от всех слов, которые заповедую вам сегодня, ни направо ни налево, чтобы пойти вслед иных богов [и] служить им.
DEUT|28|15|Если же не будешь слушать гласа Господа Бога твоего и не будешь стараться исполнять все заповеди Его и постановления Его, которые я заповедую тебе сегодня, то придут на тебя все проклятия сии и постигнут тебя.
DEUT|28|16|Проклят ты [будешь] в городе и проклят ты [будешь] на поле.
DEUT|28|17|Прокляты [будут] житницы твои и кладовые твои.
DEUT|28|18|Проклят [будет] плод чрева твоего и плод земли твоей, плод твоих волов и плод овец твоих.
DEUT|28|19|Проклят ты [будешь] при входе твоем и проклят при выходе твоем.
DEUT|28|20|Пошлет Господь на тебя проклятие, смятение и несчастье во всяком деле рук твоих, какое ни станешь ты делать, доколе не будешь истреблен, – и ты скоро погибнешь за злые дела твои, за то, что ты оставил Меня.
DEUT|28|21|Пошлет Господь на тебя моровую язву, доколе не истребит Он тебя с земли, в которую ты идешь, чтобы владеть ею.
DEUT|28|22|Поразит тебя Господь чахлостью, горячкою, лихорадкою, воспалением, засухою, палящим ветром и ржавчиною, и они будут преследовать тебя, доколе не погибнешь.
DEUT|28|23|И небеса твои, которые над головою твоею, сделаются медью, и земля под тобою железом;
DEUT|28|24|вместо дождя Господь даст земле твоей пыль, и прах с неба будет падать, падать на тебя, доколе не будешь истреблен.
DEUT|28|25|Предаст тебя Господь на поражение врагам твоим; одним путем выступишь против них, а семью путями побежишь от них; и будешь рассеян по всем царствам земли.
DEUT|28|26|И будут трупы твои пищею всем птицам небесным и зверям, и не будет отгоняющего их.
DEUT|28|27|Поразит тебя Господь проказою Египетскою, почечуем, коростою и чесоткою, от которых ты не возможешь исцелиться;
DEUT|28|28|поразит тебя Господь сумасшествием, слепотою и оцепенением сердца.
DEUT|28|29|И ты будешь ощупью ходить в полдень, как слепой ощупью ходит впотьмах, и не будешь иметь успеха в путях твоих, и будут теснить и обижать тебя всякий день, и никто не защитит тебя.
DEUT|28|30|С женою обручишься, и другой будет спать с нею; дом построишь, и не будешь жить в нем; виноградник насадишь, и не будешь пользоваться им.
DEUT|28|31|Вола твоего заколют в глазах твоих, и не будешь есть его; осла твоего уведут от тебя и не возвратят тебе; овцы твои отданы будут врагам твоим, и никто не защитит тебя.
DEUT|28|32|Сыновья твои и дочери твои будут отданы другому народу; глаза твои будут видеть и всякий день истаевать о них, и не будет силы в руках твоих.
DEUT|28|33|Плоды земли твоей и все труды твои будет есть народ, которого ты не знал; и ты будешь только притесняем и мучим во все дни.
DEUT|28|34|И сойдешь с ума от того, что будут видеть глаза твои.
DEUT|28|35|Поразит тебя Господь злою проказою на коленях и голенях, от которой ты не возможешь исцелиться, от подошвы ноги твоей до самого темени [головы] твоей.
DEUT|28|36|Отведет Господь тебя и царя твоего, которого ты поставишь над собою, к народу, которого не знал ни ты, ни отцы твои, и там будешь служить иным богам, деревянным и каменным;
DEUT|28|37|и будешь ужасом, притчею и посмешищем у всех народов, к которым отведет тебя Господь.
DEUT|28|38|Семян много вынесешь в поле, а соберешь мало, потому что поест их саранча.
DEUT|28|39|Виноградники будешь садить и возделывать, а вина не будешь пить, и не соберешь [плодов их], потому что поест их червь.
DEUT|28|40|Маслины будут у тебя во всех пределах твоих, но елеем не помажешься, потому что осыплется маслина твоя.
DEUT|28|41|Сынов и дочерей родишь, но их не будет у тебя, потому что пойдут в плен.
DEUT|28|42|Все дерева твои и плоды земли твоей погубит ржавчина.
DEUT|28|43|Пришелец, который среди тебя, будет возвышаться над тобою выше и выше, а ты опускаться будешь ниже и ниже;
DEUT|28|44|он будет давать тебе взаймы, а ты не будешь давать ему взаймы; он будет главою, а ты будешь хвостом.
DEUT|28|45|И придут на тебя все проклятия сии, и будут преследовать тебя и постигнут тебя, доколе не будешь истреблен, за то, что ты не слушал гласа Господа Бога твоего и не соблюдал заповедей Его и постановлений Его, которые Он заповедал тебе:
DEUT|28|46|они будут знамением и указанием на тебе и на семени твоем вовек.
DEUT|28|47|За то, что ты не служил Господу Богу твоему с веселием и радостью сердца, при изобилии всего,
DEUT|28|48|будешь служить врагу твоему, которого пошлет на тебя Господь, в голоде, и жажде, и наготе и во всяком недостатке; он возложит на шею твою железное ярмо, так что измучит тебя.
DEUT|28|49|Пошлет на тебя Господь народ издалека, от края земли: как орел налетит народ, которого языка ты не разумеешь,
DEUT|28|50|народ наглый, который не уважит старца и не пощадит юноши;
DEUT|28|51|и будет он есть плод скота твоего и плод земли твоей, доколе не разорит тебя, так что не оставит тебе ни хлеба, ни вина, ни елея, ни плода волов твоих, ни плода овец твоих, доколе не погубит тебя;
DEUT|28|52|и будет теснить тебя во всех жилищах твоих, доколе во всей земле твоей не разрушит высоких и крепких стен твоих, на которые ты надеешься; и будет теснить тебя во всех жилищах твоих, во всей земле твоей, которую Господь Бог твой дал тебе.
DEUT|28|53|И ты будешь есть плод чрева твоего, плоть сынов твоих и дочерей твоих, которых Господь Бог твой дал тебе, в осаде и в стеснении, в котором стеснит тебя враг твой.
DEUT|28|54|Муж, изнеженный и живший между вами в великой роскоши, безжалостным оком будет смотреть на брата своего, на жену недра своего и на остальных детей своих, которые останутся у него,
DEUT|28|55|и не даст ни одному из них плоти детей своих, которых он будет есть, потому что у него не останется ничего в осаде и в стеснении, в котором стеснит тебя враг твой во всех жилищах твоих.
DEUT|28|56|[Женщина] жившая у тебя в неге и роскоши, которая никогда ноги своей не ставила на землю по причине роскоши и изнеженности, будет безжалостным оком смотреть на мужа недра своего и на сына своего и на дочь свою
DEUT|28|57|и [не даст] им последа, выходящего из среды ног ее, и детей, которых она родит; потому что она, при недостатке во всем, тайно будет есть их, в осаде и стеснении, в котором стеснит тебя враг твой в жилищах твоих.
DEUT|28|58|Если не будешь стараться исполнять все слова закона сего, написанные в книге сей, и не будешь бояться сего славного и страшного имени Господа Бога твоего,
DEUT|28|59|то Господь поразит тебя и потомство твое необычайными язвами, язвами великими и постоянными, и болезнями злыми и постоянными;
DEUT|28|60|и наведет на тебя все язвы Египетские, которых ты боялся, и они прилипнут к тебе;
DEUT|28|61|и всякую болезнь и всякую язву, не написанную в книге закона сего, Господь наведет на тебя, доколе не будешь истреблен;
DEUT|28|62|и останется вас немного, тогда как множеством вы подобны были звездам небесным, ибо ты не слушал гласа Господа Бога твоего.
DEUT|28|63|И как радовался Господь, делая вам добро и умножая вас, так будет радоваться Господь, погубляя вас и истребляя вас, и извержены будете из земли, в которую ты идешь, чтобы владеть ею.
DEUT|28|64|И рассеет тебя Господь по всем народам, от края земли до края земли, и будешь там служить иным богам, которых не знал ни ты, ни отцы твои, дереву и камням.
DEUT|28|65|Но и между этими народами не успокоишься, и не будет места покоя для ноги твоей, и Господь даст тебе там трепещущее сердце, истаевание очей и изнывание души;
DEUT|28|66|жизнь твоя будет висеть пред тобою, и будешь трепетать ночью и днем, и не будешь уверен в жизни твоей;
DEUT|28|67|от трепета сердца твоего, которым ты будешь объят, и от того, что ты будешь видеть глазами твоими, утром ты скажешь: "о, если бы пришел вечер!", а вечером скажешь: "о, если бы наступило утро!"
DEUT|28|68|и возвратит тебя Господь в Египет на кораблях тем путем, о котором я сказал тебе: "ты более не увидишь его"; и там будете продаваться врагам вашим в рабов и в рабынь, и не будет покупающего.
DEUT|28|69|Вот слова завета, который Господь повелел Моисею поставить с сынами Израилевыми в земле Моавитской, кроме завета, который Господь поставил с ними на Хориве.
DEUT|29|1|И созвал Моисей всех [сынов] Израилевых и сказал им: вы видели все, что сделал Господь пред глазами вашими в земле Египетской с фараоном и всеми рабами его и всею землею его;
DEUT|29|2|те великие казни, которые видели глаза твои, и те великие знамения и чудеса;
DEUT|29|3|но до сего дня не дал вам Господь сердца, чтобы разуметь, очей, чтобы видеть, и ушей, чтобы слышать.
DEUT|29|4|Сорок лет водил вас по пустыне, и одежды ваши на вас не обветшали, и обувь твоя не обветшала на ноге твоей;
DEUT|29|5|хлеба вы не ели и вина и сикера не пили, дабы вы знали, что Я Господь Бог ваш.
DEUT|29|6|И когда пришли вы на место сие, выступил против нас Сигон, царь Есевонский, и Ог, царь Васанский, чтобы сразиться [с нами], и мы поразили их;
DEUT|29|7|и взяли землю их и отдали ее в удел [колену] Рувимову и Гадову и половине колена Манассиина.
DEUT|29|8|Соблюдайте же слова завета сего и исполняйте их, чтобы вам иметь успех во всем, что ни будете делать.
DEUT|29|9|Все вы сегодня стоите пред лицем Господа Бога вашего, начальники колен ваших, старейшины ваши, надзиратели ваши, все Израильтяне,
DEUT|29|10|дети ваши, жены ваши и пришельцы твои, находящиеся в стане твоем, от секущего дрова твои до черпающего воду твою,
DEUT|29|11|чтобы вступить тебе в завет Господа Бога твоего и в клятвенный договор с Ним, который Господь Бог твой сегодня поставляет с тобою,
DEUT|29|12|дабы соделать тебя сегодня Его народом, и Ему быть тебе Богом, как Он говорил тебе и как клялся отцам твоим Аврааму, Исааку и Иакову.
DEUT|29|13|Не с вами только одними я поставляю сей завет и сей клятвенный договор,
DEUT|29|14|но как с теми, которые сегодня здесь с нами стоят пред лицем Господа Бога нашего, так и с теми, которых нет здесь с нами сегодня.
DEUT|29|15|Ибо вы знаете, как мы жили в земле Египетской и как мы проходили посреди народов, чрез которые вы прошли,
DEUT|29|16|и видели мерзости их и кумиры их, деревянные и каменные, серебряные и золотые, которые у них.
DEUT|29|17|Да не будет между вами мужчины или женщины, или рода или колена, которых сердце уклонилось бы ныне от Господа Бога нашего, чтобы ходить служить богам тех народов; да не будет между вами корня, произращающего яд и полынь,
DEUT|29|18|такого человека, который, услышав слова проклятия сего, похвалялся бы в сердце своем, говоря: "я буду счастлив, несмотря на то, что буду ходить по произволу сердца моего"; и пропадет таким образом сытый с голодным;
DEUT|29|19|не простит Господь такому, но тотчас возгорится гнев Господа и ярость Его на такого человека, и падет на него все проклятие [завета сего], написанное в сей книге, и изгладит Господь имя его из поднебесной;
DEUT|29|20|и отделит его Господь на погибель от всех колен Израилевых, сообразно со всеми проклятиями завета, написанными в сей книге закона.
DEUT|29|21|И скажет последующий род, дети ваши, которые будут после вас, и чужеземец, который придет из земли дальней, увидев поражение земли сей и болезни, которыми изнурит ее Господь:
DEUT|29|22|сера и соль, пожарище – вся земля; не засевается и не произращает она, и не выходит на ней никакой травы, как по истреблении Содома, Гоморры, Адмы и Севоима, которые ниспроверг Господь во гневе Своем и в ярости Своей.
DEUT|29|23|И скажут все народы: за что Господь так поступил с сею землею? какая великая ярость гнева Его!
DEUT|29|24|И скажут: за то, что они оставили завет Господа Бога отцов своих, который Он поставил с ними, когда вывел их из земли Египетской,
DEUT|29|25|и пошли и стали служить иным богам и поклоняться им, богам, которых они не знали и [которых] Он не назначал им:
DEUT|29|26|[за то] возгорелся гнев Господа на землю сию, и навел Он на нее все проклятия [завета], написанные в сей книге;
DEUT|29|27|и извергнул их Господь из земли их в гневе, ярости и великом негодовании, и поверг их на другую землю, как ныне [видим].
DEUT|29|28|Сокрытое [принадлежит] Господу Богу нашему, а открытое – нам и сынам нашим до века, чтобы мы исполняли все слова закона сего.
DEUT|30|1|Когда придут на тебя все слова сии – благословение и проклятие, которые изложил я тебе, и примешь [их] к сердцу своему среди всех народов, в которых рассеет тебя Господь Бог твой,
DEUT|30|2|и обратишься к Господу Богу твоему и послушаешь гласа Его, как я заповедую тебе сегодня, ты и сыны твои от всего сердца твоего и от всей души твоей, –
DEUT|30|3|тогда Господь Бог твой возвратит пленных твоих и умилосердится над тобою, и опять соберет тебя от всех народов, между которыми рассеет тебя Господь Бог твой.
DEUT|30|4|Хотя бы ты был рассеян до края неба, и оттуда соберет тебя Господь Бог твой, и оттуда возьмет тебя,
DEUT|30|5|и приведет тебя Господь Бог твой в землю, которою владели отцы твои, и получишь ее во владение, и облагодетельствует тебя и размножит тебя более отцов твоих;
DEUT|30|6|и обрежет Господь Бог твой сердце твое и сердце потомства твоего, чтобы ты любил Господа Бога твоего от всего сердца твоего и от всей души твоей, дабы жить тебе;
DEUT|30|7|тогда Господь Бог твой все проклятия сии обратит на врагов твоих и ненавидящих тебя, которые гнали тебя,
DEUT|30|8|а ты обратишься и будешь слушать гласа Господа и исполнять все заповеди Его, которые заповедую тебе сегодня;
DEUT|30|9|с избытком даст тебе Господь Бог твой успех во всяком деле рук твоих, в плоде чрева твоего, в плоде скота твоего, в плоде земли твоей; ибо снова радоваться будет Господь о тебе, благодетельствуя [тебе], как Он радовался об отцах твоих,
DEUT|30|10|если будешь слушать гласа Господа Бога твоего, соблюдая заповеди Его и постановления Его, написанные в сей книге закона, и если обратишься к Господу Богу твоему всем сердцем твоим и всею душею твоею.
DEUT|30|11|Ибо заповедь сия, которую я заповедую тебе сегодня, не недоступна для тебя и не далека;
DEUT|30|12|она не на небе, чтобы можно [было] говорить: "кто взошел бы для нас на небо и принес бы ее нам, и дал бы нам услышать ее, и мы исполнили бы ее?"
DEUT|30|13|и не за морем она, чтобы можно [было] говорить: "кто сходил бы для нас за море и принес бы ее нам, и дал бы нам услышать ее, и мы исполнили бы ее?"
DEUT|30|14|но весьма близко к тебе слово сие: [оно] в устах твоих и в сердце твоем, чтобы исполнять его.
DEUT|30|15|Вот, я сегодня предложил тебе жизнь и добро, смерть и зло.
DEUT|30|16|[Я] которые заповедую тебе сегодня, любить Господа Бога твоего, ходить по путям Его и исполнять заповеди Его и постановления Его и законы Его, то будешь жить и размножишься, и благословит тебя Господь Бог твой на земле, в которую ты идешь, чтоб овладеть ею;
DEUT|30|17|если же отвратится сердце твое, и не будешь слушать, и заблудишь, и станешь поклоняться иным богам и будешь служить им,
DEUT|30|18|то я возвещаю вам сегодня, что вы погибнете и не пробудете долго на земле, для овладения которою ты переходишь Иордан.
DEUT|30|19|Во свидетели пред вами призываю сегодня небо и землю: жизнь и смерть предложил я тебе, благословение и проклятие. Избери жизнь, дабы жил ты и потомство твое,
DEUT|30|20|любил Господа Бога твоего, слушал глас Его и прилеплялся к Нему; ибо в этом жизнь твоя и долгота дней твоих, чтобы пребывать тебе на земле, которую Господь с клятвою обещал отцам твоим Аврааму, Исааку и Иакову дать им.
DEUT|31|1|И пошел Моисей, и говорил слова сии всем [сынам] Израиля,
DEUT|31|2|и сказал им: теперь мне сто двадцать лет, я не могу уже выходить и входить, и Господь сказал мне: "ты не перейдешь Иордан сей";
DEUT|31|3|Господь Бог твой Сам пойдет пред тобою; Он истребит народы сии от лица твоего, и ты овладеешь ими; Иисус пойдет пред тобою, как говорил Господь;
DEUT|31|4|и поступит Господь с ними так же, как Он поступил с Сигоном и Огом, царями Аморрейскими, и с землею их, которых он истребил;
DEUT|31|5|и предаст их Господь вам, и вы поступите с ними по всем заповедям, какие заповедал я вам;
DEUT|31|6|будьте тверды и мужественны, не бойтесь, и не страшитесь их, ибо Господь Бог твой Сам пойдет с тобою [и] не отступит от тебя и не оставит тебя.
DEUT|31|7|И призвал Моисей Иисуса и пред очами всех Израильтян сказал ему: будь тверд и мужествен, ибо ты войдешь с народом сим в землю, которую Господь клялся отцам его дать ему, и ты разделишь ее на уделы ему;
DEUT|31|8|Господь Сам пойдет пред тобою, Сам будет с тобою, не отступит от тебя и не оставит тебя, не бойся и не ужасайся.
DEUT|31|9|И написал Моисей закон сей, и отдал его священникам, сынам Левииным, носящим ковчег завета Господня, и всем старейшинам [сынов] Израилевых.
DEUT|31|10|И завещал им Моисей и сказал: по прошествии семи лет, в год отпущения, в праздник кущей,
DEUT|31|11|когда весь Израиль придет явиться пред лице Господа Бога твоего на место, которое изберет [Господь], читай сей закон пред всем Израилем вслух его;
DEUT|31|12|собери народ, мужей и жен, и детей, и пришельцев твоих, которые будут в жилищах твоих, чтоб они слушали и учились, и чтобы боялись Господа Бога вашего, и старались исполнять все слова закона сего;
DEUT|31|13|и сыны их, которые не знают [сего], услышат и научатся бояться Господа Бога вашего во все дни, доколе вы будете жить на земле, в которую вы переходите за Иордан, чтоб овладеть ею.
DEUT|31|14|И сказал Господь Моисею: вот, дни твои приблизились к смерти; призови Иисуса и станьте у скинии собрания, и Я дам ему наставления. И пришел Моисей и Иисус, и стали у скинии собрания.
DEUT|31|15|И явился Господь в скинии в столпе облачном, и стал столп облачный у входа скинии.
DEUT|31|16|И сказал Господь Моисею: вот, ты почиешь с отцами твоими, и станет народ сей блудно ходить вслед чужих богов той земли, в которую он вступает, и оставит Меня, и нарушит завет Мой, который Я поставил с ним;
DEUT|31|17|и возгорится гнев Мой на него в тот день, и Я оставлю их и сокрою лице Мое от них, и он истреблен будет, и постигнут его многие бедствия и скорби, и скажет он в тот день: "не потому ли постигли меня сии бедствия, что нет Бога моего среди меня?"
DEUT|31|18|и Я сокрою лице Мое [от него] в тот день за все беззакония его, которые он сделает, обратившись к иным богам.
DEUT|31|19|Итак напишите себе [слова] песни сей, и научи ей сынов Израилевых, и вложи ее в уста их, чтобы песнь сия была Мне свидетельством на сынов Израилевых;
DEUT|31|20|ибо Я введу их в землю, как Я клялся отцам их, где течет молоко и мед, и они будут есть и насыщаться, и утучнеют, и обратятся к иным богам, и будут служить им, а Меня отвергнут и нарушат завет Мой.
DEUT|31|21|и когда постигнут их многие бедствия и скорби, тогда песнь сия будет против них свидетельством, ибо она не выйдет из уст потомства их. Я знаю мысли их, которые они имеют ныне, прежде нежели Я ввел их в землю, о которой Я клялся.
DEUT|31|22|И написал Моисей песнь сию в тот день и научил ей сынов Израилевых.
DEUT|31|23|И заповедал Господь Иисусу, сыну Навину, и сказал [ему]: будь тверд и мужествен, ибо ты введешь сынов Израилевых в землю, о которой Я клялся им, и Я буду с тобою.
DEUT|31|24|Когда Моисей вписал в книгу все слова закона сего до конца,
DEUT|31|25|тогда Моисей повелел левитам, носящим ковчег завета Господня, сказав:
DEUT|31|26|возьмите сию книгу закона и положите ее одесную ковчега завета Господа Бога вашего, и она там будет свидетельством против тебя;
DEUT|31|27|ибо я знаю упорство твое и жестоковыйность твою: вот и теперь, когда я живу с вами ныне, вы упорны пред Господом; не тем ли более по смерти моей?
DEUT|31|28|соберите ко мне всех старейшин колен ваших и надзирателей ваших, и я скажу вслух их слова сии и призову во свидетельство на них небо и землю;
DEUT|31|29|ибо я знаю, что по смерти моей вы развратитесь и уклонитесь от пути, который я завещал вам, и в последствие времени постигнут вас бедствия за то, что вы будете делать зло пред очами Господа, раздражая Его делами рук своих.
DEUT|31|30|И изрек Моисей вслух всего собрания Израильтян слова песни сей до конца:
DEUT|32|1|Внимай, небо, я буду говорить; и слушай, земля, слова уст моих.
DEUT|32|2|Польется как дождь учение мое, как роса речь моя, как мелкий дождь на зелень, как ливень на траву.
DEUT|32|3|Имя Господа прославляю; воздайте славу Богу нашему.
DEUT|32|4|Он твердыня; совершенны дела Его, и все пути Его праведны; Бог верен, и нет неправды [в Нем]; Он праведен и истинен;
DEUT|32|5|но они развратились пред Ним, они не дети Его по своим порокам, род строптивый и развращенный.
DEUT|32|6|Сие ли воздаете вы Господу, народ глупый и несмысленный? не Он ли Отец твой, [Который] усвоил тебя, создал тебя и устроил тебя?
DEUT|32|7|Вспомни дни древние, помысли о летах прежних родов; спроси отца твоего, и он возвестит тебе, старцев твоих, и они скажут тебе.
DEUT|32|8|Когда Всевышний давал уделы народам и расселял сынов человеческих, тогда поставил пределы народов по числу сынов Израилевых;
DEUT|32|9|ибо часть Господа народ Его, Иаков наследственный удел Его.
DEUT|32|10|Он нашел его в пустыне, в степи печальной и дикой, ограждал его, смотрел за ним, хранил его, как зеницу ока Своего;
DEUT|32|11|как орел вызывает гнездо свое, носится над птенцами своими, распростирает крылья свои, берет их и носит их на перьях своих,
DEUT|32|12|так Господь один водил его, и не было с Ним чужого бога.
DEUT|32|13|Он вознес его на высоту земли и кормил произведениями полей, и питал его медом из камня и елеем из твердой скалы,
DEUT|32|14|маслом коровьим и молоком овечьим, и туком агнцев и овнов Васанских и козлов, и тучною пшеницею, и ты пил вино, кровь виноградных ягод.
DEUT|32|15|И утучнел Израиль, и стал упрям; утучнел, отолстел и разжирел; и оставил он Бога, создавшего его, и презрел твердыню спасения своего.
DEUT|32|16|[Богами] чуждыми они раздражили Его и мерзостями разгневали Его:
DEUT|32|17|приносили жертвы бесам, а не Богу, богам, которых они не знали, новым, [которые] пришли от соседей и о которых не помышляли отцы ваши.
DEUT|32|18|А Заступника, родившего тебя, ты забыл, и не помнил Бога, создавшего тебя.
DEUT|32|19|Господь увидел, и в негодовании пренебрег сынов Своих и дочерей Своих,
DEUT|32|20|и сказал: сокрою лице Мое от них [и] увижу, какой будет конец их; ибо они род развращенный; дети, в которых нет верности;
DEUT|32|21|они раздражили Меня не богом, суетными своими огорчили Меня: и Я раздражу их не народом, народом бессмысленным огорчу их;
DEUT|32|22|ибо огонь возгорелся во гневе Моем, жжет до ада преисподнего, и поядает землю и произведения ее, и попаляет основания гор;
DEUT|32|23|соберу на них бедствия и истощу на них стрелы Мои:
DEUT|32|24|[будут] истощены голодом, истреблены горячкою и лютою заразою; и пошлю на них зубы зверей и яд ползающих по земле;
DEUT|32|25|извне будет губить их меч, а в домах ужас – и юношу, и девицу, и грудного младенца, и покрытого сединою старца.
DEUT|32|26|Я сказал бы: рассею их и изглажу из среды людей память о них;
DEUT|32|27|но отложил это ради озлобления врагов, чтобы враги его не возомнили и не сказали: наша рука высока, и не Господь сделал все сие.
DEUT|32|28|Ибо они народ, потерявший рассудок, и нет в них смысла.
DEUT|32|29|О, если бы они рассудили, подумали о сем, уразумели, что с ними будет!
DEUT|32|30|Как бы мог один преследовать тысячу и двое прогонять тьму, если бы Заступник их не предал их, и Господь не отдал их!
DEUT|32|31|Ибо заступник их не таков, как наш Заступник; сами враги наши судьи в том.
DEUT|32|32|Ибо виноград их от виноградной лозы Содомской и с полей Гоморрских; ягоды их ягоды ядовитые, грозды их горькие;
DEUT|32|33|вино их яд драконов и гибельная отрава аспидов.
DEUT|32|34|Не сокрыто ли это у Меня? не запечатано ли в хранилищах Моих?
DEUT|32|35|У Меня отмщение и воздаяние, когда поколеблется нога их; ибо близок день погибели их, скоро наступит уготованное для них.
DEUT|32|36|Но Господь будет судить народ Свой и над рабами Своими умилосердится, когда Он увидит, что рука их ослабела, и не стало ни заключенных, ни оставшихся [вне].
DEUT|32|37|Тогда скажет [Господь]: где боги их, твердыня, на которую они надеялись,
DEUT|32|38|которые ели тук жертв их [и] пили вино возлияний их? пусть они восстанут и помогут вам, пусть будут для вас покровом!
DEUT|32|39|Видите ныне, что это Я, Я – и нет Бога, кроме Меня: Я умерщвляю и оживляю, Я поражаю и Я исцеляю, и никто не избавит от руки Моей.
DEUT|32|40|Я подъемлю к небесам руку Мою и говорю: живу Я во век!
DEUT|32|41|Когда изострю сверкающий меч Мой, и рука Моя приимет суд, то отмщу врагам Моим и ненавидящим Меня воздам;
DEUT|32|42|упою стрелы Мои кровью, и меч Мой насытится плотью, кровью убитых и пленных, головами начальников врага.
DEUT|32|43|Веселитесь, язычники, с народом Его; ибо Он отмстит за кровь рабов Своих, и воздаст мщение врагам Своим, и очистит землю Свою [и] народ Свой!
DEUT|32|44|И пришел Моисей [к народу] и изрек все слова песни сей вслух народа, он и Иисус, сын Навин.
DEUT|32|45|Когда Моисей изрек все слова сии всему Израилю,
DEUT|32|46|тогда сказал им: положите на сердце ваше все слова, которые я объявил вам сегодня, и завещевайте их детям своим, чтобы они старались исполнять все слова закона сего;
DEUT|32|47|ибо это не пустое для вас, но это жизнь ваша, и чрез это вы долгое время пробудете на той земле, в которую вы идете чрез Иордан, чтоб овладеть ею.
DEUT|32|48|И говорил Господь Моисею в тот же самый день и сказал:
DEUT|32|49|взойди на сию гору Аварим, на гору Нево, которая в земле Моавитской, против Иерихона, и посмотри на землю Ханаанскую, которую я даю во владение сынам Израилевым;
DEUT|32|50|и умри на горе, на которую ты взойдешь, и приложись к народу твоему, как умер Аарон, брат твой, на горе Ор, и приложился к народу своему,
DEUT|32|51|за то, что вы согрешили против Меня среди сынов Израилевых при водах Меривы в Кадесе, в пустыне Син, за то, что не явили святости Моей среди сынов Израилевых;
DEUT|32|52|пред [собою] ты увидишь землю, а не войдешь туда, в землю, которую Я даю сынам Израилевым.
DEUT|33|1|Вот благословение, которым Моисей, человек Божий, благословил сынов Израилевых пред смертью своею.
DEUT|33|2|Он сказал: Господь пришел от Синая, открылся им от Сеира, воссиял от горы Фарана и шел со тьмами святых; одесную Его огнь закона.
DEUT|33|3|Истинно Он любит народ [Свой]; все святые его в руке Твоей, и они припали к стопам Твоим, чтобы внимать словам Твоим.
DEUT|33|4|Закон дал нам Моисей, наследие обществу Иакова.
DEUT|33|5|И он был царь Израиля, когда собирались главы народа вместе с коленами Израилевыми.
DEUT|33|6|Да живет Рувим и да не умирает, и да [не] будет малочислен!
DEUT|33|7|Но об Иуде сказал сие: услыши, Господи, глас Иуды и приведи его к народу его; руками своими да защитит он себя, и Ты будь помощником против врагов его.
DEUT|33|8|И о Левии сказал: туммим Твой и урим Твой на святом муже Твоем, которого Ты искусил в Массе, с которым Ты препирался при водах Меривы,
DEUT|33|9|который говорит об отце своем и матери своей: "я на них не смотрю", и братьев своих не признает, и сыновей своих не знает; ибо они, [левиты], слова Твои хранят и завет Твой соблюдают,
DEUT|33|10|учат законам Твоим Иакова и заповедям Твоим Израиля, возлагают курение пред лице Твое и всесожжения на жертвенник Твой;
DEUT|33|11|благослови, Господи, силу его и о деле рук его благоволи, порази чресла восстающих на него и ненавидящих его, чтобы они не могли стоять.
DEUT|33|12|О Вениамине сказал: возлюбленный Господом обитает у Него безопасно, [Бог] покровительствует ему всякий день, и он покоится между раменами Его.
DEUT|33|13|Об Иосифе сказал: да благословит Господь землю его вожделенными дарами неба, росою и [дарами] бездны, лежащей внизу,
DEUT|33|14|вожделенными плодами от солнца и вожделенными произведениями луны,
DEUT|33|15|превосходнейшими произведениями гор древних и вожделенными дарами холмов вечных,
DEUT|33|16|и вожделенными дарами земли и того, что наполняет ее; благословение Явившегося в терновом кусте да приидет на главу Иосифа и на темя наилучшего из братьев своих;
DEUT|33|17|крепость его как первородного тельца, и роги его, как роги буйвола; ими избодет он народы все до пределов земли: это тьмы Ефремовы, это тысячи Манассиины.
DEUT|33|18|О Завулоне сказал: веселись, Завулон, в путях твоих, и Иссахар, в шатрах твоих;
DEUT|33|19|созывают они народ на гору, там заколают законные жертвы, ибо они питаются богатством моря и сокровищами, сокрытыми в песке.
DEUT|33|20|О Гаде сказал: благословен распространивший Гада; он покоится как лев и сокрушает и мышцу и голову;
DEUT|33|21|он избрал себе начаток [земли], там почтен уделом от законодателя, и пришел с главами народа, и исполнил правду Господа и суды с Израилем.
DEUT|33|22|О Дане сказал: Дан молодой лев, который выбегает из Васана.
DEUT|33|23|О Неффалиме сказал: Неффалим насыщен благоволением и исполнен благословения Господа; море и юг во владении [его].
DEUT|33|24|Об Асире сказал: благословен между сынами Асир, он будет любим братьями своими, и окунет в елей ногу свою;
DEUT|33|25|железо и медь – запоры твои; как дни твои, [будет умножаться] богатство твое.
DEUT|33|26|Нет подобного Богу Израилеву, Который по небесам принесся на помощь тебе и во славе Своей на облаках;
DEUT|33|27|прибежище [твое] Бог древний, и [ты] под мышцами вечными; Он прогонит врагов от лица твоего и скажет: истребляй!
DEUT|33|28|Израиль живет безопасно, один; око Иакова [видит пред] [собою] землю обильную хлебом и вином, и небеса его каплют росу.
DEUT|33|29|Блажен ты, Израиль! кто подобен тебе, народ, хранимый Господом, Который есть щит, охраняющий тебя, и меч славы твоей? Враги твои раболепствуют тебе, и ты попираешь выи их.
DEUT|34|1|И взошел Моисей с равнин Моавитских на гору Нево, на вершину Фасги, что против Иерихона, и показал ему Господь всю землю Галаад до самого Дана,
DEUT|34|2|и всю [землю] Неффалимову, и [всю] землю Ефремову и Манассиину, и всю землю Иудину, даже до самого западного моря,
DEUT|34|3|и полуденную страну и равнину долины Иерихона, город Пальм, до Сигора.
DEUT|34|4|И сказал ему Господь: вот земля, о которой Я клялся Аврааму, Исааку и Иакову, говоря: "семени твоему дам ее"; Я дал тебе увидеть ее глазами твоими, но в нее ты не войдешь.
DEUT|34|5|И умер там Моисей, раб Господень, в земле Моавитской, по слову Господню;
DEUT|34|6|и погребен на долине в земле Моавитской против Беф–Фегора, и никто не знает [места] погребения его даже до сего дня.
DEUT|34|7|Моисею было сто двадцать лет, когда он умер; но зрение его не притупилось, и крепость в нем не истощилась.
DEUT|34|8|И оплакивали Моисея сыны Израилевы на равнинах Моавитских тридцать дней. И прошли дни плача и сетования о Моисее.
DEUT|34|9|И Иисус, сын Навин, исполнился духа премудрости, потому что Моисей возложил на него руки свои, и повиновались ему сыны Израилевы и делали так, как повелел Господь Моисею.
DEUT|34|10|И не было более у Израиля пророка такого, как Моисей, которого Господь знал лицем к лицу,
DEUT|34|11|по всем знамениям и чудесам, которые послал его Господь сделать в земле Египетской над фараоном и над всеми рабами его и над всею землею его,
DEUT|34|12|и по руке сильной и по великим чудесам, которые Моисей совершил пред глазами всего Израиля.
