EXOD|1|1|А оце ймення Ізраїлевих синів, що прийшли з Яковом до Єгипту. Кожен із домом своїм прибули:
EXOD|1|2|Рувим, Симеон, Левій і Юда,
EXOD|1|3|Іссахар, Завулон і Веніямин,
EXOD|1|4|Дан і Нефталим, Ґад і Асир.
EXOD|1|5|І було всіх душ, що вийшли з стегна Якового, сімдесят душ. А Йосип був ув Єгипті.
EXOD|1|6|І вмер Йосип і всі браття його, та ввесь той рід.
EXOD|1|7|А Ізраїлеві сини плодилися сильно, і розмножувались, та й стали вони надзвичайно сильні. І наповнився ними той край.
EXOD|1|8|І став над Єгиптом новий цар, що не знав Йосипа.
EXOD|1|9|І сказав він до народу свого: Ось народ Ізраїлевих синів численніший і сильніший від нас!
EXOD|1|10|Станьмо ж мудріші за нього, щоб він не множився! Бо буде, коли нам трапиться війна, то прилучиться й він до ворогів наших, і буде воювати проти нас, і вийде з цього краю.
EXOD|1|11|І настановили над ним начальників податків, щоб його гнобити своїми тягарами. І він будував міста на запаси фараонові: Пітом і Рамесес.
EXOD|1|12|Але що більше його гнобили, то більше він множився та більше ширився. І жахалися єгиптяни через Ізраїлевих синів.
EXOD|1|13|І Єгипет змушував синів Ізраїля тяжко працювати.
EXOD|1|14|І вони огірчували їхнє життя тяжкою працею коло глини та коло цегли, і коло всякої праці на полі, кожну їхню працю, яку змушували тяжко робити.
EXOD|1|15|І звелів був єгипетський цар єврейським бабам-сповитухам, що одній ім'я Шіфра, а ім'я другій Пуа,
EXOD|1|16|і говорив: Як будете бабувати єврейок, то дивіться на порід: коли буде син, то вбийте його, а коли це дочка, то нехай живе.
EXOD|1|17|Але баби-сповитухи боялися Бога, і не робили того, як казав їм єгипетський цар. І вони лишали хлопчиків при житті.
EXOD|1|18|І покликав єгипетський цар баб-сповитух, та й сказав їм: Нащо ви робите цю річ, та лишаєте дітей при житті?
EXOD|1|19|І сказали баби-сповитухи до фараона: Бо єврейки не такі, як єгипетські жінки, бо вони самі баби-сповитухи: поки прийде до них баба-сповитуха, то вони вже й народять.
EXOD|1|20|І Бог чинив добро бабам-сповитухам, а народ розмножувався, і сильно міцнів.
EXOD|1|21|І сталося, тому, що ті баби-сповитухи боялися Бога, то Він будував їм доми.
EXOD|1|22|І наказав фараон усьому народові своєму, говорячи: Кожного народженого єврейського сина кидайте його до Річки, а кожну дочку зоставляйте при житті!
EXOD|2|1|І пішов один муж з дому Левія, і взяв собі за жінку дочку Левієву.
EXOD|2|2|І завагітніла та жінка, та й сина вродила. І побачили його, що він гарний, та й ховала його три місяці.
EXOD|2|3|Та не могла його більше ховати. І взяла йому папірусову скриньку, і виасфальтувала її асфальтом та смолою, і положила до неї дитину, та й поклала в очереті на березі Річки.
EXOD|2|4|А сестра його стояла здалека, щоб довідатися, що йому станеться.
EXOD|2|5|І зійшла фараонова дочка купатися на Річку, а служниці її ходили понад Річкою. І побачила вона ту скриньку серед очерету, і послала невільницю свою, щоб узяла її.
EXOD|2|6|І відчинила, та й побачила дитину, ось хлопчик плаче. І вона змилосердилася над ним, та й сказала: Це з єврейських дітей!
EXOD|2|7|І сказала сестра його до фараонової дочки: Чи не піти й не покликати тобі жінку-мамку з єврейок, і вона годуватиме тобі дитину?
EXOD|2|8|І сказала їй дочка фараонова: Іди. І пішла та дівчина, і покликала матір дитини.
EXOD|2|9|А дочка фараонова сказала до неї: На тобі цю дитину, та й годуй її для мене. А я дам тобі заплату. І взяла та жінка дитину, і годувала її.
EXOD|2|10|І підросло те дитя, і вона привела його до фараонової дочки, і він став їй за сина. І вона назвала йому ймення Мойсей, і сказала: бо з води я витягла його.
EXOD|2|11|І сталося за тих днів, і підріс Мойсей. І вийшов він до братів своїх, та й приглядався до їхніх терпінь. І побачив він єгиптянина, що бив єврея з братів його.
EXOD|2|12|І озирнувся він туди та сюди, і побачив, що нікого нема, та й убив єгиптянина, і заховав його в пісок.
EXOD|2|13|І вийшов він другого дня, аж ось сваряться двоє євреїв. І сказав він несправедливому: Нащо ти б'єш свого ближнього?
EXOD|2|14|А той відказав: Хто тебе настановив за начальника та за суддю над нами? Чи ти думаєш убити мене, як ти вбив був єгиптянина? І злякався Мойсей та й сказав собі: Справді, та справа стала відома!
EXOD|2|15|І почув фараон про цю справу, та й шукав, щоб убити Мойсея. І втік Мойсей від фараонового лиця, і оселився в країні Мідіян.
EXOD|2|16|А в мідіянського жерця було сім дочок. І прийшли вони, і витягали воду, і наповнили корита, щоб напоїти отару свого батька.
EXOD|2|17|І прийшли пастухи й відігнали їх. І встав Мойсей, та й оборонив їх, і напоїв їхню отару.
EXOD|2|18|І прибули вони до Реуїла, свого батька, а той поспитав: Чого ви сьогодні так скоро прийшли?.
EXOD|2|19|А ті відказали: Якийсь єгиптянин оборонив нас від руки пастухів, а також навіть натягав нам води й напоїв отару.
EXOD|2|20|І сказав він до своїх дочок: А де він? Чому ви покинули того чоловіка? Покличте його, і нехай він з'їсть хліба.
EXOD|2|21|І погодився Мойсей сидіти з тим чоловіком, а той видав за Мойсея дочку свою Ціппору.
EXOD|2|22|І породила вона сина, а він назвав ім'я йому: Ґершом, бо сказав: Я став приходьком у чужому краї.
EXOD|2|23|І сталося по довгих днях, і вмер цар Єгипту. А Ізраїлеві сини стогнали від тієї роботи та кричали. І їхній зойк через ту роботу донісся до Бога.
EXOD|2|24|І почув Бог їхній стогін. І згадав Бог Свого заповіта з Авраамом, Ісаком та Яковом.
EXOD|2|25|І Бог бачив синів Ізраїлевих, і Бог зглянувся над ними.
EXOD|3|1|А Мойсей пас отару тестя свого Їтра, жерця Мідіянського. І провадив він цю отару за пустиню, і прийшов був до Божої гори, до Хориву.
EXOD|3|2|І явився йому Ангол Господній у полум'ї огняному з-посеред тернового куща. І побачив він, що та тернина горить огнем, але не згорає кущ.
EXOD|3|3|І сказав Мойсей: Зійду но, і побачу це велике видіння, чому не згорає та тернина?
EXOD|3|4|І побачив Господь, що він зійшов подивитися. І кликнув до нього Бог з-посеред тієї тернини і сказав: Мойсею, Мойсею! А той відказав: Ось я!
EXOD|3|5|І сказав Він: Не зближайся сюди! Здійми взуття своє з ніг своїх, бо те місце, на якому стоїш ти, земля це свята!
EXOD|3|6|І сказав: Я Бог батька твого, Бог Авраама, Бог Ісака й Бог Якова! І сховав Мойсей обличчя своє, бо боявся споглянуть на Бога!
EXOD|3|7|І промовив Господь: Я справді бачив біду Свого народу, що в Єгипті, і почув його зойк перед його гнобителями, бо пізнав Я болі його.
EXOD|3|8|І Я зійшов, щоб визволити його з єгипетської руки, та щоб вивести його з цього краю до Краю доброго й широкого, до Краю, що тече молоком та медом до місця ханаанеянина, і хіттеянина, і амореянина, і періззеянина, і хіввеянина, і євусеянина.
EXOD|3|9|А тепер ось зойк Ізраїлевих синів дійшов до Мене, і Я також побачив той утиск, що ним єгиптяни їх тиснуть.
EXOD|3|10|А тепер іди ж, і Я пошлю тебе до фараона, і виведи з Єгипту народ Мій, синів Ізраїлевих!
EXOD|3|11|І сказав Мойсей до Бога: Хто я, що піду до фараона, і що виведу з Єгипту синів Ізраїлевих?
EXOD|3|12|А Він відказав: Та Я буду з тобою! А це тобі знак, що Я послав тебе: коли ти виведеш народ із Єгипту, то ви будете служити Богові на оцій горі.
EXOD|3|13|І сказав Мойсей до Бога: Ото я прийду до Ізраїлевих синів та й скажу їм: Бог ваших батьків послав мене до вас, то вони запитають мене: Яке Ім'я Його? Що я скажу їм?
EXOD|3|14|І сказав Бог Мойсеєві: Я Той, що є. І сказав: Отак скажеш Ізраїлевим синам: Сущий послав мене до вас.
EXOD|3|15|І сказав іще Бог до Мойсея: Отак скажи Ізраїлевим синам: Господь, Бог батьків ваших, Бог Авраама, Бог Ісака й Бог Якова послав мене до вас. А оце Ім'я Моє навіки, і це пам'ять про Мене з роду в рід.
EXOD|3|16|Іди, збери старших Ізраїлевих та й скажи їм: Господь, Бог батьків ваших, явився мені, Бог Авраама, Ісака та Якова, говорячи: Згадуючи, згадав Я про вас, та про заподіяне вам ув Єгипті.
EXOD|3|17|І сказав Я: Я виведу вас з єгипетської біди до Краю ханаанеянина, і хіттеянина, й амореянина, і періззеянина, і хіввеянина, і євусеянина, до Краю, що тече молоком та медом.
EXOD|3|18|І вони послухають слова твого, і прийдеш ти та старші Ізраїлеві до єгипетського царя, та й скажете йому: Господь, Бог євреїв, стрівся був нам. А тепер ми підемо в триденну дорогу в пустиню, і складемо жертви Господеві, Богові нашому!
EXOD|3|19|І Я знаю, що єгипетський цар не дасть вам піти, як не буде змушений рукою сильною.
EXOD|3|20|І Я витягну Свою руку, та й поб'ю Єгипет усіма чудами Моїми, що вчиню серед нього, а потому він відпустить вас.
EXOD|3|21|І Я дам милість цьому народові в очах Єгипту, і станеться, коли підете, не підете ви впорожні!
EXOD|3|22|Бо позичить жінка від сусідки своєї і від мешканки дому свого посуд срібний і посуд золотий та одежу, і покладете це на синів ваших та на дочок ваших, і заберете здобич від Єгипту.
EXOD|4|1|І відповів Мойсей та й сказав: Таж вони не повірять мені, і не послухають голосу мого, бо скажуть: Господь не явився тобі!
EXOD|4|2|І промовив до нього Господь: Що то в руці твоїй? Той відказав: Палиця.
EXOD|4|3|І сказав Він: Кинь її на землю! І той кинув її на землю, і вона стала вужем. І втік Мойсей від нього.
EXOD|4|4|І сказав Господь до Мойсея: Простягни свою руку, і візьми його за хвоста! І він простяг свою руку й узяв його, і той став палицею в долоні його.
EXOD|4|5|Щоб повірили, що явився тобі Господь, Бог їхніх батьків, Бог Авраама, Бог Ісака й Бог Якова.
EXOD|4|6|І сказав Господь йому ще: Засунь свою руку за пахвину свою! І засунув він руку свою за пахвину свою, і витягнув її, аж ось рука його побіліла від прокази, як сніг!
EXOD|4|7|А Він сказав: Поклади знов свою руку за пахвину свою! І він поклав знову руку свою до своєї пахвини, і витягнув її з пахвини своєї, і ось вона стала знову, як тіло його.
EXOD|4|8|І станеться, коли не повірять тобі, і не послухають голосу першої ознаки, то повірять голосу ознаки наступної.
EXOD|4|9|І станеться коли вони не повірять також обом тим ознакам, і не послухають твого голосу, то ти візьмеш води з Річки, і виллєш на суходіл. І переміниться та вода, що ти візьмеш із Річки, і станеться кров'ю на суходолі.
EXOD|4|10|Та Мойсей сказав до Господа: О Господи я не промовець ні від учора, ні від позавчора, ані відтоді, коли Ти говорив був до Свойого раба, бо я тяжкоустий та тяжкоязикий.
EXOD|4|11|І сказав йому Господь: Хто дав уста людині? Або Хто робить німим, чи глухим, чи видючим, чи темним, чи ж не Я, Господь?
EXOD|4|12|А тепер іди, а Я буду з устами твоїми, і буду навчати тебе, що ти маєш говорити.
EXOD|4|13|А він відказав: Молю Тебе, Господи, пошли іншого, кого маєш послати.
EXOD|4|14|І запалав гнів Господній на Мойсея, і Він сказав: Чи ж не Аарон твій брат, Левит? Я знаю, що він добре буде говорити. Та ось він вийде навпроти тебе, і побачить тебе, і зрадіє він у серці своїм.
EXOD|4|15|І ти будеш говорити до нього, і вкладеш слова ці в уста його, а Я буду з устами твоїми й з устами його, і буду навчати вас, що маєте робити.
EXOD|4|16|І він буде говорити за тебе до народу. І станеться, він буде тобі устами, а ти будеш йому замість Бога.
EXOD|4|17|І ти візьмеш у руку свою оцю палицю, якою ознаки чинитимеш.
EXOD|4|18|І пішов Мойсей, і вернувся до тестя свого Їтра, і сказав йому: Піду я, і вернуся до братів своїх, що в Єгипті, і побачу, чи ще живі вони. А Їтро сказав до Мойсея: Іди в мирі!
EXOD|4|19|І сказав Господь до Мойсея в Мідіяні: Іди, вернися до Єгипту, бо вимерли всі люди, що шукали твоєї душі.
EXOD|4|20|І взяв Мойсей жінку свою та синів своїх, і посадив їх на осла, та й вернувся до єгипетського краю. І взяв Мойсей палицю Божу в руку свою.
EXOD|4|21|І сказав Господь до Мойсея: Коли ти підеш, щоб вернутися до Єгипту, гляди, щоб усі чуда, які Я вклав у твою руку, ти вчинив їх перед лицем фараона, а Я ожорсточу серце його, і він не відпустить народу.
EXOD|4|22|І ти скажеш фараонові: Так сказав Господь: Син Мій, Мій перворідний то Ізраїль.
EXOD|4|23|І кажу Я тобі: Відпусти Мого сина, і нехай Мені служить. А коли ти відмовиш пустити його, то ось Я вб'ю твого сина, твого перворідного.
EXOD|4|24|І сталося в дорозі на нічлігу, стрів був його Господь і шукав, щоб убити його.
EXOD|4|25|Та Ціппора взяла кременя, і обрізала крайню плоть свого сина, і доторкнулася нею до ніг його та й сказала: Бо ти мені наречений крови!
EXOD|4|26|І пустив Він його. Тоді вона сказала: Наречений крови через обрізання.
EXOD|4|27|І сказав Господь до Аарона: Іди назустріч Мойсею в пустиню! І він пішов, і стрів його на горі Божій, і поцілував його.
EXOD|4|28|І розповів Мойсей Ааронові всі слова Господа, що послав його, і всі ті ознаки, що Він наказав був йому.
EXOD|4|29|І пішов був Мойсей та Аарон, і зібрали вони всіх старших Ізраїлевих синів.
EXOD|4|30|І переказав Аарон усі слова, що Господь говорив був Мойсеєві. А той ті ознаки чинив на очах народу.
EXOD|4|31|І повірив народ той. І почули вони, що згадав Господь Ізраїлевих синів, і що побачив біду їх, і вони схилилися, і поклонилися до землі.
EXOD|5|1|А потім прийшли Мойсей й Аарон, та й сказали до фараона: Так сказав Господь, Бог Ізраїлів: Відпусти народ Мій, і нехай вони святкують Мені на пустині!
EXOD|5|2|А фараон відказав: Хто Господь, що послухаюсь слова Його, щоб відпустити Ізраїля? Не знаю Господа, і також Ізраїля не відпущу!
EXOD|5|3|І сказали вони: Бог євреїв стрівся з нами. Нехай же ми підемо триденною дорогою на пустиню, і принесемо жертви Господеві, Богові нашому, щоб не доторкнувся Він до нас мором або мечем.
EXOD|5|4|І сказав до них цар Єгипту: Чому ви, Мойсею та Аароне, відриваєте народ від його робіт? Ідіть до своїх діл!
EXOD|5|5|І сказав фараон: Таж багато тепер цього простолюду, а ви здержуєте їх від їхніх робіт.
EXOD|5|6|І того дня фараон наказав погоничам народу та писарям, говорячи:
EXOD|5|7|Не давайте більше народові соломи, щоб робити цеглу, як учора й позавчора. Нехай ідуть самі, та збирають собі соломи.
EXOD|5|8|А призначене число цегли, що вони робили вчора й позавчора, накладете на них, не зменшуйте з нього. Вони нероби, тому кричать: Ходім, принесімо жертву нашому Богові!
EXOD|5|9|Нехай буде тяжка праця на цих людей, і нехай працюють на ній, і нехай покинуть облудні слова.
EXOD|5|10|І вийшли погоничі народу й писарі його, та й сказали до того народу, говорячи: Так сказав фараон: Я не буду давати вам соломи.
EXOD|5|11|Самі йдіть, наберіть собі соломи, де знайдете, бо нічого не зменшене з вашої роботи!.
EXOD|5|12|І розпорошився народ той по всій єгипетській землі, щоб збирати стерню на солому.
EXOD|5|13|А погоничі наставали, говорячи: Скінчіть вашу щоденну працю в час так, як коли б була солома.
EXOD|5|14|І були биті писарі синів Ізраїлевих, що їх настановили над ними фараонові погоничі, говорячи: Чому ви не скінчили свого приділу для виробу цегли й учора й сьогодні, як було дотепер?
EXOD|5|15|І прибули писарі Ізраїлевих синів, та й кричали до фараона, говорячи: Для чого ти так робиш рабам своїм?
EXOD|5|16|Соломи не дають твоїм рабам, а цеглу кажуть нам робіть! І ось раби твої биті, і грішиш ти перед народом своїм!
EXOD|5|17|А він відказав: Нероби ви, нероби! Тому ви говорите: Ходім, принесімо жертву Господеві.
EXOD|5|18|А тепер ідіть, працюйте, а соломи не дадуть вам! Але призначене число цегли ви дасте!
EXOD|5|19|І бачили Ізраїлеві писарі себе в біді, коли говорено: Не зменшуйте з цегли вашої щоденного в його часі!
EXOD|5|20|І стріли вони Мойсея та Аарона, що стояли насупроти них, як вони виходили від фараона,
EXOD|5|21|та й сказали до них: Нехай побачить вас Господь і нехай вас осудить, бо ви вчинили ненависним дух наш в очах фараона й в очах його рабів, щоб дати меча в їхню руку повбивати нас!
EXOD|5|22|І вернувся Мойсей до Господа та й сказав: Господи, чому Ти кривду вчинив цьому народові? Чому Ти послав мені це?
EXOD|5|23|Бо відколи прийшов я до фараона, щоб говорити Твоїм Ім'ям, він ще більшу кривду чинить цьому народові, а насправді Ти не визволив народу Свого!
EXOD|6|1|І сказав Господь до Мойсея: Тепер побачиш, що вчиню Я фараонові, бо він, змушений рукою сильною, їх відпустить, і, змушений рукою сильною, вижене їх із краю свого.
EXOD|6|2|І говорив Бог до Мойсея, та й сказав йому: Я Господь!
EXOD|6|3|І являвся Я Авраамові, Ісакові та Яковові Богом Всемогутнім, але Йменням Своїм Господь Я не дався їм пізнати.
EXOD|6|4|А також Я склав був із ними Свого заповіта, що дам їм землю ханаанську, землю їх мандрування, в якій вони мандрували.
EXOD|6|5|І почув Я теж стогін синів Ізраїлевих, що єгиптяни роблять їх своїми рабами, і згадав заповіта Свого.
EXOD|6|6|Тому скажи синам Ізраїлевим: Я Господь! І Я виведу вас з-під тягарів Єгипту, і визволю вас від їхньої роботи, і звільню вас витягненим раменом та великими присудами.
EXOD|6|7|І візьму вас Собі за народа, і буду вам Богом, і ви познаєте, що Я Господь, Бог ваш, що виводить вас із-під тягарів Єгипту!
EXOD|6|8|І введу вас до того Краю, що про нього Я підняв був Свою руку, щоб дати його Авраамові, Ісакові та Якову. І Я дам його вам на спадщину. Я Господь!
EXOD|6|9|І так говорив Мойсей до синів Ізраїлевих, та вони не слухали Мойсея через легкодухість та тяжку роботу.
EXOD|6|10|І казав Господь до Мойсея, говорячи:
EXOD|6|11|Увійди, говори до фараона, царя єгипетського, і нехай він відпустить Ізраїлевих синів із свого краю.
EXOD|6|12|І казав Мойсей перед лицем Господнім, говорячи: Таж Ізраїлеві сини не слухали мене, як же послухає мене фараон? А я необрізановустий!
EXOD|6|13|І казав Господь до Мойсея та до Аарона, і дав їм накази до Ізраїлевих синів та до фараона, царя єгипетського, щоб вивести Ізраїлевих синів з єгипетського краю.
EXOD|6|14|Оце голови батьківських домів їхніх. Сини Рувима, перворідного Ізраїлевого: Ханох і Паллу, Хецрон і Кармі, це родини Рувимові.
EXOD|6|15|А сини Симеонові: Ємуїл, і Ямін, і Огад, і Яхін, і Цохар, і Шаул, син ханаанеянки, це родини Симеонові.
EXOD|6|16|А оце імена синів Левієвих за їхніми родинами: Ґершон, і Кегат, і Мерарі. А літа життя Левієвого сто і тридцять і сім літ.
EXOD|6|17|Сини Ґершонові: Лівні, і Шім'ї за їхніми родинами.
EXOD|6|18|А сини Кегатові: Амрам, і Їцгар, і Хеврон, і Уззіїл. А літа життя Кегатового сто і тридцять і три роки.
EXOD|6|19|А сини Мерарі: Махлі та Муші. Оце родини Левієві за їхніми родами.
EXOD|6|20|І взяв Амрам свою тітку Йохевед собі за жінку, і вона породила йому Аарона та Мойсея. А літа життя Амрамового сто і тридцять і сім літ.
EXOD|6|21|А сини Їцгарові: Корах, і Нефеґ, і Зіхрі.
EXOD|6|22|А сини Уззіїлові: Мішаїл, і Елцафан, і Сітрі.
EXOD|6|23|І взяв Аарон Елішеву, дочку Амінадавову, сестру Нахшонову, собі за жінку, і вона породила йому Надава, і Авігу, і Елеазара, і Ітамара.
EXOD|6|24|А сини Корахові: Ассир, і Елкана, і Аваасаф, це родини Корахові.
EXOD|6|25|А Елеазар, син Ааронів, узяв собі з дочок Путіїлових за жінку, і вона породила йому Пінхаса. Оце голови батьківських домів Левітів за їхніми родинами.
EXOD|6|26|Оце Аарон і Мойсей, що Господь говорив їм: Виведіть Ізраїлевих синів з єгипетського краю за їхніми військовими відділами.
EXOD|6|27|Вони ті, що говорили до фараона, царя єгипетського, щоб вивести Ізраїлевих синів з Єгипту, це Мойсей та Аарон.
EXOD|6|28|І сталося в дні, коли Господь говорив до Мойсея в єгипетськім краї,
EXOD|6|29|то казав Господь до Мойсея, говорячи: Я Господь! Говори фараонові, цареві єгипетському, усе, що Я говорю тобі.
EXOD|6|30|І сказав Мойсей перед обличчям Господнім: Таж я необрізановустий! Як же слухати буде мене фараон?
EXOD|7|1|І сказав Господь до Мойсея: Дивись, Я поставив тебе замість Бога для фараона, а твій брат Аарон буде пророк твій.
EXOD|7|2|Ти будеш говорити все, що Я накажу тобі, а брат твій Аарон буде говорити фараонові, і нехай він відпустить Ізраїлевих синів з свого краю.
EXOD|7|3|А Я вчиню запеклим фараонове серце, і помножу ознаки мої та чуда мої в єгипетськім краї.
EXOD|7|4|І не послухає вас фараон, а Я покладу Свою руку на Єгипет, і виведу війська Свої, народ Мій, синів Ізраїлевих, з єгипетського краю великими присудами.
EXOD|7|5|І пізнають єгиптяни, що Я Господь, коли простягну Свою руку на Єгипет і виведу від них Ізраїлевих синів.
EXOD|7|6|І вчинив Мойсей та Аарон, як звелів їм Господь, так учинили вони.
EXOD|7|7|А Мойсей був віку восьмидесяти літ, а Аарон восьмидесяти і трьох літ, коли вони говорили до фараона.
EXOD|7|8|І промовив Господь до Мойсея й до Аарона, говорячи:
EXOD|7|9|Коли буде до вас говорити фараон, кажучи: Покажіть своє чудо, то скажеш Ааронові: Візьми свою палицю, та й кинь перед лицем фараоновим, нехай станеться вужем!
EXOD|7|10|І ввійшов Мойсей та Аарон до фараона, та й вчинили так, як наказав був Господь. І кинув Аарон палицю свою перед лицем фараона й перед його рабами, і вона стала вужем!
EXOD|7|11|І покликав фараон також мудреців та ворожбитів, і вчинили так само й вони, чарівники єгипетські, своїми чарами.
EXOD|7|12|І кинули кожен палицю свою, і вони поставали вужами. Та Ааронова палиця проковтнула палиці їхні.
EXOD|7|13|Та затверділо фараонове серце, і він не послухався їх, як говорив був Господь.
EXOD|7|14|І сказав Господь до Мойсея: Запекле фараонове серце, він відмовив відпустити народ!
EXOD|7|15|Піди до фараона рано вранці. Ось він вийде до води, а ти стань навпроти нього на березі Річки. А палицю, що була змінена на вужа, візьмеш у свою руку.
EXOD|7|16|І скажеш йому: Господь, Бог євреїв, послав мене до тебе, кажучи: Відпусти Мій народ, і нехай вони служать Мені на пустині! Та не послухався ти дотепер.
EXOD|7|17|Так сказав Господь: По цьому пізнаєш, що Я Господь: Ось я вдарю палицею, що в руці моїй, по воді, що в Річці, і вона зміниться на кров!
EXOD|7|18|А риба, що в Річці, погине. І засмердиться Річка, і попомучаться єгиптяни, щоб пити воду з Річки!
EXOD|7|19|І сказав Господь до Мойсея: Скажи Ааронові: Візьми свою палицю, і простягни свою руку над водою єгиптян, над їхніми річками, над їхніми потоками, і над ставами їхніми, і над кожним водозбором їхнім, і вони стануть кров'ю. І буде кров по всій єгипетській землі, і в посуді дерев'янім, і в каміннім.
EXOD|7|20|І Мойсей та Аарон зробили так, як наказав був Господь. І підняв він палицю, та й ударив воду, що в Річці, на очах фараона й на очах його рабів. І змінилася вся вода, що в Річці, на кров!
EXOD|7|21|А риби, що в Річці, погинули. І засмерділася Річка, і не могли єгиптяни пити воду з Річки. І була кров у всім єгипетськім краї.
EXOD|7|22|І так само зробили єгипетські чарівники своїми чарами. І стало запеклим фараонове серце, і він не послухався їх, як говорив був Господь.
EXOD|7|23|І повернувся фараон, і ввійшов до дому свого, і не приклав він свого серця також до цього.
EXOD|7|24|І всі єгиптяни копали біля Річки, щоб дістати води до пиття, бо не могли пити води з Річки.
EXOD|7|25|І минуло сім день по тому, як Господь ударив Річку.
EXOD|8|1|(7-26) І промовив Господь до Мойсея: Іди до фараона, та й скажи йому: Так сказав Господь: Відпусти Мій народ, і нехай вони служать Мені.
EXOD|8|2|(7-27) А коли ти відмовишся відпустити, то ось Я вдарю ввесь край твій жабами.
EXOD|8|3|(7-28) І стане Річка роїти жаби, і вони повиходять, і ввійдуть до твого дому, і до спальної кімнати твоєї, і на ліжко твоє, і до домів рабів твоїх, і до народу твого, і до печей твоїх, і до діжок твоїх.
EXOD|8|4|(7-29) І на тебе, і на народ твій, і на всіх рабів твоїх повилазять ці жаби.
EXOD|8|5|(8-1) І сказав Господь до Мойсея: Скажи Ааронові: Простягни свою руку з палицею своєю на річки, на потоки, і на ставки, і повиводь жаб на єгипетський край.
EXOD|8|6|(8-2) І простяг Аарон руку свою на єгипетські води, і вийшла жабня, та й покрила єгипетську землю.
EXOD|8|7|(8-3) Та так само зробили й єгипетські чарівники своїми чарами, і вивели жаб на єгипетську землю.
EXOD|8|8|(8-4) І покликав фараон Мойсея й Аарона, та й сказав: Благайте Господа, і нехай виведе ці жаби від мене й від народу мого, а я відпущу народ той, і нехай приносять жертви для Господа!
EXOD|8|9|(8-5) І сказав Мойсей фараонові: Накажи мені, коли маю молитися за тебе, і за слуг твоїх, і за народ твій, щоб понищити жаби від тебе й від домів твоїх, тільки в Річці вони позостануться.
EXOD|8|10|(8-6) А той відказав: На завтра. І сказав Мойсей: За словом твоїм! Щоб ти знав, що нема Такого, як Господь, Бог наш!
EXOD|8|11|(8-7) І відійдуть жаби від тебе, і від домів твоїх, і він рабів твоїх, і від народу твого, тільки в Річці вони позостануться.
EXOD|8|12|(8-8) І вийшов Мойсей та Аарон від фараона. І кликав Мойсей до Господа про ті жаби, що навів був на фараона.
EXOD|8|13|(8-9) І зробив Господь за словом Мойсея, і погинули жаби з домів, і з подвір'їв, і з піль.
EXOD|8|14|(8-10) І збирали їх цілими купами, і засмерділась земля!
EXOD|8|15|(8-11) І побачив фараон, що сталась полегша, і знову стало запеклим серце його, і не послухався їх, як говорив був Господь.
EXOD|8|16|(8-12) І сказав Господь до Мойсея: Скажи Ааронові: Простягни свою палицю, та й удар земний порох, і нехай він стане вошами в усьому єгипетському краї!
EXOD|8|17|(8-13) І зробили вони так. І простяг Аарон руку свою з палицею своєю, та й ударив земний порох, і він стався вошами на людині й на скотині. Увесь земний порох стався вошами в усьому єгипетському краї.
EXOD|8|18|(8-14) І так само робили чарівники своїми чарами, щоб навести воші, та не змогли. І була вошва на людині й на скотині.
EXOD|8|19|(8-15) І сказали чарівники фараонові: Це перст Божий! Та серце фараонове було запеклим, і він не послухався їх, як говорив був Господь.
EXOD|8|20|(8-16) І сказав Господь до Мойсея: Устань рано вранці, та й стань перед лицем фараоновим. Ось він піде до води, а ти скажи йому: Так сказав Господь: Відпусти Мій народ, і нехай вони служать Мені!
EXOD|8|21|(8-17) Бо коли ти не відпустиш народу Мого, то ось Я пошлю на тебе, і на слуг твоїх, і на народ твій, і на доми твої рої мух. І єгипетські доми будуть повні мушні, а також земля, на якій вони живуть.
EXOD|8|22|(8-18) І відділю того дня землю Ґошен, що Мій народ живе на ній, щоб не було там роїв мух, щоб ти знав, що Я Господь посеред землі!
EXOD|8|23|(8-19) І зроблю Я різницю між народом Моїм та народом твоїм. Узавтра буде це знамено!
EXOD|8|24|(8-20) І зробив Господь так. І найшла численна мушня на дім фараона, і на дім рабів його, і на всю єгипетську землю. І нищилась земля через ті рої мух!
EXOD|8|25|(8-21) І кликнув фараон до Мойсея та до Аарона, говорячи: Підіть, принесіть жертви вашому Богові в цьому краї!
EXOD|8|26|(8-22) А Мойсей відказав: Не годиться чинити так, бо то огиду для Єгипту ми приносили б у жертву Господу, Богові нашому. Тож будемо приносити в жертву огиду для єгиптян на їхніх очах, і вони не вкаменують нас?
EXOD|8|27|(8-23) Триденною дорогою ми підемо на пустиню, і принесемо жертву Господеві, Богові нашому, як скаже Він нам.
EXOD|8|28|(8-24) І сказав фараон: Я відпущу вас, і ви принесете жертву Господеві, Богові вашому на пустині. Тільки далеко не віддаляйтесь, ідучи. Моліться за мене!
EXOD|8|29|(8-25) І сказав Мойсей: Ось я виходжу від тебе, і буду благати Господа, і відступить той рій мух від фараона, і від рабів його, і від народу його взавтра. Тільки нехай більше не обманює фараон, щоб не відпустити народу принести жертву Господеві.
EXOD|8|30|(8-26) І вийшов Мойсей від фараона, і став просити Господа.
EXOD|8|31|(8-27) І зробив Господь за словом Мойсея, і відвернув рої мух від фараона, від рабів його, і від народу його. І не зосталося ані однієї.
EXOD|8|32|(8-28) А фараон зробив запеклим своє серце також і цим разом, і не відпустив він народу того!
EXOD|9|1|І сказав Господь до Мойсея: Увійди до фараона, і говори до нього: Так сказав Господь, Бог євреїв: Відпусти Мій народ, і нехай вони служать Мені!
EXOD|9|2|Бо коли ти відмовишся відпустити, і будеш держати їх ще,
EXOD|9|3|то ось Господня рука буде на худобі твоїй, що на полі, на конях, на ослах, на верблюдах, на худобі великій і дрібній, моровиця дуже тяжка.
EXOD|9|4|І відділить Господь між худобою Ізраїля й між худобою Єгипту, і не загине нічого зо всього, що належить Ізраїлевим синам.
EXOD|9|5|І призначив Господь усталений час, кажучи: Узавтра Господь зробить цю річ у цім краї.
EXOD|9|6|І зробив Господь ту річ назавтра, і вигинула вся єгипетська худоба, а з худоби Ізраїлевих синів не згинуло ані одне.
EXOD|9|7|І послав фараон довідатись, а ось не згинуло з худоби Ізраїлевої ані одне! І стало фараонове серце запеклим, і не відпустив він народу того!
EXOD|9|8|І сказав Господь до Мойсея й до Аарона: Візьміть собі повні ваші жмені сажі з печі, і нехай Мойсей кине її до неба на очах фараонових.
EXOD|9|9|І стане вона курявою над усією єгипетською землею, а на людині й скотині стане гнояками, що кинуться прищами в усьому єгипетському краї.
EXOD|9|10|І набрали вони сажі з печі, та й стали перед фараоновим лицем. І кинув її Мойсей до неба, і стали прищуваті гнояки, що кинулися на людині й на скотині.
EXOD|9|11|А чарівники не могли стати перед Мойсеєм через гнояки, бо гнояк той був на чарівниках і на всіх єгиптянах.
EXOD|9|12|І вчинив запеклим Господь фараонове серце, і він не послухався їх, як говорив був Господь до Мойсея.
EXOD|9|13|І сказав Господь до Мойсея: Устань рано вранці, і стань перед лицем фараоновим та й скажи йому: Отак сказав Господь, Бог євреїв: Відпусти Мій народ, і нехай вони служать Мені!
EXOD|9|14|Бо цим разом Я пошлю всі урази Мої на серце твоє, і на рабів твоїх, і на народ твій, щоб ти знав, що немає на всій землі Такого, як Я!
EXOD|9|15|Бо тепер, коли б Я простягнув Свою руку, то побив би тебе та народ твій мором, і ти був би вигублений із землі.
EXOD|9|16|Але Я для того залишив тебе, щоб показати тобі Мою силу, і щоб оповідали про Ймення Моє по всій землі.
EXOD|9|17|Ти ще опираєшся проти народу Мого, щоб їх не відпустити.
EXOD|9|18|Ось Я взавтра, цього саме часу, зішлю дощем тяженний град, що такого, як він, не бувало в Єгипті від дня його заложення аж до сьогодні.
EXOD|9|19|А тепер пошли, позаганяй худобу свою та все, що твоє в полі. Кожна людина й худоба, що буде застукана в полі, і не буде забрана додому, то зійде на них град, і вони повмирають!
EXOD|9|20|Хто з фараонових рабів боявся Господнього слова, той зігнав своїх рабів та свою худобу до домів.
EXOD|9|21|А хто не звернув свого серця до слова Господнього, той позалишав рабів своїх та худобу свою на полі.
EXOD|9|22|І сказав Господь до Мойсея: Простягни свою руку до неба, і нехай буде град у всьому єгипетському краї на людину, і на худобу, і на всю польову траву в єгипетській землі!
EXOD|9|23|І простяг Мойсей палицю свою до неба, і Господь дав громи та град. І зійшов на землю огонь, і Господь дощив градом на єгипетську землю.
EXOD|9|24|І був град, і огонь горів посеред тяженного граду, що не бувало такого, як він, у всім єгипетськім краї, відколи він став був народом.
EXOD|9|25|І повибивав той град у всім єгипетськім краї все, що на полі, від людини аж до худоби! І всю польову рослинність побив той град, а кожне польове дерево поламав!
EXOD|9|26|Тільки в землі Ґошен, де жили Ізраїлеві сини, не було граду.
EXOD|9|27|І послав фараон, і покликав Мойсея та Аарона, та й сказав до них: Згрішив я тим разом! Господь справедливий, а я та народ мій несправедливі!
EXOD|9|28|Благайте Господа, і досить бути Божим громам та градові! А я відпущу вас, і ви більше не залишитеся...
EXOD|9|29|І сказав до нього Мойсей: Як вийду я з міста, то простягну руки свої до Господа, громи перестануть, а граду вже не буде, щоб ти знав, що Господня ця земля!
EXOD|9|30|А ти й раби твої, знаю я, що ви ще не боїтеся перед лицем Господа Бога!
EXOD|9|31|А льон та ячмінь був побитий, бо ячмінь дозрівав, а льон цвів.
EXOD|9|32|А пшениця та жито не були вибиті, бо пізні вони.
EXOD|9|33|І вийшов Мойсей від фараона з міста, і простяг руки свої до Господа, і перестали громи та град, а дощ не лив на землю.
EXOD|9|34|І побачив фараон, що перестав дощ, і град та громи, та й далі грішив. І чинив він запеклим своє серце, він та раби його.
EXOD|9|35|І стало запеклим фараонове серце, і він не відпустив Ізраїлевих синів, як говорив був Господь через Мойсея.
EXOD|10|1|І сказав Господь до Мойсея: Увійди до фараона, бо Я зробив запеклим серце його та серце рабів його, щоб показати ці ознаки Мої серед нього,
EXOD|10|2|і щоб ти розповідав в уші сина свого та онука свого, що зробив Я в Єгипті, та про ознаки Мої, що вчинив я серед них. І ви будете знати, що Я Господь!
EXOD|10|3|І ввійшли Мойсей та Аарон до фараона, та й сказали йому: Так сказав Господь, Бог євреїв: Аж доки ти будеш відмовлятися впокоритися передо Мною? Відпусти Мій народ, і нехай вони служать Мені!
EXOD|10|4|Бо коли ти відмовишся відпустити народ Мій, то ось Я взавтра спроваджу сарану на твій край.
EXOD|10|5|І покриє вона поверхню землі, і не можна буде бачити землі. І поїсть вона решту вцілілого, позосталого вам від граду, і поїсть вона кожне дерево, що росте вам з землі.
EXOD|10|6|І переповняться нею доми ваші, і доми всіх рабів ваших, і доми всього Єгипту, чого не бачили батьки ваші та батьки батьків твоїх від дня існування їх на землі аж до сьогодні! І він відвернувся, і вийшов від фараона.
EXOD|10|7|І сказали раби фараона до нього: Аж доки цей буде нам пасткою? Відпусти цих людей, і нехай вони служать Господеві, Богові своєму. Чи ти ще не знаєш, що знищений Єгипет?
EXOD|10|8|І повернено Мойсея та Аарона до фараона, а він їм сказав: Ідіть, служіть Господеві, Богові вашому. Хто та хто піде?
EXOD|10|9|І відповів Мойсей: Ми підемо з молоддю нашою та з старими нашими, з синами нашими та з дочками нашими, з дрібною нашою худобою та з великою нашою худобою підемо, бо в нас свято Господнє.
EXOD|10|10|А він відказав: Нехай буде так Господь із вами, як я відпущу вас і дітей ваших!... Та глядіть, бо щось лихе перед вами.
EXOD|10|11|Тож нехай ідуть самі чоловіки, та й служіть Господеві, бо того ви бажаєте. І вигнано їх від лиця фараонового.
EXOD|10|12|І сказав Господь до Мойсея: Простягни свою руку на єгипетську землю сараною, і нехай вона найде на єгипетський край, і нехай поїсть усю земну траву, усе, що град позалишав.
EXOD|10|13|І простяг Мойсей свою палицю на єгипетську землю, і Господь навів східній вітер на землю, цілий день той і цілу ніч. Настав ранок, і східній вітер наніс сарани!
EXOD|10|14|І найшла сарана на всю єгипетську землю, і залягла в усім єгипетськім краї, дуже багато! Перед нею не було такої сарани, як вона, і по ній не буде такої!
EXOD|10|15|І покрила вона поверхню всієї землі, і потемніла земля! І поїла вона всю земну траву та ввесь плід дерева, що град позоставив. І не зосталось ніякої зелені ані на дереві, ані на польовій рослинності в усім єгипетськім краї!
EXOD|10|16|І поспішив фараон покликати Мойсея та Аарона, та й сказав: Згрішив я Господеві, Богові вашому, та вам!
EXOD|10|17|А тепер пробач же мій гріх тільки цього разу, і помоліться до Господа, вашого Бога, і нехай тільки відверне від мене цю смерть!
EXOD|10|18|І він вийшов від фараона й молився до Господа.
EXOD|10|19|І повернув Господь західній дуже сильний вітер назад, і він поніс сарану, та й укинув її до Червоного моря. Не позосталась жодна сарана в усім єгипетськім краї.
EXOD|10|20|Та Господь учинив запеклим фараонове серце, і він знов не відпустив Ізраїлевих синів.
EXOD|10|21|І сказав Господь до Мойсея: Простягни свою руку до Неба, і станеться темрява на єгипетській землі, і нехай буде темрява, щоб відчули її.
EXOD|10|22|І простяг Мойсей свою руку до неба, і сталася густа темрява по всій єгипетській землі три дні.
EXOD|10|23|Не бачили один одного, і ніхто не вставав з свого місця три дні! А Ізраїлевим синам було світло в їхніх садибах.
EXOD|10|24|І покликав фараон Мойсея, та й сказав: Ідіть, служіть Господеві! Тільки дрібна ваша худоба та ваша худоба велика нехай позостанеться. Також дітвора ваша нехай іде з вами!
EXOD|10|25|Та Мойсей відказав: Дай в наші руки також жертви та цілопалення, і ми спорядимо жертву Господеві, Богові нашому.
EXOD|10|26|І також худоба наша піде з нами, не зостанеться ані копита, бо з нього ми візьмемо на служення Господеві, Богові нашому. Бо ми не знаємо, поки прибудемо туди, чим будемо служити Господеві.
EXOD|10|27|І вчинив запеклим Господь фараонове серце, і він не хотів відпустити їх.
EXOD|10|28|І сказав йому фараон: Іди від мене! Стережися, щоб ти не бачив більше лиця мого, бо того дня, коли побачиш лице моє, ти помреш!
EXOD|10|29|А Мойсей відказав: Так сказав ти... Я більш уже не побачу лиця твого!
EXOD|11|1|І сказав Господь до Мойсея: Ще одну поразу наведу Я на фараона й на Єгипет. Потому він відпустить вас ізвідси. А коли він буде відпускати вас, то зовсім вас вижене звідси!
EXOD|11|2|Скажи ж у вуха народу, і нехай позичить кожен від свого ближнього, а кожна від своєї ближньої посуд срібний та посуд золотий,
EXOD|11|3|І дав Господь милість тому народові в очах Єгипту. Також і цей муж, Мойсей, був дуже великий в єгипетськім краї в очах фараонових рабів та в очах того народу.
EXOD|11|4|І промовив Мойсей: Так сказав Господь! Коло півночі Я вийду посеред Єгипту.
EXOD|11|5|І помре кожен перворідний єгипетської землі від перворідного фараона, що сидить на своїм престолі, до перворідного невільниці, що за жорнами, і все перворідне з худоби.
EXOD|11|6|І здійметься великий зойк по всій єгипетській землі, що такого, як він, не бувало, і такого, як він, більш не буде.
EXOD|11|7|А в усіх синів Ізраїлевих від людини й аж до худоби навіть пес не висуне язика свого, щоб ви знали, що відділює Господь між Єгиптом і між Ізраїлем.
EXOD|11|8|І зійдуть усі оці раби твої до мене, і поклоняться мені, кажучи: Вийди ти та ввесь народ, що слухає тебе. По цьому я вийду. І він вийшов від фараона, розпалений гнівом.
EXOD|11|9|І сказав Господь до Мойсея: Не послухав вас фараон, щоб могли помножитись чуда Мої в єгипетськім краї.
EXOD|11|10|А Мойсей та Аарон учинили всі оці чуда перед лицем фараоновим. Та зробив запеклим Господь фараонове серце, і він не відпустив Ізраїлевих синів із своєї землі.
EXOD|12|1|І сказав Господь до Мойсея й до Аарона в єгипетськім краї, говорячи:
EXOD|12|2|Оцей місяць для вас початок місяців. Він вам перший між місяцями року.
EXOD|12|3|Скажіть усій ізраїльській громаді, говорячи: У десятий день цього місяця нехай візьмуть собі кожен ягня за домом батьків, ягня на дім.
EXOD|12|4|А коли буде той дім замалий, щоб з'їсти ягня, то нехай візьме він і найближчий до його дому сусід його за числом душ. Кожен згідно з їдою своєю полічиться на те ягня.
EXOD|12|5|Ягня у вас нехай буде без вади, самець, однорічне. Візьміть його з овечок та з кіз.
EXOD|12|6|І нехай буде воно для вас пильноване аж до чотирнадцятого дня цього місяця. І заколе його цілий збір Ізраїлевої громади на смерканні.
EXOD|12|7|І нехай візьмуть тієї крови, і нехай покроплять на обидва бокові одвірки, і на одвірок верхній у тих домах, що будуть їсти його в них.
EXOD|12|8|І нехай їдять тієї ночі те м'ясо, спечене на огні, та опрісноки. Нехай їдять його на гірких травах.
EXOD|12|9|Не їжте з нього сирового та вареного, звареного в воді, бо до їди тільки спечене на огні, голова його з голінками його та з нутром його.
EXOD|12|10|І не лишайте з нього нічого до ранку, а полишене з нього до ранку спаліть на огні.
EXOD|12|11|А їсти його будете так: стегна ваші підперезані, взуття ваше на ногах ваших, а палиця ваша в руці вашій, і будете ви їсти його в поспіху. Пасха це для Господа!
EXOD|12|12|І перейду Я тієї ночі в єгипетськім краї, і повбиваю в єгипетській землі кожного перворідного від людини аж до скотини. А над усіма єгипетськими богами вчиню Я суд. Я Господь!
EXOD|12|13|І буде та кров вам знаком на тих домах, що там ви, і побачу ту кров, і обмину вас. І не буде між вами згубної порази, коли Я вбиватиму в єгипетськім краї.
EXOD|12|14|І стане той день для вас пам'яткою, і будете святкувати його, як свято для Господа на всі роди ваші! Як постанову вічну будете святкувати його!
EXOD|12|15|Сім днів будете їсти опрісноки. Але першого дня зробите, щоб не було квашеного в ваших домах, бо кожен, хто їстиме квашене, від дня першого аж до дня сьомого, то буде витята душа та з Ізраїля.
EXOD|12|16|А першого дня будуть у вас священні збори, і сьомого дня священні збори. Жодна праця не буде робитися в них, тільки що їсти кожній душі, те єдине робитимете ви.
EXOD|12|17|І ви будете додержувати опрісноків, бо саме того дня Я вивів війська ваші з єгипетського краю. І будете додержувати того дня в ваших родах, як постанови вічної.
EXOD|12|18|Першого місяця, чотирнадцятого дня місяця будете їсти опрісноки аж до вечора дня двадцять першого того ж місяця.
EXOD|12|19|Сім день квашене не буде знаходитися в ваших домах, бо кожен, хто їстиме квашене, то буде витята душа та з Ізраїльської громади, чи то серед приходьків, чи то тих, хто народився у краї.
EXOD|12|20|Жодного квашеного не будете їсти в усіх ваших оселях, будете їсти опрісноки!
EXOD|12|21|І покликав Мойсей усіх старших Ізраїлевих, та й промовив до них: Спровадьте й візьміть собі дрібну худобину за родинами вашими, і заколіть пасху.
EXOD|12|22|І візьміть в'язку ісопу й умочіть у кров, що в посудині, і доторкніться горішнього одвірка й двох одвірків бічних кров'ю, що в посудині. А ви, ніхто не вийдете з дверей дому свого аж до ранку!
EXOD|12|23|І перейде Господь ударити Єгипет, і побачить ту кров на одвірку горішнім і на двох одвірках бічних, і обмине Господь ті двері, і не дасть згубникові ввійти до ваших домів, щоб ударити.
EXOD|12|24|А ви будете дотримувати цю річ, як постанови для себе й для синів своїх аж навіки.
EXOD|12|25|І станеться, коли ви ввійдете до того Краю, що дасть вам Господь, як Він обіцяв був, то ви будете додержувати цієї служби.
EXOD|12|26|І станеться коли запитають вас ваші сини: Що то за служба ваша?
EXOD|12|27|то відкажете: Це жертва Пасха для Господа, що обминув був доми Ізраїлевих синів в Єгипті, коли побивав Єгипет, а доми наші зберіг. І схилився народ, і вклонивсь до землі.
EXOD|12|28|І пішли й учинили сини Ізраїля, як наказав був Господь Мойсеєві та Ааронові, так учинили вони.
EXOD|12|29|І сталося в половині ночі, і вдарив Господь в єгипетськім краї кожного перворідного, від перворідного фараона, що сидить на своїм престолі, аж до перворідного полоненого, що у в'язничному домі, і кожного перворідного худоби.
EXOD|12|30|І встав фараон уночі, він та всі раби його, та ввесь Єгипет. І знявся великий зойк в Єгипті, бо не було дому, щоб не було там померлого!...
EXOD|12|31|І покликав фараон Мойсея та Аарона вночі, та й сказав: Устаньте, вийдіть з-посеред народу мого, і ви, і сини Ізраїлеві. І йдіть, служіть Господеві, як ви казали!
EXOD|12|32|І дрібну вашу худобу, і худобу вашу велику візьміть, як ви казали, та й ідіть. І поблагословіть і мене!
EXOD|12|33|І квапили єгиптяни народ той, щоб спішно відпустити їх із краю, бо казали: Усі ми помремо!
EXOD|12|34|І поніс той народ тісто своє, поки воно вкисло, діжки свої, зав'язані в їхні одежі, на плечах своїх.
EXOD|12|35|І Ізраїлеві сини вчинили за словом Мойсеєвим, і позичили від єгиптян посуд срібний і посуд золотий та шати.
EXOD|12|36|А Господь дав милість тому народові в очах Єгипту, і вони позичили і забрали здобич від Єгипту.
EXOD|12|37|І вирушили Ізраїлеві сини з Рамесесу до Суккоту, близько шости сот тисяч чоловіка піхоти, крім дітей,
EXOD|12|38|а також багато різного люду піднялися з ними, і дрібна худоба й велика худоба, маєток дуже великий.
EXOD|12|39|І пекли вони те тісто, що винесли з Єгипту, на прісні коржі, бо не вкисло воно, бо вони були вигнані з Єгипту, і не могли баритися, а поживи на дорогу не приготовили собі.
EXOD|12|40|А перебування Ізраїлевих синів, що сиділи в Єгипті, чотириста років і тридцять років.
EXOD|12|41|І сталося в кінці чотирьохсот років і тридцяти років, і сталося саме того дня, вийшли всі Господні війська з єгипетського краю.
EXOD|12|42|Це ніч сторожі для Господа, бо Він вивів їх з єгипетського краю. Ця сама ніч сторожа для Господа всім синам Ізраїля на їхні покоління.
EXOD|12|43|І сказав Господь до Мойсея й до Аарона: Це постанова про Пасху: жоден чужинець не буде їсти її.
EXOD|12|44|А кожен раб людський куплений за срібло, коли обріжеш його, тоді він буде їсти її.
EXOD|12|45|Приходько та наймит не буде їсти її.
EXOD|12|46|В самому домі буде вона їстися, не винесеш із дому назовні того м'яса, а костей його не зламаєте.
EXOD|12|47|Уся громада Ізраїлева буде справляти її.
EXOD|12|48|А коли буде мешкати з тобою приходько, і схоче справляти Пасху Господеві, то нехай буде обрізаний в нього кожен чоловічої статі, а тоді він приступить справляти її, і він буде, як народжений в Краї. А кожен необрізаний не буде їсти її.
EXOD|12|49|Один закон буде для тубільця й для приходька, що мешкає серед вас.
EXOD|12|50|І вчинили всі Ізраїлеві сини, як наказав був Господь Мойсеєві та Ааронові, так учинили вони.
EXOD|12|51|І сталося того саме дня, вивів Господь Ізраїлевих синів з єгипетського краю за їхніми відділами.
EXOD|13|1|І Господь промовляв до Мойсея, говорячи:
EXOD|13|2|Посвяти Мені кожного перворідного, що розкриває всяку утробу серед Ізраїлевих синів, серед людини й серед худоби, для Мене воно!
EXOD|13|3|І сказав Мойсей до народу: Пам'ятайте той день, коли ви вийшли з Єгипту, із дому рабства! Бо силою руки Господь вивів вас ізвідти; і не будете їсти квашеного.
EXOD|13|4|Ви виходите сьогодні, у місяці авіві.
EXOD|13|5|І станеться, коли Господь уведе тебе до краю ханаанеянина, і хіттеянина, й амореянина, і хіввеянина, й євусеянина, що про нього присягнув був батькам твоїм, щоб дати тобі Край, який тече молоком та медом, то ти будеш служити ту службу того місяця.
EXOD|13|6|Сім день будеш їсти опрісноки, а дня сьомого свято для Господа!
EXOD|13|7|Опрісноки будуть їстися сім тих день, і не побачиться в тебе квашене, і не побачиться в тебе квашене в усім Краї твоїм!
EXOD|13|8|І оповіси синові своєму того дня, говорячи: Це для того, що вчинив мені Господь, коли я виходив із Єгипту.
EXOD|13|9|І буде тобі це за знака на руці твоїй, і за пам'ятку між очима твоїми, щоб Господній Закон був в устах твоїх, бо сильною рукою Господь вивів тебе із Єгипту.
EXOD|13|10|І будеш додержуватися цієї постанови в означенім часі її з року в рік.
EXOD|13|11|І станеться, коли введе тебе Господь до землі ханаанеянина, як присяг був тобі та батькам твоїм, і дасть її тобі,
EXOD|13|12|то відділиш усе, що розкриває утробу, для Господа, і все перворідне худоби, що буде в тебе, самці для Господа!
EXOD|13|13|А кожного віслюка, що розкриває утробу, викупиш овечкою; а коли не викупиш, то зламай йому шию. І кожного перворідного людського серед синів твоїх викупиш.
EXOD|13|14|І станеться, коли взавтра запитає тебе син твій, говорячи: Що то? то відповіси йому: Силою Своєї руки вивів нас Господь із Єгипту, із дому рабства.
EXOD|13|15|І сталося, коли фараон учинив запеклим своє серце, щоб не відпустити нас, то Господь повбивав усіх перворідних в єгипетськім краї, від перворідного людського й аж до перворідного худоби. Тому то я приношу в жертву Господеві все чоловічої статі, що розкриває утробу, а кожного перворідного синів своїх викупляю.
EXOD|13|16|І станеться це за знака на руці твоїй, і за пов'язку поміж очима твоїми, бо силою Своєї руки вивів нас Господь із Єгипту.
EXOD|13|17|І сталося, коли фараон відпустив був той народ, то Бог не повів їх дорогою землі филистимської, хоч була близька вона. Бо Бог сказав: Щоб не пожалкував той народ, коли він побачить війну, і не вернувся до Єгипту.
EXOD|13|18|І повів Бог той народ окружною дорогою пустині аж до Червоного моря. І вийшли Ізраїлеві сини з єгипетського краю узброєні.
EXOD|13|19|А Мойсей забрав із собою кості Йосипа, бо присягою той закляв був Ізраїлевих синів, кажучи: Напевно згадає Бог вас, і ви винесете з собою кості мої звідси.
EXOD|13|20|І вони рушили з Суккоту, і розтаборилися в Етам, на границі пустині.
EXOD|13|21|А Господь ішов перед ними вдень у стовпі хмари, щоб провадити їх дорогою, а вночі в стовпі огню, щоб світити їм, щоб ішли вдень та вночі.
EXOD|13|22|Не відступав удень стовп хмари тієї, а вночі стовп огню з-перед обличчя народу!
EXOD|14|1|І говорив Господь до Мойсея, кажучи:
EXOD|14|2|Скажи Ізраїлевим синам, і нехай вони повернуть, і нехай отаборяться перед Пі-Гахіротом, між Міґдолом і між морем, перед Баал-Цефоном. Навпроти нього отаборитесь над морем.
EXOD|14|3|І скаже фараон про Ізраїлевих синів: заблудились вони в землі цій, замкнено пустиню для них.
EXOD|14|4|І вчиню запеклим фараонове серце, і він буде гнатися за вами, а Я прославлюся через фараона та через військо його. І пізнають єгиптяни, що Я Господь! І вони вчинили так.
EXOD|14|5|І повідомлено царя єгипетського, що втік той народ. І змінилося серце фараона та рабів його до того народу, і сказали вони: Що це ми зробили, що відпустили Ізраїля від роботи нам?
EXOD|14|6|І запріг він свою колесницю, і забрав народ свій з собою.
EXOD|14|7|І взяв він шість сотень добірних колесниць, і всі колесниці Єгипту, і трійкових над усіма ними.
EXOD|14|8|І Господь учинив запеклим серце фараона, єгипетського царя, і він погнався за Ізраїлевими синами. Але Ізраїлеві сини виходили сильною рукою!
EXOD|14|9|І гналися єгиптяни за ними, уся кіннота, колесниці фараонові, і комонники його та військо його, і догнали їх, як вони отаборилися були над морем, під Пі-Гахіротом, перед Баал-Цефоном.
EXOD|14|10|А фараон наближався. І звели Ізраїлеві сини свої очі, аж ось єгиптяни женуться за ними! І дуже злякались вони... І кликали Ізраїлеві сини до Господа,
EXOD|14|11|а Мойсеєві дорікали: Чи через те, що не було гробів в Єгипті, ти забрав нас умирати в пустині? Що це вчинив ти нам, щоб вивести нас із Єгипту?
EXOD|14|12|Чи це не те саме ми говорили до тебе в Єгипті, кажучи: Позостав нас, і нехай ми робимо Єгиптові! Бо ліпше нам рабство Єгиптові, аніж помирати нам у пустині!
EXOD|14|13|І сказав Мойсей до народу: Не бійтеся! Стійте, і побачите спасіння Господа, що вчинить вам сьогодні. Бо єгиптян, яких бачите сьогодні, більше не побачите їх уже повіки!
EXOD|14|14|Господь буде воювати за вас, а ви мовчіть!
EXOD|14|15|І промовив Господь до Мойсея: Що ти до Мене кличеш? Говори до синів Ізраїлевих, нехай рушають!
EXOD|14|16|А ти підійми свою палицю, і простягни руку свою на море, і розітни його, і нехай увійдуть Ізраїлеві сини в середину моря, на суходіл.
EXOD|14|17|А Я, ось Я вчиню запеклим серце єгиптянам, і вони ввійдуть за ними. І буду Я прославлений через фараона, і через усе його військо, і через колесниці, його, і через комонників його.
EXOD|14|18|І пізнають єгиптяни, що Я Господь, коли буду Я прославлений через фараона, і через колесниці його, і через комонників його!
EXOD|14|19|І рушив Ангол Божий, що йшов перед Ізраїльським табором, і пішов за ними; і рушив стовп хмари перед ними, і став за ними,
EXOD|14|20|і ввійшов він у середину між табір Єгипту й між табір Ізраїлів. І була та хмара і темрява для Єгипту, а ніч розсвітлив він для Ізраїля. І не зближався один до одного цілу ніч.
EXOD|14|21|І простяг Мойсей руку свою на море, і Господь гнав море сильним східнім вітром цілу ніч, і зробив море суходолом, і розступилася вода.
EXOD|14|22|І ввійшли Ізраїлеві сини в середину моря, як на суходіл, а море було для них муром із правиці їхньої та з лівиці їхньої.
EXOD|14|23|А єгиптяни гналися, і ввійшли за ними всі фараонові коні й колесниці його, та його комонники до середини моря.
EXOD|14|24|І сталося за ранньої сторожі, і поглянув Господь на єгипетський табір у стовпі огня й хмари, та й привів у замішання єгипетський табір.
EXOD|14|25|І поскидав колеса з колесниць його, і вчинив, що йому було тяжко ходити. І єгиптяни сказали: Утікаймо від ізраїльтян, бо Господь воює за них з Єгиптом!
EXOD|14|26|І промовив Господь до Мойсея: Простягни свою руку на море, і нехай вернеться вода на єгиптян, на їхні колесниці й на комонників їхніх.
EXOD|14|27|І простяг Мойсей руку свою на море, і море вернулося, коли настав ранок, до сили своєї, а єгиптяни втікали навпроти нього. І кинув Господь єгиптян у середину моря!
EXOD|14|28|І вернулась вода, і позакривала колесниці та комонників усьому фараоновому військові, що ввійшло за ними в море. Ані жоден із них не зостався!
EXOD|14|29|А Ізраїлеві сини йшли суходолом у середині моря, а море було для них муром із правиці їхньої та з лівиці їхньої.
EXOD|14|30|І визволив Господь того дня Ізраїля з єгипетської руки. І бачив Ізраїль мертвих єгиптян на березі моря.
EXOD|14|31|І побачив Ізраїль сильну руку, яку виявив Господь у Єгипті, і став боятися той народ Господа! І ввірував він у Господа, та в Мойсея, раба Його.
EXOD|15|1|Тоді заспівав Мойсей та Ізраїлеві сини оцю пісню Господеві, та й проказали, говорячи: Я буду співать Господеві, бо дійсно звеличився Він, коня й верхівця його кинув до моря!
EXOD|15|2|Моя сила та пісня Господь, і Він став на спасіння мені! Це мій Бог, і прославлю Його, Він Бог батька мого, і звеличу Його!
EXOD|15|3|Господь Муж війни, Єгова Йому Ймення!
EXOD|15|4|Колесниці фараонові й військо його вкинув у море, а вибір його трійкових у Червоному морі затоплений.
EXOD|15|5|Безодні їх позакривали, зійшли до глибин, як той камінь!
EXOD|15|6|Права рука Твоя, Господи, вславлена силою, правиця Твоя трощить ворога, Господи!
EXOD|15|7|А Своєю безмірною величчю Ти розбиваєш Своїх заколотників, посилаєш палючий Свій гнів, він їх поїдає, немов ту солому!
EXOD|15|8|А подувом ніздер Твоїх вода скупчилась, вир спинився, немов та стіна, потоки загусли були в серці моря!
EXOD|15|9|Нахвалявся був ворог: Поженусь дожену! Попаюю здобичу, душа моя сповниться ними! Меча свого вихоплю я, і понищить рука моя їх!
EXOD|15|10|Та дмухнув Ти був духом Своїм і закрило їх море: вони потопились в бурхливій воді, немов оливо!
EXOD|15|11|Хто подібний Тобі серед богів, о Господи? Хто подібний Тобі, Препрославлений святістю? Ти в славі грізний, Чудотворче!
EXOD|15|12|Простягнув Ти правицю Свою і земля їх поглинула!
EXOD|15|13|Милосердям Своїм вів народ, якого Ти визволив, Своєю Ти силою ввів у мешкання Своєї святині!
EXOD|15|14|Почули народи і тремтіли, обгорнула тривога мешканців землі филистимської!
EXOD|15|15|Старшини едомські тоді побентежились, моавських вельмож обгорнуло тремтіння, розпливлися усі ханаанці!
EXOD|15|16|Напали на них страх та жах, через велич рамена Твойого замовкли, як камінь, аж поки перейде народ Твій, о Господи, аж поки перейде народ, що його Ти набув!
EXOD|15|17|Ти їх уведеш, і їх посадиш на гору спадку Твого, на місці, яке вчинив, Господи, житлом Своїм, до Святині Господньої, що поставили руки Твої,
EXOD|15|18|і Господь зацарює навіки віків!
EXOD|15|19|Бо коли ввійшов був до моря кінь фараона з колесницею його та з його комонниками, то Господь повернув на них води морські, а Ізраїлеві сини пішли суходолом у середині моря.
EXOD|15|20|І взяла бубна пророчиця Маріям, сестра Ааронова, а за нею повиходили всі жінки з бубнами та з танцями.
EXOD|15|21|І відповіла їм Маріям: Співайте для Господа, бо дійсно звеличився Він, коня й верхівця його кинув до моря!
EXOD|15|22|І повів Мойсей Ізраїля від Червоного моря, і вийшли вони до пустині Шур. І йшли вони три дні в пустині, і не знаходили води.
EXOD|15|23|І прийшли вони до Мари, і не могли пити води з Мари, бо гірка вона. Тому названо ймення їй: Мара.
EXOD|15|24|І став народ ремствувати на Мойсея, говорячи: Що ми будемо пити?
EXOD|15|25|І він кликав до Господа! І показав йому Господь дерево, і він кинув його до води, і стала вода та солодка! Там Він дав йому постанову та право, і там його випробував.
EXOD|15|26|І сказав Він: Коли дійсно будеш ти слухати голосу Господа, Бога твого, і будеш робити слушне в очах Його, і будеш слухатися заповідей Його, і будеш виконувати всі постанови Його, то всю хворобу, що Я поклав був на Єгипет, не покладу на тебе, бо Я Господь, Лікар твій!
EXOD|15|27|І прийшли вони до Єліму, а там дванадцять водних джерел та сімдесят пальм. І вони отаборилися там над водою.
EXOD|16|1|І рушили вони з Єліму, і вся громада Ізраїлевих синів прибула до пустині Сін, що між Єлімом та між Сінаєм, п'ятнадцятого дня другого місяця по виході їх з єгипетського краю.
EXOD|16|2|І стала ремствувати вся громада Ізраїлевих синів на Мойсея та на Аарона в пустині.
EXOD|16|3|І говорили їм Ізраїлеві сини: Коли б ми були повмирали від Господньої руки в єгипетськім краї, як ми сиділи над горшком м'яса, як ми їли хліба досить! Бо ви вивели нас до цієї пустині, щоб поморити голодом увесь цей збір...
EXOD|16|4|І промовив Господь до Мойсея: Ось Я спускатиму вам дощем хліб із неба, а народ виходитиме й щоденно збиратиме, скільки треба на день, щоб випробувати його, чи буде він ходити в Моєму Законі, чи ні.
EXOD|16|5|А настане шостий день, то приготують, що принесуть, і буде подвійне супроти того, що збирають день-у-день.
EXOD|16|6|І сказали Мойсей та Аарон до всіх Ізраїлевих синів: Настане вечір і ви довідаєтеся, що Господь вивів вас із єгипетського краю.
EXOD|16|7|А настане ранок, то побачите славу Господню, бо Він почув ваші ремствування на Господа. А ми що, що ви ремствуєте на нас?
EXOD|16|8|І сказав Мойсей: Довідаєтесь, як увечорі Господь дасть вам м'яса на їжу, а рано хліба на насичення, бо почув Господь ремствування ваші, що ви ремствуєте на Нього. А ми що? Не на нас ремствування ваше, а на Господа!
EXOD|16|9|І сказав Мойсей до Аарона: Скажи всій громаді Ізраїлевих синів: Наблизьтеся перед лице Господа, бо Він почув ваші ремствування!
EXOD|16|10|І сталося, коли говорив Аарон до всієї громади Ізраїлевих синів, то обернулися вони до пустині, аж ось слава Господня показалася в хмарі!
EXOD|16|11|І промовив Господь до Мойсея, говорячи:
EXOD|16|12|Я почув ремствування Ізраїлевих синів. Промовляй до них, кажучи: Під вечір будете їсти м'ясо, а рано насититесь хлібом, і познаєте, що Я Господь, Бог ваш!
EXOD|16|13|І сталося ввечорі, і знялися перепелиці, і покрили табір. А рано була верства роси навколо табору.
EXOD|16|14|І піднялася верства тієї роси, аж ось на поверхні пустині щось дрібне, вузькувате, дрібне, немов паморозь на землі.
EXOD|16|15|І побачили Ізраїлеві сини, та й казали один до одного: Ман гу?, бо не знали, що то. А Мойсей відказав їм: Це той хліб, що дав вам Господь на їжу.
EXOD|16|16|Це те, що про нього Господь наказав: Збирайте з нього кожен у міру їди своєї, гомер на голову, за числом ваших душ: візьміть кожен для того, хто в наметі його.
EXOD|16|17|І зробили так Ізраїлеві сини, і назбирали хто більше, а хто менше.
EXOD|16|18|І зміряли вони гомером, і не мав зайвого той, хто зібрав більше, а хто зібрав менше, не мав нестачі, зібрали кожен у міру своєї їди!
EXOD|16|19|І сказав до них Мойсей: Нехай ніхто не лишає з нього до ранку!
EXOD|16|20|Та не послухали вони Мойсея, і дехто позоставляли з нього до ранку, а воно зачервивіло, і стало смердюче. І розгнівався на них Мойсей!
EXOD|16|21|І збирали його щоранку, кожен у міру своєї їди. А розгрівалося сонце і воно розтавало.
EXOD|16|22|І сталося шостого дня, поназбирували вони хліба подвійно, два гомери на одного. І посходилися всі начальники громади, і розповіли Мойсеєві.
EXOD|16|23|А він сказав до них: Це те, що говорив Господь: Повний спокій, субота свята для Господа взавтра. Що будете пекти печіть, а що будете варити варіть, а все позостале покладіть собі на сховок до ранку.
EXOD|16|24|І поклали його аж до ранку, як Мойсей наказав, і не засмерділось воно, і черви не було в нім.
EXOD|16|25|І сказав Мойсей: Їжте його сьогодні, бо сьогодні субота для Господа. Сьогодні не знайдете його на полі.
EXOD|16|26|Шість день будете збирати його, а дня сьомого субота: не буде в ній того.
EXOD|16|27|І сталося сьомого дня, повиходили були з народу збирати, та не знайшли.
EXOD|16|28|І сказав Господь до Мойсея: Аж доки ви будете відмовлятися виконувати заповіді Мої та закони Мої?
EXOD|16|29|Побачте, Господь дав вам суботу, тому Він дає вам шостого дня хліба двох днів. Сидіть кожен у себе, нехай сьомого дня не виходить ніхто з свого місця!
EXOD|16|30|І сьомого дня народ відпочивав.
EXOD|16|31|І назвав Ізраїлів дім ім'я тому: манна. Вона була, як коріяндрове насіння, біла, а смак її, як тісто в меду.
EXOD|16|32|І сказав Мойсей: Оце те, що наказав Господь: Наповни нею гомер на сховок для ваших поколінь, щоб бачили той хліб, яким Я годував вас на пустині, коли Я виводив вас із єгипетського краю.
EXOD|16|33|І сказав Мойсей до Аарона: Візьми одну посудину, і поклади туди повний гомер манни, і постав її перед Господнім лицем на сховок для ваших поколінь.
EXOD|16|34|І як наказав Бог Мойсею, так поставив її Аарон перед ковчегом свідоцтва на сховок.
EXOD|16|35|А Ізраїлеві сини їли ту манну сорок літ, аж до прибуття їх до краю заселеного, їли манну аж до приходу їх до границі ханаанського Краю.
EXOD|16|36|А гомер він десята частина ефи.
EXOD|17|1|І рушила вся громада Ізраїлевих синів із пустині Сін на походи свої з наказу Господнього, і отаборилася в Рефідімі. І не було води пити народові.
EXOD|17|2|І сварився народ із Мойсеєм, і казали вони: Дайте нам води, і ми будемо пити! А Мойсей їм сказав: Чого ви сваритеся зо мною? Нащо випробовуєте Господа?
EXOD|17|3|І народ був там спраглий води. І ремствував народ на Мойсея й говорив: Нащо це ти випровадив нас із Єгипту? Щоб повбивати спраглого мене та синів моїх, та отари мої?
EXOD|17|4|І кликав Мойсей до Господа, кажучи: Що я вчиню цьому народові? Ще трохи, і вони вкаменують мене!
EXOD|17|5|І сказав Господь до Мойсея: Перейдися перед народом, і візьми з собою декого з старших Ізраїлевих, а палицю, що нею ти вдарив був Річку, візьми в свою руку, та й іди!
EXOD|17|6|Ось Я стану перед лицем твоїм там, на скелі в Хориві, а ти вдариш у скелю, і вийде із неї вода, і буде пити народ! І зробив Мойсей так на очах старших Ізраїлевих.
EXOD|17|7|І назвав він ім'я того місця: Масса та Мерива через колотнечу Ізраїлевих синів і через випробування ними Господа, коли казали: Чи є Господь серед нас, чи нема?
EXOD|17|8|І прибув Амалик, і воював з Ізраїлем у Рефідімі.
EXOD|17|9|І сказав Мойсей до Ісуса: Вибери нам людей, і вийди воюй з Амаликом. Узавтра я стану на верхів'ї гори, а Божа палиця буде в моїй руці.
EXOD|17|10|І зробив Ісус, як сказав йому Мойсей, щоб воювати з Амаликом. А Мойсей, Аарон та Хур вийшли на верхів'я гори.
EXOD|17|11|І сталося, коли Мойсей підіймав свої руки, то перемагав Ізраїль, а коли руки його опускались, то перемагав Амалик.
EXOD|17|12|А руки Мойсеєві стали тяжкі. І взяли вони каменя, і поклали під ним. І сів він на ньому, а Аарон та Хур підтримували руки йому, один із цього боку, а один із того. І були його руки сталі аж до заходу сонця.
EXOD|17|13|І переміг Ісус Амалика й народ його вістрям меча.
EXOD|17|14|І сказав Господь до Мойсея: Напиши це на пам'ятку в книзі, і поклади до вух Ісусових, що докраю зітру Я пам'ять Амаликову з-під неба.
EXOD|17|15|І збудував Мойсей жертівника, і назвав ім'я йому: Єгова-Ніссі.
EXOD|17|16|І проказав він: Бо рука на Господньому прапорі: Господеві війна з Амаликом із роду в рід!
EXOD|18|1|І почув Їтро, жрець мідіянський, Мойсеїв тесть, усе, що зробив був Бог для Мойсея та для Свого народу Ізраїлевого, що вивів Господь Ізраїля з Єгипту.
EXOD|18|2|І взяв Їтро, Мойсеїв тесть, жінку Мойсеєву Ціппору, по відісланні її,
EXOD|18|3|та обох синів її, що ймення одному Ґершом, бо сказав був: Я став приходьком у чужому краї,
EXOD|18|4|а ймення другому Еліезер, бо Бог мого батька був мені поміччю, і визволив мене від фараонового меча.
EXOD|18|5|І прибув Їтро, тесть Мойсеїв, і сини його та жінка його до Мойсея в пустиню, де він отаборився там біля Божої гори.
EXOD|18|6|І сказав він до Мойсея: Я, тесть твій Їтро, приходжу до тебе, і жінка твоя, і обидва сини її з нею.
EXOD|18|7|І вийшов Мойсей навпроти свого тестя, та й уклонився до землі, і поцілував його. І питали вони один одного про мир, і ввійшли до намету.
EXOD|18|8|І оповів Мойсей своєму тестеві про все, що зробив був Господь фараонові та Єгиптові через Ізраїля, про всі ті труднощі, які він спіткав був по дорозі, та Господь визволив їх.
EXOD|18|9|І тішився Їтро всім тим добром, що вчинив Господь для Ізраїля, що визволив його з єгипетської руки.
EXOD|18|10|І промовив Їтро: Благословенний Господь, що визволив вас з єгипетської руки та з руки фараонової, що визволив народ з-під руки єгипетської.
EXOD|18|11|Тепер я знаю, що Господь більший за всіх богів, бо зробив це за те, що єгиптяни вихвалялись над ними.
EXOD|18|12|І взяв Їтро, Мойсеїв тесть, цілопалення та жертви для Бога. І прийшов Аарон та всі старші Ізраїлеві їсти хліб з Мойсеєвим тестем перед Божим обличчям.
EXOD|18|13|І сталося назавтра, і сів Мойсей судити народ, а народ стояв навколо Мойсея від ранку аж до вечора.
EXOD|18|14|І побачив тесть Мойсеїв усе, що він робить народові, та й сказав: Що це за річ, що ти робиш народові? Для чого ти сидиш сам один, а ввесь народ стоїть навколо від ранку аж до вечора?
EXOD|18|15|А Мойсей відказав своєму тестеві: Бо народ приходить до мене питатися суду Бога.
EXOD|18|16|Бо як мають вони справу, то приходять до мене, і я суджу поміж тим і тим, та оголошую постанови Божі та закони Його.
EXOD|18|17|І сказав тесть Мойсеїв до нього: Недобра ця річ, що ти чиниш.
EXOD|18|18|Справді стомишся і ти, і народ той, що з тобою, бо ця справа тяжча за тебе. Не потрапиш ти чинити її сам один!
EXOD|18|19|Тепер послухай мого слова, пораджу тобі, і буде Бог із тобою! Стій за народ перед Богом, і принось справи до Бога.
EXOD|18|20|І ти остережеш їх за постанови та за закони, і об'явиш їм ту путь, якою вони підуть, і те діло, яке вони зроблять.
EXOD|18|21|А ти наздриш зо всього народу мужів здібних, богобоязливих, мужів справедливих, що ненавидять зиск, і настановиш їх над ними тисяцькими, сотниками, п'ятдесятниками та десятниками.
EXOD|18|22|І будуть вони судити народ кожного часу. І станеться, кожну велику справу вони принесуть до тебе, а кожну малу справу розсудять самі. Полегши собі, і нехай вони несуть тягар із тобою.
EXOD|18|23|Коли ти зробиш цю річ, а Бог тобі накаже, то ти втримаєшся, а також увесь народ цей прийде на своє місце в мирі.
EXOD|18|24|І послухався Мойсей голосу тестя свого, і зробив усе, що той був сказав.
EXOD|18|25|І вибрав Мойсей здібних мужів зо всього Ізраїля, і настановив їх начальниками над народом, тисяцькими, сотниками, п'ятдесятниками та десятниками.
EXOD|18|26|І судили вони народ кожного часу. Справу трудну приносили Мойсеєві, а кожну малу справу судили самі.
EXOD|18|27|І відпустив Мойсей тестя свого, і він пішов собі до краю свого.
EXOD|19|1|Третього місяця по виході Ізраїлевих синів із єгипетського краю, того дня прибули вони на Сінайську пустиню.
EXOD|19|2|І рушили вони з Рефідіму, і ввійшли до Сінайської пустині, та й отаборилися в пустині. І отаборився там Ізраїль навпроти гори.
EXOD|19|3|А Мойсей увійшов до Бога. І кликнув до нього Господь із гори, говорячи: Скажеш отак дому Якова, і звістиш синам Ізраїля:
EXOD|19|4|Ви бачили, що Я зробив був Єгиптові, і носив вас на крилах орлиних, і привів вас до Себе.
EXOD|19|5|А тепер, коли справді послухаєте Мого голосу, і будете дотримувати заповіту Мого, то станете Мені власністю більше всіх народів, бо вся земля то Моя!
EXOD|19|6|А ви станете Мені царством священиків та народом святим. Оце ті речі, що про них будеш казати Ізраїлевим синам.
EXOD|19|7|І прибув Мойсей, і покликав старших народніх, та й виложив перед ними всі ті слова, що Господь наказав був йому.
EXOD|19|8|І відповів увесь народ разом, та й сказав: Усе, що Господь говорив, зробимо! А Мойсей доніс слова народу до Господа.
EXOD|19|9|І промовив Господь до Мойсея: Ось Я до тебе прийду в густій хмарі, щоб чув народ, коли Я говоритиму з тобою, і щоб повірив і тобі навіки! І переповів Мойсей слова народу до Господа.
EXOD|19|10|І промовив Господь до Мойсея: Іди до людей, і освяти їх сьогодні та взавтра, і нехай вони виперуть одіж свою.
EXOD|19|11|І нехай вони будуть готові на третій день, бо третього дня зійде Господь на гору Сінай на очах усього народу.
EXOD|19|12|І обведеш границею народ довкола, говорячи: Стережіться сходити на гору й доторкуватися до краю її. Кожен, хто доторкнеться до гори, буде конче забитий!
EXOD|19|13|Нехай не доторкнеться до неї рука, бо буде конче вкаменований, або буде справді застрілений, чи то худобина, чи то людина, не буде жити вона. Як сурма засурмить протяжливо, вони вийдуть на гору.
EXOD|19|14|І зійшов Мойсей з гори до народу, і освятив народ, а вони випрали одежу свою.
EXOD|19|15|І він сказав до народу: Будьте готові на третій день; не входьте до жінок.
EXOD|19|16|І сталося третього дня, коли ранок настав, і знялися громи та блискавки, і густа хмара над горою та сильний голос сурми! І затремтів увесь народ, що був у таборі...
EXOD|19|17|І вивів Мойсей народ із табору назустріч Богові, і вони стали під горою.
EXOD|19|18|А гора Сінай уся вона димувала через те, що Господь зійшов на неї в огні! І піднявся дим її, немов дим вапнярки, і сильно затремтіла вся гора...
EXOD|19|19|І розлігся голос сурми, і він сильно все могутнів: Мойсей говорить, а Бог відповідає йому голосно...
EXOD|19|20|І зійшов Господь на гору Сінай, на верхів'я гори. І покликав Господь Мойсея на верхів'я гори. І вийшов Мойсей.
EXOD|19|21|І промовив Господь до Мойсея: Зійди, остережи народ, щоб не рвався до Господа, щоб побачити, бо багато з нього загине.
EXOD|19|22|А також священики, що будуть підходити до Господа, нехай перше освятяться, щоб Господь їх не повбивав.
EXOD|19|23|І сказав Мойсей до Господа: Не зможе народ вийти на гору Сінай, бо Ти засвідчив між нами, говорячи: Обведи границею цю гору, і освяти її.
EXOD|19|24|І промовив до нього Господь: Іди, зійди, а потім вийди ти й Аарон з тобою, а священики й народ нехай не рвуться до Господа, щоб Я не повбивав їх.
EXOD|19|25|І зійшов Мойсей до народу, і сказав їм це все.
EXOD|20|1|І Бог промовляв всі слова оці, кажучи:
EXOD|20|2|Я Господь, Бог твій, що вивів тебе з єгипетського краю з дому рабства.
EXOD|20|3|Хай не буде тобі інших богів передо Мною!
EXOD|20|4|Не роби собі різьби і всякої подоби з того, що на небі вгорі, і що на землі долі, і що в воді під землею.
EXOD|20|5|Не вклоняйся їм і не служи їм, бо Я Господь, Бог твій, Бог заздрісний, що карає за провину батьків на синах, на третіх і на четвертих поколіннях тих, хто ненавидить Мене,
EXOD|20|6|і що чинить милість тисячам поколінь тих, хто любить Мене, і хто держиться Моїх заповідей.
EXOD|20|7|Не призивай Імення Господа, Бога твого, надаремно, бо не помилує Господь того, хто призиватиме Його Ймення надаремно.
EXOD|20|8|Пам'ятай день суботній, щоб святити його!
EXOD|20|9|Шість день працюй і роби всю працю свою,
EXOD|20|10|а день сьомий субота для Господа, Бога твого: не роби жодної праці ти й син твій, та дочка твоя, раб твій та невільниця твоя, і худоба твоя, і приходько твій, що в брамах твоїх.
EXOD|20|11|Бо шість день творив Господь небо та землю, море та все, що в них, а дня сьомого спочив тому поблагословив Господь день суботній і освятив його.
EXOD|20|12|Шануй свого батька та матір свою, щоб довгі були твої дні на землі, яку Господь, Бог твій, дає тобі!
EXOD|20|13|Не вбивай!
EXOD|20|14|Не чини перелюбу!
EXOD|20|15|Не кради!
EXOD|20|16|Не свідкуй неправдиво на свого ближнього!
EXOD|20|17|Не жадай дому ближнього свого, не жадай жони ближнього свого, ані раба його, ані невільниці його, ані вола його, ані осла його, ані всього, що ближнього твого!
EXOD|20|18|І ввесь народ бачив та чув громи та полум'я, і голос сурми, і гору димлячу. І побачив народ, і всі тремтіли та й поставали здалека.
EXOD|20|19|І сказали вони до Мойсея: Говори з нами ти, і ми послухаємо, а нехай не говорить із нами Бог, щоб ми не повмирали.
EXOD|20|20|І промовив Мойсей до народу: Не бійтеся, бо Бог прибув для випробування вас, і щоб страх Його був на ваших обличчях, щоб ви не грішили.
EXOD|20|21|І став народ здалека, а Мойсей підійшов до мороку, де був Бог.
EXOD|20|22|І промовив Господь до Мойсея: Отак скажеш до Ізраїлевих синів: Ви бачили, що Я говорив з вами з небес.
EXOD|20|23|Не будете робити при Мені богів із срібла, і богів із золота не будете робити собі.
EXOD|20|24|Ти зробиш для Мене жертівника з землі, і будеш приносити на ньому свої цілопалення й свої мирні жертви, і дрібну худобу свою, і велику худобу свою. На кожному місці, де Я згадаю Ймення Своє, Я до тебе прийду й поблагословлю тебе.
EXOD|20|25|А коли зробиш Мені жертівника з каменів, то не будеш будувати його з обтесаних, бо ти підносив би над ним знаряддя своє, і занечистив би його.
EXOD|20|26|І не будеш входити до Мого жертівника ступенями, щоб не була відкрита при ньому твоя нагота.
EXOD|21|1|А оце закони, що ти викладеш перед ними:
EXOD|21|2|Коли купиш єврейського раба, нехай він працює шість років, а сьомого нехай вийде дармо на волю.
EXOD|21|3|Якщо прийде він сам один, нехай сам один і вийде; коли він має жінку, то з ним вийде й жінка його.
EXOD|21|4|Якщо пан його дасть йому жінку, і вона породить йому синів або дочок, та жінка та діти її нехай будуть для пана її, а він нехай вийде сам один.
EXOD|21|5|А якщо раб той щиро скаже: Полюбив я пана свого, жінку свою та дітей своїх, не вийду на волю,
EXOD|21|6|то нехай його пан приведе його до суддів, і підведе його до дверей або до бічних одвірків, та й проколе пан його вухо йому шилом, і він буде робити йому повіки!
EXOD|21|7|А коли хто продасть дочку свою на невільницю, не вийде вона, як виходять раби.
EXOD|21|8|Якщо вона невгодна в очах свого пана, який призначив був її собі, то нехай позволить її викупити. Не вільно йому продати її до народу чужого, коли зрадить її.
EXOD|21|9|А якщо призначить її для сина свого, то зробить їй за правом дочок.
EXOD|21|10|Якщо візьме собі іншу, то не зменшить поживи їй, одежі їй і подружнього пожиття їй.
EXOD|21|11|А коли він цих трьох речей не робитиме їй, то вона вийде дармо, без окупу.
EXOD|21|12|Хто вдарить людину, і вона вмре, той конче буде забитий.
EXOD|21|13|А хто не чатував, а Бог підвів кого в його руку, то дам тобі місце, куди той утече.
EXOD|21|14|А коли хто буде замишляти на ближнього свого, щоб забити його з хитрістю, візьмеш його від жертівника Мого на смерть.
EXOD|21|15|А хто вдарить батька свого чи матір свою, той конче буде забитий.
EXOD|21|16|А хто вкраде людину і продасть її, або буде вона знайдена в руках його, той конче буде забитий.
EXOD|21|17|І хто проклинає батька свого чи свою матір, той конче буде забитий.
EXOD|21|18|А коли будуть сваритися люди, і вдарить один одного каменем або кулаком, і той не вмре, а зляже на постелю,
EXOD|21|19|якщо встане й буде проходжуватися надворі з опертям своїм, то буде оправданий той, хто вдарив, тільки нехай дасть за прогаяння часу його та справді вилікує.
EXOD|21|20|А коли хто вдарить раба свого або невільницю свою києм, а той помре під рукою його, то конче буде покараний той.
EXOD|21|21|Тільки якщо той переживе день або два дні, то не буде покараний, бо він його гроші.
EXOD|21|22|А коли будуть битися люди, і вдарять вагітну жінку, і скине вона дитину, а іншого нещастя не станеться, то конче буде покараний, як покладе на нього чоловік тієї жінки, і він дасть за присудом суддів.
EXOD|21|23|А якщо станеться нещастя, то даси душу за душу,
EXOD|21|24|око за око, зуба за зуба, руку за руку, ногу за ногу,
EXOD|21|25|опарення за опарення, рану за рану, синяка за синяка.
EXOD|21|26|А коли хто вдарить в око раба свого, або в око невільниці своєї, і знищить його, той на волю відпустить його за око його.
EXOD|21|27|А якщо виб'є зуба раба свого, або зуба невільниці своєї, той на волю відпустить того за зуба його.
EXOD|21|28|А коли віл ударить чоловіка або жінку, а той умре, конче буде вкаменований той віл, і м'ясо його не буде їджене, а власник того вола невинний.
EXOD|21|29|А якщо віл був битливим і вчора, і третього дня, і було те засвідчене у власника його, а той його не пильнував, і заб'є той віл чоловіка або жінку, буде він укаменований, а також власник буде забитий.
EXOD|21|30|Якщо на нього буде накладений викуп, то дасть викупа за душу свою, скільки буде на нього накладене.
EXOD|21|31|Або вдарить віл сина, або вдарить дочку, буде зроблено йому за цим законом.
EXOD|21|32|Коли вдарить той віл раба або невільницю, то власник дасть панові того тридцять шеклів срібла, а віл той буде вкаменований.
EXOD|21|33|А коли хто розкриє яму, або викопає яму й не закриє її, і впаде туди віл або осел,
EXOD|21|34|власник ями відшкодує, верне гроші власникові його, а загинуле буде йому.
EXOD|21|35|А коли чийсь віл ударить вола його ближнього, і згине той, то продадуть вола живого, а гроші за нього поділять пополовині, і також загинулого поділять пополовині.
EXOD|21|36|А коли буде відоме, що віл був битливим і вчора й третього дня, а власник його не пильнував його, то конче нехай відшкодує вола за того вола, а забитий буде йому.
EXOD|22|1|(21-37) Коли хто вкраде вола або овечку, і заріже його або продасть його, то відшкодує п'ять штук великої худоби за вола того, а чотири дрібної худоби за ту овечку.
EXOD|22|2|(22-1) Коли злодій буде зловлений в підкопі, і буде побитий так, що помре, то нема провини крови на тому, хто побив.
EXOD|22|3|(22-2) Але як засвітило сонце над ним, то є на ньому провина крови. Злодій конче відшкодує, а якщо він нічого не має, то буде проданий за свою крадіжку.
EXOD|22|4|(22-3) Якщо та крадіжка справді буде знайдена в руці його живою, від вола аж до осла, до ягняти, то нехай відшкодує удвоє.
EXOD|22|5|(22-4) Коли хто випасе поле або виноградника, і пустить свою худобу й буде випасати на чужому полі, відшкодує найліпшим із поля свого й найліпшим із свого виноградника.
EXOD|22|6|(22-5) Коли вийде огонь і попаде на тернину, і буде спалена скирта, або збіжжя стояче, або поле, конче відшкодує той, хто запалив пожежу.
EXOD|22|7|(22-6) Коли хто дасть своєму ближньому срібло або посуд на збереження, а воно буде вкрадене з дому того чоловіка, якщо буде знайдений злодій, нехай відшкодує вдвоє.
EXOD|22|8|(22-7) Якщо ж злодій не буде знайдений, то власник дому буде приведений до суддів, на присягу, що не простягав своєї руки на працю свого ближнього.
EXOD|22|9|(22-8) У кожній справі провини, про вола, про осла, про овечку, про одіж, про все згублене, про яке хто скаже, що це його, нехай справа обох прийде до судді. Кого суддя визнає за винного, той відшкодує вдвоє своєму ближньому.
EXOD|22|10|(22-9) Коли хто дасть своєму ближньому на збереження осла, або вола, або овечку, чи яку іншу худобину, а вона згине, або буде скалічена, або буде заграбована, і ніхто того не бачив,
EXOD|22|11|(22-10) присяга Господня нехай буде між обома, що він не простяг своєї руки на власність свого ближнього, а власник її нехай забере, а позваний не буде відшкодувати.
EXOD|22|12|(22-11) А якщо справді буде вкрадена від нього, то нехай відшкодує власникові її.
EXOD|22|13|(22-12) Якщо дійсно буде розшарпана вона, нехай принесе її як свідоцтво, а за розшарпане він не відшкодує.
EXOD|22|14|(22-13) А коли хто позичить від свого ближнього худобину, а вона буде скалічена або згине, а власник її не був із нею, то конче відшкодує;
EXOD|22|15|(22-14) якщо ж її власник був із нею, не відшкодує. А якщо худобина була найнята, то піде та шкода в заплату її.
EXOD|22|16|(22-15) А коли хто підмовить дівчину, яка не заручена, і ляже з нею, то нехай дасть їй віно, і візьме її собі за жінку.
EXOD|22|17|(22-16) Якщо батько її справді відмовить віддати її йому, нехай відважить срібла згідно з віном дівочим.
EXOD|22|18|(22-17) Чарівниці не зоставиш при житті.
EXOD|22|19|(22-18) Кожен, хто зляжеться з худобиною, конче буде забитий.
EXOD|22|20|(22-19) Кожен, хто приносить жертву богам, крім Бога Одного, підпадає закляттю.
EXOD|22|21|(22-20) А приходька не будеш утискати та гнобити його, бо й ви були приходьками в єгипетськім краї.
EXOD|22|22|(22-21) Жодної вдови та сироти не будеш гнобити;
EXOD|22|23|(22-22) якщо ж ти справді гнобитимеш їх, то коли вони, кличучи, кликатимуть до Мене, то конче почую їхній зойк,
EXOD|22|24|(22-23) і розпалиться гнів Мій, і повбиваю вас мечем, і стануть жінки ваші вдовами, а діти ваші сиротами.
EXOD|22|25|(22-24) Якщо позичиш гроші народові Моєму, бідному, що з тобою, то не будь йому, як суворий позичальник, не покладеш на нього лихви.
EXOD|22|26|(22-25) Якщо дійсно візьмеш у заставу одежу ближнього свого, то вернеш її йому до заходу сонця,
EXOD|22|27|(22-26) бо вона єдине накриття його, вона одіж на тіло його; на чому він буде лежати? І станеться, коли буде він кликати до Мене, то почую, бо Я милосердний.
EXOD|22|28|(22-27) Бога не будеш лихословити, а начальника в народі твоїм не будеш проклинати.
EXOD|22|29|(22-28) Не будеш спізнюватися, щодо жертов, із щедрістю збіжжя та з плинами твоїми. Перворідного з синів своїх даси Мені.
EXOD|22|30|(22-29) Так зробиш волові своєму, і дрібній худобі своїй: сім день буде вона з своєю матір'ю, а восьмого дня даси її Мені.
EXOD|22|31|(22-30) І ви будете Мені святими людьми, і не будете їсти м'яса, розшарпаного в полі, псові кинете його!
EXOD|23|1|Не будеш розносити неправдивих поголосок. Не покладеш руки своєї з несправедливим, щоб бути свідком неправди.
EXOD|23|2|Не будеш з більшістю, щоб чинити зло. І не будеш висловлюватися про позов, прихиляючись до більшости, щоб перегнути правду.
EXOD|23|3|І не будеш потурати вбогому в його позові.
EXOD|23|4|Коли стрінеш вола свого ворога або осла його, що заблудив, то конче повернеш його йому.
EXOD|23|5|Коли побачиш осла свого ворога, що лежить під тягарем своїм, то не загаїшся помогти йому, конче поможеш разом із ним.
EXOD|23|6|Не перегинай суду на бік вбогого свого в його позові.
EXOD|23|7|Від неправдивої справи віддалишся, а чистого й справедливого не забий, бо Я не всправедливлю несправедливого.
EXOD|23|8|А хабара не візьмеш, бо хабар осліплює зрячих і викривляє слова справедливих.
EXOD|23|9|А приходька не будеш тиснути, бож ви познали душу приходька, бо самі були приходьками в єгипетськім краї.
EXOD|23|10|І шість літ будеш сіяти землю свою, і будеш збирати її врожай,
EXOD|23|11|а сьомого опустиш її та полишиш її, і будуть їсти вбогі народу твого, а позостале по них буде їсти польова звірина. Так само зробиш для виноградника твого, і для оливки твоєї.
EXOD|23|12|Шість день будеш робити діла свої, а сьомого дня спочинеш, щоб відпочив віл твій, і осел твій, і щоб відідхнув син невільниці твоєї й приходько.
EXOD|23|13|І все, що Я сказав вам, будете виконувати. А ймення інших богів не згадаєте, не буде почуте воно на устах твоїх.
EXOD|23|14|Три рази на рік будеш святкувати Мені.
EXOD|23|15|Будеш дотримувати свято Опрісноків; сім день будеш їсти опрісноки, як наказав тобі, окресленого часу місяця авіва, бо в нім ти був вийшов з Єгипту. І не будете являтися перед лицем Моїм з порожніми руками.
EXOD|23|16|І свято жнив первоплоду праці твоєї, що сієш на полі. І свято збирання при закінченні року, коли ти збираєш з поля працю свою.
EXOD|23|17|Три рази на рік буде являтися ввесь чоловічий рід твій перед лицем Владики Господа.
EXOD|23|18|Не будеш приносити крови жертви Моєї на квашенім, а лій Моєї святкової жертви не буде ночувати аж до ранку.
EXOD|23|19|Початки первоплоду твоєї землі принесеш до дому Господа, Бога твого. Не будеш варити ягняти в молоці його матері.
EXOD|23|20|Ось Я посилаю Ангола перед лицем твоїм, щоб він охороняв у дорозі тебе, і щоб провадив тебе до того місця, яке Я приготовив.
EXOD|23|21|Стережися перед лицем Його, і слухайся Його голосу! Не протився Йому, бо Він не пробачить вашого гріха, бо Ім'я Моє в Ньому.
EXOD|23|22|Коли ж справді послухаєш ти його голосу, і вчиниш усе, що говорю, то Я буду ворогувати проти ворогів твоїх, і буду гнобити твоїх гнобителів.
EXOD|23|23|Бо Мій Ангол ходитиме перед лицем твоїм, і запровадить тебе до амореянина, і хіттеянина, і періззеянина, і ханаанеянина, хіввеянина, і євусеянина, а Я знищу його.
EXOD|23|24|Не будеш вклонятися їхнім богам, і служити їм не будеш, і не будеш чинити за вчинками їх, бо конче порозбиваєш і конче поламаєш їхні стовпи для богів.
EXOD|23|25|І будеш служити ти Господеві, Богові своєму, і Він поблагословить твій хліб та воду твою, і з-посеред тебе усуне хворобу.
EXOD|23|26|У твоїм Краї не буде такої, що скидає плода, ані неплідної. Число твоїх днів Я доповню.
EXOD|23|27|Свій страх пошлю перед лицем твоїм, і приведу в замішання ввесь цей народ, що ти ввійдеш між нього. І всіх ворогів твоїх оберну до тебе потилицею.
EXOD|23|28|І пошлю шершня перед тобою, і він вижене перед тобою хіввеянина, ханаанеянина та хіттеянина.
EXOD|23|29|Не вижену їх перед тобою в однім році, щоб не став той Край спустошеним, і не розмножилася на тебе польова звірина.
EXOD|23|30|Помалу Я буду їх виганяти перед тобою, аж поки ти розродишся, і посядеш цей Край.
EXOD|23|31|І покладу границю твою від моря Червоного й аж до моря Филистимського, і від пустині аж до Річки, бо дам в вашу руку мешканців цього Краю, і ти виженеш їх перед собою.
EXOD|23|32|Не складай умови з ними та з їхніми богами.
EXOD|23|33|Не будуть сидіти вони в твоїм Краї, щоб не ввести тебе в гріх супроти Мене, коли будеш служити їхнім богам, бо це буде пастка тобі!
EXOD|24|1|А до Мойсея сказав Він: Вийди до Господа ти й Аарон, Надав та Авігу, та сімдесят із Ізраїлевих старших, і вклоніться здалека.
EXOD|24|2|А Мойсей нехай підійде до Господа сам, а вони не підійдуть. А народ з ним не вийде.
EXOD|24|3|І прибув Мойсей, та й оповів народові всі Господні слова та всі закони. І ввесь народ відповів одноголосно, та й сказали: Усе, про що говорив Господь, зробимо!
EXOD|24|4|І написав Мойсей всі Господні слова. І встав він рано вранці, та й збудував жертівника під горою, та дванадцять кам'яних стовпів для дванадцяти Ізраїлевих племен.
EXOD|24|5|І послав він юнаків, синів Ізраїлевих, і вони зложили цілопалення, і принесли жертви, мирні жертви для Господа, бички.
EXOD|24|6|І взяв Мойсей половину крови, і вилив до мідниць, а другу половину тієї крови вилив на жертівника.
EXOD|24|7|І взяв він книгу заповіту, та й відчитав вголос народові. А вони сказали: Усе, що говорив Господь, зробимо й послухаємо!
EXOD|24|8|І взяв Мойсей тієї крови, і покропив на народ, та й сказав: Оце кров заповіту, що Господь уклав із вами про всі оці речі!
EXOD|24|9|І вийшов Мойсей й Аарон, Надав та Авігу, та сімдесят Ізраїлевих старших,
EXOD|24|10|і вони споглядали на Ізраїлевого Бога, а під ногами Його ніби зроблене з сапфірової плити, і немов саме небо, щодо ясности.
EXOD|24|11|І він не простяг Своєї руки на достойних із синів Ізраїля. І вони споглядали на Бога, і їли й пили.
EXOD|24|12|І промовив Господь до Мойсея: Вийди до Мене на гору, і будь там. І дам тобі кам'яні таблиці, і закона та заповідь, що Я написав для навчання їх.
EXOD|24|13|І встав Мойсей та Ісус, слуга його, і вийшов Мойсей на Божу гору.
EXOD|24|14|А до старших сказав він: Сидіть нам на цім місці, аж поки ми вернемось до вас! А ось Аарон та Хур будуть із вами. Хто матиме справу, нехай прийде до них.
EXOD|24|15|І вийшов Мойсей на гору, а хмара закрила гору.
EXOD|24|16|І слава Господня спочивала на горі Сінай, а хмара закривала її шість день. А сьомого дня Він кликнув до Мойсея з середини хмари.
EXOD|24|17|А вид Господньої слави як огонь, що пожирає на верхів'ї гори, на очах Ізраїлевих синів.
EXOD|24|18|І ввійшов Мойсей у середину хмари, і вийшов на гору. І Мойсей пробував на горі сорок день та сорок ночей.
EXOD|25|1|А Господь промовляв до Мойсея, говорячи:
EXOD|25|2|Промовляй до Ізраїлевих синів, і нехай вони візьмуть для Мене приношення. Від кожного мужа, що дасть добровільно його серце, візьмете приношення для Мене.
EXOD|25|3|А оце те приношення, що візьмете від них: золото, і срібло, і мідь,
EXOD|25|4|і блакить, і пурпур, і червень, і віссон, і козина вовна,
EXOD|25|5|і шкурки баранячі, начервоно пофарбовані, і шкурки тахашеві, і дерево акацій,
EXOD|25|6|олива на освітлення, пахощі до оливи намащення, і пахощі для кадила,
EXOD|25|7|і каміння оніксове, і каміння на оправу до ефоду й до нагрудника.
EXOD|25|8|І нехай збудують Мені святиню, і перебуватиму серед них.
EXOD|25|9|Як усе, що Я покажу тобі будову скинії та будову речей її, і так зробите.
EXOD|25|10|І зроблять вони ковчега з акаційного дерева, два лікті й пів довжина його, і лікоть і пів ширина його, і лікоть і пів вишина його.
EXOD|25|11|І пообкладаєш його щирим золотом зсередини та іззовні. І зробиш вінця золотого навколо над ним.
EXOD|25|12|І виллєш для нього чотири золоті каблучки, і даси на чотирьох кутах його, дві каблучки на одному боці його, і дві каблучки на другому боці його.
EXOD|25|13|І поробиш держаки з акаційного дерева, і пообкладаєш їх золотом.
EXOD|25|14|І повсовуєш ці держаки в каблучки на боках ковчегу, щоб ними носити ковчега.
EXOD|25|15|В ковчегових каблучках будуть ці держаки; не відступлять вони від нього.
EXOD|25|16|І покладеш до ковчегу те свідоцтво, що Я тобі дам.
EXOD|25|17|І зробиш віко зо щирого золота, два лікті й пів довжина його, і лікоть і пів ширина його.
EXOD|25|18|І зробиш два золоті херувими, роботою кутою зробиш їх з обох кінців віка.
EXOD|25|19|І зроби одного херувима з кінця звідси, а одного херувима з кінця звідти. Від того віка поробите тих херувимів на обох кінцях його.
EXOD|25|20|І будуть ті херувими простягати крила догори, і затінювати своїми крильми над віком, а їхні обличчя одне до одного; до віка будуть обличчя тих херувимів.
EXOD|25|21|І покладеш те віко згори на ковчега, а до цього ковчега покладеш свідоцтво, яке Я тобі дам.
EXOD|25|22|І Я буду тобі відкриватися там, і буду говорити з тобою з-над віка з-посеред обох херувимів, що над ковчегом свідоцтва, про все, що розповім тобі для синів Ізраїлевих.
EXOD|25|23|І зробиш стола з акаційного дерева, два лікті довжина його, і лікоть ширина його, і лікоть і пів вишина його.
EXOD|25|24|І пообкладаєш його щирим золотом, і зробиш вінця золотого для нього навколо.
EXOD|25|25|І лиштву зробиш для нього в долоню навколо, і зробиш вінця золотого навколо, для лиштви його.
EXOD|25|26|І зробиш для нього чотири каблучки із золота, та й даси ці каблучки на чотирьох кінцях, що при його чотирьох ніжках.
EXOD|25|27|Навпроти лиштви будуть ці каблучки, на вкладання для держаків, щоб носити стола.
EXOD|25|28|І поробиш ті держаки з акаційного дерева, і пообкладаєш їх золотом, і на них будуть носити стола.
EXOD|25|29|І поробиш миски його, і кадильниці його, і чаші його та кухлі його, щоб ними лити, зо щирого золота їх ти поробиш.
EXOD|25|30|А на столі покладеш хліб показний, що завжди перед Моїм лицем.
EXOD|25|31|І зробиш свічника зо щирого золота, роботою кутою нехай буде зроблено цього свічника. Стовп його, і рамена його, келихи його, ґудзі його й квітки його будуть із нього.
EXOD|25|32|І шість рамен виходитимуть із боків його, три рамені свічника з одного боку його, і три рамені свічника з другого боку його.
EXOD|25|33|Три келихи мигдалоподібні в однім рамені, ґудзь і квітка, і три мигдалоподібні келихи в рамені другім, ґудзь і квітка. Так на шости раменах, що виходять із свічника.
EXOD|25|34|А на стовпі свічника чотири келихи мигдалоподібні, ґудзі його та квітки його.
EXOD|25|35|І ґудзь під двома раменами з нього, і ґудзь під іншими двома раменами з нього, і ґудзь під третіми двома раменами з нього, у шости рамен, що виходять із свічника.
EXOD|25|36|Їхні ґудзі та їхні рамена нехай будуть із нього. Увесь він одне куття щирого золота.
EXOD|25|37|І зробиш сім лямпадок до нього, і нехай засвітять його лямпадки, і нехай він світить на передню сторону його.
EXOD|25|38|А його щипчики та його лопатки на вугіль щире золото.
EXOD|25|39|З таланту щирого золота зробиш його та ввесь цей посуд.
EXOD|25|40|І дивись, і зроби за тим зразком, що тобі показувано на горі.
EXOD|26|1|А скинію зробиш із десяти покривал із суканого віссону, і блакиті, і пурпуру та з червені. Херувими мистецькою роботою зробиш ти їх.
EXOD|26|2|Довжина одного покривала двадцять і вісім ліктів, а ширина одного покривала чотири лікті. Усім покривалам міра одна.
EXOD|26|3|П'ять покривал буде поспинаних одне до одного, і п'ять покривал інших буде поспинаних одне до одного.
EXOD|26|4|І поробиш блакитні петельки на краю одного покривала з кінця в спинанні. І так само зробиш на краю кінцевого покривала в спинанні другім.
EXOD|26|5|П'ятдесят петельок поробиш у покривалі однім, і п'ятдесят петельок поробиш на кінці покривала, що в другім спинанні. Ті петельки протилеглі одна до однієї.
EXOD|26|6|І зробиш п'ятдесят золотих гачків, і поспинаєш ті покривала одне до одного тими гачками, і буде одна скинія.
EXOD|26|7|І проробиш покривала з вовни козиної на намета над внутрішньою скинією, зробиш їх одинадцять покривал.
EXOD|26|8|Довжина одного покривала тридцять ліктів, а ширина одного покривала чотири лікті. Одинадцятьом покривалам міра одна.
EXOD|26|9|І поспинаєш п'ять покривал осібно, і шість покривал осібно, а шосте покривало складеш удвоє напереді намету.
EXOD|26|10|І поробиш п'ятдесят петельок на краю одного покривала, кінцевого в спинанні, і п'ятдесят петельок на краю покривала другого спинання.
EXOD|26|11|І зробиш п'ятдесят мідяних гачків, і повсовуєш ті гачки в петельки і поспинаєш намета, і буде він один.
EXOD|26|12|А те, що звисає, лишок в наметових покривалах, половина залишку покривала, буде звисати ззаду скинії.
EXOD|26|13|І лікоть із цього, і лікоть із того боку в залишку в довжині наметового покривала буде звішений на боки скинії з цього й з того боку на покриття її.
EXOD|26|14|І зробиш накриття для скинії, баранячі начервоно пофарбовані шкурки, і накриття зверху з тахашевих шкурок.
EXOD|26|15|І поробиш для скинії стоячі дошки з акаційного дерева.
EXOD|26|16|Десять ліктів довжина дошки, і лікоть і півліктя ширина однієї дошки.
EXOD|26|17|В одній дошці дві ручки, сполучені одна до однієї. Так зробиш усім дошкам скинійним.
EXOD|26|18|І поробиш дошки для скинії, двадцять дощок на бік південний, на полудень.
EXOD|26|19|І сорок срібних підстав поробиш під тими двадцятьма дошками, дві підставі під однією дошкою для двох ручок її, і дві підставі під дошкою другою для двох ручок її.
EXOD|26|20|А для другого боку скинії, в сторону півночі двадцять дощок.
EXOD|26|21|І для них сорок срібних підстав, дві підставі під одну дошку, і дві підставі під дошку другу.
EXOD|26|22|А для заднього боку скинії на захід зробиш шість дощок.
EXOD|26|23|І дві дошки зробиш для кутів скинії на заднього бока.
EXOD|26|24|І нехай вони будуть поєднані здолу, і нехай разом будуть поєднані на верху її до однієї каблучки. Так нехай буде для обох них; нехай вони будуть для обох кутів.
EXOD|26|25|І буде вісім дощок, а їхні підстави зо срібла, шістнадцять підстав: дві підставі під одну дошку, і дві під дошку другу.
EXOD|26|26|І зробиш засуви з акаційного дерева, п'ять для дощок одного боку скинії,
EXOD|26|27|і п'ять засувів для дощок другого боку скинії, і п'ять засувів для дощок заднього боку на захід.
EXOD|26|28|А середній засув посередині дощок буде засувати від кінця до кінця.
EXOD|26|29|А ці дошки пообкладаєш золотом, а каблучки їхні, на вкладання для засувів, поробиш із золота; і ці засуви пообкладаєш золотом.
EXOD|26|30|І поставиш скинію згідно з приписами, як тобі показано на горі.
EXOD|26|31|І зробиш завісу з блакиті, і пурпуру, і червені та з суканого віссону. Мистецькою роботою зробити її з херувимами.
EXOD|26|32|І повісь її на чотирьох акаційних стовпах, пообкладаних золотом, гаки їх золоті, на чотирьох срібних підставах.
EXOD|26|33|І повісь ту завісу під гачками, і внесеш туди за завісу ковчега свідоцтва. І ця завіса буде відділяти вам між святинею й між Святеє Святих!
EXOD|26|34|І покладеш те віко на ковчега свідоцтва в Святому Святих.
EXOD|26|35|І поставиш стола назовні завіси, а свічника навпроти столу на боці скинії на південь, а стола поставиш на боці півночі.
EXOD|26|36|І зробиш заслону входу скинії з блакиті, і пурпуру, і червені та з суканого віссону, робота гаптівника.
EXOD|26|37|І зробиш для заслони п'ять акаційних стовпів, і пообкладаєш їх золотом; гаки їх золото; і виллєш для них п'ять мідяних підстав.
EXOD|27|1|І зробиш жертівника з акаційного дерева, п'ять ліктів довжина, і п'ять ліктів ширина; квадратовий нехай буде той жертівник, а вишина його три лікті.
EXOD|27|2|І поробиш роги його на чотирьох кутах його, із нього нехай будуть роги його. І пообкладаєш його міддю.
EXOD|27|3|І поробиш горшки на зсипування попелу з нього, і лопатки його, і кропильниці його, і видельця його, і його лопатки на вугіль. Для всього посуду його будеш уживати міді.
EXOD|27|4|І зробиш для нього мідяну мережу роботою сітки, а над мережею зробиш чотири мідяні каблучки на чотирьох кінцях його.
EXOD|27|5|І покладеш її здолу під лиштву жертівника, і буде та мережа аж до половини жертівника.
EXOD|27|6|І поробиш держаки для жертівника, держаки з акаційного дерева, і пообкладаєш їх міддю.
EXOD|27|7|І буде всунено держаки його в каблучки; і будуть ті держаки на двох боках жертівника при ношенні його.
EXOD|27|8|Порожнявим усередині зробиш його з дощок. Як показано було тобі на горі, так нехай зроблять.
EXOD|27|9|І зробиш скинійне подвір'я. На південну сторону, на полудень запони для подвір'я, суканий віссон; довжина першій стороні сто літків.
EXOD|27|10|А стовпів для нього двадцять, а їхніх підстав із міді двадцять. Гаки тих стовпів та обручі їхні срібло.
EXOD|27|11|І так само на сторону півночі вдовжину запони: довжина сто ліктів; а стовпів для нього двадцять, а підстав для них двадцять, із міді. Гаки тих стовпів та обручі їхні срібло.
EXOD|27|12|А ширина подвір'я в сторону заходу: запони п'ятдесят ліктів, а для них стовпів десять, а їхніх підстав десять.
EXOD|27|13|А ширина подвір'я в сторону переду, сходу, п'ятдесят ліктів.
EXOD|27|14|І на п'ятнадцять ліктів запони для боку; стовпів для них три, і підстав для них три.
EXOD|27|15|А для боку другого п'ятнадцять ліктів запони; стовпів для них три, і підстав для них три.
EXOD|27|16|А для брами подвір'я заслона на двадцять ліктів із блакиті, і пурпуру, і червені та з суканого віссону, робота гаптівника. Для них стовпів чотири, і підстав їхніх чотири.
EXOD|27|17|Усі стовпи подвір'я поспинані навколо сріблом; їхні гаки срібло, а підстави їхні мідь.
EXOD|27|18|Довжина подвір'я сто ліктів, а ширина скрізь п'ятдесят, а вишина п'ять ліктів. Запони з суканого віссону, а підстави стовпів мідь.
EXOD|27|19|Усі речі скинії для всякої служби в ній, усі кілки її й усі кілки подвір'я мідь.
EXOD|27|20|І ти накажеш Ізраїлевим синам, і нехай вони приносять тобі оливу з оливок, чисту, товчену, для освітлення, щоб завжди горіла лямпада.
EXOD|27|21|У скинії заповіту назовні завіси, що на свідоцтві, приготує її на запалення Аарон та сини його від вечора аж до ранку перед лицем Господнім. Це вічна постанова їхнім родам від Ізраїлевих синів!
EXOD|28|1|А ти візьми до себе брата свого Аарона та синів його з ним, з-поміж Ізраїлевих синів, щоб він був священиком для Мене, Аарона, Надава, і Авігу, Елеазара та Ітамара, синів Ааронових.
EXOD|28|2|І зробиш священні шати для брата свого Аарона на славу й красу.
EXOD|28|3|І ти скажеш усім мудросердим, що Я наповнив їх духом мудрости, і вони зроблять Ааронові шати для посвячення його, щоб був священиком для Мене.
EXOD|28|4|А оце ті шати, що вони зроблять: нагрудник, і ефод, і верхню шату, і хітон плетений, завій і пояс. І зробиш священні шати для брата свого Аарона та для синів його, щоб він був священиком для Мене.
EXOD|28|5|І візьмуть вони золота, і блакиті, і пурпуру, і червені та віссону,
EXOD|28|6|і зроблять ефода з золота, блакиті, і пурпуру, і червені та з віссону суканого, робота мистця.
EXOD|28|7|Два злучені нараменники будуть у нього при обох кінцях його, і буде він сполучений.
EXOD|28|8|А пояс мистецький його ефоду, що на нім, тієї ж роботи, нехай буде з нього, з золота, блакиті, і пурпуру, і червені та з суканого віссону.
EXOD|28|9|І візьмеш два оніксові камені, та й вирізьбиш на них імена Ізраїлевих синів,
EXOD|28|10|шість із їхніх імен на камені однім, а ймення шости позосталих на камені другім, за їхнім народженням.
EXOD|28|11|Роботою різьбаря каменя, різьбою печатки вирізьбиш на тих обох каменях імена Ізраїлевих синів; оточені золотими гніздами зробиш їх.
EXOD|28|12|І положиш обидва камені на нараменниках ефоду, камені пам'яти для Ізраїлевих синів. І буде носити Аарон їхні ймення перед Божим лицем на обох плечах своїх на пам'ять.
EXOD|28|13|А гнізда поробиш із золота.
EXOD|28|14|І два ланцюги зо щирого золота, плетеними поробиш їх, роботою шнурів. І даси ті плетені ланцюги на гнізда.
EXOD|28|15|І зробиш нагрудника судного, роботою мистця, як робота ефоду зробиш його, із золота, блакиті, і пурпуру, і червені та з віссону суканого зробиш його.
EXOD|28|16|Квадратовий нехай буде він, зложений удвоє, п'ядь довжина його, і п'ядь ширина його.
EXOD|28|17|І понасаджуєш на ньому каменеве насадження, чотири ряди каменя. Ряд: рубін, топаз і смарагд ряд перший.
EXOD|28|18|А ряд другий: карбункул, сапфір і яспіс.
EXOD|28|19|А ряд третій: опаль, агат і аметист.
EXOD|28|20|А четвертий ряд: хризоліт, і онікс, і берил, вони будуть вставлені в золото в своїх гніздах.
EXOD|28|21|А камені нехай будуть на ймення дванадцяти Ізраїлевих синів, на ймення їх; різьбою печатки кожен на ймення його нехай будуть для дванадцяти родів.
EXOD|28|22|І поробиш на нагруднику сукані ланцюги плетеною роботою зо щирого золота.
EXOD|28|23|І зробиш на нагруднику дві золоті каблучки, і даси ці дві каблучки на двох кінцях нагрудника.
EXOD|28|24|І даси два золоті шнури на дві ті каблучки до кінців нагрудника.
EXOD|28|25|А два кінці двох шнурів даси до двох гнізд, і даси на нараменники ефоду спереду його.
EXOD|28|26|І зробиш дві золоті каблучки, і покладеш їх на двох кінцях нагрудника на краї його, що до сторони ефоду, всередину.
EXOD|28|27|І зробиш дві золоті каблучки, та й даси їх на обидва нараменники ефоду здолу, спереду його, при сполученні його, над мистецьким поясом ефоду.
EXOD|28|28|І прив'яжуть нагрудника від каблучок його до каблучок ефоду блакитною ниткою, щоб був на мистецькім поясі ефоду, і не буде рухатись нагрудник із-над ефоду.
EXOD|28|29|І буде носити Аарон імена Ізраїлевих синів в суднім нагруднику на серці своїм, як буде входити до святині, на повсякчасну пам'ять перед Господнім лицем.
EXOD|28|30|І даси до судного нагрудника урім та туммім, і будуть вони на Аароновім серці при вході його перед Господнє лице. І буде завжди носити Аарон суд Ізраїлевих синів на своїм серці перед Господнім обличчям.
EXOD|28|31|І зробиш верхню шату для ефоду, усю блакитну.
EXOD|28|32|І нехай буде в середині її отвір для голови його; край отвору нехай буде навколо роботою ткача, як панцерний отвір буде їй, щоб їй не дертися.
EXOD|28|33|І поробиш на подолку її гранатові яблука з блакиті, і пурпуру та з червені, на подолку її навколо, і золоті дзвінки поміж ними навколо,
EXOD|28|34|золотий дзвінок і гранатове яблуко, золотий дзвінок і гранатове яблуко на подолку тієї шати навколо.
EXOD|28|35|І нехай вона буде на Ааронові для служення, і нехай буде чутий голос його при вході його до святині перед Господнє обличчя, і при виході його, щоб йому не померти.
EXOD|28|36|І зробиш квітку зо щирого золота, і вирізьбиш на ній, як різьба печатки: Святиня для Господа.
EXOD|28|37|І покладеш її на нитці з блакиті, і нехай вона буде на завої, на переді завою нехай буде вона.
EXOD|28|38|І нехай буде вона на Аароновім чолі, і нехай носить Аарон гріх тієї святощі, що Ізраїлеві сини посвятять її для всіх своїх святих дарунків. І нехай вона буде завжди на його чолі на благовоління для них перед Господнім лицем.
EXOD|28|39|І витчеш хітона з віссону, і зробиш завоя з віссону, і зробиш пояса роботою гаптяра.
EXOD|28|40|І для синів Ааронових поробиш хітони, і поробиш їм пояси, і поробиш їм покриття голови на славу й красу.
EXOD|28|41|І понадягаєш їх на брата свого Аарона та на синів його з ним. І помажеш їх, і рукоположиш їх, і посвятиш їх, і будуть вони священиками Мені.
EXOD|28|42|І пороби їм льняну спідню одіж, щоб закрити тілесну наготу, від стегон аж до голінок нехай будуть вони.
EXOD|28|43|І нехай будуть вони на Ааронові та на синах його при вході їх до скинії заповіту, або при приході їх до жертівника на служення в святині, і не понесуть вони гріха, і не помруть. Це вічна постанова йому та нащадками його по ньому!
EXOD|29|1|А оце та річ, яку ти зробиш їм для посвячення їх, щоб вони були священиками Мені. Візьми одного бичка молодого та два безвадні барани,
EXOD|29|2|і прісний хліб, і прісні калачі, змішані з оливою, і прісні коржі, помазані оливою, із ліпшої пшеничної муки поробиш їх.
EXOD|29|3|І покладеш їх до одного коша, і принесеш їх у коші, і того бичка та два ті барани.
EXOD|29|4|А Аарона та синів його приведи до входу скинії умовлення, і обмиєш їх водою.
EXOD|29|5|І візьмеш шати та й убереш Аарона в хітона, і в ефодну шату, і в ефода, і в нагрудника, і опережеш його мистецьким поясом ефоду.
EXOD|29|6|І наложиш завоя на його голову, а на завій даси вінця святости.
EXOD|29|7|І візьмеш оливу помазання, і виллєш йому на голову, та й помажеш його.
EXOD|29|8|І приведеш синів його, та й повбираєш їх у хітони.
EXOD|29|9|І попідперізуєш їх поясом, Аарона та синів його, і наложиш їм покриття голови, і буде для них священство на вічну постанову. І рукоположиш Аарона та синів його.
EXOD|29|10|І приведеш бичка до скинії заповіту, і покладе Аарон та сини його руки свої на голову того бичка.
EXOD|29|11|І заріжеш того бичка перед Господнім обличчям при вході до скинії заповіту.
EXOD|29|12|І візьмеш крови бичка, і помажеш на рогах жертівника пальцем своїм, а всю кров виллєш до основи жертівника.
EXOD|29|13|І візьмеш увесь лій, що покриває нутро, і сальника на печінці, і обидві нирки та лій, що на них, та й спалиш на жертівнику.
EXOD|29|14|А м'ясо бичка, і шкуру його та нечистоти його спалиш в огні поза табором, це жертва за гріх.
EXOD|29|15|І візьмеш одного барана, і нехай покладуть Аарон та сини його свої руки на голову того барана.
EXOD|29|16|І заріжеш того барана, і візьмеш кров його, та й покропиш жертівника навколо.
EXOD|29|17|А того барана порозтинаєш на куски його, і виполощеш нутрощі його та голінки його, і покладеш на куски його та на голову його.
EXOD|29|18|І спалиш усього барана на жертівнику, це цілопалення для Господа, пахощі любі, огняна жертва, для Господа вона.
EXOD|29|19|І візьмеш другого барана, і покладе Аарон та сини його руки свої на голову того барана.
EXOD|29|20|І заріжеш того барана, і візьмеш крови його, та й даси на пипку Ааронового вуха, і на пипку правого вуха синів його, і на великий палець правої руки їхньої, і на великий палець їхньої правої ноги. І покропиш ту кров на жертівника навколо.
EXOD|29|21|І візьмеш із крови, що на жертівнику, і з оливи помазання, та й покропиш на Аарона й на шати його, та на синів його й на шати синів його з ним. І освятиться він, і шати його та сини й шати синів його з ним!
EXOD|29|22|І візьмеш із того барана лій та курдюка, і лій, що покриває нутрощі, і сальника на печінці, й обидві нирки, і лій, що на них, і праве стегно, бо це баран посвячення.
EXOD|29|23|І один буханець хліба, і один хлібний оливний калач, і один коржик із коша з прісним, що перед лицем Господнім.
EXOD|29|24|І покладеш усе те на руку Аарона й на руки синів його, і поколихаєш його, як колихання перед Господнім лицем.
EXOD|29|25|І візьмеш його з їхньої руки, та й спалиш на жертівнику на цілопалення, на пахощі любі перед Господнім лицем, це огняна жертва для Господа.
EXOD|29|26|І візьмеш грудину з барана посвячення, що Ааронів, і поколихаєш її, як колихання перед Господнім лицем, і це буде твоя частина.
EXOD|29|27|І посвятиш грудину колихання та стегно приношення, що були колихані, і що було принесене з барана рукоположення, з того, що Ааронове, і з того, що синів його.
EXOD|29|28|І буде це Ааронові та синам його на вічну постанову від Ізраїлевих синів, бо це приношення. І буде воно приношенням від Ізраїлевих синів і мирних їхніх жертов, їхнє приношення для Господа.
EXOD|29|29|А священні шати, що Ааронові, будуть по ньому синам його на помазання в них і на рукоположення їх.
EXOD|29|30|Сім день носитиме їх той із синів його, що буде священиком замість нього, що ввійде до скинії заповіту на служення в святині.
EXOD|29|31|І візьмеш барана посвячення, і звариш м'ясо його в святім місці.
EXOD|29|32|І буде їсти Аарон та сини його м'ясо того барана, та той хліб, що в коші, при вході до скинії заповіту.
EXOD|29|33|І поїдять вони те, чим окуплено їх на рукоположення їх, на посвячення їх. А чужий не буде їсти, бо святість воно!
EXOD|29|34|А якщо позостанеться з м'яса посвячення та з того хліба до ранку, то спалиш позостале в огні, не буде те їджене, бо святість воно!
EXOD|29|35|І зробиш Ааронові та синам його так, як усе, що Я наказав був тобі. Сім день будеш посвячувати їх.
EXOD|29|36|А бичка, жертву за гріх, будеш споряджати щоденно для окуплення. І будеш очищати жертівника, коли будеш чинити окуплення його. І помажеш його на його посвячення.
EXOD|29|37|Сім день будеш складати окупа на жертівнику й освятиш його, і стане той жертівник найсвятішим. Усе, що доторкнеться до жертівника, освятиться.
EXOD|29|38|А оце те, що будеш споряджати на жертівнику: ягнята, однорічного віку, двоє на день завжди.
EXOD|29|39|Одне ягня спорядиш уранці, а друге ягня спорядиш під вечір.
EXOD|29|40|І десятину ефи пшеничної муки, мішаної в товченій оливі, чверть гіну, і на лиття чверть гіну вина на одне ягня.
EXOD|29|41|А ягня друге спорядиш під вечір; як хлібну жертву ранку й як жертву плинну її спорядиш йому, на пахощі любі, огняна жертва для Господа,
EXOD|29|42|стале цілопалення для ваших поколінь при вході до скинії заповіту перед Господнім лицем, що буду там відкриватися вам, щоб говорити до тебе там.
EXOD|29|43|І буду відкриватися там Ізраїлевим синам, і це місце буде освячене Моєю славою.
EXOD|29|44|І освячу скинію заповіту, і жертівника, і Аарона та синів його освячу, щоб вони були священиками Мені.
EXOD|29|45|І буду Я спочивати серед Ізраїлевих синів, і буду їм Богом.
EXOD|29|46|І познають вони, що Я Господь, їхній Бог, що вивів їх із єгипетського краю, щоб перебувати Мені серед них. Я Господь, їхній Бог!
EXOD|30|1|І зробиш жертівника на кадіння кадила, з акаційного дерева зробиш його.
EXOD|30|2|Лікоть довжина його, і лікоть ширина його, квадратовий нехай буде він, а два лікті вишина його. З нього виходитимуть роги його.
EXOD|30|3|І пообкладаєш його щирим золотом, дах його та стіни його навколо, та роги його. І зробиш йому вінця золотого навколо.
EXOD|30|4|І дві золоті каблучки зробиш йому під вінця його, на двох боках його зробиш, на двох сторонах, і буде це на вкладання для держаків, щоб ними носити його.
EXOD|30|5|І поробиш держаки з акаційного дерева, і пообкладаєш їх золотом.
EXOD|30|6|І поставиш його перед завісою, що над ковчегом свідоцтва, перед віком, що на свідоцтві, яким Я буду тобі відкриватися там.
EXOD|30|7|І буде Аарон кадити на ньому кадило пахощів щоранку, коли він поправлятиме лямпадки, то буде кадити його.
EXOD|30|8|І при запаленні лямпадок під вечір він буде кадити його. Це постійне кадило перед Господнім лицем на ваші покоління!
EXOD|30|9|Не запалите на ньому чужого кадила, ані цілопалення, ані жертви хлібної, і жертви рідинної не будете лити на ньому.
EXOD|30|10|І складе Аарон окупа на роги його, раз у році, з крови жертви за гріх раз у році дня Окуплення складе він окупа на нього на ваші покоління. Це найсвятіше для Господа!
EXOD|30|11|І промовив Господь до Мойсея, говорячи:
EXOD|30|12|Коли будеш робити перелік Ізраїлевих синів за тими, кого повинно лічити, то дадуть вони кожен викупа за душу свою Господеві при переліку їх, і не буде між ними моровиці при переліку їх.
EXOD|30|13|Оце дасть кожен, що переходить на переліку: половину шекля, на міру шеклем святині, двадцять ґер той шекель; половина цього шекля приношення для Господа.
EXOD|30|14|Кожен, хто переходить на переліку, від віку двадцяти літ і вище, дасть приношення для Господа.
EXOD|30|15|Багатий не побільшить, а вбогий не зменшить від половини шекля, даючи приношення Господеві для складання окупу за ваші душі.
EXOD|30|16|І візьмеш гроші окупу від Ізраїлевих синів, та й даси їх на роботу скинії заповіту. І буде воно Ізраїлевим синам на пам'ять перед Господнім обличчям для окуплення за ваші душі.
EXOD|30|17|І Господь промовляв до Мойсея, говорячи:
EXOD|30|18|І зробиш умивальницю з міді, і підстава її мідь, на вмивання. І поставиш її між скинією заповіту й між жертівником, і наллєш туди води.
EXOD|30|19|І будуть Аарон та сини його мити з неї свої руки та ноги свої.
EXOD|30|20|Коли вони входитимуть до скинії заповіту, то будуть мити в воді, щоб їм не вмерти, або коли будуть відходити до жертівника на служення, щоб спалити огняну жертву для Господа.
EXOD|30|21|І будуть вони вмивати руки свої та ноги свої, щоб їм не вмерти. І буде це для них вічна постанова, для нього й для нащадків його на їхні покоління!
EXOD|30|22|І Господь промовляв до Мойсея, говорячи:
EXOD|30|23|А ти візьми собі найкращих пахощів: самотечної мірри п'ять сотень шеклів, і запашного цинамону половину його: двісті й п'ятдесят, і запашної очеретини двісті й п'ятдесят,
EXOD|30|24|і касії п'ять сотень шеклів на міру шеклем святині, та гін оливкової оливи.
EXOD|30|25|І зробиш її миром святого помазання, масть складену, робота робітника масти. Це буде миро святого помазання.
EXOD|30|26|І намастиш ним скинію заповіту, і ковчега свідоцтва,
EXOD|30|27|і стола та всі речі його, і свічника та речі його, і жертівника кадила,
EXOD|30|28|і жертівника цілопалення та всі речі його, і вмивальницю та підставу її.
EXOD|30|29|І освятиш їх, і стануть вони найсвятішим, усе, що доторкнеться до них, освятиться!
EXOD|30|30|І помажеш Аарона та синів його, та посвятиш їх на священнослуження Мені.
EXOD|30|31|А до синів Ізраїлевих будеш говорити, кажучи: Це буде Мені миро святого помазання на ваші покоління.
EXOD|30|32|На людське тіло не буде воно лите, і за постановою про нього не буде робитися, як воно, святиня воно, воно буде святиня для вас!
EXOD|30|33|Кожен, хто сам робитиме масть, як воно, і хто дасть із нього на чужого, той буде витятий із народу свого.
EXOD|30|34|І промовив Господь до Мойсея: Візьми собі пахощів: бальзаму, і ониху, і хелбану, пахощів, та чистого ладану, кожне буде в рівній частині.
EXOD|30|35|І зробиш з цього кадило, масть, робота робітника масти, посолене, чисте, святе.
EXOD|30|36|І зітреш із неї надрібно, і даси з неї перед обличчям свідоцтва в скинії заповіту, що Я буду являтися тобі там, це буде найсвятіше для вас!
EXOD|30|37|А кадило, що зробите, за постановою про нього це зробите собі, воно буде тобі святість для Господа!
EXOD|30|38|Кожен, хто зробить, як воно, щоб нюхати з нього, той буде витятий із народу свого!
EXOD|31|1|І промовив Господь до Мойсея, говорячи:
EXOD|31|2|Дивися, Я покликав на ім'я Бецал'їла, сина Урієвого, сина Хура, Юдиного племени,
EXOD|31|3|і наповнив його Духом Божим, мудрістю, і розумуванням, і знанням, і здібністю до всякої роботи,
EXOD|31|4|на обмислення мистецьке, на роботу в золоті, і в сріблі, і в міді,
EXOD|31|5|і в обробленні каменя, щоб всаджувати, і в обробленні дерева, щоб робити в усякій роботі.
EXOD|31|6|І Я ото дав із ним Оголіява, Ахісамахового сина, Данового племени. А в серце кожного мудросердого Я дав мудрість, і зроблять вони все, що Я наказав був тобі:
EXOD|31|7|скинію заповіту, і ковчега для свідоцтва, і віко, що на ньому, і всі скинійні речі,
EXOD|31|8|і стола та речі його, і чистого свічника та всі речі його, і жертівника кадила,
EXOD|31|9|і жертівника цілопалення та всі речі його, і вмивальницю та підставу її,
EXOD|31|10|і шати служебні, і шати священні для священика Аарона, і шати синів його на священнослуження,
EXOD|31|11|і оливу помазання, і запашне кадило для святині, як усе, що Я наказав був тобі, вони зроблять.
EXOD|31|12|І промовив Господь до Мойсея, говорячи:
EXOD|31|13|А ти промовляй Ізраїлевим синам, говорячи: Тільки суботи Мої будете пильнувати, бо це знак поміж Мною та поміж вами для ваших поколінь, щоб ви познали, що Я Господь, що освячує вас!
EXOD|31|14|І будете пильнувати суботу, бо вона святість для вас. Хто опоганить її, той конче буде забитий, бо кожен, хто робить у ній роботу, то буде стята душа та з-посеред народів її!
EXOD|31|15|Шість день буде робитися праця, а дня сьомого субота відпочинку від праці, святість для Господа. Кожен, хто робить роботу за суботнього дня, той конче буде забитий!
EXOD|31|16|І будуть Ізраїлеві сини додержувати суботу, щоб зробити суботу вічним заповітом для своїх поколінь.
EXOD|31|17|Це знак навіки поміж Мною та поміж Ізраїлевими синами, бо шість день творив Господь небо та землю, а дня сьомого перервав працю та спочив.
EXOD|31|18|І дав Він Мойсеєві, коли закінчив говорити з ним на Сінайській горі, дві таблиці свідоцтва, таблиці кам'яні, писані Божим перстом.
EXOD|32|1|І побачив народ, що загаявся Мойсей зійти з гори. І зібрався народ проти Аарона, та й сказали до нього: Устань, зроби нам богів, що будуть ходити перед нами, бо той Мойсей, муж, що вивів був нас із єгипетського краю, ми не знаємо, що сталось йому.
EXOD|32|2|І сказав їм Аарон: Поздіймайте золоті сережки, що в ушах ваших жінок, ваших синів та дочок ваших, і поприносьте до мене.
EXOD|32|3|І ввесь народ поздіймав з себе золоті сережки, що в їхніх ушах, та й позносили до Аарона.
EXOD|32|4|І взяв він це з їхньої руки, і вформував його в глині, і зробив із нього лите теля. А вони сказали: Оце твої боги, Ізраїлю, що вивели тебе з єгипетського краю!
EXOD|32|5|І побачив це Аарон, і збудував жертівника перед ним. І кликнув Аарон та й сказав: Завтра свято для Господа!
EXOD|32|6|І повставали вони взавтра рано вранці, і принесли цілопалення, і привели мирну жертву. І засів народ до їди та до пиття, і встали бавитися.
EXOD|32|7|А Господь промовляв до Мойсея: Іди, зійди, бо зіпсувся народ твій, якого ти вивів із єгипетського краю.
EXOD|32|8|Зійшли вони скоро з дороги, що наказав був Я їм, зробили собі лите теля, і поклонились йому, і склали йому жертви, та й сказали: Оце твої боги, Ізраїлю, що вивели тебе з єгипетського краю!
EXOD|32|9|І промовив Господь до Мойсея: Я бачив народ той, і ось народ твердошиїй він!
EXOD|32|10|А тепер залиши Мене, і розпалиться гнів Мій на них, і Я винищу їх, а тебе зроблю великим народом.
EXOD|32|11|І Мойсей став благати лице Господа, Бога свого, та й сказав: Нащо, Господи, розпалюється гнів Твій на народ Твій, якого Ти випровадив з єгипетського краю силою великою та міцною рукою?
EXOD|32|12|Нащо будуть казати єгиптяни, говорячи: На зле ти їх вивів, щоб їх повбивати в горах, та щоб винищити їх з-поверхні землі?... Вернися з розпалу гніву Свого, та й відверни зло від Свого народу!
EXOD|32|13|Згадай про Авраама, Ісака та Ізраїля, рабів Своїх, що Ти їм присягався був Собою, та говорив їм: Помножу ваших нащадків, немов зорі небесні, і всю оту землю, що про неї казав, дам вашим нащадкам, і вони посядуть навіки.
EXOD|32|14|І відвернув Господь зло, про яке говорив, щоб зробити Своєму народові.
EXOD|32|15|І повернувся, і зійшов Мойсей із гори, а в руці його дві таблиці свідоцтва, писані з обох їхніх сторін, звідси й звідти вони були писані.
EXOD|32|16|А таблиці Божа робота вони, а письмо Боже письмо воно, вирізьблене на таблицях.
EXOD|32|17|І почув Ісус голос народу, як кричав він, та й сказав до Мойсея: Крик бою в таборі!
EXOD|32|18|А той відказав: Це не крик сили переможців і не крик слабости переможених, я чую голос співу!
EXOD|32|19|І сталося, коли він наблизився до табору, то побачив теля те та танці... І розпалився гнів Мойсеїв, і він кинув таблиці із рук своїх, та й розторощив їх під горою!...
EXOD|32|20|І схопив він теля, що зробили вони, та й спалив на огні, та змолов, аж став порох... І розсипав на поверхні води, і напоїв тим синів Ізраїлевих.
EXOD|32|21|І сказав Мойсей Ааронові: Що вчинив тобі народ цей, що ти гріх великий навів на нього?
EXOD|32|22|А Аарон відказав: Нехай не запалиться гнів мого пана! Ти знаєш народ цей, що він у злому.
EXOD|32|23|І вони сказали мені: Зроби нам богів, що будуть ходити перед нами, бо той Мойсей, муж, що вивів нас із єгипетського краю, ми не знаємо, що сталось йому.
EXOD|32|24|І сказав я до них: Хто має золото, поздіймайте з себе. І дали вони мені, а я кинув його в огонь, і вийшло те теля.
EXOD|32|25|І побачив Мойсей народ, що незагнузданий він, бо Аарон розгнуздав його на ганьбу поміж їхніми ворогами.
EXOD|32|26|І став Мойсей у брамі табору й сказав: Хто за Господа до мене! І зібралися до нього всі Левіїні сини.
EXOD|32|27|І сказав він до них: Так сказав Господь, Бог Ізраїлів: Припашіть кожен меча свого на стегно своє, перейдіть, і верніться від брами до брами в таборі, і повбивайте кожен брата свого, і кожен приятеля свого, і кожен ближнього свого.
EXOD|32|28|І зробили Левіїні сини за словом Мойсеєвим. І впало з народу того дня близько трьох тисяч чоловіка.
EXOD|32|29|І сказав Мойсей: Освятіть сьогодні себе для Господа, бо кожен мстився на сині своїм та на браті своїм, і щоб сьогодні Він дав вам благословення.
EXOD|32|30|І сталося назавтра, і сказав Мойсей до народу: Ви згрішили великим гріхом, а тепер зійду я до Господа, може складу окуплення за ваш гріх.
EXOD|32|31|І вернувся Мойсей до Господа та й сказав: О, згрішив цей народ великим гріхом, вони зробили собі золотих богів!
EXOD|32|32|А тепер, коли б Ти пробачив їм їхній гріх! А як ні, витри мене з книги Своєї, яку Ти написав...
EXOD|32|33|І промовив Господь до Мойсея: Хто згрішив Мені, того витру із книги Своєї.
EXOD|32|34|А тепер іди, провадь цей народ туди, куди казав Я тобі. Ось Мій Ангол піде перед лицем твоїм. А в день кари Моєї покараю їх за їхній гріх!
EXOD|32|35|І Господь ударив той народ за те, що вони зробили теля, яке Аарон учинив був.
EXOD|33|1|І говорив Господь до Мойсея: Іди, вийди звідси ти та той народ, що ти вивів його з єгипетського краю до того Краю, що Я присяг був його Авраамові, Ісакові та Якову, говорячи: Нащадкам твоїм дам його,
EXOD|33|2|і пошлю перед лицем твоїм Ангола, і попроганяю ханаанеянина, амореянина, і хіттеянина, і періззеянина, хіввеянина, і євусеянина,
EXOD|33|3|до Краю, що тече молоком та медом, бо Я не піду серед тебе, бо ти народ твердошиїй, щоб Я не вигубив тебе в дорозі.
EXOD|33|4|І почув народ ту лиху вістку, та й засмутився, і ніхто не поклав на себе своєї оздоби.
EXOD|33|5|Бо промовив Господь до Мойсея: Скажи Ізраїлевим синам: Ви народ твердошиїй, якщо одну хвилину піду серед тебе, то вигублю тебе! Тож тепер здійми оздобу свою з себе, Я знатиму, що вчиню тобі.
EXOD|33|6|І поздіймали Ізраїлеві сини свої оздоби під горою Хорив.
EXOD|33|7|А Мойсей узяв намета, та й нап'яв його поза табором, далеко від табору, і назвав його: скинія заповіту. І бувало, кожен, хто шукав Господа, входив до скинії заповіту, що поза табором.
EXOD|33|8|І бувало, коли виходив Мойсей до скинії, то підводився ввесь народ, і ставали кожен при вході свого намету, і дивилися за Мойсеєм, аж поки він не входив до скинії.
EXOD|33|9|І бувало, коли входив Мойсей до скинії, то сходив стовп хмари, і ставав при вході скинії, та й говорив Бог із Мойсеєм.
EXOD|33|10|І ввесь народ бачив стовпа хмари, що стояв при вході скинії. І ввесь народ підводився, та й вклонялися, кожен при вході намету свого.
EXOD|33|11|І говорив Господь до Мойсея лице в лице, як говорить хто до друга свого. І вертався він до табору, а слуга його, юнак Ісус, син Навинів, не виходив із середини скинії.
EXOD|33|12|І сказав Мойсей до Господа: Дивися, Ти говориш мені: Випровади цей народ, а Ти не дав мені знати, кого зо мною пошлеш. А Ти сказав був: Я знаю тебе на ім'я, а також знайшов ти милість в очах Моїх.
EXOD|33|13|Тож тепер, коли знайшов я милість в очах Твоїх, об'яви ж мені дорогу Свою, і я пізнаю, як знайти милість в очах Твоїх. І побач, бо цей люд то народ Твій.
EXOD|33|14|А Він відказав: Сам Я піду, і введу тебе до відпочинку.
EXOD|33|15|І сказав він до Нього: Коли сам Ти не підеш, то не виводь нас ізвідси.
EXOD|33|16|Бож чим тоді пізнається, що знайшов милість в очах Твоїх я та народ Твій? Чи ж не тим, що Ти підеш із нами? І будемо вирізнені я та народ Твій від кожного народу, що на поверхні землі.
EXOD|33|17|І промовив Господь до Мойсея: Також цю річ, про яку говорив ти, зроблю, бо ти знайшов милість в очах Моїх, і Я знаю на ім'я тебе.
EXOD|33|18|А він відказав: Покажи мені славу Свою!
EXOD|33|19|І Він промовив: Я переведу все добро Своє перед тобою, і покличу Господнім Ім'ям перед тобою. І Я помилую, до кого милостивий, і змилосерджуся, до кого милосердний.
EXOD|33|20|І Він промовив: Ти не зможеш побачити лиця Мого, бо людина не може побачити Мене і жити.
EXOD|33|21|І промовив Господь: Ось місце при Мені, і ти станеш на скелі.
EXOD|33|22|І станеться, коли буде переходити слава Моя, то Я вміщу Тебе в щілині скелі, і закрию тебе рукою Своєю, аж поки Я перейду.
EXOD|33|23|А здійму руку Свою, і ти побачиш Мене ззаду, а обличчя Моє не буде видиме.
EXOD|34|1|І промовив Господь до Мойсея: Витеши собі дві кам'яні таблиці, як перші, і Я напишу на цих таблицях слова, що були на перших таблицях, які ти розбив.
EXOD|34|2|І приготовся на рано. І вийдеш рано вранці на гору Сінай, і станеш Мені там на верхів'ї гори.
EXOD|34|3|А з тобою ніхто не вийде, і на всій горі нехай нікого не буде видно. І також дрібна худоба й худоба велика нехай не пасеться навпроти тієї гори.
EXOD|34|4|І витесав він дві кам'яні таблиці, як перші. І встав Мойсей рано вранці, та й вийшов на гору Сінай, як Господь звелів був йому. І взяв він у руку свою дві таблиці кам'яні.
EXOD|34|5|А Господь зійшов у хмарі, і став там із ним, та й покликав Ім'ям Господа.
EXOD|34|6|І перейшов Господь перед лицем його, та й викликнув: Господь, Господь, Бог милосердний, і милостивий, довготерпеливий, і многомилостивий та правдивий,
EXOD|34|7|що дотримує милість для тисяч, що вибачає провину й переступ та гріх, та певне не вважає чистим винуватого, бо карає провину батьків на дітях, і на дітях дітей, і на третіх, і на четвертих поколіннях.
EXOD|34|8|І Мойсей поквапно вклонився до землі, і впав,
EXOD|34|9|та й сказав: Якщо я знайшов милість в очах Твоїх, Владико, то нехай же Владика йде серед нас, бо народ цей твердошиїй. І Ти пробачиш нашу провину та наш гріх, і зробиш нас спадком Своїм.
EXOD|34|10|А Він відказав: Ось Я складаю заповіта перед усім народом твоїм. Я чинитиму чуда, які не були творені на всій землі і в жодного народу. І побачить увесь народ, серед якого ти знаходишся, чин Господній, що Я чиню його з тобою, який він страшний!
EXOD|34|11|Виконуй те, що Я наказую тобі сьогодні. Ось Я виганяю перед тобою амореянина, і ханаанеянина, і хіттеянина, і періззеянина, і хіввеянина, і євусеянина.
EXOD|34|12|Стережися, щоб не склав ти умови з мешканцем тієї землі, що ти входиш на неї, щоб він не став пасткою серед тебе.
EXOD|34|13|Бо ви їхні жертівники поруйнуєте, а їхні камінні стовпи для богів поторощите, а їхні дерева святі повирубуєте.
EXOD|34|14|Бо не будеш ти кланятись богові іншому, бо Господь Заздрісний ім'я Його, Бог заздрісний Він!
EXOD|34|15|Щоб не склав ти умови з мешканцем Краю, як будуть вони любодіяти вслід за богами своїми, і будуть богам своїм жертви приносити, то якщо він покличе тебе, то ти не будеш їсти із жертви його.
EXOD|34|16|І не візьмеш із дочок його для синів своїх, бо будуть вони любодіяти вслід за богами своїми, і вчинять розпусниками синів твоїх вслід за богами своїми.
EXOD|34|17|Литих богів не зробиш собі.
EXOD|34|18|Будеш виконувати свято Опрісноків. Сім день будеш їсти опрісноки, що Я наказав був тобі на умовлений час місяця авіва, бо в місяці авіві ти вийшов з Єгипту.
EXOD|34|19|Усе, що відкриває утробу то Моє, як і всяка твоя худоба, що є самець, відкриття утроби вола та вівці.
EXOD|34|20|А відкриття утроби осла викупиш ягням. А якщо його не викупиш, то заб'єш його, зламавши шию. Кожного перворідного з синів твоїх викупиш. І не будуть являтися перед обличчя Моє з порожньою рукою.
EXOD|34|21|Шість день будеш працювати, а дня сьомого спочинеш від праці; в орці й у жнива спочинеш від праці.
EXOD|34|22|І свято тижнів зробиш собі, і первоплоду жнив пшениці, і свято збору врожаю під кінець року.
EXOD|34|23|Тричі в році вся чоловіча стать буде являтися перед лице Владики Господа, Бога Ізраїлевого.
EXOD|34|24|Бо Я вижену людей перед лицем твоїм, і розширю границю твою, і ніхто не запрагне твоєї землі, коли ти ходитимеш являтися перед лице Господа, Бога твого, тричі в році.
EXOD|34|25|Не будеш приносити на квашенім крови жертви твоєї, і не переночує до рана святкова жертва Пасхи.
EXOD|34|26|Початок первоплодів твоєї землі принесеш у дім Господа, Бога твого. Не будеш варити ягняти в молоці його матері.
EXOD|34|27|І промовив Господь до Мойсея: Напиши собі слова, бо згідно з цими словами склав Я заповіта з тобою та з Ізраїлем.
EXOD|34|28|І був він там з Господом сорок день і сорок ночей, хліба не їв і води не пив. І написав на таблицях слова Заповіту, Десять Заповідей.
EXOD|34|29|І сталося, коли сходив Мойсей з гори Сінай, а обидві таблиці свідоцтва в Мойсеєвій руці при сході його з гори, що Мойсей не знав, що лице його стало променіти, бо Бог говорив з ним.
EXOD|34|30|І побачив Аарон та всі Ізраїлеві сини Мойсея, аж ось лице його променіло, і вони боялися підійти до нього!
EXOD|34|31|І кликнув до них Мойсей, і звернулися до нього Аарон та всі начальники в громаді. І Мойсей говорив до них.
EXOD|34|32|А потім попідходили всі Ізраїлеві сини, і він наказав їм усе, що Господь говорив з ним на горі Сінай.
EXOD|34|33|І скінчив Мойсей говорити з ними, і дав на лице своє покривало.
EXOD|34|34|А коли Мойсей входив перед Господнє лице на розмову з Ним, то здіймав покривало аж до свого виходу. І він виходив, і говорив до Ізраїлевих синів, що було наказано йому.
EXOD|34|35|І бачили Ізраїлеві сини лице Мойсеєве, що променіло лице Мойсеєве. І Мойсей знов накладав покривало на лице своє аж до відходу свого, щоб говорити з Ним.
EXOD|35|1|І зібрав Мойсей усю громаду Ізраїлевих синів, та й промовив до них: Ось ті речі, що Господь наказав їх чинити.
EXOD|35|2|Шість день буде робитися праця, а дня сьомого буде вам свято, субота спочинку від праці для Господа. Кожен, хто робитиме працю в нім, буде забитий!
EXOD|35|3|Не розпалите огню за суботнього дня по всіх ваших осадах.
EXOD|35|4|І сказав Мойсей до всієї громади Ізраїлевих синів, кажучи: Оце та річ, що Господь наказав, говорячи:
EXOD|35|5|Візьміть від себе приношення для Господа. Кожен за щедрим серцем своїм принесе його, приношення Господеві: золото, і срібло, і мідь,
EXOD|35|6|і блакить, і пурпур, і червень, і віссон, і вовну козину,
EXOD|35|7|і начервоно пофарбовані баранячі шкурки, і шкурки тахашеві, і акаційні дерева,
EXOD|35|8|і оливу на освітлення, і пахощі на оливу помазання, та пахощів на кадило,
EXOD|35|9|і каміння оніксове, і каміння на оправу до ефоду й до нагрудника.
EXOD|35|10|А кожен із вас мудросердий прийде та зробить, що наказав був Господь:
EXOD|35|11|скинію внутрішню та її намета зовнішнього, і покриття її, і гачки її, і дошки її, засуви її, стовпи її та підстави її;
EXOD|35|12|ковчега, і держаки його, віко й завісу заслони;
EXOD|35|13|стола, і держаки його, і всі речі його, і хліб показний;
EXOD|35|14|і свічника освітлення, і речі його, і лямпадки його, і оливу освітлення;
EXOD|35|15|і жертівника кадила, і держаки його, і оливу помазання, і кадило пахощів та заслону входу при вході;
EXOD|35|16|жертівника цілопалення, і мідяну його сітку, держаки його, і всі речі його, умивальницю й підставу її;
EXOD|35|17|запони подвір'я, стовпи його, і підстави його та заслону брами подвір'я;
EXOD|35|18|кілки скинії, і кілки подвір'я та шнури їхні;
EXOD|35|19|і шати служебні на служення в святині, священні шати для священика Аарона, та шати синів його на священнослуження.
EXOD|35|20|І вийшла вся громада Ізраїлевих синів від Мойсея.
EXOD|35|21|І приходили кожен чоловік, кого вело серце його, і кожен, кого дух його чинив щедрим, і приносили приношення Господеві для роботи скинії заповіту, і на кожну працю його, і на священні шати.
EXOD|35|22|І приходили ті чоловіки з жінками, кожен щедросердий, і приносили гачка, і носову сережку, і персня, і сережку, всякі золоті речі, та все, що людина приносила, як золото приношення для Господа.
EXOD|35|23|І кожна людина принесла, що хто мав: блакить, і пурпур, і червень, і віссон, і вовна козина, і баранячі начервоно пофарбовані шкурки, і шкурки тахашеві.
EXOD|35|24|Кожен, хто жертвував срібне та мідяне приношення, приносив Господнє приношення, і кожен, хто мав, поприносили акаційне дерево, на всяке зайняття коло тієї роботи.
EXOD|35|25|І кожна мудросерда жінка пряла руками своїми, і приносила пряжку: блакить, і пурпур, і червень, і віссон.
EXOD|35|26|І всі жінки, кого вело їхнє серце, пряли козину вовну.
EXOD|35|27|А начальники поприносили каміння оніксу, і каміння вставлення для ефоду та для нагрудника,
EXOD|35|28|і пахощі, і оливу на освітлення, і для оливи помазання, і для запашного кадила.
EXOD|35|29|Кожен чоловік та жінка, кого їхнє серце схиляло приносити для кожної праці, яку Господь наказав робити рукою Мойсея, Ізраїлеві сини приносили добровільний дар для Господа.
EXOD|35|30|І сказав Мойсей до Ізраїлевих синів: Дивіться, Господь назвав на ім'я Бецал'їла, сина Урієвого, сина Хура, Юдиного роду.
EXOD|35|31|І наповнив його Духом Божим, мудрістю, розумуванням, і знанням, і здібністю до всякої роботи
EXOD|35|32|на обмислення мистецьке, на роботу в золоті, і в сріблі, і в міді,
EXOD|35|33|і в обробленні каменя, щоб всаджувати, і в обробленні дерева, щоб робити в усякій мистецькій роботі.
EXOD|35|34|І вклав в його серце, щоб навчав, він і Оголіяв, син Ахісамаха, Данового племени.
EXOD|35|35|Він наповнив їх мудрістю серця, щоб робили вони всяку роботу обрібника, і мистця, і гаптівника в блакиті, і в пурпурі, і в червені, і в віссоні, і ткача, що роблять усяку роботу й задумують мистецькі речі.
EXOD|36|1|І зробить Бецал'їл та Оголіяв, та кожен мудросердий чоловік, кому Господь дав мудрости та розсудку, щоб уміти зробити кожну працю роботи в святині на все, що Господь наказав був.
EXOD|36|2|І покликав Мойсей Бецал'їла та Оголіява, та кожного мудросердого чоловіка, кому Господь подав мудрість у серце, кожного, кого вело серце зблизитися до тієї праці, щоб зробити її.
EXOD|36|3|І взяли вони від Мойсея все приношення, що позносили Ізраїлеві сини для праці служби святині, щоб зробити її. А вони ще приносили до нього щоранку добровільного дара.
EXOD|36|4|І прибули всі мудреці, що роблять усю роботу святині, кожен із праці своєї, яку вони роблять,
EXOD|36|5|і сказали до Мойсея, говорячи: Народ приносить більше, ніж потрібно було для праці, яку Господь звелів був зробити.
EXOD|36|6|І Мойсей наказав проголосити в таборі, говорячи: Ні чоловік, ні жінка нехай не роблять уже нічого на приношення для святині. І був стриманий народ від приносів.
EXOD|36|7|А наготовленого було досить для кожної праці, щоб зробити її, і ще зоставалось.
EXOD|36|8|І зробили кожен мудросердий із тих, що робили скинійну працю: десять покривал із суканого віссону, і блакиті, і пурпуру та з червені. Херувими мистецькою роботою він поробив їх.
EXOD|36|9|Довжина одного покривала двадцять і вісім ліктів, а ширина одного покривала чотири лікті. Усім покривалам міра одна.
EXOD|36|10|І поспинав він п'ять покривал одне до одного, і п'ять інших покривал поспинав одне до одного.
EXOD|36|11|І поробив він блакитні петельки на краю одного покривала з кінця в спинанні. Так само зробив на краю кінцевого покривала в спинанні другім.
EXOD|36|12|П'ятдесят петельок зробив він у покривалі однім, і п'ятдесят петельок зробив він на кінці покривала, що в другім спинанні. Ті петельки протилеглі одна до однієї.
EXOD|36|13|І зробив він п'ятдесят золотих гачків, і поспинав ті покривала одне до одного тими гачками, і стала одна скинія.
EXOD|36|14|І зробив він покривала з вовни козиної до намета над внутрішньою скинією, одинадцять покривал зробив таких.
EXOD|36|15|Довжина одного покривала тридцять ліктів, а ширина одного покривала чотири лікті. Одинадцятьом покривалам міра одна.
EXOD|36|16|І поспинав він п'ять покривал осібно, а шість тих покривал осібно.
EXOD|36|17|І поробив він п'ятдесят петельок на краю кінцевого покривала в спинанні, і п'ятдесят петельок поробив на краю покривала другого спинання.
EXOD|36|18|І зробив він п'ятдесят мідяних гачків на спинання скинії, щоб стала вона одна.
EXOD|36|19|І зробив він накриття для скинії, баранячі начервоно пофарбовані шкурки, і накриття зверху з тахашевих шкурок.
EXOD|36|20|І поробив він для скинії стоячі дошки з акаційного дерева.
EXOD|36|21|Десять ліктів довжина дошки, і лікоть і півліктя ширина однієї дошки.
EXOD|36|22|В одній дошці дві ручки, сполучені одна до однієї. Так він поробив усі дошки скинії.
EXOD|36|23|І поробив він дошки для скинії, двадцять дощок на бік південний, на полудень.
EXOD|36|24|І сорок срібних підстав поробив він під тими двадцятьма дошками, дві підставі під однією дошкою для ручок її, і дві підставі під дошкою другою для двох ручок її.
EXOD|36|25|А для другого боку скинії, у бік півночі зробив він двадцять дощок.
EXOD|36|26|І для них сорок срібних підстав, дві підставі під одну дошку, і дві підставі під дошку другу.
EXOD|36|27|А для заднього боку скинії на захід зробив він шість дощок.
EXOD|36|28|І дві дошки зробив він для скинійних кутів на заднього бока.
EXOD|36|29|І були вони поєднані здолу, і разом були вони поєднані на верху її до однієї каблучки. Так зробив він для них обох, для обох кутів.
EXOD|36|30|І було вісім дощок, а їхні підстави зо срібла, шістнадцять підстав: по дві підставі під одну дошку.
EXOD|36|31|І зробив він засуви з акаційного дерева, п'ять для дощок одного боку скинії,
EXOD|36|32|і п'ять засувів для дощок другого боку скинії, і п'ять засувів для дощок заднього боку на захід.
EXOD|36|33|І зробив він середнього засува, щоб засувати по середині дощок від кінця до кінця.
EXOD|36|34|А ці дошки він пообкладав золотом, а каблучки їхні, на вкладання для засувів, поробив із золота; і ці засуви він пообкладав золотом.
EXOD|36|35|І зробив він завісу з блакиті, і пурпуру, і червені та з суканого віссону. Мистецькою роботою зробив її з херувимами.
EXOD|36|36|І він зробив для неї чотири акаційні стовпи, і пообкладав їх золотом, гаки їх золоті, і вилив для них чотири срібних підставі.
EXOD|36|37|І зробив він заслону для входу скинії з блакиті, і пурпуру, і червені та з суканого віссону, робота гаптівника.
EXOD|36|38|А стовпи її п'ять, а гаки їх золоті; і він пообкладав їх верхи та їх обручі золотом; а підстави їхні п'ять із міді.
EXOD|37|1|І зробив Бецал'їл ковчега з акаційного дерева, два лікті й пів довжина його, і лікоть і пів ширина його, і лікоть і пів вишина його.
EXOD|37|2|І пообкладав він його щирим золотом зсередини та іззовні. І вінця золотого зробив навколо над ним.
EXOD|37|3|І він вилив для нього чотири золоті каблучки на чотирьох кутах його, дві каблучки на одному боці його, і дві каблучки на другому боці його.
EXOD|37|4|І він поробив держаки з акаційного дерева, і пообкладав їх золотом.
EXOD|37|5|І він повсовував ці держаки в каблучки на боках ковчегу, щоб носити ковчега.
EXOD|37|6|І віко зробив зо щирого золота, два лікті й пів довжина його, і лікоть і пів ширина його.
EXOD|37|7|І зробив два золоті херувими, роботою кутою зробив їх з обох кінців віка.
EXOD|37|8|І зробив одного херувима з кінця звідти, а одного херувима з кінця звідси. З того віка поробив тих херувимів на обох кінцях його.
EXOD|37|9|І були ті херувими з простягненими догори крилами, і затінювали своїми крилами над віком, а їхні лиця одне до одного; до віка були схилені лиця тих херувимів.
EXOD|37|10|І зробив він стола з акаційного дерева, два лікті довжина його, і лікоть ширина його, і лікоть і пів вишина його.
EXOD|37|11|І пообкладав його щирим золотом, і зробив вінця золотого для нього навколо.
EXOD|37|12|І лиштву зробив він для нього в долоню навколо, і зробив вінця золотого навколо для лиштви його.
EXOD|37|13|І він вилив для нього чотири каблучки із золота, та й дав ті каблучки на чотирьох кінцях, що при його чотирьох ніжках.
EXOD|37|14|При лиштві були ті каблучки, вкладання для держаків, щоб носити стола.
EXOD|37|15|І поробив він ті держаки з акаційного дерева, і пообкладав їх золотом, щоб носити стола.
EXOD|37|16|І поробив він ті речі, що на столі: миски його, і кадильниці його, і кухлі його та чаші його, що ними лито, золото щире.
EXOD|37|17|І зробив він свічника зо щирого золота, роботою кутою зробив він того свічника. Стовп його, і рамена його, келихи його, ґудзі його й квіти його виходили з нього.
EXOD|37|18|І шість рамен виходило з боків його, три рамені свічника з одного боку його, і три рамені свічника з другого боку його.
EXOD|37|19|Три келихи мигдалоподібні в однім рамені, ґудзь і квітка, і три мигдалоподібні келихи в рамені другім, ґудзь і квітка. Так на шости раменах, що виходять із свічника.
EXOD|37|20|А на стовпі свічника чотири келихи мигдалоподібні, ґудзі його та квітки його.
EXOD|37|21|І ґудзь під двома раменами з нього, і ґудзь під другими двома раменами з нього, і ґудзь під третіми двома раменами з нього, у шости рамен, що виходять із свічника.
EXOD|37|22|Їхні ґудзі та їхні рамена виходили з нього. Увесь він одне куття щирого золота.
EXOD|37|23|І зробив він сім лямпадок до нього; а його щипчики та його лопатки на вугіль зо щирого золота.
EXOD|37|24|З таланту щирого золота зробив він його та всі його речі.
EXOD|37|25|І зробив він кадильного жертівника з акаційного дерева, лікоть довжина його, і лікоть ширина його, квадратовий, а два лікті вишина його. З нього були його роги.
EXOD|37|26|І пообкладав він його щирим золотом, верх його та стіни його навколо, та роги його. І вінця золотого навколо зробив.
EXOD|37|27|І дві золоті каблучки зробив йому під вінця його, зробив на обох боках його, на вкладання для держаків, щоб ними носити його.
EXOD|37|28|І держаки поробив із акаційного дерева, і золотом пообкладав їх.
EXOD|37|29|І зробив він миро святого помазання, і чисте кадило пахощів, робота робітника масти.
EXOD|38|1|І зробив він жертівника з акаційного дерева, п'ять ліктів довжина його, і п'ять ліктів ширина його, квадратовий, а вишина його три лікті.
EXOD|38|2|І поробив він роги його на чотирьох кутах його, з нього були його роги. І пообкладав його міддю.
EXOD|38|3|І він поробив усі речі жертівника: горшки, і шуфлі, і кропильниці, видельця, і лопатки на вугілля. Усі речі його поробив він із міді.
EXOD|38|4|І мережу зробив він із міді для жертівника роботою сітки, під лиштву його здолу до половини його.
EXOD|38|5|І вилив він чотири каблучки на чотирьох кінцях його для мідяної мережі, на вкладання для держаків.
EXOD|38|6|І поробив він держаки з акаційного дерева, і пообкладав їх міддю.
EXOD|38|7|І повсовував він ті держаки в каблучки на боках жертівника, щоб ними носити його. Порожнявим усередині зробив його з дощок.
EXOD|38|8|І зробив він умивальницю з міді та підставу її з міді, з дзеркалами жінок, що сповняли службу при вході скинії заповіту.
EXOD|38|9|І зробив він подвір'я. На південну сторону, на полудень запони того подвір'я, суканий віссон, сто ліктів.
EXOD|38|10|А стовпів для нього двадцять, а їхніх підстав із міді двадцять. Гаки тих стовпів та обручі їхні срібло.
EXOD|38|11|А в сторону півночі сто ліктів; стовпів для них двадцять і підстав для них двадцять, із міді. Гаки тих стовпів та обручі їхні срібло.
EXOD|38|12|А в сторону заходу, запони, п'ятдесят ліктів; стовпів для них десять, і підстав для них десять. Гаки тих стовпів та обручі їхні срібло.
EXOD|38|13|А в сторону переду, сходу, п'ятдесят ліктів.
EXOD|38|14|Запони до боку п'ятнадцять ліктів; стовпів для них три, і підстав для них три.
EXOD|38|15|А для другого боку з цієї й з тієї сторони брами подвір'я запони на п'ятнадцять ліктів; стовпів для них три, і підстав для них три.
EXOD|38|16|Всі запони подвір'я навколо віссон суканий.
EXOD|38|17|А підстави для стовпів мідь, гаки стовпів та обручів їхніх срібло. А обклад верхів їх срібло, і вони всі стовпи подвір'я поспинані сріблом.
EXOD|38|18|А заслона брами подвір'я робота гаптівника: блакить, і пурпур, і червень та суканий віссон; і двадцять ліктів довжина, а вишина в ширині п'ять ліктів, відповідно запонам подвір'я.
EXOD|38|19|А стовпів для них чотири, і підстав для них чотири, із міді. Гаки їх срібло, і обклад верхів їх та їхніх обручів срібло.
EXOD|38|20|А всі кілки для скинії й для подвір'я навколо мідь.
EXOD|38|21|Оце перелік скинії, скинії свідоцтва, що був обрахований на приказ Мойсея, за допомогою Левитів під рукою Ітамара, сина Аарона, священика.
EXOD|38|22|А Бецал'їл, син Урія, сина Хура, Юдиного племени, поробив усе, що Господь наказав був Мойсеєві.
EXOD|38|23|А з ним Оголіяв, син Ахісамахів, Данового племени, оброблювач, і мистець, і гаптівник блакиттю, і пурпуром, і червенню, і віссоном.
EXOD|38|24|Усе золото, вжите для праці в усій роботі святині, то було золото колихання, двадцять і п'ять талантів та сім сотень і тридцять шеклів на міру шеклем святині.
EXOD|38|25|А срібло полічених у громаді мужів сто талантів та тисяча, і сімсот і сімдесят і п'ять шеклів на міру шеклем святині,
EXOD|38|26|на голову бека, цебто половина шекля на міру шеклем святині для кожного, хто переходив при переліку від віку двадцяти літ і вище, для шостисот тисяч і трьох тисяч і п'ятисот і п'ятидесяти.
EXOD|38|27|І було сто талантів срібла на відлиття підстав святині та підстав завіси, сотня підстав на сотню талантів, талант на підставу.
EXOD|38|28|А з тисячі й семисот і семидесяти й п'яти шеклів поробив він гаки для стовпів, і пообкладав їхні верхи та поспинав їх.
EXOD|38|29|А міді колихання було сімдесят талантів та дві тисячі й чотириста шеклів.
EXOD|38|30|І поробив він із неї підстави входу скинії заповіту, і жертівника мідяного, і його мідяну мережу, та всі речі жертівника,
EXOD|38|31|і підстави подвір'я навколо, і підстави брами подвір'я, і скинійні кілки, і всі кілки подвір'я навколо.
EXOD|39|1|А з блакиті й пурпуру та червені поробили вони службові шати для служення в святині. І поробили священні шати, що вони для Аарона, як Господь наказав був Мойсеєві.
EXOD|39|2|І зробив він ефода з золота, блакиті, і пурпуру, і червені та з суканого віссону.
EXOD|39|3|І повибивали вони золоті бляхи, та й настригли ниток на роботу серед блакиті, і серед пурпуру, і серед червені, і серед віссону, робота мистця.
EXOD|39|4|Вони зробили для нього злучені нараменники, на обох кінцях його він був сполучений.
EXOD|39|5|А пояс мистецький для накладання ефоду, що з ним з'єднаний і однакового з ним виробу, золото, блакить, і пурпур, і червень, і суканий віссон, як Господь наказав був Мойсеєві.
EXOD|39|6|І поробили вони камені оніксові, оточені золотими гніздами, вирізьблені різьбою печатки, з іменами Ізраїлевих синів.
EXOD|39|7|І він їх поклав на ефодові нараменники, камені на пам'ять для Ізраїлевих синів, як Господь наказав був Мойсеєві.
EXOD|39|8|І зробив він нагрудника, роботою мистця, як робота ефоду, золото, блакить, і пурпур, і червень, і суканий віссон.
EXOD|39|9|Квадратовий він був, складеним удвоє зробили нагрудника, п'ядь ширина його, складений удвоє.
EXOD|39|10|І понасаджували на ньому чотири ряди каменя. Ряд: рубін, топаз і смарагд ряд перший.
EXOD|39|11|А ряд другий: карбункул, сапфір і яспіс.
EXOD|39|12|А ряд третій: опаль, агат і аметист.
EXOD|39|13|А четвертий ряд: хризоліт, онікс і беріл, вони вставлені золотими насадами в своїх гніздах.
EXOD|39|14|А камені ті на ймення дванадцятьох Ізраїлевих синів вони, на ймення їх; різьбою печатки кожен на ім'я його для дванадцяти племен.
EXOD|39|15|І поробили вони на нагруднику сукані ланцюги плетеною роботою зо щирого золота.
EXOD|39|16|І зробили вони дві золоті гнізді та дві золоті каблучки, і дали ці каблучки на двох кінцях нагрудника.
EXOD|39|17|І дали два золоті шнури на дві ті каблучки до кінців нагрудника.
EXOD|39|18|А два кінці обох шнурів дали до двох гнізд, і дали на нараменники ефоду спереду його.
EXOD|39|19|І зробили дві золоті каблучки, та й поклали на обох кінцях нагрудника на краї його, що до сторони ефоду, всередину.
EXOD|39|20|І зробили вони дві золоті каблучки, та й дали їх на обидва нараменники ефоду здолу, спереду його, при сполученні його, над мистецьким поясом ефоду.
EXOD|39|21|І прив'язали нагрудника від каблучок його до каблучок ефоду блакитною ниткою, щоб був на мистецькім поясі ефоду, і не буде рухатись нагрудник із-над ефоду, як Господь наказав був Мойсеєві.
EXOD|39|22|І зробив він шату для ефоду, ткацькою роботою, всю блакитну.
EXOD|39|23|А отвір шати в середині її, як отвір панцера; край отвору її обрамований навколо, щоб не дертися їй.
EXOD|39|24|І поробили вони на подолку шати гранатові яблука з блакиті, і пурпуру та з суканої червені.
EXOD|39|25|І поробили дзвінки зо щирого золота, і дали ті дзвінки поміж гранатові яблука на подолку шати навколо, поміж ті гранатові яблука,
EXOD|39|26|дзвінок і гранатове яблуко, дзвінок і гранатове яблуко на подолку шати тієї навколо, на служення, як Господь наказав був Мойсеєві.
EXOD|39|27|І поробили вони хітони з віссону, робота ткача, для Аарона та для синів його,
EXOD|39|28|і завоя з віссону, і шапки накриття з віссону, і льняна спідня одіж із суканого віссону,
EXOD|39|29|і пояса з суканого віссону, і блакиті, і пурпура та з червені, робота гаптяра, як Господь наказав був Мойсеєві.
EXOD|39|30|І зробили квітку, вінця святости, зо щирого золота, і написали на нім письмом різьби печатки: Святиня для Господа.
EXOD|39|31|І дали на нім блакитну нитку, щоб була на завої згори, як Господь наказав був Мойсеєві.
EXOD|39|32|І скінчилася вся робота скинії, скинії заповіту. І зробили Ізраїлеві сини все, як Господь наказав був Мойсеєві, так зробили вони.
EXOD|39|33|І позносили вони до Мойсея скинію внутрішню, намета зовнішнього та всі речі її: гачки її, дошки її, засуви її, і стовпи її та підстави її,
EXOD|39|34|і накриття з баранячих начервоно пофарбованих шкурок, і накриття з тахашевих шкурок, і завісу заслони,
EXOD|39|35|ковчега свідоцтва, і держаки його, і віко,
EXOD|39|36|стола, усі речі його, і хліб показний,
EXOD|39|37|чистого свічника та лямпадки його, лямпадки розставлені, та всі речі його й оливу освітлення,
EXOD|39|38|і золотого жертівника, миро помазання, і запашне кадило, і завісу при вході скинії,
EXOD|39|39|мідяного жертівника, і його мідяну мережку, держаки його, і всі речі його, умивальницю та підставу її,
EXOD|39|40|запони подвір'я, стовпи його, і підстави його, і заслону для брами подвір'я, шнури його, і кілки його, і всі речі для служби в скинії, у скинії заповіту,
EXOD|39|41|службові шати для служення в святині, священні шати священика Аарона, і шати синів його для священнослуження.
EXOD|39|42|Усе так, як Господь наказав був Мойсеєві, так зробили Ізраїлеві сини всю ту роботу.
EXOD|39|43|І побачив Мойсей усю ту роботу, і ось вони зробили її! Як Господь наказав був, так зробили вони. І поблагословив їх Мойсей!
EXOD|40|1|А Господь промовляв до Мойсея, говорячи:
EXOD|40|2|Першого місяця, першого дня місяця поставиш намета для скинії заповіту.
EXOD|40|3|І поставиш там ковчега свідоцтва, і закриєш ковчега завісою.
EXOD|40|4|І внесеш стола, і порозкладаєш належне йому; і внесеш свічника, і запалиш його лямпадки.
EXOD|40|5|І поставиш золотого жертівника для кадила перед ковчегом свідоцтва; і повісиш заслону входу скинії.
EXOD|40|6|І поставиш жертівника цілопалення перед входом скинії, скинії заповіту.
EXOD|40|7|І поставиш умивальницю між скинією заповіту та між жертівником, і даси туди води.
EXOD|40|8|І поставиш подвір'я навколо, і даси заслону брами подвір'я.
EXOD|40|9|І візьмеш миро помазання, та й помажеш скинію та все, що в ній, і освятиш її та всі речі її, і стане вона святістю.
EXOD|40|10|І помажеш жертівника цілопалення та всі речі його, і освятиш жертівника, і стане жертівник Найсвятішим.
EXOD|40|11|І помажеш умивальницю та підставу її, і освятиш її.
EXOD|40|12|І приведеш Аарона та синів його до входу скинії заповіту, та й обмиєш їх водою.
EXOD|40|13|І зодягнеш Аарона в священні шати, і помажеш його, і освятиш його, і він буде священнослужити Мені.
EXOD|40|14|І приведеш синів його, і позодягаєш їх у хітони.
EXOD|40|15|І помажеш їх, як помазав їхнього батька, і будуть вони священнослужити Мені. І станеться, що помазання їх буде на них на вічне священство, на їхні покоління!
EXOD|40|16|І зробив Мойсей усе, як Господь наказав був йому, так він зробив.
EXOD|40|17|І сталося першого місяця другого року, першого дня місяця, була поставлена скинія!
EXOD|40|18|І поставив Мойсей скинію, і дав підстави її, і поклав дошки її, і дав засови її, і поставив стовпи її.
EXOD|40|19|І розтягнув намета над внутрішньою скинією, і поклав скинійне накриття на неї згори, як Господь наказав був Мойсеєві.
EXOD|40|20|І взяв він і поклав свідоцтво до ковчега, а на ковчега поклав держаки, і дав на ковчега віко згори.
EXOD|40|21|І вніс він ковчега до скинії, і повісив завісу заслони, і закрив ковчег свідоцтва, як Господь наказав був Мойсеєві.
EXOD|40|22|І дав він стола в скинію заповіту, на стороні скинії на північ, поза завісою.
EXOD|40|23|І порозкладав на ньому розклад хліба перед Господнім лицем, як Господь наказав був Мойсеєві.
EXOD|40|24|І поставив свічника в скинії заповіту навпроти стола, на стороні скинії на південь.
EXOD|40|25|І позасвічував лямпадки перед Господнім лицем, як Господь наказав був Мойсеєві.
EXOD|40|26|І поставив золотого жертівника в скинії заповіту перед завісою.
EXOD|40|27|І кадив він на ньому запашні кадила, як Господь наказав був Мойсеєві.
EXOD|40|28|І повісив входову заслону до скинії.
EXOD|40|29|А жертівника цілопалення поставив при вході скинії, скинії заповіту, і приніс на ньому цілопалення та жертву хлібну, як Господь наказав був Мойсеєві.
EXOD|40|30|І поставив умивальницю між скинією заповіту та між жертівником, і туди дав води на миття.
EXOD|40|31|І вмивали з нього Мойсей й Аарон та сини його руки свої та ноги свої.
EXOD|40|32|Коли вони входили до скинії заповіту, і коли зближалися до жертівника, вони обмивалися, як Господь наказав був Мойсеєві.
EXOD|40|33|І поставив подвір'я навколо скинії та жертівника, і повісив заслону брами подвір'я.
EXOD|40|34|А хмара закрила скинію заповіту, і слава Господня наповнила скинію.
EXOD|40|35|І не міг Мойсей увійти до скинії заповіту, бо хмара спочивала над нею, а слава Господня наповнила скинію.
EXOD|40|36|А коли підіймалася хмара з-над скинії, то Ізраїлеві сини рушали в усі свої подорожі.
EXOD|40|37|А якщо хмара не підіймалася, то не рушали вони аж до дня, коли вона підіймалася,
EXOD|40|38|бо над скинією вдень була хмара Господня, а вночі був огонь у ній, на очах усього Ізраїлевого дому в усіх його подорожах!
