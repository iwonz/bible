PROV|1|1|Притчи Соломона, сына Давидова, царя Израильского,
PROV|1|2|чтобы познать мудрость и наставление, понять изречения разума;
PROV|1|3|усвоить правила благоразумия, правосудия, суда и правоты;
PROV|1|4|простым дать смышленость, юноше – знание и рассудительность;
PROV|1|5|послушает мудрый – и умножит познания, и разумный найдет мудрые советы;
PROV|1|6|чтобы разуметь притчу и замысловатую речь, слова мудрецов и загадки их.
PROV|1|7|Начало мудрости – страх Господень; глупцы только презирают мудрость и наставление.
PROV|1|8|Слушай, сын мой, наставление отца твоего и не отвергай завета матери твоей,
PROV|1|9|потому что это – прекрасный венок для головы твоей и украшение для шеи твоей.
PROV|1|10|Сын мой! если будут склонять тебя грешники, не соглашайся;
PROV|1|11|если будут говорить: "иди с нами, сделаем засаду для убийства, подстережем непорочного без вины,
PROV|1|12|живых проглотим их, как преисподняя, и – целых, как нисходящих в могилу;
PROV|1|13|наберем всякого драгоценного имущества, наполним домы наши добычею;
PROV|1|14|жребий твой ты будешь бросать вместе с нами, склад один будет у всех нас", –
PROV|1|15|сын мой! не ходи в путь с ними, удержи ногу твою от стези их,
PROV|1|16|потому что ноги их бегут ко злу и спешат на пролитие крови.
PROV|1|17|В глазах всех птиц напрасно расставляется сеть,
PROV|1|18|а делают засаду для их крови и подстерегают их души.
PROV|1|19|Таковы пути всякого, кто алчет чужого добра: оно отнимает жизнь у завладевшего им.
PROV|1|20|Премудрость возглашает на улице, на площадях возвышает голос свой,
PROV|1|21|в главных местах собраний проповедует, при входах в городские ворота говорит речь свою:
PROV|1|22|"доколе, невежды, будете любить невежество? [доколе] буйные будут услаждаться буйством? доколе глупцы будут ненавидеть знание?
PROV|1|23|Обратитесь к моему обличению: вот, я изолью на вас дух мой, возвещу вам слова мои.
PROV|1|24|Я звала, и вы не послушались; простирала руку мою, и не было внимающего;
PROV|1|25|и вы отвергли все мои советы, и обличений моих не приняли.
PROV|1|26|За то и я посмеюсь вашей погибели; порадуюсь, когда придет на вас ужас;
PROV|1|27|когда придет на вас ужас, как буря, и беда, как вихрь, принесется на вас; когда постигнет вас скорбь и теснота.
PROV|1|28|Тогда будут звать меня, и я не услышу; с утра будут искать меня, и не найдут меня.
PROV|1|29|За то, что они возненавидели знание и не избрали [для себя] страха Господня,
PROV|1|30|не приняли совета моего, презрели все обличения мои;
PROV|1|31|за то и будут они вкушать от плодов путей своих и насыщаться от помыслов их.
PROV|1|32|Потому что упорство невежд убьет их, и беспечность глупцов погубит их,
PROV|1|33|а слушающий меня будет жить безопасно и спокойно, не страшась зла".
PROV|2|1|Сын мой! если ты примешь слова мои и сохранишь при себе заповеди мои,
PROV|2|2|так что ухо твое сделаешь внимательным к мудрости и наклонишь сердце твое к размышлению;
PROV|2|3|если будешь призывать знание и взывать к разуму;
PROV|2|4|если будешь искать его, как серебра, и отыскивать его, как сокровище,
PROV|2|5|то уразумеешь страх Господень и найдешь познание о Боге.
PROV|2|6|Ибо Господь дает мудрость; из уст Его – знание и разум;
PROV|2|7|Он сохраняет для праведных спасение; Он – щит для ходящих непорочно;
PROV|2|8|Он охраняет пути правды и оберегает стезю святых Своих.
PROV|2|9|Тогда ты уразумеешь правду и правосудие и прямоту, всякую добрую стезю.
PROV|2|10|Когда мудрость войдет в сердце твое, и знание будет приятно душе твоей,
PROV|2|11|тогда рассудительность будет оберегать тебя, разум будет охранять тебя,
PROV|2|12|дабы спасти тебя от пути злого, от человека, говорящего ложь,
PROV|2|13|от тех, которые оставляют стези прямые, чтобы ходить путями тьмы;
PROV|2|14|от тех, которые радуются, делая зло, восхищаются злым развратом,
PROV|2|15|которых пути кривы, и которые блуждают на стезях своих;
PROV|2|16|дабы спасти тебя от жены другого, от чужой, которая умягчает речи свои,
PROV|2|17|которая оставила руководителя юности своей и забыла завет Бога своего.
PROV|2|18|Дом ее ведет к смерти, и стези ее – к мертвецам;
PROV|2|19|никто из вошедших к ней не возвращается и не вступает на путь жизни.
PROV|2|20|Посему ходи путем добрых и держись стезей праведников,
PROV|2|21|потому что праведные будут жить на земле, и непорочные пребудут на ней;
PROV|2|22|а беззаконные будут истреблены с земли, и вероломные искоренены из нее.
PROV|3|1|Сын мой! наставления моего не забывай, и заповеди мои да хранит сердце твое;
PROV|3|2|ибо долготы дней, лет жизни и мира они приложат тебе.
PROV|3|3|Милость и истина да не оставляют тебя: обвяжи ими шею твою, напиши их на скрижали сердца твоего,
PROV|3|4|и обретешь милость и благоволение в очах Бога и людей.
PROV|3|5|Надейся на Господа всем сердцем твоим, и не полагайся на разум твой.
PROV|3|6|Во всех путях твоих познавай Его, и Он направит стези твои.
PROV|3|7|Не будь мудрецом в глазах твоих; бойся Господа и удаляйся от зла:
PROV|3|8|это будет здравием для тела твоего и питанием для костей твоих.
PROV|3|9|Чти Господа от имения твоего и от начатков всех прибытков твоих,
PROV|3|10|и наполнятся житницы твои до избытка, и точила твои будут переливаться новым вином.
PROV|3|11|Наказания Господня, сын мой, не отвергай, и не тяготись обличением Его;
PROV|3|12|ибо кого любит Господь, того наказывает и благоволит к тому, как отец к сыну своему.
PROV|3|13|Блажен человек, который снискал мудрость, и человек, который приобрел разум, –
PROV|3|14|потому что приобретение ее лучше приобретения серебра, и прибыли от нее больше, нежели от золота:
PROV|3|15|она дороже драгоценных камней; и ничто из желаемого тобою не сравнится с нею.
PROV|3|16|Долгоденствие – в правой руке ее, а в левой у нее – богатство и слава;
PROV|3|17|пути ее – пути приятные, и все стези ее – мирные.
PROV|3|18|Она – древо жизни для тех, которые приобретают ее, – и блаженны, которые сохраняют ее!
PROV|3|19|Господь премудростью основал землю, небеса утвердил разумом;
PROV|3|20|Его премудростью разверзлись бездны, и облака кропят росою.
PROV|3|21|Сын мой! не упускай их из глаз твоих; храни здравомыслие и рассудительность,
PROV|3|22|и они будут жизнью для души твоей и украшением для шеи твоей.
PROV|3|23|Тогда безопасно пойдешь по пути твоему, и нога твоя не споткнется.
PROV|3|24|Когда ляжешь спать, – не будешь бояться; и когда уснешь, – сон твой приятен будет.
PROV|3|25|Не убоишься внезапного страха и пагубы от нечестивых, когда она придет;
PROV|3|26|потому что Господь будет упованием твоим и сохранит ногу твою от уловления.
PROV|3|27|Не отказывай в благодеянии нуждающемуся, когда рука твоя в силе сделать его.
PROV|3|28|Не говори другу твоему: "пойди и приди опять, и завтра я дам", когда ты имеешь при себе.
PROV|3|29|Не замышляй против ближнего твоего зла, когда он без опасения живет с тобою.
PROV|3|30|Не ссорься с человеком без причины, когда он не сделал зла тебе.
PROV|3|31|Не соревнуй человеку, поступающему насильственно, и не избирай ни одного из путей его;
PROV|3|32|потому что мерзость пред Господом развратный, а с праведными у Него общение.
PROV|3|33|Проклятие Господне на доме нечестивого, а жилище благочестивых Он благословляет.
PROV|3|34|Если над кощунниками Он посмевается, то смиренным дает благодать.
PROV|3|35|Мудрые наследуют славу, а глупые – бесславие.
PROV|4|1|Слушайте, дети, наставление отца, и внимайте, чтобы научиться разуму,
PROV|4|2|потому что я преподал вам доброе учение. Не оставляйте заповеди моей.
PROV|4|3|Ибо и я был сын у отца моего, нежно любимый и единственный у матери моей,
PROV|4|4|и он учил меня и говорил мне: да удержит сердце твое слова мои; храни заповеди мои, и живи.
PROV|4|5|Приобретай мудрость, приобретай разум: не забывай этого и не уклоняйся от слов уст моих.
PROV|4|6|Не оставляй ее, и она будет охранять тебя; люби ее, и она будет оберегать тебя.
PROV|4|7|Главное – мудрость: приобретай мудрость, и всем имением твоим приобретай разум.
PROV|4|8|Высоко цени ее, и она возвысит тебя; она прославит тебя, если ты прилепишься к ней;
PROV|4|9|возложит на голову твою прекрасный венок, доставит тебе великолепный венец.
PROV|4|10|Слушай, сын мой, и прими слова мои, – и умножатся тебе лета жизни.
PROV|4|11|Я указываю тебе путь мудрости, веду тебя по стезям прямым.
PROV|4|12|Когда пойдешь, не будет стеснен ход твой, и когда побежишь, не споткнешься.
PROV|4|13|Крепко держись наставления, не оставляй, храни его, потому что оно – жизнь твоя.
PROV|4|14|Не вступай на стезю нечестивых и не ходи по пути злых;
PROV|4|15|оставь его, не ходи по нему, уклонись от него и пройди мимо;
PROV|4|16|потому что они не заснут, если не сделают зла; пропадает сон у них, если они не доведут кого до падения;
PROV|4|17|ибо они едят хлеб беззакония и пьют вино хищения.
PROV|4|18|Стезя праведных – как светило лучезарное, которое более и более светлеет до полного дня.
PROV|4|19|Путь же беззаконных – как тьма; они не знают, обо что споткнутся.
PROV|4|20|Сын мой! словам моим внимай, и к речам моим приклони ухо твое;
PROV|4|21|да не отходят они от глаз твоих; храни их внутри сердца твоего:
PROV|4|22|потому что они жизнь для того, кто нашел их, и здравие для всего тела его.
PROV|4|23|Больше всего хранимого храни сердце твое, потому что из него источники жизни.
PROV|4|24|Отвергни от себя лживость уст, и лукавство языка удали от себя.
PROV|4|25|Глаза твои пусть прямо смотрят, и ресницы твои да направлены будут прямо пред тобою.
PROV|4|26|Обдумай стезю для ноги твоей, и все пути твои да будут тверды.
PROV|4|27|Не уклоняйся ни направо, ни налево; удали ногу твою от зла,
PROV|4|28|[потому что пути правые наблюдает Господь, а левые – испорчены.
PROV|4|29|Он же прямыми сделает пути твои, и шествия твои в мире устроит.]
PROV|5|1|Сын мой! внимай мудрости моей, и приклони ухо твое к разуму моему,
PROV|5|2|чтобы соблюсти рассудительность, и чтобы уста твои сохранили знание.
PROV|5|3|ибо мед источают уста чужой жены, и мягче елея речь ее;
PROV|5|4|но последствия от нее горьки, как полынь, остры, как меч обоюдоострый;
PROV|5|5|ноги ее нисходят к смерти, стопы ее достигают преисподней.
PROV|5|6|Если бы ты захотел постигнуть стезю жизни ее, то пути ее непостоянны, и ты не узнаешь их.
PROV|5|7|Итак, дети, слушайте меня и не отступайте от слов уст моих.
PROV|5|8|Держи дальше от нее путь твой и не подходи близко к дверям дома ее,
PROV|5|9|чтобы здоровья твоего не отдать другим и лет твоих мучителю;
PROV|5|10|чтобы не насыщались силою твоею чужие, и труды твои не были для чужого дома.
PROV|5|11|И ты будешь стонать после, когда плоть твоя и тело твое будут истощены, –
PROV|5|12|и скажешь: "зачем я ненавидел наставление, и сердце мое пренебрегало обличением,
PROV|5|13|и я не слушал голоса учителей моих, не приклонял уха моего к наставникам моим:
PROV|5|14|едва не впал я во всякое зло среди собрания и общества!"
PROV|5|15|Пей воду из твоего водоема и текущую из твоего колодезя.
PROV|5|16|Пусть [не] разливаются источники твои по улице, потоки вод – по площадям;
PROV|5|17|пусть они будут принадлежать тебе одному, а не чужим с тобою.
PROV|5|18|Источник твой да будет благословен; и утешайся женою юности твоей,
PROV|5|19|любезною ланью и прекрасною серною: груди ее да упоявают тебя во всякое время, любовью ее услаждайся постоянно.
PROV|5|20|И для чего тебе, сын мой, увлекаться постороннею и обнимать груди чужой?
PROV|5|21|Ибо пред очами Господа пути человека, и Он измеряет все стези его.
PROV|5|22|Беззаконного уловляют собственные беззакония его, и в узах греха своего он содержится:
PROV|5|23|он умирает без наставления, и от множества безумия своего теряется.
PROV|6|1|Сын мой! если ты поручился за ближнего твоего и дал руку твою за другого, –
PROV|6|2|ты опутал себя словами уст твоих, пойман словами уст твоих.
PROV|6|3|Сделай же, сын мой, вот что, и избавь себя, так как ты попался в руки ближнего твоего: пойди, пади к ногам и умоляй ближнего твоего;
PROV|6|4|не давай сна глазам твоим и дремания веждам твоим;
PROV|6|5|спасайся, как серна из руки и как птица из руки птицелова.
PROV|6|6|Пойди к муравью, ленивец, посмотри на действия его, и будь мудрым.
PROV|6|7|Нет у него ни начальника, ни приставника, ни повелителя;
PROV|6|8|но он заготовляет летом хлеб свой, собирает во время жатвы пищу свою.
PROV|6|9|Доколе ты, ленивец, будешь спать? когда ты встанешь от сна твоего?
PROV|6|10|Немного поспишь, немного подремлешь, немного, сложив руки, полежишь:
PROV|6|11|и придет, как прохожий, бедность твоя, и нужда твоя, как разбойник.
PROV|6|12|Человек лукавый, человек нечестивый ходит со лживыми устами,
PROV|6|13|мигает глазами своими, говорит ногами своими, дает знаки пальцами своими;
PROV|6|14|коварство в сердце его: он умышляет зло во всякое время, сеет раздоры.
PROV|6|15|Зато внезапно придет погибель его, вдруг будет разбит – без исцеления.
PROV|6|16|Вот шесть, что ненавидит Господь, даже семь, что мерзость душе Его:
PROV|6|17|глаза гордые, язык лживый и руки, проливающие кровь невинную,
PROV|6|18|сердце, кующее злые замыслы, ноги, быстро бегущие к злодейству,
PROV|6|19|лжесвидетель, наговаривающий ложь и сеющий раздор между братьями.
PROV|6|20|Сын мой! храни заповедь отца твоего и не отвергай наставления матери твоей;
PROV|6|21|навяжи их навсегда на сердце твое, обвяжи ими шею твою.
PROV|6|22|Когда ты пойдешь, они будут руководить тебя; когда ляжешь спать, будут охранять тебя; когда пробудишься, будут беседовать с тобою:
PROV|6|23|ибо заповедь есть светильник, и наставление – свет, и назидательные поучения – путь к жизни,
PROV|6|24|чтобы остерегать тебя от негодной женщины, от льстивого языка чужой.
PROV|6|25|Не пожелай красоты ее в сердце твоем, и да не увлечет она тебя ресницами своими;
PROV|6|26|потому что из–за жены блудной [обнищевают] до куска хлеба, а замужняя жена уловляет дорогую душу.
PROV|6|27|Может ли кто взять себе огонь в пазуху, чтобы не прогорело платье его?
PROV|6|28|Может ли кто ходить по горящим угольям, чтобы не обжечь ног своих?
PROV|6|29|То же бывает и с тем, кто входит к жене ближнего своего: кто прикоснется к ней, не останется без вины.
PROV|6|30|Не спускают вору, если он крадет, чтобы насытить душу свою, когда он голоден;
PROV|6|31|но, будучи пойман, он заплатит всемеро, отдаст все имущество дома своего.
PROV|6|32|Кто же прелюбодействует с женщиною, у того нет ума; тот губит душу свою, кто делает это:
PROV|6|33|побои и позор найдет он, и бесчестие его не изгладится,
PROV|6|34|потому что ревность – ярость мужа, и не пощадит он в день мщения,
PROV|6|35|не примет никакого выкупа и не удовольствуется, сколько бы ты ни умножал даров.
PROV|7|1|Сын мой! храни слова мои и заповеди мои сокрой у себя.
PROV|7|2|Храни заповеди мои и живи, и учение мое, как зрачок глаз твоих.
PROV|7|3|Навяжи их на персты твои, напиши их на скрижали сердца твоего.
PROV|7|4|Скажи мудрости: "Ты сестра моя!" и разум назови родным твоим,
PROV|7|5|чтобы они охраняли тебя от жены другого, от чужой, которая умягчает слова свои.
PROV|7|6|Вот, однажды смотрел я в окно дома моего, сквозь решетку мою,
PROV|7|7|и увидел среди неопытных, заметил между молодыми людьми неразумного юношу,
PROV|7|8|переходившего площадь близ угла ее и шедшего по дороге к дому ее,
PROV|7|9|в сумерки в вечер дня, в ночной темноте и во мраке.
PROV|7|10|И вот – навстречу к нему женщина, в наряде блудницы, с коварным сердцем,
PROV|7|11|шумливая и необузданная; ноги ее не живут в доме ее:
PROV|7|12|то на улице, то на площадях, и у каждого угла строит она ковы.
PROV|7|13|Она схватила его, целовала его, и с бесстыдным лицом говорила ему:
PROV|7|14|"мирная жертва у меня: сегодня я совершила обеты мои;
PROV|7|15|поэтому и вышла навстречу тебе, чтобы отыскать тебя, и – нашла тебя;
PROV|7|16|коврами я убрала постель мою, разноцветными тканями Египетскими;
PROV|7|17|спальню мою надушила смирною, алоем и корицею;
PROV|7|18|зайди, будем упиваться нежностями до утра, насладимся любовью,
PROV|7|19|потому что мужа нет дома: он отправился в дальнюю дорогу;
PROV|7|20|кошелек серебра взял с собою; придет домой ко дню полнолуния".
PROV|7|21|Множеством ласковых слов она увлекла его, мягкостью уст своих овладела им.
PROV|7|22|Тотчас он пошел за нею, как вол идет на убой, и как олень – на выстрел,
PROV|7|23|доколе стрела не пронзит печени его; как птичка кидается в силки, и не знает, что они – на погибель ее.
PROV|7|24|Итак, дети, слушайте меня и внимайте словам уст моих.
PROV|7|25|Да не уклоняется сердце твое на пути ее, не блуждай по стезям ее,
PROV|7|26|потому что многих повергла она ранеными, и много сильных убиты ею:
PROV|7|27|дом ее – пути в преисподнюю, нисходящие во внутренние жилища смерти.
PROV|8|1|Не премудрость ли взывает? и не разум ли возвышает голос свой?
PROV|8|2|Она становится на возвышенных местах, при дороге, на распутиях;
PROV|8|3|она взывает у ворот при входе в город, при входе в двери:
PROV|8|4|"к вам, люди, взываю я, и к сынам человеческим голос мой!
PROV|8|5|Научитесь, неразумные, благоразумию, и глупые – разуму.
PROV|8|6|Слушайте, потому что я буду говорить важное, и изречение уст моих – правда;
PROV|8|7|ибо истину произнесет язык мой, и нечестие – мерзость для уст моих;
PROV|8|8|все слова уст моих справедливы; нет в них коварства и лукавства;
PROV|8|9|все они ясны для разумного и справедливы для приобретших знание.
PROV|8|10|Примите учение мое, а не серебро; лучше знание, нежели отборное золото;
PROV|8|11|потому что мудрость лучше жемчуга, и ничто из желаемого не сравнится с нею.
PROV|8|12|Я, премудрость, обитаю с разумом и ищу рассудительного знания.
PROV|8|13|Страх Господень – ненавидеть зло; гордость и высокомерие и злой путь и коварные уста я ненавижу.
PROV|8|14|У меня совет и правда; я разум, у меня сила.
PROV|8|15|Мною цари царствуют и повелители узаконяют правду;
PROV|8|16|мною начальствуют начальники и вельможи и все судьи земли.
PROV|8|17|Любящих меня я люблю, и ищущие меня найдут меня;
PROV|8|18|богатство и слава у меня, сокровище непогибающее и правда;
PROV|8|19|плоды мои лучше золота, и золота самого чистого, и пользы от меня больше, нежели от отборного серебра.
PROV|8|20|Я хожу по пути правды, по стезям правосудия,
PROV|8|21|чтобы доставить любящим меня существенное благо, и сокровищницы их я наполняю.
PROV|8|22|Господь имел меня началом пути Своего, прежде созданий Своих, искони;
PROV|8|23|от века я помазана, от начала, прежде бытия земли.
PROV|8|24|Я родилась, когда еще не существовали бездны, когда еще не было источников, обильных водою.
PROV|8|25|Я родилась прежде, нежели водружены были горы, прежде холмов,
PROV|8|26|когда еще Он не сотворил ни земли, ни полей, ни начальных пылинок вселенной.
PROV|8|27|Когда Он уготовлял небеса, [я была] там. Когда Он проводил круговую черту по лицу бездны,
PROV|8|28|когда утверждал вверху облака, когда укреплял источники бездны,
PROV|8|29|когда давал морю устав, чтобы воды не переступали пределов его, когда полагал основания земли:
PROV|8|30|тогда я была при Нем художницею, и была радостью всякий день, веселясь пред лицем Его во все время,
PROV|8|31|веселясь на земном кругу Его, и радость моя [была] с сынами человеческими.
PROV|8|32|Итак, дети, послушайте меня; и блаженны те, которые хранят пути мои!
PROV|8|33|Послушайте наставления и будьте мудры, и не отступайте [от] [него].
PROV|8|34|Блажен человек, который слушает меня, бодрствуя каждый день у ворот моих и стоя на страже у дверей моих!
PROV|8|35|потому что, кто нашел меня, тот нашел жизнь, и получит благодать от Господа;
PROV|8|36|а согрешающий против меня наносит вред душе своей: все ненавидящие меня любят смерть".
PROV|9|1|Премудрость построила себе дом, вытесала семь столбов его,
PROV|9|2|заколола жертву, растворила вино свое и приготовила у себя трапезу;
PROV|9|3|послала слуг своих провозгласить с возвышенностей городских:
PROV|9|4|"кто неразумен, обратись сюда!" И скудоумному она сказала:
PROV|9|5|"идите, ешьте хлеб мой и пейте вино, мною растворенное;
PROV|9|6|оставьте неразумие, и живите, и ходите путем разума".
PROV|9|7|Поучающий кощунника наживет себе бесславие, и обличающий нечестивого – пятно себе.
PROV|9|8|Не обличай кощунника, чтобы он не возненавидел тебя; обличай мудрого, и он возлюбит тебя;
PROV|9|9|дай [наставление] мудрому, и он будет еще мудрее; научи правдивого, и он приумножит знание.
PROV|9|10|Начало мудрости – страх Господень, и познание Святаго – разум;
PROV|9|11|потому что чрез меня умножатся дни твои, и прибавится тебе лет жизни.
PROV|9|12|если ты мудр, то мудр для себя; и если буен, то один потерпишь.
PROV|9|13|Женщина безрассудная, шумливая, глупая и ничего не знающая
PROV|9|14|садится у дверей дома своего на стуле, на возвышенных местах города,
PROV|9|15|чтобы звать проходящих дорогою, идущих прямо своими путями:
PROV|9|16|"кто глуп, обратись сюда!" и скудоумному сказала она:
PROV|9|17|"воды краденые сладки, и утаенный хлеб приятен".
PROV|9|18|И он не знает, что мертвецы там, и что в глубине преисподней зазванные ею.
PROV|10|1|Притчи Соломона. Сын мудрый радует отца, а сын глупый – огорчение для его матери.
PROV|10|2|Не доставляют пользы сокровища неправедные, правда же избавляет от смерти.
PROV|10|3|Не допустит Господь терпеть голод душе праведного, стяжание же нечестивых исторгнет.
PROV|10|4|Ленивая рука делает бедным, а рука прилежных обогащает.
PROV|10|5|Собирающий во время лета – сын разумный, спящий же во время жатвы – сын беспутный.
PROV|10|6|Благословения – на голове праведника, уста же беззаконных заградит насилие.
PROV|10|7|Память праведника пребудет благословенна, а имя нечестивых омерзеет.
PROV|10|8|Мудрый сердцем принимает заповеди, а глупый устами преткнется.
PROV|10|9|Кто ходит в непорочности, тот ходит безопасно; а кто превращает пути свои, тот будет наказан.
PROV|10|10|Кто мигает глазами, тот причиняет досаду, а глупый устами преткнется.
PROV|10|11|Уста праведника – источник жизни, уста же беззаконных заградит насилие.
PROV|10|12|Ненависть возбуждает раздоры, но любовь покрывает все грехи.
PROV|10|13|В устах разумного находится мудрость, но на теле глупого – розга.
PROV|10|14|Мудрые сберегают знание, но уста глупого – близкая погибель.
PROV|10|15|Имущество богатого – крепкий город его, беда для бедных – скудость их.
PROV|10|16|Труды праведного – к жизни, успех нечестивого – ко греху.
PROV|10|17|Кто хранит наставление, тот на пути к жизни; а отвергающий обличение – блуждает.
PROV|10|18|Кто скрывает ненависть, у того уста лживые; и кто разглашает клевету, тот глуп.
PROV|10|19|При многословии не миновать греха, а сдерживающий уста свои – разумен.
PROV|10|20|Отборное серебро – язык праведного, сердце же нечестивых – ничтожество.
PROV|10|21|Уста праведного пасут многих, а глупые умирают от недостатка разума.
PROV|10|22|Благословение Господне – оно обогащает и печали с собою не приносит.
PROV|10|23|Для глупого преступное деяние как бы забава, а человеку разумному свойственна мудрость.
PROV|10|24|Чего страшится нечестивый, то и постигнет его, а желание праведников исполнится.
PROV|10|25|Как проносится вихрь, [так] нет более нечестивого; а праведник – на вечном основании.
PROV|10|26|Что уксус для зубов и дым для глаз, то ленивый для посылающих его.
PROV|10|27|Страх Господень прибавляет дней, лета же нечестивых сократятся.
PROV|10|28|Ожидание праведников – радость, а надежда нечестивых погибнет.
PROV|10|29|Путь Господень – твердыня для непорочного и страх для делающих беззаконие.
PROV|10|30|Праведник во веки не поколеблется, нечестивые же не поживут на земле.
PROV|10|31|Уста праведника источают мудрость, а язык зловредный отсечется.
PROV|10|32|Уста праведного знают благоприятное, а уста нечестивых – развращенное.
PROV|11|1|Неверные весы – мерзость пред Господом, но правильный вес угоден Ему.
PROV|11|2|Придет гордость, придет и посрамление; но со смиренными – мудрость.
PROV|11|3|Непорочность прямодушных будет руководить их, а лукавство коварных погубит их.
PROV|11|4|Не поможет богатство в день гнева, правда же спасет от смерти.
PROV|11|5|Правда непорочного уравнивает путь его, а нечестивый падет от нечестия своего.
PROV|11|6|Правда прямодушных спасет их, а беззаконники будут уловлены беззаконием своим.
PROV|11|7|Со смертью человека нечестивого исчезает надежда, и ожидание беззаконных погибает.
PROV|11|8|Праведник спасается от беды, а вместо него попадает [в нее] нечестивый.
PROV|11|9|Устами лицемер губит ближнего своего, но праведники прозорливостью спасаются.
PROV|11|10|При благоденствии праведников веселится город, и при погибели нечестивых [бывает] торжество.
PROV|11|11|Благословением праведных возвышается город, а устами нечестивых разрушается.
PROV|11|12|Скудоумный высказывает презрение к ближнему своему; но разумный человек молчит.
PROV|11|13|Кто ходит переносчиком, тот открывает тайну; но верный человек таит дело.
PROV|11|14|При недостатке попечения падает народ, а при многих советниках благоденствует.
PROV|11|15|Зло причиняет себе, кто ручается за постороннего; а кто ненавидит ручательство, тот безопасен.
PROV|11|16|Благонравная жена приобретает славу, а трудолюбивые приобретают богатство.
PROV|11|17|Человек милосердый благотворит душе своей, а жестокосердый разрушает плоть свою.
PROV|11|18|Нечестивый делает дело ненадежное, а сеющему правду – награда верная.
PROV|11|19|Праведность [ведет] к жизни, а стремящийся к злу [стремится] к смерти своей.
PROV|11|20|Мерзость пред Господом – коварные сердцем; но благоугодны Ему непорочные в пути.
PROV|11|21|Можно поручиться, что порочный не останется ненаказанным; семя же праведных спасется.
PROV|11|22|Что золотое кольцо в носу у свиньи, то женщина красивая и – безрассудная.
PROV|11|23|Желание праведных [есть] одно добро, ожидание нечестивых – гнев.
PROV|11|24|Иной сыплет щедро, и [ему] еще прибавляется; а другой сверх меры бережлив, и однако же беднеет.
PROV|11|25|Благотворительная душа будет насыщена, и кто напояет [других], тот и сам напоен будет.
PROV|11|26|Кто удерживает у себя хлеб, того клянет народ; а на голове продающего – благословение.
PROV|11|27|Кто стремится к добру, тот ищет благоволения; а кто ищет зла, к тому оно и приходит.
PROV|11|28|Надеющийся на богатство свое упадет; а праведники, как лист, будут зеленеть.
PROV|11|29|Расстроивающий дом свой получит в удел ветер, и глупый будет рабом мудрого сердцем.
PROV|11|30|Плод праведника – древо жизни, и мудрый привлекает души.
PROV|11|31|Так праведнику воздается на земле, тем паче нечестивому и грешнику.
PROV|12|1|Кто любит наставление, тот любит знание; а кто ненавидит обличение, тот невежда.
PROV|12|2|Добрый приобретает благоволение от Господа; а человека коварного Он осудит.
PROV|12|3|Не утвердит себя человек беззаконием; корень же праведников неподвижен.
PROV|12|4|Добродетельная жена – венец для мужа своего; а позорная – как гниль в костях его.
PROV|12|5|Промышления праведных – правда, а замыслы нечестивых – коварство.
PROV|12|6|Речи нечестивых – засада для пролития крови, уста же праведных спасают их.
PROV|12|7|Коснись нечестивых несчастие – и нет их, а дом праведных стоит.
PROV|12|8|Хвалят человека по мере разума его, а развращенный сердцем будет в презрении.
PROV|12|9|Лучше простой, но работающий на себя, нежели выдающий себя за знатного, но нуждающийся в хлебе.
PROV|12|10|Праведный печется и о жизни скота своего, сердце же нечестивых жестоко.
PROV|12|11|Кто возделывает землю свою, тот будет насыщаться хлебом; а кто идет по следам празднолюбцев, тот скудоумен.
PROV|12|12|Нечестивый желает уловить в сеть зла; но корень праведных тверд.
PROV|12|13|Нечестивый уловляется грехами уст своих; но праведник выйдет из беды.
PROV|12|14|От плода уст [своих] человек насыщается добром, и воздаяние человеку – по делам рук его.
PROV|12|15|Путь глупого прямой в его глазах; но кто слушает совета, тот мудр.
PROV|12|16|У глупого тотчас же выкажется гнев его, а благоразумный скрывает оскорбление.
PROV|12|17|Кто говорит то, что знает, тот говорит правду; а у свидетеля ложного – обман.
PROV|12|18|Иной пустослов уязвляет как мечом, а язык мудрых – врачует.
PROV|12|19|Уста правдивые вечно пребывают, а лживый язык – только на мгновение.
PROV|12|20|Коварство – в сердце злоумышленников, радость – у миротворцев.
PROV|12|21|Не приключится праведнику никакого зла, нечестивые же будут преисполнены зол.
PROV|12|22|Мерзость пред Господом – уста лживые, а говорящие истину благоугодны Ему.
PROV|12|23|Человек рассудительный скрывает знание, а сердце глупых высказывает глупость.
PROV|12|24|Рука прилежных будет господствовать, а ленивая будет под данью.
PROV|12|25|Тоска на сердце человека подавляет его, а доброе слово развеселяет его.
PROV|12|26|Праведник указывает ближнему своему путь, а путь нечестивых вводит их в заблуждение.
PROV|12|27|Ленивый не жарит своей дичи; а имущество человека прилежного многоценно.
PROV|12|28|На пути правды – жизнь, и на стезе ее нет смерти.
PROV|13|1|Мудрый сын [слушает] наставление отца, а буйный не слушает обличения.
PROV|13|2|От плода уст [своих] человек вкусит добро, душа же законопреступников – зло.
PROV|13|3|Кто хранит уста свои, тот бережет душу свою; а кто широко раскрывает свой рот, тому беда.
PROV|13|4|Душа ленивого желает, но тщетно; а душа прилежных насытится.
PROV|13|5|Праведник ненавидит ложное слово, а нечестивый срамит и бесчестит [себя].
PROV|13|6|Правда хранит непорочного в пути, а нечестие губит грешника.
PROV|13|7|Иной выдает себя за богатого, а у него ничего нет; другой выдает себя за бедного, а у него богатства много.
PROV|13|8|Богатством своим человек выкупает жизнь [свою], а бедный и угрозы не слышит.
PROV|13|9|Свет праведных весело горит, светильник же нечестивых угасает.
PROV|13|10|От высокомерия происходит раздор, а у советующихся – мудрость.
PROV|13|11|Богатство от суетности истощается, а собирающий трудами умножает его.
PROV|13|12|Надежда, долго не сбывающаяся, томит сердце, а исполнившееся желание – [как] древо жизни.
PROV|13|13|Кто пренебрегает словом, тот причиняет вред себе; а кто боится заповеди, тому воздается.
PROV|13|14|[У сына лукавого ничего нет доброго, а у разумного раба дела благоуспешны, и путь его прямой.]
PROV|13|15|Учение мудрого – источник жизни, удаляющий от сетей смерти.
PROV|13|16|Добрый разум доставляет приятность, путь же беззаконных жесток.
PROV|13|17|Всякий благоразумный действует с знанием, а глупый выставляет напоказ глупость.
PROV|13|18|Худой посол попадает в беду, а верный посланник – спасение.
PROV|13|19|Нищета и посрамление отвергающему учение; а кто соблюдает наставление, будет в чести.
PROV|13|20|Желание исполнившееся – приятно для души; но несносно для глупых уклоняться от зла.
PROV|13|21|Общающийся с мудрыми будет мудр, а кто дружит с глупыми, развратится.
PROV|13|22|Грешников преследует зло, а праведникам воздается добром.
PROV|13|23|Добрый оставляет наследство [и] внукам, а богатство грешника сберегается для праведного.
PROV|13|24|Много хлеба [бывает] и на ниве бедных; но некоторые гибнут от беспорядка.
PROV|13|25|Кто жалеет розги своей, тот ненавидит сына; а кто любит, тот с детства наказывает его.
PROV|13|26|Праведник ест до сытости, а чрево беззаконных терпит лишение.
PROV|14|1|Мудрая жена устроит дом свой, а глупая разрушит его своими руками.
PROV|14|2|Идущий прямым путем боится Господа; но чьи пути кривы, тот небрежет о Нем.
PROV|14|3|В устах глупого – бич гордости; уста же мудрых охраняют их.
PROV|14|4|Где нет волов, [там] ясли пусты; а много прибыли от силы волов.
PROV|14|5|Верный свидетель не лжет, а свидетель ложный наговорит много лжи.
PROV|14|6|Распутный ищет мудрости, и не находит; а для разумного знание легко.
PROV|14|7|Отойди от человека глупого, у которого ты не замечаешь разумных уст.
PROV|14|8|Мудрость разумного – знание пути своего, глупость же безрассудных – заблуждение.
PROV|14|9|Глупые смеются над грехом, а посреди праведных – благоволение.
PROV|14|10|Сердце знает горе души своей, и в радость его не вмешается чужой.
PROV|14|11|Дом беззаконных разорится, а жилище праведных процветет.
PROV|14|12|Есть пути, которые кажутся человеку прямыми; но конец их – путь к смерти.
PROV|14|13|И при смехе [иногда] болит сердце, и концом радости бывает печаль.
PROV|14|14|Человек с развращенным сердцем насытится от путей своих, и добрый – от своих.
PROV|14|15|Глупый верит всякому слову, благоразумный же внимателен к путям своим.
PROV|14|16|Мудрый боится и удаляется от зла, а глупый раздражителен и самонадеян.
PROV|14|17|Вспыльчивый может сделать глупость; но человек, умышленно делающий зло, ненавистен.
PROV|14|18|Невежды получают в удел себе глупость, а благоразумные увенчаются знанием.
PROV|14|19|Преклонятся злые пред добрыми и нечестивые – у ворот праведника.
PROV|14|20|Бедный ненавидим бывает даже близким своим, а у богатого много друзей.
PROV|14|21|Кто презирает ближнего своего, тот грешит; а кто милосерд к бедным, тот блажен.
PROV|14|22|Не заблуждаются ли умышляющие зло? но милость и верность у благомыслящих.
PROV|14|23|От всякого труда есть прибыль, а от пустословия только ущерб.
PROV|14|24|Венец мудрых – богатство их, а глупость невежд глупость [и] [есть].
PROV|14|25|Верный свидетель спасает души, а лживый наговорит много лжи.
PROV|14|26|В страхе пред Господом – надежда твердая, и сынам Своим Он прибежище.
PROV|14|27|Страх Господень – источник жизни, удаляющий от сетей смерти.
PROV|14|28|Во множестве народа – величие царя, а при малолюдстве народа беда государю.
PROV|14|29|У терпеливого человека много разума, а раздражительный выказывает глупость.
PROV|14|30|Кроткое сердце – жизнь для тела, а зависть – гниль для костей.
PROV|14|31|Кто теснит бедного, тот хулит Творца его; чтущий же Его благотворит нуждающемуся.
PROV|14|32|За зло свое нечестивый будет отвергнут, а праведный и при смерти своей имеет надежду.
PROV|14|33|Мудрость почиет в сердце разумного, и среди глупых дает знать о себе.
PROV|14|34|Праведность возвышает народ, а беззаконие – бесчестие народов.
PROV|14|35|Благоволение царя – к рабу разумному, а гнев его – против того, кто позорит его.
PROV|15|1|Кроткий ответ отвращает гнев, а оскорбительное слово возбуждает ярость.
PROV|15|2|Язык мудрых сообщает добрые знания, а уста глупых изрыгают глупость.
PROV|15|3|На всяком месте очи Господни: они видят злых и добрых.
PROV|15|4|Кроткий язык – древо жизни, но необузданный – сокрушение духа.
PROV|15|5|Глупый пренебрегает наставлением отца своего; а кто внимает обличениям, тот благоразумен.
PROV|15|6|В доме праведника – обилие сокровищ, а в прибытке нечестивого – расстройство.
PROV|15|7|Уста мудрых распространяют знание, а сердце глупых не так.
PROV|15|8|Жертва нечестивых – мерзость пред Господом, а молитва праведных благоугодна Ему.
PROV|15|9|Мерзость пред Господом – путь нечестивого, а идущего путем правды Он любит.
PROV|15|10|Злое наказание – уклоняющемуся от пути, и ненавидящий обличение погибнет.
PROV|15|11|Преисподняя и Аваддон [открыты] пред Господом, тем более сердца сынов человеческих.
PROV|15|12|Не любит распутный обличающих его, и к мудрым не пойдет.
PROV|15|13|Веселое сердце делает лице веселым, а при сердечной скорби дух унывает.
PROV|15|14|Сердце разумного ищет знания, уста же глупых питаются глупостью.
PROV|15|15|Все дни несчастного печальны; а у кого сердце весело, у того всегда пир.
PROV|15|16|Лучше немногое при страхе Господнем, нежели большое сокровище, и при нем тревога.
PROV|15|17|Лучше блюдо зелени, и при нем любовь, нежели откормленный бык, и при нем ненависть.
PROV|15|18|Вспыльчивый человек возбуждает раздор, а терпеливый утишает распрю.
PROV|15|19|Путь ленивого – как терновый плетень, а путь праведных – гладкий.
PROV|15|20|Мудрый сын радует отца, а глупый человек пренебрегает мать свою.
PROV|15|21|Глупость – радость для малоумного, а человек разумный идет прямою дорогою.
PROV|15|22|Без совета предприятия расстроятся, а при множестве советников они состоятся.
PROV|15|23|Радость человеку в ответе уст его, и как хорошо слово вовремя!
PROV|15|24|Путь жизни мудрого вверх, чтобы уклониться от преисподней внизу.
PROV|15|25|Дом надменных разорит Господь, а межу вдовы укрепит.
PROV|15|26|Мерзость пред Господом – помышления злых, слова же непорочных угодны Ему.
PROV|15|27|Корыстолюбивый расстроит дом свой, а ненавидящий подарки будет жить.
PROV|15|28|Сердце праведного обдумывает ответ, а уста нечестивых изрыгают зло.
PROV|15|29|Далек Господь от нечестивых, а молитву праведников слышит.
PROV|15|30|Светлый взгляд радует сердце, добрая весть утучняет кости.
PROV|15|31|Ухо, внимательное к учению жизни, пребывает между мудрыми.
PROV|15|32|Отвергающий наставление нерадеет о своей душе; а кто внимает обличению, тот приобретает разум.
PROV|15|33|Страх Господень научает мудрости, и славе предшествует смирение.
PROV|16|1|Человеку [принадлежат] предположения сердца, но от Господа ответ языка.
PROV|16|2|Все пути человека чисты в его глазах, но Господь взвешивает души.
PROV|16|3|Предай Господу дела твои, и предприятия твои совершатся.
PROV|16|4|Все сделал Господь ради Себя; и даже нечестивого [блюдет] на день бедствия.
PROV|16|5|Мерзость пред Господом всякий надменный сердцем; можно поручиться, что он не останется ненаказанным.
PROV|16|6|Милосердием и правдою очищается грех, и страх Господень отводит от зла.
PROV|16|7|Когда Господу угодны пути человека, Он и врагов его примиряет с ним.
PROV|16|8|Лучше немногое с правдою, нежели множество прибытков с неправдою.
PROV|16|9|Сердце человека обдумывает свой путь, но Господь управляет шествием его.
PROV|16|10|В устах царя – слово вдохновенное; уста его не должны погрешать на суде.
PROV|16|11|Верные весы и весовые чаши – от Господа; от Него же все гири в суме.
PROV|16|12|Мерзость для царей – дело беззаконное, потому что правдою утверждается престол.
PROV|16|13|Приятны царю уста правдивые, и говорящего истину он любит.
PROV|16|14|Царский гнев – вестник смерти; но мудрый человек умилостивит его.
PROV|16|15|В светлом взоре царя – жизнь, и благоволение его – как облако с поздним дождем.
PROV|16|16|Приобретение мудрости гораздо лучше золота, и приобретение разума предпочтительнее отборного серебра.
PROV|16|17|Путь праведных – уклонение от зла: тот бережет душу свою, кто хранит путь свой.
PROV|16|18|Погибели предшествует гордость, и падению – надменность.
PROV|16|19|Лучше смиряться духом с кроткими, нежели разделять добычу с гордыми.
PROV|16|20|Кто ведет дело разумно, тот найдет благо, и кто надеется на Господа, тот блажен.
PROV|16|21|Мудрый сердцем прозовется благоразумным, и сладкая речь прибавит к учению.
PROV|16|22|Разум для имеющих его – источник жизни, а ученость глупых – глупость.
PROV|16|23|Сердце мудрого делает язык его мудрым и умножает знание в устах его.
PROV|16|24|Приятная речь – сотовый мед, сладка для души и целебна для костей.
PROV|16|25|Есть пути, которые кажутся человеку прямыми, но конец их путь к смерти.
PROV|16|26|Трудящийся трудится для себя, потому что понуждает его [к] [тому] рот его.
PROV|16|27|Человек лукавый замышляет зло, и на устах его как бы огонь палящий.
PROV|16|28|Человек коварный сеет раздор, и наушник разлучает друзей.
PROV|16|29|Человек неблагонамеренный развращает ближнего своего и ведет его на путь недобрый;
PROV|16|30|прищуривает глаза свои, чтобы придумать коварство; закусывая себе губы, совершает злодейство.
PROV|16|31|Венец славы – седина, которая находится на пути правды.
PROV|16|32|Долготерпеливый лучше храброго, и владеющий собою [лучше] завоевателя города.
PROV|16|33|В полу бросается жребий, но все решение его – от Господа.
PROV|17|1|Лучше кусок сухого хлеба, и с ним мир, нежели дом, полный заколотого скота, с раздором.
PROV|17|2|Разумный раб господствует над беспутным сыном и между братьями разделит наследство.
PROV|17|3|Плавильня – для серебра, и горнило – для золота, а сердца испытывает Господь.
PROV|17|4|Злодей внимает устам беззаконным, лжец слушается языка пагубного.
PROV|17|5|Кто ругается над нищим, тот хулит Творца его; кто радуется несчастью, тот не останется ненаказанным.
PROV|17|6|Венец стариков – сыновья сыновей, и слава детей – родители их.
PROV|17|7|Неприлична глупому важная речь, тем паче знатному – уста лживые.
PROV|17|8|Подарок – драгоценный камень в глазах владеющего им: куда ни обратится он, успеет.
PROV|17|9|Прикрывающий проступок ищет любви; а кто снова напоминает о нем, тот удаляет друга.
PROV|17|10|На разумного сильнее действует выговор, нежели на глупого сто ударов.
PROV|17|11|Возмутитель ищет только зла; поэтому жестокий ангел будет послан против него.
PROV|17|12|Лучше встретить человеку медведицу, лишенную детей, нежели глупца с его глупостью.
PROV|17|13|Кто за добро воздает злом, от дома того не отойдет зло.
PROV|17|14|Начало ссоры – как прорыв воды; оставь ссору прежде, нежели разгорелась она.
PROV|17|15|Оправдывающий нечестивого и обвиняющий праведного – оба мерзость пред Господом.
PROV|17|16|К чему сокровище в руках глупца? Для приобретения мудрости [у] [него] нет разума.
PROV|17|17|Друг любит во всякое время и, как брат, явится во время несчастья.
PROV|17|18|Человек малоумный дает руку и ручается за ближнего своего.
PROV|17|19|Кто любит ссоры, любит грех, и кто высоко поднимает ворота свои, тот ищет падения.
PROV|17|20|Коварное сердце не найдет добра, и лукавый язык попадет в беду.
PROV|17|21|Родил кто глупого, – себе на горе, и отец глупого не порадуется.
PROV|17|22|Веселое сердце благотворно, как врачевство, а унылый дух сушит кости.
PROV|17|23|Нечестивый берет подарок из пазухи, чтобы извратить пути правосудия.
PROV|17|24|Мудрость – пред лицем у разумного, а глаза глупца – на конце земли.
PROV|17|25|Глупый сын – досада отцу своему и огорчение для матери своей.
PROV|17|26|Нехорошо и обвинять правого, [и] бить вельмож за правду.
PROV|17|27|Разумный воздержан в словах своих, и благоразумный хладнокровен.
PROV|17|28|И глупец, когда молчит, может показаться мудрым, и затворяющий уста свои – благоразумным.
PROV|18|1|Прихоти ищет своенравный, восстает против всего умного.
PROV|18|2|Глупый не любит знания, а только бы выказать свой ум.
PROV|18|3|С приходом нечестивого приходит и презрение, а с бесславием – поношение.
PROV|18|4|Слова уст человеческих – глубокие воды; источник мудрости – струящийся поток.
PROV|18|5|Нехорошо быть лицеприятным к нечестивому, чтобы ниспровергнуть праведного на суде.
PROV|18|6|Уста глупого идут в ссору, и слова его вызывают побои.
PROV|18|7|Язык глупого – гибель для него, и уста его – сеть для души его.
PROV|18|8|[Ленивого низлагает страх, а души женоподобные будут голодать.]
PROV|18|9|Слова наушника – как лакомства, и они входят во внутренность чрева.
PROV|18|10|Нерадивый в работе своей – брат расточителю.
PROV|18|11|Имя Господа – крепкая башня: убегает в нее праведник – и безопасен.
PROV|18|12|Имение богатого – крепкий город его, и как высокая ограда в его воображении.
PROV|18|13|Перед падением возносится сердце человека, а смирение предшествует славе.
PROV|18|14|Кто дает ответ не выслушав, тот глуп, и стыд ему.
PROV|18|15|Дух человека переносит его немощи; а пораженный дух – кто может подкрепить его?
PROV|18|16|Сердце разумного приобретает знание, и ухо мудрых ищет знания.
PROV|18|17|Подарок у человека дает ему простор и до вельмож доведет его.
PROV|18|18|Первый в тяжбе своей прав, но приходит соперник его и исследывает его.
PROV|18|19|Жребий прекращает споры и решает между сильными.
PROV|18|20|Озлобившийся брат [неприступнее] крепкого города, и ссоры подобны запорам замка.
PROV|18|21|От плода уст человека наполняется чрево его; произведением уст своих он насыщается.
PROV|18|22|Смерть и жизнь – во власти языка, и любящие его вкусят от плодов его.
PROV|18|23|Кто нашел [добрую] жену, тот нашел благо и получил благодать от Господа.
PROV|18|24|С мольбою говорит нищий, а богатый отвечает грубо.
PROV|18|25|Кто хочет иметь друзей, тот и сам должен быть дружелюбным; и бывает друг, более привязанный, нежели брат.
PROV|19|1|Лучше бедный, ходящий в своей непорочности, нежели [богатый] со лживыми устами, и притом глупый.
PROV|19|2|Нехорошо душе без знания, и торопливый ногами оступится.
PROV|19|3|Глупость человека извращает путь его, а сердце его негодует на Господа.
PROV|19|4|Богатство прибавляет много друзей, а бедный оставляется и другом своим.
PROV|19|5|Лжесвидетель не останется ненаказанным, и кто говорит ложь, не спасется.
PROV|19|6|Многие заискивают у знатных, и всякий – друг человеку, делающему подарки.
PROV|19|7|Бедного ненавидят все братья его, тем паче друзья его удаляются от него: гонится за ними, чтобы поговорить, но и этого нет.
PROV|19|8|Кто приобретает разум, тот любит душу свою; кто наблюдает благоразумие, тот находит благо.
PROV|19|9|Лжесвидетель не останется ненаказанным, и кто говорит ложь, погибнет.
PROV|19|10|Неприлична глупцу пышность, тем паче рабу господство над князьями.
PROV|19|11|Благоразумие делает человека медленным на гнев, и слава для него – быть снисходительным к проступкам.
PROV|19|12|Гнев царя – как рев льва, а благоволение его – как роса на траву.
PROV|19|13|Глупый сын – сокрушение для отца своего, и сварливая жена – сточная труба.
PROV|19|14|Дом и имение – наследство от родителей, а разумная жена – от Господа.
PROV|19|15|Леность погружает в сонливость, и нерадивая душа будет терпеть голод.
PROV|19|16|Хранящий заповедь хранит душу свою, а нерадящий о путях своих погибнет.
PROV|19|17|Благотворящий бедному дает взаймы Господу, и Он воздаст ему за благодеяние его.
PROV|19|18|Наказывай сына своего, доколе есть надежда, и не возмущайся криком его.
PROV|19|19|Гневливый пусть терпит наказание, потому что, если пощадишь [его], придется тебе еще больше наказывать его.
PROV|19|20|Слушайся совета и принимай обличение, чтобы сделаться тебе впоследствии мудрым.
PROV|19|21|Много замыслов в сердце человека, но состоится только определенное Господом.
PROV|19|22|Радость человеку – благотворительность его, и бедный человек лучше, нежели лживый.
PROV|19|23|Страх Господень [ведет] к жизни, и [кто имеет его], всегда будет доволен, и зло не постигнет его.
PROV|19|24|Ленивый опускает руку свою в чашу, и не хочет донести ее до рта своего.
PROV|19|25|Если ты накажешь кощунника, то и простой сделается благоразумным; и [если] обличишь разумного, то он поймет наставление.
PROV|19|26|Разоряющий отца и выгоняющий мать – сын срамной и бесчестный.
PROV|19|27|Перестань, сын мой, слушать внушения об уклонении от изречений разума.
PROV|19|28|Лукавый свидетель издевается над судом, и уста беззаконных глотают неправду.
PROV|19|29|Готовы для кощунствующих суды, и побои – на тело глупых.
PROV|20|1|Вино – глумливо, сикера – буйна; и всякий, увлекающийся ими, неразумен.
PROV|20|2|Гроза царя – как бы рев льва: кто раздражает его, тот грешит против самого себя.
PROV|20|3|Честь для человека – отстать от ссоры; а всякий глупец задорен.
PROV|20|4|Ленивец зимою не пашет: поищет летом – и нет ничего.
PROV|20|5|Помыслы в сердце человека – глубокие воды, но человек разумный вычерпывает их.
PROV|20|6|Многие хвалят человека за милосердие, но правдивого человека кто находит?
PROV|20|7|Праведник ходит в своей непорочности: блаженны дети его после него!
PROV|20|8|Царь, сидящий на престоле суда, разгоняет очами своими все злое.
PROV|20|9|Кто может сказать: "я очистил мое сердце, я чист от греха моего?"
PROV|20|10|Неодинаковые весы, неодинаковая мера, то и другое – мерзость пред Господом.
PROV|20|11|Можно узнать даже отрока по занятиям его, чисто ли и правильно ли будет поведение его.
PROV|20|12|Ухо слышащее и глаз видящий – и то и другое создал Господь.
PROV|20|13|Не люби спать, чтобы тебе не обеднеть; держи открытыми глаза твои, и будешь досыта есть хлеб.
PROV|20|14|"Дурно, дурно", говорит покупатель, а когда отойдет, хвалится.
PROV|20|15|Есть золото и много жемчуга, но драгоценная утварь – уста разумные.
PROV|20|16|Возьми платье его, так как он поручился за чужого; и за стороннего возьми от него залог.
PROV|20|17|Сладок для человека хлеб, [приобретенный] неправдою; но после рот его наполнится дресвою.
PROV|20|18|Предприятия получают твердость чрез совещание, и по совещании веди войну.
PROV|20|19|Кто ходит переносчиком, тот открывает тайну; и кто широко раскрывает рот, с тем не сообщайся.
PROV|20|20|Кто злословит отца своего и свою мать, того светильник погаснет среди глубокой тьмы.
PROV|20|21|Наследство, поспешно захваченное вначале, не благословится впоследствии.
PROV|20|22|Не говори: "я отплачу за зло"; предоставь Господу, и Он сохранит тебя.
PROV|20|23|Мерзость пред Господом – неодинаковые гири, и неверные весы – не добро.
PROV|20|24|От Господа направляются шаги человека; человеку же как узнать путь свой?
PROV|20|25|Сеть для человека – поспешно давать обет, и после обета обдумывать.
PROV|20|26|Мудрый царь вывеет нечестивых и обратит на них колесо.
PROV|20|27|Светильник Господень – дух человека, испытывающий все глубины сердца.
PROV|20|28|Милость и истина охраняют царя, и милостью он поддерживает престол свой.
PROV|20|29|Слава юношей – сила их, а украшение стариков – седина.
PROV|20|30|Раны от побоев – врачевство против зла, и удары, проникающие во внутренности чрева.
PROV|21|1|Сердце царя – в руке Господа, как потоки вод: куда захочет, Он направляет его.
PROV|21|2|Всякий путь человека прям в глазах его; но Господь взвешивает сердца.
PROV|21|3|Соблюдение правды и правосудия более угодно Господу, нежели жертва.
PROV|21|4|Гордость очей и надменность сердца, отличающие нечестивых, – грех.
PROV|21|5|Помышления прилежного стремятся к изобилию, а всякий торопливый терпит лишение.
PROV|21|6|Приобретение сокровища лживым языком – мимолетное дуновение ищущих смерти.
PROV|21|7|Насилие нечестивых обрушится на них, потому что они отреклись соблюдать правду.
PROV|21|8|Превратен путь человека развращенного; а кто чист, того действие прямо.
PROV|21|9|Лучше жить в углу на кровле, нежели со сварливою женою в пространном доме.
PROV|21|10|Душа нечестивого желает зла: не найдет милости в глазах его и друг его.
PROV|21|11|Когда наказывается кощунник, простой делается мудрым; и когда вразумляется мудрый, то он приобретает знание.
PROV|21|12|Праведник наблюдает за домом нечестивого: как повергаются нечестивые в несчастие.
PROV|21|13|Кто затыкает ухо свое от вопля бедного, тот и сам будет вопить, – и не будет услышан.
PROV|21|14|Подарок тайный тушит гнев, и дар в пазуху – сильную ярость.
PROV|21|15|Соблюдение правосудия – радость для праведника и страх для делающих зло.
PROV|21|16|Человек, сбившийся с пути разума, водворится в собрании мертвецов.
PROV|21|17|Кто любит веселье, обеднеет; а кто любит вино и тук, не разбогатеет.
PROV|21|18|Выкупом будет за праведного нечестивый и за прямодушного – лукавый.
PROV|21|19|Лучше жить в земле пустынной, нежели с женою сварливою и сердитою.
PROV|21|20|Вожделенное сокровище и тук – в доме мудрого; а глупый человек расточает их.
PROV|21|21|Соблюдающий правду и милость найдет жизнь, правду и славу.
PROV|21|22|Мудрый входит в город сильных и ниспровергает крепость, на которую они надеялись.
PROV|21|23|Кто хранит уста свои и язык свой, тот хранит от бед душу свою.
PROV|21|24|Надменный злодей – кощунник имя ему – действует в пылу гордости.
PROV|21|25|Алчба ленивца убьет его, потому что руки его отказываются работать;
PROV|21|26|всякий день он сильно алчет, а праведник дает и не жалеет.
PROV|21|27|Жертва нечестивых – мерзость, особенно когда с лукавством приносят ее.
PROV|21|28|Лжесвидетель погибнет; а человек, который говорит, что знает, будет говорить всегда.
PROV|21|29|Человек нечестивый дерзок лицом своим, а праведный держит прямо путь свой.
PROV|21|30|Нет мудрости, и нет разума, и нет совета вопреки Господу.
PROV|21|31|Коня приготовляют на день битвы, но победа – от Господа.
PROV|22|1|Доброе имя лучше большого богатства, и добрая слава лучше серебра и золота.
PROV|22|2|Богатый и бедный встречаются друг с другом: того и другого создал Господь.
PROV|22|3|Благоразумный видит беду, и укрывается; а неопытные идут вперед, и наказываются.
PROV|22|4|За смирением следует страх Господень, богатство и слава и жизнь.
PROV|22|5|Терны и сети на пути коварного; кто бережет душу свою, удались от них.
PROV|22|6|Наставь юношу при начале пути его: он не уклонится от него, когда и состарится.
PROV|22|7|Богатый господствует над бедным, и должник [делается] рабом заимодавца.
PROV|22|8|Сеющий неправду пожнет беду, и трости гнева его не станет.
PROV|22|9|Милосердый будет благословляем, потому что дает бедному от хлеба своего.
PROV|22|10|Прогони кощунника, и удалится раздор, и прекратятся ссора и брань.
PROV|22|11|Кто любит чистоту сердца, у того приятность на устах, тому царь – друг.
PROV|22|12|Очи Господа охраняют знание, а слова законопреступника Он ниспровергает.
PROV|22|13|Ленивец говорит: "лев на улице! посреди площади убьют меня!"
PROV|22|14|Глубокая пропасть – уста блудниц: на кого прогневается Господь, тот упадет туда.
PROV|22|15|Глупость привязалась к сердцу юноши, но исправительная розга удалит ее от него.
PROV|22|16|Кто обижает бедного, чтобы умножить свое богатство, и кто дает богатому, тот обеднеет.
PROV|22|17|Приклони ухо твое, и слушай слова мудрых, и сердце твое обрати к моему знанию;
PROV|22|18|потому что утешительно будет, если ты будешь хранить их в сердце твоем, и они будут также в устах твоих.
PROV|22|19|Чтобы упование твое было на Господа, я учу тебя и сегодня, и ты [помни].
PROV|22|20|Не писал ли я тебе трижды в советах и наставлении,
PROV|22|21|чтобы научить тебя точным словам истины, дабы ты мог передавать слова истины посылающим тебя?
PROV|22|22|Не будь грабителем бедного, потому что он беден, и не притесняй несчастного у ворот,
PROV|22|23|потому что Господь вступится в дело их и исхитит душу у грабителей их.
PROV|22|24|Не дружись с гневливым и не сообщайся с человеком вспыльчивым,
PROV|22|25|чтобы не научиться путям его и не навлечь петли на душу твою.
PROV|22|26|Не будь из тех, которые дают руки и поручаются за долги:
PROV|22|27|если тебе нечем заплатить, то для чего доводить себя, чтобы взяли постель твою из–под тебя?
PROV|22|28|Не передвигай межи давней, которую провели отцы твои.
PROV|22|29|Видел ли ты человека проворного в своем деле? Он будет стоять перед царями, он не будет стоять перед простыми.
PROV|23|1|Когда сядешь вкушать пищу с властелином, то тщательно наблюдай, что перед тобою,
PROV|23|2|и поставь преграду в гортани твоей, если ты алчен.
PROV|23|3|Не прельщайся лакомыми яствами его; это – обманчивая пища.
PROV|23|4|Не заботься о том, чтобы нажить богатство; оставь такие мысли твои.
PROV|23|5|Устремишь глаза твои на него, и – его уже нет; потому что оно сделает себе крылья и, как орел, улетит к небу.
PROV|23|6|Не вкушай пищи у человека завистливого и не прельщайся лакомыми яствами его;
PROV|23|7|потому что, каковы мысли в душе его, таков и он; "ешь и пей", говорит он тебе, а сердце его не с тобою.
PROV|23|8|Кусок, который ты съел, изблюешь, и добрые слова твои ты потратишь напрасно.
PROV|23|9|В уши глупого не говори, потому что он презрит разумные слова твои.
PROV|23|10|Не передвигай межи давней и на поля сирот не заходи,
PROV|23|11|потому что Защитник их силен; Он вступится в дело их с тобою.
PROV|23|12|Приложи сердце твое к учению и уши твои – к умным словам.
PROV|23|13|Не оставляй юноши без наказания: если накажешь его розгою, он не умрет;
PROV|23|14|ты накажешь его розгою и спасешь душу его от преисподней.
PROV|23|15|Сын мой! если сердце твое будет мудро, то порадуется и мое сердце;
PROV|23|16|и внутренности мои будут радоваться, когда уста твои будут говорить правое.
PROV|23|17|Да не завидует сердце твое грешникам, но да пребудет оно во все дни в страхе Господнем;
PROV|23|18|потому что есть будущность, и надежда твоя не потеряна.
PROV|23|19|Слушай, сын мой, и будь мудр, и направляй сердце твое на прямой путь.
PROV|23|20|Не будь между упивающимися вином, между пресыщающимися мясом:
PROV|23|21|потому что пьяница и пресыщающийся обеднеют, и сонливость оденет в рубище.
PROV|23|22|Слушайся отца твоего: он родил тебя; и не пренебрегай матери твоей, когда она и состарится.
PROV|23|23|Купи истину и не продавай мудрости и учения и разума.
PROV|23|24|Торжествует отец праведника, и родивший мудрого радуется о нем.
PROV|23|25|Да веселится отец твой и да торжествует мать твоя, родившая тебя.
PROV|23|26|Сын мой! отдай сердце твое мне, и глаза твои да наблюдают пути мои,
PROV|23|27|потому что блудница – глубокая пропасть, и чужая жена – тесный колодезь;
PROV|23|28|она, как разбойник, сидит в засаде и умножает между людьми законопреступников.
PROV|23|29|У кого вой? у кого стон? у кого ссоры? у кого горе? у кого раны без причины? у кого багровые глаза?
PROV|23|30|У тех, которые долго сидят за вином, которые приходят отыскивать [вина] приправленного.
PROV|23|31|Не смотри на вино, как оно краснеет, как оно искрится в чаше, как оно ухаживается ровно:
PROV|23|32|впоследствии, как змей, оно укусит, и ужалит, как аспид;
PROV|23|33|глаза твои будут смотреть на чужих жен, и сердце твое заговорит развратное,
PROV|23|34|и ты будешь, как спящий среди моря и как спящий на верху мачты.
PROV|23|35|[И скажешь]: "били меня, мне не было больно; толкали меня, я не чувствовал. Когда проснусь, опять буду искать того же".
PROV|24|1|Не ревнуй злым людям и не желай быть с ними,
PROV|24|2|потому что о насилии помышляет сердце их, и о злом говорят уста их.
PROV|24|3|Мудростью устрояется дом и разумом утверждается,
PROV|24|4|и с уменьем внутренности его наполняются всяким драгоценным и прекрасным имуществом.
PROV|24|5|Человек мудрый силен, и человек разумный укрепляет силу свою.
PROV|24|6|Поэтому с обдуманностью веди войну твою, и успех [будет] при множестве совещаний.
PROV|24|7|Для глупого слишком высока мудрость; у ворот не откроет он уст своих.
PROV|24|8|Кто замышляет сделать зло, того называют злоумышленником.
PROV|24|9|Помысл глупости – грех, и кощунник – мерзость для людей.
PROV|24|10|Если ты в день бедствия оказался слабым, то бедна сила твоя.
PROV|24|11|Спасай взятых на смерть, и неужели откажешься от обреченных на убиение?
PROV|24|12|Скажешь ли: "вот, мы не знали этого"? А Испытующий сердца разве не знает? Наблюдающий над душею твоею знает это, и воздаст человеку по делам его.
PROV|24|13|Ешь, сын мой, мед, потому что он приятен, и сот, который сладок для гортани твоей:
PROV|24|14|таково и познание мудрости для души твоей. Если ты нашел [ее], то есть будущность, и надежда твоя не потеряна.
PROV|24|15|Не злоумышляй, нечестивый, против жилища праведника, не опустошай места покоя его,
PROV|24|16|ибо семь раз упадет праведник, и встанет; а нечестивые впадут в погибель.
PROV|24|17|Не радуйся, когда упадет враг твой, и да не веселится сердце твое, когда он споткнется.
PROV|24|18|Иначе, увидит Господь, и неугодно будет это в очах Его, и Он отвратит от него гнев Свой.
PROV|24|19|Не негодуй на злодеев и не завидуй нечестивым,
PROV|24|20|потому что злой не имеет будущности, – светильник нечестивых угаснет.
PROV|24|21|Бойся, сын мой, Господа и царя; с мятежниками не сообщайся,
PROV|24|22|потому что внезапно придет погибель от них, и беду от них обоих кто предузнает?
PROV|24|23|Сказано также мудрыми: иметь лицеприятие на суде – нехорошо.
PROV|24|24|Кто говорит виновному: "ты прав", того будут проклинать народы, того будут ненавидеть племена;
PROV|24|25|а обличающие будут любимы, и на них придет благословение.
PROV|24|26|В уста целует, кто отвечает словами верными.
PROV|24|27|Соверши дела твои вне дома, окончи их на поле твоем, и потом устрояй и дом твой.
PROV|24|28|Не будь лжесвидетелем на ближнего твоего: к чему тебе обманывать устами твоими?
PROV|24|29|Не говори: "как он поступил со мною, так и я поступлю с ним, воздам человеку по делам его".
PROV|24|30|Проходил я мимо поля человека ленивого и мимо виноградника человека скудоумного:
PROV|24|31|и вот, все это заросло терном, поверхность его покрылась крапивою, и каменная ограда его обрушилась.
PROV|24|32|И посмотрел я, и обратил сердце мое, и посмотрел и получил урок:
PROV|24|33|"немного поспишь, немного подремлешь, немного, сложив руки, полежишь, –
PROV|24|34|и придет, [как] прохожий, бедность твоя, и нужда твоя – как человек вооруженный".
PROV|25|1|И это притчи Соломона, которые собрали мужи Езекии, царя Иудейского.
PROV|25|2|Слава Божия – облекать тайною дело, а слава царей – исследывать дело.
PROV|25|3|Как небо в высоте и земля в глубине, так сердце царей – неисследимо.
PROV|25|4|Отдели примесь от серебра, и выйдет у серебряника сосуд:
PROV|25|5|удали неправедного от царя, и престол его утвердится правдою.
PROV|25|6|Не величайся пред лицем царя, и на месте великих не становись;
PROV|25|7|потому что лучше, когда скажут тебе: "пойди сюда повыше", нежели когда понизят тебя пред знатным, которого видели глаза твои.
PROV|25|8|Не вступай поспешно в тяжбу: иначе что будешь делать при окончании, когда соперник твой осрамит тебя?
PROV|25|9|Веди тяжбу с соперником твоим, но тайны другого не открывай,
PROV|25|10|дабы не укорил тебя услышавший это, и тогда бесчестие твое не отойдет от тебя.
PROV|25|11|Золотые яблоки в серебряных прозрачных сосудах – слово, сказанное прилично.
PROV|25|12|Золотая серьга и украшение из чистого золота – мудрый обличитель для внимательного уха.
PROV|25|13|Что прохлада от снега во время жатвы, то верный посол для посылающего его: он доставляет душе господина своего отраду.
PROV|25|14|Что тучи и ветры без дождя, то человек, хвастающий ложными подарками.
PROV|25|15|Кротостью склоняется к милости вельможа, и мягкий язык переламывает кость.
PROV|25|16|Нашел ты мед, – ешь, сколько тебе потребно, чтобы не пресытиться им и не изблевать его.
PROV|25|17|Не учащай входить в дом друга твоего, чтобы он не наскучил тобою и не возненавидел тебя.
PROV|25|18|Что молот и меч и острая стрела, то человек, произносящий ложное свидетельство против ближнего своего.
PROV|25|19|Что сломанный зуб и расслабленная нога, то надежда на ненадежного [человека] в день бедствия.
PROV|25|20|Что снимающий с себя одежду в холодный день, что уксус на рану, то поющий песни печальному сердцу.
PROV|25|21|Если голоден враг твой, накорми его хлебом; и если он жаждет, напой его водою:
PROV|25|22|ибо, [делая сие], ты собираешь горящие угли на голову его, и Господь воздаст тебе.
PROV|25|23|Северный ветер производит дождь, а тайный язык – недовольные лица.
PROV|25|24|Лучше жить в углу на кровле, нежели со сварливою женою в пространном доме.
PROV|25|25|Что холодная вода для истомленной жаждой души, то добрая весть из дальней страны.
PROV|25|26|Что возмущенный источник и поврежденный родник, то праведник, падающий пред нечестивым.
PROV|25|27|Как нехорошо есть много меду, так домогаться славы не есть слава.
PROV|25|28|Что город разрушенный, без стен, то человек, не владеющий духом своим.
PROV|26|1|Как снег летом и дождь во время жатвы, так честь неприлична глупому.
PROV|26|2|Как воробей вспорхнет, как ласточка улетит, так незаслуженное проклятие не сбудется.
PROV|26|3|Бич для коня, узда для осла, а палка для глупых.
PROV|26|4|Не отвечай глупому по глупости его, чтобы и тебе не сделаться подобным ему;
PROV|26|5|но отвечай глупому по глупости его, чтобы он не стал мудрецом в глазах своих.
PROV|26|6|Подрезывает себе ноги, терпит неприятность тот, кто дает словесное поручение глупцу.
PROV|26|7|Неровно поднимаются ноги у хромого, – и притча в устах глупцов.
PROV|26|8|Что влагающий драгоценный камень в пращу, то воздающий глупому честь.
PROV|26|9|Что [колючий] терн в руке пьяного, то притча в устах глупцов.
PROV|26|10|Сильный делает все произвольно: и глупого награждает, и всякого прохожего награждает.
PROV|26|11|Как пес возвращается на блевотину свою, так глупый повторяет глупость свою.
PROV|26|12|Видал ли ты человека, мудрого в глазах его? На глупого больше надежды, нежели на него.
PROV|26|13|Ленивец говорит: "лев на дороге! лев на площадях!"
PROV|26|14|Дверь ворочается на крючьях своих, а ленивец на постели своей.
PROV|26|15|Ленивец опускает руку свою в чашу, и ему тяжело донести ее до рта своего.
PROV|26|16|Ленивец в глазах своих мудрее семерых, отвечающих обдуманно.
PROV|26|17|Хватает пса за уши, кто, проходя мимо, вмешивается в чужую ссору.
PROV|26|18|Как притворяющийся помешанным бросает огонь, стрелы и смерть,
PROV|26|19|так – человек, который коварно вредит другу своему и потом говорит: "я только пошутил".
PROV|26|20|Где нет больше дров, огонь погасает, и где нет наушника, раздор утихает.
PROV|26|21|Уголь – для жара и дрова – для огня, а человек сварливый – для разжжения ссоры.
PROV|26|22|Слова наушника – как лакомства, и они входят во внутренность чрева.
PROV|26|23|Что нечистым серебром обложенный глиняный сосуд, то пламенные уста и сердце злобное.
PROV|26|24|Устами своими притворяется враг, а в сердце своем замышляет коварство.
PROV|26|25|Если он говорит и нежным голосом, не верь ему, потому что семь мерзостей в сердце его.
PROV|26|26|Если ненависть прикрывается наедине, то откроется злоба его в народном собрании.
PROV|26|27|Кто роет яму, тот упадет в нее, и кто покатит вверх камень, к тому он воротится.
PROV|26|28|Лживый язык ненавидит уязвляемых им, и льстивые уста готовят падение.
PROV|27|1|Не хвались завтрашним днем, потому что не знаешь, что родит тот день.
PROV|27|2|Пусть хвалит тебя другой, а не уста твои, – чужой, а не язык твой.
PROV|27|3|Тяжел камень, весок и песок; но гнев глупца тяжелее их обоих.
PROV|27|4|Жесток гнев, неукротима ярость; но кто устоит против ревности?
PROV|27|5|Лучше открытое обличение, нежели скрытая любовь.
PROV|27|6|Искренни укоризны от любящего, и лживы поцелуи ненавидящего.
PROV|27|7|Сытая душа попирает и сот, а голодной душе все горькое сладко.
PROV|27|8|Как птица, покинувшая гнездо свое, так человек, покинувший место свое.
PROV|27|9|Масть и курение радуют сердце; так сладок [всякому] друг сердечным советом своим.
PROV|27|10|Не покидай друга твоего и друга отца твоего, и в дом брата твоего не ходи в день несчастья твоего: лучше сосед вблизи, нежели брат вдали.
PROV|27|11|Будь мудр, сын мой, и радуй сердце мое; и я буду иметь, что отвечать злословящему меня.
PROV|27|12|Благоразумный видит беду и укрывается; а неопытные идут вперед [и] наказываются.
PROV|27|13|Возьми у него платье его, потому что он поручился за чужого, и за стороннего возьми от него залог.
PROV|27|14|Кто громко хвалит друга своего с раннего утра, того сочтут за злословящего.
PROV|27|15|Непрестанная капель в дождливый день и сварливая жена – равны:
PROV|27|16|кто хочет скрыть ее, тот хочет скрыть ветер и масть в правой руке своей, дающую знать о себе.
PROV|27|17|Железо железо острит, и человек изощряет взгляд друга своего.
PROV|27|18|Кто стережет смоковницу, тот будет есть плоды ее; и кто бережет господина своего, тот будет в чести.
PROV|27|19|Как в воде лицо – к лицу, так сердце человека – к человеку.
PROV|27|20|Преисподняя и Аваддон – ненасытимы; так ненасытимы и глаза человеческие.
PROV|27|21|Что плавильня – для серебра, горнило – для золота, то для человека уста, которые хвалят его.
PROV|27|22|Толки глупого в ступе пестом вместе с зерном, не отделится от него глупость его.
PROV|27|23|Хорошо наблюдай за скотом твоим, имей попечение о стадах;
PROV|27|24|потому что богатство не навек, да и власть разве из рода в род?
PROV|27|25|Прозябает трава, и является зелень, и собирают горные травы.
PROV|27|26|Овцы – на одежду тебе, и козлы – на покупку поля.
PROV|27|27|И довольно козьего молока в пищу тебе, в пищу домашним твоим и на продовольствие служанкам твоим.
PROV|28|1|Нечестивый бежит, когда никто не гонится [за ним]; а праведник смел, как лев.
PROV|28|2|Когда страна отступит от закона, тогда много в ней начальников; а при разумном и знающем муже она долговечна.
PROV|28|3|Человек бедный и притесняющий слабых [то же, что] проливной дождь, смывающий хлеб.
PROV|28|4|Отступники от закона хвалят нечестивых, а соблюдающие закон негодуют на них.
PROV|28|5|Злые люди не разумеют справедливости, а ищущие Господа разумеют все.
PROV|28|6|Лучше бедный, ходящий в своей непорочности, нежели тот, кто извращает пути свои, хотя он и богат.
PROV|28|7|Хранящий закон – сын разумный, а знающийся с расточителями срамит отца своего.
PROV|28|8|Умножающий имение свое ростом и лихвою соберет его для благотворителя бедных.
PROV|28|9|Кто отклоняет ухо свое от слушания закона, того и молитва – мерзость.
PROV|28|10|Совращающий праведных на путь зла сам упадет в свою яму, а непорочные наследуют добро.
PROV|28|11|Человек богатый – мудрец в глазах своих, но умный бедняк обличит его.
PROV|28|12|Когда торжествуют праведники, великая слава, но когда возвышаются нечестивые, люди укрываются.
PROV|28|13|Скрывающий свои преступления не будет иметь успеха; а кто сознается и оставляет их, тот будет помилован.
PROV|28|14|Блажен человек, который всегда пребывает в благоговении; а кто ожесточает сердце свое, тот попадет в беду.
PROV|28|15|Как рыкающий лев и голодный медведь, так нечестивый властелин над бедным народом.
PROV|28|16|Неразумный правитель много делает притеснений, а ненавидящий корысть продолжит дни.
PROV|28|17|Человек, виновный в пролитии человеческой крови, будет бегать до могилы, чтобы кто не схватил его.
PROV|28|18|Кто ходит непорочно, то будет невредим; а ходящий кривыми путями упадет на одном из них.
PROV|28|19|Кто возделывает землю свою, тот будет насыщаться хлебом, а кто подражает праздным, тот насытится нищетою.
PROV|28|20|Верный человек богат благословениями, а кто спешит разбогатеть, тот не останется ненаказанным.
PROV|28|21|Быть лицеприятным – нехорошо: такой человек и за кусок хлеба сделает неправду.
PROV|28|22|Спешит к богатству завистливый человек, и не думает, что нищета постигнет его.
PROV|28|23|Обличающий человека найдет после большую приязнь, нежели тот, кто льстит языком.
PROV|28|24|Кто обкрадывает отца своего и мать свою и говорит: "это не грех", тот – сообщник грабителям.
PROV|28|25|Надменный разжигает ссору, а надеющийся на Господа будет благоденствовать.
PROV|28|26|Кто надеется на себя, тот глуп; а кто ходит в мудрости, тот будет цел.
PROV|28|27|Дающий нищему не обеднеет; а кто закрывает глаза свои от него, на том много проклятий.
PROV|28|28|Когда возвышаются нечестивые, люди укрываются, а когда они падают, умножаются праведники.
PROV|29|1|Человек, который, будучи обличаем, ожесточает выю свою, внезапно сокрушится, и не будет [ему] исцеления.
PROV|29|2|Когда умножаются праведники, веселится народ, а когда господствует нечестивый, народ стенает.
PROV|29|3|Человек, любящий мудрость, радует отца своего; а кто знается с блудницами, тот расточает имение.
PROV|29|4|Царь правосудием утверждает землю, а любящий подарки разоряет ее.
PROV|29|5|Человек, льстящий другу своему, расстилает сеть ногам его.
PROV|29|6|В грехе злого человека – сеть [для него], а праведник веселится и радуется.
PROV|29|7|Праведник тщательно вникает в тяжбу бедных, а нечестивый не разбирает дела.
PROV|29|8|Люди развратные возмущают город, а мудрые утишают мятеж.
PROV|29|9|Умный человек, судясь с человеком глупым, сердится ли, смеется ли, – не имеет покоя.
PROV|29|10|Кровожадные люди ненавидят непорочного, а праведные заботятся о его жизни.
PROV|29|11|Глупый весь гнев свой изливает, а мудрый сдерживает его.
PROV|29|12|Если правитель слушает ложные речи, то и все служащие у него нечестивы.
PROV|29|13|Бедный и лихоимец встречаются друг с другом; но свет глазам того и другого дает Господь.
PROV|29|14|Если царь судит бедных по правде, то престол его навсегда утвердится.
PROV|29|15|Розга и обличение дают мудрость; но отрок, оставленный в небрежении, делает стыд своей матери.
PROV|29|16|При умножении нечестивых умножается беззаконие; но праведники увидят падение их.
PROV|29|17|Наказывай сына твоего, и он даст тебе покой, и доставит радость душе твоей.
PROV|29|18|Без откровения свыше народ необуздан, а соблюдающий закон блажен.
PROV|29|19|Словами не научится раб, потому что, хотя он понимает [их], но не слушается.
PROV|29|20|Видал ли ты человека опрометчивого в словах своих? на глупого больше надежды, нежели на него.
PROV|29|21|Если с детства воспитывать раба в неге, то впоследствии он захочет быть сыном.
PROV|29|22|Человек гневливый заводит ссору, и вспыльчивый много грешит.
PROV|29|23|Гордость человека унижает его, а смиренный духом приобретает честь.
PROV|29|24|Кто делится с вором, тот ненавидит душу свою; слышит он проклятие, но не объявляет о том.
PROV|29|25|Боязнь пред людьми ставит сеть; а надеющийся на Господа будет безопасен.
PROV|29|26|Многие ищут [благосклонного] лица правителя, но судьба человека – от Господа.
PROV|29|27|Мерзость для праведников – человек неправедный, и мерзость для нечестивого – идущий прямым путем.
PROV|30|1|Слова Агура, сына Иакеева. Вдохновенные изречения, [которые] сказал этот человек Ифиилу, Ифиилу и Укалу:
PROV|30|2|подлинно, я более невежда, нежели кто–либо из людей, и разума человеческого нет у меня,
PROV|30|3|и не научился я мудрости, и познания святых не имею.
PROV|30|4|Кто восходил на небо и нисходил? кто собрал ветер в пригоршни свои? кто завязал воду в одежду? кто поставил все пределы земли? какое имя ему? и какое имя сыну его? знаешь ли?
PROV|30|5|Всякое слово Бога чисто; Он – щит уповающим на Него.
PROV|30|6|Не прибавляй к словам Его, чтобы Он не обличил тебя, и ты не оказался лжецом.
PROV|30|7|Двух вещей я прошу у Тебя, не откажи мне, прежде нежели я умру:
PROV|30|8|суету и ложь удали от меня, нищеты и богатства не давай мне, питай меня насущным хлебом,
PROV|30|9|дабы, пресытившись, я не отрекся [Тебя] и не сказал: "кто Господь?" и чтобы, обеднев, не стал красть и употреблять имя Бога моего всуе.
PROV|30|10|Не злословь раба пред господином его, чтобы он не проклял тебя, и ты не остался виноватым.
PROV|30|11|Есть род, который проклинает отца своего и не благословляет матери своей.
PROV|30|12|Есть род, который чист в глазах своих, тогда как не омыт от нечистот своих.
PROV|30|13|Есть род – о, как высокомерны глаза его, и как подняты ресницы его!
PROV|30|14|Есть род, у которого зубы – мечи, и челюсти – ножи, чтобы пожирать бедных на земле и нищих между людьми.
PROV|30|15|У ненасытимости две дочери: "давай, давай!" Вот три ненасытимых, и четыре, которые не скажут: "довольно!"
PROV|30|16|Преисподняя и утроба бесплодная, земля, которая не насыщается водою, и огонь, который не говорит: "довольно!"
PROV|30|17|Глаз, насмехающийся над отцом и пренебрегающий покорностью к матери, выклюют вороны дольные, и сожрут птенцы орлиные!
PROV|30|18|Три вещи непостижимы для меня, и четырех я не понимаю:
PROV|30|19|пути орла на небе, пути змея на скале, пути корабля среди моря и пути мужчины к девице.
PROV|30|20|Таков путь и жены прелюбодейной; поела и обтерла рот свой, и говорит: "я ничего худого не сделала".
PROV|30|21|От трех трясется земля, четырех она не может носить:
PROV|30|22|раба, когда он делается царем; глупого, когда он досыта ест хлеб;
PROV|30|23|позорную женщину, когда она выходит замуж, и служанку, когда она занимает место госпожи своей.
PROV|30|24|Вот четыре малых на земле, но они мудрее мудрых:
PROV|30|25|муравьи – народ не сильный, но летом заготовляют пищу свою;
PROV|30|26|горные мыши – народ слабый, но ставят домы свои на скале;
PROV|30|27|у саранчи нет царя, но выступает вся она стройно;
PROV|30|28|паук лапками цепляется, но бывает в царских чертогах.
PROV|30|29|Вот трое имеют стройную походку, и четверо стройно выступают:
PROV|30|30|лев, силач между зверями, не посторонится ни перед кем;
PROV|30|31|конь и козел, и царь среди народа своего.
PROV|30|32|Если ты в заносчивости своей сделал глупость и помыслил злое, то [положи] руку на уста;
PROV|30|33|потому что, как сбивание молока производит масло, толчок в нос производит кровь, так и возбуждение гнева производит ссору.
PROV|31|1|Слова Лемуила царя. Наставление, которое преподала ему мать его:
PROV|31|2|что, сын мой? что, сын чрева моего? что, сын обетов моих?
PROV|31|3|Не отдавай женщинам сил твоих, ни путей твоих губительницам царей.
PROV|31|4|Не царям, Лемуил, не царям пить вино, и не князьям – сикеру,
PROV|31|5|чтобы, напившись, они не забыли закона и не превратили суда всех угнетаемых.
PROV|31|6|Дайте сикеру погибающему и вино огорченному душею;
PROV|31|7|пусть он выпьет и забудет бедность свою и не вспомнит больше о своем страдании.
PROV|31|8|Открывай уста твои за безгласного и для защиты всех сирот.
PROV|31|9|Открывай уста твои для правосудия и для дела бедного и нищего.
PROV|31|10|Кто найдет добродетельную жену? цена ее выше жемчугов;
PROV|31|11|уверено в ней сердце мужа ее, и он не останется без прибытка;
PROV|31|12|она воздает ему добром, а не злом, во все дни жизни своей.
PROV|31|13|Добывает шерсть и лен, и с охотою работает своими руками.
PROV|31|14|Она, как купеческие корабли, издалека добывает хлеб свой.
PROV|31|15|Она встает еще ночью и раздает пищу в доме своем и урочное служанкам своим.
PROV|31|16|Задумает она о поле, и приобретает его; от плодов рук своих насаждает виноградник.
PROV|31|17|Препоясывает силою чресла свои и укрепляет мышцы свои.
PROV|31|18|Она чувствует, что занятие ее хорошо, и – светильник ее не гаснет и ночью.
PROV|31|19|Протягивает руки свои к прялке, и персты ее берутся за веретено.
PROV|31|20|Длань свою она открывает бедному, и руку свою подает нуждающемуся.
PROV|31|21|Не боится стужи для семьи своей, потому что вся семья ее одета в двойные одежды.
PROV|31|22|Она делает себе ковры; виссон и пурпур – одежда ее.
PROV|31|23|Муж ее известен у ворот, когда сидит со старейшинами земли.
PROV|31|24|Она делает покрывала и продает, и поясы доставляет купцам Финикийским.
PROV|31|25|Крепость и красота – одежда ее, и весело смотрит она на будущее.
PROV|31|26|Уста свои открывает с мудростью, и кроткое наставление на языке ее.
PROV|31|27|Она наблюдает за хозяйством в доме своем и не ест хлеба праздности.
PROV|31|28|Встают дети и ублажают ее, – муж, и хвалит ее:
PROV|31|29|"много было жен добродетельных, но ты превзошла всех их".
PROV|31|30|Миловидность обманчива и красота суетна; но жена, боящаяся Господа, достойна хвалы.
PROV|31|31|Дайте ей от плода рук ее, и да прославят ее у ворот дела ее!
